* PEX produced on Tue Jul 15 06:06:44 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic_11.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic_11 VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 GNDA.t194 bgr_0.NFET_GATE_10uA.t5 two_stage_opamp_dummy_magic_16_0.Vb3.t4 GNDA.t193 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1 bgr_0.V_TOP.t11 VDDA.t374 VDDA.t376 VDDA.t375 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.45 ps=2.9 w=1 l=0.15
X2 VOUT-.t19 two_stage_opamp_dummy_magic_16_0.cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 VOUT+.t19 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t9 two_stage_opamp_dummy_magic_16_0.X.t25 VDDA.t159 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X5 VOUT+.t20 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 GNDA.t305 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t2 VOUT-.t17 GNDA.t304 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X7 VDDA.t117 bgr_0.V_TOP.t14 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t5 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X8 VOUT+.t21 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 two_stage_opamp_dummy_magic_16_0.V_source.t24 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t12 GNDA.t142 GNDA.t141 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X10 bgr_0.Vin+.t5 bgr_0.V_TOP.t15 VDDA.t60 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X11 VDDA.t263 two_stage_opamp_dummy_magic_16_0.Vb3.t8 two_stage_opamp_dummy_magic_16_0.VD3.t27 VDDA.t262 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X12 GNDA.t144 VDDA.t371 VDDA.t373 VDDA.t372 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X13 VDDA.t83 bgr_0.V_mir1.t17 bgr_0.1st_Vout_1.t5 VDDA.t82 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X14 VOUT+.t22 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 bgr_0.1st_Vout_2.t11 bgr_0.cap_res2.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 two_stage_opamp_dummy_magic_16_0.X.t8 two_stage_opamp_dummy_magic_16_0.Vb2.t11 two_stage_opamp_dummy_magic_16_0.VD3.t11 two_stage_opamp_dummy_magic_16_0.VD3.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X17 two_stage_opamp_dummy_magic_16_0.err_amp_mir.t3 VDDA.t368 VDDA.t370 VDDA.t369 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X18 VOUT+.t23 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X19 bgr_0.1st_Vout_2.t8 bgr_0.V_CUR_REF_REG.t3 bgr_0.V_p_2.t9 GNDA.t104 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X20 VOUT+.t24 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 VOUT+.t25 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 a_7460_23988.t0 bgr_0.Vin+.t0 GNDA.t2 sky130_fd_pr__res_xhigh_po_0p35 l=6
X23 VOUT+.t26 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X24 bgr_0.1st_Vout_2.t12 bgr_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 two_stage_opamp_dummy_magic_16_0.X.t12 two_stage_opamp_dummy_magic_16_0.Vb1.t14 two_stage_opamp_dummy_magic_16_0.VD1.t11 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X26 VDDA.t367 VDDA.t365 bgr_0.NFET_GATE_10uA.t1 VDDA.t366 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X27 GNDA.t51 a_6930_22564.t0 GNDA.t50 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X28 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t7 bgr_0.PFET_GATE_10uA.t10 VDDA.t218 VDDA.t217 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X29 VDDA.t47 bgr_0.PFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t1 VDDA.t46 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X30 VOUT-.t20 two_stage_opamp_dummy_magic_16_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 VOUT-.t21 two_stage_opamp_dummy_magic_16_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 VOUT-.t22 two_stage_opamp_dummy_magic_16_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 two_stage_opamp_dummy_magic_16_0.V_source.t1 VIN+.t0 two_stage_opamp_dummy_magic_16_0.VD2.t19 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X34 VOUT+.t27 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 bgr_0.1st_Vout_1.t11 bgr_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 bgr_0.1st_Vout_2.t0 bgr_0.V_mir2.t17 VDDA.t5 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X37 VDDA.t62 bgr_0.V_TOP.t16 bgr_0.Vin-.t6 VDDA.t61 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X38 bgr_0.1st_Vout_1.t7 bgr_0.Vin+.t6 bgr_0.V_p_1.t4 GNDA.t82 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X39 two_stage_opamp_dummy_magic_16_0.Y.t11 two_stage_opamp_dummy_magic_16_0.Vb1.t15 two_stage_opamp_dummy_magic_16_0.VD2.t0 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X40 GNDA.t152 VDDA.t415 bgr_0.V_p_2.t10 GNDA.t151 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X41 VDDA.t261 two_stage_opamp_dummy_magic_16_0.Vb3.t9 two_stage_opamp_dummy_magic_16_0.VD3.t26 VDDA.t260 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X42 VOUT+.t28 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 bgr_0.cap_res2.t0 bgr_0.PFET_GATE_10uA.t0 GNDA.t46 sky130_fd_pr__res_high_po_0p35 l=2.05
X44 bgr_0.1st_Vout_1.t12 bgr_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t9 two_stage_opamp_dummy_magic_16_0.Y.t25 VDDA.t409 GNDA.t307 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X46 two_stage_opamp_dummy_magic_16_0.V_source.t26 VIN+.t1 two_stage_opamp_dummy_magic_16_0.VD2.t18 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X47 VOUT+.t29 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X48 VOUT-.t23 two_stage_opamp_dummy_magic_16_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 two_stage_opamp_dummy_magic_16_0.V_source.t5 two_stage_opamp_dummy_magic_16_0.Vb1.t16 a_9610_2730.t0 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.6 ps=3.8 w=1.5 l=3
X50 VOUT-.t24 two_stage_opamp_dummy_magic_16_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 VOUT-.t25 two_stage_opamp_dummy_magic_16_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 VDDA.t79 bgr_0.1st_Vout_1.t13 bgr_0.V_TOP.t1 VDDA.t78 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X53 GNDA.t320 two_stage_opamp_dummy_magic_16_0.Y.t26 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t9 VDDA.t412 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X54 bgr_0.V_TOP.t17 VDDA.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 VOUT-.t26 two_stage_opamp_dummy_magic_16_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X56 GNDA.t290 GNDA.t289 two_stage_opamp_dummy_magic_16_0.X.t20 GNDA.t205 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X57 two_stage_opamp_dummy_magic_16_0.VD4.t11 VDDA.t362 VDDA.t364 VDDA.t363 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X58 GNDA.t288 GNDA.t286 bgr_0.NFET_GATE_10uA.t4 GNDA.t287 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X59 bgr_0.START_UP.t5 bgr_0.V_TOP.t18 VDDA.t187 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X60 VOUT-.t27 two_stage_opamp_dummy_magic_16_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 two_stage_opamp_dummy_magic_16_0.V_err_gate.t2 bgr_0.NFET_GATE_10uA.t6 GNDA.t192 GNDA.t191 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X62 bgr_0.1st_Vout_1.t10 bgr_0.Vin+.t7 bgr_0.V_p_1.t3 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X63 VOUT-.t28 two_stage_opamp_dummy_magic_16_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X64 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t8 two_stage_opamp_dummy_magic_16_0.X.t26 VDDA.t133 GNDA.t78 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X65 GNDA.t285 GNDA.t284 two_stage_opamp_dummy_magic_16_0.Y.t14 GNDA.t196 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X66 VOUT+.t30 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 bgr_0.1st_Vout_1.t14 bgr_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 bgr_0.V_TOP.t19 VDDA.t188 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X69 bgr_0.V_mir2.t11 bgr_0.V_mir2.t10 VDDA.t45 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X70 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t15 VDDA.t359 VDDA.t361 VDDA.t360 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X71 VOUT-.t29 two_stage_opamp_dummy_magic_16_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 VOUT-.t6 two_stage_opamp_dummy_magic_16_0.X.t27 VDDA.t135 VDDA.t134 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X73 VOUT+.t5 a_5980_2720.t0 GNDA.t130 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X74 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t13 bgr_0.PFET_GATE_10uA.t12 VDDA.t216 VDDA.t215 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X75 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t8 VDDA.t356 VDDA.t358 VDDA.t357 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X76 VDDA.t67 bgr_0.PFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t12 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X77 VOUT+.t31 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X78 bgr_0.V_TOP.t20 VDDA.t189 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 bgr_0.1st_Vout_2.t10 bgr_0.V_CUR_REF_REG.t4 bgr_0.V_p_2.t8 GNDA.t292 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X80 two_stage_opamp_dummy_magic_16_0.VD4.t37 two_stage_opamp_dummy_magic_16_0.Vb2.t12 two_stage_opamp_dummy_magic_16_0.Y.t18 two_stage_opamp_dummy_magic_16_0.VD4.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X81 VOUT+.t15 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t3 GNDA.t314 GNDA.t313 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X82 VDDA.t202 two_stage_opamp_dummy_magic_16_0.Y.t27 VOUT+.t7 VDDA.t201 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X83 VOUT-.t30 two_stage_opamp_dummy_magic_16_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 two_stage_opamp_dummy_magic_16_0.VD4.t9 two_stage_opamp_dummy_magic_16_0.Vb3.t10 VDDA.t259 VDDA.t258 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X85 VOUT-.t31 two_stage_opamp_dummy_magic_16_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X86 VOUT-.t32 two_stage_opamp_dummy_magic_16_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X87 two_stage_opamp_dummy_magic_16_0.V_err_mir_p.t2 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t7 two_stage_opamp_dummy_magic_16_0.V_err_gate.t0 VDDA.t109 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X88 VOUT-.t16 a_14010_2720.t1 GNDA.t300 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X89 bgr_0.PFET_GATE_10uA.t6 bgr_0.1st_Vout_2.t13 VDDA.t111 VDDA.t110 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X90 VOUT-.t33 two_stage_opamp_dummy_magic_16_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X91 bgr_0.V_TOP.t21 VDDA.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X92 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t9 two_stage_opamp_dummy_magic_16_0.X.t28 GNDA.t76 VDDA.t130 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X93 GNDA.t283 GNDA.t281 two_stage_opamp_dummy_magic_16_0.V_source.t32 GNDA.t282 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X94 bgr_0.START_UP_NFET1.t0 bgr_0.START_UP_NFET1 GNDA.t93 GNDA.t92 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X95 VDDA.t355 VDDA.t353 GNDA.t40 VDDA.t354 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X96 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_16_0.Vb3.t1 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t5 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X97 two_stage_opamp_dummy_magic_16_0.VD3.t9 two_stage_opamp_dummy_magic_16_0.Vb2.t13 two_stage_opamp_dummy_magic_16_0.X.t6 two_stage_opamp_dummy_magic_16_0.VD3.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X98 VOUT+.t32 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X99 two_stage_opamp_dummy_magic_16_0.V_source.t33 VIN+.t2 two_stage_opamp_dummy_magic_16_0.VD2.t17 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X100 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t8 two_stage_opamp_dummy_magic_16_0.Y.t28 VDDA.t96 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X101 two_stage_opamp_dummy_magic_16_0.V_source.t28 VIN-.t0 two_stage_opamp_dummy_magic_16_0.VD1.t14 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X102 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t9 GNDA.t279 GNDA.t280 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X103 VOUT+.t33 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X104 bgr_0.V_TOP.t22 VDDA.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 GNDA.t190 bgr_0.NFET_GATE_10uA.t7 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t13 GNDA.t189 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X106 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t12 bgr_0.NFET_GATE_10uA.t8 GNDA.t188 GNDA.t187 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X107 two_stage_opamp_dummy_magic_16_0.VD4.t35 two_stage_opamp_dummy_magic_16_0.Vb2.t14 two_stage_opamp_dummy_magic_16_0.Y.t23 two_stage_opamp_dummy_magic_16_0.VD4.t34 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X108 GNDA.t291 two_stage_opamp_dummy_magic_16_0.Y.t29 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t8 VDDA.t377 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X109 VOUT-.t34 two_stage_opamp_dummy_magic_16_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X110 VOUT-.t35 two_stage_opamp_dummy_magic_16_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 VOUT-.t36 two_stage_opamp_dummy_magic_16_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X112 VOUT-.t37 two_stage_opamp_dummy_magic_16_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 bgr_0.1st_Vout_2.t14 bgr_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 two_stage_opamp_dummy_magic_16_0.VD1.t10 two_stage_opamp_dummy_magic_16_0.Vb1.t17 two_stage_opamp_dummy_magic_16_0.X.t9 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X115 VOUT+.t34 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X116 VOUT+.t35 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X117 two_stage_opamp_dummy_magic_16_0.Vb1.t8 two_stage_opamp_dummy_magic_16_0.Vb1.t7 a_9610_2730.t4 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X118 VOUT+.t36 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 VOUT+.t37 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 VOUT+.t38 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 a_12530_23988.t1 bgr_0.Vin-.t7 GNDA.t299 sky130_fd_pr__res_xhigh_po_0p35 l=6
X122 two_stage_opamp_dummy_magic_16_0.VD3.t25 two_stage_opamp_dummy_magic_16_0.Vb3.t11 VDDA.t257 VDDA.t256 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X123 two_stage_opamp_dummy_magic_16_0.VD2.t1 two_stage_opamp_dummy_magic_16_0.Vb1.t18 two_stage_opamp_dummy_magic_16_0.Y.t10 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X124 two_stage_opamp_dummy_magic_16_0.VD3.t3 two_stage_opamp_dummy_magic_16_0.Vb2.t15 two_stage_opamp_dummy_magic_16_0.X.t1 two_stage_opamp_dummy_magic_16_0.VD3.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X125 VOUT-.t38 two_stage_opamp_dummy_magic_16_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 VOUT-.t39 two_stage_opamp_dummy_magic_16_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X127 bgr_0.1st_Vout_2.t7 bgr_0.V_mir2.t18 VDDA.t125 VDDA.t124 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X128 VOUT-.t5 two_stage_opamp_dummy_magic_16_0.X.t29 VDDA.t132 VDDA.t131 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X129 VOUT-.t40 two_stage_opamp_dummy_magic_16_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 VOUT-.t41 two_stage_opamp_dummy_magic_16_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 bgr_0.1st_Vout_2.t15 bgr_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X132 VOUT-.t42 two_stage_opamp_dummy_magic_16_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 VOUT+.t39 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 two_stage_opamp_dummy_magic_16_0.V_p_mir.t2 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t13 GNDA.t112 GNDA.t111 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X135 two_stage_opamp_dummy_magic_16_0.V_source.t23 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t14 GNDA.t116 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X136 VOUT-.t43 two_stage_opamp_dummy_magic_16_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X137 VOUT+.t40 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 VOUT+.t41 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 bgr_0.1st_Vout_1.t15 bgr_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 VOUT+.t42 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X141 bgr_0.V_mir1.t16 bgr_0.Vin-.t8 bgr_0.V_p_1.t10 GNDA.t310 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X142 bgr_0.V_mir1.t11 bgr_0.V_mir1.t10 VDDA.t25 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X143 two_stage_opamp_dummy_magic_16_0.VD3.t24 two_stage_opamp_dummy_magic_16_0.Vb3.t12 VDDA.t255 VDDA.t254 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X144 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t2 VIN+.t3 two_stage_opamp_dummy_magic_16_0.V_p_mir.t3 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X145 two_stage_opamp_dummy_magic_16_0.V_source.t0 VIN-.t1 two_stage_opamp_dummy_magic_16_0.VD1.t0 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X146 GNDA.t125 a_7580_22380.t1 GNDA.t2 sky130_fd_pr__res_xhigh_po_0p35 l=6
X147 VOUT-.t44 two_stage_opamp_dummy_magic_16_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 VOUT-.t45 two_stage_opamp_dummy_magic_16_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 VOUT+.t43 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 GNDA.t9 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t15 two_stage_opamp_dummy_magic_16_0.V_source.t22 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X151 VOUT-.t46 two_stage_opamp_dummy_magic_16_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 VOUT-.t47 two_stage_opamp_dummy_magic_16_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X153 GNDA.t114 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t16 two_stage_opamp_dummy_magic_16_0.V_source.t21 GNDA.t113 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X154 VDDA.t175 bgr_0.PFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_16_0.Vb1.t9 VDDA.t174 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X155 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t8 two_stage_opamp_dummy_magic_16_0.X.t30 GNDA.t34 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X156 VOUT-.t48 two_stage_opamp_dummy_magic_16_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 bgr_0.V_TOP.t23 VDDA.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 two_stage_opamp_dummy_magic_16_0.V_source.t40 VIN-.t2 two_stage_opamp_dummy_magic_16_0.VD1.t21 GNDA.t306 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X159 VDDA.t352 VDDA.t350 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t15 VDDA.t351 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X160 VOUT-.t49 two_stage_opamp_dummy_magic_16_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X161 VOUT-.t50 two_stage_opamp_dummy_magic_16_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 GNDA.t318 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t4 VOUT+.t16 GNDA.t317 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X163 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t13 bgr_0.PFET_GATE_10uA.t15 VDDA.t173 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X164 a_5700_5524.t0 two_stage_opamp_dummy_magic_16_0.V_tot.t0 GNDA.t39 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X165 VOUT+.t44 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 VOUT+.t45 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X167 VDDA.t253 two_stage_opamp_dummy_magic_16_0.Vb3.t13 two_stage_opamp_dummy_magic_16_0.VD4.t8 VDDA.t252 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X168 VOUT+.t17 two_stage_opamp_dummy_magic_16_0.Y.t30 VDDA.t414 VDDA.t413 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X169 GNDA.t149 VDDA.t347 VDDA.t349 VDDA.t348 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X170 bgr_0.V_mir1.t13 bgr_0.Vin-.t9 bgr_0.V_p_1.t9 GNDA.t99 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X171 VOUT+.t46 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X172 VOUT+.t47 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X173 two_stage_opamp_dummy_magic_16_0.VD3.t7 two_stage_opamp_dummy_magic_16_0.Vb2.t16 two_stage_opamp_dummy_magic_16_0.X.t4 two_stage_opamp_dummy_magic_16_0.VD3.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X174 two_stage_opamp_dummy_magic_16_0.V_err_gate.t5 two_stage_opamp_dummy_magic_16_0.V_tot.t4 two_stage_opamp_dummy_magic_16_0.V_err_mir_p.t3 VDDA.t386 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X175 GNDA.t278 GNDA.t276 two_stage_opamp_dummy_magic_16_0.err_amp_mir.t2 GNDA.t277 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X176 two_stage_opamp_dummy_magic_16_0.Vb1.t11 GNDA.t273 GNDA.t275 GNDA.t274 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X177 bgr_0.START_UP.t4 bgr_0.V_TOP.t24 VDDA.t205 VDDA.t204 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X178 VOUT-.t51 two_stage_opamp_dummy_magic_16_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X179 bgr_0.PFET_GATE_10uA.t5 bgr_0.1st_Vout_2.t16 VDDA.t20 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X180 VDDA.t185 bgr_0.V_mir1.t18 bgr_0.1st_Vout_1.t4 VDDA.t184 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X181 VOUT+.t48 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 two_stage_opamp_dummy_magic_16_0.VD2.t8 two_stage_opamp_dummy_magic_16_0.Vb1.t19 two_stage_opamp_dummy_magic_16_0.Y.t9 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X183 VOUT+.t49 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X184 VOUT-.t52 two_stage_opamp_dummy_magic_16_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 VOUT-.t53 two_stage_opamp_dummy_magic_16_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 two_stage_opamp_dummy_magic_16_0.VD2.t5 two_stage_opamp_dummy_magic_16_0.Vb1.t20 two_stage_opamp_dummy_magic_16_0.Y.t8 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X187 two_stage_opamp_dummy_magic_16_0.Vb2.t5 bgr_0.NFET_GATE_10uA.t9 GNDA.t172 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X188 VDDA.t251 two_stage_opamp_dummy_magic_16_0.Vb3.t14 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t7 VDDA.t250 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X189 GNDA.t186 bgr_0.NFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_16_0.Vb2.t4 GNDA.t185 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X190 VOUT+.t50 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 bgr_0.V_TOP.t25 VDDA.t206 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 GNDA.t184 bgr_0.NFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_16_0.Vb2.t3 GNDA.t183 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X193 two_stage_opamp_dummy_magic_16_0.Y.t17 two_stage_opamp_dummy_magic_16_0.Vb2.t17 two_stage_opamp_dummy_magic_16_0.VD4.t33 two_stage_opamp_dummy_magic_16_0.VD4.t32 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X194 VOUT+.t51 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 VOUT-.t54 two_stage_opamp_dummy_magic_16_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 VOUT-.t3 two_stage_opamp_dummy_magic_16_0.X.t31 VDDA.t77 VDDA.t76 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X197 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t7 two_stage_opamp_dummy_magic_16_0.Y.t31 GNDA.t302 VDDA.t399 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X198 VDDA.t249 two_stage_opamp_dummy_magic_16_0.Vb3.t15 two_stage_opamp_dummy_magic_16_0.VD4.t7 VDDA.t248 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X199 VOUT+.t52 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X200 VOUT+.t53 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X201 VOUT+.t54 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 VOUT+.t55 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X203 two_stage_opamp_dummy_magic_16_0.VD3.t23 two_stage_opamp_dummy_magic_16_0.Vb3.t16 VDDA.t247 VDDA.t246 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X204 VDDA.t208 bgr_0.V_TOP.t26 bgr_0.Vin+.t4 VDDA.t207 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X205 two_stage_opamp_dummy_magic_16_0.V_source.t20 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t17 GNDA.t110 GNDA.t109 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X206 bgr_0.1st_Vout_2.t1 bgr_0.V_mir2.t19 VDDA.t9 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X207 VOUT-.t55 two_stage_opamp_dummy_magic_16_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t0 a_14010_2720.t0 GNDA.t127 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X209 bgr_0.V_TOP.t13 bgr_0.1st_Vout_1.t16 VDDA.t402 VDDA.t401 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X210 bgr_0.V_CUR_REF_REG.t2 VDDA.t344 VDDA.t346 VDDA.t345 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X211 VOUT-.t56 two_stage_opamp_dummy_magic_16_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 VOUT-.t57 two_stage_opamp_dummy_magic_16_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 VOUT-.t58 two_stage_opamp_dummy_magic_16_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X214 VOUT+.t56 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X215 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t6 bgr_0.PFET_GATE_10uA.t16 VDDA.t199 VDDA.t198 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X216 VOUT-.t59 two_stage_opamp_dummy_magic_16_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 two_stage_opamp_dummy_magic_16_0.V_source.t34 VIN+.t4 two_stage_opamp_dummy_magic_16_0.VD2.t16 GNDA.t294 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X218 VDDA.t73 two_stage_opamp_dummy_magic_16_0.X.t32 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t7 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X219 two_stage_opamp_dummy_magic_16_0.X.t15 two_stage_opamp_dummy_magic_16_0.Vb2.t18 two_stage_opamp_dummy_magic_16_0.VD3.t15 two_stage_opamp_dummy_magic_16_0.VD3.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X220 VOUT+.t57 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X221 GNDA.t140 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t18 two_stage_opamp_dummy_magic_16_0.V_source.t19 GNDA.t139 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X222 VOUT+.t58 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 bgr_0.1st_Vout_2.t17 bgr_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X224 a_6810_23838.t1 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t6 GNDA.t50 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X225 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t7 two_stage_opamp_dummy_magic_16_0.X.t33 GNDA.t33 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X226 two_stage_opamp_dummy_magic_16_0.Y.t19 two_stage_opamp_dummy_magic_16_0.Vb2.t19 two_stage_opamp_dummy_magic_16_0.VD4.t31 two_stage_opamp_dummy_magic_16_0.VD4.t30 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X227 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t7 two_stage_opamp_dummy_magic_16_0.Y.t32 VDDA.t200 GNDA.t143 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X228 bgr_0.Vin+.t1 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 GNDA.t35 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X229 VDDA.t343 VDDA.t341 two_stage_opamp_dummy_magic_16_0.err_amp_out.t3 VDDA.t342 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X230 two_stage_opamp_dummy_magic_16_0.V_source.t3 VIN+.t5 two_stage_opamp_dummy_magic_16_0.VD2.t15 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X231 VOUT+.t59 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 VOUT+.t60 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X233 VOUT-.t60 two_stage_opamp_dummy_magic_16_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X234 VOUT-.t61 two_stage_opamp_dummy_magic_16_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X235 bgr_0.1st_Vout_2.t18 bgr_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 bgr_0.Vin+.t3 bgr_0.V_TOP.t27 VDDA.t141 VDDA.t140 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X237 VOUT-.t62 two_stage_opamp_dummy_magic_16_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X238 VDDA.t340 VDDA.t338 bgr_0.PFET_GATE_10uA.t9 VDDA.t339 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X239 VOUT+.t61 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 VDDA.t143 bgr_0.V_TOP.t28 bgr_0.Vin+.t2 VDDA.t142 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X241 VOUT+.t14 two_stage_opamp_dummy_magic_16_0.Y.t33 VDDA.t394 VDDA.t393 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X242 VOUT+.t62 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X243 a_5580_5524.t1 two_stage_opamp_dummy_magic_16_0.V_tot.t3 GNDA.t319 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X244 two_stage_opamp_dummy_magic_16_0.VD1.t9 two_stage_opamp_dummy_magic_16_0.Vb1.t21 two_stage_opamp_dummy_magic_16_0.X.t11 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X245 bgr_0.1st_Vout_1.t17 bgr_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 GNDA.t13 a_12410_22380.t0 GNDA.t12 sky130_fd_pr__res_xhigh_po_0p35 l=6
X247 GNDA.t182 bgr_0.NFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_16_0.Vb3.t5 GNDA.t181 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X248 VDDA.t388 two_stage_opamp_dummy_magic_16_0.V_err_gate.t6 two_stage_opamp_dummy_magic_16_0.V_err_mir_p.t1 VDDA.t387 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X249 VOUT-.t63 two_stage_opamp_dummy_magic_16_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 VOUT-.t64 two_stage_opamp_dummy_magic_16_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X251 VDDA.t245 two_stage_opamp_dummy_magic_16_0.Vb3.t17 two_stage_opamp_dummy_magic_16_0.VD3.t22 VDDA.t244 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X252 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_16_0.Y.t1 GNDA.t11 sky130_fd_pr__res_high_po_1p41 l=1.41
X253 GNDA.t118 two_stage_opamp_dummy_magic_16_0.err_amp_mir.t5 two_stage_opamp_dummy_magic_16_0.err_amp_out.t0 GNDA.t117 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X254 VOUT+.t63 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X255 bgr_0.cap_res1.t20 bgr_0.V_TOP.t3 GNDA.t74 sky130_fd_pr__res_high_po_0p35 l=2.05
X256 two_stage_opamp_dummy_magic_16_0.Vb3.t3 bgr_0.NFET_GATE_10uA.t13 GNDA.t180 GNDA.t179 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X257 bgr_0.V_mir2.t9 bgr_0.V_mir2.t8 VDDA.t88 VDDA.t87 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X258 VDDA.t337 VDDA.t335 bgr_0.V_TOP.t10 VDDA.t336 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X259 two_stage_opamp_dummy_magic_16_0.X.t0 two_stage_opamp_dummy_magic_16_0.Vb2.t20 two_stage_opamp_dummy_magic_16_0.VD3.t1 two_stage_opamp_dummy_magic_16_0.VD3.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X260 two_stage_opamp_dummy_magic_16_0.VD2.t2 two_stage_opamp_dummy_magic_16_0.Vb1.t22 two_stage_opamp_dummy_magic_16_0.Y.t7 GNDA.t306 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X261 VOUT+.t64 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 VOUT+.t65 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 bgr_0.1st_Vout_1.t18 bgr_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X264 VOUT-.t65 two_stage_opamp_dummy_magic_16_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 VOUT+.t66 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t4 bgr_0.V_TOP.t29 VDDA.t145 VDDA.t144 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X267 bgr_0.1st_Vout_2.t19 bgr_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X268 VOUT-.t0 two_stage_opamp_dummy_magic_16_0.X.t34 VDDA.t50 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X269 VOUT-.t66 two_stage_opamp_dummy_magic_16_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X270 GNDA.t298 a_13060_22630.t1 GNDA.t297 sky130_fd_pr__res_xhigh_po_0p35 l=4
X271 VOUT-.t1 two_stage_opamp_dummy_magic_16_0.X.t35 VDDA.t52 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X272 VOUT+.t67 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X273 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t6 two_stage_opamp_dummy_magic_16_0.Y.t34 GNDA.t107 VDDA.t167 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X274 VDDA.t334 VDDA.t332 GNDA.t148 VDDA.t333 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X275 bgr_0.1st_Vout_1.t3 bgr_0.V_mir1.t19 VDDA.t177 VDDA.t176 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X276 bgr_0.1st_Vout_1.t19 bgr_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 two_stage_opamp_dummy_magic_16_0.X.t18 two_stage_opamp_dummy_magic_16_0.Vb2.t21 two_stage_opamp_dummy_magic_16_0.VD3.t17 two_stage_opamp_dummy_magic_16_0.VD3.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X278 VOUT-.t67 two_stage_opamp_dummy_magic_16_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X279 two_stage_opamp_dummy_magic_16_0.V_source.t18 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t19 GNDA.t81 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X280 VDDA.t243 two_stage_opamp_dummy_magic_16_0.Vb3.t18 two_stage_opamp_dummy_magic_16_0.VD3.t21 VDDA.t242 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X281 a_9610_2730.t3 two_stage_opamp_dummy_magic_16_0.Vb1.t3 two_stage_opamp_dummy_magic_16_0.Vb1.t4 GNDA.t75 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X282 bgr_0.NFET_GATE_10uA.t0 bgr_0.PFET_GATE_10uA.t17 VDDA.t65 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X283 VDDA.t33 bgr_0.PFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t0 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X284 two_stage_opamp_dummy_magic_16_0.Y.t21 two_stage_opamp_dummy_magic_16_0.Vb2.t22 two_stage_opamp_dummy_magic_16_0.VD4.t29 two_stage_opamp_dummy_magic_16_0.VD4.t28 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X285 VOUT+.t68 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 VOUT+.t69 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X287 bgr_0.1st_Vout_1.t20 bgr_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X288 GNDA.t326 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t5 VOUT-.t18 GNDA.t325 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X289 bgr_0.V_p_2.t2 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t8 bgr_0.V_mir2.t16 GNDA.t295 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X290 VDDA.t13 two_stage_opamp_dummy_magic_16_0.X.t36 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t6 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X291 two_stage_opamp_dummy_magic_16_0.V_source.t6 VIN-.t3 two_stage_opamp_dummy_magic_16_0.VD1.t1 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X292 VDDA.t161 bgr_0.V_TOP.t30 bgr_0.START_UP.t3 VDDA.t160 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X293 VOUT+.t70 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X294 VOUT-.t68 two_stage_opamp_dummy_magic_16_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 GNDA.t103 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t20 two_stage_opamp_dummy_magic_16_0.V_source.t17 GNDA.t102 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X296 VOUT-.t69 two_stage_opamp_dummy_magic_16_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X297 a_5700_5524.t1 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t16 GNDA.t316 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X298 VOUT+.t71 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X299 VOUT+.t72 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 bgr_0.V_TOP.t31 VDDA.t162 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 bgr_0.V_TOP.t4 bgr_0.1st_Vout_1.t21 VDDA.t137 VDDA.t136 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X302 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t6 two_stage_opamp_dummy_magic_16_0.X.t37 GNDA.t7 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X303 VOUT+.t73 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 two_stage_opamp_dummy_magic_16_0.VD4.t6 two_stage_opamp_dummy_magic_16_0.Vb3.t19 VDDA.t241 VDDA.t240 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X305 two_stage_opamp_dummy_magic_16_0.V_err_p.t1 two_stage_opamp_dummy_magic_16_0.V_err_gate.t7 VDDA.t39 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X306 two_stage_opamp_dummy_magic_16_0.X.t3 two_stage_opamp_dummy_magic_16_0.Vb2.t23 two_stage_opamp_dummy_magic_16_0.VD3.t5 two_stage_opamp_dummy_magic_16_0.VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X307 GNDA.t272 GNDA.t270 VOUT-.t13 GNDA.t271 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X308 VOUT+.t8 two_stage_opamp_dummy_magic_16_0.Y.t35 VDDA.t213 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X309 VOUT-.t70 two_stage_opamp_dummy_magic_16_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 GNDA.t70 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t21 two_stage_opamp_dummy_magic_16_0.V_source.t16 GNDA.t69 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X311 two_stage_opamp_dummy_magic_16_0.VD1.t8 two_stage_opamp_dummy_magic_16_0.Vb1.t23 two_stage_opamp_dummy_magic_16_0.X.t23 GNDA.t294 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X312 VOUT-.t71 two_stage_opamp_dummy_magic_16_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 bgr_0.V_TOP.t12 bgr_0.1st_Vout_1.t22 VDDA.t390 VDDA.t389 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X314 VOUT+.t74 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 VOUT+.t75 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 VOUT+.t76 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 bgr_0.NFET_GATE_10uA.t3 bgr_0.NFET_GATE_10uA.t2 GNDA.t178 GNDA.t177 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X318 GNDA.t176 bgr_0.NFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_16_0.Vb3.t2 GNDA.t175 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X319 VOUT+.t77 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 bgr_0.V_TOP.t32 VDDA.t163 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X321 VDDA.t331 VDDA.t329 VDDA.t331 VDDA.t330 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X322 two_stage_opamp_dummy_magic_16_0.VD2.t4 two_stage_opamp_dummy_magic_16_0.Vb1.t24 two_stage_opamp_dummy_magic_16_0.Y.t6 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X323 two_stage_opamp_dummy_magic_16_0.VD4.t27 two_stage_opamp_dummy_magic_16_0.Vb2.t24 two_stage_opamp_dummy_magic_16_0.Y.t20 two_stage_opamp_dummy_magic_16_0.VD4.t26 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X324 bgr_0.1st_Vout_2.t20 bgr_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X325 VOUT-.t72 two_stage_opamp_dummy_magic_16_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X326 VOUT-.t73 two_stage_opamp_dummy_magic_16_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X327 VDDA.t68 two_stage_opamp_dummy_magic_16_0.Y.t36 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t6 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X328 VOUT-.t74 two_stage_opamp_dummy_magic_16_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X329 VOUT+.t78 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 two_stage_opamp_dummy_magic_16_0.VD4.t5 two_stage_opamp_dummy_magic_16_0.Vb3.t20 VDDA.t239 VDDA.t238 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X331 VOUT-.t15 VDDA.t326 VDDA.t328 VDDA.t327 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X332 GNDA.t269 GNDA.t268 two_stage_opamp_dummy_magic_16_0.Vb1.t10 GNDA.t57 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X333 VDDA.t7 bgr_0.PFET_GATE_10uA.t19 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t11 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X334 VDDA.t325 VDDA.t323 two_stage_opamp_dummy_magic_16_0.VD3.t29 VDDA.t324 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X335 VOUT-.t75 two_stage_opamp_dummy_magic_16_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X336 bgr_0.1st_Vout_1.t23 bgr_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X337 bgr_0.V_mir1.t9 bgr_0.V_mir1.t8 VDDA.t129 VDDA.t128 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X338 VDDA.t106 bgr_0.V_TOP.t33 bgr_0.START_UP.t2 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X339 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t5 two_stage_opamp_dummy_magic_16_0.Y.t37 GNDA.t38 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X340 VOUT-.t76 two_stage_opamp_dummy_magic_16_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X341 bgr_0.1st_Vout_2.t21 bgr_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X342 VOUT+.t79 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X343 VOUT+.t80 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X344 a_7460_23988.t1 a_7580_22380.t0 GNDA.t2 sky130_fd_pr__res_xhigh_po_0p35 l=6
X345 bgr_0.V_p_2.t7 bgr_0.V_CUR_REF_REG.t5 bgr_0.1st_Vout_2.t5 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X346 VOUT-.t77 two_stage_opamp_dummy_magic_16_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X347 two_stage_opamp_dummy_magic_16_0.V_source.t15 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t22 GNDA.t68 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X348 VOUT+.t81 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X349 two_stage_opamp_dummy_magic_16_0.VD3.t37 two_stage_opamp_dummy_magic_16_0.Vb2.t25 two_stage_opamp_dummy_magic_16_0.X.t24 two_stage_opamp_dummy_magic_16_0.VD3.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X350 VDDA.t89 two_stage_opamp_dummy_magic_16_0.X.t38 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t5 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X351 bgr_0.1st_Vout_2.t22 bgr_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X352 two_stage_opamp_dummy_magic_16_0.VD4.t25 two_stage_opamp_dummy_magic_16_0.Vb2.t26 two_stage_opamp_dummy_magic_16_0.Y.t22 two_stage_opamp_dummy_magic_16_0.VD4.t24 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X353 two_stage_opamp_dummy_magic_16_0.V_source.t2 VIN+.t6 two_stage_opamp_dummy_magic_16_0.VD2.t14 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X354 GNDA.t122 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t23 two_stage_opamp_dummy_magic_16_0.V_source.t14 GNDA.t121 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X355 bgr_0.1st_Vout_1.t9 bgr_0.Vin+.t8 bgr_0.V_p_1.t2 GNDA.t72 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X356 VDDA.t58 bgr_0.V_mir2.t20 bgr_0.1st_Vout_2.t2 VDDA.t57 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X357 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t5 two_stage_opamp_dummy_magic_16_0.X.t39 GNDA.t42 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X358 VOUT-.t78 two_stage_opamp_dummy_magic_16_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 VOUT-.t79 two_stage_opamp_dummy_magic_16_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X360 bgr_0.1st_Vout_1.t24 bgr_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X361 GNDA.t211 GNDA.t260 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X362 VOUT-.t80 two_stage_opamp_dummy_magic_16_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 bgr_0.1st_Vout_2.t23 bgr_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 two_stage_opamp_dummy_magic_16_0.V_err_p.t2 two_stage_opamp_dummy_magic_16_0.V_tot.t5 two_stage_opamp_dummy_magic_16_0.err_amp_mir.t4 VDDA.t378 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X365 GNDA.t174 bgr_0.NFET_GATE_10uA.t15 two_stage_opamp_dummy_magic_16_0.Vb2.t2 GNDA.t173 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X366 two_stage_opamp_dummy_magic_16_0.Vb2.t1 bgr_0.NFET_GATE_10uA.t16 GNDA.t170 GNDA.t169 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X367 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t14 GNDA.t265 GNDA.t267 GNDA.t266 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X368 VOUT+.t82 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X369 GNDA.t211 GNDA.t261 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X370 GNDA.t264 GNDA.t262 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t14 GNDA.t263 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X371 GNDA.t259 GNDA.t257 two_stage_opamp_dummy_magic_16_0.Vb2.t7 GNDA.t258 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X372 VOUT-.t81 two_stage_opamp_dummy_magic_16_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 VOUT+.t83 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X374 bgr_0.PFET_GATE_10uA.t8 VDDA.t320 VDDA.t322 VDDA.t321 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X375 two_stage_opamp_dummy_magic_16_0.VD3.t20 two_stage_opamp_dummy_magic_16_0.Vb3.t21 VDDA.t237 VDDA.t236 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X376 VOUT+.t84 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X377 bgr_0.1st_Vout_1.t2 bgr_0.V_mir1.t20 VDDA.t183 VDDA.t182 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X378 VOUT+.t1 two_stage_opamp_dummy_magic_16_0.Y.t38 VDDA.t29 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X379 two_stage_opamp_dummy_magic_16_0.VD1.t7 two_stage_opamp_dummy_magic_16_0.Vb1.t25 two_stage_opamp_dummy_magic_16_0.X.t21 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X380 two_stage_opamp_dummy_magic_16_0.Vb2_2.t9 two_stage_opamp_dummy_magic_16_0.Vb2.t27 VDDA.t408 VDDA.t407 sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.36 ps=2.2 w=1.8 l=0.2
X381 VOUT-.t82 two_stage_opamp_dummy_magic_16_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 VOUT-.t12 GNDA.t254 GNDA.t256 GNDA.t255 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X383 two_stage_opamp_dummy_magic_16_0.VD4.t4 two_stage_opamp_dummy_magic_16_0.Vb3.t22 VDDA.t235 VDDA.t234 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X384 bgr_0.V_p_2.t6 bgr_0.V_CUR_REF_REG.t6 bgr_0.1st_Vout_2.t3 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X385 VOUT-.t83 two_stage_opamp_dummy_magic_16_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X386 two_stage_opamp_dummy_magic_16_0.VD1.t15 VIN-.t4 two_stage_opamp_dummy_magic_16_0.V_source.t30 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X387 VOUT+.t85 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 GNDA.t211 GNDA.t241 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X389 VOUT-.t84 two_stage_opamp_dummy_magic_16_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X390 VOUT+.t86 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X391 GNDA.t211 GNDA.t240 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X392 VOUT-.t85 two_stage_opamp_dummy_magic_16_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X393 VDDA.t56 two_stage_opamp_dummy_magic_16_0.Y.t39 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t5 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X394 two_stage_opamp_dummy_magic_16_0.VD1.t13 VIN-.t5 two_stage_opamp_dummy_magic_16_0.V_source.t27 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X395 VDDA.t31 bgr_0.V_mir2.t6 bgr_0.V_mir2.t7 VDDA.t30 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X396 VOUT+.t87 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X397 VOUT+.t88 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X398 VOUT+.t89 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 VOUT+.t90 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t4 two_stage_opamp_dummy_magic_16_0.Y.t40 GNDA.t71 VDDA.t126 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X401 bgr_0.V_p_2.t5 bgr_0.V_CUR_REF_REG.t7 bgr_0.1st_Vout_2.t4 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X402 two_stage_opamp_dummy_magic_16_0.VD4.t17 two_stage_opamp_dummy_magic_16_0.VD4.t15 two_stage_opamp_dummy_magic_16_0.Y.t12 two_stage_opamp_dummy_magic_16_0.VD4.t16 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X403 VOUT+.t91 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 a_13180_23838.t1 bgr_0.V_CUR_REF_REG.t1 GNDA.t153 sky130_fd_pr__res_xhigh_po_0p35 l=4
X405 VOUT-.t86 two_stage_opamp_dummy_magic_16_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 bgr_0.V_TOP.t34 VDDA.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X407 VOUT-.t87 two_stage_opamp_dummy_magic_16_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X408 VOUT-.t88 two_stage_opamp_dummy_magic_16_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X409 VOUT-.t89 two_stage_opamp_dummy_magic_16_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 VOUT-.t90 two_stage_opamp_dummy_magic_16_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 VDDA.t157 two_stage_opamp_dummy_magic_16_0.X.t40 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t4 GNDA.t96 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X412 VOUT-.t91 two_stage_opamp_dummy_magic_16_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X413 VOUT+.t92 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 bgr_0.V_TOP.t35 VDDA.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X415 a_5580_5524.t0 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t10 GNDA.t86 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X416 VDDA.t158 two_stage_opamp_dummy_magic_16_0.X.t41 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t3 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X417 VDDA.t233 two_stage_opamp_dummy_magic_16_0.Vb3.t23 two_stage_opamp_dummy_magic_16_0.VD4.t3 VDDA.t232 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X418 VDDA.t406 bgr_0.1st_Vout_2.t24 bgr_0.PFET_GATE_10uA.t4 VDDA.t405 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X419 VDDA.t319 VDDA.t317 two_stage_opamp_dummy_magic_16_0.Vb1.t13 VDDA.t318 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X420 VOUT+.t93 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 two_stage_opamp_dummy_magic_16_0.Vb1.t12 VDDA.t314 VDDA.t316 VDDA.t315 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X422 VDDA.t152 two_stage_opamp_dummy_magic_16_0.X.t42 VOUT-.t8 VDDA.t151 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X423 VOUT-.t92 two_stage_opamp_dummy_magic_16_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X424 VDDA.t313 VDDA.t311 VOUT-.t14 VDDA.t312 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X425 VOUT+.t94 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X426 VOUT+.t95 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 VOUT+.t96 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t12 bgr_0.PFET_GATE_10uA.t20 VDDA.t211 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X429 two_stage_opamp_dummy_magic_16_0.VD3.t35 two_stage_opamp_dummy_magic_16_0.VD3.t33 two_stage_opamp_dummy_magic_16_0.X.t7 two_stage_opamp_dummy_magic_16_0.VD3.t34 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X430 VOUT-.t93 two_stage_opamp_dummy_magic_16_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 VOUT-.t94 two_stage_opamp_dummy_magic_16_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 VDDA.t121 bgr_0.PFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t11 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X433 VOUT-.t95 two_stage_opamp_dummy_magic_16_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 VOUT+.t13 two_stage_opamp_dummy_magic_16_0.Y.t41 VDDA.t385 VDDA.t384 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X435 VOUT-.t96 two_stage_opamp_dummy_magic_16_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 two_stage_opamp_dummy_magic_16_0.cap_res_X.t0 two_stage_opamp_dummy_magic_16_0.X.t13 GNDA.t85 sky130_fd_pr__res_high_po_1p41 l=1.41
X437 VOUT-.t97 two_stage_opamp_dummy_magic_16_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 bgr_0.V_TOP.t36 VDDA.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 two_stage_opamp_dummy_magic_16_0.VD1.t6 two_stage_opamp_dummy_magic_16_0.Vb1.t26 two_stage_opamp_dummy_magic_16_0.X.t2 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X440 VOUT-.t98 two_stage_opamp_dummy_magic_16_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 bgr_0.Vin-.t5 bgr_0.V_TOP.t37 VDDA.t102 VDDA.t101 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X442 two_stage_opamp_dummy_magic_16_0.Y.t16 two_stage_opamp_dummy_magic_16_0.Vb2.t28 two_stage_opamp_dummy_magic_16_0.VD4.t23 two_stage_opamp_dummy_magic_16_0.VD4.t22 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X443 VOUT-.t99 two_stage_opamp_dummy_magic_16_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X444 VDDA.t310 VDDA.t307 VDDA.t309 VDDA.t308 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0 ps=0 w=1.8 l=0.2
X445 a_14170_5524.t0 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t10 GNDA.t10 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X446 VOUT+.t97 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X447 VOUT+.t98 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X448 VDDA.t231 two_stage_opamp_dummy_magic_16_0.Vb3.t24 two_stage_opamp_dummy_magic_16_0.VD4.t2 VDDA.t230 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X449 VOUT+.t99 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X450 GNDA.t168 bgr_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t13 GNDA.t167 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X451 bgr_0.1st_Vout_1.t1 bgr_0.V_mir1.t21 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X452 two_stage_opamp_dummy_magic_16_0.Vb2.t6 GNDA.t251 GNDA.t253 GNDA.t252 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X453 VOUT+.t100 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X454 VOUT+.t101 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X455 VOUT+.t102 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 bgr_0.1st_Vout_1.t25 bgr_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X457 GNDA.t324 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t6 VOUT+.t18 GNDA.t323 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X458 VOUT-.t100 two_stage_opamp_dummy_magic_16_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 bgr_0.1st_Vout_2.t25 bgr_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 VDDA.t48 two_stage_opamp_dummy_magic_16_0.Y.t42 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t4 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X461 VOUT+.t103 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 two_stage_opamp_dummy_magic_16_0.VD2.t13 VIN+.t7 two_stage_opamp_dummy_magic_16_0.V_source.t29 GNDA.t128 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X463 VOUT-.t101 two_stage_opamp_dummy_magic_16_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X464 bgr_0.1st_Vout_1.t26 bgr_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X465 VOUT-.t102 two_stage_opamp_dummy_magic_16_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X466 VOUT-.t103 two_stage_opamp_dummy_magic_16_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X467 VOUT-.t104 two_stage_opamp_dummy_magic_16_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X468 two_stage_opamp_dummy_magic_16_0.X.t5 two_stage_opamp_dummy_magic_16_0.Vb1.t27 two_stage_opamp_dummy_magic_16_0.VD1.t5 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X469 VDDA.t229 two_stage_opamp_dummy_magic_16_0.Vb3.t25 two_stage_opamp_dummy_magic_16_0.VD4.t1 VDDA.t228 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X470 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t5 bgr_0.PFET_GATE_10uA.t22 VDDA.t195 VDDA.t194 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X471 VOUT-.t105 two_stage_opamp_dummy_magic_16_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t3 bgr_0.V_TOP.t38 VDDA.t104 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X473 VOUT+.t104 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 GNDA.t250 GNDA.t248 VOUT+.t10 GNDA.t249 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X475 VDDA.t197 bgr_0.V_mir2.t4 bgr_0.V_mir2.t5 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X476 VOUT+.t105 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X477 VDDA.t139 bgr_0.V_mir1.t6 bgr_0.V_mir1.t7 VDDA.t138 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X478 VDDA.t119 bgr_0.PFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t4 VDDA.t118 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X479 bgr_0.V_p_1.t8 bgr_0.Vin-.t10 bgr_0.V_mir1.t15 GNDA.t145 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X480 VDDA.t267 GNDA.t245 GNDA.t247 GNDA.t246 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X481 two_stage_opamp_dummy_magic_16_0.Vb2.t8 two_stage_opamp_dummy_magic_16_0.Vb2_2.t3 two_stage_opamp_dummy_magic_16_0.Vb2_2.t5 two_stage_opamp_dummy_magic_16_0.Vb2_2.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X482 two_stage_opamp_dummy_magic_16_0.Y.t5 two_stage_opamp_dummy_magic_16_0.Vb1.t28 two_stage_opamp_dummy_magic_16_0.VD2.t6 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X483 VOUT+.t106 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X484 bgr_0.1st_Vout_1.t27 bgr_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X485 bgr_0.1st_Vout_2.t26 bgr_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X486 VOUT+.t107 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X487 VOUT+.t108 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 VDDA.t154 two_stage_opamp_dummy_magic_16_0.X.t43 VOUT-.t9 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X489 bgr_0.V_TOP.t9 VDDA.t304 VDDA.t306 VDDA.t305 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X490 VOUT+.t109 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X491 bgr_0.1st_Vout_1.t28 bgr_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X492 VOUT-.t106 two_stage_opamp_dummy_magic_16_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 VDDA.t303 VDDA.t301 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t1 VDDA.t302 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X494 VDDA.t300 VDDA.t298 two_stage_opamp_dummy_magic_16_0.Vb2_2.t6 VDDA.t299 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.36 ps=2.2 w=1.8 l=0.2
X495 a_14290_5524.t0 two_stage_opamp_dummy_magic_16_0.V_tot.t2 GNDA.t56 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X496 VOUT+.t12 VDDA.t295 VDDA.t297 VDDA.t296 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X497 VDDA.t294 VDDA.t292 two_stage_opamp_dummy_magic_16_0.VD4.t10 VDDA.t293 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X498 bgr_0.V_p_1.t7 bgr_0.Vin-.t11 bgr_0.V_mir1.t14 GNDA.t105 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X499 VOUT+.t110 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X500 VOUT-.t107 two_stage_opamp_dummy_magic_16_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X501 VOUT+.t111 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X502 VOUT+.t112 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X503 VOUT+.t113 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X504 bgr_0.1st_Vout_1.t29 bgr_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X505 two_stage_opamp_dummy_magic_16_0.Vb3.t0 GNDA.t242 GNDA.t244 GNDA.t243 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X506 VOUT+.t114 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X507 two_stage_opamp_dummy_magic_16_0.V_err_gate.t4 VDDA.t289 VDDA.t291 VDDA.t290 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X508 bgr_0.Vin-.t1 bgr_0.START_UP.t6 bgr_0.V_TOP.t2 VDDA.t127 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X509 GNDA.t239 GNDA.t237 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t8 GNDA.t238 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X510 two_stage_opamp_dummy_magic_16_0.VD2.t12 VIN+.t8 two_stage_opamp_dummy_magic_16_0.V_source.t4 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X511 bgr_0.V_TOP.t0 bgr_0.START_UP.t7 bgr_0.Vin-.t0 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X512 VOUT-.t108 two_stage_opamp_dummy_magic_16_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X513 VOUT+.t115 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X514 VOUT+.t116 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X515 two_stage_opamp_dummy_magic_16_0.V_source.t13 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t24 GNDA.t62 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X516 VDDA.t411 bgr_0.1st_Vout_2.t27 bgr_0.PFET_GATE_10uA.t3 VDDA.t410 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X517 bgr_0.V_mir1.t5 bgr_0.V_mir1.t4 VDDA.t392 VDDA.t391 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X518 VOUT-.t109 two_stage_opamp_dummy_magic_16_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X519 VOUT-.t110 two_stage_opamp_dummy_magic_16_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X520 two_stage_opamp_dummy_magic_16_0.V_source.t38 two_stage_opamp_dummy_magic_16_0.err_amp_out.t4 GNDA.t312 GNDA.t311 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X521 GNDA.t43 two_stage_opamp_dummy_magic_16_0.X.t44 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t4 VDDA.t91 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X522 VOUT-.t111 two_stage_opamp_dummy_magic_16_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 GNDA.t211 GNDA.t226 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X524 bgr_0.START_UP.t1 bgr_0.START_UP.t0 bgr_0.START_UP_NFET1.t0 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X525 bgr_0.V_p_2.t3 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t9 bgr_0.V_mir2.t15 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X526 two_stage_opamp_dummy_magic_16_0.VD2.t11 VIN+.t9 two_stage_opamp_dummy_magic_16_0.V_source.t31 GNDA.t129 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X527 VDDA.t221 two_stage_opamp_dummy_magic_16_0.Y.t43 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t3 GNDA.t154 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X528 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t3 two_stage_opamp_dummy_magic_16_0.Y.t44 GNDA.t5 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X529 VDDA.t165 two_stage_opamp_dummy_magic_16_0.Y.t45 VOUT+.t3 VDDA.t164 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X530 VOUT+.t117 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X531 VOUT+.t118 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 VOUT-.t112 two_stage_opamp_dummy_magic_16_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X533 bgr_0.1st_Vout_2.t28 bgr_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X534 VDDA.t288 VDDA.t286 two_stage_opamp_dummy_magic_16_0.V_err_gate.t3 VDDA.t287 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X535 VOUT-.t113 two_stage_opamp_dummy_magic_16_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X536 VOUT+.t119 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X537 a_9610_2730.t2 two_stage_opamp_dummy_magic_16_0.Vb1.t1 two_stage_opamp_dummy_magic_16_0.Vb1.t2 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X538 VDDA.t396 bgr_0.PFET_GATE_10uA.t24 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t10 VDDA.t395 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X539 VDDA.t171 bgr_0.V_mir2.t21 bgr_0.1st_Vout_2.t9 VDDA.t170 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X540 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t11 bgr_0.PFET_GATE_10uA.t25 VDDA.t398 VDDA.t397 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X541 VOUT-.t114 two_stage_opamp_dummy_magic_16_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X542 bgr_0.V_p_1.t6 bgr_0.Vin-.t12 bgr_0.V_mir1.t12 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X543 two_stage_opamp_dummy_magic_16_0.VD4.t0 two_stage_opamp_dummy_magic_16_0.Vb3.t26 VDDA.t227 VDDA.t226 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X544 GNDA.t211 GNDA.t236 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X545 bgr_0.1st_Vout_2.t29 bgr_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X546 VOUT-.t115 two_stage_opamp_dummy_magic_16_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 VOUT-.t116 two_stage_opamp_dummy_magic_16_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X548 two_stage_opamp_dummy_magic_16_0.Y.t4 two_stage_opamp_dummy_magic_16_0.Vb1.t29 two_stage_opamp_dummy_magic_16_0.VD2.t9 GNDA.t128 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X549 VOUT+.t120 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X550 VOUT+.t9 GNDA.t233 GNDA.t235 GNDA.t234 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X551 VOUT-.t117 two_stage_opamp_dummy_magic_16_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X552 VOUT+.t121 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X553 two_stage_opamp_dummy_magic_16_0.err_amp_out.t2 GNDA.t227 GNDA.t229 GNDA.t228 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X554 bgr_0.1st_Vout_1.t30 bgr_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X555 GNDA.t231 GNDA.t230 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X556 VDDA.t93 two_stage_opamp_dummy_magic_16_0.X.t45 VOUT-.t4 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X557 a_6810_23838.t0 a_6930_22564.t1 GNDA.t50 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X558 VOUT+.t122 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X559 GNDA.t211 GNDA.t232 bgr_0.Vin-.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X560 VOUT+.t123 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 bgr_0.1st_Vout_2.t30 bgr_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X562 VDDA.t225 two_stage_opamp_dummy_magic_16_0.Vb3.t27 two_stage_opamp_dummy_magic_16_0.VD3.t19 VDDA.t224 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X563 GNDA.t120 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t25 two_stage_opamp_dummy_magic_16_0.V_source.t12 GNDA.t119 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X564 GNDA.t225 GNDA.t222 GNDA.t224 GNDA.t223 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X565 VOUT+.t6 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t7 GNDA.t136 GNDA.t135 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X566 VOUT+.t124 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X567 GNDA.t166 bgr_0.NFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_16_0.V_err_gate.t1 GNDA.t165 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X568 bgr_0.Vin-.t4 bgr_0.V_TOP.t39 VDDA.t113 VDDA.t112 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X569 a_14290_5524.t1 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t16 GNDA.t315 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X570 a_12530_23988.t0 a_12410_22380.t1 GNDA.t84 sky130_fd_pr__res_xhigh_po_0p35 l=6
X571 two_stage_opamp_dummy_magic_16_0.Vb3.t6 bgr_0.NFET_GATE_10uA.t19 GNDA.t164 GNDA.t163 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X572 bgr_0.1st_Vout_2.t31 bgr_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X573 two_stage_opamp_dummy_magic_16_0.V_p_mir.t0 VIN-.t6 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t3 GNDA.t57 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X574 two_stage_opamp_dummy_magic_16_0.VD1.t12 VIN-.t7 two_stage_opamp_dummy_magic_16_0.V_source.t25 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X575 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t2 two_stage_opamp_dummy_magic_16_0.X.t46 VDDA.t155 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X576 GNDA.t221 GNDA.t219 VDDA.t266 GNDA.t220 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X577 VOUT-.t118 two_stage_opamp_dummy_magic_16_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X578 VDDA.t11 bgr_0.V_mir2.t2 bgr_0.V_mir2.t3 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X579 two_stage_opamp_dummy_magic_16_0.V_source.t11 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t26 GNDA.t124 GNDA.t123 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X580 VOUT+.t125 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X581 bgr_0.1st_Vout_1.t31 bgr_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X582 bgr_0.1st_Vout_2.t32 bgr_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X583 bgr_0.V_p_1.t5 VDDA.t416 GNDA.t132 GNDA.t131 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X584 GNDA.t95 two_stage_opamp_dummy_magic_16_0.X.t47 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t3 VDDA.t156 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X585 VDDA.t381 two_stage_opamp_dummy_magic_16_0.Y.t46 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t2 GNDA.t293 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X586 VDDA.t285 VDDA.t283 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t14 VDDA.t284 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X587 two_stage_opamp_dummy_magic_16_0.VD1.t19 VIN-.t8 two_stage_opamp_dummy_magic_16_0.V_source.t37 GNDA.t303 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X588 VOUT+.t126 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X589 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t10 bgr_0.PFET_GATE_10uA.t26 VDDA.t54 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X590 VOUT-.t119 two_stage_opamp_dummy_magic_16_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X591 VOUT-.t120 two_stage_opamp_dummy_magic_16_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X592 a_13180_23838.t0 a_13060_22630.t0 GNDA.t55 sky130_fd_pr__res_xhigh_po_0p35 l=4
X593 VOUT+.t127 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X594 VOUT+.t128 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X595 VOUT+.t129 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X596 VDDA.t169 two_stage_opamp_dummy_magic_16_0.Y.t47 VOUT+.t4 VDDA.t168 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X597 VDDA.t273 VDDA.t271 VOUT+.t11 VDDA.t272 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X598 bgr_0.V_p_1.t1 bgr_0.Vin+.t9 bgr_0.1st_Vout_1.t8 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X599 VDDA.t3 bgr_0.V_mir1.t22 bgr_0.1st_Vout_1.t0 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X600 two_stage_opamp_dummy_magic_16_0.X.t17 two_stage_opamp_dummy_magic_16_0.Vb1.t30 two_stage_opamp_dummy_magic_16_0.VD1.t4 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X601 bgr_0.V_TOP.t40 VDDA.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X602 two_stage_opamp_dummy_magic_16_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_16_0.V_err_gate.t8 VDDA.t380 VDDA.t379 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X603 two_stage_opamp_dummy_magic_16_0.Vb2_2.t8 two_stage_opamp_dummy_magic_16_0.Vb2.t9 two_stage_opamp_dummy_magic_16_0.Vb2.t10 two_stage_opamp_dummy_magic_16_0.Vb2_2.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X604 two_stage_opamp_dummy_magic_16_0.err_amp_mir.t1 two_stage_opamp_dummy_magic_16_0.err_amp_mir.t0 GNDA.t53 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X605 VOUT-.t121 two_stage_opamp_dummy_magic_16_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X606 VOUT-.t122 two_stage_opamp_dummy_magic_16_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X607 VOUT-.t123 two_stage_opamp_dummy_magic_16_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X608 two_stage_opamp_dummy_magic_16_0.Y.t3 two_stage_opamp_dummy_magic_16_0.Vb1.t31 two_stage_opamp_dummy_magic_16_0.VD2.t3 GNDA.t129 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X609 VOUT-.t124 two_stage_opamp_dummy_magic_16_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X610 VOUT+.t130 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X611 VOUT+.t131 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X612 VDDA.t149 two_stage_opamp_dummy_magic_16_0.X.t48 VOUT-.t7 VDDA.t148 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X613 bgr_0.V_TOP.t41 VDDA.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X614 a_14170_5524.t1 two_stage_opamp_dummy_magic_16_0.V_tot.t1 GNDA.t44 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X615 bgr_0.V_p_1.t0 bgr_0.Vin+.t10 bgr_0.1st_Vout_1.t6 GNDA.t126 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X616 VDDA.t282 VDDA.t280 bgr_0.V_TOP.t8 VDDA.t281 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X617 VOUT-.t125 two_stage_opamp_dummy_magic_16_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X618 two_stage_opamp_dummy_magic_16_0.Vb2.t0 bgr_0.NFET_GATE_10uA.t20 GNDA.t162 GNDA.t161 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X619 GNDA.t160 bgr_0.NFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t11 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X620 GNDA.t29 two_stage_opamp_dummy_magic_16_0.Y.t48 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t2 VDDA.t69 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X621 VOUT-.t126 two_stage_opamp_dummy_magic_16_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X622 VOUT-.t127 two_stage_opamp_dummy_magic_16_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X623 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t12 bgr_0.NFET_GATE_10uA.t22 GNDA.t158 GNDA.t157 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X624 bgr_0.V_TOP.t42 VDDA.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X625 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t0 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t1 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0 ps=0 w=3.5 l=0.2
X626 bgr_0.V_TOP.t43 VDDA.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X627 GNDA.t66 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t27 two_stage_opamp_dummy_magic_16_0.V_source.t10 GNDA.t65 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X628 VOUT-.t128 two_stage_opamp_dummy_magic_16_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X629 two_stage_opamp_dummy_magic_16_0.Vb1.t6 two_stage_opamp_dummy_magic_16_0.Vb1.t5 a_9610_2730.t1 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X630 VOUT-.t129 two_stage_opamp_dummy_magic_16_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X631 VDDA.t123 bgr_0.V_mir2.t22 bgr_0.1st_Vout_2.t6 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X632 two_stage_opamp_dummy_magic_16_0.VD4.t21 two_stage_opamp_dummy_magic_16_0.Vb2.t29 two_stage_opamp_dummy_magic_16_0.Y.t15 two_stage_opamp_dummy_magic_16_0.VD4.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X633 VOUT-.t130 two_stage_opamp_dummy_magic_16_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X634 VDDA.t181 bgr_0.1st_Vout_1.t32 bgr_0.V_TOP.t6 VDDA.t180 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X635 VOUT+.t132 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X636 VOUT-.t131 two_stage_opamp_dummy_magic_16_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X637 VOUT-.t132 two_stage_opamp_dummy_magic_16_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X638 two_stage_opamp_dummy_magic_16_0.VD2.t21 GNDA.t217 GNDA.t218 GNDA.t208 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X639 two_stage_opamp_dummy_magic_16_0.VD2.t10 VIN+.t10 two_stage_opamp_dummy_magic_16_0.V_source.t36 GNDA.t301 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X640 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t1 two_stage_opamp_dummy_magic_16_0.X.t49 VDDA.t150 GNDA.t90 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X641 VOUT+.t133 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X642 two_stage_opamp_dummy_magic_16_0.V_source.t9 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t28 GNDA.t64 GNDA.t63 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X643 VOUT+.t134 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X644 GNDA.t30 two_stage_opamp_dummy_magic_16_0.X.t50 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t2 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X645 bgr_0.V_TOP.t44 VDDA.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X646 VDDA.t265 GNDA.t214 GNDA.t216 GNDA.t215 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X647 two_stage_opamp_dummy_magic_16_0.err_amp_out.t1 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t10 two_stage_opamp_dummy_magic_16_0.V_err_p.t3 VDDA.t400 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X648 two_stage_opamp_dummy_magic_16_0.VD2.t20 GNDA.t212 GNDA.t213 GNDA.t202 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X649 two_stage_opamp_dummy_magic_16_0.VD3.t28 VDDA.t277 VDDA.t279 VDDA.t278 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X650 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t1 a_5980_2720.t1 GNDA.t296 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X651 VOUT-.t133 two_stage_opamp_dummy_magic_16_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X652 VOUT-.t10 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t8 GNDA.t101 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X653 two_stage_opamp_dummy_magic_16_0.VD3.t13 two_stage_opamp_dummy_magic_16_0.Vb2.t30 two_stage_opamp_dummy_magic_16_0.X.t14 two_stage_opamp_dummy_magic_16_0.VD3.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X654 bgr_0.V_TOP.t45 VDDA.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X655 bgr_0.V_mir2.t1 bgr_0.V_mir2.t0 VDDA.t220 VDDA.t219 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X656 VDDA.t16 bgr_0.V_mir1.t2 bgr_0.V_mir1.t3 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X657 VDDA.t27 two_stage_opamp_dummy_magic_16_0.Y.t49 VOUT+.t0 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X658 VOUT-.t134 two_stage_opamp_dummy_magic_16_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X659 two_stage_opamp_dummy_magic_16_0.X.t16 two_stage_opamp_dummy_magic_16_0.Vb1.t32 two_stage_opamp_dummy_magic_16_0.VD1.t3 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X660 VOUT-.t135 two_stage_opamp_dummy_magic_16_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X661 VOUT-.t136 two_stage_opamp_dummy_magic_16_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X662 bgr_0.V_mir2.t14 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t11 bgr_0.V_p_2.t0 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X663 VOUT+.t135 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X664 VOUT+.t136 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X665 bgr_0.PFET_GATE_10uA.t7 VDDA.t417 GNDA.t133 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X666 two_stage_opamp_dummy_magic_16_0.Y.t2 two_stage_opamp_dummy_magic_16_0.Vb1.t33 two_stage_opamp_dummy_magic_16_0.VD2.t7 GNDA.t303 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X667 VOUT+.t137 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X668 bgr_0.1st_Vout_1.t33 bgr_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X669 VOUT-.t137 two_stage_opamp_dummy_magic_16_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X670 two_stage_opamp_dummy_magic_16_0.Vb1.t0 bgr_0.PFET_GATE_10uA.t27 VDDA.t85 VDDA.t84 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X671 VDDA.t36 bgr_0.V_TOP.t46 bgr_0.Vin-.t3 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X672 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t1 two_stage_opamp_dummy_magic_16_0.Y.t50 VDDA.t203 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X673 VOUT+.t138 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X674 VOUT-.t11 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t9 GNDA.t138 GNDA.t137 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X675 VDDA.t72 two_stage_opamp_dummy_magic_16_0.X.t51 VOUT-.t2 VDDA.t71 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X676 VOUT-.t138 two_stage_opamp_dummy_magic_16_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X677 bgr_0.PFET_GATE_10uA.t2 bgr_0.1st_Vout_2.t33 VDDA.t404 VDDA.t403 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X678 two_stage_opamp_dummy_magic_16_0.VD3.t18 two_stage_opamp_dummy_magic_16_0.Vb3.t28 VDDA.t223 VDDA.t222 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X679 VOUT+.t139 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X680 VDDA.t193 bgr_0.PFET_GATE_10uA.t28 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t10 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X681 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t14 VDDA.t274 VDDA.t276 VDDA.t275 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X682 VOUT-.t139 two_stage_opamp_dummy_magic_16_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X683 GNDA.t150 two_stage_opamp_dummy_magic_16_0.Y.t51 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t1 VDDA.t214 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X684 VOUT-.t140 two_stage_opamp_dummy_magic_16_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X685 VOUT+.t140 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X686 GNDA.t322 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t29 two_stage_opamp_dummy_magic_16_0.V_source.t8 GNDA.t321 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X687 VDDA.t18 bgr_0.1st_Vout_2.t34 bgr_0.PFET_GATE_10uA.t1 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X688 VOUT+.t141 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X689 VOUT+.t142 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X690 VOUT+.t143 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X691 VOUT+.t144 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X692 bgr_0.1st_Vout_1.t34 bgr_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X693 bgr_0.1st_Vout_2.t35 bgr_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X694 VOUT-.t141 two_stage_opamp_dummy_magic_16_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X695 bgr_0.V_mir2.t13 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t12 bgr_0.V_p_2.t1 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X696 two_stage_opamp_dummy_magic_16_0.VD1.t20 VIN-.t9 two_stage_opamp_dummy_magic_16_0.V_source.t39 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X697 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t0 two_stage_opamp_dummy_magic_16_0.X.t52 VDDA.t146 GNDA.t88 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X698 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t11 bgr_0.NFET_GATE_10uA.t23 GNDA.t156 GNDA.t155 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X699 GNDA.t89 two_stage_opamp_dummy_magic_16_0.X.t53 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t1 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X700 VOUT-.t142 two_stage_opamp_dummy_magic_16_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X701 VOUT-.t143 two_stage_opamp_dummy_magic_16_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X702 two_stage_opamp_dummy_magic_16_0.V_source.t7 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t30 GNDA.t23 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X703 GNDA.t211 GNDA.t210 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X704 VOUT-.t144 two_stage_opamp_dummy_magic_16_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X705 GNDA.t147 two_stage_opamp_dummy_magic_16_0.X.t54 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t0 VDDA.t209 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X706 VOUT+.t145 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X707 bgr_0.1st_Vout_1.t35 bgr_0.cap_res1.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X708 VOUT-.t145 two_stage_opamp_dummy_magic_16_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X709 VDDA.t179 bgr_0.1st_Vout_1.t36 bgr_0.V_TOP.t5 VDDA.t178 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X710 VDDA.t383 two_stage_opamp_dummy_magic_16_0.V_err_gate.t9 two_stage_opamp_dummy_magic_16_0.V_err_p.t0 VDDA.t382 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X711 two_stage_opamp_dummy_magic_16_0.VD1.t18 VIN-.t10 two_stage_opamp_dummy_magic_16_0.V_source.t35 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X712 GNDA.t134 VDDA.t418 bgr_0.V_TOP.t7 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X713 bgr_0.V_TOP.t47 VDDA.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X714 VOUT-.t146 two_stage_opamp_dummy_magic_16_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X715 VDDA.t98 bgr_0.V_TOP.t48 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t2 VDDA.t97 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X716 VOUT+.t146 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X717 VOUT+.t147 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X718 VDDA.t95 two_stage_opamp_dummy_magic_16_0.Y.t52 VOUT+.t2 VDDA.t94 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X719 VOUT+.t148 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X720 VOUT-.t147 two_stage_opamp_dummy_magic_16_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X721 two_stage_opamp_dummy_magic_16_0.Vb2_2.t2 two_stage_opamp_dummy_magic_16_0.Vb2_2.t0 two_stage_opamp_dummy_magic_16_0.Vb2_2.t2 two_stage_opamp_dummy_magic_16_0.Vb2_2.t1 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X722 two_stage_opamp_dummy_magic_16_0.Y.t0 two_stage_opamp_dummy_magic_16_0.VD4.t12 two_stage_opamp_dummy_magic_16_0.VD4.t14 two_stage_opamp_dummy_magic_16_0.VD4.t13 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X723 two_stage_opamp_dummy_magic_16_0.X.t19 GNDA.t207 GNDA.t209 GNDA.t208 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X724 VOUT-.t148 two_stage_opamp_dummy_magic_16_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X725 two_stage_opamp_dummy_magic_16_0.X.t22 two_stage_opamp_dummy_magic_16_0.Vb1.t34 two_stage_opamp_dummy_magic_16_0.VD1.t2 GNDA.t301 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X726 bgr_0.V_mir2.t12 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t13 bgr_0.V_p_2.t4 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X727 VOUT+.t149 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X728 VDDA.t191 bgr_0.PFET_GATE_10uA.t29 bgr_0.V_CUR_REF_REG.t0 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X729 VOUT+.t150 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X730 VOUT-.t149 two_stage_opamp_dummy_magic_16_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X731 VOUT+.t151 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X732 GNDA.t206 GNDA.t204 two_stage_opamp_dummy_magic_16_0.VD1.t17 GNDA.t205 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X733 VOUT-.t150 two_stage_opamp_dummy_magic_16_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X734 two_stage_opamp_dummy_magic_16_0.Y.t13 GNDA.t201 GNDA.t203 GNDA.t202 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X735 VOUT-.t151 two_stage_opamp_dummy_magic_16_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X736 VOUT+.t152 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X737 VOUT-.t152 two_stage_opamp_dummy_magic_16_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X738 VOUT-.t153 two_stage_opamp_dummy_magic_16_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X739 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t0 two_stage_opamp_dummy_magic_16_0.Y.t53 VDDA.t40 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X740 GNDA.t200 GNDA.t198 VDDA.t264 GNDA.t199 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X741 GNDA.t197 GNDA.t195 two_stage_opamp_dummy_magic_16_0.VD1.t16 GNDA.t196 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X742 bgr_0.V_TOP.t49 VDDA.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X743 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t0 VDDA.t268 VDDA.t270 VDDA.t269 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X744 two_stage_opamp_dummy_magic_16_0.Vb3.t7 two_stage_opamp_dummy_magic_16_0.Vb2.t31 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t10 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t9 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X745 two_stage_opamp_dummy_magic_16_0.X.t10 two_stage_opamp_dummy_magic_16_0.VD3.t30 two_stage_opamp_dummy_magic_16_0.VD3.t32 two_stage_opamp_dummy_magic_16_0.VD3.t31 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X746 VOUT+.t153 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X747 VOUT-.t154 two_stage_opamp_dummy_magic_16_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X748 VOUT+.t154 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X749 VOUT-.t155 two_stage_opamp_dummy_magic_16_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X750 bgr_0.1st_Vout_2.t36 bgr_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X751 GNDA.t106 two_stage_opamp_dummy_magic_16_0.Y.t54 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t0 VDDA.t166 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X752 VDDA.t81 bgr_0.V_mir1.t0 bgr_0.V_mir1.t1 VDDA.t80 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X753 VOUT+.t155 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X754 two_stage_opamp_dummy_magic_16_0.Y.t24 two_stage_opamp_dummy_magic_16_0.Vb2.t32 two_stage_opamp_dummy_magic_16_0.VD4.t19 two_stage_opamp_dummy_magic_16_0.VD4.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X755 VOUT+.t156 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X756 GNDA.t309 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t31 two_stage_opamp_dummy_magic_16_0.V_p_mir.t1 GNDA.t308 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X757 VOUT-.t156 two_stage_opamp_dummy_magic_16_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.t2 384.967
R1 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t10 369.534
R2 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t22 369.534
R3 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t7 369.534
R4 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t16 369.534
R5 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t12 369.534
R6 bgr_0.NFET_GATE_10uA.t2 bgr_0.NFET_GATE_10uA.n18 369.534
R7 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n20 366.553
R8 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.t9 192.8
R9 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.t17 192.8
R10 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t23 192.8
R11 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t11 192.8
R12 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t20 192.8
R13 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t21 192.8
R14 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.t8 192.8
R15 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.t15 192.8
R16 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.t19 192.8
R17 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.t5 192.8
R18 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t13 192.8
R19 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.t18 192.8
R20 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.t6 192.8
R21 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.t14 192.8
R22 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.n11 176.733
R23 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.n10 176.733
R24 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.n4 176.733
R25 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.n5 176.733
R26 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.n2 176.733
R27 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.n1 176.733
R28 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.n17 176.733
R29 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.n16 176.733
R30 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n13 169.852
R31 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n8 169.852
R32 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n14 166.133
R33 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.n0 126.877
R34 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n12 56.2338
R35 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n9 56.2338
R36 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n7 56.2338
R37 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n6 56.2338
R38 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n3 56.2338
R39 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.n15 56.2338
R40 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t1 39.4005
R41 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t0 39.4005
R42 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n19 30.6442
R43 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t4 24.0005
R44 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t3 24.0005
R45 two_stage_opamp_dummy_magic_16_0.Vb3.n25 two_stage_opamp_dummy_magic_16_0.Vb3.t14 650.511
R46 two_stage_opamp_dummy_magic_16_0.Vb3.n19 two_stage_opamp_dummy_magic_16_0.Vb3.t13 611.739
R47 two_stage_opamp_dummy_magic_16_0.Vb3.n15 two_stage_opamp_dummy_magic_16_0.Vb3.t22 611.739
R48 two_stage_opamp_dummy_magic_16_0.Vb3.n10 two_stage_opamp_dummy_magic_16_0.Vb3.t8 611.739
R49 two_stage_opamp_dummy_magic_16_0.Vb3.n6 two_stage_opamp_dummy_magic_16_0.Vb3.t16 611.739
R50 two_stage_opamp_dummy_magic_16_0.Vb3.n19 two_stage_opamp_dummy_magic_16_0.Vb3.t19 421.75
R51 two_stage_opamp_dummy_magic_16_0.Vb3.n20 two_stage_opamp_dummy_magic_16_0.Vb3.t23 421.75
R52 two_stage_opamp_dummy_magic_16_0.Vb3.n21 two_stage_opamp_dummy_magic_16_0.Vb3.t26 421.75
R53 two_stage_opamp_dummy_magic_16_0.Vb3.n22 two_stage_opamp_dummy_magic_16_0.Vb3.t25 421.75
R54 two_stage_opamp_dummy_magic_16_0.Vb3.n15 two_stage_opamp_dummy_magic_16_0.Vb3.t24 421.75
R55 two_stage_opamp_dummy_magic_16_0.Vb3.n16 two_stage_opamp_dummy_magic_16_0.Vb3.t20 421.75
R56 two_stage_opamp_dummy_magic_16_0.Vb3.n17 two_stage_opamp_dummy_magic_16_0.Vb3.t15 421.75
R57 two_stage_opamp_dummy_magic_16_0.Vb3.n18 two_stage_opamp_dummy_magic_16_0.Vb3.t10 421.75
R58 two_stage_opamp_dummy_magic_16_0.Vb3.n10 two_stage_opamp_dummy_magic_16_0.Vb3.t11 421.75
R59 two_stage_opamp_dummy_magic_16_0.Vb3.n11 two_stage_opamp_dummy_magic_16_0.Vb3.t17 421.75
R60 two_stage_opamp_dummy_magic_16_0.Vb3.n12 two_stage_opamp_dummy_magic_16_0.Vb3.t21 421.75
R61 two_stage_opamp_dummy_magic_16_0.Vb3.n13 two_stage_opamp_dummy_magic_16_0.Vb3.t27 421.75
R62 two_stage_opamp_dummy_magic_16_0.Vb3.n6 two_stage_opamp_dummy_magic_16_0.Vb3.t18 421.75
R63 two_stage_opamp_dummy_magic_16_0.Vb3.n7 two_stage_opamp_dummy_magic_16_0.Vb3.t12 421.75
R64 two_stage_opamp_dummy_magic_16_0.Vb3.n8 two_stage_opamp_dummy_magic_16_0.Vb3.t9 421.75
R65 two_stage_opamp_dummy_magic_16_0.Vb3.n9 two_stage_opamp_dummy_magic_16_0.Vb3.t28 421.75
R66 two_stage_opamp_dummy_magic_16_0.Vb3.n24 two_stage_opamp_dummy_magic_16_0.Vb3.n23 176.185
R67 two_stage_opamp_dummy_magic_16_0.Vb3.n24 two_stage_opamp_dummy_magic_16_0.Vb3.n14 175.624
R68 two_stage_opamp_dummy_magic_16_0.Vb3.n20 two_stage_opamp_dummy_magic_16_0.Vb3.n19 167.094
R69 two_stage_opamp_dummy_magic_16_0.Vb3.n21 two_stage_opamp_dummy_magic_16_0.Vb3.n20 167.094
R70 two_stage_opamp_dummy_magic_16_0.Vb3.n22 two_stage_opamp_dummy_magic_16_0.Vb3.n21 167.094
R71 two_stage_opamp_dummy_magic_16_0.Vb3.n16 two_stage_opamp_dummy_magic_16_0.Vb3.n15 167.094
R72 two_stage_opamp_dummy_magic_16_0.Vb3.n17 two_stage_opamp_dummy_magic_16_0.Vb3.n16 167.094
R73 two_stage_opamp_dummy_magic_16_0.Vb3.n18 two_stage_opamp_dummy_magic_16_0.Vb3.n17 167.094
R74 two_stage_opamp_dummy_magic_16_0.Vb3.n11 two_stage_opamp_dummy_magic_16_0.Vb3.n10 167.094
R75 two_stage_opamp_dummy_magic_16_0.Vb3.n12 two_stage_opamp_dummy_magic_16_0.Vb3.n11 167.094
R76 two_stage_opamp_dummy_magic_16_0.Vb3.n13 two_stage_opamp_dummy_magic_16_0.Vb3.n12 167.094
R77 two_stage_opamp_dummy_magic_16_0.Vb3.n7 two_stage_opamp_dummy_magic_16_0.Vb3.n6 167.094
R78 two_stage_opamp_dummy_magic_16_0.Vb3.n8 two_stage_opamp_dummy_magic_16_0.Vb3.n7 167.094
R79 two_stage_opamp_dummy_magic_16_0.Vb3.n9 two_stage_opamp_dummy_magic_16_0.Vb3.n8 167.094
R80 two_stage_opamp_dummy_magic_16_0.Vb3.n26 two_stage_opamp_dummy_magic_16_0.Vb3.n5 161.631
R81 two_stage_opamp_dummy_magic_16_0.Vb3.n2 two_stage_opamp_dummy_magic_16_0.Vb3.n0 139.639
R82 two_stage_opamp_dummy_magic_16_0.Vb3.n2 two_stage_opamp_dummy_magic_16_0.Vb3.n1 139.638
R83 two_stage_opamp_dummy_magic_16_0.Vb3.n4 two_stage_opamp_dummy_magic_16_0.Vb3.n3 134.577
R84 two_stage_opamp_dummy_magic_16_0.Vb3.n23 two_stage_opamp_dummy_magic_16_0.Vb3.n22 49.8072
R85 two_stage_opamp_dummy_magic_16_0.Vb3.n23 two_stage_opamp_dummy_magic_16_0.Vb3.n18 49.8072
R86 two_stage_opamp_dummy_magic_16_0.Vb3.n14 two_stage_opamp_dummy_magic_16_0.Vb3.n13 49.8072
R87 two_stage_opamp_dummy_magic_16_0.Vb3.n14 two_stage_opamp_dummy_magic_16_0.Vb3.n9 49.8072
R88 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_16_0.Vb3.n26 48.0943
R89 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_16_0.Vb3.n4 41.063
R90 two_stage_opamp_dummy_magic_16_0.Vb3.n3 two_stage_opamp_dummy_magic_16_0.Vb3.t4 24.0005
R91 two_stage_opamp_dummy_magic_16_0.Vb3.n3 two_stage_opamp_dummy_magic_16_0.Vb3.t3 24.0005
R92 two_stage_opamp_dummy_magic_16_0.Vb3.n1 two_stage_opamp_dummy_magic_16_0.Vb3.t5 24.0005
R93 two_stage_opamp_dummy_magic_16_0.Vb3.n1 two_stage_opamp_dummy_magic_16_0.Vb3.t0 24.0005
R94 two_stage_opamp_dummy_magic_16_0.Vb3.n0 two_stage_opamp_dummy_magic_16_0.Vb3.t2 24.0005
R95 two_stage_opamp_dummy_magic_16_0.Vb3.n0 two_stage_opamp_dummy_magic_16_0.Vb3.t6 24.0005
R96 two_stage_opamp_dummy_magic_16_0.Vb3.n25 two_stage_opamp_dummy_magic_16_0.Vb3.n24 13.7349
R97 two_stage_opamp_dummy_magic_16_0.Vb3.n5 two_stage_opamp_dummy_magic_16_0.Vb3.t1 11.2576
R98 two_stage_opamp_dummy_magic_16_0.Vb3.n5 two_stage_opamp_dummy_magic_16_0.Vb3.t7 11.2576
R99 two_stage_opamp_dummy_magic_16_0.Vb3.n4 two_stage_opamp_dummy_magic_16_0.Vb3.n2 4.5005
R100 two_stage_opamp_dummy_magic_16_0.Vb3.n26 two_stage_opamp_dummy_magic_16_0.Vb3.n25 1.438
R101 GNDA.n385 GNDA.n8 21966.8
R102 GNDA.n505 GNDA.n14 21966.8
R103 GNDA.n923 GNDA.n922 15367.3
R104 GNDA.n2582 GNDA.n8 14081.2
R105 GNDA.n507 GNDA.n12 13534.7
R106 GNDA.n10 GNDA.n9 13528.5
R107 GNDA.n11 GNDA.n7 13200
R108 GNDA.n921 GNDA.n920 12810.6
R109 GNDA.n924 GNDA.n923 11953.3
R110 GNDA.n924 GNDA.n510 11890.5
R111 GNDA.n2583 GNDA.n7 11824
R112 GNDA.n13 GNDA.n7 11671.2
R113 GNDA.n11 GNDA.n9 11178.4
R114 GNDA.n2582 GNDA.n2581 11146.8
R115 GNDA.n918 GNDA.n510 9950.42
R116 GNDA.n923 GNDA.n920 9950.42
R117 GNDA.n2581 GNDA.n9 9632.43
R118 GNDA.n919 GNDA.n918 9384.59
R119 GNDA.n920 GNDA.n919 9384.59
R120 GNDA.n2581 GNDA.n2580 9001.83
R121 GNDA.n506 GNDA.n13 7758.44
R122 GNDA.n509 GNDA.n508 7427.52
R123 GNDA.n12 GNDA.n10 4761.61
R124 GNDA.n2578 GNDA.n510 4448.89
R125 GNDA.n925 GNDA.n924 3974.19
R126 GNDA.n12 GNDA.n11 3961.87
R127 GNDA.n2580 GNDA.t11 3375.81
R128 GNDA.n919 GNDA.n508 3105.87
R129 GNDA.n2580 GNDA.n508 2321.1
R130 GNDA.n508 GNDA.n10 2315.79
R131 GNDA.n505 GNDA.t44 2006.86
R132 GNDA.n2580 GNDA.n2579 2001.83
R133 GNDA.n2583 GNDA.n2582 1965.05
R134 GNDA.n508 GNDA.n507 1779.93
R135 GNDA.n922 GNDA.n921 1460.18
R136 GNDA.n506 GNDA.t85 1440.97
R137 GNDA.n918 GNDA.n509 1440.71
R138 GNDA.n2579 GNDA.n509 1440.71
R139 GNDA.n1804 GNDA.n1803 1336.64
R140 GNDA.n2578 GNDA.t151 1258.74
R141 GNDA.n1829 GNDA.n1223 1214.72
R142 GNDA.n1835 GNDA.n1223 1214.72
R143 GNDA.n1836 GNDA.n1835 1214.72
R144 GNDA.n1836 GNDA.n1219 1214.72
R145 GNDA.n1842 GNDA.n1219 1214.72
R146 GNDA.n1844 GNDA.n1214 1214.72
R147 GNDA.n1850 GNDA.n1214 1214.72
R148 GNDA.n1851 GNDA.n1850 1214.72
R149 GNDA.n1851 GNDA.n1210 1214.72
R150 GNDA.n1857 GNDA.n1210 1214.72
R151 GNDA.n802 GNDA.n512 1212.88
R152 GNDA.n1016 GNDA.n1015 1185.07
R153 GNDA.n1017 GNDA.n1016 1185.07
R154 GNDA.n921 GNDA.n508 1167.58
R155 GNDA.n922 GNDA.t74 1012.83
R156 GNDA.n2579 GNDA.n2578 869.924
R157 GNDA.n1842 GNDA.t211 823.313
R158 GNDA.n491 GNDA.t245 762.534
R159 GNDA.n493 GNDA.t219 762.534
R160 GNDA.n367 GNDA.t198 762.534
R161 GNDA.n365 GNDA.t214 762.534
R162 GNDA.t85 GNDA.n505 702.521
R163 GNDA.n361 GNDA.n360 692.506
R164 GNDA.n377 GNDA.n376 692.506
R165 GNDA.n487 GNDA.n486 692.506
R166 GNDA.n503 GNDA.n502 692.506
R167 GNDA.n348 GNDA.n347 692.506
R168 GNDA.n287 GNDA.n284 692.506
R169 GNDA.n119 GNDA.n118 692.506
R170 GNDA.n58 GNDA.n55 692.506
R171 GNDA.n2566 GNDA.n2565 686.717
R172 GNDA.n453 GNDA.n452 686.717
R173 GNDA.n432 GNDA.n431 686.717
R174 GNDA.n382 GNDA.n381 686.717
R175 GNDA.n403 GNDA.n402 686.717
R176 GNDA.n224 GNDA.n223 686.717
R177 GNDA.n212 GNDA.n123 686.717
R178 GNDA.n153 GNDA.n152 686.717
R179 GNDA.n202 GNDA.n201 686.717
R180 GNDA.n2594 GNDA.n2593 686.717
R181 GNDA.n136 GNDA.n135 686.717
R182 GNDA.n2569 GNDA.n512 686.717
R183 GNDA.n2569 GNDA.n511 686.717
R184 GNDA.n205 GNDA.n204 686.717
R185 GNDA.n160 GNDA.n159 686.717
R186 GNDA.n475 GNDA.n468 686.717
R187 GNDA.n463 GNDA.n462 686.717
R188 GNDA.n406 GNDA.n405 686.717
R189 GNDA.n392 GNDA.n384 686.717
R190 GNDA.n439 GNDA.n438 686.717
R191 GNDA.n445 GNDA.n138 686.717
R192 GNDA.n2557 GNDA.n523 686.717
R193 GNDA.n2364 GNDA.n2353 686.717
R194 GNDA.n161 GNDA.t222 682.201
R195 GNDA.n440 GNDA.t276 674.168
R196 GNDA.n444 GNDA.t227 674.168
R197 GNDA.n1439 GNDA.n1435 669.307
R198 GNDA.n206 GNDA.t281 650.067
R199 GNDA.n2463 GNDA.n2462 585.001
R200 GNDA.n2483 GNDA.n2482 585.001
R201 GNDA.n2477 GNDA.n558 585.001
R202 GNDA.n2515 GNDA.n2514 585.001
R203 GNDA.n2525 GNDA.n2524 585.001
R204 GNDA.n2576 GNDA.n2575 585.001
R205 GNDA.n2313 GNDA.n2312 585
R206 GNDA.n2311 GNDA.n2274 585
R207 GNDA.n2310 GNDA.n2309 585
R208 GNDA.n2308 GNDA.n2307 585
R209 GNDA.n2306 GNDA.n2305 585
R210 GNDA.n2304 GNDA.n2303 585
R211 GNDA.n2302 GNDA.n2301 585
R212 GNDA.n2300 GNDA.n2299 585
R213 GNDA.n2298 GNDA.n2297 585
R214 GNDA.n2296 GNDA.n2295 585
R215 GNDA.n614 GNDA.n613 585
R216 GNDA.n2315 GNDA.n614 585
R217 GNDA.n2318 GNDA.n2317 585
R218 GNDA.n2318 GNDA.n611 585
R219 GNDA.n1505 GNDA.n1504 585
R220 GNDA.n1503 GNDA.n1502 585
R221 GNDA.n1501 GNDA.n1500 585
R222 GNDA.n1499 GNDA.n1498 585
R223 GNDA.n1497 GNDA.n1496 585
R224 GNDA.n1495 GNDA.n1494 585
R225 GNDA.n1493 GNDA.n1492 585
R226 GNDA.n1491 GNDA.n1490 585
R227 GNDA.n1489 GNDA.n1488 585
R228 GNDA.n1487 GNDA.n1486 585
R229 GNDA.n1485 GNDA.n621 585
R230 GNDA.n2315 GNDA.n621 585
R231 GNDA.n1267 GNDA.n1266 585
R232 GNDA.n1267 GNDA.n1265 585
R233 GNDA.n2315 GNDA.n2269 585
R234 GNDA.n1102 GNDA.n1101 585
R235 GNDA.n1100 GNDA.n1099 585
R236 GNDA.n1098 GNDA.n1097 585
R237 GNDA.n1096 GNDA.n1095 585
R238 GNDA.n1094 GNDA.n1093 585
R239 GNDA.n1092 GNDA.n1091 585
R240 GNDA.n1090 GNDA.n1089 585
R241 GNDA.n1088 GNDA.n1087 585
R242 GNDA.n1086 GNDA.n1085 585
R243 GNDA.n1084 GNDA.n1083 585
R244 GNDA.n1082 GNDA.n1081 585
R245 GNDA.n1856 GNDA.n1209 585
R246 GNDA.n1857 GNDA.n1856 585
R247 GNDA.n1855 GNDA.n1854 585
R248 GNDA.n1855 GNDA.n1210 585
R249 GNDA.n1853 GNDA.n1211 585
R250 GNDA.n1851 GNDA.n1211 585
R251 GNDA.n1849 GNDA.n1212 585
R252 GNDA.n1850 GNDA.n1849 585
R253 GNDA.n1848 GNDA.n1847 585
R254 GNDA.n1848 GNDA.n1214 585
R255 GNDA.n1216 GNDA.n1215 585
R256 GNDA.n1844 GNDA.n1215 585
R257 GNDA.n1841 GNDA.n1218 585
R258 GNDA.n1842 GNDA.n1841 585
R259 GNDA.n1840 GNDA.n1839 585
R260 GNDA.n1840 GNDA.n1219 585
R261 GNDA.n1838 GNDA.n1220 585
R262 GNDA.n1836 GNDA.n1220 585
R263 GNDA.n1834 GNDA.n1221 585
R264 GNDA.n1835 GNDA.n1834 585
R265 GNDA.n1833 GNDA.n1832 585
R266 GNDA.n1833 GNDA.n1223 585
R267 GNDA.n1225 GNDA.n1224 585
R268 GNDA.n1829 GNDA.n1224 585
R269 GNDA.n1830 GNDA.n1225 585
R270 GNDA.n1830 GNDA.n1829 585
R271 GNDA.n1832 GNDA.n1831 585
R272 GNDA.n1831 GNDA.n1223 585
R273 GNDA.n1222 GNDA.n1221 585
R274 GNDA.n1835 GNDA.n1222 585
R275 GNDA.n1838 GNDA.n1837 585
R276 GNDA.n1837 GNDA.n1836 585
R277 GNDA.n1839 GNDA.n1217 585
R278 GNDA.n1219 GNDA.n1217 585
R279 GNDA.n1843 GNDA.n1218 585
R280 GNDA.n1843 GNDA.n1842 585
R281 GNDA.n1845 GNDA.n1216 585
R282 GNDA.n1845 GNDA.n1844 585
R283 GNDA.n1847 GNDA.n1846 585
R284 GNDA.n1846 GNDA.n1214 585
R285 GNDA.n1213 GNDA.n1212 585
R286 GNDA.n1850 GNDA.n1213 585
R287 GNDA.n1853 GNDA.n1852 585
R288 GNDA.n1852 GNDA.n1851 585
R289 GNDA.n1854 GNDA.n1208 585
R290 GNDA.n1210 GNDA.n1208 585
R291 GNDA.n1858 GNDA.n1209 585
R292 GNDA.n1858 GNDA.n1857 585
R293 GNDA.n2189 GNDA.n1050 585
R294 GNDA.n2192 GNDA.n2191 585
R295 GNDA.n1054 GNDA.n1053 585
R296 GNDA.n1899 GNDA.n1898 585
R297 GNDA.n1900 GNDA.n1897 585
R298 GNDA.n1894 GNDA.n1893 585
R299 GNDA.n1906 GNDA.n1892 585
R300 GNDA.n1907 GNDA.n1891 585
R301 GNDA.n1908 GNDA.n1890 585
R302 GNDA.n1888 GNDA.n1887 585
R303 GNDA.n1913 GNDA.n1886 585
R304 GNDA.n1914 GNDA.n1885 585
R305 GNDA.n1915 GNDA.n1914 585
R306 GNDA.n1913 GNDA.n1912 585
R307 GNDA.n1911 GNDA.n1888 585
R308 GNDA.n1909 GNDA.n1908 585
R309 GNDA.n1907 GNDA.n1889 585
R310 GNDA.n1906 GNDA.n1905 585
R311 GNDA.n1903 GNDA.n1894 585
R312 GNDA.n1901 GNDA.n1900 585
R313 GNDA.n1899 GNDA.n1896 585
R314 GNDA.n1053 GNDA.n1052 585
R315 GNDA.n2193 GNDA.n2192 585
R316 GNDA.n2195 GNDA.n1050 585
R317 GNDA.n2185 GNDA.n2184 585
R318 GNDA.n1123 GNDA.n1079 585
R319 GNDA.n1122 GNDA.n1121 585
R320 GNDA.n1120 GNDA.n1119 585
R321 GNDA.n1118 GNDA.n1117 585
R322 GNDA.n1116 GNDA.n1115 585
R323 GNDA.n1114 GNDA.n1113 585
R324 GNDA.n1112 GNDA.n1111 585
R325 GNDA.n1110 GNDA.n1109 585
R326 GNDA.n1108 GNDA.n1107 585
R327 GNDA.n1106 GNDA.n1105 585
R328 GNDA.n1104 GNDA.n1103 585
R329 GNDA.n1884 GNDA.n1883 585
R330 GNDA.n1882 GNDA.n1881 585
R331 GNDA.n1880 GNDA.n1879 585
R332 GNDA.n1878 GNDA.n1877 585
R333 GNDA.n1876 GNDA.n1875 585
R334 GNDA.n1874 GNDA.n1873 585
R335 GNDA.n1872 GNDA.n1871 585
R336 GNDA.n1870 GNDA.n1869 585
R337 GNDA.n1868 GNDA.n1867 585
R338 GNDA.n1866 GNDA.n1865 585
R339 GNDA.n1864 GNDA.n1863 585
R340 GNDA.n1127 GNDA.n1124 585
R341 GNDA.n1939 GNDA.n1938 585
R342 GNDA.n1937 GNDA.n1936 585
R343 GNDA.n1935 GNDA.n1934 585
R344 GNDA.n1933 GNDA.n1932 585
R345 GNDA.n1931 GNDA.n1930 585
R346 GNDA.n1929 GNDA.n1928 585
R347 GNDA.n1927 GNDA.n1926 585
R348 GNDA.n1925 GNDA.n1924 585
R349 GNDA.n1923 GNDA.n1922 585
R350 GNDA.n1921 GNDA.n1920 585
R351 GNDA.n1919 GNDA.n1918 585
R352 GNDA.n1917 GNDA.n1916 585
R353 GNDA.n1654 GNDA.n1653 585
R354 GNDA.n1651 GNDA.n1264 585
R355 GNDA.n1270 GNDA.n1269 585
R356 GNDA.n1646 GNDA.n1645 585
R357 GNDA.n1644 GNDA.n1643 585
R358 GNDA.n1570 GNDA.n1274 585
R359 GNDA.n1572 GNDA.n1571 585
R360 GNDA.n1577 GNDA.n1576 585
R361 GNDA.n1575 GNDA.n1568 585
R362 GNDA.n1583 GNDA.n1582 585
R363 GNDA.n1585 GNDA.n1584 585
R364 GNDA.n1566 GNDA.n1565 585
R365 GNDA.n1860 GNDA.n1205 585
R366 GNDA.n1206 GNDA.n1205 585
R367 GNDA.n1411 GNDA.n1410 585
R368 GNDA.n1408 GNDA.n1407 585
R369 GNDA.n1406 GNDA.n1405 585
R370 GNDA.n1322 GNDA.n1298 585
R371 GNDA.n1324 GNDA.n1323 585
R372 GNDA.n1328 GNDA.n1327 585
R373 GNDA.n1330 GNDA.n1329 585
R374 GNDA.n1337 GNDA.n1336 585
R375 GNDA.n1335 GNDA.n1320 585
R376 GNDA.n1343 GNDA.n1342 585
R377 GNDA.n1345 GNDA.n1344 585
R378 GNDA.n1318 GNDA.n1317 585
R379 GNDA.n1860 GNDA.n1859 585
R380 GNDA.n1859 GNDA.n1206 585
R381 GNDA.n1733 GNDA.n1207 585
R382 GNDA.n1734 GNDA.n1670 585
R383 GNDA.n1744 GNDA.n1743 585
R384 GNDA.n1746 GNDA.n1668 585
R385 GNDA.n1749 GNDA.n1748 585
R386 GNDA.n1750 GNDA.n1664 585
R387 GNDA.n1759 GNDA.n1758 585
R388 GNDA.n1761 GNDA.n1663 585
R389 GNDA.n1764 GNDA.n1763 585
R390 GNDA.n1765 GNDA.n1657 585
R391 GNDA.n1774 GNDA.n1773 585
R392 GNDA.n1776 GNDA.n1251 585
R393 GNDA.n1806 GNDA.n1805 585
R394 GNDA.n1805 GNDA.n1804 585
R395 GNDA.n1807 GNDA.n1238 585
R396 GNDA.n1238 GNDA.n1237 585
R397 GNDA.n1809 GNDA.n1808 585
R398 GNDA.n1810 GNDA.n1809 585
R399 GNDA.n1235 GNDA.n1234 585
R400 GNDA.n1811 GNDA.n1235 585
R401 GNDA.n1814 GNDA.n1813 585
R402 GNDA.n1813 GNDA.n1812 585
R403 GNDA.n1815 GNDA.n1233 585
R404 GNDA.n1236 GNDA.n1233 585
R405 GNDA.n1817 GNDA.n1816 585
R406 GNDA.n1818 GNDA.n1817 585
R407 GNDA.n1232 GNDA.n1231 585
R408 GNDA.n1819 GNDA.n1232 585
R409 GNDA.n1822 GNDA.n1821 585
R410 GNDA.n1821 GNDA.n1820 585
R411 GNDA.n1823 GNDA.n1229 585
R412 GNDA.n1229 GNDA.n1228 585
R413 GNDA.n1825 GNDA.n1824 585
R414 GNDA.n1826 GNDA.n1825 585
R415 GNDA.n1230 GNDA.n1226 585
R416 GNDA.n1827 GNDA.n1226 585
R417 GNDA.n1440 GNDA.n1436 585
R418 GNDA.n1442 GNDA.n1441 585
R419 GNDA.t211 GNDA.n1442 585
R420 GNDA.n1449 GNDA.n1448 585
R421 GNDA.n1449 GNDA.n1227 585
R422 GNDA.n1450 GNDA.n1446 585
R423 GNDA.n1451 GNDA.n1450 585
R424 GNDA.n1454 GNDA.n1453 585
R425 GNDA.n1453 GNDA.n1452 585
R426 GNDA.n1455 GNDA.n1444 585
R427 GNDA.n1444 GNDA.n1443 585
R428 GNDA.n1457 GNDA.n1456 585
R429 GNDA.n1458 GNDA.n1457 585
R430 GNDA.n1445 GNDA.n1434 585
R431 GNDA.n1459 GNDA.n1434 585
R432 GNDA.n1462 GNDA.n1461 585
R433 GNDA.n1461 GNDA.n1460 585
R434 GNDA.n1463 GNDA.n1432 585
R435 GNDA.n1432 GNDA.n1431 585
R436 GNDA.n1465 GNDA.n1464 585
R437 GNDA.n1466 GNDA.n1465 585
R438 GNDA.n1429 GNDA.n1428 585
R439 GNDA.n1467 GNDA.n1429 585
R440 GNDA.n1470 GNDA.n1469 585
R441 GNDA.n1469 GNDA.n1468 585
R442 GNDA.n1471 GNDA.n1427 585
R443 GNDA.n1430 GNDA.n1427 585
R444 GNDA.n1529 GNDA.n1474 585
R445 GNDA.n1529 GNDA.n1528 585
R446 GNDA.n1523 GNDA.n1473 585
R447 GNDA.n1527 GNDA.n1473 585
R448 GNDA.n1525 GNDA.n1524 585
R449 GNDA.n1526 GNDA.n1525 585
R450 GNDA.n1522 GNDA.n1476 585
R451 GNDA.n1476 GNDA.n1475 585
R452 GNDA.n1521 GNDA.n1520 585
R453 GNDA.n1520 GNDA.n1519 585
R454 GNDA.n1478 GNDA.n1477 585
R455 GNDA.n1518 GNDA.n1478 585
R456 GNDA.n1516 GNDA.n1515 585
R457 GNDA.n1517 GNDA.n1516 585
R458 GNDA.n1514 GNDA.n1480 585
R459 GNDA.n1480 GNDA.n1479 585
R460 GNDA.n1513 GNDA.n1512 585
R461 GNDA.n1512 GNDA.n1511 585
R462 GNDA.n1482 GNDA.n1481 585
R463 GNDA.n1510 GNDA.n1482 585
R464 GNDA.n1508 GNDA.n1507 585
R465 GNDA.n1509 GNDA.n1508 585
R466 GNDA.n1506 GNDA.n1484 585
R467 GNDA.n1484 GNDA.n1483 585
R468 GNDA.n1563 GNDA.n1562 585
R469 GNDA.n1551 GNDA.n1295 585
R470 GNDA.n1552 GNDA.n1414 585
R471 GNDA.n1555 GNDA.n1554 585
R472 GNDA.n1417 GNDA.n1416 585
R473 GNDA.n1548 GNDA.n1547 585
R474 GNDA.n1422 GNDA.n1421 585
R475 GNDA.n1541 GNDA.n1540 585
R476 GNDA.n1539 GNDA.n1538 585
R477 GNDA.n1537 GNDA.n1426 585
R478 GNDA.n1425 GNDA.n1424 585
R479 GNDA.n1531 GNDA.n1530 585
R480 GNDA.n1564 GNDA.n1125 585
R481 GNDA.n1564 GNDA.n1206 585
R482 GNDA.n1532 GNDA.n1531 585
R483 GNDA.n1534 GNDA.n1424 585
R484 GNDA.n1537 GNDA.n1536 585
R485 GNDA.n1538 GNDA.n1423 585
R486 GNDA.n1542 GNDA.n1541 585
R487 GNDA.n1544 GNDA.n1422 585
R488 GNDA.n1547 GNDA.n1546 585
R489 GNDA.n1416 GNDA.n1415 585
R490 GNDA.n1556 GNDA.n1555 585
R491 GNDA.n1558 GNDA.n1414 585
R492 GNDA.n1559 GNDA.n1295 585
R493 GNDA.n1562 GNDA.n1561 585
R494 GNDA.n1412 GNDA.n1125 585
R495 GNDA.n1412 GNDA.n1206 585
R496 GNDA.n2161 GNDA.n1149 585
R497 GNDA.n2162 GNDA.n1147 585
R498 GNDA.n2163 GNDA.n1146 585
R499 GNDA.n1144 GNDA.n1142 585
R500 GNDA.n2169 GNDA.n1141 585
R501 GNDA.n2170 GNDA.n1139 585
R502 GNDA.n2171 GNDA.n1138 585
R503 GNDA.n1136 GNDA.n1134 585
R504 GNDA.n2176 GNDA.n1133 585
R505 GNDA.n2177 GNDA.n1131 585
R506 GNDA.n1130 GNDA.n1126 585
R507 GNDA.n2182 GNDA.n1080 585
R508 GNDA.n2182 GNDA.n2181 585
R509 GNDA.n2179 GNDA.n1126 585
R510 GNDA.n2178 GNDA.n2177 585
R511 GNDA.n2176 GNDA.n2175 585
R512 GNDA.n2174 GNDA.n1134 585
R513 GNDA.n2172 GNDA.n2171 585
R514 GNDA.n2170 GNDA.n1135 585
R515 GNDA.n2169 GNDA.n2168 585
R516 GNDA.n2166 GNDA.n1142 585
R517 GNDA.n2164 GNDA.n2163 585
R518 GNDA.n2162 GNDA.n1143 585
R519 GNDA.n2161 GNDA.n2160 585
R520 GNDA.n2487 GNDA.n2486 585
R521 GNDA.n2488 GNDA.n604 585
R522 GNDA.n2489 GNDA.n603 585
R523 GNDA.n601 GNDA.n599 585
R524 GNDA.n2495 GNDA.n598 585
R525 GNDA.n2496 GNDA.n596 585
R526 GNDA.n2497 GNDA.n595 585
R527 GNDA.n593 GNDA.n591 585
R528 GNDA.n2502 GNDA.n590 585
R529 GNDA.n2503 GNDA.n588 585
R530 GNDA.n587 GNDA.n583 585
R531 GNDA.n2508 GNDA.n579 585
R532 GNDA.n2508 GNDA.n2507 585
R533 GNDA.n2505 GNDA.n583 585
R534 GNDA.n2504 GNDA.n2503 585
R535 GNDA.n2502 GNDA.n2501 585
R536 GNDA.n2500 GNDA.n591 585
R537 GNDA.n2498 GNDA.n2497 585
R538 GNDA.n2496 GNDA.n592 585
R539 GNDA.n2495 GNDA.n2494 585
R540 GNDA.n2492 GNDA.n599 585
R541 GNDA.n2490 GNDA.n2489 585
R542 GNDA.n2488 GNDA.n600 585
R543 GNDA.n2487 GNDA.n606 585
R544 GNDA.n1025 GNDA.n745 585
R545 GNDA.n1026 GNDA.n743 585
R546 GNDA.n1027 GNDA.n742 585
R547 GNDA.n740 GNDA.n738 585
R548 GNDA.n1033 GNDA.n737 585
R549 GNDA.n1034 GNDA.n735 585
R550 GNDA.n1035 GNDA.n734 585
R551 GNDA.n732 GNDA.n730 585
R552 GNDA.n1040 GNDA.n729 585
R553 GNDA.n1041 GNDA.n727 585
R554 GNDA.n726 GNDA.n722 585
R555 GNDA.n1046 GNDA.n721 585
R556 GNDA.n1046 GNDA.n1045 585
R557 GNDA.n1043 GNDA.n722 585
R558 GNDA.n1042 GNDA.n1041 585
R559 GNDA.n1040 GNDA.n1039 585
R560 GNDA.n1038 GNDA.n730 585
R561 GNDA.n1036 GNDA.n1035 585
R562 GNDA.n1034 GNDA.n731 585
R563 GNDA.n1033 GNDA.n1032 585
R564 GNDA.n1030 GNDA.n738 585
R565 GNDA.n1028 GNDA.n1027 585
R566 GNDA.n1026 GNDA.n739 585
R567 GNDA.n1025 GNDA.n1024 585
R568 GNDA.n2511 GNDA.n2510 585
R569 GNDA.n580 GNDA.n578 585
R570 GNDA.n2277 GNDA.n2276 585
R571 GNDA.n2279 GNDA.n2278 585
R572 GNDA.n2281 GNDA.n2280 585
R573 GNDA.n2283 GNDA.n2282 585
R574 GNDA.n2285 GNDA.n2284 585
R575 GNDA.n2287 GNDA.n2286 585
R576 GNDA.n2289 GNDA.n2288 585
R577 GNDA.n2291 GNDA.n2290 585
R578 GNDA.n2293 GNDA.n2292 585
R579 GNDA.n2294 GNDA.n2275 585
R580 GNDA.n720 GNDA.n719 585
R581 GNDA.n718 GNDA.n717 585
R582 GNDA.n716 GNDA.n715 585
R583 GNDA.n714 GNDA.n713 585
R584 GNDA.n712 GNDA.n711 585
R585 GNDA.n710 GNDA.n709 585
R586 GNDA.n708 GNDA.n707 585
R587 GNDA.n706 GNDA.n705 585
R588 GNDA.n704 GNDA.n703 585
R589 GNDA.n702 GNDA.n701 585
R590 GNDA.n700 GNDA.n699 585
R591 GNDA.n584 GNDA.n581 585
R592 GNDA.n782 GNDA.n781 585
R593 GNDA.n780 GNDA.n779 585
R594 GNDA.n778 GNDA.n777 585
R595 GNDA.n776 GNDA.n775 585
R596 GNDA.n774 GNDA.n773 585
R597 GNDA.n772 GNDA.n771 585
R598 GNDA.n770 GNDA.n769 585
R599 GNDA.n768 GNDA.n767 585
R600 GNDA.n766 GNDA.n765 585
R601 GNDA.n764 GNDA.n763 585
R602 GNDA.n762 GNDA.n761 585
R603 GNDA.n723 GNDA.n698 585
R604 GNDA.n696 GNDA.n582 585
R605 GNDA.n2197 GNDA.n696 585
R606 GNDA.n2268 GNDA.n2267 585
R607 GNDA.n2265 GNDA.n2264 585
R608 GNDA.n2263 GNDA.n2262 585
R609 GNDA.n673 GNDA.n635 585
R610 GNDA.n693 GNDA.n692 585
R611 GNDA.n689 GNDA.n672 585
R612 GNDA.n676 GNDA.n675 585
R613 GNDA.n684 GNDA.n683 585
R614 GNDA.n682 GNDA.n681 585
R615 GNDA.n656 GNDA.n655 585
R616 GNDA.n2202 GNDA.n2201 585
R617 GNDA.n1150 GNDA.n657 585
R618 GNDA.n1048 GNDA.n697 585
R619 GNDA.n2197 GNDA.n697 585
R620 GNDA.n695 GNDA.n582 585
R621 GNDA.n2197 GNDA.n695 585
R622 GNDA.n2157 GNDA.n2156 585
R623 GNDA.n2154 GNDA.n2153 585
R624 GNDA.n2152 GNDA.n2151 585
R625 GNDA.n2068 GNDA.n1153 585
R626 GNDA.n2070 GNDA.n2069 585
R627 GNDA.n2074 GNDA.n2073 585
R628 GNDA.n2076 GNDA.n2075 585
R629 GNDA.n2083 GNDA.n2082 585
R630 GNDA.n2081 GNDA.n2066 585
R631 GNDA.n2089 GNDA.n2088 585
R632 GNDA.n2091 GNDA.n2090 585
R633 GNDA.n2064 GNDA.n2063 585
R634 GNDA.n2196 GNDA.n1048 585
R635 GNDA.n2197 GNDA.n2196 585
R636 GNDA.n2061 GNDA.n1049 585
R637 GNDA.n2059 GNDA.n2058 585
R638 GNDA.n2057 GNDA.n2056 585
R639 GNDA.n1973 GNDA.n1174 585
R640 GNDA.n1975 GNDA.n1974 585
R641 GNDA.n1979 GNDA.n1978 585
R642 GNDA.n1981 GNDA.n1980 585
R643 GNDA.n1988 GNDA.n1987 585
R644 GNDA.n1986 GNDA.n1971 585
R645 GNDA.n1994 GNDA.n1993 585
R646 GNDA.n1996 GNDA.n1995 585
R647 GNDA.n1969 GNDA.n1968 585
R648 GNDA.n803 GNDA.n753 585
R649 GNDA.n806 GNDA.n805 585
R650 GNDA.n805 GNDA.n804 585
R651 GNDA.n752 GNDA.n751 585
R652 GNDA.n801 GNDA.n752 585
R653 GNDA.n799 GNDA.n798 585
R654 GNDA.n800 GNDA.n799 585
R655 GNDA.n797 GNDA.n755 585
R656 GNDA.n755 GNDA.n754 585
R657 GNDA.n796 GNDA.n795 585
R658 GNDA.n795 GNDA.n526 585
R659 GNDA.n794 GNDA.n756 585
R660 GNDA.n794 GNDA.n525 585
R661 GNDA.n793 GNDA.n758 585
R662 GNDA.n793 GNDA.n792 585
R663 GNDA.n787 GNDA.n757 585
R664 GNDA.n791 GNDA.n757 585
R665 GNDA.n789 GNDA.n788 585
R666 GNDA.n790 GNDA.n789 585
R667 GNDA.n786 GNDA.n760 585
R668 GNDA.n760 GNDA.n759 585
R669 GNDA.n785 GNDA.n784 585
R670 GNDA.n784 GNDA.n783 585
R671 GNDA.n802 GNDA.n749 585
R672 GNDA.n1965 GNDA.n1964 585
R673 GNDA.n1963 GNDA.n1962 585
R674 GNDA.n1963 GNDA.n1195 585
R675 GNDA.n1961 GNDA.n1196 585
R676 GNDA.n1957 GNDA.n1196 585
R677 GNDA.n1960 GNDA.n1959 585
R678 GNDA.n1959 GNDA.n1958 585
R679 GNDA.n1198 GNDA.n1197 585
R680 GNDA.n1956 GNDA.n1198 585
R681 GNDA.n1954 GNDA.n1953 585
R682 GNDA.n1955 GNDA.n1954 585
R683 GNDA.n1952 GNDA.n1199 585
R684 GNDA.n1948 GNDA.n1199 585
R685 GNDA.n1951 GNDA.n1950 585
R686 GNDA.n1950 GNDA.n1949 585
R687 GNDA.n1201 GNDA.n1200 585
R688 GNDA.n1947 GNDA.n1201 585
R689 GNDA.n1945 GNDA.n1944 585
R690 GNDA.n1946 GNDA.n1945 585
R691 GNDA.n1943 GNDA.n1203 585
R692 GNDA.n1203 GNDA.n1202 585
R693 GNDA.n1942 GNDA.n1941 585
R694 GNDA.n1941 GNDA.n1940 585
R695 GNDA.n1967 GNDA.n1966 585
R696 GNDA.n1780 GNDA.n1779 585
R697 GNDA.n1783 GNDA.n1250 585
R698 GNDA.n1250 GNDA.n1249 585
R699 GNDA.n1785 GNDA.n1784 585
R700 GNDA.n1786 GNDA.n1785 585
R701 GNDA.n1247 GNDA.n1246 585
R702 GNDA.n1787 GNDA.n1247 585
R703 GNDA.n1790 GNDA.n1789 585
R704 GNDA.n1789 GNDA.n1788 585
R705 GNDA.n1791 GNDA.n1245 585
R706 GNDA.n1248 GNDA.n1245 585
R707 GNDA.n1793 GNDA.n1792 585
R708 GNDA.n1794 GNDA.n1793 585
R709 GNDA.n1244 GNDA.n1243 585
R710 GNDA.n1795 GNDA.n1244 585
R711 GNDA.n1798 GNDA.n1797 585
R712 GNDA.n1797 GNDA.n1796 585
R713 GNDA.n1799 GNDA.n1242 585
R714 GNDA.n1242 GNDA.n1241 585
R715 GNDA.n1801 GNDA.n1800 585
R716 GNDA.n1802 GNDA.n1801 585
R717 GNDA.n1240 GNDA.n1239 585
R718 GNDA.n1803 GNDA.n1240 585
R719 GNDA.n1778 GNDA.n1777 585
R720 GNDA.n57 GNDA.n56 585
R721 GNDA.n54 GNDA.n53 585
R722 GNDA.n53 GNDA.n17 585
R723 GNDA.n62 GNDA.n61 585
R724 GNDA.n64 GNDA.n52 585
R725 GNDA.n67 GNDA.n66 585
R726 GNDA.n50 GNDA.n49 585
R727 GNDA.n72 GNDA.n71 585
R728 GNDA.n74 GNDA.n48 585
R729 GNDA.n77 GNDA.n76 585
R730 GNDA.n46 GNDA.n45 585
R731 GNDA.n82 GNDA.n81 585
R732 GNDA.n84 GNDA.n44 585
R733 GNDA.n86 GNDA.n85 585
R734 GNDA.n85 GNDA.n17 585
R735 GNDA.n134 GNDA.n130 585
R736 GNDA.n132 GNDA.n129 585
R737 GNDA.n137 GNDA.n129 585
R738 GNDA.n2592 GNDA.n5 585
R739 GNDA.n2597 GNDA.n2596 585
R740 GNDA.n2596 GNDA.n2595 585
R741 GNDA.n200 GNDA.n195 585
R742 GNDA.n198 GNDA.n194 585
R743 GNDA.n203 GNDA.n194 585
R744 GNDA.n197 GNDA.n185 585
R745 GNDA.n151 GNDA.n150 585
R746 GNDA.n156 GNDA.n149 585
R747 GNDA.n149 GNDA.n6 585
R748 GNDA.n158 GNDA.n157 585
R749 GNDA.n33 GNDA.n32 585
R750 GNDA.n116 GNDA.n31 585
R751 GNDA.n120 GNDA.n31 585
R752 GNDA.n115 GNDA.n114 585
R753 GNDA.n113 GNDA.n112 585
R754 GNDA.n111 GNDA.n110 585
R755 GNDA.n109 GNDA.n108 585
R756 GNDA.n107 GNDA.n106 585
R757 GNDA.n105 GNDA.n104 585
R758 GNDA.n103 GNDA.n102 585
R759 GNDA.n101 GNDA.n100 585
R760 GNDA.n99 GNDA.n98 585
R761 GNDA.n97 GNDA.n96 585
R762 GNDA.n94 GNDA.n30 585
R763 GNDA.n120 GNDA.n30 585
R764 GNDA.n286 GNDA.n285 585
R765 GNDA.n283 GNDA.n282 585
R766 GNDA.n282 GNDA.n235 585
R767 GNDA.n291 GNDA.n290 585
R768 GNDA.n293 GNDA.n281 585
R769 GNDA.n296 GNDA.n295 585
R770 GNDA.n279 GNDA.n278 585
R771 GNDA.n301 GNDA.n300 585
R772 GNDA.n303 GNDA.n277 585
R773 GNDA.n306 GNDA.n305 585
R774 GNDA.n275 GNDA.n274 585
R775 GNDA.n311 GNDA.n310 585
R776 GNDA.n313 GNDA.n273 585
R777 GNDA.n315 GNDA.n314 585
R778 GNDA.n314 GNDA.n235 585
R779 GNDA.n262 GNDA.n261 585
R780 GNDA.n345 GNDA.n260 585
R781 GNDA.n349 GNDA.n260 585
R782 GNDA.n344 GNDA.n343 585
R783 GNDA.n342 GNDA.n341 585
R784 GNDA.n340 GNDA.n339 585
R785 GNDA.n338 GNDA.n337 585
R786 GNDA.n336 GNDA.n335 585
R787 GNDA.n334 GNDA.n333 585
R788 GNDA.n332 GNDA.n331 585
R789 GNDA.n330 GNDA.n329 585
R790 GNDA.n328 GNDA.n327 585
R791 GNDA.n326 GNDA.n325 585
R792 GNDA.n323 GNDA.n259 585
R793 GNDA.n349 GNDA.n259 585
R794 GNDA.n20 GNDA.n19 585
R795 GNDA.n500 GNDA.n18 585
R796 GNDA.n504 GNDA.n18 585
R797 GNDA.n499 GNDA.n498 585
R798 GNDA.n497 GNDA.n496 585
R799 GNDA.n494 GNDA.n16 585
R800 GNDA.n504 GNDA.n16 585
R801 GNDA.n211 GNDA.n210 585
R802 GNDA.n215 GNDA.n122 585
R803 GNDA.n476 GNDA.n122 585
R804 GNDA.n225 GNDA.n220 585
R805 GNDA.n227 GNDA.n226 585
R806 GNDA.n226 GNDA.n127 585
R807 GNDA.n145 GNDA.n143 585
R808 GNDA.n399 GNDA.n142 585
R809 GNDA.n404 GNDA.n142 585
R810 GNDA.n380 GNDA.n232 585
R811 GNDA.n395 GNDA.n394 585
R812 GNDA.n394 GNDA.n393 585
R813 GNDA.n479 GNDA.n478 585
R814 GNDA.n484 GNDA.n477 585
R815 GNDA.n488 GNDA.n477 585
R816 GNDA.n483 GNDA.n482 585
R817 GNDA.n481 GNDA.n24 585
R818 GNDA.n490 GNDA.n489 585
R819 GNDA.n489 GNDA.n488 585
R820 GNDA.n238 GNDA.n237 585
R821 GNDA.n374 GNDA.n236 585
R822 GNDA.n378 GNDA.n236 585
R823 GNDA.n373 GNDA.n372 585
R824 GNDA.n371 GNDA.n370 585
R825 GNDA.n368 GNDA.n234 585
R826 GNDA.n378 GNDA.n234 585
R827 GNDA.n353 GNDA.n352 585
R828 GNDA.n358 GNDA.n351 585
R829 GNDA.n362 GNDA.n351 585
R830 GNDA.n357 GNDA.n356 585
R831 GNDA.n355 GNDA.n253 585
R832 GNDA.n364 GNDA.n363 585
R833 GNDA.n363 GNDA.n362 585
R834 GNDA.n474 GNDA.n473 585
R835 GNDA.n461 GNDA.n460 585
R836 GNDA.n408 GNDA.n139 585
R837 GNDA.n391 GNDA.n390 585
R838 GNDA.n470 GNDA.n469 585
R839 GNDA.n469 GNDA.n14 585
R840 GNDA.n459 GNDA.n457 585
R841 GNDA.n457 GNDA.n456 585
R842 GNDA.n410 GNDA.n409 585
R843 GNDA.n411 GNDA.n410 585
R844 GNDA.n387 GNDA.n386 585
R845 GNDA.n386 GNDA.n385 585
R846 GNDA.n430 GNDA.n429 585
R847 GNDA.n435 GNDA.n428 585
R848 GNDA.n428 GNDA.n128 585
R849 GNDA.n437 GNDA.n436 585
R850 GNDA.n451 GNDA.n413 585
R851 GNDA.n449 GNDA.n412 585
R852 GNDA.n454 GNDA.n412 585
R853 GNDA.n448 GNDA.n447 585
R854 GNDA.n2560 GNDA.n522 585
R855 GNDA.n2563 GNDA.n2562 585
R856 GNDA.n2564 GNDA.n2563 585
R857 GNDA.n2555 GNDA.n2554 585
R858 GNDA.n2485 GNDA.n610 585
R859 GNDA.n2485 GNDA.n2484 585
R860 GNDA.n2460 GNDA.n2459 585
R861 GNDA.n2461 GNDA.n2460 585
R862 GNDA.n2457 GNDA.n612 585
R863 GNDA.n2326 GNDA.n612 585
R864 GNDA.n2324 GNDA.n2320 585
R865 GNDA.n2327 GNDA.n2324 585
R866 GNDA.n2452 GNDA.n2451 585
R867 GNDA.n2451 GNDA.n2450 585
R868 GNDA.n2329 GNDA.n2325 585
R869 GNDA.n2449 GNDA.n2325 585
R870 GNDA.n2447 GNDA.n2446 585
R871 GNDA.n2448 GNDA.n2447 585
R872 GNDA.n2372 GNDA.n2328 585
R873 GNDA.n2369 GNDA.n2328 585
R874 GNDA.n2374 GNDA.n2371 585
R875 GNDA.n2371 GNDA.n2370 585
R876 GNDA.n2380 GNDA.n2379 585
R877 GNDA.n2381 GNDA.n2380 585
R878 GNDA.n2351 GNDA.n2350 585
R879 GNDA.n2382 GNDA.n2351 585
R880 GNDA.n2386 GNDA.n2385 585
R881 GNDA.n2385 GNDA.n2384 585
R882 GNDA.n2348 GNDA.n609 585
R883 GNDA.n2383 GNDA.n609 585
R884 GNDA.n1021 GNDA.n1020 585
R885 GNDA.n1020 GNDA.n556 585
R886 GNDA.n882 GNDA.n610 585
R887 GNDA.n883 GNDA.n882 585
R888 GNDA.n887 GNDA.n885 585
R889 GNDA.n885 GNDA.n884 585
R890 GNDA.n1013 GNDA.n1012 585
R891 GNDA.n1014 GNDA.n1013 585
R892 GNDA.n889 GNDA.n886 585
R893 GNDA.n894 GNDA.n886 585
R894 GNDA.n1007 GNDA.n1006 585
R895 GNDA.n1006 GNDA.n1005 585
R896 GNDA.n896 GNDA.n893 585
R897 GNDA.n1004 GNDA.n893 585
R898 GNDA.n1002 GNDA.n1001 585
R899 GNDA.n1003 GNDA.n1002 585
R900 GNDA.n927 GNDA.n895 585
R901 GNDA.n926 GNDA.n895 585
R902 GNDA.n934 GNDA.n933 585
R903 GNDA.n935 GNDA.n934 585
R904 GNDA.n929 GNDA.n917 585
R905 GNDA.n936 GNDA.n917 585
R906 GNDA.n939 GNDA.n938 585
R907 GNDA.n938 GNDA.n937 585
R908 GNDA.n940 GNDA.n879 585
R909 GNDA.n881 GNDA.n879 585
R910 GNDA.n1019 GNDA.n880 585
R911 GNDA.n1019 GNDA.n1018 585
R912 GNDA.n1022 GNDA.n1021 585
R913 GNDA.n1022 GNDA.n553 585
R914 GNDA.n877 GNDA.n552 585
R915 GNDA.n2526 GNDA.n552 585
R916 GNDA.n2528 GNDA.n550 585
R917 GNDA.n2528 GNDA.n2527 585
R918 GNDA.n2544 GNDA.n2543 585
R919 GNDA.n2543 GNDA.n2542 585
R920 GNDA.n2531 GNDA.n2529 585
R921 GNDA.n2541 GNDA.n2529 585
R922 GNDA.n2539 GNDA.n2538 585
R923 GNDA.n2540 GNDA.n2539 585
R924 GNDA.n2534 GNDA.n527 585
R925 GNDA.n2530 GNDA.n527 585
R926 GNDA.n2552 GNDA.n2551 585
R927 GNDA.n2553 GNDA.n2552 585
R928 GNDA.n529 GNDA.n528 585
R929 GNDA.n810 GNDA.n528 585
R930 GNDA.n815 GNDA.n814 585
R931 GNDA.n816 GNDA.n815 585
R932 GNDA.n748 GNDA.n747 585
R933 GNDA.n817 GNDA.n748 585
R934 GNDA.n820 GNDA.n819 585
R935 GNDA.n819 GNDA.n818 585
R936 GNDA.n809 GNDA.n808 585
R937 GNDA.n809 GNDA.n513 585
R938 GNDA.n2367 GNDA.n2366 585
R939 GNDA.n2368 GNDA.n2367 585
R940 GNDA.n2356 GNDA.n2354 585
R941 GNDA.n2360 GNDA.n2359 585
R942 GNDA.n2362 GNDA.n2361 585
R943 GNDA.n507 GNDA.n506 519.423
R944 GNDA.n1857 GNDA.t211 512.884
R945 GNDA.n87 GNDA.t270 505.467
R946 GNDA.n322 GNDA.t233 505.467
R947 GNDA.n316 GNDA.t248 505.467
R948 GNDA.n93 GNDA.t254 505.467
R949 GNDA.n216 GNDA.t204 499.442
R950 GNDA.n396 GNDA.t212 499.442
R951 GNDA.n1 GNDA.t268 499.442
R952 GNDA.n2598 GNDA.t273 499.442
R953 GNDA.n467 GNDA.t289 489.401
R954 GNDA.n464 GNDA.t207 489.401
R955 GNDA.n141 GNDA.t284 489.401
R956 GNDA.n383 GNDA.t201 489.401
R957 GNDA.n228 GNDA.t237 475.976
R958 GNDA.n228 GNDA.t217 475.976
R959 GNDA.n147 GNDA.t195 475.976
R960 GNDA.n147 GNDA.t279 475.976
R961 GNDA.n488 GNDA.n476 445.375
R962 GNDA.n393 GNDA.n378 445.375
R963 GNDA.t151 GNDA.n511 433.382
R964 GNDA.n2464 GNDA.t257 409.067
R965 GNDA.n2481 GNDA.t265 409.067
R966 GNDA.n2478 GNDA.t286 409.067
R967 GNDA.n2516 GNDA.t242 409.067
R968 GNDA.n2523 GNDA.t262 409.067
R969 GNDA.n2574 GNDA.t251 409.067
R970 GNDA.n1844 GNDA.t211 391.411
R971 GNDA.t205 GNDA.n14 364.418
R972 GNDA.t228 GNDA.n454 364.418
R973 GNDA.n411 GNDA.t196 364.418
R974 GNDA.n385 GNDA.t202 364.418
R975 GNDA.n1060 GNDA.t211 172.876
R976 GNDA.n2188 GNDA.t211 172.876
R977 GNDA.t211 GNDA.n557 172.876
R978 GNDA.t211 GNDA.n560 172.876
R979 GNDA.n1061 GNDA.t211 172.615
R980 GNDA.n1051 GNDA.t211 172.615
R981 GNDA.t211 GNDA.n559 172.615
R982 GNDA.t211 GNDA.n524 172.615
R983 GNDA.t59 GNDA.t294 296.933
R984 GNDA.t277 GNDA.t52 296.933
R985 GNDA.t117 GNDA.t228 296.933
R986 GNDA.t196 GNDA.t79 296.933
R987 GNDA.t79 GNDA.t49 296.933
R988 GNDA.t128 GNDA.t49 296.933
R989 GNDA.t18 GNDA.t211 294.625
R990 GNDA.n59 GNDA.n58 267.125
R991 GNDA.n80 GNDA.n43 267.125
R992 GNDA.n486 GNDA.n485 267.125
R993 GNDA.n480 GNDA.n23 267.125
R994 GNDA.n502 GNDA.n501 267.125
R995 GNDA.n495 GNDA.n21 267.125
R996 GNDA.n376 GNDA.n375 267.125
R997 GNDA.n369 GNDA.n239 267.125
R998 GNDA.n360 GNDA.n359 267.125
R999 GNDA.n354 GNDA.n252 267.125
R1000 GNDA.n347 GNDA.n346 267.125
R1001 GNDA.n324 GNDA.n271 267.125
R1002 GNDA.n288 GNDA.n287 267.125
R1003 GNDA.n309 GNDA.n272 267.125
R1004 GNDA.n118 GNDA.n117 267.125
R1005 GNDA.n95 GNDA.n42 267.125
R1006 GNDA.n2316 GNDA.n2315 264.301
R1007 GNDA.n2315 GNDA.n622 264.301
R1008 GNDA.n631 GNDA.n629 264.301
R1009 GNDA.n807 GNDA.n750 264.301
R1010 GNDA.n1194 GNDA.n1193 264.301
R1011 GNDA.n1782 GNDA.n1781 264.301
R1012 GNDA.n784 GNDA.n782 259.416
R1013 GNDA.n721 GNDA.n720 259.416
R1014 GNDA.n1530 GNDA.n1529 259.416
R1015 GNDA.n2511 GNDA.n579 259.416
R1016 GNDA.n2185 GNDA.n1080 259.416
R1017 GNDA.n1941 GNDA.n1939 259.416
R1018 GNDA.n1885 GNDA.n1884 259.416
R1019 GNDA.n1805 GNDA.n1240 259.416
R1020 GNDA.n1449 GNDA.n1224 259.416
R1021 GNDA.n1622 GNDA.n1291 258.334
R1022 GNDA.n2423 GNDA.n2346 258.334
R1023 GNDA.n2241 GNDA.n2240 258.334
R1024 GNDA.n2130 GNDA.n2129 258.334
R1025 GNDA.n2035 GNDA.n2034 258.334
R1026 GNDA.n1384 GNDA.n1383 258.334
R1027 GNDA.n1718 GNDA.n1676 258.334
R1028 GNDA.n977 GNDA.n913 258.334
R1029 GNDA.n859 GNDA.n858 258.334
R1030 GNDA.t208 GNDA.n128 256.442
R1031 GNDA.n456 GNDA.t277 256.442
R1032 GNDA.t52 GNDA.n455 256.442
R1033 GNDA.n2315 GNDA.n2314 254.34
R1034 GNDA.n2315 GNDA.n2273 254.34
R1035 GNDA.n2315 GNDA.n2272 254.34
R1036 GNDA.n2315 GNDA.n2271 254.34
R1037 GNDA.n2315 GNDA.n2270 254.34
R1038 GNDA.n2315 GNDA.n616 254.34
R1039 GNDA.n2315 GNDA.n617 254.34
R1040 GNDA.n2315 GNDA.n618 254.34
R1041 GNDA.n2315 GNDA.n619 254.34
R1042 GNDA.n2315 GNDA.n620 254.34
R1043 GNDA.n2315 GNDA.n623 254.34
R1044 GNDA.n2315 GNDA.n624 254.34
R1045 GNDA.n2315 GNDA.n625 254.34
R1046 GNDA.n2315 GNDA.n626 254.34
R1047 GNDA.n2315 GNDA.n627 254.34
R1048 GNDA.n2315 GNDA.n628 254.34
R1049 GNDA.n2190 GNDA.n2188 254.34
R1050 GNDA.n2188 GNDA.n1059 254.34
R1051 GNDA.n2188 GNDA.n1058 254.34
R1052 GNDA.n2188 GNDA.n1057 254.34
R1053 GNDA.n2188 GNDA.n1056 254.34
R1054 GNDA.n2188 GNDA.n1055 254.34
R1055 GNDA.n1862 GNDA.n1051 254.34
R1056 GNDA.n1910 GNDA.n1051 254.34
R1057 GNDA.n1904 GNDA.n1051 254.34
R1058 GNDA.n1902 GNDA.n1051 254.34
R1059 GNDA.n1895 GNDA.n1051 254.34
R1060 GNDA.n2194 GNDA.n1051 254.34
R1061 GNDA.n2187 GNDA.n2186 254.34
R1062 GNDA.n2187 GNDA.n1078 254.34
R1063 GNDA.n2187 GNDA.n1077 254.34
R1064 GNDA.n2187 GNDA.n1076 254.34
R1065 GNDA.n2187 GNDA.n1075 254.34
R1066 GNDA.n2187 GNDA.n1074 254.34
R1067 GNDA.n2187 GNDA.n1073 254.34
R1068 GNDA.n2187 GNDA.n1072 254.34
R1069 GNDA.n2187 GNDA.n1071 254.34
R1070 GNDA.n2187 GNDA.n1070 254.34
R1071 GNDA.n2187 GNDA.n1069 254.34
R1072 GNDA.n2187 GNDA.n1068 254.34
R1073 GNDA.n2187 GNDA.n1067 254.34
R1074 GNDA.n2187 GNDA.n1066 254.34
R1075 GNDA.n2187 GNDA.n1065 254.34
R1076 GNDA.n2187 GNDA.n1064 254.34
R1077 GNDA.n2187 GNDA.n1063 254.34
R1078 GNDA.n2187 GNDA.n1062 254.34
R1079 GNDA.n1656 GNDA.n1655 254.34
R1080 GNDA.n1656 GNDA.n1263 254.34
R1081 GNDA.n1656 GNDA.n1262 254.34
R1082 GNDA.n1656 GNDA.n1261 254.34
R1083 GNDA.n1656 GNDA.n1260 254.34
R1084 GNDA.n1656 GNDA.n1259 254.34
R1085 GNDA.n1656 GNDA.n1258 254.34
R1086 GNDA.n1656 GNDA.n1257 254.34
R1087 GNDA.n1656 GNDA.n1256 254.34
R1088 GNDA.n1656 GNDA.n1255 254.34
R1089 GNDA.n1656 GNDA.n1254 254.34
R1090 GNDA.n1656 GNDA.n1253 254.34
R1091 GNDA.n1669 GNDA.n1656 254.34
R1092 GNDA.n1745 GNDA.n1656 254.34
R1093 GNDA.n1747 GNDA.n1656 254.34
R1094 GNDA.n1760 GNDA.n1656 254.34
R1095 GNDA.n1762 GNDA.n1656 254.34
R1096 GNDA.n1775 GNDA.n1656 254.34
R1097 GNDA.n1550 GNDA.n1294 254.34
R1098 GNDA.n1553 GNDA.n1550 254.34
R1099 GNDA.n1550 GNDA.n1549 254.34
R1100 GNDA.n1550 GNDA.n1420 254.34
R1101 GNDA.n1550 GNDA.n1419 254.34
R1102 GNDA.n1550 GNDA.n1418 254.34
R1103 GNDA.n1533 GNDA.n1413 254.34
R1104 GNDA.n1535 GNDA.n1413 254.34
R1105 GNDA.n1543 GNDA.n1413 254.34
R1106 GNDA.n1545 GNDA.n1413 254.34
R1107 GNDA.n1557 GNDA.n1413 254.34
R1108 GNDA.n1560 GNDA.n1413 254.34
R1109 GNDA.n1148 GNDA.n1060 254.34
R1110 GNDA.n1145 GNDA.n1060 254.34
R1111 GNDA.n1140 GNDA.n1060 254.34
R1112 GNDA.n1137 GNDA.n1060 254.34
R1113 GNDA.n1132 GNDA.n1060 254.34
R1114 GNDA.n1129 GNDA.n1060 254.34
R1115 GNDA.n2180 GNDA.n1061 254.34
R1116 GNDA.n1128 GNDA.n1061 254.34
R1117 GNDA.n2173 GNDA.n1061 254.34
R1118 GNDA.n2167 GNDA.n1061 254.34
R1119 GNDA.n2165 GNDA.n1061 254.34
R1120 GNDA.n2159 GNDA.n1061 254.34
R1121 GNDA.n608 GNDA.n557 254.34
R1122 GNDA.n602 GNDA.n557 254.34
R1123 GNDA.n597 GNDA.n557 254.34
R1124 GNDA.n594 GNDA.n557 254.34
R1125 GNDA.n589 GNDA.n557 254.34
R1126 GNDA.n586 GNDA.n557 254.34
R1127 GNDA.n2506 GNDA.n559 254.34
R1128 GNDA.n585 GNDA.n559 254.34
R1129 GNDA.n2499 GNDA.n559 254.34
R1130 GNDA.n2493 GNDA.n559 254.34
R1131 GNDA.n2491 GNDA.n559 254.34
R1132 GNDA.n605 GNDA.n559 254.34
R1133 GNDA.n744 GNDA.n560 254.34
R1134 GNDA.n741 GNDA.n560 254.34
R1135 GNDA.n736 GNDA.n560 254.34
R1136 GNDA.n733 GNDA.n560 254.34
R1137 GNDA.n728 GNDA.n560 254.34
R1138 GNDA.n725 GNDA.n560 254.34
R1139 GNDA.n1044 GNDA.n524 254.34
R1140 GNDA.n724 GNDA.n524 254.34
R1141 GNDA.n1037 GNDA.n524 254.34
R1142 GNDA.n1031 GNDA.n524 254.34
R1143 GNDA.n1029 GNDA.n524 254.34
R1144 GNDA.n1023 GNDA.n524 254.34
R1145 GNDA.n2513 GNDA.n2512 254.34
R1146 GNDA.n2513 GNDA.n577 254.34
R1147 GNDA.n2513 GNDA.n576 254.34
R1148 GNDA.n2513 GNDA.n575 254.34
R1149 GNDA.n2513 GNDA.n574 254.34
R1150 GNDA.n2513 GNDA.n573 254.34
R1151 GNDA.n2513 GNDA.n572 254.34
R1152 GNDA.n2513 GNDA.n571 254.34
R1153 GNDA.n2513 GNDA.n570 254.34
R1154 GNDA.n2513 GNDA.n569 254.34
R1155 GNDA.n2513 GNDA.n568 254.34
R1156 GNDA.n2513 GNDA.n567 254.34
R1157 GNDA.n2513 GNDA.n566 254.34
R1158 GNDA.n2513 GNDA.n565 254.34
R1159 GNDA.n2513 GNDA.n564 254.34
R1160 GNDA.n2513 GNDA.n563 254.34
R1161 GNDA.n2513 GNDA.n562 254.34
R1162 GNDA.n2513 GNDA.n561 254.34
R1163 GNDA.n2199 GNDA.n630 254.34
R1164 GNDA.n2199 GNDA.n634 254.34
R1165 GNDA.n2199 GNDA.n694 254.34
R1166 GNDA.n2199 GNDA.n671 254.34
R1167 GNDA.n2199 GNDA.n670 254.34
R1168 GNDA.n2200 GNDA.n2199 254.34
R1169 GNDA.n2199 GNDA.n669 254.34
R1170 GNDA.n2199 GNDA.n668 254.34
R1171 GNDA.n2199 GNDA.n667 254.34
R1172 GNDA.n2199 GNDA.n666 254.34
R1173 GNDA.n2199 GNDA.n665 254.34
R1174 GNDA.n2199 GNDA.n664 254.34
R1175 GNDA.n2199 GNDA.n663 254.34
R1176 GNDA.n2199 GNDA.n662 254.34
R1177 GNDA.n2199 GNDA.n661 254.34
R1178 GNDA.n2199 GNDA.n660 254.34
R1179 GNDA.n2199 GNDA.n659 254.34
R1180 GNDA.n2199 GNDA.n658 254.34
R1181 GNDA.t211 GNDA.n1435 250.349
R1182 GNDA.n1045 GNDA.n723 249.663
R1183 GNDA.n2507 GNDA.n584 249.663
R1184 GNDA.n1504 GNDA.n1484 249.663
R1185 GNDA.n2313 GNDA.n2275 249.663
R1186 GNDA.n1103 GNDA.n1102 249.663
R1187 GNDA.n1916 GNDA.n1915 249.663
R1188 GNDA.n2181 GNDA.n1127 249.663
R1189 GNDA.n1830 GNDA.n1226 249.663
R1190 GNDA.n1532 GNDA.n1427 249.663
R1191 GNDA.n2563 GNDA.n522 246.25
R1192 GNDA.n2563 GNDA.n2554 246.25
R1193 GNDA.n413 GNDA.n412 246.25
R1194 GNDA.n447 GNDA.n412 246.25
R1195 GNDA.n430 GNDA.n428 246.25
R1196 GNDA.n437 GNDA.n428 246.25
R1197 GNDA.n391 GNDA.n386 246.25
R1198 GNDA.n410 GNDA.n139 246.25
R1199 GNDA.n461 GNDA.n457 246.25
R1200 GNDA.n474 GNDA.n469 246.25
R1201 GNDA.n352 GNDA.n351 246.25
R1202 GNDA.n356 GNDA.n351 246.25
R1203 GNDA.n363 GNDA.n253 246.25
R1204 GNDA.n237 GNDA.n236 246.25
R1205 GNDA.n372 GNDA.n236 246.25
R1206 GNDA.n370 GNDA.n234 246.25
R1207 GNDA.n478 GNDA.n477 246.25
R1208 GNDA.n482 GNDA.n477 246.25
R1209 GNDA.n489 GNDA.n24 246.25
R1210 GNDA.n394 GNDA.n232 246.25
R1211 GNDA.n143 GNDA.n142 246.25
R1212 GNDA.n226 GNDA.n225 246.25
R1213 GNDA.n210 GNDA.n122 246.25
R1214 GNDA.n19 GNDA.n18 246.25
R1215 GNDA.n498 GNDA.n18 246.25
R1216 GNDA.n496 GNDA.n16 246.25
R1217 GNDA.n261 GNDA.n260 246.25
R1218 GNDA.n343 GNDA.n260 246.25
R1219 GNDA.n341 GNDA.n340 246.25
R1220 GNDA.n337 GNDA.n336 246.25
R1221 GNDA.n333 GNDA.n332 246.25
R1222 GNDA.n329 GNDA.n328 246.25
R1223 GNDA.n325 GNDA.n259 246.25
R1224 GNDA.n285 GNDA.n282 246.25
R1225 GNDA.n291 GNDA.n282 246.25
R1226 GNDA.n295 GNDA.n293 246.25
R1227 GNDA.n301 GNDA.n278 246.25
R1228 GNDA.n305 GNDA.n303 246.25
R1229 GNDA.n311 GNDA.n274 246.25
R1230 GNDA.n314 GNDA.n313 246.25
R1231 GNDA.n32 GNDA.n31 246.25
R1232 GNDA.n114 GNDA.n31 246.25
R1233 GNDA.n112 GNDA.n111 246.25
R1234 GNDA.n108 GNDA.n107 246.25
R1235 GNDA.n104 GNDA.n103 246.25
R1236 GNDA.n100 GNDA.n99 246.25
R1237 GNDA.n96 GNDA.n30 246.25
R1238 GNDA.n151 GNDA.n149 246.25
R1239 GNDA.n158 GNDA.n149 246.25
R1240 GNDA.n195 GNDA.n194 246.25
R1241 GNDA.n194 GNDA.n185 246.25
R1242 GNDA.n2596 GNDA.n5 246.25
R1243 GNDA.n130 GNDA.n129 246.25
R1244 GNDA.n56 GNDA.n53 246.25
R1245 GNDA.n62 GNDA.n53 246.25
R1246 GNDA.n66 GNDA.n64 246.25
R1247 GNDA.n72 GNDA.n49 246.25
R1248 GNDA.n76 GNDA.n74 246.25
R1249 GNDA.n82 GNDA.n45 246.25
R1250 GNDA.n85 GNDA.n84 246.25
R1251 GNDA.n2367 GNDA.n2354 246.25
R1252 GNDA.n2361 GNDA.n2360 246.25
R1253 GNDA.n2570 GNDA.n2569 241.643
R1254 GNDA.n55 GNDA.n17 241.643
R1255 GNDA.n63 GNDA.n17 241.643
R1256 GNDA.n65 GNDA.n17 241.643
R1257 GNDA.n73 GNDA.n17 241.643
R1258 GNDA.n75 GNDA.n17 241.643
R1259 GNDA.n83 GNDA.n17 241.643
R1260 GNDA.n137 GNDA.n136 241.643
R1261 GNDA.n2595 GNDA.n2594 241.643
R1262 GNDA.n203 GNDA.n202 241.643
R1263 GNDA.n204 GNDA.n203 241.643
R1264 GNDA.n152 GNDA.n6 241.643
R1265 GNDA.n159 GNDA.n6 241.643
R1266 GNDA.n120 GNDA.n119 241.643
R1267 GNDA.n120 GNDA.n25 241.643
R1268 GNDA.n120 GNDA.n26 241.643
R1269 GNDA.n120 GNDA.n27 241.643
R1270 GNDA.n120 GNDA.n28 241.643
R1271 GNDA.n120 GNDA.n29 241.643
R1272 GNDA.n284 GNDA.n235 241.643
R1273 GNDA.n292 GNDA.n235 241.643
R1274 GNDA.n294 GNDA.n235 241.643
R1275 GNDA.n302 GNDA.n235 241.643
R1276 GNDA.n304 GNDA.n235 241.643
R1277 GNDA.n312 GNDA.n235 241.643
R1278 GNDA.n349 GNDA.n348 241.643
R1279 GNDA.n349 GNDA.n254 241.643
R1280 GNDA.n349 GNDA.n255 241.643
R1281 GNDA.n349 GNDA.n256 241.643
R1282 GNDA.n349 GNDA.n257 241.643
R1283 GNDA.n349 GNDA.n258 241.643
R1284 GNDA.n504 GNDA.n503 241.643
R1285 GNDA.n504 GNDA.n15 241.643
R1286 GNDA.n476 GNDA.n123 241.643
R1287 GNDA.n224 GNDA.n127 241.643
R1288 GNDA.n404 GNDA.n403 241.643
R1289 GNDA.n393 GNDA.n382 241.643
R1290 GNDA.n488 GNDA.n487 241.643
R1291 GNDA.n488 GNDA.n121 241.643
R1292 GNDA.n378 GNDA.n377 241.643
R1293 GNDA.n378 GNDA.n233 241.643
R1294 GNDA.n362 GNDA.n361 241.643
R1295 GNDA.n362 GNDA.n350 241.643
R1296 GNDA.n476 GNDA.n475 241.643
R1297 GNDA.n462 GNDA.n127 241.643
R1298 GNDA.n405 GNDA.n404 241.643
R1299 GNDA.n393 GNDA.n392 241.643
R1300 GNDA.n431 GNDA.n128 241.643
R1301 GNDA.n438 GNDA.n128 241.643
R1302 GNDA.n454 GNDA.n453 241.643
R1303 GNDA.n454 GNDA.n138 241.643
R1304 GNDA.n2565 GNDA.n2564 241.643
R1305 GNDA.n2564 GNDA.n523 241.643
R1306 GNDA.n2368 GNDA.n2352 241.643
R1307 GNDA.n2368 GNDA.n2353 241.643
R1308 GNDA.n417 GNDA.n415 206.052
R1309 GNDA.n242 GNDA.n240 206.052
R1310 GNDA.n423 GNDA.n422 205.488
R1311 GNDA.n421 GNDA.n420 205.488
R1312 GNDA.n419 GNDA.n418 205.488
R1313 GNDA.n417 GNDA.n416 205.488
R1314 GNDA.n248 GNDA.n247 205.488
R1315 GNDA.n246 GNDA.n245 205.488
R1316 GNDA.n244 GNDA.n243 205.488
R1317 GNDA.n242 GNDA.n241 205.488
R1318 GNDA.n425 GNDA.n424 200.988
R1319 GNDA.n250 GNDA.n249 200.988
R1320 GNDA.n809 GNDA.n749 197
R1321 GNDA.n1020 GNDA.n1019 197
R1322 GNDA.n1565 GNDA.n1564 197
R1323 GNDA.n2485 GNDA.n609 197
R1324 GNDA.n696 GNDA.n657 197
R1325 GNDA.n1968 GNDA.n1967 197
R1326 GNDA.n2063 GNDA.n697 197
R1327 GNDA.n1777 GNDA.n1776 197
R1328 GNDA.n1317 GNDA.n1205 197
R1329 GNDA.n1442 GNDA.n1436 197
R1330 GNDA.n1022 GNDA.n552 187.249
R1331 GNDA.n885 GNDA.n882 187.249
R1332 GNDA.n1654 GNDA.n1265 187.249
R1333 GNDA.n2460 GNDA.n611 187.249
R1334 GNDA.n2269 GNDA.n2268 187.249
R1335 GNDA.n2196 GNDA.n1049 187.249
R1336 GNDA.n2156 GNDA.n695 187.249
R1337 GNDA.n1859 GNDA.n1207 187.249
R1338 GNDA.n1412 GNDA.n1411 187.249
R1339 GNDA.n2566 GNDA.n521 185
R1340 GNDA.n2558 GNDA.n2557 185
R1341 GNDA.n201 GNDA.n196 185
R1342 GNDA.n154 GNDA.n153 185
R1343 GNDA.n213 GNDA.n212 185
R1344 GNDA.n223 GNDA.n222 185
R1345 GNDA.n227 GNDA.n218 185
R1346 GNDA.n402 GNDA.n401 185
R1347 GNDA.n399 GNDA.n146 185
R1348 GNDA.n381 GNDA.n379 185
R1349 GNDA.n485 GNDA.n484 185
R1350 GNDA.n483 GNDA.n480 185
R1351 GNDA.n501 GNDA.n500 185
R1352 GNDA.n499 GNDA.n21 185
R1353 GNDA.n471 GNDA.n470 185
R1354 GNDA.n459 GNDA.n458 185
R1355 GNDA.n409 GNDA.n140 185
R1356 GNDA.n388 GNDA.n387 185
R1357 GNDA.n433 GNDA.n432 185
R1358 GNDA.n452 GNDA.n414 185
R1359 GNDA.n135 GNDA.n131 185
R1360 GNDA.n2593 GNDA.n2591 185
R1361 GNDA.n375 GNDA.n374 185
R1362 GNDA.n373 GNDA.n239 185
R1363 GNDA.n359 GNDA.n358 185
R1364 GNDA.n357 GNDA.n354 185
R1365 GNDA.n346 GNDA.n345 185
R1366 GNDA.n344 GNDA.n263 185
R1367 GNDA.n342 GNDA.n264 185
R1368 GNDA.n339 GNDA.n265 185
R1369 GNDA.n338 GNDA.n266 185
R1370 GNDA.n335 GNDA.n267 185
R1371 GNDA.n334 GNDA.n268 185
R1372 GNDA.n331 GNDA.n269 185
R1373 GNDA.n330 GNDA.n270 185
R1374 GNDA.n327 GNDA.n271 185
R1375 GNDA.n288 GNDA.n283 185
R1376 GNDA.n290 GNDA.n289 185
R1377 GNDA.n281 GNDA.n280 185
R1378 GNDA.n297 GNDA.n296 185
R1379 GNDA.n298 GNDA.n279 185
R1380 GNDA.n300 GNDA.n299 185
R1381 GNDA.n277 GNDA.n276 185
R1382 GNDA.n307 GNDA.n306 185
R1383 GNDA.n308 GNDA.n275 185
R1384 GNDA.n310 GNDA.n309 185
R1385 GNDA.n117 GNDA.n116 185
R1386 GNDA.n115 GNDA.n34 185
R1387 GNDA.n113 GNDA.n35 185
R1388 GNDA.n110 GNDA.n36 185
R1389 GNDA.n109 GNDA.n37 185
R1390 GNDA.n106 GNDA.n38 185
R1391 GNDA.n105 GNDA.n39 185
R1392 GNDA.n102 GNDA.n40 185
R1393 GNDA.n101 GNDA.n41 185
R1394 GNDA.n98 GNDA.n42 185
R1395 GNDA.n59 GNDA.n54 185
R1396 GNDA.n61 GNDA.n60 185
R1397 GNDA.n52 GNDA.n51 185
R1398 GNDA.n68 GNDA.n67 185
R1399 GNDA.n69 GNDA.n50 185
R1400 GNDA.n71 GNDA.n70 185
R1401 GNDA.n48 GNDA.n47 185
R1402 GNDA.n78 GNDA.n77 185
R1403 GNDA.n79 GNDA.n46 185
R1404 GNDA.n81 GNDA.n80 185
R1405 GNDA.n1624 GNDA.n1291 185
R1406 GNDA.n1638 GNDA.n1637 185
R1407 GNDA.n1636 GNDA.n1292 185
R1408 GNDA.n1635 GNDA.n1634 185
R1409 GNDA.n1633 GNDA.n1632 185
R1410 GNDA.n1631 GNDA.n1630 185
R1411 GNDA.n1629 GNDA.n1628 185
R1412 GNDA.n1627 GNDA.n1626 185
R1413 GNDA.n1625 GNDA.n1268 185
R1414 GNDA.n1607 GNDA.n1606 185
R1415 GNDA.n1609 GNDA.n1608 185
R1416 GNDA.n1611 GNDA.n1610 185
R1417 GNDA.n1613 GNDA.n1612 185
R1418 GNDA.n1615 GNDA.n1614 185
R1419 GNDA.n1617 GNDA.n1616 185
R1420 GNDA.n1619 GNDA.n1618 185
R1421 GNDA.n1621 GNDA.n1620 185
R1422 GNDA.n1623 GNDA.n1622 185
R1423 GNDA.n1589 GNDA.n1588 185
R1424 GNDA.n1591 GNDA.n1590 185
R1425 GNDA.n1593 GNDA.n1592 185
R1426 GNDA.n1595 GNDA.n1594 185
R1427 GNDA.n1597 GNDA.n1596 185
R1428 GNDA.n1599 GNDA.n1598 185
R1429 GNDA.n1601 GNDA.n1600 185
R1430 GNDA.n1603 GNDA.n1602 185
R1431 GNDA.n1605 GNDA.n1604 185
R1432 GNDA.n1587 GNDA.n1586 185
R1433 GNDA.n1581 GNDA.n1580 185
R1434 GNDA.n1579 GNDA.n1578 185
R1435 GNDA.n1574 GNDA.n1573 185
R1436 GNDA.n1569 GNDA.n1276 185
R1437 GNDA.n1642 GNDA.n1641 185
R1438 GNDA.n1275 GNDA.n1273 185
R1439 GNDA.n1648 GNDA.n1647 185
R1440 GNDA.n1650 GNDA.n1649 185
R1441 GNDA.n2425 GNDA.n2346 185
R1442 GNDA.n2439 GNDA.n2438 185
R1443 GNDA.n2437 GNDA.n2347 185
R1444 GNDA.n2436 GNDA.n2435 185
R1445 GNDA.n2434 GNDA.n2433 185
R1446 GNDA.n2432 GNDA.n2431 185
R1447 GNDA.n2430 GNDA.n2429 185
R1448 GNDA.n2428 GNDA.n2427 185
R1449 GNDA.n2426 GNDA.n2319 185
R1450 GNDA.n2408 GNDA.n2407 185
R1451 GNDA.n2410 GNDA.n2409 185
R1452 GNDA.n2412 GNDA.n2411 185
R1453 GNDA.n2414 GNDA.n2413 185
R1454 GNDA.n2416 GNDA.n2415 185
R1455 GNDA.n2418 GNDA.n2417 185
R1456 GNDA.n2420 GNDA.n2419 185
R1457 GNDA.n2422 GNDA.n2421 185
R1458 GNDA.n2424 GNDA.n2423 185
R1459 GNDA.n2390 GNDA.n2389 185
R1460 GNDA.n2392 GNDA.n2391 185
R1461 GNDA.n2394 GNDA.n2393 185
R1462 GNDA.n2396 GNDA.n2395 185
R1463 GNDA.n2398 GNDA.n2397 185
R1464 GNDA.n2400 GNDA.n2399 185
R1465 GNDA.n2402 GNDA.n2401 185
R1466 GNDA.n2404 GNDA.n2403 185
R1467 GNDA.n2406 GNDA.n2405 185
R1468 GNDA.n2388 GNDA.n2387 185
R1469 GNDA.n2378 GNDA.n2377 185
R1470 GNDA.n2376 GNDA.n2375 185
R1471 GNDA.n2373 GNDA.n2331 185
R1472 GNDA.n2445 GNDA.n2444 185
R1473 GNDA.n2442 GNDA.n2330 185
R1474 GNDA.n2441 GNDA.n2323 185
R1475 GNDA.n2454 GNDA.n2453 185
R1476 GNDA.n2456 GNDA.n2455 185
R1477 GNDA.n2242 GNDA.n2241 185
R1478 GNDA.n2244 GNDA.n2243 185
R1479 GNDA.n2246 GNDA.n2245 185
R1480 GNDA.n2248 GNDA.n2247 185
R1481 GNDA.n2250 GNDA.n2249 185
R1482 GNDA.n2252 GNDA.n2251 185
R1483 GNDA.n2254 GNDA.n2253 185
R1484 GNDA.n2256 GNDA.n2255 185
R1485 GNDA.n2257 GNDA.n632 185
R1486 GNDA.n2224 GNDA.n2223 185
R1487 GNDA.n2226 GNDA.n2225 185
R1488 GNDA.n2228 GNDA.n2227 185
R1489 GNDA.n2230 GNDA.n2229 185
R1490 GNDA.n2232 GNDA.n2231 185
R1491 GNDA.n2234 GNDA.n2233 185
R1492 GNDA.n2236 GNDA.n2235 185
R1493 GNDA.n2238 GNDA.n2237 185
R1494 GNDA.n2240 GNDA.n2239 185
R1495 GNDA.n2206 GNDA.n2205 185
R1496 GNDA.n2208 GNDA.n2207 185
R1497 GNDA.n2210 GNDA.n2209 185
R1498 GNDA.n2212 GNDA.n2211 185
R1499 GNDA.n2214 GNDA.n2213 185
R1500 GNDA.n2216 GNDA.n2215 185
R1501 GNDA.n2218 GNDA.n2217 185
R1502 GNDA.n2220 GNDA.n2219 185
R1503 GNDA.n2222 GNDA.n2221 185
R1504 GNDA.n2204 GNDA.n2203 185
R1505 GNDA.n680 GNDA.n679 185
R1506 GNDA.n678 GNDA.n677 185
R1507 GNDA.n686 GNDA.n685 185
R1508 GNDA.n688 GNDA.n687 185
R1509 GNDA.n691 GNDA.n690 185
R1510 GNDA.n674 GNDA.n637 185
R1511 GNDA.n2261 GNDA.n2260 185
R1512 GNDA.n636 GNDA.n633 185
R1513 GNDA.n2131 GNDA.n2130 185
R1514 GNDA.n2133 GNDA.n2132 185
R1515 GNDA.n2135 GNDA.n2134 185
R1516 GNDA.n2137 GNDA.n2136 185
R1517 GNDA.n2139 GNDA.n2138 185
R1518 GNDA.n2141 GNDA.n2140 185
R1519 GNDA.n2143 GNDA.n2142 185
R1520 GNDA.n2145 GNDA.n2144 185
R1521 GNDA.n2146 GNDA.n1151 185
R1522 GNDA.n2113 GNDA.n2112 185
R1523 GNDA.n2115 GNDA.n2114 185
R1524 GNDA.n2117 GNDA.n2116 185
R1525 GNDA.n2119 GNDA.n2118 185
R1526 GNDA.n2121 GNDA.n2120 185
R1527 GNDA.n2123 GNDA.n2122 185
R1528 GNDA.n2125 GNDA.n2124 185
R1529 GNDA.n2127 GNDA.n2126 185
R1530 GNDA.n2129 GNDA.n2128 185
R1531 GNDA.n2095 GNDA.n2094 185
R1532 GNDA.n2097 GNDA.n2096 185
R1533 GNDA.n2099 GNDA.n2098 185
R1534 GNDA.n2101 GNDA.n2100 185
R1535 GNDA.n2103 GNDA.n2102 185
R1536 GNDA.n2105 GNDA.n2104 185
R1537 GNDA.n2107 GNDA.n2106 185
R1538 GNDA.n2109 GNDA.n2108 185
R1539 GNDA.n2111 GNDA.n2110 185
R1540 GNDA.n2093 GNDA.n2092 185
R1541 GNDA.n2087 GNDA.n2086 185
R1542 GNDA.n2085 GNDA.n2084 185
R1543 GNDA.n2080 GNDA.n2079 185
R1544 GNDA.n2078 GNDA.n2077 185
R1545 GNDA.n2072 GNDA.n2071 185
R1546 GNDA.n2067 GNDA.n1155 185
R1547 GNDA.n2150 GNDA.n2149 185
R1548 GNDA.n1154 GNDA.n1152 185
R1549 GNDA.n2036 GNDA.n2035 185
R1550 GNDA.n2038 GNDA.n2037 185
R1551 GNDA.n2040 GNDA.n2039 185
R1552 GNDA.n2042 GNDA.n2041 185
R1553 GNDA.n2044 GNDA.n2043 185
R1554 GNDA.n2046 GNDA.n2045 185
R1555 GNDA.n2048 GNDA.n2047 185
R1556 GNDA.n2050 GNDA.n2049 185
R1557 GNDA.n2051 GNDA.n1172 185
R1558 GNDA.n2018 GNDA.n2017 185
R1559 GNDA.n2020 GNDA.n2019 185
R1560 GNDA.n2022 GNDA.n2021 185
R1561 GNDA.n2024 GNDA.n2023 185
R1562 GNDA.n2026 GNDA.n2025 185
R1563 GNDA.n2028 GNDA.n2027 185
R1564 GNDA.n2030 GNDA.n2029 185
R1565 GNDA.n2032 GNDA.n2031 185
R1566 GNDA.n2034 GNDA.n2033 185
R1567 GNDA.n2000 GNDA.n1999 185
R1568 GNDA.n2002 GNDA.n2001 185
R1569 GNDA.n2004 GNDA.n2003 185
R1570 GNDA.n2006 GNDA.n2005 185
R1571 GNDA.n2008 GNDA.n2007 185
R1572 GNDA.n2010 GNDA.n2009 185
R1573 GNDA.n2012 GNDA.n2011 185
R1574 GNDA.n2014 GNDA.n2013 185
R1575 GNDA.n2016 GNDA.n2015 185
R1576 GNDA.n1998 GNDA.n1997 185
R1577 GNDA.n1992 GNDA.n1991 185
R1578 GNDA.n1990 GNDA.n1989 185
R1579 GNDA.n1985 GNDA.n1984 185
R1580 GNDA.n1983 GNDA.n1982 185
R1581 GNDA.n1977 GNDA.n1976 185
R1582 GNDA.n1972 GNDA.n1176 185
R1583 GNDA.n2055 GNDA.n2054 185
R1584 GNDA.n1175 GNDA.n1173 185
R1585 GNDA.n1385 GNDA.n1384 185
R1586 GNDA.n1387 GNDA.n1386 185
R1587 GNDA.n1389 GNDA.n1388 185
R1588 GNDA.n1391 GNDA.n1390 185
R1589 GNDA.n1393 GNDA.n1392 185
R1590 GNDA.n1395 GNDA.n1394 185
R1591 GNDA.n1397 GNDA.n1396 185
R1592 GNDA.n1399 GNDA.n1398 185
R1593 GNDA.n1400 GNDA.n1296 185
R1594 GNDA.n1367 GNDA.n1366 185
R1595 GNDA.n1369 GNDA.n1368 185
R1596 GNDA.n1371 GNDA.n1370 185
R1597 GNDA.n1373 GNDA.n1372 185
R1598 GNDA.n1375 GNDA.n1374 185
R1599 GNDA.n1377 GNDA.n1376 185
R1600 GNDA.n1379 GNDA.n1378 185
R1601 GNDA.n1381 GNDA.n1380 185
R1602 GNDA.n1383 GNDA.n1382 185
R1603 GNDA.n1349 GNDA.n1348 185
R1604 GNDA.n1351 GNDA.n1350 185
R1605 GNDA.n1353 GNDA.n1352 185
R1606 GNDA.n1355 GNDA.n1354 185
R1607 GNDA.n1357 GNDA.n1356 185
R1608 GNDA.n1359 GNDA.n1358 185
R1609 GNDA.n1361 GNDA.n1360 185
R1610 GNDA.n1363 GNDA.n1362 185
R1611 GNDA.n1365 GNDA.n1364 185
R1612 GNDA.n1718 GNDA.n1717 185
R1613 GNDA.n1720 GNDA.n1675 185
R1614 GNDA.n1723 GNDA.n1722 185
R1615 GNDA.n1724 GNDA.n1674 185
R1616 GNDA.n1726 GNDA.n1725 185
R1617 GNDA.n1728 GNDA.n1673 185
R1618 GNDA.n1731 GNDA.n1730 185
R1619 GNDA.n1732 GNDA.n1672 185
R1620 GNDA.n1737 GNDA.n1736 185
R1621 GNDA.n1700 GNDA.n1680 185
R1622 GNDA.n1702 GNDA.n1701 185
R1623 GNDA.n1704 GNDA.n1679 185
R1624 GNDA.n1707 GNDA.n1706 185
R1625 GNDA.n1708 GNDA.n1678 185
R1626 GNDA.n1710 GNDA.n1709 185
R1627 GNDA.n1712 GNDA.n1677 185
R1628 GNDA.n1715 GNDA.n1714 185
R1629 GNDA.n1716 GNDA.n1676 185
R1630 GNDA.n1771 GNDA.n1770 185
R1631 GNDA.n1685 GNDA.n1659 185
R1632 GNDA.n1687 GNDA.n1686 185
R1633 GNDA.n1689 GNDA.n1683 185
R1634 GNDA.n1691 GNDA.n1690 185
R1635 GNDA.n1692 GNDA.n1682 185
R1636 GNDA.n1694 GNDA.n1693 185
R1637 GNDA.n1696 GNDA.n1681 185
R1638 GNDA.n1699 GNDA.n1698 185
R1639 GNDA.n1769 GNDA.n1658 185
R1640 GNDA.n1767 GNDA.n1766 185
R1641 GNDA.n1662 GNDA.n1661 185
R1642 GNDA.n1757 GNDA.n1756 185
R1643 GNDA.n1754 GNDA.n1665 185
R1644 GNDA.n1752 GNDA.n1751 185
R1645 GNDA.n1667 GNDA.n1666 185
R1646 GNDA.n1742 GNDA.n1741 185
R1647 GNDA.n1739 GNDA.n1671 185
R1648 GNDA.n1347 GNDA.n1346 185
R1649 GNDA.n1341 GNDA.n1340 185
R1650 GNDA.n1339 GNDA.n1338 185
R1651 GNDA.n1334 GNDA.n1333 185
R1652 GNDA.n1332 GNDA.n1331 185
R1653 GNDA.n1326 GNDA.n1325 185
R1654 GNDA.n1321 GNDA.n1300 185
R1655 GNDA.n1404 GNDA.n1403 185
R1656 GNDA.n1299 GNDA.n1297 185
R1657 GNDA.n979 GNDA.n913 185
R1658 GNDA.n994 GNDA.n993 185
R1659 GNDA.n992 GNDA.n914 185
R1660 GNDA.n991 GNDA.n990 185
R1661 GNDA.n989 GNDA.n988 185
R1662 GNDA.n987 GNDA.n986 185
R1663 GNDA.n985 GNDA.n984 185
R1664 GNDA.n983 GNDA.n982 185
R1665 GNDA.n981 GNDA.n980 185
R1666 GNDA.n962 GNDA.n961 185
R1667 GNDA.n964 GNDA.n963 185
R1668 GNDA.n966 GNDA.n965 185
R1669 GNDA.n968 GNDA.n967 185
R1670 GNDA.n970 GNDA.n969 185
R1671 GNDA.n972 GNDA.n971 185
R1672 GNDA.n974 GNDA.n973 185
R1673 GNDA.n976 GNDA.n975 185
R1674 GNDA.n978 GNDA.n977 185
R1675 GNDA.n944 GNDA.n943 185
R1676 GNDA.n946 GNDA.n945 185
R1677 GNDA.n948 GNDA.n947 185
R1678 GNDA.n950 GNDA.n949 185
R1679 GNDA.n952 GNDA.n951 185
R1680 GNDA.n954 GNDA.n953 185
R1681 GNDA.n956 GNDA.n955 185
R1682 GNDA.n958 GNDA.n957 185
R1683 GNDA.n960 GNDA.n959 185
R1684 GNDA.n942 GNDA.n941 185
R1685 GNDA.n930 GNDA.n916 185
R1686 GNDA.n932 GNDA.n931 185
R1687 GNDA.n928 GNDA.n898 185
R1688 GNDA.n1000 GNDA.n999 185
R1689 GNDA.n997 GNDA.n897 185
R1690 GNDA.n996 GNDA.n892 185
R1691 GNDA.n1009 GNDA.n1008 185
R1692 GNDA.n1011 GNDA.n1010 185
R1693 GNDA.n860 GNDA.n859 185
R1694 GNDA.n862 GNDA.n861 185
R1695 GNDA.n864 GNDA.n863 185
R1696 GNDA.n866 GNDA.n865 185
R1697 GNDA.n868 GNDA.n867 185
R1698 GNDA.n870 GNDA.n869 185
R1699 GNDA.n872 GNDA.n871 185
R1700 GNDA.n874 GNDA.n873 185
R1701 GNDA.n875 GNDA.n548 185
R1702 GNDA.n842 GNDA.n841 185
R1703 GNDA.n844 GNDA.n843 185
R1704 GNDA.n846 GNDA.n845 185
R1705 GNDA.n848 GNDA.n847 185
R1706 GNDA.n850 GNDA.n849 185
R1707 GNDA.n852 GNDA.n851 185
R1708 GNDA.n854 GNDA.n853 185
R1709 GNDA.n856 GNDA.n855 185
R1710 GNDA.n858 GNDA.n857 185
R1711 GNDA.n824 GNDA.n823 185
R1712 GNDA.n826 GNDA.n825 185
R1713 GNDA.n828 GNDA.n827 185
R1714 GNDA.n830 GNDA.n829 185
R1715 GNDA.n832 GNDA.n831 185
R1716 GNDA.n834 GNDA.n833 185
R1717 GNDA.n836 GNDA.n835 185
R1718 GNDA.n838 GNDA.n837 185
R1719 GNDA.n840 GNDA.n839 185
R1720 GNDA.n822 GNDA.n821 185
R1721 GNDA.n813 GNDA.n812 185
R1722 GNDA.n811 GNDA.n531 185
R1723 GNDA.n2550 GNDA.n2549 185
R1724 GNDA.n2533 GNDA.n530 185
R1725 GNDA.n2537 GNDA.n2536 185
R1726 GNDA.n2535 GNDA.n2532 185
R1727 GNDA.n551 GNDA.n549 185
R1728 GNDA.n2546 GNDA.n2545 185
R1729 GNDA.n2366 GNDA.n2355 185
R1730 GNDA.n2359 GNDA.n2355 185
R1731 GNDA.n2366 GNDA.n2365 185
R1732 GNDA.n2365 GNDA.n2364 185
R1733 GNDA.n1528 GNDA.t211 183.948
R1734 GNDA.n1828 GNDA.n1227 183.948
R1735 GNDA.n1430 GNDA.t211 180.013
R1736 GNDA.n1828 GNDA.n1827 180.013
R1737 GNDA.n784 GNDA.n760 175.546
R1738 GNDA.n789 GNDA.n760 175.546
R1739 GNDA.n789 GNDA.n757 175.546
R1740 GNDA.n793 GNDA.n757 175.546
R1741 GNDA.n794 GNDA.n793 175.546
R1742 GNDA.n795 GNDA.n794 175.546
R1743 GNDA.n795 GNDA.n755 175.546
R1744 GNDA.n799 GNDA.n755 175.546
R1745 GNDA.n799 GNDA.n752 175.546
R1746 GNDA.n805 GNDA.n752 175.546
R1747 GNDA.n805 GNDA.n753 175.546
R1748 GNDA.n763 GNDA.n762 175.546
R1749 GNDA.n767 GNDA.n766 175.546
R1750 GNDA.n771 GNDA.n770 175.546
R1751 GNDA.n775 GNDA.n774 175.546
R1752 GNDA.n779 GNDA.n778 175.546
R1753 GNDA.n2528 GNDA.n552 175.546
R1754 GNDA.n2543 GNDA.n2528 175.546
R1755 GNDA.n2543 GNDA.n2529 175.546
R1756 GNDA.n2539 GNDA.n2529 175.546
R1757 GNDA.n2539 GNDA.n527 175.546
R1758 GNDA.n2552 GNDA.n527 175.546
R1759 GNDA.n2552 GNDA.n528 175.546
R1760 GNDA.n815 GNDA.n528 175.546
R1761 GNDA.n815 GNDA.n748 175.546
R1762 GNDA.n819 GNDA.n748 175.546
R1763 GNDA.n819 GNDA.n809 175.546
R1764 GNDA.n1043 GNDA.n1042 175.546
R1765 GNDA.n1039 GNDA.n1038 175.546
R1766 GNDA.n1036 GNDA.n731 175.546
R1767 GNDA.n1032 GNDA.n1030 175.546
R1768 GNDA.n1028 GNDA.n739 175.546
R1769 GNDA.n727 GNDA.n726 175.546
R1770 GNDA.n732 GNDA.n729 175.546
R1771 GNDA.n735 GNDA.n734 175.546
R1772 GNDA.n740 GNDA.n737 175.546
R1773 GNDA.n743 GNDA.n742 175.546
R1774 GNDA.n701 GNDA.n700 175.546
R1775 GNDA.n705 GNDA.n704 175.546
R1776 GNDA.n709 GNDA.n708 175.546
R1777 GNDA.n713 GNDA.n712 175.546
R1778 GNDA.n717 GNDA.n716 175.546
R1779 GNDA.n1013 GNDA.n885 175.546
R1780 GNDA.n1013 GNDA.n886 175.546
R1781 GNDA.n1006 GNDA.n886 175.546
R1782 GNDA.n1006 GNDA.n893 175.546
R1783 GNDA.n1002 GNDA.n893 175.546
R1784 GNDA.n1002 GNDA.n895 175.546
R1785 GNDA.n934 GNDA.n895 175.546
R1786 GNDA.n934 GNDA.n917 175.546
R1787 GNDA.n938 GNDA.n917 175.546
R1788 GNDA.n938 GNDA.n879 175.546
R1789 GNDA.n1019 GNDA.n879 175.546
R1790 GNDA.n2505 GNDA.n2504 175.546
R1791 GNDA.n2501 GNDA.n2500 175.546
R1792 GNDA.n2498 GNDA.n592 175.546
R1793 GNDA.n2494 GNDA.n2492 175.546
R1794 GNDA.n2490 GNDA.n600 175.546
R1795 GNDA.n1426 GNDA.n1425 175.546
R1796 GNDA.n1540 GNDA.n1539 175.546
R1797 GNDA.n1548 GNDA.n1421 175.546
R1798 GNDA.n1554 GNDA.n1417 175.546
R1799 GNDA.n1552 GNDA.n1551 175.546
R1800 GNDA.n1508 GNDA.n1484 175.546
R1801 GNDA.n1508 GNDA.n1482 175.546
R1802 GNDA.n1512 GNDA.n1482 175.546
R1803 GNDA.n1512 GNDA.n1480 175.546
R1804 GNDA.n1516 GNDA.n1480 175.546
R1805 GNDA.n1516 GNDA.n1478 175.546
R1806 GNDA.n1520 GNDA.n1478 175.546
R1807 GNDA.n1520 GNDA.n1476 175.546
R1808 GNDA.n1525 GNDA.n1476 175.546
R1809 GNDA.n1525 GNDA.n1473 175.546
R1810 GNDA.n1529 GNDA.n1473 175.546
R1811 GNDA.n1269 GNDA.n1264 175.546
R1812 GNDA.n1645 GNDA.n1644 175.546
R1813 GNDA.n1571 GNDA.n1570 175.546
R1814 GNDA.n1576 GNDA.n1575 175.546
R1815 GNDA.n1584 GNDA.n1583 175.546
R1816 GNDA.n1502 GNDA.n1501 175.546
R1817 GNDA.n1498 GNDA.n1497 175.546
R1818 GNDA.n1494 GNDA.n1493 175.546
R1819 GNDA.n1490 GNDA.n1489 175.546
R1820 GNDA.n1486 GNDA.n621 175.546
R1821 GNDA.n1266 GNDA.n621 175.546
R1822 GNDA.n588 GNDA.n587 175.546
R1823 GNDA.n593 GNDA.n590 175.546
R1824 GNDA.n596 GNDA.n595 175.546
R1825 GNDA.n601 GNDA.n598 175.546
R1826 GNDA.n604 GNDA.n603 175.546
R1827 GNDA.n2292 GNDA.n2291 175.546
R1828 GNDA.n2288 GNDA.n2287 175.546
R1829 GNDA.n2284 GNDA.n2283 175.546
R1830 GNDA.n2280 GNDA.n2279 175.546
R1831 GNDA.n2276 GNDA.n578 175.546
R1832 GNDA.n2460 GNDA.n612 175.546
R1833 GNDA.n2324 GNDA.n612 175.546
R1834 GNDA.n2451 GNDA.n2324 175.546
R1835 GNDA.n2451 GNDA.n2325 175.546
R1836 GNDA.n2447 GNDA.n2325 175.546
R1837 GNDA.n2447 GNDA.n2328 175.546
R1838 GNDA.n2371 GNDA.n2328 175.546
R1839 GNDA.n2380 GNDA.n2371 175.546
R1840 GNDA.n2380 GNDA.n2351 175.546
R1841 GNDA.n2385 GNDA.n2351 175.546
R1842 GNDA.n2385 GNDA.n609 175.546
R1843 GNDA.n2309 GNDA.n2274 175.546
R1844 GNDA.n2307 GNDA.n2306 175.546
R1845 GNDA.n2303 GNDA.n2302 175.546
R1846 GNDA.n2299 GNDA.n2298 175.546
R1847 GNDA.n2295 GNDA.n614 175.546
R1848 GNDA.n2317 GNDA.n614 175.546
R1849 GNDA.n1131 GNDA.n1130 175.546
R1850 GNDA.n1136 GNDA.n1133 175.546
R1851 GNDA.n1139 GNDA.n1138 175.546
R1852 GNDA.n1144 GNDA.n1141 175.546
R1853 GNDA.n1147 GNDA.n1146 175.546
R1854 GNDA.n1107 GNDA.n1106 175.546
R1855 GNDA.n1111 GNDA.n1110 175.546
R1856 GNDA.n1115 GNDA.n1114 175.546
R1857 GNDA.n1119 GNDA.n1118 175.546
R1858 GNDA.n1121 GNDA.n1079 175.546
R1859 GNDA.n2264 GNDA.n2263 175.546
R1860 GNDA.n693 GNDA.n673 175.546
R1861 GNDA.n675 GNDA.n672 175.546
R1862 GNDA.n683 GNDA.n682 175.546
R1863 GNDA.n2201 GNDA.n656 175.546
R1864 GNDA.n1099 GNDA.n1098 175.546
R1865 GNDA.n1095 GNDA.n1094 175.546
R1866 GNDA.n1091 GNDA.n1090 175.546
R1867 GNDA.n1087 GNDA.n1086 175.546
R1868 GNDA.n1083 GNDA.n1082 175.546
R1869 GNDA.n1941 GNDA.n1203 175.546
R1870 GNDA.n1945 GNDA.n1203 175.546
R1871 GNDA.n1945 GNDA.n1201 175.546
R1872 GNDA.n1950 GNDA.n1201 175.546
R1873 GNDA.n1950 GNDA.n1199 175.546
R1874 GNDA.n1954 GNDA.n1199 175.546
R1875 GNDA.n1954 GNDA.n1198 175.546
R1876 GNDA.n1959 GNDA.n1198 175.546
R1877 GNDA.n1959 GNDA.n1196 175.546
R1878 GNDA.n1963 GNDA.n1196 175.546
R1879 GNDA.n1964 GNDA.n1963 175.546
R1880 GNDA.n1920 GNDA.n1919 175.546
R1881 GNDA.n1924 GNDA.n1923 175.546
R1882 GNDA.n1928 GNDA.n1927 175.546
R1883 GNDA.n1932 GNDA.n1931 175.546
R1884 GNDA.n1936 GNDA.n1935 175.546
R1885 GNDA.n2058 GNDA.n2057 175.546
R1886 GNDA.n1974 GNDA.n1973 175.546
R1887 GNDA.n1980 GNDA.n1979 175.546
R1888 GNDA.n1987 GNDA.n1986 175.546
R1889 GNDA.n1995 GNDA.n1994 175.546
R1890 GNDA.n1912 GNDA.n1911 175.546
R1891 GNDA.n1909 GNDA.n1889 175.546
R1892 GNDA.n1905 GNDA.n1903 175.546
R1893 GNDA.n1901 GNDA.n1896 175.546
R1894 GNDA.n2193 GNDA.n1052 175.546
R1895 GNDA.n2179 GNDA.n2178 175.546
R1896 GNDA.n2175 GNDA.n2174 175.546
R1897 GNDA.n2172 GNDA.n1135 175.546
R1898 GNDA.n2168 GNDA.n2166 175.546
R1899 GNDA.n2164 GNDA.n1143 175.546
R1900 GNDA.n1865 GNDA.n1864 175.546
R1901 GNDA.n1869 GNDA.n1868 175.546
R1902 GNDA.n1873 GNDA.n1872 175.546
R1903 GNDA.n1877 GNDA.n1876 175.546
R1904 GNDA.n1881 GNDA.n1880 175.546
R1905 GNDA.n2153 GNDA.n2152 175.546
R1906 GNDA.n2069 GNDA.n2068 175.546
R1907 GNDA.n2075 GNDA.n2074 175.546
R1908 GNDA.n2082 GNDA.n2081 175.546
R1909 GNDA.n2090 GNDA.n2089 175.546
R1910 GNDA.n1887 GNDA.n1886 175.546
R1911 GNDA.n1891 GNDA.n1890 175.546
R1912 GNDA.n1893 GNDA.n1892 175.546
R1913 GNDA.n1898 GNDA.n1897 175.546
R1914 GNDA.n2191 GNDA.n1054 175.546
R1915 GNDA.n1801 GNDA.n1240 175.546
R1916 GNDA.n1801 GNDA.n1242 175.546
R1917 GNDA.n1797 GNDA.n1242 175.546
R1918 GNDA.n1797 GNDA.n1244 175.546
R1919 GNDA.n1793 GNDA.n1244 175.546
R1920 GNDA.n1793 GNDA.n1245 175.546
R1921 GNDA.n1789 GNDA.n1245 175.546
R1922 GNDA.n1789 GNDA.n1247 175.546
R1923 GNDA.n1785 GNDA.n1247 175.546
R1924 GNDA.n1785 GNDA.n1250 175.546
R1925 GNDA.n1780 GNDA.n1250 175.546
R1926 GNDA.n1825 GNDA.n1226 175.546
R1927 GNDA.n1825 GNDA.n1229 175.546
R1928 GNDA.n1821 GNDA.n1229 175.546
R1929 GNDA.n1821 GNDA.n1232 175.546
R1930 GNDA.n1817 GNDA.n1232 175.546
R1931 GNDA.n1817 GNDA.n1233 175.546
R1932 GNDA.n1813 GNDA.n1233 175.546
R1933 GNDA.n1813 GNDA.n1235 175.546
R1934 GNDA.n1809 GNDA.n1235 175.546
R1935 GNDA.n1809 GNDA.n1238 175.546
R1936 GNDA.n1805 GNDA.n1238 175.546
R1937 GNDA.n1744 GNDA.n1670 175.546
R1938 GNDA.n1748 GNDA.n1746 175.546
R1939 GNDA.n1759 GNDA.n1664 175.546
R1940 GNDA.n1763 GNDA.n1761 175.546
R1941 GNDA.n1774 GNDA.n1657 175.546
R1942 GNDA.n1831 GNDA.n1830 175.546
R1943 GNDA.n1831 GNDA.n1222 175.546
R1944 GNDA.n1837 GNDA.n1222 175.546
R1945 GNDA.n1837 GNDA.n1217 175.546
R1946 GNDA.n1843 GNDA.n1217 175.546
R1947 GNDA.n1845 GNDA.n1843 175.546
R1948 GNDA.n1846 GNDA.n1845 175.546
R1949 GNDA.n1846 GNDA.n1213 175.546
R1950 GNDA.n1852 GNDA.n1213 175.546
R1951 GNDA.n1852 GNDA.n1208 175.546
R1952 GNDA.n1858 GNDA.n1208 175.546
R1953 GNDA.n1536 GNDA.n1534 175.546
R1954 GNDA.n1542 GNDA.n1423 175.546
R1955 GNDA.n1546 GNDA.n1544 175.546
R1956 GNDA.n1556 GNDA.n1415 175.546
R1957 GNDA.n1559 GNDA.n1558 175.546
R1958 GNDA.n1469 GNDA.n1427 175.546
R1959 GNDA.n1469 GNDA.n1429 175.546
R1960 GNDA.n1465 GNDA.n1429 175.546
R1961 GNDA.n1465 GNDA.n1432 175.546
R1962 GNDA.n1461 GNDA.n1432 175.546
R1963 GNDA.n1461 GNDA.n1434 175.546
R1964 GNDA.n1457 GNDA.n1434 175.546
R1965 GNDA.n1457 GNDA.n1444 175.546
R1966 GNDA.n1453 GNDA.n1444 175.546
R1967 GNDA.n1453 GNDA.n1450 175.546
R1968 GNDA.n1450 GNDA.n1449 175.546
R1969 GNDA.n1407 GNDA.n1406 175.546
R1970 GNDA.n1323 GNDA.n1322 175.546
R1971 GNDA.n1329 GNDA.n1328 175.546
R1972 GNDA.n1336 GNDA.n1335 175.546
R1973 GNDA.n1344 GNDA.n1343 175.546
R1974 GNDA.n1833 GNDA.n1224 175.546
R1975 GNDA.n1834 GNDA.n1833 175.546
R1976 GNDA.n1834 GNDA.n1220 175.546
R1977 GNDA.n1840 GNDA.n1220 175.546
R1978 GNDA.n1841 GNDA.n1840 175.546
R1979 GNDA.n1841 GNDA.n1215 175.546
R1980 GNDA.n1848 GNDA.n1215 175.546
R1981 GNDA.n1849 GNDA.n1848 175.546
R1982 GNDA.n1849 GNDA.n1211 175.546
R1983 GNDA.n1855 GNDA.n1211 175.546
R1984 GNDA.n1856 GNDA.n1855 175.546
R1985 GNDA.n1550 GNDA.t211 172.876
R1986 GNDA.n1413 GNDA.t211 172.615
R1987 GNDA.n1588 GNDA.n1587 163.333
R1988 GNDA.n2389 GNDA.n2388 163.333
R1989 GNDA.n2205 GNDA.n2204 163.333
R1990 GNDA.n2094 GNDA.n2093 163.333
R1991 GNDA.n1999 GNDA.n1998 163.333
R1992 GNDA.n1348 GNDA.n1347 163.333
R1993 GNDA.n1770 GNDA.n1769 163.333
R1994 GNDA.n943 GNDA.n942 163.333
R1995 GNDA.n823 GNDA.n822 163.333
R1996 GNDA.n229 GNDA.n228 152
R1997 GNDA.n398 GNDA.n147 152
R1998 GNDA.n60 GNDA.n59 150
R1999 GNDA.n60 GNDA.n51 150
R2000 GNDA.n68 GNDA.n51 150
R2001 GNDA.n69 GNDA.n68 150
R2002 GNDA.n70 GNDA.n47 150
R2003 GNDA.n78 GNDA.n47 150
R2004 GNDA.n79 GNDA.n78 150
R2005 GNDA.n80 GNDA.n79 150
R2006 GNDA.n346 GNDA.n263 150
R2007 GNDA.n264 GNDA.n263 150
R2008 GNDA.n265 GNDA.n264 150
R2009 GNDA.n266 GNDA.n265 150
R2010 GNDA.n268 GNDA.n267 150
R2011 GNDA.n269 GNDA.n268 150
R2012 GNDA.n270 GNDA.n269 150
R2013 GNDA.n271 GNDA.n270 150
R2014 GNDA.n289 GNDA.n288 150
R2015 GNDA.n289 GNDA.n280 150
R2016 GNDA.n297 GNDA.n280 150
R2017 GNDA.n298 GNDA.n297 150
R2018 GNDA.n299 GNDA.n276 150
R2019 GNDA.n307 GNDA.n276 150
R2020 GNDA.n308 GNDA.n307 150
R2021 GNDA.n309 GNDA.n308 150
R2022 GNDA.n117 GNDA.n34 150
R2023 GNDA.n35 GNDA.n34 150
R2024 GNDA.n36 GNDA.n35 150
R2025 GNDA.n37 GNDA.n36 150
R2026 GNDA.n39 GNDA.n38 150
R2027 GNDA.n40 GNDA.n39 150
R2028 GNDA.n41 GNDA.n40 150
R2029 GNDA.n42 GNDA.n41 150
R2030 GNDA.n1620 GNDA.n1619 150
R2031 GNDA.n1616 GNDA.n1615 150
R2032 GNDA.n1612 GNDA.n1611 150
R2033 GNDA.n1608 GNDA.n1607 150
R2034 GNDA.n1604 GNDA.n1603 150
R2035 GNDA.n1600 GNDA.n1599 150
R2036 GNDA.n1596 GNDA.n1595 150
R2037 GNDA.n1592 GNDA.n1591 150
R2038 GNDA.n1649 GNDA.n1648 150
R2039 GNDA.n1641 GNDA.n1275 150
R2040 GNDA.n1573 GNDA.n1276 150
R2041 GNDA.n1580 GNDA.n1579 150
R2042 GNDA.n1638 GNDA.n1292 150
R2043 GNDA.n1634 GNDA.n1633 150
R2044 GNDA.n1630 GNDA.n1629 150
R2045 GNDA.n1626 GNDA.n1625 150
R2046 GNDA.n2421 GNDA.n2420 150
R2047 GNDA.n2417 GNDA.n2416 150
R2048 GNDA.n2413 GNDA.n2412 150
R2049 GNDA.n2409 GNDA.n2408 150
R2050 GNDA.n2405 GNDA.n2404 150
R2051 GNDA.n2401 GNDA.n2400 150
R2052 GNDA.n2397 GNDA.n2396 150
R2053 GNDA.n2393 GNDA.n2392 150
R2054 GNDA.n2455 GNDA.n2454 150
R2055 GNDA.n2442 GNDA.n2441 150
R2056 GNDA.n2444 GNDA.n2331 150
R2057 GNDA.n2377 GNDA.n2376 150
R2058 GNDA.n2439 GNDA.n2347 150
R2059 GNDA.n2435 GNDA.n2434 150
R2060 GNDA.n2431 GNDA.n2430 150
R2061 GNDA.n2427 GNDA.n2426 150
R2062 GNDA.n2237 GNDA.n2236 150
R2063 GNDA.n2233 GNDA.n2232 150
R2064 GNDA.n2229 GNDA.n2228 150
R2065 GNDA.n2225 GNDA.n2224 150
R2066 GNDA.n2221 GNDA.n2220 150
R2067 GNDA.n2217 GNDA.n2216 150
R2068 GNDA.n2213 GNDA.n2212 150
R2069 GNDA.n2209 GNDA.n2208 150
R2070 GNDA.n2260 GNDA.n636 150
R2071 GNDA.n690 GNDA.n637 150
R2072 GNDA.n687 GNDA.n686 150
R2073 GNDA.n679 GNDA.n678 150
R2074 GNDA.n2245 GNDA.n2244 150
R2075 GNDA.n2249 GNDA.n2248 150
R2076 GNDA.n2253 GNDA.n2252 150
R2077 GNDA.n2257 GNDA.n2256 150
R2078 GNDA.n2126 GNDA.n2125 150
R2079 GNDA.n2122 GNDA.n2121 150
R2080 GNDA.n2118 GNDA.n2117 150
R2081 GNDA.n2114 GNDA.n2113 150
R2082 GNDA.n2110 GNDA.n2109 150
R2083 GNDA.n2106 GNDA.n2105 150
R2084 GNDA.n2102 GNDA.n2101 150
R2085 GNDA.n2098 GNDA.n2097 150
R2086 GNDA.n2149 GNDA.n1154 150
R2087 GNDA.n2071 GNDA.n1155 150
R2088 GNDA.n2079 GNDA.n2078 150
R2089 GNDA.n2086 GNDA.n2085 150
R2090 GNDA.n2134 GNDA.n2133 150
R2091 GNDA.n2138 GNDA.n2137 150
R2092 GNDA.n2142 GNDA.n2141 150
R2093 GNDA.n2146 GNDA.n2145 150
R2094 GNDA.n2031 GNDA.n2030 150
R2095 GNDA.n2027 GNDA.n2026 150
R2096 GNDA.n2023 GNDA.n2022 150
R2097 GNDA.n2019 GNDA.n2018 150
R2098 GNDA.n2015 GNDA.n2014 150
R2099 GNDA.n2011 GNDA.n2010 150
R2100 GNDA.n2007 GNDA.n2006 150
R2101 GNDA.n2003 GNDA.n2002 150
R2102 GNDA.n2054 GNDA.n1175 150
R2103 GNDA.n1976 GNDA.n1176 150
R2104 GNDA.n1984 GNDA.n1983 150
R2105 GNDA.n1991 GNDA.n1990 150
R2106 GNDA.n2039 GNDA.n2038 150
R2107 GNDA.n2043 GNDA.n2042 150
R2108 GNDA.n2047 GNDA.n2046 150
R2109 GNDA.n2051 GNDA.n2050 150
R2110 GNDA.n1380 GNDA.n1379 150
R2111 GNDA.n1376 GNDA.n1375 150
R2112 GNDA.n1372 GNDA.n1371 150
R2113 GNDA.n1368 GNDA.n1367 150
R2114 GNDA.n1364 GNDA.n1363 150
R2115 GNDA.n1360 GNDA.n1359 150
R2116 GNDA.n1356 GNDA.n1355 150
R2117 GNDA.n1352 GNDA.n1351 150
R2118 GNDA.n1403 GNDA.n1299 150
R2119 GNDA.n1325 GNDA.n1300 150
R2120 GNDA.n1333 GNDA.n1332 150
R2121 GNDA.n1340 GNDA.n1339 150
R2122 GNDA.n1388 GNDA.n1387 150
R2123 GNDA.n1392 GNDA.n1391 150
R2124 GNDA.n1396 GNDA.n1395 150
R2125 GNDA.n1400 GNDA.n1399 150
R2126 GNDA.n1714 GNDA.n1712 150
R2127 GNDA.n1710 GNDA.n1678 150
R2128 GNDA.n1706 GNDA.n1704 150
R2129 GNDA.n1702 GNDA.n1680 150
R2130 GNDA.n1698 GNDA.n1696 150
R2131 GNDA.n1694 GNDA.n1682 150
R2132 GNDA.n1690 GNDA.n1689 150
R2133 GNDA.n1687 GNDA.n1685 150
R2134 GNDA.n1741 GNDA.n1739 150
R2135 GNDA.n1752 GNDA.n1666 150
R2136 GNDA.n1756 GNDA.n1754 150
R2137 GNDA.n1767 GNDA.n1661 150
R2138 GNDA.n1722 GNDA.n1720 150
R2139 GNDA.n1726 GNDA.n1674 150
R2140 GNDA.n1730 GNDA.n1728 150
R2141 GNDA.n1737 GNDA.n1672 150
R2142 GNDA.n975 GNDA.n974 150
R2143 GNDA.n971 GNDA.n970 150
R2144 GNDA.n967 GNDA.n966 150
R2145 GNDA.n963 GNDA.n962 150
R2146 GNDA.n959 GNDA.n958 150
R2147 GNDA.n955 GNDA.n954 150
R2148 GNDA.n951 GNDA.n950 150
R2149 GNDA.n947 GNDA.n946 150
R2150 GNDA.n1010 GNDA.n1009 150
R2151 GNDA.n997 GNDA.n996 150
R2152 GNDA.n999 GNDA.n898 150
R2153 GNDA.n931 GNDA.n930 150
R2154 GNDA.n994 GNDA.n914 150
R2155 GNDA.n990 GNDA.n989 150
R2156 GNDA.n986 GNDA.n985 150
R2157 GNDA.n982 GNDA.n981 150
R2158 GNDA.n855 GNDA.n854 150
R2159 GNDA.n851 GNDA.n850 150
R2160 GNDA.n847 GNDA.n846 150
R2161 GNDA.n843 GNDA.n842 150
R2162 GNDA.n839 GNDA.n838 150
R2163 GNDA.n835 GNDA.n834 150
R2164 GNDA.n831 GNDA.n830 150
R2165 GNDA.n827 GNDA.n826 150
R2166 GNDA.n2546 GNDA.n549 150
R2167 GNDA.n2536 GNDA.n2535 150
R2168 GNDA.n2549 GNDA.n530 150
R2169 GNDA.n812 GNDA.n531 150
R2170 GNDA.n863 GNDA.n862 150
R2171 GNDA.n867 GNDA.n866 150
R2172 GNDA.n871 GNDA.n870 150
R2173 GNDA.n873 GNDA.n548 150
R2174 GNDA.t74 GNDA.t153 147.84
R2175 GNDA.t297 GNDA.t299 144.321
R2176 GNDA.n2466 GNDA.n2465 139.077
R2177 GNDA.n2468 GNDA.n2467 139.077
R2178 GNDA.n2470 GNDA.n2469 139.077
R2179 GNDA.n2476 GNDA.n2475 139.077
R2180 GNDA.n2474 GNDA.n2473 139.077
R2181 GNDA.n2472 GNDA.n2471 139.077
R2182 GNDA.n555 GNDA.n554 139.077
R2183 GNDA.n2521 GNDA.n2520 139.077
R2184 GNDA.n2519 GNDA.n2518 139.077
R2185 GNDA.n515 GNDA.n514 139.077
R2186 GNDA.t12 GNDA.t131 139.041
R2187 GNDA.n2570 GNDA.t93 135.69
R2188 GNDA.n2357 GNDA.n2355 134.268
R2189 GNDA.n2365 GNDA.n2357 134.268
R2190 GNDA.n629 GNDA.n628 132.721
R2191 GNDA.n2575 GNDA.t253 130.001
R2192 GNDA.n2524 GNDA.t264 130.001
R2193 GNDA.n2515 GNDA.t244 130.001
R2194 GNDA.n2477 GNDA.t288 130.001
R2195 GNDA.n2482 GNDA.t267 130.001
R2196 GNDA.n2463 GNDA.t259 130.001
R2197 GNDA.n1024 GNDA.n1022 124.832
R2198 GNDA.n1020 GNDA.n745 124.832
R2199 GNDA.n882 GNDA.n606 124.832
R2200 GNDA.n1564 GNDA.n1563 124.832
R2201 GNDA.n2486 GNDA.n2485 124.832
R2202 GNDA.n1149 GNDA.n696 124.832
R2203 GNDA.n2196 GNDA.n2195 124.832
R2204 GNDA.n2160 GNDA.n695 124.832
R2205 GNDA.n2189 GNDA.n697 124.832
R2206 GNDA.n1859 GNDA.n1858 124.832
R2207 GNDA.n1561 GNDA.n1412 124.832
R2208 GNDA.n1856 GNDA.n1205 124.832
R2209 GNDA.n517 GNDA.t13 115.948
R2210 GNDA.n1437 GNDA.t51 115.105
R2211 GNDA.n517 GNDA.t298 114.635
R2212 GNDA.n1438 GNDA.t125 114.635
R2213 GNDA.n456 GNDA.n128 107.975
R2214 GNDA.n454 GNDA.n411 107.975
R2215 GNDA.n476 GNDA.t205 103.665
R2216 GNDA.n393 GNDA.t202 103.665
R2217 GNDA.t243 GNDA.n556 101.942
R2218 GNDA.n2554 GNDA.n523 101.718
R2219 GNDA.n447 GNDA.n138 101.718
R2220 GNDA.n438 GNDA.n437 101.718
R2221 GNDA.n392 GNDA.n391 101.718
R2222 GNDA.n405 GNDA.n139 101.718
R2223 GNDA.n462 GNDA.n461 101.718
R2224 GNDA.n475 GNDA.n474 101.718
R2225 GNDA.n356 GNDA.n350 101.718
R2226 GNDA.n372 GNDA.n233 101.718
R2227 GNDA.n482 GNDA.n121 101.718
R2228 GNDA.n498 GNDA.n15 101.718
R2229 GNDA.n343 GNDA.n254 101.718
R2230 GNDA.n340 GNDA.n255 101.718
R2231 GNDA.n336 GNDA.n256 101.718
R2232 GNDA.n332 GNDA.n257 101.718
R2233 GNDA.n328 GNDA.n258 101.718
R2234 GNDA.n292 GNDA.n291 101.718
R2235 GNDA.n295 GNDA.n294 101.718
R2236 GNDA.n302 GNDA.n301 101.718
R2237 GNDA.n305 GNDA.n304 101.718
R2238 GNDA.n312 GNDA.n311 101.718
R2239 GNDA.n114 GNDA.n25 101.718
R2240 GNDA.n111 GNDA.n26 101.718
R2241 GNDA.n107 GNDA.n27 101.718
R2242 GNDA.n103 GNDA.n28 101.718
R2243 GNDA.n99 GNDA.n29 101.718
R2244 GNDA.n159 GNDA.n158 101.718
R2245 GNDA.n204 GNDA.n185 101.718
R2246 GNDA.n63 GNDA.n62 101.718
R2247 GNDA.n66 GNDA.n65 101.718
R2248 GNDA.n73 GNDA.n72 101.718
R2249 GNDA.n76 GNDA.n75 101.718
R2250 GNDA.n83 GNDA.n82 101.718
R2251 GNDA.n56 GNDA.n55 101.718
R2252 GNDA.n64 GNDA.n63 101.718
R2253 GNDA.n65 GNDA.n49 101.718
R2254 GNDA.n74 GNDA.n73 101.718
R2255 GNDA.n75 GNDA.n45 101.718
R2256 GNDA.n84 GNDA.n83 101.718
R2257 GNDA.n136 GNDA.n130 101.718
R2258 GNDA.n2594 GNDA.n5 101.718
R2259 GNDA.n202 GNDA.n195 101.718
R2260 GNDA.n152 GNDA.n151 101.718
R2261 GNDA.n119 GNDA.n32 101.718
R2262 GNDA.n112 GNDA.n25 101.718
R2263 GNDA.n108 GNDA.n26 101.718
R2264 GNDA.n104 GNDA.n27 101.718
R2265 GNDA.n100 GNDA.n28 101.718
R2266 GNDA.n96 GNDA.n29 101.718
R2267 GNDA.n285 GNDA.n284 101.718
R2268 GNDA.n293 GNDA.n292 101.718
R2269 GNDA.n294 GNDA.n278 101.718
R2270 GNDA.n303 GNDA.n302 101.718
R2271 GNDA.n304 GNDA.n274 101.718
R2272 GNDA.n313 GNDA.n312 101.718
R2273 GNDA.n348 GNDA.n261 101.718
R2274 GNDA.n341 GNDA.n254 101.718
R2275 GNDA.n337 GNDA.n255 101.718
R2276 GNDA.n333 GNDA.n256 101.718
R2277 GNDA.n329 GNDA.n257 101.718
R2278 GNDA.n325 GNDA.n258 101.718
R2279 GNDA.n503 GNDA.n19 101.718
R2280 GNDA.n496 GNDA.n15 101.718
R2281 GNDA.n210 GNDA.n123 101.718
R2282 GNDA.n225 GNDA.n224 101.718
R2283 GNDA.n403 GNDA.n143 101.718
R2284 GNDA.n382 GNDA.n232 101.718
R2285 GNDA.n487 GNDA.n478 101.718
R2286 GNDA.n121 GNDA.n24 101.718
R2287 GNDA.n377 GNDA.n237 101.718
R2288 GNDA.n370 GNDA.n233 101.718
R2289 GNDA.n361 GNDA.n352 101.718
R2290 GNDA.n350 GNDA.n253 101.718
R2291 GNDA.n431 GNDA.n430 101.718
R2292 GNDA.n453 GNDA.n413 101.718
R2293 GNDA.n2565 GNDA.n522 101.718
R2294 GNDA.n2354 GNDA.n2352 101.718
R2295 GNDA.n2361 GNDA.n2353 101.718
R2296 GNDA.n2360 GNDA.n2352 101.718
R2297 GNDA.n443 GNDA.n442 100.684
R2298 GNDA.n2187 GNDA.t211 47.6748
R2299 GNDA.n2513 GNDA.t211 47.6748
R2300 GNDA.n183 GNDA.n182 99.0842
R2301 GNDA.n181 GNDA.n180 99.0842
R2302 GNDA.n179 GNDA.n178 99.0842
R2303 GNDA.n177 GNDA.n176 99.0842
R2304 GNDA.n175 GNDA.n174 99.0842
R2305 GNDA.n173 GNDA.n172 99.0842
R2306 GNDA.n171 GNDA.n170 99.0842
R2307 GNDA.n169 GNDA.n168 99.0842
R2308 GNDA.n167 GNDA.n166 99.0842
R2309 GNDA.n165 GNDA.n164 99.0842
R2310 GNDA.n163 GNDA.n162 99.0842
R2311 GNDA.n783 GNDA.t211 98.9756
R2312 GNDA.n884 GNDA.n883 98.8538
R2313 GNDA.n89 GNDA.n88 94.601
R2314 GNDA.n321 GNDA.n320 94.601
R2315 GNDA.n318 GNDA.n317 94.601
R2316 GNDA.n92 GNDA.n91 94.601
R2317 GNDA.n2527 GNDA.n2526 92.6754
R2318 GNDA.t44 GNDA.t56 92.1471
R2319 GNDA.t56 GNDA.t315 92.1471
R2320 GNDA.t315 GNDA.t10 92.1471
R2321 GNDA.t127 GNDA.t300 92.1471
R2322 GNDA.n2561 GNDA.n521 91.069
R2323 GNDA.n2556 GNDA.n521 91.069
R2324 GNDA.n2558 GNDA.n520 91.069
R2325 GNDA.n2559 GNDA.n2558 91.069
R2326 GNDA.n222 GNDA.n219 91.069
R2327 GNDA.n221 GNDA.n218 91.069
R2328 GNDA.n401 GNDA.n400 91.069
R2329 GNDA.n146 GNDA.n144 91.069
R2330 GNDA.n2363 GNDA.n2355 91.069
R2331 GNDA.n2365 GNDA.n2358 91.069
R2332 GNDA.t266 GNDA.n2383 90.616
R2333 GNDA.n214 GNDA.n213 90.4158
R2334 GNDA.n199 GNDA.n196 90.2704
R2335 GNDA.n196 GNDA.n184 90.2704
R2336 GNDA.n155 GNDA.n154 90.2704
R2337 GNDA.n154 GNDA.n148 90.2704
R2338 GNDA.n379 GNDA.n231 90.2704
R2339 GNDA.n472 GNDA.n471 90.2704
R2340 GNDA.n458 GNDA.n126 90.2704
R2341 GNDA.n407 GNDA.n140 90.2704
R2342 GNDA.n389 GNDA.n388 90.2704
R2343 GNDA.n434 GNDA.n433 90.2704
R2344 GNDA.n433 GNDA.n427 90.2704
R2345 GNDA.n450 GNDA.n414 90.2704
R2346 GNDA.n446 GNDA.n414 90.2704
R2347 GNDA.n133 GNDA.n131 90.2704
R2348 GNDA.n2591 GNDA.n4 90.2704
R2349 GNDA.n1940 GNDA.t2 89.6052
R2350 GNDA.n1509 GNDA.n1483 88.5317
R2351 GNDA.n1510 GNDA.n1509 88.5317
R2352 GNDA.n1511 GNDA.n1510 88.5317
R2353 GNDA.n1511 GNDA.n1479 88.5317
R2354 GNDA.n1517 GNDA.n1479 88.5317
R2355 GNDA.n1519 GNDA.n1518 88.5317
R2356 GNDA.n1519 GNDA.n1475 88.5317
R2357 GNDA.n1526 GNDA.n1475 88.5317
R2358 GNDA.n1527 GNDA.n1526 88.5317
R2359 GNDA.n1528 GNDA.n1527 88.5317
R2360 GNDA.n1468 GNDA.n1430 88.5317
R2361 GNDA.n1468 GNDA.n1467 88.5317
R2362 GNDA.n1467 GNDA.n1466 88.5317
R2363 GNDA.n1466 GNDA.n1431 88.5317
R2364 GNDA.n1460 GNDA.n1431 88.5317
R2365 GNDA.n1459 GNDA.n1458 88.5317
R2366 GNDA.n1458 GNDA.n1443 88.5317
R2367 GNDA.n1452 GNDA.n1443 88.5317
R2368 GNDA.n1452 GNDA.n1451 88.5317
R2369 GNDA.n1451 GNDA.n1227 88.5317
R2370 GNDA.n1827 GNDA.n1826 88.5317
R2371 GNDA.n1826 GNDA.n1228 88.5317
R2372 GNDA.n1820 GNDA.n1228 88.5317
R2373 GNDA.n1820 GNDA.n1819 88.5317
R2374 GNDA.n1819 GNDA.n1818 88.5317
R2375 GNDA.n1812 GNDA.n1236 88.5317
R2376 GNDA.n1812 GNDA.n1811 88.5317
R2377 GNDA.n1811 GNDA.n1810 88.5317
R2378 GNDA.n1810 GNDA.n1237 88.5317
R2379 GNDA.n1804 GNDA.n1237 88.5317
R2380 GNDA.t300 GNDA.n504 88.3077
R2381 GNDA.t151 GNDA.n2577 85.4674
R2382 GNDA.t90 GNDA.t32 84.4682
R2383 GNDA.t88 GNDA.t6 84.4682
R2384 GNDA.t98 GNDA.t41 84.4682
R2385 GNDA.t94 GNDA.t97 84.4682
R2386 GNDA.t78 GNDA.t96 84.4682
R2387 GNDA.t307 GNDA.t24 84.4682
R2388 GNDA.t54 GNDA.t21 84.4682
R2389 GNDA.t146 GNDA.t154 84.4682
R2390 GNDA.t17 GNDA.t28 84.4682
R2391 GNDA.t143 GNDA.t293 84.4682
R2392 GNDA.n1004 GNDA.t175 84.4377
R2393 GNDA.n1436 GNDA.n1435 84.306
R2394 GNDA.t73 GNDA.t18 82.3782
R2395 GNDA.t104 GNDA.t92 82.3782
R2396 GNDA.n1829 GNDA.n1828 80.9821
R2397 GNDA.t271 GNDA.t220 80.6288
R2398 GNDA.t246 GNDA.t255 80.6288
R2399 GNDA.t249 GNDA.t199 80.6288
R2400 GNDA.t215 GNDA.t234 80.6288
R2401 GNDA.n935 GNDA.t163 80.3188
R2402 GNDA.t238 GNDA.t102 76.7893
R2403 GNDA.t87 GNDA.t141 76.7893
R2404 GNDA.t75 GNDA.t69 76.7893
R2405 GNDA.n762 GNDA.n561 76.3222
R2406 GNDA.n766 GNDA.n562 76.3222
R2407 GNDA.n770 GNDA.n563 76.3222
R2408 GNDA.n774 GNDA.n564 76.3222
R2409 GNDA.n778 GNDA.n565 76.3222
R2410 GNDA.n782 GNDA.n566 76.3222
R2411 GNDA.n1045 GNDA.n1044 76.3222
R2412 GNDA.n1042 GNDA.n724 76.3222
R2413 GNDA.n1038 GNDA.n1037 76.3222
R2414 GNDA.n1031 GNDA.n731 76.3222
R2415 GNDA.n1030 GNDA.n1029 76.3222
R2416 GNDA.n1023 GNDA.n739 76.3222
R2417 GNDA.n726 GNDA.n725 76.3222
R2418 GNDA.n729 GNDA.n728 76.3222
R2419 GNDA.n734 GNDA.n733 76.3222
R2420 GNDA.n737 GNDA.n736 76.3222
R2421 GNDA.n742 GNDA.n741 76.3222
R2422 GNDA.n745 GNDA.n744 76.3222
R2423 GNDA.n700 GNDA.n567 76.3222
R2424 GNDA.n704 GNDA.n568 76.3222
R2425 GNDA.n708 GNDA.n569 76.3222
R2426 GNDA.n712 GNDA.n570 76.3222
R2427 GNDA.n716 GNDA.n571 76.3222
R2428 GNDA.n720 GNDA.n572 76.3222
R2429 GNDA.n2507 GNDA.n2506 76.3222
R2430 GNDA.n2504 GNDA.n585 76.3222
R2431 GNDA.n2500 GNDA.n2499 76.3222
R2432 GNDA.n2493 GNDA.n592 76.3222
R2433 GNDA.n2492 GNDA.n2491 76.3222
R2434 GNDA.n605 GNDA.n600 76.3222
R2435 GNDA.n1425 GNDA.n1418 76.3222
R2436 GNDA.n1539 GNDA.n1419 76.3222
R2437 GNDA.n1421 GNDA.n1420 76.3222
R2438 GNDA.n1549 GNDA.n1417 76.3222
R2439 GNDA.n1553 GNDA.n1552 76.3222
R2440 GNDA.n1563 GNDA.n1294 76.3222
R2441 GNDA.n1655 GNDA.n1654 76.3222
R2442 GNDA.n1269 GNDA.n1263 76.3222
R2443 GNDA.n1644 GNDA.n1262 76.3222
R2444 GNDA.n1571 GNDA.n1261 76.3222
R2445 GNDA.n1575 GNDA.n1260 76.3222
R2446 GNDA.n1584 GNDA.n1259 76.3222
R2447 GNDA.n1504 GNDA.n616 76.3222
R2448 GNDA.n1501 GNDA.n617 76.3222
R2449 GNDA.n1497 GNDA.n618 76.3222
R2450 GNDA.n1493 GNDA.n619 76.3222
R2451 GNDA.n1489 GNDA.n620 76.3222
R2452 GNDA.n587 GNDA.n586 76.3222
R2453 GNDA.n590 GNDA.n589 76.3222
R2454 GNDA.n595 GNDA.n594 76.3222
R2455 GNDA.n598 GNDA.n597 76.3222
R2456 GNDA.n603 GNDA.n602 76.3222
R2457 GNDA.n2486 GNDA.n608 76.3222
R2458 GNDA.n2292 GNDA.n573 76.3222
R2459 GNDA.n2288 GNDA.n574 76.3222
R2460 GNDA.n2284 GNDA.n575 76.3222
R2461 GNDA.n2280 GNDA.n576 76.3222
R2462 GNDA.n2276 GNDA.n577 76.3222
R2463 GNDA.n2512 GNDA.n2511 76.3222
R2464 GNDA.n2314 GNDA.n2313 76.3222
R2465 GNDA.n2309 GNDA.n2273 76.3222
R2466 GNDA.n2306 GNDA.n2272 76.3222
R2467 GNDA.n2302 GNDA.n2271 76.3222
R2468 GNDA.n2298 GNDA.n2270 76.3222
R2469 GNDA.n2314 GNDA.n2274 76.3222
R2470 GNDA.n2307 GNDA.n2273 76.3222
R2471 GNDA.n2303 GNDA.n2272 76.3222
R2472 GNDA.n2299 GNDA.n2271 76.3222
R2473 GNDA.n2295 GNDA.n2270 76.3222
R2474 GNDA.n1502 GNDA.n616 76.3222
R2475 GNDA.n1498 GNDA.n617 76.3222
R2476 GNDA.n1494 GNDA.n618 76.3222
R2477 GNDA.n1490 GNDA.n619 76.3222
R2478 GNDA.n1486 GNDA.n620 76.3222
R2479 GNDA.n1130 GNDA.n1129 76.3222
R2480 GNDA.n1133 GNDA.n1132 76.3222
R2481 GNDA.n1138 GNDA.n1137 76.3222
R2482 GNDA.n1141 GNDA.n1140 76.3222
R2483 GNDA.n1146 GNDA.n1145 76.3222
R2484 GNDA.n1149 GNDA.n1148 76.3222
R2485 GNDA.n1106 GNDA.n1074 76.3222
R2486 GNDA.n1110 GNDA.n1075 76.3222
R2487 GNDA.n1114 GNDA.n1076 76.3222
R2488 GNDA.n1118 GNDA.n1077 76.3222
R2489 GNDA.n1121 GNDA.n1078 76.3222
R2490 GNDA.n2186 GNDA.n2185 76.3222
R2491 GNDA.n2268 GNDA.n630 76.3222
R2492 GNDA.n2263 GNDA.n634 76.3222
R2493 GNDA.n694 GNDA.n693 76.3222
R2494 GNDA.n675 GNDA.n671 76.3222
R2495 GNDA.n682 GNDA.n670 76.3222
R2496 GNDA.n2201 GNDA.n2200 76.3222
R2497 GNDA.n1102 GNDA.n623 76.3222
R2498 GNDA.n1098 GNDA.n624 76.3222
R2499 GNDA.n1094 GNDA.n625 76.3222
R2500 GNDA.n1090 GNDA.n626 76.3222
R2501 GNDA.n1086 GNDA.n627 76.3222
R2502 GNDA.n1082 GNDA.n628 76.3222
R2503 GNDA.n1099 GNDA.n623 76.3222
R2504 GNDA.n1095 GNDA.n624 76.3222
R2505 GNDA.n1091 GNDA.n625 76.3222
R2506 GNDA.n1087 GNDA.n626 76.3222
R2507 GNDA.n1083 GNDA.n627 76.3222
R2508 GNDA.n1919 GNDA.n1062 76.3222
R2509 GNDA.n1923 GNDA.n1063 76.3222
R2510 GNDA.n1927 GNDA.n1064 76.3222
R2511 GNDA.n1931 GNDA.n1065 76.3222
R2512 GNDA.n1935 GNDA.n1066 76.3222
R2513 GNDA.n1939 GNDA.n1067 76.3222
R2514 GNDA.n1049 GNDA.n663 76.3222
R2515 GNDA.n2057 GNDA.n662 76.3222
R2516 GNDA.n1974 GNDA.n661 76.3222
R2517 GNDA.n1980 GNDA.n660 76.3222
R2518 GNDA.n1986 GNDA.n659 76.3222
R2519 GNDA.n1995 GNDA.n658 76.3222
R2520 GNDA.n1915 GNDA.n1862 76.3222
R2521 GNDA.n1911 GNDA.n1910 76.3222
R2522 GNDA.n1904 GNDA.n1889 76.3222
R2523 GNDA.n1903 GNDA.n1902 76.3222
R2524 GNDA.n1896 GNDA.n1895 76.3222
R2525 GNDA.n2194 GNDA.n2193 76.3222
R2526 GNDA.n2181 GNDA.n2180 76.3222
R2527 GNDA.n2178 GNDA.n1128 76.3222
R2528 GNDA.n2174 GNDA.n2173 76.3222
R2529 GNDA.n2167 GNDA.n1135 76.3222
R2530 GNDA.n2166 GNDA.n2165 76.3222
R2531 GNDA.n2159 GNDA.n1143 76.3222
R2532 GNDA.n1864 GNDA.n1068 76.3222
R2533 GNDA.n1868 GNDA.n1069 76.3222
R2534 GNDA.n1872 GNDA.n1070 76.3222
R2535 GNDA.n1876 GNDA.n1071 76.3222
R2536 GNDA.n1880 GNDA.n1072 76.3222
R2537 GNDA.n1884 GNDA.n1073 76.3222
R2538 GNDA.n2156 GNDA.n669 76.3222
R2539 GNDA.n2152 GNDA.n668 76.3222
R2540 GNDA.n2069 GNDA.n667 76.3222
R2541 GNDA.n2075 GNDA.n666 76.3222
R2542 GNDA.n2081 GNDA.n665 76.3222
R2543 GNDA.n2090 GNDA.n664 76.3222
R2544 GNDA.n1886 GNDA.n1055 76.3222
R2545 GNDA.n1890 GNDA.n1056 76.3222
R2546 GNDA.n1892 GNDA.n1057 76.3222
R2547 GNDA.n1897 GNDA.n1058 76.3222
R2548 GNDA.n1059 GNDA.n1054 76.3222
R2549 GNDA.n2190 GNDA.n2189 76.3222
R2550 GNDA.n1669 GNDA.n1207 76.3222
R2551 GNDA.n1745 GNDA.n1744 76.3222
R2552 GNDA.n1748 GNDA.n1747 76.3222
R2553 GNDA.n1760 GNDA.n1759 76.3222
R2554 GNDA.n1763 GNDA.n1762 76.3222
R2555 GNDA.n1775 GNDA.n1774 76.3222
R2556 GNDA.n1533 GNDA.n1532 76.3222
R2557 GNDA.n1536 GNDA.n1535 76.3222
R2558 GNDA.n1543 GNDA.n1542 76.3222
R2559 GNDA.n1546 GNDA.n1545 76.3222
R2560 GNDA.n1557 GNDA.n1556 76.3222
R2561 GNDA.n1560 GNDA.n1559 76.3222
R2562 GNDA.n1411 GNDA.n1258 76.3222
R2563 GNDA.n1406 GNDA.n1257 76.3222
R2564 GNDA.n1323 GNDA.n1256 76.3222
R2565 GNDA.n1329 GNDA.n1255 76.3222
R2566 GNDA.n1335 GNDA.n1254 76.3222
R2567 GNDA.n1344 GNDA.n1253 76.3222
R2568 GNDA.n2191 GNDA.n2190 76.3222
R2569 GNDA.n1898 GNDA.n1059 76.3222
R2570 GNDA.n1893 GNDA.n1058 76.3222
R2571 GNDA.n1891 GNDA.n1057 76.3222
R2572 GNDA.n1887 GNDA.n1056 76.3222
R2573 GNDA.n1885 GNDA.n1055 76.3222
R2574 GNDA.n1912 GNDA.n1862 76.3222
R2575 GNDA.n1910 GNDA.n1909 76.3222
R2576 GNDA.n1905 GNDA.n1904 76.3222
R2577 GNDA.n1902 GNDA.n1901 76.3222
R2578 GNDA.n1895 GNDA.n1052 76.3222
R2579 GNDA.n2195 GNDA.n2194 76.3222
R2580 GNDA.n2186 GNDA.n1079 76.3222
R2581 GNDA.n1119 GNDA.n1078 76.3222
R2582 GNDA.n1115 GNDA.n1077 76.3222
R2583 GNDA.n1111 GNDA.n1076 76.3222
R2584 GNDA.n1107 GNDA.n1075 76.3222
R2585 GNDA.n1103 GNDA.n1074 76.3222
R2586 GNDA.n1881 GNDA.n1073 76.3222
R2587 GNDA.n1877 GNDA.n1072 76.3222
R2588 GNDA.n1873 GNDA.n1071 76.3222
R2589 GNDA.n1869 GNDA.n1070 76.3222
R2590 GNDA.n1865 GNDA.n1069 76.3222
R2591 GNDA.n1127 GNDA.n1068 76.3222
R2592 GNDA.n1936 GNDA.n1067 76.3222
R2593 GNDA.n1932 GNDA.n1066 76.3222
R2594 GNDA.n1928 GNDA.n1065 76.3222
R2595 GNDA.n1924 GNDA.n1064 76.3222
R2596 GNDA.n1920 GNDA.n1063 76.3222
R2597 GNDA.n1916 GNDA.n1062 76.3222
R2598 GNDA.n1655 GNDA.n1264 76.3222
R2599 GNDA.n1645 GNDA.n1263 76.3222
R2600 GNDA.n1570 GNDA.n1262 76.3222
R2601 GNDA.n1576 GNDA.n1261 76.3222
R2602 GNDA.n1583 GNDA.n1260 76.3222
R2603 GNDA.n1565 GNDA.n1259 76.3222
R2604 GNDA.n1407 GNDA.n1258 76.3222
R2605 GNDA.n1322 GNDA.n1257 76.3222
R2606 GNDA.n1328 GNDA.n1256 76.3222
R2607 GNDA.n1336 GNDA.n1255 76.3222
R2608 GNDA.n1343 GNDA.n1254 76.3222
R2609 GNDA.n1317 GNDA.n1253 76.3222
R2610 GNDA.n1670 GNDA.n1669 76.3222
R2611 GNDA.n1746 GNDA.n1745 76.3222
R2612 GNDA.n1747 GNDA.n1664 76.3222
R2613 GNDA.n1761 GNDA.n1760 76.3222
R2614 GNDA.n1762 GNDA.n1657 76.3222
R2615 GNDA.n1776 GNDA.n1775 76.3222
R2616 GNDA.n1551 GNDA.n1294 76.3222
R2617 GNDA.n1554 GNDA.n1553 76.3222
R2618 GNDA.n1549 GNDA.n1548 76.3222
R2619 GNDA.n1540 GNDA.n1420 76.3222
R2620 GNDA.n1426 GNDA.n1419 76.3222
R2621 GNDA.n1530 GNDA.n1418 76.3222
R2622 GNDA.n1534 GNDA.n1533 76.3222
R2623 GNDA.n1535 GNDA.n1423 76.3222
R2624 GNDA.n1544 GNDA.n1543 76.3222
R2625 GNDA.n1545 GNDA.n1415 76.3222
R2626 GNDA.n1558 GNDA.n1557 76.3222
R2627 GNDA.n1561 GNDA.n1560 76.3222
R2628 GNDA.n1148 GNDA.n1147 76.3222
R2629 GNDA.n1145 GNDA.n1144 76.3222
R2630 GNDA.n1140 GNDA.n1139 76.3222
R2631 GNDA.n1137 GNDA.n1136 76.3222
R2632 GNDA.n1132 GNDA.n1131 76.3222
R2633 GNDA.n1129 GNDA.n1080 76.3222
R2634 GNDA.n2180 GNDA.n2179 76.3222
R2635 GNDA.n2175 GNDA.n1128 76.3222
R2636 GNDA.n2173 GNDA.n2172 76.3222
R2637 GNDA.n2168 GNDA.n2167 76.3222
R2638 GNDA.n2165 GNDA.n2164 76.3222
R2639 GNDA.n2160 GNDA.n2159 76.3222
R2640 GNDA.n608 GNDA.n604 76.3222
R2641 GNDA.n602 GNDA.n601 76.3222
R2642 GNDA.n597 GNDA.n596 76.3222
R2643 GNDA.n594 GNDA.n593 76.3222
R2644 GNDA.n589 GNDA.n588 76.3222
R2645 GNDA.n586 GNDA.n579 76.3222
R2646 GNDA.n2506 GNDA.n2505 76.3222
R2647 GNDA.n2501 GNDA.n585 76.3222
R2648 GNDA.n2499 GNDA.n2498 76.3222
R2649 GNDA.n2494 GNDA.n2493 76.3222
R2650 GNDA.n2491 GNDA.n2490 76.3222
R2651 GNDA.n606 GNDA.n605 76.3222
R2652 GNDA.n744 GNDA.n743 76.3222
R2653 GNDA.n741 GNDA.n740 76.3222
R2654 GNDA.n736 GNDA.n735 76.3222
R2655 GNDA.n733 GNDA.n732 76.3222
R2656 GNDA.n728 GNDA.n727 76.3222
R2657 GNDA.n725 GNDA.n721 76.3222
R2658 GNDA.n1044 GNDA.n1043 76.3222
R2659 GNDA.n1039 GNDA.n724 76.3222
R2660 GNDA.n1037 GNDA.n1036 76.3222
R2661 GNDA.n1032 GNDA.n1031 76.3222
R2662 GNDA.n1029 GNDA.n1028 76.3222
R2663 GNDA.n1024 GNDA.n1023 76.3222
R2664 GNDA.n2512 GNDA.n578 76.3222
R2665 GNDA.n2279 GNDA.n577 76.3222
R2666 GNDA.n2283 GNDA.n576 76.3222
R2667 GNDA.n2287 GNDA.n575 76.3222
R2668 GNDA.n2291 GNDA.n574 76.3222
R2669 GNDA.n2275 GNDA.n573 76.3222
R2670 GNDA.n717 GNDA.n572 76.3222
R2671 GNDA.n713 GNDA.n571 76.3222
R2672 GNDA.n709 GNDA.n570 76.3222
R2673 GNDA.n705 GNDA.n569 76.3222
R2674 GNDA.n701 GNDA.n568 76.3222
R2675 GNDA.n584 GNDA.n567 76.3222
R2676 GNDA.n779 GNDA.n566 76.3222
R2677 GNDA.n775 GNDA.n565 76.3222
R2678 GNDA.n771 GNDA.n564 76.3222
R2679 GNDA.n767 GNDA.n563 76.3222
R2680 GNDA.n763 GNDA.n562 76.3222
R2681 GNDA.n723 GNDA.n561 76.3222
R2682 GNDA.n2264 GNDA.n630 76.3222
R2683 GNDA.n673 GNDA.n634 76.3222
R2684 GNDA.n694 GNDA.n672 76.3222
R2685 GNDA.n683 GNDA.n671 76.3222
R2686 GNDA.n670 GNDA.n656 76.3222
R2687 GNDA.n2200 GNDA.n657 76.3222
R2688 GNDA.n2153 GNDA.n669 76.3222
R2689 GNDA.n2068 GNDA.n668 76.3222
R2690 GNDA.n2074 GNDA.n667 76.3222
R2691 GNDA.n2082 GNDA.n666 76.3222
R2692 GNDA.n2089 GNDA.n665 76.3222
R2693 GNDA.n2063 GNDA.n664 76.3222
R2694 GNDA.n2058 GNDA.n663 76.3222
R2695 GNDA.n1973 GNDA.n662 76.3222
R2696 GNDA.n1979 GNDA.n661 76.3222
R2697 GNDA.n1987 GNDA.n660 76.3222
R2698 GNDA.n1994 GNDA.n659 76.3222
R2699 GNDA.n1968 GNDA.n658 76.3222
R2700 GNDA.t272 GNDA.n69 75.0005
R2701 GNDA.n70 GNDA.t272 75.0005
R2702 GNDA.n485 GNDA.t247 75.0005
R2703 GNDA.n480 GNDA.t247 75.0005
R2704 GNDA.n501 GNDA.t221 75.0005
R2705 GNDA.n21 GNDA.t221 75.0005
R2706 GNDA.n375 GNDA.t200 75.0005
R2707 GNDA.n239 GNDA.t200 75.0005
R2708 GNDA.n359 GNDA.t216 75.0005
R2709 GNDA.n354 GNDA.t216 75.0005
R2710 GNDA.t235 GNDA.n266 75.0005
R2711 GNDA.n267 GNDA.t235 75.0005
R2712 GNDA.t250 GNDA.n298 75.0005
R2713 GNDA.n299 GNDA.t250 75.0005
R2714 GNDA.t256 GNDA.n37 75.0005
R2715 GNDA.n38 GNDA.t256 75.0005
R2716 GNDA.n1607 GNDA.n1281 74.5978
R2717 GNDA.n1604 GNDA.n1281 74.5978
R2718 GNDA.n2408 GNDA.n2336 74.5978
R2719 GNDA.n2405 GNDA.n2336 74.5978
R2720 GNDA.n2224 GNDA.n643 74.5978
R2721 GNDA.n2221 GNDA.n643 74.5978
R2722 GNDA.n2113 GNDA.n1161 74.5978
R2723 GNDA.n2110 GNDA.n1161 74.5978
R2724 GNDA.n2018 GNDA.n1182 74.5978
R2725 GNDA.n2015 GNDA.n1182 74.5978
R2726 GNDA.n1367 GNDA.n1306 74.5978
R2727 GNDA.n1364 GNDA.n1306 74.5978
R2728 GNDA.n1697 GNDA.n1680 74.5978
R2729 GNDA.n1698 GNDA.n1697 74.5978
R2730 GNDA.n962 GNDA.n903 74.5978
R2731 GNDA.n959 GNDA.n903 74.5978
R2732 GNDA.n842 GNDA.n537 74.5978
R2733 GNDA.n839 GNDA.n537 74.5978
R2734 GNDA.n937 GNDA.t181 74.1404
R2735 GNDA.n894 GNDA.t177 70.0216
R2736 GNDA.n1649 GNDA.n1271 69.3109
R2737 GNDA.n1625 GNDA.n1271 69.3109
R2738 GNDA.n2455 GNDA.n2321 69.3109
R2739 GNDA.n2426 GNDA.n2321 69.3109
R2740 GNDA.n2258 GNDA.n636 69.3109
R2741 GNDA.n2258 GNDA.n2257 69.3109
R2742 GNDA.n2147 GNDA.n1154 69.3109
R2743 GNDA.n2147 GNDA.n2146 69.3109
R2744 GNDA.n2052 GNDA.n1175 69.3109
R2745 GNDA.n2052 GNDA.n2051 69.3109
R2746 GNDA.n1401 GNDA.n1299 69.3109
R2747 GNDA.n1401 GNDA.n1400 69.3109
R2748 GNDA.n1739 GNDA.n1738 69.3109
R2749 GNDA.n1738 GNDA.n1737 69.3109
R2750 GNDA.n1010 GNDA.n890 69.3109
R2751 GNDA.n981 GNDA.n890 69.3109
R2752 GNDA.n2547 GNDA.n2546 69.3109
R2753 GNDA.n2547 GNDA.n548 69.3109
R2754 GNDA.t236 GNDA.n1639 65.8183
R2755 GNDA.t236 GNDA.n1290 65.8183
R2756 GNDA.t236 GNDA.n1289 65.8183
R2757 GNDA.t236 GNDA.n1288 65.8183
R2758 GNDA.t236 GNDA.n1279 65.8183
R2759 GNDA.t236 GNDA.n1286 65.8183
R2760 GNDA.t236 GNDA.n1277 65.8183
R2761 GNDA.t236 GNDA.n1287 65.8183
R2762 GNDA.t236 GNDA.n1285 65.8183
R2763 GNDA.t236 GNDA.n1284 65.8183
R2764 GNDA.t236 GNDA.n1283 65.8183
R2765 GNDA.t236 GNDA.n1282 65.8183
R2766 GNDA.t236 GNDA.n1280 65.8183
R2767 GNDA.t236 GNDA.n1278 65.8183
R2768 GNDA.n1640 GNDA.t236 65.8183
R2769 GNDA.t236 GNDA.n1272 65.8183
R2770 GNDA.t241 GNDA.n2440 65.8183
R2771 GNDA.t241 GNDA.n2345 65.8183
R2772 GNDA.t241 GNDA.n2344 65.8183
R2773 GNDA.t241 GNDA.n2343 65.8183
R2774 GNDA.t241 GNDA.n2334 65.8183
R2775 GNDA.t241 GNDA.n2341 65.8183
R2776 GNDA.t241 GNDA.n2332 65.8183
R2777 GNDA.t241 GNDA.n2342 65.8183
R2778 GNDA.t241 GNDA.n2340 65.8183
R2779 GNDA.t241 GNDA.n2339 65.8183
R2780 GNDA.t241 GNDA.n2338 65.8183
R2781 GNDA.t241 GNDA.n2337 65.8183
R2782 GNDA.t241 GNDA.n2335 65.8183
R2783 GNDA.t241 GNDA.n2333 65.8183
R2784 GNDA.n2443 GNDA.t241 65.8183
R2785 GNDA.t241 GNDA.n2322 65.8183
R2786 GNDA.t240 GNDA.n653 65.8183
R2787 GNDA.t240 GNDA.n652 65.8183
R2788 GNDA.t240 GNDA.n651 65.8183
R2789 GNDA.t240 GNDA.n650 65.8183
R2790 GNDA.t240 GNDA.n641 65.8183
R2791 GNDA.t240 GNDA.n648 65.8183
R2792 GNDA.t240 GNDA.n638 65.8183
R2793 GNDA.t240 GNDA.n649 65.8183
R2794 GNDA.t240 GNDA.n647 65.8183
R2795 GNDA.t240 GNDA.n646 65.8183
R2796 GNDA.t240 GNDA.n645 65.8183
R2797 GNDA.t240 GNDA.n644 65.8183
R2798 GNDA.t240 GNDA.n642 65.8183
R2799 GNDA.t240 GNDA.n640 65.8183
R2800 GNDA.t240 GNDA.n639 65.8183
R2801 GNDA.n2259 GNDA.t240 65.8183
R2802 GNDA.t232 GNDA.n1171 65.8183
R2803 GNDA.t232 GNDA.n1170 65.8183
R2804 GNDA.t232 GNDA.n1169 65.8183
R2805 GNDA.t232 GNDA.n1168 65.8183
R2806 GNDA.t232 GNDA.n1159 65.8183
R2807 GNDA.t232 GNDA.n1166 65.8183
R2808 GNDA.t232 GNDA.n1156 65.8183
R2809 GNDA.t232 GNDA.n1167 65.8183
R2810 GNDA.t232 GNDA.n1165 65.8183
R2811 GNDA.t232 GNDA.n1164 65.8183
R2812 GNDA.t232 GNDA.n1163 65.8183
R2813 GNDA.t232 GNDA.n1162 65.8183
R2814 GNDA.t232 GNDA.n1160 65.8183
R2815 GNDA.t232 GNDA.n1158 65.8183
R2816 GNDA.t232 GNDA.n1157 65.8183
R2817 GNDA.n2148 GNDA.t232 65.8183
R2818 GNDA.t261 GNDA.n1192 65.8183
R2819 GNDA.t261 GNDA.n1191 65.8183
R2820 GNDA.t261 GNDA.n1190 65.8183
R2821 GNDA.t261 GNDA.n1189 65.8183
R2822 GNDA.t261 GNDA.n1180 65.8183
R2823 GNDA.t261 GNDA.n1187 65.8183
R2824 GNDA.t261 GNDA.n1177 65.8183
R2825 GNDA.t261 GNDA.n1188 65.8183
R2826 GNDA.t261 GNDA.n1186 65.8183
R2827 GNDA.t261 GNDA.n1185 65.8183
R2828 GNDA.t261 GNDA.n1184 65.8183
R2829 GNDA.t261 GNDA.n1183 65.8183
R2830 GNDA.t261 GNDA.n1181 65.8183
R2831 GNDA.t261 GNDA.n1179 65.8183
R2832 GNDA.t261 GNDA.n1178 65.8183
R2833 GNDA.n2053 GNDA.t261 65.8183
R2834 GNDA.t210 GNDA.n1316 65.8183
R2835 GNDA.t210 GNDA.n1315 65.8183
R2836 GNDA.t210 GNDA.n1314 65.8183
R2837 GNDA.t210 GNDA.n1313 65.8183
R2838 GNDA.t210 GNDA.n1304 65.8183
R2839 GNDA.t210 GNDA.n1311 65.8183
R2840 GNDA.t210 GNDA.n1301 65.8183
R2841 GNDA.t210 GNDA.n1312 65.8183
R2842 GNDA.t210 GNDA.n1310 65.8183
R2843 GNDA.t210 GNDA.n1309 65.8183
R2844 GNDA.t210 GNDA.n1308 65.8183
R2845 GNDA.t210 GNDA.n1307 65.8183
R2846 GNDA.n1719 GNDA.t226 65.8183
R2847 GNDA.n1721 GNDA.t226 65.8183
R2848 GNDA.n1727 GNDA.t226 65.8183
R2849 GNDA.n1729 GNDA.t226 65.8183
R2850 GNDA.n1703 GNDA.t226 65.8183
R2851 GNDA.n1705 GNDA.t226 65.8183
R2852 GNDA.n1711 GNDA.t226 65.8183
R2853 GNDA.n1713 GNDA.t226 65.8183
R2854 GNDA.t226 GNDA.n1660 65.8183
R2855 GNDA.n1688 GNDA.t226 65.8183
R2856 GNDA.n1684 GNDA.t226 65.8183
R2857 GNDA.n1695 GNDA.t226 65.8183
R2858 GNDA.n1768 GNDA.t226 65.8183
R2859 GNDA.n1755 GNDA.t226 65.8183
R2860 GNDA.n1753 GNDA.t226 65.8183
R2861 GNDA.n1740 GNDA.t226 65.8183
R2862 GNDA.t210 GNDA.n1305 65.8183
R2863 GNDA.t210 GNDA.n1303 65.8183
R2864 GNDA.t210 GNDA.n1302 65.8183
R2865 GNDA.n1402 GNDA.t210 65.8183
R2866 GNDA.t230 GNDA.n995 65.8183
R2867 GNDA.t230 GNDA.n912 65.8183
R2868 GNDA.t230 GNDA.n911 65.8183
R2869 GNDA.t230 GNDA.n910 65.8183
R2870 GNDA.t230 GNDA.n901 65.8183
R2871 GNDA.t230 GNDA.n908 65.8183
R2872 GNDA.t230 GNDA.n899 65.8183
R2873 GNDA.t230 GNDA.n909 65.8183
R2874 GNDA.t230 GNDA.n907 65.8183
R2875 GNDA.t230 GNDA.n906 65.8183
R2876 GNDA.t230 GNDA.n905 65.8183
R2877 GNDA.t230 GNDA.n904 65.8183
R2878 GNDA.t230 GNDA.n902 65.8183
R2879 GNDA.t230 GNDA.n900 65.8183
R2880 GNDA.n998 GNDA.t230 65.8183
R2881 GNDA.t230 GNDA.n891 65.8183
R2882 GNDA.t260 GNDA.n547 65.8183
R2883 GNDA.t260 GNDA.n546 65.8183
R2884 GNDA.t260 GNDA.n545 65.8183
R2885 GNDA.t260 GNDA.n544 65.8183
R2886 GNDA.t260 GNDA.n535 65.8183
R2887 GNDA.t260 GNDA.n542 65.8183
R2888 GNDA.t260 GNDA.n533 65.8183
R2889 GNDA.t260 GNDA.n543 65.8183
R2890 GNDA.t260 GNDA.n541 65.8183
R2891 GNDA.t260 GNDA.n540 65.8183
R2892 GNDA.t260 GNDA.n539 65.8183
R2893 GNDA.t260 GNDA.n538 65.8183
R2894 GNDA.t260 GNDA.n536 65.8183
R2895 GNDA.n2548 GNDA.t260 65.8183
R2896 GNDA.t260 GNDA.n534 65.8183
R2897 GNDA.t260 GNDA.n532 65.8183
R2898 GNDA.t3 GNDA.t26 65.7614
R2899 GNDA.t301 GNDA.t3 65.7614
R2900 GNDA.t303 GNDA.t15 65.7614
R2901 GNDA.t137 GNDA.t90 65.271
R2902 GNDA.t96 GNDA.t304 65.271
R2903 GNDA.n404 GNDA.t14 65.271
R2904 GNDA.t313 GNDA.t307 65.271
R2905 GNDA.t293 GNDA.t317 65.271
R2906 GNDA.n1966 GNDA.t211 65.0078
R2907 GNDA.t169 GNDA.n2327 63.8432
R2908 GNDA.n1005 GNDA.t191 63.8432
R2909 GNDA.n2540 GNDA.t171 63.8432
R2910 GNDA.t296 GNDA.t130 62.9326
R2911 GNDA.t316 GNDA.t86 62.9326
R2912 GNDA.t39 GNDA.t316 62.9326
R2913 GNDA.t319 GNDA.t39 62.9326
R2914 GNDA.n362 GNDA.n8 61.4316
R2915 GNDA.n2370 GNDA.t173 59.7243
R2916 GNDA.n936 GNDA.t193 59.7243
R2917 GNDA.n817 GNDA.t185 59.7243
R2918 GNDA.n2461 GNDA.t83 58.6946
R2919 GNDA.n2449 GNDA.t126 58.6946
R2920 GNDA.t310 GNDA.n2381 58.6946
R2921 GNDA.t236 GNDA.n1271 57.8461
R2922 GNDA.t241 GNDA.n2321 57.8461
R2923 GNDA.t240 GNDA.n2258 57.8461
R2924 GNDA.t232 GNDA.n2147 57.8461
R2925 GNDA.t261 GNDA.n2052 57.8461
R2926 GNDA.n1738 GNDA.t226 57.8461
R2927 GNDA.t210 GNDA.n1401 57.8461
R2928 GNDA.t230 GNDA.n890 57.8461
R2929 GNDA.t260 GNDA.n2547 57.8461
R2930 GNDA.t220 GNDA.n17 57.5921
R2931 GNDA.n120 GNDA.t246 57.5921
R2932 GNDA.t63 GNDA.n127 57.5921
R2933 GNDA.n137 GNDA.t22 57.5921
R2934 GNDA.t199 GNDA.n235 57.5921
R2935 GNDA.n349 GNDA.t215 57.5921
R2936 GNDA.n186 GNDA.n13 57.3163
R2937 GNDA.n2584 GNDA.n2583 57.3163
R2938 GNDA.t306 GNDA.n2585 56.7945
R2939 GNDA.t99 GNDA.t159 56.6352
R2940 GNDA.n1015 GNDA.t287 56.6352
R2941 GNDA.t1 GNDA.t155 56.6352
R2942 GNDA.n753 GNDA.n750 56.3995
R2943 GNDA.n1266 GNDA.n622 56.3995
R2944 GNDA.n2317 GNDA.n2316 56.3995
R2945 GNDA.n2316 GNDA.n611 56.3995
R2946 GNDA.n1265 GNDA.n622 56.3995
R2947 GNDA.n2269 GNDA.n629 56.3995
R2948 GNDA.n1964 GNDA.n1194 56.3995
R2949 GNDA.n1781 GNDA.n1780 56.3995
R2950 GNDA.n750 GNDA.n749 56.3995
R2951 GNDA.n1967 GNDA.n1194 56.3995
R2952 GNDA.n1781 GNDA.n1777 56.3995
R2953 GNDA.n2484 GNDA.n2483 55.6055
R2954 GNDA.t236 GNDA.n1281 55.2026
R2955 GNDA.t241 GNDA.n2336 55.2026
R2956 GNDA.t240 GNDA.n643 55.2026
R2957 GNDA.t232 GNDA.n1161 55.2026
R2958 GNDA.t261 GNDA.n1182 55.2026
R2959 GNDA.t210 GNDA.n1306 55.2026
R2960 GNDA.n1697 GNDA.t226 55.2026
R2961 GNDA.t230 GNDA.n903 55.2026
R2962 GNDA.t260 GNDA.n537 55.2026
R2963 GNDA.n1018 GNDA.n1017 54.5757
R2964 GNDA.n2525 GNDA.n553 54.5757
R2965 GNDA.t295 GNDA.n2541 54.5757
R2966 GNDA.n810 GNDA.t292 54.5757
R2967 GNDA.t36 GNDA.n513 54.5757
R2968 GNDA.t49 GNDA.t80 53.7527
R2969 GNDA.t179 GNDA.n936 53.546
R2970 GNDA.n1622 GNDA.n1287 53.3664
R2971 GNDA.n1619 GNDA.n1277 53.3664
R2972 GNDA.n1615 GNDA.n1286 53.3664
R2973 GNDA.n1611 GNDA.n1279 53.3664
R2974 GNDA.n1600 GNDA.n1282 53.3664
R2975 GNDA.n1596 GNDA.n1283 53.3664
R2976 GNDA.n1592 GNDA.n1284 53.3664
R2977 GNDA.n1588 GNDA.n1285 53.3664
R2978 GNDA.n1648 GNDA.n1272 53.3664
R2979 GNDA.n1641 GNDA.n1640 53.3664
R2980 GNDA.n1573 GNDA.n1278 53.3664
R2981 GNDA.n1580 GNDA.n1280 53.3664
R2982 GNDA.n1639 GNDA.n1638 53.3664
R2983 GNDA.n1292 GNDA.n1290 53.3664
R2984 GNDA.n1633 GNDA.n1289 53.3664
R2985 GNDA.n1629 GNDA.n1288 53.3664
R2986 GNDA.n1639 GNDA.n1291 53.3664
R2987 GNDA.n1634 GNDA.n1290 53.3664
R2988 GNDA.n1630 GNDA.n1289 53.3664
R2989 GNDA.n1626 GNDA.n1288 53.3664
R2990 GNDA.n1608 GNDA.n1279 53.3664
R2991 GNDA.n1612 GNDA.n1286 53.3664
R2992 GNDA.n1616 GNDA.n1277 53.3664
R2993 GNDA.n1620 GNDA.n1287 53.3664
R2994 GNDA.n1591 GNDA.n1285 53.3664
R2995 GNDA.n1595 GNDA.n1284 53.3664
R2996 GNDA.n1599 GNDA.n1283 53.3664
R2997 GNDA.n1603 GNDA.n1282 53.3664
R2998 GNDA.n1587 GNDA.n1280 53.3664
R2999 GNDA.n1579 GNDA.n1278 53.3664
R3000 GNDA.n1640 GNDA.n1276 53.3664
R3001 GNDA.n1275 GNDA.n1272 53.3664
R3002 GNDA.n2423 GNDA.n2342 53.3664
R3003 GNDA.n2420 GNDA.n2332 53.3664
R3004 GNDA.n2416 GNDA.n2341 53.3664
R3005 GNDA.n2412 GNDA.n2334 53.3664
R3006 GNDA.n2401 GNDA.n2337 53.3664
R3007 GNDA.n2397 GNDA.n2338 53.3664
R3008 GNDA.n2393 GNDA.n2339 53.3664
R3009 GNDA.n2389 GNDA.n2340 53.3664
R3010 GNDA.n2454 GNDA.n2322 53.3664
R3011 GNDA.n2443 GNDA.n2442 53.3664
R3012 GNDA.n2333 GNDA.n2331 53.3664
R3013 GNDA.n2377 GNDA.n2335 53.3664
R3014 GNDA.n2440 GNDA.n2439 53.3664
R3015 GNDA.n2347 GNDA.n2345 53.3664
R3016 GNDA.n2434 GNDA.n2344 53.3664
R3017 GNDA.n2430 GNDA.n2343 53.3664
R3018 GNDA.n2440 GNDA.n2346 53.3664
R3019 GNDA.n2435 GNDA.n2345 53.3664
R3020 GNDA.n2431 GNDA.n2344 53.3664
R3021 GNDA.n2427 GNDA.n2343 53.3664
R3022 GNDA.n2409 GNDA.n2334 53.3664
R3023 GNDA.n2413 GNDA.n2341 53.3664
R3024 GNDA.n2417 GNDA.n2332 53.3664
R3025 GNDA.n2421 GNDA.n2342 53.3664
R3026 GNDA.n2392 GNDA.n2340 53.3664
R3027 GNDA.n2396 GNDA.n2339 53.3664
R3028 GNDA.n2400 GNDA.n2338 53.3664
R3029 GNDA.n2404 GNDA.n2337 53.3664
R3030 GNDA.n2388 GNDA.n2335 53.3664
R3031 GNDA.n2376 GNDA.n2333 53.3664
R3032 GNDA.n2444 GNDA.n2443 53.3664
R3033 GNDA.n2441 GNDA.n2322 53.3664
R3034 GNDA.n2240 GNDA.n649 53.3664
R3035 GNDA.n2236 GNDA.n638 53.3664
R3036 GNDA.n2232 GNDA.n648 53.3664
R3037 GNDA.n2228 GNDA.n641 53.3664
R3038 GNDA.n2217 GNDA.n644 53.3664
R3039 GNDA.n2213 GNDA.n645 53.3664
R3040 GNDA.n2209 GNDA.n646 53.3664
R3041 GNDA.n2205 GNDA.n647 53.3664
R3042 GNDA.n2260 GNDA.n2259 53.3664
R3043 GNDA.n690 GNDA.n639 53.3664
R3044 GNDA.n686 GNDA.n640 53.3664
R3045 GNDA.n679 GNDA.n642 53.3664
R3046 GNDA.n2244 GNDA.n653 53.3664
R3047 GNDA.n2245 GNDA.n652 53.3664
R3048 GNDA.n2249 GNDA.n651 53.3664
R3049 GNDA.n2253 GNDA.n650 53.3664
R3050 GNDA.n2241 GNDA.n653 53.3664
R3051 GNDA.n2248 GNDA.n652 53.3664
R3052 GNDA.n2252 GNDA.n651 53.3664
R3053 GNDA.n2256 GNDA.n650 53.3664
R3054 GNDA.n2225 GNDA.n641 53.3664
R3055 GNDA.n2229 GNDA.n648 53.3664
R3056 GNDA.n2233 GNDA.n638 53.3664
R3057 GNDA.n2237 GNDA.n649 53.3664
R3058 GNDA.n2208 GNDA.n647 53.3664
R3059 GNDA.n2212 GNDA.n646 53.3664
R3060 GNDA.n2216 GNDA.n645 53.3664
R3061 GNDA.n2220 GNDA.n644 53.3664
R3062 GNDA.n2204 GNDA.n642 53.3664
R3063 GNDA.n678 GNDA.n640 53.3664
R3064 GNDA.n687 GNDA.n639 53.3664
R3065 GNDA.n2259 GNDA.n637 53.3664
R3066 GNDA.n2129 GNDA.n1167 53.3664
R3067 GNDA.n2125 GNDA.n1156 53.3664
R3068 GNDA.n2121 GNDA.n1166 53.3664
R3069 GNDA.n2117 GNDA.n1159 53.3664
R3070 GNDA.n2106 GNDA.n1162 53.3664
R3071 GNDA.n2102 GNDA.n1163 53.3664
R3072 GNDA.n2098 GNDA.n1164 53.3664
R3073 GNDA.n2094 GNDA.n1165 53.3664
R3074 GNDA.n2149 GNDA.n2148 53.3664
R3075 GNDA.n2071 GNDA.n1157 53.3664
R3076 GNDA.n2079 GNDA.n1158 53.3664
R3077 GNDA.n2086 GNDA.n1160 53.3664
R3078 GNDA.n2133 GNDA.n1171 53.3664
R3079 GNDA.n2134 GNDA.n1170 53.3664
R3080 GNDA.n2138 GNDA.n1169 53.3664
R3081 GNDA.n2142 GNDA.n1168 53.3664
R3082 GNDA.n2130 GNDA.n1171 53.3664
R3083 GNDA.n2137 GNDA.n1170 53.3664
R3084 GNDA.n2141 GNDA.n1169 53.3664
R3085 GNDA.n2145 GNDA.n1168 53.3664
R3086 GNDA.n2114 GNDA.n1159 53.3664
R3087 GNDA.n2118 GNDA.n1166 53.3664
R3088 GNDA.n2122 GNDA.n1156 53.3664
R3089 GNDA.n2126 GNDA.n1167 53.3664
R3090 GNDA.n2097 GNDA.n1165 53.3664
R3091 GNDA.n2101 GNDA.n1164 53.3664
R3092 GNDA.n2105 GNDA.n1163 53.3664
R3093 GNDA.n2109 GNDA.n1162 53.3664
R3094 GNDA.n2093 GNDA.n1160 53.3664
R3095 GNDA.n2085 GNDA.n1158 53.3664
R3096 GNDA.n2078 GNDA.n1157 53.3664
R3097 GNDA.n2148 GNDA.n1155 53.3664
R3098 GNDA.n2034 GNDA.n1188 53.3664
R3099 GNDA.n2030 GNDA.n1177 53.3664
R3100 GNDA.n2026 GNDA.n1187 53.3664
R3101 GNDA.n2022 GNDA.n1180 53.3664
R3102 GNDA.n2011 GNDA.n1183 53.3664
R3103 GNDA.n2007 GNDA.n1184 53.3664
R3104 GNDA.n2003 GNDA.n1185 53.3664
R3105 GNDA.n1999 GNDA.n1186 53.3664
R3106 GNDA.n2054 GNDA.n2053 53.3664
R3107 GNDA.n1976 GNDA.n1178 53.3664
R3108 GNDA.n1984 GNDA.n1179 53.3664
R3109 GNDA.n1991 GNDA.n1181 53.3664
R3110 GNDA.n2038 GNDA.n1192 53.3664
R3111 GNDA.n2039 GNDA.n1191 53.3664
R3112 GNDA.n2043 GNDA.n1190 53.3664
R3113 GNDA.n2047 GNDA.n1189 53.3664
R3114 GNDA.n2035 GNDA.n1192 53.3664
R3115 GNDA.n2042 GNDA.n1191 53.3664
R3116 GNDA.n2046 GNDA.n1190 53.3664
R3117 GNDA.n2050 GNDA.n1189 53.3664
R3118 GNDA.n2019 GNDA.n1180 53.3664
R3119 GNDA.n2023 GNDA.n1187 53.3664
R3120 GNDA.n2027 GNDA.n1177 53.3664
R3121 GNDA.n2031 GNDA.n1188 53.3664
R3122 GNDA.n2002 GNDA.n1186 53.3664
R3123 GNDA.n2006 GNDA.n1185 53.3664
R3124 GNDA.n2010 GNDA.n1184 53.3664
R3125 GNDA.n2014 GNDA.n1183 53.3664
R3126 GNDA.n1998 GNDA.n1181 53.3664
R3127 GNDA.n1990 GNDA.n1179 53.3664
R3128 GNDA.n1983 GNDA.n1178 53.3664
R3129 GNDA.n2053 GNDA.n1176 53.3664
R3130 GNDA.n1383 GNDA.n1312 53.3664
R3131 GNDA.n1379 GNDA.n1301 53.3664
R3132 GNDA.n1375 GNDA.n1311 53.3664
R3133 GNDA.n1371 GNDA.n1304 53.3664
R3134 GNDA.n1360 GNDA.n1307 53.3664
R3135 GNDA.n1356 GNDA.n1308 53.3664
R3136 GNDA.n1352 GNDA.n1309 53.3664
R3137 GNDA.n1348 GNDA.n1310 53.3664
R3138 GNDA.n1403 GNDA.n1402 53.3664
R3139 GNDA.n1325 GNDA.n1302 53.3664
R3140 GNDA.n1333 GNDA.n1303 53.3664
R3141 GNDA.n1340 GNDA.n1305 53.3664
R3142 GNDA.n1387 GNDA.n1316 53.3664
R3143 GNDA.n1388 GNDA.n1315 53.3664
R3144 GNDA.n1392 GNDA.n1314 53.3664
R3145 GNDA.n1396 GNDA.n1313 53.3664
R3146 GNDA.n1384 GNDA.n1316 53.3664
R3147 GNDA.n1391 GNDA.n1315 53.3664
R3148 GNDA.n1395 GNDA.n1314 53.3664
R3149 GNDA.n1399 GNDA.n1313 53.3664
R3150 GNDA.n1368 GNDA.n1304 53.3664
R3151 GNDA.n1372 GNDA.n1311 53.3664
R3152 GNDA.n1376 GNDA.n1301 53.3664
R3153 GNDA.n1380 GNDA.n1312 53.3664
R3154 GNDA.n1351 GNDA.n1310 53.3664
R3155 GNDA.n1355 GNDA.n1309 53.3664
R3156 GNDA.n1359 GNDA.n1308 53.3664
R3157 GNDA.n1363 GNDA.n1307 53.3664
R3158 GNDA.n1713 GNDA.n1676 53.3664
R3159 GNDA.n1712 GNDA.n1711 53.3664
R3160 GNDA.n1705 GNDA.n1678 53.3664
R3161 GNDA.n1704 GNDA.n1703 53.3664
R3162 GNDA.n1695 GNDA.n1694 53.3664
R3163 GNDA.n1690 GNDA.n1684 53.3664
R3164 GNDA.n1688 GNDA.n1687 53.3664
R3165 GNDA.n1770 GNDA.n1660 53.3664
R3166 GNDA.n1741 GNDA.n1740 53.3664
R3167 GNDA.n1753 GNDA.n1752 53.3664
R3168 GNDA.n1756 GNDA.n1755 53.3664
R3169 GNDA.n1768 GNDA.n1767 53.3664
R3170 GNDA.n1720 GNDA.n1719 53.3664
R3171 GNDA.n1722 GNDA.n1721 53.3664
R3172 GNDA.n1727 GNDA.n1726 53.3664
R3173 GNDA.n1730 GNDA.n1729 53.3664
R3174 GNDA.n1719 GNDA.n1718 53.3664
R3175 GNDA.n1721 GNDA.n1674 53.3664
R3176 GNDA.n1728 GNDA.n1727 53.3664
R3177 GNDA.n1729 GNDA.n1672 53.3664
R3178 GNDA.n1703 GNDA.n1702 53.3664
R3179 GNDA.n1706 GNDA.n1705 53.3664
R3180 GNDA.n1711 GNDA.n1710 53.3664
R3181 GNDA.n1714 GNDA.n1713 53.3664
R3182 GNDA.n1685 GNDA.n1660 53.3664
R3183 GNDA.n1689 GNDA.n1688 53.3664
R3184 GNDA.n1684 GNDA.n1682 53.3664
R3185 GNDA.n1696 GNDA.n1695 53.3664
R3186 GNDA.n1769 GNDA.n1768 53.3664
R3187 GNDA.n1755 GNDA.n1661 53.3664
R3188 GNDA.n1754 GNDA.n1753 53.3664
R3189 GNDA.n1740 GNDA.n1666 53.3664
R3190 GNDA.n1347 GNDA.n1305 53.3664
R3191 GNDA.n1339 GNDA.n1303 53.3664
R3192 GNDA.n1332 GNDA.n1302 53.3664
R3193 GNDA.n1402 GNDA.n1300 53.3664
R3194 GNDA.n977 GNDA.n909 53.3664
R3195 GNDA.n974 GNDA.n899 53.3664
R3196 GNDA.n970 GNDA.n908 53.3664
R3197 GNDA.n966 GNDA.n901 53.3664
R3198 GNDA.n955 GNDA.n904 53.3664
R3199 GNDA.n951 GNDA.n905 53.3664
R3200 GNDA.n947 GNDA.n906 53.3664
R3201 GNDA.n943 GNDA.n907 53.3664
R3202 GNDA.n1009 GNDA.n891 53.3664
R3203 GNDA.n998 GNDA.n997 53.3664
R3204 GNDA.n900 GNDA.n898 53.3664
R3205 GNDA.n930 GNDA.n902 53.3664
R3206 GNDA.n995 GNDA.n994 53.3664
R3207 GNDA.n914 GNDA.n912 53.3664
R3208 GNDA.n989 GNDA.n911 53.3664
R3209 GNDA.n985 GNDA.n910 53.3664
R3210 GNDA.n995 GNDA.n913 53.3664
R3211 GNDA.n990 GNDA.n912 53.3664
R3212 GNDA.n986 GNDA.n911 53.3664
R3213 GNDA.n982 GNDA.n910 53.3664
R3214 GNDA.n963 GNDA.n901 53.3664
R3215 GNDA.n967 GNDA.n908 53.3664
R3216 GNDA.n971 GNDA.n899 53.3664
R3217 GNDA.n975 GNDA.n909 53.3664
R3218 GNDA.n946 GNDA.n907 53.3664
R3219 GNDA.n950 GNDA.n906 53.3664
R3220 GNDA.n954 GNDA.n905 53.3664
R3221 GNDA.n958 GNDA.n904 53.3664
R3222 GNDA.n942 GNDA.n902 53.3664
R3223 GNDA.n931 GNDA.n900 53.3664
R3224 GNDA.n999 GNDA.n998 53.3664
R3225 GNDA.n996 GNDA.n891 53.3664
R3226 GNDA.n858 GNDA.n543 53.3664
R3227 GNDA.n854 GNDA.n533 53.3664
R3228 GNDA.n850 GNDA.n542 53.3664
R3229 GNDA.n846 GNDA.n535 53.3664
R3230 GNDA.n835 GNDA.n538 53.3664
R3231 GNDA.n831 GNDA.n539 53.3664
R3232 GNDA.n827 GNDA.n540 53.3664
R3233 GNDA.n823 GNDA.n541 53.3664
R3234 GNDA.n549 GNDA.n532 53.3664
R3235 GNDA.n2536 GNDA.n534 53.3664
R3236 GNDA.n2549 GNDA.n2548 53.3664
R3237 GNDA.n812 GNDA.n536 53.3664
R3238 GNDA.n862 GNDA.n547 53.3664
R3239 GNDA.n863 GNDA.n546 53.3664
R3240 GNDA.n867 GNDA.n545 53.3664
R3241 GNDA.n871 GNDA.n544 53.3664
R3242 GNDA.n859 GNDA.n547 53.3664
R3243 GNDA.n866 GNDA.n546 53.3664
R3244 GNDA.n870 GNDA.n545 53.3664
R3245 GNDA.n873 GNDA.n544 53.3664
R3246 GNDA.n843 GNDA.n535 53.3664
R3247 GNDA.n847 GNDA.n542 53.3664
R3248 GNDA.n851 GNDA.n533 53.3664
R3249 GNDA.n855 GNDA.n543 53.3664
R3250 GNDA.n826 GNDA.n541 53.3664
R3251 GNDA.n830 GNDA.n540 53.3664
R3252 GNDA.n834 GNDA.n539 53.3664
R3253 GNDA.n838 GNDA.n538 53.3664
R3254 GNDA.n822 GNDA.n536 53.3664
R3255 GNDA.n2548 GNDA.n531 53.3664
R3256 GNDA.n534 GNDA.n530 53.3664
R3257 GNDA.n2535 GNDA.n532 53.3664
R3258 GNDA.n1803 GNDA.n1802 52.7091
R3259 GNDA.n1802 GNDA.n1241 52.7091
R3260 GNDA.n1796 GNDA.n1241 52.7091
R3261 GNDA.n1796 GNDA.n1795 52.7091
R3262 GNDA.n1795 GNDA.n1794 52.7091
R3263 GNDA.n1788 GNDA.n1248 52.7091
R3264 GNDA.n1788 GNDA.n1787 52.7091
R3265 GNDA.n1787 GNDA.n1786 52.7091
R3266 GNDA.n1786 GNDA.n1249 52.7091
R3267 GNDA.n1779 GNDA.n1249 52.7091
R3268 GNDA.n1779 GNDA.n1778 52.7091
R3269 GNDA.n1778 GNDA.t46 52.7091
R3270 GNDA.n1940 GNDA.n1202 52.7091
R3271 GNDA.n1946 GNDA.n1202 52.7091
R3272 GNDA.n1947 GNDA.n1946 52.7091
R3273 GNDA.n1949 GNDA.n1947 52.7091
R3274 GNDA.n1949 GNDA.n1948 52.7091
R3275 GNDA.n1956 GNDA.n1955 52.7091
R3276 GNDA.n1958 GNDA.n1956 52.7091
R3277 GNDA.n1958 GNDA.n1957 52.7091
R3278 GNDA.n1957 GNDA.n1195 52.7091
R3279 GNDA.n1965 GNDA.n1195 52.7091
R3280 GNDA.n1966 GNDA.n1965 52.7091
R3281 GNDA.n783 GNDA.n759 52.7091
R3282 GNDA.n790 GNDA.n759 52.7091
R3283 GNDA.n791 GNDA.n790 52.7091
R3284 GNDA.n792 GNDA.n791 52.7091
R3285 GNDA.n792 GNDA.n525 52.7091
R3286 GNDA.n754 GNDA.n526 52.7091
R3287 GNDA.n800 GNDA.n754 52.7091
R3288 GNDA.n801 GNDA.n800 52.7091
R3289 GNDA.n804 GNDA.n801 52.7091
R3290 GNDA.n804 GNDA.n803 52.7091
R3291 GNDA.n803 GNDA.n802 52.7091
R3292 GNDA.t211 GNDA.n558 51.4866
R3293 GNDA.n2514 GNDA.t211 51.4866
R3294 GNDA.t325 GNDA.t88 49.9132
R3295 GNDA.t97 GNDA.t100 49.9132
R3296 GNDA.t323 GNDA.t54 49.9132
R3297 GNDA.t28 GNDA.t135 49.9132
R3298 GNDA.n1005 GNDA.t165 49.4271
R3299 GNDA.t108 GNDA.n553 48.3974
R3300 GNDA.n2484 GNDA.t77 47.3677
R3301 GNDA.t105 GNDA.t258 46.338
R3302 GNDA.t252 GNDA.t48 46.338
R3303 GNDA.t211 GNDA.n1517 46.2335
R3304 GNDA.n1460 GNDA.t211 46.2335
R3305 GNDA.n1818 GNDA.t211 46.2335
R3306 GNDA.n504 GNDA.n17 46.0738
R3307 GNDA.n488 GNDA.n120 46.0738
R3308 GNDA.t208 GNDA.t63 46.0738
R3309 GNDA.t196 GNDA.t20 46.0738
R3310 GNDA.t79 GNDA.t274 46.0738
R3311 GNDA.n378 GNDA.n235 46.0738
R3312 GNDA.n362 GNDA.n349 46.0738
R3313 GNDA.n193 GNDA.t25 44.838
R3314 GNDA.t258 GNDA.n2326 43.2488
R3315 GNDA.t165 GNDA.n894 43.2488
R3316 GNDA.n2541 GNDA.t183 43.2488
R3317 GNDA.n1518 GNDA.t211 42.2987
R3318 GNDA.t211 GNDA.n1459 42.2987
R3319 GNDA.n1236 GNDA.t211 42.2987
R3320 GNDA.t153 GNDA.t55 42.2405
R3321 GNDA.t55 GNDA.t297 42.2405
R3322 GNDA.t299 GNDA.t84 42.2405
R3323 GNDA.t84 GNDA.t12 42.2405
R3324 GNDA.n455 GNDA.t57 42.2344
R3325 GNDA.n1003 GNDA.t35 42.2191
R3326 GNDA.t91 GNDA.n2589 41.8488
R3327 GNDA.t27 GNDA.n2588 41.8488
R3328 GNDA.t45 GNDA.n2587 41.8488
R3329 GNDA.t129 GNDA.n2586 41.8488
R3330 GNDA.t128 GNDA.n2590 41.8488
R3331 GNDA.t211 GNDA.t77 41.1894
R3332 GNDA.t211 GNDA.t108 41.1894
R3333 GNDA.n455 GNDA.t117 40.4913
R3334 GNDA.t11 GNDA.t319 39.8575
R3335 GNDA.n2366 GNDA.n519 39.3903
R3336 GNDA.n2381 GNDA.t161 39.1299
R3337 GNDA.n926 GNDA.n925 39.1299
R3338 GNDA.n937 GNDA.t179 39.1299
R3339 GNDA.n818 GNDA.t252 39.1299
R3340 GNDA.t294 GNDA.t123 38.3949
R3341 GNDA.n883 GNDA.n558 38.1002
R3342 GNDA.n1017 GNDA.n881 38.1002
R3343 GNDA.n2553 GNDA.t292 38.1002
R3344 GNDA.n818 GNDA.t36 38.1002
R3345 GNDA.n2514 GNDA.n556 37.0705
R3346 GNDA.t187 GNDA.t211 36.0408
R3347 GNDA.t211 GNDA.t167 36.0408
R3348 GNDA.t60 GNDA.n191 35.8706
R3349 GNDA.t4 GNDA.n190 35.8706
R3350 GNDA.t16 GNDA.n189 35.8706
R3351 GNDA.t0 GNDA.n188 35.8706
R3352 GNDA.n186 GNDA.t205 35.8706
R3353 GNDA.t25 GNDA.n192 35.8706
R3354 GNDA.t294 GNDA.n187 35.8706
R3355 GNDA.t15 GNDA.n2584 35.8706
R3356 GNDA.n1794 GNDA.t211 35.7252
R3357 GNDA.n1948 GNDA.t211 35.7252
R3358 GNDA.t211 GNDA.n525 35.7252
R3359 GNDA.n2567 GNDA.n2566 35.3278
R3360 GNDA.t41 GNDA.t325 34.5555
R3361 GNDA.t100 GNDA.t98 34.5555
R3362 GNDA.t59 GNDA.t19 34.5555
R3363 GNDA.n455 GNDA.t121 34.5555
R3364 GNDA.t154 GNDA.t323 34.5555
R3365 GNDA.t135 GNDA.t146 34.5555
R3366 GNDA.n2326 GNDA.t83 33.9813
R3367 GNDA.t126 GNDA.n2448 33.9813
R3368 GNDA.n1015 GNDA.n1014 33.9813
R3369 GNDA.t173 GNDA.n2369 32.9516
R3370 GNDA.t193 GNDA.n935 32.9516
R3371 GNDA.t185 GNDA.n816 32.9516
R3372 GNDA.n2198 GNDA.t211 32.9056
R3373 GNDA.n1252 GNDA.t211 32.9056
R3374 GNDA.n2571 GNDA.n2570 32.3063
R3375 GNDA.t10 GNDA.t127 30.716
R3376 GNDA.t119 GNDA.t196 30.716
R3377 GNDA.t79 GNDA.t109 30.716
R3378 GNDA.t65 GNDA.t49 30.716
R3379 GNDA.t26 GNDA.n186 29.8923
R3380 GNDA.n192 GNDA.t60 29.8923
R3381 GNDA.n187 GNDA.t208 29.8923
R3382 GNDA.n191 GNDA.t4 29.8923
R3383 GNDA.n190 GNDA.t16 29.8923
R3384 GNDA.n189 GNDA.t0 29.8923
R3385 GNDA.n188 GNDA.t59 29.8923
R3386 GNDA.n2584 GNDA.t202 29.8923
R3387 GNDA.n2602 GNDA.n0 29.8047
R3388 GNDA.t92 GNDA.n511 29.2831
R3389 GNDA.n2450 GNDA.t169 28.8327
R3390 GNDA.t191 GNDA.n1004 28.8327
R3391 GNDA.t171 GNDA.n2530 28.8327
R3392 GNDA.n2450 GNDA.t99 27.803
R3393 GNDA.n2370 GNDA.t145 27.803
R3394 GNDA.n2383 GNDA.t72 27.803
R3395 GNDA.n1624 GNDA.n1623 27.5561
R3396 GNDA.n2425 GNDA.n2424 27.5561
R3397 GNDA.n2242 GNDA.n2239 27.5561
R3398 GNDA.n2131 GNDA.n2128 27.5561
R3399 GNDA.n2036 GNDA.n2033 27.5561
R3400 GNDA.n1385 GNDA.n1382 27.5561
R3401 GNDA.n1717 GNDA.n1716 27.5561
R3402 GNDA.n979 GNDA.n978 27.5561
R3403 GNDA.n860 GNDA.n857 27.5561
R3404 GNDA.t102 GNDA.n127 26.8766
R3405 GNDA.n1606 GNDA.n1605 26.6672
R3406 GNDA.n2407 GNDA.n2406 26.6672
R3407 GNDA.n2223 GNDA.n2222 26.6672
R3408 GNDA.n2112 GNDA.n2111 26.6672
R3409 GNDA.n2017 GNDA.n2016 26.6672
R3410 GNDA.n1366 GNDA.n1365 26.6672
R3411 GNDA.n1700 GNDA.n1699 26.6672
R3412 GNDA.n961 GNDA.n960 26.6672
R3413 GNDA.n841 GNDA.n840 26.6672
R3414 GNDA.t145 GNDA.t161 25.7435
R3415 GNDA.t183 GNDA.t58 25.7435
R3416 GNDA.n2357 GNDA.n2356 25.3679
R3417 GNDA.n396 GNDA.n395 24.991
R3418 GNDA.n216 GNDA.n215 24.7472
R3419 GNDA.n440 GNDA.n439 24.4576
R3420 GNDA.n445 GNDA.n444 24.4576
R3421 GNDA.n2465 GNDA.t170 24.0005
R3422 GNDA.n2465 GNDA.t160 24.0005
R3423 GNDA.n2467 GNDA.t188 24.0005
R3424 GNDA.n2467 GNDA.t174 24.0005
R3425 GNDA.n2469 GNDA.t162 24.0005
R3426 GNDA.n2469 GNDA.t190 24.0005
R3427 GNDA.n2475 GNDA.t178 24.0005
R3428 GNDA.n2475 GNDA.t166 24.0005
R3429 GNDA.n2473 GNDA.t192 24.0005
R3430 GNDA.n2473 GNDA.t176 24.0005
R3431 GNDA.n2471 GNDA.t164 24.0005
R3432 GNDA.n2471 GNDA.t194 24.0005
R3433 GNDA.n554 GNDA.t180 24.0005
R3434 GNDA.n554 GNDA.t182 24.0005
R3435 GNDA.n2520 GNDA.t158 24.0005
R3436 GNDA.n2520 GNDA.t184 24.0005
R3437 GNDA.n2518 GNDA.t172 24.0005
R3438 GNDA.n2518 GNDA.t168 24.0005
R3439 GNDA.n514 GNDA.t156 24.0005
R3440 GNDA.n514 GNDA.t186 24.0005
R3441 GNDA.n2590 GNDA.t91 23.914
R3442 GNDA.n2589 GNDA.t27 23.914
R3443 GNDA.n2588 GNDA.t45 23.914
R3444 GNDA.n2587 GNDA.t129 23.914
R3445 GNDA.n2586 GNDA.t306 23.914
R3446 GNDA.n2526 GNDA.t47 23.6841
R3447 GNDA.t58 GNDA.n2540 23.6841
R3448 GNDA.n816 GNDA.t1 23.6841
R3449 GNDA.n229 GNDA.n227 23.6611
R3450 GNDA.n399 GNDA.n398 23.6611
R3451 GNDA.n206 GNDA.n205 22.8576
R3452 GNDA.n161 GNDA.n160 22.8576
R3453 GNDA.n491 GNDA.n490 22.8576
R3454 GNDA.n494 GNDA.n493 22.8576
R3455 GNDA.n468 GNDA.n467 22.8576
R3456 GNDA.n464 GNDA.n463 22.8576
R3457 GNDA.n406 GNDA.n141 22.8576
R3458 GNDA.n384 GNDA.n383 22.8576
R3459 GNDA.n368 GNDA.n367 22.8576
R3460 GNDA.n365 GNDA.n364 22.8576
R3461 GNDA.n323 GNDA.n322 22.8576
R3462 GNDA.n316 GNDA.n315 22.8576
R3463 GNDA.n94 GNDA.n93 22.8576
R3464 GNDA.n87 GNDA.n86 22.8576
R3465 GNDA.n1014 GNDA.t177 22.6544
R3466 GNDA.n2542 GNDA.t157 22.6544
R3467 GNDA.n2577 GNDA.t92 21.084
R3468 GNDA.n1439 GNDA.n1438 21.0192
R3469 GNDA.t86 GNDA.t296 20.9779
R3470 GNDA.n193 GNDA.t301 20.9249
R3471 GNDA.n2464 GNDA.n2463 20.8233
R3472 GNDA.n2482 GNDA.n2481 20.8233
R3473 GNDA.n2478 GNDA.n2477 20.8233
R3474 GNDA.n2516 GNDA.n2515 20.8233
R3475 GNDA.n2524 GNDA.n2523 20.8233
R3476 GNDA.n2575 GNDA.n2574 20.8233
R3477 GNDA.n132 GNDA.n1 20.7243
R3478 GNDA.n2598 GNDA.n2597 20.7243
R3479 GNDA.n2368 GNDA.t211 20.5949
R3480 GNDA.t82 GNDA.n2368 20.5949
R3481 GNDA.n2483 GNDA.t72 20.5949
R3482 GNDA.t47 GNDA.n2525 20.5949
R3483 GNDA.n2564 GNDA.t37 20.5949
R3484 GNDA.n2564 GNDA.t211 20.5949
R3485 GNDA.n615 GNDA.t211 19.9378
R3486 GNDA.n424 GNDA.t42 19.7005
R3487 GNDA.n424 GNDA.t144 19.7005
R3488 GNDA.n422 GNDA.t76 19.7005
R3489 GNDA.n422 GNDA.t89 19.7005
R3490 GNDA.n420 GNDA.t7 19.7005
R3491 GNDA.n420 GNDA.t147 19.7005
R3492 GNDA.n418 GNDA.t33 19.7005
R3493 GNDA.n418 GNDA.t30 19.7005
R3494 GNDA.n416 GNDA.t34 19.7005
R3495 GNDA.n416 GNDA.t95 19.7005
R3496 GNDA.n415 GNDA.t40 19.7005
R3497 GNDA.n415 GNDA.t43 19.7005
R3498 GNDA.n249 GNDA.t148 19.7005
R3499 GNDA.n249 GNDA.t150 19.7005
R3500 GNDA.n247 GNDA.t38 19.7005
R3501 GNDA.n247 GNDA.t106 19.7005
R3502 GNDA.n245 GNDA.t71 19.7005
R3503 GNDA.n245 GNDA.t320 19.7005
R3504 GNDA.n243 GNDA.t302 19.7005
R3505 GNDA.n243 GNDA.t29 19.7005
R3506 GNDA.n241 GNDA.t107 19.7005
R3507 GNDA.n241 GNDA.t291 19.7005
R3508 GNDA.n240 GNDA.t5 19.7005
R3509 GNDA.n240 GNDA.t149 19.7005
R3510 GNDA.n1483 GNDA.t211 19.6741
R3511 GNDA.t6 GNDA.t137 19.1977
R3512 GNDA.t304 GNDA.t94 19.1977
R3513 GNDA.t31 GNDA.n137 19.1977
R3514 GNDA.n2595 GNDA.t128 19.1977
R3515 GNDA.t21 GNDA.t313 19.1977
R3516 GNDA.t317 GNDA.t17 19.1977
R3517 GNDA.n397 GNDA.n396 19.0713
R3518 GNDA.n2602 GNDA.n2601 19.008
R3519 GNDA.n1441 GNDA.n1433 18.5605
R3520 GNDA.n2382 GNDA.t189 18.5355
R3521 GNDA.t181 GNDA.n881 18.5355
R3522 GNDA.t130 GNDA.n8 18.3557
R3523 GNDA GNDA.n518 18.1546
R3524 GNDA.n493 GNDA.n492 18.1442
R3525 GNDA.n366 GNDA.n365 18.1442
R3526 GNDA.n383 GNDA.n125 17.8005
R3527 GNDA.n1942 GNDA.n1938 17.5843
R3528 GNDA.n1806 GNDA.n1239 17.5843
R3529 GNDA.n785 GNDA.n781 17.5843
R3530 GNDA.n2462 GNDA.t211 17.5058
R3531 GNDA.n2577 GNDA.n2576 17.5058
R3532 GNDA.n1248 GNDA.t211 16.9844
R3533 GNDA.n1955 GNDA.t211 16.9844
R3534 GNDA.t211 GNDA.n526 16.9844
R3535 GNDA.n1506 GNDA.n1505 16.9379
R3536 GNDA.n2312 GNDA.n2294 16.9379
R3537 GNDA.n1104 GNDA.n1101 16.9379
R3538 GNDA.n1861 GNDA.n1860 16.7709
R3539 GNDA.n1048 GNDA.n1047 16.7709
R3540 GNDA.n2183 GNDA.n1125 16.7709
R3541 GNDA.n2509 GNDA.n582 16.7709
R3542 GNDA.n251 GNDA.n250 16.5057
R3543 GNDA.n213 GNDA.t206 16.0005
R3544 GNDA.n218 GNDA.t239 16.0005
R3545 GNDA.n222 GNDA.t218 16.0005
R3546 GNDA.n146 GNDA.t197 16.0005
R3547 GNDA.n401 GNDA.t280 16.0005
R3548 GNDA.n379 GNDA.t213 16.0005
R3549 GNDA.n471 GNDA.t290 16.0005
R3550 GNDA.n458 GNDA.t209 16.0005
R3551 GNDA.n140 GNDA.t285 16.0005
R3552 GNDA.n388 GNDA.t203 16.0005
R3553 GNDA.n131 GNDA.t269 16.0005
R3554 GNDA.n2591 GNDA.t275 16.0005
R3555 GNDA.n1637 GNDA.n1624 16.0005
R3556 GNDA.n1637 GNDA.n1636 16.0005
R3557 GNDA.n1636 GNDA.n1635 16.0005
R3558 GNDA.n1635 GNDA.n1632 16.0005
R3559 GNDA.n1632 GNDA.n1631 16.0005
R3560 GNDA.n1631 GNDA.n1628 16.0005
R3561 GNDA.n1628 GNDA.n1627 16.0005
R3562 GNDA.n1627 GNDA.n1268 16.0005
R3563 GNDA.n1623 GNDA.n1621 16.0005
R3564 GNDA.n1621 GNDA.n1618 16.0005
R3565 GNDA.n1618 GNDA.n1617 16.0005
R3566 GNDA.n1617 GNDA.n1614 16.0005
R3567 GNDA.n1614 GNDA.n1613 16.0005
R3568 GNDA.n1613 GNDA.n1610 16.0005
R3569 GNDA.n1610 GNDA.n1609 16.0005
R3570 GNDA.n1609 GNDA.n1606 16.0005
R3571 GNDA.n1605 GNDA.n1602 16.0005
R3572 GNDA.n1602 GNDA.n1601 16.0005
R3573 GNDA.n1601 GNDA.n1598 16.0005
R3574 GNDA.n1598 GNDA.n1597 16.0005
R3575 GNDA.n1597 GNDA.n1594 16.0005
R3576 GNDA.n1594 GNDA.n1593 16.0005
R3577 GNDA.n1593 GNDA.n1590 16.0005
R3578 GNDA.n1590 GNDA.n1589 16.0005
R3579 GNDA.n2438 GNDA.n2425 16.0005
R3580 GNDA.n2438 GNDA.n2437 16.0005
R3581 GNDA.n2437 GNDA.n2436 16.0005
R3582 GNDA.n2436 GNDA.n2433 16.0005
R3583 GNDA.n2433 GNDA.n2432 16.0005
R3584 GNDA.n2432 GNDA.n2429 16.0005
R3585 GNDA.n2429 GNDA.n2428 16.0005
R3586 GNDA.n2428 GNDA.n2319 16.0005
R3587 GNDA.n2424 GNDA.n2422 16.0005
R3588 GNDA.n2422 GNDA.n2419 16.0005
R3589 GNDA.n2419 GNDA.n2418 16.0005
R3590 GNDA.n2418 GNDA.n2415 16.0005
R3591 GNDA.n2415 GNDA.n2414 16.0005
R3592 GNDA.n2414 GNDA.n2411 16.0005
R3593 GNDA.n2411 GNDA.n2410 16.0005
R3594 GNDA.n2410 GNDA.n2407 16.0005
R3595 GNDA.n2406 GNDA.n2403 16.0005
R3596 GNDA.n2403 GNDA.n2402 16.0005
R3597 GNDA.n2402 GNDA.n2399 16.0005
R3598 GNDA.n2399 GNDA.n2398 16.0005
R3599 GNDA.n2398 GNDA.n2395 16.0005
R3600 GNDA.n2395 GNDA.n2394 16.0005
R3601 GNDA.n2394 GNDA.n2391 16.0005
R3602 GNDA.n2391 GNDA.n2390 16.0005
R3603 GNDA.n2243 GNDA.n2242 16.0005
R3604 GNDA.n2246 GNDA.n2243 16.0005
R3605 GNDA.n2247 GNDA.n2246 16.0005
R3606 GNDA.n2250 GNDA.n2247 16.0005
R3607 GNDA.n2251 GNDA.n2250 16.0005
R3608 GNDA.n2254 GNDA.n2251 16.0005
R3609 GNDA.n2255 GNDA.n2254 16.0005
R3610 GNDA.n2255 GNDA.n632 16.0005
R3611 GNDA.n2239 GNDA.n2238 16.0005
R3612 GNDA.n2238 GNDA.n2235 16.0005
R3613 GNDA.n2235 GNDA.n2234 16.0005
R3614 GNDA.n2234 GNDA.n2231 16.0005
R3615 GNDA.n2231 GNDA.n2230 16.0005
R3616 GNDA.n2230 GNDA.n2227 16.0005
R3617 GNDA.n2227 GNDA.n2226 16.0005
R3618 GNDA.n2226 GNDA.n2223 16.0005
R3619 GNDA.n2222 GNDA.n2219 16.0005
R3620 GNDA.n2219 GNDA.n2218 16.0005
R3621 GNDA.n2218 GNDA.n2215 16.0005
R3622 GNDA.n2215 GNDA.n2214 16.0005
R3623 GNDA.n2214 GNDA.n2211 16.0005
R3624 GNDA.n2211 GNDA.n2210 16.0005
R3625 GNDA.n2210 GNDA.n2207 16.0005
R3626 GNDA.n2207 GNDA.n2206 16.0005
R3627 GNDA.n2132 GNDA.n2131 16.0005
R3628 GNDA.n2135 GNDA.n2132 16.0005
R3629 GNDA.n2136 GNDA.n2135 16.0005
R3630 GNDA.n2139 GNDA.n2136 16.0005
R3631 GNDA.n2140 GNDA.n2139 16.0005
R3632 GNDA.n2143 GNDA.n2140 16.0005
R3633 GNDA.n2144 GNDA.n2143 16.0005
R3634 GNDA.n2144 GNDA.n1151 16.0005
R3635 GNDA.n2128 GNDA.n2127 16.0005
R3636 GNDA.n2127 GNDA.n2124 16.0005
R3637 GNDA.n2124 GNDA.n2123 16.0005
R3638 GNDA.n2123 GNDA.n2120 16.0005
R3639 GNDA.n2120 GNDA.n2119 16.0005
R3640 GNDA.n2119 GNDA.n2116 16.0005
R3641 GNDA.n2116 GNDA.n2115 16.0005
R3642 GNDA.n2115 GNDA.n2112 16.0005
R3643 GNDA.n2111 GNDA.n2108 16.0005
R3644 GNDA.n2108 GNDA.n2107 16.0005
R3645 GNDA.n2107 GNDA.n2104 16.0005
R3646 GNDA.n2104 GNDA.n2103 16.0005
R3647 GNDA.n2103 GNDA.n2100 16.0005
R3648 GNDA.n2100 GNDA.n2099 16.0005
R3649 GNDA.n2099 GNDA.n2096 16.0005
R3650 GNDA.n2096 GNDA.n2095 16.0005
R3651 GNDA.n2037 GNDA.n2036 16.0005
R3652 GNDA.n2040 GNDA.n2037 16.0005
R3653 GNDA.n2041 GNDA.n2040 16.0005
R3654 GNDA.n2044 GNDA.n2041 16.0005
R3655 GNDA.n2045 GNDA.n2044 16.0005
R3656 GNDA.n2048 GNDA.n2045 16.0005
R3657 GNDA.n2049 GNDA.n2048 16.0005
R3658 GNDA.n2049 GNDA.n1172 16.0005
R3659 GNDA.n2033 GNDA.n2032 16.0005
R3660 GNDA.n2032 GNDA.n2029 16.0005
R3661 GNDA.n2029 GNDA.n2028 16.0005
R3662 GNDA.n2028 GNDA.n2025 16.0005
R3663 GNDA.n2025 GNDA.n2024 16.0005
R3664 GNDA.n2024 GNDA.n2021 16.0005
R3665 GNDA.n2021 GNDA.n2020 16.0005
R3666 GNDA.n2020 GNDA.n2017 16.0005
R3667 GNDA.n2016 GNDA.n2013 16.0005
R3668 GNDA.n2013 GNDA.n2012 16.0005
R3669 GNDA.n2012 GNDA.n2009 16.0005
R3670 GNDA.n2009 GNDA.n2008 16.0005
R3671 GNDA.n2008 GNDA.n2005 16.0005
R3672 GNDA.n2005 GNDA.n2004 16.0005
R3673 GNDA.n2004 GNDA.n2001 16.0005
R3674 GNDA.n2001 GNDA.n2000 16.0005
R3675 GNDA.n1386 GNDA.n1385 16.0005
R3676 GNDA.n1389 GNDA.n1386 16.0005
R3677 GNDA.n1390 GNDA.n1389 16.0005
R3678 GNDA.n1393 GNDA.n1390 16.0005
R3679 GNDA.n1394 GNDA.n1393 16.0005
R3680 GNDA.n1397 GNDA.n1394 16.0005
R3681 GNDA.n1398 GNDA.n1397 16.0005
R3682 GNDA.n1398 GNDA.n1296 16.0005
R3683 GNDA.n1382 GNDA.n1381 16.0005
R3684 GNDA.n1381 GNDA.n1378 16.0005
R3685 GNDA.n1378 GNDA.n1377 16.0005
R3686 GNDA.n1377 GNDA.n1374 16.0005
R3687 GNDA.n1374 GNDA.n1373 16.0005
R3688 GNDA.n1373 GNDA.n1370 16.0005
R3689 GNDA.n1370 GNDA.n1369 16.0005
R3690 GNDA.n1369 GNDA.n1366 16.0005
R3691 GNDA.n1365 GNDA.n1362 16.0005
R3692 GNDA.n1362 GNDA.n1361 16.0005
R3693 GNDA.n1361 GNDA.n1358 16.0005
R3694 GNDA.n1358 GNDA.n1357 16.0005
R3695 GNDA.n1357 GNDA.n1354 16.0005
R3696 GNDA.n1354 GNDA.n1353 16.0005
R3697 GNDA.n1353 GNDA.n1350 16.0005
R3698 GNDA.n1350 GNDA.n1349 16.0005
R3699 GNDA.n1717 GNDA.n1675 16.0005
R3700 GNDA.n1723 GNDA.n1675 16.0005
R3701 GNDA.n1724 GNDA.n1723 16.0005
R3702 GNDA.n1725 GNDA.n1724 16.0005
R3703 GNDA.n1725 GNDA.n1673 16.0005
R3704 GNDA.n1731 GNDA.n1673 16.0005
R3705 GNDA.n1732 GNDA.n1731 16.0005
R3706 GNDA.n1736 GNDA.n1732 16.0005
R3707 GNDA.n1716 GNDA.n1715 16.0005
R3708 GNDA.n1715 GNDA.n1677 16.0005
R3709 GNDA.n1709 GNDA.n1677 16.0005
R3710 GNDA.n1709 GNDA.n1708 16.0005
R3711 GNDA.n1708 GNDA.n1707 16.0005
R3712 GNDA.n1707 GNDA.n1679 16.0005
R3713 GNDA.n1701 GNDA.n1679 16.0005
R3714 GNDA.n1701 GNDA.n1700 16.0005
R3715 GNDA.n1699 GNDA.n1681 16.0005
R3716 GNDA.n1693 GNDA.n1681 16.0005
R3717 GNDA.n1693 GNDA.n1692 16.0005
R3718 GNDA.n1692 GNDA.n1691 16.0005
R3719 GNDA.n1691 GNDA.n1683 16.0005
R3720 GNDA.n1686 GNDA.n1683 16.0005
R3721 GNDA.n1686 GNDA.n1659 16.0005
R3722 GNDA.n1771 GNDA.n1659 16.0005
R3723 GNDA.n993 GNDA.n979 16.0005
R3724 GNDA.n993 GNDA.n992 16.0005
R3725 GNDA.n992 GNDA.n991 16.0005
R3726 GNDA.n991 GNDA.n988 16.0005
R3727 GNDA.n988 GNDA.n987 16.0005
R3728 GNDA.n987 GNDA.n984 16.0005
R3729 GNDA.n984 GNDA.n983 16.0005
R3730 GNDA.n983 GNDA.n980 16.0005
R3731 GNDA.n978 GNDA.n976 16.0005
R3732 GNDA.n976 GNDA.n973 16.0005
R3733 GNDA.n973 GNDA.n972 16.0005
R3734 GNDA.n972 GNDA.n969 16.0005
R3735 GNDA.n969 GNDA.n968 16.0005
R3736 GNDA.n968 GNDA.n965 16.0005
R3737 GNDA.n965 GNDA.n964 16.0005
R3738 GNDA.n964 GNDA.n961 16.0005
R3739 GNDA.n960 GNDA.n957 16.0005
R3740 GNDA.n957 GNDA.n956 16.0005
R3741 GNDA.n956 GNDA.n953 16.0005
R3742 GNDA.n953 GNDA.n952 16.0005
R3743 GNDA.n952 GNDA.n949 16.0005
R3744 GNDA.n949 GNDA.n948 16.0005
R3745 GNDA.n948 GNDA.n945 16.0005
R3746 GNDA.n945 GNDA.n944 16.0005
R3747 GNDA.n861 GNDA.n860 16.0005
R3748 GNDA.n864 GNDA.n861 16.0005
R3749 GNDA.n865 GNDA.n864 16.0005
R3750 GNDA.n868 GNDA.n865 16.0005
R3751 GNDA.n869 GNDA.n868 16.0005
R3752 GNDA.n872 GNDA.n869 16.0005
R3753 GNDA.n874 GNDA.n872 16.0005
R3754 GNDA.n875 GNDA.n874 16.0005
R3755 GNDA.n857 GNDA.n856 16.0005
R3756 GNDA.n856 GNDA.n853 16.0005
R3757 GNDA.n853 GNDA.n852 16.0005
R3758 GNDA.n852 GNDA.n849 16.0005
R3759 GNDA.n849 GNDA.n848 16.0005
R3760 GNDA.n848 GNDA.n845 16.0005
R3761 GNDA.n845 GNDA.n844 16.0005
R3762 GNDA.n844 GNDA.n841 16.0005
R3763 GNDA.n840 GNDA.n837 16.0005
R3764 GNDA.n837 GNDA.n836 16.0005
R3765 GNDA.n836 GNDA.n833 16.0005
R3766 GNDA.n833 GNDA.n832 16.0005
R3767 GNDA.n832 GNDA.n829 16.0005
R3768 GNDA.n829 GNDA.n828 16.0005
R3769 GNDA.n828 GNDA.n825 16.0005
R3770 GNDA.n825 GNDA.n824 16.0005
R3771 GNDA.n1440 GNDA.n1439 16.0005
R3772 GNDA.n1441 GNDA.n1440 16.0005
R3773 GNDA.t189 GNDA.t310 15.4463
R3774 GNDA.t157 GNDA.t295 15.4463
R3775 GNDA.n322 GNDA.n321 14.9255
R3776 GNDA.n318 GNDA.n316 14.9255
R3777 GNDA.n93 GNDA.n92 14.9255
R3778 GNDA.n89 GNDA.n87 14.9255
R3779 GNDA.n217 GNDA.n216 14.8213
R3780 GNDA.n230 GNDA.n229 14.8213
R3781 GNDA.n398 GNDA.n397 14.8213
R3782 GNDA.n2199 GNDA.n2198 14.555
R3783 GNDA.n1656 GNDA.n1252 14.555
R3784 GNDA.n444 GNDA.n443 14.4047
R3785 GNDA.n2466 GNDA.n2464 14.363
R3786 GNDA.n163 GNDA.n161 14.0818
R3787 GNDA.n2599 GNDA.n2598 14.0401
R3788 GNDA.n492 GNDA.n491 14.0193
R3789 GNDA.n367 GNDA.n366 14.0193
R3790 GNDA.n2481 GNDA.n2480 13.8005
R3791 GNDA.n2479 GNDA.n2478 13.8005
R3792 GNDA.n2517 GNDA.n2516 13.8005
R3793 GNDA.n2523 GNDA.n2522 13.8005
R3794 GNDA.n2574 GNDA.n2573 13.8005
R3795 GNDA.n207 GNDA.n206 13.8005
R3796 GNDA.n467 GNDA.n466 13.8005
R3797 GNDA.n465 GNDA.n464 13.8005
R3798 GNDA.n141 GNDA.n125 13.8005
R3799 GNDA.n441 GNDA.n440 13.8005
R3800 GNDA.n2568 GNDA.n2567 12.7542
R3801 GNDA.n319 GNDA.n3 12.6567
R3802 GNDA.n90 GNDA.n2 12.6567
R3803 GNDA.n2448 GNDA.t187 12.3572
R3804 GNDA.t163 GNDA.n926 12.3572
R3805 GNDA.t155 GNDA.n810 12.3572
R3806 GNDA.n1016 GNDA.n519 12.2193
R3807 GNDA.t46 GNDA.t50 11.7135
R3808 GNDA.n426 GNDA.n425 11.6932
R3809 GNDA.n1505 GNDA.n1503 11.6369
R3810 GNDA.n1503 GNDA.n1500 11.6369
R3811 GNDA.n1500 GNDA.n1499 11.6369
R3812 GNDA.n1499 GNDA.n1496 11.6369
R3813 GNDA.n1496 GNDA.n1495 11.6369
R3814 GNDA.n1495 GNDA.n1492 11.6369
R3815 GNDA.n1492 GNDA.n1491 11.6369
R3816 GNDA.n1491 GNDA.n1488 11.6369
R3817 GNDA.n1488 GNDA.n1487 11.6369
R3818 GNDA.n1487 GNDA.n1485 11.6369
R3819 GNDA.n2294 GNDA.n2293 11.6369
R3820 GNDA.n2293 GNDA.n2290 11.6369
R3821 GNDA.n2290 GNDA.n2289 11.6369
R3822 GNDA.n2289 GNDA.n2286 11.6369
R3823 GNDA.n2286 GNDA.n2285 11.6369
R3824 GNDA.n2285 GNDA.n2282 11.6369
R3825 GNDA.n2282 GNDA.n2281 11.6369
R3826 GNDA.n2281 GNDA.n2278 11.6369
R3827 GNDA.n2278 GNDA.n2277 11.6369
R3828 GNDA.n2277 GNDA.n580 11.6369
R3829 GNDA.n2510 GNDA.n580 11.6369
R3830 GNDA.n2312 GNDA.n2311 11.6369
R3831 GNDA.n2311 GNDA.n2310 11.6369
R3832 GNDA.n2310 GNDA.n2308 11.6369
R3833 GNDA.n2308 GNDA.n2305 11.6369
R3834 GNDA.n2305 GNDA.n2304 11.6369
R3835 GNDA.n2304 GNDA.n2301 11.6369
R3836 GNDA.n2301 GNDA.n2300 11.6369
R3837 GNDA.n2300 GNDA.n2297 11.6369
R3838 GNDA.n2297 GNDA.n2296 11.6369
R3839 GNDA.n2296 GNDA.n613 11.6369
R3840 GNDA.n1101 GNDA.n1100 11.6369
R3841 GNDA.n1100 GNDA.n1097 11.6369
R3842 GNDA.n1097 GNDA.n1096 11.6369
R3843 GNDA.n1096 GNDA.n1093 11.6369
R3844 GNDA.n1093 GNDA.n1092 11.6369
R3845 GNDA.n1092 GNDA.n1089 11.6369
R3846 GNDA.n1089 GNDA.n1088 11.6369
R3847 GNDA.n1088 GNDA.n1085 11.6369
R3848 GNDA.n1085 GNDA.n1084 11.6369
R3849 GNDA.n1084 GNDA.n1081 11.6369
R3850 GNDA.n1105 GNDA.n1104 11.6369
R3851 GNDA.n1108 GNDA.n1105 11.6369
R3852 GNDA.n1109 GNDA.n1108 11.6369
R3853 GNDA.n1112 GNDA.n1109 11.6369
R3854 GNDA.n1113 GNDA.n1112 11.6369
R3855 GNDA.n1116 GNDA.n1113 11.6369
R3856 GNDA.n1117 GNDA.n1116 11.6369
R3857 GNDA.n1120 GNDA.n1117 11.6369
R3858 GNDA.n1122 GNDA.n1120 11.6369
R3859 GNDA.n1123 GNDA.n1122 11.6369
R3860 GNDA.n2184 GNDA.n1123 11.6369
R3861 GNDA.n1943 GNDA.n1942 11.6369
R3862 GNDA.n1944 GNDA.n1943 11.6369
R3863 GNDA.n1944 GNDA.n1200 11.6369
R3864 GNDA.n1951 GNDA.n1200 11.6369
R3865 GNDA.n1952 GNDA.n1951 11.6369
R3866 GNDA.n1953 GNDA.n1952 11.6369
R3867 GNDA.n1953 GNDA.n1197 11.6369
R3868 GNDA.n1960 GNDA.n1197 11.6369
R3869 GNDA.n1961 GNDA.n1960 11.6369
R3870 GNDA.n1962 GNDA.n1961 11.6369
R3871 GNDA.n1918 GNDA.n1917 11.6369
R3872 GNDA.n1921 GNDA.n1918 11.6369
R3873 GNDA.n1922 GNDA.n1921 11.6369
R3874 GNDA.n1925 GNDA.n1922 11.6369
R3875 GNDA.n1926 GNDA.n1925 11.6369
R3876 GNDA.n1929 GNDA.n1926 11.6369
R3877 GNDA.n1930 GNDA.n1929 11.6369
R3878 GNDA.n1933 GNDA.n1930 11.6369
R3879 GNDA.n1934 GNDA.n1933 11.6369
R3880 GNDA.n1937 GNDA.n1934 11.6369
R3881 GNDA.n1938 GNDA.n1937 11.6369
R3882 GNDA.n1863 GNDA.n1124 11.6369
R3883 GNDA.n1866 GNDA.n1863 11.6369
R3884 GNDA.n1867 GNDA.n1866 11.6369
R3885 GNDA.n1870 GNDA.n1867 11.6369
R3886 GNDA.n1871 GNDA.n1870 11.6369
R3887 GNDA.n1874 GNDA.n1871 11.6369
R3888 GNDA.n1875 GNDA.n1874 11.6369
R3889 GNDA.n1878 GNDA.n1875 11.6369
R3890 GNDA.n1879 GNDA.n1878 11.6369
R3891 GNDA.n1882 GNDA.n1879 11.6369
R3892 GNDA.n1883 GNDA.n1882 11.6369
R3893 GNDA.n1824 GNDA.n1230 11.6369
R3894 GNDA.n1824 GNDA.n1823 11.6369
R3895 GNDA.n1823 GNDA.n1822 11.6369
R3896 GNDA.n1822 GNDA.n1231 11.6369
R3897 GNDA.n1816 GNDA.n1231 11.6369
R3898 GNDA.n1816 GNDA.n1815 11.6369
R3899 GNDA.n1815 GNDA.n1814 11.6369
R3900 GNDA.n1814 GNDA.n1234 11.6369
R3901 GNDA.n1808 GNDA.n1234 11.6369
R3902 GNDA.n1808 GNDA.n1807 11.6369
R3903 GNDA.n1807 GNDA.n1806 11.6369
R3904 GNDA.n1800 GNDA.n1239 11.6369
R3905 GNDA.n1800 GNDA.n1799 11.6369
R3906 GNDA.n1799 GNDA.n1798 11.6369
R3907 GNDA.n1798 GNDA.n1243 11.6369
R3908 GNDA.n1792 GNDA.n1243 11.6369
R3909 GNDA.n1792 GNDA.n1791 11.6369
R3910 GNDA.n1791 GNDA.n1790 11.6369
R3911 GNDA.n1790 GNDA.n1246 11.6369
R3912 GNDA.n1784 GNDA.n1246 11.6369
R3913 GNDA.n1784 GNDA.n1783 11.6369
R3914 GNDA.n786 GNDA.n785 11.6369
R3915 GNDA.n788 GNDA.n786 11.6369
R3916 GNDA.n788 GNDA.n787 11.6369
R3917 GNDA.n787 GNDA.n758 11.6369
R3918 GNDA.n758 GNDA.n756 11.6369
R3919 GNDA.n796 GNDA.n756 11.6369
R3920 GNDA.n797 GNDA.n796 11.6369
R3921 GNDA.n798 GNDA.n797 11.6369
R3922 GNDA.n798 GNDA.n751 11.6369
R3923 GNDA.n806 GNDA.n751 11.6369
R3924 GNDA.n761 GNDA.n698 11.6369
R3925 GNDA.n764 GNDA.n761 11.6369
R3926 GNDA.n765 GNDA.n764 11.6369
R3927 GNDA.n768 GNDA.n765 11.6369
R3928 GNDA.n769 GNDA.n768 11.6369
R3929 GNDA.n772 GNDA.n769 11.6369
R3930 GNDA.n773 GNDA.n772 11.6369
R3931 GNDA.n776 GNDA.n773 11.6369
R3932 GNDA.n777 GNDA.n776 11.6369
R3933 GNDA.n780 GNDA.n777 11.6369
R3934 GNDA.n781 GNDA.n780 11.6369
R3935 GNDA.n699 GNDA.n581 11.6369
R3936 GNDA.n702 GNDA.n699 11.6369
R3937 GNDA.n703 GNDA.n702 11.6369
R3938 GNDA.n706 GNDA.n703 11.6369
R3939 GNDA.n707 GNDA.n706 11.6369
R3940 GNDA.n710 GNDA.n707 11.6369
R3941 GNDA.n711 GNDA.n710 11.6369
R3942 GNDA.n714 GNDA.n711 11.6369
R3943 GNDA.n715 GNDA.n714 11.6369
R3944 GNDA.n718 GNDA.n715 11.6369
R3945 GNDA.n719 GNDA.n718 11.6369
R3946 GNDA.n1471 GNDA.n1470 11.6369
R3947 GNDA.n1470 GNDA.n1428 11.6369
R3948 GNDA.n1464 GNDA.n1428 11.6369
R3949 GNDA.n1464 GNDA.n1463 11.6369
R3950 GNDA.n1463 GNDA.n1462 11.6369
R3951 GNDA.n1456 GNDA.n1445 11.6369
R3952 GNDA.n1456 GNDA.n1455 11.6369
R3953 GNDA.n1455 GNDA.n1454 11.6369
R3954 GNDA.n1454 GNDA.n1446 11.6369
R3955 GNDA.n1448 GNDA.n1446 11.6369
R3956 GNDA.n1507 GNDA.n1506 11.6369
R3957 GNDA.n1507 GNDA.n1481 11.6369
R3958 GNDA.n1513 GNDA.n1481 11.6369
R3959 GNDA.n1514 GNDA.n1513 11.6369
R3960 GNDA.n1515 GNDA.n1514 11.6369
R3961 GNDA.n1515 GNDA.n1477 11.6369
R3962 GNDA.n1521 GNDA.n1477 11.6369
R3963 GNDA.n1522 GNDA.n1521 11.6369
R3964 GNDA.n1524 GNDA.n1522 11.6369
R3965 GNDA.n1524 GNDA.n1523 11.6369
R3966 GNDA.n1523 GNDA.n1474 11.6369
R3967 GNDA.t123 GNDA.t19 11.5188
R3968 GNDA.n404 GNDA.t115 11.5188
R3969 GNDA.n2595 GNDA.t80 11.5188
R3970 GNDA.n2573 GNDA.n2572 11.3792
R3971 GNDA.n251 GNDA.n3 10.8286
R3972 GNDA.n441 GNDA.n426 9.99008
R3973 GNDA.n516 GNDA.n0 9.75668
R3974 GNDA.n2365 GNDA.t132 9.6005
R3975 GNDA.n2355 GNDA.t134 9.6005
R3976 GNDA.n2558 GNDA.t152 9.6005
R3977 GNDA.n521 GNDA.t133 9.6005
R3978 GNDA.n196 GNDA.t283 9.6005
R3979 GNDA.n182 GNDA.t312 9.6005
R3980 GNDA.n182 GNDA.t114 9.6005
R3981 GNDA.n180 GNDA.t62 9.6005
R3982 GNDA.n180 GNDA.t9 9.6005
R3983 GNDA.n178 GNDA.t124 9.6005
R3984 GNDA.n178 GNDA.t140 9.6005
R3985 GNDA.n176 GNDA.t64 9.6005
R3986 GNDA.n176 GNDA.t103 9.6005
R3987 GNDA.n174 GNDA.t23 9.6005
R3988 GNDA.n174 GNDA.t122 9.6005
R3989 GNDA.n172 GNDA.t142 9.6005
R3990 GNDA.n172 GNDA.t70 9.6005
R3991 GNDA.n170 GNDA.t116 9.6005
R3992 GNDA.n170 GNDA.t120 9.6005
R3993 GNDA.n168 GNDA.t110 9.6005
R3994 GNDA.n168 GNDA.t66 9.6005
R3995 GNDA.n166 GNDA.t81 9.6005
R3996 GNDA.n166 GNDA.t322 9.6005
R3997 GNDA.n164 GNDA.t68 9.6005
R3998 GNDA.n164 GNDA.t309 9.6005
R3999 GNDA.n162 GNDA.t112 9.6005
R4000 GNDA.n162 GNDA.t224 9.6005
R4001 GNDA.n154 GNDA.t225 9.6005
R4002 GNDA.n433 GNDA.t278 9.6005
R4003 GNDA.n442 GNDA.t53 9.6005
R4004 GNDA.n442 GNDA.t118 9.6005
R4005 GNDA.n414 GNDA.t229 9.6005
R4006 GNDA.n2601 GNDA.n1 9.54008
R4007 GNDA.t2 GNDA.t211 9.37093
R4008 GNDA.n201 GNDA.n200 9.14336
R4009 GNDA.n198 GNDA.n197 9.14336
R4010 GNDA.n153 GNDA.n150 9.14336
R4011 GNDA.n157 GNDA.n156 9.14336
R4012 GNDA.n381 GNDA.n380 9.14336
R4013 GNDA.n484 GNDA.n479 9.14336
R4014 GNDA.n484 GNDA.n483 9.14336
R4015 GNDA.n483 GNDA.n481 9.14336
R4016 GNDA.n500 GNDA.n20 9.14336
R4017 GNDA.n500 GNDA.n499 9.14336
R4018 GNDA.n499 GNDA.n497 9.14336
R4019 GNDA.n473 GNDA.n470 9.14336
R4020 GNDA.n460 GNDA.n459 9.14336
R4021 GNDA.n409 GNDA.n408 9.14336
R4022 GNDA.n390 GNDA.n387 9.14336
R4023 GNDA.n432 GNDA.n429 9.14336
R4024 GNDA.n436 GNDA.n435 9.14336
R4025 GNDA.n452 GNDA.n451 9.14336
R4026 GNDA.n449 GNDA.n448 9.14336
R4027 GNDA.n135 GNDA.n134 9.14336
R4028 GNDA.n2593 GNDA.n2592 9.14336
R4029 GNDA.n374 GNDA.n238 9.14336
R4030 GNDA.n374 GNDA.n373 9.14336
R4031 GNDA.n373 GNDA.n371 9.14336
R4032 GNDA.n358 GNDA.n353 9.14336
R4033 GNDA.n358 GNDA.n357 9.14336
R4034 GNDA.n357 GNDA.n355 9.14336
R4035 GNDA.n345 GNDA.n262 9.14336
R4036 GNDA.n345 GNDA.n344 9.14336
R4037 GNDA.n344 GNDA.n342 9.14336
R4038 GNDA.n342 GNDA.n339 9.14336
R4039 GNDA.n339 GNDA.n338 9.14336
R4040 GNDA.n338 GNDA.n335 9.14336
R4041 GNDA.n335 GNDA.n334 9.14336
R4042 GNDA.n334 GNDA.n331 9.14336
R4043 GNDA.n331 GNDA.n330 9.14336
R4044 GNDA.n330 GNDA.n327 9.14336
R4045 GNDA.n327 GNDA.n326 9.14336
R4046 GNDA.n286 GNDA.n283 9.14336
R4047 GNDA.n290 GNDA.n283 9.14336
R4048 GNDA.n290 GNDA.n281 9.14336
R4049 GNDA.n296 GNDA.n281 9.14336
R4050 GNDA.n296 GNDA.n279 9.14336
R4051 GNDA.n300 GNDA.n279 9.14336
R4052 GNDA.n300 GNDA.n277 9.14336
R4053 GNDA.n306 GNDA.n277 9.14336
R4054 GNDA.n306 GNDA.n275 9.14336
R4055 GNDA.n310 GNDA.n275 9.14336
R4056 GNDA.n310 GNDA.n273 9.14336
R4057 GNDA.n116 GNDA.n33 9.14336
R4058 GNDA.n116 GNDA.n115 9.14336
R4059 GNDA.n115 GNDA.n113 9.14336
R4060 GNDA.n113 GNDA.n110 9.14336
R4061 GNDA.n110 GNDA.n109 9.14336
R4062 GNDA.n109 GNDA.n106 9.14336
R4063 GNDA.n106 GNDA.n105 9.14336
R4064 GNDA.n105 GNDA.n102 9.14336
R4065 GNDA.n102 GNDA.n101 9.14336
R4066 GNDA.n101 GNDA.n98 9.14336
R4067 GNDA.n98 GNDA.n97 9.14336
R4068 GNDA.n57 GNDA.n54 9.14336
R4069 GNDA.n61 GNDA.n54 9.14336
R4070 GNDA.n61 GNDA.n52 9.14336
R4071 GNDA.n67 GNDA.n52 9.14336
R4072 GNDA.n67 GNDA.n50 9.14336
R4073 GNDA.n71 GNDA.n50 9.14336
R4074 GNDA.n71 GNDA.n48 9.14336
R4075 GNDA.n77 GNDA.n48 9.14336
R4076 GNDA.n77 GNDA.n46 9.14336
R4077 GNDA.n81 GNDA.n46 9.14336
R4078 GNDA.n81 GNDA.n44 9.14336
R4079 GNDA.n2585 GNDA.t303 8.96839
R4080 GNDA.n2198 GNDA.n2197 8.60107
R4081 GNDA.n1252 GNDA.n1206 8.60107
R4082 GNDA.n212 GNDA.n211 8.53383
R4083 GNDA.t159 GNDA.n2449 8.23827
R4084 GNDA.t175 GNDA.n1003 8.23827
R4085 GNDA.t167 GNDA.n2553 8.23827
R4086 GNDA.n2577 GNDA.n512 8.19962
R4087 GNDA.t22 GNDA.t238 7.67938
R4088 GNDA.t121 GNDA.t31 7.67938
R4089 GNDA.t141 GNDA.t57 7.67938
R4090 GNDA.t69 GNDA.t87 7.67938
R4091 GNDA.t115 GNDA.t75 7.67938
R4092 GNDA.t14 GNDA.t119 7.67938
R4093 GNDA.t109 GNDA.t20 7.67938
R4094 GNDA.t274 GNDA.t65 7.67938
R4095 GNDA.n518 GNDA.n517 7.56675
R4096 GNDA.n1437 GNDA.n516 7.56675
R4097 GNDA.t18 GNDA.n2382 7.20855
R4098 GNDA.n2530 GNDA.t37 7.20855
R4099 GNDA.t48 GNDA.n817 7.20855
R4100 GNDA.n2576 GNDA.n513 7.20855
R4101 GNDA.n208 GNDA.n207 7.03175
R4102 GNDA.n2510 GNDA.n2509 6.72373
R4103 GNDA.n2184 GNDA.n2183 6.72373
R4104 GNDA.n1883 GNDA.n1861 6.72373
R4105 GNDA.n1047 GNDA.n719 6.72373
R4106 GNDA.n1448 GNDA.n1447 6.72373
R4107 GNDA.n1474 GNDA.n1472 6.72373
R4108 GNDA.n208 GNDA.n2 6.688
R4109 GNDA.n2600 GNDA.n2 6.28175
R4110 GNDA.n1917 GNDA.n1861 6.20656
R4111 GNDA.n2183 GNDA.n1124 6.20656
R4112 GNDA.n1447 GNDA.n1230 6.20656
R4113 GNDA.n1047 GNDA.n698 6.20656
R4114 GNDA.n2509 GNDA.n581 6.20656
R4115 GNDA.n1472 GNDA.n1471 6.20656
R4116 GNDA.t211 GNDA.t35 6.17883
R4117 GNDA.n1462 GNDA.n1433 6.07727
R4118 GNDA.n2366 GNDA.n2356 5.81868
R4119 GNDA.n2359 GNDA.n2356 5.81868
R4120 GNDA.n490 GNDA.n23 5.78934
R4121 GNDA.n495 GNDA.n494 5.78934
R4122 GNDA.n369 GNDA.n368 5.78934
R4123 GNDA.n364 GNDA.n252 5.78934
R4124 GNDA.n324 GNDA.n323 5.78934
R4125 GNDA.n315 GNDA.n272 5.78934
R4126 GNDA.n95 GNDA.n94 5.78934
R4127 GNDA.n86 GNDA.n43 5.78934
R4128 GNDA.n518 GNDA.n0 5.737
R4129 GNDA.n1445 GNDA.n1433 5.5601
R4130 GNDA.n492 GNDA.n22 5.54068
R4131 GNDA.n366 GNDA.n251 5.54068
R4132 GNDA.n1589 GNDA.n1567 5.51161
R4133 GNDA.n2390 GNDA.n2349 5.51161
R4134 GNDA.n2206 GNDA.n654 5.51161
R4135 GNDA.n2095 GNDA.n2065 5.51161
R4136 GNDA.n2000 GNDA.n1970 5.51161
R4137 GNDA.n1349 GNDA.n1319 5.51161
R4138 GNDA.n1772 GNDA.n1771 5.51161
R4139 GNDA.n944 GNDA.n915 5.51161
R4140 GNDA.n824 GNDA.n746 5.51161
R4141 GNDA.n217 GNDA.n209 5.46925
R4142 GNDA.n466 GNDA.n124 5.46925
R4143 GNDA.n1969 GNDA.n1193 5.1717
R4144 GNDA.n1782 GNDA.n1251 5.1717
R4145 GNDA.n808 GNDA.n807 5.1717
R4146 GNDA.n925 GNDA.t211 5.14911
R4147 GNDA.t263 GNDA.t104 5.14911
R4148 GNDA.n425 GNDA.n423 5.063
R4149 GNDA.n250 GNDA.n248 5.063
R4150 GNDA.n1653 GNDA.n1267 4.9157
R4151 GNDA.n2459 GNDA.n2318 4.9157
R4152 GNDA.n2267 GNDA.n631 4.9157
R4153 GNDA.n192 GNDA.t282 4.63906
R4154 GNDA.n191 GNDA.t311 4.63906
R4155 GNDA.n190 GNDA.t113 4.63906
R4156 GNDA.n189 GNDA.t61 4.63906
R4157 GNDA.n188 GNDA.t8 4.63906
R4158 GNDA.n187 GNDA.t139 4.63906
R4159 GNDA.n2601 GNDA.n2600 4.5005
R4160 GNDA.n200 GNDA.n199 4.46219
R4161 GNDA.n197 GNDA.n184 4.46219
R4162 GNDA.n199 GNDA.n198 4.46219
R4163 GNDA.n205 GNDA.n184 4.46219
R4164 GNDA.n155 GNDA.n150 4.46219
R4165 GNDA.n157 GNDA.n148 4.46219
R4166 GNDA.n156 GNDA.n155 4.46219
R4167 GNDA.n160 GNDA.n148 4.46219
R4168 GNDA.n380 GNDA.n231 4.46219
R4169 GNDA.n395 GNDA.n231 4.46219
R4170 GNDA.n473 GNDA.n472 4.46219
R4171 GNDA.n472 GNDA.n468 4.46219
R4172 GNDA.n460 GNDA.n126 4.46219
R4173 GNDA.n463 GNDA.n126 4.46219
R4174 GNDA.n408 GNDA.n407 4.46219
R4175 GNDA.n407 GNDA.n406 4.46219
R4176 GNDA.n390 GNDA.n389 4.46219
R4177 GNDA.n389 GNDA.n384 4.46219
R4178 GNDA.n434 GNDA.n429 4.46219
R4179 GNDA.n436 GNDA.n427 4.46219
R4180 GNDA.n435 GNDA.n434 4.46219
R4181 GNDA.n439 GNDA.n427 4.46219
R4182 GNDA.n451 GNDA.n450 4.46219
R4183 GNDA.n448 GNDA.n446 4.46219
R4184 GNDA.n450 GNDA.n449 4.46219
R4185 GNDA.n446 GNDA.n445 4.46219
R4186 GNDA.n134 GNDA.n133 4.46219
R4187 GNDA.n133 GNDA.n132 4.46219
R4188 GNDA.n2592 GNDA.n4 4.46219
R4189 GNDA.n2597 GNDA.n4 4.46219
R4190 GNDA.n2590 GNDA.t321 4.32986
R4191 GNDA.n2589 GNDA.t67 4.32986
R4192 GNDA.n2588 GNDA.t308 4.32986
R4193 GNDA.n2587 GNDA.t111 4.32986
R4194 GNDA.n2586 GNDA.t223 4.32986
R4195 GNDA.n1832 GNDA.n1225 4.26717
R4196 GNDA.n1832 GNDA.n1221 4.26717
R4197 GNDA.n1838 GNDA.n1221 4.26717
R4198 GNDA.n1839 GNDA.n1838 4.26717
R4199 GNDA.n1839 GNDA.n1218 4.26717
R4200 GNDA.n1218 GNDA.n1216 4.26717
R4201 GNDA.n1847 GNDA.n1216 4.26717
R4202 GNDA.n1847 GNDA.n1212 4.26717
R4203 GNDA.n1853 GNDA.n1212 4.26717
R4204 GNDA.n1854 GNDA.n1853 4.26717
R4205 GNDA.n1854 GNDA.n1209 4.26717
R4206 GNDA.n1046 GNDA.n722 4.26717
R4207 GNDA.n1041 GNDA.n722 4.26717
R4208 GNDA.n1041 GNDA.n1040 4.26717
R4209 GNDA.n1040 GNDA.n730 4.26717
R4210 GNDA.n1035 GNDA.n730 4.26717
R4211 GNDA.n1035 GNDA.n1034 4.26717
R4212 GNDA.n1034 GNDA.n1033 4.26717
R4213 GNDA.n1033 GNDA.n738 4.26717
R4214 GNDA.n1027 GNDA.n738 4.26717
R4215 GNDA.n1027 GNDA.n1026 4.26717
R4216 GNDA.n1026 GNDA.n1025 4.26717
R4217 GNDA.n1914 GNDA.n1913 4.26717
R4218 GNDA.n1913 GNDA.n1888 4.26717
R4219 GNDA.n1908 GNDA.n1888 4.26717
R4220 GNDA.n1908 GNDA.n1907 4.26717
R4221 GNDA.n1907 GNDA.n1906 4.26717
R4222 GNDA.n1906 GNDA.n1894 4.26717
R4223 GNDA.n1900 GNDA.n1894 4.26717
R4224 GNDA.n1900 GNDA.n1899 4.26717
R4225 GNDA.n1899 GNDA.n1053 4.26717
R4226 GNDA.n2192 GNDA.n1053 4.26717
R4227 GNDA.n2192 GNDA.n1050 4.26717
R4228 GNDA.n1531 GNDA.n1424 4.26717
R4229 GNDA.n1537 GNDA.n1424 4.26717
R4230 GNDA.n1538 GNDA.n1537 4.26717
R4231 GNDA.n1541 GNDA.n1538 4.26717
R4232 GNDA.n1541 GNDA.n1422 4.26717
R4233 GNDA.n1547 GNDA.n1422 4.26717
R4234 GNDA.n1547 GNDA.n1416 4.26717
R4235 GNDA.n1555 GNDA.n1416 4.26717
R4236 GNDA.n1555 GNDA.n1414 4.26717
R4237 GNDA.n1414 GNDA.n1295 4.26717
R4238 GNDA.n1562 GNDA.n1295 4.26717
R4239 GNDA.n2182 GNDA.n1126 4.26717
R4240 GNDA.n2177 GNDA.n1126 4.26717
R4241 GNDA.n2177 GNDA.n2176 4.26717
R4242 GNDA.n2176 GNDA.n1134 4.26717
R4243 GNDA.n2171 GNDA.n1134 4.26717
R4244 GNDA.n2171 GNDA.n2170 4.26717
R4245 GNDA.n2170 GNDA.n2169 4.26717
R4246 GNDA.n2169 GNDA.n1142 4.26717
R4247 GNDA.n2163 GNDA.n1142 4.26717
R4248 GNDA.n2163 GNDA.n2162 4.26717
R4249 GNDA.n2162 GNDA.n2161 4.26717
R4250 GNDA.n2508 GNDA.n583 4.26717
R4251 GNDA.n2503 GNDA.n583 4.26717
R4252 GNDA.n2503 GNDA.n2502 4.26717
R4253 GNDA.n2502 GNDA.n591 4.26717
R4254 GNDA.n2497 GNDA.n591 4.26717
R4255 GNDA.n2497 GNDA.n2496 4.26717
R4256 GNDA.n2496 GNDA.n2495 4.26717
R4257 GNDA.n2495 GNDA.n599 4.26717
R4258 GNDA.n2489 GNDA.n599 4.26717
R4259 GNDA.n2489 GNDA.n2488 4.26717
R4260 GNDA.n2488 GNDA.n2487 4.26717
R4261 GNDA.n230 GNDA.n217 4.2505
R4262 GNDA.n2599 GNDA.n3 4.21925
R4263 GNDA GNDA.n2602 4.2117
R4264 GNDA.n214 GNDA.n211 4.17148
R4265 GNDA.n215 GNDA.n214 4.17148
R4266 GNDA.n2567 GNDA.n519 4.063
R4267 GNDA.n203 GNDA.n193 4.0593
R4268 GNDA.n466 GNDA.n465 4.0005
R4269 GNDA.n1447 GNDA.n1225 3.93531
R4270 GNDA.n1047 GNDA.n1046 3.93531
R4271 GNDA.n1914 GNDA.n1861 3.93531
R4272 GNDA.n1531 GNDA.n1472 3.93531
R4273 GNDA.n2183 GNDA.n2182 3.93531
R4274 GNDA.n2509 GNDA.n2508 3.93531
R4275 GNDA.t32 GNDA.t271 3.83994
R4276 GNDA.t255 GNDA.t78 3.83994
R4277 GNDA.t24 GNDA.t249 3.83994
R4278 GNDA.t234 GNDA.t143 3.83994
R4279 GNDA.n1651 GNDA.n1650 3.7893
R4280 GNDA.n1647 GNDA.n1270 3.7893
R4281 GNDA.n1646 GNDA.n1273 3.7893
R4282 GNDA.n1643 GNDA.n1642 3.7893
R4283 GNDA.n1569 GNDA.n1274 3.7893
R4284 GNDA.n1578 GNDA.n1577 3.7893
R4285 GNDA.n1581 GNDA.n1568 3.7893
R4286 GNDA.n1586 GNDA.n1582 3.7893
R4287 GNDA.n2457 GNDA.n2456 3.7893
R4288 GNDA.n2453 GNDA.n2320 3.7893
R4289 GNDA.n2452 GNDA.n2323 3.7893
R4290 GNDA.n2330 GNDA.n2329 3.7893
R4291 GNDA.n2446 GNDA.n2445 3.7893
R4292 GNDA.n2375 GNDA.n2374 3.7893
R4293 GNDA.n2379 GNDA.n2378 3.7893
R4294 GNDA.n2387 GNDA.n2350 3.7893
R4295 GNDA.n2265 GNDA.n633 3.7893
R4296 GNDA.n2262 GNDA.n2261 3.7893
R4297 GNDA.n674 GNDA.n635 3.7893
R4298 GNDA.n692 GNDA.n691 3.7893
R4299 GNDA.n689 GNDA.n688 3.7893
R4300 GNDA.n684 GNDA.n677 3.7893
R4301 GNDA.n681 GNDA.n680 3.7893
R4302 GNDA.n2203 GNDA.n655 3.7893
R4303 GNDA.n2154 GNDA.n1152 3.7893
R4304 GNDA.n2151 GNDA.n2150 3.7893
R4305 GNDA.n2067 GNDA.n1153 3.7893
R4306 GNDA.n2072 GNDA.n2070 3.7893
R4307 GNDA.n2077 GNDA.n2073 3.7893
R4308 GNDA.n2084 GNDA.n2083 3.7893
R4309 GNDA.n2087 GNDA.n2066 3.7893
R4310 GNDA.n2092 GNDA.n2088 3.7893
R4311 GNDA.n2059 GNDA.n1173 3.7893
R4312 GNDA.n2056 GNDA.n2055 3.7893
R4313 GNDA.n1972 GNDA.n1174 3.7893
R4314 GNDA.n1977 GNDA.n1975 3.7893
R4315 GNDA.n1982 GNDA.n1978 3.7893
R4316 GNDA.n1989 GNDA.n1988 3.7893
R4317 GNDA.n1992 GNDA.n1971 3.7893
R4318 GNDA.n1997 GNDA.n1993 3.7893
R4319 GNDA.n1734 GNDA.n1671 3.7893
R4320 GNDA.n1743 GNDA.n1742 3.7893
R4321 GNDA.n1668 GNDA.n1667 3.7893
R4322 GNDA.n1751 GNDA.n1749 3.7893
R4323 GNDA.n1750 GNDA.n1665 3.7893
R4324 GNDA.n1663 GNDA.n1662 3.7893
R4325 GNDA.n1766 GNDA.n1764 3.7893
R4326 GNDA.n1765 GNDA.n1658 3.7893
R4327 GNDA.n1408 GNDA.n1297 3.7893
R4328 GNDA.n1405 GNDA.n1404 3.7893
R4329 GNDA.n1321 GNDA.n1298 3.7893
R4330 GNDA.n1326 GNDA.n1324 3.7893
R4331 GNDA.n1331 GNDA.n1327 3.7893
R4332 GNDA.n1338 GNDA.n1337 3.7893
R4333 GNDA.n1341 GNDA.n1320 3.7893
R4334 GNDA.n1346 GNDA.n1342 3.7893
R4335 GNDA.n1012 GNDA.n1011 3.7893
R4336 GNDA.n1008 GNDA.n889 3.7893
R4337 GNDA.n1007 GNDA.n892 3.7893
R4338 GNDA.n897 GNDA.n896 3.7893
R4339 GNDA.n1001 GNDA.n1000 3.7893
R4340 GNDA.n933 GNDA.n932 3.7893
R4341 GNDA.n929 GNDA.n916 3.7893
R4342 GNDA.n941 GNDA.n939 3.7893
R4343 GNDA.n2545 GNDA.n550 3.7893
R4344 GNDA.n2544 GNDA.n551 3.7893
R4345 GNDA.n2532 GNDA.n2531 3.7893
R4346 GNDA.n2538 GNDA.n2537 3.7893
R4347 GNDA.n2534 GNDA.n2533 3.7893
R4348 GNDA.n811 GNDA.n529 3.7893
R4349 GNDA.n814 GNDA.n813 3.7893
R4350 GNDA.n821 GNDA.n747 3.7893
R4351 GNDA.n1574 GNDA 3.7381
R4352 GNDA.n2373 GNDA 3.7381
R4353 GNDA.n685 GNDA 3.7381
R4354 GNDA.n2080 GNDA 3.7381
R4355 GNDA.n1985 GNDA 3.7381
R4356 GNDA GNDA.n1757 3.7381
R4357 GNDA.n1334 GNDA 3.7381
R4358 GNDA.n928 GNDA 3.7381
R4359 GNDA GNDA.n2550 3.7381
R4360 GNDA.n2572 GNDA.n516 3.51962
R4361 GNDA.n88 GNDA.t138 3.42907
R4362 GNDA.n88 GNDA.t326 3.42907
R4363 GNDA.n320 GNDA.t136 3.42907
R4364 GNDA.n320 GNDA.t318 3.42907
R4365 GNDA.n317 GNDA.t314 3.42907
R4366 GNDA.n317 GNDA.t324 3.42907
R4367 GNDA.n91 GNDA.t101 3.42907
R4368 GNDA.n91 GNDA.t305 3.42907
R4369 GNDA.n486 GNDA.n479 3.19754
R4370 GNDA.n481 GNDA.n23 3.19754
R4371 GNDA.n502 GNDA.n20 3.19754
R4372 GNDA.n497 GNDA.n495 3.19754
R4373 GNDA.n376 GNDA.n238 3.19754
R4374 GNDA.n371 GNDA.n369 3.19754
R4375 GNDA.n360 GNDA.n353 3.19754
R4376 GNDA.n355 GNDA.n252 3.19754
R4377 GNDA.n347 GNDA.n262 3.19754
R4378 GNDA.n326 GNDA.n324 3.19754
R4379 GNDA.n287 GNDA.n286 3.19754
R4380 GNDA.n273 GNDA.n272 3.19754
R4381 GNDA.n118 GNDA.n33 3.19754
R4382 GNDA.n97 GNDA.n95 3.19754
R4383 GNDA.n58 GNDA.n57 3.19754
R4384 GNDA.n44 GNDA.n43 3.19754
R4385 GNDA.n2462 GNDA.n2461 3.08966
R4386 GNDA.n2327 GNDA.t105 3.08966
R4387 GNDA.n2369 GNDA.t82 3.08966
R4388 GNDA.n2384 GNDA.t73 3.08966
R4389 GNDA.n2542 GNDA.t92 3.08966
R4390 GNDA.n2560 GNDA.n520 2.86505
R4391 GNDA.n2561 GNDA.n2560 2.86505
R4392 GNDA.n2559 GNDA.n2555 2.86505
R4393 GNDA.n2556 GNDA.n2555 2.86505
R4394 GNDA.n2562 GNDA.n2561 2.86505
R4395 GNDA.n2557 GNDA.n2556 2.86505
R4396 GNDA.n2566 GNDA.n520 2.86505
R4397 GNDA.n2562 GNDA.n2559 2.86505
R4398 GNDA.n221 GNDA.n220 2.86505
R4399 GNDA.n220 GNDA.n219 2.86505
R4400 GNDA.n227 GNDA.n219 2.86505
R4401 GNDA.n223 GNDA.n221 2.86505
R4402 GNDA.n145 GNDA.n144 2.86505
R4403 GNDA.n400 GNDA.n145 2.86505
R4404 GNDA.n400 GNDA.n399 2.86505
R4405 GNDA.n402 GNDA.n144 2.86505
R4406 GNDA.n2362 GNDA.n2358 2.86505
R4407 GNDA.n2363 GNDA.n2362 2.86505
R4408 GNDA.n2364 GNDA.n2363 2.86505
R4409 GNDA.n2359 GNDA.n2358 2.86505
R4410 GNDA.n1653 GNDA.n1652 2.6629
R4411 GNDA.n1566 GNDA.n1293 2.6629
R4412 GNDA.n2459 GNDA.n2458 2.6629
R4413 GNDA.n2348 GNDA.n607 2.6629
R4414 GNDA.n2267 GNDA.n2266 2.6629
R4415 GNDA.n2158 GNDA.n1150 2.6629
R4416 GNDA.n2157 GNDA.n2155 2.6629
R4417 GNDA.n2064 GNDA.n2062 2.6629
R4418 GNDA.n2061 GNDA.n2060 2.6629
R4419 GNDA.n1735 GNDA.n1733 2.6629
R4420 GNDA.n1410 GNDA.n1409 2.6629
R4421 GNDA.n1318 GNDA.n1204 2.6629
R4422 GNDA.n888 GNDA.n887 2.6629
R4423 GNDA.n880 GNDA.n878 2.6629
R4424 GNDA.n877 GNDA.n876 2.6629
R4425 GNDA.n209 GNDA.n208 2.53175
R4426 GNDA.n124 GNDA.n22 2.46925
R4427 GNDA.n1567 GNDA.n1566 2.4581
R4428 GNDA.n2349 GNDA.n2348 2.4581
R4429 GNDA.n1150 GNDA.n654 2.4581
R4430 GNDA.n2158 GNDA.n2157 2.4581
R4431 GNDA.n2065 GNDA.n2064 2.4581
R4432 GNDA.n2062 GNDA.n2061 2.4581
R4433 GNDA.n1970 GNDA.n1969 2.4581
R4434 GNDA.n1733 GNDA.n1204 2.4581
R4435 GNDA.n1772 GNDA.n1251 2.4581
R4436 GNDA.n1410 GNDA.n1293 2.4581
R4437 GNDA.n1319 GNDA.n1318 2.4581
R4438 GNDA.n887 GNDA.n607 2.4581
R4439 GNDA.n915 GNDA.n880 2.4581
R4440 GNDA.n878 GNDA.n877 2.4581
R4441 GNDA.n808 GNDA.n746 2.4581
R4442 GNDA.n465 GNDA.n125 2.2505
R4443 GNDA.n2585 GNDA.n6 2.20408
R4444 GNDA.n1209 GNDA.n1204 2.18124
R4445 GNDA.n1025 GNDA.n878 2.18124
R4446 GNDA.n2062 GNDA.n1050 2.18124
R4447 GNDA.n1562 GNDA.n1293 2.18124
R4448 GNDA.n2161 GNDA.n2158 2.18124
R4449 GNDA.n2487 GNDA.n607 2.18124
R4450 GNDA.n1585 GNDA.n1567 2.1509
R4451 GNDA.n2386 GNDA.n2349 2.1509
R4452 GNDA.n2202 GNDA.n654 2.1509
R4453 GNDA.n2091 GNDA.n2065 2.1509
R4454 GNDA.n1996 GNDA.n1970 2.1509
R4455 GNDA.n1773 GNDA.n1772 2.1509
R4456 GNDA.n1345 GNDA.n1319 2.1509
R4457 GNDA.n940 GNDA.n915 2.1509
R4458 GNDA.n820 GNDA.n746 2.1509
R4459 GNDA.n1652 GNDA.n1268 2.13383
R4460 GNDA.n2458 GNDA.n2319 2.13383
R4461 GNDA.n2266 GNDA.n632 2.13383
R4462 GNDA.n2155 GNDA.n1151 2.13383
R4463 GNDA.n2060 GNDA.n1172 2.13383
R4464 GNDA.n1409 GNDA.n1296 2.13383
R4465 GNDA.n1736 GNDA.n1735 2.13383
R4466 GNDA.n980 GNDA.n888 2.13383
R4467 GNDA.n876 GNDA.n875 2.13383
R4468 GNDA.n426 GNDA.n124 2.1255
R4469 GNDA.n2568 GNDA 2.09787
R4470 GNDA.n1860 GNDA.n1204 2.08643
R4471 GNDA.n1021 GNDA.n878 2.08643
R4472 GNDA.n2062 GNDA.n1048 2.08643
R4473 GNDA.n1293 GNDA.n1125 2.08643
R4474 GNDA.n2158 GNDA.n582 2.08643
R4475 GNDA.n610 GNDA.n607 2.08643
R4476 GNDA.n2384 GNDA.t266 2.05994
R4477 GNDA.n884 GNDA.t287 2.05994
R4478 GNDA.n1018 GNDA.t243 2.05994
R4479 GNDA.n2527 GNDA.t263 2.05994
R4480 GNDA.n1652 GNDA.n1651 1.9461
R4481 GNDA.n2458 GNDA.n2457 1.9461
R4482 GNDA.n2266 GNDA.n2265 1.9461
R4483 GNDA.n2155 GNDA.n2154 1.9461
R4484 GNDA.n2060 GNDA.n2059 1.9461
R4485 GNDA.n1735 GNDA.n1734 1.9461
R4486 GNDA.n1409 GNDA.n1408 1.9461
R4487 GNDA.n1012 GNDA.n888 1.9461
R4488 GNDA.n876 GNDA.n550 1.9461
R4489 GNDA.n2600 GNDA.n2599 1.938
R4490 GNDA.n1438 GNDA.n1437 1.90675
R4491 GNDA.t131 GNDA.n615 1.83728
R4492 GNDA.n397 GNDA.n230 1.7505
R4493 GNDA.n1485 GNDA.n1267 1.47392
R4494 GNDA.n2318 GNDA.n613 1.47392
R4495 GNDA.n1081 GNDA.n631 1.47392
R4496 GNDA.n1962 GNDA.n1193 1.47392
R4497 GNDA.n1783 GNDA.n1782 1.47392
R4498 GNDA.n807 GNDA.n806 1.47392
R4499 GNDA.n209 GNDA.n22 1.32862
R4500 GNDA.n2522 GNDA.n2517 0.96925
R4501 GNDA.n2480 GNDA.n2479 0.96925
R4502 GNDA.n1650 GNDA.n1270 0.8197
R4503 GNDA.n1647 GNDA.n1646 0.8197
R4504 GNDA.n1643 GNDA.n1273 0.8197
R4505 GNDA.n1642 GNDA.n1274 0.8197
R4506 GNDA.n1577 GNDA.n1574 0.8197
R4507 GNDA.n1578 GNDA.n1568 0.8197
R4508 GNDA.n1582 GNDA.n1581 0.8197
R4509 GNDA.n1586 GNDA.n1585 0.8197
R4510 GNDA.n2456 GNDA.n2320 0.8197
R4511 GNDA.n2453 GNDA.n2452 0.8197
R4512 GNDA.n2329 GNDA.n2323 0.8197
R4513 GNDA.n2446 GNDA.n2330 0.8197
R4514 GNDA.n2374 GNDA.n2373 0.8197
R4515 GNDA.n2379 GNDA.n2375 0.8197
R4516 GNDA.n2378 GNDA.n2350 0.8197
R4517 GNDA.n2387 GNDA.n2386 0.8197
R4518 GNDA.n2262 GNDA.n633 0.8197
R4519 GNDA.n2261 GNDA.n635 0.8197
R4520 GNDA.n692 GNDA.n674 0.8197
R4521 GNDA.n691 GNDA.n689 0.8197
R4522 GNDA.n685 GNDA.n684 0.8197
R4523 GNDA.n681 GNDA.n677 0.8197
R4524 GNDA.n680 GNDA.n655 0.8197
R4525 GNDA.n2203 GNDA.n2202 0.8197
R4526 GNDA.n2151 GNDA.n1152 0.8197
R4527 GNDA.n2150 GNDA.n1153 0.8197
R4528 GNDA.n2070 GNDA.n2067 0.8197
R4529 GNDA.n2073 GNDA.n2072 0.8197
R4530 GNDA.n2083 GNDA.n2080 0.8197
R4531 GNDA.n2084 GNDA.n2066 0.8197
R4532 GNDA.n2088 GNDA.n2087 0.8197
R4533 GNDA.n2092 GNDA.n2091 0.8197
R4534 GNDA.n2056 GNDA.n1173 0.8197
R4535 GNDA.n2055 GNDA.n1174 0.8197
R4536 GNDA.n1975 GNDA.n1972 0.8197
R4537 GNDA.n1978 GNDA.n1977 0.8197
R4538 GNDA.n1988 GNDA.n1985 0.8197
R4539 GNDA.n1989 GNDA.n1971 0.8197
R4540 GNDA.n1993 GNDA.n1992 0.8197
R4541 GNDA.n1997 GNDA.n1996 0.8197
R4542 GNDA.n1743 GNDA.n1671 0.8197
R4543 GNDA.n1742 GNDA.n1668 0.8197
R4544 GNDA.n1749 GNDA.n1667 0.8197
R4545 GNDA.n1751 GNDA.n1750 0.8197
R4546 GNDA.n1757 GNDA.n1663 0.8197
R4547 GNDA.n1764 GNDA.n1662 0.8197
R4548 GNDA.n1766 GNDA.n1765 0.8197
R4549 GNDA.n1773 GNDA.n1658 0.8197
R4550 GNDA.n1405 GNDA.n1297 0.8197
R4551 GNDA.n1404 GNDA.n1298 0.8197
R4552 GNDA.n1324 GNDA.n1321 0.8197
R4553 GNDA.n1327 GNDA.n1326 0.8197
R4554 GNDA.n1337 GNDA.n1334 0.8197
R4555 GNDA.n1338 GNDA.n1320 0.8197
R4556 GNDA.n1342 GNDA.n1341 0.8197
R4557 GNDA.n1346 GNDA.n1345 0.8197
R4558 GNDA.n1011 GNDA.n889 0.8197
R4559 GNDA.n1008 GNDA.n1007 0.8197
R4560 GNDA.n896 GNDA.n892 0.8197
R4561 GNDA.n1001 GNDA.n897 0.8197
R4562 GNDA.n933 GNDA.n928 0.8197
R4563 GNDA.n932 GNDA.n929 0.8197
R4564 GNDA.n939 GNDA.n916 0.8197
R4565 GNDA.n941 GNDA.n940 0.8197
R4566 GNDA.n2545 GNDA.n2544 0.8197
R4567 GNDA.n2531 GNDA.n551 0.8197
R4568 GNDA.n2538 GNDA.n2532 0.8197
R4569 GNDA.n2537 GNDA.n2534 0.8197
R4570 GNDA.n2550 GNDA.n529 0.8197
R4571 GNDA.n814 GNDA.n811 0.8197
R4572 GNDA.n813 GNDA.n747 0.8197
R4573 GNDA.n821 GNDA.n820 0.8197
R4574 GNDA.n443 GNDA.n441 0.604667
R4575 GNDA.t50 GNDA.t211 0.586152
R4576 GNDA.n2315 GNDA.n615 0.575776
R4577 GNDA GNDA.n1569 0.5637
R4578 GNDA.n2445 GNDA 0.5637
R4579 GNDA.n688 GNDA 0.5637
R4580 GNDA.n2077 GNDA 0.5637
R4581 GNDA.n1982 GNDA 0.5637
R4582 GNDA.n1665 GNDA 0.5637
R4583 GNDA.n1331 GNDA 0.5637
R4584 GNDA.n1000 GNDA 0.5637
R4585 GNDA.n2533 GNDA 0.5637
R4586 GNDA.n2573 GNDA.n515 0.563
R4587 GNDA.n2519 GNDA.n515 0.563
R4588 GNDA.n2521 GNDA.n2519 0.563
R4589 GNDA.n2522 GNDA.n2521 0.563
R4590 GNDA.n2517 GNDA.n555 0.563
R4591 GNDA.n2472 GNDA.n555 0.563
R4592 GNDA.n2474 GNDA.n2472 0.563
R4593 GNDA.n2476 GNDA.n2474 0.563
R4594 GNDA.n2479 GNDA.n2476 0.563
R4595 GNDA.n2480 GNDA.n2470 0.563
R4596 GNDA.n2470 GNDA.n2468 0.563
R4597 GNDA.n2468 GNDA.n2466 0.563
R4598 GNDA.n165 GNDA.n163 0.563
R4599 GNDA.n167 GNDA.n165 0.563
R4600 GNDA.n169 GNDA.n167 0.563
R4601 GNDA.n171 GNDA.n169 0.563
R4602 GNDA.n173 GNDA.n171 0.563
R4603 GNDA.n175 GNDA.n173 0.563
R4604 GNDA.n177 GNDA.n175 0.563
R4605 GNDA.n179 GNDA.n177 0.563
R4606 GNDA.n181 GNDA.n179 0.563
R4607 GNDA.n183 GNDA.n181 0.563
R4608 GNDA.n207 GNDA.n183 0.563
R4609 GNDA.n419 GNDA.n417 0.563
R4610 GNDA.n421 GNDA.n419 0.563
R4611 GNDA.n423 GNDA.n421 0.563
R4612 GNDA.n244 GNDA.n242 0.563
R4613 GNDA.n246 GNDA.n244 0.563
R4614 GNDA.n248 GNDA.n246 0.563
R4615 GNDA.n321 GNDA.n319 0.5005
R4616 GNDA.n319 GNDA.n318 0.5005
R4617 GNDA.n92 GNDA.n90 0.5005
R4618 GNDA.n90 GNDA.n89 0.5005
R4619 GNDA.n2571 GNDA.n2568 0.276625
R4620 GNDA.n1572 GNDA 0.2565
R4621 GNDA.n2372 GNDA 0.2565
R4622 GNDA.n676 GNDA 0.2565
R4623 GNDA GNDA.n2076 0.2565
R4624 GNDA GNDA.n1981 0.2565
R4625 GNDA.n1758 GNDA 0.2565
R4626 GNDA GNDA.n1330 0.2565
R4627 GNDA.n927 GNDA 0.2565
R4628 GNDA.n2551 GNDA 0.2565
R4629 GNDA.n2572 GNDA.n2571 0.22375
R4630 GNDA GNDA.n1572 0.0517
R4631 GNDA GNDA.n2372 0.0517
R4632 GNDA GNDA.n676 0.0517
R4633 GNDA.n2076 GNDA 0.0517
R4634 GNDA.n1981 GNDA 0.0517
R4635 GNDA.n1758 GNDA 0.0517
R4636 GNDA.n1330 GNDA 0.0517
R4637 GNDA GNDA.n927 0.0517
R4638 GNDA.n2551 GNDA 0.0517
R4639 VDDA.n345 VDDA.t295 1212.4
R4640 VDDA.n409 VDDA.t271 1212.4
R4641 VDDA.n105 VDDA.t311 1212.4
R4642 VDDA.n174 VDDA.t326 1212.4
R4643 VDDA.n418 VDDA.t300 905.125
R4644 VDDA.n417 VDDA.t310 905.125
R4645 VDDA.n202 VDDA.t289 794.668
R4646 VDDA.n206 VDDA.t286 794.668
R4647 VDDA.n186 VDDA.t368 794.668
R4648 VDDA.n231 VDDA.t341 794.668
R4649 VDDA.n526 VDDA.t340 708.125
R4650 VDDA.t340 VDDA.n482 708.125
R4651 VDDA.n503 VDDA.t282 708.125
R4652 VDDA.t282 VDDA.n485 708.125
R4653 VDDA.n415 VDDA.n414 682
R4654 VDDA.n548 VDDA.t375 676.966
R4655 VDDA.n418 VDDA.t299 672.274
R4656 VDDA.t308 VDDA.n417 672.274
R4657 VDDA.n505 VDDA.t305 660.001
R4658 VDDA.t339 VDDA.n527 657.76
R4659 VDDA.t281 VDDA.n504 657.76
R4660 VDDA.n430 VDDA.t329 652.076
R4661 VDDA.n464 VDDA.t356 652.076
R4662 VDDA.n246 VDDA.t292 652.076
R4663 VDDA.n279 VDDA.t362 652.076
R4664 VDDA.n11 VDDA.t323 652.076
R4665 VDDA.n44 VDDA.t277 652.076
R4666 VDDA.t366 VDDA.n625 645.231
R4667 VDDA.n626 VDDA.t345 645.231
R4668 VDDA.t318 VDDA.n594 643.038
R4669 VDDA.t336 VDDA.n547 643.038
R4670 VDDA.n595 VDDA.t315 643.038
R4671 VDDA.t284 VDDA.n633 643.037
R4672 VDDA.n634 VDDA.t360 643.037
R4673 VDDA.t351 VDDA.n611 643.037
R4674 VDDA.n612 VDDA.t275 643.037
R4675 VDDA.n309 VDDA.t347 624.725
R4676 VDDA.n72 VDDA.t353 624.725
R4677 VDDA.n319 VDDA.t332 601.867
R4678 VDDA.n84 VDDA.t371 601.867
R4679 VDDA.n380 VDDA.n323 587.407
R4680 VDDA.n388 VDDA.n387 587.407
R4681 VDDA.n374 VDDA.n373 587.407
R4682 VDDA.n354 VDDA.n353 587.407
R4683 VDDA.n134 VDDA.n106 587.407
R4684 VDDA.n119 VDDA.n115 587.407
R4685 VDDA.n145 VDDA.n88 587.407
R4686 VDDA.n153 VDDA.n152 587.407
R4687 VDDA.n573 VDDA.n541 587.407
R4688 VDDA.n569 VDDA.n568 587.407
R4689 VDDA.n586 VDDA.n585 587.407
R4690 VDDA.n580 VDDA.n535 587.407
R4691 VDDA.n463 VDDA.n423 585
R4692 VDDA.n445 VDDA.n444 585
R4693 VDDA.n404 VDDA.n380 585
R4694 VDDA.n403 VDDA.n381 585
R4695 VDDA.n402 VDDA.n382 585
R4696 VDDA.n399 VDDA.n383 585
R4697 VDDA.n398 VDDA.n384 585
R4698 VDDA.n395 VDDA.n385 585
R4699 VDDA.n394 VDDA.n386 585
R4700 VDDA.n391 VDDA.n387 585
R4701 VDDA.n373 VDDA.n372 585
R4702 VDDA.n369 VDDA.n347 585
R4703 VDDA.n368 VDDA.n348 585
R4704 VDDA.n365 VDDA.n349 585
R4705 VDDA.n364 VDDA.n350 585
R4706 VDDA.n361 VDDA.n351 585
R4707 VDDA.n360 VDDA.n352 585
R4708 VDDA.n357 VDDA.n353 585
R4709 VDDA.n278 VDDA.n237 585
R4710 VDDA.n260 VDDA.n259 585
R4711 VDDA.n219 VDDA.n218 585
R4712 VDDA.n216 VDDA.n215 585
R4713 VDDA.n230 VDDA.n179 585
R4714 VDDA.n201 VDDA.n188 585
R4715 VDDA.n169 VDDA.n145 585
R4716 VDDA.n168 VDDA.n146 585
R4717 VDDA.n167 VDDA.n147 585
R4718 VDDA.n164 VDDA.n148 585
R4719 VDDA.n163 VDDA.n149 585
R4720 VDDA.n160 VDDA.n150 585
R4721 VDDA.n159 VDDA.n151 585
R4722 VDDA.n156 VDDA.n152 585
R4723 VDDA.n132 VDDA.n106 585
R4724 VDDA.n131 VDDA.n130 585
R4725 VDDA.n129 VDDA.n109 585
R4726 VDDA.n128 VDDA.n127 585
R4727 VDDA.n126 VDDA.n125 585
R4728 VDDA.n124 VDDA.n114 585
R4729 VDDA.n123 VDDA.n122 585
R4730 VDDA.n121 VDDA.n115 585
R4731 VDDA.n43 VDDA.n2 585
R4732 VDDA.n25 VDDA.n24 585
R4733 VDDA.n585 VDDA.n584 585
R4734 VDDA.n583 VDDA.n580 585
R4735 VDDA.n571 VDDA.n541 585
R4736 VDDA.n570 VDDA.n569 585
R4737 VDDA.n528 VDDA.t321 540.818
R4738 VDDA.n317 VDDA.t334 464.281
R4739 VDDA.n314 VDDA.t334 464.281
R4740 VDDA.n308 VDDA.t349 464.281
R4741 VDDA.t349 VDDA.n307 464.281
R4742 VDDA.n71 VDDA.t355 464.281
R4743 VDDA.t355 VDDA.n70 464.281
R4744 VDDA.t373 VDDA.n63 464.281
R4745 VDDA.n79 VDDA.t373 464.281
R4746 VDDA.n416 VDDA.t307 447.226
R4747 VDDA.n419 VDDA.t298 447.226
R4748 VDDA.n593 VDDA.t317 419.108
R4749 VDDA.n596 VDDA.t314 419.108
R4750 VDDA.n546 VDDA.t335 413.084
R4751 VDDA.n549 VDDA.t374 413.084
R4752 VDDA.n632 VDDA.t283 409.067
R4753 VDDA.n635 VDDA.t359 409.067
R4754 VDDA.n624 VDDA.t365 409.067
R4755 VDDA.n627 VDDA.t344 409.067
R4756 VDDA.n610 VDDA.t350 409.067
R4757 VDDA.t403 VDDA.t339 407.144
R4758 VDDA.t57 VDDA.t403 407.144
R4759 VDDA.t4 VDDA.t57 407.144
R4760 VDDA.t196 VDDA.t4 407.144
R4761 VDDA.t219 VDDA.t196 407.144
R4762 VDDA.t405 VDDA.t219 407.144
R4763 VDDA.t110 VDDA.t405 407.144
R4764 VDDA.t170 VDDA.t110 407.144
R4765 VDDA.t8 VDDA.t170 407.144
R4766 VDDA.t30 VDDA.t8 407.144
R4767 VDDA.t44 VDDA.t30 407.144
R4768 VDDA.t410 VDDA.t44 407.144
R4769 VDDA.t19 VDDA.t410 407.144
R4770 VDDA.t122 VDDA.t19 407.144
R4771 VDDA.t124 VDDA.t122 407.144
R4772 VDDA.t10 VDDA.t124 407.144
R4773 VDDA.t87 VDDA.t10 407.144
R4774 VDDA.t17 VDDA.t87 407.144
R4775 VDDA.t321 VDDA.t17 407.144
R4776 VDDA.t136 VDDA.t281 407.144
R4777 VDDA.t138 VDDA.t136 407.144
R4778 VDDA.t24 VDDA.t138 407.144
R4779 VDDA.t2 VDDA.t24 407.144
R4780 VDDA.t176 VDDA.t2 407.144
R4781 VDDA.t178 VDDA.t176 407.144
R4782 VDDA.t401 VDDA.t178 407.144
R4783 VDDA.t15 VDDA.t401 407.144
R4784 VDDA.t128 VDDA.t15 407.144
R4785 VDDA.t82 VDDA.t128 407.144
R4786 VDDA.t0 VDDA.t82 407.144
R4787 VDDA.t180 VDDA.t0 407.144
R4788 VDDA.t389 VDDA.t180 407.144
R4789 VDDA.t80 VDDA.t389 407.144
R4790 VDDA.t391 VDDA.t80 407.144
R4791 VDDA.t184 VDDA.t391 407.144
R4792 VDDA.t182 VDDA.t184 407.144
R4793 VDDA.t78 VDDA.t182 407.144
R4794 VDDA.t305 VDDA.t78 407.144
R4795 VDDA.n613 VDDA.t274 390.322
R4796 VDDA.n526 VDDA.t338 379.582
R4797 VDDA.n503 VDDA.t280 379.582
R4798 VDDA.t320 VDDA.n529 379.277
R4799 VDDA.t84 VDDA.t318 373.214
R4800 VDDA.t174 VDDA.t84 373.214
R4801 VDDA.t315 VDDA.t174 373.214
R4802 VDDA.t55 VDDA.t336 373.214
R4803 VDDA.t127 VDDA.t55 373.214
R4804 VDDA.t375 VDDA.t127 373.214
R4805 VDDA.t215 VDDA.t284 373.214
R4806 VDDA.t6 VDDA.t215 373.214
R4807 VDDA.t53 VDDA.t6 373.214
R4808 VDDA.t66 VDDA.t53 373.214
R4809 VDDA.t360 VDDA.t66 373.214
R4810 VDDA.t64 VDDA.t366 373.214
R4811 VDDA.t395 VDDA.t64 373.214
R4812 VDDA.t217 VDDA.t395 373.214
R4813 VDDA.t32 VDDA.t217 373.214
R4814 VDDA.t397 VDDA.t32 373.214
R4815 VDDA.t46 VDDA.t397 373.214
R4816 VDDA.t198 VDDA.t46 373.214
R4817 VDDA.t118 VDDA.t198 373.214
R4818 VDDA.t194 VDDA.t118 373.214
R4819 VDDA.t190 VDDA.t194 373.214
R4820 VDDA.t345 VDDA.t190 373.214
R4821 VDDA.t210 VDDA.t351 373.214
R4822 VDDA.t192 VDDA.t210 373.214
R4823 VDDA.t172 VDDA.t192 373.214
R4824 VDDA.t120 VDDA.t172 373.214
R4825 VDDA.t275 VDDA.t120 373.214
R4826 VDDA.n566 VDDA.t301 360.868
R4827 VDDA.n591 VDDA.t268 360.868
R4828 VDDA.n530 VDDA.t320 358.858
R4829 VDDA.t338 VDDA.n525 358.858
R4830 VDDA.n506 VDDA.t304 358.858
R4831 VDDA.t280 VDDA.n502 358.858
R4832 VDDA.n625 VDDA.t367 354.154
R4833 VDDA.n626 VDDA.t346 354.154
R4834 VDDA.n505 VDDA.t306 354.065
R4835 VDDA.n595 VDDA.t316 354.065
R4836 VDDA.n594 VDDA.t319 354.063
R4837 VDDA.n547 VDDA.t337 354.063
R4838 VDDA.n481 VDDA.t322 351.793
R4839 VDDA.n548 VDDA.t376 347.224
R4840 VDDA.n607 VDDA.n606 345.127
R4841 VDDA.n609 VDDA.n608 345.127
R4842 VDDA.n603 VDDA.n602 344.7
R4843 VDDA.n630 VDDA.n629 344.7
R4844 VDDA.n479 VDDA.n478 341.675
R4845 VDDA.n509 VDDA.n508 341.675
R4846 VDDA.n511 VDDA.n510 341.675
R4847 VDDA.n513 VDDA.n512 341.675
R4848 VDDA.n515 VDDA.n514 341.675
R4849 VDDA.n517 VDDA.n516 341.675
R4850 VDDA.n519 VDDA.n518 341.675
R4851 VDDA.n521 VDDA.n520 341.675
R4852 VDDA.n523 VDDA.n522 341.675
R4853 VDDA.n484 VDDA.n483 341.675
R4854 VDDA.n487 VDDA.n486 341.675
R4855 VDDA.n489 VDDA.n488 341.675
R4856 VDDA.n491 VDDA.n490 341.675
R4857 VDDA.n493 VDDA.n492 341.675
R4858 VDDA.n495 VDDA.n494 341.675
R4859 VDDA.n497 VDDA.n496 341.675
R4860 VDDA.n499 VDDA.n498 341.675
R4861 VDDA.n501 VDDA.n500 341.675
R4862 VDDA.n605 VDDA.n604 339.272
R4863 VDDA.n616 VDDA.n615 339.272
R4864 VDDA.n618 VDDA.n617 339.272
R4865 VDDA.n620 VDDA.n619 339.272
R4866 VDDA.n622 VDDA.n621 339.272
R4867 VDDA.n599 VDDA.n598 334.772
R4868 VDDA.n611 VDDA.t352 332.267
R4869 VDDA.n612 VDDA.t276 332.267
R4870 VDDA.n633 VDDA.t285 332.084
R4871 VDDA.n634 VDDA.t361 332.084
R4872 VDDA.n218 VDDA.n210 291.053
R4873 VDDA.n218 VDDA.n217 291.053
R4874 VDDA.n215 VDDA.n208 291.053
R4875 VDDA.n215 VDDA.n214 291.053
R4876 VDDA.n451 VDDA.n423 290.233
R4877 VDDA.n457 VDDA.n423 290.233
R4878 VDDA.n452 VDDA.n423 290.233
R4879 VDDA.n444 VDDA.n432 290.233
R4880 VDDA.n444 VDDA.n437 290.233
R4881 VDDA.n444 VDDA.n442 290.233
R4882 VDDA.n266 VDDA.n237 290.233
R4883 VDDA.n272 VDDA.n237 290.233
R4884 VDDA.n267 VDDA.n237 290.233
R4885 VDDA.n259 VDDA.n248 290.233
R4886 VDDA.n259 VDDA.n253 290.233
R4887 VDDA.n259 VDDA.n258 290.233
R4888 VDDA.n223 VDDA.n179 290.233
R4889 VDDA.n224 VDDA.n179 290.233
R4890 VDDA.n193 VDDA.n188 290.233
R4891 VDDA.n197 VDDA.n188 290.233
R4892 VDDA.n31 VDDA.n2 290.233
R4893 VDDA.n37 VDDA.n2 290.233
R4894 VDDA.n32 VDDA.n2 290.233
R4895 VDDA.n24 VDDA.n13 290.233
R4896 VDDA.n24 VDDA.n18 290.233
R4897 VDDA.n24 VDDA.n23 290.233
R4898 VDDA.n312 VDDA.t333 267.188
R4899 VDDA.t348 VDDA.n311 267.188
R4900 VDDA.t354 VDDA.n74 267.188
R4901 VDDA.n81 VDDA.t372 267.188
R4902 VDDA.t299 VDDA.t407 259.091
R4903 VDDA.t407 VDDA.t308 259.091
R4904 VDDA.t144 VDDA.t302 251.471
R4905 VDDA.t160 VDDA.t144 251.471
R4906 VDDA.t186 VDDA.t160 251.471
R4907 VDDA.t35 VDDA.t186 251.471
R4908 VDDA.t101 VDDA.t35 251.471
R4909 VDDA.t207 VDDA.t101 251.471
R4910 VDDA.t140 VDDA.t207 251.471
R4911 VDDA.t116 VDDA.t140 251.471
R4912 VDDA.t103 VDDA.t116 251.471
R4913 VDDA.t142 VDDA.t103 251.471
R4914 VDDA.t59 VDDA.t142 251.471
R4915 VDDA.t61 VDDA.t59 251.471
R4916 VDDA.t112 VDDA.t61 251.471
R4917 VDDA.t105 VDDA.t112 251.471
R4918 VDDA.t204 VDDA.t105 251.471
R4919 VDDA.t97 VDDA.t204 251.471
R4920 VDDA.t269 VDDA.t97 251.471
R4921 VDDA.n381 VDDA.n380 246.25
R4922 VDDA.n382 VDDA.n381 246.25
R4923 VDDA.n383 VDDA.n382 246.25
R4924 VDDA.n385 VDDA.n384 246.25
R4925 VDDA.n386 VDDA.n385 246.25
R4926 VDDA.n387 VDDA.n386 246.25
R4927 VDDA.n373 VDDA.n347 246.25
R4928 VDDA.n348 VDDA.n347 246.25
R4929 VDDA.n349 VDDA.n348 246.25
R4930 VDDA.n351 VDDA.n350 246.25
R4931 VDDA.n352 VDDA.n351 246.25
R4932 VDDA.n353 VDDA.n352 246.25
R4933 VDDA.n130 VDDA.n106 246.25
R4934 VDDA.n130 VDDA.n129 246.25
R4935 VDDA.n129 VDDA.n128 246.25
R4936 VDDA.n125 VDDA.n124 246.25
R4937 VDDA.n124 VDDA.n123 246.25
R4938 VDDA.n123 VDDA.n115 246.25
R4939 VDDA.n146 VDDA.n145 246.25
R4940 VDDA.n147 VDDA.n146 246.25
R4941 VDDA.n148 VDDA.n147 246.25
R4942 VDDA.n150 VDDA.n149 246.25
R4943 VDDA.n151 VDDA.n150 246.25
R4944 VDDA.n152 VDDA.n151 246.25
R4945 VDDA.n307 VDDA.n302 243.698
R4946 VDDA.n70 VDDA.n65 243.698
R4947 VDDA.n587 VDDA.n586 243.698
R4948 VDDA.n452 VDDA.n449 242.903
R4949 VDDA.n442 VDDA.n428 242.903
R4950 VDDA.n267 VDDA.n264 242.903
R4951 VDDA.n258 VDDA.n242 242.903
R4952 VDDA.n224 VDDA.n182 242.903
R4953 VDDA.n198 VDDA.n197 242.903
R4954 VDDA.n32 VDDA.n29 242.903
R4955 VDDA.n23 VDDA.n7 242.903
R4956 VDDA.n463 VDDA.n462 238.367
R4957 VDDA.n408 VDDA.n407 238.367
R4958 VDDA.n310 VDDA.n309 238.367
R4959 VDDA.n278 VDDA.n277 238.367
R4960 VDDA.n220 VDDA.n219 238.367
R4961 VDDA.n230 VDDA.n229 238.367
R4962 VDDA.n216 VDDA.n183 238.367
R4963 VDDA.n173 VDDA.n172 238.367
R4964 VDDA.n73 VDDA.n72 238.367
R4965 VDDA.n43 VDDA.n42 238.367
R4966 VDDA.n529 VDDA.n528 238.367
R4967 VDDA.n528 VDDA.n480 238.367
R4968 VDDA.t302 VDDA.n575 237.5
R4969 VDDA.n588 VDDA.t269 237.5
R4970 VDDA.n228 VDDA.t342 221.121
R4971 VDDA.t369 VDDA.n221 221.121
R4972 VDDA.n221 VDDA.t287 221.121
R4973 VDDA.n199 VDDA.t290 221.121
R4974 VDDA.t333 VDDA.t214 217.708
R4975 VDDA.t214 VDDA.t86 217.708
R4976 VDDA.t86 VDDA.t166 217.708
R4977 VDDA.t166 VDDA.t126 217.708
R4978 VDDA.t126 VDDA.t412 217.708
R4979 VDDA.t412 VDDA.t399 217.708
R4980 VDDA.t399 VDDA.t69 217.708
R4981 VDDA.t69 VDDA.t167 217.708
R4982 VDDA.t167 VDDA.t377 217.708
R4983 VDDA.t377 VDDA.t12 217.708
R4984 VDDA.t12 VDDA.t348 217.708
R4985 VDDA.t91 VDDA.t354 217.708
R4986 VDDA.t75 VDDA.t91 217.708
R4987 VDDA.t156 VDDA.t75 217.708
R4988 VDDA.t74 VDDA.t156 217.708
R4989 VDDA.t70 VDDA.t74 217.708
R4990 VDDA.t14 VDDA.t70 217.708
R4991 VDDA.t209 VDDA.t14 217.708
R4992 VDDA.t130 VDDA.t209 217.708
R4993 VDDA.t147 VDDA.t130 217.708
R4994 VDDA.t90 VDDA.t147 217.708
R4995 VDDA.t372 VDDA.t90 217.708
R4996 VDDA.n178 VDDA.n177 213.186
R4997 VDDA.n204 VDDA.n203 213.186
R4998 VDDA.n388 VDDA.n329 190.333
R4999 VDDA.n354 VDDA.n335 190.333
R5000 VDDA.n314 VDDA.n313 190.333
R5001 VDDA.n153 VDDA.n142 190.333
R5002 VDDA.n119 VDDA.n95 190.333
R5003 VDDA.n80 VDDA.n79 190.333
R5004 VDDA.n574 VDDA.n573 190.333
R5005 VDDA.n425 VDDA.n424 185
R5006 VDDA.n460 VDDA.n459 185
R5007 VDDA.n461 VDDA.n460 185
R5008 VDDA.n458 VDDA.n450 185
R5009 VDDA.n456 VDDA.n455 185
R5010 VDDA.n454 VDDA.n453 185
R5011 VDDA.n446 VDDA.n445 185
R5012 VDDA.n447 VDDA.n446 185
R5013 VDDA.n431 VDDA.n429 185
R5014 VDDA.n434 VDDA.n433 185
R5015 VDDA.n436 VDDA.n435 185
R5016 VDDA.n439 VDDA.n438 185
R5017 VDDA.n441 VDDA.n440 185
R5018 VDDA.n379 VDDA.n324 185
R5019 VDDA.n405 VDDA.n404 185
R5020 VDDA.n406 VDDA.n405 185
R5021 VDDA.n403 VDDA.n378 185
R5022 VDDA.n402 VDDA.n401 185
R5023 VDDA.n400 VDDA.n399 185
R5024 VDDA.n398 VDDA.n397 185
R5025 VDDA.n396 VDDA.n395 185
R5026 VDDA.n394 VDDA.n393 185
R5027 VDDA.n392 VDDA.n391 185
R5028 VDDA.n390 VDDA.n389 185
R5029 VDDA.n406 VDDA.n329 185
R5030 VDDA.n376 VDDA.n375 185
R5031 VDDA.n377 VDDA.n376 185
R5032 VDDA.n346 VDDA.n336 185
R5033 VDDA.n372 VDDA.n371 185
R5034 VDDA.n370 VDDA.n369 185
R5035 VDDA.n368 VDDA.n367 185
R5036 VDDA.n366 VDDA.n365 185
R5037 VDDA.n364 VDDA.n363 185
R5038 VDDA.n362 VDDA.n361 185
R5039 VDDA.n360 VDDA.n359 185
R5040 VDDA.n358 VDDA.n357 185
R5041 VDDA.n356 VDDA.n355 185
R5042 VDDA.n377 VDDA.n335 185
R5043 VDDA.n304 VDDA.n303 185
R5044 VDDA.n306 VDDA.n305 185
R5045 VDDA.n318 VDDA.n298 185
R5046 VDDA.n312 VDDA.n298 185
R5047 VDDA.n316 VDDA.n299 185
R5048 VDDA.n315 VDDA.n300 185
R5049 VDDA.n313 VDDA.n312 185
R5050 VDDA.n239 VDDA.n238 185
R5051 VDDA.n275 VDDA.n274 185
R5052 VDDA.n276 VDDA.n275 185
R5053 VDDA.n273 VDDA.n265 185
R5054 VDDA.n271 VDDA.n270 185
R5055 VDDA.n269 VDDA.n268 185
R5056 VDDA.n261 VDDA.n260 185
R5057 VDDA.n262 VDDA.n261 185
R5058 VDDA.n247 VDDA.n243 185
R5059 VDDA.n250 VDDA.n249 185
R5060 VDDA.n252 VDDA.n251 185
R5061 VDDA.n255 VDDA.n254 185
R5062 VDDA.n257 VDDA.n256 185
R5063 VDDA.n181 VDDA.n180 185
R5064 VDDA.n227 VDDA.n226 185
R5065 VDDA.n228 VDDA.n227 185
R5066 VDDA.n225 VDDA.n222 185
R5067 VDDA.n209 VDDA.n185 185
R5068 VDDA.n213 VDDA.n184 185
R5069 VDDA.n221 VDDA.n184 185
R5070 VDDA.n212 VDDA.n211 185
R5071 VDDA.n201 VDDA.n200 185
R5072 VDDA.n200 VDDA.n199 185
R5073 VDDA.n190 VDDA.n189 185
R5074 VDDA.n195 VDDA.n194 185
R5075 VDDA.n196 VDDA.n192 185
R5076 VDDA.n144 VDDA.n89 185
R5077 VDDA.n170 VDDA.n169 185
R5078 VDDA.n171 VDDA.n170 185
R5079 VDDA.n168 VDDA.n143 185
R5080 VDDA.n167 VDDA.n166 185
R5081 VDDA.n165 VDDA.n164 185
R5082 VDDA.n163 VDDA.n162 185
R5083 VDDA.n161 VDDA.n160 185
R5084 VDDA.n159 VDDA.n158 185
R5085 VDDA.n157 VDDA.n156 185
R5086 VDDA.n155 VDDA.n154 185
R5087 VDDA.n171 VDDA.n142 185
R5088 VDDA.n136 VDDA.n135 185
R5089 VDDA.n137 VDDA.n136 185
R5090 VDDA.n133 VDDA.n96 185
R5091 VDDA.n132 VDDA.n107 185
R5092 VDDA.n131 VDDA.n108 185
R5093 VDDA.n110 VDDA.n109 185
R5094 VDDA.n127 VDDA.n111 185
R5095 VDDA.n126 VDDA.n112 185
R5096 VDDA.n114 VDDA.n113 185
R5097 VDDA.n122 VDDA.n116 185
R5098 VDDA.n121 VDDA.n117 185
R5099 VDDA.n120 VDDA.n118 185
R5100 VDDA.n137 VDDA.n95 185
R5101 VDDA.n67 VDDA.n66 185
R5102 VDDA.n69 VDDA.n68 185
R5103 VDDA.n83 VDDA.n82 185
R5104 VDDA.n82 VDDA.n81 185
R5105 VDDA.n77 VDDA.n64 185
R5106 VDDA.n78 VDDA.n76 185
R5107 VDDA.n81 VDDA.n80 185
R5108 VDDA.n4 VDDA.n3 185
R5109 VDDA.n40 VDDA.n39 185
R5110 VDDA.n41 VDDA.n40 185
R5111 VDDA.n38 VDDA.n30 185
R5112 VDDA.n36 VDDA.n35 185
R5113 VDDA.n34 VDDA.n33 185
R5114 VDDA.n26 VDDA.n25 185
R5115 VDDA.n27 VDDA.n26 185
R5116 VDDA.n12 VDDA.n8 185
R5117 VDDA.n15 VDDA.n14 185
R5118 VDDA.n17 VDDA.n16 185
R5119 VDDA.n20 VDDA.n19 185
R5120 VDDA.n22 VDDA.n21 185
R5121 VDDA.n579 VDDA.n578 185
R5122 VDDA.n584 VDDA.n577 185
R5123 VDDA.n588 VDDA.n577 185
R5124 VDDA.n583 VDDA.n582 185
R5125 VDDA.n581 VDDA.n536 185
R5126 VDDA.n590 VDDA.n589 185
R5127 VDDA.n589 VDDA.n588 185
R5128 VDDA.n575 VDDA.n574 185
R5129 VDDA.n572 VDDA.n540 185
R5130 VDDA.n571 VDDA.n542 185
R5131 VDDA.n570 VDDA.n543 185
R5132 VDDA.n545 VDDA.n544 185
R5133 VDDA.n567 VDDA.n539 185
R5134 VDDA.n575 VDDA.n539 185
R5135 VDDA.t342 VDDA.t400 180.173
R5136 VDDA.t400 VDDA.t38 180.173
R5137 VDDA.t38 VDDA.t382 180.173
R5138 VDDA.t382 VDDA.t378 180.173
R5139 VDDA.t378 VDDA.t369 180.173
R5140 VDDA.t386 VDDA.t287 180.173
R5141 VDDA.t379 VDDA.t386 180.173
R5142 VDDA.t387 VDDA.t379 180.173
R5143 VDDA.t109 VDDA.t387 180.173
R5144 VDDA.t290 VDDA.t109 180.173
R5145 VDDA.t330 VDDA.n447 170.513
R5146 VDDA.n461 VDDA.t357 170.513
R5147 VDDA.t293 VDDA.n262 170.513
R5148 VDDA.n276 VDDA.t363 170.513
R5149 VDDA.t324 VDDA.n27 170.513
R5150 VDDA.n41 VDDA.t278 170.513
R5151 VDDA.n534 VDDA.n533 168.435
R5152 VDDA.n552 VDDA.n551 168.435
R5153 VDDA.n554 VDDA.n553 168.435
R5154 VDDA.n556 VDDA.n555 168.435
R5155 VDDA.n558 VDDA.n557 168.435
R5156 VDDA.n560 VDDA.n559 168.435
R5157 VDDA.n562 VDDA.n561 168.435
R5158 VDDA.n564 VDDA.n563 168.435
R5159 VDDA.n443 VDDA.n422 159.803
R5160 VDDA.n236 VDDA.n235 159.803
R5161 VDDA.n245 VDDA.n244 159.803
R5162 VDDA.n281 VDDA.n280 159.803
R5163 VDDA.n283 VDDA.n282 159.803
R5164 VDDA.n1 VDDA.n0 159.803
R5165 VDDA.n10 VDDA.n9 159.803
R5166 VDDA.n46 VDDA.n45 159.803
R5167 VDDA.n48 VDDA.n47 159.803
R5168 VDDA.n286 VDDA.n285 155.303
R5169 VDDA.n51 VDDA.n50 155.303
R5170 VDDA.n460 VDDA.n425 150
R5171 VDDA.n460 VDDA.n450 150
R5172 VDDA.n455 VDDA.n454 150
R5173 VDDA.n446 VDDA.n429 150
R5174 VDDA.n435 VDDA.n434 150
R5175 VDDA.n440 VDDA.n439 150
R5176 VDDA.n405 VDDA.n324 150
R5177 VDDA.n405 VDDA.n378 150
R5178 VDDA.n401 VDDA.n400 150
R5179 VDDA.n397 VDDA.n396 150
R5180 VDDA.n393 VDDA.n392 150
R5181 VDDA.n389 VDDA.n329 150
R5182 VDDA.n376 VDDA.n336 150
R5183 VDDA.n371 VDDA.n370 150
R5184 VDDA.n367 VDDA.n366 150
R5185 VDDA.n363 VDDA.n362 150
R5186 VDDA.n359 VDDA.n358 150
R5187 VDDA.n355 VDDA.n335 150
R5188 VDDA.n305 VDDA.n303 150
R5189 VDDA.n299 VDDA.n298 150
R5190 VDDA.n313 VDDA.n300 150
R5191 VDDA.n275 VDDA.n239 150
R5192 VDDA.n275 VDDA.n265 150
R5193 VDDA.n270 VDDA.n269 150
R5194 VDDA.n261 VDDA.n243 150
R5195 VDDA.n251 VDDA.n250 150
R5196 VDDA.n256 VDDA.n255 150
R5197 VDDA.n185 VDDA.n184 150
R5198 VDDA.n211 VDDA.n184 150
R5199 VDDA.n227 VDDA.n181 150
R5200 VDDA.n227 VDDA.n222 150
R5201 VDDA.n200 VDDA.n190 150
R5202 VDDA.n194 VDDA.n192 150
R5203 VDDA.n170 VDDA.n89 150
R5204 VDDA.n170 VDDA.n143 150
R5205 VDDA.n166 VDDA.n165 150
R5206 VDDA.n162 VDDA.n161 150
R5207 VDDA.n158 VDDA.n157 150
R5208 VDDA.n154 VDDA.n142 150
R5209 VDDA.n136 VDDA.n96 150
R5210 VDDA.n108 VDDA.n107 150
R5211 VDDA.n111 VDDA.n110 150
R5212 VDDA.n113 VDDA.n112 150
R5213 VDDA.n117 VDDA.n116 150
R5214 VDDA.n118 VDDA.n95 150
R5215 VDDA.n68 VDDA.n66 150
R5216 VDDA.n82 VDDA.n64 150
R5217 VDDA.n80 VDDA.n76 150
R5218 VDDA.n40 VDDA.n4 150
R5219 VDDA.n40 VDDA.n30 150
R5220 VDDA.n35 VDDA.n34 150
R5221 VDDA.n26 VDDA.n8 150
R5222 VDDA.n16 VDDA.n15 150
R5223 VDDA.n21 VDDA.n20 150
R5224 VDDA.n578 VDDA.n577 150
R5225 VDDA.n582 VDDA.n577 150
R5226 VDDA.n589 VDDA.n536 150
R5227 VDDA.n574 VDDA.n540 150
R5228 VDDA.n543 VDDA.n542 150
R5229 VDDA.n544 VDDA.n539 150
R5230 VDDA.t250 VDDA.t330 146.155
R5231 VDDA.t357 VDDA.t250 146.155
R5232 VDDA.t234 VDDA.t293 146.155
R5233 VDDA.t230 VDDA.t234 146.155
R5234 VDDA.t238 VDDA.t230 146.155
R5235 VDDA.t248 VDDA.t238 146.155
R5236 VDDA.t258 VDDA.t248 146.155
R5237 VDDA.t228 VDDA.t258 146.155
R5238 VDDA.t226 VDDA.t228 146.155
R5239 VDDA.t232 VDDA.t226 146.155
R5240 VDDA.t240 VDDA.t232 146.155
R5241 VDDA.t252 VDDA.t240 146.155
R5242 VDDA.t363 VDDA.t252 146.155
R5243 VDDA.t246 VDDA.t324 146.155
R5244 VDDA.t242 VDDA.t246 146.155
R5245 VDDA.t254 VDDA.t242 146.155
R5246 VDDA.t260 VDDA.t254 146.155
R5247 VDDA.t222 VDDA.t260 146.155
R5248 VDDA.t224 VDDA.t222 146.155
R5249 VDDA.t236 VDDA.t224 146.155
R5250 VDDA.t244 VDDA.t236 146.155
R5251 VDDA.t256 VDDA.t244 146.155
R5252 VDDA.t262 VDDA.t256 146.155
R5253 VDDA.t278 VDDA.t262 146.155
R5254 VDDA.n322 VDDA.n321 145.429
R5255 VDDA.n338 VDDA.n337 145.429
R5256 VDDA.n340 VDDA.n339 145.429
R5257 VDDA.n342 VDDA.n341 145.429
R5258 VDDA.n344 VDDA.n343 145.429
R5259 VDDA.n87 VDDA.n86 145.429
R5260 VDDA.n98 VDDA.n97 145.429
R5261 VDDA.n100 VDDA.n99 145.429
R5262 VDDA.n102 VDDA.n101 145.429
R5263 VDDA.n104 VDDA.n103 145.429
R5264 VDDA.t273 VDDA.n383 123.126
R5265 VDDA.n384 VDDA.t273 123.126
R5266 VDDA.t297 VDDA.n349 123.126
R5267 VDDA.n350 VDDA.t297 123.126
R5268 VDDA.n128 VDDA.t313 123.126
R5269 VDDA.n125 VDDA.t313 123.126
R5270 VDDA.t328 VDDA.n148 123.126
R5271 VDDA.n149 VDDA.t328 123.126
R5272 VDDA.t303 VDDA.n541 123.126
R5273 VDDA.n569 VDDA.t303 123.126
R5274 VDDA.n585 VDDA.t270 123.126
R5275 VDDA.n580 VDDA.t270 123.126
R5276 VDDA.n406 VDDA.t272 100.195
R5277 VDDA.t296 VDDA.n377 100.195
R5278 VDDA.t312 VDDA.n137 100.195
R5279 VDDA.n171 VDDA.t327 100.195
R5280 VDDA.n289 VDDA.n287 97.4002
R5281 VDDA.n54 VDDA.n52 97.4002
R5282 VDDA.n297 VDDA.n296 96.8377
R5283 VDDA.n295 VDDA.n294 96.8377
R5284 VDDA.n293 VDDA.n292 96.8377
R5285 VDDA.n291 VDDA.n290 96.8377
R5286 VDDA.n289 VDDA.n288 96.8377
R5287 VDDA.n62 VDDA.n61 96.8377
R5288 VDDA.n60 VDDA.n59 96.8377
R5289 VDDA.n58 VDDA.n57 96.8377
R5290 VDDA.n56 VDDA.n55 96.8377
R5291 VDDA.n54 VDDA.n53 96.8377
R5292 VDDA.t272 VDDA.t393 81.6411
R5293 VDDA.t393 VDDA.t26 81.6411
R5294 VDDA.t26 VDDA.t212 81.6411
R5295 VDDA.t212 VDDA.t94 81.6411
R5296 VDDA.t94 VDDA.t28 81.6411
R5297 VDDA.t28 VDDA.t164 81.6411
R5298 VDDA.t164 VDDA.t413 81.6411
R5299 VDDA.t413 VDDA.t168 81.6411
R5300 VDDA.t168 VDDA.t384 81.6411
R5301 VDDA.t384 VDDA.t201 81.6411
R5302 VDDA.t201 VDDA.t296 81.6411
R5303 VDDA.t134 VDDA.t312 81.6411
R5304 VDDA.t153 VDDA.t134 81.6411
R5305 VDDA.t131 VDDA.t153 81.6411
R5306 VDDA.t92 VDDA.t131 81.6411
R5307 VDDA.t76 VDDA.t92 81.6411
R5308 VDDA.t148 VDDA.t76 81.6411
R5309 VDDA.t51 VDDA.t148 81.6411
R5310 VDDA.t151 VDDA.t51 81.6411
R5311 VDDA.t49 VDDA.t151 81.6411
R5312 VDDA.t71 VDDA.t49 81.6411
R5313 VDDA.t327 VDDA.t71 81.6411
R5314 VDDA.n462 VDDA.n461 65.8183
R5315 VDDA.n461 VDDA.n448 65.8183
R5316 VDDA.n461 VDDA.n449 65.8183
R5317 VDDA.n447 VDDA.n426 65.8183
R5318 VDDA.n447 VDDA.n427 65.8183
R5319 VDDA.n447 VDDA.n428 65.8183
R5320 VDDA.n407 VDDA.n406 65.8183
R5321 VDDA.n406 VDDA.n325 65.8183
R5322 VDDA.n406 VDDA.n326 65.8183
R5323 VDDA.n406 VDDA.n327 65.8183
R5324 VDDA.n406 VDDA.n328 65.8183
R5325 VDDA.n377 VDDA.n330 65.8183
R5326 VDDA.n377 VDDA.n331 65.8183
R5327 VDDA.n377 VDDA.n332 65.8183
R5328 VDDA.n377 VDDA.n333 65.8183
R5329 VDDA.n377 VDDA.n334 65.8183
R5330 VDDA.n311 VDDA.n310 65.8183
R5331 VDDA.n311 VDDA.n302 65.8183
R5332 VDDA.n312 VDDA.n301 65.8183
R5333 VDDA.n277 VDDA.n276 65.8183
R5334 VDDA.n276 VDDA.n263 65.8183
R5335 VDDA.n276 VDDA.n264 65.8183
R5336 VDDA.n262 VDDA.n240 65.8183
R5337 VDDA.n262 VDDA.n241 65.8183
R5338 VDDA.n262 VDDA.n242 65.8183
R5339 VDDA.n229 VDDA.n228 65.8183
R5340 VDDA.n228 VDDA.n182 65.8183
R5341 VDDA.n221 VDDA.n220 65.8183
R5342 VDDA.n221 VDDA.n183 65.8183
R5343 VDDA.n199 VDDA.n191 65.8183
R5344 VDDA.n199 VDDA.n198 65.8183
R5345 VDDA.n172 VDDA.n171 65.8183
R5346 VDDA.n171 VDDA.n138 65.8183
R5347 VDDA.n171 VDDA.n139 65.8183
R5348 VDDA.n171 VDDA.n140 65.8183
R5349 VDDA.n171 VDDA.n141 65.8183
R5350 VDDA.n137 VDDA.n90 65.8183
R5351 VDDA.n137 VDDA.n91 65.8183
R5352 VDDA.n137 VDDA.n92 65.8183
R5353 VDDA.n137 VDDA.n93 65.8183
R5354 VDDA.n137 VDDA.n94 65.8183
R5355 VDDA.n74 VDDA.n73 65.8183
R5356 VDDA.n74 VDDA.n65 65.8183
R5357 VDDA.n81 VDDA.n75 65.8183
R5358 VDDA.n42 VDDA.n41 65.8183
R5359 VDDA.n41 VDDA.n28 65.8183
R5360 VDDA.n41 VDDA.n29 65.8183
R5361 VDDA.n27 VDDA.n5 65.8183
R5362 VDDA.n27 VDDA.n6 65.8183
R5363 VDDA.n27 VDDA.n7 65.8183
R5364 VDDA.n588 VDDA.n587 65.8183
R5365 VDDA.n588 VDDA.n576 65.8183
R5366 VDDA.n575 VDDA.n537 65.8183
R5367 VDDA.n575 VDDA.n538 65.8183
R5368 VDDA.n475 VDDA.t417 59.5681
R5369 VDDA.n474 VDDA.t418 59.5681
R5370 VDDA.n450 VDDA.n448 53.3664
R5371 VDDA.n454 VDDA.n449 53.3664
R5372 VDDA.n462 VDDA.n425 53.3664
R5373 VDDA.n455 VDDA.n448 53.3664
R5374 VDDA.n429 VDDA.n426 53.3664
R5375 VDDA.n435 VDDA.n427 53.3664
R5376 VDDA.n440 VDDA.n428 53.3664
R5377 VDDA.n434 VDDA.n426 53.3664
R5378 VDDA.n439 VDDA.n427 53.3664
R5379 VDDA.n378 VDDA.n325 53.3664
R5380 VDDA.n400 VDDA.n326 53.3664
R5381 VDDA.n396 VDDA.n327 53.3664
R5382 VDDA.n392 VDDA.n328 53.3664
R5383 VDDA.n407 VDDA.n324 53.3664
R5384 VDDA.n401 VDDA.n325 53.3664
R5385 VDDA.n397 VDDA.n326 53.3664
R5386 VDDA.n393 VDDA.n327 53.3664
R5387 VDDA.n389 VDDA.n328 53.3664
R5388 VDDA.n336 VDDA.n330 53.3664
R5389 VDDA.n370 VDDA.n331 53.3664
R5390 VDDA.n366 VDDA.n332 53.3664
R5391 VDDA.n362 VDDA.n333 53.3664
R5392 VDDA.n358 VDDA.n334 53.3664
R5393 VDDA.n371 VDDA.n330 53.3664
R5394 VDDA.n367 VDDA.n331 53.3664
R5395 VDDA.n363 VDDA.n332 53.3664
R5396 VDDA.n359 VDDA.n333 53.3664
R5397 VDDA.n355 VDDA.n334 53.3664
R5398 VDDA.n310 VDDA.n303 53.3664
R5399 VDDA.n305 VDDA.n302 53.3664
R5400 VDDA.n301 VDDA.n299 53.3664
R5401 VDDA.n301 VDDA.n300 53.3664
R5402 VDDA.n265 VDDA.n263 53.3664
R5403 VDDA.n269 VDDA.n264 53.3664
R5404 VDDA.n277 VDDA.n239 53.3664
R5405 VDDA.n270 VDDA.n263 53.3664
R5406 VDDA.n243 VDDA.n240 53.3664
R5407 VDDA.n251 VDDA.n241 53.3664
R5408 VDDA.n256 VDDA.n242 53.3664
R5409 VDDA.n250 VDDA.n240 53.3664
R5410 VDDA.n255 VDDA.n241 53.3664
R5411 VDDA.n211 VDDA.n183 53.3664
R5412 VDDA.n222 VDDA.n182 53.3664
R5413 VDDA.n229 VDDA.n181 53.3664
R5414 VDDA.n220 VDDA.n185 53.3664
R5415 VDDA.n191 VDDA.n190 53.3664
R5416 VDDA.n198 VDDA.n192 53.3664
R5417 VDDA.n194 VDDA.n191 53.3664
R5418 VDDA.n143 VDDA.n138 53.3664
R5419 VDDA.n165 VDDA.n139 53.3664
R5420 VDDA.n161 VDDA.n140 53.3664
R5421 VDDA.n157 VDDA.n141 53.3664
R5422 VDDA.n172 VDDA.n89 53.3664
R5423 VDDA.n166 VDDA.n138 53.3664
R5424 VDDA.n162 VDDA.n139 53.3664
R5425 VDDA.n158 VDDA.n140 53.3664
R5426 VDDA.n154 VDDA.n141 53.3664
R5427 VDDA.n96 VDDA.n90 53.3664
R5428 VDDA.n108 VDDA.n91 53.3664
R5429 VDDA.n111 VDDA.n92 53.3664
R5430 VDDA.n113 VDDA.n93 53.3664
R5431 VDDA.n117 VDDA.n94 53.3664
R5432 VDDA.n107 VDDA.n90 53.3664
R5433 VDDA.n110 VDDA.n91 53.3664
R5434 VDDA.n112 VDDA.n92 53.3664
R5435 VDDA.n116 VDDA.n93 53.3664
R5436 VDDA.n118 VDDA.n94 53.3664
R5437 VDDA.n73 VDDA.n66 53.3664
R5438 VDDA.n68 VDDA.n65 53.3664
R5439 VDDA.n75 VDDA.n64 53.3664
R5440 VDDA.n76 VDDA.n75 53.3664
R5441 VDDA.n30 VDDA.n28 53.3664
R5442 VDDA.n34 VDDA.n29 53.3664
R5443 VDDA.n42 VDDA.n4 53.3664
R5444 VDDA.n35 VDDA.n28 53.3664
R5445 VDDA.n8 VDDA.n5 53.3664
R5446 VDDA.n16 VDDA.n6 53.3664
R5447 VDDA.n21 VDDA.n7 53.3664
R5448 VDDA.n15 VDDA.n5 53.3664
R5449 VDDA.n20 VDDA.n6 53.3664
R5450 VDDA.n582 VDDA.n576 53.3664
R5451 VDDA.n587 VDDA.n578 53.3664
R5452 VDDA.n576 VDDA.n536 53.3664
R5453 VDDA.n540 VDDA.n537 53.3664
R5454 VDDA.n543 VDDA.n538 53.3664
R5455 VDDA.n542 VDDA.n537 53.3664
R5456 VDDA.n544 VDDA.n538 53.3664
R5457 VDDA.n474 VDDA.t416 52.3888
R5458 VDDA.n231 VDDA.n230 51.6576
R5459 VDDA.n202 VDDA.n201 51.6576
R5460 VDDA.n476 VDDA.t415 48.9557
R5461 VDDA.n207 VDDA.n206 48.0005
R5462 VDDA.n207 VDDA.n186 48.0005
R5463 VDDA.n419 VDDA.n418 46.6291
R5464 VDDA.n417 VDDA.n416 46.6291
R5465 VDDA.n478 VDDA.t88 39.4005
R5466 VDDA.n478 VDDA.t18 39.4005
R5467 VDDA.n508 VDDA.t125 39.4005
R5468 VDDA.n508 VDDA.t11 39.4005
R5469 VDDA.n510 VDDA.t20 39.4005
R5470 VDDA.n510 VDDA.t123 39.4005
R5471 VDDA.n512 VDDA.t45 39.4005
R5472 VDDA.n512 VDDA.t411 39.4005
R5473 VDDA.n514 VDDA.t9 39.4005
R5474 VDDA.n514 VDDA.t31 39.4005
R5475 VDDA.n516 VDDA.t111 39.4005
R5476 VDDA.n516 VDDA.t171 39.4005
R5477 VDDA.n518 VDDA.t220 39.4005
R5478 VDDA.n518 VDDA.t406 39.4005
R5479 VDDA.n520 VDDA.t5 39.4005
R5480 VDDA.n520 VDDA.t197 39.4005
R5481 VDDA.n522 VDDA.t404 39.4005
R5482 VDDA.n522 VDDA.t58 39.4005
R5483 VDDA.n483 VDDA.t183 39.4005
R5484 VDDA.n483 VDDA.t79 39.4005
R5485 VDDA.n486 VDDA.t392 39.4005
R5486 VDDA.n486 VDDA.t185 39.4005
R5487 VDDA.n488 VDDA.t390 39.4005
R5488 VDDA.n488 VDDA.t81 39.4005
R5489 VDDA.n490 VDDA.t1 39.4005
R5490 VDDA.n490 VDDA.t181 39.4005
R5491 VDDA.n492 VDDA.t129 39.4005
R5492 VDDA.n492 VDDA.t83 39.4005
R5493 VDDA.n494 VDDA.t402 39.4005
R5494 VDDA.n494 VDDA.t16 39.4005
R5495 VDDA.n496 VDDA.t177 39.4005
R5496 VDDA.n496 VDDA.t179 39.4005
R5497 VDDA.n498 VDDA.t25 39.4005
R5498 VDDA.n498 VDDA.t3 39.4005
R5499 VDDA.n500 VDDA.t137 39.4005
R5500 VDDA.n500 VDDA.t139 39.4005
R5501 VDDA.n598 VDDA.t85 39.4005
R5502 VDDA.n598 VDDA.t175 39.4005
R5503 VDDA.n602 VDDA.t54 39.4005
R5504 VDDA.n602 VDDA.t67 39.4005
R5505 VDDA.n629 VDDA.t216 39.4005
R5506 VDDA.n629 VDDA.t7 39.4005
R5507 VDDA.n604 VDDA.t195 39.4005
R5508 VDDA.n604 VDDA.t191 39.4005
R5509 VDDA.n615 VDDA.t199 39.4005
R5510 VDDA.n615 VDDA.t119 39.4005
R5511 VDDA.n617 VDDA.t398 39.4005
R5512 VDDA.n617 VDDA.t47 39.4005
R5513 VDDA.n619 VDDA.t218 39.4005
R5514 VDDA.n619 VDDA.t33 39.4005
R5515 VDDA.n621 VDDA.t65 39.4005
R5516 VDDA.n621 VDDA.t396 39.4005
R5517 VDDA.n606 VDDA.t173 39.4005
R5518 VDDA.n606 VDDA.t121 39.4005
R5519 VDDA.n608 VDDA.t211 39.4005
R5520 VDDA.n608 VDDA.t193 39.4005
R5521 VDDA.n473 VDDA.n467 27.9413
R5522 VDDA.n635 VDDA.n634 27.2462
R5523 VDDA.n633 VDDA.n632 27.2462
R5524 VDDA.n613 VDDA.n612 27.2462
R5525 VDDA.n611 VDDA.n610 27.2462
R5526 VDDA.n594 VDDA.n593 25.087
R5527 VDDA.n596 VDDA.n595 25.087
R5528 VDDA.n627 VDDA.n626 25.0384
R5529 VDDA.n625 VDDA.n624 25.0384
R5530 VDDA.n547 VDDA.n546 22.9536
R5531 VDDA.n506 VDDA.n505 22.9536
R5532 VDDA.n464 VDDA.n463 22.8576
R5533 VDDA.n445 VDDA.n430 22.8576
R5534 VDDA.n409 VDDA.n408 22.8576
R5535 VDDA.n375 VDDA.n345 22.8576
R5536 VDDA.n319 VDDA.n318 22.8576
R5537 VDDA.n279 VDDA.n278 22.8576
R5538 VDDA.n260 VDDA.n246 22.8576
R5539 VDDA.n174 VDDA.n173 22.8576
R5540 VDDA.n135 VDDA.n105 22.8576
R5541 VDDA.n84 VDDA.n83 22.8576
R5542 VDDA.n44 VDDA.n43 22.8576
R5543 VDDA.n25 VDDA.n11 22.8576
R5544 VDDA.n591 VDDA.n590 22.8576
R5545 VDDA.n567 VDDA.n566 22.8576
R5546 VDDA.n414 VDDA.t408 21.8894
R5547 VDDA.n414 VDDA.t309 21.8894
R5548 VDDA.n467 VDDA.n466 20.883
R5549 VDDA.n530 VDDA.n480 20.7243
R5550 VDDA.n525 VDDA.n482 20.7243
R5551 VDDA.n502 VDDA.n485 20.7243
R5552 VDDA.n549 VDDA.n548 20.4312
R5553 VDDA.n473 VDDA.t115 19.9244
R5554 VDDA.n320 VDDA.n319 19.613
R5555 VDDA.n85 VDDA.n84 19.613
R5556 VDDA.n177 VDDA.t39 15.7605
R5557 VDDA.n177 VDDA.t383 15.7605
R5558 VDDA.n203 VDDA.t380 15.7605
R5559 VDDA.n203 VDDA.t388 15.7605
R5560 VDDA.n215 VDDA.t288 15.7605
R5561 VDDA.n218 VDDA.t370 15.7605
R5562 VDDA.n179 VDDA.t343 15.7605
R5563 VDDA.n188 VDDA.t291 15.7605
R5564 VDDA.n550 VDDA.n546 15.488
R5565 VDDA.n204 VDDA.n202 14.7224
R5566 VDDA.n502 VDDA.n501 14.6963
R5567 VDDA.n281 VDDA.n279 14.4255
R5568 VDDA.n246 VDDA.n245 14.4255
R5569 VDDA.n46 VDDA.n44 14.4255
R5570 VDDA.n11 VDDA.n10 14.4255
R5571 VDDA.n345 VDDA.n344 14.363
R5572 VDDA.n105 VDDA.n104 14.363
R5573 VDDA.n597 VDDA.n596 14.363
R5574 VDDA.n597 VDDA.n593 14.363
R5575 VDDA.n610 VDDA.n609 14.363
R5576 VDDA.n550 VDDA.n549 14.238
R5577 VDDA.n525 VDDA.n524 14.0713
R5578 VDDA.n531 VDDA.n530 14.0713
R5579 VDDA.n507 VDDA.n506 14.0713
R5580 VDDA.n430 VDDA.n422 14.0505
R5581 VDDA.n416 VDDA.n415 14.0505
R5582 VDDA.n465 VDDA.n464 13.8005
R5583 VDDA.n420 VDDA.n419 13.8005
R5584 VDDA.n410 VDDA.n409 13.8005
R5585 VDDA.n206 VDDA.n205 13.8005
R5586 VDDA.n187 VDDA.n186 13.8005
R5587 VDDA.n232 VDDA.n231 13.8005
R5588 VDDA.n175 VDDA.n174 13.8005
R5589 VDDA.n566 VDDA.n565 13.8005
R5590 VDDA.n592 VDDA.n591 13.8005
R5591 VDDA.n632 VDDA.n631 13.8005
R5592 VDDA.n624 VDDA.n623 13.8005
R5593 VDDA.n614 VDDA.n613 13.8005
R5594 VDDA.n628 VDDA.n627 13.8005
R5595 VDDA.n636 VDDA.n635 13.8005
R5596 VDDA.n533 VDDA.t205 13.1338
R5597 VDDA.n533 VDDA.t98 13.1338
R5598 VDDA.n551 VDDA.t113 13.1338
R5599 VDDA.n551 VDDA.t106 13.1338
R5600 VDDA.n553 VDDA.t60 13.1338
R5601 VDDA.n553 VDDA.t62 13.1338
R5602 VDDA.n555 VDDA.t104 13.1338
R5603 VDDA.n555 VDDA.t143 13.1338
R5604 VDDA.n557 VDDA.t141 13.1338
R5605 VDDA.n557 VDDA.t117 13.1338
R5606 VDDA.n559 VDDA.t102 13.1338
R5607 VDDA.n559 VDDA.t208 13.1338
R5608 VDDA.n561 VDDA.t187 13.1338
R5609 VDDA.n561 VDDA.t36 13.1338
R5610 VDDA.n563 VDDA.t145 13.1338
R5611 VDDA.n563 VDDA.t161 13.1338
R5612 VDDA.n637 VDDA.n636 11.4105
R5613 VDDA.t331 VDDA.n443 11.2576
R5614 VDDA.n443 VDDA.t251 11.2576
R5615 VDDA.n444 VDDA.t331 11.2576
R5616 VDDA.n423 VDDA.t358 11.2576
R5617 VDDA.n285 VDDA.t259 11.2576
R5618 VDDA.n285 VDDA.t229 11.2576
R5619 VDDA.n235 VDDA.t239 11.2576
R5620 VDDA.n235 VDDA.t249 11.2576
R5621 VDDA.n244 VDDA.t235 11.2576
R5622 VDDA.n244 VDDA.t231 11.2576
R5623 VDDA.n259 VDDA.t294 11.2576
R5624 VDDA.n237 VDDA.t364 11.2576
R5625 VDDA.n280 VDDA.t241 11.2576
R5626 VDDA.n280 VDDA.t253 11.2576
R5627 VDDA.n282 VDDA.t227 11.2576
R5628 VDDA.n282 VDDA.t233 11.2576
R5629 VDDA.n50 VDDA.t223 11.2576
R5630 VDDA.n50 VDDA.t225 11.2576
R5631 VDDA.n0 VDDA.t255 11.2576
R5632 VDDA.n0 VDDA.t261 11.2576
R5633 VDDA.n9 VDDA.t247 11.2576
R5634 VDDA.n9 VDDA.t243 11.2576
R5635 VDDA.n24 VDDA.t325 11.2576
R5636 VDDA.n2 VDDA.t279 11.2576
R5637 VDDA.n45 VDDA.t257 11.2576
R5638 VDDA.n45 VDDA.t263 11.2576
R5639 VDDA.n47 VDDA.t237 11.2576
R5640 VDDA.n47 VDDA.t245 11.2576
R5641 VDDA.n477 VDDA.n476 11.1572
R5642 VDDA.n85 VDDA.n62 10.938
R5643 VDDA.n320 VDDA.n297 10.9067
R5644 VDDA.n601 VDDA.n600 9.7855
R5645 VDDA.n463 VDDA.n424 9.14336
R5646 VDDA.n459 VDDA.n458 9.14336
R5647 VDDA.n456 VDDA.n453 9.14336
R5648 VDDA.n445 VDDA.n431 9.14336
R5649 VDDA.n436 VDDA.n433 9.14336
R5650 VDDA.n441 VDDA.n438 9.14336
R5651 VDDA.n404 VDDA.n379 9.14336
R5652 VDDA.n404 VDDA.n403 9.14336
R5653 VDDA.n403 VDDA.n402 9.14336
R5654 VDDA.n402 VDDA.n399 9.14336
R5655 VDDA.n399 VDDA.n398 9.14336
R5656 VDDA.n398 VDDA.n395 9.14336
R5657 VDDA.n395 VDDA.n394 9.14336
R5658 VDDA.n394 VDDA.n391 9.14336
R5659 VDDA.n391 VDDA.n390 9.14336
R5660 VDDA.n372 VDDA.n346 9.14336
R5661 VDDA.n372 VDDA.n369 9.14336
R5662 VDDA.n369 VDDA.n368 9.14336
R5663 VDDA.n368 VDDA.n365 9.14336
R5664 VDDA.n365 VDDA.n364 9.14336
R5665 VDDA.n364 VDDA.n361 9.14336
R5666 VDDA.n361 VDDA.n360 9.14336
R5667 VDDA.n360 VDDA.n357 9.14336
R5668 VDDA.n357 VDDA.n356 9.14336
R5669 VDDA.n306 VDDA.n304 9.14336
R5670 VDDA.n316 VDDA.n315 9.14336
R5671 VDDA.n278 VDDA.n238 9.14336
R5672 VDDA.n274 VDDA.n273 9.14336
R5673 VDDA.n271 VDDA.n268 9.14336
R5674 VDDA.n260 VDDA.n247 9.14336
R5675 VDDA.n252 VDDA.n249 9.14336
R5676 VDDA.n257 VDDA.n254 9.14336
R5677 VDDA.n230 VDDA.n180 9.14336
R5678 VDDA.n226 VDDA.n225 9.14336
R5679 VDDA.n201 VDDA.n189 9.14336
R5680 VDDA.n196 VDDA.n195 9.14336
R5681 VDDA.n169 VDDA.n144 9.14336
R5682 VDDA.n169 VDDA.n168 9.14336
R5683 VDDA.n168 VDDA.n167 9.14336
R5684 VDDA.n167 VDDA.n164 9.14336
R5685 VDDA.n164 VDDA.n163 9.14336
R5686 VDDA.n163 VDDA.n160 9.14336
R5687 VDDA.n160 VDDA.n159 9.14336
R5688 VDDA.n159 VDDA.n156 9.14336
R5689 VDDA.n156 VDDA.n155 9.14336
R5690 VDDA.n133 VDDA.n132 9.14336
R5691 VDDA.n132 VDDA.n131 9.14336
R5692 VDDA.n131 VDDA.n109 9.14336
R5693 VDDA.n127 VDDA.n109 9.14336
R5694 VDDA.n127 VDDA.n126 9.14336
R5695 VDDA.n126 VDDA.n114 9.14336
R5696 VDDA.n122 VDDA.n114 9.14336
R5697 VDDA.n122 VDDA.n121 9.14336
R5698 VDDA.n121 VDDA.n120 9.14336
R5699 VDDA.n69 VDDA.n67 9.14336
R5700 VDDA.n78 VDDA.n77 9.14336
R5701 VDDA.n43 VDDA.n3 9.14336
R5702 VDDA.n39 VDDA.n38 9.14336
R5703 VDDA.n36 VDDA.n33 9.14336
R5704 VDDA.n25 VDDA.n12 9.14336
R5705 VDDA.n17 VDDA.n14 9.14336
R5706 VDDA.n22 VDDA.n19 9.14336
R5707 VDDA.n584 VDDA.n579 9.14336
R5708 VDDA.n584 VDDA.n583 9.14336
R5709 VDDA.n583 VDDA.n581 9.14336
R5710 VDDA.n572 VDDA.n571 9.14336
R5711 VDDA.n571 VDDA.n570 9.14336
R5712 VDDA.n570 VDDA.n545 9.14336
R5713 VDDA.n532 VDDA.n531 8.973
R5714 VDDA.n412 VDDA.n411 8.8755
R5715 VDDA.n234 VDDA.n233 8.28175
R5716 VDDA.n233 VDDA.n232 8.21925
R5717 VDDA.n412 VDDA.n286 8.15675
R5718 VDDA.n234 VDDA.n51 8.15675
R5719 VDDA.n296 VDDA.t264 8.0005
R5720 VDDA.n296 VDDA.t56 8.0005
R5721 VDDA.n294 VDDA.t409 8.0005
R5722 VDDA.n294 VDDA.t48 8.0005
R5723 VDDA.n292 VDDA.t96 8.0005
R5724 VDDA.n292 VDDA.t221 8.0005
R5725 VDDA.n290 VDDA.t203 8.0005
R5726 VDDA.n290 VDDA.t68 8.0005
R5727 VDDA.n288 VDDA.t40 8.0005
R5728 VDDA.n288 VDDA.t381 8.0005
R5729 VDDA.n287 VDDA.t200 8.0005
R5730 VDDA.n287 VDDA.t265 8.0005
R5731 VDDA.n61 VDDA.t133 8.0005
R5732 VDDA.n61 VDDA.t267 8.0005
R5733 VDDA.n59 VDDA.t155 8.0005
R5734 VDDA.n59 VDDA.t157 8.0005
R5735 VDDA.n57 VDDA.t159 8.0005
R5736 VDDA.n57 VDDA.t158 8.0005
R5737 VDDA.n55 VDDA.t146 8.0005
R5738 VDDA.n55 VDDA.t89 8.0005
R5739 VDDA.n53 VDDA.t150 8.0005
R5740 VDDA.n53 VDDA.t13 8.0005
R5741 VDDA.n52 VDDA.t266 8.0005
R5742 VDDA.n52 VDDA.t73 8.0005
R5743 VDDA.n321 VDDA.t394 6.56717
R5744 VDDA.n321 VDDA.t27 6.56717
R5745 VDDA.n337 VDDA.t213 6.56717
R5746 VDDA.n337 VDDA.t95 6.56717
R5747 VDDA.n339 VDDA.t29 6.56717
R5748 VDDA.n339 VDDA.t165 6.56717
R5749 VDDA.n341 VDDA.t414 6.56717
R5750 VDDA.n341 VDDA.t169 6.56717
R5751 VDDA.n343 VDDA.t385 6.56717
R5752 VDDA.n343 VDDA.t202 6.56717
R5753 VDDA.n86 VDDA.t50 6.56717
R5754 VDDA.n86 VDDA.t72 6.56717
R5755 VDDA.n97 VDDA.t52 6.56717
R5756 VDDA.n97 VDDA.t152 6.56717
R5757 VDDA.n99 VDDA.t77 6.56717
R5758 VDDA.n99 VDDA.t149 6.56717
R5759 VDDA.n101 VDDA.t132 6.56717
R5760 VDDA.n101 VDDA.t93 6.56717
R5761 VDDA.n103 VDDA.t135 6.56717
R5762 VDDA.n103 VDDA.t154 6.56717
R5763 VDDA.n421 VDDA.n413 6.563
R5764 VDDA.n413 VDDA.n412 6.0005
R5765 VDDA.n413 VDDA.n234 6.0005
R5766 VDDA.n411 VDDA.n410 5.8755
R5767 VDDA.n176 VDDA.n175 5.8755
R5768 VDDA.n408 VDDA.n323 5.33286
R5769 VDDA.n375 VDDA.n374 5.33286
R5770 VDDA.n318 VDDA.n317 5.33286
R5771 VDDA.n309 VDDA.n308 5.33286
R5772 VDDA.n135 VDDA.n134 5.33286
R5773 VDDA.n173 VDDA.n88 5.33286
R5774 VDDA.n72 VDDA.n71 5.33286
R5775 VDDA.n83 VDDA.n63 5.33286
R5776 VDDA.n590 VDDA.n535 5.33286
R5777 VDDA.n568 VDDA.n567 5.33286
R5778 VDDA.n466 VDDA.n465 5.28175
R5779 VDDA.n421 VDDA.n420 5.28175
R5780 VDDA.n600 VDDA.n599 5.0005
R5781 VDDA.n411 VDDA.n320 4.90675
R5782 VDDA.n176 VDDA.n85 4.90675
R5783 VDDA.n477 VDDA.n473 4.5595
R5784 VDDA.n481 VDDA.n480 4.54311
R5785 VDDA.n529 VDDA.n481 4.54311
R5786 VDDA.n451 VDDA.n424 4.53698
R5787 VDDA.n458 VDDA.n457 4.53698
R5788 VDDA.n453 VDDA.n452 4.53698
R5789 VDDA.n459 VDDA.n451 4.53698
R5790 VDDA.n457 VDDA.n456 4.53698
R5791 VDDA.n432 VDDA.n431 4.53698
R5792 VDDA.n437 VDDA.n436 4.53698
R5793 VDDA.n442 VDDA.n441 4.53698
R5794 VDDA.n433 VDDA.n432 4.53698
R5795 VDDA.n438 VDDA.n437 4.53698
R5796 VDDA.n266 VDDA.n238 4.53698
R5797 VDDA.n273 VDDA.n272 4.53698
R5798 VDDA.n268 VDDA.n267 4.53698
R5799 VDDA.n274 VDDA.n266 4.53698
R5800 VDDA.n272 VDDA.n271 4.53698
R5801 VDDA.n248 VDDA.n247 4.53698
R5802 VDDA.n253 VDDA.n252 4.53698
R5803 VDDA.n258 VDDA.n257 4.53698
R5804 VDDA.n249 VDDA.n248 4.53698
R5805 VDDA.n254 VDDA.n253 4.53698
R5806 VDDA.n223 VDDA.n180 4.53698
R5807 VDDA.n225 VDDA.n224 4.53698
R5808 VDDA.n226 VDDA.n223 4.53698
R5809 VDDA.n193 VDDA.n189 4.53698
R5810 VDDA.n197 VDDA.n196 4.53698
R5811 VDDA.n195 VDDA.n193 4.53698
R5812 VDDA.n31 VDDA.n3 4.53698
R5813 VDDA.n38 VDDA.n37 4.53698
R5814 VDDA.n33 VDDA.n32 4.53698
R5815 VDDA.n39 VDDA.n31 4.53698
R5816 VDDA.n37 VDDA.n36 4.53698
R5817 VDDA.n13 VDDA.n12 4.53698
R5818 VDDA.n18 VDDA.n17 4.53698
R5819 VDDA.n23 VDDA.n22 4.53698
R5820 VDDA.n14 VDDA.n13 4.53698
R5821 VDDA.n19 VDDA.n18 4.53698
R5822 VDDA.n286 VDDA.n284 4.5005
R5823 VDDA.n51 VDDA.n49 4.5005
R5824 VDDA.n599 VDDA.n597 4.5005
R5825 VDDA.n527 VDDA.n482 4.48641
R5826 VDDA.n527 VDDA.n526 4.48641
R5827 VDDA.n504 VDDA.n485 4.48641
R5828 VDDA.n504 VDDA.n503 4.48641
R5829 VDDA.n475 VDDA.n474 4.12334
R5830 VDDA.n379 VDDA.n323 3.75335
R5831 VDDA.n390 VDDA.n388 3.75335
R5832 VDDA.n374 VDDA.n346 3.75335
R5833 VDDA.n356 VDDA.n354 3.75335
R5834 VDDA.n308 VDDA.n304 3.75335
R5835 VDDA.n307 VDDA.n306 3.75335
R5836 VDDA.n317 VDDA.n316 3.75335
R5837 VDDA.n315 VDDA.n314 3.75335
R5838 VDDA.n144 VDDA.n88 3.75335
R5839 VDDA.n155 VDDA.n153 3.75335
R5840 VDDA.n134 VDDA.n133 3.75335
R5841 VDDA.n120 VDDA.n119 3.75335
R5842 VDDA.n71 VDDA.n67 3.75335
R5843 VDDA.n70 VDDA.n69 3.75335
R5844 VDDA.n77 VDDA.n63 3.75335
R5845 VDDA.n79 VDDA.n78 3.75335
R5846 VDDA.n586 VDDA.n579 3.75335
R5847 VDDA.n581 VDDA.n535 3.75335
R5848 VDDA.n573 VDDA.n572 3.75335
R5849 VDDA.n568 VDDA.n545 3.75335
R5850 VDDA.n638 VDDA.n637 3.71013
R5851 VDDA.n476 VDDA.n475 3.43377
R5852 VDDA.n209 VDDA.n208 2.8957
R5853 VDDA.n210 VDDA.n209 2.8957
R5854 VDDA.n214 VDDA.n212 2.8957
R5855 VDDA.n217 VDDA.n212 2.8957
R5856 VDDA.n213 VDDA.n210 2.8957
R5857 VDDA.n217 VDDA.n216 2.8957
R5858 VDDA.n219 VDDA.n208 2.8957
R5859 VDDA.n214 VDDA.n213 2.8957
R5860 VDDA.n600 VDDA.n592 2.5005
R5861 VDDA.n219 VDDA.n207 2.32777
R5862 VDDA.n638 VDDA.n467 2.1343
R5863 VDDA VDDA.n638 2.0779
R5864 VDDA.n524 VDDA.n507 1.8755
R5865 VDDA.n565 VDDA.n550 1.84425
R5866 VDDA.n623 VDDA.n614 1.813
R5867 VDDA.n631 VDDA.n628 1.813
R5868 VDDA.n565 VDDA.n564 1.0005
R5869 VDDA.n564 VDDA.n562 1.0005
R5870 VDDA.n562 VDDA.n560 1.0005
R5871 VDDA.n560 VDDA.n558 1.0005
R5872 VDDA.n558 VDDA.n556 1.0005
R5873 VDDA.n556 VDDA.n554 1.0005
R5874 VDDA.n554 VDDA.n552 1.0005
R5875 VDDA.n552 VDDA.n534 1.0005
R5876 VDDA.n592 VDDA.n534 1.0005
R5877 VDDA.n466 VDDA.n421 0.938
R5878 VDDA.n205 VDDA.n204 0.922375
R5879 VDDA.n187 VDDA.n178 0.922375
R5880 VDDA.n232 VDDA.n178 0.922375
R5881 VDDA.n532 VDDA.n477 0.840625
R5882 VDDA.n601 VDDA.n532 0.74075
R5883 VDDA.n465 VDDA.n422 0.6255
R5884 VDDA.n420 VDDA.n415 0.6255
R5885 VDDA.n284 VDDA.n283 0.6255
R5886 VDDA.n283 VDDA.n281 0.6255
R5887 VDDA.n245 VDDA.n236 0.6255
R5888 VDDA.n284 VDDA.n236 0.6255
R5889 VDDA.n49 VDDA.n48 0.6255
R5890 VDDA.n48 VDDA.n46 0.6255
R5891 VDDA.n10 VDDA.n1 0.6255
R5892 VDDA.n49 VDDA.n1 0.6255
R5893 VDDA.n501 VDDA.n499 0.6255
R5894 VDDA.n499 VDDA.n497 0.6255
R5895 VDDA.n497 VDDA.n495 0.6255
R5896 VDDA.n495 VDDA.n493 0.6255
R5897 VDDA.n493 VDDA.n491 0.6255
R5898 VDDA.n491 VDDA.n489 0.6255
R5899 VDDA.n489 VDDA.n487 0.6255
R5900 VDDA.n487 VDDA.n484 0.6255
R5901 VDDA.n507 VDDA.n484 0.6255
R5902 VDDA.n524 VDDA.n523 0.6255
R5903 VDDA.n523 VDDA.n521 0.6255
R5904 VDDA.n521 VDDA.n519 0.6255
R5905 VDDA.n519 VDDA.n517 0.6255
R5906 VDDA.n517 VDDA.n515 0.6255
R5907 VDDA.n515 VDDA.n513 0.6255
R5908 VDDA.n513 VDDA.n511 0.6255
R5909 VDDA.n511 VDDA.n509 0.6255
R5910 VDDA.n509 VDDA.n479 0.6255
R5911 VDDA.n531 VDDA.n479 0.6255
R5912 VDDA.n344 VDDA.n342 0.563
R5913 VDDA.n342 VDDA.n340 0.563
R5914 VDDA.n340 VDDA.n338 0.563
R5915 VDDA.n338 VDDA.n322 0.563
R5916 VDDA.n410 VDDA.n322 0.563
R5917 VDDA.n291 VDDA.n289 0.563
R5918 VDDA.n293 VDDA.n291 0.563
R5919 VDDA.n295 VDDA.n293 0.563
R5920 VDDA.n297 VDDA.n295 0.563
R5921 VDDA.n104 VDDA.n102 0.563
R5922 VDDA.n102 VDDA.n100 0.563
R5923 VDDA.n100 VDDA.n98 0.563
R5924 VDDA.n98 VDDA.n87 0.563
R5925 VDDA.n175 VDDA.n87 0.563
R5926 VDDA.n56 VDDA.n54 0.563
R5927 VDDA.n58 VDDA.n56 0.563
R5928 VDDA.n60 VDDA.n58 0.563
R5929 VDDA.n62 VDDA.n60 0.563
R5930 VDDA.n609 VDDA.n607 0.563
R5931 VDDA.n614 VDDA.n607 0.563
R5932 VDDA.n623 VDDA.n622 0.563
R5933 VDDA.n622 VDDA.n620 0.563
R5934 VDDA.n620 VDDA.n618 0.563
R5935 VDDA.n618 VDDA.n616 0.563
R5936 VDDA.n616 VDDA.n605 0.563
R5937 VDDA.n628 VDDA.n605 0.563
R5938 VDDA.n631 VDDA.n630 0.563
R5939 VDDA.n630 VDDA.n603 0.563
R5940 VDDA.n636 VDDA.n603 0.563
R5941 VDDA.n233 VDDA.n176 0.46925
R5942 VDDA VDDA.n601 0.41175
R5943 VDDA.n205 VDDA.n187 0.3755
R5944 VDDA.t37 VDDA.t114 0.1603
R5945 VDDA.t23 VDDA.t63 0.1603
R5946 VDDA.t99 VDDA.t41 0.1603
R5947 VDDA.t206 VDDA.t189 0.1603
R5948 VDDA.t108 VDDA.t162 0.1603
R5949 VDDA.n469 VDDA.t163 0.159278
R5950 VDDA.n470 VDDA.t21 0.159278
R5951 VDDA.n471 VDDA.t43 0.159278
R5952 VDDA.n472 VDDA.t188 0.159278
R5953 VDDA.n472 VDDA.t107 0.1368
R5954 VDDA.n472 VDDA.t37 0.1368
R5955 VDDA.n471 VDDA.t42 0.1368
R5956 VDDA.n471 VDDA.t23 0.1368
R5957 VDDA.n470 VDDA.t100 0.1368
R5958 VDDA.n470 VDDA.t99 0.1368
R5959 VDDA.n469 VDDA.t34 0.1368
R5960 VDDA.n469 VDDA.t206 0.1368
R5961 VDDA.n468 VDDA.t22 0.1368
R5962 VDDA.n468 VDDA.t108 0.1368
R5963 VDDA.n637 VDDA 0.135625
R5964 VDDA.t163 VDDA.n468 0.00152174
R5965 VDDA.t21 VDDA.n469 0.00152174
R5966 VDDA.t43 VDDA.n470 0.00152174
R5967 VDDA.t188 VDDA.n471 0.00152174
R5968 VDDA.t115 VDDA.n472 0.00152174
R5969 bgr_0.V_TOP.n0 bgr_0.V_TOP.t29 369.534
R5970 bgr_0.V_TOP.n23 bgr_0.V_TOP.n21 339.961
R5971 bgr_0.V_TOP.n23 bgr_0.V_TOP.n22 339.272
R5972 bgr_0.V_TOP.n19 bgr_0.V_TOP.n18 339.272
R5973 bgr_0.V_TOP.n27 bgr_0.V_TOP.n26 339.272
R5974 bgr_0.V_TOP.n29 bgr_0.V_TOP.n28 339.272
R5975 bgr_0.V_TOP.n24 bgr_0.V_TOP.n20 334.772
R5976 bgr_0.V_TOP.n39 bgr_0.V_TOP.n38 224.934
R5977 bgr_0.V_TOP.n38 bgr_0.V_TOP.n37 224.934
R5978 bgr_0.V_TOP.n37 bgr_0.V_TOP.n36 224.934
R5979 bgr_0.V_TOP.n36 bgr_0.V_TOP.n35 224.934
R5980 bgr_0.V_TOP.n35 bgr_0.V_TOP.n34 224.934
R5981 bgr_0.V_TOP.n34 bgr_0.V_TOP.n33 224.934
R5982 bgr_0.V_TOP.n33 bgr_0.V_TOP.n32 224.934
R5983 bgr_0.V_TOP.n1 bgr_0.V_TOP.n0 224.934
R5984 bgr_0.V_TOP.n2 bgr_0.V_TOP.n1 224.934
R5985 bgr_0.V_TOP.n3 bgr_0.V_TOP.n2 224.934
R5986 bgr_0.V_TOP.n4 bgr_0.V_TOP.n3 224.934
R5987 bgr_0.V_TOP.n5 bgr_0.V_TOP.n4 224.934
R5988 bgr_0.V_TOP bgr_0.V_TOP.t48 214.222
R5989 bgr_0.V_TOP.n31 bgr_0.V_TOP.n30 163.175
R5990 bgr_0.V_TOP.n39 bgr_0.V_TOP.t24 144.601
R5991 bgr_0.V_TOP.n38 bgr_0.V_TOP.t33 144.601
R5992 bgr_0.V_TOP.n37 bgr_0.V_TOP.t39 144.601
R5993 bgr_0.V_TOP.n36 bgr_0.V_TOP.t16 144.601
R5994 bgr_0.V_TOP.n35 bgr_0.V_TOP.t15 144.601
R5995 bgr_0.V_TOP.n34 bgr_0.V_TOP.t28 144.601
R5996 bgr_0.V_TOP.n33 bgr_0.V_TOP.t38 144.601
R5997 bgr_0.V_TOP.n32 bgr_0.V_TOP.t14 144.601
R5998 bgr_0.V_TOP.n0 bgr_0.V_TOP.t30 144.601
R5999 bgr_0.V_TOP.n1 bgr_0.V_TOP.t18 144.601
R6000 bgr_0.V_TOP.n2 bgr_0.V_TOP.t46 144.601
R6001 bgr_0.V_TOP.n3 bgr_0.V_TOP.t37 144.601
R6002 bgr_0.V_TOP.n4 bgr_0.V_TOP.t26 144.601
R6003 bgr_0.V_TOP.n5 bgr_0.V_TOP.t27 144.601
R6004 bgr_0.V_TOP.n17 bgr_0.V_TOP.t3 108.424
R6005 bgr_0.V_TOP.n30 bgr_0.V_TOP.t7 95.4467
R6006 bgr_0.V_TOP bgr_0.V_TOP.n39 69.6227
R6007 bgr_0.V_TOP.n32 bgr_0.V_TOP.n31 69.6227
R6008 bgr_0.V_TOP.n31 bgr_0.V_TOP.n5 69.6227
R6009 bgr_0.V_TOP.n18 bgr_0.V_TOP.t8 39.4005
R6010 bgr_0.V_TOP.n18 bgr_0.V_TOP.t4 39.4005
R6011 bgr_0.V_TOP.n20 bgr_0.V_TOP.t5 39.4005
R6012 bgr_0.V_TOP.n20 bgr_0.V_TOP.t13 39.4005
R6013 bgr_0.V_TOP.n22 bgr_0.V_TOP.t2 39.4005
R6014 bgr_0.V_TOP.n22 bgr_0.V_TOP.t11 39.4005
R6015 bgr_0.V_TOP.n21 bgr_0.V_TOP.t10 39.4005
R6016 bgr_0.V_TOP.n21 bgr_0.V_TOP.t0 39.4005
R6017 bgr_0.V_TOP.n26 bgr_0.V_TOP.t6 39.4005
R6018 bgr_0.V_TOP.n26 bgr_0.V_TOP.t12 39.4005
R6019 bgr_0.V_TOP.n28 bgr_0.V_TOP.t1 39.4005
R6020 bgr_0.V_TOP.n28 bgr_0.V_TOP.t9 39.4005
R6021 bgr_0.V_TOP.n17 bgr_0.V_TOP.n16 37.1479
R6022 bgr_0.V_TOP.n19 bgr_0.V_TOP.n17 27.8371
R6023 bgr_0.V_TOP.n24 bgr_0.V_TOP.n23 8.313
R6024 bgr_0.V_TOP.n30 bgr_0.V_TOP.n29 5.188
R6025 bgr_0.V_TOP.n6 bgr_0.V_TOP.t31 4.8295
R6026 bgr_0.V_TOP.n7 bgr_0.V_TOP.t22 4.8295
R6027 bgr_0.V_TOP.n8 bgr_0.V_TOP.t20 4.8295
R6028 bgr_0.V_TOP.n9 bgr_0.V_TOP.t45 4.8295
R6029 bgr_0.V_TOP.n10 bgr_0.V_TOP.t42 4.8295
R6030 bgr_0.V_TOP.n11 bgr_0.V_TOP.t36 4.8295
R6031 bgr_0.V_TOP.n12 bgr_0.V_TOP.t17 4.8295
R6032 bgr_0.V_TOP.n13 bgr_0.V_TOP.t43 4.8295
R6033 bgr_0.V_TOP.n14 bgr_0.V_TOP.t34 4.8295
R6034 bgr_0.V_TOP.n6 bgr_0.V_TOP.t35 4.5005
R6035 bgr_0.V_TOP.n7 bgr_0.V_TOP.t32 4.5005
R6036 bgr_0.V_TOP.n8 bgr_0.V_TOP.t25 4.5005
R6037 bgr_0.V_TOP.n9 bgr_0.V_TOP.t21 4.5005
R6038 bgr_0.V_TOP.n10 bgr_0.V_TOP.t49 4.5005
R6039 bgr_0.V_TOP.n11 bgr_0.V_TOP.t44 4.5005
R6040 bgr_0.V_TOP.n12 bgr_0.V_TOP.t23 4.5005
R6041 bgr_0.V_TOP.n13 bgr_0.V_TOP.t19 4.5005
R6042 bgr_0.V_TOP.n16 bgr_0.V_TOP.t40 4.5005
R6043 bgr_0.V_TOP.n15 bgr_0.V_TOP.t47 4.5005
R6044 bgr_0.V_TOP.n14 bgr_0.V_TOP.t41 4.5005
R6045 bgr_0.V_TOP.n25 bgr_0.V_TOP.n24 4.5005
R6046 bgr_0.V_TOP.n29 bgr_0.V_TOP.n27 2.1255
R6047 bgr_0.V_TOP.n27 bgr_0.V_TOP.n25 2.1255
R6048 bgr_0.V_TOP.n25 bgr_0.V_TOP.n19 2.1255
R6049 bgr_0.V_TOP.n7 bgr_0.V_TOP.n6 0.3295
R6050 bgr_0.V_TOP.n9 bgr_0.V_TOP.n8 0.3295
R6051 bgr_0.V_TOP.n11 bgr_0.V_TOP.n10 0.3295
R6052 bgr_0.V_TOP.n13 bgr_0.V_TOP.n12 0.3295
R6053 bgr_0.V_TOP.n16 bgr_0.V_TOP.n15 0.3295
R6054 bgr_0.V_TOP.n15 bgr_0.V_TOP.n14 0.3295
R6055 bgr_0.V_TOP.n9 bgr_0.V_TOP.n7 0.2825
R6056 bgr_0.V_TOP.n11 bgr_0.V_TOP.n9 0.2825
R6057 bgr_0.V_TOP.n13 bgr_0.V_TOP.n11 0.2825
R6058 bgr_0.V_TOP.n14 bgr_0.V_TOP.n13 0.2825
R6059 VOUT-.n8 VOUT-.n0 149.19
R6060 VOUT-.n3 VOUT-.n1 149.19
R6061 VOUT-.n7 VOUT-.n6 148.626
R6062 VOUT-.n5 VOUT-.n4 148.626
R6063 VOUT-.n3 VOUT-.n2 148.626
R6064 VOUT-.n10 VOUT-.n9 144.126
R6065 VOUT-.n91 VOUT-.t16 112.184
R6066 VOUT-.n88 VOUT-.n86 98.9303
R6067 VOUT-.n90 VOUT-.n89 97.8053
R6068 VOUT-.n88 VOUT-.n87 97.8053
R6069 VOUT-.n85 VOUT-.n10 15.5682
R6070 VOUT-.n85 VOUT-.n84 11.5649
R6071 VOUT- VOUT-.n85 9.46925
R6072 VOUT-.n9 VOUT-.t9 6.56717
R6073 VOUT-.n9 VOUT-.t5 6.56717
R6074 VOUT-.n6 VOUT-.t4 6.56717
R6075 VOUT-.n6 VOUT-.t3 6.56717
R6076 VOUT-.n4 VOUT-.t7 6.56717
R6077 VOUT-.n4 VOUT-.t1 6.56717
R6078 VOUT-.n2 VOUT-.t8 6.56717
R6079 VOUT-.n2 VOUT-.t0 6.56717
R6080 VOUT-.n1 VOUT-.t2 6.56717
R6081 VOUT-.n1 VOUT-.t15 6.56717
R6082 VOUT-.n0 VOUT-.t14 6.56717
R6083 VOUT-.n0 VOUT-.t6 6.56717
R6084 VOUT-.n39 VOUT-.t68 4.8295
R6085 VOUT-.n47 VOUT-.t66 4.8295
R6086 VOUT-.n45 VOUT-.t115 4.8295
R6087 VOUT-.n43 VOUT-.t150 4.8295
R6088 VOUT-.n42 VOUT-.t132 4.8295
R6089 VOUT-.n41 VOUT-.t29 4.8295
R6090 VOUT-.n59 VOUT-.t125 4.8295
R6091 VOUT-.n60 VOUT-.t73 4.8295
R6092 VOUT-.n61 VOUT-.t23 4.8295
R6093 VOUT-.n62 VOUT-.t109 4.8295
R6094 VOUT-.n63 VOUT-.t76 4.8295
R6095 VOUT-.n64 VOUT-.t44 4.8295
R6096 VOUT-.n66 VOUT-.t37 4.8295
R6097 VOUT-.n67 VOUT-.t143 4.8295
R6098 VOUT-.n69 VOUT-.t70 4.8295
R6099 VOUT-.n70 VOUT-.t39 4.8295
R6100 VOUT-.n72 VOUT-.t32 4.8295
R6101 VOUT-.n73 VOUT-.t138 4.8295
R6102 VOUT-.n75 VOUT-.t131 4.8295
R6103 VOUT-.n76 VOUT-.t101 4.8295
R6104 VOUT-.n78 VOUT-.t28 4.8295
R6105 VOUT-.n79 VOUT-.t133 4.8295
R6106 VOUT-.n11 VOUT-.t26 4.8295
R6107 VOUT-.n13 VOUT-.t36 4.8295
R6108 VOUT-.n24 VOUT-.t140 4.8295
R6109 VOUT-.n25 VOUT-.t111 4.8295
R6110 VOUT-.n27 VOUT-.t41 4.8295
R6111 VOUT-.n28 VOUT-.t151 4.8295
R6112 VOUT-.n30 VOUT-.t80 4.8295
R6113 VOUT-.n31 VOUT-.t51 4.8295
R6114 VOUT-.n33 VOUT-.t49 4.8295
R6115 VOUT-.n34 VOUT-.t19 4.8295
R6116 VOUT-.n36 VOUT-.t85 4.8295
R6117 VOUT-.n37 VOUT-.t55 4.8295
R6118 VOUT-.n81 VOUT-.t124 4.8295
R6119 VOUT-.n49 VOUT-.t91 4.8154
R6120 VOUT-.n50 VOUT-.t69 4.8154
R6121 VOUT-.n51 VOUT-.t107 4.8154
R6122 VOUT-.n49 VOUT-.t31 4.806
R6123 VOUT-.n50 VOUT-.t149 4.806
R6124 VOUT-.n51 VOUT-.t50 4.806
R6125 VOUT-.n52 VOUT-.t144 4.806
R6126 VOUT-.n52 VOUT-.t83 4.806
R6127 VOUT-.n53 VOUT-.t120 4.806
R6128 VOUT-.n54 VOUT-.t104 4.806
R6129 VOUT-.n55 VOUT-.t137 4.806
R6130 VOUT-.n56 VOUT-.t35 4.806
R6131 VOUT-.n57 VOUT-.t156 4.806
R6132 VOUT-.n14 VOUT-.t71 4.806
R6133 VOUT-.n14 VOUT-.t113 4.806
R6134 VOUT-.n15 VOUT-.t114 4.806
R6135 VOUT-.n15 VOUT-.t24 4.806
R6136 VOUT-.n16 VOUT-.t65 4.806
R6137 VOUT-.n16 VOUT-.t62 4.806
R6138 VOUT-.n17 VOUT-.t154 4.806
R6139 VOUT-.n17 VOUT-.t95 4.806
R6140 VOUT-.n18 VOUT-.t105 4.806
R6141 VOUT-.n18 VOUT-.t126 4.806
R6142 VOUT-.n19 VOUT-.t141 4.806
R6143 VOUT-.n19 VOUT-.t38 4.806
R6144 VOUT-.n20 VOUT-.t92 4.806
R6145 VOUT-.n20 VOUT-.t74 4.806
R6146 VOUT-.n21 VOUT-.t42 4.806
R6147 VOUT-.n22 VOUT-.t82 4.806
R6148 VOUT-.n39 VOUT-.t86 4.5005
R6149 VOUT-.n40 VOUT-.t54 4.5005
R6150 VOUT-.n47 VOUT-.t77 4.5005
R6151 VOUT-.n48 VOUT-.t43 4.5005
R6152 VOUT-.n45 VOUT-.t58 4.5005
R6153 VOUT-.n46 VOUT-.t22 4.5005
R6154 VOUT-.n43 VOUT-.t94 4.5005
R6155 VOUT-.n44 VOUT-.t61 4.5005
R6156 VOUT-.n42 VOUT-.t99 4.5005
R6157 VOUT-.n41 VOUT-.t52 4.5005
R6158 VOUT-.n58 VOUT-.t155 4.5005
R6159 VOUT-.n57 VOUT-.t116 4.5005
R6160 VOUT-.n56 VOUT-.t136 4.5005
R6161 VOUT-.n55 VOUT-.t100 4.5005
R6162 VOUT-.n54 VOUT-.t64 4.5005
R6163 VOUT-.n53 VOUT-.t81 4.5005
R6164 VOUT-.n52 VOUT-.t45 4.5005
R6165 VOUT-.n51 VOUT-.t146 4.5005
R6166 VOUT-.n50 VOUT-.t108 4.5005
R6167 VOUT-.n49 VOUT-.t130 4.5005
R6168 VOUT-.n59 VOUT-.t152 4.5005
R6169 VOUT-.n60 VOUT-.t112 4.5005
R6170 VOUT-.n61 VOUT-.t47 4.5005
R6171 VOUT-.n62 VOUT-.t147 4.5005
R6172 VOUT-.n63 VOUT-.t27 4.5005
R6173 VOUT-.n65 VOUT-.t128 4.5005
R6174 VOUT-.n64 VOUT-.t97 4.5005
R6175 VOUT-.n66 VOUT-.t123 4.5005
R6176 VOUT-.n68 VOUT-.t88 4.5005
R6177 VOUT-.n67 VOUT-.t57 4.5005
R6178 VOUT-.n69 VOUT-.t20 4.5005
R6179 VOUT-.n71 VOUT-.t121 4.5005
R6180 VOUT-.n70 VOUT-.t87 4.5005
R6181 VOUT-.n72 VOUT-.t118 4.5005
R6182 VOUT-.n74 VOUT-.t84 4.5005
R6183 VOUT-.n73 VOUT-.t53 4.5005
R6184 VOUT-.n75 VOUT-.t79 4.5005
R6185 VOUT-.n77 VOUT-.t48 4.5005
R6186 VOUT-.n76 VOUT-.t153 4.5005
R6187 VOUT-.n78 VOUT-.t117 4.5005
R6188 VOUT-.n80 VOUT-.t78 4.5005
R6189 VOUT-.n79 VOUT-.t46 4.5005
R6190 VOUT-.n11 VOUT-.t119 4.5005
R6191 VOUT-.n12 VOUT-.t33 4.5005
R6192 VOUT-.n13 VOUT-.t122 4.5005
R6193 VOUT-.n23 VOUT-.t90 4.5005
R6194 VOUT-.n22 VOUT-.t56 4.5005
R6195 VOUT-.n21 VOUT-.t142 4.5005
R6196 VOUT-.n20 VOUT-.t110 4.5005
R6197 VOUT-.n19 VOUT-.t72 4.5005
R6198 VOUT-.n18 VOUT-.t25 4.5005
R6199 VOUT-.n17 VOUT-.t127 4.5005
R6200 VOUT-.n16 VOUT-.t93 4.5005
R6201 VOUT-.n15 VOUT-.t60 4.5005
R6202 VOUT-.n14 VOUT-.t148 4.5005
R6203 VOUT-.n24 VOUT-.t89 4.5005
R6204 VOUT-.n26 VOUT-.t59 4.5005
R6205 VOUT-.n25 VOUT-.t21 4.5005
R6206 VOUT-.n27 VOUT-.t129 4.5005
R6207 VOUT-.n29 VOUT-.t98 4.5005
R6208 VOUT-.n28 VOUT-.t63 4.5005
R6209 VOUT-.n30 VOUT-.t30 4.5005
R6210 VOUT-.n32 VOUT-.t134 4.5005
R6211 VOUT-.n31 VOUT-.t103 4.5005
R6212 VOUT-.n33 VOUT-.t135 4.5005
R6213 VOUT-.n35 VOUT-.t102 4.5005
R6214 VOUT-.n34 VOUT-.t67 4.5005
R6215 VOUT-.n36 VOUT-.t34 4.5005
R6216 VOUT-.n38 VOUT-.t139 4.5005
R6217 VOUT-.n37 VOUT-.t106 4.5005
R6218 VOUT-.n81 VOUT-.t75 4.5005
R6219 VOUT-.n82 VOUT-.t40 4.5005
R6220 VOUT-.n83 VOUT-.t145 4.5005
R6221 VOUT-.n84 VOUT-.t96 4.5005
R6222 VOUT-.n10 VOUT-.n8 4.5005
R6223 VOUT-.n89 VOUT-.t13 3.42907
R6224 VOUT-.n89 VOUT-.t11 3.42907
R6225 VOUT-.n87 VOUT-.t18 3.42907
R6226 VOUT-.n87 VOUT-.t10 3.42907
R6227 VOUT-.n86 VOUT-.t17 3.42907
R6228 VOUT-.n86 VOUT-.t12 3.42907
R6229 VOUT-.n91 VOUT-.n90 1.30519
R6230 VOUT- VOUT-.n91 1.24269
R6231 VOUT-.n90 VOUT-.n88 1.1255
R6232 VOUT-.n5 VOUT-.n3 0.563
R6233 VOUT-.n7 VOUT-.n5 0.563
R6234 VOUT-.n8 VOUT-.n7 0.563
R6235 VOUT-.n40 VOUT-.n39 0.3295
R6236 VOUT-.n48 VOUT-.n47 0.3295
R6237 VOUT-.n46 VOUT-.n45 0.3295
R6238 VOUT-.n44 VOUT-.n43 0.3295
R6239 VOUT-.n58 VOUT-.n41 0.3295
R6240 VOUT-.n58 VOUT-.n57 0.3295
R6241 VOUT-.n57 VOUT-.n56 0.3295
R6242 VOUT-.n56 VOUT-.n55 0.3295
R6243 VOUT-.n55 VOUT-.n54 0.3295
R6244 VOUT-.n54 VOUT-.n53 0.3295
R6245 VOUT-.n53 VOUT-.n52 0.3295
R6246 VOUT-.n52 VOUT-.n51 0.3295
R6247 VOUT-.n51 VOUT-.n50 0.3295
R6248 VOUT-.n50 VOUT-.n49 0.3295
R6249 VOUT-.n60 VOUT-.n59 0.3295
R6250 VOUT-.n62 VOUT-.n61 0.3295
R6251 VOUT-.n65 VOUT-.n63 0.3295
R6252 VOUT-.n65 VOUT-.n64 0.3295
R6253 VOUT-.n68 VOUT-.n66 0.3295
R6254 VOUT-.n68 VOUT-.n67 0.3295
R6255 VOUT-.n71 VOUT-.n69 0.3295
R6256 VOUT-.n71 VOUT-.n70 0.3295
R6257 VOUT-.n74 VOUT-.n72 0.3295
R6258 VOUT-.n74 VOUT-.n73 0.3295
R6259 VOUT-.n77 VOUT-.n75 0.3295
R6260 VOUT-.n77 VOUT-.n76 0.3295
R6261 VOUT-.n80 VOUT-.n78 0.3295
R6262 VOUT-.n80 VOUT-.n79 0.3295
R6263 VOUT-.n12 VOUT-.n11 0.3295
R6264 VOUT-.n23 VOUT-.n13 0.3295
R6265 VOUT-.n23 VOUT-.n22 0.3295
R6266 VOUT-.n22 VOUT-.n21 0.3295
R6267 VOUT-.n21 VOUT-.n20 0.3295
R6268 VOUT-.n20 VOUT-.n19 0.3295
R6269 VOUT-.n19 VOUT-.n18 0.3295
R6270 VOUT-.n18 VOUT-.n17 0.3295
R6271 VOUT-.n17 VOUT-.n16 0.3295
R6272 VOUT-.n16 VOUT-.n15 0.3295
R6273 VOUT-.n15 VOUT-.n14 0.3295
R6274 VOUT-.n26 VOUT-.n24 0.3295
R6275 VOUT-.n26 VOUT-.n25 0.3295
R6276 VOUT-.n29 VOUT-.n27 0.3295
R6277 VOUT-.n29 VOUT-.n28 0.3295
R6278 VOUT-.n32 VOUT-.n30 0.3295
R6279 VOUT-.n32 VOUT-.n31 0.3295
R6280 VOUT-.n35 VOUT-.n33 0.3295
R6281 VOUT-.n35 VOUT-.n34 0.3295
R6282 VOUT-.n38 VOUT-.n36 0.3295
R6283 VOUT-.n38 VOUT-.n37 0.3295
R6284 VOUT-.n82 VOUT-.n81 0.3295
R6285 VOUT-.n83 VOUT-.n82 0.3295
R6286 VOUT-.n84 VOUT-.n83 0.3295
R6287 VOUT-.n53 VOUT-.n48 0.306
R6288 VOUT-.n54 VOUT-.n46 0.306
R6289 VOUT-.n55 VOUT-.n44 0.306
R6290 VOUT-.n56 VOUT-.n42 0.306
R6291 VOUT-.n58 VOUT-.n40 0.2825
R6292 VOUT-.n60 VOUT-.n58 0.2825
R6293 VOUT-.n62 VOUT-.n60 0.2825
R6294 VOUT-.n65 VOUT-.n62 0.2825
R6295 VOUT-.n68 VOUT-.n65 0.2825
R6296 VOUT-.n71 VOUT-.n68 0.2825
R6297 VOUT-.n74 VOUT-.n71 0.2825
R6298 VOUT-.n77 VOUT-.n74 0.2825
R6299 VOUT-.n80 VOUT-.n77 0.2825
R6300 VOUT-.n23 VOUT-.n12 0.2825
R6301 VOUT-.n26 VOUT-.n23 0.2825
R6302 VOUT-.n29 VOUT-.n26 0.2825
R6303 VOUT-.n32 VOUT-.n29 0.2825
R6304 VOUT-.n35 VOUT-.n32 0.2825
R6305 VOUT-.n38 VOUT-.n35 0.2825
R6306 VOUT-.n82 VOUT-.n38 0.2825
R6307 VOUT-.n82 VOUT-.n80 0.2825
R6308 two_stage_opamp_dummy_magic_16_0.cap_res_X two_stage_opamp_dummy_magic_16_0.cap_res_X.t0 49.197
R6309 two_stage_opamp_dummy_magic_16_0.cap_res_X two_stage_opamp_dummy_magic_16_0.cap_res_X.t7 0.87
R6310 two_stage_opamp_dummy_magic_16_0.cap_res_X.t27 two_stage_opamp_dummy_magic_16_0.cap_res_X.t66 0.1603
R6311 two_stage_opamp_dummy_magic_16_0.cap_res_X.t49 two_stage_opamp_dummy_magic_16_0.cap_res_X.t88 0.1603
R6312 two_stage_opamp_dummy_magic_16_0.cap_res_X.t11 two_stage_opamp_dummy_magic_16_0.cap_res_X.t50 0.1603
R6313 two_stage_opamp_dummy_magic_16_0.cap_res_X.t112 two_stage_opamp_dummy_magic_16_0.cap_res_X.t13 0.1603
R6314 two_stage_opamp_dummy_magic_16_0.cap_res_X.t80 two_stage_opamp_dummy_magic_16_0.cap_res_X.t91 0.1603
R6315 two_stage_opamp_dummy_magic_16_0.cap_res_X.t114 two_stage_opamp_dummy_magic_16_0.cap_res_X.t80 0.1603
R6316 two_stage_opamp_dummy_magic_16_0.cap_res_X.t76 two_stage_opamp_dummy_magic_16_0.cap_res_X.t114 0.1603
R6317 two_stage_opamp_dummy_magic_16_0.cap_res_X.t99 two_stage_opamp_dummy_magic_16_0.cap_res_X.t42 0.1603
R6318 two_stage_opamp_dummy_magic_16_0.cap_res_X.t135 two_stage_opamp_dummy_magic_16_0.cap_res_X.t99 0.1603
R6319 two_stage_opamp_dummy_magic_16_0.cap_res_X.t93 two_stage_opamp_dummy_magic_16_0.cap_res_X.t135 0.1603
R6320 two_stage_opamp_dummy_magic_16_0.cap_res_X.t105 two_stage_opamp_dummy_magic_16_0.cap_res_X.t128 0.1603
R6321 two_stage_opamp_dummy_magic_16_0.cap_res_X.t71 two_stage_opamp_dummy_magic_16_0.cap_res_X.t89 0.1603
R6322 two_stage_opamp_dummy_magic_16_0.cap_res_X.t5 two_stage_opamp_dummy_magic_16_0.cap_res_X.t32 0.1603
R6323 two_stage_opamp_dummy_magic_16_0.cap_res_X.t110 two_stage_opamp_dummy_magic_16_0.cap_res_X.t134 0.1603
R6324 two_stage_opamp_dummy_magic_16_0.cap_res_X.t60 two_stage_opamp_dummy_magic_16_0.cap_res_X.t113 0.1603
R6325 two_stage_opamp_dummy_magic_16_0.cap_res_X.t130 two_stage_opamp_dummy_magic_16_0.cap_res_X.t81 0.1603
R6326 two_stage_opamp_dummy_magic_16_0.cap_res_X.t100 two_stage_opamp_dummy_magic_16_0.cap_res_X.t14 0.1603
R6327 two_stage_opamp_dummy_magic_16_0.cap_res_X.t34 two_stage_opamp_dummy_magic_16_0.cap_res_X.t120 0.1603
R6328 two_stage_opamp_dummy_magic_16_0.cap_res_X.t70 two_stage_opamp_dummy_magic_16_0.cap_res_X.t118 0.1603
R6329 two_stage_opamp_dummy_magic_16_0.cap_res_X.t137 two_stage_opamp_dummy_magic_16_0.cap_res_X.t87 0.1603
R6330 two_stage_opamp_dummy_magic_16_0.cap_res_X.t104 two_stage_opamp_dummy_magic_16_0.cap_res_X.t19 0.1603
R6331 two_stage_opamp_dummy_magic_16_0.cap_res_X.t39 two_stage_opamp_dummy_magic_16_0.cap_res_X.t125 0.1603
R6332 two_stage_opamp_dummy_magic_16_0.cap_res_X.t4 two_stage_opamp_dummy_magic_16_0.cap_res_X.t56 0.1603
R6333 two_stage_opamp_dummy_magic_16_0.cap_res_X.t78 two_stage_opamp_dummy_magic_16_0.cap_res_X.t26 0.1603
R6334 two_stage_opamp_dummy_magic_16_0.cap_res_X.t111 two_stage_opamp_dummy_magic_16_0.cap_res_X.t24 0.1603
R6335 two_stage_opamp_dummy_magic_16_0.cap_res_X.t40 two_stage_opamp_dummy_magic_16_0.cap_res_X.t129 0.1603
R6336 two_stage_opamp_dummy_magic_16_0.cap_res_X.t12 two_stage_opamp_dummy_magic_16_0.cap_res_X.t61 0.1603
R6337 two_stage_opamp_dummy_magic_16_0.cap_res_X.t82 two_stage_opamp_dummy_magic_16_0.cap_res_X.t33 0.1603
R6338 two_stage_opamp_dummy_magic_16_0.cap_res_X.t51 two_stage_opamp_dummy_magic_16_0.cap_res_X.t102 0.1603
R6339 two_stage_opamp_dummy_magic_16_0.cap_res_X.t123 two_stage_opamp_dummy_magic_16_0.cap_res_X.t72 0.1603
R6340 two_stage_opamp_dummy_magic_16_0.cap_res_X.t90 two_stage_opamp_dummy_magic_16_0.cap_res_X.t138 0.1603
R6341 two_stage_opamp_dummy_magic_16_0.cap_res_X.t22 two_stage_opamp_dummy_magic_16_0.cap_res_X.t108 0.1603
R6342 two_stage_opamp_dummy_magic_16_0.cap_res_X.t54 two_stage_opamp_dummy_magic_16_0.cap_res_X.t106 0.1603
R6343 two_stage_opamp_dummy_magic_16_0.cap_res_X.t127 two_stage_opamp_dummy_magic_16_0.cap_res_X.t77 0.1603
R6344 two_stage_opamp_dummy_magic_16_0.cap_res_X.t94 two_stage_opamp_dummy_magic_16_0.cap_res_X.t6 0.1603
R6345 two_stage_opamp_dummy_magic_16_0.cap_res_X.t28 two_stage_opamp_dummy_magic_16_0.cap_res_X.t116 0.1603
R6346 two_stage_opamp_dummy_magic_16_0.cap_res_X.t136 two_stage_opamp_dummy_magic_16_0.cap_res_X.t46 0.1603
R6347 two_stage_opamp_dummy_magic_16_0.cap_res_X.t68 two_stage_opamp_dummy_magic_16_0.cap_res_X.t17 0.1603
R6348 two_stage_opamp_dummy_magic_16_0.cap_res_X.t9 two_stage_opamp_dummy_magic_16_0.cap_res_X.t86 0.1603
R6349 two_stage_opamp_dummy_magic_16_0.cap_res_X.t97 two_stage_opamp_dummy_magic_16_0.cap_res_X.t43 0.1603
R6350 two_stage_opamp_dummy_magic_16_0.cap_res_X.t64 two_stage_opamp_dummy_magic_16_0.cap_res_X.t92 0.1603
R6351 two_stage_opamp_dummy_magic_16_0.cap_res_X.t30 two_stage_opamp_dummy_magic_16_0.cap_res_X.t3 0.1603
R6352 two_stage_opamp_dummy_magic_16_0.cap_res_X.t132 two_stage_opamp_dummy_magic_16_0.cap_res_X.t52 0.1603
R6353 two_stage_opamp_dummy_magic_16_0.cap_res_X.t85 two_stage_opamp_dummy_magic_16_0.cap_res_X.t16 0.1603
R6354 two_stage_opamp_dummy_magic_16_0.cap_res_X.t47 two_stage_opamp_dummy_magic_16_0.cap_res_X.t65 0.1603
R6355 two_stage_opamp_dummy_magic_16_0.cap_res_X.t15 two_stage_opamp_dummy_magic_16_0.cap_res_X.t115 0.1603
R6356 two_stage_opamp_dummy_magic_16_0.cap_res_X.t101 two_stage_opamp_dummy_magic_16_0.cap_res_X.t75 0.1603
R6357 two_stage_opamp_dummy_magic_16_0.cap_res_X.t35 two_stage_opamp_dummy_magic_16_0.cap_res_X.t121 0.1603
R6358 two_stage_opamp_dummy_magic_16_0.cap_res_X.t38 two_stage_opamp_dummy_magic_16_0.cap_res_X.t131 0.1603
R6359 two_stage_opamp_dummy_magic_16_0.cap_res_X.t58 two_stage_opamp_dummy_magic_16_0.cap_res_X.t25 0.1603
R6360 two_stage_opamp_dummy_magic_16_0.cap_res_X.t21 two_stage_opamp_dummy_magic_16_0.cap_res_X.t58 0.1603
R6361 two_stage_opamp_dummy_magic_16_0.cap_res_X.t96 two_stage_opamp_dummy_magic_16_0.cap_res_X.t57 0.1603
R6362 two_stage_opamp_dummy_magic_16_0.cap_res_X.t63 two_stage_opamp_dummy_magic_16_0.cap_res_X.t96 0.1603
R6363 two_stage_opamp_dummy_magic_16_0.cap_res_X.t7 two_stage_opamp_dummy_magic_16_0.cap_res_X.t63 0.1603
R6364 two_stage_opamp_dummy_magic_16_0.cap_res_X.n28 two_stage_opamp_dummy_magic_16_0.cap_res_X.t126 0.159278
R6365 two_stage_opamp_dummy_magic_16_0.cap_res_X.n29 two_stage_opamp_dummy_magic_16_0.cap_res_X.t8 0.159278
R6366 two_stage_opamp_dummy_magic_16_0.cap_res_X.n30 two_stage_opamp_dummy_magic_16_0.cap_res_X.t107 0.159278
R6367 two_stage_opamp_dummy_magic_16_0.cap_res_X.n31 two_stage_opamp_dummy_magic_16_0.cap_res_X.t74 0.159278
R6368 two_stage_opamp_dummy_magic_16_0.cap_res_X.n32 two_stage_opamp_dummy_magic_16_0.cap_res_X.t37 0.159278
R6369 two_stage_opamp_dummy_magic_16_0.cap_res_X.n33 two_stage_opamp_dummy_magic_16_0.cap_res_X.t53 0.159278
R6370 two_stage_opamp_dummy_magic_16_0.cap_res_X.n25 two_stage_opamp_dummy_magic_16_0.cap_res_X.t103 0.159278
R6371 two_stage_opamp_dummy_magic_16_0.cap_res_X.n0 two_stage_opamp_dummy_magic_16_0.cap_res_X.t44 0.159278
R6372 two_stage_opamp_dummy_magic_16_0.cap_res_X.n1 two_stage_opamp_dummy_magic_16_0.cap_res_X.t133 0.159278
R6373 two_stage_opamp_dummy_magic_16_0.cap_res_X.n2 two_stage_opamp_dummy_magic_16_0.cap_res_X.t95 0.159278
R6374 two_stage_opamp_dummy_magic_16_0.cap_res_X.n3 two_stage_opamp_dummy_magic_16_0.cap_res_X.t62 0.159278
R6375 two_stage_opamp_dummy_magic_16_0.cap_res_X.n4 two_stage_opamp_dummy_magic_16_0.cap_res_X.t31 0.159278
R6376 two_stage_opamp_dummy_magic_16_0.cap_res_X.n5 two_stage_opamp_dummy_magic_16_0.cap_res_X.t119 0.159278
R6377 two_stage_opamp_dummy_magic_16_0.cap_res_X.n6 two_stage_opamp_dummy_magic_16_0.cap_res_X.t83 0.159278
R6378 two_stage_opamp_dummy_magic_16_0.cap_res_X.t67 two_stage_opamp_dummy_magic_16_0.cap_res_X.n9 0.159278
R6379 two_stage_opamp_dummy_magic_16_0.cap_res_X.t98 two_stage_opamp_dummy_magic_16_0.cap_res_X.n10 0.159278
R6380 two_stage_opamp_dummy_magic_16_0.cap_res_X.t59 two_stage_opamp_dummy_magic_16_0.cap_res_X.n11 0.159278
R6381 two_stage_opamp_dummy_magic_16_0.cap_res_X.t23 two_stage_opamp_dummy_magic_16_0.cap_res_X.n12 0.159278
R6382 two_stage_opamp_dummy_magic_16_0.cap_res_X.t55 two_stage_opamp_dummy_magic_16_0.cap_res_X.n13 0.159278
R6383 two_stage_opamp_dummy_magic_16_0.cap_res_X.t18 two_stage_opamp_dummy_magic_16_0.cap_res_X.n14 0.159278
R6384 two_stage_opamp_dummy_magic_16_0.cap_res_X.t117 two_stage_opamp_dummy_magic_16_0.cap_res_X.n15 0.159278
R6385 two_stage_opamp_dummy_magic_16_0.cap_res_X.t79 two_stage_opamp_dummy_magic_16_0.cap_res_X.n16 0.159278
R6386 two_stage_opamp_dummy_magic_16_0.cap_res_X.t109 two_stage_opamp_dummy_magic_16_0.cap_res_X.n17 0.159278
R6387 two_stage_opamp_dummy_magic_16_0.cap_res_X.t73 two_stage_opamp_dummy_magic_16_0.cap_res_X.n18 0.159278
R6388 two_stage_opamp_dummy_magic_16_0.cap_res_X.t36 two_stage_opamp_dummy_magic_16_0.cap_res_X.n19 0.159278
R6389 two_stage_opamp_dummy_magic_16_0.cap_res_X.t69 two_stage_opamp_dummy_magic_16_0.cap_res_X.n20 0.159278
R6390 two_stage_opamp_dummy_magic_16_0.cap_res_X.t29 two_stage_opamp_dummy_magic_16_0.cap_res_X.n21 0.159278
R6391 two_stage_opamp_dummy_magic_16_0.cap_res_X.t10 two_stage_opamp_dummy_magic_16_0.cap_res_X.n22 0.159278
R6392 two_stage_opamp_dummy_magic_16_0.cap_res_X.t45 two_stage_opamp_dummy_magic_16_0.cap_res_X.n23 0.159278
R6393 two_stage_opamp_dummy_magic_16_0.cap_res_X.t2 two_stage_opamp_dummy_magic_16_0.cap_res_X.n24 0.159278
R6394 two_stage_opamp_dummy_magic_16_0.cap_res_X.n26 two_stage_opamp_dummy_magic_16_0.cap_res_X.t1 0.159278
R6395 two_stage_opamp_dummy_magic_16_0.cap_res_X.n27 two_stage_opamp_dummy_magic_16_0.cap_res_X.t122 0.159278
R6396 two_stage_opamp_dummy_magic_16_0.cap_res_X.n34 two_stage_opamp_dummy_magic_16_0.cap_res_X.t20 0.159278
R6397 two_stage_opamp_dummy_magic_16_0.cap_res_X.t103 two_stage_opamp_dummy_magic_16_0.cap_res_X.t71 0.137822
R6398 two_stage_opamp_dummy_magic_16_0.cap_res_X.n25 two_stage_opamp_dummy_magic_16_0.cap_res_X.t105 0.1368
R6399 two_stage_opamp_dummy_magic_16_0.cap_res_X.n24 two_stage_opamp_dummy_magic_16_0.cap_res_X.t84 0.1368
R6400 two_stage_opamp_dummy_magic_16_0.cap_res_X.n24 two_stage_opamp_dummy_magic_16_0.cap_res_X.t5 0.1368
R6401 two_stage_opamp_dummy_magic_16_0.cap_res_X.n23 two_stage_opamp_dummy_magic_16_0.cap_res_X.t48 0.1368
R6402 two_stage_opamp_dummy_magic_16_0.cap_res_X.n23 two_stage_opamp_dummy_magic_16_0.cap_res_X.t110 0.1368
R6403 two_stage_opamp_dummy_magic_16_0.cap_res_X.n22 two_stage_opamp_dummy_magic_16_0.cap_res_X.t60 0.1368
R6404 two_stage_opamp_dummy_magic_16_0.cap_res_X.n22 two_stage_opamp_dummy_magic_16_0.cap_res_X.t130 0.1368
R6405 two_stage_opamp_dummy_magic_16_0.cap_res_X.n21 two_stage_opamp_dummy_magic_16_0.cap_res_X.t100 0.1368
R6406 two_stage_opamp_dummy_magic_16_0.cap_res_X.n21 two_stage_opamp_dummy_magic_16_0.cap_res_X.t34 0.1368
R6407 two_stage_opamp_dummy_magic_16_0.cap_res_X.n20 two_stage_opamp_dummy_magic_16_0.cap_res_X.t70 0.1368
R6408 two_stage_opamp_dummy_magic_16_0.cap_res_X.n20 two_stage_opamp_dummy_magic_16_0.cap_res_X.t137 0.1368
R6409 two_stage_opamp_dummy_magic_16_0.cap_res_X.n19 two_stage_opamp_dummy_magic_16_0.cap_res_X.t104 0.1368
R6410 two_stage_opamp_dummy_magic_16_0.cap_res_X.n19 two_stage_opamp_dummy_magic_16_0.cap_res_X.t39 0.1368
R6411 two_stage_opamp_dummy_magic_16_0.cap_res_X.n18 two_stage_opamp_dummy_magic_16_0.cap_res_X.t4 0.1368
R6412 two_stage_opamp_dummy_magic_16_0.cap_res_X.n18 two_stage_opamp_dummy_magic_16_0.cap_res_X.t78 0.1368
R6413 two_stage_opamp_dummy_magic_16_0.cap_res_X.n17 two_stage_opamp_dummy_magic_16_0.cap_res_X.t111 0.1368
R6414 two_stage_opamp_dummy_magic_16_0.cap_res_X.n17 two_stage_opamp_dummy_magic_16_0.cap_res_X.t40 0.1368
R6415 two_stage_opamp_dummy_magic_16_0.cap_res_X.n16 two_stage_opamp_dummy_magic_16_0.cap_res_X.t12 0.1368
R6416 two_stage_opamp_dummy_magic_16_0.cap_res_X.n16 two_stage_opamp_dummy_magic_16_0.cap_res_X.t82 0.1368
R6417 two_stage_opamp_dummy_magic_16_0.cap_res_X.n15 two_stage_opamp_dummy_magic_16_0.cap_res_X.t51 0.1368
R6418 two_stage_opamp_dummy_magic_16_0.cap_res_X.n15 two_stage_opamp_dummy_magic_16_0.cap_res_X.t123 0.1368
R6419 two_stage_opamp_dummy_magic_16_0.cap_res_X.n14 two_stage_opamp_dummy_magic_16_0.cap_res_X.t90 0.1368
R6420 two_stage_opamp_dummy_magic_16_0.cap_res_X.n14 two_stage_opamp_dummy_magic_16_0.cap_res_X.t22 0.1368
R6421 two_stage_opamp_dummy_magic_16_0.cap_res_X.n13 two_stage_opamp_dummy_magic_16_0.cap_res_X.t54 0.1368
R6422 two_stage_opamp_dummy_magic_16_0.cap_res_X.n13 two_stage_opamp_dummy_magic_16_0.cap_res_X.t127 0.1368
R6423 two_stage_opamp_dummy_magic_16_0.cap_res_X.n12 two_stage_opamp_dummy_magic_16_0.cap_res_X.t94 0.1368
R6424 two_stage_opamp_dummy_magic_16_0.cap_res_X.n12 two_stage_opamp_dummy_magic_16_0.cap_res_X.t28 0.1368
R6425 two_stage_opamp_dummy_magic_16_0.cap_res_X.n11 two_stage_opamp_dummy_magic_16_0.cap_res_X.t136 0.1368
R6426 two_stage_opamp_dummy_magic_16_0.cap_res_X.n11 two_stage_opamp_dummy_magic_16_0.cap_res_X.t68 0.1368
R6427 two_stage_opamp_dummy_magic_16_0.cap_res_X.n10 two_stage_opamp_dummy_magic_16_0.cap_res_X.t35 0.1368
R6428 two_stage_opamp_dummy_magic_16_0.cap_res_X.n9 two_stage_opamp_dummy_magic_16_0.cap_res_X.t38 0.1368
R6429 two_stage_opamp_dummy_magic_16_0.cap_res_X.n29 two_stage_opamp_dummy_magic_16_0.cap_res_X.n28 0.1133
R6430 two_stage_opamp_dummy_magic_16_0.cap_res_X.n30 two_stage_opamp_dummy_magic_16_0.cap_res_X.n29 0.1133
R6431 two_stage_opamp_dummy_magic_16_0.cap_res_X.n31 two_stage_opamp_dummy_magic_16_0.cap_res_X.n30 0.1133
R6432 two_stage_opamp_dummy_magic_16_0.cap_res_X.n32 two_stage_opamp_dummy_magic_16_0.cap_res_X.n31 0.1133
R6433 two_stage_opamp_dummy_magic_16_0.cap_res_X.n33 two_stage_opamp_dummy_magic_16_0.cap_res_X.n32 0.1133
R6434 two_stage_opamp_dummy_magic_16_0.cap_res_X.n1 two_stage_opamp_dummy_magic_16_0.cap_res_X.n0 0.1133
R6435 two_stage_opamp_dummy_magic_16_0.cap_res_X.n2 two_stage_opamp_dummy_magic_16_0.cap_res_X.n1 0.1133
R6436 two_stage_opamp_dummy_magic_16_0.cap_res_X.n3 two_stage_opamp_dummy_magic_16_0.cap_res_X.n2 0.1133
R6437 two_stage_opamp_dummy_magic_16_0.cap_res_X.n4 two_stage_opamp_dummy_magic_16_0.cap_res_X.n3 0.1133
R6438 two_stage_opamp_dummy_magic_16_0.cap_res_X.n5 two_stage_opamp_dummy_magic_16_0.cap_res_X.n4 0.1133
R6439 two_stage_opamp_dummy_magic_16_0.cap_res_X.n6 two_stage_opamp_dummy_magic_16_0.cap_res_X.n5 0.1133
R6440 two_stage_opamp_dummy_magic_16_0.cap_res_X.n7 two_stage_opamp_dummy_magic_16_0.cap_res_X.n6 0.1133
R6441 two_stage_opamp_dummy_magic_16_0.cap_res_X.n8 two_stage_opamp_dummy_magic_16_0.cap_res_X.n7 0.1133
R6442 two_stage_opamp_dummy_magic_16_0.cap_res_X.n10 two_stage_opamp_dummy_magic_16_0.cap_res_X.n8 0.1133
R6443 two_stage_opamp_dummy_magic_16_0.cap_res_X.n26 two_stage_opamp_dummy_magic_16_0.cap_res_X.n25 0.1133
R6444 two_stage_opamp_dummy_magic_16_0.cap_res_X.n27 two_stage_opamp_dummy_magic_16_0.cap_res_X.n26 0.1133
R6445 two_stage_opamp_dummy_magic_16_0.cap_res_X.n34 two_stage_opamp_dummy_magic_16_0.cap_res_X.n27 0.1133
R6446 two_stage_opamp_dummy_magic_16_0.cap_res_X.n34 two_stage_opamp_dummy_magic_16_0.cap_res_X.n33 0.1133
R6447 two_stage_opamp_dummy_magic_16_0.cap_res_X.n28 two_stage_opamp_dummy_magic_16_0.cap_res_X.t27 0.00152174
R6448 two_stage_opamp_dummy_magic_16_0.cap_res_X.n29 two_stage_opamp_dummy_magic_16_0.cap_res_X.t49 0.00152174
R6449 two_stage_opamp_dummy_magic_16_0.cap_res_X.n30 two_stage_opamp_dummy_magic_16_0.cap_res_X.t11 0.00152174
R6450 two_stage_opamp_dummy_magic_16_0.cap_res_X.n31 two_stage_opamp_dummy_magic_16_0.cap_res_X.t112 0.00152174
R6451 two_stage_opamp_dummy_magic_16_0.cap_res_X.n32 two_stage_opamp_dummy_magic_16_0.cap_res_X.t76 0.00152174
R6452 two_stage_opamp_dummy_magic_16_0.cap_res_X.n33 two_stage_opamp_dummy_magic_16_0.cap_res_X.t93 0.00152174
R6453 two_stage_opamp_dummy_magic_16_0.cap_res_X.n0 two_stage_opamp_dummy_magic_16_0.cap_res_X.t9 0.00152174
R6454 two_stage_opamp_dummy_magic_16_0.cap_res_X.n1 two_stage_opamp_dummy_magic_16_0.cap_res_X.t97 0.00152174
R6455 two_stage_opamp_dummy_magic_16_0.cap_res_X.n2 two_stage_opamp_dummy_magic_16_0.cap_res_X.t64 0.00152174
R6456 two_stage_opamp_dummy_magic_16_0.cap_res_X.n3 two_stage_opamp_dummy_magic_16_0.cap_res_X.t30 0.00152174
R6457 two_stage_opamp_dummy_magic_16_0.cap_res_X.n4 two_stage_opamp_dummy_magic_16_0.cap_res_X.t132 0.00152174
R6458 two_stage_opamp_dummy_magic_16_0.cap_res_X.n5 two_stage_opamp_dummy_magic_16_0.cap_res_X.t85 0.00152174
R6459 two_stage_opamp_dummy_magic_16_0.cap_res_X.n6 two_stage_opamp_dummy_magic_16_0.cap_res_X.t47 0.00152174
R6460 two_stage_opamp_dummy_magic_16_0.cap_res_X.n7 two_stage_opamp_dummy_magic_16_0.cap_res_X.t15 0.00152174
R6461 two_stage_opamp_dummy_magic_16_0.cap_res_X.n8 two_stage_opamp_dummy_magic_16_0.cap_res_X.t101 0.00152174
R6462 two_stage_opamp_dummy_magic_16_0.cap_res_X.n9 two_stage_opamp_dummy_magic_16_0.cap_res_X.t124 0.00152174
R6463 two_stage_opamp_dummy_magic_16_0.cap_res_X.n10 two_stage_opamp_dummy_magic_16_0.cap_res_X.t67 0.00152174
R6464 two_stage_opamp_dummy_magic_16_0.cap_res_X.n11 two_stage_opamp_dummy_magic_16_0.cap_res_X.t98 0.00152174
R6465 two_stage_opamp_dummy_magic_16_0.cap_res_X.n12 two_stage_opamp_dummy_magic_16_0.cap_res_X.t59 0.00152174
R6466 two_stage_opamp_dummy_magic_16_0.cap_res_X.n13 two_stage_opamp_dummy_magic_16_0.cap_res_X.t23 0.00152174
R6467 two_stage_opamp_dummy_magic_16_0.cap_res_X.n14 two_stage_opamp_dummy_magic_16_0.cap_res_X.t55 0.00152174
R6468 two_stage_opamp_dummy_magic_16_0.cap_res_X.n15 two_stage_opamp_dummy_magic_16_0.cap_res_X.t18 0.00152174
R6469 two_stage_opamp_dummy_magic_16_0.cap_res_X.n16 two_stage_opamp_dummy_magic_16_0.cap_res_X.t117 0.00152174
R6470 two_stage_opamp_dummy_magic_16_0.cap_res_X.n17 two_stage_opamp_dummy_magic_16_0.cap_res_X.t79 0.00152174
R6471 two_stage_opamp_dummy_magic_16_0.cap_res_X.n18 two_stage_opamp_dummy_magic_16_0.cap_res_X.t109 0.00152174
R6472 two_stage_opamp_dummy_magic_16_0.cap_res_X.n19 two_stage_opamp_dummy_magic_16_0.cap_res_X.t73 0.00152174
R6473 two_stage_opamp_dummy_magic_16_0.cap_res_X.n20 two_stage_opamp_dummy_magic_16_0.cap_res_X.t36 0.00152174
R6474 two_stage_opamp_dummy_magic_16_0.cap_res_X.n21 two_stage_opamp_dummy_magic_16_0.cap_res_X.t69 0.00152174
R6475 two_stage_opamp_dummy_magic_16_0.cap_res_X.n22 two_stage_opamp_dummy_magic_16_0.cap_res_X.t29 0.00152174
R6476 two_stage_opamp_dummy_magic_16_0.cap_res_X.n23 two_stage_opamp_dummy_magic_16_0.cap_res_X.t10 0.00152174
R6477 two_stage_opamp_dummy_magic_16_0.cap_res_X.n24 two_stage_opamp_dummy_magic_16_0.cap_res_X.t45 0.00152174
R6478 two_stage_opamp_dummy_magic_16_0.cap_res_X.n25 two_stage_opamp_dummy_magic_16_0.cap_res_X.t2 0.00152174
R6479 two_stage_opamp_dummy_magic_16_0.cap_res_X.n26 two_stage_opamp_dummy_magic_16_0.cap_res_X.t41 0.00152174
R6480 two_stage_opamp_dummy_magic_16_0.cap_res_X.n27 two_stage_opamp_dummy_magic_16_0.cap_res_X.t21 0.00152174
R6481 two_stage_opamp_dummy_magic_16_0.cap_res_X.t57 two_stage_opamp_dummy_magic_16_0.cap_res_X.n34 0.00152174
R6482 VOUT+.n8 VOUT+.n6 149.19
R6483 VOUT+.n14 VOUT+.n13 149.19
R6484 VOUT+.n12 VOUT+.n11 148.626
R6485 VOUT+.n10 VOUT+.n9 148.626
R6486 VOUT+.n8 VOUT+.n7 148.626
R6487 VOUT+.n16 VOUT+.n15 144.126
R6488 VOUT+.n5 VOUT+.t5 112.184
R6489 VOUT+.n2 VOUT+.n0 98.9303
R6490 VOUT+.n4 VOUT+.n3 97.8053
R6491 VOUT+.n2 VOUT+.n1 97.8053
R6492 VOUT+.n91 VOUT+.n16 15.5682
R6493 VOUT+.n91 VOUT+.n90 11.5649
R6494 VOUT+ VOUT+.n91 9.2505
R6495 VOUT+.n15 VOUT+.t4 6.56717
R6496 VOUT+.n15 VOUT+.t13 6.56717
R6497 VOUT+.n13 VOUT+.t7 6.56717
R6498 VOUT+.n13 VOUT+.t12 6.56717
R6499 VOUT+.n11 VOUT+.t3 6.56717
R6500 VOUT+.n11 VOUT+.t17 6.56717
R6501 VOUT+.n9 VOUT+.t2 6.56717
R6502 VOUT+.n9 VOUT+.t1 6.56717
R6503 VOUT+.n7 VOUT+.t0 6.56717
R6504 VOUT+.n7 VOUT+.t8 6.56717
R6505 VOUT+.n6 VOUT+.t11 6.56717
R6506 VOUT+.n6 VOUT+.t14 6.56717
R6507 VOUT+.n45 VOUT+.t56 4.8295
R6508 VOUT+.n47 VOUT+.t105 4.8295
R6509 VOUT+.n48 VOUT+.t29 4.8295
R6510 VOUT+.n50 VOUT+.t60 4.8295
R6511 VOUT+.n52 VOUT+.t115 4.8295
R6512 VOUT+.n63 VOUT+.t20 4.8295
R6513 VOUT+.n66 VOUT+.t31 4.8295
R6514 VOUT+.n65 VOUT+.t121 4.8295
R6515 VOUT+.n68 VOUT+.t67 4.8295
R6516 VOUT+.n67 VOUT+.t152 4.8295
R6517 VOUT+.n69 VOUT+.t131 4.8295
R6518 VOUT+.n70 VOUT+.t118 4.8295
R6519 VOUT+.n72 VOUT+.t89 4.8295
R6520 VOUT+.n73 VOUT+.t76 4.8295
R6521 VOUT+.n75 VOUT+.t127 4.8295
R6522 VOUT+.n76 VOUT+.t110 4.8295
R6523 VOUT+.n78 VOUT+.t84 4.8295
R6524 VOUT+.n79 VOUT+.t68 4.8295
R6525 VOUT+.n81 VOUT+.t42 4.8295
R6526 VOUT+.n82 VOUT+.t30 4.8295
R6527 VOUT+.n84 VOUT+.t81 4.8295
R6528 VOUT+.n85 VOUT+.t64 4.8295
R6529 VOUT+.n17 VOUT+.t150 4.8295
R6530 VOUT+.n28 VOUT+.t75 4.8295
R6531 VOUT+.n30 VOUT+.t54 4.8295
R6532 VOUT+.n31 VOUT+.t34 4.8295
R6533 VOUT+.n33 VOUT+.t95 4.8295
R6534 VOUT+.n34 VOUT+.t79 4.8295
R6535 VOUT+.n36 VOUT+.t134 4.8295
R6536 VOUT+.n37 VOUT+.t122 4.8295
R6537 VOUT+.n39 VOUT+.t102 4.8295
R6538 VOUT+.n40 VOUT+.t82 4.8295
R6539 VOUT+.n42 VOUT+.t137 4.8295
R6540 VOUT+.n43 VOUT+.t126 4.8295
R6541 VOUT+.n87 VOUT+.t28 4.8295
R6542 VOUT+.n56 VOUT+.t57 4.8154
R6543 VOUT+.n55 VOUT+.t33 4.8154
R6544 VOUT+.n54 VOUT+.t77 4.8154
R6545 VOUT+.n62 VOUT+.t116 4.806
R6546 VOUT+.n61 VOUT+.t147 4.806
R6547 VOUT+.n60 VOUT+.t43 4.806
R6548 VOUT+.n59 VOUT+.t83 4.806
R6549 VOUT+.n58 VOUT+.t63 4.806
R6550 VOUT+.n57 VOUT+.t26 4.806
R6551 VOUT+.n57 VOUT+.t103 4.806
R6552 VOUT+.n56 VOUT+.t135 4.806
R6553 VOUT+.n55 VOUT+.t120 4.806
R6554 VOUT+.n54 VOUT+.t155 4.806
R6555 VOUT+.n27 VOUT+.t91 4.806
R6556 VOUT+.n26 VOUT+.t38 4.806
R6557 VOUT+.n25 VOUT+.t130 4.806
R6558 VOUT+.n25 VOUT+.t90 4.806
R6559 VOUT+.n24 VOUT+.t80 4.806
R6560 VOUT+.n24 VOUT+.t128 4.806
R6561 VOUT+.n23 VOUT+.t124 4.806
R6562 VOUT+.n23 VOUT+.t32 4.806
R6563 VOUT+.n22 VOUT+.t70 4.806
R6564 VOUT+.n22 VOUT+.t73 4.806
R6565 VOUT+.n21 VOUT+.t23 4.806
R6566 VOUT+.n21 VOUT+.t108 4.806
R6567 VOUT+.n20 VOUT+.t62 4.806
R6568 VOUT+.n20 VOUT+.t19 4.806
R6569 VOUT+.n19 VOUT+.t151 4.806
R6570 VOUT+.n19 VOUT+.t49 4.806
R6571 VOUT+.n46 VOUT+.t132 4.5005
R6572 VOUT+.n45 VOUT+.t96 4.5005
R6573 VOUT+.n47 VOUT+.t69 4.5005
R6574 VOUT+.n48 VOUT+.t139 4.5005
R6575 VOUT+.n49 VOUT+.t109 4.5005
R6576 VOUT+.n50 VOUT+.t37 4.5005
R6577 VOUT+.n51 VOUT+.t144 4.5005
R6578 VOUT+.n52 VOUT+.t21 4.5005
R6579 VOUT+.n53 VOUT+.t125 4.5005
R6580 VOUT+.n54 VOUT+.t119 4.5005
R6581 VOUT+.n55 VOUT+.t78 4.5005
R6582 VOUT+.n56 VOUT+.t97 4.5005
R6583 VOUT+.n57 VOUT+.t61 4.5005
R6584 VOUT+.n58 VOUT+.t27 4.5005
R6585 VOUT+.n59 VOUT+.t41 4.5005
R6586 VOUT+.n60 VOUT+.t145 4.5005
R6587 VOUT+.n61 VOUT+.t113 4.5005
R6588 VOUT+.n62 VOUT+.t72 4.5005
R6589 VOUT+.n64 VOUT+.t92 4.5005
R6590 VOUT+.n63 VOUT+.t55 4.5005
R6591 VOUT+.n66 VOUT+.t50 4.5005
R6592 VOUT+.n65 VOUT+.t156 4.5005
R6593 VOUT+.n68 VOUT+.t86 4.5005
R6594 VOUT+.n67 VOUT+.t47 4.5005
R6595 VOUT+.n69 VOUT+.t94 4.5005
R6596 VOUT+.n71 VOUT+.t39 4.5005
R6597 VOUT+.n70 VOUT+.t146 4.5005
R6598 VOUT+.n72 VOUT+.t53 4.5005
R6599 VOUT+.n74 VOUT+.t142 4.5005
R6600 VOUT+.n73 VOUT+.t112 4.5005
R6601 VOUT+.n75 VOUT+.t88 4.5005
R6602 VOUT+.n77 VOUT+.t35 4.5005
R6603 VOUT+.n76 VOUT+.t140 4.5005
R6604 VOUT+.n78 VOUT+.t46 4.5005
R6605 VOUT+.n80 VOUT+.t136 4.5005
R6606 VOUT+.n79 VOUT+.t104 4.5005
R6607 VOUT+.n81 VOUT+.t149 4.5005
R6608 VOUT+.n83 VOUT+.t99 4.5005
R6609 VOUT+.n82 VOUT+.t65 4.5005
R6610 VOUT+.n84 VOUT+.t40 4.5005
R6611 VOUT+.n86 VOUT+.t133 4.5005
R6612 VOUT+.n85 VOUT+.t98 4.5005
R6613 VOUT+.n18 VOUT+.t45 4.5005
R6614 VOUT+.n17 VOUT+.t101 4.5005
R6615 VOUT+.n19 VOUT+.t85 4.5005
R6616 VOUT+.n20 VOUT+.t48 4.5005
R6617 VOUT+.n21 VOUT+.t138 4.5005
R6618 VOUT+.n22 VOUT+.t107 4.5005
R6619 VOUT+.n23 VOUT+.t71 4.5005
R6620 VOUT+.n24 VOUT+.t25 4.5005
R6621 VOUT+.n25 VOUT+.t129 4.5005
R6622 VOUT+.n26 VOUT+.t87 4.5005
R6623 VOUT+.n27 VOUT+.t52 4.5005
R6624 VOUT+.n29 VOUT+.t141 4.5005
R6625 VOUT+.n28 VOUT+.t111 4.5005
R6626 VOUT+.n30 VOUT+.t24 4.5005
R6627 VOUT+.n32 VOUT+.t114 4.5005
R6628 VOUT+.n31 VOUT+.t74 4.5005
R6629 VOUT+.n33 VOUT+.t59 4.5005
R6630 VOUT+.n35 VOUT+.t148 4.5005
R6631 VOUT+.n34 VOUT+.t117 4.5005
R6632 VOUT+.n36 VOUT+.t100 4.5005
R6633 VOUT+.n38 VOUT+.t44 4.5005
R6634 VOUT+.n37 VOUT+.t153 4.5005
R6635 VOUT+.n39 VOUT+.t66 4.5005
R6636 VOUT+.n41 VOUT+.t154 4.5005
R6637 VOUT+.n40 VOUT+.t123 4.5005
R6638 VOUT+.n42 VOUT+.t106 4.5005
R6639 VOUT+.n44 VOUT+.t51 4.5005
R6640 VOUT+.n43 VOUT+.t22 4.5005
R6641 VOUT+.n90 VOUT+.t36 4.5005
R6642 VOUT+.n89 VOUT+.t143 4.5005
R6643 VOUT+.n88 VOUT+.t93 4.5005
R6644 VOUT+.n87 VOUT+.t58 4.5005
R6645 VOUT+.n16 VOUT+.n14 4.5005
R6646 VOUT+.n3 VOUT+.t16 3.42907
R6647 VOUT+.n3 VOUT+.t9 3.42907
R6648 VOUT+.n1 VOUT+.t18 3.42907
R6649 VOUT+.n1 VOUT+.t6 3.42907
R6650 VOUT+.n0 VOUT+.t10 3.42907
R6651 VOUT+.n0 VOUT+.t15 3.42907
R6652 VOUT+ VOUT+.n5 1.46144
R6653 VOUT+.n5 VOUT+.n4 1.30519
R6654 VOUT+.n4 VOUT+.n2 1.1255
R6655 VOUT+.n10 VOUT+.n8 0.563
R6656 VOUT+.n12 VOUT+.n10 0.563
R6657 VOUT+.n14 VOUT+.n12 0.563
R6658 VOUT+.n46 VOUT+.n45 0.3295
R6659 VOUT+.n49 VOUT+.n48 0.3295
R6660 VOUT+.n51 VOUT+.n50 0.3295
R6661 VOUT+.n53 VOUT+.n52 0.3295
R6662 VOUT+.n55 VOUT+.n54 0.3295
R6663 VOUT+.n56 VOUT+.n55 0.3295
R6664 VOUT+.n57 VOUT+.n56 0.3295
R6665 VOUT+.n58 VOUT+.n57 0.3295
R6666 VOUT+.n59 VOUT+.n58 0.3295
R6667 VOUT+.n60 VOUT+.n59 0.3295
R6668 VOUT+.n61 VOUT+.n60 0.3295
R6669 VOUT+.n62 VOUT+.n61 0.3295
R6670 VOUT+.n64 VOUT+.n62 0.3295
R6671 VOUT+.n64 VOUT+.n63 0.3295
R6672 VOUT+.n66 VOUT+.n65 0.3295
R6673 VOUT+.n68 VOUT+.n67 0.3295
R6674 VOUT+.n71 VOUT+.n69 0.3295
R6675 VOUT+.n71 VOUT+.n70 0.3295
R6676 VOUT+.n74 VOUT+.n72 0.3295
R6677 VOUT+.n74 VOUT+.n73 0.3295
R6678 VOUT+.n77 VOUT+.n75 0.3295
R6679 VOUT+.n77 VOUT+.n76 0.3295
R6680 VOUT+.n80 VOUT+.n78 0.3295
R6681 VOUT+.n80 VOUT+.n79 0.3295
R6682 VOUT+.n83 VOUT+.n81 0.3295
R6683 VOUT+.n83 VOUT+.n82 0.3295
R6684 VOUT+.n86 VOUT+.n84 0.3295
R6685 VOUT+.n86 VOUT+.n85 0.3295
R6686 VOUT+.n18 VOUT+.n17 0.3295
R6687 VOUT+.n20 VOUT+.n19 0.3295
R6688 VOUT+.n21 VOUT+.n20 0.3295
R6689 VOUT+.n22 VOUT+.n21 0.3295
R6690 VOUT+.n23 VOUT+.n22 0.3295
R6691 VOUT+.n24 VOUT+.n23 0.3295
R6692 VOUT+.n25 VOUT+.n24 0.3295
R6693 VOUT+.n26 VOUT+.n25 0.3295
R6694 VOUT+.n27 VOUT+.n26 0.3295
R6695 VOUT+.n29 VOUT+.n27 0.3295
R6696 VOUT+.n29 VOUT+.n28 0.3295
R6697 VOUT+.n32 VOUT+.n30 0.3295
R6698 VOUT+.n32 VOUT+.n31 0.3295
R6699 VOUT+.n35 VOUT+.n33 0.3295
R6700 VOUT+.n35 VOUT+.n34 0.3295
R6701 VOUT+.n38 VOUT+.n36 0.3295
R6702 VOUT+.n38 VOUT+.n37 0.3295
R6703 VOUT+.n41 VOUT+.n39 0.3295
R6704 VOUT+.n41 VOUT+.n40 0.3295
R6705 VOUT+.n44 VOUT+.n42 0.3295
R6706 VOUT+.n44 VOUT+.n43 0.3295
R6707 VOUT+.n90 VOUT+.n89 0.3295
R6708 VOUT+.n89 VOUT+.n88 0.3295
R6709 VOUT+.n88 VOUT+.n87 0.3295
R6710 VOUT+.n61 VOUT+.n47 0.306
R6711 VOUT+.n60 VOUT+.n49 0.306
R6712 VOUT+.n59 VOUT+.n51 0.306
R6713 VOUT+.n58 VOUT+.n53 0.306
R6714 VOUT+.n64 VOUT+.n46 0.2825
R6715 VOUT+.n66 VOUT+.n64 0.2825
R6716 VOUT+.n68 VOUT+.n66 0.2825
R6717 VOUT+.n71 VOUT+.n68 0.2825
R6718 VOUT+.n74 VOUT+.n71 0.2825
R6719 VOUT+.n77 VOUT+.n74 0.2825
R6720 VOUT+.n80 VOUT+.n77 0.2825
R6721 VOUT+.n83 VOUT+.n80 0.2825
R6722 VOUT+.n86 VOUT+.n83 0.2825
R6723 VOUT+.n29 VOUT+.n18 0.2825
R6724 VOUT+.n32 VOUT+.n29 0.2825
R6725 VOUT+.n35 VOUT+.n32 0.2825
R6726 VOUT+.n38 VOUT+.n35 0.2825
R6727 VOUT+.n41 VOUT+.n38 0.2825
R6728 VOUT+.n44 VOUT+.n41 0.2825
R6729 VOUT+.n88 VOUT+.n44 0.2825
R6730 VOUT+.n88 VOUT+.n86 0.2825
R6731 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t128 50.3211
R6732 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t102 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t137 0.1603
R6733 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t61 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t101 0.1603
R6734 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t1 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t36 0.1603
R6735 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t110 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t5 0.1603
R6736 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t11 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t39 0.1603
R6737 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t63 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t26 0.1603
R6738 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t45 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t81 0.1603
R6739 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t104 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t68 0.1603
R6740 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t17 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t47 0.1603
R6741 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t69 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t30 0.1603
R6742 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t53 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t89 0.1603
R6743 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t111 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t73 0.1603
R6744 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t92 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t127 0.1603
R6745 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t8 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t115 0.1603
R6746 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t93 0.1603
R6747 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t117 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t76 0.1603
R6748 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t99 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t129 0.1603
R6749 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t14 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t121 0.1603
R6750 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t135 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t31 0.1603
R6751 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t51 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t20 0.1603
R6752 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t34 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t75 0.1603
R6753 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t91 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t55 0.1603
R6754 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t4 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t35 0.1603
R6755 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t57 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t23 0.1603
R6756 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t40 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t78 0.1603
R6757 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t98 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t62 0.1603
R6758 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t83 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t123 0.1603
R6759 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t133 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t103 0.1603
R6760 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t46 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t82 0.1603
R6761 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t72 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t6 0.1603
R6762 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t109 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t95 0.1603
R6763 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t19 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t134 0.1603
R6764 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t50 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t87 0.1603
R6765 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t86 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t33 0.1603
R6766 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t132 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t77 0.1603
R6767 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t28 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t27 0.1603
R6768 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t70 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t119 0.1603
R6769 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t105 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t66 0.1603
R6770 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t56 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t7 0.1603
R6771 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t88 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t52 0.1603
R6772 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t88 0.1603
R6773 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t38 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t80 0.1603
R6774 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t79 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t124 0.1603
R6775 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t60 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t100 0.1603
R6776 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t96 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t131 0.1603
R6777 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t136 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t42 0.1603
R6778 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t32 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t136 0.1603
R6779 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t130 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t32 0.1603
R6780 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t120 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t97 0.1603
R6781 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t13 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t120 0.1603
R6782 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t116 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t13 0.1603
R6783 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t48 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t12 0.1603
R6784 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t18 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t48 0.1603
R6785 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t128 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t18 0.1603
R6786 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t25 0.159278
R6787 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t108 0.159278
R6788 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t138 0.159278
R6789 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t49 0.159278
R6790 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t84 0.159278
R6791 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t125 0.159278
R6792 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t29 0.159278
R6793 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t67 0.159278
R6794 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n15 0.159278
R6795 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t43 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n16 0.159278
R6796 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t9 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n17 0.159278
R6797 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t113 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n18 0.159278
R6798 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t3 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n19 0.159278
R6799 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t106 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n20 0.159278
R6800 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t64 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n21 0.159278
R6801 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t24 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n22 0.159278
R6802 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t58 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n23 0.159278
R6803 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t21 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n24 0.159278
R6804 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t122 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n25 0.159278
R6805 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t15 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n26 0.159278
R6806 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t118 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n27 0.159278
R6807 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t71 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n28 0.159278
R6808 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t107 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n29 0.159278
R6809 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t65 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n30 0.159278
R6810 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t41 0.159278
R6811 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t10 0.159278
R6812 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t2 0.159278
R6813 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t37 0.159278
R6814 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t22 0.159278
R6815 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t54 0.159278
R6816 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t94 0.159278
R6817 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t74 0.159278
R6818 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t114 0.159278
R6819 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t25 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t61 0.137822
R6820 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t102 0.1368
R6821 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t1 0.1368
R6822 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t126 0.1368
R6823 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t110 0.1368
R6824 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t90 0.1368
R6825 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t11 0.1368
R6826 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t63 0.1368
R6827 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t45 0.1368
R6828 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t104 0.1368
R6829 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t17 0.1368
R6830 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t69 0.1368
R6831 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t53 0.1368
R6832 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t111 0.1368
R6833 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t92 0.1368
R6834 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t8 0.1368
R6835 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t59 0.1368
R6836 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t117 0.1368
R6837 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t99 0.1368
R6838 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t14 0.1368
R6839 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t135 0.1368
R6840 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t51 0.1368
R6841 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t34 0.1368
R6842 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t91 0.1368
R6843 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t4 0.1368
R6844 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t57 0.1368
R6845 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t40 0.1368
R6846 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t98 0.1368
R6847 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t83 0.1368
R6848 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t133 0.1368
R6849 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t46 0.1368
R6850 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t56 0.1368
R6851 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n6 0.1133
R6852 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n7 0.1133
R6853 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n8 0.1133
R6854 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n9 0.1133
R6855 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n10 0.1133
R6856 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n11 0.1133
R6857 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n12 0.1133
R6858 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n13 0.1133
R6859 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n14 0.1133
R6860 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n31 0.1133
R6861 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n32 0.1133
R6862 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n0 0.1133
R6863 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n1 0.1133
R6864 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n2 0.1133
R6865 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n3 0.1133
R6866 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n4 0.1133
R6867 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n5 0.1133
R6868 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n33 0.1133
R6869 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t72 0.00152174
R6870 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t109 0.00152174
R6871 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t19 0.00152174
R6872 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t50 0.00152174
R6873 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t86 0.00152174
R6874 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t132 0.00152174
R6875 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t28 0.00152174
R6876 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t70 0.00152174
R6877 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t105 0.00152174
R6878 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t112 0.00152174
R6879 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t16 0.00152174
R6880 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t43 0.00152174
R6881 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t9 0.00152174
R6882 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t113 0.00152174
R6883 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t3 0.00152174
R6884 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t106 0.00152174
R6885 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t64 0.00152174
R6886 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t24 0.00152174
R6887 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t58 0.00152174
R6888 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t21 0.00152174
R6889 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t122 0.00152174
R6890 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t15 0.00152174
R6891 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t118 0.00152174
R6892 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t71 0.00152174
R6893 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t107 0.00152174
R6894 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t65 0.00152174
R6895 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t85 0.00152174
R6896 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t44 0.00152174
R6897 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t38 0.00152174
R6898 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t79 0.00152174
R6899 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t60 0.00152174
R6900 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t96 0.00152174
R6901 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t130 0.00152174
R6902 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t116 0.00152174
R6903 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t12 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n34 0.00152174
R6904 two_stage_opamp_dummy_magic_16_0.X.n47 two_stage_opamp_dummy_magic_16_0.X.t51 1172.87
R6905 two_stage_opamp_dummy_magic_16_0.X.n43 two_stage_opamp_dummy_magic_16_0.X.t27 1172.87
R6906 two_stage_opamp_dummy_magic_16_0.X.n50 two_stage_opamp_dummy_magic_16_0.X.t48 996.134
R6907 two_stage_opamp_dummy_magic_16_0.X.n49 two_stage_opamp_dummy_magic_16_0.X.t35 996.134
R6908 two_stage_opamp_dummy_magic_16_0.X.n48 two_stage_opamp_dummy_magic_16_0.X.t42 996.134
R6909 two_stage_opamp_dummy_magic_16_0.X.n47 two_stage_opamp_dummy_magic_16_0.X.t34 996.134
R6910 two_stage_opamp_dummy_magic_16_0.X.n43 two_stage_opamp_dummy_magic_16_0.X.t43 996.134
R6911 two_stage_opamp_dummy_magic_16_0.X.n44 two_stage_opamp_dummy_magic_16_0.X.t29 996.134
R6912 two_stage_opamp_dummy_magic_16_0.X.n45 two_stage_opamp_dummy_magic_16_0.X.t45 996.134
R6913 two_stage_opamp_dummy_magic_16_0.X.n46 two_stage_opamp_dummy_magic_16_0.X.t31 996.134
R6914 two_stage_opamp_dummy_magic_16_0.X.n25 two_stage_opamp_dummy_magic_16_0.X.t26 690.867
R6915 two_stage_opamp_dummy_magic_16_0.X.n20 two_stage_opamp_dummy_magic_16_0.X.t32 690.867
R6916 two_stage_opamp_dummy_magic_16_0.X.n16 two_stage_opamp_dummy_magic_16_0.X.t39 530.201
R6917 two_stage_opamp_dummy_magic_16_0.X.n11 two_stage_opamp_dummy_magic_16_0.X.t44 530.201
R6918 two_stage_opamp_dummy_magic_16_0.X.n25 two_stage_opamp_dummy_magic_16_0.X.t40 514.134
R6919 two_stage_opamp_dummy_magic_16_0.X.n26 two_stage_opamp_dummy_magic_16_0.X.t46 514.134
R6920 two_stage_opamp_dummy_magic_16_0.X.n27 two_stage_opamp_dummy_magic_16_0.X.t41 514.134
R6921 two_stage_opamp_dummy_magic_16_0.X.n24 two_stage_opamp_dummy_magic_16_0.X.t25 514.134
R6922 two_stage_opamp_dummy_magic_16_0.X.n23 two_stage_opamp_dummy_magic_16_0.X.t38 514.134
R6923 two_stage_opamp_dummy_magic_16_0.X.n22 two_stage_opamp_dummy_magic_16_0.X.t52 514.134
R6924 two_stage_opamp_dummy_magic_16_0.X.n21 two_stage_opamp_dummy_magic_16_0.X.t36 514.134
R6925 two_stage_opamp_dummy_magic_16_0.X.n20 two_stage_opamp_dummy_magic_16_0.X.t49 514.134
R6926 two_stage_opamp_dummy_magic_16_0.X.n18 two_stage_opamp_dummy_magic_16_0.X.t54 353.467
R6927 two_stage_opamp_dummy_magic_16_0.X.n17 two_stage_opamp_dummy_magic_16_0.X.t28 353.467
R6928 two_stage_opamp_dummy_magic_16_0.X.n16 two_stage_opamp_dummy_magic_16_0.X.t53 353.467
R6929 two_stage_opamp_dummy_magic_16_0.X.n11 two_stage_opamp_dummy_magic_16_0.X.t30 353.467
R6930 two_stage_opamp_dummy_magic_16_0.X.n12 two_stage_opamp_dummy_magic_16_0.X.t47 353.467
R6931 two_stage_opamp_dummy_magic_16_0.X.n13 two_stage_opamp_dummy_magic_16_0.X.t33 353.467
R6932 two_stage_opamp_dummy_magic_16_0.X.n14 two_stage_opamp_dummy_magic_16_0.X.t50 353.467
R6933 two_stage_opamp_dummy_magic_16_0.X.n15 two_stage_opamp_dummy_magic_16_0.X.t37 353.467
R6934 two_stage_opamp_dummy_magic_16_0.X.n50 two_stage_opamp_dummy_magic_16_0.X.n49 176.733
R6935 two_stage_opamp_dummy_magic_16_0.X.n49 two_stage_opamp_dummy_magic_16_0.X.n48 176.733
R6936 two_stage_opamp_dummy_magic_16_0.X.n48 two_stage_opamp_dummy_magic_16_0.X.n47 176.733
R6937 two_stage_opamp_dummy_magic_16_0.X.n44 two_stage_opamp_dummy_magic_16_0.X.n43 176.733
R6938 two_stage_opamp_dummy_magic_16_0.X.n45 two_stage_opamp_dummy_magic_16_0.X.n44 176.733
R6939 two_stage_opamp_dummy_magic_16_0.X.n46 two_stage_opamp_dummy_magic_16_0.X.n45 176.733
R6940 two_stage_opamp_dummy_magic_16_0.X.n18 two_stage_opamp_dummy_magic_16_0.X.n17 176.733
R6941 two_stage_opamp_dummy_magic_16_0.X.n17 two_stage_opamp_dummy_magic_16_0.X.n16 176.733
R6942 two_stage_opamp_dummy_magic_16_0.X.n12 two_stage_opamp_dummy_magic_16_0.X.n11 176.733
R6943 two_stage_opamp_dummy_magic_16_0.X.n13 two_stage_opamp_dummy_magic_16_0.X.n12 176.733
R6944 two_stage_opamp_dummy_magic_16_0.X.n14 two_stage_opamp_dummy_magic_16_0.X.n13 176.733
R6945 two_stage_opamp_dummy_magic_16_0.X.n15 two_stage_opamp_dummy_magic_16_0.X.n14 176.733
R6946 two_stage_opamp_dummy_magic_16_0.X.n27 two_stage_opamp_dummy_magic_16_0.X.n26 176.733
R6947 two_stage_opamp_dummy_magic_16_0.X.n26 two_stage_opamp_dummy_magic_16_0.X.n25 176.733
R6948 two_stage_opamp_dummy_magic_16_0.X.n21 two_stage_opamp_dummy_magic_16_0.X.n20 176.733
R6949 two_stage_opamp_dummy_magic_16_0.X.n22 two_stage_opamp_dummy_magic_16_0.X.n21 176.733
R6950 two_stage_opamp_dummy_magic_16_0.X.n23 two_stage_opamp_dummy_magic_16_0.X.n22 176.733
R6951 two_stage_opamp_dummy_magic_16_0.X.n24 two_stage_opamp_dummy_magic_16_0.X.n23 176.733
R6952 two_stage_opamp_dummy_magic_16_0.X.n52 two_stage_opamp_dummy_magic_16_0.X.n51 166.258
R6953 two_stage_opamp_dummy_magic_16_0.X.n2 two_stage_opamp_dummy_magic_16_0.X.n0 163.626
R6954 two_stage_opamp_dummy_magic_16_0.X.n8 two_stage_opamp_dummy_magic_16_0.X.n7 163.001
R6955 two_stage_opamp_dummy_magic_16_0.X.n6 two_stage_opamp_dummy_magic_16_0.X.n5 163.001
R6956 two_stage_opamp_dummy_magic_16_0.X.n4 two_stage_opamp_dummy_magic_16_0.X.n3 163.001
R6957 two_stage_opamp_dummy_magic_16_0.X.n2 two_stage_opamp_dummy_magic_16_0.X.n1 163.001
R6958 two_stage_opamp_dummy_magic_16_0.X.n29 two_stage_opamp_dummy_magic_16_0.X.n19 161.541
R6959 two_stage_opamp_dummy_magic_16_0.X.n29 two_stage_opamp_dummy_magic_16_0.X.n28 161.541
R6960 two_stage_opamp_dummy_magic_16_0.X.n10 two_stage_opamp_dummy_magic_16_0.X.n9 158.501
R6961 two_stage_opamp_dummy_magic_16_0.X.n32 two_stage_opamp_dummy_magic_16_0.X.n30 117.906
R6962 two_stage_opamp_dummy_magic_16_0.X.n40 two_stage_opamp_dummy_magic_16_0.X.n39 117.326
R6963 two_stage_opamp_dummy_magic_16_0.X.n38 two_stage_opamp_dummy_magic_16_0.X.n37 117.326
R6964 two_stage_opamp_dummy_magic_16_0.X.n36 two_stage_opamp_dummy_magic_16_0.X.n35 117.326
R6965 two_stage_opamp_dummy_magic_16_0.X.n34 two_stage_opamp_dummy_magic_16_0.X.n33 117.326
R6966 two_stage_opamp_dummy_magic_16_0.X.n32 two_stage_opamp_dummy_magic_16_0.X.n31 117.326
R6967 two_stage_opamp_dummy_magic_16_0.X.n19 two_stage_opamp_dummy_magic_16_0.X.n18 54.6272
R6968 two_stage_opamp_dummy_magic_16_0.X.n19 two_stage_opamp_dummy_magic_16_0.X.n15 54.6272
R6969 two_stage_opamp_dummy_magic_16_0.X.n28 two_stage_opamp_dummy_magic_16_0.X.n27 54.6272
R6970 two_stage_opamp_dummy_magic_16_0.X.n28 two_stage_opamp_dummy_magic_16_0.X.n24 54.6272
R6971 two_stage_opamp_dummy_magic_16_0.X.n51 two_stage_opamp_dummy_magic_16_0.X.n50 53.3126
R6972 two_stage_opamp_dummy_magic_16_0.X.n51 two_stage_opamp_dummy_magic_16_0.X.n46 53.3126
R6973 two_stage_opamp_dummy_magic_16_0.X.t13 two_stage_opamp_dummy_magic_16_0.X.n52 50.3023
R6974 two_stage_opamp_dummy_magic_16_0.X.n42 two_stage_opamp_dummy_magic_16_0.X.n10 16.8755
R6975 two_stage_opamp_dummy_magic_16_0.X.n39 two_stage_opamp_dummy_magic_16_0.X.t20 16.0005
R6976 two_stage_opamp_dummy_magic_16_0.X.n39 two_stage_opamp_dummy_magic_16_0.X.t5 16.0005
R6977 two_stage_opamp_dummy_magic_16_0.X.n37 two_stage_opamp_dummy_magic_16_0.X.t9 16.0005
R6978 two_stage_opamp_dummy_magic_16_0.X.n37 two_stage_opamp_dummy_magic_16_0.X.t22 16.0005
R6979 two_stage_opamp_dummy_magic_16_0.X.n35 two_stage_opamp_dummy_magic_16_0.X.t21 16.0005
R6980 two_stage_opamp_dummy_magic_16_0.X.n35 two_stage_opamp_dummy_magic_16_0.X.t12 16.0005
R6981 two_stage_opamp_dummy_magic_16_0.X.n33 two_stage_opamp_dummy_magic_16_0.X.t2 16.0005
R6982 two_stage_opamp_dummy_magic_16_0.X.n33 two_stage_opamp_dummy_magic_16_0.X.t17 16.0005
R6983 two_stage_opamp_dummy_magic_16_0.X.n31 two_stage_opamp_dummy_magic_16_0.X.t11 16.0005
R6984 two_stage_opamp_dummy_magic_16_0.X.n31 two_stage_opamp_dummy_magic_16_0.X.t16 16.0005
R6985 two_stage_opamp_dummy_magic_16_0.X.n30 two_stage_opamp_dummy_magic_16_0.X.t23 16.0005
R6986 two_stage_opamp_dummy_magic_16_0.X.n30 two_stage_opamp_dummy_magic_16_0.X.t19 16.0005
R6987 two_stage_opamp_dummy_magic_16_0.X.n41 two_stage_opamp_dummy_magic_16_0.X.n29 12.4067
R6988 two_stage_opamp_dummy_magic_16_0.X.n9 two_stage_opamp_dummy_magic_16_0.X.t7 11.2576
R6989 two_stage_opamp_dummy_magic_16_0.X.n9 two_stage_opamp_dummy_magic_16_0.X.t3 11.2576
R6990 two_stage_opamp_dummy_magic_16_0.X.n7 two_stage_opamp_dummy_magic_16_0.X.t4 11.2576
R6991 two_stage_opamp_dummy_magic_16_0.X.n7 two_stage_opamp_dummy_magic_16_0.X.t0 11.2576
R6992 two_stage_opamp_dummy_magic_16_0.X.n5 two_stage_opamp_dummy_magic_16_0.X.t1 11.2576
R6993 two_stage_opamp_dummy_magic_16_0.X.n5 two_stage_opamp_dummy_magic_16_0.X.t8 11.2576
R6994 two_stage_opamp_dummy_magic_16_0.X.n3 two_stage_opamp_dummy_magic_16_0.X.t14 11.2576
R6995 two_stage_opamp_dummy_magic_16_0.X.n3 two_stage_opamp_dummy_magic_16_0.X.t18 11.2576
R6996 two_stage_opamp_dummy_magic_16_0.X.n1 two_stage_opamp_dummy_magic_16_0.X.t24 11.2576
R6997 two_stage_opamp_dummy_magic_16_0.X.n1 two_stage_opamp_dummy_magic_16_0.X.t15 11.2576
R6998 two_stage_opamp_dummy_magic_16_0.X.n0 two_stage_opamp_dummy_magic_16_0.X.t6 11.2576
R6999 two_stage_opamp_dummy_magic_16_0.X.n0 two_stage_opamp_dummy_magic_16_0.X.t10 11.2576
R7000 two_stage_opamp_dummy_magic_16_0.X.n52 two_stage_opamp_dummy_magic_16_0.X.n42 7.09425
R7001 two_stage_opamp_dummy_magic_16_0.X.n41 two_stage_opamp_dummy_magic_16_0.X.n40 6.38443
R7002 two_stage_opamp_dummy_magic_16_0.X.n10 two_stage_opamp_dummy_magic_16_0.X.n8 5.1255
R7003 two_stage_opamp_dummy_magic_16_0.X.n42 two_stage_opamp_dummy_magic_16_0.X.n41 0.938
R7004 two_stage_opamp_dummy_magic_16_0.X.n4 two_stage_opamp_dummy_magic_16_0.X.n2 0.6255
R7005 two_stage_opamp_dummy_magic_16_0.X.n6 two_stage_opamp_dummy_magic_16_0.X.n4 0.6255
R7006 two_stage_opamp_dummy_magic_16_0.X.n8 two_stage_opamp_dummy_magic_16_0.X.n6 0.6255
R7007 two_stage_opamp_dummy_magic_16_0.X.n34 two_stage_opamp_dummy_magic_16_0.X.n32 0.580857
R7008 two_stage_opamp_dummy_magic_16_0.X.n36 two_stage_opamp_dummy_magic_16_0.X.n34 0.580857
R7009 two_stage_opamp_dummy_magic_16_0.X.n38 two_stage_opamp_dummy_magic_16_0.X.n36 0.580857
R7010 two_stage_opamp_dummy_magic_16_0.X.n40 two_stage_opamp_dummy_magic_16_0.X.n38 0.580857
R7011 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n0 144.827
R7012 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n1 134.577
R7013 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t10 118.986
R7014 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n3 100.6
R7015 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n10 100.038
R7016 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n8 100.038
R7017 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n6 100.038
R7018 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n4 100.038
R7019 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n12 43.284
R7020 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n2 37.4067
R7021 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t11 24.0005
R7022 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t12 24.0005
R7023 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t13 24.0005
R7024 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t14 24.0005
R7025 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t7 8.0005
R7026 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t1 8.0005
R7027 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t6 8.0005
R7028 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t0 8.0005
R7029 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t5 8.0005
R7030 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t9 8.0005
R7031 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t3 8.0005
R7032 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t2 8.0005
R7033 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t4 8.0005
R7034 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t8 8.0005
R7035 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n11 5.6255
R7036 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n5 0.563
R7037 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n7 0.563
R7038 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n9 0.563
R7039 bgr_0.V_CMFB_S2 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n13 0.047375
R7040 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t9 525.38
R7041 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t4 525.38
R7042 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t2 358.288
R7043 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t3 358.288
R7044 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t5 281.168
R7045 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t8 281.168
R7046 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t7 281.168
R7047 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t6 281.168
R7048 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n4 244.214
R7049 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n0 244.214
R7050 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n6 166.019
R7051 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n2 166.019
R7052 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t1 116.013
R7053 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t0 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n7 116.013
R7054 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n5 77.1205
R7055 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n1 77.1205
R7056 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n3 18.0005
R7057 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t11 688.859
R7058 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t10 651.343
R7059 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t7 647.968
R7060 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n2 514.134
R7061 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n4 214.056
R7062 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t8 174.726
R7063 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t13 174.726
R7064 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t9 174.726
R7065 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t12 174.726
R7066 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n6 173.591
R7067 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n9 169.216
R7068 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n7 169.216
R7069 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n1 128.534
R7070 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n3 128.534
R7071 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t6 125.736
R7072 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n11 46.6411
R7073 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t2 13.1338
R7074 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t0 13.1338
R7075 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t5 13.1338
R7076 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t3 13.1338
R7077 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t1 13.1338
R7078 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t4 13.1338
R7079 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n10 10.0317
R7080 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n8 4.3755
R7081 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n5 3.03175
R7082 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n0 1.53175
R7083 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t13 610.534
R7084 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t16 610.534
R7085 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t31 433.8
R7086 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t22 433.8
R7087 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t29 433.8
R7088 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t19 433.8
R7089 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t27 433.8
R7090 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t17 433.8
R7091 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t25 433.8
R7092 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t14 433.8
R7093 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t21 433.8
R7094 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t12 433.8
R7095 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t23 433.8
R7096 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t30 433.8
R7097 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t20 433.8
R7098 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t28 433.8
R7099 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t18 433.8
R7100 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t26 433.8
R7101 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t15 433.8
R7102 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t24 433.8
R7103 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n0 339.836
R7104 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n1 339.834
R7105 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n2 339.272
R7106 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n5 287.264
R7107 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n27 221.262
R7108 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n25 176.733
R7109 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n24 176.733
R7110 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n23 176.733
R7111 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n22 176.733
R7112 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n21 176.733
R7113 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n20 176.733
R7114 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n19 176.733
R7115 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n18 176.733
R7116 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n9 176.733
R7117 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n10 176.733
R7118 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n11 176.733
R7119 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n12 176.733
R7120 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n13 176.733
R7121 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n14 176.733
R7122 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n15 176.733
R7123 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n16 176.733
R7124 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n7 112.076
R7125 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n28 68.4678
R7126 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_16_0.V_tail_gate.n29 62.839
R7127 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n26 54.6272
R7128 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n17 54.6272
R7129 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n8 53.2453
R7130 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n4 52.01
R7131 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_16_0.V_tail_gate.n6 51.6642
R7132 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t0 39.4005
R7133 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t11 39.4005
R7134 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t1 39.4005
R7135 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t6 39.4005
R7136 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t4 39.4005
R7137 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t5 39.4005
R7138 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t10 39.4005
R7139 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t7 39.4005
R7140 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t8 16.0005
R7141 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t2 16.0005
R7142 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t3 16.0005
R7143 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t9 16.0005
R7144 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n3 0.563
R7145 two_stage_opamp_dummy_magic_16_0.V_source.n30 two_stage_opamp_dummy_magic_16_0.V_source.t5 172.933
R7146 two_stage_opamp_dummy_magic_16_0.V_source.n13 two_stage_opamp_dummy_magic_16_0.V_source.n11 117.343
R7147 two_stage_opamp_dummy_magic_16_0.V_source.n6 two_stage_opamp_dummy_magic_16_0.V_source.n4 117.343
R7148 two_stage_opamp_dummy_magic_16_0.V_source.n19 two_stage_opamp_dummy_magic_16_0.V_source.n18 116.779
R7149 two_stage_opamp_dummy_magic_16_0.V_source.n17 two_stage_opamp_dummy_magic_16_0.V_source.n16 116.779
R7150 two_stage_opamp_dummy_magic_16_0.V_source.n15 two_stage_opamp_dummy_magic_16_0.V_source.n14 116.779
R7151 two_stage_opamp_dummy_magic_16_0.V_source.n13 two_stage_opamp_dummy_magic_16_0.V_source.n12 116.779
R7152 two_stage_opamp_dummy_magic_16_0.V_source.n10 two_stage_opamp_dummy_magic_16_0.V_source.n9 116.779
R7153 two_stage_opamp_dummy_magic_16_0.V_source.n8 two_stage_opamp_dummy_magic_16_0.V_source.n7 116.779
R7154 two_stage_opamp_dummy_magic_16_0.V_source.n6 two_stage_opamp_dummy_magic_16_0.V_source.n5 116.779
R7155 two_stage_opamp_dummy_magic_16_0.V_source.n21 two_stage_opamp_dummy_magic_16_0.V_source.n3 112.272
R7156 two_stage_opamp_dummy_magic_16_0.V_source.n2 two_stage_opamp_dummy_magic_16_0.V_source.n0 102.941
R7157 two_stage_opamp_dummy_magic_16_0.V_source.n38 two_stage_opamp_dummy_magic_16_0.V_source.n37 102.285
R7158 two_stage_opamp_dummy_magic_16_0.V_source.n36 two_stage_opamp_dummy_magic_16_0.V_source.n35 102.284
R7159 two_stage_opamp_dummy_magic_16_0.V_source.n34 two_stage_opamp_dummy_magic_16_0.V_source.n33 102.284
R7160 two_stage_opamp_dummy_magic_16_0.V_source.n32 two_stage_opamp_dummy_magic_16_0.V_source.n31 102.284
R7161 two_stage_opamp_dummy_magic_16_0.V_source.n30 two_stage_opamp_dummy_magic_16_0.V_source.n29 102.284
R7162 two_stage_opamp_dummy_magic_16_0.V_source.n28 two_stage_opamp_dummy_magic_16_0.V_source.n27 102.284
R7163 two_stage_opamp_dummy_magic_16_0.V_source.n26 two_stage_opamp_dummy_magic_16_0.V_source.n25 102.284
R7164 two_stage_opamp_dummy_magic_16_0.V_source.n2 two_stage_opamp_dummy_magic_16_0.V_source.n1 102.284
R7165 two_stage_opamp_dummy_magic_16_0.V_source.n23 two_stage_opamp_dummy_magic_16_0.V_source.n22 97.7845
R7166 two_stage_opamp_dummy_magic_16_0.V_source.n18 two_stage_opamp_dummy_magic_16_0.V_source.t27 16.0005
R7167 two_stage_opamp_dummy_magic_16_0.V_source.n18 two_stage_opamp_dummy_magic_16_0.V_source.t26 16.0005
R7168 two_stage_opamp_dummy_magic_16_0.V_source.n16 two_stage_opamp_dummy_magic_16_0.V_source.t29 16.0005
R7169 two_stage_opamp_dummy_magic_16_0.V_source.n16 two_stage_opamp_dummy_magic_16_0.V_source.t28 16.0005
R7170 two_stage_opamp_dummy_magic_16_0.V_source.n14 two_stage_opamp_dummy_magic_16_0.V_source.t35 16.0005
R7171 two_stage_opamp_dummy_magic_16_0.V_source.n14 two_stage_opamp_dummy_magic_16_0.V_source.t33 16.0005
R7172 two_stage_opamp_dummy_magic_16_0.V_source.n12 two_stage_opamp_dummy_magic_16_0.V_source.t31 16.0005
R7173 two_stage_opamp_dummy_magic_16_0.V_source.n12 two_stage_opamp_dummy_magic_16_0.V_source.t40 16.0005
R7174 two_stage_opamp_dummy_magic_16_0.V_source.n11 two_stage_opamp_dummy_magic_16_0.V_source.t37 16.0005
R7175 two_stage_opamp_dummy_magic_16_0.V_source.n11 two_stage_opamp_dummy_magic_16_0.V_source.t3 16.0005
R7176 two_stage_opamp_dummy_magic_16_0.V_source.n9 two_stage_opamp_dummy_magic_16_0.V_source.t4 16.0005
R7177 two_stage_opamp_dummy_magic_16_0.V_source.n9 two_stage_opamp_dummy_magic_16_0.V_source.t0 16.0005
R7178 two_stage_opamp_dummy_magic_16_0.V_source.n7 two_stage_opamp_dummy_magic_16_0.V_source.t39 16.0005
R7179 two_stage_opamp_dummy_magic_16_0.V_source.n7 two_stage_opamp_dummy_magic_16_0.V_source.t2 16.0005
R7180 two_stage_opamp_dummy_magic_16_0.V_source.n5 two_stage_opamp_dummy_magic_16_0.V_source.t36 16.0005
R7181 two_stage_opamp_dummy_magic_16_0.V_source.n5 two_stage_opamp_dummy_magic_16_0.V_source.t6 16.0005
R7182 two_stage_opamp_dummy_magic_16_0.V_source.n4 two_stage_opamp_dummy_magic_16_0.V_source.t30 16.0005
R7183 two_stage_opamp_dummy_magic_16_0.V_source.n4 two_stage_opamp_dummy_magic_16_0.V_source.t1 16.0005
R7184 two_stage_opamp_dummy_magic_16_0.V_source.n3 two_stage_opamp_dummy_magic_16_0.V_source.t25 16.0005
R7185 two_stage_opamp_dummy_magic_16_0.V_source.n3 two_stage_opamp_dummy_magic_16_0.V_source.t34 16.0005
R7186 two_stage_opamp_dummy_magic_16_0.V_source.n35 two_stage_opamp_dummy_magic_16_0.V_source.t16 9.6005
R7187 two_stage_opamp_dummy_magic_16_0.V_source.n35 two_stage_opamp_dummy_magic_16_0.V_source.t23 9.6005
R7188 two_stage_opamp_dummy_magic_16_0.V_source.n33 two_stage_opamp_dummy_magic_16_0.V_source.t12 9.6005
R7189 two_stage_opamp_dummy_magic_16_0.V_source.n33 two_stage_opamp_dummy_magic_16_0.V_source.t20 9.6005
R7190 two_stage_opamp_dummy_magic_16_0.V_source.n31 two_stage_opamp_dummy_magic_16_0.V_source.t10 9.6005
R7191 two_stage_opamp_dummy_magic_16_0.V_source.n31 two_stage_opamp_dummy_magic_16_0.V_source.t18 9.6005
R7192 two_stage_opamp_dummy_magic_16_0.V_source.n29 two_stage_opamp_dummy_magic_16_0.V_source.t8 9.6005
R7193 two_stage_opamp_dummy_magic_16_0.V_source.n29 two_stage_opamp_dummy_magic_16_0.V_source.t15 9.6005
R7194 two_stage_opamp_dummy_magic_16_0.V_source.n27 two_stage_opamp_dummy_magic_16_0.V_source.t17 9.6005
R7195 two_stage_opamp_dummy_magic_16_0.V_source.n27 two_stage_opamp_dummy_magic_16_0.V_source.t7 9.6005
R7196 two_stage_opamp_dummy_magic_16_0.V_source.n25 two_stage_opamp_dummy_magic_16_0.V_source.t19 9.6005
R7197 two_stage_opamp_dummy_magic_16_0.V_source.n25 two_stage_opamp_dummy_magic_16_0.V_source.t9 9.6005
R7198 two_stage_opamp_dummy_magic_16_0.V_source.n22 two_stage_opamp_dummy_magic_16_0.V_source.t22 9.6005
R7199 two_stage_opamp_dummy_magic_16_0.V_source.n22 two_stage_opamp_dummy_magic_16_0.V_source.t11 9.6005
R7200 two_stage_opamp_dummy_magic_16_0.V_source.n1 two_stage_opamp_dummy_magic_16_0.V_source.t21 9.6005
R7201 two_stage_opamp_dummy_magic_16_0.V_source.n1 two_stage_opamp_dummy_magic_16_0.V_source.t13 9.6005
R7202 two_stage_opamp_dummy_magic_16_0.V_source.n0 two_stage_opamp_dummy_magic_16_0.V_source.t32 9.6005
R7203 two_stage_opamp_dummy_magic_16_0.V_source.n0 two_stage_opamp_dummy_magic_16_0.V_source.t38 9.6005
R7204 two_stage_opamp_dummy_magic_16_0.V_source.n38 two_stage_opamp_dummy_magic_16_0.V_source.t14 9.6005
R7205 two_stage_opamp_dummy_magic_16_0.V_source.t24 two_stage_opamp_dummy_magic_16_0.V_source.n38 9.6005
R7206 two_stage_opamp_dummy_magic_16_0.V_source.n21 two_stage_opamp_dummy_magic_16_0.V_source.n20 4.5005
R7207 two_stage_opamp_dummy_magic_16_0.V_source.n24 two_stage_opamp_dummy_magic_16_0.V_source.n23 4.5005
R7208 two_stage_opamp_dummy_magic_16_0.V_source.n20 two_stage_opamp_dummy_magic_16_0.V_source.n19 3.6255
R7209 two_stage_opamp_dummy_magic_16_0.V_source.n23 two_stage_opamp_dummy_magic_16_0.V_source.n21 0.774806
R7210 two_stage_opamp_dummy_magic_16_0.V_source.n32 two_stage_opamp_dummy_magic_16_0.V_source.n30 0.563
R7211 two_stage_opamp_dummy_magic_16_0.V_source.n34 two_stage_opamp_dummy_magic_16_0.V_source.n32 0.563
R7212 two_stage_opamp_dummy_magic_16_0.V_source.n36 two_stage_opamp_dummy_magic_16_0.V_source.n34 0.563
R7213 two_stage_opamp_dummy_magic_16_0.V_source.n37 two_stage_opamp_dummy_magic_16_0.V_source.n36 0.563
R7214 two_stage_opamp_dummy_magic_16_0.V_source.n15 two_stage_opamp_dummy_magic_16_0.V_source.n13 0.563
R7215 two_stage_opamp_dummy_magic_16_0.V_source.n17 two_stage_opamp_dummy_magic_16_0.V_source.n15 0.563
R7216 two_stage_opamp_dummy_magic_16_0.V_source.n19 two_stage_opamp_dummy_magic_16_0.V_source.n17 0.563
R7217 two_stage_opamp_dummy_magic_16_0.V_source.n8 two_stage_opamp_dummy_magic_16_0.V_source.n6 0.563
R7218 two_stage_opamp_dummy_magic_16_0.V_source.n10 two_stage_opamp_dummy_magic_16_0.V_source.n8 0.563
R7219 two_stage_opamp_dummy_magic_16_0.V_source.n20 two_stage_opamp_dummy_magic_16_0.V_source.n10 0.563
R7220 two_stage_opamp_dummy_magic_16_0.V_source.n24 two_stage_opamp_dummy_magic_16_0.V_source.n2 0.563
R7221 two_stage_opamp_dummy_magic_16_0.V_source.n26 two_stage_opamp_dummy_magic_16_0.V_source.n24 0.563
R7222 two_stage_opamp_dummy_magic_16_0.V_source.n28 two_stage_opamp_dummy_magic_16_0.V_source.n26 0.563
R7223 two_stage_opamp_dummy_magic_16_0.V_source.n37 two_stage_opamp_dummy_magic_16_0.V_source.n28 0.563
R7224 bgr_0.Vin+.n3 bgr_0.Vin+.n2 526.183
R7225 bgr_0.Vin+.n1 bgr_0.Vin+.n0 514.134
R7226 bgr_0.Vin+.n0 bgr_0.Vin+.t8 303.259
R7227 bgr_0.Vin+.n5 bgr_0.Vin+.n3 227.169
R7228 bgr_0.Vin+.n0 bgr_0.Vin+.t9 174.726
R7229 bgr_0.Vin+.n1 bgr_0.Vin+.t6 174.726
R7230 bgr_0.Vin+.n2 bgr_0.Vin+.t10 174.726
R7231 bgr_0.Vin+.n7 bgr_0.Vin+.n6 168.435
R7232 bgr_0.Vin+.n5 bgr_0.Vin+.n4 168.435
R7233 bgr_0.Vin+.n8 bgr_0.Vin+.t1 158.989
R7234 bgr_0.Vin+.n2 bgr_0.Vin+.n1 128.534
R7235 bgr_0.Vin+.t0 bgr_0.Vin+.n8 119.067
R7236 bgr_0.Vin+.n3 bgr_0.Vin+.t7 96.4005
R7237 bgr_0.Vin+.n8 bgr_0.Vin+.n7 35.0317
R7238 bgr_0.Vin+.n6 bgr_0.Vin+.t2 13.1338
R7239 bgr_0.Vin+.n6 bgr_0.Vin+.t5 13.1338
R7240 bgr_0.Vin+.n4 bgr_0.Vin+.t4 13.1338
R7241 bgr_0.Vin+.n4 bgr_0.Vin+.t3 13.1338
R7242 bgr_0.Vin+.n7 bgr_0.Vin+.n5 2.1255
R7243 two_stage_opamp_dummy_magic_16_0.VD3.n28 two_stage_opamp_dummy_magic_16_0.VD3.t30 652.076
R7244 two_stage_opamp_dummy_magic_16_0.VD3.n59 two_stage_opamp_dummy_magic_16_0.VD3.t33 652.076
R7245 two_stage_opamp_dummy_magic_16_0.VD3.n58 two_stage_opamp_dummy_magic_16_0.VD3.n11 585
R7246 two_stage_opamp_dummy_magic_16_0.VD3.n42 two_stage_opamp_dummy_magic_16_0.VD3.n29 585
R7247 two_stage_opamp_dummy_magic_16_0.VD3.n46 two_stage_opamp_dummy_magic_16_0.VD3.n11 290.233
R7248 two_stage_opamp_dummy_magic_16_0.VD3.n52 two_stage_opamp_dummy_magic_16_0.VD3.n11 290.233
R7249 two_stage_opamp_dummy_magic_16_0.VD3.n47 two_stage_opamp_dummy_magic_16_0.VD3.n11 290.233
R7250 two_stage_opamp_dummy_magic_16_0.VD3.n40 two_stage_opamp_dummy_magic_16_0.VD3.n29 290.233
R7251 two_stage_opamp_dummy_magic_16_0.VD3.n35 two_stage_opamp_dummy_magic_16_0.VD3.n29 290.233
R7252 two_stage_opamp_dummy_magic_16_0.VD3.n30 two_stage_opamp_dummy_magic_16_0.VD3.n29 290.233
R7253 two_stage_opamp_dummy_magic_16_0.VD3.n47 two_stage_opamp_dummy_magic_16_0.VD3.n15 242.903
R7254 two_stage_opamp_dummy_magic_16_0.VD3.n30 two_stage_opamp_dummy_magic_16_0.VD3.n18 242.903
R7255 two_stage_opamp_dummy_magic_16_0.VD3.n58 two_stage_opamp_dummy_magic_16_0.VD3.n57 238.367
R7256 two_stage_opamp_dummy_magic_16_0.VD3.n13 two_stage_opamp_dummy_magic_16_0.VD3.n12 185
R7257 two_stage_opamp_dummy_magic_16_0.VD3.n55 two_stage_opamp_dummy_magic_16_0.VD3.n54 185
R7258 two_stage_opamp_dummy_magic_16_0.VD3.n56 two_stage_opamp_dummy_magic_16_0.VD3.n55 185
R7259 two_stage_opamp_dummy_magic_16_0.VD3.n53 two_stage_opamp_dummy_magic_16_0.VD3.n45 185
R7260 two_stage_opamp_dummy_magic_16_0.VD3.n51 two_stage_opamp_dummy_magic_16_0.VD3.n50 185
R7261 two_stage_opamp_dummy_magic_16_0.VD3.n49 two_stage_opamp_dummy_magic_16_0.VD3.n48 185
R7262 two_stage_opamp_dummy_magic_16_0.VD3.n43 two_stage_opamp_dummy_magic_16_0.VD3.n42 185
R7263 two_stage_opamp_dummy_magic_16_0.VD3.n44 two_stage_opamp_dummy_magic_16_0.VD3.n43 185
R7264 two_stage_opamp_dummy_magic_16_0.VD3.n41 two_stage_opamp_dummy_magic_16_0.VD3.n19 185
R7265 two_stage_opamp_dummy_magic_16_0.VD3.n39 two_stage_opamp_dummy_magic_16_0.VD3.n38 185
R7266 two_stage_opamp_dummy_magic_16_0.VD3.n37 two_stage_opamp_dummy_magic_16_0.VD3.n36 185
R7267 two_stage_opamp_dummy_magic_16_0.VD3.n34 two_stage_opamp_dummy_magic_16_0.VD3.n33 185
R7268 two_stage_opamp_dummy_magic_16_0.VD3.n32 two_stage_opamp_dummy_magic_16_0.VD3.n31 185
R7269 two_stage_opamp_dummy_magic_16_0.VD3.n56 two_stage_opamp_dummy_magic_16_0.VD3.t34 170.513
R7270 two_stage_opamp_dummy_magic_16_0.VD3.t31 two_stage_opamp_dummy_magic_16_0.VD3.n44 170.513
R7271 two_stage_opamp_dummy_magic_16_0.VD3.n2 two_stage_opamp_dummy_magic_16_0.VD3.n0 163.626
R7272 two_stage_opamp_dummy_magic_16_0.VD3.n8 two_stage_opamp_dummy_magic_16_0.VD3.n7 163.001
R7273 two_stage_opamp_dummy_magic_16_0.VD3.n6 two_stage_opamp_dummy_magic_16_0.VD3.n5 163.001
R7274 two_stage_opamp_dummy_magic_16_0.VD3.n4 two_stage_opamp_dummy_magic_16_0.VD3.n3 163.001
R7275 two_stage_opamp_dummy_magic_16_0.VD3.n2 two_stage_opamp_dummy_magic_16_0.VD3.n1 163.001
R7276 two_stage_opamp_dummy_magic_16_0.VD3.n62 two_stage_opamp_dummy_magic_16_0.VD3.n61 162.999
R7277 two_stage_opamp_dummy_magic_16_0.VD3.n10 two_stage_opamp_dummy_magic_16_0.VD3.n9 159.803
R7278 two_stage_opamp_dummy_magic_16_0.VD3.n21 two_stage_opamp_dummy_magic_16_0.VD3.n20 159.803
R7279 two_stage_opamp_dummy_magic_16_0.VD3.n23 two_stage_opamp_dummy_magic_16_0.VD3.n22 159.803
R7280 two_stage_opamp_dummy_magic_16_0.VD3.n25 two_stage_opamp_dummy_magic_16_0.VD3.n24 159.803
R7281 two_stage_opamp_dummy_magic_16_0.VD3.n27 two_stage_opamp_dummy_magic_16_0.VD3.n26 159.803
R7282 two_stage_opamp_dummy_magic_16_0.VD3.n55 two_stage_opamp_dummy_magic_16_0.VD3.n13 150
R7283 two_stage_opamp_dummy_magic_16_0.VD3.n55 two_stage_opamp_dummy_magic_16_0.VD3.n45 150
R7284 two_stage_opamp_dummy_magic_16_0.VD3.n50 two_stage_opamp_dummy_magic_16_0.VD3.n49 150
R7285 two_stage_opamp_dummy_magic_16_0.VD3.n43 two_stage_opamp_dummy_magic_16_0.VD3.n19 150
R7286 two_stage_opamp_dummy_magic_16_0.VD3.n38 two_stage_opamp_dummy_magic_16_0.VD3.n37 150
R7287 two_stage_opamp_dummy_magic_16_0.VD3.n33 two_stage_opamp_dummy_magic_16_0.VD3.n32 150
R7288 two_stage_opamp_dummy_magic_16_0.VD3.t34 two_stage_opamp_dummy_magic_16_0.VD3.t4 146.155
R7289 two_stage_opamp_dummy_magic_16_0.VD3.t4 two_stage_opamp_dummy_magic_16_0.VD3.t6 146.155
R7290 two_stage_opamp_dummy_magic_16_0.VD3.t6 two_stage_opamp_dummy_magic_16_0.VD3.t0 146.155
R7291 two_stage_opamp_dummy_magic_16_0.VD3.t0 two_stage_opamp_dummy_magic_16_0.VD3.t2 146.155
R7292 two_stage_opamp_dummy_magic_16_0.VD3.t2 two_stage_opamp_dummy_magic_16_0.VD3.t10 146.155
R7293 two_stage_opamp_dummy_magic_16_0.VD3.t10 two_stage_opamp_dummy_magic_16_0.VD3.t12 146.155
R7294 two_stage_opamp_dummy_magic_16_0.VD3.t12 two_stage_opamp_dummy_magic_16_0.VD3.t16 146.155
R7295 two_stage_opamp_dummy_magic_16_0.VD3.t16 two_stage_opamp_dummy_magic_16_0.VD3.t36 146.155
R7296 two_stage_opamp_dummy_magic_16_0.VD3.t36 two_stage_opamp_dummy_magic_16_0.VD3.t14 146.155
R7297 two_stage_opamp_dummy_magic_16_0.VD3.t14 two_stage_opamp_dummy_magic_16_0.VD3.t8 146.155
R7298 two_stage_opamp_dummy_magic_16_0.VD3.t8 two_stage_opamp_dummy_magic_16_0.VD3.t31 146.155
R7299 two_stage_opamp_dummy_magic_16_0.VD3.n57 two_stage_opamp_dummy_magic_16_0.VD3.n56 65.8183
R7300 two_stage_opamp_dummy_magic_16_0.VD3.n56 two_stage_opamp_dummy_magic_16_0.VD3.n14 65.8183
R7301 two_stage_opamp_dummy_magic_16_0.VD3.n56 two_stage_opamp_dummy_magic_16_0.VD3.n15 65.8183
R7302 two_stage_opamp_dummy_magic_16_0.VD3.n44 two_stage_opamp_dummy_magic_16_0.VD3.n16 65.8183
R7303 two_stage_opamp_dummy_magic_16_0.VD3.n44 two_stage_opamp_dummy_magic_16_0.VD3.n17 65.8183
R7304 two_stage_opamp_dummy_magic_16_0.VD3.n44 two_stage_opamp_dummy_magic_16_0.VD3.n18 65.8183
R7305 two_stage_opamp_dummy_magic_16_0.VD3.n45 two_stage_opamp_dummy_magic_16_0.VD3.n14 53.3664
R7306 two_stage_opamp_dummy_magic_16_0.VD3.n49 two_stage_opamp_dummy_magic_16_0.VD3.n15 53.3664
R7307 two_stage_opamp_dummy_magic_16_0.VD3.n57 two_stage_opamp_dummy_magic_16_0.VD3.n13 53.3664
R7308 two_stage_opamp_dummy_magic_16_0.VD3.n50 two_stage_opamp_dummy_magic_16_0.VD3.n14 53.3664
R7309 two_stage_opamp_dummy_magic_16_0.VD3.n19 two_stage_opamp_dummy_magic_16_0.VD3.n16 53.3664
R7310 two_stage_opamp_dummy_magic_16_0.VD3.n37 two_stage_opamp_dummy_magic_16_0.VD3.n17 53.3664
R7311 two_stage_opamp_dummy_magic_16_0.VD3.n32 two_stage_opamp_dummy_magic_16_0.VD3.n18 53.3664
R7312 two_stage_opamp_dummy_magic_16_0.VD3.n38 two_stage_opamp_dummy_magic_16_0.VD3.n16 53.3664
R7313 two_stage_opamp_dummy_magic_16_0.VD3.n33 two_stage_opamp_dummy_magic_16_0.VD3.n17 53.3664
R7314 two_stage_opamp_dummy_magic_16_0.VD3.n59 two_stage_opamp_dummy_magic_16_0.VD3.n58 22.8576
R7315 two_stage_opamp_dummy_magic_16_0.VD3.n42 two_stage_opamp_dummy_magic_16_0.VD3.n28 22.8576
R7316 two_stage_opamp_dummy_magic_16_0.VD3.n28 two_stage_opamp_dummy_magic_16_0.VD3.n27 14.4255
R7317 two_stage_opamp_dummy_magic_16_0.VD3.n60 two_stage_opamp_dummy_magic_16_0.VD3.n59 13.8005
R7318 two_stage_opamp_dummy_magic_16_0.VD3.n61 two_stage_opamp_dummy_magic_16_0.VD3.n60 13.688
R7319 two_stage_opamp_dummy_magic_16_0.VD3.n9 two_stage_opamp_dummy_magic_16_0.VD3.t5 11.2576
R7320 two_stage_opamp_dummy_magic_16_0.VD3.n9 two_stage_opamp_dummy_magic_16_0.VD3.t7 11.2576
R7321 two_stage_opamp_dummy_magic_16_0.VD3.n20 two_stage_opamp_dummy_magic_16_0.VD3.t1 11.2576
R7322 two_stage_opamp_dummy_magic_16_0.VD3.n20 two_stage_opamp_dummy_magic_16_0.VD3.t3 11.2576
R7323 two_stage_opamp_dummy_magic_16_0.VD3.n22 two_stage_opamp_dummy_magic_16_0.VD3.t11 11.2576
R7324 two_stage_opamp_dummy_magic_16_0.VD3.n22 two_stage_opamp_dummy_magic_16_0.VD3.t13 11.2576
R7325 two_stage_opamp_dummy_magic_16_0.VD3.n24 two_stage_opamp_dummy_magic_16_0.VD3.t17 11.2576
R7326 two_stage_opamp_dummy_magic_16_0.VD3.n24 two_stage_opamp_dummy_magic_16_0.VD3.t37 11.2576
R7327 two_stage_opamp_dummy_magic_16_0.VD3.n26 two_stage_opamp_dummy_magic_16_0.VD3.t15 11.2576
R7328 two_stage_opamp_dummy_magic_16_0.VD3.n26 two_stage_opamp_dummy_magic_16_0.VD3.t9 11.2576
R7329 two_stage_opamp_dummy_magic_16_0.VD3.n11 two_stage_opamp_dummy_magic_16_0.VD3.t35 11.2576
R7330 two_stage_opamp_dummy_magic_16_0.VD3.n29 two_stage_opamp_dummy_magic_16_0.VD3.t32 11.2576
R7331 two_stage_opamp_dummy_magic_16_0.VD3.n7 two_stage_opamp_dummy_magic_16_0.VD3.t22 11.2576
R7332 two_stage_opamp_dummy_magic_16_0.VD3.n7 two_stage_opamp_dummy_magic_16_0.VD3.t25 11.2576
R7333 two_stage_opamp_dummy_magic_16_0.VD3.n5 two_stage_opamp_dummy_magic_16_0.VD3.t19 11.2576
R7334 two_stage_opamp_dummy_magic_16_0.VD3.n5 two_stage_opamp_dummy_magic_16_0.VD3.t20 11.2576
R7335 two_stage_opamp_dummy_magic_16_0.VD3.n3 two_stage_opamp_dummy_magic_16_0.VD3.t26 11.2576
R7336 two_stage_opamp_dummy_magic_16_0.VD3.n3 two_stage_opamp_dummy_magic_16_0.VD3.t18 11.2576
R7337 two_stage_opamp_dummy_magic_16_0.VD3.n1 two_stage_opamp_dummy_magic_16_0.VD3.t21 11.2576
R7338 two_stage_opamp_dummy_magic_16_0.VD3.n1 two_stage_opamp_dummy_magic_16_0.VD3.t24 11.2576
R7339 two_stage_opamp_dummy_magic_16_0.VD3.n0 two_stage_opamp_dummy_magic_16_0.VD3.t29 11.2576
R7340 two_stage_opamp_dummy_magic_16_0.VD3.n0 two_stage_opamp_dummy_magic_16_0.VD3.t23 11.2576
R7341 two_stage_opamp_dummy_magic_16_0.VD3.t27 two_stage_opamp_dummy_magic_16_0.VD3.n62 11.2576
R7342 two_stage_opamp_dummy_magic_16_0.VD3.n62 two_stage_opamp_dummy_magic_16_0.VD3.t28 11.2576
R7343 two_stage_opamp_dummy_magic_16_0.VD3.n58 two_stage_opamp_dummy_magic_16_0.VD3.n12 9.14336
R7344 two_stage_opamp_dummy_magic_16_0.VD3.n54 two_stage_opamp_dummy_magic_16_0.VD3.n53 9.14336
R7345 two_stage_opamp_dummy_magic_16_0.VD3.n51 two_stage_opamp_dummy_magic_16_0.VD3.n48 9.14336
R7346 two_stage_opamp_dummy_magic_16_0.VD3.n42 two_stage_opamp_dummy_magic_16_0.VD3.n41 9.14336
R7347 two_stage_opamp_dummy_magic_16_0.VD3.n39 two_stage_opamp_dummy_magic_16_0.VD3.n36 9.14336
R7348 two_stage_opamp_dummy_magic_16_0.VD3.n34 two_stage_opamp_dummy_magic_16_0.VD3.n31 9.14336
R7349 two_stage_opamp_dummy_magic_16_0.VD3.n46 two_stage_opamp_dummy_magic_16_0.VD3.n12 4.53698
R7350 two_stage_opamp_dummy_magic_16_0.VD3.n53 two_stage_opamp_dummy_magic_16_0.VD3.n52 4.53698
R7351 two_stage_opamp_dummy_magic_16_0.VD3.n48 two_stage_opamp_dummy_magic_16_0.VD3.n47 4.53698
R7352 two_stage_opamp_dummy_magic_16_0.VD3.n54 two_stage_opamp_dummy_magic_16_0.VD3.n46 4.53698
R7353 two_stage_opamp_dummy_magic_16_0.VD3.n52 two_stage_opamp_dummy_magic_16_0.VD3.n51 4.53698
R7354 two_stage_opamp_dummy_magic_16_0.VD3.n41 two_stage_opamp_dummy_magic_16_0.VD3.n40 4.53698
R7355 two_stage_opamp_dummy_magic_16_0.VD3.n36 two_stage_opamp_dummy_magic_16_0.VD3.n35 4.53698
R7356 two_stage_opamp_dummy_magic_16_0.VD3.n31 two_stage_opamp_dummy_magic_16_0.VD3.n30 4.53698
R7357 two_stage_opamp_dummy_magic_16_0.VD3.n40 two_stage_opamp_dummy_magic_16_0.VD3.n39 4.53698
R7358 two_stage_opamp_dummy_magic_16_0.VD3.n35 two_stage_opamp_dummy_magic_16_0.VD3.n34 4.53698
R7359 two_stage_opamp_dummy_magic_16_0.VD3.n27 two_stage_opamp_dummy_magic_16_0.VD3.n25 0.6255
R7360 two_stage_opamp_dummy_magic_16_0.VD3.n25 two_stage_opamp_dummy_magic_16_0.VD3.n23 0.6255
R7361 two_stage_opamp_dummy_magic_16_0.VD3.n23 two_stage_opamp_dummy_magic_16_0.VD3.n21 0.6255
R7362 two_stage_opamp_dummy_magic_16_0.VD3.n21 two_stage_opamp_dummy_magic_16_0.VD3.n10 0.6255
R7363 two_stage_opamp_dummy_magic_16_0.VD3.n60 two_stage_opamp_dummy_magic_16_0.VD3.n10 0.6255
R7364 two_stage_opamp_dummy_magic_16_0.VD3.n4 two_stage_opamp_dummy_magic_16_0.VD3.n2 0.6255
R7365 two_stage_opamp_dummy_magic_16_0.VD3.n6 two_stage_opamp_dummy_magic_16_0.VD3.n4 0.6255
R7366 two_stage_opamp_dummy_magic_16_0.VD3.n8 two_stage_opamp_dummy_magic_16_0.VD3.n6 0.6255
R7367 two_stage_opamp_dummy_magic_16_0.VD3.n61 two_stage_opamp_dummy_magic_16_0.VD3.n8 0.6255
R7368 bgr_0.V_mir1.n20 bgr_0.V_mir1.n19 325.473
R7369 bgr_0.V_mir1.n13 bgr_0.V_mir1.n12 325.473
R7370 bgr_0.V_mir1.n4 bgr_0.V_mir1.n3 325.473
R7371 bgr_0.V_mir1.n16 bgr_0.V_mir1.t19 310.488
R7372 bgr_0.V_mir1.n9 bgr_0.V_mir1.t21 310.488
R7373 bgr_0.V_mir1.n0 bgr_0.V_mir1.t20 310.488
R7374 bgr_0.V_mir1.n7 bgr_0.V_mir1.t12 278.312
R7375 bgr_0.V_mir1.n7 bgr_0.V_mir1.n6 228.939
R7376 bgr_0.V_mir1.n8 bgr_0.V_mir1.n5 224.439
R7377 bgr_0.V_mir1.n18 bgr_0.V_mir1.t6 184.097
R7378 bgr_0.V_mir1.n11 bgr_0.V_mir1.t2 184.097
R7379 bgr_0.V_mir1.n2 bgr_0.V_mir1.t0 184.097
R7380 bgr_0.V_mir1.n17 bgr_0.V_mir1.n16 167.094
R7381 bgr_0.V_mir1.n10 bgr_0.V_mir1.n9 167.094
R7382 bgr_0.V_mir1.n1 bgr_0.V_mir1.n0 167.094
R7383 bgr_0.V_mir1.n13 bgr_0.V_mir1.n11 152
R7384 bgr_0.V_mir1.n4 bgr_0.V_mir1.n2 152
R7385 bgr_0.V_mir1.n19 bgr_0.V_mir1.n18 152
R7386 bgr_0.V_mir1.n16 bgr_0.V_mir1.t22 120.501
R7387 bgr_0.V_mir1.n17 bgr_0.V_mir1.t10 120.501
R7388 bgr_0.V_mir1.n9 bgr_0.V_mir1.t17 120.501
R7389 bgr_0.V_mir1.n10 bgr_0.V_mir1.t8 120.501
R7390 bgr_0.V_mir1.n0 bgr_0.V_mir1.t18 120.501
R7391 bgr_0.V_mir1.n1 bgr_0.V_mir1.t4 120.501
R7392 bgr_0.V_mir1.n6 bgr_0.V_mir1.t15 48.0005
R7393 bgr_0.V_mir1.n6 bgr_0.V_mir1.t16 48.0005
R7394 bgr_0.V_mir1.n5 bgr_0.V_mir1.t14 48.0005
R7395 bgr_0.V_mir1.n5 bgr_0.V_mir1.t13 48.0005
R7396 bgr_0.V_mir1.n18 bgr_0.V_mir1.n17 40.7027
R7397 bgr_0.V_mir1.n11 bgr_0.V_mir1.n10 40.7027
R7398 bgr_0.V_mir1.n2 bgr_0.V_mir1.n1 40.7027
R7399 bgr_0.V_mir1.n12 bgr_0.V_mir1.t3 39.4005
R7400 bgr_0.V_mir1.n12 bgr_0.V_mir1.t9 39.4005
R7401 bgr_0.V_mir1.n3 bgr_0.V_mir1.t1 39.4005
R7402 bgr_0.V_mir1.n3 bgr_0.V_mir1.t5 39.4005
R7403 bgr_0.V_mir1.n20 bgr_0.V_mir1.t7 39.4005
R7404 bgr_0.V_mir1.t11 bgr_0.V_mir1.n20 39.4005
R7405 bgr_0.V_mir1.n15 bgr_0.V_mir1.n4 15.8005
R7406 bgr_0.V_mir1.n19 bgr_0.V_mir1.n15 15.8005
R7407 bgr_0.V_mir1.n14 bgr_0.V_mir1.n13 9.3005
R7408 bgr_0.V_mir1.n8 bgr_0.V_mir1.n7 5.8755
R7409 bgr_0.V_mir1.n15 bgr_0.V_mir1.n14 4.5005
R7410 bgr_0.V_mir1.n14 bgr_0.V_mir1.n8 0.78175
R7411 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.t13 354.854
R7412 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t21 346.8
R7413 bgr_0.1st_Vout_1.n20 bgr_0.1st_Vout_1.n19 339.522
R7414 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.n6 339.522
R7415 bgr_0.1st_Vout_1.n15 bgr_0.1st_Vout_1.n14 335.022
R7416 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t10 275.909
R7417 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.n10 227.909
R7418 bgr_0.1st_Vout_1.n13 bgr_0.1st_Vout_1.n12 222.034
R7419 bgr_0.1st_Vout_1.n17 bgr_0.1st_Vout_1.t22 184.097
R7420 bgr_0.1st_Vout_1.n17 bgr_0.1st_Vout_1.t32 184.097
R7421 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t16 184.097
R7422 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t36 184.097
R7423 bgr_0.1st_Vout_1.n18 bgr_0.1st_Vout_1.n17 166.05
R7424 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.n8 166.05
R7425 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.n4 54.2759
R7426 bgr_0.1st_Vout_1.n12 bgr_0.1st_Vout_1.t6 48.0005
R7427 bgr_0.1st_Vout_1.n12 bgr_0.1st_Vout_1.t7 48.0005
R7428 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t8 48.0005
R7429 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t9 48.0005
R7430 bgr_0.1st_Vout_1.n19 bgr_0.1st_Vout_1.t4 39.4005
R7431 bgr_0.1st_Vout_1.n19 bgr_0.1st_Vout_1.t2 39.4005
R7432 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t0 39.4005
R7433 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t3 39.4005
R7434 bgr_0.1st_Vout_1.n14 bgr_0.1st_Vout_1.t5 39.4005
R7435 bgr_0.1st_Vout_1.n14 bgr_0.1st_Vout_1.t1 39.4005
R7436 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t11 4.8295
R7437 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t29 4.8295
R7438 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t31 4.8295
R7439 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t20 4.8295
R7440 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t24 4.8295
R7441 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t14 4.8295
R7442 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t30 4.8295
R7443 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t18 4.8295
R7444 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t23 4.8295
R7445 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t15 4.5005
R7446 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t35 4.5005
R7447 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t34 4.5005
R7448 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t28 4.5005
R7449 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t27 4.5005
R7450 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t19 4.5005
R7451 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t33 4.5005
R7452 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t26 4.5005
R7453 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t25 4.5005
R7454 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t17 4.5005
R7455 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t12 4.5005
R7456 bgr_0.1st_Vout_1.n13 bgr_0.1st_Vout_1.n11 4.5005
R7457 bgr_0.1st_Vout_1.n16 bgr_0.1st_Vout_1.n15 4.5005
R7458 bgr_0.1st_Vout_1.n20 bgr_0.1st_Vout_1.n18 1.3755
R7459 bgr_0.1st_Vout_1.n16 bgr_0.1st_Vout_1.n9 1.3755
R7460 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.n5 1.188
R7461 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n2 0.8935
R7462 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.n0 0.8935
R7463 bgr_0.1st_Vout_1.n15 bgr_0.1st_Vout_1.n13 0.78175
R7464 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.n3 0.6585
R7465 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.n1 0.6585
R7466 bgr_0.1st_Vout_1.n18 bgr_0.1st_Vout_1.n16 0.6255
R7467 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.n7 0.6255
R7468 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n20 0.438
R7469 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.t33 355.293
R7470 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t34 346.8
R7471 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.n12 339.522
R7472 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n5 339.522
R7473 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n10 335.022
R7474 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t3 275.909
R7475 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.n7 227.909
R7476 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n9 222.034
R7477 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.t13 184.097
R7478 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.t24 184.097
R7479 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t16 184.097
R7480 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t27 184.097
R7481 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n11 166.05
R7482 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n6 166.05
R7483 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n4 52.9634
R7484 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.t4 48.0005
R7485 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.t10 48.0005
R7486 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t5 48.0005
R7487 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t8 48.0005
R7488 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t9 39.4005
R7489 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t1 39.4005
R7490 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t6 39.4005
R7491 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t7 39.4005
R7492 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.t2 39.4005
R7493 bgr_0.1st_Vout_2.t0 bgr_0.1st_Vout_2.n13 39.4005
R7494 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n3 5.28175
R7495 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t17 4.8295
R7496 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t35 4.8295
R7497 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t11 4.8295
R7498 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t26 4.8295
R7499 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t30 4.8295
R7500 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t19 4.8295
R7501 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t36 4.8295
R7502 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t25 4.8295
R7503 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t18 4.8295
R7504 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n8 4.5005
R7505 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t12 4.5005
R7506 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t32 4.5005
R7507 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t31 4.5005
R7508 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t23 4.5005
R7509 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t22 4.5005
R7510 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t15 4.5005
R7511 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t29 4.5005
R7512 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t21 4.5005
R7513 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t28 4.5005
R7514 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t20 4.5005
R7515 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t14 4.5005
R7516 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n0 3.188
R7517 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.n2 3.1025
R7518 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.n1 2.0005
R7519 bgr_0.cap_res2.t0 bgr_0.cap_res2.t18 121.245
R7520 bgr_0.cap_res2.t13 bgr_0.cap_res2.t7 0.1603
R7521 bgr_0.cap_res2.t6 bgr_0.cap_res2.t1 0.1603
R7522 bgr_0.cap_res2.t11 bgr_0.cap_res2.t5 0.1603
R7523 bgr_0.cap_res2.t4 bgr_0.cap_res2.t20 0.1603
R7524 bgr_0.cap_res2.t19 bgr_0.cap_res2.t16 0.1603
R7525 bgr_0.cap_res2.n1 bgr_0.cap_res2.t3 0.159278
R7526 bgr_0.cap_res2.n2 bgr_0.cap_res2.t10 0.159278
R7527 bgr_0.cap_res2.n3 bgr_0.cap_res2.t17 0.159278
R7528 bgr_0.cap_res2.n4 bgr_0.cap_res2.t12 0.159278
R7529 bgr_0.cap_res2.n4 bgr_0.cap_res2.t15 0.1368
R7530 bgr_0.cap_res2.n4 bgr_0.cap_res2.t13 0.1368
R7531 bgr_0.cap_res2.n3 bgr_0.cap_res2.t9 0.1368
R7532 bgr_0.cap_res2.n3 bgr_0.cap_res2.t6 0.1368
R7533 bgr_0.cap_res2.n2 bgr_0.cap_res2.t14 0.1368
R7534 bgr_0.cap_res2.n2 bgr_0.cap_res2.t11 0.1368
R7535 bgr_0.cap_res2.n1 bgr_0.cap_res2.t8 0.1368
R7536 bgr_0.cap_res2.n1 bgr_0.cap_res2.t4 0.1368
R7537 bgr_0.cap_res2.n0 bgr_0.cap_res2.t2 0.1368
R7538 bgr_0.cap_res2.n0 bgr_0.cap_res2.t19 0.1368
R7539 bgr_0.cap_res2.t3 bgr_0.cap_res2.n0 0.00152174
R7540 bgr_0.cap_res2.t10 bgr_0.cap_res2.n1 0.00152174
R7541 bgr_0.cap_res2.t17 bgr_0.cap_res2.n2 0.00152174
R7542 bgr_0.cap_res2.t12 bgr_0.cap_res2.n3 0.00152174
R7543 bgr_0.cap_res2.t18 bgr_0.cap_res2.n4 0.00152174
R7544 two_stage_opamp_dummy_magic_16_0.Vb2.n25 two_stage_opamp_dummy_magic_16_0.Vb2.t31 650.273
R7545 two_stage_opamp_dummy_magic_16_0.Vb2.n27 two_stage_opamp_dummy_magic_16_0.Vb2.t9 650.273
R7546 two_stage_opamp_dummy_magic_16_0.Vb2.n4 two_stage_opamp_dummy_magic_16_0.Vb2.t12 611.739
R7547 two_stage_opamp_dummy_magic_16_0.Vb2.n0 two_stage_opamp_dummy_magic_16_0.Vb2.t22 611.739
R7548 two_stage_opamp_dummy_magic_16_0.Vb2.n13 two_stage_opamp_dummy_magic_16_0.Vb2.t13 611.739
R7549 two_stage_opamp_dummy_magic_16_0.Vb2.n9 two_stage_opamp_dummy_magic_16_0.Vb2.t23 611.739
R7550 two_stage_opamp_dummy_magic_16_0.Vb2.n28 two_stage_opamp_dummy_magic_16_0.Vb2.t27 445.423
R7551 two_stage_opamp_dummy_magic_16_0.Vb2.n4 two_stage_opamp_dummy_magic_16_0.Vb2.t17 421.75
R7552 two_stage_opamp_dummy_magic_16_0.Vb2.n5 two_stage_opamp_dummy_magic_16_0.Vb2.t24 421.75
R7553 two_stage_opamp_dummy_magic_16_0.Vb2.n6 two_stage_opamp_dummy_magic_16_0.Vb2.t28 421.75
R7554 two_stage_opamp_dummy_magic_16_0.Vb2.n7 two_stage_opamp_dummy_magic_16_0.Vb2.t29 421.75
R7555 two_stage_opamp_dummy_magic_16_0.Vb2.n0 two_stage_opamp_dummy_magic_16_0.Vb2.t26 421.75
R7556 two_stage_opamp_dummy_magic_16_0.Vb2.n1 two_stage_opamp_dummy_magic_16_0.Vb2.t19 421.75
R7557 two_stage_opamp_dummy_magic_16_0.Vb2.n2 two_stage_opamp_dummy_magic_16_0.Vb2.t14 421.75
R7558 two_stage_opamp_dummy_magic_16_0.Vb2.n3 two_stage_opamp_dummy_magic_16_0.Vb2.t32 421.75
R7559 two_stage_opamp_dummy_magic_16_0.Vb2.n13 two_stage_opamp_dummy_magic_16_0.Vb2.t18 421.75
R7560 two_stage_opamp_dummy_magic_16_0.Vb2.n14 two_stage_opamp_dummy_magic_16_0.Vb2.t25 421.75
R7561 two_stage_opamp_dummy_magic_16_0.Vb2.n15 two_stage_opamp_dummy_magic_16_0.Vb2.t21 421.75
R7562 two_stage_opamp_dummy_magic_16_0.Vb2.n16 two_stage_opamp_dummy_magic_16_0.Vb2.t30 421.75
R7563 two_stage_opamp_dummy_magic_16_0.Vb2.n9 two_stage_opamp_dummy_magic_16_0.Vb2.t16 421.75
R7564 two_stage_opamp_dummy_magic_16_0.Vb2.n10 two_stage_opamp_dummy_magic_16_0.Vb2.t20 421.75
R7565 two_stage_opamp_dummy_magic_16_0.Vb2.n11 two_stage_opamp_dummy_magic_16_0.Vb2.t15 421.75
R7566 two_stage_opamp_dummy_magic_16_0.Vb2.n12 two_stage_opamp_dummy_magic_16_0.Vb2.t11 421.75
R7567 two_stage_opamp_dummy_magic_16_0.Vb2.n30 two_stage_opamp_dummy_magic_16_0.Vb2.n17 169.352
R7568 two_stage_opamp_dummy_magic_16_0.Vb2.n5 two_stage_opamp_dummy_magic_16_0.Vb2.n4 167.094
R7569 two_stage_opamp_dummy_magic_16_0.Vb2.n6 two_stage_opamp_dummy_magic_16_0.Vb2.n5 167.094
R7570 two_stage_opamp_dummy_magic_16_0.Vb2.n7 two_stage_opamp_dummy_magic_16_0.Vb2.n6 167.094
R7571 two_stage_opamp_dummy_magic_16_0.Vb2.n1 two_stage_opamp_dummy_magic_16_0.Vb2.n0 167.094
R7572 two_stage_opamp_dummy_magic_16_0.Vb2.n2 two_stage_opamp_dummy_magic_16_0.Vb2.n1 167.094
R7573 two_stage_opamp_dummy_magic_16_0.Vb2.n3 two_stage_opamp_dummy_magic_16_0.Vb2.n2 167.094
R7574 two_stage_opamp_dummy_magic_16_0.Vb2.n14 two_stage_opamp_dummy_magic_16_0.Vb2.n13 167.094
R7575 two_stage_opamp_dummy_magic_16_0.Vb2.n15 two_stage_opamp_dummy_magic_16_0.Vb2.n14 167.094
R7576 two_stage_opamp_dummy_magic_16_0.Vb2.n16 two_stage_opamp_dummy_magic_16_0.Vb2.n15 167.094
R7577 two_stage_opamp_dummy_magic_16_0.Vb2.n10 two_stage_opamp_dummy_magic_16_0.Vb2.n9 167.094
R7578 two_stage_opamp_dummy_magic_16_0.Vb2.n11 two_stage_opamp_dummy_magic_16_0.Vb2.n10 167.094
R7579 two_stage_opamp_dummy_magic_16_0.Vb2.n12 two_stage_opamp_dummy_magic_16_0.Vb2.n11 167.094
R7580 two_stage_opamp_dummy_magic_16_0.Vb2 two_stage_opamp_dummy_magic_16_0.Vb2.n8 161.477
R7581 two_stage_opamp_dummy_magic_16_0.Vb2.n27 two_stage_opamp_dummy_magic_16_0.Vb2.n26 160.06
R7582 two_stage_opamp_dummy_magic_16_0.Vb2.n20 two_stage_opamp_dummy_magic_16_0.Vb2.n18 140.857
R7583 two_stage_opamp_dummy_magic_16_0.Vb2.n22 two_stage_opamp_dummy_magic_16_0.Vb2.n21 139.608
R7584 two_stage_opamp_dummy_magic_16_0.Vb2.n24 two_stage_opamp_dummy_magic_16_0.Vb2.n23 139.608
R7585 two_stage_opamp_dummy_magic_16_0.Vb2.n20 two_stage_opamp_dummy_magic_16_0.Vb2.n19 139.608
R7586 two_stage_opamp_dummy_magic_16_0.Vb2.n25 two_stage_opamp_dummy_magic_16_0.Vb2.n24 61.3349
R7587 two_stage_opamp_dummy_magic_16_0.Vb2.n8 two_stage_opamp_dummy_magic_16_0.Vb2.n7 49.8072
R7588 two_stage_opamp_dummy_magic_16_0.Vb2.n8 two_stage_opamp_dummy_magic_16_0.Vb2.n3 49.8072
R7589 two_stage_opamp_dummy_magic_16_0.Vb2.n17 two_stage_opamp_dummy_magic_16_0.Vb2.n16 49.8072
R7590 two_stage_opamp_dummy_magic_16_0.Vb2.n17 two_stage_opamp_dummy_magic_16_0.Vb2.n12 49.8072
R7591 two_stage_opamp_dummy_magic_16_0.Vb2.n18 two_stage_opamp_dummy_magic_16_0.Vb2.t4 24.0005
R7592 two_stage_opamp_dummy_magic_16_0.Vb2.n18 two_stage_opamp_dummy_magic_16_0.Vb2.t6 24.0005
R7593 two_stage_opamp_dummy_magic_16_0.Vb2.n21 two_stage_opamp_dummy_magic_16_0.Vb2.t2 24.0005
R7594 two_stage_opamp_dummy_magic_16_0.Vb2.n21 two_stage_opamp_dummy_magic_16_0.Vb2.t0 24.0005
R7595 two_stage_opamp_dummy_magic_16_0.Vb2.n23 two_stage_opamp_dummy_magic_16_0.Vb2.t7 24.0005
R7596 two_stage_opamp_dummy_magic_16_0.Vb2.n23 two_stage_opamp_dummy_magic_16_0.Vb2.t1 24.0005
R7597 two_stage_opamp_dummy_magic_16_0.Vb2.n19 two_stage_opamp_dummy_magic_16_0.Vb2.t3 24.0005
R7598 two_stage_opamp_dummy_magic_16_0.Vb2.n19 two_stage_opamp_dummy_magic_16_0.Vb2.t5 24.0005
R7599 two_stage_opamp_dummy_magic_16_0.Vb2.n30 two_stage_opamp_dummy_magic_16_0.Vb2.n29 12.8443
R7600 two_stage_opamp_dummy_magic_16_0.Vb2.n26 two_stage_opamp_dummy_magic_16_0.Vb2.t10 11.2576
R7601 two_stage_opamp_dummy_magic_16_0.Vb2.n26 two_stage_opamp_dummy_magic_16_0.Vb2.t8 11.2576
R7602 two_stage_opamp_dummy_magic_16_0.Vb2.n22 two_stage_opamp_dummy_magic_16_0.Vb2.n20 7.563
R7603 two_stage_opamp_dummy_magic_16_0.Vb2 two_stage_opamp_dummy_magic_16_0.Vb2.n30 7.2505
R7604 two_stage_opamp_dummy_magic_16_0.Vb2.n29 two_stage_opamp_dummy_magic_16_0.Vb2.n25 4.54113
R7605 two_stage_opamp_dummy_magic_16_0.Vb2.n28 two_stage_opamp_dummy_magic_16_0.Vb2.n27 2.84425
R7606 two_stage_opamp_dummy_magic_16_0.Vb2.n24 two_stage_opamp_dummy_magic_16_0.Vb2.n22 1.2505
R7607 two_stage_opamp_dummy_magic_16_0.Vb2.n29 two_stage_opamp_dummy_magic_16_0.Vb2.n28 0.928625
R7608 two_stage_opamp_dummy_magic_16_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_16_0.err_amp_mir.t5 554.301
R7609 two_stage_opamp_dummy_magic_16_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_16_0.err_amp_mir.t0 442.837
R7610 two_stage_opamp_dummy_magic_16_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_16_0.err_amp_mir.n0 183.978
R7611 two_stage_opamp_dummy_magic_16_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_16_0.err_amp_mir.n1 173.088
R7612 two_stage_opamp_dummy_magic_16_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_16_0.err_amp_mir.n2 86.8857
R7613 two_stage_opamp_dummy_magic_16_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_16_0.err_amp_mir.t4 15.7605
R7614 two_stage_opamp_dummy_magic_16_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_16_0.err_amp_mir.t3 15.7605
R7615 two_stage_opamp_dummy_magic_16_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_16_0.err_amp_mir.t2 9.6005
R7616 two_stage_opamp_dummy_magic_16_0.err_amp_mir.t1 two_stage_opamp_dummy_magic_16_0.err_amp_mir.n3 9.6005
R7617 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.n3 526.183
R7618 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.n1 514.134
R7619 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n0 360.586
R7620 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t5 303.259
R7621 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n4 210.169
R7622 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t3 174.726
R7623 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.t7 174.726
R7624 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.t4 174.726
R7625 bgr_0.V_CUR_REF_REG.t1 bgr_0.V_CUR_REF_REG.n5 153.474
R7626 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.n2 128.534
R7627 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t6 96.4005
R7628 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t0 39.4005
R7629 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t2 39.4005
R7630 bgr_0.V_p_2.n1 bgr_0.V_p_2.n2 229.562
R7631 bgr_0.V_p_2.n1 bgr_0.V_p_2.n5 228.939
R7632 bgr_0.V_p_2.n0 bgr_0.V_p_2.n4 228.939
R7633 bgr_0.V_p_2.n0 bgr_0.V_p_2.n3 228.939
R7634 bgr_0.V_p_2.n6 bgr_0.V_p_2.n1 228.938
R7635 bgr_0.V_p_2.n0 bgr_0.V_p_2.t10 98.7279
R7636 bgr_0.V_p_2.n5 bgr_0.V_p_2.t4 48.0005
R7637 bgr_0.V_p_2.n5 bgr_0.V_p_2.t5 48.0005
R7638 bgr_0.V_p_2.n4 bgr_0.V_p_2.t8 48.0005
R7639 bgr_0.V_p_2.n4 bgr_0.V_p_2.t3 48.0005
R7640 bgr_0.V_p_2.n3 bgr_0.V_p_2.t1 48.0005
R7641 bgr_0.V_p_2.n3 bgr_0.V_p_2.t6 48.0005
R7642 bgr_0.V_p_2.n2 bgr_0.V_p_2.t0 48.0005
R7643 bgr_0.V_p_2.n2 bgr_0.V_p_2.t7 48.0005
R7644 bgr_0.V_p_2.t9 bgr_0.V_p_2.n6 48.0005
R7645 bgr_0.V_p_2.n6 bgr_0.V_p_2.t2 48.0005
R7646 bgr_0.V_p_2.n1 bgr_0.V_p_2.n0 1.8755
R7647 a_7460_23988.t0 a_7460_23988.t1 178.133
R7648 two_stage_opamp_dummy_magic_16_0.Vb1.n26 two_stage_opamp_dummy_magic_16_0.Vb1.t24 449.868
R7649 two_stage_opamp_dummy_magic_16_0.Vb1.n22 two_stage_opamp_dummy_magic_16_0.Vb1.t28 449.868
R7650 two_stage_opamp_dummy_magic_16_0.Vb1.n17 two_stage_opamp_dummy_magic_16_0.Vb1.t23 449.868
R7651 two_stage_opamp_dummy_magic_16_0.Vb1.n13 two_stage_opamp_dummy_magic_16_0.Vb1.t27 449.868
R7652 two_stage_opamp_dummy_magic_16_0.Vb1.n6 two_stage_opamp_dummy_magic_16_0.Vb1.t1 449.868
R7653 two_stage_opamp_dummy_magic_16_0.Vb1.n5 two_stage_opamp_dummy_magic_16_0.Vb1.t5 449.868
R7654 two_stage_opamp_dummy_magic_16_0.Vb1.n2 two_stage_opamp_dummy_magic_16_0.Vb1.n0 339.961
R7655 two_stage_opamp_dummy_magic_16_0.Vb1.n2 two_stage_opamp_dummy_magic_16_0.Vb1.n1 339.272
R7656 two_stage_opamp_dummy_magic_16_0.Vb1.n26 two_stage_opamp_dummy_magic_16_0.Vb1.t33 273.134
R7657 two_stage_opamp_dummy_magic_16_0.Vb1.n27 two_stage_opamp_dummy_magic_16_0.Vb1.t22 273.134
R7658 two_stage_opamp_dummy_magic_16_0.Vb1.n28 two_stage_opamp_dummy_magic_16_0.Vb1.t31 273.134
R7659 two_stage_opamp_dummy_magic_16_0.Vb1.n29 two_stage_opamp_dummy_magic_16_0.Vb1.t19 273.134
R7660 two_stage_opamp_dummy_magic_16_0.Vb1.n25 two_stage_opamp_dummy_magic_16_0.Vb1.t15 273.134
R7661 two_stage_opamp_dummy_magic_16_0.Vb1.n24 two_stage_opamp_dummy_magic_16_0.Vb1.t20 273.134
R7662 two_stage_opamp_dummy_magic_16_0.Vb1.n23 two_stage_opamp_dummy_magic_16_0.Vb1.t29 273.134
R7663 two_stage_opamp_dummy_magic_16_0.Vb1.n22 two_stage_opamp_dummy_magic_16_0.Vb1.t18 273.134
R7664 two_stage_opamp_dummy_magic_16_0.Vb1.n17 two_stage_opamp_dummy_magic_16_0.Vb1.t32 273.134
R7665 two_stage_opamp_dummy_magic_16_0.Vb1.n18 two_stage_opamp_dummy_magic_16_0.Vb1.t21 273.134
R7666 two_stage_opamp_dummy_magic_16_0.Vb1.n19 two_stage_opamp_dummy_magic_16_0.Vb1.t30 273.134
R7667 two_stage_opamp_dummy_magic_16_0.Vb1.n20 two_stage_opamp_dummy_magic_16_0.Vb1.t26 273.134
R7668 two_stage_opamp_dummy_magic_16_0.Vb1.n16 two_stage_opamp_dummy_magic_16_0.Vb1.t14 273.134
R7669 two_stage_opamp_dummy_magic_16_0.Vb1.n15 two_stage_opamp_dummy_magic_16_0.Vb1.t25 273.134
R7670 two_stage_opamp_dummy_magic_16_0.Vb1.n14 two_stage_opamp_dummy_magic_16_0.Vb1.t34 273.134
R7671 two_stage_opamp_dummy_magic_16_0.Vb1.n13 two_stage_opamp_dummy_magic_16_0.Vb1.t17 273.134
R7672 two_stage_opamp_dummy_magic_16_0.Vb1.n6 two_stage_opamp_dummy_magic_16_0.Vb1.t7 273.134
R7673 two_stage_opamp_dummy_magic_16_0.Vb1.n5 two_stage_opamp_dummy_magic_16_0.Vb1.t3 273.134
R7674 two_stage_opamp_dummy_magic_16_0.Vb1.n29 two_stage_opamp_dummy_magic_16_0.Vb1.n28 176.733
R7675 two_stage_opamp_dummy_magic_16_0.Vb1.n28 two_stage_opamp_dummy_magic_16_0.Vb1.n27 176.733
R7676 two_stage_opamp_dummy_magic_16_0.Vb1.n27 two_stage_opamp_dummy_magic_16_0.Vb1.n26 176.733
R7677 two_stage_opamp_dummy_magic_16_0.Vb1.n23 two_stage_opamp_dummy_magic_16_0.Vb1.n22 176.733
R7678 two_stage_opamp_dummy_magic_16_0.Vb1.n24 two_stage_opamp_dummy_magic_16_0.Vb1.n23 176.733
R7679 two_stage_opamp_dummy_magic_16_0.Vb1.n25 two_stage_opamp_dummy_magic_16_0.Vb1.n24 176.733
R7680 two_stage_opamp_dummy_magic_16_0.Vb1.n20 two_stage_opamp_dummy_magic_16_0.Vb1.n19 176.733
R7681 two_stage_opamp_dummy_magic_16_0.Vb1.n19 two_stage_opamp_dummy_magic_16_0.Vb1.n18 176.733
R7682 two_stage_opamp_dummy_magic_16_0.Vb1.n18 two_stage_opamp_dummy_magic_16_0.Vb1.n17 176.733
R7683 two_stage_opamp_dummy_magic_16_0.Vb1.n14 two_stage_opamp_dummy_magic_16_0.Vb1.n13 176.733
R7684 two_stage_opamp_dummy_magic_16_0.Vb1.n15 two_stage_opamp_dummy_magic_16_0.Vb1.n14 176.733
R7685 two_stage_opamp_dummy_magic_16_0.Vb1.n16 two_stage_opamp_dummy_magic_16_0.Vb1.n15 176.733
R7686 two_stage_opamp_dummy_magic_16_0.Vb1.n31 two_stage_opamp_dummy_magic_16_0.Vb1.n21 172.207
R7687 two_stage_opamp_dummy_magic_16_0.Vb1.n31 two_stage_opamp_dummy_magic_16_0.Vb1.n30 165.8
R7688 two_stage_opamp_dummy_magic_16_0.Vb1.n9 two_stage_opamp_dummy_magic_16_0.Vb1.n7 152
R7689 two_stage_opamp_dummy_magic_16_0.Vb1.n4 two_stage_opamp_dummy_magic_16_0.Vb1.n3 113.906
R7690 two_stage_opamp_dummy_magic_16_0.Vb1.n12 two_stage_opamp_dummy_magic_16_0.Vb1.n11 113.906
R7691 two_stage_opamp_dummy_magic_16_0.Vb1.n9 two_stage_opamp_dummy_magic_16_0.Vb1.n8 100.106
R7692 two_stage_opamp_dummy_magic_16_0.Vb1.n4 two_stage_opamp_dummy_magic_16_0.Vb1.t16 65.0512
R7693 two_stage_opamp_dummy_magic_16_0.Vb1.n30 two_stage_opamp_dummy_magic_16_0.Vb1.n29 54.6272
R7694 two_stage_opamp_dummy_magic_16_0.Vb1.n30 two_stage_opamp_dummy_magic_16_0.Vb1.n25 54.6272
R7695 two_stage_opamp_dummy_magic_16_0.Vb1.n21 two_stage_opamp_dummy_magic_16_0.Vb1.n20 54.6272
R7696 two_stage_opamp_dummy_magic_16_0.Vb1.n21 two_stage_opamp_dummy_magic_16_0.Vb1.n16 54.6272
R7697 two_stage_opamp_dummy_magic_16_0.Vb1.n7 two_stage_opamp_dummy_magic_16_0.Vb1.n6 45.5227
R7698 two_stage_opamp_dummy_magic_16_0.Vb1.n7 two_stage_opamp_dummy_magic_16_0.Vb1.n5 45.5227
R7699 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_16_0.Vb1.n32 44.063
R7700 two_stage_opamp_dummy_magic_16_0.Vb1.n1 two_stage_opamp_dummy_magic_16_0.Vb1.t9 39.4005
R7701 two_stage_opamp_dummy_magic_16_0.Vb1.n1 two_stage_opamp_dummy_magic_16_0.Vb1.t12 39.4005
R7702 two_stage_opamp_dummy_magic_16_0.Vb1.n0 two_stage_opamp_dummy_magic_16_0.Vb1.t13 39.4005
R7703 two_stage_opamp_dummy_magic_16_0.Vb1.n0 two_stage_opamp_dummy_magic_16_0.Vb1.t0 39.4005
R7704 two_stage_opamp_dummy_magic_16_0.Vb1.n32 two_stage_opamp_dummy_magic_16_0.Vb1.n12 17.063
R7705 two_stage_opamp_dummy_magic_16_0.Vb1.n8 two_stage_opamp_dummy_magic_16_0.Vb1.t4 16.0005
R7706 two_stage_opamp_dummy_magic_16_0.Vb1.n8 two_stage_opamp_dummy_magic_16_0.Vb1.t8 16.0005
R7707 two_stage_opamp_dummy_magic_16_0.Vb1.n3 two_stage_opamp_dummy_magic_16_0.Vb1.t10 16.0005
R7708 two_stage_opamp_dummy_magic_16_0.Vb1.n3 two_stage_opamp_dummy_magic_16_0.Vb1.t6 16.0005
R7709 two_stage_opamp_dummy_magic_16_0.Vb1.n11 two_stage_opamp_dummy_magic_16_0.Vb1.t2 16.0005
R7710 two_stage_opamp_dummy_magic_16_0.Vb1.n11 two_stage_opamp_dummy_magic_16_0.Vb1.t11 16.0005
R7711 two_stage_opamp_dummy_magic_16_0.Vb1.n10 two_stage_opamp_dummy_magic_16_0.Vb1.n9 13.8005
R7712 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_16_0.Vb1.n2 12.1255
R7713 two_stage_opamp_dummy_magic_16_0.Vb1.n32 two_stage_opamp_dummy_magic_16_0.Vb1.n31 6.92238
R7714 two_stage_opamp_dummy_magic_16_0.Vb1.n10 two_stage_opamp_dummy_magic_16_0.Vb1.n4 0.563
R7715 two_stage_opamp_dummy_magic_16_0.Vb1.n12 two_stage_opamp_dummy_magic_16_0.Vb1.n10 0.563
R7716 two_stage_opamp_dummy_magic_16_0.VD1.n3 two_stage_opamp_dummy_magic_16_0.VD1.n1 118.061
R7717 two_stage_opamp_dummy_magic_16_0.VD1.n17 two_stage_opamp_dummy_magic_16_0.VD1.n16 116.811
R7718 two_stage_opamp_dummy_magic_16_0.VD1.n19 two_stage_opamp_dummy_magic_16_0.VD1.n18 116.811
R7719 two_stage_opamp_dummy_magic_16_0.VD1.n3 two_stage_opamp_dummy_magic_16_0.VD1.n2 116.811
R7720 two_stage_opamp_dummy_magic_16_0.VD1.n11 two_stage_opamp_dummy_magic_16_0.VD1.n10 114.719
R7721 two_stage_opamp_dummy_magic_16_0.VD1.n7 two_stage_opamp_dummy_magic_16_0.VD1.n5 114.719
R7722 two_stage_opamp_dummy_magic_16_0.VD1.n7 two_stage_opamp_dummy_magic_16_0.VD1.n6 114.156
R7723 two_stage_opamp_dummy_magic_16_0.VD1.n9 two_stage_opamp_dummy_magic_16_0.VD1.n8 114.156
R7724 two_stage_opamp_dummy_magic_16_0.VD1.n14 two_stage_opamp_dummy_magic_16_0.VD1.n13 112.29
R7725 two_stage_opamp_dummy_magic_16_0.VD1 two_stage_opamp_dummy_magic_16_0.VD1.n0 112.249
R7726 two_stage_opamp_dummy_magic_16_0.VD1.n12 two_stage_opamp_dummy_magic_16_0.VD1.n4 109.639
R7727 two_stage_opamp_dummy_magic_16_0.VD1.n4 two_stage_opamp_dummy_magic_16_0.VD1.t4 16.0005
R7728 two_stage_opamp_dummy_magic_16_0.VD1.n4 two_stage_opamp_dummy_magic_16_0.VD1.t9 16.0005
R7729 two_stage_opamp_dummy_magic_16_0.VD1.n16 two_stage_opamp_dummy_magic_16_0.VD1.t16 16.0005
R7730 two_stage_opamp_dummy_magic_16_0.VD1.n16 two_stage_opamp_dummy_magic_16_0.VD1.t13 16.0005
R7731 two_stage_opamp_dummy_magic_16_0.VD1.n18 two_stage_opamp_dummy_magic_16_0.VD1.t14 16.0005
R7732 two_stage_opamp_dummy_magic_16_0.VD1.n18 two_stage_opamp_dummy_magic_16_0.VD1.t18 16.0005
R7733 two_stage_opamp_dummy_magic_16_0.VD1.n0 two_stage_opamp_dummy_magic_16_0.VD1.t21 16.0005
R7734 two_stage_opamp_dummy_magic_16_0.VD1.n0 two_stage_opamp_dummy_magic_16_0.VD1.t19 16.0005
R7735 two_stage_opamp_dummy_magic_16_0.VD1.n2 two_stage_opamp_dummy_magic_16_0.VD1.t1 16.0005
R7736 two_stage_opamp_dummy_magic_16_0.VD1.n2 two_stage_opamp_dummy_magic_16_0.VD1.t20 16.0005
R7737 two_stage_opamp_dummy_magic_16_0.VD1.n1 two_stage_opamp_dummy_magic_16_0.VD1.t17 16.0005
R7738 two_stage_opamp_dummy_magic_16_0.VD1.n1 two_stage_opamp_dummy_magic_16_0.VD1.t15 16.0005
R7739 two_stage_opamp_dummy_magic_16_0.VD1.n13 two_stage_opamp_dummy_magic_16_0.VD1.t0 16.0005
R7740 two_stage_opamp_dummy_magic_16_0.VD1.n13 two_stage_opamp_dummy_magic_16_0.VD1.t12 16.0005
R7741 two_stage_opamp_dummy_magic_16_0.VD1.n10 two_stage_opamp_dummy_magic_16_0.VD1.t3 16.0005
R7742 two_stage_opamp_dummy_magic_16_0.VD1.n10 two_stage_opamp_dummy_magic_16_0.VD1.t8 16.0005
R7743 two_stage_opamp_dummy_magic_16_0.VD1.n6 two_stage_opamp_dummy_magic_16_0.VD1.t2 16.0005
R7744 two_stage_opamp_dummy_magic_16_0.VD1.n6 two_stage_opamp_dummy_magic_16_0.VD1.t7 16.0005
R7745 two_stage_opamp_dummy_magic_16_0.VD1.n5 two_stage_opamp_dummy_magic_16_0.VD1.t5 16.0005
R7746 two_stage_opamp_dummy_magic_16_0.VD1.n5 two_stage_opamp_dummy_magic_16_0.VD1.t10 16.0005
R7747 two_stage_opamp_dummy_magic_16_0.VD1.n8 two_stage_opamp_dummy_magic_16_0.VD1.t11 16.0005
R7748 two_stage_opamp_dummy_magic_16_0.VD1.n8 two_stage_opamp_dummy_magic_16_0.VD1.t6 16.0005
R7749 two_stage_opamp_dummy_magic_16_0.VD1 two_stage_opamp_dummy_magic_16_0.VD1.n19 5.76612
R7750 two_stage_opamp_dummy_magic_16_0.VD1.n15 two_stage_opamp_dummy_magic_16_0.VD1.n14 4.5005
R7751 two_stage_opamp_dummy_magic_16_0.VD1.n12 two_stage_opamp_dummy_magic_16_0.VD1.n11 4.5005
R7752 two_stage_opamp_dummy_magic_16_0.VD1.n17 two_stage_opamp_dummy_magic_16_0.VD1.n15 3.6255
R7753 two_stage_opamp_dummy_magic_16_0.VD1.n19 two_stage_opamp_dummy_magic_16_0.VD1.n17 1.2505
R7754 two_stage_opamp_dummy_magic_16_0.VD1.n15 two_stage_opamp_dummy_magic_16_0.VD1.n3 1.2505
R7755 two_stage_opamp_dummy_magic_16_0.VD1.n11 two_stage_opamp_dummy_magic_16_0.VD1.n9 0.563
R7756 two_stage_opamp_dummy_magic_16_0.VD1.n9 two_stage_opamp_dummy_magic_16_0.VD1.n7 0.563
R7757 two_stage_opamp_dummy_magic_16_0.VD1.n14 two_stage_opamp_dummy_magic_16_0.VD1.n12 0.118871
R7758 a_6930_22564.t0 a_6930_22564.t1 178.133
R7759 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t13 369.534
R7760 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t12 369.534
R7761 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t29 369.534
R7762 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t17 369.534
R7763 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t21 369.534
R7764 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t20 369.534
R7765 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n6 341.397
R7766 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n9 339.272
R7767 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n7 339.272
R7768 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n12 334.772
R7769 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.t14 238.322
R7770 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.t27 238.322
R7771 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t26 192.8
R7772 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t19 192.8
R7773 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.t16 192.8
R7774 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.t23 192.8
R7775 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t22 192.8
R7776 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t24 192.8
R7777 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.t10 192.8
R7778 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.t18 192.8
R7779 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.t25 192.8
R7780 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.t11 192.8
R7781 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t15 192.8
R7782 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t28 192.8
R7783 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.n24 176.733
R7784 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.n23 176.733
R7785 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.n18 176.733
R7786 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.n19 176.733
R7787 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.n20 176.733
R7788 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.n21 176.733
R7789 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n2 171.321
R7790 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n5 168.166
R7791 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.n14 167.519
R7792 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n26 166.071
R7793 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.t0 137.48
R7794 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.t7 100.635
R7795 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n4 56.2338
R7796 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n3 56.2338
R7797 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n25 56.2338
R7798 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n22 56.2338
R7799 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n1 56.2338
R7800 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n0 56.2338
R7801 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t9 39.4005
R7802 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t2 39.4005
R7803 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t4 39.4005
R7804 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t6 39.4005
R7805 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t3 39.4005
R7806 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t5 39.4005
R7807 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t1 39.4005
R7808 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t8 39.4005
R7809 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n16 27.5005
R7810 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n13 9.53175
R7811 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n11 4.5005
R7812 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n17 2.34425
R7813 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n8 2.1255
R7814 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.n10 2.1255
R7815 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n15 1.688
R7816 VIN+.n9 VIN+.t5 487.051
R7817 VIN+.n4 VIN+.t3 487.051
R7818 VIN+.n3 VIN+.t4 487.051
R7819 VIN+.n7 VIN+.t9 318.656
R7820 VIN+.n7 VIN+.t2 318.656
R7821 VIN+.n5 VIN+.t7 318.656
R7822 VIN+.n5 VIN+.t1 318.656
R7823 VIN+.n1 VIN+.t8 318.656
R7824 VIN+.n1 VIN+.t6 318.656
R7825 VIN+.n0 VIN+.t10 318.656
R7826 VIN+.n0 VIN+.t0 318.656
R7827 VIN+.n2 VIN+.n0 167.05
R7828 VIN+.n8 VIN+.n7 165.8
R7829 VIN+.n6 VIN+.n5 165.8
R7830 VIN+.n2 VIN+.n1 165.8
R7831 VIN+.n6 VIN+.n4 2.35363
R7832 VIN+.n4 VIN+.n3 1.29425
R7833 VIN+.n8 VIN+.n6 1.2505
R7834 VIN+.n3 VIN+.n2 1.16612
R7835 VIN+.n9 VIN+.n8 1.16612
R7836 VIN+ VIN+.n9 0.616125
R7837 two_stage_opamp_dummy_magic_16_0.VD2.n2 two_stage_opamp_dummy_magic_16_0.VD2.n0 117.561
R7838 two_stage_opamp_dummy_magic_16_0.VD2.n19 two_stage_opamp_dummy_magic_16_0.VD2.n18 117.561
R7839 two_stage_opamp_dummy_magic_16_0.VD2.n18 two_stage_opamp_dummy_magic_16_0.VD2.n17 116.311
R7840 two_stage_opamp_dummy_magic_16_0.VD2.n16 two_stage_opamp_dummy_magic_16_0.VD2.n15 116.311
R7841 two_stage_opamp_dummy_magic_16_0.VD2.n2 two_stage_opamp_dummy_magic_16_0.VD2.n1 116.311
R7842 two_stage_opamp_dummy_magic_16_0.VD2.n7 two_stage_opamp_dummy_magic_16_0.VD2.n5 114.719
R7843 two_stage_opamp_dummy_magic_16_0.VD2.n10 two_stage_opamp_dummy_magic_16_0.VD2.n4 114.719
R7844 two_stage_opamp_dummy_magic_16_0.VD2.n9 two_stage_opamp_dummy_magic_16_0.VD2.n8 114.156
R7845 two_stage_opamp_dummy_magic_16_0.VD2.n7 two_stage_opamp_dummy_magic_16_0.VD2.n6 114.156
R7846 two_stage_opamp_dummy_magic_16_0.VD2.n13 two_stage_opamp_dummy_magic_16_0.VD2.n12 111.794
R7847 two_stage_opamp_dummy_magic_16_0.VD2.n11 two_stage_opamp_dummy_magic_16_0.VD2.n3 109.635
R7848 two_stage_opamp_dummy_magic_16_0.VD2.n17 two_stage_opamp_dummy_magic_16_0.VD2.t14 16.0005
R7849 two_stage_opamp_dummy_magic_16_0.VD2.n17 two_stage_opamp_dummy_magic_16_0.VD2.t12 16.0005
R7850 two_stage_opamp_dummy_magic_16_0.VD2.n15 two_stage_opamp_dummy_magic_16_0.VD2.t16 16.0005
R7851 two_stage_opamp_dummy_magic_16_0.VD2.n15 two_stage_opamp_dummy_magic_16_0.VD2.t21 16.0005
R7852 two_stage_opamp_dummy_magic_16_0.VD2.n8 two_stage_opamp_dummy_magic_16_0.VD2.t0 16.0005
R7853 two_stage_opamp_dummy_magic_16_0.VD2.n8 two_stage_opamp_dummy_magic_16_0.VD2.t8 16.0005
R7854 two_stage_opamp_dummy_magic_16_0.VD2.n6 two_stage_opamp_dummy_magic_16_0.VD2.t3 16.0005
R7855 two_stage_opamp_dummy_magic_16_0.VD2.n6 two_stage_opamp_dummy_magic_16_0.VD2.t2 16.0005
R7856 two_stage_opamp_dummy_magic_16_0.VD2.n5 two_stage_opamp_dummy_magic_16_0.VD2.t7 16.0005
R7857 two_stage_opamp_dummy_magic_16_0.VD2.n5 two_stage_opamp_dummy_magic_16_0.VD2.t4 16.0005
R7858 two_stage_opamp_dummy_magic_16_0.VD2.n4 two_stage_opamp_dummy_magic_16_0.VD2.t6 16.0005
R7859 two_stage_opamp_dummy_magic_16_0.VD2.n4 two_stage_opamp_dummy_magic_16_0.VD2.t1 16.0005
R7860 two_stage_opamp_dummy_magic_16_0.VD2.n3 two_stage_opamp_dummy_magic_16_0.VD2.t9 16.0005
R7861 two_stage_opamp_dummy_magic_16_0.VD2.n3 two_stage_opamp_dummy_magic_16_0.VD2.t5 16.0005
R7862 two_stage_opamp_dummy_magic_16_0.VD2.n12 two_stage_opamp_dummy_magic_16_0.VD2.t18 16.0005
R7863 two_stage_opamp_dummy_magic_16_0.VD2.n12 two_stage_opamp_dummy_magic_16_0.VD2.t13 16.0005
R7864 two_stage_opamp_dummy_magic_16_0.VD2.n1 two_stage_opamp_dummy_magic_16_0.VD2.t17 16.0005
R7865 two_stage_opamp_dummy_magic_16_0.VD2.n1 two_stage_opamp_dummy_magic_16_0.VD2.t11 16.0005
R7866 two_stage_opamp_dummy_magic_16_0.VD2.n0 two_stage_opamp_dummy_magic_16_0.VD2.t15 16.0005
R7867 two_stage_opamp_dummy_magic_16_0.VD2.n0 two_stage_opamp_dummy_magic_16_0.VD2.t20 16.0005
R7868 two_stage_opamp_dummy_magic_16_0.VD2.t19 two_stage_opamp_dummy_magic_16_0.VD2.n19 16.0005
R7869 two_stage_opamp_dummy_magic_16_0.VD2.n19 two_stage_opamp_dummy_magic_16_0.VD2.t10 16.0005
R7870 two_stage_opamp_dummy_magic_16_0.VD2.n11 two_stage_opamp_dummy_magic_16_0.VD2.n10 4.5005
R7871 two_stage_opamp_dummy_magic_16_0.VD2.n14 two_stage_opamp_dummy_magic_16_0.VD2.n13 4.5005
R7872 two_stage_opamp_dummy_magic_16_0.VD2.n16 two_stage_opamp_dummy_magic_16_0.VD2.n14 3.6255
R7873 two_stage_opamp_dummy_magic_16_0.VD2.n14 two_stage_opamp_dummy_magic_16_0.VD2.n2 1.2505
R7874 two_stage_opamp_dummy_magic_16_0.VD2.n18 two_stage_opamp_dummy_magic_16_0.VD2.n16 1.2505
R7875 two_stage_opamp_dummy_magic_16_0.VD2.n13 two_stage_opamp_dummy_magic_16_0.VD2.n11 0.618871
R7876 two_stage_opamp_dummy_magic_16_0.VD2.n9 two_stage_opamp_dummy_magic_16_0.VD2.n7 0.563
R7877 two_stage_opamp_dummy_magic_16_0.VD2.n10 two_stage_opamp_dummy_magic_16_0.VD2.n9 0.563
R7878 bgr_0.cap_res1.t20 bgr_0.cap_res1.t9 121.245
R7879 bgr_0.cap_res1.t15 bgr_0.cap_res1.t18 0.1603
R7880 bgr_0.cap_res1.t8 bgr_0.cap_res1.t14 0.1603
R7881 bgr_0.cap_res1.t13 bgr_0.cap_res1.t17 0.1603
R7882 bgr_0.cap_res1.t6 bgr_0.cap_res1.t12 0.1603
R7883 bgr_0.cap_res1.t0 bgr_0.cap_res1.t5 0.1603
R7884 bgr_0.cap_res1.n1 bgr_0.cap_res1.t16 0.159278
R7885 bgr_0.cap_res1.n2 bgr_0.cap_res1.t1 0.159278
R7886 bgr_0.cap_res1.n3 bgr_0.cap_res1.t7 0.159278
R7887 bgr_0.cap_res1.n4 bgr_0.cap_res1.t2 0.159278
R7888 bgr_0.cap_res1.n4 bgr_0.cap_res1.t15 0.1368
R7889 bgr_0.cap_res1.n4 bgr_0.cap_res1.t11 0.1368
R7890 bgr_0.cap_res1.n3 bgr_0.cap_res1.t8 0.1368
R7891 bgr_0.cap_res1.n3 bgr_0.cap_res1.t4 0.1368
R7892 bgr_0.cap_res1.n2 bgr_0.cap_res1.t13 0.1368
R7893 bgr_0.cap_res1.n2 bgr_0.cap_res1.t10 0.1368
R7894 bgr_0.cap_res1.n1 bgr_0.cap_res1.t6 0.1368
R7895 bgr_0.cap_res1.n1 bgr_0.cap_res1.t3 0.1368
R7896 bgr_0.cap_res1.n0 bgr_0.cap_res1.t0 0.1368
R7897 bgr_0.cap_res1.n0 bgr_0.cap_res1.t19 0.1368
R7898 bgr_0.cap_res1.t16 bgr_0.cap_res1.n0 0.00152174
R7899 bgr_0.cap_res1.t1 bgr_0.cap_res1.n1 0.00152174
R7900 bgr_0.cap_res1.t7 bgr_0.cap_res1.n2 0.00152174
R7901 bgr_0.cap_res1.t2 bgr_0.cap_res1.n3 0.00152174
R7902 bgr_0.cap_res1.t9 bgr_0.cap_res1.n4 0.00152174
R7903 bgr_0.V_mir2.n20 bgr_0.V_mir2.n19 325.473
R7904 bgr_0.V_mir2.n13 bgr_0.V_mir2.n12 325.473
R7905 bgr_0.V_mir2.n8 bgr_0.V_mir2.n7 325.473
R7906 bgr_0.V_mir2.n16 bgr_0.V_mir2.t21 310.488
R7907 bgr_0.V_mir2.n9 bgr_0.V_mir2.t22 310.488
R7908 bgr_0.V_mir2.n4 bgr_0.V_mir2.t20 310.488
R7909 bgr_0.V_mir2.n2 bgr_0.V_mir2.t14 278.312
R7910 bgr_0.V_mir2.n2 bgr_0.V_mir2.n1 228.939
R7911 bgr_0.V_mir2.n3 bgr_0.V_mir2.n0 224.439
R7912 bgr_0.V_mir2.n18 bgr_0.V_mir2.t10 184.097
R7913 bgr_0.V_mir2.n11 bgr_0.V_mir2.t8 184.097
R7914 bgr_0.V_mir2.n6 bgr_0.V_mir2.t0 184.097
R7915 bgr_0.V_mir2.n17 bgr_0.V_mir2.n16 167.094
R7916 bgr_0.V_mir2.n10 bgr_0.V_mir2.n9 167.094
R7917 bgr_0.V_mir2.n5 bgr_0.V_mir2.n4 167.094
R7918 bgr_0.V_mir2.n13 bgr_0.V_mir2.n11 152
R7919 bgr_0.V_mir2.n8 bgr_0.V_mir2.n6 152
R7920 bgr_0.V_mir2.n19 bgr_0.V_mir2.n18 152
R7921 bgr_0.V_mir2.n16 bgr_0.V_mir2.t19 120.501
R7922 bgr_0.V_mir2.n17 bgr_0.V_mir2.t6 120.501
R7923 bgr_0.V_mir2.n9 bgr_0.V_mir2.t18 120.501
R7924 bgr_0.V_mir2.n10 bgr_0.V_mir2.t2 120.501
R7925 bgr_0.V_mir2.n4 bgr_0.V_mir2.t17 120.501
R7926 bgr_0.V_mir2.n5 bgr_0.V_mir2.t4 120.501
R7927 bgr_0.V_mir2.n1 bgr_0.V_mir2.t16 48.0005
R7928 bgr_0.V_mir2.n1 bgr_0.V_mir2.t12 48.0005
R7929 bgr_0.V_mir2.n0 bgr_0.V_mir2.t15 48.0005
R7930 bgr_0.V_mir2.n0 bgr_0.V_mir2.t13 48.0005
R7931 bgr_0.V_mir2.n18 bgr_0.V_mir2.n17 40.7027
R7932 bgr_0.V_mir2.n11 bgr_0.V_mir2.n10 40.7027
R7933 bgr_0.V_mir2.n6 bgr_0.V_mir2.n5 40.7027
R7934 bgr_0.V_mir2.n12 bgr_0.V_mir2.t3 39.4005
R7935 bgr_0.V_mir2.n12 bgr_0.V_mir2.t9 39.4005
R7936 bgr_0.V_mir2.n7 bgr_0.V_mir2.t5 39.4005
R7937 bgr_0.V_mir2.n7 bgr_0.V_mir2.t1 39.4005
R7938 bgr_0.V_mir2.n20 bgr_0.V_mir2.t7 39.4005
R7939 bgr_0.V_mir2.t11 bgr_0.V_mir2.n20 39.4005
R7940 bgr_0.V_mir2.n14 bgr_0.V_mir2.n13 15.8005
R7941 bgr_0.V_mir2.n14 bgr_0.V_mir2.n8 15.8005
R7942 bgr_0.V_mir2.n19 bgr_0.V_mir2.n15 9.3005
R7943 bgr_0.V_mir2.n3 bgr_0.V_mir2.n2 5.8755
R7944 bgr_0.V_mir2.n15 bgr_0.V_mir2.n14 4.5005
R7945 bgr_0.V_mir2.n15 bgr_0.V_mir2.n3 0.78175
R7946 bgr_0.Vin-.n8 bgr_0.Vin-.t12 688.859
R7947 bgr_0.Vin-.n10 bgr_0.Vin-.n9 514.134
R7948 bgr_0.Vin-.n7 bgr_0.Vin-.n6 351.522
R7949 bgr_0.Vin-.n12 bgr_0.Vin-.n11 213.4
R7950 bgr_0.Vin-.n8 bgr_0.Vin-.t8 174.726
R7951 bgr_0.Vin-.n9 bgr_0.Vin-.t10 174.726
R7952 bgr_0.Vin-.n10 bgr_0.Vin-.t9 174.726
R7953 bgr_0.Vin-.n11 bgr_0.Vin-.t11 174.726
R7954 bgr_0.Vin-.n5 bgr_0.Vin-.n3 173.029
R7955 bgr_0.Vin-.n5 bgr_0.Vin-.n4 168.654
R7956 bgr_0.Vin-.n22 bgr_0.Vin-.n21 141.667
R7957 bgr_0.Vin-.n9 bgr_0.Vin-.n8 128.534
R7958 bgr_0.Vin-.n11 bgr_0.Vin-.n10 128.534
R7959 bgr_0.Vin-.n13 bgr_0.Vin-.t7 119.099
R7960 bgr_0.Vin-.n23 bgr_0.Vin-.n22 84.0884
R7961 bgr_0.Vin-.n18 bgr_0.Vin-.n17 83.5719
R7962 bgr_0.Vin-.n19 bgr_0.Vin-.n0 83.5719
R7963 bgr_0.Vin-.n20 bgr_0.Vin-.n1 83.5719
R7964 bgr_0.Vin-.n15 bgr_0.Vin-.t2 65.0299
R7965 bgr_0.Vin-.n6 bgr_0.Vin-.t0 39.4005
R7966 bgr_0.Vin-.n6 bgr_0.Vin-.t1 39.4005
R7967 bgr_0.Vin-.n14 bgr_0.Vin-.n13 28.813
R7968 bgr_0.Vin-.n19 bgr_0.Vin-.n18 26.074
R7969 bgr_0.Vin-.n20 bgr_0.Vin-.n19 26.074
R7970 bgr_0.Vin-.n22 bgr_0.Vin-.n20 26.074
R7971 bgr_0.Vin-.n13 bgr_0.Vin-.n12 16.188
R7972 bgr_0.Vin-.n4 bgr_0.Vin-.t3 13.1338
R7973 bgr_0.Vin-.n4 bgr_0.Vin-.t5 13.1338
R7974 bgr_0.Vin-.n3 bgr_0.Vin-.t6 13.1338
R7975 bgr_0.Vin-.n3 bgr_0.Vin-.t4 13.1338
R7976 bgr_0.Vin-.n12 bgr_0.Vin-.n7 11.2193
R7977 bgr_0.Vin-.n7 bgr_0.Vin-.n5 3.8755
R7978 bgr_0.Vin-.n24 bgr_0.Vin-.n23 1.56836
R7979 bgr_0.Vin-.n17 bgr_0.Vin-.n15 1.56363
R7980 bgr_0.Vin-.n25 bgr_0.Vin-.n24 1.5505
R7981 bgr_0.Vin-.n16 bgr_0.Vin-.n2 1.5505
R7982 bgr_0.Vin-.n23 bgr_0.Vin-.n1 1.14402
R7983 bgr_0.Vin-.n16 bgr_0.Vin-.n0 0.885803
R7984 bgr_0.Vin-.n17 bgr_0.Vin-.n16 0.77514
R7985 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_0.Vin-.n0 0.756696
R7986 bgr_0.Vin-.n25 bgr_0.Vin-.n1 0.701365
R7987 bgr_0.Vin-.n15 bgr_0.Vin-.n14 0.530034
R7988 bgr_0.Vin-.n18 bgr_0.Vin-.t2 0.290206
R7989 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_0.Vin-.n25 0.203382
R7990 bgr_0.Vin-.n24 bgr_0.Vin-.n2 0.0183571
R7991 bgr_0.Vin-.n14 bgr_0.Vin-.n2 0.00817857
R7992 bgr_0.V_p_1.n1 bgr_0.V_p_1.n4 229.562
R7993 bgr_0.V_p_1.n1 bgr_0.V_p_1.n5 228.939
R7994 bgr_0.V_p_1.n0 bgr_0.V_p_1.n3 228.939
R7995 bgr_0.V_p_1.n0 bgr_0.V_p_1.n2 228.939
R7996 bgr_0.V_p_1.n6 bgr_0.V_p_1.n0 228.938
R7997 bgr_0.V_p_1.n0 bgr_0.V_p_1.t5 98.7279
R7998 bgr_0.V_p_1.n5 bgr_0.V_p_1.t10 48.0005
R7999 bgr_0.V_p_1.n5 bgr_0.V_p_1.t1 48.0005
R8000 bgr_0.V_p_1.n4 bgr_0.V_p_1.t2 48.0005
R8001 bgr_0.V_p_1.n4 bgr_0.V_p_1.t6 48.0005
R8002 bgr_0.V_p_1.n3 bgr_0.V_p_1.t9 48.0005
R8003 bgr_0.V_p_1.n3 bgr_0.V_p_1.t0 48.0005
R8004 bgr_0.V_p_1.n2 bgr_0.V_p_1.t3 48.0005
R8005 bgr_0.V_p_1.n2 bgr_0.V_p_1.t7 48.0005
R8006 bgr_0.V_p_1.t4 bgr_0.V_p_1.n6 48.0005
R8007 bgr_0.V_p_1.n6 bgr_0.V_p_1.t8 48.0005
R8008 bgr_0.V_p_1.n0 bgr_0.V_p_1.n1 1.8755
R8009 two_stage_opamp_dummy_magic_16_0.Y.n47 two_stage_opamp_dummy_magic_16_0.Y.t27 1172.87
R8010 two_stage_opamp_dummy_magic_16_0.Y.n43 two_stage_opamp_dummy_magic_16_0.Y.t33 1172.87
R8011 two_stage_opamp_dummy_magic_16_0.Y.n50 two_stage_opamp_dummy_magic_16_0.Y.t45 996.134
R8012 two_stage_opamp_dummy_magic_16_0.Y.n49 two_stage_opamp_dummy_magic_16_0.Y.t30 996.134
R8013 two_stage_opamp_dummy_magic_16_0.Y.n48 two_stage_opamp_dummy_magic_16_0.Y.t47 996.134
R8014 two_stage_opamp_dummy_magic_16_0.Y.n47 two_stage_opamp_dummy_magic_16_0.Y.t41 996.134
R8015 two_stage_opamp_dummy_magic_16_0.Y.n43 two_stage_opamp_dummy_magic_16_0.Y.t49 996.134
R8016 two_stage_opamp_dummy_magic_16_0.Y.n44 two_stage_opamp_dummy_magic_16_0.Y.t35 996.134
R8017 two_stage_opamp_dummy_magic_16_0.Y.n45 two_stage_opamp_dummy_magic_16_0.Y.t52 996.134
R8018 two_stage_opamp_dummy_magic_16_0.Y.n46 two_stage_opamp_dummy_magic_16_0.Y.t38 996.134
R8019 two_stage_opamp_dummy_magic_16_0.Y.n23 two_stage_opamp_dummy_magic_16_0.Y.t32 690.867
R8020 two_stage_opamp_dummy_magic_16_0.Y.n20 two_stage_opamp_dummy_magic_16_0.Y.t39 690.867
R8021 two_stage_opamp_dummy_magic_16_0.Y.n14 two_stage_opamp_dummy_magic_16_0.Y.t44 530.201
R8022 two_stage_opamp_dummy_magic_16_0.Y.n11 two_stage_opamp_dummy_magic_16_0.Y.t51 530.201
R8023 two_stage_opamp_dummy_magic_16_0.Y.n23 two_stage_opamp_dummy_magic_16_0.Y.t46 514.134
R8024 two_stage_opamp_dummy_magic_16_0.Y.n24 two_stage_opamp_dummy_magic_16_0.Y.t53 514.134
R8025 two_stage_opamp_dummy_magic_16_0.Y.n25 two_stage_opamp_dummy_magic_16_0.Y.t36 514.134
R8026 two_stage_opamp_dummy_magic_16_0.Y.n26 two_stage_opamp_dummy_magic_16_0.Y.t50 514.134
R8027 two_stage_opamp_dummy_magic_16_0.Y.n27 two_stage_opamp_dummy_magic_16_0.Y.t43 514.134
R8028 two_stage_opamp_dummy_magic_16_0.Y.n22 two_stage_opamp_dummy_magic_16_0.Y.t28 514.134
R8029 two_stage_opamp_dummy_magic_16_0.Y.n21 two_stage_opamp_dummy_magic_16_0.Y.t42 514.134
R8030 two_stage_opamp_dummy_magic_16_0.Y.n20 two_stage_opamp_dummy_magic_16_0.Y.t25 514.134
R8031 two_stage_opamp_dummy_magic_16_0.Y.n18 two_stage_opamp_dummy_magic_16_0.Y.t26 353.467
R8032 two_stage_opamp_dummy_magic_16_0.Y.n17 two_stage_opamp_dummy_magic_16_0.Y.t31 353.467
R8033 two_stage_opamp_dummy_magic_16_0.Y.n16 two_stage_opamp_dummy_magic_16_0.Y.t48 353.467
R8034 two_stage_opamp_dummy_magic_16_0.Y.n15 two_stage_opamp_dummy_magic_16_0.Y.t34 353.467
R8035 two_stage_opamp_dummy_magic_16_0.Y.n14 two_stage_opamp_dummy_magic_16_0.Y.t29 353.467
R8036 two_stage_opamp_dummy_magic_16_0.Y.n11 two_stage_opamp_dummy_magic_16_0.Y.t37 353.467
R8037 two_stage_opamp_dummy_magic_16_0.Y.n12 two_stage_opamp_dummy_magic_16_0.Y.t54 353.467
R8038 two_stage_opamp_dummy_magic_16_0.Y.n13 two_stage_opamp_dummy_magic_16_0.Y.t40 353.467
R8039 two_stage_opamp_dummy_magic_16_0.Y.n50 two_stage_opamp_dummy_magic_16_0.Y.n49 176.733
R8040 two_stage_opamp_dummy_magic_16_0.Y.n49 two_stage_opamp_dummy_magic_16_0.Y.n48 176.733
R8041 two_stage_opamp_dummy_magic_16_0.Y.n48 two_stage_opamp_dummy_magic_16_0.Y.n47 176.733
R8042 two_stage_opamp_dummy_magic_16_0.Y.n44 two_stage_opamp_dummy_magic_16_0.Y.n43 176.733
R8043 two_stage_opamp_dummy_magic_16_0.Y.n45 two_stage_opamp_dummy_magic_16_0.Y.n44 176.733
R8044 two_stage_opamp_dummy_magic_16_0.Y.n46 two_stage_opamp_dummy_magic_16_0.Y.n45 176.733
R8045 two_stage_opamp_dummy_magic_16_0.Y.n18 two_stage_opamp_dummy_magic_16_0.Y.n17 176.733
R8046 two_stage_opamp_dummy_magic_16_0.Y.n17 two_stage_opamp_dummy_magic_16_0.Y.n16 176.733
R8047 two_stage_opamp_dummy_magic_16_0.Y.n16 two_stage_opamp_dummy_magic_16_0.Y.n15 176.733
R8048 two_stage_opamp_dummy_magic_16_0.Y.n15 two_stage_opamp_dummy_magic_16_0.Y.n14 176.733
R8049 two_stage_opamp_dummy_magic_16_0.Y.n12 two_stage_opamp_dummy_magic_16_0.Y.n11 176.733
R8050 two_stage_opamp_dummy_magic_16_0.Y.n13 two_stage_opamp_dummy_magic_16_0.Y.n12 176.733
R8051 two_stage_opamp_dummy_magic_16_0.Y.n27 two_stage_opamp_dummy_magic_16_0.Y.n26 176.733
R8052 two_stage_opamp_dummy_magic_16_0.Y.n26 two_stage_opamp_dummy_magic_16_0.Y.n25 176.733
R8053 two_stage_opamp_dummy_magic_16_0.Y.n25 two_stage_opamp_dummy_magic_16_0.Y.n24 176.733
R8054 two_stage_opamp_dummy_magic_16_0.Y.n24 two_stage_opamp_dummy_magic_16_0.Y.n23 176.733
R8055 two_stage_opamp_dummy_magic_16_0.Y.n21 two_stage_opamp_dummy_magic_16_0.Y.n20 176.733
R8056 two_stage_opamp_dummy_magic_16_0.Y.n22 two_stage_opamp_dummy_magic_16_0.Y.n21 176.733
R8057 two_stage_opamp_dummy_magic_16_0.Y.n52 two_stage_opamp_dummy_magic_16_0.Y.n51 166.258
R8058 two_stage_opamp_dummy_magic_16_0.Y.n2 two_stage_opamp_dummy_magic_16_0.Y.n0 163.626
R8059 two_stage_opamp_dummy_magic_16_0.Y.n8 two_stage_opamp_dummy_magic_16_0.Y.n7 163.001
R8060 two_stage_opamp_dummy_magic_16_0.Y.n6 two_stage_opamp_dummy_magic_16_0.Y.n5 163.001
R8061 two_stage_opamp_dummy_magic_16_0.Y.n4 two_stage_opamp_dummy_magic_16_0.Y.n3 163.001
R8062 two_stage_opamp_dummy_magic_16_0.Y.n2 two_stage_opamp_dummy_magic_16_0.Y.n1 163.001
R8063 two_stage_opamp_dummy_magic_16_0.Y.n29 two_stage_opamp_dummy_magic_16_0.Y.n19 161.541
R8064 two_stage_opamp_dummy_magic_16_0.Y.n29 two_stage_opamp_dummy_magic_16_0.Y.n28 161.541
R8065 two_stage_opamp_dummy_magic_16_0.Y.n10 two_stage_opamp_dummy_magic_16_0.Y.n9 158.501
R8066 two_stage_opamp_dummy_magic_16_0.Y.n32 two_stage_opamp_dummy_magic_16_0.Y.n30 117.906
R8067 two_stage_opamp_dummy_magic_16_0.Y.n40 two_stage_opamp_dummy_magic_16_0.Y.n39 117.326
R8068 two_stage_opamp_dummy_magic_16_0.Y.n38 two_stage_opamp_dummy_magic_16_0.Y.n37 117.326
R8069 two_stage_opamp_dummy_magic_16_0.Y.n36 two_stage_opamp_dummy_magic_16_0.Y.n35 117.326
R8070 two_stage_opamp_dummy_magic_16_0.Y.n34 two_stage_opamp_dummy_magic_16_0.Y.n33 117.326
R8071 two_stage_opamp_dummy_magic_16_0.Y.n32 two_stage_opamp_dummy_magic_16_0.Y.n31 117.326
R8072 two_stage_opamp_dummy_magic_16_0.Y.n19 two_stage_opamp_dummy_magic_16_0.Y.n18 54.6272
R8073 two_stage_opamp_dummy_magic_16_0.Y.n19 two_stage_opamp_dummy_magic_16_0.Y.n13 54.6272
R8074 two_stage_opamp_dummy_magic_16_0.Y.n28 two_stage_opamp_dummy_magic_16_0.Y.n27 54.6272
R8075 two_stage_opamp_dummy_magic_16_0.Y.n28 two_stage_opamp_dummy_magic_16_0.Y.n22 54.6272
R8076 two_stage_opamp_dummy_magic_16_0.Y.n51 two_stage_opamp_dummy_magic_16_0.Y.n50 53.3126
R8077 two_stage_opamp_dummy_magic_16_0.Y.n51 two_stage_opamp_dummy_magic_16_0.Y.n46 53.3126
R8078 two_stage_opamp_dummy_magic_16_0.Y.t1 two_stage_opamp_dummy_magic_16_0.Y.n52 50.3031
R8079 two_stage_opamp_dummy_magic_16_0.Y.n42 two_stage_opamp_dummy_magic_16_0.Y.n10 16.8755
R8080 two_stage_opamp_dummy_magic_16_0.Y.n39 two_stage_opamp_dummy_magic_16_0.Y.t6 16.0005
R8081 two_stage_opamp_dummy_magic_16_0.Y.n39 two_stage_opamp_dummy_magic_16_0.Y.t13 16.0005
R8082 two_stage_opamp_dummy_magic_16_0.Y.n37 two_stage_opamp_dummy_magic_16_0.Y.t7 16.0005
R8083 two_stage_opamp_dummy_magic_16_0.Y.n37 two_stage_opamp_dummy_magic_16_0.Y.t2 16.0005
R8084 two_stage_opamp_dummy_magic_16_0.Y.n35 two_stage_opamp_dummy_magic_16_0.Y.t9 16.0005
R8085 two_stage_opamp_dummy_magic_16_0.Y.n35 two_stage_opamp_dummy_magic_16_0.Y.t3 16.0005
R8086 two_stage_opamp_dummy_magic_16_0.Y.n33 two_stage_opamp_dummy_magic_16_0.Y.t8 16.0005
R8087 two_stage_opamp_dummy_magic_16_0.Y.n33 two_stage_opamp_dummy_magic_16_0.Y.t11 16.0005
R8088 two_stage_opamp_dummy_magic_16_0.Y.n31 two_stage_opamp_dummy_magic_16_0.Y.t10 16.0005
R8089 two_stage_opamp_dummy_magic_16_0.Y.n31 two_stage_opamp_dummy_magic_16_0.Y.t4 16.0005
R8090 two_stage_opamp_dummy_magic_16_0.Y.n30 two_stage_opamp_dummy_magic_16_0.Y.t14 16.0005
R8091 two_stage_opamp_dummy_magic_16_0.Y.n30 two_stage_opamp_dummy_magic_16_0.Y.t5 16.0005
R8092 two_stage_opamp_dummy_magic_16_0.Y.n41 two_stage_opamp_dummy_magic_16_0.Y.n29 12.4067
R8093 two_stage_opamp_dummy_magic_16_0.Y.n9 two_stage_opamp_dummy_magic_16_0.Y.t18 11.2576
R8094 two_stage_opamp_dummy_magic_16_0.Y.n9 two_stage_opamp_dummy_magic_16_0.Y.t0 11.2576
R8095 two_stage_opamp_dummy_magic_16_0.Y.n7 two_stage_opamp_dummy_magic_16_0.Y.t20 11.2576
R8096 two_stage_opamp_dummy_magic_16_0.Y.n7 two_stage_opamp_dummy_magic_16_0.Y.t17 11.2576
R8097 two_stage_opamp_dummy_magic_16_0.Y.n5 two_stage_opamp_dummy_magic_16_0.Y.t15 11.2576
R8098 two_stage_opamp_dummy_magic_16_0.Y.n5 two_stage_opamp_dummy_magic_16_0.Y.t16 11.2576
R8099 two_stage_opamp_dummy_magic_16_0.Y.n3 two_stage_opamp_dummy_magic_16_0.Y.t23 11.2576
R8100 two_stage_opamp_dummy_magic_16_0.Y.n3 two_stage_opamp_dummy_magic_16_0.Y.t24 11.2576
R8101 two_stage_opamp_dummy_magic_16_0.Y.n1 two_stage_opamp_dummy_magic_16_0.Y.t22 11.2576
R8102 two_stage_opamp_dummy_magic_16_0.Y.n1 two_stage_opamp_dummy_magic_16_0.Y.t19 11.2576
R8103 two_stage_opamp_dummy_magic_16_0.Y.n0 two_stage_opamp_dummy_magic_16_0.Y.t12 11.2576
R8104 two_stage_opamp_dummy_magic_16_0.Y.n0 two_stage_opamp_dummy_magic_16_0.Y.t21 11.2576
R8105 two_stage_opamp_dummy_magic_16_0.Y.n52 two_stage_opamp_dummy_magic_16_0.Y.n42 7.09425
R8106 two_stage_opamp_dummy_magic_16_0.Y.n41 two_stage_opamp_dummy_magic_16_0.Y.n40 6.38443
R8107 two_stage_opamp_dummy_magic_16_0.Y.n10 two_stage_opamp_dummy_magic_16_0.Y.n8 5.1255
R8108 two_stage_opamp_dummy_magic_16_0.Y.n42 two_stage_opamp_dummy_magic_16_0.Y.n41 0.938
R8109 two_stage_opamp_dummy_magic_16_0.Y.n4 two_stage_opamp_dummy_magic_16_0.Y.n2 0.6255
R8110 two_stage_opamp_dummy_magic_16_0.Y.n6 two_stage_opamp_dummy_magic_16_0.Y.n4 0.6255
R8111 two_stage_opamp_dummy_magic_16_0.Y.n8 two_stage_opamp_dummy_magic_16_0.Y.n6 0.6255
R8112 two_stage_opamp_dummy_magic_16_0.Y.n34 two_stage_opamp_dummy_magic_16_0.Y.n32 0.580857
R8113 two_stage_opamp_dummy_magic_16_0.Y.n36 two_stage_opamp_dummy_magic_16_0.Y.n34 0.580857
R8114 two_stage_opamp_dummy_magic_16_0.Y.n38 two_stage_opamp_dummy_magic_16_0.Y.n36 0.580857
R8115 two_stage_opamp_dummy_magic_16_0.Y.n40 two_stage_opamp_dummy_magic_16_0.Y.n38 0.580857
R8116 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n0 144.827
R8117 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n1 134.577
R8118 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t10 118.986
R8119 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n3 100.6
R8120 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n10 100.038
R8121 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n8 100.038
R8122 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n6 100.038
R8123 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n4 100.038
R8124 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n12 43.284
R8125 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n2 37.4067
R8126 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t13 24.0005
R8127 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t11 24.0005
R8128 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t14 24.0005
R8129 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t12 24.0005
R8130 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t2 8.0005
R8131 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t7 8.0005
R8132 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t6 8.0005
R8133 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t0 8.0005
R8134 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t3 8.0005
R8135 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t1 8.0005
R8136 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t4 8.0005
R8137 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t8 8.0005
R8138 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t5 8.0005
R8139 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t9 8.0005
R8140 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n11 5.6255
R8141 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n5 0.563
R8142 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n7 0.563
R8143 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n9 0.563
R8144 bgr_0.V_CMFB_S4 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n13 0.047375
R8145 a_9610_2730.n1 a_9610_2730.n0 114.469
R8146 a_9610_2730.n2 a_9610_2730.n1 113.906
R8147 a_9610_2730.n1 a_9610_2730.t0 96.77
R8148 a_9610_2730.n0 a_9610_2730.t4 16.0005
R8149 a_9610_2730.n0 a_9610_2730.t2 16.0005
R8150 a_9610_2730.n2 a_9610_2730.t1 16.0005
R8151 a_9610_2730.t3 a_9610_2730.n2 16.0005
R8152 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n0 345.264
R8153 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n1 344.7
R8154 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n3 292.5
R8155 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n5 209.251
R8156 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n12 208.689
R8157 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n10 208.689
R8158 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n8 208.689
R8159 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n6 208.689
R8160 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t16 120.305
R8161 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n2 52.763
R8162 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n4 51.7297
R8163 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n14 50.813
R8164 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t14 39.4005
R8165 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t13 39.4005
R8166 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t11 39.4005
R8167 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t10 39.4005
R8168 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t12 39.4005
R8169 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t15 39.4005
R8170 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t8 19.7005
R8171 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t3 19.7005
R8172 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t2 19.7005
R8173 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t6 19.7005
R8174 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t9 19.7005
R8175 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t7 19.7005
R8176 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t0 19.7005
R8177 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t4 19.7005
R8178 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t1 19.7005
R8179 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t5 19.7005
R8180 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n13 5.90675
R8181 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n7 0.563
R8182 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n9 0.563
R8183 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n11 0.563
R8184 two_stage_opamp_dummy_magic_16_0.VD4.n28 two_stage_opamp_dummy_magic_16_0.VD4.t15 652.076
R8185 two_stage_opamp_dummy_magic_16_0.VD4.n61 two_stage_opamp_dummy_magic_16_0.VD4.t12 652.076
R8186 two_stage_opamp_dummy_magic_16_0.VD4.n60 two_stage_opamp_dummy_magic_16_0.VD4.n13 585
R8187 two_stage_opamp_dummy_magic_16_0.VD4.n42 two_stage_opamp_dummy_magic_16_0.VD4.n41 585
R8188 two_stage_opamp_dummy_magic_16_0.VD4.n48 two_stage_opamp_dummy_magic_16_0.VD4.n13 290.233
R8189 two_stage_opamp_dummy_magic_16_0.VD4.n54 two_stage_opamp_dummy_magic_16_0.VD4.n13 290.233
R8190 two_stage_opamp_dummy_magic_16_0.VD4.n49 two_stage_opamp_dummy_magic_16_0.VD4.n13 290.233
R8191 two_stage_opamp_dummy_magic_16_0.VD4.n41 two_stage_opamp_dummy_magic_16_0.VD4.n30 290.233
R8192 two_stage_opamp_dummy_magic_16_0.VD4.n41 two_stage_opamp_dummy_magic_16_0.VD4.n35 290.233
R8193 two_stage_opamp_dummy_magic_16_0.VD4.n41 two_stage_opamp_dummy_magic_16_0.VD4.n40 290.233
R8194 two_stage_opamp_dummy_magic_16_0.VD4.n49 two_stage_opamp_dummy_magic_16_0.VD4.n46 242.903
R8195 two_stage_opamp_dummy_magic_16_0.VD4.n40 two_stage_opamp_dummy_magic_16_0.VD4.n18 242.903
R8196 two_stage_opamp_dummy_magic_16_0.VD4.n60 two_stage_opamp_dummy_magic_16_0.VD4.n59 238.367
R8197 two_stage_opamp_dummy_magic_16_0.VD4.n15 two_stage_opamp_dummy_magic_16_0.VD4.n14 185
R8198 two_stage_opamp_dummy_magic_16_0.VD4.n57 two_stage_opamp_dummy_magic_16_0.VD4.n56 185
R8199 two_stage_opamp_dummy_magic_16_0.VD4.n58 two_stage_opamp_dummy_magic_16_0.VD4.n57 185
R8200 two_stage_opamp_dummy_magic_16_0.VD4.n55 two_stage_opamp_dummy_magic_16_0.VD4.n47 185
R8201 two_stage_opamp_dummy_magic_16_0.VD4.n53 two_stage_opamp_dummy_magic_16_0.VD4.n52 185
R8202 two_stage_opamp_dummy_magic_16_0.VD4.n51 two_stage_opamp_dummy_magic_16_0.VD4.n50 185
R8203 two_stage_opamp_dummy_magic_16_0.VD4.n43 two_stage_opamp_dummy_magic_16_0.VD4.n42 185
R8204 two_stage_opamp_dummy_magic_16_0.VD4.n44 two_stage_opamp_dummy_magic_16_0.VD4.n43 185
R8205 two_stage_opamp_dummy_magic_16_0.VD4.n29 two_stage_opamp_dummy_magic_16_0.VD4.n19 185
R8206 two_stage_opamp_dummy_magic_16_0.VD4.n32 two_stage_opamp_dummy_magic_16_0.VD4.n31 185
R8207 two_stage_opamp_dummy_magic_16_0.VD4.n34 two_stage_opamp_dummy_magic_16_0.VD4.n33 185
R8208 two_stage_opamp_dummy_magic_16_0.VD4.n37 two_stage_opamp_dummy_magic_16_0.VD4.n36 185
R8209 two_stage_opamp_dummy_magic_16_0.VD4.n39 two_stage_opamp_dummy_magic_16_0.VD4.n38 185
R8210 two_stage_opamp_dummy_magic_16_0.VD4.t16 two_stage_opamp_dummy_magic_16_0.VD4.n44 170.513
R8211 two_stage_opamp_dummy_magic_16_0.VD4.n58 two_stage_opamp_dummy_magic_16_0.VD4.t13 170.513
R8212 two_stage_opamp_dummy_magic_16_0.VD4.n2 two_stage_opamp_dummy_magic_16_0.VD4.n0 163.626
R8213 two_stage_opamp_dummy_magic_16_0.VD4.n10 two_stage_opamp_dummy_magic_16_0.VD4.n9 163.001
R8214 two_stage_opamp_dummy_magic_16_0.VD4.n8 two_stage_opamp_dummy_magic_16_0.VD4.n7 163.001
R8215 two_stage_opamp_dummy_magic_16_0.VD4.n6 two_stage_opamp_dummy_magic_16_0.VD4.n5 163.001
R8216 two_stage_opamp_dummy_magic_16_0.VD4.n4 two_stage_opamp_dummy_magic_16_0.VD4.n3 163.001
R8217 two_stage_opamp_dummy_magic_16_0.VD4.n2 two_stage_opamp_dummy_magic_16_0.VD4.n1 163.001
R8218 two_stage_opamp_dummy_magic_16_0.VD4.n12 two_stage_opamp_dummy_magic_16_0.VD4.n11 159.804
R8219 two_stage_opamp_dummy_magic_16_0.VD4.n21 two_stage_opamp_dummy_magic_16_0.VD4.n20 159.803
R8220 two_stage_opamp_dummy_magic_16_0.VD4.n23 two_stage_opamp_dummy_magic_16_0.VD4.n22 159.803
R8221 two_stage_opamp_dummy_magic_16_0.VD4.n25 two_stage_opamp_dummy_magic_16_0.VD4.n24 159.803
R8222 two_stage_opamp_dummy_magic_16_0.VD4.n27 two_stage_opamp_dummy_magic_16_0.VD4.n26 159.803
R8223 two_stage_opamp_dummy_magic_16_0.VD4.n57 two_stage_opamp_dummy_magic_16_0.VD4.n15 150
R8224 two_stage_opamp_dummy_magic_16_0.VD4.n57 two_stage_opamp_dummy_magic_16_0.VD4.n47 150
R8225 two_stage_opamp_dummy_magic_16_0.VD4.n52 two_stage_opamp_dummy_magic_16_0.VD4.n51 150
R8226 two_stage_opamp_dummy_magic_16_0.VD4.n43 two_stage_opamp_dummy_magic_16_0.VD4.n19 150
R8227 two_stage_opamp_dummy_magic_16_0.VD4.n33 two_stage_opamp_dummy_magic_16_0.VD4.n32 150
R8228 two_stage_opamp_dummy_magic_16_0.VD4.n38 two_stage_opamp_dummy_magic_16_0.VD4.n37 150
R8229 two_stage_opamp_dummy_magic_16_0.VD4.t28 two_stage_opamp_dummy_magic_16_0.VD4.t16 146.155
R8230 two_stage_opamp_dummy_magic_16_0.VD4.t24 two_stage_opamp_dummy_magic_16_0.VD4.t28 146.155
R8231 two_stage_opamp_dummy_magic_16_0.VD4.t30 two_stage_opamp_dummy_magic_16_0.VD4.t24 146.155
R8232 two_stage_opamp_dummy_magic_16_0.VD4.t34 two_stage_opamp_dummy_magic_16_0.VD4.t30 146.155
R8233 two_stage_opamp_dummy_magic_16_0.VD4.t18 two_stage_opamp_dummy_magic_16_0.VD4.t34 146.155
R8234 two_stage_opamp_dummy_magic_16_0.VD4.t20 two_stage_opamp_dummy_magic_16_0.VD4.t18 146.155
R8235 two_stage_opamp_dummy_magic_16_0.VD4.t22 two_stage_opamp_dummy_magic_16_0.VD4.t20 146.155
R8236 two_stage_opamp_dummy_magic_16_0.VD4.t26 two_stage_opamp_dummy_magic_16_0.VD4.t22 146.155
R8237 two_stage_opamp_dummy_magic_16_0.VD4.t32 two_stage_opamp_dummy_magic_16_0.VD4.t26 146.155
R8238 two_stage_opamp_dummy_magic_16_0.VD4.t36 two_stage_opamp_dummy_magic_16_0.VD4.t32 146.155
R8239 two_stage_opamp_dummy_magic_16_0.VD4.t13 two_stage_opamp_dummy_magic_16_0.VD4.t36 146.155
R8240 two_stage_opamp_dummy_magic_16_0.VD4.n59 two_stage_opamp_dummy_magic_16_0.VD4.n58 65.8183
R8241 two_stage_opamp_dummy_magic_16_0.VD4.n58 two_stage_opamp_dummy_magic_16_0.VD4.n45 65.8183
R8242 two_stage_opamp_dummy_magic_16_0.VD4.n58 two_stage_opamp_dummy_magic_16_0.VD4.n46 65.8183
R8243 two_stage_opamp_dummy_magic_16_0.VD4.n44 two_stage_opamp_dummy_magic_16_0.VD4.n16 65.8183
R8244 two_stage_opamp_dummy_magic_16_0.VD4.n44 two_stage_opamp_dummy_magic_16_0.VD4.n17 65.8183
R8245 two_stage_opamp_dummy_magic_16_0.VD4.n44 two_stage_opamp_dummy_magic_16_0.VD4.n18 65.8183
R8246 two_stage_opamp_dummy_magic_16_0.VD4.n47 two_stage_opamp_dummy_magic_16_0.VD4.n45 53.3664
R8247 two_stage_opamp_dummy_magic_16_0.VD4.n51 two_stage_opamp_dummy_magic_16_0.VD4.n46 53.3664
R8248 two_stage_opamp_dummy_magic_16_0.VD4.n59 two_stage_opamp_dummy_magic_16_0.VD4.n15 53.3664
R8249 two_stage_opamp_dummy_magic_16_0.VD4.n52 two_stage_opamp_dummy_magic_16_0.VD4.n45 53.3664
R8250 two_stage_opamp_dummy_magic_16_0.VD4.n19 two_stage_opamp_dummy_magic_16_0.VD4.n16 53.3664
R8251 two_stage_opamp_dummy_magic_16_0.VD4.n33 two_stage_opamp_dummy_magic_16_0.VD4.n17 53.3664
R8252 two_stage_opamp_dummy_magic_16_0.VD4.n38 two_stage_opamp_dummy_magic_16_0.VD4.n18 53.3664
R8253 two_stage_opamp_dummy_magic_16_0.VD4.n32 two_stage_opamp_dummy_magic_16_0.VD4.n16 53.3664
R8254 two_stage_opamp_dummy_magic_16_0.VD4.n37 two_stage_opamp_dummy_magic_16_0.VD4.n17 53.3664
R8255 two_stage_opamp_dummy_magic_16_0.VD4.n61 two_stage_opamp_dummy_magic_16_0.VD4.n60 22.8576
R8256 two_stage_opamp_dummy_magic_16_0.VD4.n42 two_stage_opamp_dummy_magic_16_0.VD4.n28 22.8576
R8257 two_stage_opamp_dummy_magic_16_0.VD4.n28 two_stage_opamp_dummy_magic_16_0.VD4.n27 14.4255
R8258 two_stage_opamp_dummy_magic_16_0.VD4.n62 two_stage_opamp_dummy_magic_16_0.VD4.n61 13.8005
R8259 two_stage_opamp_dummy_magic_16_0.VD4.n20 two_stage_opamp_dummy_magic_16_0.VD4.t23 11.2576
R8260 two_stage_opamp_dummy_magic_16_0.VD4.n20 two_stage_opamp_dummy_magic_16_0.VD4.t27 11.2576
R8261 two_stage_opamp_dummy_magic_16_0.VD4.n22 two_stage_opamp_dummy_magic_16_0.VD4.t19 11.2576
R8262 two_stage_opamp_dummy_magic_16_0.VD4.n22 two_stage_opamp_dummy_magic_16_0.VD4.t21 11.2576
R8263 two_stage_opamp_dummy_magic_16_0.VD4.n24 two_stage_opamp_dummy_magic_16_0.VD4.t31 11.2576
R8264 two_stage_opamp_dummy_magic_16_0.VD4.n24 two_stage_opamp_dummy_magic_16_0.VD4.t35 11.2576
R8265 two_stage_opamp_dummy_magic_16_0.VD4.n26 two_stage_opamp_dummy_magic_16_0.VD4.t29 11.2576
R8266 two_stage_opamp_dummy_magic_16_0.VD4.n26 two_stage_opamp_dummy_magic_16_0.VD4.t25 11.2576
R8267 two_stage_opamp_dummy_magic_16_0.VD4.n41 two_stage_opamp_dummy_magic_16_0.VD4.t17 11.2576
R8268 two_stage_opamp_dummy_magic_16_0.VD4.n13 two_stage_opamp_dummy_magic_16_0.VD4.t14 11.2576
R8269 two_stage_opamp_dummy_magic_16_0.VD4.n9 two_stage_opamp_dummy_magic_16_0.VD4.t10 11.2576
R8270 two_stage_opamp_dummy_magic_16_0.VD4.n9 two_stage_opamp_dummy_magic_16_0.VD4.t4 11.2576
R8271 two_stage_opamp_dummy_magic_16_0.VD4.n7 two_stage_opamp_dummy_magic_16_0.VD4.t2 11.2576
R8272 two_stage_opamp_dummy_magic_16_0.VD4.n7 two_stage_opamp_dummy_magic_16_0.VD4.t5 11.2576
R8273 two_stage_opamp_dummy_magic_16_0.VD4.n5 two_stage_opamp_dummy_magic_16_0.VD4.t7 11.2576
R8274 two_stage_opamp_dummy_magic_16_0.VD4.n5 two_stage_opamp_dummy_magic_16_0.VD4.t9 11.2576
R8275 two_stage_opamp_dummy_magic_16_0.VD4.n3 two_stage_opamp_dummy_magic_16_0.VD4.t1 11.2576
R8276 two_stage_opamp_dummy_magic_16_0.VD4.n3 two_stage_opamp_dummy_magic_16_0.VD4.t0 11.2576
R8277 two_stage_opamp_dummy_magic_16_0.VD4.n1 two_stage_opamp_dummy_magic_16_0.VD4.t3 11.2576
R8278 two_stage_opamp_dummy_magic_16_0.VD4.n1 two_stage_opamp_dummy_magic_16_0.VD4.t6 11.2576
R8279 two_stage_opamp_dummy_magic_16_0.VD4.n0 two_stage_opamp_dummy_magic_16_0.VD4.t8 11.2576
R8280 two_stage_opamp_dummy_magic_16_0.VD4.n0 two_stage_opamp_dummy_magic_16_0.VD4.t11 11.2576
R8281 two_stage_opamp_dummy_magic_16_0.VD4.n11 two_stage_opamp_dummy_magic_16_0.VD4.t33 11.2576
R8282 two_stage_opamp_dummy_magic_16_0.VD4.n11 two_stage_opamp_dummy_magic_16_0.VD4.t37 11.2576
R8283 two_stage_opamp_dummy_magic_16_0.VD4.n60 two_stage_opamp_dummy_magic_16_0.VD4.n14 9.14336
R8284 two_stage_opamp_dummy_magic_16_0.VD4.n56 two_stage_opamp_dummy_magic_16_0.VD4.n55 9.14336
R8285 two_stage_opamp_dummy_magic_16_0.VD4.n53 two_stage_opamp_dummy_magic_16_0.VD4.n50 9.14336
R8286 two_stage_opamp_dummy_magic_16_0.VD4.n42 two_stage_opamp_dummy_magic_16_0.VD4.n29 9.14336
R8287 two_stage_opamp_dummy_magic_16_0.VD4.n34 two_stage_opamp_dummy_magic_16_0.VD4.n31 9.14336
R8288 two_stage_opamp_dummy_magic_16_0.VD4.n39 two_stage_opamp_dummy_magic_16_0.VD4.n36 9.14336
R8289 two_stage_opamp_dummy_magic_16_0.VD4.n63 two_stage_opamp_dummy_magic_16_0.VD4.n10 8.2505
R8290 two_stage_opamp_dummy_magic_16_0.VD4.n63 two_stage_opamp_dummy_magic_16_0.VD4.n62 5.3755
R8291 two_stage_opamp_dummy_magic_16_0.VD4.n48 two_stage_opamp_dummy_magic_16_0.VD4.n14 4.53698
R8292 two_stage_opamp_dummy_magic_16_0.VD4.n55 two_stage_opamp_dummy_magic_16_0.VD4.n54 4.53698
R8293 two_stage_opamp_dummy_magic_16_0.VD4.n50 two_stage_opamp_dummy_magic_16_0.VD4.n49 4.53698
R8294 two_stage_opamp_dummy_magic_16_0.VD4.n56 two_stage_opamp_dummy_magic_16_0.VD4.n48 4.53698
R8295 two_stage_opamp_dummy_magic_16_0.VD4.n54 two_stage_opamp_dummy_magic_16_0.VD4.n53 4.53698
R8296 two_stage_opamp_dummy_magic_16_0.VD4.n30 two_stage_opamp_dummy_magic_16_0.VD4.n29 4.53698
R8297 two_stage_opamp_dummy_magic_16_0.VD4.n35 two_stage_opamp_dummy_magic_16_0.VD4.n34 4.53698
R8298 two_stage_opamp_dummy_magic_16_0.VD4.n40 two_stage_opamp_dummy_magic_16_0.VD4.n39 4.53698
R8299 two_stage_opamp_dummy_magic_16_0.VD4.n31 two_stage_opamp_dummy_magic_16_0.VD4.n30 4.53698
R8300 two_stage_opamp_dummy_magic_16_0.VD4.n36 two_stage_opamp_dummy_magic_16_0.VD4.n35 4.53698
R8301 two_stage_opamp_dummy_magic_16_0.VD4.n4 two_stage_opamp_dummy_magic_16_0.VD4.n2 0.6255
R8302 two_stage_opamp_dummy_magic_16_0.VD4.n6 two_stage_opamp_dummy_magic_16_0.VD4.n4 0.6255
R8303 two_stage_opamp_dummy_magic_16_0.VD4.n8 two_stage_opamp_dummy_magic_16_0.VD4.n6 0.6255
R8304 two_stage_opamp_dummy_magic_16_0.VD4.n10 two_stage_opamp_dummy_magic_16_0.VD4.n8 0.6255
R8305 two_stage_opamp_dummy_magic_16_0.VD4.n62 two_stage_opamp_dummy_magic_16_0.VD4.n12 0.6255
R8306 two_stage_opamp_dummy_magic_16_0.VD4.n27 two_stage_opamp_dummy_magic_16_0.VD4.n25 0.6255
R8307 two_stage_opamp_dummy_magic_16_0.VD4.n25 two_stage_opamp_dummy_magic_16_0.VD4.n23 0.6255
R8308 two_stage_opamp_dummy_magic_16_0.VD4.n23 two_stage_opamp_dummy_magic_16_0.VD4.n21 0.6255
R8309 two_stage_opamp_dummy_magic_16_0.VD4.n21 two_stage_opamp_dummy_magic_16_0.VD4.n12 0.6255
R8310 two_stage_opamp_dummy_magic_16_0.VD4 two_stage_opamp_dummy_magic_16_0.VD4.n63 0.063
R8311 bgr_0.START_UP.n4 bgr_0.START_UP.t6 238.322
R8312 bgr_0.START_UP.n4 bgr_0.START_UP.t7 238.322
R8313 bgr_0.START_UP.n3 bgr_0.START_UP.n1 175.56
R8314 bgr_0.START_UP.n3 bgr_0.START_UP.n2 168.936
R8315 bgr_0.START_UP.n5 bgr_0.START_UP.n4 166.925
R8316 bgr_0.START_UP.n0 bgr_0.START_UP.t1 130.001
R8317 bgr_0.START_UP.n0 bgr_0.START_UP.t0 81.7074
R8318 bgr_0.START_UP bgr_0.START_UP.n0 36.9489
R8319 bgr_0.START_UP bgr_0.START_UP.n5 13.4693
R8320 bgr_0.START_UP.n1 bgr_0.START_UP.t2 13.1338
R8321 bgr_0.START_UP.n1 bgr_0.START_UP.t4 13.1338
R8322 bgr_0.START_UP.n2 bgr_0.START_UP.t3 13.1338
R8323 bgr_0.START_UP.n2 bgr_0.START_UP.t5 13.1338
R8324 bgr_0.START_UP.n5 bgr_0.START_UP.n3 4.21925
R8325 two_stage_opamp_dummy_magic_16_0.V_err_gate.n2 two_stage_opamp_dummy_magic_16_0.V_err_gate.t6 479.322
R8326 two_stage_opamp_dummy_magic_16_0.V_err_gate.n2 two_stage_opamp_dummy_magic_16_0.V_err_gate.t8 479.322
R8327 two_stage_opamp_dummy_magic_16_0.V_err_gate.n6 two_stage_opamp_dummy_magic_16_0.V_err_gate.t9 479.322
R8328 two_stage_opamp_dummy_magic_16_0.V_err_gate.n6 two_stage_opamp_dummy_magic_16_0.V_err_gate.t7 479.322
R8329 two_stage_opamp_dummy_magic_16_0.V_err_gate.n3 two_stage_opamp_dummy_magic_16_0.V_err_gate.n1 178.625
R8330 two_stage_opamp_dummy_magic_16_0.V_err_gate.n5 two_stage_opamp_dummy_magic_16_0.V_err_gate.n4 177.987
R8331 two_stage_opamp_dummy_magic_16_0.V_err_gate two_stage_opamp_dummy_magic_16_0.V_err_gate.n0 175.013
R8332 two_stage_opamp_dummy_magic_16_0.V_err_gate.n3 two_stage_opamp_dummy_magic_16_0.V_err_gate.n2 165.8
R8333 two_stage_opamp_dummy_magic_16_0.V_err_gate two_stage_opamp_dummy_magic_16_0.V_err_gate.n6 165.8
R8334 two_stage_opamp_dummy_magic_16_0.V_err_gate.n0 two_stage_opamp_dummy_magic_16_0.V_err_gate.t1 24.0005
R8335 two_stage_opamp_dummy_magic_16_0.V_err_gate.n0 two_stage_opamp_dummy_magic_16_0.V_err_gate.t2 24.0005
R8336 two_stage_opamp_dummy_magic_16_0.V_err_gate.n4 two_stage_opamp_dummy_magic_16_0.V_err_gate.t3 15.7605
R8337 two_stage_opamp_dummy_magic_16_0.V_err_gate.n4 two_stage_opamp_dummy_magic_16_0.V_err_gate.t5 15.7605
R8338 two_stage_opamp_dummy_magic_16_0.V_err_gate.n1 two_stage_opamp_dummy_magic_16_0.V_err_gate.t0 15.7605
R8339 two_stage_opamp_dummy_magic_16_0.V_err_gate.n1 two_stage_opamp_dummy_magic_16_0.V_err_gate.t4 15.7605
R8340 two_stage_opamp_dummy_magic_16_0.V_err_gate two_stage_opamp_dummy_magic_16_0.V_err_gate.n5 1.76612
R8341 two_stage_opamp_dummy_magic_16_0.V_err_gate.n5 two_stage_opamp_dummy_magic_16_0.V_err_gate.n3 0.641125
R8342 a_5980_2720.t0 a_5980_2720.t1 169.905
R8343 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t0 652.076
R8344 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t4 652.076
R8345 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n28 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n27 585
R8346 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n44 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n2 585
R8347 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n27 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n16 290.233
R8348 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n27 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n21 290.233
R8349 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n27 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n26 290.233
R8350 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n44 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n43 290.233
R8351 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n44 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n0 290.233
R8352 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n44 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n1 290.233
R8353 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n26 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n8 242.903
R8354 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n36 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n1 242.903
R8355 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n42 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n41 238.367
R8356 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n29 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n28 185
R8357 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n30 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n29 185
R8358 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n9 185
R8359 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n17 185
R8360 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n20 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n19 185
R8361 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n23 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n22 185
R8362 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n25 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n24 185
R8363 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n3 185
R8364 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n39 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n2 185
R8365 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n40 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n39 185
R8366 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n38 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n37 185
R8367 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n33 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n32 185
R8368 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n35 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n34 185
R8369 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n30 170.513
R8370 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n40 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t1 170.513
R8371 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n10 169.694
R8372 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n11 155.303
R8373 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n39 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n5 150
R8374 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n39 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n38 150
R8375 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n35 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n32 150
R8376 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n29 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n9 150
R8377 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n19 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n18 150
R8378 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n24 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n23 150
R8379 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t9 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t5 146.155
R8380 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t9 146.155
R8381 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n30 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n6 65.8183
R8382 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n30 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n7 65.8183
R8383 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n30 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n8 65.8183
R8384 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n41 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n40 65.8183
R8385 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n40 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n31 65.8183
R8386 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n40 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n36 65.8183
R8387 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n38 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n31 53.3664
R8388 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n36 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n35 53.3664
R8389 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n6 53.3664
R8390 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n19 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n7 53.3664
R8391 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n24 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n8 53.3664
R8392 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n6 53.3664
R8393 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n23 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n7 53.3664
R8394 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n41 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n5 53.3664
R8395 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n32 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n31 53.3664
R8396 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n28 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n14 22.8576
R8397 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n42 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n4 22.8576
R8398 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n13 14.4255
R8399 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n4 14.0505
R8400 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t10 11.2576
R8401 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t2 11.2576
R8402 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t7 11.2576
R8403 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t8 11.2576
R8404 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n27 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t6 11.2576
R8405 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n44 11.2576
R8406 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n28 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n15 9.14336
R8407 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n20 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n17 9.14336
R8408 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n25 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n22 9.14336
R8409 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n2 9.14336
R8410 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n37 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n2 9.14336
R8411 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n34 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n33 9.14336
R8412 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n15 4.53698
R8413 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n21 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n20 4.53698
R8414 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n26 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n25 4.53698
R8415 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n16 4.53698
R8416 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n22 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n21 4.53698
R8417 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n43 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n42 4.53698
R8418 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n37 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n0 4.53698
R8419 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n34 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n1 4.53698
R8420 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n43 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n3 4.53698
R8421 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n33 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n0 4.53698
R8422 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_16_0.Vb2_Vb3.n12 4.5005
R8423 two_stage_opamp_dummy_magic_16_0.V_err_mir_p two_stage_opamp_dummy_magic_16_0.V_err_mir_p.n0 187.315
R8424 two_stage_opamp_dummy_magic_16_0.V_err_mir_p two_stage_opamp_dummy_magic_16_0.V_err_mir_p.n1 177.755
R8425 two_stage_opamp_dummy_magic_16_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_16_0.V_err_mir_p.t3 15.7605
R8426 two_stage_opamp_dummy_magic_16_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_16_0.V_err_mir_p.t0 15.7605
R8427 two_stage_opamp_dummy_magic_16_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_16_0.V_err_mir_p.t1 15.7605
R8428 two_stage_opamp_dummy_magic_16_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_16_0.V_err_mir_p.t2 15.7605
R8429 a_14010_2720.t0 a_14010_2720.t1 169.905
R8430 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n0 344.837
R8431 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n1 344.274
R8432 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n3 292.5
R8433 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n5 209.251
R8434 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n12 208.689
R8435 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n10 208.689
R8436 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n8 208.689
R8437 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n6 208.689
R8438 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t16 120.305
R8439 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n2 52.3363
R8440 bgr_0.V_CMFB_S1 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n4 52.1563
R8441 bgr_0.V_CMFB_S1 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n14 50.813
R8442 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t11 39.4005
R8443 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t14 39.4005
R8444 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t10 39.4005
R8445 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t13 39.4005
R8446 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t15 39.4005
R8447 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t12 39.4005
R8448 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t4 19.7005
R8449 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t8 19.7005
R8450 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t3 19.7005
R8451 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t7 19.7005
R8452 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t2 19.7005
R8453 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t6 19.7005
R8454 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t0 19.7005
R8455 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t9 19.7005
R8456 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t1 19.7005
R8457 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t5 19.7005
R8458 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n13 5.90675
R8459 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n7 0.563
R8460 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n9 0.563
R8461 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n11 0.563
R8462 bgr_0.START_UP_NFET1 bgr_0.START_UP_NFET1.t0 141.653
R8463 VIN-.n1 VIN-.t4 478.096
R8464 VIN-.n5 VIN-.t5 477.303
R8465 VIN-.n4 VIN-.t6 477.303
R8466 VIN-.n8 VIN-.t8 436.36
R8467 VIN-.n2 VIN-.t7 436.36
R8468 VIN-.n6 VIN-.t10 435.382
R8469 VIN-.n0 VIN-.t9 435.382
R8470 VIN-.n6 VIN-.t0 284.24
R8471 VIN-.n0 VIN-.t3 284.24
R8472 VIN-.n8 VIN-.t2 274.106
R8473 VIN-.n2 VIN-.t1 274.106
R8474 VIN-.n7 VIN-.n6 237.055
R8475 VIN-.n1 VIN-.n0 237.055
R8476 VIN-.n9 VIN-.n8 189.309
R8477 VIN-.n3 VIN-.n2 189.309
R8478 VIN-.n4 VIN-.n3 2.46925
R8479 VIN-.n5 VIN-.n4 1.58175
R8480 VIN- VIN-.n9 1.44737
R8481 VIN-.n3 VIN-.n1 1.28175
R8482 VIN-.n9 VIN-.n7 1.28175
R8483 VIN-.n7 VIN-.n5 0.79425
R8484 a_12530_23988.t0 a_12530_23988.t1 178.133
R8485 two_stage_opamp_dummy_magic_16_0.V_p_mir.n1 two_stage_opamp_dummy_magic_16_0.V_p_mir.n0 223.127
R8486 two_stage_opamp_dummy_magic_16_0.V_p_mir.n0 two_stage_opamp_dummy_magic_16_0.V_p_mir.t3 16.0005
R8487 two_stage_opamp_dummy_magic_16_0.V_p_mir.n0 two_stage_opamp_dummy_magic_16_0.V_p_mir.t0 16.0005
R8488 two_stage_opamp_dummy_magic_16_0.V_p_mir.n1 two_stage_opamp_dummy_magic_16_0.V_p_mir.t1 9.6005
R8489 two_stage_opamp_dummy_magic_16_0.V_p_mir.t2 two_stage_opamp_dummy_magic_16_0.V_p_mir.n1 9.6005
R8490 a_7580_22380.t0 a_7580_22380.t1 178.133
R8491 a_5700_5524.t0 a_5700_5524.t1 169.905
R8492 two_stage_opamp_dummy_magic_16_0.V_tot.n2 two_stage_opamp_dummy_magic_16_0.V_tot.t4 648.25
R8493 two_stage_opamp_dummy_magic_16_0.V_tot.n1 two_stage_opamp_dummy_magic_16_0.V_tot.t5 648.25
R8494 two_stage_opamp_dummy_magic_16_0.V_tot.t0 two_stage_opamp_dummy_magic_16_0.V_tot.n3 116.546
R8495 two_stage_opamp_dummy_magic_16_0.V_tot.n0 two_stage_opamp_dummy_magic_16_0.V_tot.t2 116.546
R8496 two_stage_opamp_dummy_magic_16_0.V_tot.n3 two_stage_opamp_dummy_magic_16_0.V_tot.t3 107.328
R8497 two_stage_opamp_dummy_magic_16_0.V_tot.n0 two_stage_opamp_dummy_magic_16_0.V_tot.t1 107.328
R8498 two_stage_opamp_dummy_magic_16_0.V_tot.n1 two_stage_opamp_dummy_magic_16_0.V_tot.n0 34.9431
R8499 two_stage_opamp_dummy_magic_16_0.V_tot.n3 two_stage_opamp_dummy_magic_16_0.V_tot.n2 34.8494
R8500 two_stage_opamp_dummy_magic_16_0.V_tot.n2 two_stage_opamp_dummy_magic_16_0.V_tot.n1 1.563
R8501 a_6810_23838.t0 a_6810_23838.t1 178.133
R8502 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 195.608
R8503 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 83.5719
R8504 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 83.5719
R8505 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 83.5719
R8506 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 83.5719
R8507 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 83.5719
R8508 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 83.5719
R8509 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 83.5719
R8510 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 83.5719
R8511 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 83.5719
R8512 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 83.5719
R8513 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 83.5719
R8514 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 83.5719
R8515 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 83.5719
R8516 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 83.5719
R8517 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 83.5719
R8518 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 83.5719
R8519 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 83.5719
R8520 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 83.5719
R8521 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 83.5719
R8522 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 83.5719
R8523 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R8524 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 83.5719
R8525 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 73.8495
R8526 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 73.8495
R8527 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 73.3165
R8528 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 73.3165
R8529 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 73.3165
R8530 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 73.3165
R8531 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 73.3165
R8532 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 73.3165
R8533 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 73.19
R8534 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 73.19
R8535 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 73.19
R8536 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 73.19
R8537 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 73.19
R8538 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 73.19
R8539 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 65.0299
R8540 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 65.0299
R8541 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 26.074
R8542 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 26.074
R8543 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 26.074
R8544 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 26.074
R8545 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 26.074
R8546 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 26.074
R8547 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 26.074
R8548 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 26.074
R8549 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 25.7843
R8550 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 25.7843
R8551 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 25.7843
R8552 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 25.7843
R8553 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 25.7843
R8554 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 25.7843
R8555 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R8556 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R8557 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8558 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R8559 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R8560 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8561 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R8562 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 9.3005
R8563 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R8564 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R8565 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8566 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R8567 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 9.3005
R8568 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 9.3005
R8569 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R8570 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8571 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R8572 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R8573 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R8574 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8575 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R8576 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R8577 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R8578 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R8579 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8580 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 9.3005
R8581 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 9.3005
R8582 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 9.3005
R8583 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8584 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8585 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8586 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 9.3005
R8587 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8588 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8589 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8590 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 9.3005
R8591 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8592 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8593 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R8594 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8595 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8596 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R8597 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8598 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8599 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8600 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R8601 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8602 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8603 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 9.3005
R8604 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 9.3005
R8605 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8606 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8607 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R8608 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8609 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 4.64654
R8610 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 4.64654
R8611 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 4.64654
R8612 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 4.64654
R8613 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 4.64654
R8614 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 4.64654
R8615 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 4.64654
R8616 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 4.64654
R8617 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 4.64654
R8618 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 2.36206
R8619 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 2.36206
R8620 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 2.36206
R8621 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 2.36206
R8622 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 2.19742
R8623 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 2.19742
R8624 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 2.19742
R8625 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 2.19742
R8626 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 1.56363
R8627 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.56363
R8628 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 1.5505
R8629 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R8630 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 1.5505
R8631 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 1.5505
R8632 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 1.5505
R8633 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 1.5505
R8634 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 1.5505
R8635 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 1.5505
R8636 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 1.5505
R8637 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 1.5505
R8638 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 1.5505
R8639 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 1.5505
R8640 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 1.5505
R8641 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 1.5505
R8642 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 1.5505
R8643 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 1.5505
R8644 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 1.5505
R8645 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 1.5505
R8646 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.25468
R8647 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 1.25468
R8648 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.25468
R8649 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.25468
R8650 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 1.25468
R8651 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 1.25468
R8652 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 1.19225
R8653 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 1.19225
R8654 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 1.19225
R8655 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 1.19225
R8656 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 1.19225
R8657 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.19225
R8658 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 1.07024
R8659 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 1.07024
R8660 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 1.07024
R8661 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 1.07024
R8662 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 1.07024
R8663 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.07024
R8664 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.0237
R8665 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 1.0237
R8666 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.0237
R8667 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.0237
R8668 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 1.0237
R8669 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 1.0237
R8670 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.885803
R8671 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 0.885803
R8672 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 0.885803
R8673 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 0.885803
R8674 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.885803
R8675 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.885803
R8676 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 0.885803
R8677 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.885803
R8678 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 0.812055
R8679 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 0.812055
R8680 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.77514
R8681 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.77514
R8682 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 0.77514
R8683 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.77514
R8684 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.77514
R8685 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 0.77514
R8686 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 0.77514
R8687 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 0.77514
R8688 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.756696
R8689 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R8690 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.756696
R8691 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 0.756696
R8692 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R8693 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.756696
R8694 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R8695 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.756696
R8696 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 0.711459
R8697 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.711459
R8698 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.647417
R8699 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 0.647417
R8700 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.590702
R8701 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 0.590702
R8702 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.590702
R8703 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 0.590702
R8704 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.590702
R8705 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 0.590702
R8706 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.576566
R8707 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.576566
R8708 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 0.530034
R8709 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 0.530034
R8710 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 0.290206
R8711 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 0.290206
R8712 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 0.290206
R8713 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 0.290206
R8714 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 0.290206
R8715 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 0.290206
R8716 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 0.290206
R8717 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 0.290206
R8718 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8719 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8720 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8721 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.203382
R8722 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8723 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 0.203382
R8724 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 0.154071
R8725 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 0.154071
R8726 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 0.154071
R8727 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 0.154071
R8728 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 0.137464
R8729 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 0.137464
R8730 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 0.134964
R8731 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 0.134964
R8732 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R8733 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 0.0183571
R8734 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R8735 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R8736 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 0.0183571
R8737 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R8738 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R8739 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 0.0183571
R8740 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0183571
R8741 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R8742 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R8743 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R8744 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R8745 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 0.0183571
R8746 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R8747 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R8748 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 0.0183571
R8749 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0183571
R8750 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0106786
R8751 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0106786
R8752 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.0106786
R8753 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 0.00992001
R8754 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 0.00992001
R8755 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R8756 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 0.00992001
R8757 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R8758 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R8759 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R8760 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 0.00992001
R8761 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 0.00992001
R8762 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 0.00992001
R8763 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R8764 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 0.00992001
R8765 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R8766 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R8767 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R8768 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R8769 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 0.00992001
R8770 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R8771 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.00817857
R8772 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00817857
R8773 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 0.00817857
R8774 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 0.00817857
R8775 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.00817857
R8776 two_stage_opamp_dummy_magic_16_0.err_amp_out two_stage_opamp_dummy_magic_16_0.err_amp_out.t4 682.663
R8777 two_stage_opamp_dummy_magic_16_0.err_amp_out.n2 two_stage_opamp_dummy_magic_16_0.err_amp_out.n1 179.226
R8778 two_stage_opamp_dummy_magic_16_0.err_amp_out.n2 two_stage_opamp_dummy_magic_16_0.err_amp_out.n0 100.382
R8779 two_stage_opamp_dummy_magic_16_0.err_amp_out.n1 two_stage_opamp_dummy_magic_16_0.err_amp_out.t3 15.7605
R8780 two_stage_opamp_dummy_magic_16_0.err_amp_out.n1 two_stage_opamp_dummy_magic_16_0.err_amp_out.t1 15.7605
R8781 two_stage_opamp_dummy_magic_16_0.err_amp_out.n0 two_stage_opamp_dummy_magic_16_0.err_amp_out.t0 9.6005
R8782 two_stage_opamp_dummy_magic_16_0.err_amp_out.n0 two_stage_opamp_dummy_magic_16_0.err_amp_out.t2 9.6005
R8783 two_stage_opamp_dummy_magic_16_0.err_amp_out two_stage_opamp_dummy_magic_16_0.err_amp_out.n2 0.922375
R8784 a_5580_5524.t0 a_5580_5524.t1 262.248
R8785 a_12410_22380.t0 a_12410_22380.t1 178.133
R8786 a_13060_22630.t0 a_13060_22630.t1 178.133
R8787 two_stage_opamp_dummy_magic_16_0.V_err_p.n1 two_stage_opamp_dummy_magic_16_0.V_err_p.n0 365.07
R8788 two_stage_opamp_dummy_magic_16_0.V_err_p.n0 two_stage_opamp_dummy_magic_16_0.V_err_p.t0 15.7605
R8789 two_stage_opamp_dummy_magic_16_0.V_err_p.n0 two_stage_opamp_dummy_magic_16_0.V_err_p.t2 15.7605
R8790 two_stage_opamp_dummy_magic_16_0.V_err_p.n1 two_stage_opamp_dummy_magic_16_0.V_err_p.t3 15.7605
R8791 two_stage_opamp_dummy_magic_16_0.V_err_p.t1 two_stage_opamp_dummy_magic_16_0.V_err_p.n1 15.7605
R8792 two_stage_opamp_dummy_magic_16_0.Vb2_2.n32 two_stage_opamp_dummy_magic_16_0.Vb2_2.n31 692.967
R8793 two_stage_opamp_dummy_magic_16_0.Vb2_2.n34 two_stage_opamp_dummy_magic_16_0.Vb2_2.t0 652.076
R8794 two_stage_opamp_dummy_magic_16_0.Vb2_2.n30 two_stage_opamp_dummy_magic_16_0.Vb2_2.t3 652.076
R8795 two_stage_opamp_dummy_magic_16_0.Vb2_2.n36 two_stage_opamp_dummy_magic_16_0.Vb2_2.n0 587.407
R8796 two_stage_opamp_dummy_magic_16_0.Vb2_2.n41 two_stage_opamp_dummy_magic_16_0.Vb2_2.n2 587.407
R8797 two_stage_opamp_dummy_magic_16_0.Vb2_2.n29 two_stage_opamp_dummy_magic_16_0.Vb2_2.n11 585
R8798 two_stage_opamp_dummy_magic_16_0.Vb2_2.n3 two_stage_opamp_dummy_magic_16_0.Vb2_2.n0 585
R8799 two_stage_opamp_dummy_magic_16_0.Vb2_2.t2 two_stage_opamp_dummy_magic_16_0.Vb2_2.n44 585
R8800 two_stage_opamp_dummy_magic_16_0.Vb2_2.n43 two_stage_opamp_dummy_magic_16_0.Vb2_2.n2 585
R8801 two_stage_opamp_dummy_magic_16_0.Vb2_2.n17 two_stage_opamp_dummy_magic_16_0.Vb2_2.n11 290.233
R8802 two_stage_opamp_dummy_magic_16_0.Vb2_2.n23 two_stage_opamp_dummy_magic_16_0.Vb2_2.n11 290.233
R8803 two_stage_opamp_dummy_magic_16_0.Vb2_2.n18 two_stage_opamp_dummy_magic_16_0.Vb2_2.n11 290.233
R8804 two_stage_opamp_dummy_magic_16_0.Vb2_2.t2 two_stage_opamp_dummy_magic_16_0.Vb2_2.n0 246.25
R8805 two_stage_opamp_dummy_magic_16_0.Vb2_2.t2 two_stage_opamp_dummy_magic_16_0.Vb2_2.n2 246.25
R8806 two_stage_opamp_dummy_magic_16_0.Vb2_2.n41 two_stage_opamp_dummy_magic_16_0.Vb2_2.n40 243.698
R8807 two_stage_opamp_dummy_magic_16_0.Vb2_2.n18 two_stage_opamp_dummy_magic_16_0.Vb2_2.n15 242.903
R8808 two_stage_opamp_dummy_magic_16_0.Vb2_2.n29 two_stage_opamp_dummy_magic_16_0.Vb2_2.n28 238.367
R8809 two_stage_opamp_dummy_magic_16_0.Vb2_2.n13 two_stage_opamp_dummy_magic_16_0.Vb2_2.n12 185
R8810 two_stage_opamp_dummy_magic_16_0.Vb2_2.n26 two_stage_opamp_dummy_magic_16_0.Vb2_2.n25 185
R8811 two_stage_opamp_dummy_magic_16_0.Vb2_2.n27 two_stage_opamp_dummy_magic_16_0.Vb2_2.n26 185
R8812 two_stage_opamp_dummy_magic_16_0.Vb2_2.n24 two_stage_opamp_dummy_magic_16_0.Vb2_2.n16 185
R8813 two_stage_opamp_dummy_magic_16_0.Vb2_2.n22 two_stage_opamp_dummy_magic_16_0.Vb2_2.n21 185
R8814 two_stage_opamp_dummy_magic_16_0.Vb2_2.n20 two_stage_opamp_dummy_magic_16_0.Vb2_2.n19 185
R8815 two_stage_opamp_dummy_magic_16_0.Vb2_2.n38 two_stage_opamp_dummy_magic_16_0.Vb2_2.n37 185
R8816 two_stage_opamp_dummy_magic_16_0.Vb2_2.n39 two_stage_opamp_dummy_magic_16_0.Vb2_2.n38 185
R8817 two_stage_opamp_dummy_magic_16_0.Vb2_2.n35 two_stage_opamp_dummy_magic_16_0.Vb2_2.n10 185
R8818 two_stage_opamp_dummy_magic_16_0.Vb2_2.n7 two_stage_opamp_dummy_magic_16_0.Vb2_2.n3 185
R8819 two_stage_opamp_dummy_magic_16_0.Vb2_2.n44 two_stage_opamp_dummy_magic_16_0.Vb2_2.n4 185
R8820 two_stage_opamp_dummy_magic_16_0.Vb2_2.n43 two_stage_opamp_dummy_magic_16_0.Vb2_2.n5 185
R8821 two_stage_opamp_dummy_magic_16_0.Vb2_2.n42 two_stage_opamp_dummy_magic_16_0.Vb2_2.n6 185
R8822 two_stage_opamp_dummy_magic_16_0.Vb2_2.n39 two_stage_opamp_dummy_magic_16_0.Vb2_2.t1 170.513
R8823 two_stage_opamp_dummy_magic_16_0.Vb2_2.n27 two_stage_opamp_dummy_magic_16_0.Vb2_2.t4 170.513
R8824 two_stage_opamp_dummy_magic_16_0.Vb2_2.n32 two_stage_opamp_dummy_magic_16_0.Vb2_2.n1 155.304
R8825 two_stage_opamp_dummy_magic_16_0.Vb2_2.n26 two_stage_opamp_dummy_magic_16_0.Vb2_2.n13 150
R8826 two_stage_opamp_dummy_magic_16_0.Vb2_2.n26 two_stage_opamp_dummy_magic_16_0.Vb2_2.n16 150
R8827 two_stage_opamp_dummy_magic_16_0.Vb2_2.n21 two_stage_opamp_dummy_magic_16_0.Vb2_2.n20 150
R8828 two_stage_opamp_dummy_magic_16_0.Vb2_2.n38 two_stage_opamp_dummy_magic_16_0.Vb2_2.n10 150
R8829 two_stage_opamp_dummy_magic_16_0.Vb2_2.n7 two_stage_opamp_dummy_magic_16_0.Vb2_2.n4 150
R8830 two_stage_opamp_dummy_magic_16_0.Vb2_2.n6 two_stage_opamp_dummy_magic_16_0.Vb2_2.n5 150
R8831 two_stage_opamp_dummy_magic_16_0.Vb2_2.t7 two_stage_opamp_dummy_magic_16_0.Vb2_2.t1 146.155
R8832 two_stage_opamp_dummy_magic_16_0.Vb2_2.t4 two_stage_opamp_dummy_magic_16_0.Vb2_2.t7 146.155
R8833 two_stage_opamp_dummy_magic_16_0.Vb2_2.n28 two_stage_opamp_dummy_magic_16_0.Vb2_2.n27 65.8183
R8834 two_stage_opamp_dummy_magic_16_0.Vb2_2.n27 two_stage_opamp_dummy_magic_16_0.Vb2_2.n14 65.8183
R8835 two_stage_opamp_dummy_magic_16_0.Vb2_2.n27 two_stage_opamp_dummy_magic_16_0.Vb2_2.n15 65.8183
R8836 two_stage_opamp_dummy_magic_16_0.Vb2_2.n39 two_stage_opamp_dummy_magic_16_0.Vb2_2.n8 65.8183
R8837 two_stage_opamp_dummy_magic_16_0.Vb2_2.n39 two_stage_opamp_dummy_magic_16_0.Vb2_2.n9 65.8183
R8838 two_stage_opamp_dummy_magic_16_0.Vb2_2.n40 two_stage_opamp_dummy_magic_16_0.Vb2_2.n39 65.8183
R8839 two_stage_opamp_dummy_magic_16_0.Vb2_2.n16 two_stage_opamp_dummy_magic_16_0.Vb2_2.n14 53.3664
R8840 two_stage_opamp_dummy_magic_16_0.Vb2_2.n20 two_stage_opamp_dummy_magic_16_0.Vb2_2.n15 53.3664
R8841 two_stage_opamp_dummy_magic_16_0.Vb2_2.n28 two_stage_opamp_dummy_magic_16_0.Vb2_2.n13 53.3664
R8842 two_stage_opamp_dummy_magic_16_0.Vb2_2.n21 two_stage_opamp_dummy_magic_16_0.Vb2_2.n14 53.3664
R8843 two_stage_opamp_dummy_magic_16_0.Vb2_2.n10 two_stage_opamp_dummy_magic_16_0.Vb2_2.n8 53.3664
R8844 two_stage_opamp_dummy_magic_16_0.Vb2_2.n9 two_stage_opamp_dummy_magic_16_0.Vb2_2.n4 53.3664
R8845 two_stage_opamp_dummy_magic_16_0.Vb2_2.n40 two_stage_opamp_dummy_magic_16_0.Vb2_2.n6 53.3664
R8846 two_stage_opamp_dummy_magic_16_0.Vb2_2.n8 two_stage_opamp_dummy_magic_16_0.Vb2_2.n7 53.3664
R8847 two_stage_opamp_dummy_magic_16_0.Vb2_2.n9 two_stage_opamp_dummy_magic_16_0.Vb2_2.n5 53.3664
R8848 two_stage_opamp_dummy_magic_16_0.Vb2_2.n30 two_stage_opamp_dummy_magic_16_0.Vb2_2.n29 22.8576
R8849 two_stage_opamp_dummy_magic_16_0.Vb2_2.n37 two_stage_opamp_dummy_magic_16_0.Vb2_2.n34 22.8576
R8850 two_stage_opamp_dummy_magic_16_0.Vb2_2.n31 two_stage_opamp_dummy_magic_16_0.Vb2_2.t6 21.8894
R8851 two_stage_opamp_dummy_magic_16_0.Vb2_2.n31 two_stage_opamp_dummy_magic_16_0.Vb2_2.t9 21.8894
R8852 two_stage_opamp_dummy_magic_16_0.Vb2_2.n33 two_stage_opamp_dummy_magic_16_0.Vb2_2.n30 14.4255
R8853 two_stage_opamp_dummy_magic_16_0.Vb2_2.n34 two_stage_opamp_dummy_magic_16_0.Vb2_2.n33 14.0505
R8854 two_stage_opamp_dummy_magic_16_0.Vb2_2.n11 two_stage_opamp_dummy_magic_16_0.Vb2_2.t5 11.2576
R8855 two_stage_opamp_dummy_magic_16_0.Vb2_2.t2 two_stage_opamp_dummy_magic_16_0.Vb2_2.n1 11.2576
R8856 two_stage_opamp_dummy_magic_16_0.Vb2_2.n1 two_stage_opamp_dummy_magic_16_0.Vb2_2.t8 11.2576
R8857 two_stage_opamp_dummy_magic_16_0.Vb2_2.n29 two_stage_opamp_dummy_magic_16_0.Vb2_2.n12 9.14336
R8858 two_stage_opamp_dummy_magic_16_0.Vb2_2.n25 two_stage_opamp_dummy_magic_16_0.Vb2_2.n24 9.14336
R8859 two_stage_opamp_dummy_magic_16_0.Vb2_2.n22 two_stage_opamp_dummy_magic_16_0.Vb2_2.n19 9.14336
R8860 two_stage_opamp_dummy_magic_16_0.Vb2_2.n35 two_stage_opamp_dummy_magic_16_0.Vb2_2.n3 9.14336
R8861 two_stage_opamp_dummy_magic_16_0.Vb2_2.n44 two_stage_opamp_dummy_magic_16_0.Vb2_2.n3 9.14336
R8862 two_stage_opamp_dummy_magic_16_0.Vb2_2.n44 two_stage_opamp_dummy_magic_16_0.Vb2_2.n43 9.14336
R8863 two_stage_opamp_dummy_magic_16_0.Vb2_2.n43 two_stage_opamp_dummy_magic_16_0.Vb2_2.n42 9.14336
R8864 two_stage_opamp_dummy_magic_16_0.Vb2_2.n37 two_stage_opamp_dummy_magic_16_0.Vb2_2.n36 5.33286
R8865 two_stage_opamp_dummy_magic_16_0.Vb2_2.n17 two_stage_opamp_dummy_magic_16_0.Vb2_2.n12 4.53698
R8866 two_stage_opamp_dummy_magic_16_0.Vb2_2.n24 two_stage_opamp_dummy_magic_16_0.Vb2_2.n23 4.53698
R8867 two_stage_opamp_dummy_magic_16_0.Vb2_2.n19 two_stage_opamp_dummy_magic_16_0.Vb2_2.n18 4.53698
R8868 two_stage_opamp_dummy_magic_16_0.Vb2_2.n25 two_stage_opamp_dummy_magic_16_0.Vb2_2.n17 4.53698
R8869 two_stage_opamp_dummy_magic_16_0.Vb2_2.n23 two_stage_opamp_dummy_magic_16_0.Vb2_2.n22 4.53698
R8870 two_stage_opamp_dummy_magic_16_0.Vb2_2.n33 two_stage_opamp_dummy_magic_16_0.Vb2_2.n32 4.5005
R8871 two_stage_opamp_dummy_magic_16_0.Vb2_2.n36 two_stage_opamp_dummy_magic_16_0.Vb2_2.n35 3.75335
R8872 two_stage_opamp_dummy_magic_16_0.Vb2_2.n42 two_stage_opamp_dummy_magic_16_0.Vb2_2.n41 3.75335
R8873 a_13180_23838.t0 a_13180_23838.t1 178.133
R8874 a_14170_5524.t0 a_14170_5524.t1 298.82
R8875 a_14290_5524.t0 a_14290_5524.t1 169.905
C0 two_stage_opamp_dummy_magic_16_0.err_amp_out two_stage_opamp_dummy_magic_16_0.VD1 0.090652f
C1 bgr_0.1st_Vout_1 two_stage_opamp_dummy_magic_16_0.Vb2 0.042752f
C2 VOUT+ two_stage_opamp_dummy_magic_16_0.VD4 0.023279f
C3 bgr_0.NFET_GATE_10uA bgr_0.START_UP 1.64177f
C4 bgr_0.V_TOP two_stage_opamp_dummy_magic_16_0.V_err_amp_ref 0.583702f
C5 two_stage_opamp_dummy_magic_16_0.cap_res_X two_stage_opamp_dummy_magic_16_0.V_err_gate 0.333809f
C6 VDDA bgr_0.NFET_GATE_10uA 0.818988f
C7 VDDA two_stage_opamp_dummy_magic_16_0.V_err_gate 1.61292f
C8 bgr_0.V_TOP bgr_0.PFET_GATE_10uA 0.221314f
C9 VDDA bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.046803f
C10 VDDA bgr_0.START_UP 1.09181f
C11 VDDA two_stage_opamp_dummy_magic_16_0.cap_res_X 0.392458f
C12 m2_9370_16580# bgr_0.PFET_GATE_10uA 0.012f
C13 two_stage_opamp_dummy_magic_16_0.Vb2 two_stage_opamp_dummy_magic_16_0.VD4 1.23597f
C14 bgr_0.START_UP_NFET1 bgr_0.PFET_GATE_10uA 0.0108f
C15 m2_10730_16580# bgr_0.V_TOP 0.012f
C16 bgr_0.V_TOP bgr_0.NFET_GATE_10uA 0.052756f
C17 two_stage_opamp_dummy_magic_16_0.err_amp_out two_stage_opamp_dummy_magic_16_0.V_err_amp_ref 0.15972f
C18 VOUT+ two_stage_opamp_dummy_magic_16_0.cap_res_X 0.037134f
C19 bgr_0.V_TOP two_stage_opamp_dummy_magic_16_0.V_err_gate 0.08195f
C20 VOUT- two_stage_opamp_dummy_magic_16_0.V_err_gate 0.040291f
C21 m1_10050_19490# two_stage_opamp_dummy_magic_16_0.V_err_gate 0.091711f
C22 VDDA VOUT+ 5.84806f
C23 bgr_0.V_TOP bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.055802f
C24 bgr_0.V_TOP bgr_0.START_UP 0.792764f
C25 m1_4880_3600# m2_4880_3600# 0.016063f
C26 m1_10050_19490# bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.013969f
C27 VIN- VIN+ 0.562821f
C28 VOUT- two_stage_opamp_dummy_magic_16_0.cap_res_X 51.0174f
C29 two_stage_opamp_dummy_magic_16_0.VD4 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref 0.506178f
C30 VDDA bgr_0.V_TOP 13.2374f
C31 m2_10730_16580# bgr_0.1st_Vout_1 0.075543f
C32 VDDA VOUT- 5.85101f
C33 bgr_0.1st_Vout_1 bgr_0.NFET_GATE_10uA 0.03875f
C34 bgr_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_16_0.V_err_amp_ref 1.67032f
C35 bgr_0.1st_Vout_1 two_stage_opamp_dummy_magic_16_0.V_err_gate 0.041119f
C36 bgr_0.NFET_GATE_10uA bgr_0.START_UP_NFET1 0.351171f
C37 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_16_0.Vb2 0.538556f
C38 VIN- two_stage_opamp_dummy_magic_16_0.VD1 0.923907f
C39 two_stage_opamp_dummy_magic_16_0.V_err_mir_p two_stage_opamp_dummy_magic_16_0.V_err_amp_ref 0.047421f
C40 two_stage_opamp_dummy_magic_16_0.Vb2 two_stage_opamp_dummy_magic_16_0.V_err_gate 2.06899f
C41 bgr_0.1st_Vout_1 bgr_0.START_UP 0.04354f
C42 bgr_0.START_UP_NFET1 bgr_0.START_UP 0.145663f
C43 two_stage_opamp_dummy_magic_16_0.Vb2 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.01158f
C44 two_stage_opamp_dummy_magic_16_0.V_err_mir_p two_stage_opamp_dummy_magic_16_0.VD4 0.02057f
C45 two_stage_opamp_dummy_magic_16_0.Vb2 bgr_0.START_UP 0.08188f
C46 VDDA bgr_0.1st_Vout_1 0.896465f
C47 two_stage_opamp_dummy_magic_16_0.cap_res_X two_stage_opamp_dummy_magic_16_0.Vb2 0.615754f
C48 VIN+ two_stage_opamp_dummy_magic_16_0.VD1 0.051708f
C49 VDDA bgr_0.START_UP_NFET1 0.167059f
C50 VDDA two_stage_opamp_dummy_magic_16_0.Vb2 1.44365f
C51 VOUT+ VOUT- 0.397591f
C52 two_stage_opamp_dummy_magic_16_0.err_amp_out two_stage_opamp_dummy_magic_16_0.V_err_gate 0.055417f
C53 two_stage_opamp_dummy_magic_16_0.V_err_gate two_stage_opamp_dummy_magic_16_0.V_err_amp_ref 0.804479f
C54 VDDA two_stage_opamp_dummy_magic_16_0.err_amp_out 1.28767f
C55 bgr_0.START_UP two_stage_opamp_dummy_magic_16_0.V_err_amp_ref 1.36583f
C56 bgr_0.NFET_GATE_10uA bgr_0.PFET_GATE_10uA 0.012365f
C57 VDDA two_stage_opamp_dummy_magic_16_0.V_err_amp_ref 2.39922f
C58 two_stage_opamp_dummy_magic_16_0.V_err_mir_p two_stage_opamp_dummy_magic_16_0.V_err_gate 0.429395f
C59 VDDA two_stage_opamp_dummy_magic_16_0.VD4 4.39386f
C60 bgr_0.1st_Vout_1 bgr_0.V_TOP 2.47405f
C61 two_stage_opamp_dummy_magic_16_0.cap_res_X bgr_0.PFET_GATE_10uA 0.011459f
C62 VDDA bgr_0.PFET_GATE_10uA 7.97055f
C63 bgr_0.V_TOP two_stage_opamp_dummy_magic_16_0.Vb2 0.936691f
C64 VOUT- two_stage_opamp_dummy_magic_16_0.Vb2 0.058721f
C65 m1_10050_19490# two_stage_opamp_dummy_magic_16_0.Vb2 0.08176f
C66 VDDA two_stage_opamp_dummy_magic_16_0.V_err_mir_p 0.671539f
C67 VOUT+ two_stage_opamp_dummy_magic_16_0.V_err_amp_ref 0.042091f
C68 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_16_0.V_err_gate 3.50895f
C69 VIN+ GNDA 1.93244f
C70 VIN- GNDA 1.76634f
C71 VOUT- GNDA 15.859632f
C72 VOUT+ GNDA 15.896068f
C73 VDDA GNDA 0.120996p
C74 m2_4880_3600# GNDA 0.05269f $ **FLOATING
C75 m2_10730_16580# GNDA 0.0105f $ **FLOATING
C76 m2_9370_16580# GNDA 0.010002f $ **FLOATING
C77 m1_4880_3600# GNDA 0.059696f $ **FLOATING
C78 m1_10050_19490# GNDA 0.259273f $ **FLOATING
C79 two_stage_opamp_dummy_magic_16_0.VD1 GNDA 2.58052f
C80 two_stage_opamp_dummy_magic_16_0.cap_res_X GNDA 33.038033f
C81 two_stage_opamp_dummy_magic_16_0.err_amp_out GNDA 2.90043f
C82 two_stage_opamp_dummy_magic_16_0.V_err_mir_p GNDA 0.098443f
C83 bgr_0.1st_Vout_1 GNDA 7.823503f
C84 bgr_0.START_UP GNDA 5.877827f
C85 bgr_0.START_UP_NFET1 GNDA 4.29564f
C86 two_stage_opamp_dummy_magic_16_0.V_err_gate GNDA 7.797309f
C87 two_stage_opamp_dummy_magic_16_0.Vb2 GNDA 7.393193f
C88 bgr_0.NFET_GATE_10uA GNDA 7.92412f
C89 bgr_0.V_TOP GNDA 9.96016f
C90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA 17.8955f
C91 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref GNDA 6.835193f
C92 bgr_0.PFET_GATE_10uA GNDA 6.602193f
C93 two_stage_opamp_dummy_magic_16_0.VD4 GNDA 4.888278f
C94 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t15 GNDA 0.01637f
C95 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t12 GNDA 0.01637f
C96 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n0 GNDA 0.041034f
C97 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t10 GNDA 0.01637f
C98 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t13 GNDA 0.01637f
C99 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n1 GNDA 0.040818f
C100 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n2 GNDA 0.362787f
C101 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t11 GNDA 0.01637f
C102 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t14 GNDA 0.01637f
C103 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n3 GNDA 0.03274f
C104 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n4 GNDA 0.060887f
C105 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t16 GNDA 0.206157f
C106 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t1 GNDA 0.03274f
C107 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t5 GNDA 0.03274f
C108 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n5 GNDA 0.097293f
C109 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t0 GNDA 0.03274f
C110 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t9 GNDA 0.03274f
C111 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n6 GNDA 0.096862f
C112 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n7 GNDA 0.331325f
C113 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t2 GNDA 0.03274f
C114 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t6 GNDA 0.03274f
C115 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n8 GNDA 0.096862f
C116 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n9 GNDA 0.171607f
C117 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t3 GNDA 0.03274f
C118 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t7 GNDA 0.03274f
C119 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n10 GNDA 0.096862f
C120 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n11 GNDA 0.171607f
C121 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t4 GNDA 0.03274f
C122 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.t8 GNDA 0.03274f
C123 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n12 GNDA 0.096862f
C124 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n13 GNDA 0.239231f
C125 two_stage_opamp_dummy_magic_16_0.V_CMFB_S1.n14 GNDA 1.32734f
C126 bgr_0.V_CMFB_S1 GNDA 1.1041f
C127 two_stage_opamp_dummy_magic_16_0.V_err_gate.t1 GNDA 0.019165f
C128 two_stage_opamp_dummy_magic_16_0.V_err_gate.t2 GNDA 0.019165f
C129 two_stage_opamp_dummy_magic_16_0.V_err_gate.n0 GNDA 0.291418f
C130 two_stage_opamp_dummy_magic_16_0.V_err_gate.t0 GNDA 0.047912f
C131 two_stage_opamp_dummy_magic_16_0.V_err_gate.t4 GNDA 0.047912f
C132 two_stage_opamp_dummy_magic_16_0.V_err_gate.n1 GNDA 0.14679f
C133 two_stage_opamp_dummy_magic_16_0.V_err_gate.t8 GNDA 0.053502f
C134 two_stage_opamp_dummy_magic_16_0.V_err_gate.t6 GNDA 0.053502f
C135 two_stage_opamp_dummy_magic_16_0.V_err_gate.n2 GNDA 0.080364f
C136 two_stage_opamp_dummy_magic_16_0.V_err_gate.n3 GNDA 0.296603f
C137 two_stage_opamp_dummy_magic_16_0.V_err_gate.t3 GNDA 0.047912f
C138 two_stage_opamp_dummy_magic_16_0.V_err_gate.t5 GNDA 0.047912f
C139 two_stage_opamp_dummy_magic_16_0.V_err_gate.n4 GNDA 0.146154f
C140 two_stage_opamp_dummy_magic_16_0.V_err_gate.n5 GNDA 0.226942f
C141 two_stage_opamp_dummy_magic_16_0.V_err_gate.t7 GNDA 0.053502f
C142 two_stage_opamp_dummy_magic_16_0.V_err_gate.t9 GNDA 0.053502f
C143 two_stage_opamp_dummy_magic_16_0.V_err_gate.n6 GNDA 0.080364f
C144 bgr_0.START_UP.t0 GNDA 1.06745f
C145 bgr_0.START_UP.t1 GNDA 0.02806f
C146 bgr_0.START_UP.n0 GNDA 0.714928f
C147 bgr_0.START_UP.t2 GNDA 0.026778f
C148 bgr_0.START_UP.t4 GNDA 0.026778f
C149 bgr_0.START_UP.n1 GNDA 0.097147f
C150 bgr_0.START_UP.t3 GNDA 0.026778f
C151 bgr_0.START_UP.t5 GNDA 0.026778f
C152 bgr_0.START_UP.n2 GNDA 0.08937f
C153 bgr_0.START_UP.n3 GNDA 0.462855f
C154 bgr_0.START_UP.t7 GNDA 0.010062f
C155 bgr_0.START_UP.t6 GNDA 0.010062f
C156 bgr_0.START_UP.n4 GNDA 0.028407f
C157 bgr_0.START_UP.n5 GNDA 0.260836f
C158 two_stage_opamp_dummy_magic_16_0.VD4.t8 GNDA 0.030951f
C159 two_stage_opamp_dummy_magic_16_0.VD4.t11 GNDA 0.030951f
C160 two_stage_opamp_dummy_magic_16_0.VD4.n0 GNDA 0.108702f
C161 two_stage_opamp_dummy_magic_16_0.VD4.t3 GNDA 0.030951f
C162 two_stage_opamp_dummy_magic_16_0.VD4.t6 GNDA 0.030951f
C163 two_stage_opamp_dummy_magic_16_0.VD4.n1 GNDA 0.108329f
C164 two_stage_opamp_dummy_magic_16_0.VD4.n2 GNDA 0.202138f
C165 two_stage_opamp_dummy_magic_16_0.VD4.t1 GNDA 0.030951f
C166 two_stage_opamp_dummy_magic_16_0.VD4.t0 GNDA 0.030951f
C167 two_stage_opamp_dummy_magic_16_0.VD4.n3 GNDA 0.108329f
C168 two_stage_opamp_dummy_magic_16_0.VD4.n4 GNDA 0.104793f
C169 two_stage_opamp_dummy_magic_16_0.VD4.t7 GNDA 0.030951f
C170 two_stage_opamp_dummy_magic_16_0.VD4.t9 GNDA 0.030951f
C171 two_stage_opamp_dummy_magic_16_0.VD4.n5 GNDA 0.108329f
C172 two_stage_opamp_dummy_magic_16_0.VD4.n6 GNDA 0.104793f
C173 two_stage_opamp_dummy_magic_16_0.VD4.t2 GNDA 0.030951f
C174 two_stage_opamp_dummy_magic_16_0.VD4.t5 GNDA 0.030951f
C175 two_stage_opamp_dummy_magic_16_0.VD4.n7 GNDA 0.108329f
C176 two_stage_opamp_dummy_magic_16_0.VD4.n8 GNDA 0.104793f
C177 two_stage_opamp_dummy_magic_16_0.VD4.t10 GNDA 0.030951f
C178 two_stage_opamp_dummy_magic_16_0.VD4.t4 GNDA 0.030951f
C179 two_stage_opamp_dummy_magic_16_0.VD4.n9 GNDA 0.108329f
C180 two_stage_opamp_dummy_magic_16_0.VD4.n10 GNDA 0.153987f
C181 two_stage_opamp_dummy_magic_16_0.VD4.t33 GNDA 0.030951f
C182 two_stage_opamp_dummy_magic_16_0.VD4.t37 GNDA 0.030951f
C183 two_stage_opamp_dummy_magic_16_0.VD4.n11 GNDA 0.10726f
C184 two_stage_opamp_dummy_magic_16_0.VD4.n12 GNDA 0.104977f
C185 two_stage_opamp_dummy_magic_16_0.VD4.t14 GNDA 0.030951f
C186 two_stage_opamp_dummy_magic_16_0.VD4.n13 GNDA 0.092854f
C187 two_stage_opamp_dummy_magic_16_0.VD4.n14 GNDA 0.030951f
C188 two_stage_opamp_dummy_magic_16_0.VD4.n15 GNDA 0.017686f
C189 two_stage_opamp_dummy_magic_16_0.VD4.n18 GNDA 0.014321f
C190 two_stage_opamp_dummy_magic_16_0.VD4.n19 GNDA 0.017686f
C191 two_stage_opamp_dummy_magic_16_0.VD4.t15 GNDA 0.054268f
C192 two_stage_opamp_dummy_magic_16_0.VD4.t23 GNDA 0.030951f
C193 two_stage_opamp_dummy_magic_16_0.VD4.t27 GNDA 0.030951f
C194 two_stage_opamp_dummy_magic_16_0.VD4.n20 GNDA 0.10726f
C195 two_stage_opamp_dummy_magic_16_0.VD4.n21 GNDA 0.104977f
C196 two_stage_opamp_dummy_magic_16_0.VD4.t19 GNDA 0.030951f
C197 two_stage_opamp_dummy_magic_16_0.VD4.t21 GNDA 0.030951f
C198 two_stage_opamp_dummy_magic_16_0.VD4.n22 GNDA 0.10726f
C199 two_stage_opamp_dummy_magic_16_0.VD4.n23 GNDA 0.104977f
C200 two_stage_opamp_dummy_magic_16_0.VD4.t31 GNDA 0.030951f
C201 two_stage_opamp_dummy_magic_16_0.VD4.t35 GNDA 0.030951f
C202 two_stage_opamp_dummy_magic_16_0.VD4.n24 GNDA 0.10726f
C203 two_stage_opamp_dummy_magic_16_0.VD4.n25 GNDA 0.104977f
C204 two_stage_opamp_dummy_magic_16_0.VD4.t29 GNDA 0.030951f
C205 two_stage_opamp_dummy_magic_16_0.VD4.t25 GNDA 0.030951f
C206 two_stage_opamp_dummy_magic_16_0.VD4.n26 GNDA 0.10726f
C207 two_stage_opamp_dummy_magic_16_0.VD4.n27 GNDA 0.134403f
C208 two_stage_opamp_dummy_magic_16_0.VD4.n28 GNDA 0.046089f
C209 two_stage_opamp_dummy_magic_16_0.VD4.n29 GNDA 0.030951f
C210 two_stage_opamp_dummy_magic_16_0.VD4.n31 GNDA 0.030951f
C211 two_stage_opamp_dummy_magic_16_0.VD4.n32 GNDA 0.017686f
C212 two_stage_opamp_dummy_magic_16_0.VD4.n33 GNDA 0.017686f
C213 two_stage_opamp_dummy_magic_16_0.VD4.n34 GNDA 0.030951f
C214 two_stage_opamp_dummy_magic_16_0.VD4.n36 GNDA 0.030951f
C215 two_stage_opamp_dummy_magic_16_0.VD4.n37 GNDA 0.017686f
C216 two_stage_opamp_dummy_magic_16_0.VD4.n38 GNDA 0.017686f
C217 two_stage_opamp_dummy_magic_16_0.VD4.n39 GNDA 0.030951f
C218 two_stage_opamp_dummy_magic_16_0.VD4.n40 GNDA 0.031222f
C219 two_stage_opamp_dummy_magic_16_0.VD4.t17 GNDA 0.030951f
C220 two_stage_opamp_dummy_magic_16_0.VD4.n41 GNDA 0.092854f
C221 two_stage_opamp_dummy_magic_16_0.VD4.n42 GNDA 0.029837f
C222 two_stage_opamp_dummy_magic_16_0.VD4.n43 GNDA 0.017686f
C223 two_stage_opamp_dummy_magic_16_0.VD4.n44 GNDA 0.258664f
C224 two_stage_opamp_dummy_magic_16_0.VD4.t16 GNDA 0.224175f
C225 two_stage_opamp_dummy_magic_16_0.VD4.t28 GNDA 0.206931f
C226 two_stage_opamp_dummy_magic_16_0.VD4.t24 GNDA 0.206931f
C227 two_stage_opamp_dummy_magic_16_0.VD4.t30 GNDA 0.206931f
C228 two_stage_opamp_dummy_magic_16_0.VD4.t34 GNDA 0.206931f
C229 two_stage_opamp_dummy_magic_16_0.VD4.t18 GNDA 0.206931f
C230 two_stage_opamp_dummy_magic_16_0.VD4.t20 GNDA 0.206931f
C231 two_stage_opamp_dummy_magic_16_0.VD4.t22 GNDA 0.206931f
C232 two_stage_opamp_dummy_magic_16_0.VD4.t26 GNDA 0.206931f
C233 two_stage_opamp_dummy_magic_16_0.VD4.t32 GNDA 0.206931f
C234 two_stage_opamp_dummy_magic_16_0.VD4.t36 GNDA 0.206931f
C235 two_stage_opamp_dummy_magic_16_0.VD4.t13 GNDA 0.224175f
C236 two_stage_opamp_dummy_magic_16_0.VD4.n46 GNDA 0.014321f
C237 two_stage_opamp_dummy_magic_16_0.VD4.n47 GNDA 0.017686f
C238 two_stage_opamp_dummy_magic_16_0.VD4.n49 GNDA 0.031222f
C239 two_stage_opamp_dummy_magic_16_0.VD4.n50 GNDA 0.030951f
C240 two_stage_opamp_dummy_magic_16_0.VD4.n51 GNDA 0.017686f
C241 two_stage_opamp_dummy_magic_16_0.VD4.n52 GNDA 0.017686f
C242 two_stage_opamp_dummy_magic_16_0.VD4.n53 GNDA 0.030951f
C243 two_stage_opamp_dummy_magic_16_0.VD4.n55 GNDA 0.030951f
C244 two_stage_opamp_dummy_magic_16_0.VD4.n56 GNDA 0.030951f
C245 two_stage_opamp_dummy_magic_16_0.VD4.n57 GNDA 0.017686f
C246 two_stage_opamp_dummy_magic_16_0.VD4.n58 GNDA 0.258664f
C247 two_stage_opamp_dummy_magic_16_0.VD4.n59 GNDA 0.013727f
C248 two_stage_opamp_dummy_magic_16_0.VD4.n60 GNDA 0.033797f
C249 two_stage_opamp_dummy_magic_16_0.VD4.t12 GNDA 0.054268f
C250 two_stage_opamp_dummy_magic_16_0.VD4.n61 GNDA 0.044756f
C251 two_stage_opamp_dummy_magic_16_0.VD4.n62 GNDA 0.062101f
C252 two_stage_opamp_dummy_magic_16_0.VD4.n63 GNDA 0.087485f
C253 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t12 GNDA 0.01637f
C254 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t15 GNDA 0.01637f
C255 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n0 GNDA 0.041052f
C256 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t11 GNDA 0.01637f
C257 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t10 GNDA 0.01637f
C258 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n1 GNDA 0.040835f
C259 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n2 GNDA 0.363013f
C260 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t14 GNDA 0.01637f
C261 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t13 GNDA 0.01637f
C262 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n3 GNDA 0.03274f
C263 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n4 GNDA 0.060861f
C264 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t16 GNDA 0.206157f
C265 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t1 GNDA 0.03274f
C266 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t5 GNDA 0.03274f
C267 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n5 GNDA 0.097293f
C268 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t0 GNDA 0.03274f
C269 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t4 GNDA 0.03274f
C270 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n6 GNDA 0.096862f
C271 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n7 GNDA 0.331325f
C272 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t9 GNDA 0.03274f
C273 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t7 GNDA 0.03274f
C274 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n8 GNDA 0.096862f
C275 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n9 GNDA 0.171607f
C276 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t2 GNDA 0.03274f
C277 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t6 GNDA 0.03274f
C278 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n10 GNDA 0.096862f
C279 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n11 GNDA 0.171607f
C280 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t8 GNDA 0.03274f
C281 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.t3 GNDA 0.03274f
C282 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n12 GNDA 0.096862f
C283 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n13 GNDA 0.239231f
C284 two_stage_opamp_dummy_magic_16_0.V_CMFB_S3.n14 GNDA 1.32734f
C285 bgr_0.V_CMFB_S3 GNDA 1.10386f
C286 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t14 GNDA 0.020156f
C287 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t12 GNDA 0.020156f
C288 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n0 GNDA 0.073261f
C289 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t13 GNDA 0.020156f
C290 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t11 GNDA 0.020156f
C291 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n1 GNDA 0.060879f
C292 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n2 GNDA 1.18743f
C293 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t10 GNDA 0.247627f
C294 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t5 GNDA 0.060467f
C295 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t9 GNDA 0.060467f
C296 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n3 GNDA 0.252232f
C297 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t4 GNDA 0.060467f
C298 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t8 GNDA 0.060467f
C299 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n4 GNDA 0.251304f
C300 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n5 GNDA 0.345024f
C301 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t3 GNDA 0.060467f
C302 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t1 GNDA 0.060467f
C303 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n6 GNDA 0.251304f
C304 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n7 GNDA 0.18003f
C305 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t6 GNDA 0.060467f
C306 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t0 GNDA 0.060467f
C307 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n8 GNDA 0.251304f
C308 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n9 GNDA 0.18003f
C309 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t2 GNDA 0.060467f
C310 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.t7 GNDA 0.060467f
C311 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n10 GNDA 0.251304f
C312 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n11 GNDA 0.249769f
C313 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n12 GNDA 1.34239f
C314 two_stage_opamp_dummy_magic_16_0.V_CMFB_S4.n13 GNDA 1.98073f
C315 bgr_0.V_CMFB_S4 GNDA 0.010078f
C316 two_stage_opamp_dummy_magic_16_0.Y.t12 GNDA 0.031482f
C317 two_stage_opamp_dummy_magic_16_0.Y.t21 GNDA 0.031482f
C318 two_stage_opamp_dummy_magic_16_0.Y.n0 GNDA 0.110568f
C319 two_stage_opamp_dummy_magic_16_0.Y.t22 GNDA 0.031482f
C320 two_stage_opamp_dummy_magic_16_0.Y.t19 GNDA 0.031482f
C321 two_stage_opamp_dummy_magic_16_0.Y.n1 GNDA 0.110188f
C322 two_stage_opamp_dummy_magic_16_0.Y.n2 GNDA 0.205607f
C323 two_stage_opamp_dummy_magic_16_0.Y.t23 GNDA 0.031482f
C324 two_stage_opamp_dummy_magic_16_0.Y.t24 GNDA 0.031482f
C325 two_stage_opamp_dummy_magic_16_0.Y.n3 GNDA 0.110188f
C326 two_stage_opamp_dummy_magic_16_0.Y.n4 GNDA 0.106592f
C327 two_stage_opamp_dummy_magic_16_0.Y.t15 GNDA 0.031482f
C328 two_stage_opamp_dummy_magic_16_0.Y.t16 GNDA 0.031482f
C329 two_stage_opamp_dummy_magic_16_0.Y.n5 GNDA 0.110188f
C330 two_stage_opamp_dummy_magic_16_0.Y.n6 GNDA 0.106592f
C331 two_stage_opamp_dummy_magic_16_0.Y.t20 GNDA 0.031482f
C332 two_stage_opamp_dummy_magic_16_0.Y.t17 GNDA 0.031482f
C333 two_stage_opamp_dummy_magic_16_0.Y.n7 GNDA 0.110188f
C334 two_stage_opamp_dummy_magic_16_0.Y.n8 GNDA 0.125547f
C335 two_stage_opamp_dummy_magic_16_0.Y.t18 GNDA 0.031482f
C336 two_stage_opamp_dummy_magic_16_0.Y.t0 GNDA 0.031482f
C337 two_stage_opamp_dummy_magic_16_0.Y.n9 GNDA 0.107979f
C338 two_stage_opamp_dummy_magic_16_0.Y.n10 GNDA 0.184593f
C339 two_stage_opamp_dummy_magic_16_0.Y.t40 GNDA 0.018889f
C340 two_stage_opamp_dummy_magic_16_0.Y.t54 GNDA 0.018889f
C341 two_stage_opamp_dummy_magic_16_0.Y.t37 GNDA 0.018889f
C342 two_stage_opamp_dummy_magic_16_0.Y.t51 GNDA 0.022937f
C343 two_stage_opamp_dummy_magic_16_0.Y.n11 GNDA 0.022937f
C344 two_stage_opamp_dummy_magic_16_0.Y.n12 GNDA 0.014842f
C345 two_stage_opamp_dummy_magic_16_0.Y.n13 GNDA 0.013091f
C346 two_stage_opamp_dummy_magic_16_0.Y.t26 GNDA 0.018889f
C347 two_stage_opamp_dummy_magic_16_0.Y.t31 GNDA 0.018889f
C348 two_stage_opamp_dummy_magic_16_0.Y.t48 GNDA 0.018889f
C349 two_stage_opamp_dummy_magic_16_0.Y.t34 GNDA 0.018889f
C350 two_stage_opamp_dummy_magic_16_0.Y.t29 GNDA 0.018889f
C351 two_stage_opamp_dummy_magic_16_0.Y.t44 GNDA 0.022937f
C352 two_stage_opamp_dummy_magic_16_0.Y.n14 GNDA 0.022937f
C353 two_stage_opamp_dummy_magic_16_0.Y.n15 GNDA 0.014842f
C354 two_stage_opamp_dummy_magic_16_0.Y.n16 GNDA 0.014842f
C355 two_stage_opamp_dummy_magic_16_0.Y.n17 GNDA 0.014842f
C356 two_stage_opamp_dummy_magic_16_0.Y.n18 GNDA 0.013091f
C357 two_stage_opamp_dummy_magic_16_0.Y.n19 GNDA 0.013602f
C358 two_stage_opamp_dummy_magic_16_0.Y.t28 GNDA 0.029009f
C359 two_stage_opamp_dummy_magic_16_0.Y.t42 GNDA 0.029009f
C360 two_stage_opamp_dummy_magic_16_0.Y.t25 GNDA 0.029009f
C361 two_stage_opamp_dummy_magic_16_0.Y.t39 GNDA 0.032978f
C362 two_stage_opamp_dummy_magic_16_0.Y.n20 GNDA 0.029762f
C363 two_stage_opamp_dummy_magic_16_0.Y.n21 GNDA 0.018215f
C364 two_stage_opamp_dummy_magic_16_0.Y.n22 GNDA 0.016464f
C365 two_stage_opamp_dummy_magic_16_0.Y.t43 GNDA 0.029009f
C366 two_stage_opamp_dummy_magic_16_0.Y.t50 GNDA 0.029009f
C367 two_stage_opamp_dummy_magic_16_0.Y.t36 GNDA 0.029009f
C368 two_stage_opamp_dummy_magic_16_0.Y.t53 GNDA 0.029009f
C369 two_stage_opamp_dummy_magic_16_0.Y.t46 GNDA 0.029009f
C370 two_stage_opamp_dummy_magic_16_0.Y.t32 GNDA 0.032978f
C371 two_stage_opamp_dummy_magic_16_0.Y.n23 GNDA 0.029762f
C372 two_stage_opamp_dummy_magic_16_0.Y.n24 GNDA 0.018215f
C373 two_stage_opamp_dummy_magic_16_0.Y.n25 GNDA 0.018215f
C374 two_stage_opamp_dummy_magic_16_0.Y.n26 GNDA 0.018215f
C375 two_stage_opamp_dummy_magic_16_0.Y.n27 GNDA 0.016464f
C376 two_stage_opamp_dummy_magic_16_0.Y.n28 GNDA 0.013602f
C377 two_stage_opamp_dummy_magic_16_0.Y.n29 GNDA 0.113546f
C378 two_stage_opamp_dummy_magic_16_0.Y.t14 GNDA 0.013493f
C379 two_stage_opamp_dummy_magic_16_0.Y.t5 GNDA 0.013493f
C380 two_stage_opamp_dummy_magic_16_0.Y.n30 GNDA 0.04932f
C381 two_stage_opamp_dummy_magic_16_0.Y.t10 GNDA 0.013493f
C382 two_stage_opamp_dummy_magic_16_0.Y.t4 GNDA 0.013493f
C383 two_stage_opamp_dummy_magic_16_0.Y.n31 GNDA 0.04891f
C384 two_stage_opamp_dummy_magic_16_0.Y.n32 GNDA 0.172519f
C385 two_stage_opamp_dummy_magic_16_0.Y.t8 GNDA 0.013493f
C386 two_stage_opamp_dummy_magic_16_0.Y.t11 GNDA 0.013493f
C387 two_stage_opamp_dummy_magic_16_0.Y.n33 GNDA 0.04891f
C388 two_stage_opamp_dummy_magic_16_0.Y.n34 GNDA 0.089613f
C389 two_stage_opamp_dummy_magic_16_0.Y.t9 GNDA 0.013493f
C390 two_stage_opamp_dummy_magic_16_0.Y.t3 GNDA 0.013493f
C391 two_stage_opamp_dummy_magic_16_0.Y.n35 GNDA 0.04891f
C392 two_stage_opamp_dummy_magic_16_0.Y.n36 GNDA 0.089613f
C393 two_stage_opamp_dummy_magic_16_0.Y.t7 GNDA 0.013493f
C394 two_stage_opamp_dummy_magic_16_0.Y.t2 GNDA 0.013493f
C395 two_stage_opamp_dummy_magic_16_0.Y.n37 GNDA 0.04891f
C396 two_stage_opamp_dummy_magic_16_0.Y.n38 GNDA 0.089613f
C397 two_stage_opamp_dummy_magic_16_0.Y.t6 GNDA 0.013493f
C398 two_stage_opamp_dummy_magic_16_0.Y.t13 GNDA 0.013493f
C399 two_stage_opamp_dummy_magic_16_0.Y.n39 GNDA 0.04891f
C400 two_stage_opamp_dummy_magic_16_0.Y.n40 GNDA 0.136366f
C401 two_stage_opamp_dummy_magic_16_0.Y.n41 GNDA 0.119935f
C402 two_stage_opamp_dummy_magic_16_0.Y.n42 GNDA 0.215844f
C403 two_stage_opamp_dummy_magic_16_0.Y.t38 GNDA 0.059367f
C404 two_stage_opamp_dummy_magic_16_0.Y.t52 GNDA 0.059367f
C405 two_stage_opamp_dummy_magic_16_0.Y.t35 GNDA 0.059367f
C406 two_stage_opamp_dummy_magic_16_0.Y.t49 GNDA 0.059367f
C407 two_stage_opamp_dummy_magic_16_0.Y.t33 GNDA 0.06323f
C408 two_stage_opamp_dummy_magic_16_0.Y.n43 GNDA 0.050107f
C409 two_stage_opamp_dummy_magic_16_0.Y.n44 GNDA 0.028334f
C410 two_stage_opamp_dummy_magic_16_0.Y.n45 GNDA 0.028334f
C411 two_stage_opamp_dummy_magic_16_0.Y.n46 GNDA 0.02659f
C412 two_stage_opamp_dummy_magic_16_0.Y.t45 GNDA 0.059367f
C413 two_stage_opamp_dummy_magic_16_0.Y.t30 GNDA 0.059367f
C414 two_stage_opamp_dummy_magic_16_0.Y.t47 GNDA 0.059367f
C415 two_stage_opamp_dummy_magic_16_0.Y.t41 GNDA 0.059367f
C416 two_stage_opamp_dummy_magic_16_0.Y.t27 GNDA 0.06323f
C417 two_stage_opamp_dummy_magic_16_0.Y.n47 GNDA 0.050107f
C418 two_stage_opamp_dummy_magic_16_0.Y.n48 GNDA 0.028334f
C419 two_stage_opamp_dummy_magic_16_0.Y.n49 GNDA 0.028334f
C420 two_stage_opamp_dummy_magic_16_0.Y.n50 GNDA 0.02659f
C421 two_stage_opamp_dummy_magic_16_0.Y.n51 GNDA 0.016175f
C422 two_stage_opamp_dummy_magic_16_0.Y.n52 GNDA 0.510557f
C423 two_stage_opamp_dummy_magic_16_0.Y.t1 GNDA 0.437339f
C424 bgr_0.Vin-.n0 GNDA 0.069747f
C425 bgr_0.Vin-.n1 GNDA 0.078367f
C426 bgr_0.Vin-.n2 GNDA 0.113033f
C427 bgr_0.Vin-.t2 GNDA 0.261601f
C428 bgr_0.Vin-.t6 GNDA 0.027101f
C429 bgr_0.Vin-.t4 GNDA 0.027101f
C430 bgr_0.Vin-.n3 GNDA 0.094346f
C431 bgr_0.Vin-.t3 GNDA 0.027101f
C432 bgr_0.Vin-.t5 GNDA 0.027101f
C433 bgr_0.Vin-.n4 GNDA 0.090091f
C434 bgr_0.Vin-.n5 GNDA 0.386489f
C435 bgr_0.Vin-.n6 GNDA 0.027681f
C436 bgr_0.Vin-.n7 GNDA 0.366254f
C437 bgr_0.Vin-.t12 GNDA 0.022346f
C438 bgr_0.Vin-.n8 GNDA 0.026209f
C439 bgr_0.Vin-.n9 GNDA 0.021455f
C440 bgr_0.Vin-.n10 GNDA 0.021455f
C441 bgr_0.Vin-.n11 GNDA 0.036491f
C442 bgr_0.Vin-.n12 GNDA 0.497932f
C443 bgr_0.Vin-.t7 GNDA 0.117924f
C444 bgr_0.Vin-.n13 GNDA 0.65583f
C445 bgr_0.Vin-.n14 GNDA 1.073f
C446 bgr_0.Vin-.n15 GNDA 0.471409f
C447 bgr_0.Vin-.n16 GNDA 0.07053f
C448 bgr_0.Vin-.n17 GNDA 0.119504f
C449 bgr_0.Vin-.n18 GNDA 0.069875f
C450 bgr_0.Vin-.n19 GNDA 0.138215f
C451 bgr_0.Vin-.n20 GNDA 0.138215f
C452 bgr_0.Vin-.n21 GNDA -0.269519f
C453 bgr_0.Vin-.n22 GNDA 0.445457f
C454 bgr_0.Vin-.n23 GNDA 0.213551f
C455 bgr_0.Vin-.n24 GNDA 0.403461f
C456 bgr_0.Vin-.n25 GNDA 0.0384f
C457 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter GNDA 0.040751f
C458 bgr_0.V_mir2.t7 GNDA 0.019293f
C459 bgr_0.V_mir2.n0 GNDA 0.025223f
C460 bgr_0.V_mir2.t14 GNDA 0.041163f
C461 bgr_0.V_mir2.n1 GNDA 0.027381f
C462 bgr_0.V_mir2.n2 GNDA 0.451535f
C463 bgr_0.V_mir2.n3 GNDA 0.146338f
C464 bgr_0.V_mir2.t4 GNDA 0.023151f
C465 bgr_0.V_mir2.t17 GNDA 0.023151f
C466 bgr_0.V_mir2.t20 GNDA 0.037369f
C467 bgr_0.V_mir2.n4 GNDA 0.041731f
C468 bgr_0.V_mir2.n5 GNDA 0.028507f
C469 bgr_0.V_mir2.t0 GNDA 0.02939f
C470 bgr_0.V_mir2.n6 GNDA 0.044354f
C471 bgr_0.V_mir2.t5 GNDA 0.019293f
C472 bgr_0.V_mir2.t1 GNDA 0.019293f
C473 bgr_0.V_mir2.n7 GNDA 0.044166f
C474 bgr_0.V_mir2.n8 GNDA 0.109943f
C475 bgr_0.V_mir2.t2 GNDA 0.023151f
C476 bgr_0.V_mir2.t18 GNDA 0.023151f
C477 bgr_0.V_mir2.t22 GNDA 0.037369f
C478 bgr_0.V_mir2.n9 GNDA 0.041731f
C479 bgr_0.V_mir2.n10 GNDA 0.028507f
C480 bgr_0.V_mir2.t8 GNDA 0.02939f
C481 bgr_0.V_mir2.n11 GNDA 0.044354f
C482 bgr_0.V_mir2.t3 GNDA 0.019293f
C483 bgr_0.V_mir2.t9 GNDA 0.019293f
C484 bgr_0.V_mir2.n12 GNDA 0.044166f
C485 bgr_0.V_mir2.n13 GNDA 0.111042f
C486 bgr_0.V_mir2.n14 GNDA 0.381359f
C487 bgr_0.V_mir2.n15 GNDA 0.051125f
C488 bgr_0.V_mir2.t6 GNDA 0.023151f
C489 bgr_0.V_mir2.t19 GNDA 0.023151f
C490 bgr_0.V_mir2.t21 GNDA 0.037369f
C491 bgr_0.V_mir2.n16 GNDA 0.041731f
C492 bgr_0.V_mir2.n17 GNDA 0.028507f
C493 bgr_0.V_mir2.t10 GNDA 0.02939f
C494 bgr_0.V_mir2.n18 GNDA 0.044354f
C495 bgr_0.V_mir2.n19 GNDA 0.085095f
C496 bgr_0.V_mir2.n20 GNDA 0.044166f
C497 bgr_0.V_mir2.t11 GNDA 0.019293f
C498 bgr_0.cap_res1.t11 GNDA 0.331712f
C499 bgr_0.cap_res1.t18 GNDA 0.349187f
C500 bgr_0.cap_res1.t15 GNDA 0.350452f
C501 bgr_0.cap_res1.t4 GNDA 0.331712f
C502 bgr_0.cap_res1.t14 GNDA 0.349187f
C503 bgr_0.cap_res1.t8 GNDA 0.350452f
C504 bgr_0.cap_res1.t10 GNDA 0.331712f
C505 bgr_0.cap_res1.t17 GNDA 0.349187f
C506 bgr_0.cap_res1.t13 GNDA 0.350452f
C507 bgr_0.cap_res1.t3 GNDA 0.331712f
C508 bgr_0.cap_res1.t12 GNDA 0.349187f
C509 bgr_0.cap_res1.t6 GNDA 0.350452f
C510 bgr_0.cap_res1.t19 GNDA 0.331712f
C511 bgr_0.cap_res1.t5 GNDA 0.349187f
C512 bgr_0.cap_res1.t0 GNDA 0.350452f
C513 bgr_0.cap_res1.n0 GNDA 0.23406f
C514 bgr_0.cap_res1.t16 GNDA 0.186395f
C515 bgr_0.cap_res1.n1 GNDA 0.253961f
C516 bgr_0.cap_res1.t1 GNDA 0.186395f
C517 bgr_0.cap_res1.n2 GNDA 0.253961f
C518 bgr_0.cap_res1.t7 GNDA 0.186395f
C519 bgr_0.cap_res1.n3 GNDA 0.253961f
C520 bgr_0.cap_res1.t2 GNDA 0.186395f
C521 bgr_0.cap_res1.n4 GNDA 0.253961f
C522 bgr_0.cap_res1.t9 GNDA 0.363549f
C523 bgr_0.cap_res1.t20 GNDA 0.08421f
C524 bgr_0.PFET_GATE_10uA.t28 GNDA 0.020856f
C525 bgr_0.PFET_GATE_10uA.t20 GNDA 0.030831f
C526 bgr_0.PFET_GATE_10uA.n0 GNDA 0.033972f
C527 bgr_0.PFET_GATE_10uA.t15 GNDA 0.020856f
C528 bgr_0.PFET_GATE_10uA.t21 GNDA 0.030831f
C529 bgr_0.PFET_GATE_10uA.n1 GNDA 0.033972f
C530 bgr_0.PFET_GATE_10uA.n2 GNDA 0.040878f
C531 bgr_0.PFET_GATE_10uA.t19 GNDA 0.020856f
C532 bgr_0.PFET_GATE_10uA.t12 GNDA 0.030831f
C533 bgr_0.PFET_GATE_10uA.n3 GNDA 0.033972f
C534 bgr_0.PFET_GATE_10uA.t26 GNDA 0.020856f
C535 bgr_0.PFET_GATE_10uA.t13 GNDA 0.030831f
C536 bgr_0.PFET_GATE_10uA.n4 GNDA 0.033972f
C537 bgr_0.PFET_GATE_10uA.n5 GNDA 0.034081f
C538 bgr_0.PFET_GATE_10uA.t7 GNDA 0.312465f
C539 bgr_0.PFET_GATE_10uA.t1 GNDA 0.021391f
C540 bgr_0.PFET_GATE_10uA.t8 GNDA 0.021391f
C541 bgr_0.PFET_GATE_10uA.n6 GNDA 0.054673f
C542 bgr_0.PFET_GATE_10uA.t3 GNDA 0.021391f
C543 bgr_0.PFET_GATE_10uA.t5 GNDA 0.021391f
C544 bgr_0.PFET_GATE_10uA.n7 GNDA 0.05326f
C545 bgr_0.PFET_GATE_10uA.n8 GNDA 0.520952f
C546 bgr_0.PFET_GATE_10uA.t4 GNDA 0.021391f
C547 bgr_0.PFET_GATE_10uA.t6 GNDA 0.021391f
C548 bgr_0.PFET_GATE_10uA.n9 GNDA 0.05326f
C549 bgr_0.PFET_GATE_10uA.n10 GNDA 0.295408f
C550 bgr_0.PFET_GATE_10uA.n11 GNDA 0.603055f
C551 bgr_0.PFET_GATE_10uA.t9 GNDA 0.021391f
C552 bgr_0.PFET_GATE_10uA.t2 GNDA 0.021391f
C553 bgr_0.PFET_GATE_10uA.n12 GNDA 0.05159f
C554 bgr_0.PFET_GATE_10uA.n13 GNDA 0.275411f
C555 bgr_0.PFET_GATE_10uA.t0 GNDA 0.464967f
C556 bgr_0.PFET_GATE_10uA.t27 GNDA 0.024114f
C557 bgr_0.PFET_GATE_10uA.t14 GNDA 0.024114f
C558 bgr_0.PFET_GATE_10uA.n14 GNDA 0.069715f
C559 bgr_0.PFET_GATE_10uA.n15 GNDA 1.91969f
C560 bgr_0.PFET_GATE_10uA.n16 GNDA 0.771508f
C561 bgr_0.PFET_GATE_10uA.n17 GNDA 0.759224f
C562 bgr_0.PFET_GATE_10uA.t11 GNDA 0.020856f
C563 bgr_0.PFET_GATE_10uA.t25 GNDA 0.020856f
C564 bgr_0.PFET_GATE_10uA.t18 GNDA 0.020856f
C565 bgr_0.PFET_GATE_10uA.t10 GNDA 0.020856f
C566 bgr_0.PFET_GATE_10uA.t24 GNDA 0.020856f
C567 bgr_0.PFET_GATE_10uA.t17 GNDA 0.030831f
C568 bgr_0.PFET_GATE_10uA.n18 GNDA 0.038154f
C569 bgr_0.PFET_GATE_10uA.n19 GNDA 0.027273f
C570 bgr_0.PFET_GATE_10uA.n20 GNDA 0.027273f
C571 bgr_0.PFET_GATE_10uA.n21 GNDA 0.027273f
C572 bgr_0.PFET_GATE_10uA.n22 GNDA 0.023091f
C573 bgr_0.PFET_GATE_10uA.t16 GNDA 0.020856f
C574 bgr_0.PFET_GATE_10uA.t23 GNDA 0.020856f
C575 bgr_0.PFET_GATE_10uA.t22 GNDA 0.020856f
C576 bgr_0.PFET_GATE_10uA.t29 GNDA 0.030831f
C577 bgr_0.PFET_GATE_10uA.n23 GNDA 0.038154f
C578 bgr_0.PFET_GATE_10uA.n24 GNDA 0.027273f
C579 bgr_0.PFET_GATE_10uA.n25 GNDA 0.023091f
C580 bgr_0.PFET_GATE_10uA.n26 GNDA 0.031695f
C581 two_stage_opamp_dummy_magic_16_0.Vb1.n0 GNDA 0.016648f
C582 two_stage_opamp_dummy_magic_16_0.Vb1.n1 GNDA 0.016536f
C583 two_stage_opamp_dummy_magic_16_0.Vb1.n2 GNDA 0.181582f
C584 two_stage_opamp_dummy_magic_16_0.Vb1.t16 GNDA 0.298213f
C585 two_stage_opamp_dummy_magic_16_0.Vb1.n3 GNDA 0.035064f
C586 two_stage_opamp_dummy_magic_16_0.Vb1.n4 GNDA 0.228582f
C587 two_stage_opamp_dummy_magic_16_0.Vb1.t3 GNDA 0.010211f
C588 two_stage_opamp_dummy_magic_16_0.Vb1.t5 GNDA 0.013244f
C589 two_stage_opamp_dummy_magic_16_0.Vb1.n5 GNDA 0.013617f
C590 two_stage_opamp_dummy_magic_16_0.Vb1.t7 GNDA 0.010211f
C591 two_stage_opamp_dummy_magic_16_0.Vb1.t1 GNDA 0.013244f
C592 two_stage_opamp_dummy_magic_16_0.Vb1.n6 GNDA 0.013617f
C593 two_stage_opamp_dummy_magic_16_0.Vb1.n8 GNDA 0.030997f
C594 two_stage_opamp_dummy_magic_16_0.Vb1.n9 GNDA 0.033569f
C595 two_stage_opamp_dummy_magic_16_0.Vb1.n10 GNDA 0.027085f
C596 two_stage_opamp_dummy_magic_16_0.Vb1.n11 GNDA 0.035064f
C597 two_stage_opamp_dummy_magic_16_0.Vb1.n12 GNDA 0.183099f
C598 two_stage_opamp_dummy_magic_16_0.Vb1.t14 GNDA 0.010211f
C599 two_stage_opamp_dummy_magic_16_0.Vb1.t25 GNDA 0.010211f
C600 two_stage_opamp_dummy_magic_16_0.Vb1.t34 GNDA 0.010211f
C601 two_stage_opamp_dummy_magic_16_0.Vb1.t17 GNDA 0.010211f
C602 two_stage_opamp_dummy_magic_16_0.Vb1.t27 GNDA 0.013244f
C603 two_stage_opamp_dummy_magic_16_0.Vb1.n13 GNDA 0.0144f
C604 two_stage_opamp_dummy_magic_16_0.Vb1.t26 GNDA 0.010211f
C605 two_stage_opamp_dummy_magic_16_0.Vb1.t30 GNDA 0.010211f
C606 two_stage_opamp_dummy_magic_16_0.Vb1.t21 GNDA 0.010211f
C607 two_stage_opamp_dummy_magic_16_0.Vb1.t32 GNDA 0.010211f
C608 two_stage_opamp_dummy_magic_16_0.Vb1.t23 GNDA 0.013244f
C609 two_stage_opamp_dummy_magic_16_0.Vb1.n17 GNDA 0.0144f
C610 two_stage_opamp_dummy_magic_16_0.Vb1.n21 GNDA 0.013791f
C611 two_stage_opamp_dummy_magic_16_0.Vb1.t15 GNDA 0.010211f
C612 two_stage_opamp_dummy_magic_16_0.Vb1.t20 GNDA 0.010211f
C613 two_stage_opamp_dummy_magic_16_0.Vb1.t29 GNDA 0.010211f
C614 two_stage_opamp_dummy_magic_16_0.Vb1.t18 GNDA 0.010211f
C615 two_stage_opamp_dummy_magic_16_0.Vb1.t28 GNDA 0.013244f
C616 two_stage_opamp_dummy_magic_16_0.Vb1.n22 GNDA 0.0144f
C617 two_stage_opamp_dummy_magic_16_0.Vb1.t19 GNDA 0.010211f
C618 two_stage_opamp_dummy_magic_16_0.Vb1.t31 GNDA 0.010211f
C619 two_stage_opamp_dummy_magic_16_0.Vb1.t22 GNDA 0.010211f
C620 two_stage_opamp_dummy_magic_16_0.Vb1.t33 GNDA 0.010211f
C621 two_stage_opamp_dummy_magic_16_0.Vb1.t24 GNDA 0.013244f
C622 two_stage_opamp_dummy_magic_16_0.Vb1.n26 GNDA 0.0144f
C623 two_stage_opamp_dummy_magic_16_0.Vb1.n30 GNDA 0.010439f
C624 two_stage_opamp_dummy_magic_16_0.Vb1.n31 GNDA 0.224385f
C625 two_stage_opamp_dummy_magic_16_0.Vb1.n32 GNDA 0.53241f
C626 bgr_0.VB1_CUR_BIAS GNDA 0.377177f
C627 two_stage_opamp_dummy_magic_16_0.Vb2.t32 GNDA 0.043632f
C628 two_stage_opamp_dummy_magic_16_0.Vb2.t14 GNDA 0.043632f
C629 two_stage_opamp_dummy_magic_16_0.Vb2.t19 GNDA 0.043632f
C630 two_stage_opamp_dummy_magic_16_0.Vb2.t26 GNDA 0.043632f
C631 two_stage_opamp_dummy_magic_16_0.Vb2.t22 GNDA 0.050351f
C632 two_stage_opamp_dummy_magic_16_0.Vb2.n0 GNDA 0.04088f
C633 two_stage_opamp_dummy_magic_16_0.Vb2.n1 GNDA 0.025122f
C634 two_stage_opamp_dummy_magic_16_0.Vb2.n2 GNDA 0.025122f
C635 two_stage_opamp_dummy_magic_16_0.Vb2.n3 GNDA 0.023309f
C636 two_stage_opamp_dummy_magic_16_0.Vb2.t29 GNDA 0.043632f
C637 two_stage_opamp_dummy_magic_16_0.Vb2.t28 GNDA 0.043632f
C638 two_stage_opamp_dummy_magic_16_0.Vb2.t24 GNDA 0.043632f
C639 two_stage_opamp_dummy_magic_16_0.Vb2.t17 GNDA 0.043632f
C640 two_stage_opamp_dummy_magic_16_0.Vb2.t12 GNDA 0.050351f
C641 two_stage_opamp_dummy_magic_16_0.Vb2.n4 GNDA 0.04088f
C642 two_stage_opamp_dummy_magic_16_0.Vb2.n5 GNDA 0.025122f
C643 two_stage_opamp_dummy_magic_16_0.Vb2.n6 GNDA 0.025122f
C644 two_stage_opamp_dummy_magic_16_0.Vb2.n7 GNDA 0.023309f
C645 two_stage_opamp_dummy_magic_16_0.Vb2.n8 GNDA 0.013512f
C646 two_stage_opamp_dummy_magic_16_0.Vb2.t11 GNDA 0.043632f
C647 two_stage_opamp_dummy_magic_16_0.Vb2.t15 GNDA 0.043632f
C648 two_stage_opamp_dummy_magic_16_0.Vb2.t20 GNDA 0.043632f
C649 two_stage_opamp_dummy_magic_16_0.Vb2.t16 GNDA 0.043632f
C650 two_stage_opamp_dummy_magic_16_0.Vb2.t23 GNDA 0.050351f
C651 two_stage_opamp_dummy_magic_16_0.Vb2.n9 GNDA 0.04088f
C652 two_stage_opamp_dummy_magic_16_0.Vb2.n10 GNDA 0.025122f
C653 two_stage_opamp_dummy_magic_16_0.Vb2.n11 GNDA 0.025122f
C654 two_stage_opamp_dummy_magic_16_0.Vb2.n12 GNDA 0.023309f
C655 two_stage_opamp_dummy_magic_16_0.Vb2.t30 GNDA 0.043632f
C656 two_stage_opamp_dummy_magic_16_0.Vb2.t21 GNDA 0.043632f
C657 two_stage_opamp_dummy_magic_16_0.Vb2.t25 GNDA 0.043632f
C658 two_stage_opamp_dummy_magic_16_0.Vb2.t18 GNDA 0.043632f
C659 two_stage_opamp_dummy_magic_16_0.Vb2.t13 GNDA 0.050351f
C660 two_stage_opamp_dummy_magic_16_0.Vb2.n13 GNDA 0.04088f
C661 two_stage_opamp_dummy_magic_16_0.Vb2.n14 GNDA 0.025122f
C662 two_stage_opamp_dummy_magic_16_0.Vb2.n15 GNDA 0.025122f
C663 two_stage_opamp_dummy_magic_16_0.Vb2.n16 GNDA 0.023309f
C664 two_stage_opamp_dummy_magic_16_0.Vb2.n17 GNDA 0.016397f
C665 two_stage_opamp_dummy_magic_16_0.Vb2.n18 GNDA 0.03003f
C666 two_stage_opamp_dummy_magic_16_0.Vb2.n19 GNDA 0.029147f
C667 two_stage_opamp_dummy_magic_16_0.Vb2.n20 GNDA 0.303104f
C668 two_stage_opamp_dummy_magic_16_0.Vb2.n21 GNDA 0.029147f
C669 two_stage_opamp_dummy_magic_16_0.Vb2.n22 GNDA 0.204441f
C670 two_stage_opamp_dummy_magic_16_0.Vb2.n23 GNDA 0.029147f
C671 two_stage_opamp_dummy_magic_16_0.Vb2.n24 GNDA 0.808923f
C672 two_stage_opamp_dummy_magic_16_0.Vb2.t31 GNDA 0.053353f
C673 two_stage_opamp_dummy_magic_16_0.Vb2.n25 GNDA 0.723168f
C674 two_stage_opamp_dummy_magic_16_0.Vb2.t10 GNDA 0.030851f
C675 two_stage_opamp_dummy_magic_16_0.Vb2.t8 GNDA 0.030851f
C676 two_stage_opamp_dummy_magic_16_0.Vb2.n26 GNDA 0.107063f
C677 two_stage_opamp_dummy_magic_16_0.Vb2.t9 GNDA 0.053353f
C678 two_stage_opamp_dummy_magic_16_0.Vb2.n27 GNDA 0.18525f
C679 two_stage_opamp_dummy_magic_16_0.Vb2.t27 GNDA 0.031502f
C680 two_stage_opamp_dummy_magic_16_0.Vb2.n28 GNDA 0.094361f
C681 two_stage_opamp_dummy_magic_16_0.Vb2.n29 GNDA 0.154162f
C682 two_stage_opamp_dummy_magic_16_0.Vb2.n30 GNDA 0.287807f
C683 bgr_0.cap_res2.t7 GNDA 0.358376f
C684 bgr_0.cap_res2.t13 GNDA 0.359675f
C685 bgr_0.cap_res2.t15 GNDA 0.340442f
C686 bgr_0.cap_res2.t1 GNDA 0.358376f
C687 bgr_0.cap_res2.t6 GNDA 0.359675f
C688 bgr_0.cap_res2.t9 GNDA 0.340442f
C689 bgr_0.cap_res2.t5 GNDA 0.358376f
C690 bgr_0.cap_res2.t11 GNDA 0.359675f
C691 bgr_0.cap_res2.t14 GNDA 0.340442f
C692 bgr_0.cap_res2.t20 GNDA 0.358376f
C693 bgr_0.cap_res2.t4 GNDA 0.359675f
C694 bgr_0.cap_res2.t8 GNDA 0.340442f
C695 bgr_0.cap_res2.t16 GNDA 0.358376f
C696 bgr_0.cap_res2.t19 GNDA 0.359675f
C697 bgr_0.cap_res2.t2 GNDA 0.340442f
C698 bgr_0.cap_res2.n0 GNDA 0.24022f
C699 bgr_0.cap_res2.t3 GNDA 0.1913f
C700 bgr_0.cap_res2.n1 GNDA 0.260644f
C701 bgr_0.cap_res2.t10 GNDA 0.1913f
C702 bgr_0.cap_res2.n2 GNDA 0.260644f
C703 bgr_0.cap_res2.t17 GNDA 0.1913f
C704 bgr_0.cap_res2.n3 GNDA 0.260644f
C705 bgr_0.cap_res2.t12 GNDA 0.1913f
C706 bgr_0.cap_res2.n4 GNDA 0.260644f
C707 bgr_0.cap_res2.t18 GNDA 0.373116f
C708 bgr_0.cap_res2.t0 GNDA 0.086426f
C709 bgr_0.1st_Vout_2.n0 GNDA 0.569806f
C710 bgr_0.1st_Vout_2.n1 GNDA 0.252461f
C711 bgr_0.1st_Vout_2.n2 GNDA 1.43086f
C712 bgr_0.1st_Vout_2.n3 GNDA 0.104399f
C713 bgr_0.1st_Vout_2.n4 GNDA 1.45767f
C714 bgr_0.1st_Vout_2.t33 GNDA 0.017308f
C715 bgr_0.1st_Vout_2.t28 GNDA 0.288462f
C716 bgr_0.1st_Vout_2.t17 GNDA 0.293375f
C717 bgr_0.1st_Vout_2.t12 GNDA 0.288462f
C718 bgr_0.1st_Vout_2.t32 GNDA 0.288462f
C719 bgr_0.1st_Vout_2.t35 GNDA 0.293375f
C720 bgr_0.1st_Vout_2.t11 GNDA 0.293375f
C721 bgr_0.1st_Vout_2.t31 GNDA 0.288462f
C722 bgr_0.1st_Vout_2.t23 GNDA 0.288462f
C723 bgr_0.1st_Vout_2.t26 GNDA 0.293375f
C724 bgr_0.1st_Vout_2.t30 GNDA 0.293375f
C725 bgr_0.1st_Vout_2.t22 GNDA 0.288462f
C726 bgr_0.1st_Vout_2.t15 GNDA 0.288462f
C727 bgr_0.1st_Vout_2.t19 GNDA 0.293375f
C728 bgr_0.1st_Vout_2.t36 GNDA 0.293375f
C729 bgr_0.1st_Vout_2.t29 GNDA 0.288462f
C730 bgr_0.1st_Vout_2.t21 GNDA 0.288462f
C731 bgr_0.1st_Vout_2.t25 GNDA 0.293375f
C732 bgr_0.1st_Vout_2.t18 GNDA 0.293375f
C733 bgr_0.1st_Vout_2.t14 GNDA 0.288462f
C734 bgr_0.1st_Vout_2.t20 GNDA 0.288462f
C735 bgr_0.1st_Vout_2.t34 GNDA 0.018845f
C736 bgr_0.1st_Vout_2.n5 GNDA 0.018179f
C737 bgr_0.1st_Vout_2.t27 GNDA 0.010986f
C738 bgr_0.1st_Vout_2.t16 GNDA 0.010986f
C739 bgr_0.1st_Vout_2.n6 GNDA 0.024439f
C740 bgr_0.1st_Vout_2.n7 GNDA 0.010417f
C741 bgr_0.1st_Vout_2.t3 GNDA 0.015189f
C742 bgr_0.1st_Vout_2.n8 GNDA 0.157567f
C743 bgr_0.1st_Vout_2.n10 GNDA 0.017425f
C744 bgr_0.1st_Vout_2.t24 GNDA 0.010986f
C745 bgr_0.1st_Vout_2.t13 GNDA 0.010986f
C746 bgr_0.1st_Vout_2.n11 GNDA 0.024439f
C747 bgr_0.1st_Vout_2.n12 GNDA 0.138311f
C748 bgr_0.1st_Vout_2.n13 GNDA 0.018179f
C749 bgr_0.1st_Vout_1.n0 GNDA 0.538712f
C750 bgr_0.1st_Vout_1.n1 GNDA 0.236313f
C751 bgr_0.1st_Vout_1.n2 GNDA 0.973284f
C752 bgr_0.1st_Vout_1.n3 GNDA 0.907198f
C753 bgr_0.1st_Vout_1.n4 GNDA 0.891647f
C754 bgr_0.1st_Vout_1.t11 GNDA 0.358463f
C755 bgr_0.1st_Vout_1.t15 GNDA 0.35246f
C756 bgr_0.1st_Vout_1.t29 GNDA 0.358463f
C757 bgr_0.1st_Vout_1.t35 GNDA 0.35246f
C758 bgr_0.1st_Vout_1.t31 GNDA 0.358463f
C759 bgr_0.1st_Vout_1.t34 GNDA 0.35246f
C760 bgr_0.1st_Vout_1.t20 GNDA 0.358463f
C761 bgr_0.1st_Vout_1.t28 GNDA 0.35246f
C762 bgr_0.1st_Vout_1.t24 GNDA 0.358463f
C763 bgr_0.1st_Vout_1.t27 GNDA 0.35246f
C764 bgr_0.1st_Vout_1.t14 GNDA 0.358463f
C765 bgr_0.1st_Vout_1.t19 GNDA 0.35246f
C766 bgr_0.1st_Vout_1.t30 GNDA 0.358463f
C767 bgr_0.1st_Vout_1.t33 GNDA 0.35246f
C768 bgr_0.1st_Vout_1.t18 GNDA 0.358463f
C769 bgr_0.1st_Vout_1.t26 GNDA 0.35246f
C770 bgr_0.1st_Vout_1.t23 GNDA 0.358463f
C771 bgr_0.1st_Vout_1.t25 GNDA 0.35246f
C772 bgr_0.1st_Vout_1.t17 GNDA 0.35246f
C773 bgr_0.1st_Vout_1.t12 GNDA 0.35246f
C774 bgr_0.1st_Vout_1.t21 GNDA 0.023025f
C775 bgr_0.1st_Vout_1.n5 GNDA 0.715456f
C776 bgr_0.1st_Vout_1.n6 GNDA 0.022212f
C777 bgr_0.1st_Vout_1.n7 GNDA 0.104674f
C778 bgr_0.1st_Vout_1.t36 GNDA 0.013423f
C779 bgr_0.1st_Vout_1.t16 GNDA 0.013423f
C780 bgr_0.1st_Vout_1.n8 GNDA 0.029862f
C781 bgr_0.1st_Vout_1.n9 GNDA 0.082514f
C782 bgr_0.1st_Vout_1.t10 GNDA 0.018559f
C783 bgr_0.1st_Vout_1.n10 GNDA 0.012728f
C784 bgr_0.1st_Vout_1.n11 GNDA 0.192525f
C785 bgr_0.1st_Vout_1.n12 GNDA 0.011517f
C786 bgr_0.1st_Vout_1.n13 GNDA 0.048842f
C787 bgr_0.1st_Vout_1.n14 GNDA 0.021291f
C788 bgr_0.1st_Vout_1.n15 GNDA 0.078719f
C789 bgr_0.1st_Vout_1.n16 GNDA 0.038771f
C790 bgr_0.1st_Vout_1.t32 GNDA 0.013423f
C791 bgr_0.1st_Vout_1.t22 GNDA 0.013423f
C792 bgr_0.1st_Vout_1.n17 GNDA 0.029862f
C793 bgr_0.1st_Vout_1.n18 GNDA 0.082514f
C794 bgr_0.1st_Vout_1.n19 GNDA 0.022212f
C795 bgr_0.1st_Vout_1.n20 GNDA 0.104674f
C796 bgr_0.1st_Vout_1.t13 GNDA 0.021069f
C797 bgr_0.V_mir1.t7 GNDA 0.019293f
C798 bgr_0.V_mir1.t0 GNDA 0.02939f
C799 bgr_0.V_mir1.t4 GNDA 0.023151f
C800 bgr_0.V_mir1.t18 GNDA 0.023151f
C801 bgr_0.V_mir1.t20 GNDA 0.037369f
C802 bgr_0.V_mir1.n0 GNDA 0.041731f
C803 bgr_0.V_mir1.n1 GNDA 0.028507f
C804 bgr_0.V_mir1.n2 GNDA 0.044354f
C805 bgr_0.V_mir1.t1 GNDA 0.019293f
C806 bgr_0.V_mir1.t5 GNDA 0.019293f
C807 bgr_0.V_mir1.n3 GNDA 0.044166f
C808 bgr_0.V_mir1.n4 GNDA 0.109943f
C809 bgr_0.V_mir1.n5 GNDA 0.025223f
C810 bgr_0.V_mir1.t12 GNDA 0.041163f
C811 bgr_0.V_mir1.n6 GNDA 0.027381f
C812 bgr_0.V_mir1.n7 GNDA 0.451535f
C813 bgr_0.V_mir1.n8 GNDA 0.146338f
C814 bgr_0.V_mir1.t2 GNDA 0.02939f
C815 bgr_0.V_mir1.t8 GNDA 0.023151f
C816 bgr_0.V_mir1.t17 GNDA 0.023151f
C817 bgr_0.V_mir1.t21 GNDA 0.037369f
C818 bgr_0.V_mir1.n9 GNDA 0.041731f
C819 bgr_0.V_mir1.n10 GNDA 0.028507f
C820 bgr_0.V_mir1.n11 GNDA 0.044354f
C821 bgr_0.V_mir1.t3 GNDA 0.019293f
C822 bgr_0.V_mir1.t9 GNDA 0.019293f
C823 bgr_0.V_mir1.n12 GNDA 0.044166f
C824 bgr_0.V_mir1.n13 GNDA 0.085095f
C825 bgr_0.V_mir1.n14 GNDA 0.051125f
C826 bgr_0.V_mir1.n15 GNDA 0.381359f
C827 bgr_0.V_mir1.t6 GNDA 0.02939f
C828 bgr_0.V_mir1.t10 GNDA 0.023151f
C829 bgr_0.V_mir1.t22 GNDA 0.023151f
C830 bgr_0.V_mir1.t19 GNDA 0.037369f
C831 bgr_0.V_mir1.n16 GNDA 0.041731f
C832 bgr_0.V_mir1.n17 GNDA 0.028507f
C833 bgr_0.V_mir1.n18 GNDA 0.044354f
C834 bgr_0.V_mir1.n19 GNDA 0.111042f
C835 bgr_0.V_mir1.n20 GNDA 0.044166f
C836 bgr_0.V_mir1.t11 GNDA 0.019293f
C837 two_stage_opamp_dummy_magic_16_0.VD3.t28 GNDA 0.030951f
C838 two_stage_opamp_dummy_magic_16_0.VD3.t29 GNDA 0.030951f
C839 two_stage_opamp_dummy_magic_16_0.VD3.t23 GNDA 0.030951f
C840 two_stage_opamp_dummy_magic_16_0.VD3.n0 GNDA 0.108702f
C841 two_stage_opamp_dummy_magic_16_0.VD3.t21 GNDA 0.030951f
C842 two_stage_opamp_dummy_magic_16_0.VD3.t24 GNDA 0.030951f
C843 two_stage_opamp_dummy_magic_16_0.VD3.n1 GNDA 0.108329f
C844 two_stage_opamp_dummy_magic_16_0.VD3.n2 GNDA 0.202138f
C845 two_stage_opamp_dummy_magic_16_0.VD3.t26 GNDA 0.030951f
C846 two_stage_opamp_dummy_magic_16_0.VD3.t18 GNDA 0.030951f
C847 two_stage_opamp_dummy_magic_16_0.VD3.n3 GNDA 0.108329f
C848 two_stage_opamp_dummy_magic_16_0.VD3.n4 GNDA 0.104793f
C849 two_stage_opamp_dummy_magic_16_0.VD3.t19 GNDA 0.030951f
C850 two_stage_opamp_dummy_magic_16_0.VD3.t20 GNDA 0.030951f
C851 two_stage_opamp_dummy_magic_16_0.VD3.n5 GNDA 0.108329f
C852 two_stage_opamp_dummy_magic_16_0.VD3.n6 GNDA 0.104793f
C853 two_stage_opamp_dummy_magic_16_0.VD3.t22 GNDA 0.030951f
C854 two_stage_opamp_dummy_magic_16_0.VD3.t25 GNDA 0.030951f
C855 two_stage_opamp_dummy_magic_16_0.VD3.n7 GNDA 0.108329f
C856 two_stage_opamp_dummy_magic_16_0.VD3.n8 GNDA 0.104793f
C857 two_stage_opamp_dummy_magic_16_0.VD3.t5 GNDA 0.030951f
C858 two_stage_opamp_dummy_magic_16_0.VD3.t7 GNDA 0.030951f
C859 two_stage_opamp_dummy_magic_16_0.VD3.n9 GNDA 0.10726f
C860 two_stage_opamp_dummy_magic_16_0.VD3.n10 GNDA 0.104977f
C861 two_stage_opamp_dummy_magic_16_0.VD3.t35 GNDA 0.030951f
C862 two_stage_opamp_dummy_magic_16_0.VD3.n11 GNDA 0.092854f
C863 two_stage_opamp_dummy_magic_16_0.VD3.n12 GNDA 0.030951f
C864 two_stage_opamp_dummy_magic_16_0.VD3.n13 GNDA 0.017686f
C865 two_stage_opamp_dummy_magic_16_0.VD3.n15 GNDA 0.014321f
C866 two_stage_opamp_dummy_magic_16_0.VD3.n18 GNDA 0.014321f
C867 two_stage_opamp_dummy_magic_16_0.VD3.n19 GNDA 0.017686f
C868 two_stage_opamp_dummy_magic_16_0.VD3.t30 GNDA 0.054268f
C869 two_stage_opamp_dummy_magic_16_0.VD3.t1 GNDA 0.030951f
C870 two_stage_opamp_dummy_magic_16_0.VD3.t3 GNDA 0.030951f
C871 two_stage_opamp_dummy_magic_16_0.VD3.n20 GNDA 0.10726f
C872 two_stage_opamp_dummy_magic_16_0.VD3.n21 GNDA 0.104977f
C873 two_stage_opamp_dummy_magic_16_0.VD3.t11 GNDA 0.030951f
C874 two_stage_opamp_dummy_magic_16_0.VD3.t13 GNDA 0.030951f
C875 two_stage_opamp_dummy_magic_16_0.VD3.n22 GNDA 0.10726f
C876 two_stage_opamp_dummy_magic_16_0.VD3.n23 GNDA 0.104977f
C877 two_stage_opamp_dummy_magic_16_0.VD3.t17 GNDA 0.030951f
C878 two_stage_opamp_dummy_magic_16_0.VD3.t37 GNDA 0.030951f
C879 two_stage_opamp_dummy_magic_16_0.VD3.n24 GNDA 0.10726f
C880 two_stage_opamp_dummy_magic_16_0.VD3.n25 GNDA 0.104977f
C881 two_stage_opamp_dummy_magic_16_0.VD3.t15 GNDA 0.030951f
C882 two_stage_opamp_dummy_magic_16_0.VD3.t9 GNDA 0.030951f
C883 two_stage_opamp_dummy_magic_16_0.VD3.n26 GNDA 0.10726f
C884 two_stage_opamp_dummy_magic_16_0.VD3.n27 GNDA 0.134403f
C885 two_stage_opamp_dummy_magic_16_0.VD3.n28 GNDA 0.046089f
C886 two_stage_opamp_dummy_magic_16_0.VD3.t32 GNDA 0.030951f
C887 two_stage_opamp_dummy_magic_16_0.VD3.n29 GNDA 0.092854f
C888 two_stage_opamp_dummy_magic_16_0.VD3.n30 GNDA 0.031222f
C889 two_stage_opamp_dummy_magic_16_0.VD3.n31 GNDA 0.030951f
C890 two_stage_opamp_dummy_magic_16_0.VD3.n32 GNDA 0.017686f
C891 two_stage_opamp_dummy_magic_16_0.VD3.n33 GNDA 0.017686f
C892 two_stage_opamp_dummy_magic_16_0.VD3.n34 GNDA 0.030951f
C893 two_stage_opamp_dummy_magic_16_0.VD3.n36 GNDA 0.030951f
C894 two_stage_opamp_dummy_magic_16_0.VD3.n37 GNDA 0.017686f
C895 two_stage_opamp_dummy_magic_16_0.VD3.n38 GNDA 0.017686f
C896 two_stage_opamp_dummy_magic_16_0.VD3.n39 GNDA 0.030951f
C897 two_stage_opamp_dummy_magic_16_0.VD3.n41 GNDA 0.030951f
C898 two_stage_opamp_dummy_magic_16_0.VD3.n42 GNDA 0.029837f
C899 two_stage_opamp_dummy_magic_16_0.VD3.n43 GNDA 0.017686f
C900 two_stage_opamp_dummy_magic_16_0.VD3.n44 GNDA 0.258664f
C901 two_stage_opamp_dummy_magic_16_0.VD3.t31 GNDA 0.224175f
C902 two_stage_opamp_dummy_magic_16_0.VD3.t8 GNDA 0.206931f
C903 two_stage_opamp_dummy_magic_16_0.VD3.t14 GNDA 0.206931f
C904 two_stage_opamp_dummy_magic_16_0.VD3.t36 GNDA 0.206931f
C905 two_stage_opamp_dummy_magic_16_0.VD3.t16 GNDA 0.206931f
C906 two_stage_opamp_dummy_magic_16_0.VD3.t12 GNDA 0.206931f
C907 two_stage_opamp_dummy_magic_16_0.VD3.t10 GNDA 0.206931f
C908 two_stage_opamp_dummy_magic_16_0.VD3.t2 GNDA 0.206931f
C909 two_stage_opamp_dummy_magic_16_0.VD3.t0 GNDA 0.206931f
C910 two_stage_opamp_dummy_magic_16_0.VD3.t6 GNDA 0.206931f
C911 two_stage_opamp_dummy_magic_16_0.VD3.t4 GNDA 0.206931f
C912 two_stage_opamp_dummy_magic_16_0.VD3.t34 GNDA 0.224175f
C913 two_stage_opamp_dummy_magic_16_0.VD3.n45 GNDA 0.017686f
C914 two_stage_opamp_dummy_magic_16_0.VD3.n47 GNDA 0.031222f
C915 two_stage_opamp_dummy_magic_16_0.VD3.n48 GNDA 0.030951f
C916 two_stage_opamp_dummy_magic_16_0.VD3.n49 GNDA 0.017686f
C917 two_stage_opamp_dummy_magic_16_0.VD3.n50 GNDA 0.017686f
C918 two_stage_opamp_dummy_magic_16_0.VD3.n51 GNDA 0.030951f
C919 two_stage_opamp_dummy_magic_16_0.VD3.n53 GNDA 0.030951f
C920 two_stage_opamp_dummy_magic_16_0.VD3.n54 GNDA 0.030951f
C921 two_stage_opamp_dummy_magic_16_0.VD3.n55 GNDA 0.017686f
C922 two_stage_opamp_dummy_magic_16_0.VD3.n56 GNDA 0.258664f
C923 two_stage_opamp_dummy_magic_16_0.VD3.n57 GNDA 0.013727f
C924 two_stage_opamp_dummy_magic_16_0.VD3.n58 GNDA 0.033797f
C925 two_stage_opamp_dummy_magic_16_0.VD3.t33 GNDA 0.054268f
C926 two_stage_opamp_dummy_magic_16_0.VD3.n59 GNDA 0.044756f
C927 two_stage_opamp_dummy_magic_16_0.VD3.n60 GNDA 0.117031f
C928 two_stage_opamp_dummy_magic_16_0.VD3.n61 GNDA 0.19008f
C929 two_stage_opamp_dummy_magic_16_0.VD3.n62 GNDA 0.108328f
C930 two_stage_opamp_dummy_magic_16_0.VD3.t27 GNDA 0.030951f
C931 bgr_0.Vin+.t1 GNDA 0.173951f
C932 bgr_0.Vin+.t7 GNDA 0.010696f
C933 bgr_0.Vin+.t8 GNDA 0.025367f
C934 bgr_0.Vin+.t9 GNDA 0.01649f
C935 bgr_0.Vin+.n0 GNDA 0.054406f
C936 bgr_0.Vin+.t6 GNDA 0.01649f
C937 bgr_0.Vin+.n1 GNDA 0.042338f
C938 bgr_0.Vin+.t10 GNDA 0.01649f
C939 bgr_0.Vin+.n2 GNDA 0.042909f
C940 bgr_0.Vin+.n3 GNDA 0.130793f
C941 bgr_0.Vin+.t4 GNDA 0.05348f
C942 bgr_0.Vin+.t3 GNDA 0.05348f
C943 bgr_0.Vin+.n4 GNDA 0.176679f
C944 bgr_0.Vin+.n5 GNDA 1.27851f
C945 bgr_0.Vin+.t2 GNDA 0.05348f
C946 bgr_0.Vin+.t5 GNDA 0.05348f
C947 bgr_0.Vin+.n6 GNDA 0.176679f
C948 bgr_0.Vin+.n7 GNDA 1.06525f
C949 bgr_0.Vin+.n8 GNDA 1.7265f
C950 bgr_0.Vin+.t0 GNDA 0.232527f
C951 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t10 GNDA 0.010434f
C952 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t7 GNDA 0.010434f
C953 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n0 GNDA 0.02612f
C954 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t4 GNDA 0.010434f
C955 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t5 GNDA 0.010434f
C956 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n1 GNDA 0.02612f
C957 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t1 GNDA 0.010434f
C958 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t6 GNDA 0.010434f
C959 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n2 GNDA 0.02598f
C960 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n3 GNDA 0.17641f
C961 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n4 GNDA 0.148177f
C962 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t0 GNDA 0.010434f
C963 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t11 GNDA 0.010434f
C964 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n5 GNDA 0.020868f
C965 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n6 GNDA 0.03705f
C966 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t8 GNDA 0.015651f
C967 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t2 GNDA 0.015651f
C968 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n7 GNDA 0.053156f
C969 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t3 GNDA 0.015651f
C970 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t9 GNDA 0.015651f
C971 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n8 GNDA 0.031303f
C972 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t12 GNDA 0.027781f
C973 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t23 GNDA 0.027781f
C974 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t30 GNDA 0.027781f
C975 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t20 GNDA 0.027781f
C976 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t28 GNDA 0.027781f
C977 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t18 GNDA 0.027781f
C978 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t26 GNDA 0.027781f
C979 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t15 GNDA 0.027781f
C980 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t24 GNDA 0.027781f
C981 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t16 GNDA 0.032425f
C982 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n9 GNDA 0.030572f
C983 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n10 GNDA 0.019173f
C984 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n11 GNDA 0.019173f
C985 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n12 GNDA 0.019173f
C986 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n13 GNDA 0.019173f
C987 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n14 GNDA 0.019173f
C988 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n15 GNDA 0.019173f
C989 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n16 GNDA 0.019173f
C990 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n17 GNDA 0.017142f
C991 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t21 GNDA 0.027781f
C992 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t14 GNDA 0.027781f
C993 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t25 GNDA 0.027781f
C994 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t17 GNDA 0.027781f
C995 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t27 GNDA 0.027781f
C996 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t19 GNDA 0.027781f
C997 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t29 GNDA 0.027781f
C998 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t22 GNDA 0.027781f
C999 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t31 GNDA 0.027781f
C1000 two_stage_opamp_dummy_magic_16_0.V_tail_gate.t13 GNDA 0.032425f
C1001 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n18 GNDA 0.030572f
C1002 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n19 GNDA 0.019173f
C1003 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n20 GNDA 0.019173f
C1004 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n21 GNDA 0.019173f
C1005 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n22 GNDA 0.019173f
C1006 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n23 GNDA 0.019173f
C1007 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n24 GNDA 0.019173f
C1008 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n25 GNDA 0.019173f
C1009 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n26 GNDA 0.017142f
C1010 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n27 GNDA 0.044081f
C1011 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n28 GNDA 0.127865f
C1012 two_stage_opamp_dummy_magic_16_0.V_tail_gate.n29 GNDA 0.785356f
C1013 bgr_0.TAIL_CUR_MIR_BIAS GNDA 0.822673f
C1014 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t10 GNDA 0.042441f
C1015 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t7 GNDA 0.041727f
C1016 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n0 GNDA 0.302395f
C1017 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t6 GNDA 0.19488f
C1018 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t11 GNDA 0.030475f
C1019 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t8 GNDA 0.011396f
C1020 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n1 GNDA 0.035743f
C1021 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t13 GNDA 0.011396f
C1022 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n2 GNDA 0.029259f
C1023 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t9 GNDA 0.011396f
C1024 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n3 GNDA 0.029259f
C1025 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t12 GNDA 0.011396f
C1026 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n4 GNDA 0.050717f
C1027 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n5 GNDA 1.01397f
C1028 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t1 GNDA 0.036959f
C1029 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t4 GNDA 0.036959f
C1030 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n6 GNDA 0.130168f
C1031 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t5 GNDA 0.036959f
C1032 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t3 GNDA 0.036959f
C1033 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n7 GNDA 0.12385f
C1034 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n8 GNDA 0.578792f
C1035 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t2 GNDA 0.036959f
C1036 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.t0 GNDA 0.036959f
C1037 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n9 GNDA 0.12385f
C1038 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n10 GNDA 0.41388f
C1039 two_stage_opamp_dummy_magic_16_0.V_err_amp_ref.n11 GNDA 0.851096f
C1040 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t1 GNDA 0.105964f
C1041 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t3 GNDA 0.287618f
C1042 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t6 GNDA 0.265499f
C1043 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t7 GNDA 0.265499f
C1044 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t4 GNDA 0.315106f
C1045 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n0 GNDA 0.166436f
C1046 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n1 GNDA 0.105364f
C1047 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n2 GNDA 0.102722f
C1048 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n3 GNDA 0.485792f
C1049 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t8 GNDA 0.265499f
C1050 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t5 GNDA 0.265499f
C1051 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t9 GNDA 0.315106f
C1052 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n4 GNDA 0.166436f
C1053 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n5 GNDA 0.105364f
C1054 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t2 GNDA 0.287618f
C1055 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n6 GNDA 0.102722f
C1056 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.n7 GNDA 0.485792f
C1057 two_stage_opamp_dummy_magic_16_0.V_b_2nd_stage.t0 GNDA 0.105964f
C1058 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t13 GNDA 0.019639f
C1059 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t14 GNDA 0.019639f
C1060 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n0 GNDA 0.071382f
C1061 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t11 GNDA 0.019639f
C1062 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t12 GNDA 0.019639f
C1063 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n1 GNDA 0.059318f
C1064 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n2 GNDA 1.15698f
C1065 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t10 GNDA 0.241277f
C1066 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t4 GNDA 0.058917f
C1067 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t8 GNDA 0.058917f
C1068 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n3 GNDA 0.245765f
C1069 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t3 GNDA 0.058917f
C1070 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t2 GNDA 0.058917f
C1071 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n4 GNDA 0.244861f
C1072 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n5 GNDA 0.336177f
C1073 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t5 GNDA 0.058917f
C1074 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t9 GNDA 0.058917f
C1075 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n6 GNDA 0.244861f
C1076 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n7 GNDA 0.175414f
C1077 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t6 GNDA 0.058917f
C1078 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t0 GNDA 0.058917f
C1079 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n8 GNDA 0.244861f
C1080 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n9 GNDA 0.175414f
C1081 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t7 GNDA 0.058917f
C1082 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.t1 GNDA 0.058917f
C1083 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n10 GNDA 0.244861f
C1084 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n11 GNDA 0.243365f
C1085 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n12 GNDA 1.30797f
C1086 two_stage_opamp_dummy_magic_16_0.V_CMFB_S2.n13 GNDA 1.92994f
C1087 two_stage_opamp_dummy_magic_16_0.X.t6 GNDA 0.030949f
C1088 two_stage_opamp_dummy_magic_16_0.X.t10 GNDA 0.030949f
C1089 two_stage_opamp_dummy_magic_16_0.X.n0 GNDA 0.108693f
C1090 two_stage_opamp_dummy_magic_16_0.X.t24 GNDA 0.030949f
C1091 two_stage_opamp_dummy_magic_16_0.X.t15 GNDA 0.030949f
C1092 two_stage_opamp_dummy_magic_16_0.X.n1 GNDA 0.10832f
C1093 two_stage_opamp_dummy_magic_16_0.X.n2 GNDA 0.202123f
C1094 two_stage_opamp_dummy_magic_16_0.X.t14 GNDA 0.030949f
C1095 two_stage_opamp_dummy_magic_16_0.X.t18 GNDA 0.030949f
C1096 two_stage_opamp_dummy_magic_16_0.X.n3 GNDA 0.10832f
C1097 two_stage_opamp_dummy_magic_16_0.X.n4 GNDA 0.104785f
C1098 two_stage_opamp_dummy_magic_16_0.X.t1 GNDA 0.030949f
C1099 two_stage_opamp_dummy_magic_16_0.X.t8 GNDA 0.030949f
C1100 two_stage_opamp_dummy_magic_16_0.X.n5 GNDA 0.10832f
C1101 two_stage_opamp_dummy_magic_16_0.X.n6 GNDA 0.104785f
C1102 two_stage_opamp_dummy_magic_16_0.X.t4 GNDA 0.030949f
C1103 two_stage_opamp_dummy_magic_16_0.X.t0 GNDA 0.030949f
C1104 two_stage_opamp_dummy_magic_16_0.X.n7 GNDA 0.10832f
C1105 two_stage_opamp_dummy_magic_16_0.X.n8 GNDA 0.123419f
C1106 two_stage_opamp_dummy_magic_16_0.X.t7 GNDA 0.030949f
C1107 two_stage_opamp_dummy_magic_16_0.X.t3 GNDA 0.030949f
C1108 two_stage_opamp_dummy_magic_16_0.X.n9 GNDA 0.106149f
C1109 two_stage_opamp_dummy_magic_16_0.X.n10 GNDA 0.181464f
C1110 two_stage_opamp_dummy_magic_16_0.X.t37 GNDA 0.018569f
C1111 two_stage_opamp_dummy_magic_16_0.X.t50 GNDA 0.018569f
C1112 two_stage_opamp_dummy_magic_16_0.X.t33 GNDA 0.018569f
C1113 two_stage_opamp_dummy_magic_16_0.X.t47 GNDA 0.018569f
C1114 two_stage_opamp_dummy_magic_16_0.X.t30 GNDA 0.018569f
C1115 two_stage_opamp_dummy_magic_16_0.X.t44 GNDA 0.022549f
C1116 two_stage_opamp_dummy_magic_16_0.X.n11 GNDA 0.022549f
C1117 two_stage_opamp_dummy_magic_16_0.X.n12 GNDA 0.01459f
C1118 two_stage_opamp_dummy_magic_16_0.X.n13 GNDA 0.01459f
C1119 two_stage_opamp_dummy_magic_16_0.X.n14 GNDA 0.01459f
C1120 two_stage_opamp_dummy_magic_16_0.X.n15 GNDA 0.012869f
C1121 two_stage_opamp_dummy_magic_16_0.X.t54 GNDA 0.018569f
C1122 two_stage_opamp_dummy_magic_16_0.X.t28 GNDA 0.018569f
C1123 two_stage_opamp_dummy_magic_16_0.X.t53 GNDA 0.018569f
C1124 two_stage_opamp_dummy_magic_16_0.X.t39 GNDA 0.022549f
C1125 two_stage_opamp_dummy_magic_16_0.X.n16 GNDA 0.022549f
C1126 two_stage_opamp_dummy_magic_16_0.X.n17 GNDA 0.01459f
C1127 two_stage_opamp_dummy_magic_16_0.X.n18 GNDA 0.012869f
C1128 two_stage_opamp_dummy_magic_16_0.X.n19 GNDA 0.013372f
C1129 two_stage_opamp_dummy_magic_16_0.X.t25 GNDA 0.028517f
C1130 two_stage_opamp_dummy_magic_16_0.X.t38 GNDA 0.028517f
C1131 two_stage_opamp_dummy_magic_16_0.X.t52 GNDA 0.028517f
C1132 two_stage_opamp_dummy_magic_16_0.X.t36 GNDA 0.028517f
C1133 two_stage_opamp_dummy_magic_16_0.X.t49 GNDA 0.028517f
C1134 two_stage_opamp_dummy_magic_16_0.X.t32 GNDA 0.032419f
C1135 two_stage_opamp_dummy_magic_16_0.X.n20 GNDA 0.029258f
C1136 two_stage_opamp_dummy_magic_16_0.X.n21 GNDA 0.017906f
C1137 two_stage_opamp_dummy_magic_16_0.X.n22 GNDA 0.017906f
C1138 two_stage_opamp_dummy_magic_16_0.X.n23 GNDA 0.017906f
C1139 two_stage_opamp_dummy_magic_16_0.X.n24 GNDA 0.016185f
C1140 two_stage_opamp_dummy_magic_16_0.X.t41 GNDA 0.028517f
C1141 two_stage_opamp_dummy_magic_16_0.X.t46 GNDA 0.028517f
C1142 two_stage_opamp_dummy_magic_16_0.X.t40 GNDA 0.028517f
C1143 two_stage_opamp_dummy_magic_16_0.X.t26 GNDA 0.032419f
C1144 two_stage_opamp_dummy_magic_16_0.X.n25 GNDA 0.029258f
C1145 two_stage_opamp_dummy_magic_16_0.X.n26 GNDA 0.017906f
C1146 two_stage_opamp_dummy_magic_16_0.X.n27 GNDA 0.016185f
C1147 two_stage_opamp_dummy_magic_16_0.X.n28 GNDA 0.013372f
C1148 two_stage_opamp_dummy_magic_16_0.X.n29 GNDA 0.111621f
C1149 two_stage_opamp_dummy_magic_16_0.X.t23 GNDA 0.013264f
C1150 two_stage_opamp_dummy_magic_16_0.X.t19 GNDA 0.013264f
C1151 two_stage_opamp_dummy_magic_16_0.X.n30 GNDA 0.048484f
C1152 two_stage_opamp_dummy_magic_16_0.X.t11 GNDA 0.013264f
C1153 two_stage_opamp_dummy_magic_16_0.X.t16 GNDA 0.013264f
C1154 two_stage_opamp_dummy_magic_16_0.X.n31 GNDA 0.048081f
C1155 two_stage_opamp_dummy_magic_16_0.X.n32 GNDA 0.169595f
C1156 two_stage_opamp_dummy_magic_16_0.X.t2 GNDA 0.013264f
C1157 two_stage_opamp_dummy_magic_16_0.X.t17 GNDA 0.013264f
C1158 two_stage_opamp_dummy_magic_16_0.X.n33 GNDA 0.048081f
C1159 two_stage_opamp_dummy_magic_16_0.X.n34 GNDA 0.088094f
C1160 two_stage_opamp_dummy_magic_16_0.X.t21 GNDA 0.013264f
C1161 two_stage_opamp_dummy_magic_16_0.X.t12 GNDA 0.013264f
C1162 two_stage_opamp_dummy_magic_16_0.X.n35 GNDA 0.048081f
C1163 two_stage_opamp_dummy_magic_16_0.X.n36 GNDA 0.088094f
C1164 two_stage_opamp_dummy_magic_16_0.X.t9 GNDA 0.013264f
C1165 two_stage_opamp_dummy_magic_16_0.X.t22 GNDA 0.013264f
C1166 two_stage_opamp_dummy_magic_16_0.X.n37 GNDA 0.048081f
C1167 two_stage_opamp_dummy_magic_16_0.X.n38 GNDA 0.088094f
C1168 two_stage_opamp_dummy_magic_16_0.X.t20 GNDA 0.013264f
C1169 two_stage_opamp_dummy_magic_16_0.X.t5 GNDA 0.013264f
C1170 two_stage_opamp_dummy_magic_16_0.X.n39 GNDA 0.048081f
C1171 two_stage_opamp_dummy_magic_16_0.X.n40 GNDA 0.134054f
C1172 two_stage_opamp_dummy_magic_16_0.X.n41 GNDA 0.117902f
C1173 two_stage_opamp_dummy_magic_16_0.X.n42 GNDA 0.212185f
C1174 two_stage_opamp_dummy_magic_16_0.X.t31 GNDA 0.058361f
C1175 two_stage_opamp_dummy_magic_16_0.X.t45 GNDA 0.058361f
C1176 two_stage_opamp_dummy_magic_16_0.X.t29 GNDA 0.058361f
C1177 two_stage_opamp_dummy_magic_16_0.X.t43 GNDA 0.058361f
C1178 two_stage_opamp_dummy_magic_16_0.X.t27 GNDA 0.062158f
C1179 two_stage_opamp_dummy_magic_16_0.X.n43 GNDA 0.049258f
C1180 two_stage_opamp_dummy_magic_16_0.X.n44 GNDA 0.027854f
C1181 two_stage_opamp_dummy_magic_16_0.X.n45 GNDA 0.027854f
C1182 two_stage_opamp_dummy_magic_16_0.X.n46 GNDA 0.026139f
C1183 two_stage_opamp_dummy_magic_16_0.X.t48 GNDA 0.058361f
C1184 two_stage_opamp_dummy_magic_16_0.X.t35 GNDA 0.058361f
C1185 two_stage_opamp_dummy_magic_16_0.X.t42 GNDA 0.058361f
C1186 two_stage_opamp_dummy_magic_16_0.X.t34 GNDA 0.058361f
C1187 two_stage_opamp_dummy_magic_16_0.X.t51 GNDA 0.062158f
C1188 two_stage_opamp_dummy_magic_16_0.X.n47 GNDA 0.049258f
C1189 two_stage_opamp_dummy_magic_16_0.X.n48 GNDA 0.027854f
C1190 two_stage_opamp_dummy_magic_16_0.X.n49 GNDA 0.027854f
C1191 two_stage_opamp_dummy_magic_16_0.X.n50 GNDA 0.026139f
C1192 two_stage_opamp_dummy_magic_16_0.X.n51 GNDA 0.015901f
C1193 two_stage_opamp_dummy_magic_16_0.X.n52 GNDA 0.501906f
C1194 two_stage_opamp_dummy_magic_16_0.X.t13 GNDA 0.429924f
C1195 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t2 GNDA 0.345142f
C1196 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t80 GNDA 0.346293f
C1197 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t38 GNDA 0.186001f
C1198 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n0 GNDA 0.198613f
C1199 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t37 GNDA 0.345142f
C1200 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t124 GNDA 0.346293f
C1201 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t79 GNDA 0.186001f
C1202 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n1 GNDA 0.217197f
C1203 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t22 GNDA 0.345142f
C1204 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t100 GNDA 0.346293f
C1205 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t60 GNDA 0.186001f
C1206 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n2 GNDA 0.217197f
C1207 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t54 GNDA 0.345142f
C1208 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t131 GNDA 0.346293f
C1209 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t96 GNDA 0.186001f
C1210 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n3 GNDA 0.217197f
C1211 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t94 GNDA 0.345142f
C1212 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t42 GNDA 0.346293f
C1213 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t136 GNDA 0.364878f
C1214 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t32 GNDA 0.364878f
C1215 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t130 GNDA 0.186001f
C1216 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n4 GNDA 0.217197f
C1217 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t74 GNDA 0.345142f
C1218 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t97 GNDA 0.346293f
C1219 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t120 GNDA 0.364878f
C1220 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t13 GNDA 0.364878f
C1221 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t116 GNDA 0.186001f
C1222 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n5 GNDA 0.217197f
C1223 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t137 GNDA 0.346293f
C1224 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t102 GNDA 0.347548f
C1225 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t101 GNDA 0.346293f
C1226 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t61 GNDA 0.349008f
C1227 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t25 GNDA 0.379597f
C1228 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t126 GNDA 0.328964f
C1229 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t36 GNDA 0.346293f
C1230 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t1 GNDA 0.347548f
C1231 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t90 GNDA 0.328964f
C1232 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t5 GNDA 0.346293f
C1233 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t110 GNDA 0.347548f
C1234 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t26 GNDA 0.346293f
C1235 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t63 GNDA 0.347548f
C1236 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t39 GNDA 0.346293f
C1237 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t11 GNDA 0.347548f
C1238 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t68 GNDA 0.346293f
C1239 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t104 GNDA 0.347548f
C1240 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t81 GNDA 0.346293f
C1241 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t45 GNDA 0.347548f
C1242 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t30 GNDA 0.346293f
C1243 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t69 GNDA 0.347548f
C1244 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t47 GNDA 0.346293f
C1245 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t17 GNDA 0.347548f
C1246 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t73 GNDA 0.346293f
C1247 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t111 GNDA 0.347548f
C1248 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t89 GNDA 0.346293f
C1249 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t53 GNDA 0.347548f
C1250 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t115 GNDA 0.346293f
C1251 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t8 GNDA 0.347548f
C1252 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t127 GNDA 0.346293f
C1253 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t92 GNDA 0.347548f
C1254 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t76 GNDA 0.346293f
C1255 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t117 GNDA 0.347548f
C1256 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t93 GNDA 0.346293f
C1257 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t59 GNDA 0.347548f
C1258 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t121 GNDA 0.346293f
C1259 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t14 GNDA 0.347548f
C1260 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t129 GNDA 0.346293f
C1261 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t99 GNDA 0.347548f
C1262 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t20 GNDA 0.346293f
C1263 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t51 GNDA 0.347548f
C1264 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t31 GNDA 0.346293f
C1265 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t135 GNDA 0.347548f
C1266 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t55 GNDA 0.346293f
C1267 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t91 GNDA 0.347548f
C1268 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t75 GNDA 0.346293f
C1269 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t34 GNDA 0.347548f
C1270 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t23 GNDA 0.346293f
C1271 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t57 GNDA 0.347548f
C1272 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t35 GNDA 0.346293f
C1273 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t4 GNDA 0.347548f
C1274 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t62 GNDA 0.346293f
C1275 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t98 GNDA 0.347548f
C1276 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t78 GNDA 0.346293f
C1277 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t40 GNDA 0.347548f
C1278 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t103 GNDA 0.346293f
C1279 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t133 GNDA 0.347548f
C1280 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t123 GNDA 0.346293f
C1281 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t83 GNDA 0.347548f
C1282 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t108 GNDA 0.345142f
C1283 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t6 GNDA 0.346293f
C1284 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t72 GNDA 0.186001f
C1285 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n6 GNDA 0.198613f
C1286 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t138 GNDA 0.345142f
C1287 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t95 GNDA 0.346293f
C1288 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t109 GNDA 0.186001f
C1289 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n7 GNDA 0.217197f
C1290 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t49 GNDA 0.345142f
C1291 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t134 GNDA 0.346293f
C1292 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t19 GNDA 0.186001f
C1293 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n8 GNDA 0.217197f
C1294 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t84 GNDA 0.345142f
C1295 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t87 GNDA 0.346293f
C1296 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t50 GNDA 0.186001f
C1297 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n9 GNDA 0.217197f
C1298 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t125 GNDA 0.345142f
C1299 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t33 GNDA 0.346293f
C1300 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t86 GNDA 0.186001f
C1301 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n10 GNDA 0.217197f
C1302 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t29 GNDA 0.345142f
C1303 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t77 GNDA 0.346293f
C1304 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t132 GNDA 0.186001f
C1305 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n11 GNDA 0.217197f
C1306 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t67 GNDA 0.345142f
C1307 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t27 GNDA 0.346293f
C1308 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t28 GNDA 0.186001f
C1309 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n12 GNDA 0.217197f
C1310 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t119 GNDA 0.346293f
C1311 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t70 GNDA 0.186001f
C1312 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n13 GNDA 0.197462f
C1313 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t66 GNDA 0.346293f
C1314 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t105 GNDA 0.186001f
C1315 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n14 GNDA 0.197462f
C1316 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t82 GNDA 0.346293f
C1317 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t46 GNDA 0.347548f
C1318 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t7 GNDA 0.346293f
C1319 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t56 GNDA 0.347548f
C1320 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t112 GNDA 0.167416f
C1321 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n15 GNDA 0.215942f
C1322 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t16 GNDA 0.18485f
C1323 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n16 GNDA 0.234527f
C1324 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t43 GNDA 0.18485f
C1325 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n17 GNDA 0.251856f
C1326 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t9 GNDA 0.18485f
C1327 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n18 GNDA 0.251856f
C1328 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t113 GNDA 0.18485f
C1329 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n19 GNDA 0.251856f
C1330 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t3 GNDA 0.18485f
C1331 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n20 GNDA 0.251856f
C1332 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t106 GNDA 0.18485f
C1333 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n21 GNDA 0.251856f
C1334 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t64 GNDA 0.18485f
C1335 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n22 GNDA 0.251856f
C1336 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t24 GNDA 0.18485f
C1337 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n23 GNDA 0.251856f
C1338 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t58 GNDA 0.18485f
C1339 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n24 GNDA 0.251856f
C1340 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t21 GNDA 0.18485f
C1341 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n25 GNDA 0.251856f
C1342 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t122 GNDA 0.18485f
C1343 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n26 GNDA 0.251856f
C1344 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t15 GNDA 0.18485f
C1345 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n27 GNDA 0.251856f
C1346 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t118 GNDA 0.18485f
C1347 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n28 GNDA 0.251856f
C1348 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t71 GNDA 0.18485f
C1349 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n29 GNDA 0.251856f
C1350 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t107 GNDA 0.18485f
C1351 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n30 GNDA 0.251856f
C1352 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t65 GNDA 0.18485f
C1353 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n31 GNDA 0.234527f
C1354 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t41 GNDA 0.345142f
C1355 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t85 GNDA 0.167416f
C1356 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n32 GNDA 0.217197f
C1357 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t10 GNDA 0.345142f
C1358 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t52 GNDA 0.346293f
C1359 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t88 GNDA 0.364878f
C1360 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t44 GNDA 0.186001f
C1361 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n33 GNDA 0.217197f
C1362 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t114 GNDA 0.345142f
C1363 two_stage_opamp_dummy_magic_16_0.cap_res_Y.n34 GNDA 0.217197f
C1364 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t12 GNDA 0.186001f
C1365 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t48 GNDA 0.364878f
C1366 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t18 GNDA 0.364878f
C1367 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t128 GNDA 0.730561f
C1368 two_stage_opamp_dummy_magic_16_0.cap_res_Y.t0 GNDA 0.29977f
C1369 VOUT+.t10 GNDA 0.048668f
C1370 VOUT+.t15 GNDA 0.048668f
C1371 VOUT+.n0 GNDA 0.225914f
C1372 VOUT+.t18 GNDA 0.048668f
C1373 VOUT+.t6 GNDA 0.048668f
C1374 VOUT+.n1 GNDA 0.225185f
C1375 VOUT+.n2 GNDA 0.138481f
C1376 VOUT+.t16 GNDA 0.048668f
C1377 VOUT+.t9 GNDA 0.048668f
C1378 VOUT+.n3 GNDA 0.225185f
C1379 VOUT+.n4 GNDA 0.077142f
C1380 VOUT+.t5 GNDA 0.081011f
C1381 VOUT+.n5 GNDA 0.091611f
C1382 VOUT+.t11 GNDA 0.041716f
C1383 VOUT+.t14 GNDA 0.041716f
C1384 VOUT+.n6 GNDA 0.168663f
C1385 VOUT+.t0 GNDA 0.041716f
C1386 VOUT+.t8 GNDA 0.041716f
C1387 VOUT+.n7 GNDA 0.168362f
C1388 VOUT+.n8 GNDA 0.164256f
C1389 VOUT+.t2 GNDA 0.041716f
C1390 VOUT+.t1 GNDA 0.041716f
C1391 VOUT+.n9 GNDA 0.168362f
C1392 VOUT+.n10 GNDA 0.084712f
C1393 VOUT+.t3 GNDA 0.041716f
C1394 VOUT+.t17 GNDA 0.041716f
C1395 VOUT+.n11 GNDA 0.168362f
C1396 VOUT+.n12 GNDA 0.084712f
C1397 VOUT+.t7 GNDA 0.041716f
C1398 VOUT+.t12 GNDA 0.041716f
C1399 VOUT+.n13 GNDA 0.168663f
C1400 VOUT+.n14 GNDA 0.100402f
C1401 VOUT+.t4 GNDA 0.041716f
C1402 VOUT+.t13 GNDA 0.041716f
C1403 VOUT+.n15 GNDA 0.166369f
C1404 VOUT+.n16 GNDA 0.14091f
C1405 VOUT+.t45 GNDA 0.278104f
C1406 VOUT+.t150 GNDA 0.28284f
C1407 VOUT+.t101 GNDA 0.278104f
C1408 VOUT+.n17 GNDA 0.186459f
C1409 VOUT+.n18 GNDA 0.12167f
C1410 VOUT+.t91 GNDA 0.282247f
C1411 VOUT+.t38 GNDA 0.282247f
C1412 VOUT+.t130 GNDA 0.282247f
C1413 VOUT+.t90 GNDA 0.282247f
C1414 VOUT+.t80 GNDA 0.282247f
C1415 VOUT+.t128 GNDA 0.282247f
C1416 VOUT+.t124 GNDA 0.282247f
C1417 VOUT+.t32 GNDA 0.282247f
C1418 VOUT+.t70 GNDA 0.282247f
C1419 VOUT+.t73 GNDA 0.282247f
C1420 VOUT+.t23 GNDA 0.282247f
C1421 VOUT+.t108 GNDA 0.282247f
C1422 VOUT+.t62 GNDA 0.282247f
C1423 VOUT+.t19 GNDA 0.282247f
C1424 VOUT+.t151 GNDA 0.282247f
C1425 VOUT+.t49 GNDA 0.282247f
C1426 VOUT+.t85 GNDA 0.278104f
C1427 VOUT+.n19 GNDA 0.304579f
C1428 VOUT+.t48 GNDA 0.278104f
C1429 VOUT+.n20 GNDA 0.356724f
C1430 VOUT+.t138 GNDA 0.278104f
C1431 VOUT+.n21 GNDA 0.356724f
C1432 VOUT+.t107 GNDA 0.278104f
C1433 VOUT+.n22 GNDA 0.356724f
C1434 VOUT+.t71 GNDA 0.278104f
C1435 VOUT+.n23 GNDA 0.356724f
C1436 VOUT+.t25 GNDA 0.278104f
C1437 VOUT+.n24 GNDA 0.356724f
C1438 VOUT+.t129 GNDA 0.278104f
C1439 VOUT+.n25 GNDA 0.356724f
C1440 VOUT+.t87 GNDA 0.278104f
C1441 VOUT+.n26 GNDA 0.239197f
C1442 VOUT+.t52 GNDA 0.278104f
C1443 VOUT+.n27 GNDA 0.239197f
C1444 VOUT+.t141 GNDA 0.278104f
C1445 VOUT+.t75 GNDA 0.28284f
C1446 VOUT+.t111 GNDA 0.278104f
C1447 VOUT+.n28 GNDA 0.186459f
C1448 VOUT+.n29 GNDA 0.225959f
C1449 VOUT+.t54 GNDA 0.28284f
C1450 VOUT+.t24 GNDA 0.278104f
C1451 VOUT+.n30 GNDA 0.186459f
C1452 VOUT+.t114 GNDA 0.278104f
C1453 VOUT+.t34 GNDA 0.28284f
C1454 VOUT+.t74 GNDA 0.278104f
C1455 VOUT+.n31 GNDA 0.186459f
C1456 VOUT+.n32 GNDA 0.225959f
C1457 VOUT+.t95 GNDA 0.28284f
C1458 VOUT+.t59 GNDA 0.278104f
C1459 VOUT+.n33 GNDA 0.186459f
C1460 VOUT+.t148 GNDA 0.278104f
C1461 VOUT+.t79 GNDA 0.28284f
C1462 VOUT+.t117 GNDA 0.278104f
C1463 VOUT+.n34 GNDA 0.186459f
C1464 VOUT+.n35 GNDA 0.225959f
C1465 VOUT+.t134 GNDA 0.28284f
C1466 VOUT+.t100 GNDA 0.278104f
C1467 VOUT+.n36 GNDA 0.186459f
C1468 VOUT+.t44 GNDA 0.278104f
C1469 VOUT+.t122 GNDA 0.28284f
C1470 VOUT+.t153 GNDA 0.278104f
C1471 VOUT+.n37 GNDA 0.186459f
C1472 VOUT+.n38 GNDA 0.225959f
C1473 VOUT+.t102 GNDA 0.28284f
C1474 VOUT+.t66 GNDA 0.278104f
C1475 VOUT+.n39 GNDA 0.186459f
C1476 VOUT+.t154 GNDA 0.278104f
C1477 VOUT+.t82 GNDA 0.28284f
C1478 VOUT+.t123 GNDA 0.278104f
C1479 VOUT+.n40 GNDA 0.186459f
C1480 VOUT+.n41 GNDA 0.225959f
C1481 VOUT+.t137 GNDA 0.28284f
C1482 VOUT+.t106 GNDA 0.278104f
C1483 VOUT+.n42 GNDA 0.186459f
C1484 VOUT+.t51 GNDA 0.278104f
C1485 VOUT+.t126 GNDA 0.28284f
C1486 VOUT+.t22 GNDA 0.278104f
C1487 VOUT+.n43 GNDA 0.186459f
C1488 VOUT+.n44 GNDA 0.225959f
C1489 VOUT+.t132 GNDA 0.278104f
C1490 VOUT+.t56 GNDA 0.28284f
C1491 VOUT+.t96 GNDA 0.278104f
C1492 VOUT+.n45 GNDA 0.186459f
C1493 VOUT+.n46 GNDA 0.12167f
C1494 VOUT+.t116 GNDA 0.282247f
C1495 VOUT+.t105 GNDA 0.28284f
C1496 VOUT+.t69 GNDA 0.278104f
C1497 VOUT+.n47 GNDA 0.182114f
C1498 VOUT+.t147 GNDA 0.282247f
C1499 VOUT+.t29 GNDA 0.28284f
C1500 VOUT+.t139 GNDA 0.278104f
C1501 VOUT+.n48 GNDA 0.186459f
C1502 VOUT+.t109 GNDA 0.278104f
C1503 VOUT+.n49 GNDA 0.117325f
C1504 VOUT+.t43 GNDA 0.282247f
C1505 VOUT+.t60 GNDA 0.28284f
C1506 VOUT+.t37 GNDA 0.278104f
C1507 VOUT+.n50 GNDA 0.186459f
C1508 VOUT+.t144 GNDA 0.278104f
C1509 VOUT+.n51 GNDA 0.117325f
C1510 VOUT+.t83 GNDA 0.282247f
C1511 VOUT+.t115 GNDA 0.28284f
C1512 VOUT+.t21 GNDA 0.278104f
C1513 VOUT+.n52 GNDA 0.186459f
C1514 VOUT+.t125 GNDA 0.278104f
C1515 VOUT+.n53 GNDA 0.117325f
C1516 VOUT+.t63 GNDA 0.282247f
C1517 VOUT+.t26 GNDA 0.282247f
C1518 VOUT+.t103 GNDA 0.282247f
C1519 VOUT+.t57 GNDA 0.28248f
C1520 VOUT+.t135 GNDA 0.282247f
C1521 VOUT+.t33 GNDA 0.28248f
C1522 VOUT+.t120 GNDA 0.282247f
C1523 VOUT+.t77 GNDA 0.28248f
C1524 VOUT+.t155 GNDA 0.282247f
C1525 VOUT+.t119 GNDA 0.278104f
C1526 VOUT+.n54 GNDA 0.307823f
C1527 VOUT+.t78 GNDA 0.278104f
C1528 VOUT+.n55 GNDA 0.359967f
C1529 VOUT+.t97 GNDA 0.278104f
C1530 VOUT+.n56 GNDA 0.359967f
C1531 VOUT+.t61 GNDA 0.278104f
C1532 VOUT+.n57 GNDA 0.356724f
C1533 VOUT+.t27 GNDA 0.278104f
C1534 VOUT+.n58 GNDA 0.295687f
C1535 VOUT+.t41 GNDA 0.278104f
C1536 VOUT+.n59 GNDA 0.295687f
C1537 VOUT+.t145 GNDA 0.278104f
C1538 VOUT+.n60 GNDA 0.295687f
C1539 VOUT+.t113 GNDA 0.278104f
C1540 VOUT+.n61 GNDA 0.295687f
C1541 VOUT+.t72 GNDA 0.278104f
C1542 VOUT+.n62 GNDA 0.239197f
C1543 VOUT+.t92 GNDA 0.278104f
C1544 VOUT+.t20 GNDA 0.28284f
C1545 VOUT+.t55 GNDA 0.278104f
C1546 VOUT+.n63 GNDA 0.186459f
C1547 VOUT+.n64 GNDA 0.225959f
C1548 VOUT+.t31 GNDA 0.28284f
C1549 VOUT+.t50 GNDA 0.278104f
C1550 VOUT+.t121 GNDA 0.28284f
C1551 VOUT+.t156 GNDA 0.278104f
C1552 VOUT+.n65 GNDA 0.186459f
C1553 VOUT+.n66 GNDA 0.290748f
C1554 VOUT+.t67 GNDA 0.28284f
C1555 VOUT+.t86 GNDA 0.278104f
C1556 VOUT+.t152 GNDA 0.28284f
C1557 VOUT+.t47 GNDA 0.278104f
C1558 VOUT+.n67 GNDA 0.186459f
C1559 VOUT+.n68 GNDA 0.290748f
C1560 VOUT+.t131 GNDA 0.28284f
C1561 VOUT+.t94 GNDA 0.278104f
C1562 VOUT+.n69 GNDA 0.186459f
C1563 VOUT+.t39 GNDA 0.278104f
C1564 VOUT+.t118 GNDA 0.28284f
C1565 VOUT+.t146 GNDA 0.278104f
C1566 VOUT+.n70 GNDA 0.186459f
C1567 VOUT+.n71 GNDA 0.225959f
C1568 VOUT+.t89 GNDA 0.28284f
C1569 VOUT+.t53 GNDA 0.278104f
C1570 VOUT+.n72 GNDA 0.186459f
C1571 VOUT+.t142 GNDA 0.278104f
C1572 VOUT+.t76 GNDA 0.28284f
C1573 VOUT+.t112 GNDA 0.278104f
C1574 VOUT+.n73 GNDA 0.186459f
C1575 VOUT+.n74 GNDA 0.225959f
C1576 VOUT+.t127 GNDA 0.28284f
C1577 VOUT+.t88 GNDA 0.278104f
C1578 VOUT+.n75 GNDA 0.186459f
C1579 VOUT+.t35 GNDA 0.278104f
C1580 VOUT+.t110 GNDA 0.28284f
C1581 VOUT+.t140 GNDA 0.278104f
C1582 VOUT+.n76 GNDA 0.186459f
C1583 VOUT+.n77 GNDA 0.225959f
C1584 VOUT+.t84 GNDA 0.28284f
C1585 VOUT+.t46 GNDA 0.278104f
C1586 VOUT+.n78 GNDA 0.186459f
C1587 VOUT+.t136 GNDA 0.278104f
C1588 VOUT+.t68 GNDA 0.28284f
C1589 VOUT+.t104 GNDA 0.278104f
C1590 VOUT+.n79 GNDA 0.186459f
C1591 VOUT+.n80 GNDA 0.225959f
C1592 VOUT+.t42 GNDA 0.28284f
C1593 VOUT+.t149 GNDA 0.278104f
C1594 VOUT+.n81 GNDA 0.186459f
C1595 VOUT+.t99 GNDA 0.278104f
C1596 VOUT+.t30 GNDA 0.28284f
C1597 VOUT+.t65 GNDA 0.278104f
C1598 VOUT+.n82 GNDA 0.186459f
C1599 VOUT+.n83 GNDA 0.225959f
C1600 VOUT+.t81 GNDA 0.28284f
C1601 VOUT+.t40 GNDA 0.278104f
C1602 VOUT+.n84 GNDA 0.186459f
C1603 VOUT+.t133 GNDA 0.278104f
C1604 VOUT+.t64 GNDA 0.28284f
C1605 VOUT+.t98 GNDA 0.278104f
C1606 VOUT+.n85 GNDA 0.186459f
C1607 VOUT+.n86 GNDA 0.225959f
C1608 VOUT+.t28 GNDA 0.28284f
C1609 VOUT+.t58 GNDA 0.278104f
C1610 VOUT+.n87 GNDA 0.186459f
C1611 VOUT+.t93 GNDA 0.278104f
C1612 VOUT+.n88 GNDA 0.225959f
C1613 VOUT+.t143 GNDA 0.278104f
C1614 VOUT+.n89 GNDA 0.12167f
C1615 VOUT+.t36 GNDA 0.278104f
C1616 VOUT+.n90 GNDA 0.177423f
C1617 VOUT+.n91 GNDA 0.210673f
C1618 two_stage_opamp_dummy_magic_16_0.cap_res_X.t128 GNDA 0.346251f
C1619 two_stage_opamp_dummy_magic_16_0.cap_res_X.t105 GNDA 0.347506f
C1620 two_stage_opamp_dummy_magic_16_0.cap_res_X.t89 GNDA 0.346251f
C1621 two_stage_opamp_dummy_magic_16_0.cap_res_X.t71 GNDA 0.348966f
C1622 two_stage_opamp_dummy_magic_16_0.cap_res_X.t103 GNDA 0.379551f
C1623 two_stage_opamp_dummy_magic_16_0.cap_res_X.t32 GNDA 0.346251f
C1624 two_stage_opamp_dummy_magic_16_0.cap_res_X.t5 GNDA 0.347506f
C1625 two_stage_opamp_dummy_magic_16_0.cap_res_X.t84 GNDA 0.328924f
C1626 two_stage_opamp_dummy_magic_16_0.cap_res_X.t134 GNDA 0.346251f
C1627 two_stage_opamp_dummy_magic_16_0.cap_res_X.t110 GNDA 0.347506f
C1628 two_stage_opamp_dummy_magic_16_0.cap_res_X.t48 GNDA 0.328924f
C1629 two_stage_opamp_dummy_magic_16_0.cap_res_X.t81 GNDA 0.346251f
C1630 two_stage_opamp_dummy_magic_16_0.cap_res_X.t130 GNDA 0.347506f
C1631 two_stage_opamp_dummy_magic_16_0.cap_res_X.t113 GNDA 0.346251f
C1632 two_stage_opamp_dummy_magic_16_0.cap_res_X.t60 GNDA 0.347506f
C1633 two_stage_opamp_dummy_magic_16_0.cap_res_X.t120 GNDA 0.346251f
C1634 two_stage_opamp_dummy_magic_16_0.cap_res_X.t34 GNDA 0.347506f
C1635 two_stage_opamp_dummy_magic_16_0.cap_res_X.t14 GNDA 0.346251f
C1636 two_stage_opamp_dummy_magic_16_0.cap_res_X.t100 GNDA 0.347506f
C1637 two_stage_opamp_dummy_magic_16_0.cap_res_X.t87 GNDA 0.346251f
C1638 two_stage_opamp_dummy_magic_16_0.cap_res_X.t137 GNDA 0.347506f
C1639 two_stage_opamp_dummy_magic_16_0.cap_res_X.t118 GNDA 0.346251f
C1640 two_stage_opamp_dummy_magic_16_0.cap_res_X.t70 GNDA 0.347506f
C1641 two_stage_opamp_dummy_magic_16_0.cap_res_X.t125 GNDA 0.346251f
C1642 two_stage_opamp_dummy_magic_16_0.cap_res_X.t39 GNDA 0.347506f
C1643 two_stage_opamp_dummy_magic_16_0.cap_res_X.t19 GNDA 0.346251f
C1644 two_stage_opamp_dummy_magic_16_0.cap_res_X.t104 GNDA 0.347506f
C1645 two_stage_opamp_dummy_magic_16_0.cap_res_X.t26 GNDA 0.346251f
C1646 two_stage_opamp_dummy_magic_16_0.cap_res_X.t78 GNDA 0.347506f
C1647 two_stage_opamp_dummy_magic_16_0.cap_res_X.t56 GNDA 0.346251f
C1648 two_stage_opamp_dummy_magic_16_0.cap_res_X.t4 GNDA 0.347506f
C1649 two_stage_opamp_dummy_magic_16_0.cap_res_X.t129 GNDA 0.346251f
C1650 two_stage_opamp_dummy_magic_16_0.cap_res_X.t40 GNDA 0.347506f
C1651 two_stage_opamp_dummy_magic_16_0.cap_res_X.t24 GNDA 0.346251f
C1652 two_stage_opamp_dummy_magic_16_0.cap_res_X.t111 GNDA 0.347506f
C1653 two_stage_opamp_dummy_magic_16_0.cap_res_X.t33 GNDA 0.346251f
C1654 two_stage_opamp_dummy_magic_16_0.cap_res_X.t82 GNDA 0.347506f
C1655 two_stage_opamp_dummy_magic_16_0.cap_res_X.t61 GNDA 0.346251f
C1656 two_stage_opamp_dummy_magic_16_0.cap_res_X.t12 GNDA 0.347506f
C1657 two_stage_opamp_dummy_magic_16_0.cap_res_X.t72 GNDA 0.346251f
C1658 two_stage_opamp_dummy_magic_16_0.cap_res_X.t123 GNDA 0.347506f
C1659 two_stage_opamp_dummy_magic_16_0.cap_res_X.t102 GNDA 0.346251f
C1660 two_stage_opamp_dummy_magic_16_0.cap_res_X.t51 GNDA 0.347506f
C1661 two_stage_opamp_dummy_magic_16_0.cap_res_X.t108 GNDA 0.346251f
C1662 two_stage_opamp_dummy_magic_16_0.cap_res_X.t22 GNDA 0.347506f
C1663 two_stage_opamp_dummy_magic_16_0.cap_res_X.t138 GNDA 0.346251f
C1664 two_stage_opamp_dummy_magic_16_0.cap_res_X.t90 GNDA 0.347506f
C1665 two_stage_opamp_dummy_magic_16_0.cap_res_X.t77 GNDA 0.346251f
C1666 two_stage_opamp_dummy_magic_16_0.cap_res_X.t127 GNDA 0.347506f
C1667 two_stage_opamp_dummy_magic_16_0.cap_res_X.t106 GNDA 0.346251f
C1668 two_stage_opamp_dummy_magic_16_0.cap_res_X.t54 GNDA 0.347506f
C1669 two_stage_opamp_dummy_magic_16_0.cap_res_X.t116 GNDA 0.346251f
C1670 two_stage_opamp_dummy_magic_16_0.cap_res_X.t28 GNDA 0.347506f
C1671 two_stage_opamp_dummy_magic_16_0.cap_res_X.t6 GNDA 0.346251f
C1672 two_stage_opamp_dummy_magic_16_0.cap_res_X.t94 GNDA 0.347506f
C1673 two_stage_opamp_dummy_magic_16_0.cap_res_X.t17 GNDA 0.346251f
C1674 two_stage_opamp_dummy_magic_16_0.cap_res_X.t68 GNDA 0.347506f
C1675 two_stage_opamp_dummy_magic_16_0.cap_res_X.t46 GNDA 0.346251f
C1676 two_stage_opamp_dummy_magic_16_0.cap_res_X.t136 GNDA 0.347506f
C1677 two_stage_opamp_dummy_magic_16_0.cap_res_X.t121 GNDA 0.346251f
C1678 two_stage_opamp_dummy_magic_16_0.cap_res_X.t35 GNDA 0.347506f
C1679 two_stage_opamp_dummy_magic_16_0.cap_res_X.t44 GNDA 0.3451f
C1680 two_stage_opamp_dummy_magic_16_0.cap_res_X.t86 GNDA 0.346251f
C1681 two_stage_opamp_dummy_magic_16_0.cap_res_X.t9 GNDA 0.185978f
C1682 two_stage_opamp_dummy_magic_16_0.cap_res_X.n0 GNDA 0.198589f
C1683 two_stage_opamp_dummy_magic_16_0.cap_res_X.t133 GNDA 0.3451f
C1684 two_stage_opamp_dummy_magic_16_0.cap_res_X.t43 GNDA 0.346251f
C1685 two_stage_opamp_dummy_magic_16_0.cap_res_X.t97 GNDA 0.185978f
C1686 two_stage_opamp_dummy_magic_16_0.cap_res_X.n1 GNDA 0.217171f
C1687 two_stage_opamp_dummy_magic_16_0.cap_res_X.t95 GNDA 0.3451f
C1688 two_stage_opamp_dummy_magic_16_0.cap_res_X.t92 GNDA 0.346251f
C1689 two_stage_opamp_dummy_magic_16_0.cap_res_X.t64 GNDA 0.185978f
C1690 two_stage_opamp_dummy_magic_16_0.cap_res_X.n2 GNDA 0.217171f
C1691 two_stage_opamp_dummy_magic_16_0.cap_res_X.t62 GNDA 0.3451f
C1692 two_stage_opamp_dummy_magic_16_0.cap_res_X.t3 GNDA 0.346251f
C1693 two_stage_opamp_dummy_magic_16_0.cap_res_X.t30 GNDA 0.185978f
C1694 two_stage_opamp_dummy_magic_16_0.cap_res_X.n3 GNDA 0.217171f
C1695 two_stage_opamp_dummy_magic_16_0.cap_res_X.t31 GNDA 0.3451f
C1696 two_stage_opamp_dummy_magic_16_0.cap_res_X.t52 GNDA 0.346251f
C1697 two_stage_opamp_dummy_magic_16_0.cap_res_X.t132 GNDA 0.185978f
C1698 two_stage_opamp_dummy_magic_16_0.cap_res_X.n4 GNDA 0.217171f
C1699 two_stage_opamp_dummy_magic_16_0.cap_res_X.t119 GNDA 0.3451f
C1700 two_stage_opamp_dummy_magic_16_0.cap_res_X.t16 GNDA 0.346251f
C1701 two_stage_opamp_dummy_magic_16_0.cap_res_X.t85 GNDA 0.185978f
C1702 two_stage_opamp_dummy_magic_16_0.cap_res_X.n5 GNDA 0.217171f
C1703 two_stage_opamp_dummy_magic_16_0.cap_res_X.t83 GNDA 0.3451f
C1704 two_stage_opamp_dummy_magic_16_0.cap_res_X.t65 GNDA 0.346251f
C1705 two_stage_opamp_dummy_magic_16_0.cap_res_X.t47 GNDA 0.185978f
C1706 two_stage_opamp_dummy_magic_16_0.cap_res_X.n6 GNDA 0.217171f
C1707 two_stage_opamp_dummy_magic_16_0.cap_res_X.t115 GNDA 0.346251f
C1708 two_stage_opamp_dummy_magic_16_0.cap_res_X.t15 GNDA 0.185978f
C1709 two_stage_opamp_dummy_magic_16_0.cap_res_X.n7 GNDA 0.197438f
C1710 two_stage_opamp_dummy_magic_16_0.cap_res_X.t75 GNDA 0.346251f
C1711 two_stage_opamp_dummy_magic_16_0.cap_res_X.t101 GNDA 0.185978f
C1712 two_stage_opamp_dummy_magic_16_0.cap_res_X.n8 GNDA 0.197438f
C1713 two_stage_opamp_dummy_magic_16_0.cap_res_X.t131 GNDA 0.346251f
C1714 two_stage_opamp_dummy_magic_16_0.cap_res_X.t38 GNDA 0.347506f
C1715 two_stage_opamp_dummy_magic_16_0.cap_res_X.t124 GNDA 0.167396f
C1716 two_stage_opamp_dummy_magic_16_0.cap_res_X.n9 GNDA 0.215916f
C1717 two_stage_opamp_dummy_magic_16_0.cap_res_X.t67 GNDA 0.184828f
C1718 two_stage_opamp_dummy_magic_16_0.cap_res_X.n10 GNDA 0.234498f
C1719 two_stage_opamp_dummy_magic_16_0.cap_res_X.t98 GNDA 0.184828f
C1720 two_stage_opamp_dummy_magic_16_0.cap_res_X.n11 GNDA 0.251826f
C1721 two_stage_opamp_dummy_magic_16_0.cap_res_X.t59 GNDA 0.184828f
C1722 two_stage_opamp_dummy_magic_16_0.cap_res_X.n12 GNDA 0.251826f
C1723 two_stage_opamp_dummy_magic_16_0.cap_res_X.t23 GNDA 0.184828f
C1724 two_stage_opamp_dummy_magic_16_0.cap_res_X.n13 GNDA 0.251826f
C1725 two_stage_opamp_dummy_magic_16_0.cap_res_X.t55 GNDA 0.184828f
C1726 two_stage_opamp_dummy_magic_16_0.cap_res_X.n14 GNDA 0.251826f
C1727 two_stage_opamp_dummy_magic_16_0.cap_res_X.t18 GNDA 0.184828f
C1728 two_stage_opamp_dummy_magic_16_0.cap_res_X.n15 GNDA 0.251826f
C1729 two_stage_opamp_dummy_magic_16_0.cap_res_X.t117 GNDA 0.184828f
C1730 two_stage_opamp_dummy_magic_16_0.cap_res_X.n16 GNDA 0.251826f
C1731 two_stage_opamp_dummy_magic_16_0.cap_res_X.t79 GNDA 0.184828f
C1732 two_stage_opamp_dummy_magic_16_0.cap_res_X.n17 GNDA 0.251826f
C1733 two_stage_opamp_dummy_magic_16_0.cap_res_X.t109 GNDA 0.184828f
C1734 two_stage_opamp_dummy_magic_16_0.cap_res_X.n18 GNDA 0.251826f
C1735 two_stage_opamp_dummy_magic_16_0.cap_res_X.t73 GNDA 0.184828f
C1736 two_stage_opamp_dummy_magic_16_0.cap_res_X.n19 GNDA 0.251826f
C1737 two_stage_opamp_dummy_magic_16_0.cap_res_X.t36 GNDA 0.184828f
C1738 two_stage_opamp_dummy_magic_16_0.cap_res_X.n20 GNDA 0.251826f
C1739 two_stage_opamp_dummy_magic_16_0.cap_res_X.t69 GNDA 0.184828f
C1740 two_stage_opamp_dummy_magic_16_0.cap_res_X.n21 GNDA 0.251826f
C1741 two_stage_opamp_dummy_magic_16_0.cap_res_X.t29 GNDA 0.184828f
C1742 two_stage_opamp_dummy_magic_16_0.cap_res_X.n22 GNDA 0.251826f
C1743 two_stage_opamp_dummy_magic_16_0.cap_res_X.t10 GNDA 0.184828f
C1744 two_stage_opamp_dummy_magic_16_0.cap_res_X.n23 GNDA 0.251826f
C1745 two_stage_opamp_dummy_magic_16_0.cap_res_X.t45 GNDA 0.184828f
C1746 two_stage_opamp_dummy_magic_16_0.cap_res_X.n24 GNDA 0.251826f
C1747 two_stage_opamp_dummy_magic_16_0.cap_res_X.t2 GNDA 0.184828f
C1748 two_stage_opamp_dummy_magic_16_0.cap_res_X.n25 GNDA 0.234498f
C1749 two_stage_opamp_dummy_magic_16_0.cap_res_X.t1 GNDA 0.3451f
C1750 two_stage_opamp_dummy_magic_16_0.cap_res_X.t41 GNDA 0.167396f
C1751 two_stage_opamp_dummy_magic_16_0.cap_res_X.n26 GNDA 0.217171f
C1752 two_stage_opamp_dummy_magic_16_0.cap_res_X.t122 GNDA 0.3451f
C1753 two_stage_opamp_dummy_magic_16_0.cap_res_X.t25 GNDA 0.346251f
C1754 two_stage_opamp_dummy_magic_16_0.cap_res_X.t58 GNDA 0.364834f
C1755 two_stage_opamp_dummy_magic_16_0.cap_res_X.t21 GNDA 0.185978f
C1756 two_stage_opamp_dummy_magic_16_0.cap_res_X.n27 GNDA 0.217171f
C1757 two_stage_opamp_dummy_magic_16_0.cap_res_X.t126 GNDA 0.3451f
C1758 two_stage_opamp_dummy_magic_16_0.cap_res_X.t66 GNDA 0.346251f
C1759 two_stage_opamp_dummy_magic_16_0.cap_res_X.t27 GNDA 0.185978f
C1760 two_stage_opamp_dummy_magic_16_0.cap_res_X.n28 GNDA 0.198589f
C1761 two_stage_opamp_dummy_magic_16_0.cap_res_X.t8 GNDA 0.3451f
C1762 two_stage_opamp_dummy_magic_16_0.cap_res_X.t88 GNDA 0.346251f
C1763 two_stage_opamp_dummy_magic_16_0.cap_res_X.t49 GNDA 0.185978f
C1764 two_stage_opamp_dummy_magic_16_0.cap_res_X.n29 GNDA 0.217171f
C1765 two_stage_opamp_dummy_magic_16_0.cap_res_X.t107 GNDA 0.3451f
C1766 two_stage_opamp_dummy_magic_16_0.cap_res_X.t50 GNDA 0.346251f
C1767 two_stage_opamp_dummy_magic_16_0.cap_res_X.t11 GNDA 0.185978f
C1768 two_stage_opamp_dummy_magic_16_0.cap_res_X.n30 GNDA 0.217171f
C1769 two_stage_opamp_dummy_magic_16_0.cap_res_X.t74 GNDA 0.3451f
C1770 two_stage_opamp_dummy_magic_16_0.cap_res_X.t13 GNDA 0.346251f
C1771 two_stage_opamp_dummy_magic_16_0.cap_res_X.t112 GNDA 0.185978f
C1772 two_stage_opamp_dummy_magic_16_0.cap_res_X.n31 GNDA 0.217171f
C1773 two_stage_opamp_dummy_magic_16_0.cap_res_X.t37 GNDA 0.3451f
C1774 two_stage_opamp_dummy_magic_16_0.cap_res_X.t91 GNDA 0.346251f
C1775 two_stage_opamp_dummy_magic_16_0.cap_res_X.t80 GNDA 0.364834f
C1776 two_stage_opamp_dummy_magic_16_0.cap_res_X.t114 GNDA 0.364834f
C1777 two_stage_opamp_dummy_magic_16_0.cap_res_X.t76 GNDA 0.185978f
C1778 two_stage_opamp_dummy_magic_16_0.cap_res_X.n32 GNDA 0.217171f
C1779 two_stage_opamp_dummy_magic_16_0.cap_res_X.t53 GNDA 0.3451f
C1780 two_stage_opamp_dummy_magic_16_0.cap_res_X.t42 GNDA 0.346251f
C1781 two_stage_opamp_dummy_magic_16_0.cap_res_X.t99 GNDA 0.364834f
C1782 two_stage_opamp_dummy_magic_16_0.cap_res_X.t135 GNDA 0.364834f
C1783 two_stage_opamp_dummy_magic_16_0.cap_res_X.t93 GNDA 0.185978f
C1784 two_stage_opamp_dummy_magic_16_0.cap_res_X.n33 GNDA 0.217171f
C1785 two_stage_opamp_dummy_magic_16_0.cap_res_X.t20 GNDA 0.3451f
C1786 two_stage_opamp_dummy_magic_16_0.cap_res_X.n34 GNDA 0.217171f
C1787 two_stage_opamp_dummy_magic_16_0.cap_res_X.t57 GNDA 0.185978f
C1788 two_stage_opamp_dummy_magic_16_0.cap_res_X.t96 GNDA 0.364834f
C1789 two_stage_opamp_dummy_magic_16_0.cap_res_X.t63 GNDA 0.364834f
C1790 two_stage_opamp_dummy_magic_16_0.cap_res_X.t7 GNDA 0.430822f
C1791 two_stage_opamp_dummy_magic_16_0.cap_res_X.t0 GNDA 0.292647f
C1792 VOUT-.t14 GNDA 0.041786f
C1793 VOUT-.t6 GNDA 0.041786f
C1794 VOUT-.n0 GNDA 0.16895f
C1795 VOUT-.t2 GNDA 0.041786f
C1796 VOUT-.t15 GNDA 0.041786f
C1797 VOUT-.n1 GNDA 0.168949f
C1798 VOUT-.t8 GNDA 0.041786f
C1799 VOUT-.t0 GNDA 0.041786f
C1800 VOUT-.n2 GNDA 0.168648f
C1801 VOUT-.n3 GNDA 0.164536f
C1802 VOUT-.t7 GNDA 0.041786f
C1803 VOUT-.t1 GNDA 0.041786f
C1804 VOUT-.n4 GNDA 0.168648f
C1805 VOUT-.n5 GNDA 0.084856f
C1806 VOUT-.t4 GNDA 0.041786f
C1807 VOUT-.t3 GNDA 0.041786f
C1808 VOUT-.n6 GNDA 0.168648f
C1809 VOUT-.n7 GNDA 0.084856f
C1810 VOUT-.n8 GNDA 0.100572f
C1811 VOUT-.t9 GNDA 0.041786f
C1812 VOUT-.t5 GNDA 0.041786f
C1813 VOUT-.n9 GNDA 0.166651f
C1814 VOUT-.n10 GNDA 0.141149f
C1815 VOUT-.t26 GNDA 0.283321f
C1816 VOUT-.t119 GNDA 0.278576f
C1817 VOUT-.n11 GNDA 0.186776f
C1818 VOUT-.t33 GNDA 0.278576f
C1819 VOUT-.n12 GNDA 0.121877f
C1820 VOUT-.t36 GNDA 0.283321f
C1821 VOUT-.t122 GNDA 0.278576f
C1822 VOUT-.n13 GNDA 0.186776f
C1823 VOUT-.t90 GNDA 0.278576f
C1824 VOUT-.t82 GNDA 0.282727f
C1825 VOUT-.t42 GNDA 0.282727f
C1826 VOUT-.t92 GNDA 0.282727f
C1827 VOUT-.t74 GNDA 0.282727f
C1828 VOUT-.t141 GNDA 0.282727f
C1829 VOUT-.t38 GNDA 0.282727f
C1830 VOUT-.t105 GNDA 0.282727f
C1831 VOUT-.t126 GNDA 0.282727f
C1832 VOUT-.t154 GNDA 0.282727f
C1833 VOUT-.t95 GNDA 0.282727f
C1834 VOUT-.t65 GNDA 0.282727f
C1835 VOUT-.t62 GNDA 0.282727f
C1836 VOUT-.t114 GNDA 0.282727f
C1837 VOUT-.t24 GNDA 0.282727f
C1838 VOUT-.t71 GNDA 0.282727f
C1839 VOUT-.t113 GNDA 0.282727f
C1840 VOUT-.t148 GNDA 0.278576f
C1841 VOUT-.n14 GNDA 0.305096f
C1842 VOUT-.t60 GNDA 0.278576f
C1843 VOUT-.n15 GNDA 0.357329f
C1844 VOUT-.t93 GNDA 0.278576f
C1845 VOUT-.n16 GNDA 0.357329f
C1846 VOUT-.t127 GNDA 0.278576f
C1847 VOUT-.n17 GNDA 0.357329f
C1848 VOUT-.t25 GNDA 0.278576f
C1849 VOUT-.n18 GNDA 0.357329f
C1850 VOUT-.t72 GNDA 0.278576f
C1851 VOUT-.n19 GNDA 0.357329f
C1852 VOUT-.t110 GNDA 0.278576f
C1853 VOUT-.n20 GNDA 0.357329f
C1854 VOUT-.t142 GNDA 0.278576f
C1855 VOUT-.n21 GNDA 0.239603f
C1856 VOUT-.t56 GNDA 0.278576f
C1857 VOUT-.n22 GNDA 0.239603f
C1858 VOUT-.n23 GNDA 0.226343f
C1859 VOUT-.t140 GNDA 0.283321f
C1860 VOUT-.t89 GNDA 0.278576f
C1861 VOUT-.n24 GNDA 0.186776f
C1862 VOUT-.t59 GNDA 0.278576f
C1863 VOUT-.t111 GNDA 0.283321f
C1864 VOUT-.t21 GNDA 0.278576f
C1865 VOUT-.n25 GNDA 0.186776f
C1866 VOUT-.n26 GNDA 0.226343f
C1867 VOUT-.t41 GNDA 0.283321f
C1868 VOUT-.t129 GNDA 0.278576f
C1869 VOUT-.n27 GNDA 0.186776f
C1870 VOUT-.t98 GNDA 0.278576f
C1871 VOUT-.t151 GNDA 0.283321f
C1872 VOUT-.t63 GNDA 0.278576f
C1873 VOUT-.n28 GNDA 0.186776f
C1874 VOUT-.n29 GNDA 0.226343f
C1875 VOUT-.t80 GNDA 0.283321f
C1876 VOUT-.t30 GNDA 0.278576f
C1877 VOUT-.n30 GNDA 0.186776f
C1878 VOUT-.t134 GNDA 0.278576f
C1879 VOUT-.t51 GNDA 0.283321f
C1880 VOUT-.t103 GNDA 0.278576f
C1881 VOUT-.n31 GNDA 0.186776f
C1882 VOUT-.n32 GNDA 0.226343f
C1883 VOUT-.t49 GNDA 0.283321f
C1884 VOUT-.t135 GNDA 0.278576f
C1885 VOUT-.n33 GNDA 0.186776f
C1886 VOUT-.t102 GNDA 0.278576f
C1887 VOUT-.t19 GNDA 0.283321f
C1888 VOUT-.t67 GNDA 0.278576f
C1889 VOUT-.n34 GNDA 0.186776f
C1890 VOUT-.n35 GNDA 0.226343f
C1891 VOUT-.t85 GNDA 0.283321f
C1892 VOUT-.t34 GNDA 0.278576f
C1893 VOUT-.n36 GNDA 0.186776f
C1894 VOUT-.t139 GNDA 0.278576f
C1895 VOUT-.t55 GNDA 0.283321f
C1896 VOUT-.t106 GNDA 0.278576f
C1897 VOUT-.n37 GNDA 0.186776f
C1898 VOUT-.n38 GNDA 0.226343f
C1899 VOUT-.t68 GNDA 0.283321f
C1900 VOUT-.t86 GNDA 0.278576f
C1901 VOUT-.n39 GNDA 0.186776f
C1902 VOUT-.t54 GNDA 0.278576f
C1903 VOUT-.n40 GNDA 0.121877f
C1904 VOUT-.t29 GNDA 0.283321f
C1905 VOUT-.t52 GNDA 0.278576f
C1906 VOUT-.n41 GNDA 0.186776f
C1907 VOUT-.t155 GNDA 0.278576f
C1908 VOUT-.t156 GNDA 0.282727f
C1909 VOUT-.t132 GNDA 0.283321f
C1910 VOUT-.t99 GNDA 0.278576f
C1911 VOUT-.n42 GNDA 0.182423f
C1912 VOUT-.t35 GNDA 0.282727f
C1913 VOUT-.t150 GNDA 0.283321f
C1914 VOUT-.t94 GNDA 0.278576f
C1915 VOUT-.n43 GNDA 0.186776f
C1916 VOUT-.t61 GNDA 0.278576f
C1917 VOUT-.n44 GNDA 0.117524f
C1918 VOUT-.t137 GNDA 0.282727f
C1919 VOUT-.t115 GNDA 0.283321f
C1920 VOUT-.t58 GNDA 0.278576f
C1921 VOUT-.n45 GNDA 0.186776f
C1922 VOUT-.t22 GNDA 0.278576f
C1923 VOUT-.n46 GNDA 0.117524f
C1924 VOUT-.t104 GNDA 0.282727f
C1925 VOUT-.t66 GNDA 0.283321f
C1926 VOUT-.t77 GNDA 0.278576f
C1927 VOUT-.n47 GNDA 0.186776f
C1928 VOUT-.t43 GNDA 0.278576f
C1929 VOUT-.n48 GNDA 0.117524f
C1930 VOUT-.t120 GNDA 0.282727f
C1931 VOUT-.t144 GNDA 0.282727f
C1932 VOUT-.t83 GNDA 0.282727f
C1933 VOUT-.t107 GNDA 0.28296f
C1934 VOUT-.t50 GNDA 0.282727f
C1935 VOUT-.t69 GNDA 0.28296f
C1936 VOUT-.t149 GNDA 0.282727f
C1937 VOUT-.t91 GNDA 0.28296f
C1938 VOUT-.t31 GNDA 0.282727f
C1939 VOUT-.t130 GNDA 0.278576f
C1940 VOUT-.n49 GNDA 0.308345f
C1941 VOUT-.t108 GNDA 0.278576f
C1942 VOUT-.n50 GNDA 0.360578f
C1943 VOUT-.t146 GNDA 0.278576f
C1944 VOUT-.n51 GNDA 0.360578f
C1945 VOUT-.t45 GNDA 0.278576f
C1946 VOUT-.n52 GNDA 0.357329f
C1947 VOUT-.t81 GNDA 0.278576f
C1948 VOUT-.n53 GNDA 0.296189f
C1949 VOUT-.t64 GNDA 0.278576f
C1950 VOUT-.n54 GNDA 0.296189f
C1951 VOUT-.t100 GNDA 0.278576f
C1952 VOUT-.n55 GNDA 0.296189f
C1953 VOUT-.t136 GNDA 0.278576f
C1954 VOUT-.n56 GNDA 0.296189f
C1955 VOUT-.t116 GNDA 0.278576f
C1956 VOUT-.n57 GNDA 0.239603f
C1957 VOUT-.n58 GNDA 0.226343f
C1958 VOUT-.t125 GNDA 0.283321f
C1959 VOUT-.t152 GNDA 0.278576f
C1960 VOUT-.n59 GNDA 0.186776f
C1961 VOUT-.t112 GNDA 0.278576f
C1962 VOUT-.t73 GNDA 0.283321f
C1963 VOUT-.n60 GNDA 0.291242f
C1964 VOUT-.t23 GNDA 0.283321f
C1965 VOUT-.t47 GNDA 0.278576f
C1966 VOUT-.n61 GNDA 0.186776f
C1967 VOUT-.t147 GNDA 0.278576f
C1968 VOUT-.t109 GNDA 0.283321f
C1969 VOUT-.n62 GNDA 0.291242f
C1970 VOUT-.t76 GNDA 0.283321f
C1971 VOUT-.t27 GNDA 0.278576f
C1972 VOUT-.n63 GNDA 0.186776f
C1973 VOUT-.t128 GNDA 0.278576f
C1974 VOUT-.t44 GNDA 0.283321f
C1975 VOUT-.t97 GNDA 0.278576f
C1976 VOUT-.n64 GNDA 0.186776f
C1977 VOUT-.n65 GNDA 0.226343f
C1978 VOUT-.t37 GNDA 0.283321f
C1979 VOUT-.t123 GNDA 0.278576f
C1980 VOUT-.n66 GNDA 0.186776f
C1981 VOUT-.t88 GNDA 0.278576f
C1982 VOUT-.t143 GNDA 0.283321f
C1983 VOUT-.t57 GNDA 0.278576f
C1984 VOUT-.n67 GNDA 0.186776f
C1985 VOUT-.n68 GNDA 0.226343f
C1986 VOUT-.t70 GNDA 0.283321f
C1987 VOUT-.t20 GNDA 0.278576f
C1988 VOUT-.n69 GNDA 0.186776f
C1989 VOUT-.t121 GNDA 0.278576f
C1990 VOUT-.t39 GNDA 0.283321f
C1991 VOUT-.t87 GNDA 0.278576f
C1992 VOUT-.n70 GNDA 0.186776f
C1993 VOUT-.n71 GNDA 0.226343f
C1994 VOUT-.t32 GNDA 0.283321f
C1995 VOUT-.t118 GNDA 0.278576f
C1996 VOUT-.n72 GNDA 0.186776f
C1997 VOUT-.t84 GNDA 0.278576f
C1998 VOUT-.t138 GNDA 0.283321f
C1999 VOUT-.t53 GNDA 0.278576f
C2000 VOUT-.n73 GNDA 0.186776f
C2001 VOUT-.n74 GNDA 0.226343f
C2002 VOUT-.t131 GNDA 0.283321f
C2003 VOUT-.t79 GNDA 0.278576f
C2004 VOUT-.n75 GNDA 0.186776f
C2005 VOUT-.t48 GNDA 0.278576f
C2006 VOUT-.t101 GNDA 0.283321f
C2007 VOUT-.t153 GNDA 0.278576f
C2008 VOUT-.n76 GNDA 0.186776f
C2009 VOUT-.n77 GNDA 0.226343f
C2010 VOUT-.t28 GNDA 0.283321f
C2011 VOUT-.t117 GNDA 0.278576f
C2012 VOUT-.n78 GNDA 0.186776f
C2013 VOUT-.t78 GNDA 0.278576f
C2014 VOUT-.t133 GNDA 0.283321f
C2015 VOUT-.t46 GNDA 0.278576f
C2016 VOUT-.n79 GNDA 0.186776f
C2017 VOUT-.n80 GNDA 0.226343f
C2018 VOUT-.t124 GNDA 0.283321f
C2019 VOUT-.t75 GNDA 0.278576f
C2020 VOUT-.n81 GNDA 0.186776f
C2021 VOUT-.t40 GNDA 0.278576f
C2022 VOUT-.n82 GNDA 0.226343f
C2023 VOUT-.t145 GNDA 0.278576f
C2024 VOUT-.n83 GNDA 0.121877f
C2025 VOUT-.t96 GNDA 0.278576f
C2026 VOUT-.n84 GNDA 0.177725f
C2027 VOUT-.n85 GNDA 0.212227f
C2028 VOUT-.t17 GNDA 0.048751f
C2029 VOUT-.t12 GNDA 0.048751f
C2030 VOUT-.n86 GNDA 0.226297f
C2031 VOUT-.t18 GNDA 0.048751f
C2032 VOUT-.t10 GNDA 0.048751f
C2033 VOUT-.n87 GNDA 0.225568f
C2034 VOUT-.n88 GNDA 0.138716f
C2035 VOUT-.t13 GNDA 0.048751f
C2036 VOUT-.t11 GNDA 0.048751f
C2037 VOUT-.n89 GNDA 0.225568f
C2038 VOUT-.n90 GNDA 0.077273f
C2039 VOUT-.t16 GNDA 0.081149f
C2040 VOUT-.n91 GNDA 0.089317f
C2041 bgr_0.V_TOP.t24 GNDA 0.095448f
C2042 bgr_0.V_TOP.t33 GNDA 0.095448f
C2043 bgr_0.V_TOP.t39 GNDA 0.095448f
C2044 bgr_0.V_TOP.t16 GNDA 0.095448f
C2045 bgr_0.V_TOP.t15 GNDA 0.095448f
C2046 bgr_0.V_TOP.t28 GNDA 0.095448f
C2047 bgr_0.V_TOP.t38 GNDA 0.095448f
C2048 bgr_0.V_TOP.t14 GNDA 0.095448f
C2049 bgr_0.V_TOP.t27 GNDA 0.095448f
C2050 bgr_0.V_TOP.t26 GNDA 0.095448f
C2051 bgr_0.V_TOP.t37 GNDA 0.095448f
C2052 bgr_0.V_TOP.t46 GNDA 0.095448f
C2053 bgr_0.V_TOP.t18 GNDA 0.095448f
C2054 bgr_0.V_TOP.t30 GNDA 0.095448f
C2055 bgr_0.V_TOP.t29 GNDA 0.124774f
C2056 bgr_0.V_TOP.n0 GNDA 0.069758f
C2057 bgr_0.V_TOP.n1 GNDA 0.050905f
C2058 bgr_0.V_TOP.n2 GNDA 0.050905f
C2059 bgr_0.V_TOP.n3 GNDA 0.050905f
C2060 bgr_0.V_TOP.n4 GNDA 0.050905f
C2061 bgr_0.V_TOP.n5 GNDA 0.04747f
C2062 bgr_0.V_TOP.t7 GNDA 0.122745f
C2063 bgr_0.V_TOP.t40 GNDA 0.36361f
C2064 bgr_0.V_TOP.t31 GNDA 0.369803f
C2065 bgr_0.V_TOP.t35 GNDA 0.36361f
C2066 bgr_0.V_TOP.n6 GNDA 0.243789f
C2067 bgr_0.V_TOP.t32 GNDA 0.36361f
C2068 bgr_0.V_TOP.t22 GNDA 0.369803f
C2069 bgr_0.V_TOP.n7 GNDA 0.311966f
C2070 bgr_0.V_TOP.t20 GNDA 0.369803f
C2071 bgr_0.V_TOP.t25 GNDA 0.36361f
C2072 bgr_0.V_TOP.n8 GNDA 0.243789f
C2073 bgr_0.V_TOP.t21 GNDA 0.36361f
C2074 bgr_0.V_TOP.t45 GNDA 0.369803f
C2075 bgr_0.V_TOP.n9 GNDA 0.380142f
C2076 bgr_0.V_TOP.t42 GNDA 0.369803f
C2077 bgr_0.V_TOP.t49 GNDA 0.36361f
C2078 bgr_0.V_TOP.n10 GNDA 0.243789f
C2079 bgr_0.V_TOP.t44 GNDA 0.36361f
C2080 bgr_0.V_TOP.t36 GNDA 0.369803f
C2081 bgr_0.V_TOP.n11 GNDA 0.380142f
C2082 bgr_0.V_TOP.t17 GNDA 0.369803f
C2083 bgr_0.V_TOP.t23 GNDA 0.36361f
C2084 bgr_0.V_TOP.n12 GNDA 0.243789f
C2085 bgr_0.V_TOP.t19 GNDA 0.36361f
C2086 bgr_0.V_TOP.t43 GNDA 0.369803f
C2087 bgr_0.V_TOP.n13 GNDA 0.380142f
C2088 bgr_0.V_TOP.t34 GNDA 0.369803f
C2089 bgr_0.V_TOP.t41 GNDA 0.36361f
C2090 bgr_0.V_TOP.n14 GNDA 0.311966f
C2091 bgr_0.V_TOP.t47 GNDA 0.36361f
C2092 bgr_0.V_TOP.n15 GNDA 0.159079f
C2093 bgr_0.V_TOP.n16 GNDA 0.544408f
C2094 bgr_0.V_TOP.t3 GNDA 0.102288f
C2095 bgr_0.V_TOP.n17 GNDA 0.724299f
C2096 bgr_0.V_TOP.n18 GNDA 0.022634f
C2097 bgr_0.V_TOP.n19 GNDA 0.414649f
C2098 bgr_0.V_TOP.n20 GNDA 0.021924f
C2099 bgr_0.V_TOP.n21 GNDA 0.022786f
C2100 bgr_0.V_TOP.n22 GNDA 0.022634f
C2101 bgr_0.V_TOP.n23 GNDA 0.209756f
C2102 bgr_0.V_TOP.n24 GNDA 0.127416f
C2103 bgr_0.V_TOP.n25 GNDA 0.072722f
C2104 bgr_0.V_TOP.n26 GNDA 0.022634f
C2105 bgr_0.V_TOP.n27 GNDA 0.125537f
C2106 bgr_0.V_TOP.n28 GNDA 0.022634f
C2107 bgr_0.V_TOP.n29 GNDA 0.124344f
C2108 bgr_0.V_TOP.n30 GNDA 0.273328f
C2109 bgr_0.V_TOP.n31 GNDA 0.019234f
C2110 bgr_0.V_TOP.n32 GNDA 0.04747f
C2111 bgr_0.V_TOP.n33 GNDA 0.050905f
C2112 bgr_0.V_TOP.n34 GNDA 0.050905f
C2113 bgr_0.V_TOP.n35 GNDA 0.050905f
C2114 bgr_0.V_TOP.n36 GNDA 0.050905f
C2115 bgr_0.V_TOP.n37 GNDA 0.050905f
C2116 bgr_0.V_TOP.n38 GNDA 0.050905f
C2117 bgr_0.V_TOP.n39 GNDA 0.04747f
C2118 bgr_0.V_TOP.t48 GNDA 0.109989f
C2119 VDDA.t255 GNDA 0.021275f
C2120 VDDA.t261 GNDA 0.021275f
C2121 VDDA.n0 GNDA 0.073729f
C2122 VDDA.n1 GNDA 0.072159f
C2123 VDDA.t279 GNDA 0.021275f
C2124 VDDA.n2 GNDA 0.063826f
C2125 VDDA.n3 GNDA 0.021275f
C2126 VDDA.n4 GNDA 0.012157f
C2127 VDDA.n8 GNDA 0.012157f
C2128 VDDA.t323 GNDA 0.037303f
C2129 VDDA.t247 GNDA 0.021275f
C2130 VDDA.t243 GNDA 0.021275f
C2131 VDDA.n9 GNDA 0.073729f
C2132 VDDA.n10 GNDA 0.092386f
C2133 VDDA.n11 GNDA 0.031681f
C2134 VDDA.n12 GNDA 0.021275f
C2135 VDDA.n14 GNDA 0.021275f
C2136 VDDA.n15 GNDA 0.012157f
C2137 VDDA.n16 GNDA 0.012157f
C2138 VDDA.n17 GNDA 0.021275f
C2139 VDDA.n19 GNDA 0.021275f
C2140 VDDA.n20 GNDA 0.012157f
C2141 VDDA.n21 GNDA 0.012157f
C2142 VDDA.n22 GNDA 0.021275f
C2143 VDDA.n23 GNDA 0.021461f
C2144 VDDA.t325 GNDA 0.021275f
C2145 VDDA.n24 GNDA 0.063826f
C2146 VDDA.n25 GNDA 0.020509f
C2147 VDDA.n26 GNDA 0.012157f
C2148 VDDA.n27 GNDA 0.177801f
C2149 VDDA.t324 GNDA 0.154094f
C2150 VDDA.t246 GNDA 0.142241f
C2151 VDDA.t242 GNDA 0.142241f
C2152 VDDA.t254 GNDA 0.142241f
C2153 VDDA.t260 GNDA 0.142241f
C2154 VDDA.t222 GNDA 0.142241f
C2155 VDDA.t224 GNDA 0.142241f
C2156 VDDA.t236 GNDA 0.142241f
C2157 VDDA.t244 GNDA 0.142241f
C2158 VDDA.t256 GNDA 0.142241f
C2159 VDDA.t262 GNDA 0.142241f
C2160 VDDA.t278 GNDA 0.154094f
C2161 VDDA.n30 GNDA 0.012157f
C2162 VDDA.n32 GNDA 0.021461f
C2163 VDDA.n33 GNDA 0.021275f
C2164 VDDA.n34 GNDA 0.012157f
C2165 VDDA.n35 GNDA 0.012157f
C2166 VDDA.n36 GNDA 0.021275f
C2167 VDDA.n38 GNDA 0.021275f
C2168 VDDA.n39 GNDA 0.021275f
C2169 VDDA.n40 GNDA 0.012157f
C2170 VDDA.n41 GNDA 0.177801f
C2171 VDDA.n43 GNDA 0.023231f
C2172 VDDA.t277 GNDA 0.037303f
C2173 VDDA.n44 GNDA 0.031681f
C2174 VDDA.t257 GNDA 0.021275f
C2175 VDDA.t263 GNDA 0.021275f
C2176 VDDA.n45 GNDA 0.073729f
C2177 VDDA.n46 GNDA 0.092386f
C2178 VDDA.t237 GNDA 0.021275f
C2179 VDDA.t245 GNDA 0.021275f
C2180 VDDA.n47 GNDA 0.073729f
C2181 VDDA.n48 GNDA 0.072159f
C2182 VDDA.n49 GNDA 0.019452f
C2183 VDDA.t223 GNDA 0.021275f
C2184 VDDA.t225 GNDA 0.021275f
C2185 VDDA.n50 GNDA 0.072202f
C2186 VDDA.n51 GNDA 0.083176f
C2187 VDDA.t266 GNDA 0.018236f
C2188 VDDA.t73 GNDA 0.018236f
C2189 VDDA.n52 GNDA 0.075413f
C2190 VDDA.t150 GNDA 0.018236f
C2191 VDDA.t13 GNDA 0.018236f
C2192 VDDA.n53 GNDA 0.075124f
C2193 VDDA.n54 GNDA 0.104159f
C2194 VDDA.t146 GNDA 0.018236f
C2195 VDDA.t89 GNDA 0.018236f
C2196 VDDA.n55 GNDA 0.075124f
C2197 VDDA.n56 GNDA 0.054352f
C2198 VDDA.t159 GNDA 0.018236f
C2199 VDDA.t158 GNDA 0.018236f
C2200 VDDA.n57 GNDA 0.075124f
C2201 VDDA.n58 GNDA 0.054352f
C2202 VDDA.t155 GNDA 0.018236f
C2203 VDDA.t157 GNDA 0.018236f
C2204 VDDA.n59 GNDA 0.075124f
C2205 VDDA.n60 GNDA 0.054352f
C2206 VDDA.t133 GNDA 0.018236f
C2207 VDDA.t267 GNDA 0.018236f
C2208 VDDA.n61 GNDA 0.075124f
C2209 VDDA.n62 GNDA 0.110331f
C2210 VDDA.t371 GNDA 0.018376f
C2211 VDDA.n64 GNDA 0.012157f
C2212 VDDA.n66 GNDA 0.012157f
C2213 VDDA.t353 GNDA 0.019205f
C2214 VDDA.n67 GNDA 0.021275f
C2215 VDDA.n68 GNDA 0.012157f
C2216 VDDA.n69 GNDA 0.021275f
C2217 VDDA.n70 GNDA 0.029601f
C2218 VDDA.t355 GNDA 0.032052f
C2219 VDDA.n72 GNDA 0.048665f
C2220 VDDA.n74 GNDA 0.107592f
C2221 VDDA.t354 GNDA 0.089356f
C2222 VDDA.t91 GNDA 0.080238f
C2223 VDDA.t75 GNDA 0.080238f
C2224 VDDA.t156 GNDA 0.080238f
C2225 VDDA.t74 GNDA 0.080238f
C2226 VDDA.t70 GNDA 0.080238f
C2227 VDDA.t14 GNDA 0.080238f
C2228 VDDA.t209 GNDA 0.080238f
C2229 VDDA.t130 GNDA 0.080238f
C2230 VDDA.t147 GNDA 0.080238f
C2231 VDDA.t90 GNDA 0.080238f
C2232 VDDA.t372 GNDA 0.089356f
C2233 VDDA.n76 GNDA 0.012157f
C2234 VDDA.n77 GNDA 0.021275f
C2235 VDDA.n78 GNDA 0.021275f
C2236 VDDA.t373 GNDA 0.032052f
C2237 VDDA.n79 GNDA 0.026799f
C2238 VDDA.n80 GNDA 0.012795f
C2239 VDDA.n81 GNDA 0.107592f
C2240 VDDA.n82 GNDA 0.012157f
C2241 VDDA.n83 GNDA 0.024111f
C2242 VDDA.n84 GNDA 0.038962f
C2243 VDDA.n85 GNDA 0.171778f
C2244 VDDA.t50 GNDA 0.036472f
C2245 VDDA.t72 GNDA 0.036472f
C2246 VDDA.n86 GNDA 0.146321f
C2247 VDDA.n87 GNDA 0.074335f
C2248 VDDA.n89 GNDA 0.012157f
C2249 VDDA.n95 GNDA 0.012795f
C2250 VDDA.n96 GNDA 0.012157f
C2251 VDDA.t311 GNDA 0.044192f
C2252 VDDA.t52 GNDA 0.036472f
C2253 VDDA.t152 GNDA 0.036472f
C2254 VDDA.n97 GNDA 0.146321f
C2255 VDDA.n98 GNDA 0.074335f
C2256 VDDA.t77 GNDA 0.036472f
C2257 VDDA.t149 GNDA 0.036472f
C2258 VDDA.n99 GNDA 0.146321f
C2259 VDDA.n100 GNDA 0.074335f
C2260 VDDA.t132 GNDA 0.036472f
C2261 VDDA.t93 GNDA 0.036472f
C2262 VDDA.n101 GNDA 0.146321f
C2263 VDDA.n102 GNDA 0.074335f
C2264 VDDA.t135 GNDA 0.036472f
C2265 VDDA.t154 GNDA 0.036472f
C2266 VDDA.n103 GNDA 0.146321f
C2267 VDDA.n104 GNDA 0.094066f
C2268 VDDA.n105 GNDA 0.036381f
C2269 VDDA.n106 GNDA 0.024187f
C2270 VDDA.n107 GNDA 0.012157f
C2271 VDDA.n108 GNDA 0.012157f
C2272 VDDA.n109 GNDA 0.021275f
C2273 VDDA.n110 GNDA 0.012157f
C2274 VDDA.n111 GNDA 0.012157f
C2275 VDDA.n112 GNDA 0.012157f
C2276 VDDA.n113 GNDA 0.012157f
C2277 VDDA.n114 GNDA 0.021275f
C2278 VDDA.n115 GNDA 0.024187f
C2279 VDDA.n116 GNDA 0.012157f
C2280 VDDA.n117 GNDA 0.012157f
C2281 VDDA.n118 GNDA 0.012157f
C2282 VDDA.n119 GNDA 0.030795f
C2283 VDDA.n120 GNDA 0.021275f
C2284 VDDA.n121 GNDA 0.021275f
C2285 VDDA.n122 GNDA 0.021275f
C2286 VDDA.n123 GNDA 0.012157f
C2287 VDDA.n124 GNDA 0.012157f
C2288 VDDA.n126 GNDA 0.021275f
C2289 VDDA.n127 GNDA 0.021275f
C2290 VDDA.n129 GNDA 0.012157f
C2291 VDDA.n130 GNDA 0.012157f
C2292 VDDA.n131 GNDA 0.021275f
C2293 VDDA.n132 GNDA 0.021275f
C2294 VDDA.n133 GNDA 0.021275f
C2295 VDDA.n135 GNDA 0.024111f
C2296 VDDA.n136 GNDA 0.012157f
C2297 VDDA.n137 GNDA 0.286913f
C2298 VDDA.t312 GNDA 0.238283f
C2299 VDDA.t134 GNDA 0.213969f
C2300 VDDA.t153 GNDA 0.213969f
C2301 VDDA.t131 GNDA 0.213969f
C2302 VDDA.t92 GNDA 0.213969f
C2303 VDDA.t76 GNDA 0.213969f
C2304 VDDA.t148 GNDA 0.213969f
C2305 VDDA.t51 GNDA 0.213969f
C2306 VDDA.t151 GNDA 0.213969f
C2307 VDDA.t49 GNDA 0.213969f
C2308 VDDA.t71 GNDA 0.213969f
C2309 VDDA.t327 GNDA 0.238283f
C2310 VDDA.n142 GNDA 0.012795f
C2311 VDDA.n143 GNDA 0.012157f
C2312 VDDA.n144 GNDA 0.021275f
C2313 VDDA.n145 GNDA 0.024187f
C2314 VDDA.n146 GNDA 0.012157f
C2315 VDDA.n147 GNDA 0.012157f
C2316 VDDA.n150 GNDA 0.012157f
C2317 VDDA.n151 GNDA 0.012157f
C2318 VDDA.n152 GNDA 0.024187f
C2319 VDDA.n153 GNDA 0.030795f
C2320 VDDA.n154 GNDA 0.012157f
C2321 VDDA.n155 GNDA 0.021275f
C2322 VDDA.n156 GNDA 0.021275f
C2323 VDDA.n157 GNDA 0.012157f
C2324 VDDA.n158 GNDA 0.012157f
C2325 VDDA.n159 GNDA 0.021275f
C2326 VDDA.n160 GNDA 0.021275f
C2327 VDDA.n161 GNDA 0.012157f
C2328 VDDA.n162 GNDA 0.012157f
C2329 VDDA.n163 GNDA 0.021275f
C2330 VDDA.n164 GNDA 0.021275f
C2331 VDDA.n165 GNDA 0.012157f
C2332 VDDA.n166 GNDA 0.012157f
C2333 VDDA.n167 GNDA 0.021275f
C2334 VDDA.n168 GNDA 0.021275f
C2335 VDDA.n169 GNDA 0.021275f
C2336 VDDA.n170 GNDA 0.012157f
C2337 VDDA.n171 GNDA 0.286913f
C2338 VDDA.n173 GNDA 0.026833f
C2339 VDDA.t326 GNDA 0.044192f
C2340 VDDA.n174 GNDA 0.035577f
C2341 VDDA.n175 GNDA 0.049454f
C2342 VDDA.n176 GNDA 0.064692f
C2343 VDDA.t39 GNDA 0.015197f
C2344 VDDA.t383 GNDA 0.015197f
C2345 VDDA.n177 GNDA 0.0524f
C2346 VDDA.n178 GNDA 0.067761f
C2347 VDDA.t343 GNDA 0.015197f
C2348 VDDA.n179 GNDA 0.04559f
C2349 VDDA.n180 GNDA 0.021275f
C2350 VDDA.n181 GNDA 0.012157f
C2351 VDDA.t287 GNDA 0.107972f
C2352 VDDA.n184 GNDA 0.012157f
C2353 VDDA.n185 GNDA 0.012157f
C2354 VDDA.t368 GNDA 0.022836f
C2355 VDDA.n186 GNDA 0.031153f
C2356 VDDA.n187 GNDA 0.026408f
C2357 VDDA.t289 GNDA 0.022836f
C2358 VDDA.t291 GNDA 0.015197f
C2359 VDDA.n188 GNDA 0.04559f
C2360 VDDA.n189 GNDA 0.021275f
C2361 VDDA.n190 GNDA 0.012157f
C2362 VDDA.t386 GNDA 0.096955f
C2363 VDDA.t379 GNDA 0.096955f
C2364 VDDA.t387 GNDA 0.096955f
C2365 VDDA.t109 GNDA 0.096955f
C2366 VDDA.t290 GNDA 0.107972f
C2367 VDDA.n192 GNDA 0.012157f
C2368 VDDA.n194 GNDA 0.012157f
C2369 VDDA.n195 GNDA 0.021275f
C2370 VDDA.n196 GNDA 0.021275f
C2371 VDDA.n197 GNDA 0.021461f
C2372 VDDA.n199 GNDA 0.130007f
C2373 VDDA.n200 GNDA 0.012157f
C2374 VDDA.n201 GNDA 0.023309f
C2375 VDDA.n202 GNDA 0.033295f
C2376 VDDA.t380 GNDA 0.015197f
C2377 VDDA.t388 GNDA 0.015197f
C2378 VDDA.n203 GNDA 0.0524f
C2379 VDDA.n204 GNDA 0.090237f
C2380 VDDA.n205 GNDA 0.026408f
C2381 VDDA.t286 GNDA 0.022836f
C2382 VDDA.n206 GNDA 0.031153f
C2383 VDDA.n207 GNDA 0.016291f
C2384 VDDA.t370 GNDA 0.015197f
C2385 VDDA.n209 GNDA 0.033433f
C2386 VDDA.n211 GNDA 0.012157f
C2387 VDDA.n212 GNDA 0.033433f
C2388 VDDA.n213 GNDA 0.033433f
C2389 VDDA.t288 GNDA 0.015197f
C2390 VDDA.n215 GNDA 0.04559f
C2391 VDDA.n216 GNDA 0.032811f
C2392 VDDA.n218 GNDA 0.04559f
C2393 VDDA.n219 GNDA 0.026125f
C2394 VDDA.n221 GNDA 0.11899f
C2395 VDDA.t369 GNDA 0.107972f
C2396 VDDA.t378 GNDA 0.096955f
C2397 VDDA.t382 GNDA 0.096955f
C2398 VDDA.t38 GNDA 0.096955f
C2399 VDDA.t400 GNDA 0.096955f
C2400 VDDA.t342 GNDA 0.107972f
C2401 VDDA.n222 GNDA 0.012157f
C2402 VDDA.n224 GNDA 0.021461f
C2403 VDDA.n225 GNDA 0.021275f
C2404 VDDA.n226 GNDA 0.021275f
C2405 VDDA.n227 GNDA 0.012157f
C2406 VDDA.n228 GNDA 0.130007f
C2407 VDDA.n230 GNDA 0.02603f
C2408 VDDA.t341 GNDA 0.022836f
C2409 VDDA.n231 GNDA 0.031794f
C2410 VDDA.n232 GNDA 0.083391f
C2411 VDDA.n233 GNDA 0.093453f
C2412 VDDA.n234 GNDA 0.144311f
C2413 VDDA.t239 GNDA 0.021275f
C2414 VDDA.t249 GNDA 0.021275f
C2415 VDDA.n235 GNDA 0.073729f
C2416 VDDA.n236 GNDA 0.072159f
C2417 VDDA.t364 GNDA 0.021275f
C2418 VDDA.n237 GNDA 0.063826f
C2419 VDDA.n238 GNDA 0.021275f
C2420 VDDA.n239 GNDA 0.012157f
C2421 VDDA.n243 GNDA 0.012157f
C2422 VDDA.t292 GNDA 0.037303f
C2423 VDDA.t235 GNDA 0.021275f
C2424 VDDA.t231 GNDA 0.021275f
C2425 VDDA.n244 GNDA 0.073729f
C2426 VDDA.n245 GNDA 0.092386f
C2427 VDDA.n246 GNDA 0.031681f
C2428 VDDA.n247 GNDA 0.021275f
C2429 VDDA.n249 GNDA 0.021275f
C2430 VDDA.n250 GNDA 0.012157f
C2431 VDDA.n251 GNDA 0.012157f
C2432 VDDA.n252 GNDA 0.021275f
C2433 VDDA.n254 GNDA 0.021275f
C2434 VDDA.n255 GNDA 0.012157f
C2435 VDDA.n256 GNDA 0.012157f
C2436 VDDA.n257 GNDA 0.021275f
C2437 VDDA.n258 GNDA 0.021461f
C2438 VDDA.t294 GNDA 0.021275f
C2439 VDDA.n259 GNDA 0.063826f
C2440 VDDA.n260 GNDA 0.020509f
C2441 VDDA.n261 GNDA 0.012157f
C2442 VDDA.n262 GNDA 0.177801f
C2443 VDDA.t293 GNDA 0.154094f
C2444 VDDA.t234 GNDA 0.142241f
C2445 VDDA.t230 GNDA 0.142241f
C2446 VDDA.t238 GNDA 0.142241f
C2447 VDDA.t248 GNDA 0.142241f
C2448 VDDA.t258 GNDA 0.142241f
C2449 VDDA.t228 GNDA 0.142241f
C2450 VDDA.t226 GNDA 0.142241f
C2451 VDDA.t232 GNDA 0.142241f
C2452 VDDA.t240 GNDA 0.142241f
C2453 VDDA.t252 GNDA 0.142241f
C2454 VDDA.t363 GNDA 0.154094f
C2455 VDDA.n265 GNDA 0.012157f
C2456 VDDA.n267 GNDA 0.021461f
C2457 VDDA.n268 GNDA 0.021275f
C2458 VDDA.n269 GNDA 0.012157f
C2459 VDDA.n270 GNDA 0.012157f
C2460 VDDA.n271 GNDA 0.021275f
C2461 VDDA.n273 GNDA 0.021275f
C2462 VDDA.n274 GNDA 0.021275f
C2463 VDDA.n275 GNDA 0.012157f
C2464 VDDA.n276 GNDA 0.177801f
C2465 VDDA.n278 GNDA 0.023231f
C2466 VDDA.t362 GNDA 0.037303f
C2467 VDDA.n279 GNDA 0.031681f
C2468 VDDA.t241 GNDA 0.021275f
C2469 VDDA.t253 GNDA 0.021275f
C2470 VDDA.n280 GNDA 0.073729f
C2471 VDDA.n281 GNDA 0.092386f
C2472 VDDA.t227 GNDA 0.021275f
C2473 VDDA.t233 GNDA 0.021275f
C2474 VDDA.n282 GNDA 0.073729f
C2475 VDDA.n283 GNDA 0.072159f
C2476 VDDA.n284 GNDA 0.019452f
C2477 VDDA.t259 GNDA 0.021275f
C2478 VDDA.t229 GNDA 0.021275f
C2479 VDDA.n285 GNDA 0.072202f
C2480 VDDA.n286 GNDA 0.083176f
C2481 VDDA.t200 GNDA 0.018236f
C2482 VDDA.t265 GNDA 0.018236f
C2483 VDDA.n287 GNDA 0.075413f
C2484 VDDA.t40 GNDA 0.018236f
C2485 VDDA.t381 GNDA 0.018236f
C2486 VDDA.n288 GNDA 0.075124f
C2487 VDDA.n289 GNDA 0.104159f
C2488 VDDA.t203 GNDA 0.018236f
C2489 VDDA.t68 GNDA 0.018236f
C2490 VDDA.n290 GNDA 0.075124f
C2491 VDDA.n291 GNDA 0.054352f
C2492 VDDA.t96 GNDA 0.018236f
C2493 VDDA.t221 GNDA 0.018236f
C2494 VDDA.n292 GNDA 0.075124f
C2495 VDDA.n293 GNDA 0.054352f
C2496 VDDA.t409 GNDA 0.018236f
C2497 VDDA.t48 GNDA 0.018236f
C2498 VDDA.n294 GNDA 0.075124f
C2499 VDDA.n295 GNDA 0.054352f
C2500 VDDA.t264 GNDA 0.018236f
C2501 VDDA.t56 GNDA 0.018236f
C2502 VDDA.n296 GNDA 0.075124f
C2503 VDDA.n297 GNDA 0.1101f
C2504 VDDA.t332 GNDA 0.018376f
C2505 VDDA.n298 GNDA 0.012157f
C2506 VDDA.t334 GNDA 0.032052f
C2507 VDDA.n299 GNDA 0.012157f
C2508 VDDA.n300 GNDA 0.012157f
C2509 VDDA.n303 GNDA 0.012157f
C2510 VDDA.t347 GNDA 0.019205f
C2511 VDDA.n304 GNDA 0.021275f
C2512 VDDA.n305 GNDA 0.012157f
C2513 VDDA.n306 GNDA 0.021275f
C2514 VDDA.n307 GNDA 0.029601f
C2515 VDDA.t349 GNDA 0.032052f
C2516 VDDA.n309 GNDA 0.048665f
C2517 VDDA.n311 GNDA 0.107592f
C2518 VDDA.t348 GNDA 0.089356f
C2519 VDDA.t12 GNDA 0.080238f
C2520 VDDA.t377 GNDA 0.080238f
C2521 VDDA.t167 GNDA 0.080238f
C2522 VDDA.t69 GNDA 0.080238f
C2523 VDDA.t399 GNDA 0.080238f
C2524 VDDA.t412 GNDA 0.080238f
C2525 VDDA.t126 GNDA 0.080238f
C2526 VDDA.t166 GNDA 0.080238f
C2527 VDDA.t86 GNDA 0.080238f
C2528 VDDA.t214 GNDA 0.080238f
C2529 VDDA.t333 GNDA 0.089356f
C2530 VDDA.n312 GNDA 0.107592f
C2531 VDDA.n313 GNDA 0.012795f
C2532 VDDA.n314 GNDA 0.026799f
C2533 VDDA.n315 GNDA 0.021275f
C2534 VDDA.n316 GNDA 0.021275f
C2535 VDDA.n318 GNDA 0.024111f
C2536 VDDA.n319 GNDA 0.038962f
C2537 VDDA.n320 GNDA 0.171401f
C2538 VDDA.t394 GNDA 0.036472f
C2539 VDDA.t27 GNDA 0.036472f
C2540 VDDA.n321 GNDA 0.146321f
C2541 VDDA.n322 GNDA 0.074335f
C2542 VDDA.n324 GNDA 0.012157f
C2543 VDDA.n329 GNDA 0.012795f
C2544 VDDA.n335 GNDA 0.012795f
C2545 VDDA.n336 GNDA 0.012157f
C2546 VDDA.t295 GNDA 0.044192f
C2547 VDDA.t213 GNDA 0.036472f
C2548 VDDA.t95 GNDA 0.036472f
C2549 VDDA.n337 GNDA 0.146321f
C2550 VDDA.n338 GNDA 0.074335f
C2551 VDDA.t29 GNDA 0.036472f
C2552 VDDA.t165 GNDA 0.036472f
C2553 VDDA.n339 GNDA 0.146321f
C2554 VDDA.n340 GNDA 0.074335f
C2555 VDDA.t414 GNDA 0.036472f
C2556 VDDA.t169 GNDA 0.036472f
C2557 VDDA.n341 GNDA 0.146321f
C2558 VDDA.n342 GNDA 0.074335f
C2559 VDDA.t385 GNDA 0.036472f
C2560 VDDA.t202 GNDA 0.036472f
C2561 VDDA.n343 GNDA 0.146321f
C2562 VDDA.n344 GNDA 0.094066f
C2563 VDDA.n345 GNDA 0.036381f
C2564 VDDA.n346 GNDA 0.021275f
C2565 VDDA.n347 GNDA 0.012157f
C2566 VDDA.n348 GNDA 0.012157f
C2567 VDDA.n351 GNDA 0.012157f
C2568 VDDA.n352 GNDA 0.012157f
C2569 VDDA.n353 GNDA 0.024187f
C2570 VDDA.n354 GNDA 0.030795f
C2571 VDDA.n355 GNDA 0.012157f
C2572 VDDA.n356 GNDA 0.021275f
C2573 VDDA.n357 GNDA 0.021275f
C2574 VDDA.n358 GNDA 0.012157f
C2575 VDDA.n359 GNDA 0.012157f
C2576 VDDA.n360 GNDA 0.021275f
C2577 VDDA.n361 GNDA 0.021275f
C2578 VDDA.n362 GNDA 0.012157f
C2579 VDDA.n363 GNDA 0.012157f
C2580 VDDA.n364 GNDA 0.021275f
C2581 VDDA.n365 GNDA 0.021275f
C2582 VDDA.n366 GNDA 0.012157f
C2583 VDDA.n367 GNDA 0.012157f
C2584 VDDA.n368 GNDA 0.021275f
C2585 VDDA.n369 GNDA 0.021275f
C2586 VDDA.n370 GNDA 0.012157f
C2587 VDDA.n371 GNDA 0.012157f
C2588 VDDA.n372 GNDA 0.021275f
C2589 VDDA.n373 GNDA 0.024187f
C2590 VDDA.n375 GNDA 0.024111f
C2591 VDDA.n376 GNDA 0.012157f
C2592 VDDA.n377 GNDA 0.286913f
C2593 VDDA.t296 GNDA 0.238283f
C2594 VDDA.t201 GNDA 0.213969f
C2595 VDDA.t384 GNDA 0.213969f
C2596 VDDA.t168 GNDA 0.213969f
C2597 VDDA.t413 GNDA 0.213969f
C2598 VDDA.t164 GNDA 0.213969f
C2599 VDDA.t28 GNDA 0.213969f
C2600 VDDA.t94 GNDA 0.213969f
C2601 VDDA.t212 GNDA 0.213969f
C2602 VDDA.t26 GNDA 0.213969f
C2603 VDDA.t393 GNDA 0.213969f
C2604 VDDA.t272 GNDA 0.238283f
C2605 VDDA.n378 GNDA 0.012157f
C2606 VDDA.n379 GNDA 0.021275f
C2607 VDDA.n380 GNDA 0.024187f
C2608 VDDA.n381 GNDA 0.012157f
C2609 VDDA.n382 GNDA 0.012157f
C2610 VDDA.n385 GNDA 0.012157f
C2611 VDDA.n386 GNDA 0.012157f
C2612 VDDA.n387 GNDA 0.024187f
C2613 VDDA.n388 GNDA 0.030795f
C2614 VDDA.n389 GNDA 0.012157f
C2615 VDDA.n390 GNDA 0.021275f
C2616 VDDA.n391 GNDA 0.021275f
C2617 VDDA.n392 GNDA 0.012157f
C2618 VDDA.n393 GNDA 0.012157f
C2619 VDDA.n394 GNDA 0.021275f
C2620 VDDA.n395 GNDA 0.021275f
C2621 VDDA.n396 GNDA 0.012157f
C2622 VDDA.n397 GNDA 0.012157f
C2623 VDDA.n398 GNDA 0.021275f
C2624 VDDA.n399 GNDA 0.021275f
C2625 VDDA.n400 GNDA 0.012157f
C2626 VDDA.n401 GNDA 0.012157f
C2627 VDDA.n402 GNDA 0.021275f
C2628 VDDA.n403 GNDA 0.021275f
C2629 VDDA.n404 GNDA 0.021275f
C2630 VDDA.n405 GNDA 0.012157f
C2631 VDDA.n406 GNDA 0.286913f
C2632 VDDA.n408 GNDA 0.026833f
C2633 VDDA.t271 GNDA 0.044192f
C2634 VDDA.n409 GNDA 0.035577f
C2635 VDDA.n410 GNDA 0.049454f
C2636 VDDA.n411 GNDA 0.128574f
C2637 VDDA.n412 GNDA 0.148804f
C2638 VDDA.n413 GNDA 0.132984f
C2639 VDDA.t408 GNDA 0.010942f
C2640 VDDA.t309 GNDA 0.010942f
C2641 VDDA.n414 GNDA 0.025388f
C2642 VDDA.n415 GNDA 0.082369f
C2643 VDDA.t300 GNDA 0.038822f
C2644 VDDA.t307 GNDA 0.022445f
C2645 VDDA.n416 GNDA 0.044399f
C2646 VDDA.t310 GNDA 0.038822f
C2647 VDDA.n417 GNDA 0.072884f
C2648 VDDA.t308 GNDA 0.130082f
C2649 VDDA.t407 GNDA 0.080238f
C2650 VDDA.t299 GNDA 0.130082f
C2651 VDDA.n418 GNDA 0.072884f
C2652 VDDA.t298 GNDA 0.022445f
C2653 VDDA.n419 GNDA 0.044088f
C2654 VDDA.n420 GNDA 0.041251f
C2655 VDDA.n421 GNDA 0.058445f
C2656 VDDA.n422 GNDA 0.085697f
C2657 VDDA.t358 GNDA 0.021275f
C2658 VDDA.n423 GNDA 0.063826f
C2659 VDDA.n424 GNDA 0.021275f
C2660 VDDA.n425 GNDA 0.012157f
C2661 VDDA.n429 GNDA 0.012157f
C2662 VDDA.t329 GNDA 0.037303f
C2663 VDDA.n430 GNDA 0.031076f
C2664 VDDA.n431 GNDA 0.021275f
C2665 VDDA.n433 GNDA 0.021275f
C2666 VDDA.n434 GNDA 0.012157f
C2667 VDDA.n435 GNDA 0.012157f
C2668 VDDA.n436 GNDA 0.021275f
C2669 VDDA.n438 GNDA 0.021275f
C2670 VDDA.n439 GNDA 0.012157f
C2671 VDDA.n440 GNDA 0.012157f
C2672 VDDA.n441 GNDA 0.021275f
C2673 VDDA.n442 GNDA 0.021461f
C2674 VDDA.t251 GNDA 0.021275f
C2675 VDDA.n443 GNDA 0.073729f
C2676 VDDA.t331 GNDA 0.042551f
C2677 VDDA.n444 GNDA 0.063826f
C2678 VDDA.n445 GNDA 0.020509f
C2679 VDDA.n446 GNDA 0.012157f
C2680 VDDA.n447 GNDA 0.177801f
C2681 VDDA.t330 GNDA 0.154094f
C2682 VDDA.t250 GNDA 0.142241f
C2683 VDDA.t357 GNDA 0.154094f
C2684 VDDA.n450 GNDA 0.012157f
C2685 VDDA.n452 GNDA 0.021461f
C2686 VDDA.n453 GNDA 0.021275f
C2687 VDDA.n454 GNDA 0.012157f
C2688 VDDA.n455 GNDA 0.012157f
C2689 VDDA.n456 GNDA 0.021275f
C2690 VDDA.n458 GNDA 0.021275f
C2691 VDDA.n459 GNDA 0.021275f
C2692 VDDA.n460 GNDA 0.012157f
C2693 VDDA.n461 GNDA 0.177801f
C2694 VDDA.n463 GNDA 0.023231f
C2695 VDDA.t356 GNDA 0.037303f
C2696 VDDA.n464 GNDA 0.030765f
C2697 VDDA.n465 GNDA 0.041251f
C2698 VDDA.n466 GNDA 0.172485f
C2699 VDDA.n467 GNDA 3.26626f
C2700 VDDA.t114 GNDA 0.339797f
C2701 VDDA.t37 GNDA 0.341029f
C2702 VDDA.t107 GNDA 0.322793f
C2703 VDDA.t63 GNDA 0.339797f
C2704 VDDA.t23 GNDA 0.341029f
C2705 VDDA.t42 GNDA 0.322793f
C2706 VDDA.t41 GNDA 0.339797f
C2707 VDDA.t99 GNDA 0.341029f
C2708 VDDA.t100 GNDA 0.322793f
C2709 VDDA.t189 GNDA 0.339797f
C2710 VDDA.t206 GNDA 0.341029f
C2711 VDDA.t34 GNDA 0.322793f
C2712 VDDA.t162 GNDA 0.339797f
C2713 VDDA.t108 GNDA 0.341029f
C2714 VDDA.t22 GNDA 0.322793f
C2715 VDDA.n468 GNDA 0.227766f
C2716 VDDA.t163 GNDA 0.181382f
C2717 VDDA.n469 GNDA 0.247132f
C2718 VDDA.t21 GNDA 0.181382f
C2719 VDDA.n470 GNDA 0.247132f
C2720 VDDA.t43 GNDA 0.181382f
C2721 VDDA.n471 GNDA 0.247132f
C2722 VDDA.t188 GNDA 0.181382f
C2723 VDDA.n472 GNDA 0.247132f
C2724 VDDA.t115 GNDA 0.317752f
C2725 VDDA.n473 GNDA 2.82193f
C2726 VDDA.t415 GNDA 0.672021f
C2727 VDDA.t417 GNDA 0.716246f
C2728 VDDA.t418 GNDA 0.715966f
C2729 VDDA.t416 GNDA 0.689013f
C2730 VDDA.n474 GNDA 0.479624f
C2731 VDDA.n475 GNDA 0.235533f
C2732 VDDA.n476 GNDA 0.342366f
C2733 VDDA.n477 GNDA 0.624948f
C2734 VDDA.n478 GNDA 0.015289f
C2735 VDDA.n479 GNDA 0.06191f
C2736 VDDA.n480 GNDA 0.025708f
C2737 VDDA.t322 GNDA 0.021144f
C2738 VDDA.n482 GNDA 0.025708f
C2739 VDDA.n483 GNDA 0.015289f
C2740 VDDA.n484 GNDA 0.06191f
C2741 VDDA.t306 GNDA 0.021291f
C2742 VDDA.n485 GNDA 0.025708f
C2743 VDDA.n486 GNDA 0.015289f
C2744 VDDA.n487 GNDA 0.06191f
C2745 VDDA.n488 GNDA 0.015289f
C2746 VDDA.n489 GNDA 0.06191f
C2747 VDDA.n490 GNDA 0.015289f
C2748 VDDA.n491 GNDA 0.06191f
C2749 VDDA.n492 GNDA 0.015289f
C2750 VDDA.n493 GNDA 0.06191f
C2751 VDDA.n494 GNDA 0.015289f
C2752 VDDA.n495 GNDA 0.06191f
C2753 VDDA.n496 GNDA 0.015289f
C2754 VDDA.n497 GNDA 0.06191f
C2755 VDDA.n498 GNDA 0.015289f
C2756 VDDA.n499 GNDA 0.06191f
C2757 VDDA.n500 GNDA 0.015289f
C2758 VDDA.n501 GNDA 0.088968f
C2759 VDDA.n502 GNDA 0.023571f
C2760 VDDA.t280 GNDA 0.022439f
C2761 VDDA.t282 GNDA 0.021144f
C2762 VDDA.n503 GNDA 0.040529f
C2763 VDDA.n504 GNDA 0.061608f
C2764 VDDA.t281 GNDA 0.076405f
C2765 VDDA.t136 GNDA 0.051061f
C2766 VDDA.t138 GNDA 0.051061f
C2767 VDDA.t24 GNDA 0.051061f
C2768 VDDA.t2 GNDA 0.051061f
C2769 VDDA.t176 GNDA 0.051061f
C2770 VDDA.t178 GNDA 0.051061f
C2771 VDDA.t401 GNDA 0.051061f
C2772 VDDA.t15 GNDA 0.051061f
C2773 VDDA.t128 GNDA 0.051061f
C2774 VDDA.t82 GNDA 0.051061f
C2775 VDDA.t0 GNDA 0.051061f
C2776 VDDA.t180 GNDA 0.051061f
C2777 VDDA.t389 GNDA 0.051061f
C2778 VDDA.t80 GNDA 0.051061f
C2779 VDDA.t391 GNDA 0.051061f
C2780 VDDA.t184 GNDA 0.051061f
C2781 VDDA.t182 GNDA 0.051061f
C2782 VDDA.t78 GNDA 0.051061f
C2783 VDDA.t305 GNDA 0.077886f
C2784 VDDA.n505 GNDA 0.1109f
C2785 VDDA.t304 GNDA 0.015047f
C2786 VDDA.n506 GNDA 0.024866f
C2787 VDDA.n507 GNDA 0.04528f
C2788 VDDA.n508 GNDA 0.015289f
C2789 VDDA.n509 GNDA 0.06191f
C2790 VDDA.n510 GNDA 0.015289f
C2791 VDDA.n511 GNDA 0.06191f
C2792 VDDA.n512 GNDA 0.015289f
C2793 VDDA.n513 GNDA 0.06191f
C2794 VDDA.n514 GNDA 0.015289f
C2795 VDDA.n515 GNDA 0.06191f
C2796 VDDA.n516 GNDA 0.015289f
C2797 VDDA.n517 GNDA 0.06191f
C2798 VDDA.n518 GNDA 0.015289f
C2799 VDDA.n519 GNDA 0.06191f
C2800 VDDA.n520 GNDA 0.015289f
C2801 VDDA.n521 GNDA 0.06191f
C2802 VDDA.n522 GNDA 0.015289f
C2803 VDDA.n523 GNDA 0.06191f
C2804 VDDA.n524 GNDA 0.04528f
C2805 VDDA.n525 GNDA 0.022369f
C2806 VDDA.t338 GNDA 0.022439f
C2807 VDDA.t340 GNDA 0.021144f
C2808 VDDA.n526 GNDA 0.040529f
C2809 VDDA.n527 GNDA 0.061608f
C2810 VDDA.t339 GNDA 0.076405f
C2811 VDDA.t403 GNDA 0.051061f
C2812 VDDA.t57 GNDA 0.051061f
C2813 VDDA.t4 GNDA 0.051061f
C2814 VDDA.t196 GNDA 0.051061f
C2815 VDDA.t219 GNDA 0.051061f
C2816 VDDA.t405 GNDA 0.051061f
C2817 VDDA.t110 GNDA 0.051061f
C2818 VDDA.t170 GNDA 0.051061f
C2819 VDDA.t8 GNDA 0.051061f
C2820 VDDA.t30 GNDA 0.051061f
C2821 VDDA.t44 GNDA 0.051061f
C2822 VDDA.t410 GNDA 0.051061f
C2823 VDDA.t19 GNDA 0.051061f
C2824 VDDA.t122 GNDA 0.051061f
C2825 VDDA.t124 GNDA 0.051061f
C2826 VDDA.t10 GNDA 0.051061f
C2827 VDDA.t87 GNDA 0.051061f
C2828 VDDA.t17 GNDA 0.051061f
C2829 VDDA.t321 GNDA 0.063083f
C2830 VDDA.n528 GNDA 0.074929f
C2831 VDDA.n529 GNDA 0.040693f
C2832 VDDA.t320 GNDA 0.022428f
C2833 VDDA.n530 GNDA 0.022369f
C2834 VDDA.n531 GNDA 0.10494f
C2835 VDDA.n532 GNDA 0.202331f
C2836 VDDA.t205 GNDA 0.018236f
C2837 VDDA.t98 GNDA 0.018236f
C2838 VDDA.n533 GNDA 0.060246f
C2839 VDDA.n534 GNDA 0.077739f
C2840 VDDA.n536 GNDA 0.012157f
C2841 VDDA.n539 GNDA 0.012157f
C2842 VDDA.n540 GNDA 0.012157f
C2843 VDDA.n541 GNDA 0.021148f
C2844 VDDA.n542 GNDA 0.012157f
C2845 VDDA.n543 GNDA 0.012157f
C2846 VDDA.n544 GNDA 0.012157f
C2847 VDDA.n545 GNDA 0.021275f
C2848 VDDA.t301 GNDA 0.086957f
C2849 VDDA.t335 GNDA 0.011524f
C2850 VDDA.n546 GNDA 0.029861f
C2851 VDDA.t376 GNDA 0.02427f
C2852 VDDA.t337 GNDA 0.021291f
C2853 VDDA.n547 GNDA 0.106516f
C2854 VDDA.t336 GNDA 0.07376f
C2855 VDDA.t55 GNDA 0.046806f
C2856 VDDA.t127 GNDA 0.046806f
C2857 VDDA.t375 GNDA 0.075384f
C2858 VDDA.n548 GNDA 0.111556f
C2859 VDDA.t374 GNDA 0.011524f
C2860 VDDA.n549 GNDA 0.029634f
C2861 VDDA.n550 GNDA 0.089143f
C2862 VDDA.t113 GNDA 0.018236f
C2863 VDDA.t106 GNDA 0.018236f
C2864 VDDA.n551 GNDA 0.060246f
C2865 VDDA.n552 GNDA 0.077739f
C2866 VDDA.t60 GNDA 0.018236f
C2867 VDDA.t62 GNDA 0.018236f
C2868 VDDA.n553 GNDA 0.060246f
C2869 VDDA.n554 GNDA 0.077739f
C2870 VDDA.t104 GNDA 0.018236f
C2871 VDDA.t143 GNDA 0.018236f
C2872 VDDA.n555 GNDA 0.060246f
C2873 VDDA.n556 GNDA 0.077739f
C2874 VDDA.t141 GNDA 0.018236f
C2875 VDDA.t117 GNDA 0.018236f
C2876 VDDA.n557 GNDA 0.060246f
C2877 VDDA.n558 GNDA 0.077739f
C2878 VDDA.t102 GNDA 0.018236f
C2879 VDDA.t208 GNDA 0.018236f
C2880 VDDA.n559 GNDA 0.060246f
C2881 VDDA.n560 GNDA 0.077739f
C2882 VDDA.t187 GNDA 0.018236f
C2883 VDDA.t36 GNDA 0.018236f
C2884 VDDA.n561 GNDA 0.060246f
C2885 VDDA.n562 GNDA 0.077739f
C2886 VDDA.t145 GNDA 0.018236f
C2887 VDDA.t161 GNDA 0.018236f
C2888 VDDA.n563 GNDA 0.060246f
C2889 VDDA.n564 GNDA 0.077739f
C2890 VDDA.n565 GNDA 0.041507f
C2891 VDDA.n566 GNDA 0.032475f
C2892 VDDA.n567 GNDA 0.024111f
C2893 VDDA.n569 GNDA 0.021148f
C2894 VDDA.n570 GNDA 0.021275f
C2895 VDDA.n571 GNDA 0.021275f
C2896 VDDA.n572 GNDA 0.021275f
C2897 VDDA.n573 GNDA 0.030795f
C2898 VDDA.n574 GNDA 0.012795f
C2899 VDDA.n575 GNDA 0.170506f
C2900 VDDA.t302 GNDA 0.18084f
C2901 VDDA.t144 GNDA 0.186007f
C2902 VDDA.t160 GNDA 0.186007f
C2903 VDDA.t186 GNDA 0.186007f
C2904 VDDA.t35 GNDA 0.186007f
C2905 VDDA.t101 GNDA 0.186007f
C2906 VDDA.t207 GNDA 0.186007f
C2907 VDDA.t140 GNDA 0.186007f
C2908 VDDA.t116 GNDA 0.186007f
C2909 VDDA.t103 GNDA 0.186007f
C2910 VDDA.t142 GNDA 0.186007f
C2911 VDDA.t59 GNDA 0.186007f
C2912 VDDA.t61 GNDA 0.186007f
C2913 VDDA.t112 GNDA 0.186007f
C2914 VDDA.t105 GNDA 0.186007f
C2915 VDDA.t204 GNDA 0.186007f
C2916 VDDA.t97 GNDA 0.186007f
C2917 VDDA.t269 GNDA 0.18084f
C2918 VDDA.n577 GNDA 0.012157f
C2919 VDDA.n578 GNDA 0.012157f
C2920 VDDA.n579 GNDA 0.021275f
C2921 VDDA.n580 GNDA 0.021148f
C2922 VDDA.n581 GNDA 0.021275f
C2923 VDDA.n582 GNDA 0.012157f
C2924 VDDA.n583 GNDA 0.021275f
C2925 VDDA.n584 GNDA 0.021275f
C2926 VDDA.n585 GNDA 0.021148f
C2927 VDDA.n586 GNDA 0.033597f
C2928 VDDA.n588 GNDA 0.170506f
C2929 VDDA.n589 GNDA 0.012157f
C2930 VDDA.n590 GNDA 0.024111f
C2931 VDDA.t268 GNDA 0.086957f
C2932 VDDA.n591 GNDA 0.032475f
C2933 VDDA.n592 GNDA 0.047889f
C2934 VDDA.t317 GNDA 0.011226f
C2935 VDDA.n593 GNDA 0.023987f
C2936 VDDA.t316 GNDA 0.021291f
C2937 VDDA.t319 GNDA 0.021291f
C2938 VDDA.n594 GNDA 0.105916f
C2939 VDDA.t318 GNDA 0.07376f
C2940 VDDA.t84 GNDA 0.046806f
C2941 VDDA.t174 GNDA 0.046806f
C2942 VDDA.t315 GNDA 0.07376f
C2943 VDDA.n595 GNDA 0.105916f
C2944 VDDA.t314 GNDA 0.011226f
C2945 VDDA.n596 GNDA 0.023987f
C2946 VDDA.n597 GNDA 0.057698f
C2947 VDDA.n598 GNDA 0.01466f
C2948 VDDA.n599 GNDA 0.051475f
C2949 VDDA.n600 GNDA 0.119522f
C2950 VDDA.n601 GNDA 0.165081f
C2951 VDDA.n602 GNDA 0.015163f
C2952 VDDA.n603 GNDA 0.053525f
C2953 VDDA.t361 GNDA 0.022162f
C2954 VDDA.t285 GNDA 0.022162f
C2955 VDDA.t283 GNDA 0.011971f
C2956 VDDA.n604 GNDA 0.015135f
C2957 VDDA.n605 GNDA 0.053554f
C2958 VDDA.t365 GNDA 0.011971f
C2959 VDDA.n606 GNDA 0.01517f
C2960 VDDA.n607 GNDA 0.053519f
C2961 VDDA.t276 GNDA 0.022173f
C2962 VDDA.t352 GNDA 0.022173f
C2963 VDDA.t350 GNDA 0.011971f
C2964 VDDA.n608 GNDA 0.01517f
C2965 VDDA.n609 GNDA 0.07325f
C2966 VDDA.n610 GNDA 0.025424f
C2967 VDDA.n611 GNDA 0.063275f
C2968 VDDA.t351 GNDA 0.066683f
C2969 VDDA.t210 GNDA 0.046806f
C2970 VDDA.t192 GNDA 0.046806f
C2971 VDDA.t172 GNDA 0.046806f
C2972 VDDA.t120 GNDA 0.046806f
C2973 VDDA.t275 GNDA 0.066683f
C2974 VDDA.n612 GNDA 0.063275f
C2975 VDDA.t274 GNDA 0.012351f
C2976 VDDA.n613 GNDA 0.025f
C2977 VDDA.n614 GNDA 0.036948f
C2978 VDDA.n615 GNDA 0.015135f
C2979 VDDA.n616 GNDA 0.053554f
C2980 VDDA.n617 GNDA 0.015135f
C2981 VDDA.n618 GNDA 0.053554f
C2982 VDDA.n619 GNDA 0.015135f
C2983 VDDA.n620 GNDA 0.053554f
C2984 VDDA.n621 GNDA 0.015135f
C2985 VDDA.n622 GNDA 0.053554f
C2986 VDDA.n623 GNDA 0.036948f
C2987 VDDA.n624 GNDA 0.02365f
C2988 VDDA.t367 GNDA 0.021248f
C2989 VDDA.n625 GNDA 0.064999f
C2990 VDDA.t366 GNDA 0.066854f
C2991 VDDA.t64 GNDA 0.046806f
C2992 VDDA.t395 GNDA 0.046806f
C2993 VDDA.t217 GNDA 0.046806f
C2994 VDDA.t32 GNDA 0.046806f
C2995 VDDA.t397 GNDA 0.046806f
C2996 VDDA.t46 GNDA 0.046806f
C2997 VDDA.t198 GNDA 0.046806f
C2998 VDDA.t118 GNDA 0.046806f
C2999 VDDA.t194 GNDA 0.046806f
C3000 VDDA.t190 GNDA 0.046806f
C3001 VDDA.t345 GNDA 0.066854f
C3002 VDDA.t346 GNDA 0.021248f
C3003 VDDA.n626 GNDA 0.064999f
C3004 VDDA.t344 GNDA 0.011971f
C3005 VDDA.n627 GNDA 0.02365f
C3006 VDDA.n628 GNDA 0.036948f
C3007 VDDA.n629 GNDA 0.015163f
C3008 VDDA.n630 GNDA 0.053525f
C3009 VDDA.n631 GNDA 0.036948f
C3010 VDDA.n632 GNDA 0.02462f
C3011 VDDA.n633 GNDA 0.063286f
C3012 VDDA.t284 GNDA 0.066683f
C3013 VDDA.t215 GNDA 0.046806f
C3014 VDDA.t6 GNDA 0.046806f
C3015 VDDA.t53 GNDA 0.046806f
C3016 VDDA.t66 GNDA 0.046806f
C3017 VDDA.t360 GNDA 0.066683f
C3018 VDDA.n634 GNDA 0.063286f
C3019 VDDA.t359 GNDA 0.011971f
C3020 VDDA.n635 GNDA 0.02462f
C3021 VDDA.n636 GNDA 0.122923f
C3022 VDDA.n637 GNDA 0.143507f
C3023 VDDA.n638 GNDA 0.68414f
C3024 two_stage_opamp_dummy_magic_16_0.Vb3.t2 GNDA 0.014599f
C3025 two_stage_opamp_dummy_magic_16_0.Vb3.t6 GNDA 0.014599f
C3026 two_stage_opamp_dummy_magic_16_0.Vb3.n0 GNDA 0.047024f
C3027 two_stage_opamp_dummy_magic_16_0.Vb3.t5 GNDA 0.014599f
C3028 two_stage_opamp_dummy_magic_16_0.Vb3.t0 GNDA 0.014599f
C3029 two_stage_opamp_dummy_magic_16_0.Vb3.n1 GNDA 0.047024f
C3030 two_stage_opamp_dummy_magic_16_0.Vb3.n2 GNDA 0.25924f
C3031 two_stage_opamp_dummy_magic_16_0.Vb3.t4 GNDA 0.014599f
C3032 two_stage_opamp_dummy_magic_16_0.Vb3.t3 GNDA 0.014599f
C3033 two_stage_opamp_dummy_magic_16_0.Vb3.n3 GNDA 0.044094f
C3034 two_stage_opamp_dummy_magic_16_0.Vb3.n4 GNDA 0.785193f
C3035 two_stage_opamp_dummy_magic_16_0.Vb3.t1 GNDA 0.051095f
C3036 two_stage_opamp_dummy_magic_16_0.Vb3.t7 GNDA 0.051095f
C3037 two_stage_opamp_dummy_magic_16_0.Vb3.n5 GNDA 0.180135f
C3038 two_stage_opamp_dummy_magic_16_0.Vb3.t28 GNDA 0.072263f
C3039 two_stage_opamp_dummy_magic_16_0.Vb3.t9 GNDA 0.072263f
C3040 two_stage_opamp_dummy_magic_16_0.Vb3.t12 GNDA 0.072263f
C3041 two_stage_opamp_dummy_magic_16_0.Vb3.t18 GNDA 0.072263f
C3042 two_stage_opamp_dummy_magic_16_0.Vb3.t16 GNDA 0.083391f
C3043 two_stage_opamp_dummy_magic_16_0.Vb3.n6 GNDA 0.067705f
C3044 two_stage_opamp_dummy_magic_16_0.Vb3.n7 GNDA 0.041606f
C3045 two_stage_opamp_dummy_magic_16_0.Vb3.n8 GNDA 0.041606f
C3046 two_stage_opamp_dummy_magic_16_0.Vb3.n9 GNDA 0.038604f
C3047 two_stage_opamp_dummy_magic_16_0.Vb3.t27 GNDA 0.072263f
C3048 two_stage_opamp_dummy_magic_16_0.Vb3.t21 GNDA 0.072263f
C3049 two_stage_opamp_dummy_magic_16_0.Vb3.t17 GNDA 0.072263f
C3050 two_stage_opamp_dummy_magic_16_0.Vb3.t11 GNDA 0.072263f
C3051 two_stage_opamp_dummy_magic_16_0.Vb3.t8 GNDA 0.083391f
C3052 two_stage_opamp_dummy_magic_16_0.Vb3.n10 GNDA 0.067705f
C3053 two_stage_opamp_dummy_magic_16_0.Vb3.n11 GNDA 0.041606f
C3054 two_stage_opamp_dummy_magic_16_0.Vb3.n12 GNDA 0.041606f
C3055 two_stage_opamp_dummy_magic_16_0.Vb3.n13 GNDA 0.038604f
C3056 two_stage_opamp_dummy_magic_16_0.Vb3.n14 GNDA 0.040946f
C3057 two_stage_opamp_dummy_magic_16_0.Vb3.t10 GNDA 0.072263f
C3058 two_stage_opamp_dummy_magic_16_0.Vb3.t15 GNDA 0.072263f
C3059 two_stage_opamp_dummy_magic_16_0.Vb3.t20 GNDA 0.072263f
C3060 two_stage_opamp_dummy_magic_16_0.Vb3.t24 GNDA 0.072263f
C3061 two_stage_opamp_dummy_magic_16_0.Vb3.t22 GNDA 0.083391f
C3062 two_stage_opamp_dummy_magic_16_0.Vb3.n15 GNDA 0.067705f
C3063 two_stage_opamp_dummy_magic_16_0.Vb3.n16 GNDA 0.041606f
C3064 two_stage_opamp_dummy_magic_16_0.Vb3.n17 GNDA 0.041606f
C3065 two_stage_opamp_dummy_magic_16_0.Vb3.n18 GNDA 0.038604f
C3066 two_stage_opamp_dummy_magic_16_0.Vb3.t25 GNDA 0.072263f
C3067 two_stage_opamp_dummy_magic_16_0.Vb3.t26 GNDA 0.072263f
C3068 two_stage_opamp_dummy_magic_16_0.Vb3.t23 GNDA 0.072263f
C3069 two_stage_opamp_dummy_magic_16_0.Vb3.t19 GNDA 0.072263f
C3070 two_stage_opamp_dummy_magic_16_0.Vb3.t13 GNDA 0.083391f
C3071 two_stage_opamp_dummy_magic_16_0.Vb3.n19 GNDA 0.067705f
C3072 two_stage_opamp_dummy_magic_16_0.Vb3.n20 GNDA 0.041606f
C3073 two_stage_opamp_dummy_magic_16_0.Vb3.n21 GNDA 0.041606f
C3074 two_stage_opamp_dummy_magic_16_0.Vb3.n22 GNDA 0.038604f
C3075 two_stage_opamp_dummy_magic_16_0.Vb3.n23 GNDA 0.04262f
C3076 two_stage_opamp_dummy_magic_16_0.Vb3.n24 GNDA 1.17334f
C3077 two_stage_opamp_dummy_magic_16_0.Vb3.t14 GNDA 0.08858f
C3078 two_stage_opamp_dummy_magic_16_0.Vb3.n25 GNDA 0.307922f
C3079 two_stage_opamp_dummy_magic_16_0.Vb3.n26 GNDA 0.912484f
C3080 bgr_0.VB3_CUR_BIAS GNDA 1.63375f
C3081 bgr_0.NFET_GATE_10uA.t4 GNDA 0.01496f
C3082 bgr_0.NFET_GATE_10uA.t3 GNDA 0.01496f
C3083 bgr_0.NFET_GATE_10uA.n0 GNDA 0.042091f
C3084 bgr_0.NFET_GATE_10uA.t18 GNDA 0.014586f
C3085 bgr_0.NFET_GATE_10uA.t6 GNDA 0.014586f
C3086 bgr_0.NFET_GATE_10uA.t14 GNDA 0.014586f
C3087 bgr_0.NFET_GATE_10uA.t19 GNDA 0.014586f
C3088 bgr_0.NFET_GATE_10uA.t5 GNDA 0.014586f
C3089 bgr_0.NFET_GATE_10uA.t13 GNDA 0.014586f
C3090 bgr_0.NFET_GATE_10uA.t12 GNDA 0.021563f
C3091 bgr_0.NFET_GATE_10uA.n1 GNDA 0.026685f
C3092 bgr_0.NFET_GATE_10uA.n2 GNDA 0.019075f
C3093 bgr_0.NFET_GATE_10uA.n3 GNDA 0.016149f
C3094 bgr_0.NFET_GATE_10uA.t15 GNDA 0.014586f
C3095 bgr_0.NFET_GATE_10uA.t8 GNDA 0.014586f
C3096 bgr_0.NFET_GATE_10uA.t21 GNDA 0.014586f
C3097 bgr_0.NFET_GATE_10uA.t16 GNDA 0.021563f
C3098 bgr_0.NFET_GATE_10uA.n4 GNDA 0.026685f
C3099 bgr_0.NFET_GATE_10uA.n5 GNDA 0.019075f
C3100 bgr_0.NFET_GATE_10uA.n6 GNDA 0.016149f
C3101 bgr_0.NFET_GATE_10uA.t20 GNDA 0.014586f
C3102 bgr_0.NFET_GATE_10uA.t7 GNDA 0.021563f
C3103 bgr_0.NFET_GATE_10uA.n7 GNDA 0.02376f
C3104 bgr_0.NFET_GATE_10uA.n8 GNDA 0.026114f
C3105 bgr_0.NFET_GATE_10uA.t11 GNDA 0.014586f
C3106 bgr_0.NFET_GATE_10uA.t22 GNDA 0.021563f
C3107 bgr_0.NFET_GATE_10uA.n9 GNDA 0.02376f
C3108 bgr_0.NFET_GATE_10uA.t9 GNDA 0.014586f
C3109 bgr_0.NFET_GATE_10uA.t17 GNDA 0.014586f
C3110 bgr_0.NFET_GATE_10uA.t23 GNDA 0.014586f
C3111 bgr_0.NFET_GATE_10uA.t10 GNDA 0.021563f
C3112 bgr_0.NFET_GATE_10uA.n10 GNDA 0.026685f
C3113 bgr_0.NFET_GATE_10uA.n11 GNDA 0.019075f
C3114 bgr_0.NFET_GATE_10uA.n12 GNDA 0.016149f
C3115 bgr_0.NFET_GATE_10uA.n13 GNDA 0.026114f
C3116 bgr_0.NFET_GATE_10uA.n14 GNDA 0.605807f
C3117 bgr_0.NFET_GATE_10uA.n15 GNDA 0.022264f
C3118 bgr_0.NFET_GATE_10uA.n16 GNDA 0.016149f
C3119 bgr_0.NFET_GATE_10uA.n17 GNDA 0.019075f
C3120 bgr_0.NFET_GATE_10uA.n18 GNDA 0.026685f
C3121 bgr_0.NFET_GATE_10uA.t2 GNDA 0.034164f
C3122 bgr_0.NFET_GATE_10uA.n19 GNDA 0.327308f
C3123 bgr_0.NFET_GATE_10uA.t1 GNDA 0.01496f
C3124 bgr_0.NFET_GATE_10uA.t0 GNDA 0.01496f
C3125 bgr_0.NFET_GATE_10uA.n20 GNDA 0.088541f
.ends

