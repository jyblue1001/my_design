* NGSPICE file created from two_stage_opamp_dummy_magic_24.ext - technology: sky130A

.subckt two_stage_opamp_dummy_magic_24 V_CMFB_S1 V_CMFB_S3 Vb3 Vb2 V_CMFB_S2 V_CMFB_S4
+ VOUT- VOUT+ V_tail_gate V_err_amp_ref V_err_gate
X0 VD4 Vb2 Y VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1 w_109520_3890# V_err_gate V_err_mir_p w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X2 a_109560_2850# a_112630_1380# V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X3 w_109520_3890# Vb3 VD3 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X4 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 a_109560_2850# a_109560_2850# w_109520_3890# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X7 VD2 Vb1 Y a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X8 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X11 VD1 Vb1 X a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X12 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X14 w_109520_3890# X VOUT- w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X15 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 a_109560_2850# Y V_CMFB_S3 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X19 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 w_109520_3890# w_109520_3890# VD3 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X21 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X23 V_p_mir a_112630_1380# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X24 w_109520_3890# Y V_CMFB_S4 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X25 Y Vb1 VD2 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X26 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 a_118250_3658# V_CMFB_S2 a_109560_2850# sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X28 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X29 w_109520_3890# X V_CMFB_S2 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X30 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 a_109560_2850# a_109560_2850# err_amp_out a_109560_2850# sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X34 a_109560_2850# w_109520_3890# w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X35 VD2 VIN+ V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X36 VD4 Vb2 Y VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X37 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 w_109520_3890# w_109520_3890# a_109560_2850# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X40 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X41 VD1 VIN- V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X42 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 w_109520_3890# w_109520_3890# a_109560_2850# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X46 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 VOUT+ a_109200_146# a_109560_2850# sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X48 V_CMFB_S4 Y w_109520_3890# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X49 a_108920_3658# V_CMFB_S4 a_109560_2850# sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X50 V_err_gate w_109520_3890# w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X51 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 Vb1 Vb1 a_113080_300# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X53 VD3 Vb2 X VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X54 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 V_CMFB_S2 X w_109520_3890# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X56 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X57 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X58 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 VD1 Vb1 X a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X60 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X62 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X63 w_109520_3890# X VOUT- w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X64 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X65 a_109560_2850# Y V_CMFB_S3 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X66 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X69 V_source Vb1 a_113080_300# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.6 ps=3.8 w=1.5 l=3
X70 a_109560_2850# X V_CMFB_S1 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X71 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 V_source a_112630_1380# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X73 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 w_109520_3890# Vb3 VD4 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X75 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X77 a_109560_2850# V_b_2nd_stage VOUT- a_109560_2850# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X78 a_109560_2850# err_amp_mir err_amp_mir a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X79 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X80 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X81 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X82 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X86 VD2 VIN+ V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X87 VD1 VIN- V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X88 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 VD1 VIN- V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X90 V_CMFB_S3 Y a_109560_2850# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X91 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X92 cap_res_Y Y a_109560_2850# sky130_fd_pr__res_high_po_1p41 l=1.41
X93 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X94 a_109560_2850# a_112630_1380# V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X95 V_CMFB_S1 X a_109560_2850# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X96 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X98 w_109520_3890# w_109520_3890# err_amp_out w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X99 Vb2_Vb3 Vb2_Vb3 Vb2_Vb3 Vb2_Vb3 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=5.6 ps=31.2 w=3.5 l=0.2
X100 V_CMFB_S2 X w_109520_3890# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X101 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X102 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X103 VD1 Vb1 X a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X104 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X106 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 VOUT- a_109560_2850# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X109 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X110 V_source VIN+ VD2 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X111 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X112 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 w_109520_3890# X VOUT- w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X114 Vb1 Vb1 a_113080_300# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X115 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X116 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X117 a_118370_3658# V_CMFB_S1 a_109560_2850# sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X118 V_source a_112630_1380# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X119 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 Vb2_Vb3 w_109520_3890# w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X121 Y Vb1 VD2 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X122 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X127 X VD3 VD3 VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X128 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 VD2 a_109560_2850# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X130 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 Vb2_Vb3 Vb2_Vb3 Vb3 Vb2_Vb3 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X132 VD1 VIN- V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X133 w_109520_3890# Vb3 VD4 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X134 VOUT+ V_b_2nd_stage a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X135 a_109560_2850# a_112630_1380# V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X136 V_CMFB_S1 X a_109560_2850# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X137 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 V_err_p V_err_gate w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X139 V_CMFB_S2 X w_109520_3890# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X140 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X141 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X142 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X143 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X146 a_108920_3658# V_tot a_109560_2850# sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X147 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 w_109520_3890# Y VOUT+ w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X149 a_118250_3658# V_tot a_109560_2850# sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X150 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X153 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X155 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X156 VD4 Vb3 w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X157 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 w_109520_3890# Y VOUT+ w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X159 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X160 Y Vb1 VD2 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X161 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X163 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X167 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X168 VD1 VIN- V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X169 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X170 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 Vb3 Vb2 Vb2_Vb3 Vb2_Vb3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X172 V_CMFB_S1 X a_109560_2850# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X173 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 a_109560_2850# a_112630_1380# V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X175 X Vb2 VD3 VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X176 a_109560_2850# a_112630_1380# V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X177 V_err_p V_tot err_amp_mir w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X178 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X179 V_CMFB_S2 X w_109520_3890# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X180 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X184 w_109520_3890# Y VOUT+ w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X185 a_109560_2850# a_109560_2850# VD2 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X186 VD4 Vb3 w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X187 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 VD4 Vb2 Y VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X190 w_109520_3890# X VOUT- w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X191 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 a_118370_3658# V_tot a_109560_2850# sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X193 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X194 w_109520_3890# w_109520_3890# V_err_gate w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X195 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 V_source err_amp_out a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X197 w_109520_3890# Vb3 Vb2_Vb3 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X198 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 Y Vb1 VD2 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X200 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X201 VD3 Vb2 X VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X202 X Vb1 VD1 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X203 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X204 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X205 VOUT+ Y w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X206 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 VD4 Vb3 w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X210 VOUT- X w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X211 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X214 VD1 a_109560_2850# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X215 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 V_CMFB_S1 X a_109560_2850# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X217 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X218 a_109560_2850# a_112630_1380# V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X219 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X220 V_CMFB_S4 Y w_109520_3890# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X221 Vb2_2 Vb2 w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.36 ps=2.2 w=1.8 l=0.2
X222 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 a_109560_2850# a_112630_1380# V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X224 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X225 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X226 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X227 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X228 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 VOUT+ V_b_2nd_stage a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X231 w_109520_3890# Y VOUT+ w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X232 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X233 V_tail_gate VIN- V_p_mir a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X234 V_source VIN+ VD2 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X235 V_CMFB_S4 Y w_109520_3890# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X236 w_109520_3890# Vb3 VD4 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X237 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X238 VD3 Vb2 X VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X239 Y VD4 VD4 VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X240 V_err_mir_p V_err_gate w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X241 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X242 VD3 w_109520_3890# w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X243 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 V_source a_112630_1380# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X245 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 Y Vb1 VD2 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X248 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X249 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 X Vb1 VD1 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X251 X Vb1 VD1 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X252 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 VOUT+ Y w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X255 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 VOUT- X w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X257 V_CMFB_S3 Y a_109560_2850# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X258 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X259 VD3 Vb2 X VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X260 VD3 Vb3 w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X261 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 a_109560_2850# a_112630_1380# V_p_mir a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X263 V_CMFB_S4 Y w_109520_3890# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X264 VD2 Vb1 Y a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X265 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X267 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X268 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 V_CMFB_S2 X w_109520_3890# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X270 w_109520_3890# w_109520_3890# w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=68.76 ps=379 w=1.8 l=0.2
X271 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X272 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X273 w_109520_3890# Vb3 VD4 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X274 V_CMFB_S3 Y a_109560_2850# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X275 V_source VIN+ VD2 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X276 Y Vb2 VD4 VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X277 V_tail_gate a_109560_2850# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X278 a_109560_2850# a_109560_2850# VD1 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X279 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X280 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X281 a_109560_2850# a_109560_2850# Vb1 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X282 w_109520_3890# w_109520_3890# w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X283 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X285 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 w_109520_3890# Y V_CMFB_S4 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X287 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X288 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X289 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X290 VOUT- V_b_2nd_stage a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X291 V_err_mir_p V_err_amp_ref V_err_gate w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X292 err_amp_mir w_109520_3890# w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X293 X Vb2 VD3 VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X294 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X296 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X297 w_109520_3890# X V_CMFB_S2 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X298 VOUT+ a_109560_2850# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X299 Y a_109560_2850# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X300 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 X Vb1 VD1 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X303 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X305 Vb2 Vb2_2 Vb2_2 Vb2_2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X306 w_109520_3890# w_109520_3890# VD4 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X307 Vb1 a_109560_2850# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X308 Y Vb2 VD4 VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X309 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X311 VOUT- X w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X312 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 V_CMFB_S3 Y a_109560_2850# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X314 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 w_109520_3890# w_109520_3890# Vb2_2 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.36 ps=2.2 w=1.8 l=0.2
X318 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 V_CMFB_S1 X a_109560_2850# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X320 a_109560_2850# a_109560_2850# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=50.4 ps=284 w=2.5 l=0.15
X321 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X322 V_CMFB_S4 Y w_109520_3890# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X323 a_109560_2850# V_b_2nd_stage VOUT- a_109560_2850# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X324 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X325 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X326 err_amp_out err_amp_mir a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X327 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 V_source VIN+ VD2 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X329 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 V_source VIN- VD1 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X331 X Vb2 VD3 VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X332 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X333 a_109560_2850# Y V_CMFB_S3 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X334 V_source VIN- VD1 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X335 w_109520_3890# Vb3 VD3 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X336 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X337 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X338 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X339 V_source a_112630_1380# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X340 w_109520_3890# Y V_CMFB_S4 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X341 a_109560_2850# X V_CMFB_S1 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X342 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X343 w_109520_3890# X V_CMFB_S2 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X344 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 X Vb1 VD1 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X346 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X347 a_113080_300# Vb1 Vb1 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X348 a_109560_2850# a_109560_2850# VOUT+ a_109560_2850# sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X349 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X352 X Vb2 VD3 VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X353 VOUT- X w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X354 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X355 w_109520_3890# Vb3 VD3 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X356 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X357 V_CMFB_S3 Y a_109560_2850# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X358 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X360 a_109560_2850# a_112630_1380# V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X361 cap_res_X X a_109560_2850# sky130_fd_pr__res_high_po_1p41 l=1.41
X362 a_109560_2850# a_109560_2850# Y a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X363 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 VD4 Vb3 w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X365 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X366 VD4 Vb2 Y VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X367 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X368 err_amp_mir a_109560_2850# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X369 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X370 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X371 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X374 V_source VIN+ VD2 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X375 V_source VIN- VD1 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X376 a_109560_2850# Y V_CMFB_S3 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X377 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X378 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 V_source a_112630_1380# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X380 a_109560_2850# X V_CMFB_S1 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X381 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 err_amp_out V_err_amp_ref V_err_p w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X383 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X384 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X385 Vb2_2 Vb2 Vb2 Vb2_2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X386 w_109520_3890# X V_CMFB_S2 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X387 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 VD4 Vb2 Y VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X389 w_109520_3890# Vb3 VD3 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X390 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X391 X a_109560_2850# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X392 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X393 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 VD2 VIN+ V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X395 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X396 VOUT- w_109520_3890# w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X397 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X398 VOUT- V_b_2nd_stage a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X399 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 VD4 w_109520_3890# w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X402 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 a_113080_300# Vb1 Vb1 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X404 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X405 VOUT+ Y w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X406 VD2 Vb1 Y a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X407 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X408 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X409 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 a_109040_3658# V_tot a_109560_2850# sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X412 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X413 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 VD3 Vb2 X VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X415 VD3 Vb3 w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X416 V_source VIN- VD1 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X417 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X418 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X419 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X420 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X422 VD4 VD4 Y VD4 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X423 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X424 VOUT- a_118210_146# a_109560_2850# sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X425 a_109560_2850# X V_CMFB_S1 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X426 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 V_source a_112630_1380# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X428 V_source a_112630_1380# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X429 w_109520_3890# V_err_gate V_err_p w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X430 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 w_109520_3890# X V_CMFB_S2 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X432 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 VD3 VD3 X VD3 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X436 VOUT+ Y w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X437 VD3 Vb3 w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X438 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X442 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X443 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X444 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 a_109560_2850# a_109560_2850# V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X446 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X447 w_109520_3890# Vb3 VD4 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X448 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X449 VD2 Vb1 Y a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X450 Y Vb2 VD4 VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X451 VD3 Vb3 w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X452 VOUT+ w_109520_3890# w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X453 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X454 a_109560_2850# V_b_2nd_stage VOUT+ a_109560_2850# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X455 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 a_109560_2850# a_109560_2850# X a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X457 w_109520_3890# w_109520_3890# VOUT+ w_109520_3890# sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X458 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 w_109520_3890# w_109520_3890# VOUT- w_109520_3890# sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X461 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 V_source VIN- VD1 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X464 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X465 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X466 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X467 a_109560_2850# X V_CMFB_S1 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X468 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X469 Vb2_2 Vb2_2 Vb2_2 Vb2_2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=4.92 ps=27.8 w=3.5 l=0.2
X470 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X471 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 V_source a_112630_1380# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X473 Y Vb2 VD4 VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X474 w_109520_3890# a_109560_2850# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X475 VD3 Vb3 w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X476 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X477 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X478 V_b_2nd_stage a_109200_146# a_109560_2850# sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X479 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X480 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X481 VOUT+ Y w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X482 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X484 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X485 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X486 a_109560_2850# a_109560_2850# V_tail_gate a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X487 VD2 VIN+ V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X488 w_109520_3890# Y V_CMFB_S4 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X489 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 Y Vb2 VD4 VD4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X491 VOUT- X w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X492 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X494 V_err_gate V_tot V_err_mir_p w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X495 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X496 a_109560_2850# a_112630_1380# V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X497 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 a_109040_3658# V_CMFB_S3 a_109560_2850# sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X499 VD2 Vb1 Y a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X500 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X501 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X502 X Vb2 VD3 VD3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X503 VD1 Vb1 X a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X504 VD1 Vb1 X a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X505 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X506 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X507 w_109520_3890# Vb3 VD3 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X508 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X509 w_109520_3890# Y VOUT+ w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X510 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 VOUT- cap_res_X sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X512 a_109560_2850# a_109560_2850# VOUT- a_109560_2850# sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X513 w_109520_3890# X VOUT- w_109520_3890# sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X514 a_109560_2850# V_b_2nd_stage VOUT+ a_109560_2850# sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X515 a_109560_2850# w_109520_3890# w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X516 V_source a_112630_1380# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X517 w_109520_3890# Y V_CMFB_S4 a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X518 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X519 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X520 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X521 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X522 a_109560_2850# Y V_CMFB_S3 w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X523 V_b_2nd_stage a_118210_146# a_109560_2850# sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X524 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 V_p_mir VIN+ V_tail_gate a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X526 VD2 VIN+ V_source a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X527 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 w_109520_3890# a_109560_2850# a_109560_2850# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X529 VD4 Vb3 w_109520_3890# w_109520_3890# sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X530 VOUT+ cap_res_Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X531 a_109560_2850# a_109560_2850# w_109520_3890# a_109560_2850# sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
.ends

