* NGSPICE file created from pfd_3.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

**.subckt pfd_3 F_REF F_VCO QA QB VDDA GNDA
Xsky130_fd_sc_hd__inv_1_4 sky130_fd_sc_hd__inv_1_4/A GNDA VSUBS sky130_fd_sc_hd__inv_1_4/VPB
+ VDDA sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__nor2_1_1 sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__nor2_1_2/A
+ GNDA VSUBS sky130_fd_sc_hd__inv_1_4/VPB VDDA QB sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_0 F_VCO QB GNDA VSUBS sky130_fd_sc_hd__inv_1_4/VPB VDDA sky130_fd_sc_hd__nor2_1_2/A
+ sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_2 sky130_fd_sc_hd__nor2_1_2/A sky130_fd_sc_hd__nor2_1_3/Y
+ GNDA VSUBS sky130_fd_sc_hd__inv_1_4/VPB VDDA sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_3 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__nor2_1_3/B
+ GNDA VSUBS sky130_fd_sc_hd__inv_1_4/VPB VDDA sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_4 F_REF QA GNDA VSUBS sky130_fd_sc_hd__inv_1_4/VPB VDDA sky130_fd_sc_hd__nor2_1_7/B
+ sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_5 sky130_fd_sc_hd__nor2_1_7/B sky130_fd_sc_hd__nor2_1_6/Y
+ GNDA VSUBS sky130_fd_sc_hd__inv_1_4/VPB VDDA sky130_fd_sc_hd__nor2_1_7/A sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_6 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__nor2_1_7/A
+ GNDA VSUBS sky130_fd_sc_hd__inv_1_4/VPB VDDA sky130_fd_sc_hd__nor2_1_6/Y sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_7 sky130_fd_sc_hd__nor2_1_7/A sky130_fd_sc_hd__nor2_1_7/B
+ GNDA VSUBS sky130_fd_sc_hd__inv_1_4/VPB VDDA QA sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nand2_1_1 QA QB GNDA VSUBS sky130_fd_sc_hd__inv_1_4/VPB VDDA sky130_fd_sc_hd__inv_1_2/A
+ sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__inv_1_0 sky130_fd_sc_hd__inv_1_4/Y GNDA VSUBS sky130_fd_sc_hd__inv_1_4/VPB
+ VDDA sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_1 sky130_fd_sc_hd__inv_1_1/A GNDA VSUBS sky130_fd_sc_hd__inv_1_4/VPB
+ VDDA sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_2 sky130_fd_sc_hd__inv_1_2/A GNDA VSUBS sky130_fd_sc_hd__inv_1_4/VPB
+ VDDA sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_3 sky130_fd_sc_hd__inv_1_3/A GNDA VSUBS sky130_fd_sc_hd__inv_1_4/VPB
+ VDDA sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1
**.ends

