** sch_path: /foss/designs/my_design/projects/opamp/xschem_ngspice/tb_bgr_opamp_dummy_magic.sch
**.subckt tb_bgr_opamp_dummy_magic
VDD VDD GND pwl(0 0 1us 0 2us 1.8)
V2 VIN- GND sin(1.24 -0.001 100k)
V1 VIN+ GND sin(1.24 0.001 100k)
XC1 VOUT+ GND sky130_fd_pr__cap_mim_m3_1 W=23 L=23 MF=1 m=1
XC2 VOUT- GND sky130_fd_pr__cap_mim_m3_1 W=23 L=23 MF=1 m=1
x2 VDD GND VOUT+ VOUT- VIN+ VIN- bgr_opamp_dummy_magic
**** begin user architecture code
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt




.include /foss/designs/my_design/projects/opamp/xschem_ngspice/bgr_opamp_dummy_magic.spice
* .include /foss/designs/my_design/projects/opamp/xschem_ngspice/two_stage_opamp_dummy_magic.spice
* .include /foss/designs/my_design/projects/opamp/xschem_ngspice/ref_volt_cur_gen_dummy_magic.spice


.option method=gear
.option wnflag=1
.option savecurrents

.save
+v(vout+)
+v(vout-)
+v(vin+)
+v(vin-)
+v(x2.two_stage_opamp_dummy_magic_0.v_cmfb_s1.t0)
+v(x2.two_stage_opamp_dummy_magic_0.v_cmfb_s2.t0)
+v(x2.two_stage_opamp_dummy_magic_0.v_cmfb_s3.t0)
+v(x2.two_stage_opamp_dummy_magic_0.v_cmfb_s4.t0)
+v(x2.two_stage_opamp_dummy_magic_0.x.t0)
+v(x2.two_stage_opamp_dummy_magic_0.y.t0)
+v(x2.two_stage_opamp_dummy_magic_0.v_tot.t0)
+v(x2.two_stage_opamp_dummy_magic_0.v_err_amp_ref.t0)


* .ic v(v_top) = 1.8

.control

  * let runs=3
  * let run=1

  * dowhile run <= runs
    * save v(vout+) v(vout-) v(vin+) v(vin-) v(v_err_amp_ref) v(x2.x) v(x2.y) v(x2.vb1) v(x2.vb2) v(x2.vb3) v(x2.v_tot)
    save all
    remzerovec
    set appendwrite
    * dc temp -40 120 10 VDD 0 4.0 0.2
    * dc VDD 0 2.0 0.02 temp -40 120 40
    * dc V5 0 0.01 0.0001
    tran 2n 30u
    * tran 10n 150u
    * tran 1p 3n
    * tran 0.1ns 30us
    * ac dec 40 1 10T
    * write tb_bgr_opamp_dummy_magic.raw
    * write tb_bgr_opamp_dummy_magic_2.raw
    * write tb_bgr_opamp_dummy_magic_3.raw
    * write tb_bgr_opamp_dummy_magic_4.raw
    * write tb_bgr_opamp_dummy_magic_5.raw
    * write tb_bgr_opamp_dummy_magic_6.raw
    * write tb_bgr_opamp_dummy_magic_7.raw
    * write tb_bgr_opamp_dummy_magic_8.raw
    * write tb_bgr_opamp_dummy_magic_9.raw
    * write tb_bgr_opamp_dummy_magic_10.raw
    * write tb_bgr_opamp_dummy_magic_11.raw
    * write tb_bgr_opamp_dummy_magic_12.raw
    * write tb_bgr_opamp_dummy_magic_13.raw
    * write tb_bgr_opamp_dummy_magic_14.raw
    * write tb_bgr_opamp_dummy_magic_15.raw
    * write tb_bgr_opamp_dummy_magic_16.raw
    * write tb_bgr_opamp_dummy_magic_17.raw
    * write tb_bgr_opamp_dummy_magic_18.raw
    * write tb_bgr_opamp_dummy_magic_19.raw
    * write tb_bgr_opamp_dummy_magic_20.raw
    * write tb_bgr_opamp_dummy_magic_21.raw
    * write tb_bgr_opamp_dummy_magic_22.raw
    * write tb_bgr_opamp_dummy_magic_23.raw
    * write tb_bgr_opamp_dummy_magic_24.raw
    * write tb_bgr_opamp_dummy_magic_25.raw
    * write tb_bgr_opamp_dummy_magic_26.raw
    write tb_bgr_opamp_dummy_magic_27.raw
    * write tb_bgr_opamp_dummy_magic_mc.raw
    * write tb_bgr_opamp_dummy_magic_tt_mm.raw
    * write tb_bgr_opamp_dummy_magic_AC.raw
    * reset
    * let run = run + 1
  * end
.endc



**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
