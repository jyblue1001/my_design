* PEX produced on Mon Feb 17 02:31:51 PM CET 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from charge_pump_cell_4.ext - technology: sky130A

.subckt charge_pump_cell_4 VDDA GNDA x vout UP_b DOWN I_IN UP_input DOWN_input opamp_out
X0 UP_input.t0 UP_b.t0 sky130_fd_pr__cap_mim_m3_1 l=6.3 w=8.75
X1 GNDA.t3 I_IN.t0 I_IN.t1 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=2 pd=9 as=2 ps=9 w=4 l=0.6
X2 VDDA.t3 UP_input.t1 vout.t0 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=4 pd=17 as=4 ps=17 w=8 l=0.6
X3 GNDA.t5 DOWN_input.t0 vout.t1 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=2 pd=9 as=2 ps=9 w=4 l=0.6
X4 x.t0 opamp_out.t0 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=3.6 pd=16.9 as=4 ps=17 w=8 l=0.6
X5 x.t1 I_IN.t2 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=2 pd=9 as=2 ps=9 w=4 l=0.6
X6 DOWN_input.t1 DOWN.t0 sky130_fd_pr__cap_mim_m3_1 l=2.6 w=3.1
R0 UP_input UP_input.t1 333.384
R1 UP_input UP_input.t0 326.658
R2 UP_b UP_b.t0 10.2459
R3 I_IN.t0 I_IN.t2 879.65
R4 I_IN.n0 I_IN.t0 388.983
R5 I_IN I_IN.n0 80.0005
R6 I_IN.n0 I_IN.t1 79.5157
R7 GNDA.t2 GNDA.n39 34765
R8 GNDA.t4 GNDA.t0 972.093
R9 GNDA.n38 GNDA.n37 669.307
R10 GNDA.n16 GNDA.n3 669.307
R11 GNDA.n50 GNDA.n1 669.307
R12 GNDA.n36 GNDA.n22 585
R13 GNDA.n34 GNDA.n21 585
R14 GNDA.n39 GNDA.n21 585
R15 GNDA.n33 GNDA.n32 585
R16 GNDA.n30 GNDA.n29 585
R17 GNDA.n28 GNDA.n27 585
R18 GNDA.n25 GNDA.n24 585
R19 GNDA.n20 GNDA.n0 585
R20 GNDA.n39 GNDA.n20 585
R21 GNDA.n15 GNDA.n14 585
R22 GNDA.n13 GNDA.n11 585
R23 GNDA.n43 GNDA.n42 585
R24 GNDA.n12 GNDA.n9 585
R25 GNDA.n47 GNDA.n8 585
R26 GNDA.n7 GNDA.n6 585
R27 GNDA.n39 GNDA.t4 537.21
R28 GNDA.n40 GNDA.t0 537.21
R29 GNDA.n40 GNDA.t2 537.21
R30 GNDA.n39 GNDA.n38 250.349
R31 GNDA.n39 GNDA.n18 250.349
R32 GNDA.n39 GNDA.n19 250.349
R33 GNDA.n41 GNDA.n40 250.349
R34 GNDA.n40 GNDA.n17 250.349
R35 GNDA.n40 GNDA.n1 250.349
R36 GNDA.n40 GNDA.n16 250.349
R37 GNDA.n22 GNDA.n21 197
R38 GNDA.n32 GNDA.n21 197
R39 GNDA.n29 GNDA.n28 197
R40 GNDA.n24 GNDA.n20 197
R41 GNDA.n15 GNDA.n13 197
R42 GNDA.n42 GNDA.n12 197
R43 GNDA.n8 GNDA.n7 197
R44 GNDA.n37 GNDA.n23 185
R45 GNDA.n23 GNDA.n0 185
R46 GNDA.n50 GNDA.n49 185
R47 GNDA.n49 GNDA.n3 185
R48 GNDA.n45 GNDA.n44 91.3721
R49 GNDA.n46 GNDA.n45 91.3721
R50 GNDA.n45 GNDA.n2 91.3721
R51 GNDA.n45 GNDA.n10 91.3721
R52 GNDA.n49 GNDA.n4 91.3721
R53 GNDA.n49 GNDA.n5 91.3721
R54 GNDA.n49 GNDA.n48 91.3721
R55 GNDA.n35 GNDA.n23 90.7567
R56 GNDA.n31 GNDA.n23 90.7567
R57 GNDA.n26 GNDA.n23 90.7567
R58 GNDA.n32 GNDA.n18 84.306
R59 GNDA.n28 GNDA.n19 84.306
R60 GNDA.n38 GNDA.n22 84.306
R61 GNDA.n29 GNDA.n18 84.306
R62 GNDA.n24 GNDA.n19 84.306
R63 GNDA.n41 GNDA.n13 84.306
R64 GNDA.n17 GNDA.n12 84.306
R65 GNDA.n7 GNDA.n1 84.306
R66 GNDA.n16 GNDA.n15 84.306
R67 GNDA.n42 GNDA.n41 84.306
R68 GNDA.n17 GNDA.n8 84.306
R69 GNDA.n51 GNDA.n0 37.9505
R70 GNDA.n51 GNDA.n50 34.4485
R71 GNDA.n49 GNDA.t3 7.5005
R72 GNDA.n23 GNDA.t5 7.5005
R73 GNDA.n45 GNDA.t1 7.5005
R74 GNDA.n37 GNDA.n36 7.11161
R75 GNDA.n34 GNDA.n33 7.11161
R76 GNDA.n30 GNDA.n27 7.11161
R77 GNDA.n25 GNDA.n0 7.11161
R78 GNDA.n36 GNDA.n35 3.48951
R79 GNDA.n33 GNDA.n31 3.48951
R80 GNDA.n27 GNDA.n26 3.48951
R81 GNDA.n35 GNDA.n34 3.48951
R82 GNDA.n31 GNDA.n30 3.48951
R83 GNDA.n26 GNDA.n25 3.48951
R84 GNDA.n10 GNDA.n3 2.25882
R85 GNDA.n11 GNDA.n4 2.25882
R86 GNDA.n44 GNDA.n11 2.25882
R87 GNDA.n9 GNDA.n5 2.25882
R88 GNDA.n46 GNDA.n9 2.25882
R89 GNDA.n48 GNDA.n6 2.25882
R90 GNDA.n6 GNDA.n2 2.25882
R91 GNDA.n14 GNDA.n10 2.25882
R92 GNDA.n44 GNDA.n43 2.25882
R93 GNDA.n47 GNDA.n46 2.25882
R94 GNDA.n50 GNDA.n2 2.25882
R95 GNDA.n14 GNDA.n4 2.25882
R96 GNDA.n43 GNDA.n5 2.25882
R97 GNDA.n48 GNDA.n47 2.25882
R98 GNDA GNDA.n51 0.75146
R99 vout vout.t0 150.468
R100 vout vout.t1 95.5157
R101 VDDA.n43 VDDA.n0 585
R102 VDDA.n43 VDDA.n42 585
R103 VDDA.n89 VDDA.n88 290.733
R104 VDDA.n88 VDDA.n52 290.733
R105 VDDA.n88 VDDA.n53 290.733
R106 VDDA.n88 VDDA.n54 290.733
R107 VDDA.n88 VDDA.n55 290.733
R108 VDDA.n88 VDDA.n56 290.733
R109 VDDA.n88 VDDA.n87 290.733
R110 VDDA.n88 VDDA.n1 290.733
R111 VDDA.n44 VDDA.n43 290.733
R112 VDDA.n43 VDDA.n14 290.733
R113 VDDA.n43 VDDA.n19 290.733
R114 VDDA.n43 VDDA.n24 290.733
R115 VDDA.n43 VDDA.n29 290.733
R116 VDDA.n43 VDDA.n34 290.733
R117 VDDA.n43 VDDA.n39 290.733
R118 VDDA.n87 VDDA.n86 233.841
R119 VDDA.n94 VDDA.n93 230.308
R120 VDDA.t0 VDDA.t2 202.81
R121 VDDA.n92 VDDA.n91 185
R122 VDDA.n90 VDDA.n50 185
R123 VDDA.n60 VDDA.n51 185
R124 VDDA.n62 VDDA.n61 185
R125 VDDA.n65 VDDA.n64 185
R126 VDDA.n67 VDDA.n66 185
R127 VDDA.n70 VDDA.n69 185
R128 VDDA.n72 VDDA.n71 185
R129 VDDA.n75 VDDA.n74 185
R130 VDDA.n77 VDDA.n76 185
R131 VDDA.n80 VDDA.n79 185
R132 VDDA.n82 VDDA.n81 185
R133 VDDA.n84 VDDA.n58 185
R134 VDDA.n85 VDDA.n57 185
R135 VDDA.n47 VDDA.n0 185
R136 VDDA.n48 VDDA.n47 185
R137 VDDA.n46 VDDA.n45 185
R138 VDDA.n11 VDDA.n10 185
R139 VDDA.n13 VDDA.n12 185
R140 VDDA.n16 VDDA.n15 185
R141 VDDA.n18 VDDA.n17 185
R142 VDDA.n21 VDDA.n20 185
R143 VDDA.n23 VDDA.n22 185
R144 VDDA.n26 VDDA.n25 185
R145 VDDA.n28 VDDA.n27 185
R146 VDDA.n31 VDDA.n30 185
R147 VDDA.n33 VDDA.n32 185
R148 VDDA.n36 VDDA.n35 185
R149 VDDA.n38 VDDA.n37 185
R150 VDDA.n41 VDDA.n40 185
R151 VDDA.n42 VDDA.n9 185
R152 VDDA.n48 VDDA.n9 185
R153 VDDA.n92 VDDA.n50 120.001
R154 VDDA.n62 VDDA.n60 120.001
R155 VDDA.n67 VDDA.n64 120.001
R156 VDDA.n72 VDDA.n69 120.001
R157 VDDA.n77 VDDA.n74 120.001
R158 VDDA.n82 VDDA.n79 120.001
R159 VDDA.n85 VDDA.n84 120.001
R160 VDDA.n47 VDDA.n46 120.001
R161 VDDA.n12 VDDA.n11 120.001
R162 VDDA.n17 VDDA.n16 120.001
R163 VDDA.n22 VDDA.n21 120.001
R164 VDDA.n27 VDDA.n26 120.001
R165 VDDA.n32 VDDA.n31 120.001
R166 VDDA.n37 VDDA.n36 120.001
R167 VDDA.n40 VDDA.n9 120.001
R168 VDDA.t2 VDDA.n48 112.079
R169 VDDA.n49 VDDA.t0 112.079
R170 VDDA.n93 VDDA.n49 69.8479
R171 VDDA.n59 VDDA.n49 69.8479
R172 VDDA.n63 VDDA.n49 69.8479
R173 VDDA.n68 VDDA.n49 69.8479
R174 VDDA.n73 VDDA.n49 69.8479
R175 VDDA.n78 VDDA.n49 69.8479
R176 VDDA.n83 VDDA.n49 69.8479
R177 VDDA.n86 VDDA.n49 69.8479
R178 VDDA.n48 VDDA.n2 69.8479
R179 VDDA.n48 VDDA.n3 69.8479
R180 VDDA.n48 VDDA.n4 69.8479
R181 VDDA.n48 VDDA.n5 69.8479
R182 VDDA.n48 VDDA.n6 69.8479
R183 VDDA.n48 VDDA.n7 69.8479
R184 VDDA.n48 VDDA.n8 69.8479
R185 VDDA.n93 VDDA.n92 45.3071
R186 VDDA.n59 VDDA.n50 45.3071
R187 VDDA.n63 VDDA.n62 45.3071
R188 VDDA.n68 VDDA.n67 45.3071
R189 VDDA.n73 VDDA.n72 45.3071
R190 VDDA.n78 VDDA.n77 45.3071
R191 VDDA.n83 VDDA.n82 45.3071
R192 VDDA.n86 VDDA.n85 45.3071
R193 VDDA.n60 VDDA.n59 45.3071
R194 VDDA.n64 VDDA.n63 45.3071
R195 VDDA.n69 VDDA.n68 45.3071
R196 VDDA.n74 VDDA.n73 45.3071
R197 VDDA.n79 VDDA.n78 45.3071
R198 VDDA.n84 VDDA.n83 45.3071
R199 VDDA.n46 VDDA.n2 45.3071
R200 VDDA.n12 VDDA.n3 45.3071
R201 VDDA.n17 VDDA.n4 45.3071
R202 VDDA.n22 VDDA.n5 45.3071
R203 VDDA.n27 VDDA.n6 45.3071
R204 VDDA.n32 VDDA.n7 45.3071
R205 VDDA.n37 VDDA.n8 45.3071
R206 VDDA.n11 VDDA.n2 45.3071
R207 VDDA.n16 VDDA.n3 45.3071
R208 VDDA.n21 VDDA.n4 45.3071
R209 VDDA.n26 VDDA.n5 45.3071
R210 VDDA.n31 VDDA.n6 45.3071
R211 VDDA.n36 VDDA.n7 45.3071
R212 VDDA.n40 VDDA.n8 45.3071
R213 VDDA.n95 VDDA.n0 41.4847
R214 VDDA.n95 VDDA.n94 38.3476
R215 VDDA.n91 VDDA.n90 7.11161
R216 VDDA.n61 VDDA.n51 7.11161
R217 VDDA.n66 VDDA.n65 7.11161
R218 VDDA.n71 VDDA.n70 7.11161
R219 VDDA.n76 VDDA.n75 7.11161
R220 VDDA.n81 VDDA.n80 7.11161
R221 VDDA.n58 VDDA.n57 7.11161
R222 VDDA.n45 VDDA.n0 7.11161
R223 VDDA.n13 VDDA.n10 7.11161
R224 VDDA.n18 VDDA.n15 7.11161
R225 VDDA.n23 VDDA.n20 7.11161
R226 VDDA.n28 VDDA.n25 7.11161
R227 VDDA.n33 VDDA.n30 7.11161
R228 VDDA.n38 VDDA.n35 7.11161
R229 VDDA.n42 VDDA.n41 7.11161
R230 VDDA.n43 VDDA.t3 6.15675
R231 VDDA.n88 VDDA.t1 6.15675
R232 VDDA.n94 VDDA.n1 3.53508
R233 VDDA.n90 VDDA.n89 3.53508
R234 VDDA.n61 VDDA.n52 3.53508
R235 VDDA.n66 VDDA.n53 3.53508
R236 VDDA.n71 VDDA.n54 3.53508
R237 VDDA.n76 VDDA.n55 3.53508
R238 VDDA.n81 VDDA.n56 3.53508
R239 VDDA.n87 VDDA.n57 3.53508
R240 VDDA.n91 VDDA.n1 3.53508
R241 VDDA.n89 VDDA.n51 3.53508
R242 VDDA.n65 VDDA.n52 3.53508
R243 VDDA.n70 VDDA.n53 3.53508
R244 VDDA.n75 VDDA.n54 3.53508
R245 VDDA.n80 VDDA.n55 3.53508
R246 VDDA.n58 VDDA.n56 3.53508
R247 VDDA.n45 VDDA.n44 3.53508
R248 VDDA.n14 VDDA.n13 3.53508
R249 VDDA.n19 VDDA.n18 3.53508
R250 VDDA.n24 VDDA.n23 3.53508
R251 VDDA.n29 VDDA.n28 3.53508
R252 VDDA.n34 VDDA.n33 3.53508
R253 VDDA.n39 VDDA.n38 3.53508
R254 VDDA.n44 VDDA.n10 3.53508
R255 VDDA.n15 VDDA.n14 3.53508
R256 VDDA.n20 VDDA.n19 3.53508
R257 VDDA.n25 VDDA.n24 3.53508
R258 VDDA.n30 VDDA.n29 3.53508
R259 VDDA.n35 VDDA.n34 3.53508
R260 VDDA.n41 VDDA.n39 3.53508
R261 VDDA VDDA.n95 0.939041
R262 DOWN_input.t0 DOWN_input.n0 494.05
R263 DOWN_input DOWN_input.t1 326.658
R264 DOWN_input DOWN_input.t0 172.718
R265 opamp_out opamp_out.t0 369.534
R266 x x.t0 147.425
R267 x x.t1 109.915
R268 DOWN DOWN.t0 10.2215
C0 DOWN I_IN 0.022543f
C1 opamp_out VDDA 0.323172f
C2 UP_b opamp_out 0.022669f
C3 UP_b DOWN 0.039793f
C4 VDDA UP_input 0.484285f
C5 DOWN_input vout 0.261437f
C6 UP_b UP_input 0.222182f
C7 x vout 0.715241f
C8 DOWN DOWN_input 0.202326f
C9 opamp_out x 0.218577f
C10 DOWN_input UP_input 0.102282f
C11 vout UP_input 0.38509f
C12 UP_b VDDA 0.557519f
C13 I_IN DOWN_input 0.013941f
C14 I_IN x 0.119536f
C15 VDDA vout 0.356465f
C16 UP_b vout 0.012981f
C17 VDDA x 0.359776f
C18 DOWN GNDA 1.91849f
C19 UP_b GNDA 2.91095f
C20 DOWN_input GNDA 1.01941f
C21 I_IN GNDA 1.67577f
C22 vout GNDA 0.410407f
C23 x GNDA 0.316274f
C24 UP_input GNDA 0.638409f
C25 opamp_out GNDA 0.117526f
C26 VDDA GNDA 6.29776f
.ends

