magic
tech sky130A
timestamp 1749008454
<< nwell >>
rect 2545 1880 5285 2950
<< pwell >>
rect -45 1685 130 1725
rect 3165 1615 3805 1665
rect 4205 1615 4845 1665
rect 11030 1565 11730 1715
rect 11770 1565 12030 1715
rect 12070 1565 12770 1715
rect 2835 1205 3955 1455
rect 4055 1205 5175 1455
rect 2945 975 5065 1075
rect 11205 1025 12620 1275
rect 2995 780 5015 880
<< nmos >>
rect 3205 1615 3225 1665
rect 3265 1615 3285 1665
rect 3325 1615 3345 1665
rect 3385 1615 3405 1665
rect 3445 1615 3465 1665
rect 3505 1615 3525 1665
rect 3565 1615 3585 1665
rect 3625 1615 3645 1665
rect 3685 1615 3705 1665
rect 3745 1615 3765 1665
rect 4245 1615 4265 1665
rect 4305 1615 4325 1665
rect 4365 1615 4385 1665
rect 4425 1615 4445 1665
rect 4485 1615 4505 1665
rect 4545 1615 4565 1665
rect 4605 1615 4625 1665
rect 4665 1615 4685 1665
rect 4725 1615 4745 1665
rect 4785 1615 4805 1665
rect 11070 1565 11085 1715
rect 11125 1565 11140 1715
rect 11180 1565 11195 1715
rect 11235 1565 11250 1715
rect 11290 1565 11305 1715
rect 11345 1565 11360 1715
rect 11400 1565 11415 1715
rect 11455 1565 11470 1715
rect 11510 1565 11525 1715
rect 11565 1565 11580 1715
rect 11620 1565 11635 1715
rect 11675 1565 11690 1715
rect 11810 1565 11825 1715
rect 11865 1565 11880 1715
rect 11920 1565 11935 1715
rect 11975 1565 11990 1715
rect 12110 1565 12125 1715
rect 12165 1565 12180 1715
rect 12220 1565 12235 1715
rect 12275 1565 12290 1715
rect 12330 1565 12345 1715
rect 12385 1565 12400 1715
rect 12440 1565 12455 1715
rect 12495 1565 12510 1715
rect 12550 1565 12565 1715
rect 12605 1565 12620 1715
rect 12660 1565 12675 1715
rect 12715 1565 12730 1715
rect 2875 1205 3375 1455
rect 3415 1205 3915 1455
rect 4095 1205 4595 1455
rect 4635 1205 5135 1455
rect 2985 975 3985 1075
rect 4025 975 5025 1075
rect 11245 1025 11260 1275
rect 11300 1025 11315 1275
rect 11355 1025 11370 1275
rect 11410 1025 11425 1275
rect 11465 1025 11480 1275
rect 11520 1025 11535 1275
rect 11575 1025 11590 1275
rect 11630 1025 11645 1275
rect 11685 1025 11700 1275
rect 11740 1025 11755 1275
rect 11795 1025 11810 1275
rect 11850 1025 11865 1275
rect 11905 1025 11920 1275
rect 11960 1025 11975 1275
rect 12015 1025 12030 1275
rect 12070 1025 12085 1275
rect 12125 1025 12140 1275
rect 12180 1025 12195 1275
rect 12235 1025 12250 1275
rect 12290 1025 12305 1275
rect 12345 1025 12360 1275
rect 12400 1025 12415 1275
rect 12455 1025 12470 1275
rect 12510 1025 12525 1275
rect 12565 1025 12580 1275
rect 3035 780 3085 880
rect 3125 780 3175 880
rect 3215 780 3265 880
rect 3305 780 3355 880
rect 3395 780 3445 880
rect 3485 780 3535 880
rect 3575 780 3625 880
rect 3665 780 3715 880
rect 3755 780 3805 880
rect 3845 780 3895 880
rect 3935 780 3985 880
rect 4025 780 4075 880
rect 4115 780 4165 880
rect 4205 780 4255 880
rect 4295 780 4345 880
rect 4385 780 4435 880
rect 4475 780 4525 880
rect 4565 780 4615 880
rect 4655 780 4705 880
rect 4745 780 4795 880
rect 4835 780 4885 880
rect 4925 780 4975 880
<< pmos >>
rect 3035 2830 3085 2930
rect 3125 2830 3175 2930
rect 3215 2830 3265 2930
rect 3305 2830 3355 2930
rect 3395 2830 3445 2930
rect 3485 2830 3535 2930
rect 3575 2830 3625 2930
rect 3665 2830 3715 2930
rect 3755 2830 3805 2930
rect 3845 2830 3895 2930
rect 3935 2830 3985 2930
rect 4025 2830 4075 2930
rect 4115 2830 4165 2930
rect 4205 2830 4255 2930
rect 4295 2830 4345 2930
rect 4385 2830 4435 2930
rect 4475 2830 4525 2930
rect 4565 2830 4615 2930
rect 4655 2830 4705 2930
rect 4745 2830 4795 2930
rect 4835 2830 4885 2930
rect 4925 2830 4975 2930
rect 3215 2400 3265 2700
rect 3305 2400 3355 2700
rect 3395 2400 3445 2700
rect 3485 2400 3535 2700
rect 3575 2400 3625 2700
rect 3665 2400 3715 2700
rect 3755 2400 3805 2700
rect 3845 2400 3895 2700
rect 3935 2400 3985 2700
rect 4025 2400 4075 2700
rect 4115 2400 4165 2700
rect 4205 2400 4255 2700
rect 4295 2400 4345 2700
rect 4385 2400 4435 2700
rect 4475 2400 4525 2700
rect 4565 2400 4615 2700
rect 4655 2400 4705 2700
rect 4745 2400 4795 2700
rect 2605 1900 2620 2000
rect 2660 1900 2675 2000
rect 2785 1900 2805 2000
rect 2845 1900 2865 2000
rect 2905 1900 2925 2000
rect 2965 1900 2985 2000
rect 3025 1900 3045 2000
rect 3085 1900 3105 2000
rect 3145 1900 3165 2000
rect 3205 1900 3225 2000
rect 3265 1900 3285 2000
rect 3325 1900 3345 2000
rect 3385 1900 3405 2000
rect 3445 1900 3465 2000
rect 3505 1900 3525 2000
rect 3565 1900 3585 2000
rect 3625 1900 3645 2000
rect 3685 1900 3705 2000
rect 3745 1900 3765 2000
rect 3805 1900 3825 2000
rect 3865 1900 3885 2000
rect 3925 1900 3945 2000
rect 4065 1900 4085 2000
rect 4125 1900 4145 2000
rect 4185 1900 4205 2000
rect 4245 1900 4265 2000
rect 4305 1900 4325 2000
rect 4365 1900 4385 2000
rect 4425 1900 4445 2000
rect 4485 1900 4505 2000
rect 4545 1900 4565 2000
rect 4605 1900 4625 2000
rect 4665 1900 4685 2000
rect 4725 1900 4745 2000
rect 4785 1900 4805 2000
rect 4845 1900 4865 2000
rect 4905 1900 4925 2000
rect 4965 1900 4985 2000
rect 5025 1900 5045 2000
rect 5085 1900 5105 2000
rect 5145 1900 5165 2000
rect 5205 1900 5225 2000
<< ndiff >>
rect 11030 1700 11070 1715
rect 11030 1680 11040 1700
rect 11060 1680 11070 1700
rect 3165 1650 3205 1665
rect 3165 1630 3175 1650
rect 3195 1630 3205 1650
rect 3165 1615 3205 1630
rect 3225 1650 3265 1665
rect 3225 1630 3235 1650
rect 3255 1630 3265 1650
rect 3225 1615 3265 1630
rect 3285 1650 3325 1665
rect 3285 1630 3295 1650
rect 3315 1630 3325 1650
rect 3285 1615 3325 1630
rect 3345 1650 3385 1665
rect 3345 1630 3355 1650
rect 3375 1630 3385 1650
rect 3345 1615 3385 1630
rect 3405 1650 3445 1665
rect 3405 1630 3415 1650
rect 3435 1630 3445 1650
rect 3405 1615 3445 1630
rect 3465 1650 3505 1665
rect 3465 1630 3475 1650
rect 3495 1630 3505 1650
rect 3465 1615 3505 1630
rect 3525 1650 3565 1665
rect 3525 1630 3535 1650
rect 3555 1630 3565 1650
rect 3525 1615 3565 1630
rect 3585 1650 3625 1665
rect 3585 1630 3595 1650
rect 3615 1630 3625 1650
rect 3585 1615 3625 1630
rect 3645 1650 3685 1665
rect 3645 1630 3655 1650
rect 3675 1630 3685 1650
rect 3645 1615 3685 1630
rect 3705 1650 3745 1665
rect 3705 1630 3715 1650
rect 3735 1630 3745 1650
rect 3705 1615 3745 1630
rect 3765 1650 3805 1665
rect 3765 1630 3775 1650
rect 3795 1630 3805 1650
rect 3765 1615 3805 1630
rect 4205 1650 4245 1665
rect 4205 1630 4215 1650
rect 4235 1630 4245 1650
rect 4205 1615 4245 1630
rect 4265 1650 4305 1665
rect 4265 1630 4275 1650
rect 4295 1630 4305 1650
rect 4265 1615 4305 1630
rect 4325 1650 4365 1665
rect 4325 1630 4335 1650
rect 4355 1630 4365 1650
rect 4325 1615 4365 1630
rect 4385 1650 4425 1665
rect 4385 1630 4395 1650
rect 4415 1630 4425 1650
rect 4385 1615 4425 1630
rect 4445 1650 4485 1665
rect 4445 1630 4455 1650
rect 4475 1630 4485 1650
rect 4445 1615 4485 1630
rect 4505 1650 4545 1665
rect 4505 1630 4515 1650
rect 4535 1630 4545 1650
rect 4505 1615 4545 1630
rect 4565 1650 4605 1665
rect 4565 1630 4575 1650
rect 4595 1630 4605 1650
rect 4565 1615 4605 1630
rect 4625 1650 4665 1665
rect 4625 1630 4635 1650
rect 4655 1630 4665 1650
rect 4625 1615 4665 1630
rect 4685 1650 4725 1665
rect 4685 1630 4695 1650
rect 4715 1630 4725 1650
rect 4685 1615 4725 1630
rect 4745 1650 4785 1665
rect 4745 1630 4755 1650
rect 4775 1630 4785 1650
rect 4745 1615 4785 1630
rect 4805 1650 4845 1665
rect 4805 1630 4815 1650
rect 4835 1630 4845 1650
rect 4805 1615 4845 1630
rect 11030 1650 11070 1680
rect 11030 1630 11040 1650
rect 11060 1630 11070 1650
rect 11030 1600 11070 1630
rect 11030 1580 11040 1600
rect 11060 1580 11070 1600
rect 11030 1565 11070 1580
rect 11085 1700 11125 1715
rect 11085 1680 11095 1700
rect 11115 1680 11125 1700
rect 11085 1650 11125 1680
rect 11085 1630 11095 1650
rect 11115 1630 11125 1650
rect 11085 1600 11125 1630
rect 11085 1580 11095 1600
rect 11115 1580 11125 1600
rect 11085 1565 11125 1580
rect 11140 1700 11180 1715
rect 11140 1680 11150 1700
rect 11170 1680 11180 1700
rect 11140 1650 11180 1680
rect 11140 1630 11150 1650
rect 11170 1630 11180 1650
rect 11140 1600 11180 1630
rect 11140 1580 11150 1600
rect 11170 1580 11180 1600
rect 11140 1565 11180 1580
rect 11195 1700 11235 1715
rect 11195 1680 11205 1700
rect 11225 1680 11235 1700
rect 11195 1650 11235 1680
rect 11195 1630 11205 1650
rect 11225 1630 11235 1650
rect 11195 1600 11235 1630
rect 11195 1580 11205 1600
rect 11225 1580 11235 1600
rect 11195 1565 11235 1580
rect 11250 1700 11290 1715
rect 11250 1680 11260 1700
rect 11280 1680 11290 1700
rect 11250 1650 11290 1680
rect 11250 1630 11260 1650
rect 11280 1630 11290 1650
rect 11250 1600 11290 1630
rect 11250 1580 11260 1600
rect 11280 1580 11290 1600
rect 11250 1565 11290 1580
rect 11305 1700 11345 1715
rect 11305 1680 11315 1700
rect 11335 1680 11345 1700
rect 11305 1650 11345 1680
rect 11305 1630 11315 1650
rect 11335 1630 11345 1650
rect 11305 1600 11345 1630
rect 11305 1580 11315 1600
rect 11335 1580 11345 1600
rect 11305 1565 11345 1580
rect 11360 1700 11400 1715
rect 11360 1680 11370 1700
rect 11390 1680 11400 1700
rect 11360 1650 11400 1680
rect 11360 1630 11370 1650
rect 11390 1630 11400 1650
rect 11360 1600 11400 1630
rect 11360 1580 11370 1600
rect 11390 1580 11400 1600
rect 11360 1565 11400 1580
rect 11415 1700 11455 1715
rect 11415 1680 11425 1700
rect 11445 1680 11455 1700
rect 11415 1650 11455 1680
rect 11415 1630 11425 1650
rect 11445 1630 11455 1650
rect 11415 1600 11455 1630
rect 11415 1580 11425 1600
rect 11445 1580 11455 1600
rect 11415 1565 11455 1580
rect 11470 1700 11510 1715
rect 11470 1680 11480 1700
rect 11500 1680 11510 1700
rect 11470 1650 11510 1680
rect 11470 1630 11480 1650
rect 11500 1630 11510 1650
rect 11470 1600 11510 1630
rect 11470 1580 11480 1600
rect 11500 1580 11510 1600
rect 11470 1565 11510 1580
rect 11525 1700 11565 1715
rect 11525 1680 11535 1700
rect 11555 1680 11565 1700
rect 11525 1650 11565 1680
rect 11525 1630 11535 1650
rect 11555 1630 11565 1650
rect 11525 1600 11565 1630
rect 11525 1580 11535 1600
rect 11555 1580 11565 1600
rect 11525 1565 11565 1580
rect 11580 1700 11620 1715
rect 11580 1680 11590 1700
rect 11610 1680 11620 1700
rect 11580 1650 11620 1680
rect 11580 1630 11590 1650
rect 11610 1630 11620 1650
rect 11580 1600 11620 1630
rect 11580 1580 11590 1600
rect 11610 1580 11620 1600
rect 11580 1565 11620 1580
rect 11635 1700 11675 1715
rect 11635 1680 11645 1700
rect 11665 1680 11675 1700
rect 11635 1650 11675 1680
rect 11635 1630 11645 1650
rect 11665 1630 11675 1650
rect 11635 1600 11675 1630
rect 11635 1580 11645 1600
rect 11665 1580 11675 1600
rect 11635 1565 11675 1580
rect 11690 1700 11730 1715
rect 11770 1700 11810 1715
rect 11690 1680 11700 1700
rect 11720 1680 11730 1700
rect 11770 1680 11780 1700
rect 11800 1680 11810 1700
rect 11690 1650 11730 1680
rect 11770 1650 11810 1680
rect 11690 1630 11700 1650
rect 11720 1630 11730 1650
rect 11770 1630 11780 1650
rect 11800 1630 11810 1650
rect 11690 1600 11730 1630
rect 11770 1600 11810 1630
rect 11690 1580 11700 1600
rect 11720 1580 11730 1600
rect 11770 1580 11780 1600
rect 11800 1580 11810 1600
rect 11690 1565 11730 1580
rect 11770 1565 11810 1580
rect 11825 1700 11865 1715
rect 11825 1680 11835 1700
rect 11855 1680 11865 1700
rect 11825 1650 11865 1680
rect 11825 1630 11835 1650
rect 11855 1630 11865 1650
rect 11825 1600 11865 1630
rect 11825 1580 11835 1600
rect 11855 1580 11865 1600
rect 11825 1565 11865 1580
rect 11880 1700 11920 1715
rect 11880 1680 11890 1700
rect 11910 1680 11920 1700
rect 11880 1650 11920 1680
rect 11880 1630 11890 1650
rect 11910 1630 11920 1650
rect 11880 1600 11920 1630
rect 11880 1580 11890 1600
rect 11910 1580 11920 1600
rect 11880 1565 11920 1580
rect 11935 1700 11975 1715
rect 11935 1680 11945 1700
rect 11965 1680 11975 1700
rect 11935 1650 11975 1680
rect 11935 1630 11945 1650
rect 11965 1630 11975 1650
rect 11935 1600 11975 1630
rect 11935 1580 11945 1600
rect 11965 1580 11975 1600
rect 11935 1565 11975 1580
rect 11990 1700 12030 1715
rect 12070 1700 12110 1715
rect 11990 1680 12000 1700
rect 12020 1680 12030 1700
rect 12070 1680 12080 1700
rect 12100 1680 12110 1700
rect 11990 1650 12030 1680
rect 12070 1650 12110 1680
rect 11990 1630 12000 1650
rect 12020 1630 12030 1650
rect 12070 1630 12080 1650
rect 12100 1630 12110 1650
rect 11990 1600 12030 1630
rect 12070 1600 12110 1630
rect 11990 1580 12000 1600
rect 12020 1580 12030 1600
rect 12070 1580 12080 1600
rect 12100 1580 12110 1600
rect 11990 1565 12030 1580
rect 12070 1565 12110 1580
rect 12125 1700 12165 1715
rect 12125 1680 12135 1700
rect 12155 1680 12165 1700
rect 12125 1650 12165 1680
rect 12125 1630 12135 1650
rect 12155 1630 12165 1650
rect 12125 1600 12165 1630
rect 12125 1580 12135 1600
rect 12155 1580 12165 1600
rect 12125 1565 12165 1580
rect 12180 1700 12220 1715
rect 12180 1680 12190 1700
rect 12210 1680 12220 1700
rect 12180 1650 12220 1680
rect 12180 1630 12190 1650
rect 12210 1630 12220 1650
rect 12180 1600 12220 1630
rect 12180 1580 12190 1600
rect 12210 1580 12220 1600
rect 12180 1565 12220 1580
rect 12235 1700 12275 1715
rect 12235 1680 12245 1700
rect 12265 1680 12275 1700
rect 12235 1650 12275 1680
rect 12235 1630 12245 1650
rect 12265 1630 12275 1650
rect 12235 1600 12275 1630
rect 12235 1580 12245 1600
rect 12265 1580 12275 1600
rect 12235 1565 12275 1580
rect 12290 1700 12330 1715
rect 12290 1680 12300 1700
rect 12320 1680 12330 1700
rect 12290 1650 12330 1680
rect 12290 1630 12300 1650
rect 12320 1630 12330 1650
rect 12290 1600 12330 1630
rect 12290 1580 12300 1600
rect 12320 1580 12330 1600
rect 12290 1565 12330 1580
rect 12345 1700 12385 1715
rect 12345 1680 12355 1700
rect 12375 1680 12385 1700
rect 12345 1650 12385 1680
rect 12345 1630 12355 1650
rect 12375 1630 12385 1650
rect 12345 1600 12385 1630
rect 12345 1580 12355 1600
rect 12375 1580 12385 1600
rect 12345 1565 12385 1580
rect 12400 1700 12440 1715
rect 12400 1680 12410 1700
rect 12430 1680 12440 1700
rect 12400 1650 12440 1680
rect 12400 1630 12410 1650
rect 12430 1630 12440 1650
rect 12400 1600 12440 1630
rect 12400 1580 12410 1600
rect 12430 1580 12440 1600
rect 12400 1565 12440 1580
rect 12455 1700 12495 1715
rect 12455 1680 12465 1700
rect 12485 1680 12495 1700
rect 12455 1650 12495 1680
rect 12455 1630 12465 1650
rect 12485 1630 12495 1650
rect 12455 1600 12495 1630
rect 12455 1580 12465 1600
rect 12485 1580 12495 1600
rect 12455 1565 12495 1580
rect 12510 1700 12550 1715
rect 12510 1680 12520 1700
rect 12540 1680 12550 1700
rect 12510 1650 12550 1680
rect 12510 1630 12520 1650
rect 12540 1630 12550 1650
rect 12510 1600 12550 1630
rect 12510 1580 12520 1600
rect 12540 1580 12550 1600
rect 12510 1565 12550 1580
rect 12565 1700 12605 1715
rect 12565 1680 12575 1700
rect 12595 1680 12605 1700
rect 12565 1650 12605 1680
rect 12565 1630 12575 1650
rect 12595 1630 12605 1650
rect 12565 1600 12605 1630
rect 12565 1580 12575 1600
rect 12595 1580 12605 1600
rect 12565 1565 12605 1580
rect 12620 1700 12660 1715
rect 12620 1680 12630 1700
rect 12650 1680 12660 1700
rect 12620 1650 12660 1680
rect 12620 1630 12630 1650
rect 12650 1630 12660 1650
rect 12620 1600 12660 1630
rect 12620 1580 12630 1600
rect 12650 1580 12660 1600
rect 12620 1565 12660 1580
rect 12675 1700 12715 1715
rect 12675 1680 12685 1700
rect 12705 1680 12715 1700
rect 12675 1650 12715 1680
rect 12675 1630 12685 1650
rect 12705 1630 12715 1650
rect 12675 1600 12715 1630
rect 12675 1580 12685 1600
rect 12705 1580 12715 1600
rect 12675 1565 12715 1580
rect 12730 1700 12770 1715
rect 12730 1680 12740 1700
rect 12760 1680 12770 1700
rect 12730 1650 12770 1680
rect 12730 1630 12740 1650
rect 12760 1630 12770 1650
rect 12730 1600 12770 1630
rect 12730 1580 12740 1600
rect 12760 1580 12770 1600
rect 12730 1565 12770 1580
rect 2835 1440 2875 1455
rect 2835 1420 2845 1440
rect 2865 1420 2875 1440
rect 2835 1390 2875 1420
rect 2835 1370 2845 1390
rect 2865 1370 2875 1390
rect 2835 1340 2875 1370
rect 2835 1320 2845 1340
rect 2865 1320 2875 1340
rect 2835 1290 2875 1320
rect 2835 1270 2845 1290
rect 2865 1270 2875 1290
rect 2835 1240 2875 1270
rect 2835 1220 2845 1240
rect 2865 1220 2875 1240
rect 2835 1205 2875 1220
rect 3375 1440 3415 1455
rect 3375 1420 3385 1440
rect 3405 1420 3415 1440
rect 3375 1390 3415 1420
rect 3375 1370 3385 1390
rect 3405 1370 3415 1390
rect 3375 1340 3415 1370
rect 3375 1320 3385 1340
rect 3405 1320 3415 1340
rect 3375 1290 3415 1320
rect 3375 1270 3385 1290
rect 3405 1270 3415 1290
rect 3375 1240 3415 1270
rect 3375 1220 3385 1240
rect 3405 1220 3415 1240
rect 3375 1205 3415 1220
rect 3915 1440 3955 1455
rect 3915 1420 3925 1440
rect 3945 1420 3955 1440
rect 3915 1390 3955 1420
rect 3915 1370 3925 1390
rect 3945 1370 3955 1390
rect 3915 1340 3955 1370
rect 3915 1320 3925 1340
rect 3945 1320 3955 1340
rect 3915 1290 3955 1320
rect 3915 1270 3925 1290
rect 3945 1270 3955 1290
rect 3915 1240 3955 1270
rect 3915 1220 3925 1240
rect 3945 1220 3955 1240
rect 3915 1205 3955 1220
rect 4055 1440 4095 1455
rect 4055 1420 4065 1440
rect 4085 1420 4095 1440
rect 4055 1390 4095 1420
rect 4055 1370 4065 1390
rect 4085 1370 4095 1390
rect 4055 1340 4095 1370
rect 4055 1320 4065 1340
rect 4085 1320 4095 1340
rect 4055 1290 4095 1320
rect 4055 1270 4065 1290
rect 4085 1270 4095 1290
rect 4055 1240 4095 1270
rect 4055 1220 4065 1240
rect 4085 1220 4095 1240
rect 4055 1205 4095 1220
rect 4595 1440 4635 1455
rect 4595 1420 4605 1440
rect 4625 1420 4635 1440
rect 4595 1390 4635 1420
rect 4595 1370 4605 1390
rect 4625 1370 4635 1390
rect 4595 1340 4635 1370
rect 4595 1320 4605 1340
rect 4625 1320 4635 1340
rect 4595 1290 4635 1320
rect 4595 1270 4605 1290
rect 4625 1270 4635 1290
rect 4595 1240 4635 1270
rect 4595 1220 4605 1240
rect 4625 1220 4635 1240
rect 4595 1205 4635 1220
rect 5135 1440 5175 1455
rect 5135 1420 5145 1440
rect 5165 1420 5175 1440
rect 5135 1390 5175 1420
rect 5135 1370 5145 1390
rect 5165 1370 5175 1390
rect 5135 1340 5175 1370
rect 5135 1320 5145 1340
rect 5165 1320 5175 1340
rect 5135 1290 5175 1320
rect 5135 1270 5145 1290
rect 5165 1270 5175 1290
rect 5135 1240 5175 1270
rect 5135 1220 5145 1240
rect 5165 1220 5175 1240
rect 5135 1205 5175 1220
rect 11205 1260 11245 1275
rect 11205 1240 11215 1260
rect 11235 1240 11245 1260
rect 11205 1210 11245 1240
rect 11205 1190 11215 1210
rect 11235 1190 11245 1210
rect 11205 1160 11245 1190
rect 11205 1140 11215 1160
rect 11235 1140 11245 1160
rect 11205 1110 11245 1140
rect 11205 1090 11215 1110
rect 11235 1090 11245 1110
rect 2945 1060 2985 1075
rect 2945 1040 2955 1060
rect 2975 1040 2985 1060
rect 2945 1010 2985 1040
rect 2945 990 2955 1010
rect 2975 990 2985 1010
rect 2945 975 2985 990
rect 3985 1060 4025 1075
rect 3985 1040 3995 1060
rect 4015 1040 4025 1060
rect 3985 1010 4025 1040
rect 3985 990 3995 1010
rect 4015 990 4025 1010
rect 3985 975 4025 990
rect 5025 1060 5065 1075
rect 5025 1040 5035 1060
rect 5055 1040 5065 1060
rect 5025 1010 5065 1040
rect 11205 1060 11245 1090
rect 11205 1040 11215 1060
rect 11235 1040 11245 1060
rect 11205 1025 11245 1040
rect 11260 1260 11300 1275
rect 11260 1240 11270 1260
rect 11290 1240 11300 1260
rect 11260 1210 11300 1240
rect 11260 1190 11270 1210
rect 11290 1190 11300 1210
rect 11260 1160 11300 1190
rect 11260 1140 11270 1160
rect 11290 1140 11300 1160
rect 11260 1110 11300 1140
rect 11260 1090 11270 1110
rect 11290 1090 11300 1110
rect 11260 1060 11300 1090
rect 11260 1040 11270 1060
rect 11290 1040 11300 1060
rect 11260 1025 11300 1040
rect 11315 1260 11355 1275
rect 11315 1240 11325 1260
rect 11345 1240 11355 1260
rect 11315 1210 11355 1240
rect 11315 1190 11325 1210
rect 11345 1190 11355 1210
rect 11315 1160 11355 1190
rect 11315 1140 11325 1160
rect 11345 1140 11355 1160
rect 11315 1110 11355 1140
rect 11315 1090 11325 1110
rect 11345 1090 11355 1110
rect 11315 1060 11355 1090
rect 11315 1040 11325 1060
rect 11345 1040 11355 1060
rect 11315 1025 11355 1040
rect 11370 1260 11410 1275
rect 11370 1240 11380 1260
rect 11400 1240 11410 1260
rect 11370 1210 11410 1240
rect 11370 1190 11380 1210
rect 11400 1190 11410 1210
rect 11370 1160 11410 1190
rect 11370 1140 11380 1160
rect 11400 1140 11410 1160
rect 11370 1110 11410 1140
rect 11370 1090 11380 1110
rect 11400 1090 11410 1110
rect 11370 1060 11410 1090
rect 11370 1040 11380 1060
rect 11400 1040 11410 1060
rect 11370 1025 11410 1040
rect 11425 1260 11465 1275
rect 11425 1240 11435 1260
rect 11455 1240 11465 1260
rect 11425 1210 11465 1240
rect 11425 1190 11435 1210
rect 11455 1190 11465 1210
rect 11425 1160 11465 1190
rect 11425 1140 11435 1160
rect 11455 1140 11465 1160
rect 11425 1110 11465 1140
rect 11425 1090 11435 1110
rect 11455 1090 11465 1110
rect 11425 1060 11465 1090
rect 11425 1040 11435 1060
rect 11455 1040 11465 1060
rect 11425 1025 11465 1040
rect 11480 1260 11520 1275
rect 11480 1240 11490 1260
rect 11510 1240 11520 1260
rect 11480 1210 11520 1240
rect 11480 1190 11490 1210
rect 11510 1190 11520 1210
rect 11480 1160 11520 1190
rect 11480 1140 11490 1160
rect 11510 1140 11520 1160
rect 11480 1110 11520 1140
rect 11480 1090 11490 1110
rect 11510 1090 11520 1110
rect 11480 1060 11520 1090
rect 11480 1040 11490 1060
rect 11510 1040 11520 1060
rect 11480 1025 11520 1040
rect 11535 1260 11575 1275
rect 11535 1240 11545 1260
rect 11565 1240 11575 1260
rect 11535 1210 11575 1240
rect 11535 1190 11545 1210
rect 11565 1190 11575 1210
rect 11535 1160 11575 1190
rect 11535 1140 11545 1160
rect 11565 1140 11575 1160
rect 11535 1110 11575 1140
rect 11535 1090 11545 1110
rect 11565 1090 11575 1110
rect 11535 1060 11575 1090
rect 11535 1040 11545 1060
rect 11565 1040 11575 1060
rect 11535 1025 11575 1040
rect 11590 1260 11630 1275
rect 11590 1240 11600 1260
rect 11620 1240 11630 1260
rect 11590 1210 11630 1240
rect 11590 1190 11600 1210
rect 11620 1190 11630 1210
rect 11590 1160 11630 1190
rect 11590 1140 11600 1160
rect 11620 1140 11630 1160
rect 11590 1110 11630 1140
rect 11590 1090 11600 1110
rect 11620 1090 11630 1110
rect 11590 1060 11630 1090
rect 11590 1040 11600 1060
rect 11620 1040 11630 1060
rect 11590 1025 11630 1040
rect 11645 1260 11685 1275
rect 11645 1240 11655 1260
rect 11675 1240 11685 1260
rect 11645 1210 11685 1240
rect 11645 1190 11655 1210
rect 11675 1190 11685 1210
rect 11645 1160 11685 1190
rect 11645 1140 11655 1160
rect 11675 1140 11685 1160
rect 11645 1110 11685 1140
rect 11645 1090 11655 1110
rect 11675 1090 11685 1110
rect 11645 1060 11685 1090
rect 11645 1040 11655 1060
rect 11675 1040 11685 1060
rect 11645 1025 11685 1040
rect 11700 1260 11740 1275
rect 11700 1240 11710 1260
rect 11730 1240 11740 1260
rect 11700 1210 11740 1240
rect 11700 1190 11710 1210
rect 11730 1190 11740 1210
rect 11700 1160 11740 1190
rect 11700 1140 11710 1160
rect 11730 1140 11740 1160
rect 11700 1110 11740 1140
rect 11700 1090 11710 1110
rect 11730 1090 11740 1110
rect 11700 1060 11740 1090
rect 11700 1040 11710 1060
rect 11730 1040 11740 1060
rect 11700 1025 11740 1040
rect 11755 1260 11795 1275
rect 11755 1240 11765 1260
rect 11785 1240 11795 1260
rect 11755 1210 11795 1240
rect 11755 1190 11765 1210
rect 11785 1190 11795 1210
rect 11755 1160 11795 1190
rect 11755 1140 11765 1160
rect 11785 1140 11795 1160
rect 11755 1110 11795 1140
rect 11755 1090 11765 1110
rect 11785 1090 11795 1110
rect 11755 1060 11795 1090
rect 11755 1040 11765 1060
rect 11785 1040 11795 1060
rect 11755 1025 11795 1040
rect 11810 1260 11850 1275
rect 11810 1240 11820 1260
rect 11840 1240 11850 1260
rect 11810 1210 11850 1240
rect 11810 1190 11820 1210
rect 11840 1190 11850 1210
rect 11810 1160 11850 1190
rect 11810 1140 11820 1160
rect 11840 1140 11850 1160
rect 11810 1110 11850 1140
rect 11810 1090 11820 1110
rect 11840 1090 11850 1110
rect 11810 1060 11850 1090
rect 11810 1040 11820 1060
rect 11840 1040 11850 1060
rect 11810 1025 11850 1040
rect 11865 1260 11905 1275
rect 11865 1240 11875 1260
rect 11895 1240 11905 1260
rect 11865 1210 11905 1240
rect 11865 1190 11875 1210
rect 11895 1190 11905 1210
rect 11865 1160 11905 1190
rect 11865 1140 11875 1160
rect 11895 1140 11905 1160
rect 11865 1110 11905 1140
rect 11865 1090 11875 1110
rect 11895 1090 11905 1110
rect 11865 1060 11905 1090
rect 11865 1040 11875 1060
rect 11895 1040 11905 1060
rect 11865 1025 11905 1040
rect 11920 1260 11960 1275
rect 11920 1240 11930 1260
rect 11950 1240 11960 1260
rect 11920 1210 11960 1240
rect 11920 1190 11930 1210
rect 11950 1190 11960 1210
rect 11920 1160 11960 1190
rect 11920 1140 11930 1160
rect 11950 1140 11960 1160
rect 11920 1110 11960 1140
rect 11920 1090 11930 1110
rect 11950 1090 11960 1110
rect 11920 1060 11960 1090
rect 11920 1040 11930 1060
rect 11950 1040 11960 1060
rect 11920 1025 11960 1040
rect 11975 1260 12015 1275
rect 11975 1240 11985 1260
rect 12005 1240 12015 1260
rect 11975 1210 12015 1240
rect 11975 1190 11985 1210
rect 12005 1190 12015 1210
rect 11975 1160 12015 1190
rect 11975 1140 11985 1160
rect 12005 1140 12015 1160
rect 11975 1110 12015 1140
rect 11975 1090 11985 1110
rect 12005 1090 12015 1110
rect 11975 1060 12015 1090
rect 11975 1040 11985 1060
rect 12005 1040 12015 1060
rect 11975 1025 12015 1040
rect 12030 1260 12070 1275
rect 12030 1240 12040 1260
rect 12060 1240 12070 1260
rect 12030 1210 12070 1240
rect 12030 1190 12040 1210
rect 12060 1190 12070 1210
rect 12030 1160 12070 1190
rect 12030 1140 12040 1160
rect 12060 1140 12070 1160
rect 12030 1110 12070 1140
rect 12030 1090 12040 1110
rect 12060 1090 12070 1110
rect 12030 1060 12070 1090
rect 12030 1040 12040 1060
rect 12060 1040 12070 1060
rect 12030 1025 12070 1040
rect 12085 1260 12125 1275
rect 12085 1240 12095 1260
rect 12115 1240 12125 1260
rect 12085 1210 12125 1240
rect 12085 1190 12095 1210
rect 12115 1190 12125 1210
rect 12085 1160 12125 1190
rect 12085 1140 12095 1160
rect 12115 1140 12125 1160
rect 12085 1110 12125 1140
rect 12085 1090 12095 1110
rect 12115 1090 12125 1110
rect 12085 1060 12125 1090
rect 12085 1040 12095 1060
rect 12115 1040 12125 1060
rect 12085 1025 12125 1040
rect 12140 1260 12180 1275
rect 12140 1240 12150 1260
rect 12170 1240 12180 1260
rect 12140 1210 12180 1240
rect 12140 1190 12150 1210
rect 12170 1190 12180 1210
rect 12140 1160 12180 1190
rect 12140 1140 12150 1160
rect 12170 1140 12180 1160
rect 12140 1110 12180 1140
rect 12140 1090 12150 1110
rect 12170 1090 12180 1110
rect 12140 1060 12180 1090
rect 12140 1040 12150 1060
rect 12170 1040 12180 1060
rect 12140 1025 12180 1040
rect 12195 1260 12235 1275
rect 12195 1240 12205 1260
rect 12225 1240 12235 1260
rect 12195 1210 12235 1240
rect 12195 1190 12205 1210
rect 12225 1190 12235 1210
rect 12195 1160 12235 1190
rect 12195 1140 12205 1160
rect 12225 1140 12235 1160
rect 12195 1110 12235 1140
rect 12195 1090 12205 1110
rect 12225 1090 12235 1110
rect 12195 1060 12235 1090
rect 12195 1040 12205 1060
rect 12225 1040 12235 1060
rect 12195 1025 12235 1040
rect 12250 1260 12290 1275
rect 12250 1240 12260 1260
rect 12280 1240 12290 1260
rect 12250 1210 12290 1240
rect 12250 1190 12260 1210
rect 12280 1190 12290 1210
rect 12250 1160 12290 1190
rect 12250 1140 12260 1160
rect 12280 1140 12290 1160
rect 12250 1110 12290 1140
rect 12250 1090 12260 1110
rect 12280 1090 12290 1110
rect 12250 1060 12290 1090
rect 12250 1040 12260 1060
rect 12280 1040 12290 1060
rect 12250 1025 12290 1040
rect 12305 1260 12345 1275
rect 12305 1240 12315 1260
rect 12335 1240 12345 1260
rect 12305 1210 12345 1240
rect 12305 1190 12315 1210
rect 12335 1190 12345 1210
rect 12305 1160 12345 1190
rect 12305 1140 12315 1160
rect 12335 1140 12345 1160
rect 12305 1110 12345 1140
rect 12305 1090 12315 1110
rect 12335 1090 12345 1110
rect 12305 1060 12345 1090
rect 12305 1040 12315 1060
rect 12335 1040 12345 1060
rect 12305 1025 12345 1040
rect 12360 1260 12400 1275
rect 12360 1240 12370 1260
rect 12390 1240 12400 1260
rect 12360 1210 12400 1240
rect 12360 1190 12370 1210
rect 12390 1190 12400 1210
rect 12360 1160 12400 1190
rect 12360 1140 12370 1160
rect 12390 1140 12400 1160
rect 12360 1110 12400 1140
rect 12360 1090 12370 1110
rect 12390 1090 12400 1110
rect 12360 1060 12400 1090
rect 12360 1040 12370 1060
rect 12390 1040 12400 1060
rect 12360 1025 12400 1040
rect 12415 1260 12455 1275
rect 12415 1240 12425 1260
rect 12445 1240 12455 1260
rect 12415 1210 12455 1240
rect 12415 1190 12425 1210
rect 12445 1190 12455 1210
rect 12415 1160 12455 1190
rect 12415 1140 12425 1160
rect 12445 1140 12455 1160
rect 12415 1110 12455 1140
rect 12415 1090 12425 1110
rect 12445 1090 12455 1110
rect 12415 1060 12455 1090
rect 12415 1040 12425 1060
rect 12445 1040 12455 1060
rect 12415 1025 12455 1040
rect 12470 1260 12510 1275
rect 12470 1240 12480 1260
rect 12500 1240 12510 1260
rect 12470 1210 12510 1240
rect 12470 1190 12480 1210
rect 12500 1190 12510 1210
rect 12470 1160 12510 1190
rect 12470 1140 12480 1160
rect 12500 1140 12510 1160
rect 12470 1110 12510 1140
rect 12470 1090 12480 1110
rect 12500 1090 12510 1110
rect 12470 1060 12510 1090
rect 12470 1040 12480 1060
rect 12500 1040 12510 1060
rect 12470 1025 12510 1040
rect 12525 1260 12565 1275
rect 12525 1240 12535 1260
rect 12555 1240 12565 1260
rect 12525 1210 12565 1240
rect 12525 1190 12535 1210
rect 12555 1190 12565 1210
rect 12525 1160 12565 1190
rect 12525 1140 12535 1160
rect 12555 1140 12565 1160
rect 12525 1110 12565 1140
rect 12525 1090 12535 1110
rect 12555 1090 12565 1110
rect 12525 1060 12565 1090
rect 12525 1040 12535 1060
rect 12555 1040 12565 1060
rect 12525 1025 12565 1040
rect 12580 1260 12620 1275
rect 12580 1240 12590 1260
rect 12610 1240 12620 1260
rect 12580 1210 12620 1240
rect 12580 1190 12590 1210
rect 12610 1190 12620 1210
rect 12580 1160 12620 1190
rect 12580 1140 12590 1160
rect 12610 1140 12620 1160
rect 12580 1110 12620 1140
rect 12580 1090 12590 1110
rect 12610 1090 12620 1110
rect 12580 1060 12620 1090
rect 12580 1040 12590 1060
rect 12610 1040 12620 1060
rect 12580 1025 12620 1040
rect 5025 990 5035 1010
rect 5055 990 5065 1010
rect 5025 975 5065 990
rect 2995 865 3035 880
rect 2995 845 3005 865
rect 3025 845 3035 865
rect 2995 815 3035 845
rect 2995 795 3005 815
rect 3025 795 3035 815
rect 2995 780 3035 795
rect 3085 865 3125 880
rect 3085 845 3095 865
rect 3115 845 3125 865
rect 3085 815 3125 845
rect 3085 795 3095 815
rect 3115 795 3125 815
rect 3085 780 3125 795
rect 3175 865 3215 880
rect 3175 845 3185 865
rect 3205 845 3215 865
rect 3175 815 3215 845
rect 3175 795 3185 815
rect 3205 795 3215 815
rect 3175 780 3215 795
rect 3265 865 3305 880
rect 3265 845 3275 865
rect 3295 845 3305 865
rect 3265 815 3305 845
rect 3265 795 3275 815
rect 3295 795 3305 815
rect 3265 780 3305 795
rect 3355 865 3395 880
rect 3355 845 3365 865
rect 3385 845 3395 865
rect 3355 815 3395 845
rect 3355 795 3365 815
rect 3385 795 3395 815
rect 3355 780 3395 795
rect 3445 865 3485 880
rect 3445 845 3455 865
rect 3475 845 3485 865
rect 3445 815 3485 845
rect 3445 795 3455 815
rect 3475 795 3485 815
rect 3445 780 3485 795
rect 3535 865 3575 880
rect 3535 845 3545 865
rect 3565 845 3575 865
rect 3535 815 3575 845
rect 3535 795 3545 815
rect 3565 795 3575 815
rect 3535 780 3575 795
rect 3625 865 3665 880
rect 3625 845 3635 865
rect 3655 845 3665 865
rect 3625 815 3665 845
rect 3625 795 3635 815
rect 3655 795 3665 815
rect 3625 780 3665 795
rect 3715 865 3755 880
rect 3715 845 3725 865
rect 3745 845 3755 865
rect 3715 815 3755 845
rect 3715 795 3725 815
rect 3745 795 3755 815
rect 3715 780 3755 795
rect 3805 865 3845 880
rect 3805 845 3815 865
rect 3835 845 3845 865
rect 3805 815 3845 845
rect 3805 795 3815 815
rect 3835 795 3845 815
rect 3805 780 3845 795
rect 3895 865 3935 880
rect 3895 845 3905 865
rect 3925 845 3935 865
rect 3895 815 3935 845
rect 3895 795 3905 815
rect 3925 795 3935 815
rect 3895 780 3935 795
rect 3985 865 4025 880
rect 3985 845 3995 865
rect 4015 845 4025 865
rect 3985 815 4025 845
rect 3985 795 3995 815
rect 4015 795 4025 815
rect 3985 780 4025 795
rect 4075 865 4115 880
rect 4075 845 4085 865
rect 4105 845 4115 865
rect 4075 815 4115 845
rect 4075 795 4085 815
rect 4105 795 4115 815
rect 4075 780 4115 795
rect 4165 865 4205 880
rect 4165 845 4175 865
rect 4195 845 4205 865
rect 4165 815 4205 845
rect 4165 795 4175 815
rect 4195 795 4205 815
rect 4165 780 4205 795
rect 4255 865 4295 880
rect 4255 845 4265 865
rect 4285 845 4295 865
rect 4255 815 4295 845
rect 4255 795 4265 815
rect 4285 795 4295 815
rect 4255 780 4295 795
rect 4345 865 4385 880
rect 4345 845 4355 865
rect 4375 845 4385 865
rect 4345 815 4385 845
rect 4345 795 4355 815
rect 4375 795 4385 815
rect 4345 780 4385 795
rect 4435 865 4475 880
rect 4435 845 4445 865
rect 4465 845 4475 865
rect 4435 815 4475 845
rect 4435 795 4445 815
rect 4465 795 4475 815
rect 4435 780 4475 795
rect 4525 865 4565 880
rect 4525 845 4535 865
rect 4555 845 4565 865
rect 4525 815 4565 845
rect 4525 795 4535 815
rect 4555 795 4565 815
rect 4525 780 4565 795
rect 4615 865 4655 880
rect 4615 845 4625 865
rect 4645 845 4655 865
rect 4615 815 4655 845
rect 4615 795 4625 815
rect 4645 795 4655 815
rect 4615 780 4655 795
rect 4705 865 4745 880
rect 4705 845 4715 865
rect 4735 845 4745 865
rect 4705 815 4745 845
rect 4705 795 4715 815
rect 4735 795 4745 815
rect 4705 780 4745 795
rect 4795 865 4835 880
rect 4795 845 4805 865
rect 4825 845 4835 865
rect 4795 815 4835 845
rect 4795 795 4805 815
rect 4825 795 4835 815
rect 4795 780 4835 795
rect 4885 865 4925 880
rect 4885 845 4895 865
rect 4915 845 4925 865
rect 4885 815 4925 845
rect 4885 795 4895 815
rect 4915 795 4925 815
rect 4885 780 4925 795
rect 4975 865 5015 880
rect 4975 845 4985 865
rect 5005 845 5015 865
rect 4975 815 5015 845
rect 4975 795 4985 815
rect 5005 795 5015 815
rect 4975 780 5015 795
<< pdiff >>
rect 2995 2915 3035 2930
rect 2995 2895 3005 2915
rect 3025 2895 3035 2915
rect 2995 2865 3035 2895
rect 2995 2845 3005 2865
rect 3025 2845 3035 2865
rect 2995 2830 3035 2845
rect 3085 2915 3125 2930
rect 3085 2895 3095 2915
rect 3115 2895 3125 2915
rect 3085 2865 3125 2895
rect 3085 2845 3095 2865
rect 3115 2845 3125 2865
rect 3085 2830 3125 2845
rect 3175 2915 3215 2930
rect 3175 2895 3185 2915
rect 3205 2895 3215 2915
rect 3175 2865 3215 2895
rect 3175 2845 3185 2865
rect 3205 2845 3215 2865
rect 3175 2830 3215 2845
rect 3265 2915 3305 2930
rect 3265 2895 3275 2915
rect 3295 2895 3305 2915
rect 3265 2865 3305 2895
rect 3265 2845 3275 2865
rect 3295 2845 3305 2865
rect 3265 2830 3305 2845
rect 3355 2915 3395 2930
rect 3355 2895 3365 2915
rect 3385 2895 3395 2915
rect 3355 2865 3395 2895
rect 3355 2845 3365 2865
rect 3385 2845 3395 2865
rect 3355 2830 3395 2845
rect 3445 2915 3485 2930
rect 3445 2895 3455 2915
rect 3475 2895 3485 2915
rect 3445 2865 3485 2895
rect 3445 2845 3455 2865
rect 3475 2845 3485 2865
rect 3445 2830 3485 2845
rect 3535 2915 3575 2930
rect 3535 2895 3545 2915
rect 3565 2895 3575 2915
rect 3535 2865 3575 2895
rect 3535 2845 3545 2865
rect 3565 2845 3575 2865
rect 3535 2830 3575 2845
rect 3625 2915 3665 2930
rect 3625 2895 3635 2915
rect 3655 2895 3665 2915
rect 3625 2865 3665 2895
rect 3625 2845 3635 2865
rect 3655 2845 3665 2865
rect 3625 2830 3665 2845
rect 3715 2915 3755 2930
rect 3715 2895 3725 2915
rect 3745 2895 3755 2915
rect 3715 2865 3755 2895
rect 3715 2845 3725 2865
rect 3745 2845 3755 2865
rect 3715 2830 3755 2845
rect 3805 2915 3845 2930
rect 3805 2895 3815 2915
rect 3835 2895 3845 2915
rect 3805 2865 3845 2895
rect 3805 2845 3815 2865
rect 3835 2845 3845 2865
rect 3805 2830 3845 2845
rect 3895 2915 3935 2930
rect 3895 2895 3905 2915
rect 3925 2895 3935 2915
rect 3895 2865 3935 2895
rect 3895 2845 3905 2865
rect 3925 2845 3935 2865
rect 3895 2830 3935 2845
rect 3985 2915 4025 2930
rect 3985 2895 3995 2915
rect 4015 2895 4025 2915
rect 3985 2865 4025 2895
rect 3985 2845 3995 2865
rect 4015 2845 4025 2865
rect 3985 2830 4025 2845
rect 4075 2915 4115 2930
rect 4075 2895 4085 2915
rect 4105 2895 4115 2915
rect 4075 2865 4115 2895
rect 4075 2845 4085 2865
rect 4105 2845 4115 2865
rect 4075 2830 4115 2845
rect 4165 2915 4205 2930
rect 4165 2895 4175 2915
rect 4195 2895 4205 2915
rect 4165 2865 4205 2895
rect 4165 2845 4175 2865
rect 4195 2845 4205 2865
rect 4165 2830 4205 2845
rect 4255 2915 4295 2930
rect 4255 2895 4265 2915
rect 4285 2895 4295 2915
rect 4255 2865 4295 2895
rect 4255 2845 4265 2865
rect 4285 2845 4295 2865
rect 4255 2830 4295 2845
rect 4345 2915 4385 2930
rect 4345 2895 4355 2915
rect 4375 2895 4385 2915
rect 4345 2865 4385 2895
rect 4345 2845 4355 2865
rect 4375 2845 4385 2865
rect 4345 2830 4385 2845
rect 4435 2915 4475 2930
rect 4435 2895 4445 2915
rect 4465 2895 4475 2915
rect 4435 2865 4475 2895
rect 4435 2845 4445 2865
rect 4465 2845 4475 2865
rect 4435 2830 4475 2845
rect 4525 2915 4565 2930
rect 4525 2895 4535 2915
rect 4555 2895 4565 2915
rect 4525 2865 4565 2895
rect 4525 2845 4535 2865
rect 4555 2845 4565 2865
rect 4525 2830 4565 2845
rect 4615 2915 4655 2930
rect 4615 2895 4625 2915
rect 4645 2895 4655 2915
rect 4615 2865 4655 2895
rect 4615 2845 4625 2865
rect 4645 2845 4655 2865
rect 4615 2830 4655 2845
rect 4705 2915 4745 2930
rect 4705 2895 4715 2915
rect 4735 2895 4745 2915
rect 4705 2865 4745 2895
rect 4705 2845 4715 2865
rect 4735 2845 4745 2865
rect 4705 2830 4745 2845
rect 4795 2915 4835 2930
rect 4795 2895 4805 2915
rect 4825 2895 4835 2915
rect 4795 2865 4835 2895
rect 4795 2845 4805 2865
rect 4825 2845 4835 2865
rect 4795 2830 4835 2845
rect 4885 2915 4925 2930
rect 4885 2895 4895 2915
rect 4915 2895 4925 2915
rect 4885 2865 4925 2895
rect 4885 2845 4895 2865
rect 4915 2845 4925 2865
rect 4885 2830 4925 2845
rect 4975 2915 5015 2930
rect 4975 2895 4985 2915
rect 5005 2895 5015 2915
rect 4975 2865 5015 2895
rect 4975 2845 4985 2865
rect 5005 2845 5015 2865
rect 4975 2830 5015 2845
rect 3175 2685 3215 2700
rect 3175 2665 3185 2685
rect 3205 2665 3215 2685
rect 3175 2635 3215 2665
rect 3175 2615 3185 2635
rect 3205 2615 3215 2635
rect 3175 2585 3215 2615
rect 3175 2565 3185 2585
rect 3205 2565 3215 2585
rect 3175 2535 3215 2565
rect 3175 2515 3185 2535
rect 3205 2515 3215 2535
rect 3175 2485 3215 2515
rect 3175 2465 3185 2485
rect 3205 2465 3215 2485
rect 3175 2435 3215 2465
rect 3175 2415 3185 2435
rect 3205 2415 3215 2435
rect 3175 2400 3215 2415
rect 3265 2685 3305 2700
rect 3265 2665 3275 2685
rect 3295 2665 3305 2685
rect 3265 2635 3305 2665
rect 3265 2615 3275 2635
rect 3295 2615 3305 2635
rect 3265 2585 3305 2615
rect 3265 2565 3275 2585
rect 3295 2565 3305 2585
rect 3265 2535 3305 2565
rect 3265 2515 3275 2535
rect 3295 2515 3305 2535
rect 3265 2485 3305 2515
rect 3265 2465 3275 2485
rect 3295 2465 3305 2485
rect 3265 2435 3305 2465
rect 3265 2415 3275 2435
rect 3295 2415 3305 2435
rect 3265 2400 3305 2415
rect 3355 2685 3395 2700
rect 3355 2665 3365 2685
rect 3385 2665 3395 2685
rect 3355 2635 3395 2665
rect 3355 2615 3365 2635
rect 3385 2615 3395 2635
rect 3355 2585 3395 2615
rect 3355 2565 3365 2585
rect 3385 2565 3395 2585
rect 3355 2535 3395 2565
rect 3355 2515 3365 2535
rect 3385 2515 3395 2535
rect 3355 2485 3395 2515
rect 3355 2465 3365 2485
rect 3385 2465 3395 2485
rect 3355 2435 3395 2465
rect 3355 2415 3365 2435
rect 3385 2415 3395 2435
rect 3355 2400 3395 2415
rect 3445 2685 3485 2700
rect 3445 2665 3455 2685
rect 3475 2665 3485 2685
rect 3445 2635 3485 2665
rect 3445 2615 3455 2635
rect 3475 2615 3485 2635
rect 3445 2585 3485 2615
rect 3445 2565 3455 2585
rect 3475 2565 3485 2585
rect 3445 2535 3485 2565
rect 3445 2515 3455 2535
rect 3475 2515 3485 2535
rect 3445 2485 3485 2515
rect 3445 2465 3455 2485
rect 3475 2465 3485 2485
rect 3445 2435 3485 2465
rect 3445 2415 3455 2435
rect 3475 2415 3485 2435
rect 3445 2400 3485 2415
rect 3535 2685 3575 2700
rect 3535 2665 3545 2685
rect 3565 2665 3575 2685
rect 3535 2635 3575 2665
rect 3535 2615 3545 2635
rect 3565 2615 3575 2635
rect 3535 2585 3575 2615
rect 3535 2565 3545 2585
rect 3565 2565 3575 2585
rect 3535 2535 3575 2565
rect 3535 2515 3545 2535
rect 3565 2515 3575 2535
rect 3535 2485 3575 2515
rect 3535 2465 3545 2485
rect 3565 2465 3575 2485
rect 3535 2435 3575 2465
rect 3535 2415 3545 2435
rect 3565 2415 3575 2435
rect 3535 2400 3575 2415
rect 3625 2685 3665 2700
rect 3625 2665 3635 2685
rect 3655 2665 3665 2685
rect 3625 2635 3665 2665
rect 3625 2615 3635 2635
rect 3655 2615 3665 2635
rect 3625 2585 3665 2615
rect 3625 2565 3635 2585
rect 3655 2565 3665 2585
rect 3625 2535 3665 2565
rect 3625 2515 3635 2535
rect 3655 2515 3665 2535
rect 3625 2485 3665 2515
rect 3625 2465 3635 2485
rect 3655 2465 3665 2485
rect 3625 2435 3665 2465
rect 3625 2415 3635 2435
rect 3655 2415 3665 2435
rect 3625 2400 3665 2415
rect 3715 2685 3755 2700
rect 3715 2665 3725 2685
rect 3745 2665 3755 2685
rect 3715 2635 3755 2665
rect 3715 2615 3725 2635
rect 3745 2615 3755 2635
rect 3715 2585 3755 2615
rect 3715 2565 3725 2585
rect 3745 2565 3755 2585
rect 3715 2535 3755 2565
rect 3715 2515 3725 2535
rect 3745 2515 3755 2535
rect 3715 2485 3755 2515
rect 3715 2465 3725 2485
rect 3745 2465 3755 2485
rect 3715 2435 3755 2465
rect 3715 2415 3725 2435
rect 3745 2415 3755 2435
rect 3715 2400 3755 2415
rect 3805 2685 3845 2700
rect 3805 2665 3815 2685
rect 3835 2665 3845 2685
rect 3805 2635 3845 2665
rect 3805 2615 3815 2635
rect 3835 2615 3845 2635
rect 3805 2585 3845 2615
rect 3805 2565 3815 2585
rect 3835 2565 3845 2585
rect 3805 2535 3845 2565
rect 3805 2515 3815 2535
rect 3835 2515 3845 2535
rect 3805 2485 3845 2515
rect 3805 2465 3815 2485
rect 3835 2465 3845 2485
rect 3805 2435 3845 2465
rect 3805 2415 3815 2435
rect 3835 2415 3845 2435
rect 3805 2400 3845 2415
rect 3895 2685 3935 2700
rect 3895 2665 3905 2685
rect 3925 2665 3935 2685
rect 3895 2635 3935 2665
rect 3895 2615 3905 2635
rect 3925 2615 3935 2635
rect 3895 2585 3935 2615
rect 3895 2565 3905 2585
rect 3925 2565 3935 2585
rect 3895 2535 3935 2565
rect 3895 2515 3905 2535
rect 3925 2515 3935 2535
rect 3895 2485 3935 2515
rect 3895 2465 3905 2485
rect 3925 2465 3935 2485
rect 3895 2435 3935 2465
rect 3895 2415 3905 2435
rect 3925 2415 3935 2435
rect 3895 2400 3935 2415
rect 3985 2685 4025 2700
rect 3985 2665 3995 2685
rect 4015 2665 4025 2685
rect 3985 2635 4025 2665
rect 3985 2615 3995 2635
rect 4015 2615 4025 2635
rect 3985 2585 4025 2615
rect 3985 2565 3995 2585
rect 4015 2565 4025 2585
rect 3985 2535 4025 2565
rect 3985 2515 3995 2535
rect 4015 2515 4025 2535
rect 3985 2485 4025 2515
rect 3985 2465 3995 2485
rect 4015 2465 4025 2485
rect 3985 2435 4025 2465
rect 3985 2415 3995 2435
rect 4015 2415 4025 2435
rect 3985 2400 4025 2415
rect 4075 2685 4115 2700
rect 4075 2665 4085 2685
rect 4105 2665 4115 2685
rect 4075 2635 4115 2665
rect 4075 2615 4085 2635
rect 4105 2615 4115 2635
rect 4075 2585 4115 2615
rect 4075 2565 4085 2585
rect 4105 2565 4115 2585
rect 4075 2535 4115 2565
rect 4075 2515 4085 2535
rect 4105 2515 4115 2535
rect 4075 2485 4115 2515
rect 4075 2465 4085 2485
rect 4105 2465 4115 2485
rect 4075 2435 4115 2465
rect 4075 2415 4085 2435
rect 4105 2415 4115 2435
rect 4075 2400 4115 2415
rect 4165 2685 4205 2700
rect 4165 2665 4175 2685
rect 4195 2665 4205 2685
rect 4165 2635 4205 2665
rect 4165 2615 4175 2635
rect 4195 2615 4205 2635
rect 4165 2585 4205 2615
rect 4165 2565 4175 2585
rect 4195 2565 4205 2585
rect 4165 2535 4205 2565
rect 4165 2515 4175 2535
rect 4195 2515 4205 2535
rect 4165 2485 4205 2515
rect 4165 2465 4175 2485
rect 4195 2465 4205 2485
rect 4165 2435 4205 2465
rect 4165 2415 4175 2435
rect 4195 2415 4205 2435
rect 4165 2400 4205 2415
rect 4255 2685 4295 2700
rect 4255 2665 4265 2685
rect 4285 2665 4295 2685
rect 4255 2635 4295 2665
rect 4255 2615 4265 2635
rect 4285 2615 4295 2635
rect 4255 2585 4295 2615
rect 4255 2565 4265 2585
rect 4285 2565 4295 2585
rect 4255 2535 4295 2565
rect 4255 2515 4265 2535
rect 4285 2515 4295 2535
rect 4255 2485 4295 2515
rect 4255 2465 4265 2485
rect 4285 2465 4295 2485
rect 4255 2435 4295 2465
rect 4255 2415 4265 2435
rect 4285 2415 4295 2435
rect 4255 2400 4295 2415
rect 4345 2685 4385 2700
rect 4345 2665 4355 2685
rect 4375 2665 4385 2685
rect 4345 2635 4385 2665
rect 4345 2615 4355 2635
rect 4375 2615 4385 2635
rect 4345 2585 4385 2615
rect 4345 2565 4355 2585
rect 4375 2565 4385 2585
rect 4345 2535 4385 2565
rect 4345 2515 4355 2535
rect 4375 2515 4385 2535
rect 4345 2485 4385 2515
rect 4345 2465 4355 2485
rect 4375 2465 4385 2485
rect 4345 2435 4385 2465
rect 4345 2415 4355 2435
rect 4375 2415 4385 2435
rect 4345 2400 4385 2415
rect 4435 2685 4475 2700
rect 4435 2665 4445 2685
rect 4465 2665 4475 2685
rect 4435 2635 4475 2665
rect 4435 2615 4445 2635
rect 4465 2615 4475 2635
rect 4435 2585 4475 2615
rect 4435 2565 4445 2585
rect 4465 2565 4475 2585
rect 4435 2535 4475 2565
rect 4435 2515 4445 2535
rect 4465 2515 4475 2535
rect 4435 2485 4475 2515
rect 4435 2465 4445 2485
rect 4465 2465 4475 2485
rect 4435 2435 4475 2465
rect 4435 2415 4445 2435
rect 4465 2415 4475 2435
rect 4435 2400 4475 2415
rect 4525 2685 4565 2700
rect 4525 2665 4535 2685
rect 4555 2665 4565 2685
rect 4525 2635 4565 2665
rect 4525 2615 4535 2635
rect 4555 2615 4565 2635
rect 4525 2585 4565 2615
rect 4525 2565 4535 2585
rect 4555 2565 4565 2585
rect 4525 2535 4565 2565
rect 4525 2515 4535 2535
rect 4555 2515 4565 2535
rect 4525 2485 4565 2515
rect 4525 2465 4535 2485
rect 4555 2465 4565 2485
rect 4525 2435 4565 2465
rect 4525 2415 4535 2435
rect 4555 2415 4565 2435
rect 4525 2400 4565 2415
rect 4615 2685 4655 2700
rect 4615 2665 4625 2685
rect 4645 2665 4655 2685
rect 4615 2635 4655 2665
rect 4615 2615 4625 2635
rect 4645 2615 4655 2635
rect 4615 2585 4655 2615
rect 4615 2565 4625 2585
rect 4645 2565 4655 2585
rect 4615 2535 4655 2565
rect 4615 2515 4625 2535
rect 4645 2515 4655 2535
rect 4615 2485 4655 2515
rect 4615 2465 4625 2485
rect 4645 2465 4655 2485
rect 4615 2435 4655 2465
rect 4615 2415 4625 2435
rect 4645 2415 4655 2435
rect 4615 2400 4655 2415
rect 4705 2685 4745 2700
rect 4705 2665 4715 2685
rect 4735 2665 4745 2685
rect 4705 2635 4745 2665
rect 4705 2615 4715 2635
rect 4735 2615 4745 2635
rect 4705 2585 4745 2615
rect 4705 2565 4715 2585
rect 4735 2565 4745 2585
rect 4705 2535 4745 2565
rect 4705 2515 4715 2535
rect 4735 2515 4745 2535
rect 4705 2485 4745 2515
rect 4705 2465 4715 2485
rect 4735 2465 4745 2485
rect 4705 2435 4745 2465
rect 4705 2415 4715 2435
rect 4735 2415 4745 2435
rect 4705 2400 4745 2415
rect 4795 2685 4835 2700
rect 4795 2665 4805 2685
rect 4825 2665 4835 2685
rect 4795 2635 4835 2665
rect 4795 2615 4805 2635
rect 4825 2615 4835 2635
rect 4795 2585 4835 2615
rect 4795 2565 4805 2585
rect 4825 2565 4835 2585
rect 4795 2535 4835 2565
rect 4795 2515 4805 2535
rect 4825 2515 4835 2535
rect 4795 2485 4835 2515
rect 4795 2465 4805 2485
rect 4825 2465 4835 2485
rect 4795 2435 4835 2465
rect 4795 2415 4805 2435
rect 4825 2415 4835 2435
rect 4795 2400 4835 2415
rect 2565 1985 2605 2000
rect 2565 1965 2575 1985
rect 2595 1965 2605 1985
rect 2565 1935 2605 1965
rect 2565 1915 2575 1935
rect 2595 1915 2605 1935
rect 2565 1900 2605 1915
rect 2620 1985 2660 2000
rect 2620 1965 2630 1985
rect 2650 1965 2660 1985
rect 2620 1935 2660 1965
rect 2620 1915 2630 1935
rect 2650 1915 2660 1935
rect 2620 1900 2660 1915
rect 2675 1985 2715 2000
rect 2675 1965 2685 1985
rect 2705 1965 2715 1985
rect 2675 1935 2715 1965
rect 2675 1915 2685 1935
rect 2705 1915 2715 1935
rect 2675 1900 2715 1915
rect 2745 1985 2785 2000
rect 2745 1965 2755 1985
rect 2775 1965 2785 1985
rect 2745 1935 2785 1965
rect 2745 1915 2755 1935
rect 2775 1915 2785 1935
rect 2745 1900 2785 1915
rect 2805 1985 2845 2000
rect 2805 1965 2815 1985
rect 2835 1965 2845 1985
rect 2805 1935 2845 1965
rect 2805 1915 2815 1935
rect 2835 1915 2845 1935
rect 2805 1900 2845 1915
rect 2865 1985 2905 2000
rect 2865 1965 2875 1985
rect 2895 1965 2905 1985
rect 2865 1935 2905 1965
rect 2865 1915 2875 1935
rect 2895 1915 2905 1935
rect 2865 1900 2905 1915
rect 2925 1985 2965 2000
rect 2925 1965 2935 1985
rect 2955 1965 2965 1985
rect 2925 1935 2965 1965
rect 2925 1915 2935 1935
rect 2955 1915 2965 1935
rect 2925 1900 2965 1915
rect 2985 1985 3025 2000
rect 2985 1965 2995 1985
rect 3015 1965 3025 1985
rect 2985 1935 3025 1965
rect 2985 1915 2995 1935
rect 3015 1915 3025 1935
rect 2985 1900 3025 1915
rect 3045 1985 3085 2000
rect 3045 1965 3055 1985
rect 3075 1965 3085 1985
rect 3045 1935 3085 1965
rect 3045 1915 3055 1935
rect 3075 1915 3085 1935
rect 3045 1900 3085 1915
rect 3105 1985 3145 2000
rect 3105 1965 3115 1985
rect 3135 1965 3145 1985
rect 3105 1935 3145 1965
rect 3105 1915 3115 1935
rect 3135 1915 3145 1935
rect 3105 1900 3145 1915
rect 3165 1985 3205 2000
rect 3165 1965 3175 1985
rect 3195 1965 3205 1985
rect 3165 1935 3205 1965
rect 3165 1915 3175 1935
rect 3195 1915 3205 1935
rect 3165 1900 3205 1915
rect 3225 1985 3265 2000
rect 3225 1965 3235 1985
rect 3255 1965 3265 1985
rect 3225 1935 3265 1965
rect 3225 1915 3235 1935
rect 3255 1915 3265 1935
rect 3225 1900 3265 1915
rect 3285 1985 3325 2000
rect 3285 1965 3295 1985
rect 3315 1965 3325 1985
rect 3285 1935 3325 1965
rect 3285 1915 3295 1935
rect 3315 1915 3325 1935
rect 3285 1900 3325 1915
rect 3345 1985 3385 2000
rect 3345 1965 3355 1985
rect 3375 1965 3385 1985
rect 3345 1935 3385 1965
rect 3345 1915 3355 1935
rect 3375 1915 3385 1935
rect 3345 1900 3385 1915
rect 3405 1985 3445 2000
rect 3405 1965 3415 1985
rect 3435 1965 3445 1985
rect 3405 1935 3445 1965
rect 3405 1915 3415 1935
rect 3435 1915 3445 1935
rect 3405 1900 3445 1915
rect 3465 1985 3505 2000
rect 3465 1965 3475 1985
rect 3495 1965 3505 1985
rect 3465 1935 3505 1965
rect 3465 1915 3475 1935
rect 3495 1915 3505 1935
rect 3465 1900 3505 1915
rect 3525 1985 3565 2000
rect 3525 1965 3535 1985
rect 3555 1965 3565 1985
rect 3525 1935 3565 1965
rect 3525 1915 3535 1935
rect 3555 1915 3565 1935
rect 3525 1900 3565 1915
rect 3585 1985 3625 2000
rect 3585 1965 3595 1985
rect 3615 1965 3625 1985
rect 3585 1935 3625 1965
rect 3585 1915 3595 1935
rect 3615 1915 3625 1935
rect 3585 1900 3625 1915
rect 3645 1985 3685 2000
rect 3645 1965 3655 1985
rect 3675 1965 3685 1985
rect 3645 1935 3685 1965
rect 3645 1915 3655 1935
rect 3675 1915 3685 1935
rect 3645 1900 3685 1915
rect 3705 1985 3745 2000
rect 3705 1965 3715 1985
rect 3735 1965 3745 1985
rect 3705 1935 3745 1965
rect 3705 1915 3715 1935
rect 3735 1915 3745 1935
rect 3705 1900 3745 1915
rect 3765 1985 3805 2000
rect 3765 1965 3775 1985
rect 3795 1965 3805 1985
rect 3765 1935 3805 1965
rect 3765 1915 3775 1935
rect 3795 1915 3805 1935
rect 3765 1900 3805 1915
rect 3825 1985 3865 2000
rect 3825 1965 3835 1985
rect 3855 1965 3865 1985
rect 3825 1935 3865 1965
rect 3825 1915 3835 1935
rect 3855 1915 3865 1935
rect 3825 1900 3865 1915
rect 3885 1985 3925 2000
rect 3885 1965 3895 1985
rect 3915 1965 3925 1985
rect 3885 1935 3925 1965
rect 3885 1915 3895 1935
rect 3915 1915 3925 1935
rect 3885 1900 3925 1915
rect 3945 1985 3985 2000
rect 4025 1985 4065 2000
rect 3945 1965 3955 1985
rect 3975 1965 3985 1985
rect 4025 1965 4035 1985
rect 4055 1965 4065 1985
rect 3945 1935 3985 1965
rect 4025 1935 4065 1965
rect 3945 1915 3955 1935
rect 3975 1915 3985 1935
rect 4025 1915 4035 1935
rect 4055 1915 4065 1935
rect 3945 1900 3985 1915
rect 4025 1900 4065 1915
rect 4085 1985 4125 2000
rect 4085 1965 4095 1985
rect 4115 1965 4125 1985
rect 4085 1935 4125 1965
rect 4085 1915 4095 1935
rect 4115 1915 4125 1935
rect 4085 1900 4125 1915
rect 4145 1985 4185 2000
rect 4145 1965 4155 1985
rect 4175 1965 4185 1985
rect 4145 1935 4185 1965
rect 4145 1915 4155 1935
rect 4175 1915 4185 1935
rect 4145 1900 4185 1915
rect 4205 1985 4245 2000
rect 4205 1965 4215 1985
rect 4235 1965 4245 1985
rect 4205 1935 4245 1965
rect 4205 1915 4215 1935
rect 4235 1915 4245 1935
rect 4205 1900 4245 1915
rect 4265 1985 4305 2000
rect 4265 1965 4275 1985
rect 4295 1965 4305 1985
rect 4265 1935 4305 1965
rect 4265 1915 4275 1935
rect 4295 1915 4305 1935
rect 4265 1900 4305 1915
rect 4325 1985 4365 2000
rect 4325 1965 4335 1985
rect 4355 1965 4365 1985
rect 4325 1935 4365 1965
rect 4325 1915 4335 1935
rect 4355 1915 4365 1935
rect 4325 1900 4365 1915
rect 4385 1985 4425 2000
rect 4385 1965 4395 1985
rect 4415 1965 4425 1985
rect 4385 1935 4425 1965
rect 4385 1915 4395 1935
rect 4415 1915 4425 1935
rect 4385 1900 4425 1915
rect 4445 1985 4485 2000
rect 4445 1965 4455 1985
rect 4475 1965 4485 1985
rect 4445 1935 4485 1965
rect 4445 1915 4455 1935
rect 4475 1915 4485 1935
rect 4445 1900 4485 1915
rect 4505 1985 4545 2000
rect 4505 1965 4515 1985
rect 4535 1965 4545 1985
rect 4505 1935 4545 1965
rect 4505 1915 4515 1935
rect 4535 1915 4545 1935
rect 4505 1900 4545 1915
rect 4565 1985 4605 2000
rect 4565 1965 4575 1985
rect 4595 1965 4605 1985
rect 4565 1935 4605 1965
rect 4565 1915 4575 1935
rect 4595 1915 4605 1935
rect 4565 1900 4605 1915
rect 4625 1985 4665 2000
rect 4625 1965 4635 1985
rect 4655 1965 4665 1985
rect 4625 1935 4665 1965
rect 4625 1915 4635 1935
rect 4655 1915 4665 1935
rect 4625 1900 4665 1915
rect 4685 1985 4725 2000
rect 4685 1965 4695 1985
rect 4715 1965 4725 1985
rect 4685 1935 4725 1965
rect 4685 1915 4695 1935
rect 4715 1915 4725 1935
rect 4685 1900 4725 1915
rect 4745 1985 4785 2000
rect 4745 1965 4755 1985
rect 4775 1965 4785 1985
rect 4745 1935 4785 1965
rect 4745 1915 4755 1935
rect 4775 1915 4785 1935
rect 4745 1900 4785 1915
rect 4805 1985 4845 2000
rect 4805 1965 4815 1985
rect 4835 1965 4845 1985
rect 4805 1935 4845 1965
rect 4805 1915 4815 1935
rect 4835 1915 4845 1935
rect 4805 1900 4845 1915
rect 4865 1985 4905 2000
rect 4865 1965 4875 1985
rect 4895 1965 4905 1985
rect 4865 1935 4905 1965
rect 4865 1915 4875 1935
rect 4895 1915 4905 1935
rect 4865 1900 4905 1915
rect 4925 1985 4965 2000
rect 4925 1965 4935 1985
rect 4955 1965 4965 1985
rect 4925 1935 4965 1965
rect 4925 1915 4935 1935
rect 4955 1915 4965 1935
rect 4925 1900 4965 1915
rect 4985 1985 5025 2000
rect 4985 1965 4995 1985
rect 5015 1965 5025 1985
rect 4985 1935 5025 1965
rect 4985 1915 4995 1935
rect 5015 1915 5025 1935
rect 4985 1900 5025 1915
rect 5045 1985 5085 2000
rect 5045 1965 5055 1985
rect 5075 1965 5085 1985
rect 5045 1935 5085 1965
rect 5045 1915 5055 1935
rect 5075 1915 5085 1935
rect 5045 1900 5085 1915
rect 5105 1985 5145 2000
rect 5105 1965 5115 1985
rect 5135 1965 5145 1985
rect 5105 1935 5145 1965
rect 5105 1915 5115 1935
rect 5135 1915 5145 1935
rect 5105 1900 5145 1915
rect 5165 1985 5205 2000
rect 5165 1965 5175 1985
rect 5195 1965 5205 1985
rect 5165 1935 5205 1965
rect 5165 1915 5175 1935
rect 5195 1915 5205 1935
rect 5165 1900 5205 1915
rect 5225 1985 5265 2000
rect 5225 1965 5235 1985
rect 5255 1965 5265 1985
rect 5225 1935 5265 1965
rect 5225 1915 5235 1935
rect 5255 1915 5265 1935
rect 5225 1900 5265 1915
<< ndiffc >>
rect 11040 1680 11060 1700
rect 3175 1630 3195 1650
rect 3235 1630 3255 1650
rect 3295 1630 3315 1650
rect 3355 1630 3375 1650
rect 3415 1630 3435 1650
rect 3475 1630 3495 1650
rect 3535 1630 3555 1650
rect 3595 1630 3615 1650
rect 3655 1630 3675 1650
rect 3715 1630 3735 1650
rect 3775 1630 3795 1650
rect 4215 1630 4235 1650
rect 4275 1630 4295 1650
rect 4335 1630 4355 1650
rect 4395 1630 4415 1650
rect 4455 1630 4475 1650
rect 4515 1630 4535 1650
rect 4575 1630 4595 1650
rect 4635 1630 4655 1650
rect 4695 1630 4715 1650
rect 4755 1630 4775 1650
rect 4815 1630 4835 1650
rect 11040 1630 11060 1650
rect 11040 1580 11060 1600
rect 11095 1680 11115 1700
rect 11095 1630 11115 1650
rect 11095 1580 11115 1600
rect 11150 1680 11170 1700
rect 11150 1630 11170 1650
rect 11150 1580 11170 1600
rect 11205 1680 11225 1700
rect 11205 1630 11225 1650
rect 11205 1580 11225 1600
rect 11260 1680 11280 1700
rect 11260 1630 11280 1650
rect 11260 1580 11280 1600
rect 11315 1680 11335 1700
rect 11315 1630 11335 1650
rect 11315 1580 11335 1600
rect 11370 1680 11390 1700
rect 11370 1630 11390 1650
rect 11370 1580 11390 1600
rect 11425 1680 11445 1700
rect 11425 1630 11445 1650
rect 11425 1580 11445 1600
rect 11480 1680 11500 1700
rect 11480 1630 11500 1650
rect 11480 1580 11500 1600
rect 11535 1680 11555 1700
rect 11535 1630 11555 1650
rect 11535 1580 11555 1600
rect 11590 1680 11610 1700
rect 11590 1630 11610 1650
rect 11590 1580 11610 1600
rect 11645 1680 11665 1700
rect 11645 1630 11665 1650
rect 11645 1580 11665 1600
rect 11700 1680 11720 1700
rect 11780 1680 11800 1700
rect 11700 1630 11720 1650
rect 11780 1630 11800 1650
rect 11700 1580 11720 1600
rect 11780 1580 11800 1600
rect 11835 1680 11855 1700
rect 11835 1630 11855 1650
rect 11835 1580 11855 1600
rect 11890 1680 11910 1700
rect 11890 1630 11910 1650
rect 11890 1580 11910 1600
rect 11945 1680 11965 1700
rect 11945 1630 11965 1650
rect 11945 1580 11965 1600
rect 12000 1680 12020 1700
rect 12080 1680 12100 1700
rect 12000 1630 12020 1650
rect 12080 1630 12100 1650
rect 12000 1580 12020 1600
rect 12080 1580 12100 1600
rect 12135 1680 12155 1700
rect 12135 1630 12155 1650
rect 12135 1580 12155 1600
rect 12190 1680 12210 1700
rect 12190 1630 12210 1650
rect 12190 1580 12210 1600
rect 12245 1680 12265 1700
rect 12245 1630 12265 1650
rect 12245 1580 12265 1600
rect 12300 1680 12320 1700
rect 12300 1630 12320 1650
rect 12300 1580 12320 1600
rect 12355 1680 12375 1700
rect 12355 1630 12375 1650
rect 12355 1580 12375 1600
rect 12410 1680 12430 1700
rect 12410 1630 12430 1650
rect 12410 1580 12430 1600
rect 12465 1680 12485 1700
rect 12465 1630 12485 1650
rect 12465 1580 12485 1600
rect 12520 1680 12540 1700
rect 12520 1630 12540 1650
rect 12520 1580 12540 1600
rect 12575 1680 12595 1700
rect 12575 1630 12595 1650
rect 12575 1580 12595 1600
rect 12630 1680 12650 1700
rect 12630 1630 12650 1650
rect 12630 1580 12650 1600
rect 12685 1680 12705 1700
rect 12685 1630 12705 1650
rect 12685 1580 12705 1600
rect 12740 1680 12760 1700
rect 12740 1630 12760 1650
rect 12740 1580 12760 1600
rect 2845 1420 2865 1440
rect 2845 1370 2865 1390
rect 2845 1320 2865 1340
rect 2845 1270 2865 1290
rect 2845 1220 2865 1240
rect 3385 1420 3405 1440
rect 3385 1370 3405 1390
rect 3385 1320 3405 1340
rect 3385 1270 3405 1290
rect 3385 1220 3405 1240
rect 3925 1420 3945 1440
rect 3925 1370 3945 1390
rect 3925 1320 3945 1340
rect 3925 1270 3945 1290
rect 3925 1220 3945 1240
rect 4065 1420 4085 1440
rect 4065 1370 4085 1390
rect 4065 1320 4085 1340
rect 4065 1270 4085 1290
rect 4065 1220 4085 1240
rect 4605 1420 4625 1440
rect 4605 1370 4625 1390
rect 4605 1320 4625 1340
rect 4605 1270 4625 1290
rect 4605 1220 4625 1240
rect 5145 1420 5165 1440
rect 5145 1370 5165 1390
rect 5145 1320 5165 1340
rect 5145 1270 5165 1290
rect 5145 1220 5165 1240
rect 11215 1240 11235 1260
rect 11215 1190 11235 1210
rect 11215 1140 11235 1160
rect 11215 1090 11235 1110
rect 2955 1040 2975 1060
rect 2955 990 2975 1010
rect 3995 1040 4015 1060
rect 3995 990 4015 1010
rect 5035 1040 5055 1060
rect 11215 1040 11235 1060
rect 11270 1240 11290 1260
rect 11270 1190 11290 1210
rect 11270 1140 11290 1160
rect 11270 1090 11290 1110
rect 11270 1040 11290 1060
rect 11325 1240 11345 1260
rect 11325 1190 11345 1210
rect 11325 1140 11345 1160
rect 11325 1090 11345 1110
rect 11325 1040 11345 1060
rect 11380 1240 11400 1260
rect 11380 1190 11400 1210
rect 11380 1140 11400 1160
rect 11380 1090 11400 1110
rect 11380 1040 11400 1060
rect 11435 1240 11455 1260
rect 11435 1190 11455 1210
rect 11435 1140 11455 1160
rect 11435 1090 11455 1110
rect 11435 1040 11455 1060
rect 11490 1240 11510 1260
rect 11490 1190 11510 1210
rect 11490 1140 11510 1160
rect 11490 1090 11510 1110
rect 11490 1040 11510 1060
rect 11545 1240 11565 1260
rect 11545 1190 11565 1210
rect 11545 1140 11565 1160
rect 11545 1090 11565 1110
rect 11545 1040 11565 1060
rect 11600 1240 11620 1260
rect 11600 1190 11620 1210
rect 11600 1140 11620 1160
rect 11600 1090 11620 1110
rect 11600 1040 11620 1060
rect 11655 1240 11675 1260
rect 11655 1190 11675 1210
rect 11655 1140 11675 1160
rect 11655 1090 11675 1110
rect 11655 1040 11675 1060
rect 11710 1240 11730 1260
rect 11710 1190 11730 1210
rect 11710 1140 11730 1160
rect 11710 1090 11730 1110
rect 11710 1040 11730 1060
rect 11765 1240 11785 1260
rect 11765 1190 11785 1210
rect 11765 1140 11785 1160
rect 11765 1090 11785 1110
rect 11765 1040 11785 1060
rect 11820 1240 11840 1260
rect 11820 1190 11840 1210
rect 11820 1140 11840 1160
rect 11820 1090 11840 1110
rect 11820 1040 11840 1060
rect 11875 1240 11895 1260
rect 11875 1190 11895 1210
rect 11875 1140 11895 1160
rect 11875 1090 11895 1110
rect 11875 1040 11895 1060
rect 11930 1240 11950 1260
rect 11930 1190 11950 1210
rect 11930 1140 11950 1160
rect 11930 1090 11950 1110
rect 11930 1040 11950 1060
rect 11985 1240 12005 1260
rect 11985 1190 12005 1210
rect 11985 1140 12005 1160
rect 11985 1090 12005 1110
rect 11985 1040 12005 1060
rect 12040 1240 12060 1260
rect 12040 1190 12060 1210
rect 12040 1140 12060 1160
rect 12040 1090 12060 1110
rect 12040 1040 12060 1060
rect 12095 1240 12115 1260
rect 12095 1190 12115 1210
rect 12095 1140 12115 1160
rect 12095 1090 12115 1110
rect 12095 1040 12115 1060
rect 12150 1240 12170 1260
rect 12150 1190 12170 1210
rect 12150 1140 12170 1160
rect 12150 1090 12170 1110
rect 12150 1040 12170 1060
rect 12205 1240 12225 1260
rect 12205 1190 12225 1210
rect 12205 1140 12225 1160
rect 12205 1090 12225 1110
rect 12205 1040 12225 1060
rect 12260 1240 12280 1260
rect 12260 1190 12280 1210
rect 12260 1140 12280 1160
rect 12260 1090 12280 1110
rect 12260 1040 12280 1060
rect 12315 1240 12335 1260
rect 12315 1190 12335 1210
rect 12315 1140 12335 1160
rect 12315 1090 12335 1110
rect 12315 1040 12335 1060
rect 12370 1240 12390 1260
rect 12370 1190 12390 1210
rect 12370 1140 12390 1160
rect 12370 1090 12390 1110
rect 12370 1040 12390 1060
rect 12425 1240 12445 1260
rect 12425 1190 12445 1210
rect 12425 1140 12445 1160
rect 12425 1090 12445 1110
rect 12425 1040 12445 1060
rect 12480 1240 12500 1260
rect 12480 1190 12500 1210
rect 12480 1140 12500 1160
rect 12480 1090 12500 1110
rect 12480 1040 12500 1060
rect 12535 1240 12555 1260
rect 12535 1190 12555 1210
rect 12535 1140 12555 1160
rect 12535 1090 12555 1110
rect 12535 1040 12555 1060
rect 12590 1240 12610 1260
rect 12590 1190 12610 1210
rect 12590 1140 12610 1160
rect 12590 1090 12610 1110
rect 12590 1040 12610 1060
rect 5035 990 5055 1010
rect 3005 845 3025 865
rect 3005 795 3025 815
rect 3095 845 3115 865
rect 3095 795 3115 815
rect 3185 845 3205 865
rect 3185 795 3205 815
rect 3275 845 3295 865
rect 3275 795 3295 815
rect 3365 845 3385 865
rect 3365 795 3385 815
rect 3455 845 3475 865
rect 3455 795 3475 815
rect 3545 845 3565 865
rect 3545 795 3565 815
rect 3635 845 3655 865
rect 3635 795 3655 815
rect 3725 845 3745 865
rect 3725 795 3745 815
rect 3815 845 3835 865
rect 3815 795 3835 815
rect 3905 845 3925 865
rect 3905 795 3925 815
rect 3995 845 4015 865
rect 3995 795 4015 815
rect 4085 845 4105 865
rect 4085 795 4105 815
rect 4175 845 4195 865
rect 4175 795 4195 815
rect 4265 845 4285 865
rect 4265 795 4285 815
rect 4355 845 4375 865
rect 4355 795 4375 815
rect 4445 845 4465 865
rect 4445 795 4465 815
rect 4535 845 4555 865
rect 4535 795 4555 815
rect 4625 845 4645 865
rect 4625 795 4645 815
rect 4715 845 4735 865
rect 4715 795 4735 815
rect 4805 845 4825 865
rect 4805 795 4825 815
rect 4895 845 4915 865
rect 4895 795 4915 815
rect 4985 845 5005 865
rect 4985 795 5005 815
<< pdiffc >>
rect 3005 2895 3025 2915
rect 3005 2845 3025 2865
rect 3095 2895 3115 2915
rect 3095 2845 3115 2865
rect 3185 2895 3205 2915
rect 3185 2845 3205 2865
rect 3275 2895 3295 2915
rect 3275 2845 3295 2865
rect 3365 2895 3385 2915
rect 3365 2845 3385 2865
rect 3455 2895 3475 2915
rect 3455 2845 3475 2865
rect 3545 2895 3565 2915
rect 3545 2845 3565 2865
rect 3635 2895 3655 2915
rect 3635 2845 3655 2865
rect 3725 2895 3745 2915
rect 3725 2845 3745 2865
rect 3815 2895 3835 2915
rect 3815 2845 3835 2865
rect 3905 2895 3925 2915
rect 3905 2845 3925 2865
rect 3995 2895 4015 2915
rect 3995 2845 4015 2865
rect 4085 2895 4105 2915
rect 4085 2845 4105 2865
rect 4175 2895 4195 2915
rect 4175 2845 4195 2865
rect 4265 2895 4285 2915
rect 4265 2845 4285 2865
rect 4355 2895 4375 2915
rect 4355 2845 4375 2865
rect 4445 2895 4465 2915
rect 4445 2845 4465 2865
rect 4535 2895 4555 2915
rect 4535 2845 4555 2865
rect 4625 2895 4645 2915
rect 4625 2845 4645 2865
rect 4715 2895 4735 2915
rect 4715 2845 4735 2865
rect 4805 2895 4825 2915
rect 4805 2845 4825 2865
rect 4895 2895 4915 2915
rect 4895 2845 4915 2865
rect 4985 2895 5005 2915
rect 4985 2845 5005 2865
rect 3185 2665 3205 2685
rect 3185 2615 3205 2635
rect 3185 2565 3205 2585
rect 3185 2515 3205 2535
rect 3185 2465 3205 2485
rect 3185 2415 3205 2435
rect 3275 2665 3295 2685
rect 3275 2615 3295 2635
rect 3275 2565 3295 2585
rect 3275 2515 3295 2535
rect 3275 2465 3295 2485
rect 3275 2415 3295 2435
rect 3365 2665 3385 2685
rect 3365 2615 3385 2635
rect 3365 2565 3385 2585
rect 3365 2515 3385 2535
rect 3365 2465 3385 2485
rect 3365 2415 3385 2435
rect 3455 2665 3475 2685
rect 3455 2615 3475 2635
rect 3455 2565 3475 2585
rect 3455 2515 3475 2535
rect 3455 2465 3475 2485
rect 3455 2415 3475 2435
rect 3545 2665 3565 2685
rect 3545 2615 3565 2635
rect 3545 2565 3565 2585
rect 3545 2515 3565 2535
rect 3545 2465 3565 2485
rect 3545 2415 3565 2435
rect 3635 2665 3655 2685
rect 3635 2615 3655 2635
rect 3635 2565 3655 2585
rect 3635 2515 3655 2535
rect 3635 2465 3655 2485
rect 3635 2415 3655 2435
rect 3725 2665 3745 2685
rect 3725 2615 3745 2635
rect 3725 2565 3745 2585
rect 3725 2515 3745 2535
rect 3725 2465 3745 2485
rect 3725 2415 3745 2435
rect 3815 2665 3835 2685
rect 3815 2615 3835 2635
rect 3815 2565 3835 2585
rect 3815 2515 3835 2535
rect 3815 2465 3835 2485
rect 3815 2415 3835 2435
rect 3905 2665 3925 2685
rect 3905 2615 3925 2635
rect 3905 2565 3925 2585
rect 3905 2515 3925 2535
rect 3905 2465 3925 2485
rect 3905 2415 3925 2435
rect 3995 2665 4015 2685
rect 3995 2615 4015 2635
rect 3995 2565 4015 2585
rect 3995 2515 4015 2535
rect 3995 2465 4015 2485
rect 3995 2415 4015 2435
rect 4085 2665 4105 2685
rect 4085 2615 4105 2635
rect 4085 2565 4105 2585
rect 4085 2515 4105 2535
rect 4085 2465 4105 2485
rect 4085 2415 4105 2435
rect 4175 2665 4195 2685
rect 4175 2615 4195 2635
rect 4175 2565 4195 2585
rect 4175 2515 4195 2535
rect 4175 2465 4195 2485
rect 4175 2415 4195 2435
rect 4265 2665 4285 2685
rect 4265 2615 4285 2635
rect 4265 2565 4285 2585
rect 4265 2515 4285 2535
rect 4265 2465 4285 2485
rect 4265 2415 4285 2435
rect 4355 2665 4375 2685
rect 4355 2615 4375 2635
rect 4355 2565 4375 2585
rect 4355 2515 4375 2535
rect 4355 2465 4375 2485
rect 4355 2415 4375 2435
rect 4445 2665 4465 2685
rect 4445 2615 4465 2635
rect 4445 2565 4465 2585
rect 4445 2515 4465 2535
rect 4445 2465 4465 2485
rect 4445 2415 4465 2435
rect 4535 2665 4555 2685
rect 4535 2615 4555 2635
rect 4535 2565 4555 2585
rect 4535 2515 4555 2535
rect 4535 2465 4555 2485
rect 4535 2415 4555 2435
rect 4625 2665 4645 2685
rect 4625 2615 4645 2635
rect 4625 2565 4645 2585
rect 4625 2515 4645 2535
rect 4625 2465 4645 2485
rect 4625 2415 4645 2435
rect 4715 2665 4735 2685
rect 4715 2615 4735 2635
rect 4715 2565 4735 2585
rect 4715 2515 4735 2535
rect 4715 2465 4735 2485
rect 4715 2415 4735 2435
rect 4805 2665 4825 2685
rect 4805 2615 4825 2635
rect 4805 2565 4825 2585
rect 4805 2515 4825 2535
rect 4805 2465 4825 2485
rect 4805 2415 4825 2435
rect 2575 1965 2595 1985
rect 2575 1915 2595 1935
rect 2630 1965 2650 1985
rect 2630 1915 2650 1935
rect 2685 1965 2705 1985
rect 2685 1915 2705 1935
rect 2755 1965 2775 1985
rect 2755 1915 2775 1935
rect 2815 1965 2835 1985
rect 2815 1915 2835 1935
rect 2875 1965 2895 1985
rect 2875 1915 2895 1935
rect 2935 1965 2955 1985
rect 2935 1915 2955 1935
rect 2995 1965 3015 1985
rect 2995 1915 3015 1935
rect 3055 1965 3075 1985
rect 3055 1915 3075 1935
rect 3115 1965 3135 1985
rect 3115 1915 3135 1935
rect 3175 1965 3195 1985
rect 3175 1915 3195 1935
rect 3235 1965 3255 1985
rect 3235 1915 3255 1935
rect 3295 1965 3315 1985
rect 3295 1915 3315 1935
rect 3355 1965 3375 1985
rect 3355 1915 3375 1935
rect 3415 1965 3435 1985
rect 3415 1915 3435 1935
rect 3475 1965 3495 1985
rect 3475 1915 3495 1935
rect 3535 1965 3555 1985
rect 3535 1915 3555 1935
rect 3595 1965 3615 1985
rect 3595 1915 3615 1935
rect 3655 1965 3675 1985
rect 3655 1915 3675 1935
rect 3715 1965 3735 1985
rect 3715 1915 3735 1935
rect 3775 1965 3795 1985
rect 3775 1915 3795 1935
rect 3835 1965 3855 1985
rect 3835 1915 3855 1935
rect 3895 1965 3915 1985
rect 3895 1915 3915 1935
rect 3955 1965 3975 1985
rect 4035 1965 4055 1985
rect 3955 1915 3975 1935
rect 4035 1915 4055 1935
rect 4095 1965 4115 1985
rect 4095 1915 4115 1935
rect 4155 1965 4175 1985
rect 4155 1915 4175 1935
rect 4215 1965 4235 1985
rect 4215 1915 4235 1935
rect 4275 1965 4295 1985
rect 4275 1915 4295 1935
rect 4335 1965 4355 1985
rect 4335 1915 4355 1935
rect 4395 1965 4415 1985
rect 4395 1915 4415 1935
rect 4455 1965 4475 1985
rect 4455 1915 4475 1935
rect 4515 1965 4535 1985
rect 4515 1915 4535 1935
rect 4575 1965 4595 1985
rect 4575 1915 4595 1935
rect 4635 1965 4655 1985
rect 4635 1915 4655 1935
rect 4695 1965 4715 1985
rect 4695 1915 4715 1935
rect 4755 1965 4775 1985
rect 4755 1915 4775 1935
rect 4815 1965 4835 1985
rect 4815 1915 4835 1935
rect 4875 1965 4895 1985
rect 4875 1915 4895 1935
rect 4935 1965 4955 1985
rect 4935 1915 4955 1935
rect 4995 1965 5015 1985
rect 4995 1915 5015 1935
rect 5055 1965 5075 1985
rect 5055 1915 5075 1935
rect 5115 1965 5135 1985
rect 5115 1915 5135 1935
rect 5175 1965 5195 1985
rect 5175 1915 5195 1935
rect 5235 1965 5255 1985
rect 5235 1915 5255 1935
<< psubdiff >>
rect 905 2910 1125 2920
rect 905 2880 920 2910
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1125 2910
rect 905 2870 1125 2880
rect -50 1715 100 1730
rect -50 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 100 1715
rect -50 1680 100 1695
rect 10990 1700 11030 1715
rect 10990 1680 11000 1700
rect 11020 1680 11030 1700
rect 3980 1650 4030 1665
rect 3980 1630 3995 1650
rect 4015 1630 4030 1650
rect 3980 1615 4030 1630
rect 10990 1650 11030 1680
rect 10990 1630 11000 1650
rect 11020 1630 11030 1650
rect 10990 1600 11030 1630
rect 10990 1580 11000 1600
rect 11020 1580 11030 1600
rect 10990 1565 11030 1580
rect 11730 1700 11770 1715
rect 11730 1680 11740 1700
rect 11760 1680 11770 1700
rect 11730 1650 11770 1680
rect 11730 1630 11740 1650
rect 11760 1630 11770 1650
rect 11730 1600 11770 1630
rect 11730 1580 11740 1600
rect 11760 1580 11770 1600
rect 11730 1565 11770 1580
rect 12030 1700 12070 1715
rect 12030 1680 12040 1700
rect 12060 1680 12070 1700
rect 12030 1650 12070 1680
rect 12030 1630 12040 1650
rect 12060 1630 12070 1650
rect 12030 1600 12070 1630
rect 12030 1580 12040 1600
rect 12060 1580 12070 1600
rect 12030 1565 12070 1580
rect 12770 1700 12810 1715
rect 12770 1680 12780 1700
rect 12800 1680 12810 1700
rect 12770 1650 12810 1680
rect 12770 1630 12780 1650
rect 12800 1630 12810 1650
rect 12770 1600 12810 1630
rect 12770 1580 12780 1600
rect 12800 1580 12810 1600
rect 12770 1565 12810 1580
rect 11165 1260 11205 1275
rect 11165 1240 11175 1260
rect 11195 1240 11205 1260
rect 11165 1210 11205 1240
rect 11165 1190 11175 1210
rect 11195 1190 11205 1210
rect 11165 1160 11205 1190
rect 11165 1140 11175 1160
rect 11195 1140 11205 1160
rect 11165 1110 11205 1140
rect 11165 1090 11175 1110
rect 11195 1090 11205 1110
rect 5065 1060 5105 1075
rect 5065 1040 5075 1060
rect 5095 1040 5105 1060
rect 5065 1010 5105 1040
rect 11165 1060 11205 1090
rect 11165 1040 11175 1060
rect 11195 1040 11205 1060
rect 11165 1025 11205 1040
rect 12620 1260 12660 1275
rect 12620 1240 12630 1260
rect 12650 1240 12660 1260
rect 12620 1210 12660 1240
rect 12620 1190 12630 1210
rect 12650 1190 12660 1210
rect 12620 1160 12660 1190
rect 12620 1140 12630 1160
rect 12650 1140 12660 1160
rect 12620 1110 12660 1140
rect 12620 1090 12630 1110
rect 12650 1090 12660 1110
rect 12620 1060 12660 1090
rect 12620 1040 12630 1060
rect 12650 1040 12660 1060
rect 12620 1025 12660 1040
rect 5065 990 5075 1010
rect 5095 990 5105 1010
rect 5065 975 5105 990
rect 2955 865 2995 880
rect 2955 845 2965 865
rect 2985 845 2995 865
rect 2955 815 2995 845
rect 2955 795 2965 815
rect 2985 795 2995 815
rect 2955 780 2995 795
rect 5015 865 5055 880
rect 5015 845 5025 865
rect 5045 845 5055 865
rect 5015 815 5055 845
rect 5015 795 5025 815
rect 5045 795 5055 815
rect 5015 780 5055 795
<< nsubdiff >>
rect 2955 2915 2995 2930
rect 2955 2895 2965 2915
rect 2985 2895 2995 2915
rect 2955 2865 2995 2895
rect 2955 2845 2965 2865
rect 2985 2845 2995 2865
rect 2955 2830 2995 2845
rect 5015 2915 5055 2930
rect 5015 2895 5025 2915
rect 5045 2895 5055 2915
rect 5015 2865 5055 2895
rect 5015 2845 5025 2865
rect 5045 2845 5055 2865
rect 5015 2830 5055 2845
rect 3135 2685 3175 2700
rect 3135 2665 3145 2685
rect 3165 2665 3175 2685
rect 3135 2635 3175 2665
rect 3135 2615 3145 2635
rect 3165 2615 3175 2635
rect 3135 2585 3175 2615
rect 3135 2565 3145 2585
rect 3165 2565 3175 2585
rect 3135 2535 3175 2565
rect 3135 2515 3145 2535
rect 3165 2515 3175 2535
rect 3135 2485 3175 2515
rect 3135 2465 3145 2485
rect 3165 2465 3175 2485
rect 3135 2435 3175 2465
rect 3135 2415 3145 2435
rect 3165 2415 3175 2435
rect 3135 2400 3175 2415
rect 4835 2685 4875 2700
rect 4835 2665 4845 2685
rect 4865 2665 4875 2685
rect 4835 2635 4875 2665
rect 4835 2615 4845 2635
rect 4865 2615 4875 2635
rect 4835 2585 4875 2615
rect 4835 2565 4845 2585
rect 4865 2565 4875 2585
rect 4835 2535 4875 2565
rect 4835 2515 4845 2535
rect 4865 2515 4875 2535
rect 4835 2485 4875 2515
rect 4835 2465 4845 2485
rect 4865 2465 4875 2485
rect 4835 2435 4875 2465
rect 4835 2415 4845 2435
rect 4865 2415 4875 2435
rect 4835 2400 4875 2415
rect 3985 1985 4025 2000
rect 3985 1965 3995 1985
rect 4015 1965 4025 1985
rect 3985 1935 4025 1965
rect 3985 1915 3995 1935
rect 4015 1915 4025 1935
rect 3985 1900 4025 1915
<< psubdiffcont >>
rect 920 2880 950 2910
rect 1000 2880 1030 2910
rect 1080 2880 1110 2910
rect -35 1695 -15 1715
rect 15 1695 35 1715
rect 65 1695 85 1715
rect 11000 1680 11020 1700
rect 3995 1630 4015 1650
rect 11000 1630 11020 1650
rect 11000 1580 11020 1600
rect 11740 1680 11760 1700
rect 11740 1630 11760 1650
rect 11740 1580 11760 1600
rect 12040 1680 12060 1700
rect 12040 1630 12060 1650
rect 12040 1580 12060 1600
rect 12780 1680 12800 1700
rect 12780 1630 12800 1650
rect 12780 1580 12800 1600
rect 11175 1240 11195 1260
rect 11175 1190 11195 1210
rect 11175 1140 11195 1160
rect 11175 1090 11195 1110
rect 5075 1040 5095 1060
rect 11175 1040 11195 1060
rect 12630 1240 12650 1260
rect 12630 1190 12650 1210
rect 12630 1140 12650 1160
rect 12630 1090 12650 1110
rect 12630 1040 12650 1060
rect 5075 990 5095 1010
rect 2965 845 2985 865
rect 2965 795 2985 815
rect 5025 845 5045 865
rect 5025 795 5045 815
<< nsubdiffcont >>
rect 2965 2895 2985 2915
rect 2965 2845 2985 2865
rect 5025 2895 5045 2915
rect 5025 2845 5045 2865
rect 3145 2665 3165 2685
rect 3145 2615 3165 2635
rect 3145 2565 3165 2585
rect 3145 2515 3165 2535
rect 3145 2465 3165 2485
rect 3145 2415 3165 2435
rect 4845 2665 4865 2685
rect 4845 2615 4865 2635
rect 4845 2565 4865 2585
rect 4845 2515 4865 2535
rect 4845 2465 4865 2485
rect 4845 2415 4865 2435
rect 3995 1965 4015 1985
rect 3995 1915 4015 1935
<< poly >>
rect 3140 2975 3175 2985
rect 3140 2955 3145 2975
rect 3165 2955 3175 2975
rect 3140 2945 3175 2955
rect 4835 2975 4870 2985
rect 4835 2955 4845 2975
rect 4865 2955 4870 2975
rect 4835 2945 4870 2955
rect 3035 2930 3085 2945
rect 3125 2930 3175 2945
rect 3215 2930 3265 2945
rect 3305 2930 3355 2945
rect 3395 2930 3445 2945
rect 3485 2930 3535 2945
rect 3575 2930 3625 2945
rect 3665 2930 3715 2945
rect 3755 2930 3805 2945
rect 3845 2930 3895 2945
rect 3935 2930 3985 2945
rect 4025 2930 4075 2945
rect 4115 2930 4165 2945
rect 4205 2930 4255 2945
rect 4295 2930 4345 2945
rect 4385 2930 4435 2945
rect 4475 2930 4525 2945
rect 4565 2930 4615 2945
rect 4655 2930 4705 2945
rect 4745 2930 4795 2945
rect 4835 2930 4885 2945
rect 4925 2930 4975 2945
rect 3035 2815 3085 2830
rect 2995 2805 3085 2815
rect 3125 2820 3175 2830
rect 3215 2820 3265 2830
rect 3305 2820 3355 2830
rect 3395 2820 3445 2830
rect 3485 2820 3535 2830
rect 3575 2820 3625 2830
rect 3665 2820 3715 2830
rect 3755 2820 3805 2830
rect 3845 2820 3895 2830
rect 3935 2820 3985 2830
rect 4025 2820 4075 2830
rect 4115 2820 4165 2830
rect 4205 2820 4255 2830
rect 4295 2820 4345 2830
rect 4385 2820 4435 2830
rect 4475 2820 4525 2830
rect 4565 2820 4615 2830
rect 4655 2820 4705 2830
rect 4745 2820 4795 2830
rect 4835 2820 4885 2830
rect 3125 2805 4885 2820
rect 4925 2815 4975 2830
rect 4925 2805 5015 2815
rect 2995 2785 3005 2805
rect 3025 2800 3085 2805
rect 4925 2800 4985 2805
rect 3025 2785 3035 2800
rect 2995 2775 3035 2785
rect 4975 2785 4985 2800
rect 5005 2785 5015 2805
rect 4975 2775 5015 2785
rect 3175 2745 3215 2755
rect 3175 2725 3185 2745
rect 3205 2730 3215 2745
rect 4795 2745 4835 2755
rect 4795 2730 4805 2745
rect 3205 2725 3265 2730
rect 3175 2715 3265 2725
rect 4745 2725 4805 2730
rect 4825 2725 4835 2745
rect 4745 2715 4835 2725
rect 3215 2700 3265 2715
rect 3305 2700 3355 2715
rect 3395 2700 3445 2715
rect 3485 2700 3535 2715
rect 3575 2700 3625 2715
rect 3665 2700 3715 2715
rect 3755 2700 3805 2715
rect 3845 2700 3895 2715
rect 3935 2700 3985 2715
rect 4025 2700 4075 2715
rect 4115 2700 4165 2715
rect 4205 2700 4255 2715
rect 4295 2700 4345 2715
rect 4385 2700 4435 2715
rect 4475 2700 4525 2715
rect 4565 2700 4615 2715
rect 4655 2700 4705 2715
rect 4745 2700 4795 2715
rect 3215 2385 3265 2400
rect 3305 2390 3355 2400
rect 3395 2390 3445 2400
rect 3485 2390 3535 2400
rect 3575 2390 3625 2400
rect 3665 2390 3715 2400
rect 3755 2390 3805 2400
rect 3845 2390 3895 2400
rect 3935 2390 3985 2400
rect 4025 2390 4075 2400
rect 4115 2390 4165 2400
rect 4205 2390 4255 2400
rect 4295 2390 4345 2400
rect 4385 2390 4435 2400
rect 4475 2390 4525 2400
rect 4565 2390 4615 2400
rect 4655 2390 4705 2400
rect 3305 2375 4705 2390
rect 4745 2385 4795 2400
rect 3355 2370 3395 2375
rect 3355 2350 3365 2370
rect 3385 2350 3395 2370
rect 3355 2340 3395 2350
rect 3885 2355 3895 2375
rect 3915 2355 3925 2375
rect 3885 2345 3925 2355
rect 2605 2000 2620 2015
rect 2660 2000 2675 2015
rect 2785 2000 2805 2015
rect 2845 2000 2865 2015
rect 2905 2000 2925 2015
rect 2965 2000 2985 2015
rect 3025 2000 3045 2015
rect 3085 2000 3105 2015
rect 3145 2000 3165 2015
rect 3205 2000 3225 2015
rect 3265 2000 3285 2015
rect 3325 2000 3345 2015
rect 3385 2000 3405 2015
rect 3445 2000 3465 2015
rect 3505 2000 3525 2015
rect 3565 2000 3585 2015
rect 3625 2000 3645 2015
rect 3685 2000 3705 2015
rect 3745 2000 3765 2015
rect 3805 2000 3825 2015
rect 3865 2000 3885 2015
rect 3925 2000 3945 2015
rect 4065 2000 4085 2015
rect 4125 2000 4145 2015
rect 4185 2000 4205 2015
rect 4245 2000 4265 2015
rect 4305 2000 4325 2015
rect 4365 2000 4385 2015
rect 4425 2000 4445 2015
rect 4485 2000 4505 2015
rect 4545 2000 4565 2015
rect 4605 2000 4625 2015
rect 4665 2000 4685 2015
rect 4725 2000 4745 2015
rect 4785 2000 4805 2015
rect 4845 2000 4865 2015
rect 4905 2000 4925 2015
rect 4965 2000 4985 2015
rect 5025 2000 5045 2015
rect 5085 2000 5105 2015
rect 5145 2000 5165 2015
rect 5205 2000 5225 2015
rect 2605 1890 2620 1900
rect 2660 1890 2675 1900
rect 2605 1875 2675 1890
rect 2785 1885 2805 1900
rect 2845 1885 2865 1900
rect 2905 1890 2925 1900
rect 2965 1890 2985 1900
rect 3025 1890 3045 1900
rect 3085 1890 3105 1900
rect 2765 1875 2805 1885
rect 2620 1855 2630 1875
rect 2650 1855 2660 1875
rect 2620 1845 2660 1855
rect 2765 1855 2775 1875
rect 2795 1855 2805 1875
rect 2765 1845 2805 1855
rect 2835 1875 2875 1885
rect 2905 1875 3105 1890
rect 3145 1890 3165 1900
rect 3205 1890 3225 1900
rect 3145 1875 3225 1890
rect 3265 1890 3285 1900
rect 3325 1890 3345 1900
rect 3385 1890 3405 1900
rect 3445 1890 3465 1900
rect 3265 1875 3465 1890
rect 3505 1890 3525 1900
rect 3565 1890 3585 1900
rect 3505 1875 3585 1890
rect 3625 1890 3645 1900
rect 3685 1890 3705 1900
rect 3745 1890 3765 1900
rect 3805 1890 3825 1900
rect 3625 1875 3825 1890
rect 3865 1885 3885 1900
rect 3925 1890 3945 1900
rect 4065 1890 4085 1900
rect 3855 1875 3895 1885
rect 3925 1875 4085 1890
rect 4125 1885 4145 1900
rect 4185 1890 4205 1900
rect 4245 1890 4265 1900
rect 4305 1890 4325 1900
rect 4365 1890 4385 1900
rect 4115 1875 4155 1885
rect 4185 1875 4385 1890
rect 4425 1890 4445 1900
rect 4485 1890 4505 1900
rect 4425 1875 4505 1890
rect 4545 1890 4565 1900
rect 4605 1890 4625 1900
rect 4665 1890 4685 1900
rect 4725 1890 4745 1900
rect 4545 1875 4745 1890
rect 4785 1890 4805 1900
rect 4845 1890 4865 1900
rect 4785 1875 4865 1890
rect 4905 1890 4925 1900
rect 4965 1890 4985 1900
rect 5025 1890 5045 1900
rect 5085 1890 5105 1900
rect 4905 1875 5105 1890
rect 5145 1885 5165 1900
rect 5205 1885 5225 1900
rect 5135 1875 5175 1885
rect 2835 1855 2845 1875
rect 2865 1855 2875 1875
rect 2835 1845 2875 1855
rect 2925 1855 2935 1875
rect 2955 1855 2965 1875
rect 2925 1845 2965 1855
rect 3165 1855 3175 1875
rect 3195 1855 3205 1875
rect 3165 1845 3205 1855
rect 3285 1855 3295 1875
rect 3315 1855 3325 1875
rect 3285 1845 3325 1855
rect 3525 1855 3535 1875
rect 3555 1855 3565 1875
rect 3525 1845 3565 1855
rect 3645 1855 3655 1875
rect 3675 1855 3685 1875
rect 3645 1845 3685 1855
rect 3855 1855 3865 1875
rect 3885 1855 3895 1875
rect 3855 1845 3895 1855
rect 3985 1870 4025 1875
rect 3985 1850 3995 1870
rect 4015 1850 4025 1870
rect 3985 1840 4025 1850
rect 4115 1855 4125 1875
rect 4145 1855 4155 1875
rect 4115 1845 4155 1855
rect 4325 1855 4335 1875
rect 4355 1855 4365 1875
rect 4325 1845 4365 1855
rect 4445 1855 4455 1875
rect 4475 1855 4485 1875
rect 4445 1845 4485 1855
rect 4685 1855 4695 1875
rect 4715 1855 4725 1875
rect 4685 1845 4725 1855
rect 4805 1855 4815 1875
rect 4835 1855 4845 1875
rect 4805 1845 4845 1855
rect 5045 1855 5055 1875
rect 5075 1855 5085 1875
rect 5045 1845 5085 1855
rect 5135 1855 5145 1875
rect 5165 1855 5175 1875
rect 5135 1845 5175 1855
rect 5205 1875 5245 1885
rect 5205 1855 5215 1875
rect 5235 1855 5245 1875
rect 5205 1845 5245 1855
rect 3225 1755 3265 1765
rect 3225 1735 3235 1755
rect 3255 1735 3265 1755
rect 3225 1720 3265 1735
rect 4745 1755 4785 1765
rect 4745 1735 4755 1755
rect 4775 1735 4785 1755
rect 11237 1760 11269 1770
rect 11237 1740 11243 1760
rect 11260 1740 11269 1760
rect 11457 1760 11489 1770
rect 11457 1740 11463 1760
rect 11480 1740 11489 1760
rect 4745 1720 4785 1735
rect 11180 1730 11269 1740
rect 11400 1730 11489 1740
rect 11601 1760 11635 1770
rect 11601 1740 11610 1760
rect 11627 1740 11635 1760
rect 11867 1760 11899 1770
rect 11867 1745 11876 1760
rect 11601 1730 11635 1740
rect 11865 1740 11876 1745
rect 11893 1740 11899 1760
rect 12277 1760 12309 1770
rect 12277 1740 12283 1760
rect 12300 1740 12309 1760
rect 12497 1760 12529 1770
rect 12497 1740 12503 1760
rect 12520 1740 12529 1760
rect 11865 1730 11899 1740
rect 12220 1730 12309 1740
rect 12440 1730 12529 1740
rect 12641 1760 12675 1770
rect 12641 1740 12650 1760
rect 12667 1740 12675 1760
rect 12641 1730 12675 1740
rect 3225 1705 3765 1720
rect 3205 1665 3225 1680
rect 3265 1665 3285 1705
rect 3325 1665 3345 1705
rect 3385 1665 3405 1680
rect 3445 1665 3465 1680
rect 3505 1665 3525 1705
rect 3565 1665 3585 1705
rect 3625 1665 3645 1680
rect 3685 1665 3705 1680
rect 3745 1665 3765 1705
rect 4245 1705 4785 1720
rect 11070 1715 11085 1730
rect 11125 1715 11140 1730
rect 11180 1725 11250 1730
rect 11180 1715 11195 1725
rect 11235 1715 11250 1725
rect 11290 1715 11305 1730
rect 11345 1715 11360 1730
rect 11400 1725 11470 1730
rect 11400 1715 11415 1725
rect 11455 1715 11470 1725
rect 11510 1715 11525 1730
rect 11565 1715 11580 1730
rect 11620 1715 11635 1730
rect 11675 1715 11690 1730
rect 11810 1715 11825 1730
rect 11865 1715 11880 1730
rect 11920 1715 11935 1730
rect 11975 1715 11990 1730
rect 12110 1715 12125 1730
rect 12165 1715 12180 1730
rect 12220 1725 12290 1730
rect 12220 1715 12235 1725
rect 12275 1715 12290 1725
rect 12330 1715 12345 1730
rect 12385 1715 12400 1730
rect 12440 1725 12510 1730
rect 12440 1715 12455 1725
rect 12495 1715 12510 1725
rect 12550 1715 12565 1730
rect 12605 1715 12620 1730
rect 12660 1715 12675 1730
rect 12715 1715 12730 1730
rect 4245 1665 4265 1705
rect 4305 1665 4325 1680
rect 4365 1665 4385 1680
rect 4425 1665 4445 1705
rect 4485 1665 4505 1705
rect 4545 1665 4565 1680
rect 4605 1665 4625 1680
rect 4665 1665 4685 1705
rect 4725 1665 4745 1705
rect 4785 1665 4805 1680
rect 3205 1600 3225 1615
rect 3265 1600 3285 1615
rect 3325 1600 3345 1615
rect 3165 1590 3225 1600
rect 3165 1570 3175 1590
rect 3195 1575 3225 1590
rect 3385 1575 3405 1615
rect 3445 1575 3465 1615
rect 3505 1600 3525 1615
rect 3565 1600 3585 1615
rect 3625 1575 3645 1615
rect 3685 1575 3705 1615
rect 3745 1600 3765 1615
rect 4245 1600 4265 1615
rect 3195 1570 3705 1575
rect 3165 1560 3705 1570
rect 4305 1575 4325 1615
rect 4365 1575 4385 1615
rect 4425 1600 4445 1615
rect 4485 1600 4505 1615
rect 4545 1575 4565 1615
rect 4605 1575 4625 1615
rect 4665 1600 4685 1615
rect 4725 1600 4745 1615
rect 4785 1600 4805 1615
rect 4785 1590 4845 1600
rect 4785 1575 4815 1590
rect 4305 1570 4815 1575
rect 4835 1570 4845 1590
rect 4305 1560 4845 1570
rect 11070 1555 11085 1565
rect 10990 1540 11085 1555
rect 11125 1550 11140 1565
rect 11180 1550 11195 1565
rect 11235 1550 11250 1565
rect 11290 1555 11305 1565
rect 11345 1555 11360 1565
rect 11106 1540 11140 1550
rect 11290 1540 11360 1555
rect 11400 1550 11415 1565
rect 11455 1550 11470 1565
rect 11510 1555 11525 1565
rect 11565 1555 11580 1565
rect 11510 1540 11580 1555
rect 11620 1550 11635 1565
rect 11675 1555 11690 1565
rect 11810 1555 11825 1565
rect 11675 1540 11825 1555
rect 11865 1550 11880 1565
rect 11920 1550 11935 1565
rect 11975 1555 11990 1565
rect 12110 1555 12125 1565
rect 11920 1540 11954 1550
rect 11975 1540 12125 1555
rect 12165 1550 12180 1565
rect 12220 1550 12235 1565
rect 12275 1550 12290 1565
rect 12330 1555 12345 1565
rect 12385 1555 12400 1565
rect 12146 1540 12180 1550
rect 12330 1540 12400 1555
rect 12440 1550 12455 1565
rect 12495 1550 12510 1565
rect 12550 1555 12565 1565
rect 12605 1555 12620 1565
rect 12550 1540 12620 1555
rect 12660 1550 12675 1565
rect 12715 1555 12730 1565
rect 12715 1540 12810 1555
rect 10990 1520 11000 1540
rect 11020 1520 11030 1540
rect 10990 1510 11030 1520
rect 11106 1520 11112 1540
rect 11129 1520 11138 1540
rect 11106 1510 11138 1520
rect 11305 1520 11315 1540
rect 11335 1520 11345 1540
rect 11305 1510 11345 1520
rect 11525 1520 11535 1540
rect 11555 1520 11565 1540
rect 11525 1510 11565 1520
rect 11730 1520 11740 1540
rect 11760 1520 11770 1540
rect 11730 1510 11770 1520
rect 11922 1520 11928 1540
rect 11945 1520 11954 1540
rect 11922 1510 11954 1520
rect 12030 1520 12040 1540
rect 12060 1520 12070 1540
rect 12030 1510 12070 1520
rect 12146 1520 12152 1540
rect 12169 1520 12178 1540
rect 12146 1510 12178 1520
rect 12345 1520 12355 1540
rect 12375 1520 12385 1540
rect 12345 1510 12385 1520
rect 12565 1520 12575 1540
rect 12595 1520 12605 1540
rect 12565 1510 12605 1520
rect 12770 1520 12780 1540
rect 12800 1520 12810 1540
rect 12770 1510 12810 1520
rect 2925 1495 2965 1505
rect 2925 1475 2935 1495
rect 2955 1475 2965 1495
rect 2925 1470 2965 1475
rect 3045 1495 3085 1505
rect 3045 1475 3055 1495
rect 3075 1475 3085 1495
rect 3045 1470 3085 1475
rect 3165 1495 3205 1505
rect 3165 1475 3175 1495
rect 3195 1475 3205 1495
rect 3165 1470 3205 1475
rect 3285 1495 3325 1505
rect 3285 1475 3295 1495
rect 3315 1475 3325 1495
rect 3285 1470 3325 1475
rect 3525 1495 3565 1505
rect 3525 1475 3535 1495
rect 3555 1475 3565 1495
rect 3525 1470 3565 1475
rect 3645 1495 3685 1505
rect 3645 1475 3655 1495
rect 3675 1475 3685 1495
rect 3645 1470 3685 1475
rect 3765 1495 3805 1505
rect 3765 1475 3775 1495
rect 3795 1475 3805 1495
rect 3765 1470 3805 1475
rect 4205 1495 4245 1505
rect 4205 1475 4215 1495
rect 4235 1475 4245 1495
rect 4205 1470 4245 1475
rect 4325 1495 4365 1505
rect 4325 1475 4335 1495
rect 4355 1475 4365 1495
rect 4325 1470 4365 1475
rect 4445 1495 4485 1505
rect 4445 1475 4455 1495
rect 4475 1475 4485 1495
rect 4445 1470 4485 1475
rect 4685 1495 4725 1505
rect 4685 1475 4695 1495
rect 4715 1475 4725 1495
rect 4685 1470 4725 1475
rect 4805 1495 4845 1505
rect 4805 1475 4815 1495
rect 4835 1475 4845 1495
rect 4805 1470 4845 1475
rect 4925 1495 4965 1505
rect 4925 1475 4935 1495
rect 4955 1475 4965 1495
rect 4925 1470 4965 1475
rect 5045 1495 5085 1505
rect 5045 1475 5055 1495
rect 5075 1475 5085 1495
rect 5045 1470 5085 1475
rect 2875 1455 3375 1470
rect 3415 1455 3915 1470
rect 4095 1455 4595 1470
rect 4635 1455 5135 1470
rect 11815 1320 11845 1330
rect 11815 1300 11820 1320
rect 11840 1300 11845 1320
rect 12510 1315 12595 1330
rect 11245 1275 11260 1290
rect 11300 1285 12360 1300
rect 11300 1275 11315 1285
rect 11355 1275 11370 1285
rect 11410 1275 11425 1285
rect 11465 1275 11480 1285
rect 11520 1275 11535 1285
rect 11575 1275 11590 1285
rect 11630 1275 11645 1285
rect 11685 1275 11700 1285
rect 11740 1275 11755 1285
rect 11795 1275 11810 1285
rect 11850 1275 11865 1285
rect 11905 1275 11920 1285
rect 11960 1275 11975 1285
rect 12015 1275 12030 1285
rect 12070 1275 12085 1285
rect 12125 1275 12140 1285
rect 12180 1275 12195 1285
rect 12235 1275 12250 1285
rect 12290 1275 12305 1285
rect 12345 1275 12360 1285
rect 12400 1285 12470 1300
rect 12400 1275 12415 1285
rect 12455 1275 12470 1285
rect 12510 1275 12525 1315
rect 12565 1275 12580 1290
rect 2875 1190 3375 1205
rect 3415 1190 3915 1205
rect 4095 1190 4595 1205
rect 4635 1190 5135 1205
rect 3025 1120 3065 1130
rect 3025 1100 3035 1120
rect 3055 1100 3065 1120
rect 3025 1090 3065 1100
rect 3105 1120 3145 1130
rect 3105 1100 3115 1120
rect 3135 1100 3145 1120
rect 3105 1090 3145 1100
rect 3185 1120 3225 1130
rect 3185 1100 3195 1120
rect 3215 1100 3225 1120
rect 3185 1090 3225 1100
rect 3265 1120 3305 1130
rect 3265 1100 3275 1120
rect 3295 1100 3305 1120
rect 3265 1090 3305 1100
rect 3345 1120 3385 1130
rect 3345 1100 3355 1120
rect 3375 1100 3385 1120
rect 3345 1090 3385 1100
rect 3425 1120 3465 1130
rect 3425 1100 3435 1120
rect 3455 1100 3465 1120
rect 3425 1090 3465 1100
rect 3505 1120 3545 1130
rect 3505 1100 3515 1120
rect 3535 1100 3545 1120
rect 3505 1090 3545 1100
rect 3585 1120 3625 1130
rect 3585 1100 3595 1120
rect 3615 1100 3625 1120
rect 3585 1090 3625 1100
rect 3665 1120 3705 1130
rect 3665 1100 3675 1120
rect 3695 1100 3705 1120
rect 3665 1090 3705 1100
rect 3745 1120 3785 1130
rect 3745 1100 3755 1120
rect 3775 1100 3785 1120
rect 3745 1090 3785 1100
rect 3825 1120 3865 1130
rect 3825 1100 3835 1120
rect 3855 1100 3865 1120
rect 3825 1090 3865 1100
rect 3905 1120 3945 1130
rect 3905 1100 3915 1120
rect 3935 1100 3945 1120
rect 3905 1090 3945 1100
rect 4065 1120 4105 1130
rect 4065 1100 4075 1120
rect 4095 1100 4105 1120
rect 4065 1090 4105 1100
rect 4145 1120 4185 1130
rect 4145 1100 4155 1120
rect 4175 1100 4185 1120
rect 4145 1090 4185 1100
rect 4225 1120 4265 1130
rect 4225 1100 4235 1120
rect 4255 1100 4265 1120
rect 4225 1090 4265 1100
rect 4305 1120 4345 1130
rect 4305 1100 4315 1120
rect 4335 1100 4345 1120
rect 4305 1090 4345 1100
rect 4385 1120 4425 1130
rect 4385 1100 4395 1120
rect 4415 1100 4425 1120
rect 4385 1090 4425 1100
rect 4465 1120 4505 1130
rect 4465 1100 4475 1120
rect 4495 1100 4505 1120
rect 4465 1090 4505 1100
rect 4545 1120 4585 1130
rect 4545 1100 4555 1120
rect 4575 1100 4585 1120
rect 4545 1090 4585 1100
rect 4625 1120 4665 1130
rect 4625 1100 4635 1120
rect 4655 1100 4665 1120
rect 4625 1090 4665 1100
rect 4705 1120 4745 1130
rect 4705 1100 4715 1120
rect 4735 1100 4745 1120
rect 4705 1090 4745 1100
rect 4785 1120 4825 1130
rect 4785 1100 4795 1120
rect 4815 1100 4825 1120
rect 4785 1090 4825 1100
rect 4865 1120 4905 1130
rect 4865 1100 4875 1120
rect 4895 1100 4905 1120
rect 4865 1090 4905 1100
rect 4945 1120 4985 1130
rect 4945 1100 4955 1120
rect 4975 1100 4985 1120
rect 4945 1090 4985 1100
rect 2985 1075 3985 1090
rect 4025 1075 5025 1090
rect 11245 1010 11260 1025
rect 11300 1010 11315 1025
rect 11355 1010 11370 1025
rect 11410 1010 11425 1025
rect 11465 1010 11480 1025
rect 11520 1010 11535 1025
rect 11575 1010 11590 1025
rect 11630 1010 11645 1025
rect 11685 1010 11700 1025
rect 11740 1010 11755 1025
rect 11795 1010 11810 1025
rect 11850 1010 11865 1025
rect 11905 1010 11920 1025
rect 11960 1010 11975 1025
rect 12015 1010 12030 1025
rect 12070 1010 12085 1025
rect 12125 1010 12140 1025
rect 12180 1010 12195 1025
rect 12235 1010 12250 1025
rect 12290 1010 12305 1025
rect 12345 1010 12360 1025
rect 12400 1010 12415 1025
rect 12455 1010 12470 1025
rect 12510 1010 12525 1025
rect 12565 1010 12580 1025
rect 11165 1000 11260 1010
rect 11165 980 11175 1000
rect 11195 995 11260 1000
rect 12565 1000 12660 1010
rect 12565 995 12630 1000
rect 11195 980 11205 995
rect 2985 960 3985 975
rect 4025 960 5025 975
rect 11165 970 11205 980
rect 12620 980 12630 995
rect 12650 980 12660 1000
rect 12620 970 12660 980
rect 2995 925 3035 935
rect 2995 905 3005 925
rect 3025 905 3035 925
rect 4975 925 5015 935
rect 4975 905 4985 925
rect 5005 905 5015 925
rect 2995 890 3085 905
rect 3035 880 3085 890
rect 3125 890 4885 905
rect 3125 880 3175 890
rect 3215 880 3265 890
rect 3305 880 3355 890
rect 3395 880 3445 890
rect 3485 880 3535 890
rect 3575 880 3625 890
rect 3665 880 3715 890
rect 3755 880 3805 890
rect 3845 880 3895 890
rect 3935 880 3985 890
rect 4025 880 4075 890
rect 4115 880 4165 890
rect 4205 880 4255 890
rect 4295 880 4345 890
rect 4385 880 4435 890
rect 4475 880 4525 890
rect 4565 880 4615 890
rect 4655 880 4705 890
rect 4745 880 4795 890
rect 4835 880 4885 890
rect 4925 890 5015 905
rect 4925 880 4975 890
rect 3035 765 3085 780
rect 3125 755 3175 780
rect 3215 765 3265 780
rect 3305 765 3355 780
rect 3395 765 3445 780
rect 3485 765 3535 780
rect 3575 765 3625 780
rect 3665 765 3715 780
rect 3755 765 3805 780
rect 3845 765 3895 780
rect 3935 765 3985 780
rect 4025 765 4075 780
rect 4115 765 4165 780
rect 4205 765 4255 780
rect 4295 765 4345 780
rect 4385 765 4435 780
rect 4475 765 4525 780
rect 4565 765 4615 780
rect 4655 765 4705 780
rect 4745 765 4795 780
rect 4835 765 4885 780
rect 4925 765 4975 780
rect 3125 750 3140 755
rect 3130 735 3140 750
rect 3160 750 3175 755
rect 3160 735 3170 750
rect 3130 725 3170 735
<< polycont >>
rect 3145 2955 3165 2975
rect 4845 2955 4865 2975
rect 3005 2785 3025 2805
rect 4985 2785 5005 2805
rect 3185 2725 3205 2745
rect 4805 2725 4825 2745
rect 3365 2350 3385 2370
rect 3895 2355 3915 2375
rect 2630 1855 2650 1875
rect 2775 1855 2795 1875
rect 2845 1855 2865 1875
rect 2935 1855 2955 1875
rect 3175 1855 3195 1875
rect 3295 1855 3315 1875
rect 3535 1855 3555 1875
rect 3655 1855 3675 1875
rect 3865 1855 3885 1875
rect 3995 1850 4015 1870
rect 4125 1855 4145 1875
rect 4335 1855 4355 1875
rect 4455 1855 4475 1875
rect 4695 1855 4715 1875
rect 4815 1855 4835 1875
rect 5055 1855 5075 1875
rect 5145 1855 5165 1875
rect 5215 1855 5235 1875
rect 3235 1735 3255 1755
rect 4755 1735 4775 1755
rect 11243 1740 11260 1760
rect 11463 1740 11480 1760
rect 11610 1740 11627 1760
rect 11876 1740 11893 1760
rect 12283 1740 12300 1760
rect 12503 1740 12520 1760
rect 12650 1740 12667 1760
rect 3175 1570 3195 1590
rect 4815 1570 4835 1590
rect 11000 1520 11020 1540
rect 11112 1520 11129 1540
rect 11315 1520 11335 1540
rect 11535 1520 11555 1540
rect 11740 1520 11760 1540
rect 11928 1520 11945 1540
rect 12040 1520 12060 1540
rect 12152 1520 12169 1540
rect 12355 1520 12375 1540
rect 12575 1520 12595 1540
rect 12780 1520 12800 1540
rect 2935 1475 2955 1495
rect 3055 1475 3075 1495
rect 3175 1475 3195 1495
rect 3295 1475 3315 1495
rect 3535 1475 3555 1495
rect 3655 1475 3675 1495
rect 3775 1475 3795 1495
rect 4215 1475 4235 1495
rect 4335 1475 4355 1495
rect 4455 1475 4475 1495
rect 4695 1475 4715 1495
rect 4815 1475 4835 1495
rect 4935 1475 4955 1495
rect 5055 1475 5075 1495
rect 11820 1300 11840 1320
rect 3035 1100 3055 1120
rect 3115 1100 3135 1120
rect 3195 1100 3215 1120
rect 3275 1100 3295 1120
rect 3355 1100 3375 1120
rect 3435 1100 3455 1120
rect 3515 1100 3535 1120
rect 3595 1100 3615 1120
rect 3675 1100 3695 1120
rect 3755 1100 3775 1120
rect 3835 1100 3855 1120
rect 3915 1100 3935 1120
rect 4075 1100 4095 1120
rect 4155 1100 4175 1120
rect 4235 1100 4255 1120
rect 4315 1100 4335 1120
rect 4395 1100 4415 1120
rect 4475 1100 4495 1120
rect 4555 1100 4575 1120
rect 4635 1100 4655 1120
rect 4715 1100 4735 1120
rect 4795 1100 4815 1120
rect 4875 1100 4895 1120
rect 4955 1100 4975 1120
rect 11175 980 11195 1000
rect 12630 980 12650 1000
rect 3005 905 3025 925
rect 4985 905 5005 925
rect 3140 735 3160 755
<< xpolycontact >>
rect 91 3170 311 3205
rect 925 3170 1145 3205
rect 1306 3165 1526 3200
rect 2110 3165 2330 3200
rect 91 3110 311 3145
rect 925 3110 1145 3145
rect 1306 3105 1526 3140
rect 2110 3105 2330 3140
rect 91 3030 311 3065
rect 895 3030 1115 3065
rect 1306 3045 1526 3080
rect 2110 3045 2330 3080
rect 91 2970 311 3005
rect 895 2970 1115 3005
rect 1306 2985 1526 3020
rect 2110 2985 2330 3020
rect 1306 2925 1526 2960
rect 2110 2925 2330 2960
rect 1306 2865 1526 2900
rect 2110 2865 2330 2900
rect 96 2820 315 2855
rect 504 2820 724 2855
rect 1306 2805 1526 2840
rect 1740 2805 1960 2840
rect 96 2760 315 2795
rect 504 2760 724 2795
<< ppolyres >>
rect 315 2820 504 2855
rect 315 2760 504 2795
<< xpolyres >>
rect 311 3170 925 3205
rect 1526 3165 2110 3200
rect 311 3110 925 3145
rect 1526 3105 2110 3140
rect 311 3030 895 3065
rect 1526 3045 2110 3080
rect 311 2970 895 3005
rect 1526 2985 2110 3020
rect 1526 2925 2110 2960
rect 1526 2865 2110 2900
rect 1526 2805 1740 2840
<< locali >>
rect 1266 3495 1296 3525
rect 4445 3465 4475 3495
rect -10 3415 20 3445
rect 945 3415 975 3445
rect 1645 3415 1675 3445
rect 2475 3420 2505 3450
rect 5145 3415 5175 3445
rect -55 3360 -25 3390
rect 2695 3360 2725 3390
rect 1210 3310 1240 3340
rect 3140 3310 3170 3340
rect 3395 3305 3425 3335
rect 5365 3305 5395 3335
rect 1165 3255 1195 3285
rect 4890 3255 4920 3285
rect 5415 3255 5445 3285
rect 2740 3210 2770 3240
rect 46 3200 91 3205
rect 46 3175 56 3200
rect 81 3175 91 3200
rect 46 3170 91 3175
rect 1110 3145 1145 3170
rect 1261 3195 1306 3200
rect 1261 3170 1271 3195
rect 1296 3170 1306 3195
rect 1261 3165 1306 3170
rect 2330 3165 2370 3200
rect 46 3140 91 3145
rect 46 3115 56 3140
rect 81 3115 91 3140
rect 46 3110 91 3115
rect 1261 3135 1306 3140
rect 1261 3110 1271 3135
rect 1296 3110 1306 3135
rect 1261 3105 1306 3110
rect 1165 3070 1195 3100
rect 2295 3080 2330 3105
rect 46 3060 91 3065
rect 46 3035 56 3060
rect 81 3035 91 3060
rect 46 3030 91 3035
rect 1080 3005 1115 3030
rect 46 3000 91 3005
rect 46 2975 56 3000
rect 81 2975 91 3000
rect 46 2970 91 2975
rect 1266 3045 1306 3080
rect 910 2910 1120 2915
rect 910 2880 920 2910
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1120 2910
rect 910 2875 1120 2880
rect 1266 2900 1286 3045
rect 2350 3020 2370 3165
rect 2625 3155 2655 3185
rect 4445 3155 4475 3185
rect 3140 3110 3170 3140
rect 4840 3110 4870 3140
rect 5320 3110 5350 3140
rect 3990 3050 4020 3080
rect 2330 2985 2370 3020
rect 3450 3005 3480 3035
rect 3810 3005 3840 3035
rect 4350 3005 4380 3035
rect 4710 3005 4740 3035
rect 1306 2960 1341 2985
rect 2330 2955 2375 2960
rect 2330 2930 2340 2955
rect 2365 2930 2375 2955
rect 2330 2925 2375 2930
rect 2430 2925 2460 2955
rect 2520 2945 2560 2985
rect 3080 2975 3120 2985
rect 3080 2955 3090 2975
rect 3110 2955 3120 2975
rect 3080 2945 3120 2955
rect 3140 2975 3175 2985
rect 3140 2955 3145 2975
rect 3165 2955 3175 2975
rect 3140 2945 3175 2955
rect 3265 2975 3305 2985
rect 3265 2955 3275 2975
rect 3295 2955 3305 2975
rect 3265 2945 3305 2955
rect 3445 2975 3485 2985
rect 3445 2955 3455 2975
rect 3475 2955 3485 2975
rect 3445 2945 3485 2955
rect 3625 2975 3665 2985
rect 3625 2955 3635 2975
rect 3655 2955 3665 2975
rect 3625 2945 3665 2955
rect 3805 2975 3845 2985
rect 3805 2955 3815 2975
rect 3835 2955 3845 2975
rect 3805 2945 3845 2955
rect 3985 2975 4025 2985
rect 3985 2955 3995 2975
rect 4015 2955 4025 2975
rect 3985 2945 4025 2955
rect 4165 2975 4205 2985
rect 4165 2955 4175 2975
rect 4195 2955 4205 2975
rect 4165 2945 4205 2955
rect 4345 2975 4385 2985
rect 4345 2955 4355 2975
rect 4375 2955 4385 2975
rect 4345 2945 4385 2955
rect 4525 2975 4565 2985
rect 4525 2955 4535 2975
rect 4555 2955 4565 2975
rect 4525 2945 4565 2955
rect 4705 2975 4745 2985
rect 4705 2955 4715 2975
rect 4735 2955 4745 2975
rect 4705 2945 4745 2955
rect 4835 2975 4870 2985
rect 4835 2955 4845 2975
rect 4865 2955 4870 2975
rect 4835 2945 4870 2955
rect 4890 2975 4925 2985
rect 4890 2955 4895 2975
rect 4915 2955 4925 2975
rect 4890 2945 4925 2955
rect 3095 2925 3115 2945
rect 3275 2925 3295 2945
rect 3455 2925 3475 2945
rect 3635 2925 3655 2945
rect 3815 2925 3835 2945
rect 3995 2925 4015 2945
rect 4175 2925 4195 2945
rect 4355 2925 4375 2945
rect 4535 2925 4555 2945
rect 4715 2925 4735 2945
rect 4895 2925 4915 2945
rect 2960 2915 3030 2925
rect 1266 2865 1306 2900
rect 2330 2895 2375 2905
rect 2330 2870 2340 2895
rect 2365 2870 2375 2895
rect 2330 2860 2375 2870
rect 2960 2895 2965 2915
rect 2985 2895 3005 2915
rect 3025 2895 3030 2915
rect 2960 2865 3030 2895
rect -55 2825 -25 2855
rect 51 2850 96 2855
rect 51 2825 61 2850
rect 86 2825 96 2850
rect 51 2820 96 2825
rect 724 2850 769 2855
rect 724 2825 734 2850
rect 759 2825 769 2850
rect 724 2820 769 2825
rect 1210 2820 1240 2850
rect 2960 2845 2965 2865
rect 2985 2845 3005 2865
rect 3025 2845 3030 2865
rect 1261 2835 1306 2840
rect 1261 2810 1271 2835
rect 1296 2810 1306 2835
rect 1261 2805 1306 2810
rect 1960 2835 2005 2840
rect 1960 2810 1970 2835
rect 1995 2810 2005 2835
rect 1960 2805 2005 2810
rect 2330 2800 2370 2840
rect 2960 2835 3030 2845
rect 3090 2915 3120 2925
rect 3090 2895 3095 2915
rect 3115 2895 3120 2915
rect 3090 2865 3120 2895
rect 3090 2845 3095 2865
rect 3115 2845 3120 2865
rect 3090 2835 3120 2845
rect 3180 2915 3210 2925
rect 3180 2895 3185 2915
rect 3205 2895 3210 2915
rect 3180 2865 3210 2895
rect 3180 2845 3185 2865
rect 3205 2845 3210 2865
rect 3180 2835 3210 2845
rect 3270 2915 3300 2925
rect 3270 2895 3275 2915
rect 3295 2895 3300 2915
rect 3270 2865 3300 2895
rect 3270 2845 3275 2865
rect 3295 2845 3300 2865
rect 3270 2835 3300 2845
rect 3360 2915 3390 2925
rect 3360 2895 3365 2915
rect 3385 2895 3390 2915
rect 3360 2865 3390 2895
rect 3360 2845 3365 2865
rect 3385 2845 3390 2865
rect 3360 2835 3390 2845
rect 3450 2915 3480 2925
rect 3450 2895 3455 2915
rect 3475 2895 3480 2915
rect 3450 2865 3480 2895
rect 3450 2845 3455 2865
rect 3475 2845 3480 2865
rect 3450 2835 3480 2845
rect 3540 2915 3570 2925
rect 3540 2895 3545 2915
rect 3565 2895 3570 2915
rect 3540 2865 3570 2895
rect 3540 2845 3545 2865
rect 3565 2845 3570 2865
rect 3540 2835 3570 2845
rect 3630 2915 3660 2925
rect 3630 2895 3635 2915
rect 3655 2895 3660 2915
rect 3630 2865 3660 2895
rect 3630 2845 3635 2865
rect 3655 2845 3660 2865
rect 3630 2835 3660 2845
rect 3720 2915 3750 2925
rect 3720 2895 3725 2915
rect 3745 2895 3750 2915
rect 3720 2865 3750 2895
rect 3720 2845 3725 2865
rect 3745 2845 3750 2865
rect 3720 2835 3750 2845
rect 3810 2915 3840 2925
rect 3810 2895 3815 2915
rect 3835 2895 3840 2915
rect 3810 2865 3840 2895
rect 3810 2845 3815 2865
rect 3835 2845 3840 2865
rect 3810 2835 3840 2845
rect 3900 2915 3930 2925
rect 3900 2895 3905 2915
rect 3925 2895 3930 2915
rect 3900 2865 3930 2895
rect 3900 2845 3905 2865
rect 3925 2845 3930 2865
rect 3900 2835 3930 2845
rect 3990 2915 4020 2925
rect 3990 2895 3995 2915
rect 4015 2895 4020 2915
rect 3990 2865 4020 2895
rect 3990 2845 3995 2865
rect 4015 2845 4020 2865
rect 3990 2835 4020 2845
rect 4080 2915 4110 2925
rect 4080 2895 4085 2915
rect 4105 2895 4110 2915
rect 4080 2865 4110 2895
rect 4080 2845 4085 2865
rect 4105 2845 4110 2865
rect 4080 2835 4110 2845
rect 4170 2915 4200 2925
rect 4170 2895 4175 2915
rect 4195 2895 4200 2915
rect 4170 2865 4200 2895
rect 4170 2845 4175 2865
rect 4195 2845 4200 2865
rect 4170 2835 4200 2845
rect 4260 2915 4290 2925
rect 4260 2895 4265 2915
rect 4285 2895 4290 2915
rect 4260 2865 4290 2895
rect 4260 2845 4265 2865
rect 4285 2845 4290 2865
rect 4260 2835 4290 2845
rect 4350 2915 4380 2925
rect 4350 2895 4355 2915
rect 4375 2895 4380 2915
rect 4350 2865 4380 2895
rect 4350 2845 4355 2865
rect 4375 2845 4380 2865
rect 4350 2835 4380 2845
rect 4440 2915 4470 2925
rect 4440 2895 4445 2915
rect 4465 2895 4470 2915
rect 4440 2865 4470 2895
rect 4440 2845 4445 2865
rect 4465 2845 4470 2865
rect 4440 2835 4470 2845
rect 4530 2915 4560 2925
rect 4530 2895 4535 2915
rect 4555 2895 4560 2915
rect 4530 2865 4560 2895
rect 4530 2845 4535 2865
rect 4555 2845 4560 2865
rect 4530 2835 4560 2845
rect 4620 2915 4650 2925
rect 4620 2895 4625 2915
rect 4645 2895 4650 2915
rect 4620 2865 4650 2895
rect 4620 2845 4625 2865
rect 4645 2845 4650 2865
rect 4620 2835 4650 2845
rect 4710 2915 4740 2925
rect 4710 2895 4715 2915
rect 4735 2895 4740 2915
rect 4710 2865 4740 2895
rect 4710 2845 4715 2865
rect 4735 2845 4740 2865
rect 4710 2835 4740 2845
rect 4800 2915 4830 2925
rect 4800 2895 4805 2915
rect 4825 2895 4830 2915
rect 4800 2865 4830 2895
rect 4800 2845 4805 2865
rect 4825 2845 4830 2865
rect 4800 2835 4830 2845
rect 4890 2915 4920 2925
rect 4890 2895 4895 2915
rect 4915 2895 4920 2915
rect 4890 2865 4920 2895
rect 4890 2845 4895 2865
rect 4915 2845 4920 2865
rect 4890 2835 4920 2845
rect 4980 2915 5050 2925
rect 4980 2895 4985 2915
rect 5005 2895 5025 2915
rect 5045 2895 5050 2915
rect 4980 2865 5050 2895
rect 4980 2845 4985 2865
rect 5005 2845 5025 2865
rect 5045 2845 5050 2865
rect 4980 2835 5050 2845
rect 3005 2815 3025 2835
rect 3185 2815 3205 2835
rect 3365 2815 3385 2835
rect 3545 2815 3565 2835
rect 3725 2815 3745 2835
rect 3905 2815 3925 2835
rect 4085 2815 4105 2835
rect 4265 2815 4285 2835
rect 4445 2815 4465 2835
rect 4625 2815 4645 2835
rect 4805 2815 4825 2835
rect 4985 2815 5005 2835
rect 2995 2805 3035 2815
rect -10 2765 20 2795
rect 51 2790 96 2795
rect 51 2765 61 2790
rect 86 2765 96 2790
rect 51 2760 96 2765
rect 724 2790 769 2795
rect 724 2765 734 2790
rect 759 2765 769 2790
rect 724 2760 769 2765
rect 2620 2755 2660 2795
rect 2995 2785 3005 2805
rect 3025 2785 3035 2805
rect 2995 2775 3035 2785
rect 3175 2805 3215 2815
rect 3175 2785 3185 2805
rect 3205 2785 3215 2805
rect 3175 2775 3215 2785
rect 3355 2805 3395 2815
rect 3355 2785 3365 2805
rect 3385 2785 3395 2805
rect 3355 2775 3395 2785
rect 3535 2805 3575 2815
rect 3535 2785 3545 2805
rect 3565 2785 3575 2805
rect 3535 2775 3575 2785
rect 3715 2805 3755 2815
rect 3715 2785 3725 2805
rect 3745 2785 3755 2805
rect 3715 2775 3755 2785
rect 3895 2805 3935 2815
rect 3895 2785 3905 2805
rect 3925 2785 3935 2805
rect 3895 2775 3935 2785
rect 4075 2805 4115 2815
rect 4075 2785 4085 2805
rect 4105 2785 4115 2805
rect 4075 2775 4115 2785
rect 4255 2805 4295 2815
rect 4255 2785 4265 2805
rect 4285 2785 4295 2805
rect 4255 2775 4295 2785
rect 4435 2805 4475 2815
rect 4435 2785 4445 2805
rect 4465 2785 4475 2805
rect 4435 2775 4475 2785
rect 4615 2805 4655 2815
rect 4615 2785 4625 2805
rect 4645 2785 4655 2805
rect 4615 2775 4655 2785
rect 4795 2805 4835 2815
rect 4795 2785 4805 2805
rect 4825 2785 4835 2805
rect 4795 2775 4835 2785
rect 4975 2805 5015 2815
rect 4975 2785 4985 2805
rect 5005 2785 5015 2805
rect 4975 2775 5015 2785
rect 1266 2715 1296 2745
rect 2150 2710 2190 2750
rect 3175 2745 3215 2755
rect 3175 2725 3185 2745
rect 3205 2725 3215 2745
rect 3175 2715 3215 2725
rect 3355 2745 3395 2755
rect 3355 2725 3365 2745
rect 3385 2725 3395 2745
rect 3355 2715 3395 2725
rect 3535 2745 3575 2755
rect 3535 2725 3545 2745
rect 3565 2725 3575 2745
rect 3535 2715 3575 2725
rect 3715 2745 3755 2755
rect 3715 2725 3725 2745
rect 3745 2725 3755 2745
rect 3715 2715 3755 2725
rect 3895 2745 3935 2755
rect 3895 2725 3905 2745
rect 3925 2725 3935 2745
rect 3895 2715 3935 2725
rect 4075 2745 4115 2755
rect 4075 2725 4085 2745
rect 4105 2725 4115 2745
rect 4075 2715 4115 2725
rect 4255 2745 4295 2755
rect 4255 2725 4265 2745
rect 4285 2725 4295 2745
rect 4255 2715 4295 2725
rect 4435 2745 4475 2755
rect 4435 2725 4445 2745
rect 4465 2725 4475 2745
rect 4435 2715 4475 2725
rect 4615 2745 4655 2755
rect 4615 2725 4625 2745
rect 4645 2725 4655 2745
rect 4615 2715 4655 2725
rect 4795 2745 4835 2755
rect 4795 2725 4805 2745
rect 4825 2725 4835 2745
rect 4795 2715 4835 2725
rect 650 2055 775 2700
rect 1330 2055 1455 2700
rect 2010 2055 2135 2700
rect 3185 2695 3205 2715
rect 3365 2695 3385 2715
rect 3545 2695 3565 2715
rect 3725 2695 3745 2715
rect 3905 2695 3925 2715
rect 4085 2695 4105 2715
rect 4265 2695 4285 2715
rect 4445 2695 4465 2715
rect 4625 2695 4645 2715
rect 4805 2695 4825 2715
rect 3140 2685 3210 2695
rect 3140 2665 3145 2685
rect 3165 2665 3185 2685
rect 3205 2665 3210 2685
rect 3140 2635 3210 2665
rect 3140 2615 3145 2635
rect 3165 2615 3185 2635
rect 3205 2615 3210 2635
rect 3140 2585 3210 2615
rect 3140 2565 3145 2585
rect 3165 2565 3185 2585
rect 3205 2565 3210 2585
rect 3140 2535 3210 2565
rect 3140 2515 3145 2535
rect 3165 2515 3185 2535
rect 3205 2515 3210 2535
rect 3140 2485 3210 2515
rect 3140 2465 3145 2485
rect 3165 2465 3185 2485
rect 3205 2465 3210 2485
rect 3140 2435 3210 2465
rect 3140 2415 3145 2435
rect 3165 2415 3185 2435
rect 3205 2415 3210 2435
rect 3140 2405 3210 2415
rect 3270 2685 3300 2695
rect 3270 2665 3275 2685
rect 3295 2665 3300 2685
rect 3270 2635 3300 2665
rect 3270 2615 3275 2635
rect 3295 2615 3300 2635
rect 3270 2585 3300 2615
rect 3270 2565 3275 2585
rect 3295 2565 3300 2585
rect 3270 2535 3300 2565
rect 3270 2515 3275 2535
rect 3295 2515 3300 2535
rect 3270 2485 3300 2515
rect 3270 2465 3275 2485
rect 3295 2465 3300 2485
rect 3270 2435 3300 2465
rect 3270 2415 3275 2435
rect 3295 2415 3300 2435
rect 3270 2405 3300 2415
rect 3360 2685 3390 2695
rect 3360 2665 3365 2685
rect 3385 2665 3390 2685
rect 3360 2635 3390 2665
rect 3360 2615 3365 2635
rect 3385 2615 3390 2635
rect 3360 2585 3390 2615
rect 3360 2565 3365 2585
rect 3385 2565 3390 2585
rect 3360 2535 3390 2565
rect 3360 2515 3365 2535
rect 3385 2515 3390 2535
rect 3360 2485 3390 2515
rect 3360 2465 3365 2485
rect 3385 2465 3390 2485
rect 3360 2435 3390 2465
rect 3360 2415 3365 2435
rect 3385 2415 3390 2435
rect 3360 2405 3390 2415
rect 3450 2685 3480 2695
rect 3450 2665 3455 2685
rect 3475 2665 3480 2685
rect 3450 2635 3480 2665
rect 3450 2615 3455 2635
rect 3475 2615 3480 2635
rect 3450 2585 3480 2615
rect 3450 2565 3455 2585
rect 3475 2565 3480 2585
rect 3450 2535 3480 2565
rect 3450 2515 3455 2535
rect 3475 2515 3480 2535
rect 3450 2485 3480 2515
rect 3450 2465 3455 2485
rect 3475 2465 3480 2485
rect 3450 2435 3480 2465
rect 3450 2415 3455 2435
rect 3475 2415 3480 2435
rect 3450 2405 3480 2415
rect 3540 2685 3570 2695
rect 3540 2665 3545 2685
rect 3565 2665 3570 2685
rect 3540 2635 3570 2665
rect 3540 2615 3545 2635
rect 3565 2615 3570 2635
rect 3540 2585 3570 2615
rect 3540 2565 3545 2585
rect 3565 2565 3570 2585
rect 3540 2535 3570 2565
rect 3540 2515 3545 2535
rect 3565 2515 3570 2535
rect 3540 2485 3570 2515
rect 3540 2465 3545 2485
rect 3565 2465 3570 2485
rect 3540 2435 3570 2465
rect 3540 2415 3545 2435
rect 3565 2415 3570 2435
rect 3540 2405 3570 2415
rect 3630 2685 3660 2695
rect 3630 2665 3635 2685
rect 3655 2665 3660 2685
rect 3630 2635 3660 2665
rect 3630 2615 3635 2635
rect 3655 2615 3660 2635
rect 3630 2585 3660 2615
rect 3630 2565 3635 2585
rect 3655 2565 3660 2585
rect 3630 2535 3660 2565
rect 3630 2515 3635 2535
rect 3655 2515 3660 2535
rect 3630 2485 3660 2515
rect 3630 2465 3635 2485
rect 3655 2465 3660 2485
rect 3630 2435 3660 2465
rect 3630 2415 3635 2435
rect 3655 2415 3660 2435
rect 3630 2405 3660 2415
rect 3720 2685 3750 2695
rect 3720 2665 3725 2685
rect 3745 2665 3750 2685
rect 3720 2635 3750 2665
rect 3720 2615 3725 2635
rect 3745 2615 3750 2635
rect 3720 2585 3750 2615
rect 3720 2565 3725 2585
rect 3745 2565 3750 2585
rect 3720 2535 3750 2565
rect 3720 2515 3725 2535
rect 3745 2515 3750 2535
rect 3720 2485 3750 2515
rect 3720 2465 3725 2485
rect 3745 2465 3750 2485
rect 3720 2435 3750 2465
rect 3720 2415 3725 2435
rect 3745 2415 3750 2435
rect 3720 2405 3750 2415
rect 3810 2685 3840 2695
rect 3810 2665 3815 2685
rect 3835 2665 3840 2685
rect 3810 2635 3840 2665
rect 3810 2615 3815 2635
rect 3835 2615 3840 2635
rect 3810 2585 3840 2615
rect 3810 2565 3815 2585
rect 3835 2565 3840 2585
rect 3810 2535 3840 2565
rect 3810 2515 3815 2535
rect 3835 2515 3840 2535
rect 3810 2485 3840 2515
rect 3810 2465 3815 2485
rect 3835 2465 3840 2485
rect 3810 2435 3840 2465
rect 3810 2415 3815 2435
rect 3835 2415 3840 2435
rect 3810 2405 3840 2415
rect 3900 2685 3930 2695
rect 3900 2665 3905 2685
rect 3925 2665 3930 2685
rect 3900 2635 3930 2665
rect 3900 2615 3905 2635
rect 3925 2615 3930 2635
rect 3900 2585 3930 2615
rect 3900 2565 3905 2585
rect 3925 2565 3930 2585
rect 3900 2535 3930 2565
rect 3900 2515 3905 2535
rect 3925 2515 3930 2535
rect 3900 2485 3930 2515
rect 3900 2465 3905 2485
rect 3925 2465 3930 2485
rect 3900 2435 3930 2465
rect 3900 2415 3905 2435
rect 3925 2415 3930 2435
rect 3900 2405 3930 2415
rect 3990 2685 4020 2695
rect 3990 2665 3995 2685
rect 4015 2665 4020 2685
rect 3990 2635 4020 2665
rect 3990 2615 3995 2635
rect 4015 2615 4020 2635
rect 3990 2585 4020 2615
rect 3990 2565 3995 2585
rect 4015 2565 4020 2585
rect 3990 2535 4020 2565
rect 3990 2515 3995 2535
rect 4015 2515 4020 2535
rect 3990 2485 4020 2515
rect 3990 2465 3995 2485
rect 4015 2465 4020 2485
rect 3990 2435 4020 2465
rect 3990 2415 3995 2435
rect 4015 2415 4020 2435
rect 3990 2405 4020 2415
rect 4080 2685 4110 2695
rect 4080 2665 4085 2685
rect 4105 2665 4110 2685
rect 4080 2635 4110 2665
rect 4080 2615 4085 2635
rect 4105 2615 4110 2635
rect 4080 2585 4110 2615
rect 4080 2565 4085 2585
rect 4105 2565 4110 2585
rect 4080 2535 4110 2565
rect 4080 2515 4085 2535
rect 4105 2515 4110 2535
rect 4080 2485 4110 2515
rect 4080 2465 4085 2485
rect 4105 2465 4110 2485
rect 4080 2435 4110 2465
rect 4080 2415 4085 2435
rect 4105 2415 4110 2435
rect 4080 2405 4110 2415
rect 4170 2685 4200 2695
rect 4170 2665 4175 2685
rect 4195 2665 4200 2685
rect 4170 2635 4200 2665
rect 4170 2615 4175 2635
rect 4195 2615 4200 2635
rect 4170 2585 4200 2615
rect 4170 2565 4175 2585
rect 4195 2565 4200 2585
rect 4170 2535 4200 2565
rect 4170 2515 4175 2535
rect 4195 2515 4200 2535
rect 4170 2485 4200 2515
rect 4170 2465 4175 2485
rect 4195 2465 4200 2485
rect 4170 2435 4200 2465
rect 4170 2415 4175 2435
rect 4195 2415 4200 2435
rect 4170 2405 4200 2415
rect 4260 2685 4290 2695
rect 4260 2665 4265 2685
rect 4285 2665 4290 2685
rect 4260 2635 4290 2665
rect 4260 2615 4265 2635
rect 4285 2615 4290 2635
rect 4260 2585 4290 2615
rect 4260 2565 4265 2585
rect 4285 2565 4290 2585
rect 4260 2535 4290 2565
rect 4260 2515 4265 2535
rect 4285 2515 4290 2535
rect 4260 2485 4290 2515
rect 4260 2465 4265 2485
rect 4285 2465 4290 2485
rect 4260 2435 4290 2465
rect 4260 2415 4265 2435
rect 4285 2415 4290 2435
rect 4260 2405 4290 2415
rect 4350 2685 4380 2695
rect 4350 2665 4355 2685
rect 4375 2665 4380 2685
rect 4350 2635 4380 2665
rect 4350 2615 4355 2635
rect 4375 2615 4380 2635
rect 4350 2585 4380 2615
rect 4350 2565 4355 2585
rect 4375 2565 4380 2585
rect 4350 2535 4380 2565
rect 4350 2515 4355 2535
rect 4375 2515 4380 2535
rect 4350 2485 4380 2515
rect 4350 2465 4355 2485
rect 4375 2465 4380 2485
rect 4350 2435 4380 2465
rect 4350 2415 4355 2435
rect 4375 2415 4380 2435
rect 4350 2405 4380 2415
rect 4440 2685 4470 2695
rect 4440 2665 4445 2685
rect 4465 2665 4470 2685
rect 4440 2635 4470 2665
rect 4440 2615 4445 2635
rect 4465 2615 4470 2635
rect 4440 2585 4470 2615
rect 4440 2565 4445 2585
rect 4465 2565 4470 2585
rect 4440 2535 4470 2565
rect 4440 2515 4445 2535
rect 4465 2515 4470 2535
rect 4440 2485 4470 2515
rect 4440 2465 4445 2485
rect 4465 2465 4470 2485
rect 4440 2435 4470 2465
rect 4440 2415 4445 2435
rect 4465 2415 4470 2435
rect 4440 2405 4470 2415
rect 4530 2685 4560 2695
rect 4530 2665 4535 2685
rect 4555 2665 4560 2685
rect 4530 2635 4560 2665
rect 4530 2615 4535 2635
rect 4555 2615 4560 2635
rect 4530 2585 4560 2615
rect 4530 2565 4535 2585
rect 4555 2565 4560 2585
rect 4530 2535 4560 2565
rect 4530 2515 4535 2535
rect 4555 2515 4560 2535
rect 4530 2485 4560 2515
rect 4530 2465 4535 2485
rect 4555 2465 4560 2485
rect 4530 2435 4560 2465
rect 4530 2415 4535 2435
rect 4555 2415 4560 2435
rect 4530 2405 4560 2415
rect 4620 2685 4650 2695
rect 4620 2665 4625 2685
rect 4645 2665 4650 2685
rect 4620 2635 4650 2665
rect 4620 2615 4625 2635
rect 4645 2615 4650 2635
rect 4620 2585 4650 2615
rect 4620 2565 4625 2585
rect 4645 2565 4650 2585
rect 4620 2535 4650 2565
rect 4620 2515 4625 2535
rect 4645 2515 4650 2535
rect 4620 2485 4650 2515
rect 4620 2465 4625 2485
rect 4645 2465 4650 2485
rect 4620 2435 4650 2465
rect 4620 2415 4625 2435
rect 4645 2415 4650 2435
rect 4620 2405 4650 2415
rect 4710 2685 4740 2695
rect 4710 2665 4715 2685
rect 4735 2665 4740 2685
rect 4710 2635 4740 2665
rect 4710 2615 4715 2635
rect 4735 2615 4740 2635
rect 4710 2585 4740 2615
rect 4710 2565 4715 2585
rect 4735 2565 4740 2585
rect 4710 2535 4740 2565
rect 4710 2515 4715 2535
rect 4735 2515 4740 2535
rect 4710 2485 4740 2515
rect 4710 2465 4715 2485
rect 4735 2465 4740 2485
rect 4710 2435 4740 2465
rect 4710 2415 4715 2435
rect 4735 2415 4740 2435
rect 4710 2405 4740 2415
rect 4800 2685 4870 2695
rect 4800 2665 4805 2685
rect 4825 2665 4845 2685
rect 4865 2665 4870 2685
rect 4800 2635 4870 2665
rect 4800 2615 4805 2635
rect 4825 2615 4845 2635
rect 4865 2615 4870 2635
rect 4800 2585 4870 2615
rect 4800 2565 4805 2585
rect 4825 2565 4845 2585
rect 4865 2565 4870 2585
rect 4800 2535 4870 2565
rect 4800 2515 4805 2535
rect 4825 2515 4845 2535
rect 4865 2515 4870 2535
rect 4800 2485 4870 2515
rect 4800 2465 4805 2485
rect 4825 2465 4845 2485
rect 4865 2465 4870 2485
rect 4800 2435 4870 2465
rect 4800 2415 4805 2435
rect 4825 2415 4845 2435
rect 4865 2415 4870 2435
rect 4800 2405 4870 2415
rect 3275 2385 3295 2405
rect 3455 2385 3475 2405
rect 3265 2375 3305 2385
rect 3265 2355 3275 2375
rect 3295 2355 3305 2375
rect 3265 2345 3305 2355
rect 3355 2370 3395 2380
rect 3355 2350 3365 2370
rect 3385 2350 3395 2370
rect 2625 2315 2655 2345
rect 3355 2340 3395 2350
rect 3445 2375 3485 2385
rect 3445 2355 3455 2375
rect 3475 2355 3485 2375
rect 3445 2345 3485 2355
rect 3635 2340 3655 2405
rect 3815 2385 3835 2405
rect 3995 2385 4015 2405
rect 4175 2385 4195 2405
rect 3805 2375 3845 2385
rect 3805 2355 3815 2375
rect 3835 2355 3845 2375
rect 3805 2345 3845 2355
rect 3885 2375 3925 2385
rect 3885 2355 3895 2375
rect 3915 2355 3925 2375
rect 3885 2345 3925 2355
rect 3985 2375 4025 2385
rect 3985 2355 3995 2375
rect 4015 2355 4025 2375
rect 3985 2345 4025 2355
rect 4165 2375 4205 2385
rect 4165 2355 4175 2375
rect 4195 2355 4205 2375
rect 4165 2345 4205 2355
rect 4355 2340 4375 2405
rect 4535 2385 4555 2405
rect 4715 2385 4735 2405
rect 4525 2375 4565 2385
rect 4525 2355 4535 2375
rect 4555 2355 4565 2375
rect 4525 2345 4565 2355
rect 4705 2375 4745 2385
rect 4705 2355 4715 2375
rect 4735 2355 4745 2375
rect 4705 2345 4745 2355
rect 3625 2330 3665 2340
rect 3625 2310 3635 2330
rect 3655 2310 3665 2330
rect 3625 2300 3665 2310
rect 4345 2330 4385 2340
rect 4345 2310 4355 2330
rect 4375 2310 4385 2330
rect 4345 2300 4385 2310
rect 2740 2260 2770 2290
rect 3445 2285 3485 2295
rect 3445 2265 3455 2285
rect 3475 2265 3485 2285
rect 3445 2255 3485 2265
rect 4525 2285 4565 2295
rect 4525 2265 4535 2285
rect 4555 2265 4565 2285
rect 4525 2255 4565 2265
rect 5275 2260 5305 2290
rect 2430 2215 2460 2245
rect 3810 2215 3840 2245
rect 2335 2170 2365 2200
rect 2385 2120 2415 2150
rect 3630 2120 3660 2150
rect 4090 2115 4120 2145
rect 5320 2115 5350 2145
rect 2745 2090 2785 2100
rect 2745 2070 2755 2090
rect 2775 2070 2785 2090
rect 2745 2060 2785 2070
rect 2865 2090 2905 2100
rect 2865 2070 2875 2090
rect 2895 2070 2905 2090
rect 2865 2060 2905 2070
rect 2985 2090 3025 2100
rect 2985 2070 2995 2090
rect 3015 2070 3025 2090
rect 2985 2060 3025 2070
rect 3105 2090 3145 2100
rect 3105 2070 3115 2090
rect 3135 2070 3145 2090
rect 3105 2060 3145 2070
rect 3225 2090 3265 2100
rect 3225 2070 3235 2090
rect 3255 2070 3265 2090
rect 3225 2060 3265 2070
rect 3345 2090 3385 2100
rect 3345 2070 3355 2090
rect 3375 2070 3385 2090
rect 3345 2060 3385 2070
rect 3465 2090 3505 2100
rect 3465 2070 3475 2090
rect 3495 2070 3505 2090
rect 3465 2060 3505 2070
rect 3585 2090 3625 2100
rect 3585 2070 3595 2090
rect 3615 2070 3625 2090
rect 3585 2060 3625 2070
rect 3705 2090 3745 2100
rect 3705 2070 3715 2090
rect 3735 2070 3745 2090
rect 3705 2060 3745 2070
rect 3825 2090 3865 2100
rect 3825 2070 3835 2090
rect 3855 2070 3865 2090
rect 3825 2060 3865 2070
rect 3985 2090 4025 2100
rect 3985 2070 3995 2090
rect 4015 2070 4025 2090
rect 3985 2060 4025 2070
rect 4145 2090 4185 2100
rect 4145 2070 4155 2090
rect 4175 2070 4185 2090
rect 4145 2060 4185 2070
rect 4265 2090 4305 2100
rect 4265 2070 4275 2090
rect 4295 2070 4305 2090
rect 4265 2060 4305 2070
rect 4385 2090 4425 2100
rect 4385 2070 4395 2090
rect 4415 2070 4425 2090
rect 4385 2060 4425 2070
rect 4505 2090 4545 2100
rect 4505 2070 4515 2090
rect 4535 2070 4545 2090
rect 4505 2060 4545 2070
rect 4625 2090 4665 2100
rect 4625 2070 4635 2090
rect 4655 2070 4665 2090
rect 4625 2060 4665 2070
rect 4745 2090 4785 2100
rect 4745 2070 4755 2090
rect 4775 2070 4785 2090
rect 4745 2060 4785 2070
rect 4865 2090 4905 2100
rect 4865 2070 4875 2090
rect 4895 2070 4905 2090
rect 4865 2060 4905 2070
rect 4985 2090 5025 2100
rect 4985 2070 4995 2090
rect 5015 2070 5025 2090
rect 4985 2060 5025 2070
rect 5105 2090 5145 2100
rect 5105 2070 5115 2090
rect 5135 2070 5145 2090
rect 5105 2060 5145 2070
rect 5225 2090 5265 2100
rect 5225 2070 5235 2090
rect 5255 2070 5265 2090
rect 5225 2060 5265 2070
rect 125 2015 2135 2055
rect 2620 2045 2660 2055
rect 2620 2025 2630 2045
rect 2650 2025 2660 2045
rect 2620 2015 2660 2025
rect -45 1715 130 1725
rect -45 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 130 1715
rect -45 1685 130 1695
rect 650 1375 775 2015
rect 1330 1375 1455 2015
rect 2010 1375 2135 2015
rect 2630 1995 2650 2015
rect 2755 1995 2775 2060
rect 2805 2045 2845 2055
rect 2805 2025 2815 2045
rect 2835 2025 2845 2045
rect 2805 2015 2845 2025
rect 2815 1995 2835 2015
rect 2875 1995 2895 2060
rect 2995 1995 3015 2060
rect 3115 1995 3135 2060
rect 3165 2045 3205 2055
rect 3165 2025 3175 2045
rect 3195 2025 3205 2045
rect 3165 2015 3205 2025
rect 3175 1995 3195 2015
rect 3235 1995 3255 2060
rect 3355 1995 3375 2060
rect 3475 1995 3495 2060
rect 3525 2045 3565 2055
rect 3525 2025 3535 2045
rect 3555 2025 3565 2045
rect 3525 2015 3565 2025
rect 3535 1995 3555 2015
rect 3595 1995 3615 2060
rect 3715 1995 3735 2060
rect 3835 1995 3855 2060
rect 3885 2045 3925 2055
rect 3885 2025 3895 2045
rect 3915 2025 3925 2045
rect 3885 2015 3925 2025
rect 3895 1995 3915 2015
rect 3995 1995 4015 2060
rect 4085 2045 4125 2055
rect 4085 2025 4095 2045
rect 4115 2025 4125 2045
rect 4085 2015 4125 2025
rect 4095 1995 4115 2015
rect 4155 1995 4175 2060
rect 4275 1995 4295 2060
rect 4395 1995 4415 2060
rect 4445 2045 4485 2055
rect 4445 2025 4455 2045
rect 4475 2025 4485 2045
rect 4445 2015 4485 2025
rect 4455 1995 4475 2015
rect 4515 1995 4535 2060
rect 4635 1995 4655 2060
rect 4755 1995 4775 2060
rect 4805 2045 4845 2055
rect 4805 2025 4815 2045
rect 4835 2025 4845 2045
rect 4805 2015 4845 2025
rect 4815 1995 4835 2015
rect 4875 1995 4895 2060
rect 4995 1995 5015 2060
rect 5115 1995 5135 2060
rect 5165 2045 5205 2055
rect 5165 2025 5175 2045
rect 5195 2025 5205 2045
rect 5165 2015 5205 2025
rect 5175 1995 5195 2015
rect 5235 1995 5255 2060
rect 2570 1985 2600 1995
rect 2570 1965 2575 1985
rect 2595 1965 2600 1985
rect 2570 1935 2600 1965
rect 2570 1915 2575 1935
rect 2595 1915 2600 1935
rect 2570 1905 2600 1915
rect 2625 1985 2655 1995
rect 2625 1965 2630 1985
rect 2650 1965 2655 1985
rect 2625 1935 2655 1965
rect 2625 1915 2630 1935
rect 2650 1915 2655 1935
rect 2625 1905 2655 1915
rect 2680 1985 2710 1995
rect 2680 1965 2685 1985
rect 2705 1965 2710 1985
rect 2680 1935 2710 1965
rect 2680 1915 2685 1935
rect 2705 1915 2710 1935
rect 2680 1905 2710 1915
rect 2750 1985 2780 1995
rect 2750 1965 2755 1985
rect 2775 1965 2780 1985
rect 2750 1935 2780 1965
rect 2750 1915 2755 1935
rect 2775 1915 2780 1935
rect 2750 1905 2780 1915
rect 2810 1985 2840 1995
rect 2810 1965 2815 1985
rect 2835 1965 2840 1985
rect 2810 1935 2840 1965
rect 2810 1915 2815 1935
rect 2835 1915 2840 1935
rect 2810 1905 2840 1915
rect 2870 1985 2900 1995
rect 2870 1965 2875 1985
rect 2895 1965 2900 1985
rect 2870 1935 2900 1965
rect 2870 1915 2875 1935
rect 2895 1915 2900 1935
rect 2870 1905 2900 1915
rect 2930 1985 2960 1995
rect 2930 1965 2935 1985
rect 2955 1965 2960 1985
rect 2930 1935 2960 1965
rect 2930 1915 2935 1935
rect 2955 1915 2960 1935
rect 2930 1905 2960 1915
rect 2990 1985 3020 1995
rect 2990 1965 2995 1985
rect 3015 1965 3020 1985
rect 2990 1935 3020 1965
rect 2990 1915 2995 1935
rect 3015 1915 3020 1935
rect 2990 1905 3020 1915
rect 3050 1985 3080 1995
rect 3050 1965 3055 1985
rect 3075 1965 3080 1985
rect 3050 1935 3080 1965
rect 3050 1915 3055 1935
rect 3075 1915 3080 1935
rect 3050 1905 3080 1915
rect 3110 1985 3140 1995
rect 3110 1965 3115 1985
rect 3135 1965 3140 1985
rect 3110 1935 3140 1965
rect 3110 1915 3115 1935
rect 3135 1915 3140 1935
rect 3110 1905 3140 1915
rect 3170 1985 3200 1995
rect 3170 1965 3175 1985
rect 3195 1965 3200 1985
rect 3170 1935 3200 1965
rect 3170 1915 3175 1935
rect 3195 1915 3200 1935
rect 3170 1905 3200 1915
rect 3230 1985 3260 1995
rect 3230 1965 3235 1985
rect 3255 1965 3260 1985
rect 3230 1935 3260 1965
rect 3230 1915 3235 1935
rect 3255 1915 3260 1935
rect 3230 1905 3260 1915
rect 3290 1985 3320 1995
rect 3290 1965 3295 1985
rect 3315 1965 3320 1985
rect 3290 1935 3320 1965
rect 3290 1915 3295 1935
rect 3315 1915 3320 1935
rect 3290 1905 3320 1915
rect 3350 1985 3380 1995
rect 3350 1965 3355 1985
rect 3375 1965 3380 1985
rect 3350 1935 3380 1965
rect 3350 1915 3355 1935
rect 3375 1915 3380 1935
rect 3350 1905 3380 1915
rect 3410 1985 3440 1995
rect 3410 1965 3415 1985
rect 3435 1965 3440 1985
rect 3410 1935 3440 1965
rect 3410 1915 3415 1935
rect 3435 1915 3440 1935
rect 3410 1905 3440 1915
rect 3470 1985 3500 1995
rect 3470 1965 3475 1985
rect 3495 1965 3500 1985
rect 3470 1935 3500 1965
rect 3470 1915 3475 1935
rect 3495 1915 3500 1935
rect 3470 1905 3500 1915
rect 3530 1985 3560 1995
rect 3530 1965 3535 1985
rect 3555 1965 3560 1985
rect 3530 1935 3560 1965
rect 3530 1915 3535 1935
rect 3555 1915 3560 1935
rect 3530 1905 3560 1915
rect 3590 1985 3620 1995
rect 3590 1965 3595 1985
rect 3615 1965 3620 1985
rect 3590 1935 3620 1965
rect 3590 1915 3595 1935
rect 3615 1915 3620 1935
rect 3590 1905 3620 1915
rect 3650 1985 3680 1995
rect 3650 1965 3655 1985
rect 3675 1965 3680 1985
rect 3650 1935 3680 1965
rect 3650 1915 3655 1935
rect 3675 1915 3680 1935
rect 3650 1905 3680 1915
rect 3710 1985 3740 1995
rect 3710 1965 3715 1985
rect 3735 1965 3740 1985
rect 3710 1935 3740 1965
rect 3710 1915 3715 1935
rect 3735 1915 3740 1935
rect 3710 1905 3740 1915
rect 3770 1985 3800 1995
rect 3770 1965 3775 1985
rect 3795 1965 3800 1985
rect 3770 1935 3800 1965
rect 3770 1915 3775 1935
rect 3795 1915 3800 1935
rect 3770 1905 3800 1915
rect 3830 1985 3860 1995
rect 3830 1965 3835 1985
rect 3855 1965 3860 1985
rect 3830 1935 3860 1965
rect 3830 1915 3835 1935
rect 3855 1915 3860 1935
rect 3830 1905 3860 1915
rect 3890 1985 3920 1995
rect 3890 1965 3895 1985
rect 3915 1965 3920 1985
rect 3890 1935 3920 1965
rect 3890 1915 3895 1935
rect 3915 1915 3920 1935
rect 3890 1905 3920 1915
rect 3950 1985 4060 1995
rect 3950 1965 3955 1985
rect 3975 1965 3995 1985
rect 4015 1965 4035 1985
rect 4055 1965 4060 1985
rect 3950 1935 4060 1965
rect 3950 1915 3955 1935
rect 3975 1915 3995 1935
rect 4015 1915 4035 1935
rect 4055 1915 4060 1935
rect 3950 1905 4060 1915
rect 4090 1985 4120 1995
rect 4090 1965 4095 1985
rect 4115 1965 4120 1985
rect 4090 1935 4120 1965
rect 4090 1915 4095 1935
rect 4115 1915 4120 1935
rect 4090 1905 4120 1915
rect 4150 1985 4180 1995
rect 4150 1965 4155 1985
rect 4175 1965 4180 1985
rect 4150 1935 4180 1965
rect 4150 1915 4155 1935
rect 4175 1915 4180 1935
rect 4150 1905 4180 1915
rect 4210 1985 4240 1995
rect 4210 1965 4215 1985
rect 4235 1965 4240 1985
rect 4210 1935 4240 1965
rect 4210 1915 4215 1935
rect 4235 1915 4240 1935
rect 4210 1905 4240 1915
rect 4270 1985 4300 1995
rect 4270 1965 4275 1985
rect 4295 1965 4300 1985
rect 4270 1935 4300 1965
rect 4270 1915 4275 1935
rect 4295 1915 4300 1935
rect 4270 1905 4300 1915
rect 4330 1985 4360 1995
rect 4330 1965 4335 1985
rect 4355 1965 4360 1985
rect 4330 1935 4360 1965
rect 4330 1915 4335 1935
rect 4355 1915 4360 1935
rect 4330 1905 4360 1915
rect 4390 1985 4420 1995
rect 4390 1965 4395 1985
rect 4415 1965 4420 1985
rect 4390 1935 4420 1965
rect 4390 1915 4395 1935
rect 4415 1915 4420 1935
rect 4390 1905 4420 1915
rect 4450 1985 4480 1995
rect 4450 1965 4455 1985
rect 4475 1965 4480 1985
rect 4450 1935 4480 1965
rect 4450 1915 4455 1935
rect 4475 1915 4480 1935
rect 4450 1905 4480 1915
rect 4510 1985 4540 1995
rect 4510 1965 4515 1985
rect 4535 1965 4540 1985
rect 4510 1935 4540 1965
rect 4510 1915 4515 1935
rect 4535 1915 4540 1935
rect 4510 1905 4540 1915
rect 4570 1985 4600 1995
rect 4570 1965 4575 1985
rect 4595 1965 4600 1985
rect 4570 1935 4600 1965
rect 4570 1915 4575 1935
rect 4595 1915 4600 1935
rect 4570 1905 4600 1915
rect 4630 1985 4660 1995
rect 4630 1965 4635 1985
rect 4655 1965 4660 1985
rect 4630 1935 4660 1965
rect 4630 1915 4635 1935
rect 4655 1915 4660 1935
rect 4630 1905 4660 1915
rect 4690 1985 4720 1995
rect 4690 1965 4695 1985
rect 4715 1965 4720 1985
rect 4690 1935 4720 1965
rect 4690 1915 4695 1935
rect 4715 1915 4720 1935
rect 4690 1905 4720 1915
rect 4750 1985 4780 1995
rect 4750 1965 4755 1985
rect 4775 1965 4780 1985
rect 4750 1935 4780 1965
rect 4750 1915 4755 1935
rect 4775 1915 4780 1935
rect 4750 1905 4780 1915
rect 4810 1985 4840 1995
rect 4810 1965 4815 1985
rect 4835 1965 4840 1985
rect 4810 1935 4840 1965
rect 4810 1915 4815 1935
rect 4835 1915 4840 1935
rect 4810 1905 4840 1915
rect 4870 1985 4900 1995
rect 4870 1965 4875 1985
rect 4895 1965 4900 1985
rect 4870 1935 4900 1965
rect 4870 1915 4875 1935
rect 4895 1915 4900 1935
rect 4870 1905 4900 1915
rect 4930 1985 4960 1995
rect 4930 1965 4935 1985
rect 4955 1965 4960 1985
rect 4930 1935 4960 1965
rect 4930 1915 4935 1935
rect 4955 1915 4960 1935
rect 4930 1905 4960 1915
rect 4990 1985 5020 1995
rect 4990 1965 4995 1985
rect 5015 1965 5020 1985
rect 4990 1935 5020 1965
rect 4990 1915 4995 1935
rect 5015 1915 5020 1935
rect 4990 1905 5020 1915
rect 5050 1985 5080 1995
rect 5050 1965 5055 1985
rect 5075 1965 5080 1985
rect 5050 1935 5080 1965
rect 5050 1915 5055 1935
rect 5075 1915 5080 1935
rect 5050 1905 5080 1915
rect 5110 1985 5140 1995
rect 5110 1965 5115 1985
rect 5135 1965 5140 1985
rect 5110 1935 5140 1965
rect 5110 1915 5115 1935
rect 5135 1915 5140 1935
rect 5110 1905 5140 1915
rect 5170 1985 5200 1995
rect 5170 1965 5175 1985
rect 5195 1965 5200 1985
rect 5170 1935 5200 1965
rect 5170 1915 5175 1935
rect 5195 1915 5200 1935
rect 5170 1905 5200 1915
rect 5230 1985 5260 1995
rect 5230 1965 5235 1985
rect 5255 1965 5260 1985
rect 5230 1935 5260 1965
rect 5230 1915 5235 1935
rect 5255 1915 5260 1935
rect 5230 1905 5260 1915
rect 2575 1885 2595 1905
rect 2685 1885 2705 1905
rect 2755 1885 2775 1905
rect 2935 1885 2955 1905
rect 3055 1885 3075 1905
rect 3295 1885 3315 1905
rect 3415 1885 3435 1905
rect 3655 1885 3675 1905
rect 3775 1885 3795 1905
rect 2565 1875 2600 1885
rect 2565 1855 2575 1875
rect 2595 1855 2600 1875
rect 2565 1845 2600 1855
rect 2620 1875 2660 1885
rect 2620 1855 2630 1875
rect 2650 1855 2660 1875
rect 2620 1845 2660 1855
rect 2680 1875 2715 1885
rect 2680 1855 2685 1875
rect 2705 1855 2715 1875
rect 2680 1845 2715 1855
rect 2755 1875 2805 1885
rect 2755 1855 2775 1875
rect 2795 1855 2805 1875
rect 2755 1845 2805 1855
rect 2835 1875 2875 1885
rect 2835 1855 2845 1875
rect 2865 1855 2875 1875
rect 2835 1845 2875 1855
rect 2925 1875 2965 1885
rect 2925 1855 2935 1875
rect 2955 1855 2965 1875
rect 2925 1845 2965 1855
rect 3045 1875 3085 1885
rect 3045 1855 3055 1875
rect 3075 1855 3085 1875
rect 3045 1845 3085 1855
rect 3165 1875 3205 1885
rect 3165 1855 3175 1875
rect 3195 1855 3205 1875
rect 3165 1845 3205 1855
rect 3285 1875 3325 1885
rect 3285 1855 3295 1875
rect 3315 1855 3325 1875
rect 3285 1845 3325 1855
rect 3405 1875 3445 1885
rect 3405 1855 3415 1875
rect 3435 1855 3445 1875
rect 3405 1845 3445 1855
rect 3525 1875 3565 1885
rect 3525 1855 3535 1875
rect 3555 1855 3565 1875
rect 3525 1845 3565 1855
rect 3645 1875 3685 1885
rect 3645 1855 3655 1875
rect 3675 1855 3685 1875
rect 3645 1845 3685 1855
rect 3765 1875 3805 1885
rect 3765 1855 3775 1875
rect 3795 1855 3805 1875
rect 3765 1845 3805 1855
rect 3855 1875 3895 1885
rect 3995 1880 4015 1905
rect 4215 1885 4235 1905
rect 4335 1885 4355 1905
rect 4575 1885 4595 1905
rect 4695 1885 4715 1905
rect 4935 1885 4955 1905
rect 5055 1885 5075 1905
rect 5235 1885 5255 1905
rect 3855 1855 3865 1875
rect 3885 1855 3895 1875
rect 3855 1845 3895 1855
rect 3985 1870 4025 1880
rect 3985 1850 3995 1870
rect 4015 1850 4025 1870
rect 3985 1840 4025 1850
rect 4115 1875 4155 1885
rect 4115 1855 4125 1875
rect 4145 1855 4155 1875
rect 4115 1845 4155 1855
rect 4205 1875 4245 1885
rect 4205 1855 4215 1875
rect 4235 1855 4245 1875
rect 4205 1845 4245 1855
rect 4325 1875 4365 1885
rect 4325 1855 4335 1875
rect 4355 1855 4365 1875
rect 4325 1845 4365 1855
rect 4445 1875 4485 1885
rect 4445 1855 4455 1875
rect 4475 1855 4485 1875
rect 4445 1845 4485 1855
rect 4565 1875 4605 1885
rect 4565 1855 4575 1875
rect 4595 1855 4605 1875
rect 4565 1845 4605 1855
rect 4685 1875 4725 1885
rect 4685 1855 4695 1875
rect 4715 1855 4725 1875
rect 4685 1845 4725 1855
rect 4805 1875 4845 1885
rect 4805 1855 4815 1875
rect 4835 1855 4845 1875
rect 4805 1845 4845 1855
rect 4925 1875 4965 1885
rect 4925 1855 4935 1875
rect 4955 1855 4965 1875
rect 4925 1845 4965 1855
rect 5045 1875 5085 1885
rect 5045 1855 5055 1875
rect 5075 1855 5085 1875
rect 5045 1845 5085 1855
rect 5135 1875 5175 1885
rect 5135 1855 5145 1875
rect 5165 1855 5175 1875
rect 5135 1845 5175 1855
rect 5205 1875 5255 1885
rect 5205 1855 5215 1875
rect 5235 1855 5255 1875
rect 5205 1845 5255 1855
rect 2475 1790 2505 1820
rect 2835 1785 2875 1825
rect 3045 1815 3085 1825
rect 3045 1795 3055 1815
rect 3075 1795 3085 1815
rect 3045 1785 3085 1795
rect 3165 1785 3205 1825
rect 3405 1815 3445 1825
rect 3405 1795 3415 1815
rect 3435 1795 3445 1815
rect 3405 1785 3445 1795
rect 3525 1785 3565 1825
rect 3765 1815 3805 1825
rect 3765 1795 3775 1815
rect 3795 1795 3805 1815
rect 3765 1785 3805 1795
rect 3855 1785 3895 1825
rect 4115 1785 4155 1825
rect 4205 1815 4245 1825
rect 4205 1795 4215 1815
rect 4235 1795 4245 1815
rect 4205 1785 4245 1795
rect 4445 1785 4485 1825
rect 4565 1815 4605 1825
rect 4565 1795 4575 1815
rect 4595 1795 4605 1815
rect 4565 1785 4605 1795
rect 4805 1785 4845 1825
rect 4925 1815 4965 1825
rect 4925 1795 4935 1815
rect 4955 1795 4965 1815
rect 4925 1785 4965 1795
rect 5135 1785 5175 1825
rect 11190 1820 11230 1830
rect 5365 1790 5395 1820
rect 11085 1805 11125 1815
rect 11085 1785 11095 1805
rect 11115 1785 11125 1805
rect 11190 1800 11200 1820
rect 11220 1800 11230 1820
rect 11410 1820 11450 1830
rect 11190 1790 11230 1800
rect 11305 1805 11345 1815
rect 11085 1775 11125 1785
rect 2430 1730 2460 1760
rect 2570 1730 2600 1760
rect 2680 1730 2710 1760
rect 2805 1735 2835 1765
rect 3225 1755 3265 1765
rect 3225 1735 3235 1755
rect 3255 1735 3265 1755
rect 3225 1725 3265 1735
rect 3285 1755 3325 1765
rect 3285 1735 3295 1755
rect 3315 1735 3325 1755
rect 3285 1725 3325 1735
rect 3525 1755 3565 1765
rect 3525 1735 3535 1755
rect 3555 1735 3565 1755
rect 3525 1725 3565 1735
rect 3765 1755 3805 1765
rect 3765 1735 3775 1755
rect 3795 1735 3805 1755
rect 3765 1725 3805 1735
rect 4205 1755 4245 1765
rect 4205 1735 4215 1755
rect 4235 1735 4245 1755
rect 4205 1725 4245 1735
rect 4445 1755 4485 1765
rect 4445 1735 4455 1755
rect 4475 1735 4485 1755
rect 4445 1725 4485 1735
rect 4685 1755 4725 1765
rect 4685 1735 4695 1755
rect 4715 1735 4725 1755
rect 4685 1725 4725 1735
rect 4745 1755 4785 1765
rect 4745 1735 4755 1755
rect 4775 1735 4785 1755
rect 4745 1725 4785 1735
rect 5275 1730 5305 1760
rect 3165 1710 3205 1720
rect 2805 1680 2835 1710
rect 3165 1690 3175 1710
rect 3195 1690 3205 1710
rect 3165 1680 3205 1690
rect 2385 1635 2415 1665
rect 2625 1635 2655 1665
rect 3175 1660 3195 1680
rect 3295 1660 3315 1725
rect 3405 1710 3445 1720
rect 3405 1690 3415 1710
rect 3435 1690 3445 1710
rect 3405 1680 3445 1690
rect 3415 1660 3435 1680
rect 3535 1660 3555 1725
rect 3645 1710 3685 1720
rect 3645 1690 3655 1710
rect 3675 1690 3685 1710
rect 3645 1680 3685 1690
rect 3655 1660 3675 1680
rect 3775 1660 3795 1725
rect 4215 1660 4235 1725
rect 4325 1710 4365 1720
rect 4325 1690 4335 1710
rect 4355 1690 4365 1710
rect 4325 1680 4365 1690
rect 4335 1660 4355 1680
rect 4455 1660 4475 1725
rect 4565 1710 4605 1720
rect 4565 1690 4575 1710
rect 4595 1690 4605 1710
rect 4565 1680 4605 1690
rect 4575 1660 4595 1680
rect 4695 1660 4715 1725
rect 4805 1710 4845 1720
rect 11095 1710 11115 1775
rect 11200 1710 11220 1790
rect 11305 1785 11315 1805
rect 11335 1785 11345 1805
rect 11410 1800 11420 1820
rect 11440 1800 11450 1820
rect 11640 1820 11680 1830
rect 11410 1790 11450 1800
rect 11525 1805 11565 1815
rect 11305 1775 11345 1785
rect 11237 1760 11269 1770
rect 11237 1740 11243 1760
rect 11260 1740 11269 1760
rect 11237 1730 11269 1740
rect 11315 1710 11335 1775
rect 11420 1710 11440 1790
rect 11525 1785 11535 1805
rect 11555 1785 11565 1805
rect 11640 1800 11650 1820
rect 11670 1800 11680 1820
rect 12230 1820 12270 1830
rect 11640 1790 11680 1800
rect 12125 1805 12165 1815
rect 11525 1775 11565 1785
rect 11457 1760 11489 1770
rect 11457 1740 11463 1760
rect 11480 1740 11489 1760
rect 11457 1730 11489 1740
rect 11535 1710 11555 1775
rect 11601 1760 11633 1770
rect 11601 1740 11610 1760
rect 11627 1740 11633 1760
rect 11601 1730 11633 1740
rect 11650 1710 11670 1790
rect 12125 1785 12135 1805
rect 12155 1785 12165 1805
rect 12230 1800 12240 1820
rect 12260 1800 12270 1820
rect 12450 1820 12490 1830
rect 12230 1790 12270 1800
rect 12345 1805 12385 1815
rect 12125 1775 12165 1785
rect 11820 1760 11850 1770
rect 11820 1740 11825 1760
rect 11845 1740 11850 1760
rect 11820 1730 11850 1740
rect 11867 1760 11899 1770
rect 11867 1740 11876 1760
rect 11893 1740 11899 1760
rect 11867 1730 11899 1740
rect 11950 1760 11980 1770
rect 11950 1740 11955 1760
rect 11975 1740 11980 1760
rect 11950 1730 11980 1740
rect 11830 1710 11850 1730
rect 11950 1710 11970 1730
rect 12135 1710 12155 1775
rect 12240 1710 12260 1790
rect 12345 1785 12355 1805
rect 12375 1785 12385 1805
rect 12450 1800 12460 1820
rect 12480 1800 12490 1820
rect 12680 1820 12720 1830
rect 12450 1790 12490 1800
rect 12565 1805 12605 1815
rect 12345 1775 12385 1785
rect 12277 1760 12309 1770
rect 12277 1740 12283 1760
rect 12300 1740 12309 1760
rect 12277 1730 12309 1740
rect 12355 1710 12375 1775
rect 12460 1710 12480 1790
rect 12565 1785 12575 1805
rect 12595 1785 12605 1805
rect 12680 1800 12690 1820
rect 12710 1800 12720 1820
rect 12680 1790 12720 1800
rect 12565 1775 12605 1785
rect 12497 1760 12529 1770
rect 12497 1740 12503 1760
rect 12520 1740 12529 1760
rect 12497 1730 12529 1740
rect 12575 1710 12595 1775
rect 12641 1760 12673 1770
rect 12641 1740 12650 1760
rect 12667 1740 12673 1760
rect 12641 1730 12673 1740
rect 12690 1710 12710 1790
rect 4805 1690 4815 1710
rect 4835 1690 4845 1710
rect 4805 1680 4845 1690
rect 10990 1700 11065 1710
rect 10990 1680 11000 1700
rect 11020 1680 11040 1700
rect 11060 1680 11065 1700
rect 4815 1660 4835 1680
rect 3170 1650 3200 1660
rect 3170 1630 3175 1650
rect 3195 1630 3200 1650
rect 3170 1620 3200 1630
rect 3230 1650 3260 1660
rect 3230 1630 3235 1650
rect 3255 1630 3260 1650
rect 3230 1620 3260 1630
rect 3290 1650 3320 1660
rect 3290 1630 3295 1650
rect 3315 1630 3320 1650
rect 3290 1620 3320 1630
rect 3350 1650 3380 1660
rect 3350 1630 3355 1650
rect 3375 1630 3380 1650
rect 3350 1620 3380 1630
rect 3410 1650 3440 1660
rect 3410 1630 3415 1650
rect 3435 1630 3440 1650
rect 3410 1620 3440 1630
rect 3470 1650 3500 1660
rect 3470 1630 3475 1650
rect 3495 1630 3500 1650
rect 3470 1620 3500 1630
rect 3530 1650 3560 1660
rect 3530 1630 3535 1650
rect 3555 1630 3560 1650
rect 3530 1620 3560 1630
rect 3590 1650 3620 1660
rect 3590 1630 3595 1650
rect 3615 1630 3620 1650
rect 3590 1620 3620 1630
rect 3650 1650 3680 1660
rect 3650 1630 3655 1650
rect 3675 1630 3680 1650
rect 3650 1620 3680 1630
rect 3710 1650 3740 1660
rect 3710 1630 3715 1650
rect 3735 1630 3740 1650
rect 3710 1620 3740 1630
rect 3770 1650 3800 1660
rect 3770 1630 3775 1650
rect 3795 1630 3800 1650
rect 3770 1620 3800 1630
rect 3985 1650 4025 1660
rect 3985 1630 3995 1650
rect 4015 1630 4025 1650
rect 3985 1620 4025 1630
rect 4210 1650 4240 1660
rect 4210 1630 4215 1650
rect 4235 1630 4240 1650
rect 4210 1620 4240 1630
rect 4270 1650 4300 1660
rect 4270 1630 4275 1650
rect 4295 1630 4300 1650
rect 4270 1620 4300 1630
rect 4330 1650 4360 1660
rect 4330 1630 4335 1650
rect 4355 1630 4360 1650
rect 4330 1620 4360 1630
rect 4390 1650 4420 1660
rect 4390 1630 4395 1650
rect 4415 1630 4420 1650
rect 4390 1620 4420 1630
rect 4450 1650 4480 1660
rect 4450 1630 4455 1650
rect 4475 1630 4480 1650
rect 4450 1620 4480 1630
rect 4510 1650 4540 1660
rect 4510 1630 4515 1650
rect 4535 1630 4540 1650
rect 4510 1620 4540 1630
rect 4570 1650 4600 1660
rect 4570 1630 4575 1650
rect 4595 1630 4600 1650
rect 4570 1620 4600 1630
rect 4630 1650 4660 1660
rect 4630 1630 4635 1650
rect 4655 1630 4660 1650
rect 4630 1620 4660 1630
rect 4690 1650 4720 1660
rect 4690 1630 4695 1650
rect 4715 1630 4720 1650
rect 4690 1620 4720 1630
rect 4750 1650 4780 1660
rect 4750 1630 4755 1650
rect 4775 1630 4780 1650
rect 4750 1620 4780 1630
rect 4810 1650 4840 1660
rect 4810 1630 4815 1650
rect 4835 1630 4840 1650
rect 4810 1620 4840 1630
rect 10990 1650 11065 1680
rect 10990 1630 11000 1650
rect 11020 1630 11040 1650
rect 11060 1630 11065 1650
rect 2335 1565 2365 1595
rect 3165 1590 3205 1600
rect 3165 1570 3175 1590
rect 3195 1570 3205 1590
rect 3165 1560 3205 1570
rect 3235 1550 3255 1620
rect 3355 1550 3375 1620
rect 3475 1550 3495 1620
rect 3595 1550 3615 1620
rect 3715 1550 3735 1620
rect 4275 1550 4295 1620
rect 4395 1550 4415 1620
rect 4515 1550 4535 1620
rect 4635 1550 4655 1620
rect 4755 1550 4775 1620
rect 10990 1600 11065 1630
rect 4805 1590 4845 1600
rect 4805 1570 4815 1590
rect 4835 1570 4845 1590
rect 4805 1560 4845 1570
rect 5415 1565 5445 1595
rect 10990 1580 11000 1600
rect 11020 1580 11040 1600
rect 11060 1580 11065 1600
rect 10990 1570 11065 1580
rect 11090 1700 11120 1710
rect 11090 1680 11095 1700
rect 11115 1680 11120 1700
rect 11090 1650 11120 1680
rect 11090 1630 11095 1650
rect 11115 1630 11120 1650
rect 11090 1600 11120 1630
rect 11090 1580 11095 1600
rect 11115 1580 11120 1600
rect 11090 1570 11120 1580
rect 11145 1700 11175 1710
rect 11145 1680 11150 1700
rect 11170 1680 11175 1700
rect 11145 1650 11175 1680
rect 11145 1630 11150 1650
rect 11170 1630 11175 1650
rect 11145 1600 11175 1630
rect 11145 1580 11150 1600
rect 11170 1580 11175 1600
rect 11145 1570 11175 1580
rect 11200 1700 11230 1710
rect 11200 1680 11205 1700
rect 11225 1680 11230 1700
rect 11200 1650 11230 1680
rect 11200 1630 11205 1650
rect 11225 1630 11230 1650
rect 11200 1600 11230 1630
rect 11200 1580 11205 1600
rect 11225 1580 11230 1600
rect 11200 1570 11230 1580
rect 11255 1700 11285 1710
rect 11255 1680 11260 1700
rect 11280 1680 11285 1700
rect 11255 1650 11285 1680
rect 11255 1630 11260 1650
rect 11280 1630 11285 1650
rect 11255 1600 11285 1630
rect 11255 1580 11260 1600
rect 11280 1580 11285 1600
rect 11255 1570 11285 1580
rect 11310 1700 11340 1710
rect 11310 1680 11315 1700
rect 11335 1680 11340 1700
rect 11310 1650 11340 1680
rect 11310 1630 11315 1650
rect 11335 1630 11340 1650
rect 11310 1600 11340 1630
rect 11310 1580 11315 1600
rect 11335 1580 11340 1600
rect 11310 1570 11340 1580
rect 11365 1700 11395 1710
rect 11365 1680 11370 1700
rect 11390 1680 11395 1700
rect 11365 1650 11395 1680
rect 11365 1630 11370 1650
rect 11390 1630 11395 1650
rect 11365 1600 11395 1630
rect 11365 1580 11370 1600
rect 11390 1580 11395 1600
rect 11365 1570 11395 1580
rect 11420 1700 11450 1710
rect 11420 1680 11425 1700
rect 11445 1680 11450 1700
rect 11420 1650 11450 1680
rect 11420 1630 11425 1650
rect 11445 1630 11450 1650
rect 11420 1600 11450 1630
rect 11420 1580 11425 1600
rect 11445 1580 11450 1600
rect 11420 1570 11450 1580
rect 11475 1700 11505 1710
rect 11475 1680 11480 1700
rect 11500 1680 11505 1700
rect 11475 1650 11505 1680
rect 11475 1630 11480 1650
rect 11500 1630 11505 1650
rect 11475 1600 11505 1630
rect 11475 1580 11480 1600
rect 11500 1580 11505 1600
rect 11475 1570 11505 1580
rect 11530 1700 11560 1710
rect 11530 1680 11535 1700
rect 11555 1680 11560 1700
rect 11530 1650 11560 1680
rect 11530 1630 11535 1650
rect 11555 1630 11560 1650
rect 11530 1600 11560 1630
rect 11530 1580 11535 1600
rect 11555 1580 11560 1600
rect 11530 1570 11560 1580
rect 11585 1700 11615 1710
rect 11585 1680 11590 1700
rect 11610 1680 11615 1700
rect 11585 1650 11615 1680
rect 11585 1630 11590 1650
rect 11610 1630 11615 1650
rect 11585 1600 11615 1630
rect 11585 1580 11590 1600
rect 11610 1580 11615 1600
rect 11585 1570 11615 1580
rect 11640 1700 11670 1710
rect 11640 1680 11645 1700
rect 11665 1680 11670 1700
rect 11640 1650 11670 1680
rect 11640 1630 11645 1650
rect 11665 1630 11670 1650
rect 11640 1600 11670 1630
rect 11640 1580 11645 1600
rect 11665 1580 11670 1600
rect 11640 1570 11670 1580
rect 11695 1700 11805 1710
rect 11695 1680 11700 1700
rect 11720 1680 11740 1700
rect 11760 1680 11780 1700
rect 11800 1680 11805 1700
rect 11695 1650 11805 1680
rect 11695 1630 11700 1650
rect 11720 1630 11740 1650
rect 11760 1630 11780 1650
rect 11800 1630 11805 1650
rect 11695 1600 11805 1630
rect 11695 1580 11700 1600
rect 11720 1580 11740 1600
rect 11760 1580 11780 1600
rect 11800 1580 11805 1600
rect 11695 1570 11805 1580
rect 11830 1700 11860 1710
rect 11830 1680 11835 1700
rect 11855 1680 11860 1700
rect 11830 1650 11860 1680
rect 11830 1630 11835 1650
rect 11855 1630 11860 1650
rect 11830 1600 11860 1630
rect 11830 1580 11835 1600
rect 11855 1580 11860 1600
rect 11830 1570 11860 1580
rect 11885 1700 11915 1710
rect 11885 1680 11890 1700
rect 11910 1680 11915 1700
rect 11885 1650 11915 1680
rect 11885 1630 11890 1650
rect 11910 1630 11915 1650
rect 11885 1600 11915 1630
rect 11885 1580 11890 1600
rect 11910 1580 11915 1600
rect 11885 1570 11915 1580
rect 11940 1700 11970 1710
rect 11940 1680 11945 1700
rect 11965 1680 11970 1700
rect 11940 1650 11970 1680
rect 11940 1630 11945 1650
rect 11965 1630 11970 1650
rect 11940 1600 11970 1630
rect 11940 1580 11945 1600
rect 11965 1580 11970 1600
rect 11940 1570 11970 1580
rect 11995 1700 12105 1710
rect 11995 1680 12000 1700
rect 12020 1680 12040 1700
rect 12060 1680 12080 1700
rect 12100 1680 12105 1700
rect 11995 1650 12105 1680
rect 11995 1630 12000 1650
rect 12020 1630 12040 1650
rect 12060 1630 12080 1650
rect 12100 1630 12105 1650
rect 11995 1600 12105 1630
rect 11995 1580 12000 1600
rect 12020 1580 12040 1600
rect 12060 1580 12080 1600
rect 12100 1580 12105 1600
rect 11995 1570 12105 1580
rect 12130 1700 12160 1710
rect 12130 1680 12135 1700
rect 12155 1680 12160 1700
rect 12130 1650 12160 1680
rect 12130 1630 12135 1650
rect 12155 1630 12160 1650
rect 12130 1600 12160 1630
rect 12130 1580 12135 1600
rect 12155 1580 12160 1600
rect 12130 1570 12160 1580
rect 12185 1700 12215 1710
rect 12185 1680 12190 1700
rect 12210 1680 12215 1700
rect 12185 1650 12215 1680
rect 12185 1630 12190 1650
rect 12210 1630 12215 1650
rect 12185 1600 12215 1630
rect 12185 1580 12190 1600
rect 12210 1580 12215 1600
rect 12185 1570 12215 1580
rect 12240 1700 12270 1710
rect 12240 1680 12245 1700
rect 12265 1680 12270 1700
rect 12240 1650 12270 1680
rect 12240 1630 12245 1650
rect 12265 1630 12270 1650
rect 12240 1600 12270 1630
rect 12240 1580 12245 1600
rect 12265 1580 12270 1600
rect 12240 1570 12270 1580
rect 12295 1700 12325 1710
rect 12295 1680 12300 1700
rect 12320 1680 12325 1700
rect 12295 1650 12325 1680
rect 12295 1630 12300 1650
rect 12320 1630 12325 1650
rect 12295 1600 12325 1630
rect 12295 1580 12300 1600
rect 12320 1580 12325 1600
rect 12295 1570 12325 1580
rect 12350 1700 12380 1710
rect 12350 1680 12355 1700
rect 12375 1680 12380 1700
rect 12350 1650 12380 1680
rect 12350 1630 12355 1650
rect 12375 1630 12380 1650
rect 12350 1600 12380 1630
rect 12350 1580 12355 1600
rect 12375 1580 12380 1600
rect 12350 1570 12380 1580
rect 12405 1700 12435 1710
rect 12405 1680 12410 1700
rect 12430 1680 12435 1700
rect 12405 1650 12435 1680
rect 12405 1630 12410 1650
rect 12430 1630 12435 1650
rect 12405 1600 12435 1630
rect 12405 1580 12410 1600
rect 12430 1580 12435 1600
rect 12405 1570 12435 1580
rect 12460 1700 12490 1710
rect 12460 1680 12465 1700
rect 12485 1680 12490 1700
rect 12460 1650 12490 1680
rect 12460 1630 12465 1650
rect 12485 1630 12490 1650
rect 12460 1600 12490 1630
rect 12460 1580 12465 1600
rect 12485 1580 12490 1600
rect 12460 1570 12490 1580
rect 12515 1700 12545 1710
rect 12515 1680 12520 1700
rect 12540 1680 12545 1700
rect 12515 1650 12545 1680
rect 12515 1630 12520 1650
rect 12540 1630 12545 1650
rect 12515 1600 12545 1630
rect 12515 1580 12520 1600
rect 12540 1580 12545 1600
rect 12515 1570 12545 1580
rect 12570 1700 12600 1710
rect 12570 1680 12575 1700
rect 12595 1680 12600 1700
rect 12570 1650 12600 1680
rect 12570 1630 12575 1650
rect 12595 1630 12600 1650
rect 12570 1600 12600 1630
rect 12570 1580 12575 1600
rect 12595 1580 12600 1600
rect 12570 1570 12600 1580
rect 12625 1700 12655 1710
rect 12625 1680 12630 1700
rect 12650 1680 12655 1700
rect 12625 1650 12655 1680
rect 12625 1630 12630 1650
rect 12650 1630 12655 1650
rect 12625 1600 12655 1630
rect 12625 1580 12630 1600
rect 12650 1580 12655 1600
rect 12625 1570 12655 1580
rect 12680 1700 12710 1710
rect 12680 1680 12685 1700
rect 12705 1680 12710 1700
rect 12680 1650 12710 1680
rect 12680 1630 12685 1650
rect 12705 1630 12710 1650
rect 12680 1600 12710 1630
rect 12680 1580 12685 1600
rect 12705 1580 12710 1600
rect 12680 1570 12710 1580
rect 12735 1700 12810 1710
rect 12735 1680 12740 1700
rect 12760 1680 12780 1700
rect 12800 1680 12810 1700
rect 12735 1650 12810 1680
rect 12735 1630 12740 1650
rect 12760 1630 12780 1650
rect 12800 1630 12810 1650
rect 12735 1600 12810 1630
rect 12735 1580 12740 1600
rect 12760 1580 12780 1600
rect 12800 1580 12810 1600
rect 12735 1570 12810 1580
rect 11000 1550 11020 1570
rect 3225 1540 3265 1550
rect 3225 1520 3235 1540
rect 3255 1520 3265 1540
rect 3225 1510 3265 1520
rect 3345 1540 3385 1550
rect 3345 1520 3355 1540
rect 3375 1520 3385 1540
rect 3345 1510 3385 1520
rect 3465 1540 3505 1550
rect 3465 1520 3475 1540
rect 3495 1520 3505 1540
rect 3465 1510 3505 1520
rect 3585 1540 3625 1550
rect 3585 1520 3595 1540
rect 3615 1520 3625 1540
rect 3585 1510 3625 1520
rect 3705 1540 3745 1550
rect 3705 1520 3715 1540
rect 3735 1520 3745 1540
rect 3705 1510 3745 1520
rect 4265 1540 4305 1550
rect 4265 1520 4275 1540
rect 4295 1520 4305 1540
rect 4265 1510 4305 1520
rect 4385 1540 4425 1550
rect 4385 1520 4395 1540
rect 4415 1520 4425 1540
rect 4385 1510 4425 1520
rect 4505 1540 4545 1550
rect 4505 1520 4515 1540
rect 4535 1520 4545 1540
rect 4505 1510 4545 1520
rect 4625 1540 4665 1550
rect 4625 1520 4635 1540
rect 4655 1520 4665 1540
rect 4625 1510 4665 1520
rect 4745 1540 4785 1550
rect 4745 1520 4755 1540
rect 4775 1520 4785 1540
rect 4745 1510 4785 1520
rect 10990 1540 11030 1550
rect 10990 1520 11000 1540
rect 11020 1520 11030 1540
rect 10990 1510 11030 1520
rect 11106 1540 11138 1550
rect 11106 1520 11112 1540
rect 11129 1520 11138 1540
rect 11106 1510 11138 1520
rect 2925 1495 2965 1505
rect 2835 1480 2875 1490
rect 2835 1460 2845 1480
rect 2865 1460 2875 1480
rect 2925 1475 2935 1495
rect 2955 1475 2965 1495
rect 2925 1465 2965 1475
rect 3045 1495 3085 1505
rect 3045 1475 3055 1495
rect 3075 1475 3085 1495
rect 3045 1465 3085 1475
rect 3165 1495 3205 1505
rect 3165 1475 3175 1495
rect 3195 1475 3205 1495
rect 3165 1465 3205 1475
rect 3285 1495 3325 1505
rect 3285 1475 3295 1495
rect 3315 1475 3325 1495
rect 3285 1465 3325 1475
rect 3525 1495 3565 1505
rect 3525 1475 3535 1495
rect 3555 1475 3565 1495
rect 3525 1465 3565 1475
rect 3645 1495 3685 1505
rect 3645 1475 3655 1495
rect 3675 1475 3685 1495
rect 3645 1465 3685 1475
rect 3765 1495 3805 1505
rect 3765 1475 3775 1495
rect 3795 1475 3805 1495
rect 4205 1495 4245 1505
rect 3765 1465 3805 1475
rect 3915 1480 3955 1490
rect 2835 1450 2875 1460
rect 3915 1460 3925 1480
rect 3945 1460 3955 1480
rect 3915 1450 3955 1460
rect 4055 1480 4095 1490
rect 4055 1460 4065 1480
rect 4085 1460 4095 1480
rect 4205 1475 4215 1495
rect 4235 1475 4245 1495
rect 4205 1465 4245 1475
rect 4325 1495 4365 1505
rect 4325 1475 4335 1495
rect 4355 1475 4365 1495
rect 4325 1465 4365 1475
rect 4445 1495 4485 1505
rect 4445 1475 4455 1495
rect 4475 1475 4485 1495
rect 4445 1465 4485 1475
rect 4685 1495 4725 1505
rect 4685 1475 4695 1495
rect 4715 1475 4725 1495
rect 4685 1465 4725 1475
rect 4805 1495 4845 1505
rect 4805 1475 4815 1495
rect 4835 1475 4845 1495
rect 4805 1465 4845 1475
rect 4925 1495 4965 1505
rect 4925 1475 4935 1495
rect 4955 1475 4965 1495
rect 4925 1465 4965 1475
rect 5045 1495 5085 1505
rect 5045 1475 5055 1495
rect 5075 1475 5085 1495
rect 11155 1490 11175 1570
rect 11260 1490 11280 1570
rect 11305 1540 11345 1550
rect 11305 1520 11315 1540
rect 11335 1520 11345 1540
rect 11305 1510 11345 1520
rect 11370 1490 11390 1570
rect 11480 1490 11500 1570
rect 11525 1540 11565 1550
rect 11525 1520 11535 1540
rect 11555 1520 11565 1540
rect 11525 1510 11565 1520
rect 11590 1490 11610 1570
rect 11740 1550 11760 1570
rect 11830 1550 11850 1570
rect 11885 1550 11905 1570
rect 12040 1550 12060 1570
rect 11730 1540 11770 1550
rect 11730 1520 11740 1540
rect 11760 1520 11770 1540
rect 11730 1510 11770 1520
rect 11825 1540 11855 1550
rect 11825 1520 11830 1540
rect 11850 1520 11855 1540
rect 11825 1510 11855 1520
rect 11875 1540 11905 1550
rect 11875 1520 11880 1540
rect 11900 1520 11905 1540
rect 11875 1510 11905 1520
rect 11922 1540 11954 1550
rect 11922 1520 11928 1540
rect 11945 1520 11954 1540
rect 11922 1510 11954 1520
rect 12030 1540 12070 1550
rect 12030 1520 12040 1540
rect 12060 1520 12070 1540
rect 12030 1510 12070 1520
rect 12146 1540 12178 1550
rect 12146 1520 12152 1540
rect 12169 1520 12178 1540
rect 12146 1510 12178 1520
rect 12195 1490 12215 1570
rect 12300 1490 12320 1570
rect 12345 1540 12385 1550
rect 12345 1520 12355 1540
rect 12375 1520 12385 1540
rect 12345 1510 12385 1520
rect 12410 1490 12430 1570
rect 12520 1490 12540 1570
rect 12565 1540 12605 1550
rect 12565 1520 12575 1540
rect 12595 1520 12605 1540
rect 12565 1510 12605 1520
rect 12630 1490 12650 1570
rect 12780 1550 12800 1570
rect 12770 1540 12810 1550
rect 12770 1520 12780 1540
rect 12800 1520 12810 1540
rect 12770 1510 12810 1520
rect 5045 1465 5085 1475
rect 5135 1480 5175 1490
rect 4055 1450 4095 1460
rect 5135 1460 5145 1480
rect 5165 1460 5175 1480
rect 5135 1450 5175 1460
rect 11145 1480 11185 1490
rect 11145 1460 11155 1480
rect 11175 1460 11185 1480
rect 11145 1450 11185 1460
rect 11250 1480 11290 1490
rect 11250 1460 11260 1480
rect 11280 1460 11290 1480
rect 11250 1450 11290 1460
rect 11360 1480 11400 1490
rect 11360 1460 11370 1480
rect 11390 1460 11400 1480
rect 11360 1450 11400 1460
rect 11470 1480 11510 1490
rect 11470 1460 11480 1480
rect 11500 1460 11510 1480
rect 11470 1450 11510 1460
rect 11580 1480 11620 1490
rect 11580 1460 11590 1480
rect 11610 1460 11620 1480
rect 11580 1450 11620 1460
rect 12185 1480 12225 1490
rect 12185 1460 12195 1480
rect 12215 1460 12225 1480
rect 12185 1450 12225 1460
rect 12290 1480 12330 1490
rect 12290 1460 12300 1480
rect 12320 1460 12330 1480
rect 12290 1450 12330 1460
rect 12400 1480 12440 1490
rect 12400 1460 12410 1480
rect 12430 1460 12440 1480
rect 12400 1450 12440 1460
rect 12510 1480 12550 1490
rect 12510 1460 12520 1480
rect 12540 1460 12550 1480
rect 12510 1450 12550 1460
rect 12620 1480 12660 1490
rect 12620 1460 12630 1480
rect 12650 1460 12660 1480
rect 12620 1450 12660 1460
rect 125 1335 2135 1375
rect 650 690 775 1335
rect 1330 690 1455 1335
rect 2010 695 2135 1335
rect 2840 1440 2870 1450
rect 2840 1420 2845 1440
rect 2865 1420 2870 1440
rect 2840 1390 2870 1420
rect 2840 1370 2845 1390
rect 2865 1370 2870 1390
rect 2840 1340 2870 1370
rect 2840 1320 2845 1340
rect 2865 1320 2870 1340
rect 2840 1290 2870 1320
rect 2840 1270 2845 1290
rect 2865 1270 2870 1290
rect 2840 1240 2870 1270
rect 2840 1220 2845 1240
rect 2865 1220 2870 1240
rect 2840 1210 2870 1220
rect 3380 1440 3410 1450
rect 3380 1420 3385 1440
rect 3405 1420 3410 1440
rect 3380 1390 3410 1420
rect 3380 1370 3385 1390
rect 3405 1370 3410 1390
rect 3380 1340 3410 1370
rect 3380 1320 3385 1340
rect 3405 1320 3410 1340
rect 3380 1290 3410 1320
rect 3380 1270 3385 1290
rect 3405 1270 3410 1290
rect 3380 1240 3410 1270
rect 3380 1220 3385 1240
rect 3405 1220 3410 1240
rect 3380 1210 3410 1220
rect 3920 1440 3950 1450
rect 3920 1420 3925 1440
rect 3945 1420 3950 1440
rect 3920 1390 3950 1420
rect 3920 1370 3925 1390
rect 3945 1370 3950 1390
rect 3920 1340 3950 1370
rect 3920 1320 3925 1340
rect 3945 1320 3950 1340
rect 3920 1290 3950 1320
rect 3920 1270 3925 1290
rect 3945 1270 3950 1290
rect 3920 1240 3950 1270
rect 3920 1220 3925 1240
rect 3945 1220 3950 1240
rect 3920 1210 3950 1220
rect 4060 1440 4090 1450
rect 4060 1420 4065 1440
rect 4085 1420 4090 1440
rect 4060 1390 4090 1420
rect 4060 1370 4065 1390
rect 4085 1370 4090 1390
rect 4060 1340 4090 1370
rect 4060 1320 4065 1340
rect 4085 1320 4090 1340
rect 4060 1290 4090 1320
rect 4060 1270 4065 1290
rect 4085 1270 4090 1290
rect 4060 1240 4090 1270
rect 4060 1220 4065 1240
rect 4085 1220 4090 1240
rect 4060 1210 4090 1220
rect 4600 1440 4630 1450
rect 4600 1420 4605 1440
rect 4625 1420 4630 1440
rect 4600 1390 4630 1420
rect 4600 1370 4605 1390
rect 4625 1370 4630 1390
rect 4600 1340 4630 1370
rect 4600 1320 4605 1340
rect 4625 1320 4630 1340
rect 4600 1290 4630 1320
rect 4600 1270 4605 1290
rect 4625 1270 4630 1290
rect 4600 1240 4630 1270
rect 4600 1220 4605 1240
rect 4625 1220 4630 1240
rect 4600 1210 4630 1220
rect 5140 1440 5170 1450
rect 5140 1420 5145 1440
rect 5165 1420 5170 1440
rect 5140 1390 5170 1420
rect 11810 1400 11850 1440
rect 5140 1370 5145 1390
rect 5165 1370 5170 1390
rect 5140 1340 5170 1370
rect 11315 1350 11355 1390
rect 11880 1350 11920 1390
rect 5140 1320 5145 1340
rect 5165 1320 5170 1340
rect 5140 1290 5170 1320
rect 11315 1320 11355 1330
rect 11315 1300 11325 1320
rect 11345 1300 11355 1320
rect 11315 1290 11355 1300
rect 11425 1320 11465 1330
rect 11425 1300 11435 1320
rect 11455 1300 11465 1320
rect 11425 1290 11465 1300
rect 11535 1320 11575 1330
rect 11535 1300 11545 1320
rect 11565 1300 11575 1320
rect 11535 1290 11575 1300
rect 11645 1320 11685 1330
rect 11645 1300 11655 1320
rect 11675 1300 11685 1320
rect 11645 1290 11685 1300
rect 11755 1320 11795 1330
rect 11755 1300 11765 1320
rect 11785 1300 11795 1320
rect 11755 1290 11795 1300
rect 11815 1320 11845 1330
rect 11815 1300 11820 1320
rect 11840 1300 11845 1320
rect 11815 1290 11845 1300
rect 11865 1320 11905 1330
rect 11865 1300 11875 1320
rect 11895 1300 11905 1320
rect 11865 1290 11905 1300
rect 11975 1320 12015 1330
rect 11975 1300 11985 1320
rect 12005 1300 12015 1320
rect 11975 1290 12015 1300
rect 12085 1320 12125 1330
rect 12085 1300 12095 1320
rect 12115 1300 12125 1320
rect 12085 1290 12125 1300
rect 12195 1320 12235 1330
rect 12195 1300 12205 1320
rect 12225 1300 12235 1320
rect 12195 1290 12235 1300
rect 12305 1320 12345 1330
rect 12305 1300 12315 1320
rect 12335 1300 12345 1320
rect 12305 1290 12345 1300
rect 12415 1320 12455 1330
rect 12415 1300 12425 1320
rect 12445 1300 12455 1320
rect 12415 1290 12455 1300
rect 12525 1320 12565 1330
rect 12525 1300 12535 1320
rect 12555 1300 12565 1320
rect 12525 1290 12565 1300
rect 5140 1270 5145 1290
rect 5165 1270 5170 1290
rect 11325 1270 11345 1290
rect 11435 1270 11455 1290
rect 11545 1270 11565 1290
rect 11655 1270 11675 1290
rect 11765 1270 11785 1290
rect 11875 1270 11895 1290
rect 11985 1270 12005 1290
rect 12095 1270 12115 1290
rect 12205 1270 12225 1290
rect 12315 1270 12335 1290
rect 12425 1270 12445 1290
rect 12535 1270 12555 1290
rect 5140 1240 5170 1270
rect 5140 1220 5145 1240
rect 5165 1220 5170 1240
rect 5140 1210 5170 1220
rect 11170 1260 11240 1270
rect 11170 1240 11175 1260
rect 11195 1240 11215 1260
rect 11235 1240 11240 1260
rect 11170 1210 11240 1240
rect 3385 1190 3405 1210
rect 4605 1190 4625 1210
rect 11170 1190 11175 1210
rect 11195 1190 11215 1210
rect 11235 1190 11240 1210
rect 3375 1180 3415 1190
rect 3375 1160 3385 1180
rect 3405 1160 3415 1180
rect 3375 1150 3415 1160
rect 3990 1155 4020 1185
rect 4595 1180 4635 1190
rect 4595 1160 4605 1180
rect 4625 1160 4635 1180
rect 4595 1150 4635 1160
rect 11170 1160 11240 1190
rect 11170 1140 11175 1160
rect 11195 1140 11215 1160
rect 11235 1140 11240 1160
rect 2945 1120 2985 1130
rect 2945 1100 2955 1120
rect 2975 1100 2985 1120
rect 2945 1090 2985 1100
rect 3025 1120 3065 1130
rect 3025 1100 3035 1120
rect 3055 1100 3065 1120
rect 3025 1090 3065 1100
rect 3105 1120 3145 1130
rect 3105 1100 3115 1120
rect 3135 1100 3145 1120
rect 3105 1090 3145 1100
rect 3185 1120 3225 1130
rect 3185 1100 3195 1120
rect 3215 1100 3225 1120
rect 3185 1090 3225 1100
rect 3265 1120 3305 1130
rect 3265 1100 3275 1120
rect 3295 1100 3305 1120
rect 3265 1090 3305 1100
rect 3345 1120 3385 1130
rect 3345 1100 3355 1120
rect 3375 1100 3385 1120
rect 3345 1090 3385 1100
rect 3425 1120 3465 1130
rect 3425 1100 3435 1120
rect 3455 1100 3465 1120
rect 3425 1090 3465 1100
rect 3505 1120 3545 1130
rect 3505 1100 3515 1120
rect 3535 1100 3545 1120
rect 3505 1090 3545 1100
rect 3585 1120 3625 1130
rect 3585 1100 3595 1120
rect 3615 1100 3625 1120
rect 3585 1090 3625 1100
rect 3665 1120 3705 1130
rect 3665 1100 3675 1120
rect 3695 1100 3705 1120
rect 3665 1090 3705 1100
rect 3745 1120 3785 1130
rect 3745 1100 3755 1120
rect 3775 1100 3785 1120
rect 3745 1090 3785 1100
rect 3825 1120 3865 1130
rect 3825 1100 3835 1120
rect 3855 1100 3865 1120
rect 3825 1090 3865 1100
rect 3905 1120 3945 1130
rect 3905 1100 3915 1120
rect 3935 1100 3945 1120
rect 3905 1090 3945 1100
rect 3985 1120 4025 1130
rect 3985 1100 3995 1120
rect 4015 1100 4025 1120
rect 3985 1090 4025 1100
rect 4065 1120 4105 1130
rect 4065 1100 4075 1120
rect 4095 1100 4105 1120
rect 4065 1090 4105 1100
rect 4145 1120 4185 1130
rect 4145 1100 4155 1120
rect 4175 1100 4185 1120
rect 4145 1090 4185 1100
rect 4225 1120 4265 1130
rect 4225 1100 4235 1120
rect 4255 1100 4265 1120
rect 4225 1090 4265 1100
rect 4305 1120 4345 1130
rect 4305 1100 4315 1120
rect 4335 1100 4345 1120
rect 4305 1090 4345 1100
rect 4385 1120 4425 1130
rect 4385 1100 4395 1120
rect 4415 1100 4425 1120
rect 4385 1090 4425 1100
rect 4465 1120 4505 1130
rect 4465 1100 4475 1120
rect 4495 1100 4505 1120
rect 4465 1090 4505 1100
rect 4545 1120 4585 1130
rect 4545 1100 4555 1120
rect 4575 1100 4585 1120
rect 4545 1090 4585 1100
rect 4625 1120 4665 1130
rect 4625 1100 4635 1120
rect 4655 1100 4665 1120
rect 4625 1090 4665 1100
rect 4705 1120 4745 1130
rect 4705 1100 4715 1120
rect 4735 1100 4745 1120
rect 4705 1090 4745 1100
rect 4785 1120 4825 1130
rect 4785 1100 4795 1120
rect 4815 1100 4825 1120
rect 4785 1090 4825 1100
rect 4865 1120 4905 1130
rect 4865 1100 4875 1120
rect 4895 1100 4905 1120
rect 4865 1090 4905 1100
rect 4945 1120 4985 1130
rect 4945 1100 4955 1120
rect 4975 1100 4985 1120
rect 4945 1090 4985 1100
rect 11170 1110 11240 1140
rect 11170 1090 11175 1110
rect 11195 1090 11215 1110
rect 11235 1090 11240 1110
rect 2955 1070 2975 1090
rect 3995 1070 4015 1090
rect 2950 1060 2980 1070
rect 2950 1045 2955 1060
rect 2935 1040 2955 1045
rect 2975 1040 2980 1060
rect 2625 1010 2655 1040
rect 2910 1035 2980 1040
rect 2910 1015 2915 1035
rect 2935 1015 2980 1035
rect 2910 1010 2980 1015
rect 2935 1005 2955 1010
rect 2950 990 2955 1005
rect 2975 990 2980 1010
rect 2950 980 2980 990
rect 3990 1060 4020 1070
rect 3990 1040 3995 1060
rect 4015 1040 4020 1060
rect 3990 1010 4020 1040
rect 3990 990 3995 1010
rect 4015 990 4020 1010
rect 3990 980 4020 990
rect 5030 1060 5100 1070
rect 5030 1040 5035 1060
rect 5055 1040 5075 1060
rect 5095 1045 5100 1060
rect 11170 1060 11240 1090
rect 5095 1040 5150 1045
rect 5030 1035 5150 1040
rect 5030 1015 5120 1035
rect 5140 1015 5150 1035
rect 11170 1040 11175 1060
rect 11195 1040 11215 1060
rect 11235 1040 11240 1060
rect 11170 1030 11240 1040
rect 11265 1260 11295 1270
rect 11265 1240 11270 1260
rect 11290 1240 11295 1260
rect 11265 1210 11295 1240
rect 11265 1190 11270 1210
rect 11290 1190 11295 1210
rect 11265 1160 11295 1190
rect 11265 1140 11270 1160
rect 11290 1140 11295 1160
rect 11265 1110 11295 1140
rect 11265 1090 11270 1110
rect 11290 1090 11295 1110
rect 11265 1060 11295 1090
rect 11265 1040 11270 1060
rect 11290 1040 11295 1060
rect 11265 1030 11295 1040
rect 11320 1260 11350 1270
rect 11320 1240 11325 1260
rect 11345 1240 11350 1260
rect 11320 1210 11350 1240
rect 11320 1190 11325 1210
rect 11345 1190 11350 1210
rect 11320 1160 11350 1190
rect 11320 1140 11325 1160
rect 11345 1140 11350 1160
rect 11320 1110 11350 1140
rect 11320 1090 11325 1110
rect 11345 1090 11350 1110
rect 11320 1060 11350 1090
rect 11320 1040 11325 1060
rect 11345 1040 11350 1060
rect 11320 1030 11350 1040
rect 11375 1260 11405 1270
rect 11375 1240 11380 1260
rect 11400 1240 11405 1260
rect 11375 1210 11405 1240
rect 11375 1190 11380 1210
rect 11400 1190 11405 1210
rect 11375 1160 11405 1190
rect 11375 1140 11380 1160
rect 11400 1140 11405 1160
rect 11375 1110 11405 1140
rect 11375 1090 11380 1110
rect 11400 1090 11405 1110
rect 11375 1060 11405 1090
rect 11375 1040 11380 1060
rect 11400 1040 11405 1060
rect 11375 1030 11405 1040
rect 11430 1260 11460 1270
rect 11430 1240 11435 1260
rect 11455 1240 11460 1260
rect 11430 1210 11460 1240
rect 11430 1190 11435 1210
rect 11455 1190 11460 1210
rect 11430 1160 11460 1190
rect 11430 1140 11435 1160
rect 11455 1140 11460 1160
rect 11430 1110 11460 1140
rect 11430 1090 11435 1110
rect 11455 1090 11460 1110
rect 11430 1060 11460 1090
rect 11430 1040 11435 1060
rect 11455 1040 11460 1060
rect 11430 1030 11460 1040
rect 11485 1260 11515 1270
rect 11485 1240 11490 1260
rect 11510 1240 11515 1260
rect 11485 1210 11515 1240
rect 11485 1190 11490 1210
rect 11510 1190 11515 1210
rect 11485 1160 11515 1190
rect 11485 1140 11490 1160
rect 11510 1140 11515 1160
rect 11485 1110 11515 1140
rect 11485 1090 11490 1110
rect 11510 1090 11515 1110
rect 11485 1060 11515 1090
rect 11485 1040 11490 1060
rect 11510 1040 11515 1060
rect 11485 1030 11515 1040
rect 11540 1260 11570 1270
rect 11540 1240 11545 1260
rect 11565 1240 11570 1260
rect 11540 1210 11570 1240
rect 11540 1190 11545 1210
rect 11565 1190 11570 1210
rect 11540 1160 11570 1190
rect 11540 1140 11545 1160
rect 11565 1140 11570 1160
rect 11540 1110 11570 1140
rect 11540 1090 11545 1110
rect 11565 1090 11570 1110
rect 11540 1060 11570 1090
rect 11540 1040 11545 1060
rect 11565 1040 11570 1060
rect 11540 1030 11570 1040
rect 11595 1260 11625 1270
rect 11595 1240 11600 1260
rect 11620 1240 11625 1260
rect 11595 1210 11625 1240
rect 11595 1190 11600 1210
rect 11620 1190 11625 1210
rect 11595 1160 11625 1190
rect 11595 1140 11600 1160
rect 11620 1140 11625 1160
rect 11595 1110 11625 1140
rect 11595 1090 11600 1110
rect 11620 1090 11625 1110
rect 11595 1060 11625 1090
rect 11595 1040 11600 1060
rect 11620 1040 11625 1060
rect 11595 1030 11625 1040
rect 11650 1260 11680 1270
rect 11650 1240 11655 1260
rect 11675 1240 11680 1260
rect 11650 1210 11680 1240
rect 11650 1190 11655 1210
rect 11675 1190 11680 1210
rect 11650 1160 11680 1190
rect 11650 1140 11655 1160
rect 11675 1140 11680 1160
rect 11650 1110 11680 1140
rect 11650 1090 11655 1110
rect 11675 1090 11680 1110
rect 11650 1060 11680 1090
rect 11650 1040 11655 1060
rect 11675 1040 11680 1060
rect 11650 1030 11680 1040
rect 11705 1260 11735 1270
rect 11705 1240 11710 1260
rect 11730 1240 11735 1260
rect 11705 1210 11735 1240
rect 11705 1190 11710 1210
rect 11730 1190 11735 1210
rect 11705 1160 11735 1190
rect 11705 1140 11710 1160
rect 11730 1140 11735 1160
rect 11705 1110 11735 1140
rect 11705 1090 11710 1110
rect 11730 1090 11735 1110
rect 11705 1060 11735 1090
rect 11705 1040 11710 1060
rect 11730 1040 11735 1060
rect 11705 1030 11735 1040
rect 11760 1260 11790 1270
rect 11760 1240 11765 1260
rect 11785 1240 11790 1260
rect 11760 1210 11790 1240
rect 11760 1190 11765 1210
rect 11785 1190 11790 1210
rect 11760 1160 11790 1190
rect 11760 1140 11765 1160
rect 11785 1140 11790 1160
rect 11760 1110 11790 1140
rect 11760 1090 11765 1110
rect 11785 1090 11790 1110
rect 11760 1060 11790 1090
rect 11760 1040 11765 1060
rect 11785 1040 11790 1060
rect 11760 1030 11790 1040
rect 11815 1260 11845 1270
rect 11815 1240 11820 1260
rect 11840 1240 11845 1260
rect 11815 1210 11845 1240
rect 11815 1190 11820 1210
rect 11840 1190 11845 1210
rect 11815 1160 11845 1190
rect 11815 1140 11820 1160
rect 11840 1140 11845 1160
rect 11815 1110 11845 1140
rect 11815 1090 11820 1110
rect 11840 1090 11845 1110
rect 11815 1060 11845 1090
rect 11815 1040 11820 1060
rect 11840 1040 11845 1060
rect 11815 1030 11845 1040
rect 11870 1260 11900 1270
rect 11870 1240 11875 1260
rect 11895 1240 11900 1260
rect 11870 1210 11900 1240
rect 11870 1190 11875 1210
rect 11895 1190 11900 1210
rect 11870 1160 11900 1190
rect 11870 1140 11875 1160
rect 11895 1140 11900 1160
rect 11870 1110 11900 1140
rect 11870 1090 11875 1110
rect 11895 1090 11900 1110
rect 11870 1060 11900 1090
rect 11870 1040 11875 1060
rect 11895 1040 11900 1060
rect 11870 1030 11900 1040
rect 11925 1260 11955 1270
rect 11925 1240 11930 1260
rect 11950 1240 11955 1260
rect 11925 1210 11955 1240
rect 11925 1190 11930 1210
rect 11950 1190 11955 1210
rect 11925 1160 11955 1190
rect 11925 1140 11930 1160
rect 11950 1140 11955 1160
rect 11925 1110 11955 1140
rect 11925 1090 11930 1110
rect 11950 1090 11955 1110
rect 11925 1060 11955 1090
rect 11925 1040 11930 1060
rect 11950 1040 11955 1060
rect 11925 1030 11955 1040
rect 11980 1260 12010 1270
rect 11980 1240 11985 1260
rect 12005 1240 12010 1260
rect 11980 1210 12010 1240
rect 11980 1190 11985 1210
rect 12005 1190 12010 1210
rect 11980 1160 12010 1190
rect 11980 1140 11985 1160
rect 12005 1140 12010 1160
rect 11980 1110 12010 1140
rect 11980 1090 11985 1110
rect 12005 1090 12010 1110
rect 11980 1060 12010 1090
rect 11980 1040 11985 1060
rect 12005 1040 12010 1060
rect 11980 1030 12010 1040
rect 12035 1260 12065 1270
rect 12035 1240 12040 1260
rect 12060 1240 12065 1260
rect 12035 1210 12065 1240
rect 12035 1190 12040 1210
rect 12060 1190 12065 1210
rect 12035 1160 12065 1190
rect 12035 1140 12040 1160
rect 12060 1140 12065 1160
rect 12035 1110 12065 1140
rect 12035 1090 12040 1110
rect 12060 1090 12065 1110
rect 12035 1060 12065 1090
rect 12035 1040 12040 1060
rect 12060 1040 12065 1060
rect 12035 1030 12065 1040
rect 12090 1260 12120 1270
rect 12090 1240 12095 1260
rect 12115 1240 12120 1260
rect 12090 1210 12120 1240
rect 12090 1190 12095 1210
rect 12115 1190 12120 1210
rect 12090 1160 12120 1190
rect 12090 1140 12095 1160
rect 12115 1140 12120 1160
rect 12090 1110 12120 1140
rect 12090 1090 12095 1110
rect 12115 1090 12120 1110
rect 12090 1060 12120 1090
rect 12090 1040 12095 1060
rect 12115 1040 12120 1060
rect 12090 1030 12120 1040
rect 12145 1260 12175 1270
rect 12145 1240 12150 1260
rect 12170 1240 12175 1260
rect 12145 1210 12175 1240
rect 12145 1190 12150 1210
rect 12170 1190 12175 1210
rect 12145 1160 12175 1190
rect 12145 1140 12150 1160
rect 12170 1140 12175 1160
rect 12145 1110 12175 1140
rect 12145 1090 12150 1110
rect 12170 1090 12175 1110
rect 12145 1060 12175 1090
rect 12145 1040 12150 1060
rect 12170 1040 12175 1060
rect 12145 1030 12175 1040
rect 12200 1260 12230 1270
rect 12200 1240 12205 1260
rect 12225 1240 12230 1260
rect 12200 1210 12230 1240
rect 12200 1190 12205 1210
rect 12225 1190 12230 1210
rect 12200 1160 12230 1190
rect 12200 1140 12205 1160
rect 12225 1140 12230 1160
rect 12200 1110 12230 1140
rect 12200 1090 12205 1110
rect 12225 1090 12230 1110
rect 12200 1060 12230 1090
rect 12200 1040 12205 1060
rect 12225 1040 12230 1060
rect 12200 1030 12230 1040
rect 12255 1260 12285 1270
rect 12255 1240 12260 1260
rect 12280 1240 12285 1260
rect 12255 1210 12285 1240
rect 12255 1190 12260 1210
rect 12280 1190 12285 1210
rect 12255 1160 12285 1190
rect 12255 1140 12260 1160
rect 12280 1140 12285 1160
rect 12255 1110 12285 1140
rect 12255 1090 12260 1110
rect 12280 1090 12285 1110
rect 12255 1060 12285 1090
rect 12255 1040 12260 1060
rect 12280 1040 12285 1060
rect 12255 1030 12285 1040
rect 12310 1260 12340 1270
rect 12310 1240 12315 1260
rect 12335 1240 12340 1260
rect 12310 1210 12340 1240
rect 12310 1190 12315 1210
rect 12335 1190 12340 1210
rect 12310 1160 12340 1190
rect 12310 1140 12315 1160
rect 12335 1140 12340 1160
rect 12310 1110 12340 1140
rect 12310 1090 12315 1110
rect 12335 1090 12340 1110
rect 12310 1060 12340 1090
rect 12310 1040 12315 1060
rect 12335 1040 12340 1060
rect 12310 1030 12340 1040
rect 12365 1260 12395 1270
rect 12365 1240 12370 1260
rect 12390 1240 12395 1260
rect 12365 1210 12395 1240
rect 12365 1190 12370 1210
rect 12390 1190 12395 1210
rect 12365 1160 12395 1190
rect 12365 1140 12370 1160
rect 12390 1140 12395 1160
rect 12365 1110 12395 1140
rect 12365 1090 12370 1110
rect 12390 1090 12395 1110
rect 12365 1060 12395 1090
rect 12365 1040 12370 1060
rect 12390 1040 12395 1060
rect 12365 1030 12395 1040
rect 12420 1260 12450 1270
rect 12420 1240 12425 1260
rect 12445 1240 12450 1260
rect 12420 1210 12450 1240
rect 12420 1190 12425 1210
rect 12445 1190 12450 1210
rect 12420 1160 12450 1190
rect 12420 1140 12425 1160
rect 12445 1140 12450 1160
rect 12420 1110 12450 1140
rect 12420 1090 12425 1110
rect 12445 1090 12450 1110
rect 12420 1060 12450 1090
rect 12420 1040 12425 1060
rect 12445 1040 12450 1060
rect 12420 1030 12450 1040
rect 12475 1260 12505 1270
rect 12475 1240 12480 1260
rect 12500 1240 12505 1260
rect 12475 1210 12505 1240
rect 12475 1190 12480 1210
rect 12500 1190 12505 1210
rect 12475 1160 12505 1190
rect 12475 1140 12480 1160
rect 12500 1140 12505 1160
rect 12475 1110 12505 1140
rect 12475 1090 12480 1110
rect 12500 1090 12505 1110
rect 12475 1060 12505 1090
rect 12475 1040 12480 1060
rect 12500 1040 12505 1060
rect 12475 1030 12505 1040
rect 12530 1260 12560 1270
rect 12530 1240 12535 1260
rect 12555 1240 12560 1260
rect 12530 1210 12560 1240
rect 12530 1190 12535 1210
rect 12555 1190 12560 1210
rect 12530 1160 12560 1190
rect 12530 1140 12535 1160
rect 12555 1140 12560 1160
rect 12530 1110 12560 1140
rect 12530 1090 12535 1110
rect 12555 1090 12560 1110
rect 12530 1060 12560 1090
rect 12530 1040 12535 1060
rect 12555 1040 12560 1060
rect 12530 1030 12560 1040
rect 12585 1260 12655 1270
rect 12585 1240 12590 1260
rect 12610 1240 12630 1260
rect 12650 1240 12655 1260
rect 12585 1210 12655 1240
rect 12585 1190 12590 1210
rect 12610 1190 12630 1210
rect 12650 1190 12655 1210
rect 12585 1160 12655 1190
rect 12585 1140 12590 1160
rect 12610 1140 12630 1160
rect 12650 1140 12655 1160
rect 12585 1110 12655 1140
rect 12585 1090 12590 1110
rect 12610 1090 12630 1110
rect 12650 1090 12655 1110
rect 12585 1060 12655 1090
rect 12585 1040 12590 1060
rect 12610 1040 12630 1060
rect 12650 1040 12655 1060
rect 12585 1030 12655 1040
rect 5030 1010 5150 1015
rect 11175 1010 11195 1030
rect 11270 1010 11290 1030
rect 11380 1010 11400 1030
rect 11490 1010 11510 1030
rect 11600 1010 11620 1030
rect 11710 1010 11730 1030
rect 11820 1010 11840 1030
rect 11930 1010 11950 1030
rect 12040 1010 12060 1030
rect 12150 1010 12170 1030
rect 12260 1010 12280 1030
rect 12370 1010 12390 1030
rect 12480 1010 12500 1030
rect 12630 1010 12650 1030
rect 5030 990 5035 1010
rect 5055 990 5075 1010
rect 5095 1005 5150 1010
rect 5095 990 5100 1005
rect 5030 980 5100 990
rect 11165 1000 11205 1010
rect 11165 980 11175 1000
rect 11195 980 11205 1000
rect 11165 970 11205 980
rect 11260 1000 11300 1010
rect 11260 980 11270 1000
rect 11290 980 11300 1000
rect 11260 970 11300 980
rect 11370 1000 11410 1010
rect 11370 980 11380 1000
rect 11400 980 11410 1000
rect 11370 970 11410 980
rect 11480 1000 11520 1010
rect 11480 980 11490 1000
rect 11510 980 11520 1000
rect 11480 970 11520 980
rect 11590 1000 11630 1010
rect 11590 980 11600 1000
rect 11620 980 11630 1000
rect 11590 970 11630 980
rect 11700 1000 11740 1010
rect 11700 980 11710 1000
rect 11730 980 11740 1000
rect 11700 970 11740 980
rect 11810 1000 11850 1010
rect 11810 980 11820 1000
rect 11840 980 11850 1000
rect 11810 970 11850 980
rect 11920 1000 11960 1010
rect 11920 980 11930 1000
rect 11950 980 11960 1000
rect 11920 970 11960 980
rect 12030 1000 12070 1010
rect 12030 980 12040 1000
rect 12060 980 12070 1000
rect 12030 970 12070 980
rect 12140 1000 12180 1010
rect 12140 980 12150 1000
rect 12170 980 12180 1000
rect 12140 970 12180 980
rect 12250 1000 12290 1010
rect 12250 980 12260 1000
rect 12280 980 12290 1000
rect 12250 970 12290 980
rect 12360 1000 12400 1010
rect 12360 980 12370 1000
rect 12390 980 12400 1000
rect 12360 970 12400 980
rect 12470 1000 12510 1010
rect 12470 980 12480 1000
rect 12500 980 12510 1000
rect 12470 970 12510 980
rect 12620 1000 12660 1010
rect 12620 980 12630 1000
rect 12650 980 12660 1000
rect 12620 970 12660 980
rect 2995 925 3035 935
rect 2995 905 3005 925
rect 3025 905 3035 925
rect 2995 895 3035 905
rect 3175 925 3215 935
rect 3175 905 3185 925
rect 3205 905 3215 925
rect 3175 895 3215 905
rect 3355 925 3395 935
rect 3355 905 3365 925
rect 3385 905 3395 925
rect 3355 895 3395 905
rect 3535 925 3575 935
rect 3535 905 3545 925
rect 3565 905 3575 925
rect 3535 895 3575 905
rect 3715 925 3755 935
rect 3715 905 3725 925
rect 3745 905 3755 925
rect 3715 895 3755 905
rect 3895 925 3935 935
rect 3895 905 3905 925
rect 3925 905 3935 925
rect 3895 895 3935 905
rect 4075 925 4115 935
rect 4075 905 4085 925
rect 4105 905 4115 925
rect 4075 895 4115 905
rect 4255 925 4295 935
rect 4255 905 4265 925
rect 4285 905 4295 925
rect 4255 895 4295 905
rect 4435 925 4475 935
rect 4435 905 4445 925
rect 4465 905 4475 925
rect 4435 895 4475 905
rect 4615 925 4655 935
rect 4615 905 4625 925
rect 4645 905 4655 925
rect 4615 895 4655 905
rect 4795 925 4835 935
rect 4795 905 4805 925
rect 4825 905 4835 925
rect 4795 895 4835 905
rect 4975 925 5015 935
rect 4975 905 4985 925
rect 5005 905 5015 925
rect 4975 895 5015 905
rect 3005 875 3025 895
rect 3185 875 3205 895
rect 3365 875 3385 895
rect 3545 875 3565 895
rect 3725 875 3745 895
rect 3905 875 3925 895
rect 4085 875 4105 895
rect 4265 875 4285 895
rect 4445 875 4465 895
rect 4625 875 4645 895
rect 4805 875 4825 895
rect 4985 875 5005 895
rect 2960 865 3030 875
rect 2960 845 2965 865
rect 2985 845 3005 865
rect 3025 845 3030 865
rect 2960 815 3030 845
rect 2960 795 2965 815
rect 2985 795 3005 815
rect 3025 795 3030 815
rect 2960 785 3030 795
rect 3090 865 3120 875
rect 3090 845 3095 865
rect 3115 845 3120 865
rect 3090 815 3120 845
rect 3090 795 3095 815
rect 3115 795 3120 815
rect 3090 785 3120 795
rect 3180 865 3210 875
rect 3180 845 3185 865
rect 3205 845 3210 865
rect 3180 815 3210 845
rect 3180 795 3185 815
rect 3205 795 3210 815
rect 3180 785 3210 795
rect 3270 865 3300 875
rect 3270 845 3275 865
rect 3295 845 3300 865
rect 3270 815 3300 845
rect 3270 795 3275 815
rect 3295 795 3300 815
rect 3270 785 3300 795
rect 3360 865 3390 875
rect 3360 845 3365 865
rect 3385 845 3390 865
rect 3360 815 3390 845
rect 3360 795 3365 815
rect 3385 795 3390 815
rect 3360 785 3390 795
rect 3450 865 3480 875
rect 3450 845 3455 865
rect 3475 845 3480 865
rect 3450 815 3480 845
rect 3450 795 3455 815
rect 3475 795 3480 815
rect 3450 785 3480 795
rect 3540 865 3570 875
rect 3540 845 3545 865
rect 3565 845 3570 865
rect 3540 815 3570 845
rect 3540 795 3545 815
rect 3565 795 3570 815
rect 3540 785 3570 795
rect 3630 865 3660 875
rect 3630 845 3635 865
rect 3655 845 3660 865
rect 3630 815 3660 845
rect 3630 795 3635 815
rect 3655 795 3660 815
rect 3630 785 3660 795
rect 3720 865 3750 875
rect 3720 845 3725 865
rect 3745 845 3750 865
rect 3720 815 3750 845
rect 3720 795 3725 815
rect 3745 795 3750 815
rect 3720 785 3750 795
rect 3810 865 3840 875
rect 3810 845 3815 865
rect 3835 845 3840 865
rect 3810 815 3840 845
rect 3810 795 3815 815
rect 3835 795 3840 815
rect 3810 785 3840 795
rect 3900 865 3930 875
rect 3900 845 3905 865
rect 3925 845 3930 865
rect 3900 815 3930 845
rect 3900 795 3905 815
rect 3925 795 3930 815
rect 3900 785 3930 795
rect 3990 865 4020 875
rect 3990 845 3995 865
rect 4015 845 4020 865
rect 3990 815 4020 845
rect 3990 795 3995 815
rect 4015 795 4020 815
rect 3990 785 4020 795
rect 4080 865 4110 875
rect 4080 845 4085 865
rect 4105 845 4110 865
rect 4080 815 4110 845
rect 4080 795 4085 815
rect 4105 795 4110 815
rect 4080 785 4110 795
rect 4170 865 4200 875
rect 4170 845 4175 865
rect 4195 845 4200 865
rect 4170 815 4200 845
rect 4170 795 4175 815
rect 4195 795 4200 815
rect 4170 785 4200 795
rect 4260 865 4290 875
rect 4260 845 4265 865
rect 4285 845 4290 865
rect 4260 815 4290 845
rect 4260 795 4265 815
rect 4285 795 4290 815
rect 4260 785 4290 795
rect 4350 865 4380 875
rect 4350 845 4355 865
rect 4375 845 4380 865
rect 4350 815 4380 845
rect 4350 795 4355 815
rect 4375 795 4380 815
rect 4350 785 4380 795
rect 4440 865 4470 875
rect 4440 845 4445 865
rect 4465 845 4470 865
rect 4440 815 4470 845
rect 4440 795 4445 815
rect 4465 795 4470 815
rect 4440 785 4470 795
rect 4530 865 4560 875
rect 4530 845 4535 865
rect 4555 845 4560 865
rect 4530 815 4560 845
rect 4530 795 4535 815
rect 4555 795 4560 815
rect 4530 785 4560 795
rect 4620 865 4650 875
rect 4620 845 4625 865
rect 4645 845 4650 865
rect 4620 815 4650 845
rect 4620 795 4625 815
rect 4645 795 4650 815
rect 4620 785 4650 795
rect 4710 865 4740 875
rect 4710 845 4715 865
rect 4735 845 4740 865
rect 4710 815 4740 845
rect 4710 795 4715 815
rect 4735 795 4740 815
rect 4710 785 4740 795
rect 4800 865 4830 875
rect 4800 845 4805 865
rect 4825 845 4830 865
rect 4800 815 4830 845
rect 4800 795 4805 815
rect 4825 795 4830 815
rect 4800 785 4830 795
rect 4890 865 4920 875
rect 4890 845 4895 865
rect 4915 845 4920 865
rect 4890 815 4920 845
rect 4890 795 4895 815
rect 4915 795 4920 815
rect 4890 785 4920 795
rect 4980 865 5050 875
rect 4980 845 4985 865
rect 5005 845 5025 865
rect 5045 845 5050 865
rect 4980 815 5050 845
rect 4980 795 4985 815
rect 5005 795 5025 815
rect 5045 795 5050 815
rect 4980 785 5050 795
rect 3095 765 3115 785
rect 3275 765 3295 785
rect 3455 765 3475 785
rect 3635 765 3655 785
rect 3815 765 3835 785
rect 3995 765 4015 785
rect 4175 765 4195 785
rect 4355 765 4375 785
rect 4535 765 4555 785
rect 4715 765 4735 785
rect 4895 765 4915 785
rect 2525 730 2555 760
rect 3095 755 3170 765
rect 3095 745 3140 755
rect 3130 735 3140 745
rect 3160 735 3170 755
rect 3130 725 3170 735
rect 3265 755 3305 765
rect 3265 735 3275 755
rect 3295 735 3305 755
rect 3265 725 3305 735
rect 3445 755 3485 765
rect 3445 735 3455 755
rect 3475 735 3485 755
rect 3445 725 3485 735
rect 3625 755 3665 765
rect 3625 735 3635 755
rect 3655 735 3665 755
rect 3625 725 3665 735
rect 3805 755 3845 765
rect 3805 735 3815 755
rect 3835 735 3845 755
rect 3805 725 3845 735
rect 3985 755 4025 765
rect 3985 735 3995 755
rect 4015 735 4025 755
rect 3985 725 4025 735
rect 4165 755 4205 765
rect 4165 735 4175 755
rect 4195 735 4205 755
rect 4165 725 4205 735
rect 4345 755 4385 765
rect 4345 735 4355 755
rect 4375 735 4385 755
rect 4345 725 4385 735
rect 4525 755 4565 765
rect 4525 735 4535 755
rect 4555 735 4565 755
rect 4525 725 4565 735
rect 4705 755 4745 765
rect 4705 735 4715 755
rect 4735 735 4745 755
rect 4705 725 4745 735
rect 4885 755 4925 765
rect 4885 735 4895 755
rect 4915 735 4925 755
rect 4885 725 4925 735
rect 3450 675 3480 705
rect 3810 675 3840 705
rect 4170 675 4200 705
<< viali >>
rect 56 3175 81 3200
rect 1271 3170 1296 3195
rect 56 3115 81 3140
rect 1271 3110 1296 3135
rect 56 3035 81 3060
rect 56 2975 81 3000
rect 920 2880 950 2910
rect 1000 2880 1030 2910
rect 1080 2880 1110 2910
rect 2340 2930 2365 2955
rect 3090 2955 3110 2975
rect 3145 2955 3165 2975
rect 3275 2955 3295 2975
rect 3455 2955 3475 2975
rect 3635 2955 3655 2975
rect 3815 2955 3835 2975
rect 3995 2955 4015 2975
rect 4175 2955 4195 2975
rect 4355 2955 4375 2975
rect 4535 2955 4555 2975
rect 4715 2955 4735 2975
rect 4845 2955 4865 2975
rect 4895 2955 4915 2975
rect 2340 2870 2365 2895
rect 61 2825 86 2850
rect 734 2825 759 2850
rect 1271 2810 1296 2835
rect 1970 2810 1995 2835
rect 61 2765 86 2790
rect 734 2765 759 2790
rect 3005 2785 3025 2805
rect 3185 2785 3205 2805
rect 3365 2785 3385 2805
rect 3545 2785 3565 2805
rect 3725 2785 3745 2805
rect 3905 2785 3925 2805
rect 4085 2785 4105 2805
rect 4265 2785 4285 2805
rect 4445 2785 4465 2805
rect 4625 2785 4645 2805
rect 4805 2785 4825 2805
rect 4985 2785 5005 2805
rect 3185 2725 3205 2745
rect 3365 2725 3385 2745
rect 3545 2725 3565 2745
rect 3725 2725 3745 2745
rect 3905 2725 3925 2745
rect 4085 2725 4105 2745
rect 4265 2725 4285 2745
rect 4445 2725 4465 2745
rect 4625 2725 4645 2745
rect 4805 2725 4825 2745
rect 3275 2355 3295 2375
rect 3365 2350 3385 2370
rect 3455 2355 3475 2375
rect 3815 2355 3835 2375
rect 3895 2355 3915 2375
rect 3995 2355 4015 2375
rect 4175 2355 4195 2375
rect 4535 2355 4555 2375
rect 4715 2355 4735 2375
rect 3635 2310 3655 2330
rect 4355 2310 4375 2330
rect 3455 2265 3475 2285
rect 4535 2265 4555 2285
rect 2755 2070 2775 2090
rect 2875 2070 2895 2090
rect 2995 2070 3015 2090
rect 3115 2070 3135 2090
rect 3235 2070 3255 2090
rect 3355 2070 3375 2090
rect 3475 2070 3495 2090
rect 3595 2070 3615 2090
rect 3715 2070 3735 2090
rect 3835 2070 3855 2090
rect 3995 2070 4015 2090
rect 4155 2070 4175 2090
rect 4275 2070 4295 2090
rect 4395 2070 4415 2090
rect 4515 2070 4535 2090
rect 4635 2070 4655 2090
rect 4755 2070 4775 2090
rect 4875 2070 4895 2090
rect 4995 2070 5015 2090
rect 5115 2070 5135 2090
rect 5235 2070 5255 2090
rect 2630 2025 2650 2045
rect -35 1695 -15 1715
rect 2815 2025 2835 2045
rect 3175 2025 3195 2045
rect 3535 2025 3555 2045
rect 3895 2025 3915 2045
rect 4095 2025 4115 2045
rect 4455 2025 4475 2045
rect 4815 2025 4835 2045
rect 5175 2025 5195 2045
rect 2575 1855 2595 1875
rect 2630 1855 2650 1875
rect 2685 1855 2705 1875
rect 2845 1855 2865 1875
rect 2935 1855 2955 1875
rect 3055 1855 3075 1875
rect 3175 1855 3195 1875
rect 3295 1855 3315 1875
rect 3415 1855 3435 1875
rect 3535 1855 3555 1875
rect 3655 1855 3675 1875
rect 3775 1855 3795 1875
rect 3865 1855 3885 1875
rect 4125 1855 4145 1875
rect 4215 1855 4235 1875
rect 4335 1855 4355 1875
rect 4455 1855 4475 1875
rect 4575 1855 4595 1875
rect 4695 1855 4715 1875
rect 4815 1855 4835 1875
rect 4935 1855 4955 1875
rect 5055 1855 5075 1875
rect 5145 1855 5165 1875
rect 3055 1795 3075 1815
rect 3415 1795 3435 1815
rect 3775 1795 3795 1815
rect 4215 1795 4235 1815
rect 4575 1795 4595 1815
rect 4935 1795 4955 1815
rect 11095 1785 11115 1805
rect 11200 1800 11220 1820
rect 3235 1735 3255 1755
rect 3295 1735 3315 1755
rect 3535 1735 3555 1755
rect 3775 1735 3795 1755
rect 4215 1735 4235 1755
rect 4455 1735 4475 1755
rect 4695 1735 4715 1755
rect 4755 1735 4775 1755
rect 3175 1690 3195 1710
rect 3415 1690 3435 1710
rect 3655 1690 3675 1710
rect 4335 1690 4355 1710
rect 4575 1690 4595 1710
rect 11315 1785 11335 1805
rect 11420 1800 11440 1820
rect 11243 1740 11260 1760
rect 11535 1785 11555 1805
rect 11650 1800 11670 1820
rect 11463 1740 11480 1760
rect 11610 1740 11627 1760
rect 12135 1785 12155 1805
rect 12240 1800 12260 1820
rect 11825 1740 11845 1760
rect 11876 1740 11893 1760
rect 11955 1740 11975 1760
rect 12355 1785 12375 1805
rect 12460 1800 12480 1820
rect 12283 1740 12300 1760
rect 12575 1785 12595 1805
rect 12690 1800 12710 1820
rect 12503 1740 12520 1760
rect 12650 1740 12667 1760
rect 4815 1690 4835 1710
rect 3995 1630 4015 1650
rect 3175 1570 3195 1590
rect 4815 1570 4835 1590
rect 3235 1520 3255 1540
rect 3355 1520 3375 1540
rect 3475 1520 3495 1540
rect 3595 1520 3615 1540
rect 3715 1520 3735 1540
rect 4275 1520 4295 1540
rect 4395 1520 4415 1540
rect 4515 1520 4535 1540
rect 4635 1520 4655 1540
rect 4755 1520 4775 1540
rect 11112 1520 11129 1540
rect 2845 1460 2865 1480
rect 2935 1475 2955 1495
rect 3055 1475 3075 1495
rect 3175 1475 3195 1495
rect 3295 1475 3315 1495
rect 3535 1475 3555 1495
rect 3655 1475 3675 1495
rect 3775 1475 3795 1495
rect 3925 1460 3945 1480
rect 4065 1460 4085 1480
rect 4215 1475 4235 1495
rect 4335 1475 4355 1495
rect 4455 1475 4475 1495
rect 4695 1475 4715 1495
rect 4815 1475 4835 1495
rect 4935 1475 4955 1495
rect 5055 1475 5075 1495
rect 11315 1520 11335 1540
rect 11535 1520 11555 1540
rect 11830 1520 11850 1540
rect 11880 1520 11900 1540
rect 11928 1520 11945 1540
rect 12152 1520 12169 1540
rect 12355 1520 12375 1540
rect 12575 1520 12595 1540
rect 5145 1460 5165 1480
rect 11155 1460 11175 1480
rect 11260 1460 11280 1480
rect 11370 1460 11390 1480
rect 11480 1460 11500 1480
rect 11590 1460 11610 1480
rect 12195 1460 12215 1480
rect 12300 1460 12320 1480
rect 12410 1460 12430 1480
rect 12520 1460 12540 1480
rect 12630 1460 12650 1480
rect 11325 1300 11345 1320
rect 11435 1300 11455 1320
rect 11545 1300 11565 1320
rect 11655 1300 11675 1320
rect 11765 1300 11785 1320
rect 11820 1300 11840 1320
rect 11875 1300 11895 1320
rect 11985 1300 12005 1320
rect 12095 1300 12115 1320
rect 12205 1300 12225 1320
rect 12315 1300 12335 1320
rect 12425 1300 12445 1320
rect 12535 1300 12555 1320
rect 3385 1160 3405 1180
rect 4605 1160 4625 1180
rect 2955 1100 2975 1120
rect 3035 1100 3055 1120
rect 3115 1100 3135 1120
rect 3195 1100 3215 1120
rect 3275 1100 3295 1120
rect 3355 1100 3375 1120
rect 3435 1100 3455 1120
rect 3515 1100 3535 1120
rect 3595 1100 3615 1120
rect 3675 1100 3695 1120
rect 3755 1100 3775 1120
rect 3835 1100 3855 1120
rect 3915 1100 3935 1120
rect 3995 1100 4015 1120
rect 4075 1100 4095 1120
rect 4155 1100 4175 1120
rect 4235 1100 4255 1120
rect 4315 1100 4335 1120
rect 4395 1100 4415 1120
rect 4475 1100 4495 1120
rect 4555 1100 4575 1120
rect 4635 1100 4655 1120
rect 4715 1100 4735 1120
rect 4795 1100 4815 1120
rect 4875 1100 4895 1120
rect 4955 1100 4975 1120
rect 2915 1015 2935 1035
rect 5120 1015 5140 1035
rect 11175 980 11195 1000
rect 11270 980 11290 1000
rect 11380 980 11400 1000
rect 11490 980 11510 1000
rect 11600 980 11620 1000
rect 11710 980 11730 1000
rect 11820 980 11840 1000
rect 11930 980 11950 1000
rect 12040 980 12060 1000
rect 12150 980 12170 1000
rect 12260 980 12280 1000
rect 12370 980 12390 1000
rect 12480 980 12500 1000
rect 12630 980 12650 1000
rect 3005 905 3025 925
rect 3185 905 3205 925
rect 3365 905 3385 925
rect 3545 905 3565 925
rect 3725 905 3745 925
rect 3905 905 3925 925
rect 4085 905 4105 925
rect 4265 905 4285 925
rect 4445 905 4465 925
rect 4625 905 4645 925
rect 4805 905 4825 925
rect 4985 905 5005 925
rect 3140 735 3160 755
rect 3275 735 3295 755
rect 3455 735 3475 755
rect 3635 735 3655 755
rect 3815 735 3835 755
rect 3995 735 4015 755
rect 4175 735 4195 755
rect 4355 735 4375 755
rect 4535 735 4555 755
rect 4715 735 4735 755
rect 4895 735 4915 755
<< metal1 >>
rect 1261 3525 1301 3530
rect 1261 3495 1266 3525
rect 1296 3495 1301 3525
rect 1261 3490 1301 3495
rect 4440 3495 4480 3500
rect -15 3445 25 3450
rect -15 3415 -10 3445
rect 20 3415 25 3445
rect -15 3410 25 3415
rect 940 3445 980 3450
rect 940 3415 945 3445
rect 975 3415 980 3445
rect 940 3410 980 3415
rect -60 3390 -20 3395
rect -60 3360 -55 3390
rect -25 3360 -20 3390
rect -60 3355 -20 3360
rect -50 2860 -30 3355
rect -60 2855 -20 2860
rect -60 2825 -55 2855
rect -25 2825 -20 2855
rect -60 2820 -20 2825
rect -5 2800 15 3410
rect 1205 3340 1245 3345
rect 1205 3310 1210 3340
rect 1240 3310 1245 3340
rect 1205 3305 1245 3310
rect 1160 3285 1200 3290
rect 1160 3255 1165 3285
rect 1195 3255 1200 3285
rect 1160 3250 1200 3255
rect 46 3170 51 3205
rect 86 3170 91 3205
rect 46 3110 51 3145
rect 86 3110 91 3145
rect 1170 3105 1190 3250
rect 1160 3100 1200 3105
rect 1160 3070 1165 3100
rect 1195 3070 1200 3100
rect 1160 3065 1200 3070
rect 46 3030 51 3065
rect 86 3030 91 3065
rect 46 2970 51 3005
rect 86 2970 91 3005
rect 905 2910 1125 2920
rect 905 2880 920 2910
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1125 2910
rect 905 2870 1125 2880
rect 1215 2855 1235 3305
rect 1271 3200 1291 3490
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect 1635 3445 1685 3455
rect 1635 3415 1645 3445
rect 1675 3415 1685 3445
rect 2470 3450 2510 3455
rect 2470 3420 2475 3450
rect 2505 3420 2510 3450
rect 2470 3415 2510 3420
rect 1635 3405 1685 3415
rect 1261 3165 1266 3200
rect 1301 3165 1306 3200
rect 1271 3140 1291 3165
rect 1261 3105 1266 3140
rect 1301 3105 1306 3140
rect 2330 2925 2335 2960
rect 2370 2925 2375 2960
rect 2425 2955 2465 2960
rect 2425 2925 2430 2955
rect 2460 2925 2465 2955
rect 2425 2920 2465 2925
rect 2330 2900 2375 2905
rect 2330 2865 2335 2900
rect 2370 2865 2375 2900
rect 2330 2860 2375 2865
rect 51 2820 56 2855
rect 91 2820 96 2855
rect 724 2820 729 2855
rect 764 2820 769 2855
rect 1205 2850 1245 2855
rect 1205 2820 1210 2850
rect 1240 2820 1245 2850
rect 2340 2840 2360 2860
rect 1205 2815 1245 2820
rect 1261 2805 1266 2840
rect 1301 2805 1306 2840
rect 1960 2805 1965 2840
rect 2000 2805 2005 2840
rect 2330 2835 2370 2840
rect 2330 2805 2335 2835
rect 2365 2805 2370 2835
rect -15 2795 25 2800
rect -15 2765 -10 2795
rect 20 2765 25 2795
rect -15 2760 25 2765
rect 51 2760 56 2795
rect 91 2760 96 2795
rect 724 2760 729 2795
rect 764 2760 769 2795
rect 1271 2750 1291 2805
rect 2330 2800 2370 2805
rect 1261 2745 1301 2750
rect 1261 2715 1266 2745
rect 1296 2715 1301 2745
rect 1261 2710 1301 2715
rect 2150 2745 2190 2750
rect 2150 2715 2155 2745
rect 2185 2715 2190 2745
rect 2150 2710 2190 2715
rect 275 2200 1985 2550
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1715 -70 1720
rect -45 1720 -5 1725
rect -45 1715 -40 1720
rect -75 1695 -40 1715
rect -75 1690 -70 1695
rect -110 1685 -70 1690
rect -45 1690 -40 1695
rect -10 1690 -5 1720
rect -45 1685 -5 1690
rect 275 1190 625 2200
rect 952 1710 1302 1870
rect 952 1680 1270 1710
rect 1297 1680 1302 1710
rect 952 1520 1302 1680
rect 1330 1190 1455 1345
rect 1635 1190 1985 2200
rect 2160 1190 2180 2710
rect 2340 2205 2360 2800
rect 2435 2250 2455 2920
rect 2425 2245 2465 2250
rect 2425 2215 2430 2245
rect 2460 2215 2465 2245
rect 2425 2210 2465 2215
rect 2330 2200 2370 2205
rect 2330 2170 2335 2200
rect 2365 2170 2370 2200
rect 2330 2165 2370 2170
rect 2340 1600 2360 2165
rect 2380 2150 2420 2155
rect 2380 2120 2385 2150
rect 2415 2120 2420 2150
rect 2380 2115 2420 2120
rect 2390 1670 2410 2115
rect 2435 1765 2455 2210
rect 2480 1825 2500 3415
rect 2690 3390 2730 3395
rect 2690 3360 2695 3390
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 3135 3340 3175 3345
rect 3135 3310 3140 3340
rect 3170 3310 3175 3340
rect 3135 3305 3175 3310
rect 3385 3335 3435 3345
rect 3385 3305 3395 3335
rect 3425 3305 3435 3335
rect 2735 3240 2775 3245
rect 2735 3210 2740 3240
rect 2770 3210 2775 3240
rect 2735 3205 2775 3210
rect 2620 3185 2660 3190
rect 2620 3155 2625 3185
rect 2655 3155 2660 3185
rect 2620 3150 2660 3155
rect 2520 2980 2560 2985
rect 2520 2950 2525 2980
rect 2555 2950 2560 2980
rect 2520 2945 2560 2950
rect 2470 1820 2510 1825
rect 2470 1790 2475 1820
rect 2505 1790 2510 1820
rect 2470 1785 2510 1790
rect 2425 1760 2465 1765
rect 2425 1730 2430 1760
rect 2460 1730 2465 1760
rect 2425 1725 2465 1730
rect 2380 1665 2420 1670
rect 2380 1635 2385 1665
rect 2415 1635 2420 1665
rect 2380 1630 2420 1635
rect 2330 1595 2370 1600
rect 2330 1565 2335 1595
rect 2365 1565 2370 1595
rect 2330 1560 2370 1565
rect 275 840 2180 1190
rect 2530 765 2550 2945
rect 2630 2795 2650 3150
rect 2620 2790 2660 2795
rect 2620 2760 2625 2790
rect 2655 2760 2660 2790
rect 2620 2755 2660 2760
rect 2630 2350 2650 2755
rect 2620 2345 2660 2350
rect 2620 2315 2625 2345
rect 2655 2315 2660 2345
rect 2620 2310 2660 2315
rect 2630 2055 2650 2310
rect 2745 2295 2765 3205
rect 3145 3145 3165 3305
rect 3385 3295 3435 3305
rect 4450 3190 4470 3460
rect 5135 3445 5185 3455
rect 5135 3415 5145 3445
rect 5175 3415 5185 3445
rect 5135 3405 5185 3415
rect 5360 3335 5400 3340
rect 5360 3305 5365 3335
rect 5395 3305 5400 3335
rect 5360 3300 5400 3305
rect 4885 3285 4925 3290
rect 4885 3255 4890 3285
rect 4920 3255 4925 3285
rect 4885 3250 4925 3255
rect 4440 3185 4480 3190
rect 4440 3155 4445 3185
rect 4475 3155 4480 3185
rect 4440 3150 4480 3155
rect 3135 3140 3175 3145
rect 3135 3110 3140 3140
rect 3170 3110 3175 3140
rect 3135 3105 3175 3110
rect 4835 3140 4875 3145
rect 4835 3110 4840 3140
rect 4870 3110 4875 3140
rect 4835 3105 4875 3110
rect 3145 2985 3165 3105
rect 3985 3080 4025 3085
rect 3985 3050 3990 3080
rect 4020 3050 4025 3080
rect 3985 3045 4025 3050
rect 3445 3035 3485 3040
rect 3445 3005 3450 3035
rect 3480 3005 3485 3035
rect 3445 3000 3485 3005
rect 3805 3035 3845 3040
rect 3805 3005 3810 3035
rect 3840 3005 3845 3035
rect 3805 3000 3845 3005
rect 3455 2985 3475 3000
rect 3815 2985 3835 3000
rect 3995 2985 4015 3045
rect 4345 3035 4385 3040
rect 4345 3005 4350 3035
rect 4380 3005 4385 3035
rect 4345 3000 4385 3005
rect 4705 3035 4745 3040
rect 4705 3005 4710 3035
rect 4740 3005 4745 3035
rect 4705 3000 4745 3005
rect 4355 2985 4375 3000
rect 4715 2985 4735 3000
rect 4845 2985 4865 3105
rect 4895 2985 4915 3250
rect 5315 3140 5355 3145
rect 5315 3110 5320 3140
rect 5350 3110 5355 3140
rect 5315 3105 5355 3110
rect 3080 2980 3120 2985
rect 3080 2950 3085 2980
rect 3115 2950 3120 2980
rect 3080 2945 3120 2950
rect 3140 2975 3175 2985
rect 3140 2955 3145 2975
rect 3165 2955 3175 2975
rect 3140 2945 3175 2955
rect 3265 2980 3305 2985
rect 3265 2950 3270 2980
rect 3300 2950 3305 2980
rect 3265 2945 3305 2950
rect 3445 2975 3485 2985
rect 3445 2955 3455 2975
rect 3475 2955 3485 2975
rect 3445 2945 3485 2955
rect 3625 2980 3665 2985
rect 3625 2950 3630 2980
rect 3660 2950 3665 2980
rect 3625 2945 3665 2950
rect 3805 2975 3845 2985
rect 3805 2955 3815 2975
rect 3835 2955 3845 2975
rect 3805 2945 3845 2955
rect 3985 2975 4025 2985
rect 3985 2955 3995 2975
rect 4015 2955 4025 2975
rect 3985 2945 4025 2955
rect 4165 2980 4205 2985
rect 4165 2950 4170 2980
rect 4200 2950 4205 2980
rect 4165 2945 4205 2950
rect 4345 2975 4385 2985
rect 4345 2955 4355 2975
rect 4375 2955 4385 2975
rect 4345 2945 4385 2955
rect 4525 2980 4565 2985
rect 4525 2950 4530 2980
rect 4560 2950 4565 2980
rect 4525 2945 4565 2950
rect 4705 2975 4745 2985
rect 4705 2955 4715 2975
rect 4735 2955 4745 2975
rect 4705 2945 4745 2955
rect 4835 2975 4870 2985
rect 4835 2955 4845 2975
rect 4865 2955 4870 2975
rect 4835 2945 4870 2955
rect 4890 2975 4925 2985
rect 4890 2955 4895 2975
rect 4915 2955 4925 2975
rect 4890 2945 4925 2955
rect 2995 2810 3035 2815
rect 2995 2780 3000 2810
rect 3030 2780 3035 2810
rect 2995 2775 3035 2780
rect 3175 2810 3215 2815
rect 3175 2780 3180 2810
rect 3210 2780 3215 2810
rect 3175 2775 3215 2780
rect 3355 2810 3395 2815
rect 3355 2780 3360 2810
rect 3390 2780 3395 2810
rect 3355 2775 3395 2780
rect 3535 2810 3575 2815
rect 3535 2780 3540 2810
rect 3570 2780 3575 2810
rect 3535 2775 3575 2780
rect 3715 2810 3755 2815
rect 3715 2780 3720 2810
rect 3750 2780 3755 2810
rect 3715 2775 3755 2780
rect 3895 2810 3935 2815
rect 3895 2780 3900 2810
rect 3930 2780 3935 2810
rect 3895 2775 3935 2780
rect 4075 2810 4115 2815
rect 4075 2780 4080 2810
rect 4110 2780 4115 2810
rect 4075 2775 4115 2780
rect 4255 2810 4295 2815
rect 4255 2780 4260 2810
rect 4290 2780 4295 2810
rect 4255 2775 4295 2780
rect 4435 2810 4475 2815
rect 4435 2780 4440 2810
rect 4470 2780 4475 2810
rect 4435 2775 4475 2780
rect 4615 2810 4655 2815
rect 4615 2780 4620 2810
rect 4650 2780 4655 2810
rect 4615 2775 4655 2780
rect 4795 2810 4835 2815
rect 4795 2780 4800 2810
rect 4830 2780 4835 2810
rect 4795 2775 4835 2780
rect 4975 2810 5015 2815
rect 4975 2780 4980 2810
rect 5010 2780 5015 2810
rect 4975 2775 5015 2780
rect 4805 2755 4825 2775
rect 3175 2750 3215 2755
rect 3175 2720 3180 2750
rect 3210 2720 3215 2750
rect 3175 2715 3215 2720
rect 3355 2750 3395 2755
rect 3355 2720 3360 2750
rect 3390 2720 3395 2750
rect 3355 2715 3395 2720
rect 3535 2750 3575 2755
rect 3535 2720 3540 2750
rect 3570 2720 3575 2750
rect 3535 2715 3575 2720
rect 3715 2750 3755 2755
rect 3715 2720 3720 2750
rect 3750 2720 3755 2750
rect 3715 2715 3755 2720
rect 3895 2750 3935 2755
rect 3895 2720 3900 2750
rect 3930 2720 3935 2750
rect 3895 2715 3935 2720
rect 4075 2750 4115 2755
rect 4075 2720 4080 2750
rect 4110 2720 4115 2750
rect 4075 2715 4115 2720
rect 4255 2750 4295 2755
rect 4255 2720 4260 2750
rect 4290 2720 4295 2750
rect 4255 2715 4295 2720
rect 4435 2750 4475 2755
rect 4435 2720 4440 2750
rect 4470 2720 4475 2750
rect 4435 2715 4475 2720
rect 4615 2750 4655 2755
rect 4615 2720 4620 2750
rect 4650 2720 4655 2750
rect 4615 2715 4655 2720
rect 4795 2750 4835 2755
rect 4795 2720 4800 2750
rect 4830 2720 4835 2750
rect 4795 2715 4835 2720
rect 3265 2375 3305 2385
rect 3265 2355 3275 2375
rect 3295 2355 3305 2375
rect 3265 2345 3305 2355
rect 3355 2375 3395 2380
rect 3355 2345 3360 2375
rect 3390 2345 3395 2375
rect 3445 2375 3485 2385
rect 3445 2355 3455 2375
rect 3475 2355 3485 2375
rect 3445 2345 3485 2355
rect 3805 2380 3845 2385
rect 3805 2350 3810 2380
rect 3840 2350 3845 2380
rect 3805 2345 3845 2350
rect 3885 2375 3925 2385
rect 3885 2355 3895 2375
rect 3915 2355 3925 2375
rect 3885 2345 3925 2355
rect 3985 2375 4025 2385
rect 3985 2355 3995 2375
rect 4015 2355 4025 2375
rect 3985 2345 4025 2355
rect 4165 2380 4205 2385
rect 4165 2350 4170 2380
rect 4200 2350 4205 2380
rect 4165 2345 4205 2350
rect 4525 2375 4565 2385
rect 4525 2355 4535 2375
rect 4555 2355 4565 2375
rect 4525 2345 4565 2355
rect 4705 2375 4745 2385
rect 4705 2355 4715 2375
rect 4735 2355 4745 2375
rect 4705 2345 4745 2355
rect 2735 2290 2775 2295
rect 2735 2260 2740 2290
rect 2770 2260 2775 2290
rect 2735 2255 2775 2260
rect 3275 2205 3295 2345
rect 3355 2340 3395 2345
rect 3455 2295 3475 2345
rect 3625 2335 3665 2340
rect 3625 2305 3630 2335
rect 3660 2305 3665 2335
rect 3625 2300 3665 2305
rect 3445 2290 3485 2295
rect 3445 2260 3450 2290
rect 3480 2260 3485 2290
rect 3445 2255 3485 2260
rect 3265 2200 3305 2205
rect 3265 2170 3270 2200
rect 3300 2170 3305 2200
rect 3265 2165 3305 2170
rect 3635 2155 3655 2300
rect 3815 2250 3835 2345
rect 3805 2245 3845 2250
rect 3805 2215 3810 2245
rect 3840 2215 3845 2245
rect 3805 2210 3845 2215
rect 3625 2150 3665 2155
rect 3625 2120 3630 2150
rect 3660 2120 3665 2150
rect 3625 2115 3665 2120
rect 2745 2095 2785 2100
rect 2745 2065 2750 2095
rect 2780 2065 2785 2095
rect 2745 2060 2785 2065
rect 2865 2095 2905 2100
rect 2865 2065 2870 2095
rect 2900 2065 2905 2095
rect 2865 2060 2905 2065
rect 2985 2095 3025 2100
rect 2985 2065 2990 2095
rect 3020 2065 3025 2095
rect 2985 2060 3025 2065
rect 3105 2095 3145 2100
rect 3105 2065 3110 2095
rect 3140 2065 3145 2095
rect 3105 2060 3145 2065
rect 3225 2095 3265 2100
rect 3225 2065 3230 2095
rect 3260 2065 3265 2095
rect 3225 2060 3265 2065
rect 3345 2095 3385 2100
rect 3345 2065 3350 2095
rect 3380 2065 3385 2095
rect 3345 2060 3385 2065
rect 3465 2095 3505 2100
rect 3465 2065 3470 2095
rect 3500 2065 3505 2095
rect 3465 2060 3505 2065
rect 3585 2095 3625 2100
rect 3585 2065 3590 2095
rect 3620 2065 3625 2095
rect 3585 2060 3625 2065
rect 3705 2095 3745 2100
rect 3705 2065 3710 2095
rect 3740 2065 3745 2095
rect 3705 2060 3745 2065
rect 3825 2095 3865 2100
rect 3825 2065 3830 2095
rect 3860 2065 3865 2095
rect 3825 2060 3865 2065
rect 3895 2055 3915 2345
rect 3995 2205 4015 2345
rect 4345 2335 4385 2340
rect 4345 2305 4350 2335
rect 4380 2305 4385 2335
rect 4345 2300 4385 2305
rect 4535 2295 4555 2345
rect 4525 2290 4565 2295
rect 4525 2260 4530 2290
rect 4560 2260 4565 2290
rect 4525 2255 4565 2260
rect 4715 2205 4735 2345
rect 5270 2290 5310 2295
rect 5270 2260 5275 2290
rect 5305 2260 5310 2290
rect 5270 2255 5310 2260
rect 3985 2200 4025 2205
rect 3985 2170 3990 2200
rect 4020 2170 4025 2200
rect 3985 2165 4025 2170
rect 4705 2200 4745 2205
rect 4705 2170 4710 2200
rect 4740 2170 4745 2200
rect 4705 2165 4745 2170
rect 4085 2145 4125 2150
rect 4085 2115 4090 2145
rect 4120 2115 4125 2145
rect 4085 2110 4125 2115
rect 3985 2095 4025 2100
rect 3985 2065 3990 2095
rect 4020 2065 4025 2095
rect 3985 2060 4025 2065
rect 4095 2055 4115 2110
rect 4145 2095 4185 2100
rect 4145 2065 4150 2095
rect 4180 2065 4185 2095
rect 4145 2060 4185 2065
rect 4265 2095 4305 2100
rect 4265 2065 4270 2095
rect 4300 2065 4305 2095
rect 4265 2060 4305 2065
rect 4385 2095 4425 2100
rect 4385 2065 4390 2095
rect 4420 2065 4425 2095
rect 4385 2060 4425 2065
rect 4505 2095 4545 2100
rect 4505 2065 4510 2095
rect 4540 2065 4545 2095
rect 4505 2060 4545 2065
rect 4625 2095 4665 2100
rect 4625 2065 4630 2095
rect 4660 2065 4665 2095
rect 4625 2060 4665 2065
rect 4745 2095 4785 2100
rect 4745 2065 4750 2095
rect 4780 2065 4785 2095
rect 4745 2060 4785 2065
rect 4865 2095 4905 2100
rect 4865 2065 4870 2095
rect 4900 2065 4905 2095
rect 4865 2060 4905 2065
rect 4985 2095 5025 2100
rect 4985 2065 4990 2095
rect 5020 2065 5025 2095
rect 4985 2060 5025 2065
rect 5105 2095 5145 2100
rect 5105 2065 5110 2095
rect 5140 2065 5145 2095
rect 5105 2060 5145 2065
rect 5225 2095 5265 2100
rect 5225 2065 5230 2095
rect 5260 2065 5265 2095
rect 5225 2060 5265 2065
rect 2620 2050 2660 2055
rect 2620 2020 2625 2050
rect 2655 2020 2660 2050
rect 2620 2015 2660 2020
rect 2805 2050 2845 2055
rect 2805 2020 2810 2050
rect 2840 2020 2845 2050
rect 2805 2015 2845 2020
rect 3165 2050 3205 2055
rect 3165 2020 3170 2050
rect 3200 2020 3205 2050
rect 3165 2015 3205 2020
rect 3525 2050 3565 2055
rect 3525 2020 3530 2050
rect 3560 2020 3565 2050
rect 3525 2015 3565 2020
rect 3885 2050 3925 2055
rect 3885 2020 3890 2050
rect 3920 2045 3925 2050
rect 4085 2050 4125 2055
rect 4085 2045 4090 2050
rect 3920 2020 3945 2045
rect 3885 2015 3945 2020
rect 2565 1875 2600 1885
rect 2565 1855 2575 1875
rect 2595 1855 2600 1875
rect 2565 1845 2600 1855
rect 2620 1875 2660 1885
rect 2620 1855 2630 1875
rect 2650 1855 2660 1875
rect 2620 1845 2660 1855
rect 2680 1875 2715 1885
rect 2680 1855 2685 1875
rect 2705 1855 2715 1875
rect 2680 1845 2715 1855
rect 2835 1875 2875 1885
rect 2835 1855 2845 1875
rect 2865 1855 2875 1875
rect 2835 1845 2875 1855
rect 2925 1880 2965 1885
rect 2925 1850 2930 1880
rect 2960 1850 2965 1880
rect 2925 1845 2965 1850
rect 3045 1875 3085 1885
rect 3045 1855 3055 1875
rect 3075 1855 3085 1875
rect 3045 1845 3085 1855
rect 3165 1875 3205 1885
rect 3165 1855 3175 1875
rect 3195 1855 3205 1875
rect 3165 1845 3205 1855
rect 3285 1880 3325 1885
rect 3285 1850 3290 1880
rect 3320 1850 3325 1880
rect 3285 1845 3325 1850
rect 3405 1875 3445 1885
rect 3405 1855 3415 1875
rect 3435 1855 3445 1875
rect 3405 1845 3445 1855
rect 3525 1875 3565 1885
rect 3525 1855 3535 1875
rect 3555 1855 3565 1875
rect 3525 1845 3565 1855
rect 3645 1880 3685 1885
rect 3645 1850 3650 1880
rect 3680 1850 3685 1880
rect 3645 1845 3685 1850
rect 3765 1875 3805 1885
rect 3765 1855 3775 1875
rect 3795 1855 3805 1875
rect 3765 1845 3805 1855
rect 3855 1875 3895 1885
rect 3855 1855 3865 1875
rect 3885 1855 3895 1875
rect 3855 1845 3895 1855
rect 2575 1765 2595 1845
rect 2565 1760 2605 1765
rect 2565 1730 2570 1760
rect 2600 1730 2605 1760
rect 2565 1725 2605 1730
rect 2630 1670 2650 1845
rect 2685 1765 2705 1845
rect 2845 1825 2865 1845
rect 3055 1825 3075 1845
rect 3175 1825 3195 1845
rect 2835 1820 2875 1825
rect 2835 1790 2840 1820
rect 2870 1790 2875 1820
rect 2835 1785 2875 1790
rect 3045 1820 3085 1825
rect 3045 1790 3050 1820
rect 3080 1790 3085 1820
rect 3045 1785 3085 1790
rect 3165 1820 3205 1825
rect 3165 1790 3170 1820
rect 3200 1790 3205 1820
rect 3165 1785 3205 1790
rect 2800 1765 2840 1770
rect 3295 1765 3315 1845
rect 3415 1825 3435 1845
rect 3535 1825 3555 1845
rect 3775 1825 3795 1845
rect 3865 1825 3885 1845
rect 3405 1820 3445 1825
rect 3405 1790 3410 1820
rect 3440 1790 3445 1820
rect 3405 1785 3445 1790
rect 3525 1820 3565 1825
rect 3525 1790 3530 1820
rect 3560 1790 3565 1820
rect 3525 1785 3565 1790
rect 3765 1820 3805 1825
rect 3765 1790 3770 1820
rect 3800 1790 3805 1820
rect 3765 1785 3805 1790
rect 3855 1820 3895 1825
rect 3855 1790 3860 1820
rect 3890 1790 3895 1820
rect 3855 1785 3895 1790
rect 2675 1760 2715 1765
rect 2675 1730 2680 1760
rect 2710 1730 2715 1760
rect 2800 1735 2805 1765
rect 2835 1735 2840 1765
rect 2800 1730 2840 1735
rect 3225 1760 3265 1765
rect 3225 1730 3230 1760
rect 3260 1730 3265 1760
rect 2675 1725 2715 1730
rect 2810 1715 2830 1730
rect 3225 1725 3265 1730
rect 3285 1760 3325 1765
rect 3285 1730 3290 1760
rect 3320 1730 3325 1760
rect 3285 1725 3325 1730
rect 3415 1720 3435 1785
rect 3525 1760 3565 1765
rect 3525 1730 3530 1760
rect 3560 1730 3565 1760
rect 3525 1725 3565 1730
rect 3765 1760 3805 1765
rect 3765 1730 3770 1760
rect 3800 1730 3805 1760
rect 3765 1725 3805 1730
rect 3165 1715 3205 1720
rect 2800 1710 2840 1715
rect 2800 1680 2805 1710
rect 2835 1680 2840 1710
rect 3165 1685 3170 1715
rect 3200 1685 3205 1715
rect 3165 1680 3205 1685
rect 3405 1715 3445 1720
rect 3405 1685 3410 1715
rect 3440 1685 3445 1715
rect 3405 1680 3445 1685
rect 3645 1715 3685 1720
rect 3645 1685 3650 1715
rect 3680 1685 3685 1715
rect 3645 1680 3685 1685
rect 2800 1675 2840 1680
rect 2620 1665 2660 1670
rect 2620 1635 2625 1665
rect 2655 1635 2660 1665
rect 2620 1630 2660 1635
rect 2630 1045 2650 1630
rect 3165 1595 3205 1600
rect 3165 1565 3170 1595
rect 3200 1565 3205 1595
rect 3165 1560 3205 1565
rect 2835 1545 2875 1550
rect 2835 1515 2840 1545
rect 2870 1515 2875 1545
rect 2835 1510 2875 1515
rect 3225 1545 3265 1550
rect 3225 1515 3230 1545
rect 3260 1515 3265 1545
rect 3225 1510 3265 1515
rect 3345 1545 3385 1550
rect 3345 1515 3350 1545
rect 3380 1515 3385 1545
rect 3345 1510 3385 1515
rect 3465 1545 3505 1550
rect 3465 1515 3470 1545
rect 3500 1515 3505 1545
rect 3465 1510 3505 1515
rect 3585 1545 3625 1550
rect 3585 1515 3590 1545
rect 3620 1515 3625 1545
rect 3585 1510 3625 1515
rect 3705 1545 3745 1550
rect 3705 1515 3710 1545
rect 3740 1515 3745 1545
rect 3705 1510 3745 1515
rect 2845 1490 2865 1510
rect 2925 1500 2965 1505
rect 2835 1480 2875 1490
rect 2835 1460 2845 1480
rect 2865 1460 2875 1480
rect 2925 1470 2930 1500
rect 2960 1470 2965 1500
rect 2925 1465 2965 1470
rect 3045 1500 3085 1505
rect 3045 1470 3050 1500
rect 3080 1470 3085 1500
rect 3045 1465 3085 1470
rect 3165 1500 3205 1505
rect 3165 1470 3170 1500
rect 3200 1470 3205 1500
rect 3165 1465 3205 1470
rect 3285 1500 3325 1505
rect 3285 1470 3290 1500
rect 3320 1470 3325 1500
rect 3285 1465 3325 1470
rect 3525 1500 3565 1505
rect 3525 1470 3530 1500
rect 3560 1470 3565 1500
rect 3525 1465 3565 1470
rect 3645 1500 3685 1505
rect 3645 1470 3650 1500
rect 3680 1470 3685 1500
rect 3645 1465 3685 1470
rect 3765 1500 3805 1505
rect 3765 1470 3770 1500
rect 3800 1470 3805 1500
rect 3925 1490 3945 2015
rect 4065 2020 4090 2045
rect 4120 2020 4125 2050
rect 4065 2015 4125 2020
rect 4445 2050 4485 2055
rect 4445 2020 4450 2050
rect 4480 2020 4485 2050
rect 4445 2015 4485 2020
rect 4805 2050 4845 2055
rect 4805 2020 4810 2050
rect 4840 2020 4845 2050
rect 4805 2015 4845 2020
rect 5165 2050 5205 2055
rect 5165 2020 5170 2050
rect 5200 2020 5205 2050
rect 5165 2015 5205 2020
rect 3985 1650 4025 1660
rect 3985 1630 3995 1650
rect 4015 1630 4025 1650
rect 3985 1620 4025 1630
rect 3765 1465 3805 1470
rect 3915 1480 3955 1490
rect 2835 1450 2875 1460
rect 3915 1460 3925 1480
rect 3945 1460 3955 1480
rect 3915 1450 3955 1460
rect 3995 1190 4015 1620
rect 4065 1490 4085 2015
rect 4115 1875 4155 1885
rect 4115 1855 4125 1875
rect 4145 1855 4155 1875
rect 4115 1845 4155 1855
rect 4205 1875 4245 1885
rect 4205 1855 4215 1875
rect 4235 1855 4245 1875
rect 4205 1845 4245 1855
rect 4325 1880 4365 1885
rect 4325 1850 4330 1880
rect 4360 1850 4365 1880
rect 4325 1845 4365 1850
rect 4445 1875 4485 1885
rect 4445 1855 4455 1875
rect 4475 1855 4485 1875
rect 4445 1845 4485 1855
rect 4565 1875 4605 1885
rect 4565 1855 4575 1875
rect 4595 1855 4605 1875
rect 4565 1845 4605 1855
rect 4685 1880 4725 1885
rect 4685 1850 4690 1880
rect 4720 1850 4725 1880
rect 4685 1845 4725 1850
rect 4805 1875 4845 1885
rect 4805 1855 4815 1875
rect 4835 1855 4845 1875
rect 4805 1845 4845 1855
rect 4925 1875 4965 1885
rect 4925 1855 4935 1875
rect 4955 1855 4965 1875
rect 4925 1845 4965 1855
rect 5045 1880 5085 1885
rect 5045 1850 5050 1880
rect 5080 1850 5085 1880
rect 5045 1845 5085 1850
rect 5135 1875 5175 1885
rect 5135 1855 5145 1875
rect 5165 1855 5175 1875
rect 5135 1845 5175 1855
rect 4125 1825 4145 1845
rect 4215 1825 4235 1845
rect 4455 1825 4475 1845
rect 4575 1825 4595 1845
rect 4115 1820 4155 1825
rect 4115 1790 4120 1820
rect 4150 1790 4155 1820
rect 4115 1785 4155 1790
rect 4205 1820 4245 1825
rect 4205 1790 4210 1820
rect 4240 1790 4245 1820
rect 4205 1785 4245 1790
rect 4445 1820 4485 1825
rect 4445 1790 4450 1820
rect 4480 1790 4485 1820
rect 4445 1785 4485 1790
rect 4565 1820 4605 1825
rect 4565 1790 4570 1820
rect 4600 1790 4605 1820
rect 4565 1785 4605 1790
rect 4205 1760 4245 1765
rect 4205 1730 4210 1760
rect 4240 1730 4245 1760
rect 4205 1725 4245 1730
rect 4445 1760 4485 1765
rect 4445 1730 4450 1760
rect 4480 1730 4485 1760
rect 4445 1725 4485 1730
rect 4575 1720 4595 1785
rect 4695 1765 4715 1845
rect 4815 1825 4835 1845
rect 4935 1825 4955 1845
rect 5145 1825 5165 1845
rect 4805 1820 4845 1825
rect 4805 1790 4810 1820
rect 4840 1790 4845 1820
rect 4805 1785 4845 1790
rect 4925 1820 4965 1825
rect 4925 1790 4930 1820
rect 4960 1790 4965 1820
rect 4925 1785 4965 1790
rect 5135 1820 5175 1825
rect 5135 1790 5140 1820
rect 5170 1790 5175 1820
rect 5135 1785 5175 1790
rect 5280 1765 5300 2255
rect 5325 2150 5345 3105
rect 5315 2145 5355 2150
rect 5315 2115 5320 2145
rect 5350 2115 5355 2145
rect 5315 2110 5355 2115
rect 5370 1825 5390 3300
rect 5410 3285 5450 3290
rect 5410 3255 5415 3285
rect 5445 3255 5450 3285
rect 5410 3250 5450 3255
rect 5360 1820 5400 1825
rect 5360 1790 5365 1820
rect 5395 1790 5400 1820
rect 5360 1785 5400 1790
rect 4685 1760 4725 1765
rect 4685 1730 4690 1760
rect 4720 1730 4725 1760
rect 4685 1725 4725 1730
rect 4745 1760 4785 1765
rect 4745 1730 4750 1760
rect 4780 1730 4785 1760
rect 4745 1725 4785 1730
rect 5270 1760 5310 1765
rect 5270 1730 5275 1760
rect 5305 1730 5310 1760
rect 5270 1725 5310 1730
rect 4325 1715 4365 1720
rect 4325 1685 4330 1715
rect 4360 1685 4365 1715
rect 4325 1680 4365 1685
rect 4565 1715 4605 1720
rect 4565 1685 4570 1715
rect 4600 1685 4605 1715
rect 4565 1680 4605 1685
rect 4805 1715 4845 1720
rect 4805 1685 4810 1715
rect 4840 1685 4845 1715
rect 4805 1680 4845 1685
rect 5420 1600 5440 3250
rect 11190 1900 11230 1905
rect 11190 1870 11195 1900
rect 11225 1870 11230 1900
rect 11190 1865 11230 1870
rect 11410 1900 11450 1905
rect 11410 1870 11415 1900
rect 11445 1870 11450 1900
rect 11410 1865 11450 1870
rect 11640 1900 11680 1905
rect 11640 1870 11645 1900
rect 11675 1870 11680 1900
rect 11640 1865 11680 1870
rect 12230 1900 12270 1905
rect 12230 1870 12235 1900
rect 12265 1870 12270 1900
rect 12230 1865 12270 1870
rect 12450 1900 12490 1905
rect 12450 1870 12455 1900
rect 12485 1870 12490 1900
rect 12450 1865 12490 1870
rect 12680 1900 12720 1905
rect 12680 1870 12685 1900
rect 12715 1870 12720 1900
rect 12680 1865 12720 1870
rect 11200 1830 11220 1865
rect 11420 1830 11440 1865
rect 11650 1830 11670 1865
rect 11820 1855 11860 1860
rect 11190 1820 11230 1830
rect 11085 1810 11125 1815
rect 11085 1780 11090 1810
rect 11120 1780 11125 1810
rect 11190 1800 11200 1820
rect 11220 1800 11230 1820
rect 11410 1820 11450 1830
rect 11190 1790 11230 1800
rect 11305 1810 11345 1815
rect 11085 1775 11125 1780
rect 11305 1780 11310 1810
rect 11340 1780 11345 1810
rect 11410 1800 11420 1820
rect 11440 1800 11450 1820
rect 11640 1820 11680 1830
rect 11820 1825 11825 1855
rect 11855 1825 11860 1855
rect 11820 1820 11860 1825
rect 11940 1855 11980 1860
rect 11940 1825 11945 1855
rect 11975 1825 11980 1855
rect 12240 1830 12260 1865
rect 12460 1830 12480 1865
rect 12690 1830 12710 1865
rect 11940 1820 11980 1825
rect 12230 1820 12270 1830
rect 11410 1790 11450 1800
rect 11525 1810 11565 1815
rect 11305 1775 11345 1780
rect 11525 1780 11530 1810
rect 11560 1780 11565 1810
rect 11640 1800 11650 1820
rect 11670 1800 11680 1820
rect 11640 1790 11680 1800
rect 11525 1775 11565 1780
rect 11830 1770 11850 1820
rect 11950 1770 11970 1820
rect 12125 1810 12165 1815
rect 12125 1780 12130 1810
rect 12160 1780 12165 1810
rect 12230 1800 12240 1820
rect 12260 1800 12270 1820
rect 12450 1820 12490 1830
rect 12230 1790 12270 1800
rect 12345 1810 12385 1815
rect 12125 1775 12165 1780
rect 12345 1780 12350 1810
rect 12380 1780 12385 1810
rect 12450 1800 12460 1820
rect 12480 1800 12490 1820
rect 12680 1820 12720 1830
rect 12450 1790 12490 1800
rect 12565 1810 12605 1815
rect 12345 1775 12385 1780
rect 12565 1780 12570 1810
rect 12600 1780 12605 1810
rect 12680 1800 12690 1820
rect 12710 1800 12720 1820
rect 12680 1790 12720 1800
rect 12565 1775 12605 1780
rect 11237 1765 11269 1770
rect 11237 1735 11240 1765
rect 11266 1735 11269 1765
rect 11237 1730 11269 1735
rect 11457 1765 11489 1770
rect 11457 1735 11460 1765
rect 11486 1735 11489 1765
rect 11457 1730 11489 1735
rect 11601 1765 11633 1770
rect 11601 1735 11604 1765
rect 11630 1735 11633 1765
rect 11601 1730 11633 1735
rect 11820 1760 11850 1770
rect 11820 1740 11825 1760
rect 11845 1740 11850 1760
rect 11820 1730 11850 1740
rect 11867 1765 11899 1770
rect 11867 1735 11870 1765
rect 11896 1735 11899 1765
rect 11867 1730 11899 1735
rect 11950 1760 11980 1770
rect 11950 1740 11955 1760
rect 11975 1740 11980 1760
rect 11950 1730 11980 1740
rect 12277 1765 12309 1770
rect 12277 1735 12280 1765
rect 12306 1735 12309 1765
rect 12277 1730 12309 1735
rect 12497 1765 12529 1770
rect 12497 1735 12500 1765
rect 12526 1735 12529 1765
rect 12497 1730 12529 1735
rect 12641 1765 12673 1770
rect 12641 1735 12644 1765
rect 12670 1735 12673 1765
rect 12641 1730 12673 1735
rect 4805 1595 4845 1600
rect 4805 1565 4810 1595
rect 4840 1565 4845 1595
rect 4805 1560 4845 1565
rect 5410 1595 5450 1600
rect 5410 1565 5415 1595
rect 5445 1565 5450 1595
rect 5410 1560 5450 1565
rect 4265 1545 4305 1550
rect 4265 1515 4270 1545
rect 4300 1515 4305 1545
rect 4265 1510 4305 1515
rect 4385 1545 4425 1550
rect 4385 1515 4390 1545
rect 4420 1515 4425 1545
rect 4385 1510 4425 1515
rect 4505 1545 4545 1550
rect 4505 1515 4510 1545
rect 4540 1515 4545 1545
rect 4505 1510 4545 1515
rect 4625 1545 4665 1550
rect 4625 1515 4630 1545
rect 4660 1515 4665 1545
rect 4625 1510 4665 1515
rect 4745 1545 4785 1550
rect 4745 1515 4750 1545
rect 4780 1515 4785 1545
rect 4745 1510 4785 1515
rect 5135 1545 5175 1550
rect 5135 1515 5140 1545
rect 5170 1515 5175 1545
rect 5135 1510 5175 1515
rect 11106 1545 11138 1550
rect 11106 1515 11109 1545
rect 11135 1515 11138 1545
rect 11106 1510 11138 1515
rect 11305 1545 11345 1550
rect 11305 1515 11310 1545
rect 11340 1515 11345 1545
rect 11305 1510 11345 1515
rect 11525 1545 11565 1550
rect 11525 1515 11530 1545
rect 11560 1515 11565 1545
rect 11525 1510 11565 1515
rect 11825 1540 11855 1550
rect 11825 1520 11830 1540
rect 11850 1520 11855 1540
rect 11825 1510 11855 1520
rect 11875 1540 11905 1550
rect 11875 1520 11880 1540
rect 11900 1520 11905 1540
rect 11875 1510 11905 1520
rect 11922 1545 11954 1550
rect 11922 1515 11925 1545
rect 11951 1515 11954 1545
rect 11922 1510 11954 1515
rect 12146 1545 12178 1550
rect 12146 1515 12149 1545
rect 12175 1515 12178 1545
rect 12146 1510 12178 1515
rect 12345 1545 12385 1550
rect 12345 1515 12350 1545
rect 12380 1515 12385 1545
rect 12345 1510 12385 1515
rect 12565 1545 12605 1550
rect 12565 1515 12570 1545
rect 12600 1515 12605 1545
rect 12565 1510 12605 1515
rect 4205 1500 4245 1505
rect 4055 1480 4095 1490
rect 4055 1460 4065 1480
rect 4085 1460 4095 1480
rect 4205 1470 4210 1500
rect 4240 1470 4245 1500
rect 4205 1465 4245 1470
rect 4325 1500 4365 1505
rect 4325 1470 4330 1500
rect 4360 1470 4365 1500
rect 4325 1465 4365 1470
rect 4445 1500 4485 1505
rect 4445 1470 4450 1500
rect 4480 1470 4485 1500
rect 4445 1465 4485 1470
rect 4685 1500 4725 1505
rect 4685 1470 4690 1500
rect 4720 1470 4725 1500
rect 4685 1465 4725 1470
rect 4805 1500 4845 1505
rect 4805 1470 4810 1500
rect 4840 1470 4845 1500
rect 4805 1465 4845 1470
rect 4925 1500 4965 1505
rect 4925 1470 4930 1500
rect 4960 1470 4965 1500
rect 4925 1465 4965 1470
rect 5045 1500 5085 1505
rect 5045 1470 5050 1500
rect 5080 1470 5085 1500
rect 5145 1490 5165 1510
rect 5045 1465 5085 1470
rect 5135 1480 5175 1490
rect 4055 1450 4095 1460
rect 5135 1460 5145 1480
rect 5165 1460 5175 1480
rect 5135 1450 5175 1460
rect 11145 1485 11185 1490
rect 11145 1455 11150 1485
rect 11180 1455 11185 1485
rect 11145 1450 11185 1455
rect 11250 1485 11290 1490
rect 11250 1455 11255 1485
rect 11285 1455 11290 1485
rect 11250 1450 11290 1455
rect 11360 1485 11400 1490
rect 11360 1455 11365 1485
rect 11395 1455 11400 1485
rect 11360 1450 11400 1455
rect 11470 1485 11510 1490
rect 11470 1455 11475 1485
rect 11505 1455 11510 1485
rect 11470 1450 11510 1455
rect 11580 1485 11620 1490
rect 11580 1455 11585 1485
rect 11615 1455 11620 1485
rect 11580 1450 11620 1455
rect 11830 1440 11850 1510
rect 11810 1435 11850 1440
rect 11810 1405 11815 1435
rect 11845 1405 11850 1435
rect 11810 1400 11850 1405
rect 11315 1385 11355 1390
rect 11315 1355 11320 1385
rect 11350 1355 11355 1385
rect 11315 1350 11355 1355
rect 11325 1330 11345 1350
rect 11820 1330 11840 1400
rect 11880 1390 11900 1510
rect 12185 1485 12225 1490
rect 12185 1455 12190 1485
rect 12220 1455 12225 1485
rect 12185 1450 12225 1455
rect 12290 1485 12330 1490
rect 12290 1455 12295 1485
rect 12325 1455 12330 1485
rect 12290 1450 12330 1455
rect 12400 1485 12440 1490
rect 12400 1455 12405 1485
rect 12435 1455 12440 1485
rect 12400 1450 12440 1455
rect 12510 1485 12550 1490
rect 12510 1455 12515 1485
rect 12545 1455 12550 1485
rect 12510 1450 12550 1455
rect 12620 1485 12660 1490
rect 12620 1455 12625 1485
rect 12655 1455 12660 1485
rect 12620 1450 12660 1455
rect 11880 1385 11920 1390
rect 11880 1355 11885 1385
rect 11915 1355 11920 1385
rect 11880 1350 11920 1355
rect 11315 1320 11355 1330
rect 11315 1300 11325 1320
rect 11345 1300 11355 1320
rect 11315 1290 11355 1300
rect 11425 1325 11465 1330
rect 11425 1295 11430 1325
rect 11460 1295 11465 1325
rect 11425 1290 11465 1295
rect 11535 1325 11575 1330
rect 11535 1295 11540 1325
rect 11570 1295 11575 1325
rect 11535 1290 11575 1295
rect 11645 1325 11685 1330
rect 11645 1295 11650 1325
rect 11680 1295 11685 1325
rect 11645 1290 11685 1295
rect 11755 1325 11795 1330
rect 11755 1295 11760 1325
rect 11790 1295 11795 1325
rect 11755 1290 11795 1295
rect 11815 1320 11845 1330
rect 11815 1300 11820 1320
rect 11840 1300 11845 1320
rect 11815 1290 11845 1300
rect 11865 1325 11905 1330
rect 11865 1295 11870 1325
rect 11900 1295 11905 1325
rect 11865 1290 11905 1295
rect 11975 1325 12015 1330
rect 11975 1295 11980 1325
rect 12010 1295 12015 1325
rect 11975 1290 12015 1295
rect 12085 1325 12125 1330
rect 12085 1295 12090 1325
rect 12120 1295 12125 1325
rect 12085 1290 12125 1295
rect 12195 1325 12235 1330
rect 12195 1295 12200 1325
rect 12230 1295 12235 1325
rect 12195 1290 12235 1295
rect 12305 1325 12345 1330
rect 12305 1295 12310 1325
rect 12340 1295 12345 1325
rect 12305 1290 12345 1295
rect 12415 1325 12455 1330
rect 12415 1295 12420 1325
rect 12450 1295 12455 1325
rect 12415 1290 12455 1295
rect 12525 1325 12565 1330
rect 12525 1295 12530 1325
rect 12560 1295 12565 1325
rect 12525 1290 12565 1295
rect 3375 1185 3415 1190
rect 3375 1155 3380 1185
rect 3410 1155 3415 1185
rect 3375 1150 3415 1155
rect 3985 1185 4025 1190
rect 3985 1155 3990 1185
rect 4020 1155 4025 1185
rect 3985 1150 4025 1155
rect 4595 1185 4635 1190
rect 4595 1155 4600 1185
rect 4630 1155 4635 1185
rect 4595 1150 4635 1155
rect 2945 1125 2985 1130
rect 2945 1095 2950 1125
rect 2980 1095 2985 1125
rect 2945 1090 2985 1095
rect 3025 1125 3065 1130
rect 3025 1095 3030 1125
rect 3060 1095 3065 1125
rect 3025 1090 3065 1095
rect 3105 1125 3145 1130
rect 3105 1095 3110 1125
rect 3140 1095 3145 1125
rect 3105 1090 3145 1095
rect 3185 1125 3225 1130
rect 3185 1095 3190 1125
rect 3220 1095 3225 1125
rect 3185 1090 3225 1095
rect 3265 1125 3305 1130
rect 3265 1095 3270 1125
rect 3300 1095 3305 1125
rect 3265 1090 3305 1095
rect 3345 1125 3385 1130
rect 3345 1095 3350 1125
rect 3380 1095 3385 1125
rect 3345 1090 3385 1095
rect 3425 1125 3465 1130
rect 3425 1095 3430 1125
rect 3460 1095 3465 1125
rect 3425 1090 3465 1095
rect 3505 1125 3545 1130
rect 3505 1095 3510 1125
rect 3540 1095 3545 1125
rect 3505 1090 3545 1095
rect 3585 1125 3625 1130
rect 3585 1095 3590 1125
rect 3620 1095 3625 1125
rect 3585 1090 3625 1095
rect 3665 1125 3705 1130
rect 3665 1095 3670 1125
rect 3700 1095 3705 1125
rect 3665 1090 3705 1095
rect 3745 1125 3785 1130
rect 3745 1095 3750 1125
rect 3780 1095 3785 1125
rect 3745 1090 3785 1095
rect 3825 1125 3865 1130
rect 3825 1095 3830 1125
rect 3860 1095 3865 1125
rect 3825 1090 3865 1095
rect 3905 1125 3945 1130
rect 3905 1095 3910 1125
rect 3940 1095 3945 1125
rect 3905 1090 3945 1095
rect 3985 1125 4025 1130
rect 3985 1095 3990 1125
rect 4020 1095 4025 1125
rect 3985 1090 4025 1095
rect 4065 1125 4105 1130
rect 4065 1095 4070 1125
rect 4100 1095 4105 1125
rect 4065 1090 4105 1095
rect 4145 1125 4185 1130
rect 4145 1095 4150 1125
rect 4180 1095 4185 1125
rect 4145 1090 4185 1095
rect 4225 1125 4265 1130
rect 4225 1095 4230 1125
rect 4260 1095 4265 1125
rect 4225 1090 4265 1095
rect 4305 1125 4345 1130
rect 4305 1095 4310 1125
rect 4340 1095 4345 1125
rect 4305 1090 4345 1095
rect 4385 1125 4425 1130
rect 4385 1095 4390 1125
rect 4420 1095 4425 1125
rect 4385 1090 4425 1095
rect 4465 1125 4505 1130
rect 4465 1095 4470 1125
rect 4500 1095 4505 1125
rect 4465 1090 4505 1095
rect 4545 1125 4585 1130
rect 4545 1095 4550 1125
rect 4580 1095 4585 1125
rect 4545 1090 4585 1095
rect 4625 1125 4665 1130
rect 4625 1095 4630 1125
rect 4660 1095 4665 1125
rect 4625 1090 4665 1095
rect 4705 1125 4745 1130
rect 4705 1095 4710 1125
rect 4740 1095 4745 1125
rect 4705 1090 4745 1095
rect 4785 1125 4825 1130
rect 4785 1095 4790 1125
rect 4820 1095 4825 1125
rect 4785 1090 4825 1095
rect 4865 1125 4905 1130
rect 4865 1095 4870 1125
rect 4900 1095 4905 1125
rect 4865 1090 4905 1095
rect 4945 1125 4985 1130
rect 4945 1095 4950 1125
rect 4980 1095 4985 1125
rect 4945 1090 4985 1095
rect 2620 1040 2660 1045
rect 2620 1010 2625 1040
rect 2655 1010 2660 1040
rect 2620 1005 2660 1010
rect 2905 1040 2945 1045
rect 2905 1010 2910 1040
rect 2940 1010 2945 1040
rect 2905 1005 2945 1010
rect 5110 1040 5150 1045
rect 5110 1010 5115 1040
rect 5145 1010 5150 1040
rect 5110 1005 5150 1010
rect 11165 1005 11205 1010
rect 11165 975 11170 1005
rect 11200 975 11205 1005
rect 11165 970 11205 975
rect 11260 1005 11300 1010
rect 11260 975 11265 1005
rect 11295 975 11300 1005
rect 11260 970 11300 975
rect 11370 1005 11410 1010
rect 11370 975 11375 1005
rect 11405 975 11410 1005
rect 11370 970 11410 975
rect 11480 1005 11520 1010
rect 11480 975 11485 1005
rect 11515 975 11520 1005
rect 11480 970 11520 975
rect 11590 1005 11630 1010
rect 11590 975 11595 1005
rect 11625 975 11630 1005
rect 11590 970 11630 975
rect 11700 1005 11740 1010
rect 11700 975 11705 1005
rect 11735 975 11740 1005
rect 11700 970 11740 975
rect 11810 1005 11850 1010
rect 11810 975 11815 1005
rect 11845 975 11850 1005
rect 11810 970 11850 975
rect 11920 1005 11960 1010
rect 11920 975 11925 1005
rect 11955 975 11960 1005
rect 11920 970 11960 975
rect 12030 1005 12070 1010
rect 12030 975 12035 1005
rect 12065 975 12070 1005
rect 12030 970 12070 975
rect 12140 1005 12180 1010
rect 12140 975 12145 1005
rect 12175 975 12180 1005
rect 12140 970 12180 975
rect 12250 1005 12290 1010
rect 12250 975 12255 1005
rect 12285 975 12290 1005
rect 12250 970 12290 975
rect 12360 1005 12400 1010
rect 12360 975 12365 1005
rect 12395 975 12400 1005
rect 12360 970 12400 975
rect 12470 1005 12510 1010
rect 12470 975 12475 1005
rect 12505 975 12510 1005
rect 12470 970 12510 975
rect 12620 1005 12660 1010
rect 12620 975 12625 1005
rect 12655 975 12660 1005
rect 12620 970 12660 975
rect 2995 930 3035 935
rect 2995 900 3000 930
rect 3030 900 3035 930
rect 2995 895 3035 900
rect 3175 930 3215 935
rect 3175 900 3180 930
rect 3210 900 3215 930
rect 3175 895 3215 900
rect 3355 930 3395 935
rect 3355 900 3360 930
rect 3390 900 3395 930
rect 3355 895 3395 900
rect 3535 930 3575 935
rect 3535 900 3540 930
rect 3570 900 3575 930
rect 3535 895 3575 900
rect 3715 930 3755 935
rect 3715 900 3720 930
rect 3750 900 3755 930
rect 3715 895 3755 900
rect 3895 930 3935 935
rect 3895 900 3900 930
rect 3930 900 3935 930
rect 3895 895 3935 900
rect 4075 930 4115 935
rect 4075 900 4080 930
rect 4110 900 4115 930
rect 4075 895 4115 900
rect 4255 930 4295 935
rect 4255 900 4260 930
rect 4290 900 4295 930
rect 4255 895 4295 900
rect 4435 930 4475 935
rect 4435 900 4440 930
rect 4470 900 4475 930
rect 4435 895 4475 900
rect 4615 930 4655 935
rect 4615 900 4620 930
rect 4650 900 4655 930
rect 4615 895 4655 900
rect 4795 930 4835 935
rect 4795 900 4800 930
rect 4830 900 4835 930
rect 4795 895 4835 900
rect 4975 930 5015 935
rect 4975 900 4980 930
rect 5010 900 5015 930
rect 4975 895 5015 900
rect 2520 760 2560 765
rect 2520 730 2525 760
rect 2555 730 2560 760
rect 2520 725 2560 730
rect 3130 760 3170 765
rect 3130 730 3135 760
rect 3165 730 3170 760
rect 3130 725 3170 730
rect 3265 755 3305 765
rect 3265 735 3275 755
rect 3295 735 3305 755
rect 3265 725 3305 735
rect 3445 755 3485 765
rect 3445 735 3455 755
rect 3475 735 3485 755
rect 3445 725 3485 735
rect 3625 760 3665 765
rect 3625 730 3630 760
rect 3660 730 3665 760
rect 3625 725 3665 730
rect 3805 755 3845 765
rect 3805 735 3815 755
rect 3835 735 3845 755
rect 3805 725 3845 735
rect 3985 760 4025 765
rect 3985 730 3990 760
rect 4020 730 4025 760
rect 3985 725 4025 730
rect 4165 755 4205 765
rect 4165 735 4175 755
rect 4195 735 4205 755
rect 4165 725 4205 735
rect 4345 760 4385 765
rect 4345 730 4350 760
rect 4380 730 4385 760
rect 4345 725 4385 730
rect 4525 760 4565 765
rect 4525 730 4530 760
rect 4560 730 4565 760
rect 4525 725 4565 730
rect 4705 760 4745 765
rect 4705 730 4710 760
rect 4740 730 4745 760
rect 4705 725 4745 730
rect 4885 760 4925 765
rect 4885 730 4890 760
rect 4920 730 4925 760
rect 4885 725 4925 730
rect 3275 295 3295 725
rect 3455 710 3475 725
rect 3815 710 3835 725
rect 3445 705 3485 710
rect 3445 675 3450 705
rect 3480 675 3485 705
rect 3445 670 3485 675
rect 3805 705 3845 710
rect 3805 675 3810 705
rect 3840 675 3845 705
rect 3805 670 3845 675
rect 3815 295 3835 670
rect 3995 295 4015 725
rect 4175 710 4195 725
rect 4165 705 4205 710
rect 4165 675 4170 705
rect 4200 675 4205 705
rect 4165 670 4205 675
rect 4715 295 4735 725
<< via1 >>
rect 1266 3495 1296 3525
rect -10 3415 20 3445
rect 945 3415 975 3445
rect -55 3360 -25 3390
rect -55 2825 -25 2855
rect 1210 3310 1240 3340
rect 1165 3255 1195 3285
rect 51 3200 86 3205
rect 51 3175 56 3200
rect 56 3175 81 3200
rect 81 3175 86 3200
rect 51 3170 86 3175
rect 51 3140 86 3145
rect 51 3115 56 3140
rect 56 3115 81 3140
rect 81 3115 86 3140
rect 51 3110 86 3115
rect 1165 3070 1195 3100
rect 51 3060 86 3065
rect 51 3035 56 3060
rect 56 3035 81 3060
rect 81 3035 86 3060
rect 51 3030 86 3035
rect 51 3000 86 3005
rect 51 2975 56 3000
rect 56 2975 81 3000
rect 81 2975 86 3000
rect 51 2970 86 2975
rect 920 2880 950 2910
rect 1000 2880 1030 2910
rect 1080 2880 1110 2910
rect 4445 3465 4475 3495
rect 1645 3415 1675 3445
rect 2475 3420 2505 3450
rect 1266 3195 1301 3200
rect 1266 3170 1271 3195
rect 1271 3170 1296 3195
rect 1296 3170 1301 3195
rect 1266 3165 1301 3170
rect 1266 3135 1301 3140
rect 1266 3110 1271 3135
rect 1271 3110 1296 3135
rect 1296 3110 1301 3135
rect 1266 3105 1301 3110
rect 2335 2955 2370 2960
rect 2335 2930 2340 2955
rect 2340 2930 2365 2955
rect 2365 2930 2370 2955
rect 2335 2925 2370 2930
rect 2430 2925 2460 2955
rect 2335 2895 2370 2900
rect 2335 2870 2340 2895
rect 2340 2870 2365 2895
rect 2365 2870 2370 2895
rect 2335 2865 2370 2870
rect 56 2850 91 2855
rect 56 2825 61 2850
rect 61 2825 86 2850
rect 86 2825 91 2850
rect 56 2820 91 2825
rect 729 2850 764 2855
rect 729 2825 734 2850
rect 734 2825 759 2850
rect 759 2825 764 2850
rect 729 2820 764 2825
rect 1210 2820 1240 2850
rect 1266 2835 1301 2840
rect 1266 2810 1271 2835
rect 1271 2810 1296 2835
rect 1296 2810 1301 2835
rect 1266 2805 1301 2810
rect 1965 2835 2000 2840
rect 1965 2810 1970 2835
rect 1970 2810 1995 2835
rect 1995 2810 2000 2835
rect 1965 2805 2000 2810
rect 2335 2805 2365 2835
rect -10 2765 20 2795
rect 56 2790 91 2795
rect 56 2765 61 2790
rect 61 2765 86 2790
rect 86 2765 91 2790
rect 56 2760 91 2765
rect 729 2790 764 2795
rect 729 2765 734 2790
rect 734 2765 759 2790
rect 759 2765 764 2790
rect 729 2760 764 2765
rect 1266 2715 1296 2745
rect 2155 2715 2185 2745
rect -105 1690 -75 1720
rect -40 1715 -10 1720
rect -40 1695 -35 1715
rect -35 1695 -15 1715
rect -15 1695 -10 1715
rect -40 1690 -10 1695
rect 1270 1680 1297 1710
rect 2430 2215 2460 2245
rect 2335 2170 2365 2200
rect 2385 2120 2415 2150
rect 2695 3360 2725 3390
rect 3140 3310 3170 3340
rect 3395 3305 3425 3335
rect 2740 3210 2770 3240
rect 2625 3155 2655 3185
rect 2525 2950 2555 2980
rect 2475 1790 2505 1820
rect 2430 1730 2460 1760
rect 2385 1635 2415 1665
rect 2335 1565 2365 1595
rect 2625 2760 2655 2790
rect 2625 2315 2655 2345
rect 5145 3415 5175 3445
rect 5365 3305 5395 3335
rect 4890 3255 4920 3285
rect 4445 3155 4475 3185
rect 3140 3110 3170 3140
rect 4840 3110 4870 3140
rect 3990 3050 4020 3080
rect 3450 3005 3480 3035
rect 3810 3005 3840 3035
rect 4350 3005 4380 3035
rect 4710 3005 4740 3035
rect 5320 3110 5350 3140
rect 3085 2975 3115 2980
rect 3085 2955 3090 2975
rect 3090 2955 3110 2975
rect 3110 2955 3115 2975
rect 3085 2950 3115 2955
rect 3270 2975 3300 2980
rect 3270 2955 3275 2975
rect 3275 2955 3295 2975
rect 3295 2955 3300 2975
rect 3270 2950 3300 2955
rect 3630 2975 3660 2980
rect 3630 2955 3635 2975
rect 3635 2955 3655 2975
rect 3655 2955 3660 2975
rect 3630 2950 3660 2955
rect 4170 2975 4200 2980
rect 4170 2955 4175 2975
rect 4175 2955 4195 2975
rect 4195 2955 4200 2975
rect 4170 2950 4200 2955
rect 4530 2975 4560 2980
rect 4530 2955 4535 2975
rect 4535 2955 4555 2975
rect 4555 2955 4560 2975
rect 4530 2950 4560 2955
rect 3000 2805 3030 2810
rect 3000 2785 3005 2805
rect 3005 2785 3025 2805
rect 3025 2785 3030 2805
rect 3000 2780 3030 2785
rect 3180 2805 3210 2810
rect 3180 2785 3185 2805
rect 3185 2785 3205 2805
rect 3205 2785 3210 2805
rect 3180 2780 3210 2785
rect 3360 2805 3390 2810
rect 3360 2785 3365 2805
rect 3365 2785 3385 2805
rect 3385 2785 3390 2805
rect 3360 2780 3390 2785
rect 3540 2805 3570 2810
rect 3540 2785 3545 2805
rect 3545 2785 3565 2805
rect 3565 2785 3570 2805
rect 3540 2780 3570 2785
rect 3720 2805 3750 2810
rect 3720 2785 3725 2805
rect 3725 2785 3745 2805
rect 3745 2785 3750 2805
rect 3720 2780 3750 2785
rect 3900 2805 3930 2810
rect 3900 2785 3905 2805
rect 3905 2785 3925 2805
rect 3925 2785 3930 2805
rect 3900 2780 3930 2785
rect 4080 2805 4110 2810
rect 4080 2785 4085 2805
rect 4085 2785 4105 2805
rect 4105 2785 4110 2805
rect 4080 2780 4110 2785
rect 4260 2805 4290 2810
rect 4260 2785 4265 2805
rect 4265 2785 4285 2805
rect 4285 2785 4290 2805
rect 4260 2780 4290 2785
rect 4440 2805 4470 2810
rect 4440 2785 4445 2805
rect 4445 2785 4465 2805
rect 4465 2785 4470 2805
rect 4440 2780 4470 2785
rect 4620 2805 4650 2810
rect 4620 2785 4625 2805
rect 4625 2785 4645 2805
rect 4645 2785 4650 2805
rect 4620 2780 4650 2785
rect 4800 2805 4830 2810
rect 4800 2785 4805 2805
rect 4805 2785 4825 2805
rect 4825 2785 4830 2805
rect 4800 2780 4830 2785
rect 4980 2805 5010 2810
rect 4980 2785 4985 2805
rect 4985 2785 5005 2805
rect 5005 2785 5010 2805
rect 4980 2780 5010 2785
rect 3180 2745 3210 2750
rect 3180 2725 3185 2745
rect 3185 2725 3205 2745
rect 3205 2725 3210 2745
rect 3180 2720 3210 2725
rect 3360 2745 3390 2750
rect 3360 2725 3365 2745
rect 3365 2725 3385 2745
rect 3385 2725 3390 2745
rect 3360 2720 3390 2725
rect 3540 2745 3570 2750
rect 3540 2725 3545 2745
rect 3545 2725 3565 2745
rect 3565 2725 3570 2745
rect 3540 2720 3570 2725
rect 3720 2745 3750 2750
rect 3720 2725 3725 2745
rect 3725 2725 3745 2745
rect 3745 2725 3750 2745
rect 3720 2720 3750 2725
rect 3900 2745 3930 2750
rect 3900 2725 3905 2745
rect 3905 2725 3925 2745
rect 3925 2725 3930 2745
rect 3900 2720 3930 2725
rect 4080 2745 4110 2750
rect 4080 2725 4085 2745
rect 4085 2725 4105 2745
rect 4105 2725 4110 2745
rect 4080 2720 4110 2725
rect 4260 2745 4290 2750
rect 4260 2725 4265 2745
rect 4265 2725 4285 2745
rect 4285 2725 4290 2745
rect 4260 2720 4290 2725
rect 4440 2745 4470 2750
rect 4440 2725 4445 2745
rect 4445 2725 4465 2745
rect 4465 2725 4470 2745
rect 4440 2720 4470 2725
rect 4620 2745 4650 2750
rect 4620 2725 4625 2745
rect 4625 2725 4645 2745
rect 4645 2725 4650 2745
rect 4620 2720 4650 2725
rect 4800 2745 4830 2750
rect 4800 2725 4805 2745
rect 4805 2725 4825 2745
rect 4825 2725 4830 2745
rect 4800 2720 4830 2725
rect 3360 2370 3390 2375
rect 3360 2350 3365 2370
rect 3365 2350 3385 2370
rect 3385 2350 3390 2370
rect 3360 2345 3390 2350
rect 3810 2375 3840 2380
rect 3810 2355 3815 2375
rect 3815 2355 3835 2375
rect 3835 2355 3840 2375
rect 3810 2350 3840 2355
rect 4170 2375 4200 2380
rect 4170 2355 4175 2375
rect 4175 2355 4195 2375
rect 4195 2355 4200 2375
rect 4170 2350 4200 2355
rect 2740 2260 2770 2290
rect 3630 2330 3660 2335
rect 3630 2310 3635 2330
rect 3635 2310 3655 2330
rect 3655 2310 3660 2330
rect 3630 2305 3660 2310
rect 3450 2285 3480 2290
rect 3450 2265 3455 2285
rect 3455 2265 3475 2285
rect 3475 2265 3480 2285
rect 3450 2260 3480 2265
rect 3270 2170 3300 2200
rect 3810 2215 3840 2245
rect 3630 2120 3660 2150
rect 2750 2090 2780 2095
rect 2750 2070 2755 2090
rect 2755 2070 2775 2090
rect 2775 2070 2780 2090
rect 2750 2065 2780 2070
rect 2870 2090 2900 2095
rect 2870 2070 2875 2090
rect 2875 2070 2895 2090
rect 2895 2070 2900 2090
rect 2870 2065 2900 2070
rect 2990 2090 3020 2095
rect 2990 2070 2995 2090
rect 2995 2070 3015 2090
rect 3015 2070 3020 2090
rect 2990 2065 3020 2070
rect 3110 2090 3140 2095
rect 3110 2070 3115 2090
rect 3115 2070 3135 2090
rect 3135 2070 3140 2090
rect 3110 2065 3140 2070
rect 3230 2090 3260 2095
rect 3230 2070 3235 2090
rect 3235 2070 3255 2090
rect 3255 2070 3260 2090
rect 3230 2065 3260 2070
rect 3350 2090 3380 2095
rect 3350 2070 3355 2090
rect 3355 2070 3375 2090
rect 3375 2070 3380 2090
rect 3350 2065 3380 2070
rect 3470 2090 3500 2095
rect 3470 2070 3475 2090
rect 3475 2070 3495 2090
rect 3495 2070 3500 2090
rect 3470 2065 3500 2070
rect 3590 2090 3620 2095
rect 3590 2070 3595 2090
rect 3595 2070 3615 2090
rect 3615 2070 3620 2090
rect 3590 2065 3620 2070
rect 3710 2090 3740 2095
rect 3710 2070 3715 2090
rect 3715 2070 3735 2090
rect 3735 2070 3740 2090
rect 3710 2065 3740 2070
rect 3830 2090 3860 2095
rect 3830 2070 3835 2090
rect 3835 2070 3855 2090
rect 3855 2070 3860 2090
rect 3830 2065 3860 2070
rect 4350 2330 4380 2335
rect 4350 2310 4355 2330
rect 4355 2310 4375 2330
rect 4375 2310 4380 2330
rect 4350 2305 4380 2310
rect 4530 2285 4560 2290
rect 4530 2265 4535 2285
rect 4535 2265 4555 2285
rect 4555 2265 4560 2285
rect 4530 2260 4560 2265
rect 5275 2260 5305 2290
rect 3990 2170 4020 2200
rect 4710 2170 4740 2200
rect 4090 2115 4120 2145
rect 3990 2090 4020 2095
rect 3990 2070 3995 2090
rect 3995 2070 4015 2090
rect 4015 2070 4020 2090
rect 3990 2065 4020 2070
rect 4150 2090 4180 2095
rect 4150 2070 4155 2090
rect 4155 2070 4175 2090
rect 4175 2070 4180 2090
rect 4150 2065 4180 2070
rect 4270 2090 4300 2095
rect 4270 2070 4275 2090
rect 4275 2070 4295 2090
rect 4295 2070 4300 2090
rect 4270 2065 4300 2070
rect 4390 2090 4420 2095
rect 4390 2070 4395 2090
rect 4395 2070 4415 2090
rect 4415 2070 4420 2090
rect 4390 2065 4420 2070
rect 4510 2090 4540 2095
rect 4510 2070 4515 2090
rect 4515 2070 4535 2090
rect 4535 2070 4540 2090
rect 4510 2065 4540 2070
rect 4630 2090 4660 2095
rect 4630 2070 4635 2090
rect 4635 2070 4655 2090
rect 4655 2070 4660 2090
rect 4630 2065 4660 2070
rect 4750 2090 4780 2095
rect 4750 2070 4755 2090
rect 4755 2070 4775 2090
rect 4775 2070 4780 2090
rect 4750 2065 4780 2070
rect 4870 2090 4900 2095
rect 4870 2070 4875 2090
rect 4875 2070 4895 2090
rect 4895 2070 4900 2090
rect 4870 2065 4900 2070
rect 4990 2090 5020 2095
rect 4990 2070 4995 2090
rect 4995 2070 5015 2090
rect 5015 2070 5020 2090
rect 4990 2065 5020 2070
rect 5110 2090 5140 2095
rect 5110 2070 5115 2090
rect 5115 2070 5135 2090
rect 5135 2070 5140 2090
rect 5110 2065 5140 2070
rect 5230 2090 5260 2095
rect 5230 2070 5235 2090
rect 5235 2070 5255 2090
rect 5255 2070 5260 2090
rect 5230 2065 5260 2070
rect 2625 2045 2655 2050
rect 2625 2025 2630 2045
rect 2630 2025 2650 2045
rect 2650 2025 2655 2045
rect 2625 2020 2655 2025
rect 2810 2045 2840 2050
rect 2810 2025 2815 2045
rect 2815 2025 2835 2045
rect 2835 2025 2840 2045
rect 2810 2020 2840 2025
rect 3170 2045 3200 2050
rect 3170 2025 3175 2045
rect 3175 2025 3195 2045
rect 3195 2025 3200 2045
rect 3170 2020 3200 2025
rect 3530 2045 3560 2050
rect 3530 2025 3535 2045
rect 3535 2025 3555 2045
rect 3555 2025 3560 2045
rect 3530 2020 3560 2025
rect 3890 2045 3920 2050
rect 4090 2045 4120 2050
rect 3890 2025 3895 2045
rect 3895 2025 3915 2045
rect 3915 2025 3920 2045
rect 3890 2020 3920 2025
rect 2930 1875 2960 1880
rect 2930 1855 2935 1875
rect 2935 1855 2955 1875
rect 2955 1855 2960 1875
rect 2930 1850 2960 1855
rect 3290 1875 3320 1880
rect 3290 1855 3295 1875
rect 3295 1855 3315 1875
rect 3315 1855 3320 1875
rect 3290 1850 3320 1855
rect 3650 1875 3680 1880
rect 3650 1855 3655 1875
rect 3655 1855 3675 1875
rect 3675 1855 3680 1875
rect 3650 1850 3680 1855
rect 2570 1730 2600 1760
rect 2840 1790 2870 1820
rect 3050 1815 3080 1820
rect 3050 1795 3055 1815
rect 3055 1795 3075 1815
rect 3075 1795 3080 1815
rect 3050 1790 3080 1795
rect 3170 1790 3200 1820
rect 3410 1815 3440 1820
rect 3410 1795 3415 1815
rect 3415 1795 3435 1815
rect 3435 1795 3440 1815
rect 3410 1790 3440 1795
rect 3530 1790 3560 1820
rect 3770 1815 3800 1820
rect 3770 1795 3775 1815
rect 3775 1795 3795 1815
rect 3795 1795 3800 1815
rect 3770 1790 3800 1795
rect 3860 1790 3890 1820
rect 2680 1730 2710 1760
rect 2805 1735 2835 1765
rect 3230 1755 3260 1760
rect 3230 1735 3235 1755
rect 3235 1735 3255 1755
rect 3255 1735 3260 1755
rect 3230 1730 3260 1735
rect 3290 1755 3320 1760
rect 3290 1735 3295 1755
rect 3295 1735 3315 1755
rect 3315 1735 3320 1755
rect 3290 1730 3320 1735
rect 3530 1755 3560 1760
rect 3530 1735 3535 1755
rect 3535 1735 3555 1755
rect 3555 1735 3560 1755
rect 3530 1730 3560 1735
rect 3770 1755 3800 1760
rect 3770 1735 3775 1755
rect 3775 1735 3795 1755
rect 3795 1735 3800 1755
rect 3770 1730 3800 1735
rect 2805 1680 2835 1710
rect 3170 1710 3200 1715
rect 3170 1690 3175 1710
rect 3175 1690 3195 1710
rect 3195 1690 3200 1710
rect 3170 1685 3200 1690
rect 3410 1710 3440 1715
rect 3410 1690 3415 1710
rect 3415 1690 3435 1710
rect 3435 1690 3440 1710
rect 3410 1685 3440 1690
rect 3650 1710 3680 1715
rect 3650 1690 3655 1710
rect 3655 1690 3675 1710
rect 3675 1690 3680 1710
rect 3650 1685 3680 1690
rect 2625 1635 2655 1665
rect 3170 1590 3200 1595
rect 3170 1570 3175 1590
rect 3175 1570 3195 1590
rect 3195 1570 3200 1590
rect 3170 1565 3200 1570
rect 2840 1515 2870 1545
rect 3230 1540 3260 1545
rect 3230 1520 3235 1540
rect 3235 1520 3255 1540
rect 3255 1520 3260 1540
rect 3230 1515 3260 1520
rect 3350 1540 3380 1545
rect 3350 1520 3355 1540
rect 3355 1520 3375 1540
rect 3375 1520 3380 1540
rect 3350 1515 3380 1520
rect 3470 1540 3500 1545
rect 3470 1520 3475 1540
rect 3475 1520 3495 1540
rect 3495 1520 3500 1540
rect 3470 1515 3500 1520
rect 3590 1540 3620 1545
rect 3590 1520 3595 1540
rect 3595 1520 3615 1540
rect 3615 1520 3620 1540
rect 3590 1515 3620 1520
rect 3710 1540 3740 1545
rect 3710 1520 3715 1540
rect 3715 1520 3735 1540
rect 3735 1520 3740 1540
rect 3710 1515 3740 1520
rect 2930 1495 2960 1500
rect 2930 1475 2935 1495
rect 2935 1475 2955 1495
rect 2955 1475 2960 1495
rect 2930 1470 2960 1475
rect 3050 1495 3080 1500
rect 3050 1475 3055 1495
rect 3055 1475 3075 1495
rect 3075 1475 3080 1495
rect 3050 1470 3080 1475
rect 3170 1495 3200 1500
rect 3170 1475 3175 1495
rect 3175 1475 3195 1495
rect 3195 1475 3200 1495
rect 3170 1470 3200 1475
rect 3290 1495 3320 1500
rect 3290 1475 3295 1495
rect 3295 1475 3315 1495
rect 3315 1475 3320 1495
rect 3290 1470 3320 1475
rect 3530 1495 3560 1500
rect 3530 1475 3535 1495
rect 3535 1475 3555 1495
rect 3555 1475 3560 1495
rect 3530 1470 3560 1475
rect 3650 1495 3680 1500
rect 3650 1475 3655 1495
rect 3655 1475 3675 1495
rect 3675 1475 3680 1495
rect 3650 1470 3680 1475
rect 3770 1495 3800 1500
rect 3770 1475 3775 1495
rect 3775 1475 3795 1495
rect 3795 1475 3800 1495
rect 3770 1470 3800 1475
rect 4090 2025 4095 2045
rect 4095 2025 4115 2045
rect 4115 2025 4120 2045
rect 4090 2020 4120 2025
rect 4450 2045 4480 2050
rect 4450 2025 4455 2045
rect 4455 2025 4475 2045
rect 4475 2025 4480 2045
rect 4450 2020 4480 2025
rect 4810 2045 4840 2050
rect 4810 2025 4815 2045
rect 4815 2025 4835 2045
rect 4835 2025 4840 2045
rect 4810 2020 4840 2025
rect 5170 2045 5200 2050
rect 5170 2025 5175 2045
rect 5175 2025 5195 2045
rect 5195 2025 5200 2045
rect 5170 2020 5200 2025
rect 4330 1875 4360 1880
rect 4330 1855 4335 1875
rect 4335 1855 4355 1875
rect 4355 1855 4360 1875
rect 4330 1850 4360 1855
rect 4690 1875 4720 1880
rect 4690 1855 4695 1875
rect 4695 1855 4715 1875
rect 4715 1855 4720 1875
rect 4690 1850 4720 1855
rect 5050 1875 5080 1880
rect 5050 1855 5055 1875
rect 5055 1855 5075 1875
rect 5075 1855 5080 1875
rect 5050 1850 5080 1855
rect 4120 1790 4150 1820
rect 4210 1815 4240 1820
rect 4210 1795 4215 1815
rect 4215 1795 4235 1815
rect 4235 1795 4240 1815
rect 4210 1790 4240 1795
rect 4450 1790 4480 1820
rect 4570 1815 4600 1820
rect 4570 1795 4575 1815
rect 4575 1795 4595 1815
rect 4595 1795 4600 1815
rect 4570 1790 4600 1795
rect 4210 1755 4240 1760
rect 4210 1735 4215 1755
rect 4215 1735 4235 1755
rect 4235 1735 4240 1755
rect 4210 1730 4240 1735
rect 4450 1755 4480 1760
rect 4450 1735 4455 1755
rect 4455 1735 4475 1755
rect 4475 1735 4480 1755
rect 4450 1730 4480 1735
rect 4810 1790 4840 1820
rect 4930 1815 4960 1820
rect 4930 1795 4935 1815
rect 4935 1795 4955 1815
rect 4955 1795 4960 1815
rect 4930 1790 4960 1795
rect 5140 1790 5170 1820
rect 5320 2115 5350 2145
rect 5415 3255 5445 3285
rect 5365 1790 5395 1820
rect 4690 1755 4720 1760
rect 4690 1735 4695 1755
rect 4695 1735 4715 1755
rect 4715 1735 4720 1755
rect 4690 1730 4720 1735
rect 4750 1755 4780 1760
rect 4750 1735 4755 1755
rect 4755 1735 4775 1755
rect 4775 1735 4780 1755
rect 4750 1730 4780 1735
rect 5275 1730 5305 1760
rect 4330 1710 4360 1715
rect 4330 1690 4335 1710
rect 4335 1690 4355 1710
rect 4355 1690 4360 1710
rect 4330 1685 4360 1690
rect 4570 1710 4600 1715
rect 4570 1690 4575 1710
rect 4575 1690 4595 1710
rect 4595 1690 4600 1710
rect 4570 1685 4600 1690
rect 4810 1710 4840 1715
rect 4810 1690 4815 1710
rect 4815 1690 4835 1710
rect 4835 1690 4840 1710
rect 4810 1685 4840 1690
rect 11195 1870 11225 1900
rect 11415 1870 11445 1900
rect 11645 1870 11675 1900
rect 12235 1870 12265 1900
rect 12455 1870 12485 1900
rect 12685 1870 12715 1900
rect 11090 1805 11120 1810
rect 11090 1785 11095 1805
rect 11095 1785 11115 1805
rect 11115 1785 11120 1805
rect 11090 1780 11120 1785
rect 11310 1805 11340 1810
rect 11310 1785 11315 1805
rect 11315 1785 11335 1805
rect 11335 1785 11340 1805
rect 11310 1780 11340 1785
rect 11825 1825 11855 1855
rect 11945 1825 11975 1855
rect 11530 1805 11560 1810
rect 11530 1785 11535 1805
rect 11535 1785 11555 1805
rect 11555 1785 11560 1805
rect 11530 1780 11560 1785
rect 12130 1805 12160 1810
rect 12130 1785 12135 1805
rect 12135 1785 12155 1805
rect 12155 1785 12160 1805
rect 12130 1780 12160 1785
rect 12350 1805 12380 1810
rect 12350 1785 12355 1805
rect 12355 1785 12375 1805
rect 12375 1785 12380 1805
rect 12350 1780 12380 1785
rect 12570 1805 12600 1810
rect 12570 1785 12575 1805
rect 12575 1785 12595 1805
rect 12595 1785 12600 1805
rect 12570 1780 12600 1785
rect 11240 1760 11266 1765
rect 11240 1740 11243 1760
rect 11243 1740 11260 1760
rect 11260 1740 11266 1760
rect 11240 1735 11266 1740
rect 11460 1760 11486 1765
rect 11460 1740 11463 1760
rect 11463 1740 11480 1760
rect 11480 1740 11486 1760
rect 11460 1735 11486 1740
rect 11604 1760 11630 1765
rect 11604 1740 11610 1760
rect 11610 1740 11627 1760
rect 11627 1740 11630 1760
rect 11604 1735 11630 1740
rect 11870 1760 11896 1765
rect 11870 1740 11876 1760
rect 11876 1740 11893 1760
rect 11893 1740 11896 1760
rect 11870 1735 11896 1740
rect 12280 1760 12306 1765
rect 12280 1740 12283 1760
rect 12283 1740 12300 1760
rect 12300 1740 12306 1760
rect 12280 1735 12306 1740
rect 12500 1760 12526 1765
rect 12500 1740 12503 1760
rect 12503 1740 12520 1760
rect 12520 1740 12526 1760
rect 12500 1735 12526 1740
rect 12644 1760 12670 1765
rect 12644 1740 12650 1760
rect 12650 1740 12667 1760
rect 12667 1740 12670 1760
rect 12644 1735 12670 1740
rect 4810 1590 4840 1595
rect 4810 1570 4815 1590
rect 4815 1570 4835 1590
rect 4835 1570 4840 1590
rect 4810 1565 4840 1570
rect 5415 1565 5445 1595
rect 4270 1540 4300 1545
rect 4270 1520 4275 1540
rect 4275 1520 4295 1540
rect 4295 1520 4300 1540
rect 4270 1515 4300 1520
rect 4390 1540 4420 1545
rect 4390 1520 4395 1540
rect 4395 1520 4415 1540
rect 4415 1520 4420 1540
rect 4390 1515 4420 1520
rect 4510 1540 4540 1545
rect 4510 1520 4515 1540
rect 4515 1520 4535 1540
rect 4535 1520 4540 1540
rect 4510 1515 4540 1520
rect 4630 1540 4660 1545
rect 4630 1520 4635 1540
rect 4635 1520 4655 1540
rect 4655 1520 4660 1540
rect 4630 1515 4660 1520
rect 4750 1540 4780 1545
rect 4750 1520 4755 1540
rect 4755 1520 4775 1540
rect 4775 1520 4780 1540
rect 4750 1515 4780 1520
rect 5140 1515 5170 1545
rect 11109 1540 11135 1545
rect 11109 1520 11112 1540
rect 11112 1520 11129 1540
rect 11129 1520 11135 1540
rect 11109 1515 11135 1520
rect 11310 1540 11340 1545
rect 11310 1520 11315 1540
rect 11315 1520 11335 1540
rect 11335 1520 11340 1540
rect 11310 1515 11340 1520
rect 11530 1540 11560 1545
rect 11530 1520 11535 1540
rect 11535 1520 11555 1540
rect 11555 1520 11560 1540
rect 11530 1515 11560 1520
rect 11925 1540 11951 1545
rect 11925 1520 11928 1540
rect 11928 1520 11945 1540
rect 11945 1520 11951 1540
rect 11925 1515 11951 1520
rect 12149 1540 12175 1545
rect 12149 1520 12152 1540
rect 12152 1520 12169 1540
rect 12169 1520 12175 1540
rect 12149 1515 12175 1520
rect 12350 1540 12380 1545
rect 12350 1520 12355 1540
rect 12355 1520 12375 1540
rect 12375 1520 12380 1540
rect 12350 1515 12380 1520
rect 12570 1540 12600 1545
rect 12570 1520 12575 1540
rect 12575 1520 12595 1540
rect 12595 1520 12600 1540
rect 12570 1515 12600 1520
rect 4210 1495 4240 1500
rect 4210 1475 4215 1495
rect 4215 1475 4235 1495
rect 4235 1475 4240 1495
rect 4210 1470 4240 1475
rect 4330 1495 4360 1500
rect 4330 1475 4335 1495
rect 4335 1475 4355 1495
rect 4355 1475 4360 1495
rect 4330 1470 4360 1475
rect 4450 1495 4480 1500
rect 4450 1475 4455 1495
rect 4455 1475 4475 1495
rect 4475 1475 4480 1495
rect 4450 1470 4480 1475
rect 4690 1495 4720 1500
rect 4690 1475 4695 1495
rect 4695 1475 4715 1495
rect 4715 1475 4720 1495
rect 4690 1470 4720 1475
rect 4810 1495 4840 1500
rect 4810 1475 4815 1495
rect 4815 1475 4835 1495
rect 4835 1475 4840 1495
rect 4810 1470 4840 1475
rect 4930 1495 4960 1500
rect 4930 1475 4935 1495
rect 4935 1475 4955 1495
rect 4955 1475 4960 1495
rect 4930 1470 4960 1475
rect 5050 1495 5080 1500
rect 5050 1475 5055 1495
rect 5055 1475 5075 1495
rect 5075 1475 5080 1495
rect 5050 1470 5080 1475
rect 11150 1480 11180 1485
rect 11150 1460 11155 1480
rect 11155 1460 11175 1480
rect 11175 1460 11180 1480
rect 11150 1455 11180 1460
rect 11255 1480 11285 1485
rect 11255 1460 11260 1480
rect 11260 1460 11280 1480
rect 11280 1460 11285 1480
rect 11255 1455 11285 1460
rect 11365 1480 11395 1485
rect 11365 1460 11370 1480
rect 11370 1460 11390 1480
rect 11390 1460 11395 1480
rect 11365 1455 11395 1460
rect 11475 1480 11505 1485
rect 11475 1460 11480 1480
rect 11480 1460 11500 1480
rect 11500 1460 11505 1480
rect 11475 1455 11505 1460
rect 11585 1480 11615 1485
rect 11585 1460 11590 1480
rect 11590 1460 11610 1480
rect 11610 1460 11615 1480
rect 11585 1455 11615 1460
rect 11815 1405 11845 1435
rect 11320 1355 11350 1385
rect 12190 1480 12220 1485
rect 12190 1460 12195 1480
rect 12195 1460 12215 1480
rect 12215 1460 12220 1480
rect 12190 1455 12220 1460
rect 12295 1480 12325 1485
rect 12295 1460 12300 1480
rect 12300 1460 12320 1480
rect 12320 1460 12325 1480
rect 12295 1455 12325 1460
rect 12405 1480 12435 1485
rect 12405 1460 12410 1480
rect 12410 1460 12430 1480
rect 12430 1460 12435 1480
rect 12405 1455 12435 1460
rect 12515 1480 12545 1485
rect 12515 1460 12520 1480
rect 12520 1460 12540 1480
rect 12540 1460 12545 1480
rect 12515 1455 12545 1460
rect 12625 1480 12655 1485
rect 12625 1460 12630 1480
rect 12630 1460 12650 1480
rect 12650 1460 12655 1480
rect 12625 1455 12655 1460
rect 11885 1355 11915 1385
rect 11430 1320 11460 1325
rect 11430 1300 11435 1320
rect 11435 1300 11455 1320
rect 11455 1300 11460 1320
rect 11430 1295 11460 1300
rect 11540 1320 11570 1325
rect 11540 1300 11545 1320
rect 11545 1300 11565 1320
rect 11565 1300 11570 1320
rect 11540 1295 11570 1300
rect 11650 1320 11680 1325
rect 11650 1300 11655 1320
rect 11655 1300 11675 1320
rect 11675 1300 11680 1320
rect 11650 1295 11680 1300
rect 11760 1320 11790 1325
rect 11760 1300 11765 1320
rect 11765 1300 11785 1320
rect 11785 1300 11790 1320
rect 11760 1295 11790 1300
rect 11870 1320 11900 1325
rect 11870 1300 11875 1320
rect 11875 1300 11895 1320
rect 11895 1300 11900 1320
rect 11870 1295 11900 1300
rect 11980 1320 12010 1325
rect 11980 1300 11985 1320
rect 11985 1300 12005 1320
rect 12005 1300 12010 1320
rect 11980 1295 12010 1300
rect 12090 1320 12120 1325
rect 12090 1300 12095 1320
rect 12095 1300 12115 1320
rect 12115 1300 12120 1320
rect 12090 1295 12120 1300
rect 12200 1320 12230 1325
rect 12200 1300 12205 1320
rect 12205 1300 12225 1320
rect 12225 1300 12230 1320
rect 12200 1295 12230 1300
rect 12310 1320 12340 1325
rect 12310 1300 12315 1320
rect 12315 1300 12335 1320
rect 12335 1300 12340 1320
rect 12310 1295 12340 1300
rect 12420 1320 12450 1325
rect 12420 1300 12425 1320
rect 12425 1300 12445 1320
rect 12445 1300 12450 1320
rect 12420 1295 12450 1300
rect 12530 1320 12560 1325
rect 12530 1300 12535 1320
rect 12535 1300 12555 1320
rect 12555 1300 12560 1320
rect 12530 1295 12560 1300
rect 3380 1180 3410 1185
rect 3380 1160 3385 1180
rect 3385 1160 3405 1180
rect 3405 1160 3410 1180
rect 3380 1155 3410 1160
rect 3990 1155 4020 1185
rect 4600 1180 4630 1185
rect 4600 1160 4605 1180
rect 4605 1160 4625 1180
rect 4625 1160 4630 1180
rect 4600 1155 4630 1160
rect 2950 1120 2980 1125
rect 2950 1100 2955 1120
rect 2955 1100 2975 1120
rect 2975 1100 2980 1120
rect 2950 1095 2980 1100
rect 3030 1120 3060 1125
rect 3030 1100 3035 1120
rect 3035 1100 3055 1120
rect 3055 1100 3060 1120
rect 3030 1095 3060 1100
rect 3110 1120 3140 1125
rect 3110 1100 3115 1120
rect 3115 1100 3135 1120
rect 3135 1100 3140 1120
rect 3110 1095 3140 1100
rect 3190 1120 3220 1125
rect 3190 1100 3195 1120
rect 3195 1100 3215 1120
rect 3215 1100 3220 1120
rect 3190 1095 3220 1100
rect 3270 1120 3300 1125
rect 3270 1100 3275 1120
rect 3275 1100 3295 1120
rect 3295 1100 3300 1120
rect 3270 1095 3300 1100
rect 3350 1120 3380 1125
rect 3350 1100 3355 1120
rect 3355 1100 3375 1120
rect 3375 1100 3380 1120
rect 3350 1095 3380 1100
rect 3430 1120 3460 1125
rect 3430 1100 3435 1120
rect 3435 1100 3455 1120
rect 3455 1100 3460 1120
rect 3430 1095 3460 1100
rect 3510 1120 3540 1125
rect 3510 1100 3515 1120
rect 3515 1100 3535 1120
rect 3535 1100 3540 1120
rect 3510 1095 3540 1100
rect 3590 1120 3620 1125
rect 3590 1100 3595 1120
rect 3595 1100 3615 1120
rect 3615 1100 3620 1120
rect 3590 1095 3620 1100
rect 3670 1120 3700 1125
rect 3670 1100 3675 1120
rect 3675 1100 3695 1120
rect 3695 1100 3700 1120
rect 3670 1095 3700 1100
rect 3750 1120 3780 1125
rect 3750 1100 3755 1120
rect 3755 1100 3775 1120
rect 3775 1100 3780 1120
rect 3750 1095 3780 1100
rect 3830 1120 3860 1125
rect 3830 1100 3835 1120
rect 3835 1100 3855 1120
rect 3855 1100 3860 1120
rect 3830 1095 3860 1100
rect 3910 1120 3940 1125
rect 3910 1100 3915 1120
rect 3915 1100 3935 1120
rect 3935 1100 3940 1120
rect 3910 1095 3940 1100
rect 3990 1120 4020 1125
rect 3990 1100 3995 1120
rect 3995 1100 4015 1120
rect 4015 1100 4020 1120
rect 3990 1095 4020 1100
rect 4070 1120 4100 1125
rect 4070 1100 4075 1120
rect 4075 1100 4095 1120
rect 4095 1100 4100 1120
rect 4070 1095 4100 1100
rect 4150 1120 4180 1125
rect 4150 1100 4155 1120
rect 4155 1100 4175 1120
rect 4175 1100 4180 1120
rect 4150 1095 4180 1100
rect 4230 1120 4260 1125
rect 4230 1100 4235 1120
rect 4235 1100 4255 1120
rect 4255 1100 4260 1120
rect 4230 1095 4260 1100
rect 4310 1120 4340 1125
rect 4310 1100 4315 1120
rect 4315 1100 4335 1120
rect 4335 1100 4340 1120
rect 4310 1095 4340 1100
rect 4390 1120 4420 1125
rect 4390 1100 4395 1120
rect 4395 1100 4415 1120
rect 4415 1100 4420 1120
rect 4390 1095 4420 1100
rect 4470 1120 4500 1125
rect 4470 1100 4475 1120
rect 4475 1100 4495 1120
rect 4495 1100 4500 1120
rect 4470 1095 4500 1100
rect 4550 1120 4580 1125
rect 4550 1100 4555 1120
rect 4555 1100 4575 1120
rect 4575 1100 4580 1120
rect 4550 1095 4580 1100
rect 4630 1120 4660 1125
rect 4630 1100 4635 1120
rect 4635 1100 4655 1120
rect 4655 1100 4660 1120
rect 4630 1095 4660 1100
rect 4710 1120 4740 1125
rect 4710 1100 4715 1120
rect 4715 1100 4735 1120
rect 4735 1100 4740 1120
rect 4710 1095 4740 1100
rect 4790 1120 4820 1125
rect 4790 1100 4795 1120
rect 4795 1100 4815 1120
rect 4815 1100 4820 1120
rect 4790 1095 4820 1100
rect 4870 1120 4900 1125
rect 4870 1100 4875 1120
rect 4875 1100 4895 1120
rect 4895 1100 4900 1120
rect 4870 1095 4900 1100
rect 4950 1120 4980 1125
rect 4950 1100 4955 1120
rect 4955 1100 4975 1120
rect 4975 1100 4980 1120
rect 4950 1095 4980 1100
rect 2625 1010 2655 1040
rect 2910 1035 2940 1040
rect 2910 1015 2915 1035
rect 2915 1015 2935 1035
rect 2935 1015 2940 1035
rect 2910 1010 2940 1015
rect 5115 1035 5145 1040
rect 5115 1015 5120 1035
rect 5120 1015 5140 1035
rect 5140 1015 5145 1035
rect 5115 1010 5145 1015
rect 11170 1000 11200 1005
rect 11170 980 11175 1000
rect 11175 980 11195 1000
rect 11195 980 11200 1000
rect 11170 975 11200 980
rect 11265 1000 11295 1005
rect 11265 980 11270 1000
rect 11270 980 11290 1000
rect 11290 980 11295 1000
rect 11265 975 11295 980
rect 11375 1000 11405 1005
rect 11375 980 11380 1000
rect 11380 980 11400 1000
rect 11400 980 11405 1000
rect 11375 975 11405 980
rect 11485 1000 11515 1005
rect 11485 980 11490 1000
rect 11490 980 11510 1000
rect 11510 980 11515 1000
rect 11485 975 11515 980
rect 11595 1000 11625 1005
rect 11595 980 11600 1000
rect 11600 980 11620 1000
rect 11620 980 11625 1000
rect 11595 975 11625 980
rect 11705 1000 11735 1005
rect 11705 980 11710 1000
rect 11710 980 11730 1000
rect 11730 980 11735 1000
rect 11705 975 11735 980
rect 11815 1000 11845 1005
rect 11815 980 11820 1000
rect 11820 980 11840 1000
rect 11840 980 11845 1000
rect 11815 975 11845 980
rect 11925 1000 11955 1005
rect 11925 980 11930 1000
rect 11930 980 11950 1000
rect 11950 980 11955 1000
rect 11925 975 11955 980
rect 12035 1000 12065 1005
rect 12035 980 12040 1000
rect 12040 980 12060 1000
rect 12060 980 12065 1000
rect 12035 975 12065 980
rect 12145 1000 12175 1005
rect 12145 980 12150 1000
rect 12150 980 12170 1000
rect 12170 980 12175 1000
rect 12145 975 12175 980
rect 12255 1000 12285 1005
rect 12255 980 12260 1000
rect 12260 980 12280 1000
rect 12280 980 12285 1000
rect 12255 975 12285 980
rect 12365 1000 12395 1005
rect 12365 980 12370 1000
rect 12370 980 12390 1000
rect 12390 980 12395 1000
rect 12365 975 12395 980
rect 12475 1000 12505 1005
rect 12475 980 12480 1000
rect 12480 980 12500 1000
rect 12500 980 12505 1000
rect 12475 975 12505 980
rect 12625 1000 12655 1005
rect 12625 980 12630 1000
rect 12630 980 12650 1000
rect 12650 980 12655 1000
rect 12625 975 12655 980
rect 3000 925 3030 930
rect 3000 905 3005 925
rect 3005 905 3025 925
rect 3025 905 3030 925
rect 3000 900 3030 905
rect 3180 925 3210 930
rect 3180 905 3185 925
rect 3185 905 3205 925
rect 3205 905 3210 925
rect 3180 900 3210 905
rect 3360 925 3390 930
rect 3360 905 3365 925
rect 3365 905 3385 925
rect 3385 905 3390 925
rect 3360 900 3390 905
rect 3540 925 3570 930
rect 3540 905 3545 925
rect 3545 905 3565 925
rect 3565 905 3570 925
rect 3540 900 3570 905
rect 3720 925 3750 930
rect 3720 905 3725 925
rect 3725 905 3745 925
rect 3745 905 3750 925
rect 3720 900 3750 905
rect 3900 925 3930 930
rect 3900 905 3905 925
rect 3905 905 3925 925
rect 3925 905 3930 925
rect 3900 900 3930 905
rect 4080 925 4110 930
rect 4080 905 4085 925
rect 4085 905 4105 925
rect 4105 905 4110 925
rect 4080 900 4110 905
rect 4260 925 4290 930
rect 4260 905 4265 925
rect 4265 905 4285 925
rect 4285 905 4290 925
rect 4260 900 4290 905
rect 4440 925 4470 930
rect 4440 905 4445 925
rect 4445 905 4465 925
rect 4465 905 4470 925
rect 4440 900 4470 905
rect 4620 925 4650 930
rect 4620 905 4625 925
rect 4625 905 4645 925
rect 4645 905 4650 925
rect 4620 900 4650 905
rect 4800 925 4830 930
rect 4800 905 4805 925
rect 4805 905 4825 925
rect 4825 905 4830 925
rect 4800 900 4830 905
rect 4980 925 5010 930
rect 4980 905 4985 925
rect 4985 905 5005 925
rect 5005 905 5010 925
rect 4980 900 5010 905
rect 2525 730 2555 760
rect 3135 755 3165 760
rect 3135 735 3140 755
rect 3140 735 3160 755
rect 3160 735 3165 755
rect 3135 730 3165 735
rect 3630 755 3660 760
rect 3630 735 3635 755
rect 3635 735 3655 755
rect 3655 735 3660 755
rect 3630 730 3660 735
rect 3990 755 4020 760
rect 3990 735 3995 755
rect 3995 735 4015 755
rect 4015 735 4020 755
rect 3990 730 4020 735
rect 4350 755 4380 760
rect 4350 735 4355 755
rect 4355 735 4375 755
rect 4375 735 4380 755
rect 4350 730 4380 735
rect 4530 755 4560 760
rect 4530 735 4535 755
rect 4535 735 4555 755
rect 4555 735 4560 755
rect 4530 730 4560 735
rect 4710 755 4740 760
rect 4710 735 4715 755
rect 4715 735 4735 755
rect 4735 735 4740 755
rect 4710 730 4740 735
rect 4890 755 4920 760
rect 4890 735 4895 755
rect 4895 735 4915 755
rect 4915 735 4920 755
rect 4890 730 4920 735
rect 3450 675 3480 705
rect 3810 675 3840 705
rect 4170 675 4200 705
<< metal2 >>
rect -195 4990 -155 4995
rect -195 4960 -190 4990
rect -160 4960 -155 4990
rect -195 4955 -155 4960
rect 5550 4990 5590 4995
rect 5550 4960 5555 4990
rect 5585 4960 5590 4990
rect 5550 4955 5590 4960
rect -110 3525 -70 3530
rect -110 3495 -105 3525
rect -75 3520 -70 3525
rect 1261 3525 1301 3530
rect 1261 3520 1266 3525
rect -75 3500 1266 3520
rect -75 3495 -70 3500
rect -110 3490 -70 3495
rect 1261 3495 1266 3500
rect 1296 3495 1301 3525
rect 1261 3490 1301 3495
rect 4440 3495 4480 3500
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect -15 3445 25 3450
rect -15 3415 -10 3445
rect 20 3440 25 3445
rect 940 3445 980 3450
rect 940 3440 945 3445
rect 20 3420 945 3440
rect 20 3415 25 3420
rect -15 3410 25 3415
rect 940 3415 945 3420
rect 975 3415 980 3445
rect 940 3410 980 3415
rect 1635 3445 1685 3455
rect 2470 3450 2510 3455
rect 2470 3445 2475 3450
rect 1635 3415 1645 3445
rect 1675 3425 2475 3445
rect 1675 3415 1685 3425
rect 2470 3420 2475 3425
rect 2505 3420 2510 3450
rect 2470 3415 2510 3420
rect 5135 3445 5185 3455
rect 5135 3415 5145 3445
rect 5175 3440 5185 3445
rect 5550 3445 5590 3450
rect 5550 3440 5555 3445
rect 5175 3420 5555 3440
rect 5175 3415 5185 3420
rect 1635 3405 1685 3415
rect 5135 3405 5185 3415
rect 5550 3415 5555 3420
rect 5585 3415 5590 3445
rect 5550 3410 5590 3415
rect -60 3390 -20 3395
rect -60 3360 -55 3390
rect -25 3385 -20 3390
rect 2690 3390 2730 3395
rect 2690 3385 2695 3390
rect -25 3365 2695 3385
rect -25 3360 -20 3365
rect -60 3355 -20 3360
rect 2690 3360 2695 3365
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 1205 3340 1245 3345
rect 1205 3310 1210 3340
rect 1240 3335 1245 3340
rect 3135 3340 3175 3345
rect 3135 3335 3140 3340
rect 1240 3315 3140 3335
rect 1240 3310 1245 3315
rect 1205 3305 1245 3310
rect 3135 3310 3140 3315
rect 3170 3310 3175 3340
rect 3135 3305 3175 3310
rect 3385 3335 3435 3345
rect 3385 3305 3395 3335
rect 3425 3330 3435 3335
rect 5360 3335 5400 3340
rect 5360 3330 5365 3335
rect 3425 3310 5365 3330
rect 3425 3305 3435 3310
rect 3385 3295 3435 3305
rect 5360 3305 5365 3310
rect 5395 3305 5400 3335
rect 5360 3300 5400 3305
rect 1160 3285 1200 3290
rect 1160 3255 1165 3285
rect 1195 3280 1200 3285
rect 4885 3285 4925 3290
rect 4885 3280 4890 3285
rect 1195 3260 4890 3280
rect 1195 3255 1200 3260
rect 1160 3250 1200 3255
rect 4885 3255 4890 3260
rect 4920 3280 4925 3285
rect 5410 3285 5450 3290
rect 5410 3280 5415 3285
rect 4920 3260 5415 3280
rect 4920 3255 4925 3260
rect 4885 3250 4925 3255
rect 5410 3255 5415 3260
rect 5445 3255 5450 3285
rect 5410 3250 5450 3255
rect 2735 3240 2775 3245
rect 2735 3235 2740 3240
rect 46 3215 2740 3235
rect 46 3205 91 3215
rect 2735 3210 2740 3215
rect 2770 3210 2775 3240
rect 2735 3205 2775 3210
rect 46 3170 51 3205
rect 86 3170 91 3205
rect 1261 3165 1266 3200
rect 1301 3165 1306 3200
rect 2620 3185 2660 3190
rect 2620 3155 2625 3185
rect 2655 3180 2660 3185
rect 4440 3185 4480 3190
rect 4440 3180 4445 3185
rect 2655 3160 4445 3180
rect 2655 3155 2660 3160
rect 2620 3150 2660 3155
rect 4440 3155 4445 3160
rect 4475 3155 4480 3185
rect 4440 3150 4480 3155
rect -110 3140 -70 3145
rect -110 3110 -105 3140
rect -75 3135 -70 3140
rect 46 3135 51 3145
rect -75 3115 51 3135
rect -75 3110 -70 3115
rect 46 3110 51 3115
rect 86 3110 91 3145
rect 3135 3140 3175 3145
rect -110 3105 -70 3110
rect 1261 3105 1266 3140
rect 1301 3105 1306 3140
rect 3135 3110 3140 3140
rect 3170 3135 3175 3140
rect 4835 3140 4875 3145
rect 4835 3135 4840 3140
rect 3170 3115 4840 3135
rect 3170 3110 3175 3115
rect 3135 3105 3175 3110
rect 4835 3110 4840 3115
rect 4870 3135 4875 3140
rect 5315 3140 5355 3145
rect 5315 3135 5320 3140
rect 4870 3115 5320 3135
rect 4870 3110 4875 3115
rect 4835 3105 4875 3110
rect 5315 3110 5320 3115
rect 5350 3110 5355 3140
rect 5315 3105 5355 3110
rect 1160 3100 1200 3105
rect 1160 3095 1165 3100
rect 46 3075 1165 3095
rect 46 3065 91 3075
rect 1160 3070 1165 3075
rect 1195 3070 1200 3100
rect 1160 3065 1200 3070
rect 3985 3080 4025 3085
rect 46 3030 51 3065
rect 86 3030 91 3065
rect 3985 3050 3990 3080
rect 4020 3075 4025 3080
rect 4020 3055 6100 3075
rect 4020 3050 4025 3055
rect 3985 3045 4025 3050
rect 3445 3035 3485 3040
rect 3445 3005 3450 3035
rect 3480 3030 3485 3035
rect 3805 3035 3845 3040
rect 3805 3030 3810 3035
rect 3480 3010 3810 3030
rect 3480 3005 3485 3010
rect -110 3000 -70 3005
rect -110 2970 -105 3000
rect -75 2995 -70 3000
rect 46 2995 51 3005
rect -75 2975 51 2995
rect -75 2970 -70 2975
rect 46 2970 51 2975
rect 86 2970 91 3005
rect 3445 3000 3485 3005
rect 3805 3005 3810 3010
rect 3840 3030 3845 3035
rect 4345 3035 4385 3040
rect 4345 3030 4350 3035
rect 3840 3010 4350 3030
rect 3840 3005 3845 3010
rect 3805 3000 3845 3005
rect 4345 3005 4350 3010
rect 4380 3030 4385 3035
rect 4705 3035 4745 3040
rect 4705 3030 4710 3035
rect 4380 3010 4710 3030
rect 4380 3005 4385 3010
rect 4345 3000 4385 3005
rect 4705 3005 4710 3010
rect 4740 3030 4745 3035
rect 4740 3010 6100 3030
rect 4740 3005 4745 3010
rect 4705 3000 4745 3005
rect 2520 2980 2560 2985
rect -110 2965 -70 2970
rect 2330 2925 2335 2960
rect 2370 2950 2375 2960
rect 2425 2955 2465 2960
rect 2425 2950 2430 2955
rect 2370 2930 2430 2950
rect 2370 2925 2375 2930
rect 2425 2925 2430 2930
rect 2460 2925 2465 2955
rect 2520 2950 2525 2980
rect 2555 2975 2560 2980
rect 3080 2980 3120 2985
rect 3080 2975 3085 2980
rect 2555 2955 3085 2975
rect 2555 2950 2560 2955
rect 2520 2945 2560 2950
rect 3080 2950 3085 2955
rect 3115 2950 3120 2980
rect 3080 2945 3120 2950
rect 3265 2980 3305 2985
rect 3265 2950 3270 2980
rect 3300 2975 3305 2980
rect 3625 2980 3665 2985
rect 3625 2975 3630 2980
rect 3300 2955 3630 2975
rect 3300 2950 3305 2955
rect 3265 2945 3305 2950
rect 3625 2950 3630 2955
rect 3660 2975 3665 2980
rect 4165 2980 4205 2985
rect 4165 2975 4170 2980
rect 3660 2955 4170 2975
rect 3660 2950 3665 2955
rect 3625 2945 3665 2950
rect 4165 2950 4170 2955
rect 4200 2975 4205 2980
rect 4525 2980 4565 2985
rect 4525 2975 4530 2980
rect 4200 2955 4530 2975
rect 4200 2950 4205 2955
rect 4165 2945 4205 2950
rect 4525 2950 4530 2955
rect 4560 2975 4565 2980
rect 4560 2955 6100 2975
rect 4560 2950 4565 2955
rect 4525 2945 4565 2950
rect 2425 2920 2465 2925
rect -110 2910 -70 2915
rect -110 2880 -105 2910
rect -75 2905 -70 2910
rect 905 2910 1125 2920
rect 905 2905 920 2910
rect -75 2885 920 2905
rect -75 2880 -70 2885
rect -110 2875 -70 2880
rect 905 2880 920 2885
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1125 2910
rect 905 2870 1125 2880
rect 2330 2900 2375 2905
rect 2330 2865 2335 2900
rect 2370 2865 2375 2900
rect 2330 2860 2375 2865
rect -60 2855 -20 2860
rect -60 2825 -55 2855
rect -25 2850 -20 2855
rect 51 2850 56 2855
rect -25 2830 56 2850
rect -25 2825 -20 2830
rect -60 2820 -20 2825
rect 51 2820 56 2830
rect 91 2820 96 2855
rect 724 2820 729 2855
rect 764 2845 769 2855
rect 1205 2850 1245 2855
rect 1205 2845 1210 2850
rect 764 2825 1210 2845
rect 764 2820 769 2825
rect 1205 2820 1210 2825
rect 1240 2820 1245 2850
rect 1205 2815 1245 2820
rect 1261 2805 1266 2840
rect 1301 2805 1306 2840
rect 1960 2805 1965 2840
rect 2000 2830 2005 2840
rect 2330 2835 2370 2840
rect 2330 2830 2335 2835
rect 2000 2810 2335 2830
rect 2000 2805 2005 2810
rect 2330 2805 2335 2810
rect 2365 2805 2370 2835
rect 2330 2800 2370 2805
rect 2995 2810 3035 2815
rect -15 2795 25 2800
rect -15 2765 -10 2795
rect 20 2785 25 2795
rect 51 2785 56 2795
rect 20 2765 56 2785
rect -15 2760 25 2765
rect 51 2760 56 2765
rect 91 2760 96 2795
rect 724 2760 729 2795
rect 764 2785 769 2795
rect 2620 2790 2660 2795
rect 2620 2785 2625 2790
rect 764 2765 2625 2785
rect 764 2760 769 2765
rect 2620 2760 2625 2765
rect 2655 2760 2660 2790
rect 2995 2780 3000 2810
rect 3030 2805 3035 2810
rect 3175 2810 3215 2815
rect 3175 2805 3180 2810
rect 3030 2785 3180 2805
rect 3030 2780 3035 2785
rect 2995 2775 3035 2780
rect 3175 2780 3180 2785
rect 3210 2805 3215 2810
rect 3355 2810 3395 2815
rect 3355 2805 3360 2810
rect 3210 2785 3360 2805
rect 3210 2780 3215 2785
rect 3175 2775 3215 2780
rect 3355 2780 3360 2785
rect 3390 2805 3395 2810
rect 3535 2810 3575 2815
rect 3535 2805 3540 2810
rect 3390 2785 3540 2805
rect 3390 2780 3395 2785
rect 3355 2775 3395 2780
rect 3535 2780 3540 2785
rect 3570 2805 3575 2810
rect 3715 2810 3755 2815
rect 3715 2805 3720 2810
rect 3570 2785 3720 2805
rect 3570 2780 3575 2785
rect 3535 2775 3575 2780
rect 3715 2780 3720 2785
rect 3750 2805 3755 2810
rect 3895 2810 3935 2815
rect 3895 2805 3900 2810
rect 3750 2785 3900 2805
rect 3750 2780 3755 2785
rect 3715 2775 3755 2780
rect 3895 2780 3900 2785
rect 3930 2805 3935 2810
rect 4075 2810 4115 2815
rect 4075 2805 4080 2810
rect 3930 2785 4080 2805
rect 3930 2780 3935 2785
rect 3895 2775 3935 2780
rect 4075 2780 4080 2785
rect 4110 2805 4115 2810
rect 4255 2810 4295 2815
rect 4255 2805 4260 2810
rect 4110 2785 4260 2805
rect 4110 2780 4115 2785
rect 4075 2775 4115 2780
rect 4255 2780 4260 2785
rect 4290 2805 4295 2810
rect 4435 2810 4475 2815
rect 4435 2805 4440 2810
rect 4290 2785 4440 2805
rect 4290 2780 4295 2785
rect 4255 2775 4295 2780
rect 4435 2780 4440 2785
rect 4470 2805 4475 2810
rect 4615 2810 4655 2815
rect 4615 2805 4620 2810
rect 4470 2785 4620 2805
rect 4470 2780 4475 2785
rect 4435 2775 4475 2780
rect 4615 2780 4620 2785
rect 4650 2805 4655 2810
rect 4795 2810 4835 2815
rect 4795 2805 4800 2810
rect 4650 2785 4800 2805
rect 4650 2780 4655 2785
rect 4615 2775 4655 2780
rect 4795 2780 4800 2785
rect 4830 2805 4835 2810
rect 4975 2810 5015 2815
rect 4975 2805 4980 2810
rect 4830 2785 4980 2805
rect 4830 2780 4835 2785
rect 4795 2775 4835 2780
rect 4975 2780 4980 2785
rect 5010 2805 5015 2810
rect 5550 2810 5590 2815
rect 5550 2805 5555 2810
rect 5010 2785 5555 2805
rect 5010 2780 5015 2785
rect 4975 2775 5015 2780
rect 5550 2780 5555 2785
rect 5585 2780 5590 2810
rect 5550 2775 5590 2780
rect 2620 2755 2660 2760
rect 3175 2750 3215 2755
rect 1261 2745 1301 2750
rect 1261 2715 1266 2745
rect 1296 2740 1301 2745
rect 2150 2745 2190 2750
rect 2150 2740 2155 2745
rect 1296 2720 2155 2740
rect 1296 2715 1301 2720
rect 1261 2710 1301 2715
rect 2150 2715 2155 2720
rect 2185 2715 2190 2745
rect 3175 2720 3180 2750
rect 3210 2745 3215 2750
rect 3355 2750 3395 2755
rect 3355 2745 3360 2750
rect 3210 2725 3360 2745
rect 3210 2720 3215 2725
rect 3175 2715 3215 2720
rect 3355 2720 3360 2725
rect 3390 2745 3395 2750
rect 3535 2750 3575 2755
rect 3535 2745 3540 2750
rect 3390 2725 3540 2745
rect 3390 2720 3395 2725
rect 3355 2715 3395 2720
rect 3535 2720 3540 2725
rect 3570 2745 3575 2750
rect 3715 2750 3755 2755
rect 3715 2745 3720 2750
rect 3570 2725 3720 2745
rect 3570 2720 3575 2725
rect 3535 2715 3575 2720
rect 3715 2720 3720 2725
rect 3750 2745 3755 2750
rect 3895 2750 3935 2755
rect 3895 2745 3900 2750
rect 3750 2725 3900 2745
rect 3750 2720 3755 2725
rect 3715 2715 3755 2720
rect 3895 2720 3900 2725
rect 3930 2745 3935 2750
rect 4075 2750 4115 2755
rect 4075 2745 4080 2750
rect 3930 2725 4080 2745
rect 3930 2720 3935 2725
rect 3895 2715 3935 2720
rect 4075 2720 4080 2725
rect 4110 2745 4115 2750
rect 4255 2750 4295 2755
rect 4255 2745 4260 2750
rect 4110 2725 4260 2745
rect 4110 2720 4115 2725
rect 4075 2715 4115 2720
rect 4255 2720 4260 2725
rect 4290 2745 4295 2750
rect 4435 2750 4475 2755
rect 4435 2745 4440 2750
rect 4290 2725 4440 2745
rect 4290 2720 4295 2725
rect 4255 2715 4295 2720
rect 4435 2720 4440 2725
rect 4470 2745 4475 2750
rect 4615 2750 4655 2755
rect 4615 2745 4620 2750
rect 4470 2725 4620 2745
rect 4470 2720 4475 2725
rect 4435 2715 4475 2720
rect 4615 2720 4620 2725
rect 4650 2745 4655 2750
rect 4795 2750 4835 2755
rect 4795 2745 4800 2750
rect 4650 2725 4800 2745
rect 4650 2720 4655 2725
rect 4615 2715 4655 2720
rect 4795 2720 4800 2725
rect 4830 2720 4835 2750
rect 4795 2715 4835 2720
rect 2150 2710 2190 2715
rect 3805 2380 3845 2385
rect 3355 2375 3395 2380
rect 2620 2345 2660 2350
rect 2620 2315 2625 2345
rect 2655 2340 2660 2345
rect 3355 2345 3360 2375
rect 3390 2345 3395 2375
rect 3805 2350 3810 2380
rect 3840 2375 3845 2380
rect 4165 2380 4205 2385
rect 4165 2375 4170 2380
rect 3840 2355 4170 2375
rect 3840 2350 3845 2355
rect 3805 2345 3845 2350
rect 4165 2350 4170 2355
rect 4200 2350 4205 2380
rect 4165 2345 4205 2350
rect 3355 2340 3395 2345
rect 2655 2320 3395 2340
rect 3625 2335 3665 2340
rect 2655 2315 2660 2320
rect 2620 2310 2660 2315
rect 3625 2305 3630 2335
rect 3660 2330 3665 2335
rect 4345 2335 4385 2340
rect 4345 2330 4350 2335
rect 3660 2310 4350 2330
rect 3660 2305 3665 2310
rect 3625 2300 3665 2305
rect 4345 2305 4350 2310
rect 4380 2305 4385 2335
rect 4345 2300 4385 2305
rect 2735 2290 2775 2295
rect 2735 2260 2740 2290
rect 2770 2285 2775 2290
rect 3445 2290 3485 2295
rect 3445 2285 3450 2290
rect 2770 2265 3450 2285
rect 2770 2260 2775 2265
rect 2735 2255 2775 2260
rect 3445 2260 3450 2265
rect 3480 2285 3485 2290
rect 4525 2290 4565 2295
rect 4525 2285 4530 2290
rect 3480 2265 4530 2285
rect 3480 2260 3485 2265
rect 3445 2255 3485 2260
rect 4525 2260 4530 2265
rect 4560 2285 4565 2290
rect 5270 2290 5310 2295
rect 5270 2285 5275 2290
rect 4560 2265 5275 2285
rect 4560 2260 4565 2265
rect 4525 2255 4565 2260
rect 5270 2260 5275 2265
rect 5305 2260 5310 2290
rect 5270 2255 5310 2260
rect 2425 2245 2465 2250
rect 2425 2215 2430 2245
rect 2460 2240 2465 2245
rect 3805 2245 3845 2250
rect 3805 2240 3810 2245
rect 2460 2220 3810 2240
rect 2460 2215 2465 2220
rect 2425 2210 2465 2215
rect 3805 2215 3810 2220
rect 3840 2215 3845 2245
rect 3805 2210 3845 2215
rect 2330 2200 2370 2205
rect 2330 2170 2335 2200
rect 2365 2195 2370 2200
rect 3265 2200 3305 2205
rect 3265 2195 3270 2200
rect 2365 2175 3270 2195
rect 2365 2170 2370 2175
rect 2330 2165 2370 2170
rect 3265 2170 3270 2175
rect 3300 2195 3305 2200
rect 3985 2200 4025 2205
rect 3985 2195 3990 2200
rect 3300 2175 3990 2195
rect 3300 2170 3305 2175
rect 3265 2165 3305 2170
rect 3985 2170 3990 2175
rect 4020 2195 4025 2200
rect 4705 2200 4745 2205
rect 4705 2195 4710 2200
rect 4020 2175 4710 2195
rect 4020 2170 4025 2175
rect 3985 2165 4025 2170
rect 4705 2170 4710 2175
rect 4740 2170 4745 2200
rect 4705 2165 4745 2170
rect 2380 2150 2420 2155
rect 2380 2120 2385 2150
rect 2415 2145 2420 2150
rect 3625 2150 3665 2155
rect 3625 2145 3630 2150
rect 2415 2125 3630 2145
rect 2415 2120 2420 2125
rect 2380 2115 2420 2120
rect 3625 2120 3630 2125
rect 3660 2120 3665 2150
rect 3625 2115 3665 2120
rect 4085 2145 4125 2150
rect 4085 2115 4090 2145
rect 4120 2140 4125 2145
rect 5315 2145 5355 2150
rect 5315 2140 5320 2145
rect 4120 2120 5320 2140
rect 4120 2115 4125 2120
rect 4085 2110 4125 2115
rect 5315 2115 5320 2120
rect 5350 2115 5355 2145
rect 5315 2110 5355 2115
rect 2745 2095 2785 2100
rect 2745 2065 2750 2095
rect 2780 2090 2785 2095
rect 2865 2095 2905 2100
rect 2865 2090 2870 2095
rect 2780 2070 2870 2090
rect 2780 2065 2785 2070
rect 2745 2060 2785 2065
rect 2865 2065 2870 2070
rect 2900 2090 2905 2095
rect 2985 2095 3025 2100
rect 2985 2090 2990 2095
rect 2900 2070 2990 2090
rect 2900 2065 2905 2070
rect 2865 2060 2905 2065
rect 2985 2065 2990 2070
rect 3020 2090 3025 2095
rect 3105 2095 3145 2100
rect 3105 2090 3110 2095
rect 3020 2070 3110 2090
rect 3020 2065 3025 2070
rect 2985 2060 3025 2065
rect 3105 2065 3110 2070
rect 3140 2090 3145 2095
rect 3225 2095 3265 2100
rect 3225 2090 3230 2095
rect 3140 2070 3230 2090
rect 3140 2065 3145 2070
rect 3105 2060 3145 2065
rect 3225 2065 3230 2070
rect 3260 2090 3265 2095
rect 3345 2095 3385 2100
rect 3345 2090 3350 2095
rect 3260 2070 3350 2090
rect 3260 2065 3265 2070
rect 3225 2060 3265 2065
rect 3345 2065 3350 2070
rect 3380 2090 3385 2095
rect 3465 2095 3505 2100
rect 3465 2090 3470 2095
rect 3380 2070 3470 2090
rect 3380 2065 3385 2070
rect 3345 2060 3385 2065
rect 3465 2065 3470 2070
rect 3500 2090 3505 2095
rect 3585 2095 3625 2100
rect 3585 2090 3590 2095
rect 3500 2070 3590 2090
rect 3500 2065 3505 2070
rect 3465 2060 3505 2065
rect 3585 2065 3590 2070
rect 3620 2090 3625 2095
rect 3705 2095 3745 2100
rect 3705 2090 3710 2095
rect 3620 2070 3710 2090
rect 3620 2065 3625 2070
rect 3585 2060 3625 2065
rect 3705 2065 3710 2070
rect 3740 2090 3745 2095
rect 3825 2095 3865 2100
rect 3825 2090 3830 2095
rect 3740 2070 3830 2090
rect 3740 2065 3745 2070
rect 3705 2060 3745 2065
rect 3825 2065 3830 2070
rect 3860 2090 3865 2095
rect 3985 2095 4025 2100
rect 3985 2090 3990 2095
rect 3860 2070 3990 2090
rect 3860 2065 3865 2070
rect 3825 2060 3865 2065
rect 3985 2065 3990 2070
rect 4020 2090 4025 2095
rect 4145 2095 4185 2100
rect 4145 2090 4150 2095
rect 4020 2070 4150 2090
rect 4020 2065 4025 2070
rect 3985 2060 4025 2065
rect 4145 2065 4150 2070
rect 4180 2090 4185 2095
rect 4265 2095 4305 2100
rect 4265 2090 4270 2095
rect 4180 2070 4270 2090
rect 4180 2065 4185 2070
rect 4145 2060 4185 2065
rect 4265 2065 4270 2070
rect 4300 2090 4305 2095
rect 4385 2095 4425 2100
rect 4385 2090 4390 2095
rect 4300 2070 4390 2090
rect 4300 2065 4305 2070
rect 4265 2060 4305 2065
rect 4385 2065 4390 2070
rect 4420 2090 4425 2095
rect 4505 2095 4545 2100
rect 4505 2090 4510 2095
rect 4420 2070 4510 2090
rect 4420 2065 4425 2070
rect 4385 2060 4425 2065
rect 4505 2065 4510 2070
rect 4540 2090 4545 2095
rect 4625 2095 4665 2100
rect 4625 2090 4630 2095
rect 4540 2070 4630 2090
rect 4540 2065 4545 2070
rect 4505 2060 4545 2065
rect 4625 2065 4630 2070
rect 4660 2090 4665 2095
rect 4745 2095 4785 2100
rect 4745 2090 4750 2095
rect 4660 2070 4750 2090
rect 4660 2065 4665 2070
rect 4625 2060 4665 2065
rect 4745 2065 4750 2070
rect 4780 2090 4785 2095
rect 4865 2095 4905 2100
rect 4865 2090 4870 2095
rect 4780 2070 4870 2090
rect 4780 2065 4785 2070
rect 4745 2060 4785 2065
rect 4865 2065 4870 2070
rect 4900 2090 4905 2095
rect 4985 2095 5025 2100
rect 4985 2090 4990 2095
rect 4900 2070 4990 2090
rect 4900 2065 4905 2070
rect 4865 2060 4905 2065
rect 4985 2065 4990 2070
rect 5020 2090 5025 2095
rect 5105 2095 5145 2100
rect 5105 2090 5110 2095
rect 5020 2070 5110 2090
rect 5020 2065 5025 2070
rect 4985 2060 5025 2065
rect 5105 2065 5110 2070
rect 5140 2090 5145 2095
rect 5225 2095 5265 2100
rect 5225 2090 5230 2095
rect 5140 2070 5230 2090
rect 5140 2065 5145 2070
rect 5105 2060 5145 2065
rect 5225 2065 5230 2070
rect 5260 2090 5265 2095
rect 5550 2095 5590 2100
rect 5550 2090 5555 2095
rect 5260 2070 5555 2090
rect 5260 2065 5265 2070
rect 5225 2060 5265 2065
rect 5550 2065 5555 2070
rect 5585 2065 5590 2095
rect 5550 2060 5590 2065
rect 2620 2050 2660 2055
rect 2620 2020 2625 2050
rect 2655 2020 2660 2050
rect 2620 2015 2660 2020
rect 2805 2050 2845 2055
rect 2805 2020 2810 2050
rect 2840 2045 2845 2050
rect 3165 2050 3205 2055
rect 3165 2045 3170 2050
rect 2840 2025 3170 2045
rect 2840 2020 2845 2025
rect 2805 2015 2845 2020
rect 3165 2020 3170 2025
rect 3200 2045 3205 2050
rect 3525 2050 3565 2055
rect 3525 2045 3530 2050
rect 3200 2025 3530 2045
rect 3200 2020 3205 2025
rect 3165 2015 3205 2020
rect 3525 2020 3530 2025
rect 3560 2045 3565 2050
rect 3885 2050 3925 2055
rect 3885 2045 3890 2050
rect 3560 2025 3890 2045
rect 3560 2020 3565 2025
rect 3525 2015 3565 2020
rect 3885 2020 3890 2025
rect 3920 2020 3925 2050
rect 3885 2015 3925 2020
rect 4085 2050 4125 2055
rect 4085 2020 4090 2050
rect 4120 2045 4125 2050
rect 4445 2050 4485 2055
rect 4445 2045 4450 2050
rect 4120 2025 4450 2045
rect 4120 2020 4125 2025
rect 4085 2015 4125 2020
rect 4445 2020 4450 2025
rect 4480 2045 4485 2050
rect 4805 2050 4845 2055
rect 4805 2045 4810 2050
rect 4480 2025 4810 2045
rect 4480 2020 4485 2025
rect 4445 2015 4485 2020
rect 4805 2020 4810 2025
rect 4840 2045 4845 2050
rect 5165 2050 5205 2055
rect 5165 2045 5170 2050
rect 4840 2025 5170 2045
rect 4840 2020 4845 2025
rect 4805 2015 4845 2020
rect 5165 2020 5170 2025
rect 5200 2020 5205 2050
rect 5165 2015 5205 2020
rect 11190 1900 11230 1905
rect 2925 1880 2965 1885
rect 2925 1850 2930 1880
rect 2960 1875 2965 1880
rect 3045 1875 3085 1885
rect 3285 1880 3325 1885
rect 3285 1875 3290 1880
rect 2960 1855 3290 1875
rect 2960 1850 2965 1855
rect 2925 1845 2965 1850
rect 3045 1845 3085 1855
rect 3285 1850 3290 1855
rect 3320 1875 3325 1880
rect 3405 1875 3445 1885
rect 3645 1880 3685 1885
rect 3645 1875 3650 1880
rect 3320 1855 3650 1875
rect 3320 1850 3325 1855
rect 3285 1845 3325 1850
rect 3405 1845 3445 1855
rect 3645 1850 3650 1855
rect 3680 1850 3685 1880
rect 3645 1845 3685 1850
rect 3765 1845 3805 1885
rect 4205 1845 4245 1885
rect 4325 1880 4365 1885
rect 4325 1850 4330 1880
rect 4360 1875 4365 1880
rect 4565 1875 4605 1885
rect 4685 1880 4725 1885
rect 4685 1875 4690 1880
rect 4360 1855 4690 1875
rect 4360 1850 4365 1855
rect 4325 1845 4365 1850
rect 4565 1845 4605 1855
rect 4685 1850 4690 1855
rect 4720 1875 4725 1880
rect 4925 1875 4965 1885
rect 5045 1880 5085 1885
rect 5045 1875 5050 1880
rect 4720 1855 5050 1875
rect 4720 1850 4725 1855
rect 4685 1845 4725 1850
rect 4925 1845 4965 1855
rect 5045 1850 5050 1855
rect 5080 1875 5085 1880
rect 5080 1855 5175 1875
rect 11190 1870 11195 1900
rect 11225 1895 11230 1900
rect 11410 1900 11450 1905
rect 11410 1895 11415 1900
rect 11225 1875 11415 1895
rect 11225 1870 11230 1875
rect 11190 1865 11230 1870
rect 11410 1870 11415 1875
rect 11445 1895 11450 1900
rect 11640 1900 11680 1905
rect 11640 1895 11645 1900
rect 11445 1875 11645 1895
rect 11445 1870 11450 1875
rect 11410 1865 11450 1870
rect 11640 1870 11645 1875
rect 11675 1895 11680 1900
rect 12230 1900 12270 1905
rect 12230 1895 12235 1900
rect 11675 1875 12235 1895
rect 11675 1870 11680 1875
rect 11640 1865 11680 1870
rect 12230 1870 12235 1875
rect 12265 1895 12270 1900
rect 12450 1900 12490 1905
rect 12450 1895 12455 1900
rect 12265 1875 12455 1895
rect 12265 1870 12270 1875
rect 12230 1865 12270 1870
rect 12450 1870 12455 1875
rect 12485 1895 12490 1900
rect 12680 1900 12720 1905
rect 12680 1895 12685 1900
rect 12485 1875 12685 1895
rect 12485 1870 12490 1875
rect 12450 1865 12490 1870
rect 12680 1870 12685 1875
rect 12715 1870 12720 1900
rect 12680 1865 12720 1870
rect 11820 1855 11860 1860
rect 5080 1850 5085 1855
rect 5045 1845 5085 1850
rect 11820 1825 11825 1855
rect 11855 1850 11860 1855
rect 11940 1855 11980 1860
rect 11940 1850 11945 1855
rect 11855 1830 11945 1850
rect 11855 1825 11860 1830
rect 2470 1820 2510 1825
rect 2470 1790 2475 1820
rect 2505 1815 2510 1820
rect 2835 1820 2875 1825
rect 2835 1815 2840 1820
rect 2505 1795 2840 1815
rect 2505 1790 2510 1795
rect 2470 1785 2510 1790
rect 2835 1790 2840 1795
rect 2870 1815 2875 1820
rect 3045 1820 3085 1825
rect 3045 1815 3050 1820
rect 2870 1795 3050 1815
rect 2870 1790 2875 1795
rect 2835 1785 2875 1790
rect 3045 1790 3050 1795
rect 3080 1815 3085 1820
rect 3165 1820 3205 1825
rect 3165 1815 3170 1820
rect 3080 1795 3170 1815
rect 3080 1790 3085 1795
rect 3045 1785 3085 1790
rect 3165 1790 3170 1795
rect 3200 1815 3205 1820
rect 3405 1820 3445 1825
rect 3405 1815 3410 1820
rect 3200 1795 3410 1815
rect 3200 1790 3205 1795
rect 3165 1785 3205 1790
rect 3405 1790 3410 1795
rect 3440 1815 3445 1820
rect 3525 1820 3565 1825
rect 3525 1815 3530 1820
rect 3440 1795 3530 1815
rect 3440 1790 3445 1795
rect 3405 1785 3445 1790
rect 3525 1790 3530 1795
rect 3560 1815 3565 1820
rect 3765 1820 3805 1825
rect 3765 1815 3770 1820
rect 3560 1795 3770 1815
rect 3560 1790 3565 1795
rect 3525 1785 3565 1790
rect 3765 1790 3770 1795
rect 3800 1815 3805 1820
rect 3855 1820 3895 1825
rect 3855 1815 3860 1820
rect 3800 1795 3860 1815
rect 3800 1790 3805 1795
rect 3765 1785 3805 1790
rect 3855 1790 3860 1795
rect 3890 1790 3895 1820
rect 3855 1785 3895 1790
rect 4115 1820 4155 1825
rect 4115 1790 4120 1820
rect 4150 1815 4155 1820
rect 4205 1820 4245 1825
rect 4205 1815 4210 1820
rect 4150 1795 4210 1815
rect 4150 1790 4155 1795
rect 4115 1785 4155 1790
rect 4205 1790 4210 1795
rect 4240 1815 4245 1820
rect 4445 1820 4485 1825
rect 4445 1815 4450 1820
rect 4240 1795 4450 1815
rect 4240 1790 4245 1795
rect 4205 1785 4245 1790
rect 4445 1790 4450 1795
rect 4480 1815 4485 1820
rect 4565 1820 4605 1825
rect 4565 1815 4570 1820
rect 4480 1795 4570 1815
rect 4480 1790 4485 1795
rect 4445 1785 4485 1790
rect 4565 1790 4570 1795
rect 4600 1815 4605 1820
rect 4805 1820 4845 1825
rect 4805 1815 4810 1820
rect 4600 1795 4810 1815
rect 4600 1790 4605 1795
rect 4565 1785 4605 1790
rect 4805 1790 4810 1795
rect 4840 1815 4845 1820
rect 4925 1820 4965 1825
rect 4925 1815 4930 1820
rect 4840 1795 4930 1815
rect 4840 1790 4845 1795
rect 4805 1785 4845 1790
rect 4925 1790 4930 1795
rect 4960 1815 4965 1820
rect 5135 1820 5175 1825
rect 5135 1815 5140 1820
rect 4960 1795 5140 1815
rect 4960 1790 4965 1795
rect 4925 1785 4965 1790
rect 5135 1790 5140 1795
rect 5170 1815 5175 1820
rect 5360 1820 5400 1825
rect 11820 1820 11860 1825
rect 11940 1825 11945 1830
rect 11975 1825 11980 1855
rect 11940 1820 11980 1825
rect 5360 1815 5365 1820
rect 5170 1795 5365 1815
rect 5170 1790 5175 1795
rect 5135 1785 5175 1790
rect 5360 1790 5365 1795
rect 5395 1790 5400 1820
rect 5360 1785 5400 1790
rect 11085 1810 11125 1815
rect 11085 1780 11090 1810
rect 11120 1805 11125 1810
rect 11305 1810 11345 1815
rect 11305 1805 11310 1810
rect 11120 1785 11310 1805
rect 11120 1780 11125 1785
rect 11085 1775 11125 1780
rect 11305 1780 11310 1785
rect 11340 1805 11345 1810
rect 11525 1810 11565 1815
rect 11525 1805 11530 1810
rect 11340 1785 11530 1805
rect 11340 1780 11345 1785
rect 11305 1775 11345 1780
rect 11525 1780 11530 1785
rect 11560 1805 11565 1810
rect 12125 1810 12165 1815
rect 12125 1805 12130 1810
rect 11560 1785 12130 1805
rect 11560 1780 11565 1785
rect 11525 1775 11565 1780
rect 12125 1780 12130 1785
rect 12160 1805 12165 1810
rect 12345 1810 12385 1815
rect 12345 1805 12350 1810
rect 12160 1785 12350 1805
rect 12160 1780 12165 1785
rect 12125 1775 12165 1780
rect 12345 1780 12350 1785
rect 12380 1805 12385 1810
rect 12565 1810 12605 1815
rect 12565 1805 12570 1810
rect 12380 1785 12570 1805
rect 12380 1780 12385 1785
rect 12345 1775 12385 1780
rect 12565 1780 12570 1785
rect 12600 1780 12605 1810
rect 12565 1775 12605 1780
rect 2800 1765 2840 1770
rect 11237 1765 11269 1770
rect 2425 1760 2465 1765
rect 2425 1730 2430 1760
rect 2460 1755 2465 1760
rect 2565 1760 2605 1765
rect 2565 1755 2570 1760
rect 2460 1735 2570 1755
rect 2460 1730 2465 1735
rect 2425 1725 2465 1730
rect 2565 1730 2570 1735
rect 2600 1755 2605 1760
rect 2675 1760 2715 1765
rect 2675 1755 2680 1760
rect 2600 1735 2680 1755
rect 2600 1730 2605 1735
rect 2565 1725 2605 1730
rect 2675 1730 2680 1735
rect 2710 1755 2715 1760
rect 2800 1755 2805 1765
rect 2710 1735 2805 1755
rect 2835 1755 2840 1765
rect 3225 1760 3265 1765
rect 3225 1755 3230 1760
rect 2835 1735 3230 1755
rect 2710 1730 2715 1735
rect 2800 1730 2840 1735
rect 3225 1730 3230 1735
rect 3260 1730 3265 1760
rect 2675 1725 2715 1730
rect 3225 1725 3265 1730
rect 3285 1760 3325 1765
rect 3285 1730 3290 1760
rect 3320 1755 3325 1760
rect 3525 1760 3565 1765
rect 3525 1755 3530 1760
rect 3320 1735 3530 1755
rect 3320 1730 3325 1735
rect 3285 1725 3325 1730
rect 3525 1730 3530 1735
rect 3560 1755 3565 1760
rect 3765 1760 3805 1765
rect 3765 1755 3770 1760
rect 3560 1735 3770 1755
rect 3560 1730 3565 1735
rect 3525 1725 3565 1730
rect 3765 1730 3770 1735
rect 3800 1730 3805 1760
rect 3765 1725 3805 1730
rect 4205 1760 4245 1765
rect 4205 1730 4210 1760
rect 4240 1755 4245 1760
rect 4445 1760 4485 1765
rect 4445 1755 4450 1760
rect 4240 1735 4450 1755
rect 4240 1730 4245 1735
rect 4205 1725 4245 1730
rect 4445 1730 4450 1735
rect 4480 1755 4485 1760
rect 4685 1760 4725 1765
rect 4685 1755 4690 1760
rect 4480 1735 4690 1755
rect 4480 1730 4485 1735
rect 4445 1725 4485 1730
rect 4685 1730 4690 1735
rect 4720 1730 4725 1760
rect 4685 1725 4725 1730
rect 4745 1760 4785 1765
rect 4745 1730 4750 1760
rect 4780 1755 4785 1760
rect 5270 1760 5310 1765
rect 11237 1760 11240 1765
rect 5270 1755 5275 1760
rect 4780 1735 5275 1755
rect 4780 1730 4785 1735
rect 4745 1725 4785 1730
rect 5270 1730 5275 1735
rect 5305 1755 5310 1760
rect 5305 1735 6100 1755
rect 10805 1740 11240 1760
rect 11237 1735 11240 1740
rect 11266 1760 11269 1765
rect 11457 1765 11489 1770
rect 11457 1760 11460 1765
rect 11266 1740 11460 1760
rect 11266 1735 11269 1740
rect 5305 1730 5310 1735
rect 11237 1730 11269 1735
rect 11457 1735 11460 1740
rect 11486 1760 11489 1765
rect 11601 1765 11633 1770
rect 11601 1760 11604 1765
rect 11486 1740 11604 1760
rect 11486 1735 11489 1740
rect 11457 1730 11489 1735
rect 11601 1735 11604 1740
rect 11630 1760 11633 1765
rect 11867 1765 11899 1770
rect 11867 1760 11870 1765
rect 11630 1740 11870 1760
rect 11630 1735 11633 1740
rect 11601 1730 11633 1735
rect 11867 1735 11870 1740
rect 11896 1760 11899 1765
rect 12277 1765 12309 1770
rect 12277 1760 12280 1765
rect 11896 1740 12280 1760
rect 11896 1735 11899 1740
rect 11867 1730 11899 1735
rect 12277 1735 12280 1740
rect 12306 1760 12309 1765
rect 12497 1765 12529 1770
rect 12497 1760 12500 1765
rect 12306 1740 12500 1760
rect 12306 1735 12309 1740
rect 12277 1730 12309 1735
rect 12497 1735 12500 1740
rect 12526 1760 12529 1765
rect 12641 1765 12673 1770
rect 12641 1760 12644 1765
rect 12526 1740 12644 1760
rect 12526 1735 12529 1740
rect 12497 1730 12529 1735
rect 12641 1735 12644 1740
rect 12670 1735 12673 1765
rect 12641 1730 12673 1735
rect 5270 1725 5310 1730
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 1685 -70 1690
rect -45 1720 -5 1725
rect -45 1690 -40 1720
rect -10 1690 -5 1720
rect 3165 1715 3205 1720
rect -45 1685 -5 1690
rect 1262 1710 1302 1715
rect 1262 1680 1270 1710
rect 1297 1705 1302 1710
rect 2800 1710 2840 1715
rect 2800 1705 2805 1710
rect 1297 1685 2805 1705
rect 1297 1680 1302 1685
rect 1262 1675 1302 1680
rect 2800 1680 2805 1685
rect 2835 1680 2840 1710
rect 3165 1685 3170 1715
rect 3200 1710 3205 1715
rect 3405 1715 3445 1720
rect 3405 1710 3410 1715
rect 3200 1690 3410 1710
rect 3200 1685 3205 1690
rect 3165 1680 3205 1685
rect 3405 1685 3410 1690
rect 3440 1710 3445 1715
rect 3645 1715 3685 1720
rect 3645 1710 3650 1715
rect 3440 1690 3650 1710
rect 3440 1685 3445 1690
rect 3405 1680 3445 1685
rect 3645 1685 3650 1690
rect 3680 1685 3685 1715
rect 3645 1680 3685 1685
rect 4325 1715 4365 1720
rect 4325 1685 4330 1715
rect 4360 1710 4365 1715
rect 4565 1715 4605 1720
rect 4565 1710 4570 1715
rect 4360 1690 4570 1710
rect 4360 1685 4365 1690
rect 4325 1680 4365 1685
rect 4565 1685 4570 1690
rect 4600 1710 4605 1715
rect 4805 1715 4845 1720
rect 4805 1710 4810 1715
rect 4600 1690 4810 1710
rect 4600 1685 4605 1690
rect 4565 1680 4605 1685
rect 4805 1685 4810 1690
rect 4840 1685 4845 1715
rect 4805 1680 4845 1685
rect 2800 1675 2840 1680
rect 2380 1665 2420 1670
rect 2380 1635 2385 1665
rect 2415 1660 2420 1665
rect 2620 1665 2660 1670
rect 2620 1660 2625 1665
rect 2415 1640 2625 1660
rect 2415 1635 2420 1640
rect 2380 1630 2420 1635
rect 2620 1635 2625 1640
rect 2655 1635 2660 1665
rect 2620 1630 2660 1635
rect 2330 1595 2370 1600
rect 2330 1565 2335 1595
rect 2365 1590 2370 1595
rect 3165 1595 3205 1600
rect 3165 1590 3170 1595
rect 2365 1570 3170 1590
rect 2365 1565 2370 1570
rect 2330 1560 2370 1565
rect 3165 1565 3170 1570
rect 3200 1565 3205 1595
rect 3165 1560 3205 1565
rect 4805 1595 4845 1600
rect 4805 1565 4810 1595
rect 4840 1590 4845 1595
rect 5410 1595 5450 1600
rect 5410 1590 5415 1595
rect 4840 1570 5415 1590
rect 4840 1565 4845 1570
rect 4805 1560 4845 1565
rect 5410 1565 5415 1570
rect 5445 1565 5450 1595
rect 5410 1560 5450 1565
rect 2835 1545 2875 1550
rect 2835 1515 2840 1545
rect 2870 1540 2875 1545
rect 3225 1545 3265 1550
rect 3225 1540 3230 1545
rect 2870 1520 3230 1540
rect 2870 1515 2875 1520
rect 2835 1510 2875 1515
rect 3225 1515 3230 1520
rect 3260 1540 3265 1545
rect 3345 1545 3385 1550
rect 3345 1540 3350 1545
rect 3260 1520 3350 1540
rect 3260 1515 3265 1520
rect 3225 1510 3265 1515
rect 3345 1515 3350 1520
rect 3380 1540 3385 1545
rect 3465 1545 3505 1550
rect 3465 1540 3470 1545
rect 3380 1520 3470 1540
rect 3380 1515 3385 1520
rect 3345 1510 3385 1515
rect 3465 1515 3470 1520
rect 3500 1540 3505 1545
rect 3585 1545 3625 1550
rect 3585 1540 3590 1545
rect 3500 1520 3590 1540
rect 3500 1515 3505 1520
rect 3465 1510 3505 1515
rect 3585 1515 3590 1520
rect 3620 1540 3625 1545
rect 3705 1545 3745 1550
rect 3705 1540 3710 1545
rect 3620 1520 3710 1540
rect 3620 1515 3625 1520
rect 3585 1510 3625 1515
rect 3705 1515 3710 1520
rect 3740 1515 3745 1545
rect 3705 1510 3745 1515
rect 4265 1545 4305 1550
rect 4265 1515 4270 1545
rect 4300 1540 4305 1545
rect 4385 1545 4425 1550
rect 4385 1540 4390 1545
rect 4300 1520 4390 1540
rect 4300 1515 4305 1520
rect 4265 1510 4305 1515
rect 4385 1515 4390 1520
rect 4420 1540 4425 1545
rect 4505 1545 4545 1550
rect 4505 1540 4510 1545
rect 4420 1520 4510 1540
rect 4420 1515 4425 1520
rect 4385 1510 4425 1515
rect 4505 1515 4510 1520
rect 4540 1540 4545 1545
rect 4625 1545 4665 1550
rect 4625 1540 4630 1545
rect 4540 1520 4630 1540
rect 4540 1515 4545 1520
rect 4505 1510 4545 1515
rect 4625 1515 4630 1520
rect 4660 1540 4665 1545
rect 4745 1545 4785 1550
rect 4745 1540 4750 1545
rect 4660 1520 4750 1540
rect 4660 1515 4665 1520
rect 4625 1510 4665 1515
rect 4745 1515 4750 1520
rect 4780 1540 4785 1545
rect 5135 1545 5175 1550
rect 5135 1540 5140 1545
rect 4780 1520 5140 1540
rect 4780 1515 4785 1520
rect 4745 1510 4785 1515
rect 5135 1515 5140 1520
rect 5170 1515 5175 1545
rect 11106 1545 11138 1550
rect 11106 1540 11109 1545
rect 10805 1520 11109 1540
rect 5135 1510 5175 1515
rect 11106 1515 11109 1520
rect 11135 1540 11138 1545
rect 11305 1545 11345 1550
rect 11305 1540 11310 1545
rect 11135 1520 11310 1540
rect 11135 1515 11138 1520
rect 11106 1510 11138 1515
rect 11305 1515 11310 1520
rect 11340 1540 11345 1545
rect 11525 1545 11565 1550
rect 11525 1540 11530 1545
rect 11340 1520 11530 1540
rect 11340 1515 11345 1520
rect 11305 1510 11345 1515
rect 11525 1515 11530 1520
rect 11560 1540 11565 1545
rect 11922 1545 11954 1550
rect 11922 1540 11925 1545
rect 11560 1520 11925 1540
rect 11560 1515 11565 1520
rect 11525 1510 11565 1515
rect 11922 1515 11925 1520
rect 11951 1540 11954 1545
rect 12146 1545 12178 1550
rect 12146 1540 12149 1545
rect 11951 1520 12149 1540
rect 11951 1515 11954 1520
rect 11922 1510 11954 1515
rect 12146 1515 12149 1520
rect 12175 1540 12178 1545
rect 12345 1545 12385 1550
rect 12345 1540 12350 1545
rect 12175 1520 12350 1540
rect 12175 1515 12178 1520
rect 12146 1510 12178 1515
rect 12345 1515 12350 1520
rect 12380 1540 12385 1545
rect 12565 1545 12605 1550
rect 12565 1540 12570 1545
rect 12380 1520 12570 1540
rect 12380 1515 12385 1520
rect 12345 1510 12385 1515
rect 12565 1515 12570 1520
rect 12600 1515 12605 1545
rect 12565 1510 12605 1515
rect 2925 1500 2965 1505
rect 2925 1470 2930 1500
rect 2960 1495 2965 1500
rect 3045 1500 3085 1505
rect 3045 1495 3050 1500
rect 2960 1475 3050 1495
rect 2960 1470 2965 1475
rect 2925 1465 2965 1470
rect 3045 1470 3050 1475
rect 3080 1495 3085 1500
rect 3165 1500 3205 1505
rect 3165 1495 3170 1500
rect 3080 1475 3170 1495
rect 3080 1470 3085 1475
rect 3045 1465 3085 1470
rect 3165 1470 3170 1475
rect 3200 1495 3205 1500
rect 3285 1500 3325 1505
rect 3285 1495 3290 1500
rect 3200 1475 3290 1495
rect 3200 1470 3205 1475
rect 3165 1465 3205 1470
rect 3285 1470 3290 1475
rect 3320 1495 3325 1500
rect 3525 1500 3565 1505
rect 3525 1495 3530 1500
rect 3320 1475 3530 1495
rect 3320 1470 3325 1475
rect 3285 1465 3325 1470
rect 3525 1470 3530 1475
rect 3560 1495 3565 1500
rect 3645 1500 3685 1505
rect 3645 1495 3650 1500
rect 3560 1475 3650 1495
rect 3560 1470 3565 1475
rect 3525 1465 3565 1470
rect 3645 1470 3650 1475
rect 3680 1495 3685 1500
rect 3765 1500 3805 1505
rect 3765 1495 3770 1500
rect 3680 1475 3770 1495
rect 3680 1470 3685 1475
rect 3645 1465 3685 1470
rect 3765 1470 3770 1475
rect 3800 1495 3805 1500
rect 4205 1500 4245 1505
rect 4205 1495 4210 1500
rect 3800 1475 4210 1495
rect 3800 1470 3805 1475
rect 3765 1465 3805 1470
rect 4205 1470 4210 1475
rect 4240 1495 4245 1500
rect 4325 1500 4365 1505
rect 4325 1495 4330 1500
rect 4240 1475 4330 1495
rect 4240 1470 4245 1475
rect 4205 1465 4245 1470
rect 4325 1470 4330 1475
rect 4360 1495 4365 1500
rect 4445 1500 4485 1505
rect 4445 1495 4450 1500
rect 4360 1475 4450 1495
rect 4360 1470 4365 1475
rect 4325 1465 4365 1470
rect 4445 1470 4450 1475
rect 4480 1495 4485 1500
rect 4685 1500 4725 1505
rect 4685 1495 4690 1500
rect 4480 1475 4690 1495
rect 4480 1470 4485 1475
rect 4445 1465 4485 1470
rect 4685 1470 4690 1475
rect 4720 1495 4725 1500
rect 4805 1500 4845 1505
rect 4805 1495 4810 1500
rect 4720 1475 4810 1495
rect 4720 1470 4725 1475
rect 4685 1465 4725 1470
rect 4805 1470 4810 1475
rect 4840 1495 4845 1500
rect 4925 1500 4965 1505
rect 4925 1495 4930 1500
rect 4840 1475 4930 1495
rect 4840 1470 4845 1475
rect 4805 1465 4845 1470
rect 4925 1470 4930 1475
rect 4960 1495 4965 1500
rect 5045 1500 5085 1505
rect 5045 1495 5050 1500
rect 4960 1475 5050 1495
rect 4960 1470 4965 1475
rect 4925 1465 4965 1470
rect 5045 1470 5050 1475
rect 5080 1495 5085 1500
rect 5550 1500 5590 1505
rect 5550 1495 5555 1500
rect 5080 1475 5555 1495
rect 5080 1470 5085 1475
rect 5045 1465 5085 1470
rect 5550 1470 5555 1475
rect 5585 1470 5590 1500
rect 5550 1465 5590 1470
rect 11145 1485 11185 1490
rect 11145 1455 11150 1485
rect 11180 1480 11185 1485
rect 11250 1485 11290 1490
rect 11250 1480 11255 1485
rect 11180 1460 11255 1480
rect 11180 1455 11185 1460
rect 11145 1450 11185 1455
rect 11250 1455 11255 1460
rect 11285 1480 11290 1485
rect 11360 1485 11400 1490
rect 11360 1480 11365 1485
rect 11285 1460 11365 1480
rect 11285 1455 11290 1460
rect 11250 1450 11290 1455
rect 11360 1455 11365 1460
rect 11395 1480 11400 1485
rect 11470 1485 11510 1490
rect 11470 1480 11475 1485
rect 11395 1460 11475 1480
rect 11395 1455 11400 1460
rect 11360 1450 11400 1455
rect 11470 1455 11475 1460
rect 11505 1480 11510 1485
rect 11580 1485 11620 1490
rect 11580 1480 11585 1485
rect 11505 1460 11585 1480
rect 11505 1455 11510 1460
rect 11470 1450 11510 1455
rect 11580 1455 11585 1460
rect 11615 1480 11620 1485
rect 12185 1485 12225 1490
rect 12185 1480 12190 1485
rect 11615 1460 12190 1480
rect 11615 1455 11620 1460
rect 11580 1450 11620 1455
rect 12185 1455 12190 1460
rect 12220 1480 12225 1485
rect 12290 1485 12330 1490
rect 12290 1480 12295 1485
rect 12220 1460 12295 1480
rect 12220 1455 12225 1460
rect 12185 1450 12225 1455
rect 12290 1455 12295 1460
rect 12325 1480 12330 1485
rect 12400 1485 12440 1490
rect 12400 1480 12405 1485
rect 12325 1460 12405 1480
rect 12325 1455 12330 1460
rect 12290 1450 12330 1455
rect 12400 1455 12405 1460
rect 12435 1480 12440 1485
rect 12510 1485 12550 1490
rect 12510 1480 12515 1485
rect 12435 1460 12515 1480
rect 12435 1455 12440 1460
rect 12400 1450 12440 1455
rect 12510 1455 12515 1460
rect 12545 1480 12550 1485
rect 12620 1485 12660 1490
rect 12620 1480 12625 1485
rect 12545 1460 12625 1480
rect 12545 1455 12550 1460
rect 12510 1450 12550 1455
rect 12620 1455 12625 1460
rect 12655 1455 12660 1485
rect 12620 1450 12660 1455
rect 11810 1435 11850 1440
rect 11810 1405 11815 1435
rect 11845 1405 11850 1435
rect 11810 1400 11850 1405
rect 11315 1385 11355 1390
rect 11315 1355 11320 1385
rect 11350 1380 11355 1385
rect 11880 1385 11920 1390
rect 11880 1380 11885 1385
rect 11350 1360 11885 1380
rect 11350 1355 11355 1360
rect 11315 1350 11355 1355
rect 11880 1355 11885 1360
rect 11915 1355 11920 1385
rect 11880 1350 11920 1355
rect 11425 1325 11465 1330
rect 11425 1295 11430 1325
rect 11460 1320 11465 1325
rect 11535 1325 11575 1330
rect 11535 1320 11540 1325
rect 11460 1300 11540 1320
rect 11460 1295 11465 1300
rect 11425 1290 11465 1295
rect 11535 1295 11540 1300
rect 11570 1320 11575 1325
rect 11645 1325 11685 1330
rect 11645 1320 11650 1325
rect 11570 1300 11650 1320
rect 11570 1295 11575 1300
rect 11535 1290 11575 1295
rect 11645 1295 11650 1300
rect 11680 1320 11685 1325
rect 11755 1325 11795 1330
rect 11755 1320 11760 1325
rect 11680 1300 11760 1320
rect 11680 1295 11685 1300
rect 11645 1290 11685 1295
rect 11755 1295 11760 1300
rect 11790 1320 11795 1325
rect 11865 1325 11905 1330
rect 11865 1320 11870 1325
rect 11790 1300 11870 1320
rect 11790 1295 11795 1300
rect 11755 1290 11795 1295
rect 11865 1295 11870 1300
rect 11900 1320 11905 1325
rect 11975 1325 12015 1330
rect 11975 1320 11980 1325
rect 11900 1300 11980 1320
rect 11900 1295 11905 1300
rect 11865 1290 11905 1295
rect 11975 1295 11980 1300
rect 12010 1320 12015 1325
rect 12085 1325 12125 1330
rect 12085 1320 12090 1325
rect 12010 1300 12090 1320
rect 12010 1295 12015 1300
rect 11975 1290 12015 1295
rect 12085 1295 12090 1300
rect 12120 1320 12125 1325
rect 12195 1325 12235 1330
rect 12195 1320 12200 1325
rect 12120 1300 12200 1320
rect 12120 1295 12125 1300
rect 12085 1290 12125 1295
rect 12195 1295 12200 1300
rect 12230 1320 12235 1325
rect 12305 1325 12345 1330
rect 12305 1320 12310 1325
rect 12230 1300 12310 1320
rect 12230 1295 12235 1300
rect 12195 1290 12235 1295
rect 12305 1295 12310 1300
rect 12340 1320 12345 1325
rect 12415 1325 12455 1330
rect 12415 1320 12420 1325
rect 12340 1300 12420 1320
rect 12340 1295 12345 1300
rect 12305 1290 12345 1295
rect 12415 1295 12420 1300
rect 12450 1320 12455 1325
rect 12525 1325 12565 1330
rect 12525 1320 12530 1325
rect 12450 1300 12530 1320
rect 12450 1295 12455 1300
rect 12415 1290 12455 1295
rect 12525 1295 12530 1300
rect 12560 1295 12565 1325
rect 12525 1290 12565 1295
rect 3375 1185 3415 1190
rect 3375 1155 3380 1185
rect 3410 1180 3415 1185
rect 3985 1185 4025 1190
rect 3985 1180 3990 1185
rect 3410 1160 3990 1180
rect 3410 1155 3415 1160
rect 3375 1150 3415 1155
rect 3985 1155 3990 1160
rect 4020 1180 4025 1185
rect 4595 1185 4635 1190
rect 4595 1180 4600 1185
rect 4020 1160 4600 1180
rect 4020 1155 4025 1160
rect 3985 1150 4025 1155
rect 4595 1155 4600 1160
rect 4630 1180 4635 1185
rect 5465 1185 5505 1190
rect 5465 1180 5470 1185
rect 4630 1160 5470 1180
rect 4630 1155 4635 1160
rect 4595 1150 4635 1155
rect 5465 1155 5470 1160
rect 5500 1155 5505 1185
rect 5465 1150 5505 1155
rect 2945 1125 2985 1130
rect 2945 1095 2950 1125
rect 2980 1120 2985 1125
rect 3025 1125 3065 1130
rect 3025 1120 3030 1125
rect 2980 1100 3030 1120
rect 2980 1095 2985 1100
rect 2945 1090 2985 1095
rect 3025 1095 3030 1100
rect 3060 1120 3065 1125
rect 3105 1125 3145 1130
rect 3105 1120 3110 1125
rect 3060 1100 3110 1120
rect 3060 1095 3065 1100
rect 3025 1090 3065 1095
rect 3105 1095 3110 1100
rect 3140 1120 3145 1125
rect 3185 1125 3225 1130
rect 3185 1120 3190 1125
rect 3140 1100 3190 1120
rect 3140 1095 3145 1100
rect 3105 1090 3145 1095
rect 3185 1095 3190 1100
rect 3220 1120 3225 1125
rect 3265 1125 3305 1130
rect 3265 1120 3270 1125
rect 3220 1100 3270 1120
rect 3220 1095 3225 1100
rect 3185 1090 3225 1095
rect 3265 1095 3270 1100
rect 3300 1120 3305 1125
rect 3345 1125 3385 1130
rect 3345 1120 3350 1125
rect 3300 1100 3350 1120
rect 3300 1095 3305 1100
rect 3265 1090 3305 1095
rect 3345 1095 3350 1100
rect 3380 1120 3385 1125
rect 3425 1125 3465 1130
rect 3425 1120 3430 1125
rect 3380 1100 3430 1120
rect 3380 1095 3385 1100
rect 3345 1090 3385 1095
rect 3425 1095 3430 1100
rect 3460 1120 3465 1125
rect 3505 1125 3545 1130
rect 3505 1120 3510 1125
rect 3460 1100 3510 1120
rect 3460 1095 3465 1100
rect 3425 1090 3465 1095
rect 3505 1095 3510 1100
rect 3540 1120 3545 1125
rect 3585 1125 3625 1130
rect 3585 1120 3590 1125
rect 3540 1100 3590 1120
rect 3540 1095 3545 1100
rect 3505 1090 3545 1095
rect 3585 1095 3590 1100
rect 3620 1120 3625 1125
rect 3665 1125 3705 1130
rect 3665 1120 3670 1125
rect 3620 1100 3670 1120
rect 3620 1095 3625 1100
rect 3585 1090 3625 1095
rect 3665 1095 3670 1100
rect 3700 1120 3705 1125
rect 3745 1125 3785 1130
rect 3745 1120 3750 1125
rect 3700 1100 3750 1120
rect 3700 1095 3705 1100
rect 3665 1090 3705 1095
rect 3745 1095 3750 1100
rect 3780 1120 3785 1125
rect 3825 1125 3865 1130
rect 3825 1120 3830 1125
rect 3780 1100 3830 1120
rect 3780 1095 3785 1100
rect 3745 1090 3785 1095
rect 3825 1095 3830 1100
rect 3860 1120 3865 1125
rect 3905 1125 3945 1130
rect 3905 1120 3910 1125
rect 3860 1100 3910 1120
rect 3860 1095 3865 1100
rect 3825 1090 3865 1095
rect 3905 1095 3910 1100
rect 3940 1095 3945 1125
rect 3905 1090 3945 1095
rect 3985 1125 4025 1130
rect 3985 1095 3990 1125
rect 4020 1120 4025 1125
rect 4065 1125 4105 1130
rect 4065 1120 4070 1125
rect 4020 1100 4070 1120
rect 4020 1095 4025 1100
rect 3985 1090 4025 1095
rect 4065 1095 4070 1100
rect 4100 1120 4105 1125
rect 4145 1125 4185 1130
rect 4145 1120 4150 1125
rect 4100 1100 4150 1120
rect 4100 1095 4105 1100
rect 4065 1090 4105 1095
rect 4145 1095 4150 1100
rect 4180 1120 4185 1125
rect 4225 1125 4265 1130
rect 4225 1120 4230 1125
rect 4180 1100 4230 1120
rect 4180 1095 4185 1100
rect 4145 1090 4185 1095
rect 4225 1095 4230 1100
rect 4260 1120 4265 1125
rect 4305 1125 4345 1130
rect 4305 1120 4310 1125
rect 4260 1100 4310 1120
rect 4260 1095 4265 1100
rect 4225 1090 4265 1095
rect 4305 1095 4310 1100
rect 4340 1120 4345 1125
rect 4385 1125 4425 1130
rect 4385 1120 4390 1125
rect 4340 1100 4390 1120
rect 4340 1095 4345 1100
rect 4305 1090 4345 1095
rect 4385 1095 4390 1100
rect 4420 1120 4425 1125
rect 4465 1125 4505 1130
rect 4465 1120 4470 1125
rect 4420 1100 4470 1120
rect 4420 1095 4425 1100
rect 4385 1090 4425 1095
rect 4465 1095 4470 1100
rect 4500 1120 4505 1125
rect 4545 1125 4585 1130
rect 4545 1120 4550 1125
rect 4500 1100 4550 1120
rect 4500 1095 4505 1100
rect 4465 1090 4505 1095
rect 4545 1095 4550 1100
rect 4580 1120 4585 1125
rect 4625 1125 4665 1130
rect 4625 1120 4630 1125
rect 4580 1100 4630 1120
rect 4580 1095 4585 1100
rect 4545 1090 4585 1095
rect 4625 1095 4630 1100
rect 4660 1120 4665 1125
rect 4705 1125 4745 1130
rect 4705 1120 4710 1125
rect 4660 1100 4710 1120
rect 4660 1095 4665 1100
rect 4625 1090 4665 1095
rect 4705 1095 4710 1100
rect 4740 1120 4745 1125
rect 4785 1125 4825 1130
rect 4785 1120 4790 1125
rect 4740 1100 4790 1120
rect 4740 1095 4745 1100
rect 4705 1090 4745 1095
rect 4785 1095 4790 1100
rect 4820 1120 4825 1125
rect 4865 1125 4905 1130
rect 4865 1120 4870 1125
rect 4820 1100 4870 1120
rect 4820 1095 4825 1100
rect 4785 1090 4825 1095
rect 4865 1095 4870 1100
rect 4900 1120 4905 1125
rect 4945 1125 4985 1130
rect 4945 1120 4950 1125
rect 4900 1100 4950 1120
rect 4900 1095 4905 1100
rect 4865 1090 4905 1095
rect 4945 1095 4950 1100
rect 4980 1095 4985 1125
rect 4945 1090 4985 1095
rect 2620 1040 2660 1045
rect 2620 1010 2625 1040
rect 2655 1035 2660 1040
rect 2905 1040 2945 1045
rect 2905 1035 2910 1040
rect 2655 1015 2910 1035
rect 2655 1010 2660 1015
rect 2620 1005 2660 1010
rect 2905 1010 2910 1015
rect 2940 1010 2945 1040
rect 2905 1005 2945 1010
rect 5110 1040 5150 1045
rect 5110 1010 5115 1040
rect 5145 1035 5150 1040
rect 5465 1040 5505 1045
rect 5465 1035 5470 1040
rect 5145 1015 5470 1035
rect 5145 1010 5150 1015
rect 5110 1005 5150 1010
rect 5465 1010 5470 1015
rect 5500 1010 5505 1040
rect 5465 1005 5505 1010
rect 11165 1005 11205 1010
rect 11165 975 11170 1005
rect 11200 1000 11205 1005
rect 11260 1005 11300 1010
rect 11260 1000 11265 1005
rect 11200 980 11265 1000
rect 11200 975 11205 980
rect 11165 970 11205 975
rect 11260 975 11265 980
rect 11295 1000 11300 1005
rect 11370 1005 11410 1010
rect 11370 1000 11375 1005
rect 11295 980 11375 1000
rect 11295 975 11300 980
rect 11260 970 11300 975
rect 11370 975 11375 980
rect 11405 1000 11410 1005
rect 11480 1005 11520 1010
rect 11480 1000 11485 1005
rect 11405 980 11485 1000
rect 11405 975 11410 980
rect 11370 970 11410 975
rect 11480 975 11485 980
rect 11515 1000 11520 1005
rect 11590 1005 11630 1010
rect 11590 1000 11595 1005
rect 11515 980 11595 1000
rect 11515 975 11520 980
rect 11480 970 11520 975
rect 11590 975 11595 980
rect 11625 1000 11630 1005
rect 11700 1005 11740 1010
rect 11700 1000 11705 1005
rect 11625 980 11705 1000
rect 11625 975 11630 980
rect 11590 970 11630 975
rect 11700 975 11705 980
rect 11735 1000 11740 1005
rect 11810 1005 11850 1010
rect 11810 1000 11815 1005
rect 11735 980 11815 1000
rect 11735 975 11740 980
rect 11700 970 11740 975
rect 11810 975 11815 980
rect 11845 1000 11850 1005
rect 11920 1005 11960 1010
rect 11920 1000 11925 1005
rect 11845 980 11925 1000
rect 11845 975 11850 980
rect 11810 970 11850 975
rect 11920 975 11925 980
rect 11955 1000 11960 1005
rect 12030 1005 12070 1010
rect 12030 1000 12035 1005
rect 11955 980 12035 1000
rect 11955 975 11960 980
rect 11920 970 11960 975
rect 12030 975 12035 980
rect 12065 1000 12070 1005
rect 12140 1005 12180 1010
rect 12140 1000 12145 1005
rect 12065 980 12145 1000
rect 12065 975 12070 980
rect 12030 970 12070 975
rect 12140 975 12145 980
rect 12175 1000 12180 1005
rect 12250 1005 12290 1010
rect 12250 1000 12255 1005
rect 12175 980 12255 1000
rect 12175 975 12180 980
rect 12140 970 12180 975
rect 12250 975 12255 980
rect 12285 1000 12290 1005
rect 12360 1005 12400 1010
rect 12360 1000 12365 1005
rect 12285 980 12365 1000
rect 12285 975 12290 980
rect 12250 970 12290 975
rect 12360 975 12365 980
rect 12395 1000 12400 1005
rect 12470 1005 12510 1010
rect 12470 1000 12475 1005
rect 12395 980 12475 1000
rect 12395 975 12400 980
rect 12360 970 12400 975
rect 12470 975 12475 980
rect 12505 1000 12510 1005
rect 12620 1005 12660 1010
rect 12620 1000 12625 1005
rect 12505 980 12625 1000
rect 12505 975 12510 980
rect 12470 970 12510 975
rect 12620 975 12625 980
rect 12655 975 12660 1005
rect 12620 970 12660 975
rect 2995 930 3035 935
rect 2995 900 3000 930
rect 3030 925 3035 930
rect 3175 930 3215 935
rect 3175 925 3180 930
rect 3030 905 3180 925
rect 3030 900 3035 905
rect 2995 895 3035 900
rect 3175 900 3180 905
rect 3210 925 3215 930
rect 3355 930 3395 935
rect 3355 925 3360 930
rect 3210 905 3360 925
rect 3210 900 3215 905
rect 3175 895 3215 900
rect 3355 900 3360 905
rect 3390 925 3395 930
rect 3535 930 3575 935
rect 3535 925 3540 930
rect 3390 905 3540 925
rect 3390 900 3395 905
rect 3355 895 3395 900
rect 3535 900 3540 905
rect 3570 925 3575 930
rect 3715 930 3755 935
rect 3715 925 3720 930
rect 3570 905 3720 925
rect 3570 900 3575 905
rect 3535 895 3575 900
rect 3715 900 3720 905
rect 3750 925 3755 930
rect 3895 930 3935 935
rect 3895 925 3900 930
rect 3750 905 3900 925
rect 3750 900 3755 905
rect 3715 895 3755 900
rect 3895 900 3900 905
rect 3930 925 3935 930
rect 4075 930 4115 935
rect 4075 925 4080 930
rect 3930 905 4080 925
rect 3930 900 3935 905
rect 3895 895 3935 900
rect 4075 900 4080 905
rect 4110 925 4115 930
rect 4255 930 4295 935
rect 4255 925 4260 930
rect 4110 905 4260 925
rect 4110 900 4115 905
rect 4075 895 4115 900
rect 4255 900 4260 905
rect 4290 925 4295 930
rect 4435 930 4475 935
rect 4435 925 4440 930
rect 4290 905 4440 925
rect 4290 900 4295 905
rect 4255 895 4295 900
rect 4435 900 4440 905
rect 4470 925 4475 930
rect 4615 930 4655 935
rect 4615 925 4620 930
rect 4470 905 4620 925
rect 4470 900 4475 905
rect 4435 895 4475 900
rect 4615 900 4620 905
rect 4650 925 4655 930
rect 4795 930 4835 935
rect 4795 925 4800 930
rect 4650 905 4800 925
rect 4650 900 4655 905
rect 4615 895 4655 900
rect 4795 900 4800 905
rect 4830 925 4835 930
rect 4975 930 5015 935
rect 4975 925 4980 930
rect 4830 905 4980 925
rect 4830 900 4835 905
rect 4795 895 4835 900
rect 4975 900 4980 905
rect 5010 925 5015 930
rect 5465 930 5505 935
rect 5465 925 5470 930
rect 5010 905 5470 925
rect 5010 900 5015 905
rect 4975 895 5015 900
rect 5465 900 5470 905
rect 5500 900 5505 930
rect 5465 895 5505 900
rect 2520 760 2560 765
rect 2520 730 2525 760
rect 2555 755 2560 760
rect 3130 760 3170 765
rect 3130 755 3135 760
rect 2555 735 3135 755
rect 2555 730 2560 735
rect 2520 725 2560 730
rect 3130 730 3135 735
rect 3165 730 3170 760
rect 3130 725 3170 730
rect 3625 760 3665 765
rect 3625 730 3630 760
rect 3660 755 3665 760
rect 3985 760 4025 765
rect 3985 755 3990 760
rect 3660 735 3990 755
rect 3660 730 3665 735
rect 3625 725 3665 730
rect 3985 730 3990 735
rect 4020 755 4025 760
rect 4345 760 4385 765
rect 4345 755 4350 760
rect 4020 735 4350 755
rect 4020 730 4025 735
rect 3985 725 4025 730
rect 4345 730 4350 735
rect 4380 730 4385 760
rect 4345 725 4385 730
rect 4525 760 4565 765
rect 4525 730 4530 760
rect 4560 755 4565 760
rect 4705 760 4745 765
rect 4705 755 4710 760
rect 4560 735 4710 755
rect 4560 730 4565 735
rect 4525 725 4565 730
rect 4705 730 4710 735
rect 4740 755 4745 760
rect 4885 760 4925 765
rect 4885 755 4890 760
rect 4740 735 4890 755
rect 4740 730 4745 735
rect 4705 725 4745 730
rect 4885 730 4890 735
rect 4920 730 4925 760
rect 4885 725 4925 730
rect 3445 705 3485 710
rect 3445 675 3450 705
rect 3480 700 3485 705
rect 3805 705 3845 710
rect 3805 700 3810 705
rect 3480 680 3810 700
rect 3480 675 3485 680
rect 3445 670 3485 675
rect 3805 675 3810 680
rect 3840 700 3845 705
rect 4165 705 4205 710
rect 4165 700 4170 705
rect 3840 680 4170 700
rect 3840 675 3845 680
rect 3805 670 3845 675
rect 4165 675 4170 680
rect 4200 675 4205 705
rect 4165 670 4205 675
rect -195 575 -155 580
rect -195 545 -190 575
rect -160 545 -155 575
rect -195 540 -155 545
<< via2 >>
rect -190 4960 -160 4990
rect 5555 4960 5585 4990
rect -105 3495 -75 3525
rect 4445 3465 4475 3495
rect 945 3415 975 3445
rect 1645 3415 1675 3445
rect 5145 3415 5175 3445
rect 5555 3415 5585 3445
rect 2695 3360 2725 3390
rect 3395 3305 3425 3335
rect -105 3110 -75 3140
rect -105 2970 -75 3000
rect -105 2880 -75 2910
rect 5555 2780 5585 2810
rect 5555 2065 5585 2095
rect -105 1690 -75 1720
rect 5555 1470 5585 1500
rect 5470 1155 5500 1185
rect 5470 1010 5500 1040
rect 5470 900 5500 930
rect -190 545 -160 575
<< metal3 >>
rect -200 4995 -150 5000
rect -200 4955 -195 4995
rect -155 4955 -150 4995
rect -200 4950 -150 4955
rect 5545 4995 5595 5000
rect 5545 4955 5550 4995
rect 5590 4955 5595 4995
rect 5545 4950 5595 4955
rect -195 585 -155 4950
rect -115 4910 -65 4915
rect -115 4870 -110 4910
rect -70 4870 -65 4910
rect -115 4865 -65 4870
rect 5460 4910 5510 4915
rect 5460 4870 5465 4910
rect 5505 4870 5510 4910
rect 5460 4865 5510 4870
rect -110 3525 -70 4865
rect 145 4770 375 4855
rect 495 4770 725 4855
rect 845 4770 1075 4855
rect 1195 4770 1425 4855
rect 1545 4770 1775 4855
rect 145 4720 1775 4770
rect 145 4625 375 4720
rect 495 4625 725 4720
rect 845 4625 1075 4720
rect 1195 4625 1425 4720
rect 1545 4625 1775 4720
rect 1895 4770 2125 4855
rect 2245 4770 2475 4855
rect 2595 4770 2825 4855
rect 2945 4770 3175 4855
rect 3295 4770 3525 4855
rect 1895 4720 3525 4770
rect 1895 4625 2125 4720
rect 2245 4625 2475 4720
rect 2595 4625 2825 4720
rect 2945 4625 3175 4720
rect 3295 4625 3525 4720
rect 3645 4770 3875 4855
rect 3995 4770 4225 4855
rect 4345 4770 4575 4855
rect 4695 4770 4925 4855
rect 5045 4770 5275 4855
rect 3645 4720 5275 4770
rect 3645 4625 3875 4720
rect 3995 4625 4225 4720
rect 4345 4625 4575 4720
rect 4695 4625 4925 4720
rect 5045 4625 5275 4720
rect 935 4505 985 4625
rect 2685 4505 2735 4625
rect 4435 4505 4485 4625
rect 145 4420 375 4505
rect 495 4420 725 4505
rect 845 4420 1075 4505
rect 1195 4420 1425 4505
rect 1545 4420 1775 4505
rect 145 4370 1775 4420
rect 145 4275 375 4370
rect 495 4275 725 4370
rect 845 4275 1075 4370
rect 1195 4275 1425 4370
rect 1545 4275 1775 4370
rect 1895 4420 2125 4505
rect 2245 4420 2475 4505
rect 2595 4420 2825 4505
rect 2945 4420 3175 4505
rect 3295 4420 3525 4505
rect 1895 4370 3525 4420
rect 1895 4275 2125 4370
rect 2245 4275 2475 4370
rect 2595 4275 2825 4370
rect 2945 4275 3175 4370
rect 3295 4275 3525 4370
rect 3645 4420 3875 4505
rect 3995 4420 4225 4505
rect 4345 4420 4575 4505
rect 4695 4420 4925 4505
rect 5045 4420 5275 4505
rect 3645 4370 5275 4420
rect 3645 4275 3875 4370
rect 3995 4275 4225 4370
rect 4345 4275 4575 4370
rect 4695 4275 4925 4370
rect 5045 4275 5275 4370
rect 935 4155 985 4275
rect 2685 4155 2735 4275
rect 4435 4155 4485 4275
rect 145 4070 375 4155
rect 495 4070 725 4155
rect 845 4070 1075 4155
rect 1195 4070 1425 4155
rect 1545 4070 1775 4155
rect 145 4020 1775 4070
rect 145 3925 375 4020
rect 495 3925 725 4020
rect 845 3925 1075 4020
rect 1195 3925 1425 4020
rect 1545 3925 1775 4020
rect 1895 4070 2125 4155
rect 2245 4070 2475 4155
rect 2595 4070 2825 4155
rect 2945 4070 3175 4155
rect 3295 4070 3525 4155
rect 1895 4020 3525 4070
rect 1895 3925 2125 4020
rect 2245 3925 2475 4020
rect 2595 3925 2825 4020
rect 2945 3925 3175 4020
rect 3295 3925 3525 4020
rect 3645 4070 3875 4155
rect 3995 4070 4225 4155
rect 4345 4070 4575 4155
rect 4695 4070 4925 4155
rect 5045 4070 5275 4155
rect 3645 4020 5275 4070
rect 3645 3925 3875 4020
rect 3995 3925 4225 4020
rect 4345 3925 4575 4020
rect 4695 3925 4925 4020
rect 5045 3925 5275 4020
rect 935 3805 985 3925
rect 2685 3805 2735 3925
rect 4435 3805 4485 3925
rect 145 3720 375 3805
rect 495 3720 725 3805
rect 845 3720 1075 3805
rect 1195 3720 1425 3805
rect 1545 3720 1775 3805
rect 145 3670 1775 3720
rect 145 3575 375 3670
rect 495 3575 725 3670
rect 845 3575 1075 3670
rect 1195 3575 1425 3670
rect 1545 3575 1775 3670
rect 1895 3720 2125 3805
rect 2245 3720 2475 3805
rect 2595 3720 2825 3805
rect 2945 3720 3175 3805
rect 3295 3720 3525 3805
rect 1895 3670 3525 3720
rect 1895 3575 2125 3670
rect 2245 3575 2475 3670
rect 2595 3575 2825 3670
rect 2945 3575 3175 3670
rect 3295 3575 3525 3670
rect 3645 3720 3875 3805
rect 3995 3720 4225 3805
rect 4345 3720 4575 3805
rect 4695 3720 4925 3805
rect 5045 3720 5275 3805
rect 3645 3670 5275 3720
rect 3645 3575 3875 3670
rect 3995 3575 4225 3670
rect 4345 3575 4575 3670
rect 4695 3575 4925 3670
rect 5045 3575 5275 3670
rect -110 3495 -105 3525
rect -75 3495 -70 3525
rect -110 3140 -70 3495
rect 940 3445 980 3575
rect 940 3415 945 3445
rect 975 3415 980 3445
rect 940 3410 980 3415
rect 1635 3450 1685 3455
rect 1635 3410 1640 3450
rect 1680 3410 1685 3450
rect 1635 3405 1685 3410
rect 2690 3390 2730 3575
rect 4440 3495 4480 3575
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect 5135 3450 5185 3455
rect 5135 3410 5140 3450
rect 5180 3410 5185 3450
rect 5135 3405 5185 3410
rect 2690 3360 2695 3390
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 3385 3340 3435 3345
rect 3385 3300 3390 3340
rect 3430 3300 3435 3340
rect 3385 3295 3435 3300
rect -110 3110 -105 3140
rect -75 3110 -70 3140
rect -110 3000 -70 3110
rect -110 2970 -105 3000
rect -75 2970 -70 3000
rect -110 2910 -70 2970
rect -110 2880 -105 2910
rect -75 2880 -70 2910
rect -110 1720 -70 2880
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 665 -70 1690
rect 5465 1185 5505 4865
rect 5465 1155 5470 1185
rect 5500 1155 5505 1185
rect 5465 1040 5505 1155
rect 5465 1010 5470 1040
rect 5500 1010 5505 1040
rect 5465 930 5505 1010
rect 5465 900 5470 930
rect 5500 900 5505 930
rect 5465 665 5505 900
rect 5550 3445 5590 4950
rect 5550 3415 5555 3445
rect 5585 3415 5590 3445
rect 5550 2810 5590 3415
rect 5550 2780 5555 2810
rect 5585 2780 5590 2810
rect 5550 2095 5590 2780
rect 5550 2065 5555 2095
rect 5585 2065 5590 2095
rect 5550 1500 5590 2065
rect 5550 1470 5555 1500
rect 5585 1470 5590 1500
rect -115 660 -65 665
rect -115 620 -110 660
rect -70 620 -65 660
rect -115 615 -65 620
rect 5460 660 5510 665
rect 5460 620 5465 660
rect 5505 620 5510 660
rect 5460 615 5510 620
rect 5550 585 5590 1470
rect -200 580 -150 585
rect -200 540 -195 580
rect -155 540 -150 580
rect -200 535 -150 540
rect 5545 580 5595 585
rect 5545 540 5550 580
rect 5590 540 5595 580
rect 5545 535 5595 540
<< via3 >>
rect -195 4990 -155 4995
rect -195 4960 -190 4990
rect -190 4960 -160 4990
rect -160 4960 -155 4990
rect -195 4955 -155 4960
rect 5550 4990 5590 4995
rect 5550 4960 5555 4990
rect 5555 4960 5585 4990
rect 5585 4960 5590 4990
rect 5550 4955 5590 4960
rect -110 4870 -70 4910
rect 5465 4870 5505 4910
rect 1640 3445 1680 3450
rect 1640 3415 1645 3445
rect 1645 3415 1675 3445
rect 1675 3415 1680 3445
rect 1640 3410 1680 3415
rect 5140 3445 5180 3450
rect 5140 3415 5145 3445
rect 5145 3415 5175 3445
rect 5175 3415 5180 3445
rect 5140 3410 5180 3415
rect 3390 3335 3430 3340
rect 3390 3305 3395 3335
rect 3395 3305 3425 3335
rect 3425 3305 3430 3335
rect 3390 3300 3430 3305
rect -110 620 -70 660
rect 5465 620 5505 660
rect -195 575 -155 580
rect -195 545 -190 575
rect -190 545 -160 575
rect -160 545 -155 575
rect -195 540 -155 545
rect 5550 540 5590 580
<< mimcap >>
rect 160 4765 360 4840
rect 160 4725 240 4765
rect 280 4725 360 4765
rect 160 4640 360 4725
rect 510 4765 710 4840
rect 510 4725 590 4765
rect 630 4725 710 4765
rect 510 4640 710 4725
rect 860 4765 1060 4840
rect 860 4725 940 4765
rect 980 4725 1060 4765
rect 860 4640 1060 4725
rect 1210 4765 1410 4840
rect 1210 4725 1290 4765
rect 1330 4725 1410 4765
rect 1210 4640 1410 4725
rect 1560 4765 1760 4840
rect 1560 4725 1640 4765
rect 1680 4725 1760 4765
rect 1560 4640 1760 4725
rect 1910 4765 2110 4840
rect 1910 4725 1990 4765
rect 2030 4725 2110 4765
rect 1910 4640 2110 4725
rect 2260 4765 2460 4840
rect 2260 4725 2340 4765
rect 2380 4725 2460 4765
rect 2260 4640 2460 4725
rect 2610 4765 2810 4840
rect 2610 4725 2690 4765
rect 2730 4725 2810 4765
rect 2610 4640 2810 4725
rect 2960 4765 3160 4840
rect 2960 4725 3040 4765
rect 3080 4725 3160 4765
rect 2960 4640 3160 4725
rect 3310 4765 3510 4840
rect 3310 4725 3390 4765
rect 3430 4725 3510 4765
rect 3310 4640 3510 4725
rect 3660 4765 3860 4840
rect 3660 4725 3740 4765
rect 3780 4725 3860 4765
rect 3660 4640 3860 4725
rect 4010 4765 4210 4840
rect 4010 4725 4090 4765
rect 4130 4725 4210 4765
rect 4010 4640 4210 4725
rect 4360 4765 4560 4840
rect 4360 4725 4440 4765
rect 4480 4725 4560 4765
rect 4360 4640 4560 4725
rect 4710 4765 4910 4840
rect 4710 4725 4790 4765
rect 4830 4725 4910 4765
rect 4710 4640 4910 4725
rect 5060 4765 5260 4840
rect 5060 4725 5140 4765
rect 5180 4725 5260 4765
rect 5060 4640 5260 4725
rect 160 4415 360 4490
rect 160 4375 240 4415
rect 280 4375 360 4415
rect 160 4290 360 4375
rect 510 4415 710 4490
rect 510 4375 590 4415
rect 630 4375 710 4415
rect 510 4290 710 4375
rect 860 4415 1060 4490
rect 860 4375 940 4415
rect 980 4375 1060 4415
rect 860 4290 1060 4375
rect 1210 4415 1410 4490
rect 1210 4375 1290 4415
rect 1330 4375 1410 4415
rect 1210 4290 1410 4375
rect 1560 4415 1760 4490
rect 1560 4375 1640 4415
rect 1680 4375 1760 4415
rect 1560 4290 1760 4375
rect 1910 4415 2110 4490
rect 1910 4375 1990 4415
rect 2030 4375 2110 4415
rect 1910 4290 2110 4375
rect 2260 4415 2460 4490
rect 2260 4375 2340 4415
rect 2380 4375 2460 4415
rect 2260 4290 2460 4375
rect 2610 4415 2810 4490
rect 2610 4375 2690 4415
rect 2730 4375 2810 4415
rect 2610 4290 2810 4375
rect 2960 4415 3160 4490
rect 2960 4375 3040 4415
rect 3080 4375 3160 4415
rect 2960 4290 3160 4375
rect 3310 4415 3510 4490
rect 3310 4375 3390 4415
rect 3430 4375 3510 4415
rect 3310 4290 3510 4375
rect 3660 4415 3860 4490
rect 3660 4375 3740 4415
rect 3780 4375 3860 4415
rect 3660 4290 3860 4375
rect 4010 4415 4210 4490
rect 4010 4375 4090 4415
rect 4130 4375 4210 4415
rect 4010 4290 4210 4375
rect 4360 4415 4560 4490
rect 4360 4375 4440 4415
rect 4480 4375 4560 4415
rect 4360 4290 4560 4375
rect 4710 4415 4910 4490
rect 4710 4375 4790 4415
rect 4830 4375 4910 4415
rect 4710 4290 4910 4375
rect 5060 4415 5260 4490
rect 5060 4375 5140 4415
rect 5180 4375 5260 4415
rect 5060 4290 5260 4375
rect 160 4065 360 4140
rect 160 4025 240 4065
rect 280 4025 360 4065
rect 160 3940 360 4025
rect 510 4065 710 4140
rect 510 4025 590 4065
rect 630 4025 710 4065
rect 510 3940 710 4025
rect 860 4065 1060 4140
rect 860 4025 940 4065
rect 980 4025 1060 4065
rect 860 3940 1060 4025
rect 1210 4065 1410 4140
rect 1210 4025 1290 4065
rect 1330 4025 1410 4065
rect 1210 3940 1410 4025
rect 1560 4065 1760 4140
rect 1560 4025 1640 4065
rect 1680 4025 1760 4065
rect 1560 3940 1760 4025
rect 1910 4065 2110 4140
rect 1910 4025 1990 4065
rect 2030 4025 2110 4065
rect 1910 3940 2110 4025
rect 2260 4065 2460 4140
rect 2260 4025 2340 4065
rect 2380 4025 2460 4065
rect 2260 3940 2460 4025
rect 2610 4065 2810 4140
rect 2610 4025 2690 4065
rect 2730 4025 2810 4065
rect 2610 3940 2810 4025
rect 2960 4065 3160 4140
rect 2960 4025 3040 4065
rect 3080 4025 3160 4065
rect 2960 3940 3160 4025
rect 3310 4065 3510 4140
rect 3310 4025 3390 4065
rect 3430 4025 3510 4065
rect 3310 3940 3510 4025
rect 3660 4065 3860 4140
rect 3660 4025 3740 4065
rect 3780 4025 3860 4065
rect 3660 3940 3860 4025
rect 4010 4065 4210 4140
rect 4010 4025 4090 4065
rect 4130 4025 4210 4065
rect 4010 3940 4210 4025
rect 4360 4065 4560 4140
rect 4360 4025 4440 4065
rect 4480 4025 4560 4065
rect 4360 3940 4560 4025
rect 4710 4065 4910 4140
rect 4710 4025 4790 4065
rect 4830 4025 4910 4065
rect 4710 3940 4910 4025
rect 5060 4065 5260 4140
rect 5060 4025 5140 4065
rect 5180 4025 5260 4065
rect 5060 3940 5260 4025
rect 160 3715 360 3790
rect 160 3675 240 3715
rect 280 3675 360 3715
rect 160 3590 360 3675
rect 510 3715 710 3790
rect 510 3675 590 3715
rect 630 3675 710 3715
rect 510 3590 710 3675
rect 860 3715 1060 3790
rect 860 3675 940 3715
rect 980 3675 1060 3715
rect 860 3590 1060 3675
rect 1210 3715 1410 3790
rect 1210 3675 1290 3715
rect 1330 3675 1410 3715
rect 1210 3590 1410 3675
rect 1560 3715 1760 3790
rect 1560 3675 1640 3715
rect 1680 3675 1760 3715
rect 1560 3590 1760 3675
rect 1910 3715 2110 3790
rect 1910 3675 1990 3715
rect 2030 3675 2110 3715
rect 1910 3590 2110 3675
rect 2260 3715 2460 3790
rect 2260 3675 2340 3715
rect 2380 3675 2460 3715
rect 2260 3590 2460 3675
rect 2610 3715 2810 3790
rect 2610 3675 2690 3715
rect 2730 3675 2810 3715
rect 2610 3590 2810 3675
rect 2960 3715 3160 3790
rect 2960 3675 3040 3715
rect 3080 3675 3160 3715
rect 2960 3590 3160 3675
rect 3310 3715 3510 3790
rect 3310 3675 3390 3715
rect 3430 3675 3510 3715
rect 3310 3590 3510 3675
rect 3660 3715 3860 3790
rect 3660 3675 3740 3715
rect 3780 3675 3860 3715
rect 3660 3590 3860 3675
rect 4010 3715 4210 3790
rect 4010 3675 4090 3715
rect 4130 3675 4210 3715
rect 4010 3590 4210 3675
rect 4360 3715 4560 3790
rect 4360 3675 4440 3715
rect 4480 3675 4560 3715
rect 4360 3590 4560 3675
rect 4710 3715 4910 3790
rect 4710 3675 4790 3715
rect 4830 3675 4910 3715
rect 4710 3590 4910 3675
rect 5060 3715 5260 3790
rect 5060 3675 5140 3715
rect 5180 3675 5260 3715
rect 5060 3590 5260 3675
<< mimcapcontact >>
rect 240 4725 280 4765
rect 590 4725 630 4765
rect 940 4725 980 4765
rect 1290 4725 1330 4765
rect 1640 4725 1680 4765
rect 1990 4725 2030 4765
rect 2340 4725 2380 4765
rect 2690 4725 2730 4765
rect 3040 4725 3080 4765
rect 3390 4725 3430 4765
rect 3740 4725 3780 4765
rect 4090 4725 4130 4765
rect 4440 4725 4480 4765
rect 4790 4725 4830 4765
rect 5140 4725 5180 4765
rect 240 4375 280 4415
rect 590 4375 630 4415
rect 940 4375 980 4415
rect 1290 4375 1330 4415
rect 1640 4375 1680 4415
rect 1990 4375 2030 4415
rect 2340 4375 2380 4415
rect 2690 4375 2730 4415
rect 3040 4375 3080 4415
rect 3390 4375 3430 4415
rect 3740 4375 3780 4415
rect 4090 4375 4130 4415
rect 4440 4375 4480 4415
rect 4790 4375 4830 4415
rect 5140 4375 5180 4415
rect 240 4025 280 4065
rect 590 4025 630 4065
rect 940 4025 980 4065
rect 1290 4025 1330 4065
rect 1640 4025 1680 4065
rect 1990 4025 2030 4065
rect 2340 4025 2380 4065
rect 2690 4025 2730 4065
rect 3040 4025 3080 4065
rect 3390 4025 3430 4065
rect 3740 4025 3780 4065
rect 4090 4025 4130 4065
rect 4440 4025 4480 4065
rect 4790 4025 4830 4065
rect 5140 4025 5180 4065
rect 240 3675 280 3715
rect 590 3675 630 3715
rect 940 3675 980 3715
rect 1290 3675 1330 3715
rect 1640 3675 1680 3715
rect 1990 3675 2030 3715
rect 2340 3675 2380 3715
rect 2690 3675 2730 3715
rect 3040 3675 3080 3715
rect 3390 3675 3430 3715
rect 3740 3675 3780 3715
rect 4090 3675 4130 3715
rect 4440 3675 4480 3715
rect 4790 3675 4830 3715
rect 5140 3675 5180 3715
<< metal4 >>
rect -200 4995 5595 5000
rect -200 4955 -195 4995
rect -155 4955 5550 4995
rect 5590 4955 5595 4995
rect -200 4950 5595 4955
rect -115 4910 5510 4915
rect -115 4870 -110 4910
rect -70 4870 5465 4910
rect 5505 4870 5510 4910
rect -115 4865 5510 4870
rect 235 4765 1685 4770
rect 235 4725 240 4765
rect 280 4725 590 4765
rect 630 4725 940 4765
rect 980 4725 1290 4765
rect 1330 4725 1640 4765
rect 1680 4725 1685 4765
rect 235 4720 1685 4725
rect 1985 4765 3435 4770
rect 1985 4725 1990 4765
rect 2030 4725 2340 4765
rect 2380 4725 2690 4765
rect 2730 4725 3040 4765
rect 3080 4725 3390 4765
rect 3430 4725 3435 4765
rect 1985 4720 3435 4725
rect 3735 4765 5185 4770
rect 3735 4725 3740 4765
rect 3780 4725 4090 4765
rect 4130 4725 4440 4765
rect 4480 4725 4790 4765
rect 4830 4725 5140 4765
rect 5180 4725 5185 4765
rect 3735 4720 5185 4725
rect 935 4420 985 4720
rect 2685 4420 2735 4720
rect 4435 4420 4485 4720
rect 235 4415 1685 4420
rect 235 4375 240 4415
rect 280 4375 590 4415
rect 630 4375 940 4415
rect 980 4375 1290 4415
rect 1330 4375 1640 4415
rect 1680 4375 1685 4415
rect 235 4370 1685 4375
rect 1985 4415 3435 4420
rect 1985 4375 1990 4415
rect 2030 4375 2340 4415
rect 2380 4375 2690 4415
rect 2730 4375 3040 4415
rect 3080 4375 3390 4415
rect 3430 4375 3435 4415
rect 1985 4370 3435 4375
rect 3735 4415 5185 4420
rect 3735 4375 3740 4415
rect 3780 4375 4090 4415
rect 4130 4375 4440 4415
rect 4480 4375 4790 4415
rect 4830 4375 5140 4415
rect 5180 4375 5185 4415
rect 3735 4370 5185 4375
rect 935 4070 985 4370
rect 2685 4070 2735 4370
rect 4435 4070 4485 4370
rect 235 4065 1685 4070
rect 235 4025 240 4065
rect 280 4025 590 4065
rect 630 4025 940 4065
rect 980 4025 1290 4065
rect 1330 4025 1640 4065
rect 1680 4025 1685 4065
rect 235 4020 1685 4025
rect 1985 4065 3435 4070
rect 1985 4025 1990 4065
rect 2030 4025 2340 4065
rect 2380 4025 2690 4065
rect 2730 4025 3040 4065
rect 3080 4025 3390 4065
rect 3430 4025 3435 4065
rect 1985 4020 3435 4025
rect 3735 4065 5185 4070
rect 3735 4025 3740 4065
rect 3780 4025 4090 4065
rect 4130 4025 4440 4065
rect 4480 4025 4790 4065
rect 4830 4025 5140 4065
rect 5180 4025 5185 4065
rect 3735 4020 5185 4025
rect 935 3720 985 4020
rect 2685 3720 2735 4020
rect 4435 3720 4485 4020
rect 235 3715 1685 3720
rect 235 3675 240 3715
rect 280 3675 590 3715
rect 630 3675 940 3715
rect 980 3675 1290 3715
rect 1330 3675 1640 3715
rect 1680 3675 1685 3715
rect 235 3670 1685 3675
rect 1985 3715 3435 3720
rect 1985 3675 1990 3715
rect 2030 3675 2340 3715
rect 2380 3675 2690 3715
rect 2730 3675 3040 3715
rect 3080 3675 3390 3715
rect 3430 3675 3435 3715
rect 1985 3670 3435 3675
rect 3735 3715 5185 3720
rect 3735 3675 3740 3715
rect 3780 3675 4090 3715
rect 4130 3675 4440 3715
rect 4480 3675 4790 3715
rect 4830 3675 5140 3715
rect 5180 3675 5185 3715
rect 3735 3670 5185 3675
rect 1635 3450 1685 3670
rect 1635 3410 1640 3450
rect 1680 3410 1685 3450
rect 1635 3405 1685 3410
rect 3385 3340 3435 3670
rect 5135 3450 5185 3670
rect 5135 3410 5140 3450
rect 5180 3410 5185 3450
rect 5135 3405 5185 3410
rect 3385 3300 3390 3340
rect 3430 3300 3435 3340
rect 3385 3295 3435 3300
rect -115 660 5510 665
rect -115 620 -110 660
rect -70 620 5465 660
rect 5505 620 5510 660
rect -115 615 5510 620
rect -200 580 5595 585
rect -200 540 -195 580
rect -155 540 5550 580
rect 5590 540 5595 580
rect -200 535 5595 540
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 795 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1723858470
transform 1 0 795 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1723858470
transform 1 0 795 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1723858470
transform 1 0 115 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1723858470
transform 1 0 115 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1723858470
transform 1 0 115 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1723858470
transform 1 0 1475 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1723858470
transform 1 0 1475 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1723858470
transform 1 0 1475 0 1 1360
box 0 0 670 670
<< labels >>
flabel metal2 2950 1735 2950 1735 5 FreeSans 400 0 0 -80 Vin-
flabel metal2 2955 1590 2955 1590 1 FreeSans 400 0 0 80 Vin+
flabel metal2 2945 1845 2945 1845 5 FreeSans 400 0 0 -40 V_mir1
flabel metal2 3745 1530 3745 1530 3 FreeSans 400 0 40 0 V_p1
flabel metal1 2650 1155 2650 1155 3 FreeSans 400 0 200 0 START_UP
flabel metal2 3785 1785 3785 1785 5 FreeSans 400 0 0 -40 1st_Vout1
flabel metal2 455 3440 455 3440 1 FreeSans 400 0 0 40 cap_res1
flabel metal3 2730 3375 2730 3375 3 FreeSans 400 0 40 0 cap_res2
flabel metal1 2550 845 2550 845 3 FreeSans 400 0 40 0 NFET_GATE_10uA
flabel metal2 5120 1590 5120 1590 1 FreeSans 400 0 0 80 V_CUR_REF_REG
flabel metal2 4225 1785 4225 1785 5 FreeSans 400 0 0 -40 1st_Vout2
flabel metal2 5065 1845 5065 1845 5 FreeSans 400 0 0 -40 V_mir2
flabel metal2 4265 1530 4265 1530 7 FreeSans 400 0 -40 0 V_p2
flabel metal1 3275 350 3275 350 7 FreeSans 400 0 -400 0 CMFB_NFET_CUR_BIAS
port 8 w
flabel metal1 3825 295 3825 295 5 FreeSans 400 0 0 -200 VB2_CUR_BIAS
port 5 s
flabel metal1 4015 350 4015 350 3 FreeSans 400 0 200 0 ERR_AMP_CUR_BIAS
port 7 e
flabel metal1 4725 295 4725 295 5 FreeSans 400 0 0 -200 VB3_CUR_BIAS
port 6 s
flabel metal1 4985 1110 4985 1110 3 FreeSans 400 0 200 0 START_UP_NFET1
flabel metal2 4115 3135 4115 3135 1 FreeSans 400 0 0 40 PFET_GATE_10uA
flabel metal2 6080 3075 6080 3075 1 FreeSans 400 0 0 200 VB1_CUR_BIAS
port 1 n
flabel metal2 6100 3020 6100 3020 3 FreeSans 400 0 200 0 TAIL_CUR_MIR_BIAS
port 9 e
flabel metal2 6080 2955 6080 2955 5 FreeSans 400 0 0 -200 CMFB_PFET_CUR_BIAS
port 10 s
flabel metal2 6100 1745 6100 1745 3 FreeSans 400 0 200 0 ERR_AMP_REF
port 3 e
flabel metal3 5590 4400 5590 4400 3 FreeSans 800 0 80 0 VDDA
port 4 e
flabel metal3 5505 4175 5505 4175 3 FreeSans 800 0 80 0 GNDA
port 2 e
flabel metal1 2180 1010 2180 1010 3 FreeSans 400 0 40 0 Vbe2
flabel poly 4635 2375 4635 2375 5 FreeSans 400 0 0 -40 V_TOP
<< end >>
