* NGSPICE file created from low_volt_BGR_11.ext - technology: sky130A

** .subckt sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 Emitter Collector Base m=1
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
.ends

** .subckt low_volt_BGR_11 VDDA V_out GNDA
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
+ GNDA GNDA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
+ GNDA GNDA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6 Vin- GNDA GNDA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
+ GNDA GNDA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
+ GNDA GNDA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
+ GNDA GNDA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
+ GNDA GNDA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
X0 GNDA a_4938_4530# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X1 VDDA V_TOP Vin- VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X2 VDDA V_TOP V_out VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X3 V_mirror V_mirror VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X4 GNDA a_4938_4770# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X5 VDDA V_TOP Vin- VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X6 1st_Vout V_mirror VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X7 V_out VDDA VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=0.6
X8 GNDA start_up start_up GNDA sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=10
X9 Vin+ V_TOP VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X10 Vin- start_up V_TOP VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X11 VDDA V_TOP start_up VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X12 Vin- V_TOP VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X13 GNDA GNDA V_mirror GNDA sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.6
X14 V_TOP V_TOP GNDA GNDA sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=1.6 ps=8.8 w=4 l=4
X15 VDDA V_mirror V_mirror VDDA sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X16 V_mirror Vin- V_p GNDA sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.6
X17 VDDA VDDA V_TOP VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.6
X18 1st_Vout Vin+ V_p GNDA sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.6
X19 V_TOP 1st_Vout VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X20 Vin+ a_4938_3210# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X21 VDDA V_TOP Vin+ VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X22 1st_Vout V_mirror VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X23 V_p Vin- V_mirror GNDA sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.6
X24 V_out a_4938_2970# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X25 VDDA VDDA V_out VDDA sky130_fd_pr__pfet_01v8 ad=1.6 pd=8.8 as=0.8 ps=4.4 w=4 l=0.6
X26 VDDA 1st_Vout V_TOP VDDA sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X27 a_3410_3330# a_4938_3210# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X28 V_out V_TOP VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X29 VDDA V_mirror V_mirror VDDA sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X30 Vin- V_TOP VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X31 a_3410_3450# a_4938_3810# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X32 a_3410_3450# a_4938_3090# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X33 Vin- a_4938_3090# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X34 VDDA V_TOP V_out VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X35 VDDA V_TOP Vin+ VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X36 a_3410_3330# a_4938_3930# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X37 a_3410_3570# a_4938_2970# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X38 V_mirror Vin- V_p GNDA sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.6
X39 a_3410_3570# a_4938_3690# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X40 a_3410_4410# a_4938_3690# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X41 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter Vin+ GNDA sky130_fd_pr__res_xhigh_po_0p35 l=3.5
X42 V_p Vin+ 1st_Vout GNDA sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.6
X43 GNDA V_p V_p GNDA sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=1.6 ps=8.8 w=4 l=4
X44 V_mirror V_mirror VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X45 V_p Vin- V_mirror GNDA sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.6
X46 a_3410_4410# a_4938_4530# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X47 a_3410_4170# a_4938_3930# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X48 V_TOP 1st_Vout VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X49 V_p Vin+ 1st_Vout GNDA sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.6
X50 a_3410_4290# a_4938_4650# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X51 VDDA V_mirror 1st_Vout VDDA sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X52 V_mirror GNDA GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.6
X53 Vin+ V_TOP VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X54 a_3410_4290# a_4938_3810# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X55 VDDA 1st_Vout V_TOP VDDA sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X56 1st_Vout Vin+ V_p GNDA sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.6
X57 GNDA a_4938_4650# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X58 V_out V_TOP VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.6
X59 VDDA V_mirror 1st_Vout VDDA sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.6
X60 a_3410_4170# a_4938_4770# GNDA sky130_fd_pr__res_xhigh_po_0p35 l=5.6
X61 V_TOP VDDA VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.6
.ends

