* PEX produced on Thu Feb 20 03:15:05 PM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from VCO_FD.ext - technology: sky130A

.subckt VCO_FD VDDA GNDA V_CONT V_OUT120
X0 a_2046_966.t2 a_110_1544.t3 VDDA.t83 VDDA.t82 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=1.5
X1 GNDA.t105 div120_0.div5_0.E.t2 div120_0.div5_0.I.t2 GNDA.t104 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X2 div120_0.div3_2_0.D.t0 div120_0.div3_2_0.C.t4 GNDA.t67 GNDA.t66 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X3 div120_0.div2_3_1.CLK.t1 V_OSC.t2 VDDA.t44 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X4 div120_0.div5_0.G.t0 V_OUT120.t2 div120_0.div5_0.F.t0 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X5 div120_0.div3_2_0.H.t2 div120_0.div3_2_0.CLK.t3 GNDA.t89 GNDA.t88 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X6 div120_0.div24.t1 div120_0.div3_2_0.I.t2 VDDA.t50 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X7 a_2046_228.t0 V_CONT.t0 GNDA.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X8 div120_0.div3_2_0.C.t3 div120_0.div3_2_0.A.t2 VDDA.t75 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X9 GNDA.t57 V_OSC.t3 div120_0.div2_3_1.CLK.t2 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X10 div120_0.div2_3_2.CLK.t1 div120_0.div2.t2 VDDA.t39 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X11 a_2046_228.t2 VDDA.t94 GNDA.t103 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.15
X12 a_1492_228.t1 V_CONT.t1 GNDA.t8 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X13 V_OUT120.t0 div120_0.div5_0.M.t4 GNDA.t42 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X14 div120_0.div5_0.H.t0 div120_0.div24.t3 div120_0.div5_0.G.t2 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X15 VDDA.t18 div120_0.div5_0.Q2_b.t2 div120_0.div5_0.G.t1 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X16 a_938_228.t0 V_CONT.t2 GNDA.t29 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X17 div120_0.div5_0.Q2_b.t1 div120_0.div5_0.J.t4 GNDA.t114 GNDA.t113 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X18 div120_0.div2_3_2.C.t3 div120_0.div2_3_2.CLK.t3 GNDA.t3 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X19 VDDA.t34 div120_0.div5_0.A.t3 div120_0.div5_0.B.t0 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X20 div120_0.div3_2_0.C.t2 div120_0.div3_2_0.CLK.t4 GNDA.t87 GNDA.t86 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X21 a_1492_228.t2 VDDA.t95 GNDA.t102 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.15
X22 div120_0.div2_3_2.B.t0 div120_0.div4.t2 GNDA.t91 GNDA.t90 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X23 div120_0.div5_0.E.t1 div120_0.div24.t4 VDDA.t87 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X24 a_938_228.t2 VDDA.t96 GNDA.t101 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.15
X25 GNDA.t23 div120_0.div2_3_0.CLK.t3 div120_0.div2_3_0.C.t2 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X26 div120_0.div5_0.L.t0 V_OUT120.t3 GNDA.t73 GNDA.t72 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X27 GNDA.t64 div120_0.div2_3_1.CLK.t3 div120_0.div2_3_1.C.t3 GNDA.t63 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X28 VDDA.t81 a_110_1544.t1 a_110_1544.t2 VDDA.t80 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=1.5
X29 div120_0.div5_0.M.t3 div120_0.div5_0.Q2_b.t3 GNDA.t112 GNDA.t111 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X30 div120_0.div5_0.J.t3 div120_0.div24.t5 GNDA.t38 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X31 GNDA.t95 div120_0.div3_2_0.I.t3 div120_0.div3_2_0.G.t1 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X32 a_2046_966.t1 GNDA.t118 VDDA.t48 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.15
X33 div120_0.div4.t0 div120_0.div2_3_2.C.t4 GNDA.t44 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X34 div120_0.div5_0.E.t0 div120_0.div5_0.D.t4 GNDA.t40 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X35 div120_0.div24.t2 div120_0.div3_2_0.I.t4 GNDA.t69 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X36 GNDA.t25 div120_0.div2_3_0.CLK.t4 div120_0.div2_3_0.C.t1 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X37 div120_0.div5_0.A.t1 div120_0.div5_0.Q2_b.t4 VDDA.t26 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X38 GNDA.t62 div120_0.div2_3_1.CLK.t4 div120_0.div2_3_1.C.t2 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X39 VDDA.t93 div120_0.div4.t3 div120_0.div2_3_0.CLK.t1 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X40 div120_0.div3_2_0.A.t0 div120_0.div3_2_0.CLK.t5 div120_0.div3_2_0.B.t0 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X41 div120_0.div2_3_2.A.t1 div120_0.div2_3_2.CLK.t4 div120_0.div2_3_2.B.t1 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X42 div120_0.div3_2_0.F.t0 div120_0.div3_2_0.CLK.t6 div120_0.div3_2_0.E.t0 GNDA.t84 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X43 div120_0.div3_2_0.I.t0 div120_0.div3_2_0.CLK.t7 VDDA.t71 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X44 div120_0.div5_0.M.t1 div120_0.div5_0.K.t2 VDDA.t30 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X45 VDDA.t32 div120_0.div8.t2 div120_0.div3_2_0.CLK.t2 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X46 div120_0.div5_0.C.t0 div120_0.div5_0.A.t4 GNDA.t48 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X47 a_938_966.t2 GNDA.t119 VDDA.t28 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.15
X48 div120_0.div5_0.D.t3 div120_0.div24.t6 GNDA.t27 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X49 div120_0.div3_2_0.E.t2 div120_0.div3_2_0.I.t5 VDDA.t7 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X50 a_2046_966.t0 V_OSC.t4 a_1460_718.t1 VDDA.t42 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.16
X51 div120_0.div5_0.I.t0 V_OUT120.t4 GNDA.t71 GNDA.t70 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X52 GNDA.t19 div120_0.div8.t3 div120_0.div3_2_0.CLK.t1 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X53 VDDA.t85 div120_0.div4.t4 div120_0.div2_3_2.A.t0 VDDA.t84 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X54 a_1492_966.t1 a_110_1544.t4 VDDA.t79 VDDA.t78 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=1.5
X55 GNDA.t16 V_CONT.t3 a_110_1544.t0 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X56 GNDA.t83 div120_0.div3_2_0.CLK.t8 div120_0.div3_2_0.H.t1 GNDA.t82 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X57 a_938_966.t1 a_110_1544.t5 VDDA.t77 VDDA.t76 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=1.5
X58 VDDA.t63 div120_0.div5_0.G.t3 div120_0.div5_0.J.t0 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X59 div120_0.div3_2_0.D.t1 div120_0.div3_2_0.CLK.t9 VDDA.t69 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X60 a_1492_966.t0 a_1460_718.t2 a_906_718.t0 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.16
X61 VDDA.t5 div120_0.div3_2_0.I.t6 div120_0.div24.t0 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X62 a_938_966.t0 a_906_718.t2 V_OSC.t1 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.16
X63 div120_0.div2_3_0.CLK.t0 div120_0.div4.t5 VDDA.t9 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X64 div120_0.div2_3_1.B.t1 div120_0.div2.t3 GNDA.t99 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X65 div120_0.div2_3_0.B.t1 div120_0.div8.t4 GNDA.t36 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X66 a_2046_228.t1 V_OSC.t5 a_1460_718.t0 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.16
X67 VDDA.t73 div120_0.div8.t5 div120_0.div2_3_0.A.t1 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X68 div120_0.div5_0.I.t1 div120_0.div5_0.Q2_b.t5 div120_0.div5_0.H.t1 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X69 div120_0.div5_0.F.t1 div120_0.div5_0.E.t3 VDDA.t52 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X70 VDDA.t41 V_OSC.t6 div120_0.div2_3_1.CLK.t0 VDDA.t40 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X71 GNDA.t1 div120_0.div2_3_2.CLK.t5 div120_0.div2_3_2.C.t2 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X72 GNDA.t81 div120_0.div3_2_0.CLK.t10 div120_0.div3_2_0.C.t1 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X73 div120_0.div2_3_1.C.t0 div120_0.div2_3_1.A.t2 VDDA.t16 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X74 GNDA.t14 div120_0.div24.t7 div120_0.div5_0.D.t2 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X75 GNDA.t79 div120_0.div3_2_0.CLK.t11 div120_0.div3_2_0.H.t0 GNDA.t78 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X76 div120_0.div5_0.D.t0 div120_0.div5_0.B.t2 VDDA.t20 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X77 a_1492_228.t0 a_1460_718.t3 a_906_718.t1 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.16
X78 a_938_228.t1 a_906_718.t3 V_OSC.t0 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.16
X79 div120_0.div5_0.A.t2 div120_0.div5_0.Q2_b.t6 GNDA.t117 GNDA.t116 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X80 VDDA.t3 div120_0.div24.t8 div120_0.div3_2_0.A.t1 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X81 VDDA.t1 div120_0.div2.t4 div120_0.div2_3_2.CLK.t0 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X82 div120_0.div8.t1 div120_0.div2_3_0.C.t4 GNDA.t93 GNDA.t92 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X83 div120_0.div5_0.K.t1 div120_0.div5_0.Q2_b.t7 div120_0.div5_0.L.t1 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X84 div120_0.div2.t0 div120_0.div2_3_1.C.t4 GNDA.t10 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X85 div120_0.div2.t1 div120_0.div2_3_1.CLK.t5 VDDA.t46 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X86 GNDA.t50 div120_0.div5_0.Q2_b.t8 div120_0.div5_0.M.t2 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X87 GNDA.t31 div120_0.div24.t9 div120_0.div5_0.J.t2 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X88 GNDA.t75 div120_0.div2_3_2.CLK.t6 div120_0.div2_3_2.C.t1 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X89 GNDA.t97 div120_0.div2.t5 div120_0.div2_3_2.CLK.t2 GNDA.t96 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X90 div120_0.div4.t1 div120_0.div2_3_2.CLK.t7 VDDA.t61 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X91 div120_0.div2_3_0.C.t0 div120_0.div2_3_0.CLK.t5 GNDA.t21 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X92 div120_0.div2_3_1.C.t1 div120_0.div2_3_1.CLK.t6 GNDA.t60 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X93 GNDA.t46 div120_0.div5_0.Q2_b.t9 div120_0.div5_0.M.t0 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X94 VDDA.t22 div120_0.div2.t6 div120_0.div2_3_1.A.t1 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X95 GNDA.t110 div120_0.div24.t10 div120_0.div5_0.J.t1 GNDA.t109 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X96 div120_0.div3_2_0.G.t0 div120_0.div3_2_0.D.t2 div120_0.div3_2_0.F.t1 GNDA.t65 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X97 div120_0.div8.t0 div120_0.div2_3_0.CLK.t6 VDDA.t14 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X98 GNDA.t54 div120_0.div4.t6 div120_0.div2_3_0.CLK.t2 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X99 VDDA.t89 div120_0.div5_0.Q2_b.t10 div120_0.div5_0.A.t0 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X100 div120_0.div3_2_0.CLK.t0 div120_0.div8.t6 VDDA.t11 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X101 div120_0.div5_0.B.t1 div120_0.div24.t11 div120_0.div5_0.C.t1 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X102 VDDA.t56 div120_0.div3_2_0.E.t3 div120_0.div3_2_0.H.t3 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X103 div120_0.div3_2_0.B.t1 div120_0.div24.t12 GNDA.t34 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X104 V_OUT120.t1 div120_0.div5_0.Q2_b.t11 VDDA.t91 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X105 a_1492_966.t2 GNDA.t120 VDDA.t24 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.15
X106 div120_0.div2_3_2.C.t0 div120_0.div2_3_2.A.t2 VDDA.t54 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X107 div120_0.div3_2_0.I.t1 div120_0.div3_2_0.H.t4 GNDA.t12 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X108 VDDA.t65 V_OUT120.t5 div120_0.div5_0.K.t0 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X109 GNDA.t77 div120_0.div3_2_0.CLK.t12 div120_0.div3_2_0.C.t0 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X110 div120_0.div5_0.Q2_b.t0 div120_0.div24.t13 VDDA.t37 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X111 GNDA.t107 div120_0.div24.t14 div120_0.div5_0.D.t1 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X112 div120_0.div2_3_1.A.t0 div120_0.div2_3_1.CLK.t7 div120_0.div2_3_1.B.t0 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X113 VDDA.t58 div120_0.div3_2_0.D.t3 div120_0.div3_2_0.E.t1 VDDA.t57 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X114 div120_0.div2_3_0.A.t0 div120_0.div2_3_0.CLK.t7 div120_0.div2_3_0.B.t0 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X115 div120_0.div2_3_0.C.t3 div120_0.div2_3_0.A.t2 VDDA.t67 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
R0 a_110_1544.t0 a_110_1544.n2 466.82
R1 a_110_1544.n2 a_110_1544.t1 225.869
R2 a_110_1544.n2 a_110_1544.t2 225.786
R3 a_110_1544.t1 a_110_1544.n1 188.501
R4 a_110_1544.n0 a_110_1544.t3 188.501
R5 a_110_1544.n1 a_110_1544.n0 107.442
R6 a_110_1544.n1 a_110_1544.t5 81.0592
R7 a_110_1544.n0 a_110_1544.t4 81.0592
R8 VDDA.t17 VDDA.t86 2804.76
R9 VDDA.t64 VDDA.t36 2533.33
R10 VDDA.t68 VDDA.t57 2307.14
R11 VDDA.t70 VDDA.t49 2126.19
R12 VDDA.t31 VDDA.t13 2080.95
R13 VDDA.t60 VDDA.t92 2080.95
R14 VDDA.t0 VDDA.t45 2080.95
R15 VDDA.t25 VDDA.t33 1538.1
R16 VDDA.t62 VDDA.t59 1492.86
R17 VDDA.t6 VDDA.t55 1492.86
R18 VDDA.t47 VDDA.t40 1406.73
R19 VDDA.n10 VDDA.t29 1289.29
R20 VDDA.t19 VDDA.n31 1289.29
R21 VDDA.t4 VDDA.t88 1130.95
R22 VDDA.t2 VDDA.t10 1130.95
R23 VDDA.t8 VDDA.t72 1130.95
R24 VDDA.t84 VDDA.t38 1130.95
R25 VDDA.t43 VDDA.t21 1130.95
R26 VDDA.n1 VDDA.t94 1007.38
R27 VDDA.n32 VDDA.t74 927.381
R28 VDDA.t66 VDDA.n46 927.381
R29 VDDA.n47 VDDA.t53 927.381
R30 VDDA.t15 VDDA.n62 927.381
R31 VDDA.n23 VDDA.t50 673.101
R32 VDDA.n24 VDDA.t5 673.101
R33 VDDA.n11 VDDA.t91 667.62
R34 VDDA.n3 VDDA.t46 663.801
R35 VDDA.n5 VDDA.t61 663.801
R36 VDDA.n6 VDDA.t14 663.801
R37 VDDA.n8 VDDA.t69 663.801
R38 VDDA.n9 VDDA.t87 663.801
R39 VDDA.n2 VDDA.t96 618.567
R40 VDDA.n10 VDDA.t90 610.715
R41 VDDA.n31 VDDA.t86 610.715
R42 VDDA.n32 VDDA.t68 610.715
R43 VDDA.n46 VDDA.t13 610.715
R44 VDDA.n47 VDDA.t60 610.715
R45 VDDA.n62 VDDA.t45 610.715
R46 VDDA.n57 VDDA.n56 594.301
R47 VDDA.n59 VDDA.n58 594.301
R48 VDDA.n53 VDDA.n52 594.301
R49 VDDA.n51 VDDA.n50 594.301
R50 VDDA.n41 VDDA.n40 594.301
R51 VDDA.n43 VDDA.n42 594.301
R52 VDDA.n38 VDDA.n37 594.301
R53 VDDA.n36 VDDA.n35 594.301
R54 VDDA.n20 VDDA.n19 594.301
R55 VDDA.n22 VDDA.n21 594.301
R56 VDDA.n26 VDDA.n25 594.301
R57 VDDA.n28 VDDA.n27 594.301
R58 VDDA.n17 VDDA.n16 594.301
R59 VDDA.n15 VDDA.n14 594.301
R60 VDDA.n13 VDDA.n12 594.301
R61 VDDA.t29 VDDA.t64 497.62
R62 VDDA.t36 VDDA.t62 497.62
R63 VDDA.t59 VDDA.t51 497.62
R64 VDDA.t51 VDDA.t17 497.62
R65 VDDA.t33 VDDA.t19 497.62
R66 VDDA.t88 VDDA.t25 497.62
R67 VDDA.t49 VDDA.t4 497.62
R68 VDDA.t55 VDDA.t70 497.62
R69 VDDA.t57 VDDA.t6 497.62
R70 VDDA.t74 VDDA.t2 497.62
R71 VDDA.t10 VDDA.t31 497.62
R72 VDDA.t72 VDDA.t66 497.62
R73 VDDA.t92 VDDA.t8 497.62
R74 VDDA.t53 VDDA.t84 497.62
R75 VDDA.t38 VDDA.t0 497.62
R76 VDDA.t21 VDDA.t15 497.62
R77 VDDA.t40 VDDA.t43 497.62
R78 VDDA.t76 VDDA.t80 488.219
R79 VDDA.t23 VDDA.t82 480.288
R80 VDDA.n11 VDDA.n10 373.781
R81 VDDA.n31 VDDA.n30 370
R82 VDDA.n33 VDDA.n32 370
R83 VDDA.n46 VDDA.n45 370
R84 VDDA.n48 VDDA.n47 370
R85 VDDA.n62 VDDA.n61 370
R86 VDDA.n64 VDDA.n2 357.406
R87 VDDA.n67 VDDA.t28 354.418
R88 VDDA.n55 VDDA.t48 354.418
R89 VDDA.n64 VDDA.t24 349.767
R90 VDDA.n63 VDDA.t27 341.048
R91 VDDA.n2 VDDA.n1 308.481
R92 VDDA.n64 VDDA.n63 185
R93 VDDA.n69 VDDA.t81 143.486
R94 VDDA.n68 VDDA.t77 143.486
R95 VDDA.n66 VDDA.t79 143.486
R96 VDDA.n0 VDDA.t83 143.486
R97 VDDA.n63 VDDA.t78 139.239
R98 VDDA.n1 VDDA.t95 117.287
R99 VDDA.n56 VDDA.t44 78.8005
R100 VDDA.n56 VDDA.t41 78.8005
R101 VDDA.n58 VDDA.t16 78.8005
R102 VDDA.n58 VDDA.t22 78.8005
R103 VDDA.n52 VDDA.t39 78.8005
R104 VDDA.n52 VDDA.t1 78.8005
R105 VDDA.n50 VDDA.t54 78.8005
R106 VDDA.n50 VDDA.t85 78.8005
R107 VDDA.n40 VDDA.t9 78.8005
R108 VDDA.n40 VDDA.t93 78.8005
R109 VDDA.n42 VDDA.t67 78.8005
R110 VDDA.n42 VDDA.t73 78.8005
R111 VDDA.n37 VDDA.t11 78.8005
R112 VDDA.n37 VDDA.t32 78.8005
R113 VDDA.n35 VDDA.t75 78.8005
R114 VDDA.n35 VDDA.t3 78.8005
R115 VDDA.n19 VDDA.t7 78.8005
R116 VDDA.n19 VDDA.t58 78.8005
R117 VDDA.n21 VDDA.t71 78.8005
R118 VDDA.n21 VDDA.t56 78.8005
R119 VDDA.n25 VDDA.t26 78.8005
R120 VDDA.n25 VDDA.t89 78.8005
R121 VDDA.n27 VDDA.t20 78.8005
R122 VDDA.n27 VDDA.t34 78.8005
R123 VDDA.n16 VDDA.t52 78.8005
R124 VDDA.n16 VDDA.t18 78.8005
R125 VDDA.n14 VDDA.t37 78.8005
R126 VDDA.n14 VDDA.t63 78.8005
R127 VDDA.n12 VDDA.t30 78.8005
R128 VDDA.n12 VDDA.t65 78.8005
R129 VDDA.n61 VDDA.n3 12.8005
R130 VDDA.n48 VDDA.n5 12.8005
R131 VDDA.n45 VDDA.n6 12.8005
R132 VDDA.n33 VDDA.n8 12.8005
R133 VDDA.n30 VDDA.n9 12.8005
R134 VDDA.n18 VDDA.n9 9.3005
R135 VDDA.n30 VDDA.n29 9.3005
R136 VDDA.n8 VDDA.n7 9.3005
R137 VDDA.n34 VDDA.n33 9.3005
R138 VDDA.n39 VDDA.n6 9.3005
R139 VDDA.n45 VDDA.n44 9.3005
R140 VDDA.n5 VDDA.n4 9.3005
R141 VDDA.n49 VDDA.n48 9.3005
R142 VDDA.n54 VDDA.n3 9.3005
R143 VDDA.n61 VDDA.n60 9.3005
R144 VDDA.t82 VDDA.t42 7.05059
R145 VDDA.t78 VDDA.t12 7.05059
R146 VDDA.t35 VDDA.t76 7.05059
R147 VDDA.n13 VDDA.n11 3.20124
R148 VDDA.n65 VDDA.n64 2.32108
R149 VDDA.n18 VDDA.n17 0.913
R150 VDDA.t42 VDDA.t47 0.881762
R151 VDDA.t12 VDDA.t23 0.881762
R152 VDDA.t27 VDDA.t35 0.881762
R153 VDDA.n15 VDDA.n13 0.838
R154 VDDA.n20 VDDA.n7 0.7755
R155 VDDA.n17 VDDA.n15 0.688
R156 VDDA.n23 VDDA.n22 0.588
R157 VDDA.n28 VDDA.n26 0.563
R158 VDDA.n22 VDDA.n20 0.5505
R159 VDDA.n39 VDDA 0.4755
R160 VDDA VDDA.n4 0.4755
R161 VDDA.n54 VDDA 0.4755
R162 VDDA.n38 VDDA.n36 0.4505
R163 VDDA.n43 VDDA.n41 0.4505
R164 VDDA.n53 VDDA.n51 0.4505
R165 VDDA.n59 VDDA.n57 0.4505
R166 VDDA.n29 VDDA.n28 0.4255
R167 VDDA.n36 VDDA.n34 0.3255
R168 VDDA.n44 VDDA.n43 0.3255
R169 VDDA.n51 VDDA.n49 0.3255
R170 VDDA.n60 VDDA.n59 0.3255
R171 VDDA.n24 VDDA.n23 0.2755
R172 VDDA VDDA.n55 0.268714
R173 VDDA.n26 VDDA 0.238
R174 VDDA VDDA.n38 0.238
R175 VDDA.n41 VDDA 0.238
R176 VDDA VDDA.n53 0.238
R177 VDDA.n57 VDDA 0.238
R178 VDDA.n29 VDDA.n18 0.1005
R179 VDDA.n34 VDDA.n7 0.1005
R180 VDDA.n44 VDDA.n39 0.1005
R181 VDDA.n49 VDDA.n4 0.1005
R182 VDDA.n60 VDDA.n54 0.1005
R183 VDDA.n65 VDDA.n0 0.0901819
R184 VDDA VDDA.n69 0.0875743
R185 VDDA.n67 VDDA.n66 0.0798344
R186 VDDA VDDA.n24 0.0755
R187 VDDA.n69 VDDA.n68 0.0302988
R188 VDDA.n55 VDDA.n0 0.0283638
R189 VDDA.n68 VDDA.n67 0.0283638
R190 VDDA.n66 VDDA.n65 0.0189745
R191 a_2046_966.n0 a_2046_966.t0 398.087
R192 a_2046_966.t1 a_2046_966.n0 349.767
R193 a_2046_966.n0 a_2046_966.t2 212.364
R194 div120_0.div5_0.E.n0 div120_0.div5_0.E.t3 1207.57
R195 div120_0.div5_0.E.n0 div120_0.div5_0.E.t1 723
R196 div120_0.div5_0.E.t3 div120_0.div5_0.E.t2 514.134
R197 div120_0.div5_0.E.t0 div120_0.div5_0.E.n0 314.921
R198 div120_0.div5_0.I.t0 div120_0.div5_0.I.n0 531.067
R199 div120_0.div5_0.I.n0 div120_0.div5_0.I.t2 48.0005
R200 div120_0.div5_0.I.n0 div120_0.div5_0.I.t1 48.0005
R201 GNDA.t52 GNDA.t15 2694.17
R202 GNDA.t51 GNDA.t28 2627.65
R203 GNDA.t4 GNDA.t56 2472.44
R204 GNDA.n64 GNDA.t7 1848.38
R205 GNDA.t68 GNDA.t116 1619.63
R206 GNDA.t39 GNDA.t32 1574.64
R207 GNDA.t113 GNDA.t72 1529.65
R208 GNDA.t70 GNDA.t109 1484.66
R209 GNDA.t84 GNDA.t66 1484.66
R210 GNDA.t76 GNDA.t85 1484.66
R211 GNDA.t17 GNDA.t24 1484.66
R212 GNDA.t74 GNDA.t6 1484.66
R213 GNDA.t58 GNDA.t61 1484.66
R214 GNDA.t116 GNDA.n29 1417.18
R215 GNDA.n47 GNDA.n46 1179.3
R216 GNDA.n49 GNDA.n48 1179.3
R217 GNDA.n63 GNDA.n62 1179.3
R218 GNDA.n65 GNDA.n64 1170
R219 GNDA.n31 GNDA.n30 1170
R220 GNDA.n29 GNDA.n28 1170
R221 GNDA.t115 GNDA.t45 1124.74
R222 GNDA.t108 GNDA.t106 1124.74
R223 GNDA.t11 GNDA.t68 1124.74
R224 GNDA.n2 GNDA.t119 1076.47
R225 GNDA.n30 GNDA.t78 877.302
R226 GNDA.n47 GNDA.t18 877.302
R227 GNDA.t92 GNDA.n47 877.302
R228 GNDA.n48 GNDA.t53 877.302
R229 GNDA.n48 GNDA.t43 877.302
R230 GNDA.n63 GNDA.t96 877.302
R231 GNDA.t9 GNDA.n63 877.302
R232 GNDA.n64 GNDA.t55 779.266
R233 GNDA.n29 GNDA.t47 607.362
R234 GNDA.n30 GNDA.t94 607.362
R235 GNDA.n3 GNDA.n2 504.493
R236 GNDA.t49 GNDA.t41 494.889
R237 GNDA.t111 GNDA.t49 494.889
R238 GNDA.t45 GNDA.t111 494.889
R239 GNDA.t72 GNDA.t115 494.889
R240 GNDA.t30 GNDA.t113 494.889
R241 GNDA.t37 GNDA.t30 494.889
R242 GNDA.t109 GNDA.t37 494.889
R243 GNDA.t104 GNDA.t70 494.889
R244 GNDA.t100 GNDA.t104 494.889
R245 GNDA.t32 GNDA.t100 494.889
R246 GNDA.t13 GNDA.t39 494.889
R247 GNDA.t26 GNDA.t13 494.889
R248 GNDA.t106 GNDA.t26 494.889
R249 GNDA.t47 GNDA.t108 494.889
R250 GNDA.t82 GNDA.t11 494.889
R251 GNDA.t88 GNDA.t82 494.889
R252 GNDA.t78 GNDA.t88 494.889
R253 GNDA.t94 GNDA.t65 494.889
R254 GNDA.t65 GNDA.t84 494.889
R255 GNDA.t66 GNDA.t80 494.889
R256 GNDA.t80 GNDA.t86 494.889
R257 GNDA.t86 GNDA.t76 494.889
R258 GNDA.t85 GNDA.t33 494.889
R259 GNDA.t33 GNDA.t18 494.889
R260 GNDA.t22 GNDA.t92 494.889
R261 GNDA.t20 GNDA.t22 494.889
R262 GNDA.t24 GNDA.t20 494.889
R263 GNDA.t35 GNDA.t17 494.889
R264 GNDA.t53 GNDA.t35 494.889
R265 GNDA.t43 GNDA.t0 494.889
R266 GNDA.t0 GNDA.t2 494.889
R267 GNDA.t2 GNDA.t74 494.889
R268 GNDA.t6 GNDA.t90 494.889
R269 GNDA.t90 GNDA.t96 494.889
R270 GNDA.t63 GNDA.t9 494.889
R271 GNDA.t59 GNDA.t63 494.889
R272 GNDA.t61 GNDA.t59 494.889
R273 GNDA.t98 GNDA.t58 494.889
R274 GNDA.t56 GNDA.t98 494.889
R275 GNDA.n3 GNDA.t118 491.64
R276 GNDA.n65 GNDA.n3 352.723
R277 GNDA.n68 GNDA.t101 264.067
R278 GNDA.n67 GNDA.t102 264.067
R279 GNDA.n1 GNDA.t103 254.768
R280 GNDA.n25 GNDA.t69 242.3
R281 GNDA.n26 GNDA.t117 242.3
R282 GNDA.n9 GNDA.t73 242.3
R283 GNDA.n32 GNDA.t95 233
R284 GNDA.n5 GNDA.t48 233
R285 GNDA.n8 GNDA.n6 194.576
R286 GNDA.n57 GNDA.n56 194.3
R287 GNDA.n59 GNDA.n58 194.3
R288 GNDA.n61 GNDA.n60 194.3
R289 GNDA.n55 GNDA.n54 194.3
R290 GNDA.n53 GNDA.n52 194.3
R291 GNDA.n51 GNDA.n50 194.3
R292 GNDA.n41 GNDA.n40 194.3
R293 GNDA.n43 GNDA.n42 194.3
R294 GNDA.n45 GNDA.n44 194.3
R295 GNDA.n39 GNDA.n38 194.3
R296 GNDA.n37 GNDA.n36 194.3
R297 GNDA.n35 GNDA.n34 194.3
R298 GNDA.n22 GNDA.n21 194.3
R299 GNDA.n24 GNDA.n23 194.3
R300 GNDA.n19 GNDA.n18 194.3
R301 GNDA.n17 GNDA.n16 194.3
R302 GNDA.n15 GNDA.n14 194.3
R303 GNDA.n13 GNDA.n12 194.3
R304 GNDA.n11 GNDA.n10 194.3
R305 GNDA.n8 GNDA.n7 194.3
R306 GNDA.n2 GNDA.t120 186.374
R307 GNDA.n69 GNDA.t16 127.15
R308 GNDA.n68 GNDA.t29 127.15
R309 GNDA.n67 GNDA.t8 127.15
R310 GNDA.n0 GNDA.t5 127.15
R311 GNDA.n56 GNDA.t99 48.0005
R312 GNDA.n56 GNDA.t57 48.0005
R313 GNDA.n58 GNDA.t60 48.0005
R314 GNDA.n58 GNDA.t62 48.0005
R315 GNDA.n60 GNDA.t10 48.0005
R316 GNDA.n60 GNDA.t64 48.0005
R317 GNDA.n54 GNDA.t91 48.0005
R318 GNDA.n54 GNDA.t97 48.0005
R319 GNDA.n52 GNDA.t3 48.0005
R320 GNDA.n52 GNDA.t75 48.0005
R321 GNDA.n50 GNDA.t44 48.0005
R322 GNDA.n50 GNDA.t1 48.0005
R323 GNDA.n40 GNDA.t36 48.0005
R324 GNDA.n40 GNDA.t54 48.0005
R325 GNDA.n42 GNDA.t21 48.0005
R326 GNDA.n42 GNDA.t25 48.0005
R327 GNDA.n44 GNDA.t93 48.0005
R328 GNDA.n44 GNDA.t23 48.0005
R329 GNDA.n38 GNDA.t34 48.0005
R330 GNDA.n38 GNDA.t19 48.0005
R331 GNDA.n36 GNDA.t87 48.0005
R332 GNDA.n36 GNDA.t77 48.0005
R333 GNDA.n34 GNDA.t67 48.0005
R334 GNDA.n34 GNDA.t81 48.0005
R335 GNDA.n21 GNDA.t89 48.0005
R336 GNDA.n21 GNDA.t79 48.0005
R337 GNDA.n23 GNDA.t12 48.0005
R338 GNDA.n23 GNDA.t83 48.0005
R339 GNDA.n18 GNDA.t27 48.0005
R340 GNDA.n18 GNDA.t107 48.0005
R341 GNDA.n16 GNDA.t40 48.0005
R342 GNDA.n16 GNDA.t14 48.0005
R343 GNDA.n14 GNDA.t71 48.0005
R344 GNDA.n14 GNDA.t105 48.0005
R345 GNDA.n12 GNDA.t38 48.0005
R346 GNDA.n12 GNDA.t110 48.0005
R347 GNDA.n10 GNDA.t114 48.0005
R348 GNDA.n10 GNDA.t31 48.0005
R349 GNDA.n7 GNDA.t112 48.0005
R350 GNDA.n7 GNDA.t46 48.0005
R351 GNDA.n6 GNDA.t42 48.0005
R352 GNDA.n6 GNDA.t50 48.0005
R353 GNDA.n65 GNDA.n1 14.8842
R354 GNDA.n32 GNDA.n31 12.8005
R355 GNDA.n28 GNDA.n5 12.8005
R356 GNDA.n20 GNDA.n5 9.3005
R357 GNDA.n28 GNDA.n27 9.3005
R358 GNDA.n31 GNDA.n4 9.3005
R359 GNDA.n33 GNDA.n32 9.3005
R360 GNDA.n1 GNDA.n0 9.3005
R361 GNDA.n66 GNDA.n65 9.3005
R362 GNDA.t55 GNDA.t4 4.75212
R363 GNDA.t7 GNDA.t51 4.75212
R364 GNDA.t28 GNDA.t52 4.75212
R365 GNDA.n17 GNDA.n15 0.8505
R366 GNDA.n35 GNDA.n33 0.8255
R367 GNDA.n39 GNDA.n37 0.688
R368 GNDA.n43 GNDA.n41 0.688
R369 GNDA.n55 GNDA.n53 0.688
R370 GNDA.n59 GNDA.n57 0.688
R371 GNDA.n9 GNDA.n8 0.588
R372 GNDA.n20 GNDA.n19 0.588
R373 GNDA.n15 GNDA.n13 0.5505
R374 GNDA.n27 GNDA.n26 0.463
R375 GNDA.n11 GNDA.n9 0.4255
R376 GNDA GNDA.n25 0.3505
R377 GNDA.n25 GNDA.n24 0.313
R378 GNDA.n22 GNDA.n4 0.313
R379 GNDA.n46 GNDA.n45 0.313
R380 GNDA.n51 GNDA.n49 0.313
R381 GNDA.n62 GNDA.n61 0.313
R382 GNDA.n13 GNDA.n11 0.2755
R383 GNDA.n19 GNDA.n17 0.2755
R384 GNDA.n24 GNDA.n22 0.2755
R385 GNDA.n37 GNDA.n35 0.2755
R386 GNDA.n45 GNDA.n43 0.2755
R387 GNDA.n53 GNDA.n51 0.2755
R388 GNDA.n61 GNDA.n59 0.2755
R389 GNDA GNDA.n39 0.238
R390 GNDA.n41 GNDA 0.238
R391 GNDA GNDA.n55 0.238
R392 GNDA.n57 GNDA 0.238
R393 GNDA.n68 GNDA.n67 0.192861
R394 GNDA GNDA.n0 0.177962
R395 GNDA.n67 GNDA.n66 0.158139
R396 GNDA.n69 GNDA.n68 0.152583
R397 GNDA.n27 GNDA.n20 0.1005
R398 GNDA.n26 GNDA 0.1005
R399 GNDA.n33 GNDA.n4 0.1005
R400 GNDA.n46 GNDA 0.0755
R401 GNDA.n49 GNDA 0.0755
R402 GNDA.n62 GNDA 0.0755
R403 GNDA GNDA.n69 0.063
R404 GNDA.n66 GNDA.n0 0.0352222
R405 div120_0.div3_2_0.C.n2 div120_0.div3_2_0.C.t3 721.4
R406 div120_0.div3_2_0.C.n1 div120_0.div3_2_0.C.t4 350.349
R407 div120_0.div3_2_0.C.t0 div120_0.div3_2_0.C.n2 276.733
R408 div120_0.div3_2_0.C.n1 div120_0.div3_2_0.C.n0 206.333
R409 div120_0.div3_2_0.C.n0 div120_0.div3_2_0.C.t1 48.0005
R410 div120_0.div3_2_0.C.n0 div120_0.div3_2_0.C.t2 48.0005
R411 div120_0.div3_2_0.C.n2 div120_0.div3_2_0.C.n1 48.0005
R412 div120_0.div3_2_0.D.n1 div120_0.div3_2_0.D.n0 701.467
R413 div120_0.div3_2_0.D.n1 div120_0.div3_2_0.D.t1 694.201
R414 div120_0.div3_2_0.D.n0 div120_0.div3_2_0.D.t2 321.334
R415 div120_0.div3_2_0.D.t0 div120_0.div3_2_0.D.n1 314.921
R416 div120_0.div3_2_0.D.n0 div120_0.div3_2_0.D.t3 144.601
R417 V_OSC.n3 V_OSC.n2 2160.31
R418 V_OSC.t6 V_OSC.t2 401.668
R419 V_OSC.n2 V_OSC.t1 374.728
R420 V_OSC.n2 V_OSC.t0 271.567
R421 V_OSC.n0 V_OSC.t6 257.067
R422 div120_0.div2_3_1.VIN V_OSC.n0 216.9
R423 V_OSC.n0 V_OSC.t3 208.868
R424 V_OSC.n1 V_OSC.t4 199.686
R425 vco2_2_0.V_OSC div120_0.VIN 182.5
R426 V_OSC.n3 V_OSC.n1 181.013
R427 V_OSC.n1 V_OSC.t5 128.893
R428 vco2_2_0.V_OSC V_OSC.n3 44.8005
R429 div120_0.VIN div120_0.div2_3_1.VIN 32.1338
R430 div120_0.div2_3_1.CLK.n4 div120_0.div2_3_1.CLK.t0 723.534
R431 div120_0.div2_3_1.CLK.t1 div120_0.div2_3_1.CLK.n5 723.534
R432 div120_0.div2_3_1.CLK.n0 div120_0.div2_3_1.CLK.t5 369.534
R433 div120_0.div2_3_1.CLK.n3 div120_0.div2_3_1.CLK.n2 366.856
R434 div120_0.div2_3_1.CLK.n4 div120_0.div2_3_1.CLK.t2 254.333
R435 div120_0.div2_3_1.CLK.n3 div120_0.div2_3_1.CLK.t7 190.123
R436 div120_0.div2_3_1.CLK.n5 div120_0.div2_3_1.CLK.n3 187.201
R437 div120_0.div2_3_1.CLK.n1 div120_0.div2_3_1.CLK.n0 176.733
R438 div120_0.div2_3_1.CLK.n2 div120_0.div2_3_1.CLK.n1 176.733
R439 div120_0.div2_3_1.CLK.n0 div120_0.div2_3_1.CLK.t3 112.468
R440 div120_0.div2_3_1.CLK.n2 div120_0.div2_3_1.CLK.t4 112.468
R441 div120_0.div2_3_1.CLK.n1 div120_0.div2_3_1.CLK.t6 112.468
R442 div120_0.div2_3_1.CLK.n5 div120_0.div2_3_1.CLK.n4 70.4005
R443 V_OUT120.n2 V_OUT120.n1 2120.39
R444 V_OUT120.n1 V_OUT120.t2 1992.27
R445 V_OUT120.n3 V_OUT120.t1 751.801
R446 V_OUT120.t2 V_OUT120.t4 514.134
R447 V_OUT120.n0 V_OUT120.t3 289.2
R448 V_OUT120.n2 V_OUT120.t0 233
R449 V_OUT120.n1 V_OUT120.n0 208.868
R450 V_OUT120.n0 V_OUT120.t5 176.733
R451 V_OUT120.n3 V_OUT120.n2 40.3205
R452 V_OUT120 V_OUT120.n3 32.0005
R453 div120_0.div5_0.F.t0 div120_0.div5_0.F.t1 157.601
R454 div120_0.div5_0.G.n0 div120_0.div5_0.G.t0 685.134
R455 div120_0.div5_0.G.n1 div120_0.div5_0.G.t1 685.134
R456 div120_0.div5_0.G.n0 div120_0.div5_0.G.t3 534.268
R457 div120_0.div5_0.G.t2 div120_0.div5_0.G.n1 340.521
R458 div120_0.div5_0.G.n1 div120_0.div5_0.G.n0 105.6
R459 div120_0.div3_2_0.CLK.n3 div120_0.div3_2_0.CLK.n2 742.51
R460 div120_0.div3_2_0.CLK.n9 div120_0.div3_2_0.CLK.t2 723.534
R461 div120_0.div3_2_0.CLK.n8 div120_0.div3_2_0.CLK.t0 723.534
R462 div120_0.div3_2_0.CLK.n2 div120_0.div3_2_0.CLK.n1 684.806
R463 div120_0.div3_2_0.CLK.n7 div120_0.div3_2_0.CLK.n6 366.856
R464 div120_0.div3_2_0.CLK.n0 div120_0.div3_2_0.CLK.t7 337.401
R465 div120_0.div3_2_0.CLK.n0 div120_0.div3_2_0.CLK.t8 305.267
R466 div120_0.div3_2_0.CLK.t1 div120_0.div3_2_0.CLK.n9 254.333
R467 div120_0.div3_2_0.CLK.n4 div120_0.div3_2_0.CLK.n3 224.934
R468 div120_0.div3_2_0.CLK.n7 div120_0.div3_2_0.CLK.t5 190.123
R469 div120_0.div3_2_0.CLK.n8 div120_0.div3_2_0.CLK.n7 187.201
R470 div120_0.div3_2_0.CLK.n1 div120_0.div3_2_0.CLK.n0 176.733
R471 div120_0.div3_2_0.CLK.n5 div120_0.div3_2_0.CLK.n4 176.733
R472 div120_0.div3_2_0.CLK.n6 div120_0.div3_2_0.CLK.n5 176.733
R473 div120_0.div3_2_0.CLK.n3 div120_0.div3_2_0.CLK.t9 144.601
R474 div120_0.div3_2_0.CLK.n2 div120_0.div3_2_0.CLK.t6 131.976
R475 div120_0.div3_2_0.CLK.n0 div120_0.div3_2_0.CLK.t3 128.534
R476 div120_0.div3_2_0.CLK.n1 div120_0.div3_2_0.CLK.t11 128.534
R477 div120_0.div3_2_0.CLK.n4 div120_0.div3_2_0.CLK.t10 112.468
R478 div120_0.div3_2_0.CLK.n6 div120_0.div3_2_0.CLK.t12 112.468
R479 div120_0.div3_2_0.CLK.n5 div120_0.div3_2_0.CLK.t4 112.468
R480 div120_0.div3_2_0.CLK.n9 div120_0.div3_2_0.CLK.n8 70.4005
R481 div120_0.div3_2_0.H.n0 div120_0.div3_2_0.H.t3 723.534
R482 div120_0.div3_2_0.H.n1 div120_0.div3_2_0.H.t4 553.534
R483 div120_0.div3_2_0.H.n0 div120_0.div3_2_0.H.t0 254.333
R484 div120_0.div3_2_0.H.n2 div120_0.div3_2_0.H.n1 206.333
R485 div120_0.div3_2_0.H.n1 div120_0.div3_2_0.H.n0 70.4005
R486 div120_0.div3_2_0.H.n2 div120_0.div3_2_0.H.t1 48.0005
R487 div120_0.div3_2_0.H.t2 div120_0.div3_2_0.H.n2 48.0005
R488 div120_0.div3_2_0.I.n0 div120_0.div3_2_0.I.t0 663.801
R489 div120_0.div3_2_0.I.n0 div120_0.div3_2_0.I.t5 568.067
R490 div120_0.div3_2_0.I.t5 div120_0.div3_2_0.I.t3 514.134
R491 div120_0.div3_2_0.I.n3 div120_0.div3_2_0.I.n2 344.8
R492 div120_0.div3_2_0.I.n1 div120_0.div3_2_0.I.t6 289.2
R493 div120_0.div3_2_0.I.t1 div120_0.div3_2_0.I.n3 275.454
R494 div120_0.div3_2_0.I.n2 div120_0.div3_2_0.I.t4 241
R495 div120_0.div3_2_0.I.n1 div120_0.div3_2_0.I.t2 112.468
R496 div120_0.div3_2_0.I.n3 div120_0.div3_2_0.I.n0 97.9205
R497 div120_0.div3_2_0.I.n2 div120_0.div3_2_0.I.n1 64.2672
R498 div120_0.div24.n10 div120_0.div24.t12 4546.23
R499 div120_0.div24.n3 div120_0.div24.n2 919.244
R500 div120_0.div3_2_0.VOUT div120_0.div24.n7 886.702
R501 div120_0.div24.t12 div120_0.div24.t8 819.4
R502 div120_0.div24.n2 div120_0.div24.n1 758.606
R503 div120_0.div24.n9 div120_0.div24.n8 628.734
R504 div120_0.div24.n7 div120_0.div24.n6 364.178
R505 div120_0.div24.n0 div120_0.div24.t13 337.401
R506 div120_0.div24.n0 div120_0.div24.t9 305.267
R507 div120_0.div24.n9 div120_0.div24.t2 257.534
R508 div120_0.div24.n4 div120_0.div24.t7 192.8
R509 div120_0.div24.n1 div120_0.div24.n0 176.733
R510 div120_0.div24.n6 div120_0.div24.n5 176.733
R511 div120_0.div24.n4 div120_0.div24.n3 160.667
R512 div120_0.div24.n3 div120_0.div24.t4 144.601
R513 div120_0.div24.n2 div120_0.div24.t3 131.976
R514 div120_0.div24.n0 div120_0.div24.t5 128.534
R515 div120_0.div24.n1 div120_0.div24.t10 128.534
R516 div120_0.div24.n6 div120_0.div24.t14 112.468
R517 div120_0.div24.n5 div120_0.div24.t6 112.468
R518 div120_0.div24.n7 div120_0.div24.t11 112.468
R519 div120_0.div24.n5 div120_0.div24.n4 96.4005
R520 div120_0.div24.n8 div120_0.div24.t0 78.8005
R521 div120_0.div24.n8 div120_0.div24.t1 78.8005
R522 div120_0.div5_0.VIN div120_0.div24.n10 28.8005
R523 div120_0.div24.n10 div120_0.div24.n9 9.6005
R524 div120_0.div5_0.VIN div120_0.div3_2_0.VOUT 6.4005
R525 V_CONT V_CONT.t3 570.367
R526 V_CONT.t3 V_CONT.n1 488.83
R527 V_CONT.n0 V_CONT.t0 486.271
R528 V_CONT.n1 V_CONT.t2 384.967
R529 V_CONT.n0 V_CONT.t1 384.967
R530 V_CONT.n1 V_CONT.n0 101.303
R531 a_2046_228.n0 a_2046_228.t1 289.967
R532 a_2046_228.n0 a_2046_228.t2 254.768
R533 a_2046_228.t0 a_2046_228.n0 161.701
R534 div120_0.div3_2_0.A.n0 div120_0.div3_2_0.A.t1 713.933
R535 div120_0.div3_2_0.A.n0 div120_0.div3_2_0.A.t2 314.233
R536 div120_0.div3_2_0.A.t0 div120_0.div3_2_0.A.n0 308.2
R537 div120_0.div2.t6 div120_0.div2.t3 819.4
R538 div120_0.div2.n0 div120_0.div2.t1 663.801
R539 div120_0.div2.n0 div120_0.div2.t6 489.168
R540 div120_0.div2.t4 div120_0.div2.t2 401.668
R541 div120_0.div2.n1 div120_0.div2.t0 270.12
R542 div120_0.div2.n2 div120_0.div2.t4 257.067
R543 div120_0.div2_3_2.VIN div120_0.div2.n2 216.9
R544 div120_0.div2.n2 div120_0.div2.t5 208.868
R545 div120_0.div2.n3 div120_0.div2_3_2.VIN 192.167
R546 div120_0.div2.n1 div120_0.div2.n0 67.2005
R547 div120_0.div2.n3 div120_0.div2.n1 25.6005
R548 div120_0.div2_3_1.VOUT div120_0.div2.n3 4.8005
R549 div120_0.div2_3_2.CLK.n4 div120_0.div2_3_2.CLK.t0 723.534
R550 div120_0.div2_3_2.CLK.t1 div120_0.div2_3_2.CLK.n5 723.534
R551 div120_0.div2_3_2.CLK.n0 div120_0.div2_3_2.CLK.t7 369.534
R552 div120_0.div2_3_2.CLK.n3 div120_0.div2_3_2.CLK.n2 366.856
R553 div120_0.div2_3_2.CLK.n4 div120_0.div2_3_2.CLK.t2 254.333
R554 div120_0.div2_3_2.CLK.n3 div120_0.div2_3_2.CLK.t4 190.123
R555 div120_0.div2_3_2.CLK.n5 div120_0.div2_3_2.CLK.n3 187.201
R556 div120_0.div2_3_2.CLK.n1 div120_0.div2_3_2.CLK.n0 176.733
R557 div120_0.div2_3_2.CLK.n2 div120_0.div2_3_2.CLK.n1 176.733
R558 div120_0.div2_3_2.CLK.n0 div120_0.div2_3_2.CLK.t5 112.468
R559 div120_0.div2_3_2.CLK.n2 div120_0.div2_3_2.CLK.t6 112.468
R560 div120_0.div2_3_2.CLK.n1 div120_0.div2_3_2.CLK.t3 112.468
R561 div120_0.div2_3_2.CLK.n5 div120_0.div2_3_2.CLK.n4 70.4005
R562 a_1492_228.n0 a_1492_228.t0 289.967
R563 a_1492_228.n0 a_1492_228.t2 254.768
R564 a_1492_228.t1 a_1492_228.n0 161.701
R565 div120_0.div5_0.M.n2 div120_0.div5_0.M.t1 761.4
R566 div120_0.div5_0.M.n1 div120_0.div5_0.M.t4 349.433
R567 div120_0.div5_0.M.t0 div120_0.div5_0.M.n2 254.333
R568 div120_0.div5_0.M.n1 div120_0.div5_0.M.n0 206.333
R569 div120_0.div5_0.M.n2 div120_0.div5_0.M.n1 70.4005
R570 div120_0.div5_0.M.n0 div120_0.div5_0.M.t2 48.0005
R571 div120_0.div5_0.M.n0 div120_0.div5_0.M.t3 48.0005
R572 div120_0.div5_0.H.t0 div120_0.div5_0.H.t1 96.0005
R573 div120_0.div5_0.Q2_b.n6 div120_0.div5_0.Q2_b.t6 2779.53
R574 div120_0.div5_0.Q2_b.n7 div120_0.div5_0.Q2_b.n6 1206
R575 div120_0.div5_0.Q2_b.n4 div120_0.div5_0.Q2_b.t0 777.4
R576 div120_0.div5_0.Q2_b.t5 div120_0.div5_0.Q2_b.t2 514.134
R577 div120_0.div5_0.Q2_b.n3 div120_0.div5_0.Q2_b.n2 364.178
R578 div120_0.div5_0.Q2_b.n0 div120_0.div5_0.Q2_b.t11 353.467
R579 div120_0.div5_0.Q2_b.t6 div120_0.div5_0.Q2_b.n5 353.467
R580 div120_0.div5_0.Q2_b.n5 div120_0.div5_0.Q2_b.t4 289.2
R581 div120_0.div5_0.Q2_b.n4 div120_0.div5_0.Q2_b.n3 257.079
R582 div120_0.div5_0.Q2_b.t1 div120_0.div5_0.Q2_b.n7 233
R583 div120_0.div5_0.Q2_b.n6 div120_0.div5_0.Q2_b.t5 208.868
R584 div120_0.div5_0.Q2_b.n0 div120_0.div5_0.Q2_b.t8 192.8
R585 div120_0.div5_0.Q2_b.n2 div120_0.div5_0.Q2_b.n1 176.733
R586 div120_0.div5_0.Q2_b.n2 div120_0.div5_0.Q2_b.t9 112.468
R587 div120_0.div5_0.Q2_b.n1 div120_0.div5_0.Q2_b.t3 112.468
R588 div120_0.div5_0.Q2_b.n3 div120_0.div5_0.Q2_b.t7 112.468
R589 div120_0.div5_0.Q2_b.n5 div120_0.div5_0.Q2_b.t10 112.468
R590 div120_0.div5_0.Q2_b.n1 div120_0.div5_0.Q2_b.n0 96.4005
R591 div120_0.div5_0.Q2_b.n7 div120_0.div5_0.Q2_b.n4 21.3338
R592 a_938_228.n0 a_938_228.t1 289.967
R593 a_938_228.n0 a_938_228.t2 254.768
R594 a_938_228.t0 a_938_228.n0 161.701
R595 div120_0.div5_0.J.n0 div120_0.div5_0.J.t0 723.534
R596 div120_0.div5_0.J.n1 div120_0.div5_0.J.t4 553.534
R597 div120_0.div5_0.J.n0 div120_0.div5_0.J.t1 254.333
R598 div120_0.div5_0.J.n2 div120_0.div5_0.J.n1 206.333
R599 div120_0.div5_0.J.n1 div120_0.div5_0.J.n0 70.4005
R600 div120_0.div5_0.J.n2 div120_0.div5_0.J.t2 48.0005
R601 div120_0.div5_0.J.t3 div120_0.div5_0.J.n2 48.0005
R602 div120_0.div2_3_2.C.n0 div120_0.div2_3_2.C.t0 721.4
R603 div120_0.div2_3_2.C.n1 div120_0.div2_3_2.C.t4 349.433
R604 div120_0.div2_3_2.C.n0 div120_0.div2_3_2.C.t1 276.733
R605 div120_0.div2_3_2.C.n2 div120_0.div2_3_2.C.n1 206.333
R606 div120_0.div2_3_2.C.n1 div120_0.div2_3_2.C.n0 48.0005
R607 div120_0.div2_3_2.C.n2 div120_0.div2_3_2.C.t2 48.0005
R608 div120_0.div2_3_2.C.t3 div120_0.div2_3_2.C.n2 48.0005
R609 div120_0.div5_0.A.n2 div120_0.div5_0.A.t0 755.534
R610 div120_0.div5_0.A.t1 div120_0.div5_0.A.n2 685.134
R611 div120_0.div5_0.A.n1 div120_0.div5_0.A.n0 389.733
R612 div120_0.div5_0.A.n1 div120_0.div5_0.A.t2 340.2
R613 div120_0.div5_0.A.n0 div120_0.div5_0.A.t4 321.334
R614 div120_0.div5_0.A.n0 div120_0.div5_0.A.t3 144.601
R615 div120_0.div5_0.A.n2 div120_0.div5_0.A.n1 19.2005
R616 div120_0.div5_0.B.n0 div120_0.div5_0.B.t0 663.801
R617 div120_0.div5_0.B.n0 div120_0.div5_0.B.t2 380.368
R618 div120_0.div5_0.B div120_0.div5_0.B.t1 282.921
R619 div120_0.div5_0.B div120_0.div5_0.B.n0 114.133
R620 div120_0.div4.t4 div120_0.div4.t2 819.4
R621 div120_0.div4.n0 div120_0.div4.t1 663.801
R622 div120_0.div4.n0 div120_0.div4.t4 489.168
R623 div120_0.div4.t3 div120_0.div4.t5 401.668
R624 div120_0.div4.n1 div120_0.div4.t0 270.12
R625 div120_0.div4.n2 div120_0.div4.t3 257.067
R626 div120_0.div2_3_0.VIN div120_0.div4.n2 216.9
R627 div120_0.div4.n2 div120_0.div4.t6 208.868
R628 div120_0.div4.n3 div120_0.div2_3_0.VIN 192.167
R629 div120_0.div4.n1 div120_0.div4.n0 67.2005
R630 div120_0.div4.n3 div120_0.div4.n1 25.6005
R631 div120_0.div2_3_2.VOUT div120_0.div4.n3 4.8005
R632 div120_0.div2_3_2.B.t0 div120_0.div2_3_2.B.t1 96.0005
R633 div120_0.div2_3_0.CLK.n4 div120_0.div2_3_0.CLK.t0 723.534
R634 div120_0.div2_3_0.CLK.t1 div120_0.div2_3_0.CLK.n5 723.534
R635 div120_0.div2_3_0.CLK.n0 div120_0.div2_3_0.CLK.t6 369.534
R636 div120_0.div2_3_0.CLK.n3 div120_0.div2_3_0.CLK.n2 366.856
R637 div120_0.div2_3_0.CLK.n5 div120_0.div2_3_0.CLK.t2 254.333
R638 div120_0.div2_3_0.CLK.n3 div120_0.div2_3_0.CLK.t7 190.123
R639 div120_0.div2_3_0.CLK.n4 div120_0.div2_3_0.CLK.n3 187.201
R640 div120_0.div2_3_0.CLK.n1 div120_0.div2_3_0.CLK.n0 176.733
R641 div120_0.div2_3_0.CLK.n2 div120_0.div2_3_0.CLK.n1 176.733
R642 div120_0.div2_3_0.CLK.n0 div120_0.div2_3_0.CLK.t3 112.468
R643 div120_0.div2_3_0.CLK.n2 div120_0.div2_3_0.CLK.t4 112.468
R644 div120_0.div2_3_0.CLK.n1 div120_0.div2_3_0.CLK.t5 112.468
R645 div120_0.div2_3_0.CLK.n5 div120_0.div2_3_0.CLK.n4 70.4005
R646 div120_0.div2_3_0.C.n0 div120_0.div2_3_0.C.t3 721.4
R647 div120_0.div2_3_0.C.n1 div120_0.div2_3_0.C.t4 349.433
R648 div120_0.div2_3_0.C.n0 div120_0.div2_3_0.C.t1 276.733
R649 div120_0.div2_3_0.C.n2 div120_0.div2_3_0.C.n1 206.333
R650 div120_0.div2_3_0.C.n1 div120_0.div2_3_0.C.n0 48.0005
R651 div120_0.div2_3_0.C.t2 div120_0.div2_3_0.C.n2 48.0005
R652 div120_0.div2_3_0.C.n2 div120_0.div2_3_0.C.t0 48.0005
R653 div120_0.div5_0.L.t0 div120_0.div5_0.L.t1 96.0005
R654 div120_0.div2_3_1.C.n0 div120_0.div2_3_1.C.t0 721.4
R655 div120_0.div2_3_1.C.n1 div120_0.div2_3_1.C.t4 349.433
R656 div120_0.div2_3_1.C.n0 div120_0.div2_3_1.C.t2 276.733
R657 div120_0.div2_3_1.C.n2 div120_0.div2_3_1.C.n1 206.333
R658 div120_0.div2_3_1.C.n1 div120_0.div2_3_1.C.n0 48.0005
R659 div120_0.div2_3_1.C.t3 div120_0.div2_3_1.C.n2 48.0005
R660 div120_0.div2_3_1.C.n2 div120_0.div2_3_1.C.t1 48.0005
R661 div120_0.div3_2_0.G.t0 div120_0.div3_2_0.G.t1 96.0005
R662 div120_0.div5_0.D.n0 div120_0.div5_0.D.t0 761.4
R663 div120_0.div5_0.D.n1 div120_0.div5_0.D.t4 350.349
R664 div120_0.div5_0.D.n0 div120_0.div5_0.D.t1 254.333
R665 div120_0.div5_0.D.n2 div120_0.div5_0.D.n1 206.333
R666 div120_0.div5_0.D.n1 div120_0.div5_0.D.n0 70.4005
R667 div120_0.div5_0.D.n2 div120_0.div5_0.D.t2 48.0005
R668 div120_0.div5_0.D.t3 div120_0.div5_0.D.n2 48.0005
R669 div120_0.div3_2_0.B.t0 div120_0.div3_2_0.B.t1 96.0005
R670 div120_0.div2_3_2.A.n0 div120_0.div2_3_2.A.t0 713.933
R671 div120_0.div2_3_2.A.n0 div120_0.div2_3_2.A.t2 314.233
R672 div120_0.div2_3_2.A.t1 div120_0.div2_3_2.A.n0 308.2
R673 div120_0.div3_2_0.E.n0 div120_0.div3_2_0.E.t2 685.134
R674 div120_0.div3_2_0.E.n1 div120_0.div3_2_0.E.t1 663.801
R675 div120_0.div3_2_0.E.n0 div120_0.div3_2_0.E.t3 534.268
R676 div120_0.div3_2_0.E.t0 div120_0.div3_2_0.E.n1 362.921
R677 div120_0.div3_2_0.E.n1 div120_0.div3_2_0.E.n0 91.7338
R678 div120_0.div3_2_0.F.t0 div120_0.div3_2_0.F.t1 96.0005
R679 div120_0.div5_0.K.n0 div120_0.div5_0.K.t0 663.801
R680 div120_0.div5_0.K.t1 div120_0.div5_0.K.n0 397.053
R681 div120_0.div5_0.K.n0 div120_0.div5_0.K.t2 380.368
R682 div120_0.div8.t5 div120_0.div8.t4 819.4
R683 div120_0.div8.n0 div120_0.div8.t0 663.801
R684 div120_0.div8.n0 div120_0.div8.t5 489.168
R685 div120_0.div8.t2 div120_0.div8.t6 401.668
R686 div120_0.div8.n1 div120_0.div8.t1 270.12
R687 div120_0.div8.n2 div120_0.div8.t2 257.067
R688 div120_0.div3_2_0.VIN div120_0.div8.n2 216.9
R689 div120_0.div8.n2 div120_0.div8.t3 208.868
R690 div120_0.div8.n3 div120_0.div3_2_0.VIN 192.167
R691 div120_0.div8.n1 div120_0.div8.n0 67.2005
R692 div120_0.div8.n3 div120_0.div8.n1 25.6005
R693 div120_0.div2_3_0.VOUT div120_0.div8.n3 4.8005
R694 div120_0.div5_0.C.t0 div120_0.div5_0.C.t1 96.0005
R695 a_938_966.n0 a_938_966.t0 398.087
R696 a_938_966.t2 a_938_966.n0 349.767
R697 a_938_966.n0 a_938_966.t1 212.364
R698 a_1460_718.n1 a_1460_718.n0 791.453
R699 a_1460_718.t1 a_1460_718.n1 374.728
R700 a_1460_718.n1 a_1460_718.t0 271.567
R701 a_1460_718.n0 a_1460_718.t2 186.775
R702 a_1460_718.n0 a_1460_718.t3 115.981
R703 a_1492_966.n0 a_1492_966.t0 398.087
R704 a_1492_966.t2 a_1492_966.n0 349.767
R705 a_1492_966.n0 a_1492_966.t1 212.364
R706 a_906_718.n1 a_906_718.n0 785.028
R707 a_906_718.t0 a_906_718.n1 374.728
R708 a_906_718.n1 a_906_718.t1 271.567
R709 a_906_718.n0 a_906_718.t2 186.775
R710 a_906_718.n0 a_906_718.t3 115.981
R711 div120_0.div2_3_1.B.t0 div120_0.div2_3_1.B.t1 96.0005
R712 div120_0.div2_3_0.B.t0 div120_0.div2_3_0.B.t1 96.0005
R713 div120_0.div2_3_0.A.n0 div120_0.div2_3_0.A.t1 713.933
R714 div120_0.div2_3_0.A.n0 div120_0.div2_3_0.A.t2 314.233
R715 div120_0.div2_3_0.A.t0 div120_0.div2_3_0.A.n0 308.2
R716 div120_0.div2_3_1.A.n0 div120_0.div2_3_1.A.t1 713.933
R717 div120_0.div2_3_1.A.n0 div120_0.div2_3_1.A.t2 314.233
R718 div120_0.div2_3_1.A.t0 div120_0.div2_3_1.A.n0 308.2
C0 VDDA V_OUT120 0.659192f
C1 div120_0.div5_0.B VDDA 0.308332f
C2 VDDA V_CONT 0.065461f
C3 V_OUT120 GNDA 1.8905f
C4 V_CONT GNDA 1.55223f
C5 VDDA GNDA 20.72292f
C6 div120_0.div5_0.B GNDA 0.250854f
C7 VDDA.t83 GNDA 0.012818f
C8 VDDA.n0 GNDA 0.085326f
C9 VDDA.t45 GNDA 0.022708f
C10 VDDA.t13 GNDA 0.022708f
C11 VDDA.n7 GNDA 0.012721f
C12 VDDA.t86 GNDA 0.028814f
C13 VDDA.t90 GNDA 0.033012f
C14 VDDA.t17 GNDA 0.02786f
C15 VDDA.t59 GNDA 0.016792f
C16 VDDA.t62 GNDA 0.016792f
C17 VDDA.t36 GNDA 0.02557f
C18 VDDA.t64 GNDA 0.02557f
C19 VDDA.t29 GNDA 0.015075f
C20 VDDA.n10 GNDA 0.014581f
C21 VDDA.n13 GNDA 0.041037f
C22 VDDA.n15 GNDA 0.023889f
C23 VDDA.n17 GNDA 0.024979f
C24 VDDA.n18 GNDA 0.01472f
C25 VDDA.n20 GNDA 0.020981f
C26 VDDA.n22 GNDA 0.018255f
C27 VDDA.n23 GNDA 0.014515f
C28 VDDA.n26 GNDA 0.013348f
C29 VDDA.n28 GNDA 0.016074f
C30 VDDA.n31 GNDA 0.014575f
C31 VDDA.t19 GNDA 0.015075f
C32 VDDA.t33 GNDA 0.017174f
C33 VDDA.t25 GNDA 0.017174f
C34 VDDA.t88 GNDA 0.013739f
C35 VDDA.t4 GNDA 0.013739f
C36 VDDA.t49 GNDA 0.022135f
C37 VDDA.t70 GNDA 0.022135f
C38 VDDA.t55 GNDA 0.016792f
C39 VDDA.t6 GNDA 0.016792f
C40 VDDA.t57 GNDA 0.023662f
C41 VDDA.t68 GNDA 0.024616f
C42 VDDA.t31 GNDA 0.021753f
C43 VDDA.t10 GNDA 0.013739f
C44 VDDA.t2 GNDA 0.013739f
C45 VDDA.t74 GNDA 0.012022f
C46 VDDA.n32 GNDA 0.011522f
C47 VDDA.n36 GNDA 0.012985f
C48 VDDA.n38 GNDA 0.011713f
C49 VDDA.n41 GNDA 0.011713f
C50 VDDA.n43 GNDA 0.012985f
C51 VDDA.n46 GNDA 0.011522f
C52 VDDA.t66 GNDA 0.012022f
C53 VDDA.t72 GNDA 0.013739f
C54 VDDA.t8 GNDA 0.013739f
C55 VDDA.t92 GNDA 0.021753f
C56 VDDA.t60 GNDA 0.022708f
C57 VDDA.t0 GNDA 0.021753f
C58 VDDA.t38 GNDA 0.013739f
C59 VDDA.t84 GNDA 0.013739f
C60 VDDA.t53 GNDA 0.012022f
C61 VDDA.n47 GNDA 0.011522f
C62 VDDA.n51 GNDA 0.012985f
C63 VDDA.n53 GNDA 0.011713f
C64 VDDA.n55 GNDA 0.114508f
C65 VDDA.n57 GNDA 0.011713f
C66 VDDA.n59 GNDA 0.012985f
C67 VDDA.n62 GNDA 0.011522f
C68 VDDA.t15 GNDA 0.012022f
C69 VDDA.t21 GNDA 0.013739f
C70 VDDA.t43 GNDA 0.013739f
C71 VDDA.t40 GNDA 0.025125f
C72 VDDA.t47 GNDA 0.107419f
C73 VDDA.t82 GNDA 0.108338f
C74 VDDA.t23 GNDA 0.106966f
C75 VDDA.t78 GNDA 0.032521f
C76 VDDA.t80 GNDA 0.249588f
C77 VDDA.t76 GNDA 0.110101f
C78 VDDA.t27 GNDA 0.076013f
C79 VDDA.n63 GNDA 0.103644f
C80 VDDA.n64 GNDA 0.013211f
C81 VDDA.n65 GNDA 0.06061f
C82 VDDA.t79 GNDA 0.012818f
C83 VDDA.n66 GNDA 0.075885f
C84 VDDA.n67 GNDA 0.066142f
C85 VDDA.t77 GNDA 0.012818f
C86 VDDA.n68 GNDA 0.048337f
C87 VDDA.t81 GNDA 0.012818f
C88 VDDA.n69 GNDA 0.084261f
C89 a_110_1544.t2 GNDA 0.159497f
C90 a_110_1544.t3 GNDA 0.482598f
C91 a_110_1544.t4 GNDA 0.378972f
C92 a_110_1544.n0 GNDA 0.287213f
C93 a_110_1544.t5 GNDA 0.378972f
C94 a_110_1544.n1 GNDA 0.286839f
C95 a_110_1544.t1 GNDA 0.537461f
C96 a_110_1544.n2 GNDA 0.24614f
C97 a_110_1544.t0 GNDA 0.142309f
.ends

