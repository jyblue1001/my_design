* PEX produced on Mon Jun 30 03:14:22 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from two_stage_opamp_dummy_magic.ext - technology: sky130A

.subckt two_stage_opamp_dummy_magic VDDA V_CMFB_S1 V_CMFB_S3 Vb3 Vb2 Vb1 V_CMFB_S2
+ V_CMFB_S4 VOUT- VOUT+ V_tail_gate V_err_amp_ref V_err_gate VIN+ VIN- GNDA
X0 VOUT-.t19 cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1 VOUT-.t20 cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2 VOUT-.t21 cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 V_p.t34 V_tail_gate.t4 GNDA.t153 GNDA.t152 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X4 V_p.t33 V_tail_gate.t5 GNDA.t151 GNDA.t150 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X5 V_err_gate.t8 V_err_amp_ref.t0 V_err_mir_p.t12 VDDA.t233 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X6 VD4.t25 VDDA.t177 VDDA.t179 VDDA.t178 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X7 VDDA.t76 X.t25 VOUT-.t10 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X8 GNDA.t89 VDDA.t174 VDDA.t176 VDDA.t175 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X9 VOUT+.t19 cap_res_Y.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 VOUT+.t20 cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X11 VOUT+.t21 cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 err_amp_mir.t16 err_amp_mir.t15 GNDA.t66 GNDA.t65 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X13 VOUT+.t22 cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X14 VOUT-.t22 cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 VOUT-.t23 cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 VOUT-.t24 cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 VDDA.t109 Y.t25 V_CMFB_S4.t9 GNDA.t111 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X18 a_58940_5092.t1 V_CMFB_S2.t0 GNDA.t113 sky130_fd_pr__res_xhigh_po_0p35 l=4.07
X19 VOUT-.t25 cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 VD1.t20 Vb1.t2 Y.t22 GNDA.t243 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X21 Vb3.t7 Vb2.t3 Vb2_Vb3.t23 Vb2_Vb3.t22 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1 as=0.12 ps=1 w=0.6 l=0.2
X22 VDDA.t219 V_err_gate.t12 V_err_mir_p.t19 VDDA.t218 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X23 VDDA.t217 V_err_gate.t13 V_err_mir_p.t7 VDDA.t216 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X24 err_amp_mir.t4 V_tot.t4 V_err_p.t4 VDDA.t69 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X25 VOUT-.t26 cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X26 VOUT-.t27 cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 VOUT+.t23 cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X28 V_p.t36 VIN+.t0 VD2.t9 GNDA.t233 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X29 VOUT+.t24 cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 VOUT+.t25 cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 VDDA.t223 GNDA.t223 GNDA.t225 GNDA.t224 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X32 V_CMFB_S3.t10 Y.t26 GNDA.t70 VDDA.t65 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X33 VOUT+.t26 cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 VOUT+.t27 cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 VOUT+.t13 VDDA.t171 VDDA.t173 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X36 V_CMFB_S1.t10 X.t26 GNDA.t227 VDDA.t237 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X37 VOUT-.t28 cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 VOUT+.t28 cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 GNDA.t40 err_amp_mir.t13 err_amp_mir.t14 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X40 VDDA.t170 VDDA.t168 Vb2_Vb3.t11 VDDA.t169 sky130_fd_pr__pfet_01v8 ad=0.32 pd=2.4 as=0.16 ps=1.2 w=0.8 l=0.2
X41 VOUT+.t29 cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 VOUT+.t30 cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 VOUT-.t29 cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 V_err_p.t16 V_err_gate.t14 VDDA.t215 VDDA.t214 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X45 VOUT+.t31 cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 VOUT+.t32 cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 VOUT+.t33 cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X48 VOUT-.t30 cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 GNDA.t222 GNDA.t221 V_tail_gate.t0 GNDA.t102 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X50 VD1.t8 VIN-.t0 V_p.t12 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X51 Y.t24 VD4.t35 VD4.t37 VD4.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X52 VOUT+.t34 cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X53 VOUT+.t35 cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X54 V_err_gate.t7 V_err_amp_ref.t1 V_err_mir_p.t15 VDDA.t232 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X55 VOUT+.t36 cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X56 VOUT+.t37 cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X57 V_p.t32 V_tail_gate.t6 GNDA.t149 GNDA.t148 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X58 cap_res_Y.t0 Y.t2 GNDA.t7 sky130_fd_pr__res_high_po_1p41 l=1.41
X59 VDDA.t14 Y.t27 VOUT+.t0 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X60 X.t8 Vb1.t3 VD2.t21 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X61 VOUT+.t38 cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X62 VOUT-.t31 cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X63 VOUT+.t39 cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X64 VDDA.t46 X.t27 VOUT-.t5 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X65 Vb3.t6 Vb2.t4 Vb2_Vb3.t21 Vb2_Vb3.t20 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1 as=0.12 ps=1 w=0.6 l=0.2
X66 VOUT+.t40 cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 err_amp_out.t11 err_amp_mir.t17 GNDA.t107 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X68 VDDA.t39 Y.t28 V_CMFB_S4.t8 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X69 VOUT+.t41 cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X70 VOUT-.t32 cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X71 VDDA.t213 V_err_gate.t15 V_err_mir_p.t1 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X72 VOUT-.t33 cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X73 VOUT+.t42 cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 GNDA.t220 GNDA.t218 VOUT-.t9 GNDA.t219 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X75 a_59060_4632.t0 V_CMFB_S1.t0 GNDA.t10 sky130_fd_pr__res_xhigh_po_0p35 l=1.77
X76 VOUT-.t34 cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X77 VD4.t31 Vb3.t8 VDDA.t255 VDDA.t254 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X78 VD1.t19 Vb1.t4 Y.t17 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X79 VDDA.t211 V_err_gate.t16 V_err_p.t15 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X80 VOUT+.t43 cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X81 VOUT-.t35 cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X82 err_amp_out.t6 V_err_amp_ref.t2 V_err_p.t17 VDDA.t231 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X83 VOUT-.t36 cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 VOUT+.t44 cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 GNDA.t147 V_tail_gate.t7 V_p.t31 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X86 V_CMFB_S3.t9 Y.t29 GNDA.t20 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X87 VOUT-.t37 cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 VDDA.t167 VDDA.t165 GNDA.t63 VDDA.t166 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X89 V_CMFB_S1.t9 X.t28 GNDA.t230 VDDA.t240 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X90 GNDA.t87 err_amp_mir.t18 err_amp_out.t10 GNDA.t86 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X91 V_CMFB_S2.t10 X.t29 VDDA.t90 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X92 VDDA.t85 Vb3.t9 VD3.t15 VDDA.t84 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X93 GNDA.t217 GNDA.t215 VDDA.t222 GNDA.t216 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X94 VOUT+.t45 cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 VOUT-.t38 cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X96 VOUT+.t46 cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 V_err_mir_p.t3 V_err_gate.t17 VDDA.t209 VDDA.t208 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X98 VOUT+.t47 cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X99 VOUT-.t39 cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 VOUT+.t48 cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X101 V_err_p.t18 V_err_amp_ref.t3 err_amp_out.t5 VDDA.t230 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X102 V_p_mir.t0 VIN-.t1 V_tail_gate.t1 GNDA.t109 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X103 VD2.t8 VIN+.t1 V_p.t14 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X104 VOUT+.t49 cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 VOUT+.t10 V_b_2nd_stage.t2 GNDA.t98 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X106 VDDA.t55 Vb3.t10 VD4.t12 VDDA.t54 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X107 V_err_gate.t3 V_tot.t5 V_err_mir_p.t9 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X108 V_p.t30 V_tail_gate.t8 GNDA.t145 GNDA.t144 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X109 Vb2_Vb3.t10 VDDA.t162 VDDA.t164 VDDA.t163 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.2 as=0.32 ps=2.4 w=0.8 l=0.2
X110 VDDA.t30 Y.t30 VOUT+.t4 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X111 VDDA.t161 VDDA.t159 VOUT+.t12 VDDA.t160 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X112 X.t10 Vb1.t5 VD2.t20 GNDA.t72 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X113 VDDA.t97 X.t30 VOUT-.t16 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X114 VOUT-.t40 cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 Y.t5 Vb2.t5 VD4.t4 VD4.t3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X116 VOUT-.t41 cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X117 VOUT-.t42 cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X118 VOUT-.t43 cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 VOUT+.t50 cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 VDDA.t18 Y.t31 V_CMFB_S4.t7 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X121 VDDA.t203 V_err_gate.t18 V_err_p.t14 VDDA.t202 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X122 VOUT+.t51 cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 VOUT-.t44 cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 VOUT-.t17 GNDA.t212 GNDA.t214 GNDA.t213 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X125 err_amp_mir.t5 VDDA.t156 VDDA.t158 VDDA.t157 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X126 VOUT-.t45 cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X127 VOUT-.t46 cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 GNDA.t143 V_tail_gate.t9 V_p.t29 GNDA.t142 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X129 GNDA.t141 V_tail_gate.t10 V_p.t28 GNDA.t140 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X130 VD3.t37 Vb2.t6 X.t14 VD3.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X131 VOUT-.t47 cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X132 V_CMFB_S3.t8 Y.t32 GNDA.t44 VDDA.t40 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X133 VOUT-.t48 cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 VOUT-.t49 cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X135 VOUT-.t50 cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X136 V_CMFB_S2.t9 X.t31 VDDA.t101 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X137 VOUT-.t51 cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 VOUT+.t52 cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 VOUT-.t4 V_b_2nd_stage.t3 GNDA.t38 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X140 VDDA.t242 Vb3.t11 VD4.t26 VDDA.t241 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X141 VD3.t17 VDDA.t153 VDDA.t155 VDDA.t154 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X142 VD4.t18 Vb2.t7 Y.t15 VD4.t17 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X143 VD2.t7 VIN+.t2 V_p.t13 GNDA.t90 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X144 V_err_p.t3 V_tot.t6 err_amp_mir.t0 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X145 VD1.t1 VIN-.t2 V_p.t1 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X146 VOUT-.t52 cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 Vb2_Vb3.t19 Vb2.t8 Vb3.t5 Vb2_Vb3.t18 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1 as=0.12 ps=1 w=0.6 l=0.2
X148 V_err_gate.t6 V_err_amp_ref.t4 V_err_mir_p.t11 VDDA.t229 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X149 X.t6 Vb1.t6 VD2.t19 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X150 VOUT-.t8 V_b_2nd_stage.t4 GNDA.t78 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X151 VOUT-.t53 cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 VDDA.t235 Y.t33 VOUT+.t16 VDDA.t234 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X153 X.t23 Vb1.t7 VD2.t18 GNDA.t237 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X154 VOUT+.t53 cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X155 VOUT+.t54 cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X156 VOUT-.t54 cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 VOUT+.t55 cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 VOUT+.t56 cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 VDDA.t98 Y.t34 V_CMFB_S4.t6 GNDA.t101 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X160 VOUT-.t55 cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X161 VDDA.t87 Vb3.t12 VD4.t14 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X162 VOUT+.t57 cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X163 GNDA.t30 V_b_2nd_stage.t5 VOUT+.t3 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X164 VOUT-.t56 cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 VOUT-.t57 cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 VOUT+.t58 cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X167 VOUT-.t58 cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X168 VOUT-.t59 cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X169 GNDA.t139 V_tail_gate.t11 V_p.t27 GNDA.t138 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X170 VOUT-.t60 cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 Vb2.t2 Vb2.t1 VDDA.t103 VDDA.t102 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.03 as=0.126 ps=1.03 w=0.63 l=0.2
X172 VOUT-.t61 cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X173 V_b_2nd_stage.t1 a_67950_1836.t0 GNDA.t100 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X174 VD3.t14 Vb3.t13 VDDA.t52 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X175 VOUT+.t59 cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 VOUT-.t62 cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 V_CMFB_S3.t7 Y.t35 GNDA.t22 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X178 VOUT-.t63 cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X179 VOUT-.t64 cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X180 GNDA.t103 err_amp_mir.t11 err_amp_mir.t12 GNDA.t102 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X181 VD4.t23 Vb2.t9 Y.t18 VD4.t22 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X182 GNDA.t211 GNDA.t209 err_amp_out.t1 GNDA.t210 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X183 X.t4 VD3.t3 VD3.t5 VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X184 VOUT+.t60 cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 GNDA.t61 V_b_2nd_stage.t6 VOUT+.t6 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X186 V_CMFB_S2.t8 X.t32 VDDA.t80 GNDA.t82 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X187 Y.t20 GNDA.t206 GNDA.t208 GNDA.t207 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X188 Y.t12 Vb1.t8 VD1.t18 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X189 V_err_p.t13 V_err_gate.t19 VDDA.t207 VDDA.t206 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X190 Y.t13 Vb1.t9 VD1.t17 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X191 VOUT+.t61 cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 VOUT-.t65 cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X193 VOUT+.t62 cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X194 VD1.t5 VIN-.t3 V_p.t5 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X195 VD4.t7 Vb3.t14 VDDA.t48 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X196 VOUT-.t66 cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 VDDA.t152 VDDA.t150 err_amp_out.t0 VDDA.t151 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X198 VOUT+.t63 cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 VD1.t6 VIN-.t4 V_p.t7 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X200 VD2.t6 VIN+.t3 V_p.t8 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X201 VOUT-.t67 cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 VOUT+.t64 cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X203 V_p_mir.t3 V_tail_gate.t12 GNDA.t137 GNDA.t136 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X204 V_err_gate.t9 VDDA.t143 VDDA.t145 VDDA.t144 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X205 VOUT+.t65 cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X206 VOUT-.t68 cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 V_err_gate.t2 V_tot.t7 V_err_mir_p.t8 VDDA.t104 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X208 VD3.t13 Vb3.t15 VDDA.t44 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X209 X.t5 Vb1.t10 VD2.t17 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X210 GNDA.t81 X.t33 V_CMFB_S1.t8 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X211 VOUT-.t69 cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 VOUT+.t66 cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 VOUT+.t67 cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X214 VDDA.t26 Y.t36 VOUT+.t1 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X215 VD4.t9 Vb2.t10 Y.t7 VD4.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X216 VDDA.t221 GNDA.t203 GNDA.t205 GNDA.t204 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X217 VOUT+.t68 cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X218 VOUT-.t70 cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X219 VOUT-.t71 cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X220 VOUT-.t72 cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X221 GNDA.t202 GNDA.t200 GNDA.t202 GNDA.t201 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0 ps=0 w=1 l=0.15
X222 V_p.t4 VIN-.t5 VD1.t4 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X223 VDDA.t205 V_err_gate.t20 V_err_p.t12 VDDA.t204 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X224 VOUT-.t73 cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X225 VOUT+.t69 cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X226 VOUT+.t70 cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X227 VOUT+.t71 cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X228 GNDA.t135 V_tail_gate.t13 V_p.t26 GNDA.t134 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X229 X.t3 Vb2.t11 VD3.t35 VD3.t34 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X230 VOUT-.t74 cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X231 GNDA.t133 V_tail_gate.t14 V_p.t25 GNDA.t132 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X232 VOUT-.t14 X.t34 VDDA.t94 VDDA.t93 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X233 VOUT-.t75 cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X234 VOUT-.t76 cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X235 VDDA.t149 VDDA.t146 VDDA.t148 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.06 as=0 ps=0 w=0.63 l=0.2
X236 VD4.t30 Vb3.t16 VDDA.t253 VDDA.t252 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X237 V_CMFB_S4.t5 Y.t37 VDDA.t42 GNDA.t50 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X238 V_CMFB_S2.t7 X.t35 VDDA.t73 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X239 VOUT-.t77 cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 VOUT-.t78 cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 Y.t16 Vb2.t12 VD4.t20 VD4.t19 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X242 VOUT+.t72 cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X243 VOUT-.t79 cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 VOUT+.t73 cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 VOUT+.t74 cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 V_err_mir_p.t0 V_err_gate.t21 VDDA.t201 VDDA.t200 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X247 VOUT-.t80 cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X248 Y.t10 Vb1.t11 VD1.t16 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X249 VOUT+.t75 cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 VD2.t11 GNDA.t197 GNDA.t199 GNDA.t198 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X251 V_err_p.t2 V_tot.t8 err_amp_mir.t3 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X252 VOUT-.t81 cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 VD2.t5 VIN+.t4 V_p.t40 GNDA.t246 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X254 X.t22 Vb2.t13 VD3.t33 VD3.t32 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X255 VOUT-.t82 cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 VDDA.t61 Vb3.t17 Vb2_Vb3.t7 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.2 as=0.16 ps=1.2 w=0.8 l=0.2
X257 VOUT+.t76 cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 GNDA.t23 X.t36 V_CMFB_S1.t7 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X259 X.t21 GNDA.t194 GNDA.t196 GNDA.t195 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X260 VOUT-.t83 cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X261 VD4.t13 Vb3.t18 VDDA.t59 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X262 VOUT-.t84 cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 a_68230_5092.t0 V_CMFB_S4.t10 GNDA.t234 sky130_fd_pr__res_xhigh_po_0p35 l=4.07
X264 VOUT+.t77 cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 VOUT+.t78 cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 VOUT+.t79 cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X267 VOUT+.t80 cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X268 VOUT-.t85 cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 VOUT+.t81 cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X270 VOUT+.t82 cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 V_p.t35 GNDA.t191 GNDA.t193 GNDA.t192 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X272 VDDA.t142 VDDA.t140 Vb2.t0 VDDA.t141 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.06 as=0.126 ps=1.03 w=0.63 l=0.2
X273 a_58940_5092.t0 V_tot.t2 GNDA.t84 sky130_fd_pr__res_xhigh_po_0p35 l=4.07
X274 GNDA.t131 V_tail_gate.t15 V_p.t24 GNDA.t130 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X275 VDDA.t244 Vb3.t19 VD3.t12 VDDA.t243 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X276 VOUT-.t86 cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 VOUT+.t83 cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X278 VDDA.t139 VDDA.t137 V_err_gate.t10 VDDA.t138 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X279 Y.t14 Vb2.t14 VD4.t16 VD4.t15 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X280 VOUT-.t1 X.t37 VDDA.t6 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X281 V_CMFB_S3.t6 Y.t38 GNDA.t21 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X282 V_p.t37 Vb1.t0 Vb1.t1 GNDA.t235 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=2.3
X283 VOUT-.t87 cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 VOUT+.t84 cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X285 VOUT-.t88 cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 VOUT+.t85 cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X287 VOUT+.t86 cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X288 VOUT-.t89 cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X289 GNDA.t42 err_amp_mir.t9 err_amp_mir.t10 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X290 V_CMFB_S4.t4 Y.t39 VDDA.t64 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X291 VOUT-.t90 cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 GNDA.t190 GNDA.t188 VDDA.t220 GNDA.t189 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X293 V_CMFB_S2.t6 X.t38 VDDA.t238 GNDA.t228 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X294 VOUT+.t87 cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 V_err_p.t11 V_err_gate.t22 VDDA.t199 VDDA.t198 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X296 Y.t8 Vb1.t12 VD1.t15 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X297 V_err_p.t10 V_err_gate.t23 VDDA.t197 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X298 VOUT+.t88 cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X299 VOUT+.t89 cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 VD1.t21 VIN-.t6 V_p.t39 GNDA.t240 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X301 VDDA.t248 Vb3.t20 VD3.t11 VDDA.t247 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X302 VOUT-.t91 cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 Y.t0 Vb2.t15 VD4.t1 VD4.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X304 VDDA.t63 Y.t40 VOUT+.t7 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X305 GNDA.t229 X.t39 V_CMFB_S1.t6 VDDA.t239 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X306 VOUT-.t92 cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X307 err_amp_out.t9 err_amp_mir.t19 GNDA.t14 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X308 VOUT+.t90 cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 cap_res_X.t0 X.t1 GNDA.t2 sky130_fd_pr__res_high_po_1p41 l=1.41
X310 VOUT+.t91 cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X311 VOUT+.t92 cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X312 VD1.t14 Vb1.t13 Y.t9 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X313 VDDA.t136 VDDA.t134 V_err_p.t6 VDDA.t135 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X314 GNDA.t187 GNDA.t185 VD1.t10 GNDA.t186 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X315 VD3.t31 Vb2.t16 X.t19 VD3.t30 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X316 VOUT-.t93 cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 VOUT+.t93 cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 VOUT-.t94 cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 VOUT+.t94 cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 GNDA.t129 V_tail_gate.t16 V_p_mir.t2 GNDA.t128 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X321 V_err_mir_p.t13 V_err_amp_ref.t5 V_err_gate.t5 VDDA.t228 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X322 VOUT-.t95 cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 GNDA.t127 V_tail_gate.t17 V_p.t23 GNDA.t126 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X324 VOUT-.t96 cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X325 V_err_mir_p.t4 V_tot.t9 V_err_gate.t0 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X326 VDDA.t251 Vb3.t21 VD4.t29 VDDA.t250 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X327 GNDA.t184 GNDA.t182 X.t20 GNDA.t183 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X328 VOUT-.t97 cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X329 VOUT-.t11 X.t40 VDDA.t79 VDDA.t78 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X330 VOUT-.t98 cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X331 GNDA.t105 err_amp_mir.t20 err_amp_out.t8 GNDA.t104 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X332 V_b_2nd_stage.t0 a_59460_1836.t0 GNDA.t33 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X333 V_CMFB_S4.t3 Y.t41 VDDA.t110 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X334 VDDA.t133 VDDA.t131 VD3.t16 VDDA.t132 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X335 Y.t3 Vb1.t14 VD1.t13 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X336 V_err_mir_p.t17 V_err_gate.t24 VDDA.t195 VDDA.t194 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X337 VD3.t29 Vb2.t17 X.t16 VD3.t28 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X338 VOUT+.t95 cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X339 VOUT+.t96 cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X340 VOUT-.t99 cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X341 VOUT-.t100 cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X342 VOUT-.t101 cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X343 V_err_p.t21 V_err_amp_ref.t6 err_amp_out.t4 VDDA.t227 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X344 Vb2_Vb3.t8 Vb3.t22 VDDA.t67 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.2 as=0.16 ps=1.2 w=0.8 l=0.2
X345 VOUT-.t102 cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X346 V_p.t22 V_tail_gate.t18 GNDA.t123 GNDA.t122 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X347 VD2.t10 GNDA.t179 GNDA.t181 GNDA.t180 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X348 VOUT+.t97 cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X349 VOUT-.t103 cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 VDDA.t130 VDDA.t128 VD4.t24 VDDA.t129 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X351 GNDA.t25 Y.t42 V_CMFB_S3.t5 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X352 a_68350_4632.t1 V_CMFB_S3.t0 GNDA.t94 sky130_fd_pr__res_xhigh_po_0p35 l=1.77
X353 GNDA.t3 X.t41 V_CMFB_S1.t5 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X354 VOUT-.t104 cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X355 VOUT+.t98 cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X356 VOUT+.t99 cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X357 err_amp_mir.t8 err_amp_mir.t7 GNDA.t232 GNDA.t231 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X358 GNDA.t80 X.t42 V_CMFB_S1.t4 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X359 VOUT-.t105 cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X360 VOUT-.t106 cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X361 VOUT+.t100 cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X362 VDDA.t193 V_err_gate.t25 V_err_mir_p.t10 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X363 VOUT-.t107 cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 VOUT-.t108 cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X365 VOUT+.t101 cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X366 VOUT-.t109 cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X367 V_tail_gate.t3 VIN+.t5 V_p_mir.t1 GNDA.t162 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X368 V_p.t11 VIN+.t6 VD2.t4 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X369 VD3.t10 Vb3.t23 VDDA.t32 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X370 VD4.t11 Vb2.t18 Y.t11 VD4.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X371 VOUT+.t102 cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 V_err_mir_p.t6 V_tot.t10 V_err_gate.t1 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X373 VOUT+.t103 cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X374 GNDA.t125 V_tail_gate.t19 V_p.t21 GNDA.t124 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X375 VOUT+.t8 Y.t43 VDDA.t71 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X376 VD2.t16 Vb1.t15 X.t13 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X377 VOUT-.t110 cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X378 VOUT-.t18 X.t43 VDDA.t258 VDDA.t257 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X379 VOUT+.t104 cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X380 VOUT-.t6 X.t44 VDDA.t57 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X381 VD3.t2 VD3.t0 X.t17 VD3.t1 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X382 VOUT-.t111 cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 VOUT-.t112 cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X384 V_CMFB_S4.t2 Y.t44 VDDA.t33 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X385 VOUT-.t113 cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X386 VOUT+.t105 cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X387 VOUT+.t106 cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 V_err_mir_p.t2 V_err_gate.t26 VDDA.t191 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X389 VOUT-.t114 cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X390 VOUT-.t115 cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X391 VOUT+.t107 cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X392 VD3.t9 Vb3.t24 VDDA.t24 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X393 V_err_p.t1 V_tot.t11 err_amp_mir.t1 VDDA.t50 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X394 VOUT-.t116 cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X395 VD4.t34 VD4.t32 Y.t23 VD4.t33 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X396 VOUT-.t117 cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X397 V_p.t20 V_tail_gate.t20 GNDA.t121 GNDA.t120 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X398 VOUT-.t118 cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 GNDA.t178 GNDA.t176 GNDA.t178 GNDA.t177 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0 ps=0 w=2.5 l=0.15
X400 VOUT+.t108 cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 GNDA.t245 Y.t45 V_CMFB_S3.t4 VDDA.t256 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X402 GNDA.t175 GNDA.t173 VOUT+.t15 GNDA.t174 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X403 VOUT-.t119 cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 err_amp_out.t7 err_amp_mir.t21 GNDA.t57 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X405 VOUT-.t120 cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 VDDA.t1 X.t45 V_CMFB_S2.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X407 VD3.t8 Vb3.t25 VDDA.t8 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X408 VOUT+.t109 cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X409 VOUT-.t121 cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 VOUT-.t122 cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 X.t18 Vb2.t19 VD3.t27 VD3.t26 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X412 VOUT+.t110 cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X413 VOUT+.t111 cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 VOUT-.t123 cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X415 VOUT+.t112 cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 VDDA.t183 V_err_gate.t27 V_err_p.t9 VDDA.t182 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X417 V_p.t15 VIN+.t7 VD2.t3 GNDA.t92 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X418 err_amp_out.t3 V_err_amp_ref.t7 V_err_p.t19 VDDA.t226 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X419 V_tail_gate.t2 GNDA.t158 GNDA.t160 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X420 GNDA.t236 VDDA.t125 VDDA.t127 VDDA.t126 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X421 VOUT+.t113 cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X422 GNDA.t172 GNDA.t170 VD1.t9 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X423 VD4.t2 Vb3.t26 VDDA.t17 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X424 VOUT+.t114 cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X425 Vb3.t1 Vb2_Vb3.t4 Vb2_Vb3.t6 Vb2_Vb3.t5 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1 as=0.24 ps=2 w=0.6 l=0.2
X426 VOUT+.t115 cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 V_err_mir_p.t14 V_err_amp_ref.t8 V_err_gate.t4 VDDA.t225 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X428 VOUT-.t124 cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X429 GNDA.t36 V_b_2nd_stage.t7 VOUT-.t3 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X430 VD2.t15 Vb1.t16 X.t24 GNDA.t247 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X431 VOUT-.t15 a_59460_1836.t1 GNDA.t96 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X432 VOUT+.t9 Y.t46 VDDA.t89 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X433 VOUT+.t116 cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 VOUT+.t117 cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 VOUT+.t118 cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 VOUT-.t125 cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 VOUT+.t119 cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 VOUT-.t126 cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 VOUT+.t120 cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 VOUT+.t121 cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 VOUT+.t122 cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X442 X.t12 Vb2.t20 VD3.t25 VD3.t24 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X443 V_err_p.t5 VDDA.t122 VDDA.t124 VDDA.t123 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X444 VOUT+.t123 cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 VDDA.t37 Vb3.t27 Vb2_Vb3.t0 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.2 as=0.16 ps=1.2 w=0.8 l=0.2
X446 GNDA.t76 V_b_2nd_stage.t8 VOUT-.t7 GNDA.t75 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X447 VOUT-.t12 VDDA.t119 VDDA.t121 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X448 VOUT-.t127 cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X449 a_68350_4632.t0 V_tot.t1 GNDA.t69 sky130_fd_pr__res_xhigh_po_0p35 l=1.77
X450 Vb3.t4 Vb2.t21 Vb2_Vb3.t17 Vb2_Vb3.t16 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1 as=0.12 ps=1 w=0.6 l=0.2
X451 V_p.t19 V_tail_gate.t21 GNDA.t119 GNDA.t118 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X452 VOUT-.t128 cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X453 X.t2 Vb2.t22 VD3.t23 VD3.t22 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X454 VOUT+.t124 cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X455 VOUT+.t125 cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 GNDA.t45 Y.t47 V_CMFB_S3.t3 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X457 VOUT-.t129 cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X458 VOUT+.t126 cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 VOUT+.t127 cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 VOUT+.t128 cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 VOUT+.t14 GNDA.t167 GNDA.t169 GNDA.t168 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X462 VDDA.t12 X.t46 V_CMFB_S2.t4 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X463 VOUT+.t129 cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X464 VOUT-.t130 cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X465 VDDA.t83 Vb3.t28 VD3.t7 VDDA.t82 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X466 GNDA.t166 GNDA.t164 Y.t19 GNDA.t165 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X467 Y.t21 Vb2.t23 VD4.t28 VD4.t27 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X468 VOUT+.t130 cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X469 V_p.t10 VIN-.t7 VD1.t7 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X470 V_p.t0 VIN-.t8 VD1.t0 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X471 VOUT-.t131 cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 VOUT+.t131 cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X473 VOUT+.t132 cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 V_p.t9 VIN+.t8 VD2.t2 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X475 VOUT-.t132 cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X476 VOUT+.t133 cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X477 VOUT+.t2 V_b_2nd_stage.t9 GNDA.t28 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X478 V_err_mir_p.t18 V_tot.t12 V_err_gate.t11 VDDA.t249 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X479 V_CMFB_S1.t3 X.t47 GNDA.t5 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X480 VD2.t14 Vb1.t17 X.t0 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X481 VOUT+.t134 cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 VOUT-.t133 cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 VOUT+.t135 cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X484 VOUT+.t136 cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X485 VOUT+.t18 a_67950_1836.t1 GNDA.t242 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X486 VOUT+.t5 Y.t48 VDDA.t35 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X487 VDDA.t118 VDDA.t116 GNDA.t244 VDDA.t117 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X488 VD2.t13 Vb1.t18 X.t15 GNDA.t88 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X489 VOUT+.t137 cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 V_CMFB_S4.t1 Y.t49 VDDA.t259 GNDA.t248 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X491 V_err_mir_p.t16 V_err_gate.t28 VDDA.t189 VDDA.t188 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X492 VOUT+.t138 cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 VOUT+.t139 cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X494 VOUT-.t134 cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X495 VOUT+.t140 cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X496 VOUT-.t135 cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X497 VOUT+.t141 cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 V_p.t18 V_tail_gate.t22 GNDA.t117 GNDA.t116 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X499 VDDA.t3 X.t48 VOUT-.t0 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X500 VOUT+.t142 cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X501 VDDA.t115 VDDA.t113 VOUT-.t13 VDDA.t114 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X502 VDDA.t100 Vb3.t29 VD3.t6 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X503 err_amp_mir.t6 GNDA.t161 GNDA.t163 GNDA.t162 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X504 GNDA.t110 Y.t50 V_CMFB_S3.t2 VDDA.t108 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X505 VD3.t21 Vb2.t24 X.t9 VD3.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X506 VDDA.t260 X.t49 V_CMFB_S2.t3 GNDA.t249 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X507 VOUT-.t136 cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X508 VOUT+.t143 cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X509 VOUT-.t137 cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 VOUT+.t144 cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 VDDA.t187 V_err_gate.t29 V_err_mir_p.t5 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X512 VOUT-.t138 cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X513 VOUT-.t139 cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X514 VD1.t12 Vb1.t19 Y.t1 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X515 VDDA.t107 Vb3.t30 VD4.t21 VDDA.t106 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X516 VOUT-.t140 cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X517 V_p.t16 VIN+.t9 VD2.t1 GNDA.t95 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X518 err_amp_out.t2 V_err_amp_ref.t9 V_err_p.t20 VDDA.t224 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X519 V_p.t6 VIN+.t10 VD2.t0 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X520 Vb2_Vb3.t15 Vb2.t25 Vb3.t3 Vb2_Vb3.t14 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1 as=0.12 ps=1 w=0.6 l=0.2
X521 GNDA.t157 GNDA.t154 GNDA.t156 GNDA.t155 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X522 V_CMFB_S1.t2 X.t50 GNDA.t226 VDDA.t236 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X523 VD2.t12 Vb1.t20 X.t7 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X524 VOUT+.t17 Y.t51 VDDA.t246 VDDA.t245 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X525 VOUT-.t141 cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X526 Vb2_Vb3.t9 Vb3.t31 VDDA.t92 VDDA.t91 sky130_fd_pr__pfet_01v8 ad=0.16 pd=1.2 as=0.16 ps=1.2 w=0.8 l=0.2
X527 VOUT-.t142 cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 GNDA.t239 err_amp_out.t12 V_p.t38 GNDA.t238 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X529 VD1.t3 VIN-.t9 V_p.t3 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X530 V_err_p.t8 V_err_gate.t30 VDDA.t185 VDDA.t184 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X531 VOUT+.t145 cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 Vb2_Vb3.t3 Vb2_Vb3.t1 Vb3.t0 Vb2_Vb3.t2 sky130_fd_pr__pfet_01v8 ad=0.24 pd=2 as=0.12 ps=1 w=0.6 l=0.2
X533 a_68230_5092.t1 V_tot.t3 GNDA.t241 sky130_fd_pr__res_xhigh_po_0p35 l=4.07
X534 VD3.t19 Vb2.t26 X.t11 VD3.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X535 V_p.t17 V_tail_gate.t23 GNDA.t115 GNDA.t114 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X536 VOUT+.t146 cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X537 VOUT-.t143 cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X538 VDDA.t10 X.t51 VOUT-.t2 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X539 GNDA.t26 Y.t52 V_CMFB_S3.t1 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X540 VOUT-.t144 cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X541 VOUT-.t145 cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X542 VDDA.t15 Y.t53 V_CMFB_S4.t0 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X543 Vb2_Vb3.t13 Vb2.t27 Vb3.t2 Vb2_Vb3.t12 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1 as=0.12 ps=1 w=0.6 l=0.2
X544 VDDA.t81 X.t52 V_CMFB_S2.t2 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X545 VOUT+.t147 cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X546 VOUT+.t148 cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 VDDA.t95 X.t53 V_CMFB_S2.t1 GNDA.t99 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X548 VOUT-.t146 cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X549 VOUT-.t147 cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X550 VOUT-.t148 cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X551 VD4.t6 Vb2.t28 Y.t6 VD4.t5 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X552 VOUT-.t149 cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X553 VOUT+.t149 cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X554 VDDA.t181 V_err_gate.t31 V_err_p.t7 VDDA.t180 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X555 VOUT+.t150 cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X556 VD1.t11 Vb1.t21 Y.t4 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X557 err_amp_mir.t2 V_tot.t13 V_err_p.t0 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X558 a_59060_4632.t1 V_tot.t0 GNDA.t18 sky130_fd_pr__res_xhigh_po_0p35 l=1.77
X559 V_p.t2 VIN-.t10 VD1.t2 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X560 VOUT-.t150 cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 VOUT-.t151 cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X562 VOUT+.t151 cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X563 V_CMFB_S1.t1 X.t54 GNDA.t8 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X564 VOUT-.t152 cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X565 VOUT+.t11 Y.t54 VDDA.t112 VDDA.t111 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X566 VOUT+.t152 cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X567 VOUT+.t153 cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X568 VOUT-.t153 cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X569 VOUT-.t154 cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 VOUT-.t155 cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X571 VOUT+.t154 cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X572 VOUT-.t156 cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X573 VOUT+.t155 cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X574 VOUT+.t156 cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 VOUT-.n14 VOUT-.n6 145.989
R1 VOUT-.n9 VOUT-.n7 145.989
R2 VOUT-.n13 VOUT-.n12 145.427
R3 VOUT-.n11 VOUT-.n10 145.427
R4 VOUT-.n9 VOUT-.n8 145.427
R5 VOUT-.n16 VOUT-.n15 140.927
R6 VOUT-.n5 VOUT-.t15 113.192
R7 VOUT-.n2 VOUT-.n0 95.7303
R8 VOUT-.n4 VOUT-.n3 94.6053
R9 VOUT-.n2 VOUT-.n1 94.6053
R10 VOUT-.n100 VOUT-.n16 20.5943
R11 VOUT-.n100 VOUT-.n99 11.7059
R12 VOUT- VOUT-.n100 7.813
R13 VOUT-.n15 VOUT-.t0 6.56717
R14 VOUT-.n15 VOUT-.t14 6.56717
R15 VOUT-.n12 VOUT-.t2 6.56717
R16 VOUT-.n12 VOUT-.t1 6.56717
R17 VOUT-.n10 VOUT-.t10 6.56717
R18 VOUT-.n10 VOUT-.t11 6.56717
R19 VOUT-.n8 VOUT-.t5 6.56717
R20 VOUT-.n8 VOUT-.t18 6.56717
R21 VOUT-.n7 VOUT-.t16 6.56717
R22 VOUT-.n7 VOUT-.t12 6.56717
R23 VOUT-.n6 VOUT-.t13 6.56717
R24 VOUT-.n6 VOUT-.t6 6.56717
R25 VOUT-.n46 VOUT-.t74 4.8295
R26 VOUT-.n48 VOUT-.t80 4.8295
R27 VOUT-.n51 VOUT-.t114 4.8295
R28 VOUT-.n54 VOUT-.t22 4.8295
R29 VOUT-.n57 VOUT-.t123 4.8295
R30 VOUT-.n70 VOUT-.t31 4.8295
R31 VOUT-.n72 VOUT-.t89 4.8295
R32 VOUT-.n73 VOUT-.t70 4.8295
R33 VOUT-.n75 VOUT-.t125 4.8295
R34 VOUT-.n76 VOUT-.t106 4.8295
R35 VOUT-.n78 VOUT-.t85 4.8295
R36 VOUT-.n79 VOUT-.t65 4.8295
R37 VOUT-.n81 VOUT-.t39 4.8295
R38 VOUT-.n82 VOUT-.t27 4.8295
R39 VOUT-.n84 VOUT-.t79 4.8295
R40 VOUT-.n85 VOUT-.t57 4.8295
R41 VOUT-.n87 VOUT-.t35 4.8295
R42 VOUT-.n88 VOUT-.t21 4.8295
R43 VOUT-.n90 VOUT-.t135 4.8295
R44 VOUT-.n91 VOUT-.t124 4.8295
R45 VOUT-.n93 VOUT-.t96 4.8295
R46 VOUT-.n94 VOUT-.t84 4.8295
R47 VOUT-.n17 VOUT-.t121 4.8295
R48 VOUT-.n29 VOUT-.t36 4.8295
R49 VOUT-.n31 VOUT-.t105 4.8295
R50 VOUT-.n32 VOUT-.t76 4.8295
R51 VOUT-.n34 VOUT-.t42 4.8295
R52 VOUT-.n35 VOUT-.t30 4.8295
R53 VOUT-.n37 VOUT-.t88 4.8295
R54 VOUT-.n38 VOUT-.t72 4.8295
R55 VOUT-.n40 VOUT-.t51 4.8295
R56 VOUT-.n41 VOUT-.t33 4.8295
R57 VOUT-.n43 VOUT-.t92 4.8295
R58 VOUT-.n44 VOUT-.t77 4.8295
R59 VOUT-.n96 VOUT-.t119 4.8295
R60 VOUT-.n69 VOUT-.t129 4.806
R61 VOUT-.n68 VOUT-.t26 4.806
R62 VOUT-.n67 VOUT-.t64 4.806
R63 VOUT-.n66 VOUT-.t101 4.806
R64 VOUT-.n65 VOUT-.t82 4.806
R65 VOUT-.n64 VOUT-.t56 4.806
R66 VOUT-.n63 VOUT-.t98 4.806
R67 VOUT-.n62 VOUT-.t78 4.806
R68 VOUT-.n61 VOUT-.t118 4.806
R69 VOUT-.n60 VOUT-.t149 4.806
R70 VOUT-.n28 VOUT-.t97 4.806
R71 VOUT-.n27 VOUT-.t133 4.806
R72 VOUT-.n26 VOUT-.t28 4.806
R73 VOUT-.n25 VOUT-.t63 4.806
R74 VOUT-.n24 VOUT-.t117 4.806
R75 VOUT-.n23 VOUT-.t69 4.806
R76 VOUT-.n22 VOUT-.t104 4.806
R77 VOUT-.n21 VOUT-.t150 4.806
R78 VOUT-.n20 VOUT-.t46 4.806
R79 VOUT-.n19 VOUT-.t86 4.806
R80 VOUT-.n47 VOUT-.t143 4.5005
R81 VOUT-.n46 VOUT-.t113 4.5005
R82 VOUT-.n48 VOUT-.t122 4.5005
R83 VOUT-.n49 VOUT-.t154 4.5005
R84 VOUT-.n50 VOUT-.t126 4.5005
R85 VOUT-.n51 VOUT-.t148 4.5005
R86 VOUT-.n52 VOUT-.t49 4.5005
R87 VOUT-.n53 VOUT-.t155 4.5005
R88 VOUT-.n54 VOUT-.t62 4.5005
R89 VOUT-.n55 VOUT-.t103 4.5005
R90 VOUT-.n56 VOUT-.t68 4.5005
R91 VOUT-.n57 VOUT-.t156 4.5005
R92 VOUT-.n58 VOUT-.t54 4.5005
R93 VOUT-.n59 VOUT-.t23 4.5005
R94 VOUT-.n60 VOUT-.t115 4.5005
R95 VOUT-.n61 VOUT-.t75 4.5005
R96 VOUT-.n62 VOUT-.t34 4.5005
R97 VOUT-.n63 VOUT-.t55 4.5005
R98 VOUT-.n64 VOUT-.t20 4.5005
R99 VOUT-.n65 VOUT-.t37 4.5005
R100 VOUT-.n66 VOUT-.t59 4.5005
R101 VOUT-.n67 VOUT-.t24 4.5005
R102 VOUT-.n68 VOUT-.t127 4.5005
R103 VOUT-.n69 VOUT-.t90 4.5005
R104 VOUT-.n71 VOUT-.t110 4.5005
R105 VOUT-.n70 VOUT-.t73 4.5005
R106 VOUT-.n72 VOUT-.t50 4.5005
R107 VOUT-.n74 VOUT-.t139 4.5005
R108 VOUT-.n73 VOUT-.t109 4.5005
R109 VOUT-.n75 VOUT-.t87 4.5005
R110 VOUT-.n77 VOUT-.t32 4.5005
R111 VOUT-.n76 VOUT-.t137 4.5005
R112 VOUT-.n78 VOUT-.t41 4.5005
R113 VOUT-.n80 VOUT-.t134 4.5005
R114 VOUT-.n79 VOUT-.t99 4.5005
R115 VOUT-.n81 VOUT-.t142 4.5005
R116 VOUT-.n83 VOUT-.t94 4.5005
R117 VOUT-.n82 VOUT-.t58 4.5005
R118 VOUT-.n84 VOUT-.t38 4.5005
R119 VOUT-.n86 VOUT-.t131 4.5005
R120 VOUT-.n85 VOUT-.t93 4.5005
R121 VOUT-.n87 VOUT-.t140 4.5005
R122 VOUT-.n89 VOUT-.t91 4.5005
R123 VOUT-.n88 VOUT-.t52 4.5005
R124 VOUT-.n90 VOUT-.t102 4.5005
R125 VOUT-.n92 VOUT-.t47 4.5005
R126 VOUT-.n91 VOUT-.t152 4.5005
R127 VOUT-.n93 VOUT-.t60 4.5005
R128 VOUT-.n95 VOUT-.t145 4.5005
R129 VOUT-.n94 VOUT-.t120 4.5005
R130 VOUT-.n18 VOUT-.t43 4.5005
R131 VOUT-.n17 VOUT-.t147 4.5005
R132 VOUT-.n19 VOUT-.t29 4.5005
R133 VOUT-.n20 VOUT-.t81 4.5005
R134 VOUT-.n21 VOUT-.t128 4.5005
R135 VOUT-.n22 VOUT-.t136 4.5005
R136 VOUT-.n23 VOUT-.t44 4.5005
R137 VOUT-.n24 VOUT-.t45 4.5005
R138 VOUT-.n25 VOUT-.t61 4.5005
R139 VOUT-.n26 VOUT-.t111 4.5005
R140 VOUT-.n27 VOUT-.t19 4.5005
R141 VOUT-.n28 VOUT-.t67 4.5005
R142 VOUT-.n30 VOUT-.t83 4.5005
R143 VOUT-.n29 VOUT-.t130 4.5005
R144 VOUT-.n31 VOUT-.t151 4.5005
R145 VOUT-.n33 VOUT-.t116 4.5005
R146 VOUT-.n32 VOUT-.t25 4.5005
R147 VOUT-.n34 VOUT-.t146 4.5005
R148 VOUT-.n36 VOUT-.t100 4.5005
R149 VOUT-.n35 VOUT-.t66 4.5005
R150 VOUT-.n37 VOUT-.t48 4.5005
R151 VOUT-.n39 VOUT-.t138 4.5005
R152 VOUT-.n38 VOUT-.t108 4.5005
R153 VOUT-.n40 VOUT-.t153 4.5005
R154 VOUT-.n42 VOUT-.t107 4.5005
R155 VOUT-.n41 VOUT-.t71 4.5005
R156 VOUT-.n43 VOUT-.t53 4.5005
R157 VOUT-.n45 VOUT-.t141 4.5005
R158 VOUT-.n44 VOUT-.t112 4.5005
R159 VOUT-.n99 VOUT-.t132 4.5005
R160 VOUT-.n98 VOUT-.t95 4.5005
R161 VOUT-.n97 VOUT-.t40 4.5005
R162 VOUT-.n96 VOUT-.t144 4.5005
R163 VOUT-.n16 VOUT-.n14 4.5005
R164 VOUT-.n3 VOUT-.t3 3.42907
R165 VOUT-.n3 VOUT-.t17 3.42907
R166 VOUT-.n1 VOUT-.t7 3.42907
R167 VOUT-.n1 VOUT-.t4 3.42907
R168 VOUT-.n0 VOUT-.t9 3.42907
R169 VOUT-.n0 VOUT-.t8 3.42907
R170 VOUT- VOUT-.n5 2.84425
R171 VOUT-.n5 VOUT-.n4 2.03175
R172 VOUT-.n4 VOUT-.n2 1.1255
R173 VOUT-.n11 VOUT-.n9 0.563
R174 VOUT-.n13 VOUT-.n11 0.563
R175 VOUT-.n14 VOUT-.n13 0.563
R176 VOUT-.n47 VOUT-.n46 0.3295
R177 VOUT-.n50 VOUT-.n49 0.3295
R178 VOUT-.n49 VOUT-.n48 0.3295
R179 VOUT-.n53 VOUT-.n52 0.3295
R180 VOUT-.n52 VOUT-.n51 0.3295
R181 VOUT-.n56 VOUT-.n55 0.3295
R182 VOUT-.n55 VOUT-.n54 0.3295
R183 VOUT-.n59 VOUT-.n58 0.3295
R184 VOUT-.n58 VOUT-.n57 0.3295
R185 VOUT-.n61 VOUT-.n60 0.3295
R186 VOUT-.n62 VOUT-.n61 0.3295
R187 VOUT-.n63 VOUT-.n62 0.3295
R188 VOUT-.n64 VOUT-.n63 0.3295
R189 VOUT-.n65 VOUT-.n64 0.3295
R190 VOUT-.n66 VOUT-.n65 0.3295
R191 VOUT-.n67 VOUT-.n66 0.3295
R192 VOUT-.n68 VOUT-.n67 0.3295
R193 VOUT-.n69 VOUT-.n68 0.3295
R194 VOUT-.n71 VOUT-.n69 0.3295
R195 VOUT-.n71 VOUT-.n70 0.3295
R196 VOUT-.n74 VOUT-.n72 0.3295
R197 VOUT-.n74 VOUT-.n73 0.3295
R198 VOUT-.n77 VOUT-.n75 0.3295
R199 VOUT-.n77 VOUT-.n76 0.3295
R200 VOUT-.n80 VOUT-.n78 0.3295
R201 VOUT-.n80 VOUT-.n79 0.3295
R202 VOUT-.n83 VOUT-.n81 0.3295
R203 VOUT-.n83 VOUT-.n82 0.3295
R204 VOUT-.n86 VOUT-.n84 0.3295
R205 VOUT-.n86 VOUT-.n85 0.3295
R206 VOUT-.n89 VOUT-.n87 0.3295
R207 VOUT-.n89 VOUT-.n88 0.3295
R208 VOUT-.n92 VOUT-.n90 0.3295
R209 VOUT-.n92 VOUT-.n91 0.3295
R210 VOUT-.n95 VOUT-.n93 0.3295
R211 VOUT-.n95 VOUT-.n94 0.3295
R212 VOUT-.n18 VOUT-.n17 0.3295
R213 VOUT-.n20 VOUT-.n19 0.3295
R214 VOUT-.n21 VOUT-.n20 0.3295
R215 VOUT-.n22 VOUT-.n21 0.3295
R216 VOUT-.n23 VOUT-.n22 0.3295
R217 VOUT-.n24 VOUT-.n23 0.3295
R218 VOUT-.n25 VOUT-.n24 0.3295
R219 VOUT-.n26 VOUT-.n25 0.3295
R220 VOUT-.n27 VOUT-.n26 0.3295
R221 VOUT-.n28 VOUT-.n27 0.3295
R222 VOUT-.n30 VOUT-.n28 0.3295
R223 VOUT-.n30 VOUT-.n29 0.3295
R224 VOUT-.n33 VOUT-.n31 0.3295
R225 VOUT-.n33 VOUT-.n32 0.3295
R226 VOUT-.n36 VOUT-.n34 0.3295
R227 VOUT-.n36 VOUT-.n35 0.3295
R228 VOUT-.n39 VOUT-.n37 0.3295
R229 VOUT-.n39 VOUT-.n38 0.3295
R230 VOUT-.n42 VOUT-.n40 0.3295
R231 VOUT-.n42 VOUT-.n41 0.3295
R232 VOUT-.n45 VOUT-.n43 0.3295
R233 VOUT-.n45 VOUT-.n44 0.3295
R234 VOUT-.n99 VOUT-.n98 0.3295
R235 VOUT-.n98 VOUT-.n97 0.3295
R236 VOUT-.n97 VOUT-.n96 0.3295
R237 VOUT-.n67 VOUT-.n50 0.306
R238 VOUT-.n66 VOUT-.n53 0.306
R239 VOUT-.n65 VOUT-.n56 0.306
R240 VOUT-.n64 VOUT-.n59 0.306
R241 VOUT-.n71 VOUT-.n47 0.2825
R242 VOUT-.n74 VOUT-.n71 0.2825
R243 VOUT-.n77 VOUT-.n74 0.2825
R244 VOUT-.n80 VOUT-.n77 0.2825
R245 VOUT-.n83 VOUT-.n80 0.2825
R246 VOUT-.n86 VOUT-.n83 0.2825
R247 VOUT-.n89 VOUT-.n86 0.2825
R248 VOUT-.n92 VOUT-.n89 0.2825
R249 VOUT-.n95 VOUT-.n92 0.2825
R250 VOUT-.n30 VOUT-.n18 0.2825
R251 VOUT-.n33 VOUT-.n30 0.2825
R252 VOUT-.n36 VOUT-.n33 0.2825
R253 VOUT-.n39 VOUT-.n36 0.2825
R254 VOUT-.n42 VOUT-.n39 0.2825
R255 VOUT-.n45 VOUT-.n42 0.2825
R256 VOUT-.n97 VOUT-.n45 0.2825
R257 VOUT-.n97 VOUT-.n95 0.2825
R258 cap_res_X cap_res_X.t0 49.083
R259 cap_res_X.t84 cap_res_X.t126 0.1603
R260 cap_res_X.t44 cap_res_X.t83 0.1603
R261 cap_res_X.t48 cap_res_X.t87 0.1603
R262 cap_res_X.t107 cap_res_X.t68 0.1603
R263 cap_res_X.t20 cap_res_X.t51 0.1603
R264 cap_res_X.t70 cap_res_X.t32 0.1603
R265 cap_res_X.t58 cap_res_X.t92 0.1603
R266 cap_res_X.t116 cap_res_X.t72 0.1603
R267 cap_res_X.t99 cap_res_X.t130 0.1603
R268 cap_res_X.t15 cap_res_X.t118 0.1603
R269 cap_res_X.t64 cap_res_X.t100 0.1603
R270 cap_res_X.t119 cap_res_X.t78 0.1603
R271 cap_res_X.t105 cap_res_X.t136 0.1603
R272 cap_res_X.t17 cap_res_X.t122 0.1603
R273 cap_res_X.t5 cap_res_X.t33 0.1603
R274 cap_res_X.t55 cap_res_X.t22 0.1603
R275 cap_res_X.t37 cap_res_X.t73 0.1603
R276 cap_res_X.t97 cap_res_X.t61 0.1603
R277 cap_res_X.t13 cap_res_X.t38 0.1603
R278 cap_res_X.t62 cap_res_X.t25 0.1603
R279 cap_res_X.t45 cap_res_X.t80 0.1603
R280 cap_res_X.t104 cap_res_X.t65 0.1603
R281 cap_res_X.t86 cap_res_X.t124 0.1603
R282 cap_res_X.t4 cap_res_X.t106 0.1603
R283 cap_res_X.t49 cap_res_X.t85 0.1603
R284 cap_res_X.t109 cap_res_X.t69 0.1603
R285 cap_res_X.t91 cap_res_X.t127 0.1603
R286 cap_res_X.t11 cap_res_X.t115 0.1603
R287 cap_res_X.t132 cap_res_X.t81 0.1603
R288 cap_res_X.t6 cap_res_X.t52 0.1603
R289 cap_res_X.t27 cap_res_X.t121 0.1603
R290 cap_res_X.t128 cap_res_X.t71 0.1603
R291 cap_res_X.t76 cap_res_X.t111 0.1603
R292 cap_res_X.t29 cap_res_X.t7 0.1603
R293 cap_res_X.t21 cap_res_X.t53 0.1603
R294 cap_res_X.t113 cap_res_X.t88 0.1603
R295 cap_res_X.t112 cap_res_X.t40 0.1603
R296 cap_res_X.t96 cap_res_X.t94 0.1603
R297 cap_res_X.t46 cap_res_X.t129 0.1603
R298 cap_res_X.t138 cap_res_X.t24 0.1603
R299 cap_res_X.t90 cap_res_X.t60 0.1603
R300 cap_res_X.t10 cap_res_X.t36 0.1603
R301 cap_res_X.t35 cap_res_X.t77 0.1603
R302 cap_res_X.t3 cap_res_X.t35 0.1603
R303 cap_res_X.t31 cap_res_X.t3 0.1603
R304 cap_res_X.t133 cap_res_X.t31 0.1603
R305 cap_res_X.t1 cap_res_X.t34 0.1603
R306 cap_res_X.t103 cap_res_X.t1 0.1603
R307 cap_res_X.t134 cap_res_X.t103 0.1603
R308 cap_res_X.t137 cap_res_X.t134 0.1603
R309 cap_res_X.t95 cap_res_X.t135 0.1603
R310 cap_res_X.t54 cap_res_X.t95 0.1603
R311 cap_res_X.t89 cap_res_X.t54 0.1603
R312 cap_res_X.t120 cap_res_X.t89 0.1603
R313 cap_res_X.t2 cap_res_X.t98 0.1603
R314 cap_res_X.t108 cap_res_X.t2 0.1603
R315 cap_res_X.t9 cap_res_X.t108 0.1603
R316 cap_res_X.t43 cap_res_X.t9 0.1603
R317 cap_res_X.n31 cap_res_X.t14 0.159278
R318 cap_res_X.t74 cap_res_X.n15 0.159278
R319 cap_res_X.t41 cap_res_X.n16 0.159278
R320 cap_res_X.t57 cap_res_X.n17 0.159278
R321 cap_res_X.t19 cap_res_X.n18 0.159278
R322 cap_res_X.t50 cap_res_X.n19 0.159278
R323 cap_res_X.t16 cap_res_X.n20 0.159278
R324 cap_res_X.t117 cap_res_X.n21 0.159278
R325 cap_res_X.t12 cap_res_X.n22 0.159278
R326 cap_res_X.t110 cap_res_X.n23 0.159278
R327 cap_res_X.t66 cap_res_X.n24 0.159278
R328 cap_res_X.t26 cap_res_X.n25 0.159278
R329 cap_res_X.t63 cap_res_X.n26 0.159278
R330 cap_res_X.t23 cap_res_X.n27 0.159278
R331 cap_res_X.t125 cap_res_X.n28 0.159278
R332 cap_res_X.t18 cap_res_X.n29 0.159278
R333 cap_res_X.t47 cap_res_X.n30 0.159278
R334 cap_res_X.n32 cap_res_X.t28 0.159278
R335 cap_res_X.n33 cap_res_X.t131 0.159278
R336 cap_res_X.n34 cap_res_X.t93 0.159278
R337 cap_res_X.n0 cap_res_X.t8 0.159278
R338 cap_res_X.n1 cap_res_X.t39 0.159278
R339 cap_res_X.n2 cap_res_X.t79 0.159278
R340 cap_res_X.n3 cap_res_X.t59 0.159278
R341 cap_res_X.n4 cap_res_X.t101 0.159278
R342 cap_res_X.n5 cap_res_X.t75 0.159278
R343 cap_res_X.n35 cap_res_X.t56 0.159278
R344 cap_res_X.t14 cap_res_X.t44 0.137822
R345 cap_res_X.n31 cap_res_X.t84 0.1368
R346 cap_res_X.n30 cap_res_X.t48 0.1368
R347 cap_res_X.n30 cap_res_X.t107 0.1368
R348 cap_res_X.n29 cap_res_X.t20 0.1368
R349 cap_res_X.n29 cap_res_X.t70 0.1368
R350 cap_res_X.n28 cap_res_X.t58 0.1368
R351 cap_res_X.n28 cap_res_X.t116 0.1368
R352 cap_res_X.n27 cap_res_X.t99 0.1368
R353 cap_res_X.n27 cap_res_X.t15 0.1368
R354 cap_res_X.n26 cap_res_X.t64 0.1368
R355 cap_res_X.n26 cap_res_X.t119 0.1368
R356 cap_res_X.n25 cap_res_X.t105 0.1368
R357 cap_res_X.n25 cap_res_X.t17 0.1368
R358 cap_res_X.n24 cap_res_X.t5 0.1368
R359 cap_res_X.n24 cap_res_X.t55 0.1368
R360 cap_res_X.n23 cap_res_X.t37 0.1368
R361 cap_res_X.n23 cap_res_X.t97 0.1368
R362 cap_res_X.n22 cap_res_X.t13 0.1368
R363 cap_res_X.n22 cap_res_X.t62 0.1368
R364 cap_res_X.n21 cap_res_X.t45 0.1368
R365 cap_res_X.n21 cap_res_X.t104 0.1368
R366 cap_res_X.n20 cap_res_X.t86 0.1368
R367 cap_res_X.n20 cap_res_X.t4 0.1368
R368 cap_res_X.n19 cap_res_X.t49 0.1368
R369 cap_res_X.n19 cap_res_X.t109 0.1368
R370 cap_res_X.n18 cap_res_X.t91 0.1368
R371 cap_res_X.n18 cap_res_X.t11 0.1368
R372 cap_res_X.n17 cap_res_X.t132 0.1368
R373 cap_res_X.n17 cap_res_X.t6 0.1368
R374 cap_res_X.n16 cap_res_X.t27 0.1368
R375 cap_res_X.n15 cap_res_X.t10 0.1368
R376 cap_res_X cap_res_X.t43 0.118
R377 cap_res_X.n6 cap_res_X.t128 0.114322
R378 cap_res_X.n7 cap_res_X.n6 0.1133
R379 cap_res_X.n8 cap_res_X.n7 0.1133
R380 cap_res_X.n9 cap_res_X.n8 0.1133
R381 cap_res_X.n10 cap_res_X.n9 0.1133
R382 cap_res_X.n11 cap_res_X.n10 0.1133
R383 cap_res_X.n12 cap_res_X.n11 0.1133
R384 cap_res_X.n13 cap_res_X.n12 0.1133
R385 cap_res_X.n14 cap_res_X.n13 0.1133
R386 cap_res_X.n16 cap_res_X.n14 0.1133
R387 cap_res_X.n32 cap_res_X.n31 0.1133
R388 cap_res_X.n33 cap_res_X.n32 0.1133
R389 cap_res_X.n34 cap_res_X.n33 0.1133
R390 cap_res_X.n1 cap_res_X.n0 0.1133
R391 cap_res_X.n2 cap_res_X.n1 0.1133
R392 cap_res_X.n3 cap_res_X.n2 0.1133
R393 cap_res_X.n4 cap_res_X.n3 0.1133
R394 cap_res_X.n5 cap_res_X.n4 0.1133
R395 cap_res_X.n35 cap_res_X.n5 0.1133
R396 cap_res_X.n35 cap_res_X.n34 0.1133
R397 cap_res_X.n6 cap_res_X.t76 0.00152174
R398 cap_res_X.n7 cap_res_X.t29 0.00152174
R399 cap_res_X.n8 cap_res_X.t21 0.00152174
R400 cap_res_X.n9 cap_res_X.t113 0.00152174
R401 cap_res_X.n10 cap_res_X.t112 0.00152174
R402 cap_res_X.n11 cap_res_X.t96 0.00152174
R403 cap_res_X.n12 cap_res_X.t46 0.00152174
R404 cap_res_X.n13 cap_res_X.t138 0.00152174
R405 cap_res_X.n14 cap_res_X.t90 0.00152174
R406 cap_res_X.n15 cap_res_X.t114 0.00152174
R407 cap_res_X.n16 cap_res_X.t74 0.00152174
R408 cap_res_X.n17 cap_res_X.t41 0.00152174
R409 cap_res_X.n18 cap_res_X.t57 0.00152174
R410 cap_res_X.n19 cap_res_X.t19 0.00152174
R411 cap_res_X.n20 cap_res_X.t50 0.00152174
R412 cap_res_X.n21 cap_res_X.t16 0.00152174
R413 cap_res_X.n22 cap_res_X.t117 0.00152174
R414 cap_res_X.n23 cap_res_X.t12 0.00152174
R415 cap_res_X.n24 cap_res_X.t110 0.00152174
R416 cap_res_X.n25 cap_res_X.t66 0.00152174
R417 cap_res_X.n26 cap_res_X.t26 0.00152174
R418 cap_res_X.n27 cap_res_X.t63 0.00152174
R419 cap_res_X.n28 cap_res_X.t23 0.00152174
R420 cap_res_X.n29 cap_res_X.t125 0.00152174
R421 cap_res_X.n30 cap_res_X.t18 0.00152174
R422 cap_res_X.n31 cap_res_X.t47 0.00152174
R423 cap_res_X.n32 cap_res_X.t67 0.00152174
R424 cap_res_X.n33 cap_res_X.t30 0.00152174
R425 cap_res_X.n34 cap_res_X.t133 0.00152174
R426 cap_res_X.n0 cap_res_X.t42 0.00152174
R427 cap_res_X.n1 cap_res_X.t82 0.00152174
R428 cap_res_X.n2 cap_res_X.t123 0.00152174
R429 cap_res_X.n3 cap_res_X.t102 0.00152174
R430 cap_res_X.n4 cap_res_X.t137 0.00152174
R431 cap_res_X.n5 cap_res_X.t120 0.00152174
R432 cap_res_X.t98 cap_res_X.n35 0.00152174
R433 V_tail_gate.n10 V_tail_gate.t12 610.534
R434 V_tail_gate.n3 V_tail_gate.t9 610.534
R435 V_tail_gate.n10 V_tail_gate.t16 433.8
R436 V_tail_gate.n11 V_tail_gate.t4 433.8
R437 V_tail_gate.n12 V_tail_gate.t15 433.8
R438 V_tail_gate.n13 V_tail_gate.t23 433.8
R439 V_tail_gate.n14 V_tail_gate.t13 433.8
R440 V_tail_gate.n15 V_tail_gate.t8 433.8
R441 V_tail_gate.n16 V_tail_gate.t19 433.8
R442 V_tail_gate.n17 V_tail_gate.t6 433.8
R443 V_tail_gate.n18 V_tail_gate.t17 433.8
R444 V_tail_gate.n19 V_tail_gate.t5 433.8
R445 V_tail_gate.n20 V_tail_gate.t10 433.8
R446 V_tail_gate.n9 V_tail_gate.t20 433.8
R447 V_tail_gate.n8 V_tail_gate.t7 433.8
R448 V_tail_gate.n7 V_tail_gate.t18 433.8
R449 V_tail_gate.n6 V_tail_gate.t14 433.8
R450 V_tail_gate.n5 V_tail_gate.t22 433.8
R451 V_tail_gate.n4 V_tail_gate.t11 433.8
R452 V_tail_gate.n3 V_tail_gate.t21 433.8
R453 V_tail_gate.n2 V_tail_gate.n0 183.029
R454 V_tail_gate.n20 V_tail_gate.n19 176.733
R455 V_tail_gate.n19 V_tail_gate.n18 176.733
R456 V_tail_gate.n18 V_tail_gate.n17 176.733
R457 V_tail_gate.n17 V_tail_gate.n16 176.733
R458 V_tail_gate.n16 V_tail_gate.n15 176.733
R459 V_tail_gate.n15 V_tail_gate.n14 176.733
R460 V_tail_gate.n14 V_tail_gate.n13 176.733
R461 V_tail_gate.n13 V_tail_gate.n12 176.733
R462 V_tail_gate.n12 V_tail_gate.n11 176.733
R463 V_tail_gate.n11 V_tail_gate.n10 176.733
R464 V_tail_gate.n4 V_tail_gate.n3 176.733
R465 V_tail_gate.n5 V_tail_gate.n4 176.733
R466 V_tail_gate.n6 V_tail_gate.n5 176.733
R467 V_tail_gate.n7 V_tail_gate.n6 176.733
R468 V_tail_gate.n8 V_tail_gate.n7 176.733
R469 V_tail_gate.n9 V_tail_gate.n8 176.733
R470 V_tail_gate V_tail_gate.n21 161.633
R471 V_tail_gate V_tail_gate.n2 59.6601
R472 V_tail_gate.n21 V_tail_gate.n20 56.2338
R473 V_tail_gate.n21 V_tail_gate.n9 56.2338
R474 V_tail_gate.n2 V_tail_gate.n1 53.2453
R475 V_tail_gate.n1 V_tail_gate.t1 16.0005
R476 V_tail_gate.n1 V_tail_gate.t2 16.0005
R477 V_tail_gate.n0 V_tail_gate.t0 16.0005
R478 V_tail_gate.n0 V_tail_gate.t3 16.0005
R479 GNDA.n148 GNDA.n147 41223.8
R480 GNDA.n152 GNDA.n47 40376.5
R481 GNDA.n51 GNDA.n50 40376.5
R482 GNDA.n149 GNDA.n24 32661.5
R483 GNDA.n245 GNDA.n24 32661.5
R484 GNDA.n48 GNDA.n47 30739.1
R485 GNDA.n50 GNDA.n48 30739.1
R486 GNDA.n49 GNDA.n47 29723.7
R487 GNDA.n148 GNDA.n52 28430.8
R488 GNDA.n246 GNDA.n45 28430.8
R489 GNDA.n151 GNDA.n150 28372.4
R490 GNDA.n152 GNDA.n151 27462.1
R491 GNDA.n50 GNDA.n49 25662.2
R492 GNDA.n152 GNDA.n46 25233.2
R493 GNDA.n51 GNDA.n46 24115.4
R494 GNDA.n151 GNDA.n24 19630.8
R495 GNDA.n297 GNDA.n24 19630.8
R496 GNDA.n150 GNDA.n149 14773.1
R497 GNDA.n245 GNDA.n244 14714.3
R498 GNDA.n298 GNDA.n23 10835
R499 GNDA.n296 GNDA.n23 10835
R500 GNDA.n296 GNDA.n22 10835
R501 GNDA.n298 GNDA.n22 10835
R502 GNDA.n247 GNDA.n246 10371.4
R503 GNDA.n151 GNDA.n48 9476.92
R504 GNDA.n55 GNDA.n6 9308.25
R505 GNDA.n302 GNDA.n6 9308.25
R506 GNDA.n55 GNDA.n7 9308.25
R507 GNDA.n302 GNDA.n7 9308.25
R508 GNDA.n255 GNDA.n250 9259
R509 GNDA.n257 GNDA.n250 8914.25
R510 GNDA.n49 GNDA.n46 8677.78
R511 GNDA.n255 GNDA.n43 8175.5
R512 GNDA.n257 GNDA.n43 7830.75
R513 GNDA.n120 GNDA.n61 7732.25
R514 GNDA.n120 GNDA.n62 7732.25
R515 GNDA.n122 GNDA.n61 7732.25
R516 GNDA.n122 GNDA.n62 7732.25
R517 GNDA.n203 GNDA.n163 7732.25
R518 GNDA.n234 GNDA.n163 7732.25
R519 GNDA.n203 GNDA.n171 7732.25
R520 GNDA.n234 GNDA.n171 7732.25
R521 GNDA.n100 GNDA.n78 7338.25
R522 GNDA.n182 GNDA.n153 7338.25
R523 GNDA.n242 GNDA.n153 7289
R524 GNDA.n95 GNDA.n78 7092
R525 GNDA.n111 GNDA.n69 6057.75
R526 GNDA.n113 GNDA.n111 6057.75
R527 GNDA.n69 GNDA.n66 6057.75
R528 GNDA.n113 GNDA.n66 6057.75
R529 GNDA.n168 GNDA.n161 6057.75
R530 GNDA.n237 GNDA.n161 6057.75
R531 GNDA.n168 GNDA.n162 6057.75
R532 GNDA.n237 GNDA.n162 6057.75
R533 GNDA.n244 GNDA.n243 5592.24
R534 GNDA.n100 GNDA.n79 5319
R535 GNDA.n182 GNDA.n154 5319
R536 GNDA.n95 GNDA.n79 5269.75
R537 GNDA.n242 GNDA.n154 5269.75
R538 GNDA.n107 GNDA.n73 5171.25
R539 GNDA.n196 GNDA.n176 5171.25
R540 GNDA.n103 GNDA.n73 5122
R541 GNDA.n178 GNDA.n176 5122
R542 GNDA.n107 GNDA.n74 4944.7
R543 GNDA.n196 GNDA.n195 4944.7
R544 GNDA.n269 GNDA.n25 4925
R545 GNDA.n283 GNDA.n25 4925
R546 GNDA.n103 GNDA.n74 4895.45
R547 GNDA.n195 GNDA.n178 4895.45
R548 GNDA.n269 GNDA.n26 4728
R549 GNDA.n283 GNDA.n26 4728
R550 GNDA.n150 GNDA.n52 4727.03
R551 GNDA.n144 GNDA.n32 3595.25
R552 GNDA.n266 GNDA.n32 3595.25
R553 GNDA.n144 GNDA.n33 3250.5
R554 GNDA.n266 GNDA.n33 3250.5
R555 GNDA.n251 GNDA.n5 3053.5
R556 GNDA.n305 GNDA.n5 3004.25
R557 GNDA.n251 GNDA.n3 2955
R558 GNDA.n246 GNDA.n245 2933.33
R559 GNDA.n149 GNDA.n148 2933.33
R560 GNDA.n305 GNDA.n3 2905.75
R561 GNDA.n93 GNDA.n84 2326.02
R562 GNDA.n86 GNDA.n84 2326.02
R563 GNDA.n192 GNDA.n179 2326.02
R564 GNDA.n185 GNDA.n179 2326.02
R565 GNDA.n89 GNDA.n84 1114.8
R566 GNDA.n189 GNDA.n179 1114.8
R567 GNDA.n158 GNDA.t223 734.418
R568 GNDA.n164 GNDA.t215 734.418
R569 GNDA.n67 GNDA.t203 734.418
R570 GNDA.n70 GNDA.t188 734.418
R571 GNDA.n295 GNDA.n289 704
R572 GNDA.n295 GNDA.n294 697.601
R573 GNDA.n225 GNDA.t154 682.201
R574 GNDA.n260 GNDA.t176 666.134
R575 GNDA.n52 GNDA.n51 624.324
R576 GNDA.n191 GNDA.n180 617.601
R577 GNDA.n92 GNDA.n87 617.601
R578 GNDA.n254 GNDA.n253 601.601
R579 GNDA.n301 GNDA.n300 598.4
R580 GNDA.n300 GNDA.n17 598.4
R581 GNDA.n172 GNDA.t212 535.191
R582 GNDA.n199 GNDA.t218 535.191
R583 GNDA.n63 GNDA.t173 535.191
R584 GNDA.n117 GNDA.t167 535.191
R585 GNDA.n254 GNDA.n39 531.201
R586 GNDA.n232 GNDA.n204 496
R587 GNDA.n123 GNDA.n60 496
R588 GNDA.n8 GNDA.t194 493.418
R589 GNDA.n12 GNDA.t182 493.418
R590 GNDA.n11 GNDA.t206 493.418
R591 GNDA.n10 GNDA.t164 493.418
R592 GNDA.n290 GNDA.t197 493.418
R593 GNDA.n291 GNDA.t185 493.418
R594 GNDA.n20 GNDA.t158 493.418
R595 GNDA.n18 GNDA.t221 493.418
R596 GNDA.n286 GNDA.t179 493.418
R597 GNDA.n285 GNDA.t170 493.418
R598 GNDA.n233 GNDA.n232 489.601
R599 GNDA.n123 GNDA.n59 489.601
R600 GNDA.n157 GNDA.n156 476.8
R601 GNDA.n99 GNDA.n80 476.8
R602 GNDA.n241 GNDA.n155 448
R603 GNDA.n96 GNDA.n81 448
R604 GNDA.n263 GNDA.t191 441.2
R605 GNDA.n258 GNDA.n40 428.8
R606 GNDA.n141 GNDA.t200 425.134
R607 GNDA.n16 GNDA.n15 422.401
R608 GNDA.n13 GNDA.n9 422.401
R609 GNDA.n293 GNDA.n292 422.401
R610 GNDA.n288 GNDA.n287 422.401
R611 GNDA.n95 GNDA.t241 402.776
R612 GNDA.n167 GNDA.n160 387.2
R613 GNDA.n115 GNDA.n114 387.2
R614 GNDA.n238 GNDA.n160 380.8
R615 GNDA.n115 GNDA.n65 380.8
R616 GNDA.n259 GNDA.n258 355.2
R617 GNDA.n241 GNDA.n240 342.401
R618 GNDA.n97 GNDA.n96 342.401
R619 GNDA.n177 GNDA.n174 332.8
R620 GNDA.n104 GNDA.n76 332.8
R621 GNDA.n27 GNDA.t161 332.75
R622 GNDA.n29 GNDA.t209 332.75
R623 GNDA.n197 GNDA.n175 321.281
R624 GNDA.n106 GNDA.n105 321.281
R625 GNDA.n177 GNDA.n175 318.08
R626 GNDA.n105 GNDA.n104 318.08
R627 GNDA.n204 GNDA.n202 310.401
R628 GNDA.n118 GNDA.n60 310.401
R629 GNDA.n233 GNDA.n173 304
R630 GNDA.n64 GNDA.n59 304
R631 GNDA.n282 GNDA.n281 300.8
R632 GNDA.n281 GNDA.n270 300.8
R633 GNDA.n198 GNDA.n174 300.8
R634 GNDA.n76 GNDA.n75 300.8
R635 GNDA.n191 GNDA.n190 296
R636 GNDA.n90 GNDA.n87 296
R637 GNDA.n238 GNDA.n237 292.5
R638 GNDA.n237 GNDA.n236 292.5
R639 GNDA.n162 GNDA.n160 292.5
R640 GNDA.t37 GNDA.n162 292.5
R641 GNDA.n168 GNDA.n167 292.5
R642 GNDA.n169 GNDA.n168 292.5
R643 GNDA.n165 GNDA.n161 292.5
R644 GNDA.t37 GNDA.n161 292.5
R645 GNDA.n242 GNDA.n241 292.5
R646 GNDA.n243 GNDA.n242 292.5
R647 GNDA.n240 GNDA.n154 292.5
R648 GNDA.n187 GNDA.n154 292.5
R649 GNDA.n182 GNDA.n157 292.5
R650 GNDA.n183 GNDA.n182 292.5
R651 GNDA.n156 GNDA.n153 292.5
R652 GNDA.n187 GNDA.n153 292.5
R653 GNDA.n190 GNDA.n189 292.5
R654 GNDA.n189 GNDA.n188 292.5
R655 GNDA.n176 GNDA.n174 292.5
R656 GNDA.n194 GNDA.n176 292.5
R657 GNDA.n178 GNDA.n177 292.5
R658 GNDA.n184 GNDA.n178 292.5
R659 GNDA.n195 GNDA.n175 292.5
R660 GNDA.n195 GNDA.n194 292.5
R661 GNDA.n197 GNDA.n196 292.5
R662 GNDA.n196 GNDA.n45 292.5
R663 GNDA.n234 GNDA.n233 292.5
R664 GNDA.n235 GNDA.n234 292.5
R665 GNDA.n201 GNDA.n163 292.5
R666 GNDA.n170 GNDA.n163 292.5
R667 GNDA.n204 GNDA.n203 292.5
R668 GNDA.n203 GNDA.n44 292.5
R669 GNDA.n232 GNDA.n171 292.5
R670 GNDA.n171 GNDA.n170 292.5
R671 GNDA.n107 GNDA.n106 292.5
R672 GNDA.n108 GNDA.n107 292.5
R673 GNDA.n105 GNDA.n74 292.5
R674 GNDA.n77 GNDA.n74 292.5
R675 GNDA.n104 GNDA.n103 292.5
R676 GNDA.n103 GNDA.n102 292.5
R677 GNDA.n76 GNDA.n73 292.5
R678 GNDA.n77 GNDA.n73 292.5
R679 GNDA.n62 GNDA.n60 292.5
R680 GNDA.n62 GNDA.n53 292.5
R681 GNDA.n123 GNDA.n122 292.5
R682 GNDA.n122 GNDA.n121 292.5
R683 GNDA.n61 GNDA.n59 292.5
R684 GNDA.n110 GNDA.n61 292.5
R685 GNDA.n120 GNDA.n119 292.5
R686 GNDA.n121 GNDA.n120 292.5
R687 GNDA.n114 GNDA.n113 292.5
R688 GNDA.n113 GNDA.n112 292.5
R689 GNDA.n115 GNDA.n66 292.5
R690 GNDA.t60 GNDA.n66 292.5
R691 GNDA.n69 GNDA.n65 292.5
R692 GNDA.n109 GNDA.n69 292.5
R693 GNDA.n111 GNDA.n72 292.5
R694 GNDA.n111 GNDA.t60 292.5
R695 GNDA.n100 GNDA.n99 292.5
R696 GNDA.n101 GNDA.n100 292.5
R697 GNDA.n97 GNDA.n79 292.5
R698 GNDA.n82 GNDA.n79 292.5
R699 GNDA.n96 GNDA.n95 292.5
R700 GNDA.n80 GNDA.n78 292.5
R701 GNDA.n83 GNDA.n78 292.5
R702 GNDA.n90 GNDA.n89 292.5
R703 GNDA.n89 GNDA.n88 292.5
R704 GNDA.n283 GNDA.n282 292.5
R705 GNDA.n284 GNDA.n283 292.5
R706 GNDA.n281 GNDA.n26 292.5
R707 GNDA.n41 GNDA.n26 292.5
R708 GNDA.n270 GNDA.n269 292.5
R709 GNDA.n269 GNDA.n268 292.5
R710 GNDA.n30 GNDA.n25 292.5
R711 GNDA.n41 GNDA.n25 292.5
R712 GNDA.n306 GNDA.n305 292.5
R713 GNDA.n305 GNDA.n304 292.5
R714 GNDA.n307 GNDA.n3 292.5
R715 GNDA.t235 GNDA.n3 292.5
R716 GNDA.n251 GNDA.n2 292.5
R717 GNDA.n252 GNDA.n251 292.5
R718 GNDA.n5 GNDA.n4 292.5
R719 GNDA.t235 GNDA.n5 292.5
R720 GNDA.n266 GNDA.n265 292.5
R721 GNDA.n267 GNDA.n266 292.5
R722 GNDA.n35 GNDA.n33 292.5
R723 GNDA.n54 GNDA.n33 292.5
R724 GNDA.n144 GNDA.n143 292.5
R725 GNDA.n145 GNDA.n144 292.5
R726 GNDA.n34 GNDA.n32 292.5
R727 GNDA.n54 GNDA.n32 292.5
R728 GNDA.n253 GNDA.n250 292.5
R729 GNDA.n250 GNDA.n249 292.5
R730 GNDA.n258 GNDA.n257 292.5
R731 GNDA.n257 GNDA.n256 292.5
R732 GNDA.n43 GNDA.n39 292.5
R733 GNDA.n43 GNDA.n42 292.5
R734 GNDA.n255 GNDA.n254 292.5
R735 GNDA.n256 GNDA.n255 292.5
R736 GNDA.n302 GNDA.n301 292.5
R737 GNDA.n303 GNDA.n302 292.5
R738 GNDA.n14 GNDA.n6 292.5
R739 GNDA.n297 GNDA.n6 292.5
R740 GNDA.n55 GNDA.n17 292.5
R741 GNDA.n56 GNDA.n55 292.5
R742 GNDA.n300 GNDA.n7 292.5
R743 GNDA.n297 GNDA.n7 292.5
R744 GNDA.n299 GNDA.n298 292.5
R745 GNDA.n298 GNDA.n297 292.5
R746 GNDA.n289 GNDA.n22 292.5
R747 GNDA.n146 GNDA.n22 292.5
R748 GNDA.n296 GNDA.n295 292.5
R749 GNDA.n297 GNDA.n296 292.5
R750 GNDA.n294 GNDA.n23 292.5
R751 GNDA.n248 GNDA.n23 292.5
R752 GNDA.n27 GNDA.t163 258.601
R753 GNDA.n29 GNDA.t211 258.601
R754 GNDA.n240 GNDA.n239 246.4
R755 GNDA.n98 GNDA.n97 246.4
R756 GNDA.n181 GNDA.n180 238.4
R757 GNDA.n92 GNDA.n91 238.4
R758 GNDA.n244 GNDA.n152 235.249
R759 GNDA.n143 GNDA.n34 233.601
R760 GNDA.n265 GNDA.n34 233.601
R761 GNDA.n276 GNDA.n274 227.096
R762 GNDA.n273 GNDA.n271 227.096
R763 GNDA.n276 GNDA.n275 226.534
R764 GNDA.n273 GNDA.n272 226.534
R765 GNDA.n172 GNDA.t214 224.525
R766 GNDA.n199 GNDA.t220 224.525
R767 GNDA.n63 GNDA.t175 224.525
R768 GNDA.n117 GNDA.t169 224.525
R769 GNDA.n279 GNDA.n278 222.034
R770 GNDA.n31 GNDA.n30 211.201
R771 GNDA.n30 GNDA.n28 211.201
R772 GNDA.n166 GNDA.n165 211.201
R773 GNDA.n165 GNDA.n159 211.201
R774 GNDA.n72 GNDA.n71 211.201
R775 GNDA.n72 GNDA.n68 211.201
R776 GNDA.n311 GNDA.n309 206.052
R777 GNDA.n129 GNDA.n127 206.052
R778 GNDA.n319 GNDA.n318 205.488
R779 GNDA.n317 GNDA.n316 205.488
R780 GNDA.n315 GNDA.n314 205.488
R781 GNDA.n313 GNDA.n312 205.488
R782 GNDA.n311 GNDA.n310 205.488
R783 GNDA.n137 GNDA.n136 205.488
R784 GNDA.n135 GNDA.n134 205.488
R785 GNDA.n133 GNDA.n132 205.488
R786 GNDA.n131 GNDA.n130 205.488
R787 GNDA.n129 GNDA.n128 205.488
R788 GNDA.n4 GNDA.n2 198.4
R789 GNDA.n306 GNDA.n4 195.201
R790 GNDA.n192 GNDA.n191 195
R791 GNDA.n193 GNDA.n192 195
R792 GNDA.n185 GNDA.n180 195
R793 GNDA.n186 GNDA.n185 195
R794 GNDA.n87 GNDA.n86 195
R795 GNDA.n86 GNDA.n85 195
R796 GNDA.n93 GNDA.n92 195
R797 GNDA.n94 GNDA.n93 195
R798 GNDA.n202 GNDA.n201 192
R799 GNDA.n119 GNDA.n118 192
R800 GNDA.n307 GNDA.n2 185.601
R801 GNDA.n307 GNDA.n306 182.4
R802 GNDA.n167 GNDA.n166 182.4
R803 GNDA.n114 GNDA.n68 182.4
R804 GNDA.n248 GNDA.n247 179.363
R805 GNDA.n238 GNDA.n159 176
R806 GNDA.n71 GNDA.n65 176
R807 GNDA.n247 GNDA.n44 171.817
R808 GNDA.n249 GNDA.n248 164.906
R809 GNDA.n263 GNDA.t193 162.857
R810 GNDA.n141 GNDA.t202 162.857
R811 GNDA.n301 GNDA.n9 160
R812 GNDA.n17 GNDA.n16 160
R813 GNDA.n289 GNDA.n288 160
R814 GNDA.n143 GNDA.n142 156.8
R815 GNDA.n259 GNDA.n39 153.601
R816 GNDA.n200 GNDA.n173 153.601
R817 GNDA.n116 GNDA.n64 153.601
R818 GNDA.n294 GNDA.n293 153.601
R819 GNDA.n158 GNDA.t225 152.994
R820 GNDA.n164 GNDA.t217 152.994
R821 GNDA.n67 GNDA.t205 152.994
R822 GNDA.n70 GNDA.t190 152.994
R823 GNDA.n265 GNDA.n264 150.4
R824 GNDA.n253 GNDA.n40 150.4
R825 GNDA.n85 GNDA.n52 150.329
R826 GNDA.n57 GNDA.n36 139.077
R827 GNDA.t216 GNDA.n169 130.731
R828 GNDA.n112 GNDA.t204 130.731
R829 GNDA.n147 GNDA.n146 127.249
R830 GNDA.n236 GNDA.n235 119.525
R831 GNDA.n110 GNDA.n109 119.525
R832 GNDA.n108 GNDA.t242 115.79
R833 GNDA.n8 GNDA.t196 113.974
R834 GNDA.n12 GNDA.t184 113.974
R835 GNDA.n11 GNDA.t208 113.974
R836 GNDA.n10 GNDA.t166 113.974
R837 GNDA.n290 GNDA.t199 113.974
R838 GNDA.n291 GNDA.t187 113.974
R839 GNDA.n20 GNDA.t160 113.974
R840 GNDA.n18 GNDA.t222 113.974
R841 GNDA.n286 GNDA.t181 113.974
R842 GNDA.n285 GNDA.t172 113.974
R843 GNDA.n102 GNDA.n101 112.055
R844 GNDA.n282 GNDA.n28 108.8
R845 GNDA.n270 GNDA.n31 108.8
R846 GNDA.n145 GNDA.t171 101.194
R847 GNDA.n85 GNDA.t234 101.183
R848 GNDA.n38 GNDA.n37 99.0842
R849 GNDA.n206 GNDA.n205 99.0842
R850 GNDA.n208 GNDA.n207 99.0842
R851 GNDA.n210 GNDA.n209 99.0842
R852 GNDA.n212 GNDA.n211 99.0842
R853 GNDA.n214 GNDA.n213 99.0842
R854 GNDA.n216 GNDA.n215 99.0842
R855 GNDA.n218 GNDA.n217 99.0842
R856 GNDA.n220 GNDA.n219 99.0842
R857 GNDA.n222 GNDA.n221 99.0842
R858 GNDA.n224 GNDA.n223 99.0842
R859 GNDA.n231 GNDA.n230 95.101
R860 GNDA.n124 GNDA.n58 95.101
R861 GNDA.n225 GNDA.t157 94.8842
R862 GNDA.n260 GNDA.t178 94.8842
R863 GNDA.n126 GNDA.n125 94.601
R864 GNDA.n229 GNDA.n228 94.601
R865 GNDA.n94 GNDA.n83 92.5103
R866 GNDA.n146 GNDA.n145 89.9494
R867 GNDA.t241 GNDA.t69 89.644
R868 GNDA.t94 GNDA.t234 89.644
R869 GNDA.n239 GNDA.n157 86.4005
R870 GNDA.n99 GNDA.n98 86.4005
R871 GNDA.t4 GNDA.t85 82.1737
R872 GNDA.t82 GNDA.t249 82.1737
R873 GNDA.t79 GNDA.t83 82.1737
R874 GNDA.t228 GNDA.t224 82.1737
R875 GNDA.t111 GNDA.t189 82.1737
R876 GNDA.t43 GNDA.t112 82.1737
R877 GNDA.t19 GNDA.t32 82.1737
R878 GNDA.t101 GNDA.t67 82.1737
R879 GNDA.t96 GNDA.n45 78.6626
R880 GNDA.n243 GNDA.t84 78.6626
R881 GNDA.t99 GNDA.t219 78.4385
R882 GNDA.t168 GNDA.t248 78.4385
R883 GNDA.n184 GNDA.n183 76.1251
R884 GNDA.t77 GNDA.t99 70.9682
R885 GNDA.t213 GNDA.t228 70.9682
R886 GNDA.t174 GNDA.t111 70.9682
R887 GNDA.t248 GNDA.t29 70.9682
R888 GNDA.n299 GNDA.n21 64.0005
R889 GNDA.n299 GNDA.n19 64.0005
R890 GNDA.n264 GNDA.n35 60.8005
R891 GNDA.t34 GNDA.t155 59.9664
R892 GNDA.t7 GNDA.n83 57.241
R893 GNDA.t75 GNDA.t4 56.0277
R894 GNDA.t35 GNDA.t79 56.0277
R895 GNDA.t97 GNDA.t43 56.0277
R896 GNDA.t67 GNDA.t27 56.0277
R897 GNDA.n142 GNDA.n35 54.4005
R898 GNDA.t18 GNDA.n186 53.2877
R899 GNDA.t12 GNDA.t106 52.4707
R900 GNDA.t93 GNDA.t102 52.4707
R901 GNDA.t207 GNDA.t162 52.4707
R902 GNDA.n292 GNDA.n21 51.2005
R903 GNDA.n287 GNDA.n19 51.2005
R904 GNDA.n88 GNDA.t234 49.1464
R905 GNDA.n170 GNDA.t108 48.5574
R906 GNDA.n82 GNDA.t94 48.5574
R907 GNDA.n77 GNDA.t242 48.5574
R908 GNDA.n121 GNDA.t11 48.5574
R909 GNDA.n278 GNDA.t57 48.0005
R910 GNDA.n278 GNDA.t42 48.0005
R911 GNDA.n275 GNDA.t66 48.0005
R912 GNDA.n275 GNDA.t105 48.0005
R913 GNDA.n274 GNDA.t107 48.0005
R914 GNDA.n274 GNDA.t103 48.0005
R915 GNDA.n272 GNDA.t232 48.0005
R916 GNDA.n272 GNDA.t87 48.0005
R917 GNDA.n271 GNDA.t14 48.0005
R918 GNDA.n271 GNDA.t40 48.0005
R919 GNDA.t73 GNDA.t126 44.9749
R920 GNDA.t72 GNDA.t148 44.9749
R921 GNDA.t237 GNDA.t144 44.9749
R922 GNDA.t88 GNDA.t134 44.9749
R923 GNDA.t47 GNDA.t114 44.9749
R924 GNDA.t0 GNDA.t130 44.9749
R925 GNDA.t46 GNDA.t152 44.9749
R926 GNDA.t49 GNDA.t128 44.9749
R927 GNDA.n236 GNDA.n45 44.8222
R928 GNDA.n109 GNDA.n108 44.8222
R929 GNDA.n190 GNDA.n181 44.8005
R930 GNDA.n91 GNDA.n90 44.8005
R931 GNDA.n188 GNDA.t113 43.1378
R932 GNDA.n56 GNDA.t16 41.2271
R933 GNDA.n297 GNDA.t109 41.2271
R934 GNDA.n256 GNDA.t150 41.2271
R935 GNDA.t95 GNDA.n303 41.2271
R936 GNDA.n303 GNDA.t198 41.2271
R937 GNDA.t9 GNDA.t37 41.0871
R938 GNDA.t37 GNDA.t82 41.0871
R939 GNDA.t69 GNDA.n82 41.0871
R940 GNDA.t100 GNDA.n77 41.0871
R941 GNDA.t60 GNDA.t19 41.0871
R942 GNDA.t60 GNDA.t50 41.0871
R943 GNDA.t171 GNDA.t201 37.4792
R944 GNDA.t54 GNDA.t192 37.4792
R945 GNDA.t53 GNDA.t210 37.4792
R946 GNDA.t39 GNDA.t51 37.4792
R947 GNDA.t246 GNDA.t86 37.4792
R948 GNDA.t17 GNDA.t56 37.4792
R949 GNDA.t240 GNDA.t41 37.4792
R950 GNDA.t233 GNDA.t65 37.4792
R951 GNDA.t180 GNDA.t104 37.4792
R952 GNDA.t52 GNDA.t140 37.4792
R953 GNDA.t150 GNDA.t73 37.4792
R954 GNDA.n320 GNDA.n319 36.9067
R955 GNDA.n138 GNDA.n137 36.6567
R956 GNDA.t16 GNDA.n54 33.7313
R957 GNDA.n268 GNDA.t238 33.7313
R958 GNDA.n267 GNDA.t13 33.7313
R959 GNDA.n42 GNDA.t231 33.7313
R960 GNDA.t120 GNDA.n284 33.7313
R961 GNDA.n304 GNDA.t195 33.7313
R962 GNDA.n170 GNDA.t9 33.6168
R963 GNDA.n121 GNDA.t50 33.6168
R964 GNDA.n194 GNDA.t96 32.9878
R965 GNDA.t10 GNDA.n187 32.9878
R966 GNDA.t192 GNDA.t165 29.9835
R967 GNDA.t210 GNDA.t71 29.9835
R968 GNDA.t58 GNDA.t13 29.9835
R969 GNDA.t62 GNDA.t39 29.9835
R970 GNDA.t231 GNDA.t1 29.9835
R971 GNDA.t159 GNDA.t183 29.9835
R972 GNDA.n169 GNDA.n44 29.8817
R973 GNDA.n112 GNDA.n53 29.8817
R974 GNDA.n239 GNDA.n238 28.413
R975 GNDA.n98 GNDA.n65 28.413
R976 GNDA.n233 GNDA.n198 28.038
R977 GNDA.n75 GNDA.n59 28.038
R978 GNDA.n187 GNDA.t18 27.9128
R979 GNDA.n297 GNDA.t146 26.2356
R980 GNDA.n252 GNDA.t124 26.2356
R981 GNDA.n249 GNDA.t198 26.2356
R982 GNDA.t108 GNDA.t75 26.1465
R983 GNDA.t249 GNDA.t35 26.1465
R984 GNDA.t32 GNDA.t97 26.1465
R985 GNDA.t27 GNDA.t11 26.1465
R986 GNDA.n201 GNDA.n200 25.6005
R987 GNDA.n119 GNDA.n116 25.6005
R988 GNDA.t202 GNDA.n57 24.0005
R989 GNDA.n57 GNDA.t239 24.0005
R990 GNDA.n294 GNDA.n0 23.488
R991 GNDA.t126 GNDA.t186 22.4877
R992 GNDA.t148 GNDA.t74 22.4877
R993 GNDA.t124 GNDA.t68 22.4877
R994 GNDA.t144 GNDA.t91 22.4877
R995 GNDA.t134 GNDA.t31 22.4877
R996 GNDA.t114 GNDA.t24 22.4877
R997 GNDA.t130 GNDA.t92 22.4877
R998 GNDA.t152 GNDA.t90 22.4877
R999 GNDA.t128 GNDA.t64 22.4877
R1000 GNDA.t136 GNDA.t34 22.4877
R1001 GNDA.t155 GNDA.t95 22.4877
R1002 GNDA.n142 GNDA.n141 22.4005
R1003 GNDA.n264 GNDA.n263 22.4005
R1004 GNDA.n260 GNDA.n259 22.4005
R1005 GNDA.n225 GNDA.n40 22.4005
R1006 GNDA.n198 GNDA.n197 22.4005
R1007 GNDA.n106 GNDA.n75 22.4005
R1008 GNDA.n15 GNDA.n14 22.4005
R1009 GNDA.n14 GNDA.n13 22.4005
R1010 GNDA.n28 GNDA.n27 21.3338
R1011 GNDA.n31 GNDA.n29 21.3338
R1012 GNDA.n159 GNDA.n158 21.3338
R1013 GNDA.n166 GNDA.n164 21.3338
R1014 GNDA.n173 GNDA.n172 21.3338
R1015 GNDA.n202 GNDA.n199 21.3338
R1016 GNDA.n68 GNDA.n67 21.3338
R1017 GNDA.n71 GNDA.n70 21.3338
R1018 GNDA.n64 GNDA.n63 21.3338
R1019 GNDA.n118 GNDA.n117 21.3338
R1020 GNDA.n9 GNDA.n8 21.3338
R1021 GNDA.n13 GNDA.n12 21.3338
R1022 GNDA.n15 GNDA.n11 21.3338
R1023 GNDA.n16 GNDA.n10 21.3338
R1024 GNDA.n293 GNDA.n290 21.3338
R1025 GNDA.n292 GNDA.n291 21.3338
R1026 GNDA.n21 GNDA.n20 21.3338
R1027 GNDA.n19 GNDA.n18 21.3338
R1028 GNDA.n287 GNDA.n286 21.3338
R1029 GNDA.n288 GNDA.n285 21.3338
R1030 GNDA GNDA.n321 21.221
R1031 GNDA.n194 GNDA.n193 20.3004
R1032 GNDA.n318 GNDA.t230 19.7005
R1033 GNDA.n318 GNDA.t236 19.7005
R1034 GNDA.n316 GNDA.t227 19.7005
R1035 GNDA.n316 GNDA.t3 19.7005
R1036 GNDA.n314 GNDA.t8 19.7005
R1037 GNDA.n314 GNDA.t229 19.7005
R1038 GNDA.n312 GNDA.t226 19.7005
R1039 GNDA.n312 GNDA.t23 19.7005
R1040 GNDA.n310 GNDA.t5 19.7005
R1041 GNDA.n310 GNDA.t81 19.7005
R1042 GNDA.n309 GNDA.t244 19.7005
R1043 GNDA.n309 GNDA.t80 19.7005
R1044 GNDA.n136 GNDA.t63 19.7005
R1045 GNDA.n136 GNDA.t245 19.7005
R1046 GNDA.n134 GNDA.t44 19.7005
R1047 GNDA.n134 GNDA.t45 19.7005
R1048 GNDA.n132 GNDA.t22 19.7005
R1049 GNDA.n132 GNDA.t110 19.7005
R1050 GNDA.n130 GNDA.t70 19.7005
R1051 GNDA.n130 GNDA.t25 19.7005
R1052 GNDA.n128 GNDA.t20 19.7005
R1053 GNDA.n128 GNDA.t26 19.7005
R1054 GNDA.n127 GNDA.t21 19.7005
R1055 GNDA.n127 GNDA.t89 19.7005
R1056 GNDA.n181 GNDA.n155 19.3505
R1057 GNDA.n91 GNDA.n81 19.3505
R1058 GNDA.n300 GNDA.n299 19.288
R1059 GNDA.n200 GNDA.n160 19.1005
R1060 GNDA.n116 GNDA.n115 19.1005
R1061 GNDA.t247 GNDA.n252 18.7399
R1062 GNDA.t2 GNDA.t10 17.2554
R1063 GNDA.t165 GNDA.t53 14.992
R1064 GNDA.t71 GNDA.t6 14.992
R1065 GNDA.t51 GNDA.t58 14.992
R1066 GNDA.t48 GNDA.t62 14.992
R1067 GNDA.t1 GNDA.t246 14.992
R1068 GNDA.t86 GNDA.t177 14.992
R1069 GNDA.t177 GNDA.t59 14.992
R1070 GNDA.t59 GNDA.t17 14.992
R1071 GNDA.t56 GNDA.t142 14.992
R1072 GNDA.t142 GNDA.t15 14.992
R1073 GNDA.t41 GNDA.t118 14.992
R1074 GNDA.t118 GNDA.t55 14.992
R1075 GNDA.t55 GNDA.t233 14.992
R1076 GNDA.t65 GNDA.t138 14.992
R1077 GNDA.t138 GNDA.t243 14.992
R1078 GNDA.t243 GNDA.t180 14.992
R1079 GNDA.t104 GNDA.t116 14.992
R1080 GNDA.t116 GNDA.t12 14.992
R1081 GNDA.t106 GNDA.t132 14.992
R1082 GNDA.t132 GNDA.t93 14.992
R1083 GNDA.t102 GNDA.t122 14.992
R1084 GNDA.t122 GNDA.t207 14.992
R1085 GNDA.t162 GNDA.t146 14.992
R1086 GNDA.t109 GNDA.t120 14.992
R1087 GNDA.t140 GNDA.t159 14.992
R1088 GNDA.t186 GNDA.t72 14.992
R1089 GNDA.t74 GNDA.t247 14.992
R1090 GNDA.t68 GNDA.t237 14.992
R1091 GNDA.t91 GNDA.t88 14.992
R1092 GNDA.t31 GNDA.t47 14.992
R1093 GNDA.t92 GNDA.t46 14.992
R1094 GNDA.t90 GNDA.t49 14.992
R1095 GNDA.t64 GNDA.t195 14.992
R1096 GNDA.n147 GNDA.n53 14.9411
R1097 GNDA.n232 GNDA.n231 14.0505
R1098 GNDA.n124 GNDA.n123 14.0505
R1099 GNDA.n308 GNDA.n307 14.0193
R1100 GNDA.n263 GNDA.n262 13.8005
R1101 GNDA.n226 GNDA.n225 13.8005
R1102 GNDA.n261 GNDA.n260 13.8005
R1103 GNDA.n141 GNDA.n140 13.8005
R1104 GNDA.n156 GNDA.n155 12.8005
R1105 GNDA.n81 GNDA.n80 12.8005
R1106 GNDA.n139 GNDA.n138 11.6255
R1107 GNDA.n268 GNDA.t54 11.2441
R1108 GNDA.t15 GNDA.n41 11.2441
R1109 GNDA.t235 GNDA.t0 11.2441
R1110 GNDA.n304 GNDA.t136 11.2441
R1111 GNDA.t85 GNDA.t77 11.2059
R1112 GNDA.t83 GNDA.t213 11.2059
R1113 GNDA.n235 GNDA.t224 11.2059
R1114 GNDA.t189 GNDA.n110 11.2059
R1115 GNDA.t112 GNDA.t174 11.2059
R1116 GNDA.t29 GNDA.t101 11.2059
R1117 GNDA.t178 GNDA.n38 9.6005
R1118 GNDA.n38 GNDA.t143 9.6005
R1119 GNDA.n205 GNDA.t119 9.6005
R1120 GNDA.n205 GNDA.t139 9.6005
R1121 GNDA.n207 GNDA.t117 9.6005
R1122 GNDA.n207 GNDA.t133 9.6005
R1123 GNDA.n209 GNDA.t123 9.6005
R1124 GNDA.n209 GNDA.t147 9.6005
R1125 GNDA.n211 GNDA.t121 9.6005
R1126 GNDA.n211 GNDA.t141 9.6005
R1127 GNDA.n213 GNDA.t151 9.6005
R1128 GNDA.n213 GNDA.t127 9.6005
R1129 GNDA.n215 GNDA.t149 9.6005
R1130 GNDA.n215 GNDA.t125 9.6005
R1131 GNDA.n217 GNDA.t145 9.6005
R1132 GNDA.n217 GNDA.t135 9.6005
R1133 GNDA.n219 GNDA.t115 9.6005
R1134 GNDA.n219 GNDA.t131 9.6005
R1135 GNDA.n221 GNDA.t153 9.6005
R1136 GNDA.n221 GNDA.t129 9.6005
R1137 GNDA.n223 GNDA.t137 9.6005
R1138 GNDA.n223 GNDA.t156 9.6005
R1139 GNDA.n281 GNDA.n280 9.3005
R1140 GNDA.t241 GNDA.n94 8.6733
R1141 GNDA.n193 GNDA.t33 7.61296
R1142 GNDA.n186 GNDA.t84 7.61296
R1143 GNDA.n308 GNDA.n1 5.03175
R1144 GNDA.n138 GNDA.n1 4.90675
R1145 GNDA.n280 GNDA.n1 4.7505
R1146 GNDA.n279 GNDA.n277 4.5005
R1147 GNDA.n227 GNDA.n0 4.5005
R1148 GNDA.n321 GNDA.n320 4.5005
R1149 GNDA.t201 GNDA.n56 3.74837
R1150 GNDA.n54 GNDA.t238 3.74837
R1151 GNDA.t6 GNDA.n267 3.74837
R1152 GNDA.n42 GNDA.t48 3.74837
R1153 GNDA.n41 GNDA.t240 3.74837
R1154 GNDA.n284 GNDA.t183 3.74837
R1155 GNDA.n256 GNDA.t52 3.74837
R1156 GNDA.t24 GNDA.t235 3.74837
R1157 GNDA.t219 GNDA.t216 3.73564
R1158 GNDA.n102 GNDA.t234 3.73564
R1159 GNDA.n101 GNDA.t100 3.73564
R1160 GNDA.t204 GNDA.t168 3.73564
R1161 GNDA.n320 GNDA.n308 3.6255
R1162 GNDA.n125 GNDA.t28 3.42907
R1163 GNDA.n125 GNDA.t30 3.42907
R1164 GNDA.n228 GNDA.t78 3.42907
R1165 GNDA.n228 GNDA.t76 3.42907
R1166 GNDA.n230 GNDA.t38 3.42907
R1167 GNDA.n230 GNDA.t36 3.42907
R1168 GNDA.n58 GNDA.t98 3.42907
R1169 GNDA.n58 GNDA.t61 3.42907
R1170 GNDA.n183 GNDA.t33 2.53799
R1171 GNDA.t113 GNDA.n184 2.53799
R1172 GNDA.n321 GNDA.n0 2.5005
R1173 GNDA.n229 GNDA.n227 2.063
R1174 GNDA.n139 GNDA.n126 1.813
R1175 GNDA.n227 GNDA.n226 1.78175
R1176 GNDA.n140 GNDA.n139 1.78175
R1177 GNDA.n262 GNDA.n261 1.21925
R1178 GNDA.n262 GNDA.n36 0.6255
R1179 GNDA.n88 GNDA.t7 0.578687
R1180 GNDA.n277 GNDA.n276 0.563
R1181 GNDA.n277 GNDA.n273 0.563
R1182 GNDA.n313 GNDA.n311 0.563
R1183 GNDA.n315 GNDA.n313 0.563
R1184 GNDA.n317 GNDA.n315 0.563
R1185 GNDA.n319 GNDA.n317 0.563
R1186 GNDA.n131 GNDA.n129 0.563
R1187 GNDA.n133 GNDA.n131 0.563
R1188 GNDA.n135 GNDA.n133 0.563
R1189 GNDA.n137 GNDA.n135 0.563
R1190 GNDA.n224 GNDA.n222 0.563
R1191 GNDA.n222 GNDA.n220 0.563
R1192 GNDA.n220 GNDA.n218 0.563
R1193 GNDA.n218 GNDA.n216 0.563
R1194 GNDA.n216 GNDA.n214 0.563
R1195 GNDA.n214 GNDA.n212 0.563
R1196 GNDA.n212 GNDA.n210 0.563
R1197 GNDA.n210 GNDA.n208 0.563
R1198 GNDA.n208 GNDA.n206 0.563
R1199 GNDA.n206 GNDA.n37 0.563
R1200 GNDA.n188 GNDA.t2 0.507997
R1201 GNDA.n231 GNDA.n229 0.5005
R1202 GNDA.n126 GNDA.n124 0.5005
R1203 GNDA.n226 GNDA.n224 0.28175
R1204 GNDA.n280 GNDA.n279 0.2505
R1205 GNDA.n261 GNDA.n37 0.2505
R1206 GNDA.n140 GNDA.n36 0.2505
R1207 V_p.n22 V_p.n0 237.327
R1208 V_p.n32 V_p.t37 202.407
R1209 V_p.n11 V_p.n9 118.168
R1210 V_p.n4 V_p.n2 117.831
R1211 V_p.n17 V_p.n16 117.269
R1212 V_p.n15 V_p.n14 117.269
R1213 V_p.n13 V_p.n12 117.269
R1214 V_p.n11 V_p.n10 117.269
R1215 V_p.n8 V_p.n7 117.269
R1216 V_p.n6 V_p.n5 117.269
R1217 V_p.n4 V_p.n3 117.269
R1218 V_p.n19 V_p.n1 113.136
R1219 V_p.n38 V_p.n37 99.6482
R1220 V_p.n37 V_p.n36 99.0845
R1221 V_p.n35 V_p.n34 99.0845
R1222 V_p.n30 V_p.n29 99.0845
R1223 V_p.n28 V_p.n27 99.0845
R1224 V_p.n26 V_p.n25 99.0845
R1225 V_p.n24 V_p.n23 99.0845
R1226 V_p.n32 V_p.n31 94.5845
R1227 V_p.n21 V_p.n20 94.5845
R1228 V_p.n0 V_p.t38 24.0005
R1229 V_p.n0 V_p.t35 24.0005
R1230 V_p.n16 V_p.t12 16.0005
R1231 V_p.n16 V_p.t11 16.0005
R1232 V_p.n14 V_p.t14 16.0005
R1233 V_p.n14 V_p.t4 16.0005
R1234 V_p.n12 V_p.t3 16.0005
R1235 V_p.n12 V_p.t15 16.0005
R1236 V_p.n10 V_p.t13 16.0005
R1237 V_p.n10 V_p.t10 16.0005
R1238 V_p.n9 V_p.t5 16.0005
R1239 V_p.n9 V_p.t16 16.0005
R1240 V_p.n7 V_p.t40 16.0005
R1241 V_p.n7 V_p.t2 16.0005
R1242 V_p.n5 V_p.t7 16.0005
R1243 V_p.n5 V_p.t6 16.0005
R1244 V_p.n3 V_p.t8 16.0005
R1245 V_p.n3 V_p.t0 16.0005
R1246 V_p.n2 V_p.t1 16.0005
R1247 V_p.n2 V_p.t9 16.0005
R1248 V_p.n1 V_p.t39 16.0005
R1249 V_p.n1 V_p.t36 16.0005
R1250 V_p.n36 V_p.t26 9.6005
R1251 V_p.n36 V_p.t17 9.6005
R1252 V_p.n34 V_p.t21 9.6005
R1253 V_p.n34 V_p.t30 9.6005
R1254 V_p.n31 V_p.t23 9.6005
R1255 V_p.n31 V_p.t32 9.6005
R1256 V_p.n29 V_p.t28 9.6005
R1257 V_p.n29 V_p.t33 9.6005
R1258 V_p.n27 V_p.t31 9.6005
R1259 V_p.n27 V_p.t20 9.6005
R1260 V_p.n25 V_p.t25 9.6005
R1261 V_p.n25 V_p.t22 9.6005
R1262 V_p.n23 V_p.t27 9.6005
R1263 V_p.n23 V_p.t18 9.6005
R1264 V_p.n20 V_p.t29 9.6005
R1265 V_p.n20 V_p.t19 9.6005
R1266 V_p.n38 V_p.t24 9.6005
R1267 V_p.t34 V_p.n38 9.6005
R1268 V_p.n19 V_p.n18 4.5005
R1269 V_p.n22 V_p.n21 4.5005
R1270 V_p.n33 V_p.n32 4.5005
R1271 V_p.n18 V_p.n17 3.65675
R1272 V_p.n21 V_p.n19 1.28175
R1273 V_p.n13 V_p.n11 0.563
R1274 V_p.n15 V_p.n13 0.563
R1275 V_p.n17 V_p.n15 0.563
R1276 V_p.n6 V_p.n4 0.563
R1277 V_p.n8 V_p.n6 0.563
R1278 V_p.n24 V_p.n22 0.563
R1279 V_p.n26 V_p.n24 0.563
R1280 V_p.n28 V_p.n26 0.563
R1281 V_p.n30 V_p.n28 0.563
R1282 V_p.n33 V_p.n30 0.563
R1283 V_p.n35 V_p.n33 0.563
R1284 V_p.n37 V_p.n35 0.563
R1285 V_p.n18 V_p.n8 0.53175
R1286 V_err_amp_ref.n1 V_err_amp_ref.t9 323.491
R1287 V_err_amp_ref.n4 V_err_amp_ref.t0 322.692
R1288 V_err_amp_ref.n7 V_err_amp_ref.t4 270.591
R1289 V_err_amp_ref.n5 V_err_amp_ref.t1 270.591
R1290 V_err_amp_ref.n2 V_err_amp_ref.t2 270.591
R1291 V_err_amp_ref.n0 V_err_amp_ref.t7 270.591
R1292 V_err_amp_ref.n8 V_err_amp_ref.n7 233.374
R1293 V_err_amp_ref.n6 V_err_amp_ref.n5 233.374
R1294 V_err_amp_ref.n3 V_err_amp_ref.n2 233.374
R1295 V_err_amp_ref.n1 V_err_amp_ref.n0 233.374
R1296 V_err_amp_ref.n7 V_err_amp_ref.t8 129.24
R1297 V_err_amp_ref.n5 V_err_amp_ref.t5 129.24
R1298 V_err_amp_ref.n2 V_err_amp_ref.t6 129.24
R1299 V_err_amp_ref.n0 V_err_amp_ref.t3 129.24
R1300 V_err_amp_ref.n4 V_err_amp_ref.n3 3.688
R1301 V_err_amp_ref V_err_amp_ref.n8 3.2505
R1302 V_err_amp_ref.n3 V_err_amp_ref.n1 1.2755
R1303 V_err_amp_ref.n8 V_err_amp_ref.n6 1.2755
R1304 V_err_amp_ref.n6 V_err_amp_ref.n4 0.8005
R1305 V_err_mir_p.n1 V_err_mir_p.n8 632.186
R1306 V_err_mir_p.n1 V_err_mir_p.n11 630.264
R1307 V_err_mir_p.n1 V_err_mir_p.n10 630.264
R1308 V_err_mir_p.n1 V_err_mir_p.n9 630.264
R1309 V_err_mir_p.n0 V_err_mir_p.n5 628.003
R1310 V_err_mir_p.n0 V_err_mir_p.n3 628.003
R1311 V_err_mir_p.n0 V_err_mir_p.n4 626.753
R1312 V_err_mir_p.n12 V_err_mir_p.n0 626.753
R1313 V_err_mir_p.n2 V_err_mir_p.n7 625.756
R1314 V_err_mir_p.n2 V_err_mir_p.n6 622.231
R1315 V_err_mir_p.n6 V_err_mir_p.t19 78.8005
R1316 V_err_mir_p.n6 V_err_mir_p.t16 78.8005
R1317 V_err_mir_p.n11 V_err_mir_p.t8 78.8005
R1318 V_err_mir_p.n11 V_err_mir_p.t13 78.8005
R1319 V_err_mir_p.n10 V_err_mir_p.t15 78.8005
R1320 V_err_mir_p.n10 V_err_mir_p.t6 78.8005
R1321 V_err_mir_p.n9 V_err_mir_p.t9 78.8005
R1322 V_err_mir_p.n9 V_err_mir_p.t14 78.8005
R1323 V_err_mir_p.n8 V_err_mir_p.t11 78.8005
R1324 V_err_mir_p.n8 V_err_mir_p.t18 78.8005
R1325 V_err_mir_p.n7 V_err_mir_p.t12 78.8005
R1326 V_err_mir_p.n7 V_err_mir_p.t4 78.8005
R1327 V_err_mir_p.n5 V_err_mir_p.t1 78.8005
R1328 V_err_mir_p.n5 V_err_mir_p.t2 78.8005
R1329 V_err_mir_p.n4 V_err_mir_p.t7 78.8005
R1330 V_err_mir_p.n4 V_err_mir_p.t17 78.8005
R1331 V_err_mir_p.n3 V_err_mir_p.t10 78.8005
R1332 V_err_mir_p.n3 V_err_mir_p.t3 78.8005
R1333 V_err_mir_p.n12 V_err_mir_p.t5 78.8005
R1334 V_err_mir_p.t0 V_err_mir_p.n12 78.8005
R1335 V_err_mir_p.n0 V_err_mir_p.n2 7.94147
R1336 V_err_mir_p.n2 V_err_mir_p.n1 6.188
R1337 V_err_gate.n21 V_err_gate.n19 630.857
R1338 V_err_gate.n24 V_err_gate.n22 627.316
R1339 V_err_gate.n26 V_err_gate.n25 626.784
R1340 V_err_gate.n24 V_err_gate.n23 626.784
R1341 V_err_gate.n21 V_err_gate.n20 626.784
R1342 V_err_gate.n29 V_err_gate.n28 585
R1343 V_err_gate.n16 V_err_gate.t18 289.2
R1344 V_err_gate.n0 V_err_gate.t14 289.2
R1345 V_err_gate.n17 V_err_gate.n16 176.733
R1346 V_err_gate.n1 V_err_gate.n0 176.733
R1347 V_err_gate.n2 V_err_gate.n1 176.733
R1348 V_err_gate.n3 V_err_gate.n2 176.733
R1349 V_err_gate.n4 V_err_gate.n3 176.733
R1350 V_err_gate.n5 V_err_gate.n4 176.733
R1351 V_err_gate.n6 V_err_gate.n5 176.733
R1352 V_err_gate.n7 V_err_gate.n6 176.733
R1353 V_err_gate.n8 V_err_gate.n7 176.733
R1354 V_err_gate.n9 V_err_gate.n8 176.733
R1355 V_err_gate.n10 V_err_gate.n9 176.733
R1356 V_err_gate.n11 V_err_gate.n10 176.733
R1357 V_err_gate.n12 V_err_gate.n11 176.733
R1358 V_err_gate.n13 V_err_gate.n12 176.733
R1359 V_err_gate.n14 V_err_gate.n13 176.733
R1360 V_err_gate.n15 V_err_gate.n14 176.733
R1361 V_err_gate V_err_gate.n18 162.214
R1362 V_err_gate.n17 V_err_gate.t15 112.468
R1363 V_err_gate.n16 V_err_gate.t26 112.468
R1364 V_err_gate.n0 V_err_gate.t25 112.468
R1365 V_err_gate.n1 V_err_gate.t17 112.468
R1366 V_err_gate.n2 V_err_gate.t27 112.468
R1367 V_err_gate.n3 V_err_gate.t23 112.468
R1368 V_err_gate.n4 V_err_gate.t13 112.468
R1369 V_err_gate.n5 V_err_gate.t24 112.468
R1370 V_err_gate.n6 V_err_gate.t16 112.468
R1371 V_err_gate.n7 V_err_gate.t19 112.468
R1372 V_err_gate.n8 V_err_gate.t29 112.468
R1373 V_err_gate.n9 V_err_gate.t21 112.468
R1374 V_err_gate.n10 V_err_gate.t31 112.468
R1375 V_err_gate.n11 V_err_gate.t22 112.468
R1376 V_err_gate.n12 V_err_gate.t12 112.468
R1377 V_err_gate.n13 V_err_gate.t28 112.468
R1378 V_err_gate.n14 V_err_gate.t20 112.468
R1379 V_err_gate.n15 V_err_gate.t30 112.468
R1380 V_err_gate.n28 V_err_gate.t5 78.8005
R1381 V_err_gate.n28 V_err_gate.t7 78.8005
R1382 V_err_gate.n25 V_err_gate.t1 78.8005
R1383 V_err_gate.n25 V_err_gate.t3 78.8005
R1384 V_err_gate.n23 V_err_gate.t4 78.8005
R1385 V_err_gate.n23 V_err_gate.t6 78.8005
R1386 V_err_gate.n22 V_err_gate.t11 78.8005
R1387 V_err_gate.n22 V_err_gate.t9 78.8005
R1388 V_err_gate.n20 V_err_gate.t0 78.8005
R1389 V_err_gate.n20 V_err_gate.t2 78.8005
R1390 V_err_gate.n19 V_err_gate.t10 78.8005
R1391 V_err_gate.n19 V_err_gate.t8 78.8005
R1392 V_err_gate.n18 V_err_gate.n17 49.8072
R1393 V_err_gate.n18 V_err_gate.n15 49.8072
R1394 V_err_gate.n29 V_err_gate.n27 41.7838
R1395 V_err_gate V_err_gate.n29 39.8443
R1396 V_err_gate.n26 V_err_gate.n24 0.59425
R1397 V_err_gate.n27 V_err_gate.n21 0.59425
R1398 V_err_gate.n27 V_err_gate.n26 0.53175
R1399 VDDA.n141 VDDA.n137 4605
R1400 VDDA.n141 VDDA.n138 4605
R1401 VDDA.n42 VDDA.n28 4605
R1402 VDDA.n44 VDDA.n28 4605
R1403 VDDA.n206 VDDA.n182 4590
R1404 VDDA.n208 VDDA.n182 4590
R1405 VDDA.n208 VDDA.n183 4590
R1406 VDDA.n206 VDDA.n183 4590
R1407 VDDA.n143 VDDA.n137 4575
R1408 VDDA.n143 VDDA.n138 4575
R1409 VDDA.n42 VDDA.n29 4575
R1410 VDDA.n44 VDDA.n29 4575
R1411 VDDA.n101 VDDA.n94 4020
R1412 VDDA.n103 VDDA.n94 4020
R1413 VDDA.n101 VDDA.n100 4020
R1414 VDDA.n103 VDDA.n100 4020
R1415 VDDA.n77 VDDA.n70 4020
R1416 VDDA.n79 VDDA.n70 4020
R1417 VDDA.n77 VDDA.n76 4020
R1418 VDDA.n79 VDDA.n76 4020
R1419 VDDA.n121 VDDA.n114 3390
R1420 VDDA.n123 VDDA.n114 3390
R1421 VDDA.n121 VDDA.n120 3390
R1422 VDDA.n123 VDDA.n120 3390
R1423 VDDA.n21 VDDA.n14 3390
R1424 VDDA.n23 VDDA.n14 3390
R1425 VDDA.n21 VDDA.n20 3390
R1426 VDDA.n23 VDDA.n20 3390
R1427 VDDA.n230 VDDA.n221 3060
R1428 VDDA.n230 VDDA.n222 2970
R1429 VDDA.n163 VDDA.n157 2940
R1430 VDDA.n165 VDDA.n157 2940
R1431 VDDA.n165 VDDA.n162 2940
R1432 VDDA.n163 VDDA.n162 2940
R1433 VDDA.n171 VDDA.n152 2940
R1434 VDDA.n173 VDDA.n152 2940
R1435 VDDA.n173 VDDA.n170 2940
R1436 VDDA.n171 VDDA.n170 2940
R1437 VDDA.n232 VDDA.n221 2820
R1438 VDDA.n232 VDDA.n222 2730
R1439 VDDA.n135 VDDA.t119 1216.42
R1440 VDDA.n146 VDDA.t113 1216.42
R1441 VDDA.n39 VDDA.t159 1216.42
R1442 VDDA.n47 VDDA.t171 1216.42
R1443 VDDA.n159 VDDA.t152 689.4
R1444 VDDA.n158 VDDA.t158 689.4
R1445 VDDA.n154 VDDA.t139 689.4
R1446 VDDA.n153 VDDA.t145 689.4
R1447 VDDA.n218 VDDA.t142 675.274
R1448 VDDA.n219 VDDA.t149 675.274
R1449 VDDA.n202 VDDA.t136 663.801
R1450 VDDA.n212 VDDA.t124 663.801
R1451 VDDA.n97 VDDA.t131 660.109
R1452 VDDA.n95 VDDA.t153 660.109
R1453 VDDA.n73 VDDA.t128 660.109
R1454 VDDA.n71 VDDA.t177 660.109
R1455 VDDA.n223 VDDA.t170 634.25
R1456 VDDA.n238 VDDA.t164 634.25
R1457 VDDA.n216 VDDA.n215 632.933
R1458 VDDA.n225 VDDA.n224 632.933
R1459 VDDA.n241 VDDA.n240 631.227
R1460 VDDA.n179 VDDA.n178 626.534
R1461 VDDA.n185 VDDA.n184 626.534
R1462 VDDA.n187 VDDA.n186 626.534
R1463 VDDA.n189 VDDA.n188 626.534
R1464 VDDA.n191 VDDA.n190 626.534
R1465 VDDA.n193 VDDA.n192 626.534
R1466 VDDA.n195 VDDA.n194 626.534
R1467 VDDA.n197 VDDA.n196 626.534
R1468 VDDA.n199 VDDA.n198 626.534
R1469 VDDA.n201 VDDA.n200 626.534
R1470 VDDA.n117 VDDA.t116 573.75
R1471 VDDA.n115 VDDA.t125 573.75
R1472 VDDA.n17 VDDA.t165 573.75
R1473 VDDA.n15 VDDA.t174 573.75
R1474 VDDA.n140 VDDA.n112 491.2
R1475 VDDA.n140 VDDA.n139 491.2
R1476 VDDA.n45 VDDA.n27 491.2
R1477 VDDA.n41 VDDA.n27 491.2
R1478 VDDA.n205 VDDA.n181 489.601
R1479 VDDA.n209 VDDA.n181 489.601
R1480 VDDA.n105 VDDA.n104 428.8
R1481 VDDA.n105 VDDA.n93 428.8
R1482 VDDA.n81 VDDA.n80 428.8
R1483 VDDA.n81 VDDA.n69 428.8
R1484 VDDA.t141 VDDA.t163 392.065
R1485 VDDA.t135 VDDA.n206 389.375
R1486 VDDA.n208 VDDA.t123 389.375
R1487 VDDA.t138 VDDA.n170 389.375
R1488 VDDA.t144 VDDA.n152 389.375
R1489 VDDA.n204 VDDA.n180 387.2
R1490 VDDA.n210 VDDA.n180 387.2
R1491 VDDA.t151 VDDA.n162 384.168
R1492 VDDA.t157 VDDA.n157 384.168
R1493 VDDA.t169 VDDA.n230 363.93
R1494 VDDA.n232 VDDA.t147 363.93
R1495 VDDA.n125 VDDA.n124 355.2
R1496 VDDA.n125 VDDA.n113 355.2
R1497 VDDA.n25 VDDA.n24 355.2
R1498 VDDA.n25 VDDA.n13 355.2
R1499 VDDA.n227 VDDA.t168 334.759
R1500 VDDA.n237 VDDA.t162 334.759
R1501 VDDA.n203 VDDA.t134 332.75
R1502 VDDA.n211 VDDA.t122 332.75
R1503 VDDA.n159 VDDA.t150 332.75
R1504 VDDA.n158 VDDA.t156 332.75
R1505 VDDA.n154 VDDA.t137 332.75
R1506 VDDA.n153 VDDA.t143 332.75
R1507 VDDA.t168 VDDA.n226 326.726
R1508 VDDA.n229 VDDA.n220 326.401
R1509 VDDA.n218 VDDA.t140 314.274
R1510 VDDA.n219 VDDA.t146 314.274
R1511 VDDA.n161 VDDA.n156 313.601
R1512 VDDA.n168 VDDA.n156 307.2
R1513 VDDA.n176 VDDA.n151 307.2
R1514 VDDA.n169 VDDA.n151 307.2
R1515 VDDA.n233 VDDA.n220 300.8
R1516 VDDA.t117 VDDA.n121 285.815
R1517 VDDA.n123 VDDA.t126 285.815
R1518 VDDA.t166 VDDA.n21 285.815
R1519 VDDA.n23 VDDA.t175 285.815
R1520 VDDA.n117 VDDA.t118 277.916
R1521 VDDA.n115 VDDA.t127 277.916
R1522 VDDA.n17 VDDA.t167 277.916
R1523 VDDA.n15 VDDA.t176 277.916
R1524 VDDA.n145 VDDA.n112 276.8
R1525 VDDA.n139 VDDA.n136 276.8
R1526 VDDA.n46 VDDA.n45 276.8
R1527 VDDA.n41 VDDA.n40 276.8
R1528 VDDA.t132 VDDA.n101 239.915
R1529 VDDA.n103 VDDA.t154 239.915
R1530 VDDA.t129 VDDA.n77 239.915
R1531 VDDA.n79 VDDA.t178 239.915
R1532 VDDA.n99 VDDA.n98 230.4
R1533 VDDA.n99 VDDA.n96 230.4
R1534 VDDA.n75 VDDA.n74 230.4
R1535 VDDA.n75 VDDA.n72 230.4
R1536 VDDA.n166 VDDA.n160 211.201
R1537 VDDA.n167 VDDA.n166 211.201
R1538 VDDA.n175 VDDA.n174 211.201
R1539 VDDA.n119 VDDA.n118 211.201
R1540 VDDA.n119 VDDA.n116 211.201
R1541 VDDA.n19 VDDA.n18 211.201
R1542 VDDA.n19 VDDA.n16 211.201
R1543 VDDA.n228 VDDA.n217 208
R1544 VDDA.n145 VDDA.n144 204.8
R1545 VDDA.n144 VDDA.n136 204.8
R1546 VDDA.n40 VDDA.n26 204.8
R1547 VDDA.n46 VDDA.n26 204.8
R1548 VDDA.n174 VDDA.n155 202.971
R1549 VDDA.n104 VDDA.n96 198.4
R1550 VDDA.n98 VDDA.n93 198.4
R1551 VDDA.n80 VDDA.n72 198.4
R1552 VDDA.n74 VDDA.n69 198.4
R1553 VDDA.t214 VDDA.t135 186.607
R1554 VDDA.t192 VDDA.t214 186.607
R1555 VDDA.t208 VDDA.t192 186.607
R1556 VDDA.t182 VDDA.t208 186.607
R1557 VDDA.t196 VDDA.t182 186.607
R1558 VDDA.t216 VDDA.t196 186.607
R1559 VDDA.t194 VDDA.t216 186.607
R1560 VDDA.t210 VDDA.t194 186.607
R1561 VDDA.t206 VDDA.t210 186.607
R1562 VDDA.t186 VDDA.t206 186.607
R1563 VDDA.t180 VDDA.t200 186.607
R1564 VDDA.t198 VDDA.t180 186.607
R1565 VDDA.t218 VDDA.t198 186.607
R1566 VDDA.t188 VDDA.t218 186.607
R1567 VDDA.t204 VDDA.t188 186.607
R1568 VDDA.t184 VDDA.t204 186.607
R1569 VDDA.t212 VDDA.t184 186.607
R1570 VDDA.t190 VDDA.t212 186.607
R1571 VDDA.t202 VDDA.t190 186.607
R1572 VDDA.t123 VDDA.t202 186.607
R1573 VDDA.t233 VDDA.t138 186.607
R1574 VDDA.t38 VDDA.t233 186.607
R1575 VDDA.t104 VDDA.t38 186.607
R1576 VDDA.t228 VDDA.t104 186.607
R1577 VDDA.t232 VDDA.t228 186.607
R1578 VDDA.t72 VDDA.t105 186.607
R1579 VDDA.t105 VDDA.t225 186.607
R1580 VDDA.t225 VDDA.t229 186.607
R1581 VDDA.t229 VDDA.t249 186.607
R1582 VDDA.t249 VDDA.t144 186.607
R1583 VDDA.t224 VDDA.t151 183.333
R1584 VDDA.t68 VDDA.t224 183.333
R1585 VDDA.t53 VDDA.t68 183.333
R1586 VDDA.t230 VDDA.t53 183.333
R1587 VDDA.t226 VDDA.t230 183.333
R1588 VDDA.t49 VDDA.t69 183.333
R1589 VDDA.t69 VDDA.t227 183.333
R1590 VDDA.t227 VDDA.t231 183.333
R1591 VDDA.t231 VDDA.t50 183.333
R1592 VDDA.t50 VDDA.t157 183.333
R1593 VDDA.t91 VDDA.t169 180.952
R1594 VDDA.t36 VDDA.t91 180.952
R1595 VDDA.t66 VDDA.t36 180.952
R1596 VDDA.t60 VDDA.t66 180.952
R1597 VDDA.t102 VDDA.t141 180.952
R1598 VDDA.t147 VDDA.t102 180.952
R1599 VDDA.n134 VDDA.t121 178.124
R1600 VDDA.n147 VDDA.t115 178.124
R1601 VDDA.n38 VDDA.t161 178.124
R1602 VDDA.n48 VDDA.t173 178.124
R1603 VDDA.n231 VDDA.t60 165.874
R1604 VDDA.t114 VDDA.n137 161.817
R1605 VDDA.t120 VDDA.n138 161.817
R1606 VDDA.t160 VDDA.n42 161.817
R1607 VDDA.n44 VDDA.t172 161.817
R1608 VDDA.n91 VDDA.n89 160.428
R1609 VDDA.n88 VDDA.n86 160.428
R1610 VDDA.n67 VDDA.n65 160.428
R1611 VDDA.n64 VDDA.n62 160.428
R1612 VDDA.n91 VDDA.n90 159.803
R1613 VDDA.n88 VDDA.n87 159.803
R1614 VDDA.n67 VDDA.n66 159.803
R1615 VDDA.n64 VDDA.n63 159.803
R1616 VDDA.n97 VDDA.t133 155.125
R1617 VDDA.n95 VDDA.t155 155.125
R1618 VDDA.n73 VDDA.t130 155.125
R1619 VDDA.n71 VDDA.t179 155.125
R1620 VDDA.n134 VDDA.n133 151.882
R1621 VDDA.n38 VDDA.n37 151.882
R1622 VDDA.n148 VDDA.n147 151.321
R1623 VDDA.n49 VDDA.n48 151.321
R1624 VDDA.n124 VDDA.n116 150.4
R1625 VDDA.n118 VDDA.n113 150.4
R1626 VDDA.n24 VDDA.n16 150.4
R1627 VDDA.n18 VDDA.n13 150.4
R1628 VDDA.n107 VDDA.n106 146.002
R1629 VDDA.n83 VDDA.n82 146.002
R1630 VDDA.n111 VDDA.n110 145.429
R1631 VDDA.n127 VDDA.n126 145.429
R1632 VDDA.n129 VDDA.n128 145.429
R1633 VDDA.n131 VDDA.n130 145.429
R1634 VDDA.n133 VDDA.n132 145.429
R1635 VDDA.n12 VDDA.n11 145.429
R1636 VDDA.n31 VDDA.n30 145.429
R1637 VDDA.n33 VDDA.n32 145.429
R1638 VDDA.n35 VDDA.n34 145.429
R1639 VDDA.n37 VDDA.n36 145.429
R1640 VDDA.n147 VDDA.n146 135.387
R1641 VDDA.n135 VDDA.n134 135.387
R1642 VDDA.n48 VDDA.n47 135.387
R1643 VDDA.n39 VDDA.n38 135.387
R1644 VDDA.t74 VDDA.t117 121.513
R1645 VDDA.t4 VDDA.t74 121.513
R1646 VDDA.t77 VDDA.t4 121.513
R1647 VDDA.t236 VDDA.t77 121.513
R1648 VDDA.t22 VDDA.t236 121.513
R1649 VDDA.t239 VDDA.t11 121.513
R1650 VDDA.t237 VDDA.t239 121.513
R1651 VDDA.t0 VDDA.t237 121.513
R1652 VDDA.t240 VDDA.t0 121.513
R1653 VDDA.t126 VDDA.t240 121.513
R1654 VDDA.t256 VDDA.t166 121.513
R1655 VDDA.t40 VDDA.t256 121.513
R1656 VDDA.t41 VDDA.t40 121.513
R1657 VDDA.t21 VDDA.t41 121.513
R1658 VDDA.t108 VDDA.t21 121.513
R1659 VDDA.t27 VDDA.t65 121.513
R1660 VDDA.t19 VDDA.t27 121.513
R1661 VDDA.t28 VDDA.t19 121.513
R1662 VDDA.t20 VDDA.t28 121.513
R1663 VDDA.t175 VDDA.t20 121.513
R1664 VDDA.n235 VDDA.n234 115.201
R1665 VDDA.n229 VDDA.n228 108.8
R1666 VDDA.n234 VDDA.n233 108.8
R1667 VDDA.n205 VDDA.n204 102.4
R1668 VDDA.n210 VDDA.n209 102.4
R1669 VDDA.n161 VDDA.n160 102.4
R1670 VDDA.t23 VDDA.t132 98.2764
R1671 VDDA.t247 VDDA.t23 98.2764
R1672 VDDA.t43 VDDA.t247 98.2764
R1673 VDDA.t99 VDDA.t43 98.2764
R1674 VDDA.t7 VDDA.t99 98.2764
R1675 VDDA.t31 VDDA.t82 98.2764
R1676 VDDA.t243 VDDA.t31 98.2764
R1677 VDDA.t51 VDDA.t243 98.2764
R1678 VDDA.t84 VDDA.t51 98.2764
R1679 VDDA.t154 VDDA.t84 98.2764
R1680 VDDA.t58 VDDA.t129 98.2764
R1681 VDDA.t86 VDDA.t58 98.2764
R1682 VDDA.t254 VDDA.t86 98.2764
R1683 VDDA.t106 VDDA.t254 98.2764
R1684 VDDA.t16 VDDA.t106 98.2764
R1685 VDDA.t252 VDDA.t250 98.2764
R1686 VDDA.t241 VDDA.t252 98.2764
R1687 VDDA.t47 VDDA.t241 98.2764
R1688 VDDA.t54 VDDA.t47 98.2764
R1689 VDDA.t178 VDDA.t54 98.2764
R1690 VDDA.n52 VDDA.n50 97.4034
R1691 VDDA.n2 VDDA.n0 97.4034
R1692 VDDA.n60 VDDA.n59 96.8409
R1693 VDDA.n58 VDDA.n57 96.8409
R1694 VDDA.n56 VDDA.n55 96.8409
R1695 VDDA.n54 VDDA.n53 96.8409
R1696 VDDA.n52 VDDA.n51 96.8409
R1697 VDDA.n10 VDDA.n9 96.8409
R1698 VDDA.n8 VDDA.n7 96.8409
R1699 VDDA.n6 VDDA.n5 96.8409
R1700 VDDA.n4 VDDA.n3 96.8409
R1701 VDDA.n2 VDDA.n1 96.8409
R1702 VDDA.n168 VDDA.n167 96.0005
R1703 VDDA.n169 VDDA.n155 96.0005
R1704 VDDA.n176 VDDA.n175 96.0005
R1705 VDDA.n207 VDDA.t186 93.3041
R1706 VDDA.t200 VDDA.n207 93.3041
R1707 VDDA.n172 VDDA.t232 93.3041
R1708 VDDA.n172 VDDA.t72 93.3041
R1709 VDDA.n230 VDDA.n229 92.5005
R1710 VDDA.n221 VDDA.n220 92.5005
R1711 VDDA.n231 VDDA.n221 92.5005
R1712 VDDA.n233 VDDA.n232 92.5005
R1713 VDDA.n222 VDDA.n217 92.5005
R1714 VDDA.n231 VDDA.n222 92.5005
R1715 VDDA.n206 VDDA.n205 92.5005
R1716 VDDA.n182 VDDA.n181 92.5005
R1717 VDDA.n207 VDDA.n182 92.5005
R1718 VDDA.n209 VDDA.n208 92.5005
R1719 VDDA.n183 VDDA.n180 92.5005
R1720 VDDA.n207 VDDA.n183 92.5005
R1721 VDDA.n163 VDDA.n156 92.5005
R1722 VDDA.n164 VDDA.n163 92.5005
R1723 VDDA.n162 VDDA.n161 92.5005
R1724 VDDA.n166 VDDA.n165 92.5005
R1725 VDDA.n165 VDDA.n164 92.5005
R1726 VDDA.n168 VDDA.n157 92.5005
R1727 VDDA.n171 VDDA.n151 92.5005
R1728 VDDA.n172 VDDA.n171 92.5005
R1729 VDDA.n170 VDDA.n169 92.5005
R1730 VDDA.n174 VDDA.n173 92.5005
R1731 VDDA.n173 VDDA.n172 92.5005
R1732 VDDA.n176 VDDA.n152 92.5005
R1733 VDDA.n124 VDDA.n123 92.5005
R1734 VDDA.n120 VDDA.n119 92.5005
R1735 VDDA.n122 VDDA.n120 92.5005
R1736 VDDA.n121 VDDA.n113 92.5005
R1737 VDDA.n125 VDDA.n114 92.5005
R1738 VDDA.n122 VDDA.n114 92.5005
R1739 VDDA.n144 VDDA.n143 92.5005
R1740 VDDA.n143 VDDA.n142 92.5005
R1741 VDDA.n141 VDDA.n140 92.5005
R1742 VDDA.n142 VDDA.n141 92.5005
R1743 VDDA.n104 VDDA.n103 92.5005
R1744 VDDA.n100 VDDA.n99 92.5005
R1745 VDDA.n102 VDDA.n100 92.5005
R1746 VDDA.n101 VDDA.n93 92.5005
R1747 VDDA.n105 VDDA.n94 92.5005
R1748 VDDA.n102 VDDA.n94 92.5005
R1749 VDDA.n80 VDDA.n79 92.5005
R1750 VDDA.n76 VDDA.n75 92.5005
R1751 VDDA.n78 VDDA.n76 92.5005
R1752 VDDA.n77 VDDA.n69 92.5005
R1753 VDDA.n81 VDDA.n70 92.5005
R1754 VDDA.n78 VDDA.n70 92.5005
R1755 VDDA.n24 VDDA.n23 92.5005
R1756 VDDA.n20 VDDA.n19 92.5005
R1757 VDDA.n22 VDDA.n20 92.5005
R1758 VDDA.n21 VDDA.n13 92.5005
R1759 VDDA.n25 VDDA.n14 92.5005
R1760 VDDA.n22 VDDA.n14 92.5005
R1761 VDDA.n29 VDDA.n26 92.5005
R1762 VDDA.n43 VDDA.n29 92.5005
R1763 VDDA.n28 VDDA.n27 92.5005
R1764 VDDA.n43 VDDA.n28 92.5005
R1765 VDDA.n164 VDDA.t226 91.6672
R1766 VDDA.n164 VDDA.t49 91.6672
R1767 VDDA.n178 VDDA.t191 78.8005
R1768 VDDA.n178 VDDA.t203 78.8005
R1769 VDDA.n184 VDDA.t185 78.8005
R1770 VDDA.n184 VDDA.t213 78.8005
R1771 VDDA.n186 VDDA.t189 78.8005
R1772 VDDA.n186 VDDA.t205 78.8005
R1773 VDDA.n188 VDDA.t199 78.8005
R1774 VDDA.n188 VDDA.t219 78.8005
R1775 VDDA.n190 VDDA.t201 78.8005
R1776 VDDA.n190 VDDA.t181 78.8005
R1777 VDDA.n192 VDDA.t207 78.8005
R1778 VDDA.n192 VDDA.t187 78.8005
R1779 VDDA.n194 VDDA.t195 78.8005
R1780 VDDA.n194 VDDA.t211 78.8005
R1781 VDDA.n196 VDDA.t197 78.8005
R1782 VDDA.n196 VDDA.t217 78.8005
R1783 VDDA.n198 VDDA.t209 78.8005
R1784 VDDA.n198 VDDA.t183 78.8005
R1785 VDDA.n200 VDDA.t215 78.8005
R1786 VDDA.n200 VDDA.t193 78.8005
R1787 VDDA.t56 VDDA.t114 62.9523
R1788 VDDA.t2 VDDA.t56 62.9523
R1789 VDDA.t93 VDDA.t2 62.9523
R1790 VDDA.t9 VDDA.t93 62.9523
R1791 VDDA.t5 VDDA.t9 62.9523
R1792 VDDA.t75 VDDA.t78 62.9523
R1793 VDDA.t78 VDDA.t45 62.9523
R1794 VDDA.t45 VDDA.t257 62.9523
R1795 VDDA.t257 VDDA.t96 62.9523
R1796 VDDA.t96 VDDA.t120 62.9523
R1797 VDDA.t88 VDDA.t160 62.9523
R1798 VDDA.t234 VDDA.t88 62.9523
R1799 VDDA.t34 VDDA.t234 62.9523
R1800 VDDA.t25 VDDA.t34 62.9523
R1801 VDDA.t245 VDDA.t25 62.9523
R1802 VDDA.t70 VDDA.t13 62.9523
R1803 VDDA.t29 VDDA.t70 62.9523
R1804 VDDA.t111 VDDA.t29 62.9523
R1805 VDDA.t62 VDDA.t111 62.9523
R1806 VDDA.t172 VDDA.t62 62.9523
R1807 VDDA.n240 VDDA.t103 62.5402
R1808 VDDA.n240 VDDA.t148 62.5402
R1809 VDDA.n137 VDDA.n112 61.6672
R1810 VDDA.n139 VDDA.n138 61.6672
R1811 VDDA.n45 VDDA.n44 61.6672
R1812 VDDA.n42 VDDA.n41 61.6672
R1813 VDDA.n122 VDDA.t22 60.7563
R1814 VDDA.t11 VDDA.n122 60.7563
R1815 VDDA.n22 VDDA.t108 60.7563
R1816 VDDA.t65 VDDA.n22 60.7563
R1817 VDDA.n215 VDDA.t67 49.2505
R1818 VDDA.n215 VDDA.t61 49.2505
R1819 VDDA.n224 VDDA.t92 49.2505
R1820 VDDA.n224 VDDA.t37 49.2505
R1821 VDDA.n102 VDDA.t7 49.1384
R1822 VDDA.t82 VDDA.n102 49.1384
R1823 VDDA.n78 VDDA.t16 49.1384
R1824 VDDA.t250 VDDA.n78 49.1384
R1825 VDDA.n239 VDDA.n238 47.9338
R1826 VDDA.n236 VDDA.n235 44.8005
R1827 VDDA.n202 VDDA.n201 42.0963
R1828 VDDA.n213 VDDA.n212 41.5338
R1829 VDDA.n226 VDDA.n223 34.1338
R1830 VDDA.n238 VDDA.n237 32.0005
R1831 VDDA.n227 VDDA.n223 32.0005
R1832 VDDA.n142 VDDA.t5 31.4764
R1833 VDDA.n142 VDDA.t75 31.4764
R1834 VDDA.n43 VDDA.t245 31.4764
R1835 VDDA.t13 VDDA.n43 31.4764
R1836 VDDA.n169 VDDA.n168 28.663
R1837 VDDA.n212 VDDA.n211 25.6005
R1838 VDDA.n203 VDDA.n202 25.6005
R1839 VDDA.n237 VDDA.n236 24.5338
R1840 VDDA.n235 VDDA.n218 24.5338
R1841 VDDA.n234 VDDA.n219 24.5338
R1842 VDDA.n228 VDDA.n227 24.5338
R1843 VDDA VDDA.n242 23.1273
R1844 VDDA.n236 VDDA.n217 22.4005
R1845 VDDA.n211 VDDA.n210 21.3338
R1846 VDDA.n204 VDDA.n203 21.3338
R1847 VDDA.n160 VDDA.n159 21.3338
R1848 VDDA.n167 VDDA.n158 21.3338
R1849 VDDA.n155 VDDA.n154 21.3338
R1850 VDDA.n175 VDDA.n153 21.3338
R1851 VDDA.n118 VDDA.n117 21.3338
R1852 VDDA.n116 VDDA.n115 21.3338
R1853 VDDA.n146 VDDA.n145 21.3338
R1854 VDDA.n136 VDDA.n135 21.3338
R1855 VDDA.n98 VDDA.n97 21.3338
R1856 VDDA.n96 VDDA.n95 21.3338
R1857 VDDA.n74 VDDA.n73 21.3338
R1858 VDDA.n72 VDDA.n71 21.3338
R1859 VDDA.n18 VDDA.n17 21.3338
R1860 VDDA.n16 VDDA.n15 21.3338
R1861 VDDA.n47 VDDA.n46 21.3338
R1862 VDDA.n40 VDDA.n39 21.3338
R1863 VDDA.n61 VDDA.n60 21.1567
R1864 VDDA.n177 VDDA.n176 19.5505
R1865 VDDA.n144 VDDA.n125 19.538
R1866 VDDA.n26 VDDA.n25 19.538
R1867 VDDA.n107 VDDA.n105 19.2005
R1868 VDDA.n83 VDDA.n81 19.2005
R1869 VDDA.n150 VDDA.n10 16.8443
R1870 VDDA.t163 VDDA.n231 15.0799
R1871 VDDA.n226 VDDA.n225 14.4255
R1872 VDDA.n106 VDDA.t8 11.2576
R1873 VDDA.n106 VDDA.t83 11.2576
R1874 VDDA.n90 VDDA.t32 11.2576
R1875 VDDA.n90 VDDA.t244 11.2576
R1876 VDDA.n89 VDDA.t52 11.2576
R1877 VDDA.n89 VDDA.t85 11.2576
R1878 VDDA.n87 VDDA.t44 11.2576
R1879 VDDA.n87 VDDA.t100 11.2576
R1880 VDDA.n86 VDDA.t24 11.2576
R1881 VDDA.n86 VDDA.t248 11.2576
R1882 VDDA.n82 VDDA.t17 11.2576
R1883 VDDA.n82 VDDA.t251 11.2576
R1884 VDDA.n66 VDDA.t253 11.2576
R1885 VDDA.n66 VDDA.t242 11.2576
R1886 VDDA.n65 VDDA.t48 11.2576
R1887 VDDA.n65 VDDA.t55 11.2576
R1888 VDDA.n63 VDDA.t255 11.2576
R1889 VDDA.n63 VDDA.t107 11.2576
R1890 VDDA.n62 VDDA.t59 11.2576
R1891 VDDA.n62 VDDA.t87 11.2576
R1892 VDDA.n108 VDDA.n107 9.3005
R1893 VDDA.n84 VDDA.n83 9.3005
R1894 VDDA.n59 VDDA.t259 8.0005
R1895 VDDA.n59 VDDA.t221 8.0005
R1896 VDDA.n57 VDDA.t64 8.0005
R1897 VDDA.n57 VDDA.t98 8.0005
R1898 VDDA.n55 VDDA.t42 8.0005
R1899 VDDA.n55 VDDA.t15 8.0005
R1900 VDDA.n53 VDDA.t33 8.0005
R1901 VDDA.n53 VDDA.t18 8.0005
R1902 VDDA.n51 VDDA.t110 8.0005
R1903 VDDA.n51 VDDA.t39 8.0005
R1904 VDDA.n50 VDDA.t220 8.0005
R1905 VDDA.n50 VDDA.t109 8.0005
R1906 VDDA.n9 VDDA.t222 8.0005
R1907 VDDA.n9 VDDA.t95 8.0005
R1908 VDDA.n7 VDDA.t90 8.0005
R1909 VDDA.n7 VDDA.t1 8.0005
R1910 VDDA.n5 VDDA.t101 8.0005
R1911 VDDA.n5 VDDA.t12 8.0005
R1912 VDDA.n3 VDDA.t80 8.0005
R1913 VDDA.n3 VDDA.t260 8.0005
R1914 VDDA.n1 VDDA.t73 8.0005
R1915 VDDA.n1 VDDA.t81 8.0005
R1916 VDDA.n0 VDDA.t238 8.0005
R1917 VDDA.n0 VDDA.t223 8.0005
R1918 VDDA.n214 VDDA.n213 7.438
R1919 VDDA.n242 VDDA.n241 7.03175
R1920 VDDA.n110 VDDA.t57 6.56717
R1921 VDDA.n110 VDDA.t3 6.56717
R1922 VDDA.n126 VDDA.t94 6.56717
R1923 VDDA.n126 VDDA.t10 6.56717
R1924 VDDA.n128 VDDA.t6 6.56717
R1925 VDDA.n128 VDDA.t76 6.56717
R1926 VDDA.n130 VDDA.t79 6.56717
R1927 VDDA.n130 VDDA.t46 6.56717
R1928 VDDA.n132 VDDA.t258 6.56717
R1929 VDDA.n132 VDDA.t97 6.56717
R1930 VDDA.n11 VDDA.t112 6.56717
R1931 VDDA.n11 VDDA.t63 6.56717
R1932 VDDA.n30 VDDA.t71 6.56717
R1933 VDDA.n30 VDDA.t30 6.56717
R1934 VDDA.n32 VDDA.t246 6.56717
R1935 VDDA.n32 VDDA.t14 6.56717
R1936 VDDA.n34 VDDA.t35 6.56717
R1937 VDDA.n34 VDDA.t26 6.56717
R1938 VDDA.n36 VDDA.t89 6.56717
R1939 VDDA.n36 VDDA.t235 6.56717
R1940 VDDA.n109 VDDA.n85 6.313
R1941 VDDA.n109 VDDA.n108 5.063
R1942 VDDA.n85 VDDA.n84 5.063
R1943 VDDA.n108 VDDA.n92 4.5005
R1944 VDDA.n84 VDDA.n68 4.5005
R1945 VDDA.n150 VDDA.n149 4.5005
R1946 VDDA.n85 VDDA.n61 3.688
R1947 VDDA.n149 VDDA.n109 3.5005
R1948 VDDA.n214 VDDA.n177 2.813
R1949 VDDA.n242 VDDA.n214 2.563
R1950 VDDA.n177 VDDA.n150 1.46925
R1951 VDDA.n241 VDDA.n239 1.063
R1952 VDDA.n149 VDDA.n148 0.938
R1953 VDDA.n61 VDDA.n49 0.7505
R1954 VDDA.n225 VDDA.n216 0.6255
R1955 VDDA.n239 VDDA.n216 0.6255
R1956 VDDA.n92 VDDA.n91 0.6255
R1957 VDDA.n92 VDDA.n88 0.6255
R1958 VDDA.n68 VDDA.n67 0.6255
R1959 VDDA.n68 VDDA.n64 0.6255
R1960 VDDA.n201 VDDA.n199 0.563
R1961 VDDA.n199 VDDA.n197 0.563
R1962 VDDA.n197 VDDA.n195 0.563
R1963 VDDA.n195 VDDA.n193 0.563
R1964 VDDA.n193 VDDA.n191 0.563
R1965 VDDA.n191 VDDA.n189 0.563
R1966 VDDA.n189 VDDA.n187 0.563
R1967 VDDA.n187 VDDA.n185 0.563
R1968 VDDA.n185 VDDA.n179 0.563
R1969 VDDA.n213 VDDA.n179 0.563
R1970 VDDA.n133 VDDA.n131 0.563
R1971 VDDA.n131 VDDA.n129 0.563
R1972 VDDA.n129 VDDA.n127 0.563
R1973 VDDA.n127 VDDA.n111 0.563
R1974 VDDA.n148 VDDA.n111 0.563
R1975 VDDA.n54 VDDA.n52 0.563
R1976 VDDA.n56 VDDA.n54 0.563
R1977 VDDA.n58 VDDA.n56 0.563
R1978 VDDA.n60 VDDA.n58 0.563
R1979 VDDA.n37 VDDA.n35 0.563
R1980 VDDA.n35 VDDA.n33 0.563
R1981 VDDA.n33 VDDA.n31 0.563
R1982 VDDA.n31 VDDA.n12 0.563
R1983 VDDA.n49 VDDA.n12 0.563
R1984 VDDA.n4 VDDA.n2 0.563
R1985 VDDA.n6 VDDA.n4 0.563
R1986 VDDA.n8 VDDA.n6 0.563
R1987 VDDA.n10 VDDA.n8 0.563
R1988 VD4.n28 VD4.n23 4020
R1989 VD4.n30 VD4.n23 4020
R1990 VD4.n30 VD4.n24 4020
R1991 VD4.n28 VD4.n24 4020
R1992 VD4.n33 VD4.t35 660.109
R1993 VD4.n25 VD4.t32 660.109
R1994 VD4.n27 VD4.n22 428.8
R1995 VD4.n31 VD4.n22 428.8
R1996 VD4.t33 VD4.n28 239.915
R1997 VD4.n30 VD4.t36 239.915
R1998 VD4.n26 VD4.n0 230.4
R1999 VD4.n32 VD4.n0 230.4
R2000 VD4.n27 VD4.n26 198.4
R2001 VD4.n32 VD4.n31 198.4
R2002 VD4.n19 VD4.n17 160.428
R2003 VD4.n6 VD4.n4 160.427
R2004 VD4.n11 VD4.n3 160.427
R2005 VD4.n14 VD4.n2 160.053
R2006 VD4.n19 VD4.n18 159.803
R2007 VD4.n16 VD4.n15 159.803
R2008 VD4.n10 VD4.n9 159.802
R2009 VD4.n8 VD4.n7 159.802
R2010 VD4.n6 VD4.n5 159.802
R2011 VD4.n13 VD4.n12 155.302
R2012 VD4.n25 VD4.t34 155.125
R2013 VD4.t37 VD4.n33 155.125
R2014 VD4.n21 VD4.n1 146.002
R2015 VD4.t0 VD4.t33 98.2764
R2016 VD4.t8 VD4.t0 98.2764
R2017 VD4.t3 VD4.t8 98.2764
R2018 VD4.t5 VD4.t3 98.2764
R2019 VD4.t27 VD4.t5 98.2764
R2020 VD4.t15 VD4.t10 98.2764
R2021 VD4.t22 VD4.t15 98.2764
R2022 VD4.t19 VD4.t22 98.2764
R2023 VD4.t17 VD4.t19 98.2764
R2024 VD4.t36 VD4.t17 98.2764
R2025 VD4.n28 VD4.n27 92.5005
R2026 VD4.n23 VD4.n22 92.5005
R2027 VD4.n29 VD4.n23 92.5005
R2028 VD4.n31 VD4.n30 92.5005
R2029 VD4.n24 VD4.n0 92.5005
R2030 VD4.n29 VD4.n24 92.5005
R2031 VD4.n29 VD4.t27 49.1384
R2032 VD4.t10 VD4.n29 49.1384
R2033 VD4.n26 VD4.n25 21.3338
R2034 VD4.n33 VD4.n32 21.3338
R2035 VD4.n22 VD4.n21 19.2005
R2036 VD4.n21 VD4.n20 13.8005
R2037 VD4.n18 VD4.t16 11.2576
R2038 VD4.n18 VD4.t23 11.2576
R2039 VD4.n17 VD4.t20 11.2576
R2040 VD4.n17 VD4.t18 11.2576
R2041 VD4.n15 VD4.t4 11.2576
R2042 VD4.n15 VD4.t6 11.2576
R2043 VD4.n12 VD4.t14 11.2576
R2044 VD4.n12 VD4.t31 11.2576
R2045 VD4.n9 VD4.t21 11.2576
R2046 VD4.n9 VD4.t2 11.2576
R2047 VD4.n7 VD4.t29 11.2576
R2048 VD4.n7 VD4.t30 11.2576
R2049 VD4.n5 VD4.t26 11.2576
R2050 VD4.n5 VD4.t7 11.2576
R2051 VD4.n4 VD4.t12 11.2576
R2052 VD4.n4 VD4.t25 11.2576
R2053 VD4.n3 VD4.t24 11.2576
R2054 VD4.n3 VD4.t13 11.2576
R2055 VD4.n2 VD4.t1 11.2576
R2056 VD4.n2 VD4.t9 11.2576
R2057 VD4.n1 VD4.t28 11.2576
R2058 VD4.n1 VD4.t11 11.2576
R2059 VD4.n14 VD4.n13 6.188
R2060 VD4.n13 VD4.n11 4.5005
R2061 VD4.n20 VD4.n19 0.6255
R2062 VD4.n8 VD4.n6 0.6255
R2063 VD4.n10 VD4.n8 0.6255
R2064 VD4.n11 VD4.n10 0.6255
R2065 VD4.n20 VD4.n16 0.6255
R2066 VD4.n16 VD4.n14 0.2505
R2067 X.n49 X.t30 1172.87
R2068 X.n43 X.t44 1172.87
R2069 X.n50 X.t27 996.134
R2070 X.n49 X.t43 996.134
R2071 X.n43 X.t48 996.134
R2072 X.n44 X.t34 996.134
R2073 X.n45 X.t51 996.134
R2074 X.n46 X.t37 996.134
R2075 X.n47 X.t25 996.134
R2076 X.n48 X.t40 996.134
R2077 X.n33 X.t38 690.867
R2078 X.n32 X.t53 690.867
R2079 X.n24 X.t28 530.201
R2080 X.n23 X.t42 530.201
R2081 X.n33 X.t52 514.134
R2082 X.n34 X.t35 514.134
R2083 X.n35 X.t49 514.134
R2084 X.n36 X.t32 514.134
R2085 X.n37 X.t46 514.134
R2086 X.n38 X.t31 514.134
R2087 X.n39 X.t45 514.134
R2088 X.n32 X.t29 514.134
R2089 X.n30 X.t33 353.467
R2090 X.n29 X.t50 353.467
R2091 X.n28 X.t36 353.467
R2092 X.n27 X.t54 353.467
R2093 X.n26 X.t39 353.467
R2094 X.n25 X.t26 353.467
R2095 X.n24 X.t41 353.467
R2096 X.n23 X.t47 353.467
R2097 X.n50 X.n49 176.733
R2098 X.n44 X.n43 176.733
R2099 X.n45 X.n44 176.733
R2100 X.n46 X.n45 176.733
R2101 X.n47 X.n46 176.733
R2102 X.n48 X.n47 176.733
R2103 X.n30 X.n29 176.733
R2104 X.n29 X.n28 176.733
R2105 X.n28 X.n27 176.733
R2106 X.n27 X.n26 176.733
R2107 X.n26 X.n25 176.733
R2108 X.n25 X.n24 176.733
R2109 X.n39 X.n38 176.733
R2110 X.n38 X.n37 176.733
R2111 X.n37 X.n36 176.733
R2112 X.n36 X.n35 176.733
R2113 X.n35 X.n34 176.733
R2114 X.n34 X.n33 176.733
R2115 X.n52 X.n51 166.436
R2116 X.n41 X.n31 161.875
R2117 X.n41 X.n40 161.686
R2118 X.n2 X.n0 160.427
R2119 X.n8 X.n7 159.802
R2120 X.n6 X.n5 159.802
R2121 X.n4 X.n3 159.802
R2122 X.n2 X.n1 159.802
R2123 X.n10 X.n9 155.302
R2124 X.n15 X.n13 114.689
R2125 X.n20 X.n12 114.689
R2126 X.n19 X.n18 114.126
R2127 X.n17 X.n16 114.126
R2128 X.n15 X.n14 114.126
R2129 X.n21 X.n11 109.626
R2130 X.n51 X.n50 51.9494
R2131 X.n51 X.n48 51.9494
R2132 X.n31 X.n30 51.9494
R2133 X.n31 X.n23 51.9494
R2134 X.n40 X.n39 51.9494
R2135 X.n40 X.n32 51.9494
R2136 X.t1 X.n52 49.3036
R2137 X.n18 X.t24 16.0005
R2138 X.n18 X.t23 16.0005
R2139 X.n16 X.t15 16.0005
R2140 X.n16 X.t6 16.0005
R2141 X.n14 X.t0 16.0005
R2142 X.n14 X.t5 16.0005
R2143 X.n13 X.t7 16.0005
R2144 X.n13 X.t21 16.0005
R2145 X.n12 X.t20 16.0005
R2146 X.n12 X.t8 16.0005
R2147 X.n11 X.t13 16.0005
R2148 X.n11 X.t10 16.0005
R2149 X.n52 X.n42 15.7193
R2150 X.n9 X.t17 11.2576
R2151 X.n9 X.t12 11.2576
R2152 X.n7 X.t16 11.2576
R2153 X.n7 X.t22 11.2576
R2154 X.n5 X.t11 11.2576
R2155 X.n5 X.t2 11.2576
R2156 X.n3 X.t9 11.2576
R2157 X.n3 X.t18 11.2576
R2158 X.n1 X.t19 11.2576
R2159 X.n1 X.t3 11.2576
R2160 X.n0 X.t14 11.2576
R2161 X.n0 X.t4 11.2576
R2162 X.n42 X.n22 10.188
R2163 X.n42 X.n41 6.188
R2164 X.n10 X.n8 5.1255
R2165 X.n21 X.n20 4.5005
R2166 X.n4 X.n2 0.6255
R2167 X.n6 X.n4 0.6255
R2168 X.n8 X.n6 0.6255
R2169 X.n17 X.n15 0.563
R2170 X.n19 X.n17 0.563
R2171 X.n20 X.n19 0.563
R2172 X.n22 X.n10 0.5005
R2173 X.n22 X.n21 0.438
R2174 VOUT+.n2 VOUT+.n0 145.989
R2175 VOUT+.n8 VOUT+.n7 145.989
R2176 VOUT+.n6 VOUT+.n5 145.427
R2177 VOUT+.n4 VOUT+.n3 145.427
R2178 VOUT+.n2 VOUT+.n1 145.427
R2179 VOUT+.n10 VOUT+.n9 140.927
R2180 VOUT+.n100 VOUT+.t18 113.192
R2181 VOUT+.n97 VOUT+.n95 95.7303
R2182 VOUT+.n99 VOUT+.n98 94.6053
R2183 VOUT+.n97 VOUT+.n96 94.6053
R2184 VOUT+.n94 VOUT+.n10 20.5943
R2185 VOUT+.n94 VOUT+.n93 11.7059
R2186 VOUT+ VOUT+.n94 7.813
R2187 VOUT+.n9 VOUT+.t4 6.56717
R2188 VOUT+.n9 VOUT+.t11 6.56717
R2189 VOUT+.n7 VOUT+.t7 6.56717
R2190 VOUT+.n7 VOUT+.t13 6.56717
R2191 VOUT+.n5 VOUT+.t0 6.56717
R2192 VOUT+.n5 VOUT+.t8 6.56717
R2193 VOUT+.n3 VOUT+.t1 6.56717
R2194 VOUT+.n3 VOUT+.t17 6.56717
R2195 VOUT+.n1 VOUT+.t16 6.56717
R2196 VOUT+.n1 VOUT+.t5 6.56717
R2197 VOUT+.n0 VOUT+.t12 6.56717
R2198 VOUT+.n0 VOUT+.t9 6.56717
R2199 VOUT+.n40 VOUT+.t67 4.8295
R2200 VOUT+.n52 VOUT+.t58 4.8295
R2201 VOUT+.n49 VOUT+.t93 4.8295
R2202 VOUT+.n46 VOUT+.t131 4.8295
R2203 VOUT+.n43 VOUT+.t46 4.8295
R2204 VOUT+.n42 VOUT+.t30 4.8295
R2205 VOUT+.n66 VOUT+.t56 4.8295
R2206 VOUT+.n67 VOUT+.t119 4.8295
R2207 VOUT+.n69 VOUT+.t90 4.8295
R2208 VOUT+.n70 VOUT+.t153 4.8295
R2209 VOUT+.n72 VOUT+.t52 4.8295
R2210 VOUT+.n73 VOUT+.t109 4.8295
R2211 VOUT+.n75 VOUT+.t150 4.8295
R2212 VOUT+.n76 VOUT+.t73 4.8295
R2213 VOUT+.n78 VOUT+.t51 4.8295
R2214 VOUT+.n79 VOUT+.t105 4.8295
R2215 VOUT+.n81 VOUT+.t145 4.8295
R2216 VOUT+.n82 VOUT+.t69 4.8295
R2217 VOUT+.n84 VOUT+.t102 4.8295
R2218 VOUT+.n85 VOUT+.t34 4.8295
R2219 VOUT+.n87 VOUT+.t65 4.8295
R2220 VOUT+.n88 VOUT+.t133 4.8295
R2221 VOUT+.n11 VOUT+.t98 4.8295
R2222 VOUT+.n13 VOUT+.t146 4.8295
R2223 VOUT+.n25 VOUT+.t123 4.8295
R2224 VOUT+.n26 VOUT+.t104 4.8295
R2225 VOUT+.n28 VOUT+.t156 4.8295
R2226 VOUT+.n29 VOUT+.t79 4.8295
R2227 VOUT+.n31 VOUT+.t55 4.8295
R2228 VOUT+.n32 VOUT+.t117 4.8295
R2229 VOUT+.n34 VOUT+.t22 4.8295
R2230 VOUT+.n35 VOUT+.t84 4.8295
R2231 VOUT+.n37 VOUT+.t59 4.8295
R2232 VOUT+.n38 VOUT+.t124 4.8295
R2233 VOUT+.n90 VOUT+.t97 4.8295
R2234 VOUT+.n55 VOUT+.t130 4.806
R2235 VOUT+.n56 VOUT+.t28 4.806
R2236 VOUT+.n57 VOUT+.t62 4.806
R2237 VOUT+.n58 VOUT+.t99 4.806
R2238 VOUT+.n59 VOUT+.t81 4.806
R2239 VOUT+.n60 VOUT+.t114 4.806
R2240 VOUT+.n61 VOUT+.t155 4.806
R2241 VOUT+.n62 VOUT+.t140 4.806
R2242 VOUT+.n63 VOUT+.t39 4.806
R2243 VOUT+.n64 VOUT+.t151 4.806
R2244 VOUT+.n14 VOUT+.t138 4.806
R2245 VOUT+.n15 VOUT+.t31 4.806
R2246 VOUT+.n16 VOUT+.t61 4.806
R2247 VOUT+.n17 VOUT+.t95 4.806
R2248 VOUT+.n18 VOUT+.t148 4.806
R2249 VOUT+.n19 VOUT+.t50 4.806
R2250 VOUT+.n20 VOUT+.t80 4.806
R2251 VOUT+.n21 VOUT+.t135 4.806
R2252 VOUT+.n22 VOUT+.t27 4.806
R2253 VOUT+.n23 VOUT+.t121 4.806
R2254 VOUT+.n40 VOUT+.t33 4.5005
R2255 VOUT+.n41 VOUT+.t136 4.5005
R2256 VOUT+.n52 VOUT+.t96 4.5005
R2257 VOUT+.n53 VOUT+.t143 4.5005
R2258 VOUT+.n54 VOUT+.t100 4.5005
R2259 VOUT+.n49 VOUT+.t139 4.5005
R2260 VOUT+.n50 VOUT+.t41 4.5005
R2261 VOUT+.n51 VOUT+.t144 4.5005
R2262 VOUT+.n46 VOUT+.t32 4.5005
R2263 VOUT+.n47 VOUT+.t68 4.5005
R2264 VOUT+.n48 VOUT+.t42 4.5005
R2265 VOUT+.n43 VOUT+.t77 4.5005
R2266 VOUT+.n44 VOUT+.t116 4.5005
R2267 VOUT+.n45 VOUT+.t86 4.5005
R2268 VOUT+.n42 VOUT+.t132 4.5005
R2269 VOUT+.n65 VOUT+.t92 4.5005
R2270 VOUT+.n64 VOUT+.t108 4.5005
R2271 VOUT+.n63 VOUT+.t137 4.5005
R2272 VOUT+.n62 VOUT+.t94 4.5005
R2273 VOUT+.n61 VOUT+.t112 4.5005
R2274 VOUT+.n60 VOUT+.t76 4.5005
R2275 VOUT+.n59 VOUT+.t48 4.5005
R2276 VOUT+.n58 VOUT+.t60 4.5005
R2277 VOUT+.n57 VOUT+.t23 4.5005
R2278 VOUT+.n56 VOUT+.t129 4.5005
R2279 VOUT+.n55 VOUT+.t89 4.5005
R2280 VOUT+.n66 VOUT+.t21 4.5005
R2281 VOUT+.n68 VOUT+.t127 4.5005
R2282 VOUT+.n67 VOUT+.t74 4.5005
R2283 VOUT+.n69 VOUT+.t54 4.5005
R2284 VOUT+.n71 VOUT+.t20 4.5005
R2285 VOUT+.n70 VOUT+.t106 4.5005
R2286 VOUT+.n72 VOUT+.t154 4.5005
R2287 VOUT+.n74 VOUT+.t122 4.5005
R2288 VOUT+.n73 VOUT+.t70 4.5005
R2289 VOUT+.n75 VOUT+.t111 4.5005
R2290 VOUT+.n77 VOUT+.t82 4.5005
R2291 VOUT+.n76 VOUT+.t35 4.5005
R2292 VOUT+.n78 VOUT+.t149 4.5005
R2293 VOUT+.n80 VOUT+.t110 4.5005
R2294 VOUT+.n79 VOUT+.t63 4.5005
R2295 VOUT+.n81 VOUT+.t107 4.5005
R2296 VOUT+.n83 VOUT+.t75 4.5005
R2297 VOUT+.n82 VOUT+.t25 4.5005
R2298 VOUT+.n84 VOUT+.t71 4.5005
R2299 VOUT+.n86 VOUT+.t44 4.5005
R2300 VOUT+.n85 VOUT+.t125 4.5005
R2301 VOUT+.n87 VOUT+.t37 4.5005
R2302 VOUT+.n89 VOUT+.t141 4.5005
R2303 VOUT+.n88 VOUT+.t85 4.5005
R2304 VOUT+.n11 VOUT+.t66 4.5005
R2305 VOUT+.n12 VOUT+.t38 4.5005
R2306 VOUT+.n13 VOUT+.t53 4.5005
R2307 VOUT+.n24 VOUT+.t101 4.5005
R2308 VOUT+.n23 VOUT+.t113 4.5005
R2309 VOUT+.n22 VOUT+.t115 4.5005
R2310 VOUT+.n21 VOUT+.t29 4.5005
R2311 VOUT+.n20 VOUT+.t45 4.5005
R2312 VOUT+.n19 VOUT+.t88 4.5005
R2313 VOUT+.n18 VOUT+.t142 4.5005
R2314 VOUT+.n17 VOUT+.t147 4.5005
R2315 VOUT+.n16 VOUT+.t57 4.5005
R2316 VOUT+.n15 VOUT+.t103 4.5005
R2317 VOUT+.n14 VOUT+.t152 4.5005
R2318 VOUT+.n25 VOUT+.t40 4.5005
R2319 VOUT+.n27 VOUT+.t83 4.5005
R2320 VOUT+.n26 VOUT+.t49 4.5005
R2321 VOUT+.n28 VOUT+.t120 4.5005
R2322 VOUT+.n30 VOUT+.t87 4.5005
R2323 VOUT+.n29 VOUT+.t43 4.5005
R2324 VOUT+.n31 VOUT+.t19 4.5005
R2325 VOUT+.n33 VOUT+.t126 4.5005
R2326 VOUT+.n32 VOUT+.t72 4.5005
R2327 VOUT+.n34 VOUT+.t128 4.5005
R2328 VOUT+.n36 VOUT+.t91 4.5005
R2329 VOUT+.n35 VOUT+.t47 4.5005
R2330 VOUT+.n37 VOUT+.t26 4.5005
R2331 VOUT+.n39 VOUT+.t134 4.5005
R2332 VOUT+.n38 VOUT+.t78 4.5005
R2333 VOUT+.n90 VOUT+.t64 4.5005
R2334 VOUT+.n91 VOUT+.t36 4.5005
R2335 VOUT+.n92 VOUT+.t118 4.5005
R2336 VOUT+.n93 VOUT+.t24 4.5005
R2337 VOUT+.n10 VOUT+.n8 4.5005
R2338 VOUT+.n98 VOUT+.t15 3.42907
R2339 VOUT+.n98 VOUT+.t10 3.42907
R2340 VOUT+.n96 VOUT+.t6 3.42907
R2341 VOUT+.n96 VOUT+.t2 3.42907
R2342 VOUT+.n95 VOUT+.t3 3.42907
R2343 VOUT+.n95 VOUT+.t14 3.42907
R2344 VOUT+ VOUT+.n100 2.84425
R2345 VOUT+.n100 VOUT+.n99 2.03175
R2346 VOUT+.n99 VOUT+.n97 1.1255
R2347 VOUT+.n4 VOUT+.n2 0.563
R2348 VOUT+.n6 VOUT+.n4 0.563
R2349 VOUT+.n8 VOUT+.n6 0.563
R2350 VOUT+.n41 VOUT+.n40 0.3295
R2351 VOUT+.n54 VOUT+.n53 0.3295
R2352 VOUT+.n53 VOUT+.n52 0.3295
R2353 VOUT+.n51 VOUT+.n50 0.3295
R2354 VOUT+.n50 VOUT+.n49 0.3295
R2355 VOUT+.n48 VOUT+.n47 0.3295
R2356 VOUT+.n47 VOUT+.n46 0.3295
R2357 VOUT+.n45 VOUT+.n44 0.3295
R2358 VOUT+.n44 VOUT+.n43 0.3295
R2359 VOUT+.n65 VOUT+.n42 0.3295
R2360 VOUT+.n65 VOUT+.n64 0.3295
R2361 VOUT+.n64 VOUT+.n63 0.3295
R2362 VOUT+.n63 VOUT+.n62 0.3295
R2363 VOUT+.n62 VOUT+.n61 0.3295
R2364 VOUT+.n61 VOUT+.n60 0.3295
R2365 VOUT+.n60 VOUT+.n59 0.3295
R2366 VOUT+.n59 VOUT+.n58 0.3295
R2367 VOUT+.n58 VOUT+.n57 0.3295
R2368 VOUT+.n57 VOUT+.n56 0.3295
R2369 VOUT+.n56 VOUT+.n55 0.3295
R2370 VOUT+.n68 VOUT+.n66 0.3295
R2371 VOUT+.n68 VOUT+.n67 0.3295
R2372 VOUT+.n71 VOUT+.n69 0.3295
R2373 VOUT+.n71 VOUT+.n70 0.3295
R2374 VOUT+.n74 VOUT+.n72 0.3295
R2375 VOUT+.n74 VOUT+.n73 0.3295
R2376 VOUT+.n77 VOUT+.n75 0.3295
R2377 VOUT+.n77 VOUT+.n76 0.3295
R2378 VOUT+.n80 VOUT+.n78 0.3295
R2379 VOUT+.n80 VOUT+.n79 0.3295
R2380 VOUT+.n83 VOUT+.n81 0.3295
R2381 VOUT+.n83 VOUT+.n82 0.3295
R2382 VOUT+.n86 VOUT+.n84 0.3295
R2383 VOUT+.n86 VOUT+.n85 0.3295
R2384 VOUT+.n89 VOUT+.n87 0.3295
R2385 VOUT+.n89 VOUT+.n88 0.3295
R2386 VOUT+.n12 VOUT+.n11 0.3295
R2387 VOUT+.n24 VOUT+.n13 0.3295
R2388 VOUT+.n24 VOUT+.n23 0.3295
R2389 VOUT+.n23 VOUT+.n22 0.3295
R2390 VOUT+.n22 VOUT+.n21 0.3295
R2391 VOUT+.n21 VOUT+.n20 0.3295
R2392 VOUT+.n20 VOUT+.n19 0.3295
R2393 VOUT+.n19 VOUT+.n18 0.3295
R2394 VOUT+.n18 VOUT+.n17 0.3295
R2395 VOUT+.n17 VOUT+.n16 0.3295
R2396 VOUT+.n16 VOUT+.n15 0.3295
R2397 VOUT+.n15 VOUT+.n14 0.3295
R2398 VOUT+.n27 VOUT+.n25 0.3295
R2399 VOUT+.n27 VOUT+.n26 0.3295
R2400 VOUT+.n30 VOUT+.n28 0.3295
R2401 VOUT+.n30 VOUT+.n29 0.3295
R2402 VOUT+.n33 VOUT+.n31 0.3295
R2403 VOUT+.n33 VOUT+.n32 0.3295
R2404 VOUT+.n36 VOUT+.n34 0.3295
R2405 VOUT+.n36 VOUT+.n35 0.3295
R2406 VOUT+.n39 VOUT+.n37 0.3295
R2407 VOUT+.n39 VOUT+.n38 0.3295
R2408 VOUT+.n91 VOUT+.n90 0.3295
R2409 VOUT+.n92 VOUT+.n91 0.3295
R2410 VOUT+.n93 VOUT+.n92 0.3295
R2411 VOUT+.n59 VOUT+.n54 0.306
R2412 VOUT+.n60 VOUT+.n51 0.306
R2413 VOUT+.n61 VOUT+.n48 0.306
R2414 VOUT+.n62 VOUT+.n45 0.306
R2415 VOUT+.n65 VOUT+.n41 0.2825
R2416 VOUT+.n68 VOUT+.n65 0.2825
R2417 VOUT+.n71 VOUT+.n68 0.2825
R2418 VOUT+.n74 VOUT+.n71 0.2825
R2419 VOUT+.n77 VOUT+.n74 0.2825
R2420 VOUT+.n80 VOUT+.n77 0.2825
R2421 VOUT+.n83 VOUT+.n80 0.2825
R2422 VOUT+.n86 VOUT+.n83 0.2825
R2423 VOUT+.n89 VOUT+.n86 0.2825
R2424 VOUT+.n24 VOUT+.n12 0.2825
R2425 VOUT+.n27 VOUT+.n24 0.2825
R2426 VOUT+.n30 VOUT+.n27 0.2825
R2427 VOUT+.n33 VOUT+.n30 0.2825
R2428 VOUT+.n36 VOUT+.n33 0.2825
R2429 VOUT+.n39 VOUT+.n36 0.2825
R2430 VOUT+.n91 VOUT+.n39 0.2825
R2431 VOUT+.n91 VOUT+.n89 0.2825
R2432 cap_res_Y.t0 cap_res_Y.t26 49.2006
R2433 cap_res_Y.t61 cap_res_Y.t99 0.1603
R2434 cap_res_Y.t14 cap_res_Y.t61 0.1603
R2435 cap_res_Y.t57 cap_res_Y.t14 0.1603
R2436 cap_res_Y.t109 cap_res_Y.t57 0.1603
R2437 cap_res_Y.t18 cap_res_Y.t64 0.1603
R2438 cap_res_Y.t116 cap_res_Y.t18 0.1603
R2439 cap_res_Y.t13 cap_res_Y.t116 0.1603
R2440 cap_res_Y.t81 cap_res_Y.t13 0.1603
R2441 cap_res_Y.t25 cap_res_Y.t127 0.1603
R2442 cap_res_Y.t124 cap_res_Y.t90 0.1603
R2443 cap_res_Y.t83 cap_res_Y.t38 0.1603
R2444 cap_res_Y.t136 cap_res_Y.t101 0.1603
R2445 cap_res_Y.t51 cap_res_Y.t4 0.1603
R2446 cap_res_Y.t103 cap_res_Y.t67 0.1603
R2447 cap_res_Y.t87 cap_res_Y.t48 0.1603
R2448 cap_res_Y.t3 cap_res_Y.t105 0.1603
R2449 cap_res_Y.t122 cap_res_Y.t84 0.1603
R2450 cap_res_Y.t46 cap_res_Y.t7 0.1603
R2451 cap_res_Y.t94 cap_res_Y.t52 0.1603
R2452 cap_res_Y.t8 cap_res_Y.t106 0.1603
R2453 cap_res_Y.t132 cap_res_Y.t88 0.1603
R2454 cap_res_Y.t50 cap_res_Y.t12 0.1603
R2455 cap_res_Y.t32 cap_res_Y.t123 0.1603
R2456 cap_res_Y.t86 cap_res_Y.t55 0.1603
R2457 cap_res_Y.t72 cap_res_Y.t24 0.1603
R2458 cap_res_Y.t120 cap_res_Y.t92 0.1603
R2459 cap_res_Y.t39 cap_res_Y.t133 0.1603
R2460 cap_res_Y.t93 cap_res_Y.t60 0.1603
R2461 cap_res_Y.t79 cap_res_Y.t33 0.1603
R2462 cap_res_Y.t131 cap_res_Y.t98 0.1603
R2463 cap_res_Y.t110 cap_res_Y.t73 0.1603
R2464 cap_res_Y.t29 cap_res_Y.t135 0.1603
R2465 cap_res_Y.t85 cap_res_Y.t40 0.1603
R2466 cap_res_Y.t138 cap_res_Y.t102 0.1603
R2467 cap_res_Y.t114 cap_res_Y.t78 0.1603
R2468 cap_res_Y.t37 cap_res_Y.t1 0.1603
R2469 cap_res_Y.t108 cap_res_Y.t53 0.1603
R2470 cap_res_Y.t117 cap_res_Y.t34 0.1603
R2471 cap_res_Y.t5 cap_res_Y.t19 0.1603
R2472 cap_res_Y.t54 cap_res_Y.t126 0.1603
R2473 cap_res_Y.t100 cap_res_Y.t96 0.1603
R2474 cap_res_Y.t10 cap_res_Y.t62 0.1603
R2475 cap_res_Y.t15 cap_res_Y.t9 0.1603
R2476 cap_res_Y.t69 cap_res_Y.t107 0.1603
R2477 cap_res_Y.t112 cap_res_Y.t77 0.1603
R2478 cap_res_Y.t128 cap_res_Y.t22 0.1603
R2479 cap_res_Y.t42 cap_res_Y.t130 0.1603
R2480 cap_res_Y.t44 cap_res_Y.t36 0.1603
R2481 cap_res_Y.t104 cap_res_Y.t11 0.1603
R2482 cap_res_Y.t91 cap_res_Y.t59 0.1603
R2483 cap_res_Y.t80 cap_res_Y.t111 0.1603
R2484 cap_res_Y.t41 cap_res_Y.t80 0.1603
R2485 cap_res_Y.t71 cap_res_Y.t41 0.1603
R2486 cap_res_Y.t63 cap_res_Y.t71 0.1603
R2487 cap_res_Y.t115 cap_res_Y.t45 0.1603
R2488 cap_res_Y.t89 cap_res_Y.t115 0.1603
R2489 cap_res_Y.t125 cap_res_Y.t89 0.1603
R2490 cap_res_Y.t26 cap_res_Y.t125 0.1603
R2491 cap_res_Y.n29 cap_res_Y.t27 0.159278
R2492 cap_res_Y.n30 cap_res_Y.t129 0.159278
R2493 cap_res_Y.n31 cap_res_Y.t95 0.159278
R2494 cap_res_Y.n32 cap_res_Y.t58 0.159278
R2495 cap_res_Y.n33 cap_res_Y.t76 0.159278
R2496 cap_res_Y.n34 cap_res_Y.t43 0.159278
R2497 cap_res_Y.n25 cap_res_Y.t21 0.159278
R2498 cap_res_Y.t56 cap_res_Y.n9 0.159278
R2499 cap_res_Y.t74 cap_res_Y.n10 0.159278
R2500 cap_res_Y.t70 cap_res_Y.n11 0.159278
R2501 cap_res_Y.t31 cap_res_Y.n12 0.159278
R2502 cap_res_Y.t66 cap_res_Y.n13 0.159278
R2503 cap_res_Y.t23 cap_res_Y.n14 0.159278
R2504 cap_res_Y.t121 cap_res_Y.n15 0.159278
R2505 cap_res_Y.t16 cap_res_Y.n16 0.159278
R2506 cap_res_Y.t113 cap_res_Y.n17 0.159278
R2507 cap_res_Y.t82 cap_res_Y.n18 0.159278
R2508 cap_res_Y.t47 cap_res_Y.n19 0.159278
R2509 cap_res_Y.t75 cap_res_Y.n20 0.159278
R2510 cap_res_Y.t35 cap_res_Y.n21 0.159278
R2511 cap_res_Y.t137 cap_res_Y.n22 0.159278
R2512 cap_res_Y.t30 cap_res_Y.n23 0.159278
R2513 cap_res_Y.t65 cap_res_Y.n24 0.159278
R2514 cap_res_Y.n26 cap_res_Y.t6 0.159278
R2515 cap_res_Y.n27 cap_res_Y.t118 0.159278
R2516 cap_res_Y.n28 cap_res_Y.t17 0.159278
R2517 cap_res_Y.n35 cap_res_Y.t2 0.159278
R2518 cap_res_Y.t21 cap_res_Y.t124 0.137822
R2519 cap_res_Y.n25 cap_res_Y.t25 0.1368
R2520 cap_res_Y.n24 cap_res_Y.t83 0.1368
R2521 cap_res_Y.n24 cap_res_Y.t136 0.1368
R2522 cap_res_Y.n23 cap_res_Y.t51 0.1368
R2523 cap_res_Y.n23 cap_res_Y.t103 0.1368
R2524 cap_res_Y.n22 cap_res_Y.t87 0.1368
R2525 cap_res_Y.n22 cap_res_Y.t3 0.1368
R2526 cap_res_Y.n21 cap_res_Y.t122 0.1368
R2527 cap_res_Y.n21 cap_res_Y.t46 0.1368
R2528 cap_res_Y.n20 cap_res_Y.t94 0.1368
R2529 cap_res_Y.n20 cap_res_Y.t8 0.1368
R2530 cap_res_Y.n19 cap_res_Y.t132 0.1368
R2531 cap_res_Y.n19 cap_res_Y.t50 0.1368
R2532 cap_res_Y.n18 cap_res_Y.t32 0.1368
R2533 cap_res_Y.n18 cap_res_Y.t86 0.1368
R2534 cap_res_Y.n17 cap_res_Y.t72 0.1368
R2535 cap_res_Y.n17 cap_res_Y.t120 0.1368
R2536 cap_res_Y.n16 cap_res_Y.t39 0.1368
R2537 cap_res_Y.n16 cap_res_Y.t93 0.1368
R2538 cap_res_Y.n15 cap_res_Y.t79 0.1368
R2539 cap_res_Y.n15 cap_res_Y.t131 0.1368
R2540 cap_res_Y.n14 cap_res_Y.t110 0.1368
R2541 cap_res_Y.n14 cap_res_Y.t29 0.1368
R2542 cap_res_Y.n13 cap_res_Y.t85 0.1368
R2543 cap_res_Y.n13 cap_res_Y.t138 0.1368
R2544 cap_res_Y.n12 cap_res_Y.t114 0.1368
R2545 cap_res_Y.n12 cap_res_Y.t37 0.1368
R2546 cap_res_Y.n11 cap_res_Y.t108 0.1368
R2547 cap_res_Y.n11 cap_res_Y.t117 0.1368
R2548 cap_res_Y.n10 cap_res_Y.t104 0.1368
R2549 cap_res_Y.n9 cap_res_Y.t91 0.1368
R2550 cap_res_Y.n0 cap_res_Y.t5 0.114322
R2551 cap_res_Y.n30 cap_res_Y.n29 0.1133
R2552 cap_res_Y.n31 cap_res_Y.n30 0.1133
R2553 cap_res_Y.n32 cap_res_Y.n31 0.1133
R2554 cap_res_Y.n33 cap_res_Y.n32 0.1133
R2555 cap_res_Y.n34 cap_res_Y.n33 0.1133
R2556 cap_res_Y.n1 cap_res_Y.n0 0.1133
R2557 cap_res_Y.n2 cap_res_Y.n1 0.1133
R2558 cap_res_Y.n3 cap_res_Y.n2 0.1133
R2559 cap_res_Y.n4 cap_res_Y.n3 0.1133
R2560 cap_res_Y.n5 cap_res_Y.n4 0.1133
R2561 cap_res_Y.n6 cap_res_Y.n5 0.1133
R2562 cap_res_Y.n7 cap_res_Y.n6 0.1133
R2563 cap_res_Y.n8 cap_res_Y.n7 0.1133
R2564 cap_res_Y.n10 cap_res_Y.n8 0.1133
R2565 cap_res_Y.n26 cap_res_Y.n25 0.1133
R2566 cap_res_Y.n27 cap_res_Y.n26 0.1133
R2567 cap_res_Y.n28 cap_res_Y.n27 0.1133
R2568 cap_res_Y.n35 cap_res_Y.n28 0.1133
R2569 cap_res_Y.n35 cap_res_Y.n34 0.1133
R2570 cap_res_Y.n29 cap_res_Y.t68 0.00152174
R2571 cap_res_Y.n30 cap_res_Y.t28 0.00152174
R2572 cap_res_Y.n31 cap_res_Y.t134 0.00152174
R2573 cap_res_Y.n32 cap_res_Y.t97 0.00152174
R2574 cap_res_Y.n33 cap_res_Y.t109 0.00152174
R2575 cap_res_Y.n34 cap_res_Y.t81 0.00152174
R2576 cap_res_Y.n0 cap_res_Y.t54 0.00152174
R2577 cap_res_Y.n1 cap_res_Y.t100 0.00152174
R2578 cap_res_Y.n2 cap_res_Y.t10 0.00152174
R2579 cap_res_Y.n3 cap_res_Y.t15 0.00152174
R2580 cap_res_Y.n4 cap_res_Y.t69 0.00152174
R2581 cap_res_Y.n5 cap_res_Y.t112 0.00152174
R2582 cap_res_Y.n6 cap_res_Y.t128 0.00152174
R2583 cap_res_Y.n7 cap_res_Y.t42 0.00152174
R2584 cap_res_Y.n8 cap_res_Y.t44 0.00152174
R2585 cap_res_Y.n9 cap_res_Y.t119 0.00152174
R2586 cap_res_Y.n10 cap_res_Y.t56 0.00152174
R2587 cap_res_Y.n11 cap_res_Y.t74 0.00152174
R2588 cap_res_Y.n12 cap_res_Y.t70 0.00152174
R2589 cap_res_Y.n13 cap_res_Y.t31 0.00152174
R2590 cap_res_Y.n14 cap_res_Y.t66 0.00152174
R2591 cap_res_Y.n15 cap_res_Y.t23 0.00152174
R2592 cap_res_Y.n16 cap_res_Y.t121 0.00152174
R2593 cap_res_Y.n17 cap_res_Y.t16 0.00152174
R2594 cap_res_Y.n18 cap_res_Y.t113 0.00152174
R2595 cap_res_Y.n19 cap_res_Y.t82 0.00152174
R2596 cap_res_Y.n20 cap_res_Y.t47 0.00152174
R2597 cap_res_Y.n21 cap_res_Y.t75 0.00152174
R2598 cap_res_Y.n22 cap_res_Y.t35 0.00152174
R2599 cap_res_Y.n23 cap_res_Y.t137 0.00152174
R2600 cap_res_Y.n24 cap_res_Y.t30 0.00152174
R2601 cap_res_Y.n25 cap_res_Y.t65 0.00152174
R2602 cap_res_Y.n26 cap_res_Y.t49 0.00152174
R2603 cap_res_Y.n27 cap_res_Y.t20 0.00152174
R2604 cap_res_Y.n28 cap_res_Y.t63 0.00152174
R2605 cap_res_Y.t45 cap_res_Y.n35 0.00152174
R2606 err_amp_mir.n2 err_amp_mir.n0 628.034
R2607 err_amp_mir.n4 err_amp_mir.n3 626.784
R2608 err_amp_mir.n2 err_amp_mir.n1 626.784
R2609 err_amp_mir.n7 err_amp_mir.t11 289.2
R2610 err_amp_mir.n6 err_amp_mir.t19 289.2
R2611 err_amp_mir.n12 err_amp_mir.n11 228.252
R2612 err_amp_mir.n13 err_amp_mir.n10 212.733
R2613 err_amp_mir.n21 err_amp_mir.n20 212.733
R2614 err_amp_mir.n9 err_amp_mir.n8 176.733
R2615 err_amp_mir.n8 err_amp_mir.n7 176.733
R2616 err_amp_mir.n18 err_amp_mir.n17 176.733
R2617 err_amp_mir.n17 err_amp_mir.n16 176.733
R2618 err_amp_mir.n16 err_amp_mir.n15 176.733
R2619 err_amp_mir.n14 err_amp_mir.n13 152
R2620 err_amp_mir.n20 err_amp_mir.n19 152
R2621 err_amp_mir.n7 err_amp_mir.t17 112.468
R2622 err_amp_mir.n8 err_amp_mir.t20 112.468
R2623 err_amp_mir.n9 err_amp_mir.t15 112.468
R2624 err_amp_mir.n6 err_amp_mir.t13 112.468
R2625 err_amp_mir.n15 err_amp_mir.t9 112.468
R2626 err_amp_mir.n16 err_amp_mir.t21 112.468
R2627 err_amp_mir.n17 err_amp_mir.t18 112.468
R2628 err_amp_mir.n18 err_amp_mir.t7 112.468
R2629 err_amp_mir.n3 err_amp_mir.t3 78.8005
R2630 err_amp_mir.n3 err_amp_mir.t2 78.8005
R2631 err_amp_mir.n1 err_amp_mir.t0 78.8005
R2632 err_amp_mir.n1 err_amp_mir.t4 78.8005
R2633 err_amp_mir.n0 err_amp_mir.t1 78.8005
R2634 err_amp_mir.n0 err_amp_mir.t5 78.8005
R2635 err_amp_mir.n10 err_amp_mir.t10 48.0005
R2636 err_amp_mir.n10 err_amp_mir.t16 48.0005
R2637 err_amp_mir.n11 err_amp_mir.t12 48.0005
R2638 err_amp_mir.n11 err_amp_mir.t6 48.0005
R2639 err_amp_mir.t14 err_amp_mir.n21 48.0005
R2640 err_amp_mir.n21 err_amp_mir.t8 48.0005
R2641 err_amp_mir.n14 err_amp_mir.n9 45.5227
R2642 err_amp_mir.n19 err_amp_mir.n6 45.5227
R2643 err_amp_mir.n19 err_amp_mir.n18 45.5227
R2644 err_amp_mir.n15 err_amp_mir.n14 45.5227
R2645 err_amp_mir.n5 err_amp_mir.n4 33.8443
R2646 err_amp_mir.n13 err_amp_mir.n12 14.2693
R2647 err_amp_mir.n20 err_amp_mir.n5 14.2693
R2648 err_amp_mir.n12 err_amp_mir.n5 1.2505
R2649 err_amp_mir.n4 err_amp_mir.n2 1.2505
R2650 Y.n43 Y.t40 1172.87
R2651 Y.n41 Y.t46 1172.87
R2652 Y.n48 Y.t36 996.134
R2653 Y.n47 Y.t51 996.134
R2654 Y.n46 Y.t27 996.134
R2655 Y.n45 Y.t43 996.134
R2656 Y.n44 Y.t30 996.134
R2657 Y.n43 Y.t54 996.134
R2658 Y.n41 Y.t33 996.134
R2659 Y.n42 Y.t48 996.134
R2660 Y.n38 Y.t49 690.867
R2661 Y.n31 Y.t25 690.867
R2662 Y.n29 Y.t38 530.201
R2663 Y.n22 Y.t45 530.201
R2664 Y.n38 Y.t34 514.134
R2665 Y.n37 Y.t39 514.134
R2666 Y.n36 Y.t53 514.134
R2667 Y.n35 Y.t37 514.134
R2668 Y.n34 Y.t31 514.134
R2669 Y.n33 Y.t44 514.134
R2670 Y.n32 Y.t28 514.134
R2671 Y.n31 Y.t41 514.134
R2672 Y.n29 Y.t52 353.467
R2673 Y.n22 Y.t32 353.467
R2674 Y.n23 Y.t47 353.467
R2675 Y.n24 Y.t35 353.467
R2676 Y.n25 Y.t50 353.467
R2677 Y.n26 Y.t26 353.467
R2678 Y.n27 Y.t42 353.467
R2679 Y.n28 Y.t29 353.467
R2680 Y.n48 Y.n47 176.733
R2681 Y.n47 Y.n46 176.733
R2682 Y.n46 Y.n45 176.733
R2683 Y.n45 Y.n44 176.733
R2684 Y.n44 Y.n43 176.733
R2685 Y.n42 Y.n41 176.733
R2686 Y.n23 Y.n22 176.733
R2687 Y.n24 Y.n23 176.733
R2688 Y.n25 Y.n24 176.733
R2689 Y.n26 Y.n25 176.733
R2690 Y.n27 Y.n26 176.733
R2691 Y.n28 Y.n27 176.733
R2692 Y.n32 Y.n31 176.733
R2693 Y.n33 Y.n32 176.733
R2694 Y.n34 Y.n33 176.733
R2695 Y.n35 Y.n34 176.733
R2696 Y.n36 Y.n35 176.733
R2697 Y.n37 Y.n36 176.733
R2698 Y.n50 Y.n49 166.375
R2699 Y.n40 Y.n30 161.875
R2700 Y.n40 Y.n39 161.686
R2701 Y.n2 Y.n0 160.427
R2702 Y.n8 Y.n7 159.802
R2703 Y.n6 Y.n5 159.802
R2704 Y.n4 Y.n3 159.802
R2705 Y.n2 Y.n1 159.802
R2706 Y.n10 Y.n9 155.302
R2707 Y.n20 Y.n19 114.689
R2708 Y.n14 Y.n12 114.689
R2709 Y.n18 Y.n17 114.126
R2710 Y.n16 Y.n15 114.126
R2711 Y.n14 Y.n13 114.126
R2712 Y.n21 Y.n11 109.626
R2713 Y.n49 Y.n48 51.9494
R2714 Y.n49 Y.n42 51.9494
R2715 Y.n30 Y.n29 51.9494
R2716 Y.n30 Y.n28 51.9494
R2717 Y.n39 Y.n38 51.9494
R2718 Y.n39 Y.n37 51.9494
R2719 Y.n50 Y.t2 49.2412
R2720 Y.n19 Y.t17 16.0005
R2721 Y.n19 Y.t20 16.0005
R2722 Y.n17 Y.t4 16.0005
R2723 Y.n17 Y.t8 16.0005
R2724 Y.n15 Y.t1 16.0005
R2725 Y.n15 Y.t10 16.0005
R2726 Y.n13 Y.t9 16.0005
R2727 Y.n13 Y.t12 16.0005
R2728 Y.n12 Y.t19 16.0005
R2729 Y.n12 Y.t13 16.0005
R2730 Y.n11 Y.t22 16.0005
R2731 Y.n11 Y.t3 16.0005
R2732 Y.n51 Y.n50 15.6567
R2733 Y.n9 Y.t15 11.2576
R2734 Y.n9 Y.t24 11.2576
R2735 Y.n7 Y.t18 11.2576
R2736 Y.n7 Y.t16 11.2576
R2737 Y.n5 Y.t11 11.2576
R2738 Y.n5 Y.t14 11.2576
R2739 Y.n3 Y.t6 11.2576
R2740 Y.n3 Y.t21 11.2576
R2741 Y.n1 Y.t7 11.2576
R2742 Y.n1 Y.t5 11.2576
R2743 Y.n0 Y.t23 11.2576
R2744 Y.n0 Y.t0 11.2576
R2745 Y Y.n51 10.313
R2746 Y.n51 Y.n40 6.063
R2747 Y.n10 Y.n8 5.1255
R2748 Y.n21 Y.n20 4.5005
R2749 Y.n4 Y.n2 0.6255
R2750 Y.n6 Y.n4 0.6255
R2751 Y.n8 Y.n6 0.6255
R2752 Y.n16 Y.n14 0.563
R2753 Y.n18 Y.n16 0.563
R2754 Y.n20 Y.n18 0.563
R2755 Y Y.n10 0.5005
R2756 Y Y.n21 0.438
R2757 V_CMFB_S4 V_CMFB_S4.t10 125.129
R2758 V_CMFB_S4.n2 V_CMFB_S4.n1 96.9009
R2759 V_CMFB_S4.n4 V_CMFB_S4.n3 96.8384
R2760 V_CMFB_S4.n6 V_CMFB_S4.n5 96.8384
R2761 V_CMFB_S4.n8 V_CMFB_S4.n7 96.8384
R2762 V_CMFB_S4.n10 V_CMFB_S4.n9 96.8384
R2763 V_CMFB_S4.n1 V_CMFB_S4.t6 8.0005
R2764 V_CMFB_S4.n1 V_CMFB_S4.t1 8.0005
R2765 V_CMFB_S4.n3 V_CMFB_S4.t0 8.0005
R2766 V_CMFB_S4.n3 V_CMFB_S4.t4 8.0005
R2767 V_CMFB_S4.n5 V_CMFB_S4.t7 8.0005
R2768 V_CMFB_S4.n5 V_CMFB_S4.t5 8.0005
R2769 V_CMFB_S4.n7 V_CMFB_S4.t8 8.0005
R2770 V_CMFB_S4.n7 V_CMFB_S4.t2 8.0005
R2771 V_CMFB_S4.n9 V_CMFB_S4.t9 8.0005
R2772 V_CMFB_S4.n9 V_CMFB_S4.t3 8.0005
R2773 V_CMFB_S4.n2 V_CMFB_S4.n0 2.04738
R2774 V_CMFB_S4 V_CMFB_S4.n10 1.34425
R2775 V_CMFB_S4.n10 V_CMFB_S4.n8 0.563
R2776 V_CMFB_S4.n8 V_CMFB_S4.n6 0.563
R2777 V_CMFB_S4.n6 V_CMFB_S4.n4 0.563
R2778 V_CMFB_S4.n4 V_CMFB_S4.n2 0.5005
R2779 a_58940_5092.t0 a_58940_5092.t1 291.822
R2780 V_CMFB_S2 V_CMFB_S2.t0 125.16
R2781 V_CMFB_S2.n2 V_CMFB_S2.n0 97.4009
R2782 V_CMFB_S2.n8 V_CMFB_S2.n7 96.8384
R2783 V_CMFB_S2.n6 V_CMFB_S2.n5 96.8384
R2784 V_CMFB_S2.n4 V_CMFB_S2.n3 96.8384
R2785 V_CMFB_S2.n2 V_CMFB_S2.n1 96.8384
R2786 V_CMFB_S2.n7 V_CMFB_S2.t2 8.0005
R2787 V_CMFB_S2.n7 V_CMFB_S2.t6 8.0005
R2788 V_CMFB_S2.n5 V_CMFB_S2.t3 8.0005
R2789 V_CMFB_S2.n5 V_CMFB_S2.t7 8.0005
R2790 V_CMFB_S2.n3 V_CMFB_S2.t4 8.0005
R2791 V_CMFB_S2.n3 V_CMFB_S2.t8 8.0005
R2792 V_CMFB_S2.n1 V_CMFB_S2.t5 8.0005
R2793 V_CMFB_S2.n1 V_CMFB_S2.t9 8.0005
R2794 V_CMFB_S2.n0 V_CMFB_S2.t1 8.0005
R2795 V_CMFB_S2.n0 V_CMFB_S2.t10 8.0005
R2796 V_CMFB_S2 V_CMFB_S2.n8 1.313
R2797 V_CMFB_S2.n4 V_CMFB_S2.n2 0.563
R2798 V_CMFB_S2.n6 V_CMFB_S2.n4 0.563
R2799 V_CMFB_S2.n8 V_CMFB_S2.n6 0.563
R2800 Vb1.n14 Vb1.t20 449.868
R2801 Vb1.n10 Vb1.t3 449.868
R2802 Vb1.n5 Vb1.t4 449.868
R2803 Vb1.n1 Vb1.t9 449.868
R2804 Vb1.n14 Vb1.t10 273.134
R2805 Vb1.n15 Vb1.t17 273.134
R2806 Vb1.n16 Vb1.t6 273.134
R2807 Vb1.n17 Vb1.t18 273.134
R2808 Vb1.n13 Vb1.t7 273.134
R2809 Vb1.n12 Vb1.t16 273.134
R2810 Vb1.n11 Vb1.t5 273.134
R2811 Vb1.n10 Vb1.t15 273.134
R2812 Vb1.n5 Vb1.t14 273.134
R2813 Vb1.n6 Vb1.t2 273.134
R2814 Vb1.n7 Vb1.t12 273.134
R2815 Vb1.n8 Vb1.t21 273.134
R2816 Vb1.n4 Vb1.t11 273.134
R2817 Vb1.n3 Vb1.t19 273.134
R2818 Vb1.n2 Vb1.t8 273.134
R2819 Vb1.n1 Vb1.t13 273.134
R2820 Vb1.n0 Vb1.t1 184.498
R2821 Vb1.n17 Vb1.n16 176.733
R2822 Vb1.n16 Vb1.n15 176.733
R2823 Vb1.n15 Vb1.n14 176.733
R2824 Vb1.n11 Vb1.n10 176.733
R2825 Vb1.n12 Vb1.n11 176.733
R2826 Vb1.n13 Vb1.n12 176.733
R2827 Vb1.n8 Vb1.n7 176.733
R2828 Vb1.n7 Vb1.n6 176.733
R2829 Vb1.n6 Vb1.n5 176.733
R2830 Vb1.n2 Vb1.n1 176.733
R2831 Vb1.n3 Vb1.n2 176.733
R2832 Vb1.n4 Vb1.n3 176.733
R2833 Vb1.n19 Vb1.n9 170.269
R2834 Vb1.n19 Vb1.n18 165.8
R2835 Vb1.n0 Vb1.t0 58.5723
R2836 Vb1.n18 Vb1.n17 56.2338
R2837 Vb1.n18 Vb1.n13 56.2338
R2838 Vb1.n9 Vb1.n8 56.2338
R2839 Vb1.n9 Vb1.n4 56.2338
R2840 Vb1.n20 Vb1.n0 20.7804
R2841 Vb1.n20 Vb1.n19 8.67238
R2842 Vb1 Vb1.n20 0.063
R2843 VD1.n9 VD1.n7 114.719
R2844 VD1.n6 VD1.n4 114.719
R2845 VD1.n6 VD1.n5 114.156
R2846 VD1.n9 VD1.n8 114.156
R2847 VD1.n2 VD1.n0 113.081
R2848 VD1.n16 VD1.n15 111.769
R2849 VD1.n18 VD1.n17 111.769
R2850 VD1 VD1.n19 111.769
R2851 VD1.n2 VD1.n1 111.769
R2852 VD1.n11 VD1.n3 109.656
R2853 VD1.n13 VD1.n12 107.269
R2854 VD1.n7 VD1.t13 16.0005
R2855 VD1.n7 VD1.t19 16.0005
R2856 VD1.n3 VD1.t16 16.0005
R2857 VD1.n3 VD1.t11 16.0005
R2858 VD1.n15 VD1.t10 16.0005
R2859 VD1.n15 VD1.t8 16.0005
R2860 VD1.n17 VD1.t4 16.0005
R2861 VD1.n17 VD1.t3 16.0005
R2862 VD1.n19 VD1.t7 16.0005
R2863 VD1.n19 VD1.t5 16.0005
R2864 VD1.n1 VD1.t0 16.0005
R2865 VD1.n1 VD1.t6 16.0005
R2866 VD1.n0 VD1.t9 16.0005
R2867 VD1.n0 VD1.t1 16.0005
R2868 VD1.n12 VD1.t2 16.0005
R2869 VD1.n12 VD1.t21 16.0005
R2870 VD1.n5 VD1.t18 16.0005
R2871 VD1.n5 VD1.t12 16.0005
R2872 VD1.n4 VD1.t17 16.0005
R2873 VD1.n4 VD1.t14 16.0005
R2874 VD1.n8 VD1.t15 16.0005
R2875 VD1.n8 VD1.t20 16.0005
R2876 VD1.n14 VD1.n13 4.5005
R2877 VD1.n11 VD1.n10 4.5005
R2878 VD1.n16 VD1.n14 3.563
R2879 VD1.n18 VD1.n16 1.313
R2880 VD1.n14 VD1.n2 1.2505
R2881 VD1 VD1.n18 1.2505
R2882 VD1.n10 VD1.n6 0.563
R2883 VD1.n10 VD1.n9 0.563
R2884 VD1.n13 VD1.n11 0.21925
R2885 Vb2.n6 Vb2.n5 621.268
R2886 Vb2.n21 Vb2.t6 611.739
R2887 Vb2.n17 Vb2.t20 611.739
R2888 Vb2.n12 Vb2.t7 611.739
R2889 Vb2.n8 Vb2.t15 611.739
R2890 Vb2.n21 Vb2.t11 421.75
R2891 Vb2.n22 Vb2.t16 421.75
R2892 Vb2.n23 Vb2.t19 421.75
R2893 Vb2.n24 Vb2.t24 421.75
R2894 Vb2.n17 Vb2.t17 421.75
R2895 Vb2.n18 Vb2.t13 421.75
R2896 Vb2.n19 Vb2.t26 421.75
R2897 Vb2.n20 Vb2.t22 421.75
R2898 Vb2.n12 Vb2.t12 421.75
R2899 Vb2.n13 Vb2.t9 421.75
R2900 Vb2.n14 Vb2.t14 421.75
R2901 Vb2.n15 Vb2.t18 421.75
R2902 Vb2.n8 Vb2.t10 421.75
R2903 Vb2.n9 Vb2.t5 421.75
R2904 Vb2.n10 Vb2.t28 421.75
R2905 Vb2.n11 Vb2.t23 421.75
R2906 Vb2.n6 Vb2.t1 288.166
R2907 Vb2.n0 Vb2.t21 262.288
R2908 Vb2.n7 Vb2.n4 172.811
R2909 Vb2.n26 Vb2.n25 169.125
R2910 Vb2.n26 Vb2.n16 169.125
R2911 Vb2.n22 Vb2.n21 167.094
R2912 Vb2.n23 Vb2.n22 167.094
R2913 Vb2.n24 Vb2.n23 167.094
R2914 Vb2.n18 Vb2.n17 167.094
R2915 Vb2.n19 Vb2.n18 167.094
R2916 Vb2.n20 Vb2.n19 167.094
R2917 Vb2.n13 Vb2.n12 167.094
R2918 Vb2.n14 Vb2.n13 167.094
R2919 Vb2.n15 Vb2.n14 167.094
R2920 Vb2.n9 Vb2.n8 167.094
R2921 Vb2.n10 Vb2.n9 167.094
R2922 Vb2.n11 Vb2.n10 167.094
R2923 Vb2.n1 Vb2.n0 167.094
R2924 Vb2.n2 Vb2.n1 167.094
R2925 Vb2.n3 Vb2.n2 167.094
R2926 Vb2.n4 Vb2.t25 142.325
R2927 Vb2.n0 Vb2.t8 72.3005
R2928 Vb2.n1 Vb2.t4 72.3005
R2929 Vb2.n2 Vb2.t27 72.3005
R2930 Vb2.n3 Vb2.t3 72.3005
R2931 Vb2.n5 Vb2.t0 62.5402
R2932 Vb2.n5 Vb2.t2 62.5402
R2933 Vb2.n25 Vb2.n24 47.1294
R2934 Vb2.n25 Vb2.n20 47.1294
R2935 Vb2.n16 Vb2.n15 47.1294
R2936 Vb2.n16 Vb2.n11 47.1294
R2937 Vb2.n4 Vb2.n3 47.1294
R2938 Vb2.n27 Vb2.n7 34.938
R2939 Vb2.n7 Vb2.n6 14.6443
R2940 Vb2.n27 Vb2.n26 4.5005
R2941 Vb2 Vb2.n27 0.063
R2942 Vb2_Vb3.n12 Vb2_Vb3.n7 2445
R2943 Vb2_Vb3.n14 Vb2_Vb3.n6 2430
R2944 Vb2_Vb3.n14 Vb2_Vb3.n7 2430
R2945 Vb2_Vb3.n12 Vb2_Vb3.n6 2415
R2946 Vb2_Vb3.n8 Vb2_Vb3.t3 650.668
R2947 Vb2_Vb3.n18 Vb2_Vb3.t6 650.668
R2948 Vb2_Vb3.n0 Vb2_Vb3.n22 637.288
R2949 Vb2_Vb3.n0 Vb2_Vb3.n23 636.663
R2950 Vb2_Vb3.n0 Vb2_Vb3.n24 636.663
R2951 Vb2_Vb3.n2 Vb2_Vb3.n3 628.668
R2952 Vb2_Vb3.n1 Vb2_Vb3.n19 628.668
R2953 Vb2_Vb3.n21 Vb2_Vb3.n20 624.168
R2954 Vb2_Vb3.n14 Vb2_Vb3.t5 387.329
R2955 Vb2_Vb3.t2 Vb2_Vb3.n12 356.495
R2956 Vb2_Vb3.n9 Vb2_Vb3.t1 310.659
R2957 Vb2_Vb3.n17 Vb2_Vb3.t4 310.659
R2958 Vb2_Vb3.n15 Vb2_Vb3.n5 259.2
R2959 Vb2_Vb3.n11 Vb2_Vb3.n5 257.601
R2960 Vb2_Vb3.t16 Vb2_Vb3.t2 196.553
R2961 Vb2_Vb3.t18 Vb2_Vb3.t16 196.553
R2962 Vb2_Vb3.t20 Vb2_Vb3.t18 196.553
R2963 Vb2_Vb3.t22 Vb2_Vb3.t12 196.553
R2964 Vb2_Vb3.t14 Vb2_Vb3.t22 196.553
R2965 Vb2_Vb3.t5 Vb2_Vb3.t14 196.553
R2966 Vb2_Vb3.n10 Vb2_Vb3.n4 153.601
R2967 Vb2_Vb3.n16 Vb2_Vb3.n4 153.601
R2968 Vb2_Vb3.n11 Vb2_Vb3.n10 107.201
R2969 Vb2_Vb3.n16 Vb2_Vb3.n15 105.6
R2970 Vb2_Vb3.n13 Vb2_Vb3.t20 98.2764
R2971 Vb2_Vb3.t12 Vb2_Vb3.n13 98.2764
R2972 Vb2_Vb3.n6 Vb2_Vb3.n5 92.5005
R2973 Vb2_Vb3.n13 Vb2_Vb3.n6 92.5005
R2974 Vb2_Vb3.n15 Vb2_Vb3.n14 92.5005
R2975 Vb2_Vb3.n7 Vb2_Vb3.n4 92.5005
R2976 Vb2_Vb3.n13 Vb2_Vb3.n7 92.5005
R2977 Vb2_Vb3.n20 Vb2_Vb3.t21 65.6672
R2978 Vb2_Vb3.n20 Vb2_Vb3.t13 65.6672
R2979 Vb2_Vb3.n3 Vb2_Vb3.t17 65.6672
R2980 Vb2_Vb3.n3 Vb2_Vb3.t19 65.6672
R2981 Vb2_Vb3.n19 Vb2_Vb3.t23 65.6672
R2982 Vb2_Vb3.n19 Vb2_Vb3.t15 65.6672
R2983 Vb2_Vb3.n12 Vb2_Vb3.n11 61.6672
R2984 Vb2_Vb3.n23 Vb2_Vb3.t0 49.2505
R2985 Vb2_Vb3.n23 Vb2_Vb3.t8 49.2505
R2986 Vb2_Vb3.n22 Vb2_Vb3.t7 49.2505
R2987 Vb2_Vb3.n22 Vb2_Vb3.t10 49.2505
R2988 Vb2_Vb3.n24 Vb2_Vb3.t11 49.2505
R2989 Vb2_Vb3.n24 Vb2_Vb3.t9 49.2505
R2990 Vb2_Vb3.n1 Vb2_Vb3.n18 44.2922
R2991 Vb2_Vb3.n8 Vb2_Vb3.n2 44.2922
R2992 Vb2_Vb3.n18 Vb2_Vb3.n17 27.7338
R2993 Vb2_Vb3.n9 Vb2_Vb3.n8 27.7338
R2994 Vb2_Vb3.n17 Vb2_Vb3.n16 21.3338
R2995 Vb2_Vb3.n10 Vb2_Vb3.n9 21.3338
R2996 Vb2_Vb3 Vb2_Vb3.n21 7.188
R2997 Vb2_Vb3.n21 Vb2_Vb3.n2 4.5005
R2998 Vb2_Vb3 Vb2_Vb3.n0 2.313
R2999 Vb2_Vb3.n2 Vb2_Vb3.n1 1.2505
R3000 Vb3.n11 Vb3.n9 629.293
R3001 Vb3.n15 Vb3.n14 628.668
R3002 Vb3.n13 Vb3.n12 628.668
R3003 Vb3.n11 Vb3.n10 628.668
R3004 Vb3.n24 Vb3.t9 611.739
R3005 Vb3.n20 Vb3.t24 611.739
R3006 Vb3.n4 Vb3.t10 611.739
R3007 Vb3.n0 Vb3.t18 611.739
R3008 Vb3.n24 Vb3.t13 421.75
R3009 Vb3.n25 Vb3.t19 421.75
R3010 Vb3.n26 Vb3.t23 421.75
R3011 Vb3.n27 Vb3.t28 421.75
R3012 Vb3.n20 Vb3.t20 421.75
R3013 Vb3.n21 Vb3.t15 421.75
R3014 Vb3.n22 Vb3.t29 421.75
R3015 Vb3.n23 Vb3.t25 421.75
R3016 Vb3.n4 Vb3.t14 421.75
R3017 Vb3.n5 Vb3.t11 421.75
R3018 Vb3.n6 Vb3.t16 421.75
R3019 Vb3.n7 Vb3.t21 421.75
R3020 Vb3.n0 Vb3.t12 421.75
R3021 Vb3.n1 Vb3.t8 421.75
R3022 Vb3.n2 Vb3.t30 421.75
R3023 Vb3.n3 Vb3.t26 421.75
R3024 Vb3.n17 Vb3.t17 286.389
R3025 Vb3.n16 Vb3.t31 286.389
R3026 Vb3.n30 Vb3.n8 169.343
R3027 Vb3.n25 Vb3.n24 167.094
R3028 Vb3.n26 Vb3.n25 167.094
R3029 Vb3.n27 Vb3.n26 167.094
R3030 Vb3.n21 Vb3.n20 167.094
R3031 Vb3.n22 Vb3.n21 167.094
R3032 Vb3.n23 Vb3.n22 167.094
R3033 Vb3.n5 Vb3.n4 167.094
R3034 Vb3.n6 Vb3.n5 167.094
R3035 Vb3.n7 Vb3.n6 167.094
R3036 Vb3.n1 Vb3.n0 167.094
R3037 Vb3.n2 Vb3.n1 167.094
R3038 Vb3.n3 Vb3.n2 167.094
R3039 Vb3.n29 Vb3.n28 166.25
R3040 Vb3.n19 Vb3.n18 165.8
R3041 Vb3.n17 Vb3.t22 96.4005
R3042 Vb3.n16 Vb3.t27 96.4005
R3043 Vb3.n14 Vb3.t3 65.6672
R3044 Vb3.n14 Vb3.t1 65.6672
R3045 Vb3.n12 Vb3.t2 65.6672
R3046 Vb3.n12 Vb3.t7 65.6672
R3047 Vb3.n10 Vb3.t5 65.6672
R3048 Vb3.n10 Vb3.t6 65.6672
R3049 Vb3.n9 Vb3.t0 65.6672
R3050 Vb3.n9 Vb3.t4 65.6672
R3051 Vb3.n28 Vb3.n27 47.1294
R3052 Vb3.n28 Vb3.n23 47.1294
R3053 Vb3.n8 Vb3.n7 47.1294
R3054 Vb3.n8 Vb3.n3 47.1294
R3055 Vb3.n18 Vb3.n17 38.5605
R3056 Vb3.n18 Vb3.n16 38.5605
R3057 Vb3.n29 Vb3.n19 26.8755
R3058 Vb3 Vb3.n30 4.563
R3059 Vb3.n19 Vb3.n15 3.688
R3060 Vb3.n30 Vb3.n29 3.09425
R3061 Vb3.n13 Vb3.n11 0.6255
R3062 Vb3.n15 Vb3.n13 0.6255
R3063 V_tot.n1 V_tot.t12 327.623
R3064 V_tot.n4 V_tot.t11 326.365
R3065 V_tot.n0 V_tot.t5 168.701
R3066 V_tot.n0 V_tot.t10 168.701
R3067 V_tot.n8 V_tot.n7 165.8
R3068 V_tot.n6 V_tot.n5 165.8
R3069 V_tot.n3 V_tot.n2 165.8
R3070 V_tot.n1 V_tot.n0 165.8
R3071 V_tot.n7 V_tot.t13 157.989
R3072 V_tot.n7 V_tot.t8 157.989
R3073 V_tot.n5 V_tot.t4 157.989
R3074 V_tot.n5 V_tot.t6 157.989
R3075 V_tot.n2 V_tot.t7 157.989
R3076 V_tot.n2 V_tot.t9 157.989
R3077 V_tot.n9 V_tot.t1 117.591
R3078 V_tot.t0 V_tot.n11 117.591
R3079 V_tot.n11 V_tot.t2 108.424
R3080 V_tot.n9 V_tot.t3 108.424
R3081 V_tot.n11 V_tot.n10 42.6121
R3082 V_tot.n10 V_tot.n9 21.2996
R3083 V_tot.n10 V_tot.n8 17.0005
R3084 V_tot.n4 V_tot.n3 3.31612
R3085 V_tot.n3 V_tot.n1 1.26612
R3086 V_tot.n8 V_tot.n6 1.2505
R3087 V_tot.n6 V_tot.n4 1.15363
R3088 V_err_p.n11 V_err_p.n9 630.827
R3089 V_err_p.n15 V_err_p.n14 630.264
R3090 V_err_p.n13 V_err_p.n12 630.264
R3091 V_err_p.n11 V_err_p.n10 630.264
R3092 V_err_p.n2 V_err_p.n0 627.784
R3093 V_err_p.n19 V_err_p.n18 627.784
R3094 V_err_p.n16 V_err_p.n8 627.168
R3095 V_err_p.n6 V_err_p.n5 626.534
R3096 V_err_p.n4 V_err_p.n3 626.534
R3097 V_err_p.n2 V_err_p.n1 626.534
R3098 V_err_p.n17 V_err_p.n7 622.034
R3099 V_err_p.n7 V_err_p.t9 78.8005
R3100 V_err_p.n7 V_err_p.t10 78.8005
R3101 V_err_p.n14 V_err_p.t4 78.8005
R3102 V_err_p.n14 V_err_p.t21 78.8005
R3103 V_err_p.n12 V_err_p.t19 78.8005
R3104 V_err_p.n12 V_err_p.t3 78.8005
R3105 V_err_p.n10 V_err_p.t0 78.8005
R3106 V_err_p.n10 V_err_p.t18 78.8005
R3107 V_err_p.n9 V_err_p.t20 78.8005
R3108 V_err_p.n9 V_err_p.t2 78.8005
R3109 V_err_p.n8 V_err_p.t17 78.8005
R3110 V_err_p.n8 V_err_p.t1 78.8005
R3111 V_err_p.n5 V_err_p.t15 78.8005
R3112 V_err_p.n5 V_err_p.t13 78.8005
R3113 V_err_p.n3 V_err_p.t7 78.8005
R3114 V_err_p.n3 V_err_p.t11 78.8005
R3115 V_err_p.n1 V_err_p.t12 78.8005
R3116 V_err_p.n1 V_err_p.t8 78.8005
R3117 V_err_p.n0 V_err_p.t14 78.8005
R3118 V_err_p.n0 V_err_p.t5 78.8005
R3119 V_err_p.n19 V_err_p.t6 78.8005
R3120 V_err_p.t16 V_err_p.n19 78.8005
R3121 V_err_p.n16 V_err_p.n15 5.0005
R3122 V_err_p.n18 V_err_p.n17 4.5005
R3123 V_err_p.n17 V_err_p.n16 1.3272
R3124 V_err_p.n4 V_err_p.n2 1.2505
R3125 V_err_p.n6 V_err_p.n4 1.2505
R3126 V_err_p.n18 V_err_p.n6 1.2505
R3127 V_err_p.n13 V_err_p.n11 0.563
R3128 V_err_p.n15 V_err_p.n13 0.563
R3129 VIN+.n9 VIN+.t9 485.127
R3130 VIN+.n4 VIN+.t5 485.127
R3131 VIN+.n3 VIN+.t0 485.127
R3132 VIN+.n7 VIN+.t2 318.656
R3133 VIN+.n7 VIN+.t7 318.656
R3134 VIN+.n5 VIN+.t1 318.656
R3135 VIN+.n5 VIN+.t6 318.656
R3136 VIN+.n1 VIN+.t4 318.656
R3137 VIN+.n1 VIN+.t10 318.656
R3138 VIN+.n0 VIN+.t3 318.656
R3139 VIN+.n0 VIN+.t8 318.656
R3140 VIN+.n2 VIN+.n0 167.05
R3141 VIN+.n8 VIN+.n7 165.8
R3142 VIN+.n6 VIN+.n5 165.8
R3143 VIN+.n2 VIN+.n1 165.8
R3144 VIN+.n6 VIN+.n4 2.34425
R3145 VIN+.n4 VIN+.n3 1.3005
R3146 VIN+.n8 VIN+.n6 1.2505
R3147 VIN+ VIN+.n9 1.213
R3148 VIN+.n3 VIN+.n2 1.15675
R3149 VIN+.n9 VIN+.n8 1.15675
R3150 VD2.n12 VD2.n10 114.719
R3151 VD2.n9 VD2.n7 114.719
R3152 VD2.n12 VD2.n11 114.156
R3153 VD2.n9 VD2.n8 114.156
R3154 VD2.n5 VD2.n3 112.456
R3155 VD2.n2 VD2.n0 112.456
R3156 VD2.n5 VD2.n4 111.206
R3157 VD2.n2 VD2.n1 111.206
R3158 VD2.n19 VD2.n18 111.204
R3159 VD2.n14 VD2.n6 109.656
R3160 VD2.n16 VD2.n15 106.706
R3161 VD2.n11 VD2.t19 16.0005
R3162 VD2.n11 VD2.t14 16.0005
R3163 VD2.n10 VD2.t17 16.0005
R3164 VD2.n10 VD2.t12 16.0005
R3165 VD2.n8 VD2.t20 16.0005
R3166 VD2.n8 VD2.t15 16.0005
R3167 VD2.n7 VD2.t21 16.0005
R3168 VD2.n7 VD2.t16 16.0005
R3169 VD2.n6 VD2.t18 16.0005
R3170 VD2.n6 VD2.t13 16.0005
R3171 VD2.n15 VD2.t4 16.0005
R3172 VD2.n15 VD2.t8 16.0005
R3173 VD2.n4 VD2.t3 16.0005
R3174 VD2.n4 VD2.t7 16.0005
R3175 VD2.n3 VD2.t1 16.0005
R3176 VD2.n3 VD2.t11 16.0005
R3177 VD2.n1 VD2.t0 16.0005
R3178 VD2.n1 VD2.t5 16.0005
R3179 VD2.n0 VD2.t2 16.0005
R3180 VD2.n0 VD2.t6 16.0005
R3181 VD2.t9 VD2.n19 16.0005
R3182 VD2.n19 VD2.t10 16.0005
R3183 VD2.n14 VD2.n13 4.5005
R3184 VD2.n17 VD2.n16 4.5005
R3185 VD2.n18 VD2.n17 3.6255
R3186 VD2.n17 VD2.n5 1.2505
R3187 VD2.n18 VD2.n2 1.2505
R3188 VD2.n16 VD2.n14 0.78175
R3189 VD2.n13 VD2.n12 0.563
R3190 VD2.n13 VD2.n9 0.563
R3191 V_CMFB_S3.n2 V_CMFB_S3.n1 205.552
R3192 V_CMFB_S3.n4 V_CMFB_S3.n3 205.488
R3193 V_CMFB_S3.n6 V_CMFB_S3.n5 205.488
R3194 V_CMFB_S3.n8 V_CMFB_S3.n7 205.488
R3195 V_CMFB_S3.n10 V_CMFB_S3.n9 205.488
R3196 V_CMFB_S3 V_CMFB_S3.t0 126.974
R3197 V_CMFB_S3.n1 V_CMFB_S3.t1 19.7005
R3198 V_CMFB_S3.n1 V_CMFB_S3.t6 19.7005
R3199 V_CMFB_S3.n3 V_CMFB_S3.t5 19.7005
R3200 V_CMFB_S3.n3 V_CMFB_S3.t9 19.7005
R3201 V_CMFB_S3.n5 V_CMFB_S3.t2 19.7005
R3202 V_CMFB_S3.n5 V_CMFB_S3.t10 19.7005
R3203 V_CMFB_S3.n7 V_CMFB_S3.t3 19.7005
R3204 V_CMFB_S3.n7 V_CMFB_S3.t7 19.7005
R3205 V_CMFB_S3.n9 V_CMFB_S3.t4 19.7005
R3206 V_CMFB_S3.n9 V_CMFB_S3.t8 19.7005
R3207 V_CMFB_S3.n2 V_CMFB_S3.n0 2.188
R3208 V_CMFB_S3 V_CMFB_S3.n10 1.6255
R3209 V_CMFB_S3.n10 V_CMFB_S3.n8 0.563
R3210 V_CMFB_S3.n8 V_CMFB_S3.n6 0.563
R3211 V_CMFB_S3.n6 V_CMFB_S3.n4 0.563
R3212 V_CMFB_S3.n4 V_CMFB_S3.n2 0.5005
R3213 V_CMFB_S1.n2 V_CMFB_S1.n0 206.052
R3214 V_CMFB_S1.n8 V_CMFB_S1.n7 205.488
R3215 V_CMFB_S1.n6 V_CMFB_S1.n5 205.488
R3216 V_CMFB_S1.n4 V_CMFB_S1.n3 205.488
R3217 V_CMFB_S1.n2 V_CMFB_S1.n1 205.488
R3218 V_CMFB_S1 V_CMFB_S1.t0 127.004
R3219 V_CMFB_S1.n7 V_CMFB_S1.t5 19.7005
R3220 V_CMFB_S1.n7 V_CMFB_S1.t9 19.7005
R3221 V_CMFB_S1.n5 V_CMFB_S1.t6 19.7005
R3222 V_CMFB_S1.n5 V_CMFB_S1.t10 19.7005
R3223 V_CMFB_S1.n3 V_CMFB_S1.t7 19.7005
R3224 V_CMFB_S1.n3 V_CMFB_S1.t1 19.7005
R3225 V_CMFB_S1.n1 V_CMFB_S1.t8 19.7005
R3226 V_CMFB_S1.n1 V_CMFB_S1.t2 19.7005
R3227 V_CMFB_S1.n0 V_CMFB_S1.t4 19.7005
R3228 V_CMFB_S1.n0 V_CMFB_S1.t3 19.7005
R3229 V_CMFB_S1 V_CMFB_S1.n8 1.59425
R3230 V_CMFB_S1.n4 V_CMFB_S1.n2 0.563
R3231 V_CMFB_S1.n6 V_CMFB_S1.n4 0.563
R3232 V_CMFB_S1.n8 V_CMFB_S1.n6 0.563
R3233 VIN-.n4 VIN-.t1 485.021
R3234 VIN-.n1 VIN-.t2 484.159
R3235 VIN-.n5 VIN-.t0 483.358
R3236 VIN-.n8 VIN-.t3 431.536
R3237 VIN-.n2 VIN-.t6 431.536
R3238 VIN-.n6 VIN-.t9 431.257
R3239 VIN-.n0 VIN-.t4 431.257
R3240 VIN-.n6 VIN-.t5 289.908
R3241 VIN-.n0 VIN-.t8 289.908
R3242 VIN-.n8 VIN-.t7 279.183
R3243 VIN-.n2 VIN-.t10 279.183
R3244 VIN-.n7 VIN-.n6 233.374
R3245 VIN-.n1 VIN-.n0 233.374
R3246 VIN-.n9 VIN-.n8 188.989
R3247 VIN-.n3 VIN-.n2 188.989
R3248 VIN-.n4 VIN-.n3 2.463
R3249 VIN- VIN-.n9 2.03175
R3250 VIN-.n5 VIN-.n4 1.563
R3251 VIN-.n3 VIN-.n1 1.2755
R3252 VIN-.n9 VIN-.n7 1.2755
R3253 VIN-.n7 VIN-.n5 0.8005
R3254 err_amp_out.n7 err_amp_out.n6 630.607
R3255 err_amp_out.n9 err_amp_out.n8 627.128
R3256 err_amp_out err_amp_out.n10 627.128
R3257 err_amp_out.n5 err_amp_out.t12 410.666
R3258 err_amp_out.n2 err_amp_out.n0 227.784
R3259 err_amp_out.n2 err_amp_out.n1 226.534
R3260 err_amp_out.n4 err_amp_out.n3 226.534
R3261 err_amp_out.n6 err_amp_out.t0 78.8005
R3262 err_amp_out.n6 err_amp_out.t2 78.8005
R3263 err_amp_out.n8 err_amp_out.t5 78.8005
R3264 err_amp_out.n8 err_amp_out.t3 78.8005
R3265 err_amp_out.n10 err_amp_out.t4 78.8005
R3266 err_amp_out.n10 err_amp_out.t6 78.8005
R3267 err_amp_out.n1 err_amp_out.t10 48.0005
R3268 err_amp_out.n1 err_amp_out.t7 48.0005
R3269 err_amp_out.n3 err_amp_out.t1 48.0005
R3270 err_amp_out.n3 err_amp_out.t9 48.0005
R3271 err_amp_out.n0 err_amp_out.t8 48.0005
R3272 err_amp_out.n0 err_amp_out.t11 48.0005
R3273 err_amp_out.n7 err_amp_out.n5 21.1255
R3274 err_amp_out.n5 err_amp_out.n4 10.8755
R3275 err_amp_out.n9 err_amp_out.n7 1.3755
R3276 err_amp_out.n4 err_amp_out.n2 1.2505
R3277 err_amp_out err_amp_out.n9 1.2505
R3278 a_59060_4632.t0 a_59060_4632.t1 169.905
R3279 VD3.n22 VD3.n15 4020
R3280 VD3.n24 VD3.n15 4020
R3281 VD3.n22 VD3.n21 4020
R3282 VD3.n24 VD3.n21 4020
R3283 VD3.n18 VD3.t0 660.109
R3284 VD3.n16 VD3.t3 660.109
R3285 VD3.n26 VD3.n25 428.8
R3286 VD3.n26 VD3.n14 428.8
R3287 VD3.t1 VD3.n22 239.915
R3288 VD3.n24 VD3.t4 239.915
R3289 VD3.n20 VD3.n19 230.4
R3290 VD3.n20 VD3.n17 230.4
R3291 VD3.n25 VD3.n17 198.4
R3292 VD3.n19 VD3.n14 198.4
R3293 VD3.n13 VD3.n11 160.428
R3294 VD3.n8 VD3.n7 160.427
R3295 VD3.n2 VD3.n0 160.427
R3296 VD3.n33 VD3.n32 160.054
R3297 VD3.n31 VD3.n30 159.803
R3298 VD3.n13 VD3.n12 159.803
R3299 VD3.n6 VD3.n5 159.802
R3300 VD3.n4 VD3.n3 159.802
R3301 VD3.n2 VD3.n1 159.802
R3302 VD3.n10 VD3.n9 155.302
R3303 VD3.n18 VD3.t2 155.125
R3304 VD3.n16 VD3.t5 155.125
R3305 VD3.n28 VD3.n27 146.002
R3306 VD3.t24 VD3.t1 98.2764
R3307 VD3.t28 VD3.t24 98.2764
R3308 VD3.t32 VD3.t28 98.2764
R3309 VD3.t18 VD3.t32 98.2764
R3310 VD3.t22 VD3.t18 98.2764
R3311 VD3.t26 VD3.t20 98.2764
R3312 VD3.t30 VD3.t26 98.2764
R3313 VD3.t34 VD3.t30 98.2764
R3314 VD3.t36 VD3.t34 98.2764
R3315 VD3.t4 VD3.t36 98.2764
R3316 VD3.n25 VD3.n24 92.5005
R3317 VD3.n21 VD3.n20 92.5005
R3318 VD3.n23 VD3.n21 92.5005
R3319 VD3.n22 VD3.n14 92.5005
R3320 VD3.n26 VD3.n15 92.5005
R3321 VD3.n23 VD3.n15 92.5005
R3322 VD3.n23 VD3.t22 49.1384
R3323 VD3.t20 VD3.n23 49.1384
R3324 VD3.n19 VD3.n18 21.3338
R3325 VD3.n17 VD3.n16 21.3338
R3326 VD3.n28 VD3.n26 19.2005
R3327 VD3.n29 VD3.n28 13.8005
R3328 VD3.n9 VD3.t12 11.2576
R3329 VD3.n9 VD3.t14 11.2576
R3330 VD3.n7 VD3.t15 11.2576
R3331 VD3.n7 VD3.t17 11.2576
R3332 VD3.n5 VD3.t7 11.2576
R3333 VD3.n5 VD3.t10 11.2576
R3334 VD3.n3 VD3.t6 11.2576
R3335 VD3.n3 VD3.t8 11.2576
R3336 VD3.n1 VD3.t11 11.2576
R3337 VD3.n1 VD3.t13 11.2576
R3338 VD3.n0 VD3.t16 11.2576
R3339 VD3.n0 VD3.t9 11.2576
R3340 VD3.n30 VD3.t27 11.2576
R3341 VD3.n30 VD3.t31 11.2576
R3342 VD3.n27 VD3.t23 11.2576
R3343 VD3.n27 VD3.t21 11.2576
R3344 VD3.n12 VD3.t33 11.2576
R3345 VD3.n12 VD3.t19 11.2576
R3346 VD3.n11 VD3.t25 11.2576
R3347 VD3.n11 VD3.t29 11.2576
R3348 VD3.n32 VD3.t35 11.2576
R3349 VD3.n32 VD3.t37 11.2576
R3350 VD3 VD3.n33 5.40675
R3351 VD3.n10 VD3.n8 4.5005
R3352 VD3 VD3.n10 0.78175
R3353 VD3.n4 VD3.n2 0.6255
R3354 VD3.n6 VD3.n4 0.6255
R3355 VD3.n8 VD3.n6 0.6255
R3356 VD3.n29 VD3.n13 0.6255
R3357 VD3.n31 VD3.n29 0.6255
R3358 VD3.n33 VD3.n31 0.2505
R3359 V_p_mir.n1 V_p_mir.n0 220.678
R3360 V_p_mir.n0 V_p_mir.t1 16.0005
R3361 V_p_mir.n0 V_p_mir.t0 16.0005
R3362 V_p_mir.t2 V_p_mir.n1 9.6005
R3363 V_p_mir.n1 V_p_mir.t3 9.6005
R3364 V_b_2nd_stage.n4 V_b_2nd_stage.t7 525.38
R3365 V_b_2nd_stage.n0 V_b_2nd_stage.t2 525.38
R3366 V_b_2nd_stage.n6 V_b_2nd_stage.t4 366.856
R3367 V_b_2nd_stage.n2 V_b_2nd_stage.t5 366.856
R3368 V_b_2nd_stage.n4 V_b_2nd_stage.t3 281.168
R3369 V_b_2nd_stage.n5 V_b_2nd_stage.t8 281.168
R3370 V_b_2nd_stage.n0 V_b_2nd_stage.t6 281.168
R3371 V_b_2nd_stage.n1 V_b_2nd_stage.t9 281.168
R3372 V_b_2nd_stage.n5 V_b_2nd_stage.n4 244.214
R3373 V_b_2nd_stage.n1 V_b_2nd_stage.n0 244.214
R3374 V_b_2nd_stage.n7 V_b_2nd_stage.n6 166.03
R3375 V_b_2nd_stage.n3 V_b_2nd_stage.n2 166.03
R3376 V_b_2nd_stage.n3 V_b_2nd_stage.t1 117.849
R3377 V_b_2nd_stage.t0 V_b_2nd_stage.n7 117.849
R3378 V_b_2nd_stage.n6 V_b_2nd_stage.n5 85.6894
R3379 V_b_2nd_stage.n2 V_b_2nd_stage.n1 85.6894
R3380 V_b_2nd_stage.n7 V_b_2nd_stage.n3 39.5005
R3381 a_67950_1836.t0 a_67950_1836.t1 169.905
R3382 a_68230_5092.t0 a_68230_5092.t1 291.183
R3383 a_59460_1836.t0 a_59460_1836.t1 169.905
R3384 a_68350_4632.t0 a_68350_4632.t1 169.905
C0 Vb2_Vb3 VOUT+ 0.03526f
C1 Vb2_Vb3 VDDA 1.65337f
C2 Vb2 V_err_gate 0.045935f
C3 VDDA V_CMFB_S4 2.27197f
C4 Vb2_Vb3 Vb3 1.18941f
C5 VD3 VDDA 3.78008f
C6 Vb2 V_err_amp_ref 0.039506f
C7 Vb2_Vb3 cap_res_X 0.014914f
C8 VOUT- VOUT+ 0.210644f
C9 VDDA VOUT- 6.76964f
C10 VIN- VIN+ 0.555219f
C11 VD3 Vb3 1.2438f
C12 V_err_gate V_err_amp_ref 1.21744f
C13 VOUT- V_CMFB_S1 0.063238f
C14 Vb3 VOUT- 0.012148f
C15 VDDA VOUT+ 6.69701f
C16 V_CMFB_S3 V_CMFB_S4 1.19888f
C17 cap_res_X VOUT- 50.7541f
C18 VDDA err_amp_out 1.00936f
C19 V_CMFB_S2 VDDA 2.27175f
C20 VDDA V_CMFB_S1 0.593809f
C21 VDDA Vb3 6.3346f
C22 cap_res_X VOUT+ 0.020189f
C23 VDDA cap_res_X 0.659054f
C24 VD3 Vb1 0.028096f
C25 Vb2_Vb3 Vb2 0.795916f
C26 V_tail_gate VIN- 0.230373f
C27 Y V_CMFB_S4 0.715786f
C28 V_CMFB_S3 VOUT+ 0.061977f
C29 Vb1 VOUT- 0.013066f
C30 V_CMFB_S2 V_CMFB_S1 1.20062f
C31 V_CMFB_S3 VDDA 0.592955f
C32 Vb1 VIN- 0.038504f
C33 Vb3 cap_res_X 0.012315f
C34 Vb2_Vb3 V_err_gate 0.012774f
C35 V_tail_gate VIN+ 0.107855f
C36 VD3 Vb2 2.18512f
C37 Vb1 VDDA 0.335789f
C38 VOUT- Vb2 0.011026f
C39 Vb1 VIN+ 0.021067f
C40 VD1 VIN- 0.881219f
C41 Y VOUT+ 2.11549f
C42 VDDA Y 4.15645f
C43 VD3 V_err_gate 0.011317f
C44 Y err_amp_out 0.040365f
C45 VDDA Vb2 1.6078f
C46 Vb1 cap_res_X 0.027198f
C47 VD1 VIN+ 0.057219f
C48 err_amp_out VD1 0.017581f
C49 Vb3 Y 0.010233f
C50 VDDA V_err_gate 3.27456f
C51 Vb3 Vb2 2.95326f
C52 Vb1 V_tail_gate 0.015387f
C53 V_CMFB_S3 Y 0.629597f
C54 Vb3 V_err_gate 0.019752f
C55 VDDA V_err_amp_ref 2.09177f
C56 Vb1 Y 0.840154f
C57 err_amp_out V_err_amp_ref 0.406563f
C58 V_tail_gate VD1 0.213374f
C59 Vb1 Vb2 0.056219f
C60 Vb1 VD1 0.395378f
C61 Vb3 V_err_amp_ref 0.051187f
C62 Y Vb2 1.51102f
C63 Y VD1 1.06369f
C64 V_tail_gate GNDA 3.86357f
C65 VIN+ GNDA 2.09054f
C66 VIN- GNDA 2.185862f
C67 V_CMFB_S4 GNDA 1.652507f
C68 Vb1 GNDA 5.64729f
C69 V_CMFB_S3 GNDA 2.3321f
C70 V_CMFB_S2 GNDA 1.660983f
C71 V_CMFB_S1 GNDA 2.32262f
C72 VOUT+ GNDA 17.930159f
C73 VOUT- GNDA 17.928366f
C74 V_err_amp_ref GNDA 0.557195f
C75 V_err_gate GNDA 1.075647f
C76 Vb2 GNDA 2.33068f
C77 Vb3 GNDA 1.674793f
C78 VDDA GNDA 72.25549f
C79 VD1 GNDA 2.41268f
C80 Y GNDA 4.986685f
C81 cap_res_X GNDA 33.82925f
C82 err_amp_out GNDA 3.001013f
C83 VD3 GNDA 6.547144f
C84 Vb2_Vb3 GNDA 3.42409f
C85 V_b_2nd_stage.t1 GNDA 0.163765f
C86 V_b_2nd_stage.t9 GNDA 0.409099f
C87 V_b_2nd_stage.t6 GNDA 0.409099f
C88 V_b_2nd_stage.t2 GNDA 0.485537f
C89 V_b_2nd_stage.n0 GNDA 0.256456f
C90 V_b_2nd_stage.n1 GNDA 0.162306f
C91 V_b_2nd_stage.t5 GNDA 0.446073f
C92 V_b_2nd_stage.n2 GNDA 0.149996f
C93 V_b_2nd_stage.n3 GNDA 0.917914f
C94 V_b_2nd_stage.t4 GNDA 0.446073f
C95 V_b_2nd_stage.t8 GNDA 0.409099f
C96 V_b_2nd_stage.t3 GNDA 0.409099f
C97 V_b_2nd_stage.t7 GNDA 0.485537f
C98 V_b_2nd_stage.n4 GNDA 0.256456f
C99 V_b_2nd_stage.n5 GNDA 0.162306f
C100 V_b_2nd_stage.n6 GNDA 0.149996f
C101 V_b_2nd_stage.n7 GNDA 0.917423f
C102 V_b_2nd_stage.t0 GNDA 0.163765f
C103 VD3.t16 GNDA 0.032109f
C104 VD3.t9 GNDA 0.032109f
C105 VD3.n0 GNDA 0.111667f
C106 VD3.t11 GNDA 0.032109f
C107 VD3.t13 GNDA 0.032109f
C108 VD3.n1 GNDA 0.111271f
C109 VD3.n2 GNDA 0.210069f
C110 VD3.t6 GNDA 0.032109f
C111 VD3.t8 GNDA 0.032109f
C112 VD3.n3 GNDA 0.111271f
C113 VD3.n4 GNDA 0.108902f
C114 VD3.t7 GNDA 0.032109f
C115 VD3.t10 GNDA 0.032109f
C116 VD3.n5 GNDA 0.111271f
C117 VD3.n6 GNDA 0.108902f
C118 VD3.t15 GNDA 0.032109f
C119 VD3.t17 GNDA 0.032109f
C120 VD3.n7 GNDA 0.111667f
C121 VD3.n8 GNDA 0.130524f
C122 VD3.t12 GNDA 0.032109f
C123 VD3.t14 GNDA 0.032109f
C124 VD3.n9 GNDA 0.108966f
C125 VD3.n10 GNDA 0.091263f
C126 VD3.t25 GNDA 0.032109f
C127 VD3.t29 GNDA 0.032109f
C128 VD3.n11 GNDA 0.111667f
C129 VD3.t33 GNDA 0.032109f
C130 VD3.t19 GNDA 0.032109f
C131 VD3.n12 GNDA 0.111271f
C132 VD3.n13 GNDA 0.210069f
C133 VD3.n14 GNDA 0.091409f
C134 VD3.n15 GNDA 0.124299f
C135 VD3.t5 GNDA 0.158399f
C136 VD3.t3 GNDA 0.055912f
C137 VD3.n16 GNDA 0.103335f
C138 VD3.n17 GNDA 0.066614f
C139 VD3.t2 GNDA 0.158399f
C140 VD3.t0 GNDA 0.055912f
C141 VD3.n18 GNDA 0.103335f
C142 VD3.n19 GNDA 0.066614f
C143 VD3.n20 GNDA 0.066052f
C144 VD3.n21 GNDA 0.124299f
C145 VD3.n22 GNDA 0.370433f
C146 VD3.t1 GNDA 0.552924f
C147 VD3.t24 GNDA 0.319251f
C148 VD3.t28 GNDA 0.319251f
C149 VD3.t32 GNDA 0.319251f
C150 VD3.t18 GNDA 0.319251f
C151 VD3.t22 GNDA 0.239438f
C152 VD3.n23 GNDA 0.159625f
C153 VD3.t20 GNDA 0.239438f
C154 VD3.t26 GNDA 0.319251f
C155 VD3.t30 GNDA 0.319251f
C156 VD3.t34 GNDA 0.319251f
C157 VD3.t36 GNDA 0.319251f
C158 VD3.t4 GNDA 0.552924f
C159 VD3.n24 GNDA 0.370433f
C160 VD3.n25 GNDA 0.091409f
C161 VD3.n26 GNDA 0.127969f
C162 VD3.t23 GNDA 0.032109f
C163 VD3.t21 GNDA 0.032109f
C164 VD3.n27 GNDA 0.104687f
C165 VD3.n28 GNDA 0.076237f
C166 VD3.n29 GNDA 0.039248f
C167 VD3.t27 GNDA 0.032109f
C168 VD3.t31 GNDA 0.032109f
C169 VD3.n30 GNDA 0.111271f
C170 VD3.n31 GNDA 0.103398f
C171 VD3.t35 GNDA 0.032109f
C172 VD3.t37 GNDA 0.032109f
C173 VD3.n32 GNDA 0.111421f
C174 VD3.n33 GNDA 0.118607f
C175 err_amp_out.t8 GNDA 0.013323f
C176 err_amp_out.t11 GNDA 0.013323f
C177 err_amp_out.n0 GNDA 0.038344f
C178 err_amp_out.t10 GNDA 0.013323f
C179 err_amp_out.t7 GNDA 0.013323f
C180 err_amp_out.n1 GNDA 0.037203f
C181 err_amp_out.n2 GNDA 0.462683f
C182 err_amp_out.t1 GNDA 0.013323f
C183 err_amp_out.t9 GNDA 0.013323f
C184 err_amp_out.n3 GNDA 0.037203f
C185 err_amp_out.n4 GNDA 0.493922f
C186 err_amp_out.t12 GNDA 0.059015f
C187 err_amp_out.n5 GNDA 1.65781f
C188 err_amp_out.t0 GNDA 0.013323f
C189 err_amp_out.t2 GNDA 0.013323f
C190 err_amp_out.n6 GNDA 0.030943f
C191 err_amp_out.n7 GNDA 0.914249f
C192 err_amp_out.t5 GNDA 0.013323f
C193 err_amp_out.t3 GNDA 0.013323f
C194 err_amp_out.n8 GNDA 0.031191f
C195 err_amp_out.n9 GNDA 0.349833f
C196 err_amp_out.t4 GNDA 0.013323f
C197 err_amp_out.t6 GNDA 0.013323f
C198 err_amp_out.n10 GNDA 0.031191f
C199 VIN-.t2 GNDA 0.050642f
C200 VIN-.t8 GNDA 0.033412f
C201 VIN-.t4 GNDA 0.041251f
C202 VIN-.n0 GNDA 0.059274f
C203 VIN-.n1 GNDA 0.280478f
C204 VIN-.t10 GNDA 0.032863f
C205 VIN-.t6 GNDA 0.041265f
C206 VIN-.n2 GNDA 0.064892f
C207 VIN-.n3 GNDA 0.200879f
C208 VIN-.t1 GNDA 0.050078f
C209 VIN-.n4 GNDA 0.236241f
C210 VIN-.t0 GNDA 0.050425f
C211 VIN-.n5 GNDA 0.180621f
C212 VIN-.t5 GNDA 0.033412f
C213 VIN-.t9 GNDA 0.041251f
C214 VIN-.n6 GNDA 0.059274f
C215 VIN-.n7 GNDA 0.149629f
C216 VIN-.t7 GNDA 0.032863f
C217 VIN-.t3 GNDA 0.041265f
C218 VIN-.n8 GNDA 0.064892f
C219 VIN-.n9 GNDA 0.186141f
C220 VD2.t10 GNDA 0.013877f
C221 VD2.t2 GNDA 0.013877f
C222 VD2.t6 GNDA 0.013877f
C223 VD2.n0 GNDA 0.048872f
C224 VD2.t0 GNDA 0.013877f
C225 VD2.t5 GNDA 0.013877f
C226 VD2.n1 GNDA 0.047884f
C227 VD2.n2 GNDA 0.193373f
C228 VD2.t1 GNDA 0.013877f
C229 VD2.t11 GNDA 0.013877f
C230 VD2.n3 GNDA 0.048872f
C231 VD2.t3 GNDA 0.013877f
C232 VD2.t7 GNDA 0.013877f
C233 VD2.n4 GNDA 0.047884f
C234 VD2.n5 GNDA 0.193373f
C235 VD2.t18 GNDA 0.013877f
C236 VD2.t13 GNDA 0.013877f
C237 VD2.n6 GNDA 0.04687f
C238 VD2.t21 GNDA 0.013877f
C239 VD2.t16 GNDA 0.013877f
C240 VD2.n7 GNDA 0.050131f
C241 VD2.t20 GNDA 0.013877f
C242 VD2.t15 GNDA 0.013877f
C243 VD2.n8 GNDA 0.04969f
C244 VD2.n9 GNDA 0.186051f
C245 VD2.t17 GNDA 0.013877f
C246 VD2.t12 GNDA 0.013877f
C247 VD2.n10 GNDA 0.050131f
C248 VD2.t19 GNDA 0.013877f
C249 VD2.t14 GNDA 0.013877f
C250 VD2.n11 GNDA 0.04969f
C251 VD2.n12 GNDA 0.186051f
C252 VD2.n13 GNDA 0.027755f
C253 VD2.n14 GNDA 0.081264f
C254 VD2.t4 GNDA 0.013877f
C255 VD2.t8 GNDA 0.013877f
C256 VD2.n15 GNDA 0.045463f
C257 VD2.n16 GNDA 0.069533f
C258 VD2.n17 GNDA 0.083264f
C259 VD2.n18 GNDA 0.140662f
C260 VD2.n19 GNDA 0.047884f
C261 VD2.t9 GNDA 0.013877f
C262 VIN+.t8 GNDA 0.041803f
C263 VIN+.t3 GNDA 0.041803f
C264 VIN+.n0 GNDA 0.086391f
C265 VIN+.t10 GNDA 0.041803f
C266 VIN+.t4 GNDA 0.041803f
C267 VIN+.n1 GNDA 0.085194f
C268 VIN+.n2 GNDA 0.359761f
C269 VIN+.t0 GNDA 0.058811f
C270 VIN+.n3 GNDA 0.215335f
C271 VIN+.t5 GNDA 0.058811f
C272 VIN+.n4 GNDA 0.262589f
C273 VIN+.t6 GNDA 0.041803f
C274 VIN+.t1 GNDA 0.041803f
C275 VIN+.n5 GNDA 0.085194f
C276 VIN+.n6 GNDA 0.248358f
C277 VIN+.t7 GNDA 0.041803f
C278 VIN+.t2 GNDA 0.041803f
C279 VIN+.n7 GNDA 0.085194f
C280 VIN+.n8 GNDA 0.200956f
C281 VIN+.t9 GNDA 0.058811f
C282 VIN+.n9 GNDA 0.211601f
C283 V_err_p.n0 GNDA 0.02127f
C284 V_err_p.n1 GNDA 0.020976f
C285 V_err_p.n2 GNDA 0.328367f
C286 V_err_p.n3 GNDA 0.020976f
C287 V_err_p.n4 GNDA 0.180843f
C288 V_err_p.n5 GNDA 0.020976f
C289 V_err_p.n6 GNDA 0.180843f
C290 V_err_p.n7 GNDA 0.020358f
C291 V_err_p.n8 GNDA 0.020407f
C292 V_err_p.n9 GNDA 0.021244f
C293 V_err_p.n10 GNDA 0.021116f
C294 V_err_p.n11 GNDA 0.299998f
C295 V_err_p.n12 GNDA 0.021116f
C296 V_err_p.n13 GNDA 0.156484f
C297 V_err_p.n14 GNDA 0.021116f
C298 V_err_p.n15 GNDA 0.190977f
C299 V_err_p.n16 GNDA 0.153542f
C300 V_err_p.n17 GNDA 0.133374f
C301 V_err_p.n18 GNDA 0.242929f
C302 V_err_p.n19 GNDA 0.02127f
C303 V_tot.t2 GNDA 0.092891f
C304 V_tot.t12 GNDA 0.011218f
C305 V_tot.n0 GNDA 0.018267f
C306 V_tot.n1 GNDA 0.106822f
C307 V_tot.n2 GNDA 0.021464f
C308 V_tot.n3 GNDA 0.095301f
C309 V_tot.t11 GNDA 0.011144f
C310 V_tot.n4 GNDA 0.091464f
C311 V_tot.n5 GNDA 0.021464f
C312 V_tot.n6 GNDA 0.066547f
C313 V_tot.n7 GNDA 0.021464f
C314 V_tot.n8 GNDA 0.204094f
C315 V_tot.t1 GNDA 0.098951f
C316 V_tot.t3 GNDA 0.092891f
C317 V_tot.n9 GNDA 0.321853f
C318 V_tot.n10 GNDA 0.772935f
C319 V_tot.n11 GNDA 0.513063f
C320 V_tot.t0 GNDA 0.098962f
C321 Vb3.t26 GNDA 0.142488f
C322 Vb3.t30 GNDA 0.142488f
C323 Vb3.t8 GNDA 0.142488f
C324 Vb3.t12 GNDA 0.142488f
C325 Vb3.t18 GNDA 0.16443f
C326 Vb3.n0 GNDA 0.133499f
C327 Vb3.n1 GNDA 0.082038f
C328 Vb3.n2 GNDA 0.082038f
C329 Vb3.n3 GNDA 0.076818f
C330 Vb3.t21 GNDA 0.142488f
C331 Vb3.t16 GNDA 0.142488f
C332 Vb3.t11 GNDA 0.142488f
C333 Vb3.t14 GNDA 0.142488f
C334 Vb3.t10 GNDA 0.16443f
C335 Vb3.n4 GNDA 0.133499f
C336 Vb3.n5 GNDA 0.082038f
C337 Vb3.n6 GNDA 0.082038f
C338 Vb3.n7 GNDA 0.076818f
C339 Vb3.n8 GNDA 0.052403f
C340 Vb3.t0 GNDA 0.017271f
C341 Vb3.t4 GNDA 0.017271f
C342 Vb3.n9 GNDA 0.039513f
C343 Vb3.t5 GNDA 0.017271f
C344 Vb3.t6 GNDA 0.017271f
C345 Vb3.n10 GNDA 0.039304f
C346 Vb3.n11 GNDA 0.445078f
C347 Vb3.t2 GNDA 0.017271f
C348 Vb3.t7 GNDA 0.017271f
C349 Vb3.n12 GNDA 0.039304f
C350 Vb3.n13 GNDA 0.234158f
C351 Vb3.t3 GNDA 0.017271f
C352 Vb3.t1 GNDA 0.017271f
C353 Vb3.n14 GNDA 0.039304f
C354 Vb3.n15 GNDA 0.375207f
C355 Vb3.t27 GNDA 0.025907f
C356 Vb3.t31 GNDA 0.046996f
C357 Vb3.n16 GNDA 0.053393f
C358 Vb3.t22 GNDA 0.025907f
C359 Vb3.t17 GNDA 0.046996f
C360 Vb3.n17 GNDA 0.053393f
C361 Vb3.n18 GNDA 0.05186f
C362 Vb3.n19 GNDA 1.21196f
C363 Vb3.t25 GNDA 0.142488f
C364 Vb3.t29 GNDA 0.142488f
C365 Vb3.t15 GNDA 0.142488f
C366 Vb3.t20 GNDA 0.142488f
C367 Vb3.t24 GNDA 0.16443f
C368 Vb3.n20 GNDA 0.133499f
C369 Vb3.n21 GNDA 0.082038f
C370 Vb3.n22 GNDA 0.082038f
C371 Vb3.n23 GNDA 0.076818f
C372 Vb3.t28 GNDA 0.142488f
C373 Vb3.t23 GNDA 0.142488f
C374 Vb3.t19 GNDA 0.142488f
C375 Vb3.t13 GNDA 0.142488f
C376 Vb3.t9 GNDA 0.16443f
C377 Vb3.n24 GNDA 0.133499f
C378 Vb3.n25 GNDA 0.082038f
C379 Vb3.n26 GNDA 0.082038f
C380 Vb3.n27 GNDA 0.076818f
C381 Vb3.n28 GNDA 0.046387f
C382 Vb3.n29 GNDA 1.21075f
C383 Vb3.n30 GNDA 0.643317f
C384 Vb2.t21 GNDA 0.021274f
C385 Vb2.n0 GNDA 0.028404f
C386 Vb2.n1 GNDA 0.022435f
C387 Vb2.n2 GNDA 0.022435f
C388 Vb2.n3 GNDA 0.019529f
C389 Vb2.t25 GNDA 0.01528f
C390 Vb2.n4 GNDA 0.045624f
C391 Vb2.t0 GNDA 0.010096f
C392 Vb2.t2 GNDA 0.010096f
C393 Vb2.n5 GNDA 0.021923f
C394 Vb2.t1 GNDA 0.031354f
C395 Vb2.n6 GNDA 0.106311f
C396 Vb2.n7 GNDA 1.12036f
C397 Vb2.t23 GNDA 0.079325f
C398 Vb2.t28 GNDA 0.079325f
C399 Vb2.t5 GNDA 0.079325f
C400 Vb2.t10 GNDA 0.079325f
C401 Vb2.t15 GNDA 0.09154f
C402 Vb2.n8 GNDA 0.07432f
C403 Vb2.n9 GNDA 0.045672f
C404 Vb2.n10 GNDA 0.045672f
C405 Vb2.n11 GNDA 0.042765f
C406 Vb2.t18 GNDA 0.079325f
C407 Vb2.t14 GNDA 0.079325f
C408 Vb2.t9 GNDA 0.079325f
C409 Vb2.t12 GNDA 0.079325f
C410 Vb2.t7 GNDA 0.09154f
C411 Vb2.n12 GNDA 0.07432f
C412 Vb2.n13 GNDA 0.045672f
C413 Vb2.n14 GNDA 0.045672f
C414 Vb2.n15 GNDA 0.042765f
C415 Vb2.n16 GNDA 0.028605f
C416 Vb2.t22 GNDA 0.079325f
C417 Vb2.t26 GNDA 0.079325f
C418 Vb2.t13 GNDA 0.079325f
C419 Vb2.t17 GNDA 0.079325f
C420 Vb2.t20 GNDA 0.09154f
C421 Vb2.n17 GNDA 0.07432f
C422 Vb2.n18 GNDA 0.045672f
C423 Vb2.n19 GNDA 0.045672f
C424 Vb2.n20 GNDA 0.042765f
C425 Vb2.t24 GNDA 0.079325f
C426 Vb2.t19 GNDA 0.079325f
C427 Vb2.t16 GNDA 0.079325f
C428 Vb2.t11 GNDA 0.079325f
C429 Vb2.t6 GNDA 0.09154f
C430 Vb2.n21 GNDA 0.07432f
C431 Vb2.n22 GNDA 0.045672f
C432 Vb2.n23 GNDA 0.045672f
C433 Vb2.n24 GNDA 0.042765f
C434 Vb2.n25 GNDA 0.028605f
C435 Vb2.n26 GNDA 0.516578f
C436 Vb2.n27 GNDA 0.63715f
C437 V_CMFB_S2.t1 GNDA 0.039423f
C438 V_CMFB_S2.t10 GNDA 0.039423f
C439 V_CMFB_S2.n0 GNDA 0.163029f
C440 V_CMFB_S2.t5 GNDA 0.039423f
C441 V_CMFB_S2.t9 GNDA 0.039423f
C442 V_CMFB_S2.n1 GNDA 0.162404f
C443 V_CMFB_S2.n2 GNDA 0.225173f
C444 V_CMFB_S2.t4 GNDA 0.039423f
C445 V_CMFB_S2.t8 GNDA 0.039423f
C446 V_CMFB_S2.n3 GNDA 0.162404f
C447 V_CMFB_S2.n4 GNDA 0.117499f
C448 V_CMFB_S2.t3 GNDA 0.039423f
C449 V_CMFB_S2.t7 GNDA 0.039423f
C450 V_CMFB_S2.n5 GNDA 0.162404f
C451 V_CMFB_S2.n6 GNDA 0.117499f
C452 V_CMFB_S2.t2 GNDA 0.039423f
C453 V_CMFB_S2.t6 GNDA 0.039423f
C454 V_CMFB_S2.n7 GNDA 0.162404f
C455 V_CMFB_S2.n8 GNDA 0.133268f
C456 V_CMFB_S2.t0 GNDA 0.174042f
C457 V_CMFB_S4.n0 GNDA -0.172147f
C458 V_CMFB_S4.t6 GNDA 0.039423f
C459 V_CMFB_S4.t1 GNDA 0.039423f
C460 V_CMFB_S4.n1 GNDA 0.162465f
C461 V_CMFB_S4.n2 GNDA 0.282193f
C462 V_CMFB_S4.t0 GNDA 0.039423f
C463 V_CMFB_S4.t4 GNDA 0.039423f
C464 V_CMFB_S4.n3 GNDA 0.162404f
C465 V_CMFB_S4.n4 GNDA 0.115692f
C466 V_CMFB_S4.t7 GNDA 0.039423f
C467 V_CMFB_S4.t5 GNDA 0.039423f
C468 V_CMFB_S4.n5 GNDA 0.162404f
C469 V_CMFB_S4.n6 GNDA 0.117499f
C470 V_CMFB_S4.t8 GNDA 0.039423f
C471 V_CMFB_S4.t2 GNDA 0.039423f
C472 V_CMFB_S4.n7 GNDA 0.162404f
C473 V_CMFB_S4.n8 GNDA 0.117499f
C474 V_CMFB_S4.t9 GNDA 0.039423f
C475 V_CMFB_S4.t3 GNDA 0.039423f
C476 V_CMFB_S4.n9 GNDA 0.162404f
C477 V_CMFB_S4.n10 GNDA 0.133925f
C478 V_CMFB_S4.t10 GNDA 0.173892f
C479 Y.t23 GNDA 0.053187f
C480 Y.t0 GNDA 0.053187f
C481 Y.n0 GNDA 0.184972f
C482 Y.t7 GNDA 0.053187f
C483 Y.t5 GNDA 0.053187f
C484 Y.n1 GNDA 0.184316f
C485 Y.n2 GNDA 0.347971f
C486 Y.t6 GNDA 0.053187f
C487 Y.t21 GNDA 0.053187f
C488 Y.n3 GNDA 0.184316f
C489 Y.n4 GNDA 0.180392f
C490 Y.t11 GNDA 0.053187f
C491 Y.t14 GNDA 0.053187f
C492 Y.n5 GNDA 0.184316f
C493 Y.n6 GNDA 0.180392f
C494 Y.t18 GNDA 0.053187f
C495 Y.t16 GNDA 0.053187f
C496 Y.n7 GNDA 0.184316f
C497 Y.n8 GNDA 0.212415f
C498 Y.t15 GNDA 0.053187f
C499 Y.t24 GNDA 0.053187f
C500 Y.n9 GNDA 0.180498f
C501 Y.n10 GNDA 0.149147f
C502 Y.t22 GNDA 0.022794f
C503 Y.t3 GNDA 0.022794f
C504 Y.n11 GNDA 0.076959f
C505 Y.t19 GNDA 0.022794f
C506 Y.t13 GNDA 0.022794f
C507 Y.n12 GNDA 0.082252f
C508 Y.t9 GNDA 0.022794f
C509 Y.t12 GNDA 0.022794f
C510 Y.n13 GNDA 0.081534f
C511 Y.n14 GNDA 0.302737f
C512 Y.t1 GNDA 0.022794f
C513 Y.t10 GNDA 0.022794f
C514 Y.n15 GNDA 0.081534f
C515 Y.n16 GNDA 0.157046f
C516 Y.t4 GNDA 0.022794f
C517 Y.t8 GNDA 0.022794f
C518 Y.n17 GNDA 0.081534f
C519 Y.n18 GNDA 0.157046f
C520 Y.t17 GNDA 0.022794f
C521 Y.t20 GNDA 0.022794f
C522 Y.n19 GNDA 0.082252f
C523 Y.n20 GNDA 0.191279f
C524 Y.n21 GNDA 0.123631f
C525 Y.t29 GNDA 0.031912f
C526 Y.t42 GNDA 0.031912f
C527 Y.t26 GNDA 0.031912f
C528 Y.t50 GNDA 0.031912f
C529 Y.t35 GNDA 0.031912f
C530 Y.t47 GNDA 0.031912f
C531 Y.t32 GNDA 0.031912f
C532 Y.t45 GNDA 0.03875f
C533 Y.n22 GNDA 0.03875f
C534 Y.n23 GNDA 0.025074f
C535 Y.n24 GNDA 0.025074f
C536 Y.n25 GNDA 0.025074f
C537 Y.n26 GNDA 0.025074f
C538 Y.n27 GNDA 0.025074f
C539 Y.n28 GNDA 0.022459f
C540 Y.t52 GNDA 0.031912f
C541 Y.t38 GNDA 0.03875f
C542 Y.n29 GNDA 0.036135f
C543 Y.n30 GNDA 0.022101f
C544 Y.t39 GNDA 0.049008f
C545 Y.t53 GNDA 0.049008f
C546 Y.t37 GNDA 0.049008f
C547 Y.t31 GNDA 0.049008f
C548 Y.t44 GNDA 0.049008f
C549 Y.t28 GNDA 0.049008f
C550 Y.t41 GNDA 0.049008f
C551 Y.t25 GNDA 0.055713f
C552 Y.n31 GNDA 0.05028f
C553 Y.n32 GNDA 0.030772f
C554 Y.n33 GNDA 0.030772f
C555 Y.n34 GNDA 0.030772f
C556 Y.n35 GNDA 0.030772f
C557 Y.n36 GNDA 0.030772f
C558 Y.n37 GNDA 0.028157f
C559 Y.t34 GNDA 0.049008f
C560 Y.t49 GNDA 0.055713f
C561 Y.n38 GNDA 0.047665f
C562 Y.n39 GNDA 0.022031f
C563 Y.n40 GNDA 0.153015f
C564 Y.t2 GNDA 0.741299f
C565 Y.t48 GNDA 0.100295f
C566 Y.t33 GNDA 0.100295f
C567 Y.t46 GNDA 0.106821f
C568 Y.n41 GNDA 0.084651f
C569 Y.n42 GNDA 0.045253f
C570 Y.t36 GNDA 0.100295f
C571 Y.t51 GNDA 0.100295f
C572 Y.t27 GNDA 0.100295f
C573 Y.t43 GNDA 0.100295f
C574 Y.t30 GNDA 0.100295f
C575 Y.t54 GNDA 0.100295f
C576 Y.t40 GNDA 0.106821f
C577 Y.n43 GNDA 0.084651f
C578 Y.n44 GNDA 0.047868f
C579 Y.n45 GNDA 0.047868f
C580 Y.n46 GNDA 0.047868f
C581 Y.n47 GNDA 0.047868f
C582 Y.n48 GNDA 0.045253f
C583 Y.n49 GNDA 0.024415f
C584 Y.n50 GNDA 1.03694f
C585 Y.n51 GNDA 0.458663f
C586 err_amp_mir.t8 GNDA 0.020233f
C587 err_amp_mir.t1 GNDA 0.020233f
C588 err_amp_mir.t5 GNDA 0.020233f
C589 err_amp_mir.n0 GNDA 0.047731f
C590 err_amp_mir.t0 GNDA 0.020233f
C591 err_amp_mir.t4 GNDA 0.020233f
C592 err_amp_mir.n1 GNDA 0.046922f
C593 err_amp_mir.n2 GNDA 0.884615f
C594 err_amp_mir.t3 GNDA 0.020233f
C595 err_amp_mir.t2 GNDA 0.020233f
C596 err_amp_mir.n3 GNDA 0.046922f
C597 err_amp_mir.n4 GNDA 2.10658f
C598 err_amp_mir.n5 GNDA 1.98101f
C599 err_amp_mir.t13 GNDA 0.016692f
C600 err_amp_mir.t19 GNDA 0.036166f
C601 err_amp_mir.n6 GNDA 0.051623f
C602 err_amp_mir.t7 GNDA 0.016692f
C603 err_amp_mir.t18 GNDA 0.016692f
C604 err_amp_mir.t21 GNDA 0.016692f
C605 err_amp_mir.t9 GNDA 0.016692f
C606 err_amp_mir.t15 GNDA 0.016692f
C607 err_amp_mir.t20 GNDA 0.016692f
C608 err_amp_mir.t17 GNDA 0.016692f
C609 err_amp_mir.t11 GNDA 0.036166f
C610 err_amp_mir.n7 GNDA 0.056399f
C611 err_amp_mir.n8 GNDA 0.044006f
C612 err_amp_mir.n9 GNDA 0.039231f
C613 err_amp_mir.t10 GNDA 0.020233f
C614 err_amp_mir.t16 GNDA 0.020233f
C615 err_amp_mir.n10 GNDA 0.04777f
C616 err_amp_mir.t12 GNDA 0.020233f
C617 err_amp_mir.t6 GNDA 0.020233f
C618 err_amp_mir.n11 GNDA 0.061393f
C619 err_amp_mir.n12 GNDA 0.746838f
C620 err_amp_mir.n13 GNDA 0.17992f
C621 err_amp_mir.n14 GNDA 0.05811f
C622 err_amp_mir.n15 GNDA 0.039231f
C623 err_amp_mir.n16 GNDA 0.044006f
C624 err_amp_mir.n17 GNDA 0.044006f
C625 err_amp_mir.n18 GNDA 0.039231f
C626 err_amp_mir.n19 GNDA 0.05811f
C627 err_amp_mir.n20 GNDA 0.17992f
C628 err_amp_mir.n21 GNDA 0.04777f
C629 err_amp_mir.t14 GNDA 0.020233f
C630 cap_res_Y.t127 GNDA 0.345114f
C631 cap_res_Y.t25 GNDA 0.346365f
C632 cap_res_Y.t90 GNDA 0.345114f
C633 cap_res_Y.t124 GNDA 0.34782f
C634 cap_res_Y.t21 GNDA 0.378304f
C635 cap_res_Y.t101 GNDA 0.345114f
C636 cap_res_Y.t136 GNDA 0.346365f
C637 cap_res_Y.t38 GNDA 0.345114f
C638 cap_res_Y.t83 GNDA 0.346365f
C639 cap_res_Y.t67 GNDA 0.345114f
C640 cap_res_Y.t103 GNDA 0.346365f
C641 cap_res_Y.t4 GNDA 0.345114f
C642 cap_res_Y.t51 GNDA 0.346365f
C643 cap_res_Y.t105 GNDA 0.345114f
C644 cap_res_Y.t3 GNDA 0.346365f
C645 cap_res_Y.t48 GNDA 0.345114f
C646 cap_res_Y.t87 GNDA 0.346365f
C647 cap_res_Y.t7 GNDA 0.345114f
C648 cap_res_Y.t46 GNDA 0.346365f
C649 cap_res_Y.t84 GNDA 0.345114f
C650 cap_res_Y.t122 GNDA 0.346365f
C651 cap_res_Y.t106 GNDA 0.345114f
C652 cap_res_Y.t8 GNDA 0.346365f
C653 cap_res_Y.t52 GNDA 0.345114f
C654 cap_res_Y.t94 GNDA 0.346365f
C655 cap_res_Y.t12 GNDA 0.345114f
C656 cap_res_Y.t50 GNDA 0.346365f
C657 cap_res_Y.t88 GNDA 0.345114f
C658 cap_res_Y.t132 GNDA 0.346365f
C659 cap_res_Y.t55 GNDA 0.345114f
C660 cap_res_Y.t86 GNDA 0.346365f
C661 cap_res_Y.t123 GNDA 0.345114f
C662 cap_res_Y.t32 GNDA 0.346365f
C663 cap_res_Y.t92 GNDA 0.345114f
C664 cap_res_Y.t120 GNDA 0.346365f
C665 cap_res_Y.t24 GNDA 0.345114f
C666 cap_res_Y.t72 GNDA 0.346365f
C667 cap_res_Y.t60 GNDA 0.345114f
C668 cap_res_Y.t93 GNDA 0.346365f
C669 cap_res_Y.t133 GNDA 0.345114f
C670 cap_res_Y.t39 GNDA 0.346365f
C671 cap_res_Y.t98 GNDA 0.345114f
C672 cap_res_Y.t131 GNDA 0.346365f
C673 cap_res_Y.t33 GNDA 0.345114f
C674 cap_res_Y.t79 GNDA 0.346365f
C675 cap_res_Y.t135 GNDA 0.345114f
C676 cap_res_Y.t29 GNDA 0.346365f
C677 cap_res_Y.t73 GNDA 0.345114f
C678 cap_res_Y.t110 GNDA 0.346365f
C679 cap_res_Y.t102 GNDA 0.345114f
C680 cap_res_Y.t138 GNDA 0.346365f
C681 cap_res_Y.t40 GNDA 0.345114f
C682 cap_res_Y.t85 GNDA 0.346365f
C683 cap_res_Y.t1 GNDA 0.345114f
C684 cap_res_Y.t37 GNDA 0.346365f
C685 cap_res_Y.t78 GNDA 0.345114f
C686 cap_res_Y.t114 GNDA 0.346365f
C687 cap_res_Y.t34 GNDA 0.345114f
C688 cap_res_Y.t117 GNDA 0.346365f
C689 cap_res_Y.t53 GNDA 0.345114f
C690 cap_res_Y.t108 GNDA 0.346365f
C691 cap_res_Y.t11 GNDA 0.345114f
C692 cap_res_Y.t104 GNDA 0.346365f
C693 cap_res_Y.t19 GNDA 0.345114f
C694 cap_res_Y.t5 GNDA 0.362035f
C695 cap_res_Y.t126 GNDA 0.345114f
C696 cap_res_Y.t54 GNDA 0.185368f
C697 cap_res_Y.n0 GNDA 0.198389f
C698 cap_res_Y.t96 GNDA 0.345114f
C699 cap_res_Y.t100 GNDA 0.185368f
C700 cap_res_Y.n1 GNDA 0.196789f
C701 cap_res_Y.t62 GNDA 0.345114f
C702 cap_res_Y.t10 GNDA 0.185368f
C703 cap_res_Y.n2 GNDA 0.196789f
C704 cap_res_Y.t9 GNDA 0.345114f
C705 cap_res_Y.t15 GNDA 0.185368f
C706 cap_res_Y.n3 GNDA 0.196789f
C707 cap_res_Y.t107 GNDA 0.345114f
C708 cap_res_Y.t69 GNDA 0.185368f
C709 cap_res_Y.n4 GNDA 0.196789f
C710 cap_res_Y.t77 GNDA 0.345114f
C711 cap_res_Y.t112 GNDA 0.185368f
C712 cap_res_Y.n5 GNDA 0.196789f
C713 cap_res_Y.t22 GNDA 0.345114f
C714 cap_res_Y.t128 GNDA 0.185368f
C715 cap_res_Y.n6 GNDA 0.196789f
C716 cap_res_Y.t130 GNDA 0.345114f
C717 cap_res_Y.t42 GNDA 0.185368f
C718 cap_res_Y.n7 GNDA 0.196789f
C719 cap_res_Y.t36 GNDA 0.345114f
C720 cap_res_Y.t44 GNDA 0.185368f
C721 cap_res_Y.n8 GNDA 0.196789f
C722 cap_res_Y.t59 GNDA 0.345114f
C723 cap_res_Y.t91 GNDA 0.346365f
C724 cap_res_Y.t119 GNDA 0.166846f
C725 cap_res_Y.n9 GNDA 0.215207f
C726 cap_res_Y.t56 GNDA 0.18422f
C727 cap_res_Y.n10 GNDA 0.233728f
C728 cap_res_Y.t74 GNDA 0.18422f
C729 cap_res_Y.n11 GNDA 0.250999f
C730 cap_res_Y.t70 GNDA 0.18422f
C731 cap_res_Y.n12 GNDA 0.250999f
C732 cap_res_Y.t31 GNDA 0.18422f
C733 cap_res_Y.n13 GNDA 0.250999f
C734 cap_res_Y.t66 GNDA 0.18422f
C735 cap_res_Y.n14 GNDA 0.250999f
C736 cap_res_Y.t23 GNDA 0.18422f
C737 cap_res_Y.n15 GNDA 0.250999f
C738 cap_res_Y.t121 GNDA 0.18422f
C739 cap_res_Y.n16 GNDA 0.250999f
C740 cap_res_Y.t16 GNDA 0.18422f
C741 cap_res_Y.n17 GNDA 0.250999f
C742 cap_res_Y.t113 GNDA 0.18422f
C743 cap_res_Y.n18 GNDA 0.250999f
C744 cap_res_Y.t82 GNDA 0.18422f
C745 cap_res_Y.n19 GNDA 0.250999f
C746 cap_res_Y.t47 GNDA 0.18422f
C747 cap_res_Y.n20 GNDA 0.250999f
C748 cap_res_Y.t75 GNDA 0.18422f
C749 cap_res_Y.n21 GNDA 0.250999f
C750 cap_res_Y.t35 GNDA 0.18422f
C751 cap_res_Y.n22 GNDA 0.250999f
C752 cap_res_Y.t137 GNDA 0.18422f
C753 cap_res_Y.n23 GNDA 0.250999f
C754 cap_res_Y.t30 GNDA 0.18422f
C755 cap_res_Y.n24 GNDA 0.250999f
C756 cap_res_Y.t65 GNDA 0.18422f
C757 cap_res_Y.n25 GNDA 0.233728f
C758 cap_res_Y.t6 GNDA 0.343967f
C759 cap_res_Y.t49 GNDA 0.166846f
C760 cap_res_Y.n26 GNDA 0.216458f
C761 cap_res_Y.t118 GNDA 0.343967f
C762 cap_res_Y.t20 GNDA 0.166846f
C763 cap_res_Y.n27 GNDA 0.216458f
C764 cap_res_Y.t17 GNDA 0.343967f
C765 cap_res_Y.t111 GNDA 0.345114f
C766 cap_res_Y.t80 GNDA 0.363635f
C767 cap_res_Y.t41 GNDA 0.363635f
C768 cap_res_Y.t71 GNDA 0.363635f
C769 cap_res_Y.t63 GNDA 0.185368f
C770 cap_res_Y.n28 GNDA 0.216458f
C771 cap_res_Y.t27 GNDA 0.343967f
C772 cap_res_Y.t68 GNDA 0.166846f
C773 cap_res_Y.n29 GNDA 0.197936f
C774 cap_res_Y.t129 GNDA 0.343967f
C775 cap_res_Y.t28 GNDA 0.166846f
C776 cap_res_Y.n30 GNDA 0.216458f
C777 cap_res_Y.t95 GNDA 0.343967f
C778 cap_res_Y.t134 GNDA 0.166846f
C779 cap_res_Y.n31 GNDA 0.216458f
C780 cap_res_Y.t58 GNDA 0.343967f
C781 cap_res_Y.t97 GNDA 0.166846f
C782 cap_res_Y.n32 GNDA 0.216458f
C783 cap_res_Y.t76 GNDA 0.343967f
C784 cap_res_Y.t99 GNDA 0.345114f
C785 cap_res_Y.t61 GNDA 0.363635f
C786 cap_res_Y.t14 GNDA 0.363635f
C787 cap_res_Y.t57 GNDA 0.363635f
C788 cap_res_Y.t109 GNDA 0.185368f
C789 cap_res_Y.n33 GNDA 0.216458f
C790 cap_res_Y.t43 GNDA 0.343967f
C791 cap_res_Y.t64 GNDA 0.345114f
C792 cap_res_Y.t18 GNDA 0.363635f
C793 cap_res_Y.t116 GNDA 0.363635f
C794 cap_res_Y.t13 GNDA 0.363635f
C795 cap_res_Y.t81 GNDA 0.185368f
C796 cap_res_Y.n34 GNDA 0.216458f
C797 cap_res_Y.t2 GNDA 0.343967f
C798 cap_res_Y.n35 GNDA 0.216458f
C799 cap_res_Y.t45 GNDA 0.185368f
C800 cap_res_Y.t115 GNDA 0.363635f
C801 cap_res_Y.t89 GNDA 0.363635f
C802 cap_res_Y.t125 GNDA 0.363635f
C803 cap_res_Y.t26 GNDA 0.602274f
C804 cap_res_Y.t0 GNDA 0.298233f
C805 VOUT+.t12 GNDA 0.043577f
C806 VOUT+.t9 GNDA 0.043577f
C807 VOUT+.n0 GNDA 0.175148f
C808 VOUT+.t16 GNDA 0.043577f
C809 VOUT+.t5 GNDA 0.043577f
C810 VOUT+.n1 GNDA 0.174825f
C811 VOUT+.n2 GNDA 0.172223f
C812 VOUT+.t1 GNDA 0.043577f
C813 VOUT+.t17 GNDA 0.043577f
C814 VOUT+.n3 GNDA 0.174825f
C815 VOUT+.n4 GNDA 0.088815f
C816 VOUT+.t0 GNDA 0.043577f
C817 VOUT+.t8 GNDA 0.043577f
C818 VOUT+.n5 GNDA 0.174825f
C819 VOUT+.n6 GNDA 0.088815f
C820 VOUT+.t7 GNDA 0.043577f
C821 VOUT+.t13 GNDA 0.043577f
C822 VOUT+.n7 GNDA 0.175148f
C823 VOUT+.n8 GNDA 0.105197f
C824 VOUT+.t4 GNDA 0.043577f
C825 VOUT+.t11 GNDA 0.043577f
C826 VOUT+.n9 GNDA 0.172685f
C827 VOUT+.n10 GNDA 0.210763f
C828 VOUT+.t98 GNDA 0.295461f
C829 VOUT+.t66 GNDA 0.290513f
C830 VOUT+.n11 GNDA 0.194779f
C831 VOUT+.t38 GNDA 0.290513f
C832 VOUT+.n12 GNDA 0.127099f
C833 VOUT+.t146 GNDA 0.295461f
C834 VOUT+.t53 GNDA 0.290513f
C835 VOUT+.n13 GNDA 0.194779f
C836 VOUT+.t101 GNDA 0.290513f
C837 VOUT+.t121 GNDA 0.294841f
C838 VOUT+.t27 GNDA 0.294841f
C839 VOUT+.t135 GNDA 0.294841f
C840 VOUT+.t80 GNDA 0.294841f
C841 VOUT+.t50 GNDA 0.294841f
C842 VOUT+.t148 GNDA 0.294841f
C843 VOUT+.t95 GNDA 0.294841f
C844 VOUT+.t61 GNDA 0.294841f
C845 VOUT+.t31 GNDA 0.294841f
C846 VOUT+.t138 GNDA 0.294841f
C847 VOUT+.t152 GNDA 0.290513f
C848 VOUT+.n14 GNDA 0.195399f
C849 VOUT+.t103 GNDA 0.290513f
C850 VOUT+.n15 GNDA 0.24987f
C851 VOUT+.t57 GNDA 0.290513f
C852 VOUT+.n16 GNDA 0.24987f
C853 VOUT+.t147 GNDA 0.290513f
C854 VOUT+.n17 GNDA 0.24987f
C855 VOUT+.t142 GNDA 0.290513f
C856 VOUT+.n18 GNDA 0.24987f
C857 VOUT+.t88 GNDA 0.290513f
C858 VOUT+.n19 GNDA 0.24987f
C859 VOUT+.t45 GNDA 0.290513f
C860 VOUT+.n20 GNDA 0.24987f
C861 VOUT+.t29 GNDA 0.290513f
C862 VOUT+.n21 GNDA 0.24987f
C863 VOUT+.t115 GNDA 0.290513f
C864 VOUT+.n22 GNDA 0.24987f
C865 VOUT+.t113 GNDA 0.290513f
C866 VOUT+.n23 GNDA 0.24987f
C867 VOUT+.n24 GNDA 0.236042f
C868 VOUT+.t123 GNDA 0.295461f
C869 VOUT+.t40 GNDA 0.290513f
C870 VOUT+.n25 GNDA 0.194779f
C871 VOUT+.t83 GNDA 0.290513f
C872 VOUT+.t104 GNDA 0.295461f
C873 VOUT+.t49 GNDA 0.290513f
C874 VOUT+.n26 GNDA 0.194779f
C875 VOUT+.n27 GNDA 0.236042f
C876 VOUT+.t156 GNDA 0.295461f
C877 VOUT+.t120 GNDA 0.290513f
C878 VOUT+.n28 GNDA 0.194779f
C879 VOUT+.t87 GNDA 0.290513f
C880 VOUT+.t79 GNDA 0.295461f
C881 VOUT+.t43 GNDA 0.290513f
C882 VOUT+.n29 GNDA 0.194779f
C883 VOUT+.n30 GNDA 0.236042f
C884 VOUT+.t55 GNDA 0.295461f
C885 VOUT+.t19 GNDA 0.290513f
C886 VOUT+.n31 GNDA 0.194779f
C887 VOUT+.t126 GNDA 0.290513f
C888 VOUT+.t117 GNDA 0.295461f
C889 VOUT+.t72 GNDA 0.290513f
C890 VOUT+.n32 GNDA 0.194779f
C891 VOUT+.n33 GNDA 0.236042f
C892 VOUT+.t22 GNDA 0.295461f
C893 VOUT+.t128 GNDA 0.290513f
C894 VOUT+.n34 GNDA 0.194779f
C895 VOUT+.t91 GNDA 0.290513f
C896 VOUT+.t84 GNDA 0.295461f
C897 VOUT+.t47 GNDA 0.290513f
C898 VOUT+.n35 GNDA 0.194779f
C899 VOUT+.n36 GNDA 0.236042f
C900 VOUT+.t59 GNDA 0.295461f
C901 VOUT+.t26 GNDA 0.290513f
C902 VOUT+.n37 GNDA 0.194779f
C903 VOUT+.t134 GNDA 0.290513f
C904 VOUT+.t124 GNDA 0.295337f
C905 VOUT+.t78 GNDA 0.290513f
C906 VOUT+.n38 GNDA 0.193087f
C907 VOUT+.n39 GNDA 0.236042f
C908 VOUT+.t67 GNDA 0.295461f
C909 VOUT+.t33 GNDA 0.290513f
C910 VOUT+.n40 GNDA 0.194779f
C911 VOUT+.t136 GNDA 0.290513f
C912 VOUT+.n41 GNDA 0.127099f
C913 VOUT+.t30 GNDA 0.295461f
C914 VOUT+.t132 GNDA 0.290513f
C915 VOUT+.n42 GNDA 0.194779f
C916 VOUT+.t92 GNDA 0.290513f
C917 VOUT+.t151 GNDA 0.294841f
C918 VOUT+.t39 GNDA 0.294841f
C919 VOUT+.t46 GNDA 0.295461f
C920 VOUT+.t77 GNDA 0.290513f
C921 VOUT+.n43 GNDA 0.194779f
C922 VOUT+.t116 GNDA 0.290513f
C923 VOUT+.n44 GNDA 0.127099f
C924 VOUT+.t86 GNDA 0.290513f
C925 VOUT+.n45 GNDA 0.12256f
C926 VOUT+.t140 GNDA 0.294841f
C927 VOUT+.t131 GNDA 0.295461f
C928 VOUT+.t32 GNDA 0.290513f
C929 VOUT+.n46 GNDA 0.194779f
C930 VOUT+.t68 GNDA 0.290513f
C931 VOUT+.n47 GNDA 0.127099f
C932 VOUT+.t42 GNDA 0.290513f
C933 VOUT+.n48 GNDA 0.12256f
C934 VOUT+.t155 GNDA 0.294841f
C935 VOUT+.t93 GNDA 0.295461f
C936 VOUT+.t139 GNDA 0.290513f
C937 VOUT+.n49 GNDA 0.194779f
C938 VOUT+.t41 GNDA 0.290513f
C939 VOUT+.n50 GNDA 0.127099f
C940 VOUT+.t144 GNDA 0.290513f
C941 VOUT+.n51 GNDA 0.12256f
C942 VOUT+.t114 GNDA 0.294841f
C943 VOUT+.t58 GNDA 0.295461f
C944 VOUT+.t96 GNDA 0.290513f
C945 VOUT+.n52 GNDA 0.194779f
C946 VOUT+.t143 GNDA 0.290513f
C947 VOUT+.n53 GNDA 0.127099f
C948 VOUT+.t100 GNDA 0.290513f
C949 VOUT+.n54 GNDA 0.12256f
C950 VOUT+.t81 GNDA 0.294841f
C951 VOUT+.t99 GNDA 0.294841f
C952 VOUT+.t62 GNDA 0.294841f
C953 VOUT+.t28 GNDA 0.294841f
C954 VOUT+.t130 GNDA 0.294841f
C955 VOUT+.t89 GNDA 0.290513f
C956 VOUT+.n55 GNDA 0.195399f
C957 VOUT+.t129 GNDA 0.290513f
C958 VOUT+.n56 GNDA 0.24987f
C959 VOUT+.t23 GNDA 0.290513f
C960 VOUT+.n57 GNDA 0.24987f
C961 VOUT+.t60 GNDA 0.290513f
C962 VOUT+.n58 GNDA 0.24987f
C963 VOUT+.t48 GNDA 0.290513f
C964 VOUT+.n59 GNDA 0.30888f
C965 VOUT+.t76 GNDA 0.290513f
C966 VOUT+.n60 GNDA 0.30888f
C967 VOUT+.t112 GNDA 0.290513f
C968 VOUT+.n61 GNDA 0.30888f
C969 VOUT+.t94 GNDA 0.290513f
C970 VOUT+.n62 GNDA 0.30888f
C971 VOUT+.t137 GNDA 0.290513f
C972 VOUT+.n63 GNDA 0.24987f
C973 VOUT+.t108 GNDA 0.290513f
C974 VOUT+.n64 GNDA 0.24987f
C975 VOUT+.n65 GNDA 0.236042f
C976 VOUT+.t56 GNDA 0.295461f
C977 VOUT+.t21 GNDA 0.290513f
C978 VOUT+.n66 GNDA 0.194779f
C979 VOUT+.t127 GNDA 0.290513f
C980 VOUT+.t119 GNDA 0.295461f
C981 VOUT+.t74 GNDA 0.290513f
C982 VOUT+.n67 GNDA 0.194779f
C983 VOUT+.n68 GNDA 0.236042f
C984 VOUT+.t90 GNDA 0.295461f
C985 VOUT+.t54 GNDA 0.290513f
C986 VOUT+.n69 GNDA 0.194779f
C987 VOUT+.t20 GNDA 0.290513f
C988 VOUT+.t153 GNDA 0.295461f
C989 VOUT+.t106 GNDA 0.290513f
C990 VOUT+.n70 GNDA 0.194779f
C991 VOUT+.n71 GNDA 0.236042f
C992 VOUT+.t52 GNDA 0.295461f
C993 VOUT+.t154 GNDA 0.290513f
C994 VOUT+.n72 GNDA 0.194779f
C995 VOUT+.t122 GNDA 0.290513f
C996 VOUT+.t109 GNDA 0.295461f
C997 VOUT+.t70 GNDA 0.290513f
C998 VOUT+.n73 GNDA 0.194779f
C999 VOUT+.n74 GNDA 0.236042f
C1000 VOUT+.t150 GNDA 0.295461f
C1001 VOUT+.t111 GNDA 0.290513f
C1002 VOUT+.n75 GNDA 0.194779f
C1003 VOUT+.t82 GNDA 0.290513f
C1004 VOUT+.t73 GNDA 0.295461f
C1005 VOUT+.t35 GNDA 0.290513f
C1006 VOUT+.n76 GNDA 0.194779f
C1007 VOUT+.n77 GNDA 0.236042f
C1008 VOUT+.t51 GNDA 0.295461f
C1009 VOUT+.t149 GNDA 0.290513f
C1010 VOUT+.n78 GNDA 0.194779f
C1011 VOUT+.t110 GNDA 0.290513f
C1012 VOUT+.t105 GNDA 0.295461f
C1013 VOUT+.t63 GNDA 0.290513f
C1014 VOUT+.n79 GNDA 0.194779f
C1015 VOUT+.n80 GNDA 0.236042f
C1016 VOUT+.t145 GNDA 0.295461f
C1017 VOUT+.t107 GNDA 0.290513f
C1018 VOUT+.n81 GNDA 0.194779f
C1019 VOUT+.t75 GNDA 0.290513f
C1020 VOUT+.t69 GNDA 0.295461f
C1021 VOUT+.t25 GNDA 0.290513f
C1022 VOUT+.n82 GNDA 0.194779f
C1023 VOUT+.n83 GNDA 0.236042f
C1024 VOUT+.t102 GNDA 0.295461f
C1025 VOUT+.t71 GNDA 0.290513f
C1026 VOUT+.n84 GNDA 0.194779f
C1027 VOUT+.t44 GNDA 0.290513f
C1028 VOUT+.t34 GNDA 0.295461f
C1029 VOUT+.t125 GNDA 0.290513f
C1030 VOUT+.n85 GNDA 0.194779f
C1031 VOUT+.n86 GNDA 0.236042f
C1032 VOUT+.t65 GNDA 0.295461f
C1033 VOUT+.t37 GNDA 0.290513f
C1034 VOUT+.n87 GNDA 0.194779f
C1035 VOUT+.t141 GNDA 0.290513f
C1036 VOUT+.t133 GNDA 0.295461f
C1037 VOUT+.t85 GNDA 0.290513f
C1038 VOUT+.n88 GNDA 0.194779f
C1039 VOUT+.n89 GNDA 0.236042f
C1040 VOUT+.t97 GNDA 0.295461f
C1041 VOUT+.t64 GNDA 0.290513f
C1042 VOUT+.n90 GNDA 0.194779f
C1043 VOUT+.t36 GNDA 0.290513f
C1044 VOUT+.n91 GNDA 0.236042f
C1045 VOUT+.t118 GNDA 0.290513f
C1046 VOUT+.n92 GNDA 0.127099f
C1047 VOUT+.t24 GNDA 0.290513f
C1048 VOUT+.n93 GNDA 0.238016f
C1049 VOUT+.n94 GNDA 0.268648f
C1050 VOUT+.t3 GNDA 0.05084f
C1051 VOUT+.t14 GNDA 0.05084f
C1052 VOUT+.n95 GNDA 0.235187f
C1053 VOUT+.t6 GNDA 0.05084f
C1054 VOUT+.t2 GNDA 0.05084f
C1055 VOUT+.n96 GNDA 0.2344f
C1056 VOUT+.n97 GNDA 0.144847f
C1057 VOUT+.t15 GNDA 0.05084f
C1058 VOUT+.t10 GNDA 0.05084f
C1059 VOUT+.n98 GNDA 0.2344f
C1060 VOUT+.n99 GNDA 0.089159f
C1061 VOUT+.t18 GNDA 0.084056f
C1062 VOUT+.n100 GNDA 0.119121f
C1063 X.t14 GNDA 0.052601f
C1064 X.t4 GNDA 0.052601f
C1065 X.n0 GNDA 0.182935f
C1066 X.t19 GNDA 0.052601f
C1067 X.t3 GNDA 0.052601f
C1068 X.n1 GNDA 0.182287f
C1069 X.n2 GNDA 0.344139f
C1070 X.t9 GNDA 0.052601f
C1071 X.t18 GNDA 0.052601f
C1072 X.n3 GNDA 0.182287f
C1073 X.n4 GNDA 0.178405f
C1074 X.t11 GNDA 0.052601f
C1075 X.t2 GNDA 0.052601f
C1076 X.n5 GNDA 0.182287f
C1077 X.n6 GNDA 0.178405f
C1078 X.t16 GNDA 0.052601f
C1079 X.t22 GNDA 0.052601f
C1080 X.n7 GNDA 0.182287f
C1081 X.n8 GNDA 0.210076f
C1082 X.t17 GNDA 0.052601f
C1083 X.t12 GNDA 0.052601f
C1084 X.n9 GNDA 0.178511f
C1085 X.n10 GNDA 0.147505f
C1086 X.t13 GNDA 0.022543f
C1087 X.t10 GNDA 0.022543f
C1088 X.n11 GNDA 0.076111f
C1089 X.t20 GNDA 0.022543f
C1090 X.t8 GNDA 0.022543f
C1091 X.n12 GNDA 0.081346f
C1092 X.t7 GNDA 0.022543f
C1093 X.t21 GNDA 0.022543f
C1094 X.n13 GNDA 0.081346f
C1095 X.t0 GNDA 0.022543f
C1096 X.t5 GNDA 0.022543f
C1097 X.n14 GNDA 0.080636f
C1098 X.n15 GNDA 0.299403f
C1099 X.t15 GNDA 0.022543f
C1100 X.t6 GNDA 0.022543f
C1101 X.n16 GNDA 0.080636f
C1102 X.n17 GNDA 0.155317f
C1103 X.t24 GNDA 0.022543f
C1104 X.t23 GNDA 0.022543f
C1105 X.n18 GNDA 0.080636f
C1106 X.n19 GNDA 0.155317f
C1107 X.n20 GNDA 0.189173f
C1108 X.n21 GNDA 0.122269f
C1109 X.n22 GNDA 0.128676f
C1110 X.t47 GNDA 0.03156f
C1111 X.t42 GNDA 0.038324f
C1112 X.n23 GNDA 0.035737f
C1113 X.t33 GNDA 0.03156f
C1114 X.t50 GNDA 0.03156f
C1115 X.t36 GNDA 0.03156f
C1116 X.t54 GNDA 0.03156f
C1117 X.t39 GNDA 0.03156f
C1118 X.t26 GNDA 0.03156f
C1119 X.t41 GNDA 0.03156f
C1120 X.t28 GNDA 0.038324f
C1121 X.n24 GNDA 0.038324f
C1122 X.n25 GNDA 0.024798f
C1123 X.n26 GNDA 0.024798f
C1124 X.n27 GNDA 0.024798f
C1125 X.n28 GNDA 0.024798f
C1126 X.n29 GNDA 0.024798f
C1127 X.n30 GNDA 0.022211f
C1128 X.n31 GNDA 0.021857f
C1129 X.t29 GNDA 0.048468f
C1130 X.t53 GNDA 0.0551f
C1131 X.n32 GNDA 0.04714f
C1132 X.t45 GNDA 0.048468f
C1133 X.t31 GNDA 0.048468f
C1134 X.t46 GNDA 0.048468f
C1135 X.t32 GNDA 0.048468f
C1136 X.t49 GNDA 0.048468f
C1137 X.t35 GNDA 0.048468f
C1138 X.t52 GNDA 0.048468f
C1139 X.t38 GNDA 0.0551f
C1140 X.n33 GNDA 0.049726f
C1141 X.n34 GNDA 0.030433f
C1142 X.n35 GNDA 0.030433f
C1143 X.n36 GNDA 0.030433f
C1144 X.n37 GNDA 0.030433f
C1145 X.n38 GNDA 0.030433f
C1146 X.n39 GNDA 0.027847f
C1147 X.n40 GNDA 0.021789f
C1148 X.n41 GNDA 0.153028f
C1149 X.n42 GNDA 0.454714f
C1150 X.t40 GNDA 0.09919f
C1151 X.t25 GNDA 0.09919f
C1152 X.t37 GNDA 0.09919f
C1153 X.t51 GNDA 0.09919f
C1154 X.t34 GNDA 0.09919f
C1155 X.t48 GNDA 0.09919f
C1156 X.t44 GNDA 0.105644f
C1157 X.n43 GNDA 0.083719f
C1158 X.n44 GNDA 0.047341f
C1159 X.n45 GNDA 0.047341f
C1160 X.n46 GNDA 0.047341f
C1161 X.n47 GNDA 0.047341f
C1162 X.n48 GNDA 0.044755f
C1163 X.t27 GNDA 0.09919f
C1164 X.t43 GNDA 0.09919f
C1165 X.t30 GNDA 0.105644f
C1166 X.n49 GNDA 0.083719f
C1167 X.n50 GNDA 0.044755f
C1168 X.n51 GNDA 0.024251f
C1169 X.n52 GNDA 1.03308f
C1170 X.t1 GNDA 0.734227f
C1171 VD4.n0 GNDA 0.050227f
C1172 VD4.t28 GNDA 0.024416f
C1173 VD4.t11 GNDA 0.024416f
C1174 VD4.n1 GNDA 0.079606f
C1175 VD4.t1 GNDA 0.024416f
C1176 VD4.t9 GNDA 0.024416f
C1177 VD4.n2 GNDA 0.084727f
C1178 VD4.t24 GNDA 0.024416f
C1179 VD4.t13 GNDA 0.024416f
C1180 VD4.n3 GNDA 0.084913f
C1181 VD4.t12 GNDA 0.024416f
C1182 VD4.t25 GNDA 0.024416f
C1183 VD4.n4 GNDA 0.084913f
C1184 VD4.t26 GNDA 0.024416f
C1185 VD4.t7 GNDA 0.024416f
C1186 VD4.n5 GNDA 0.084613f
C1187 VD4.n6 GNDA 0.15974f
C1188 VD4.t29 GNDA 0.024416f
C1189 VD4.t30 GNDA 0.024416f
C1190 VD4.n7 GNDA 0.084613f
C1191 VD4.n8 GNDA 0.082811f
C1192 VD4.t21 GNDA 0.024416f
C1193 VD4.t2 GNDA 0.024416f
C1194 VD4.n9 GNDA 0.084613f
C1195 VD4.n10 GNDA 0.082811f
C1196 VD4.n11 GNDA 0.099252f
C1197 VD4.t14 GNDA 0.024416f
C1198 VD4.t31 GNDA 0.024416f
C1199 VD4.n12 GNDA 0.08286f
C1200 VD4.n13 GNDA 0.100481f
C1201 VD4.n14 GNDA 0.094683f
C1202 VD4.t4 GNDA 0.024416f
C1203 VD4.t6 GNDA 0.024416f
C1204 VD4.n15 GNDA 0.084612f
C1205 VD4.n16 GNDA 0.078625f
C1206 VD4.t20 GNDA 0.024416f
C1207 VD4.t18 GNDA 0.024416f
C1208 VD4.n17 GNDA 0.084913f
C1209 VD4.t16 GNDA 0.024416f
C1210 VD4.t23 GNDA 0.024416f
C1211 VD4.n18 GNDA 0.084612f
C1212 VD4.n19 GNDA 0.15974f
C1213 VD4.n20 GNDA 0.029845f
C1214 VD4.n21 GNDA 0.057972f
C1215 VD4.n22 GNDA 0.097309f
C1216 VD4.n23 GNDA 0.094519f
C1217 VD4.n24 GNDA 0.094519f
C1218 VD4.t34 GNDA 0.120449f
C1219 VD4.t32 GNDA 0.042516f
C1220 VD4.n25 GNDA 0.078578f
C1221 VD4.n26 GNDA 0.050655f
C1222 VD4.n27 GNDA 0.069509f
C1223 VD4.n28 GNDA 0.281683f
C1224 VD4.t33 GNDA 0.420453f
C1225 VD4.t0 GNDA 0.242764f
C1226 VD4.t8 GNDA 0.242764f
C1227 VD4.t3 GNDA 0.242764f
C1228 VD4.t5 GNDA 0.242764f
C1229 VD4.t27 GNDA 0.182073f
C1230 VD4.n29 GNDA 0.121382f
C1231 VD4.t10 GNDA 0.182073f
C1232 VD4.t15 GNDA 0.242764f
C1233 VD4.t22 GNDA 0.242764f
C1234 VD4.t19 GNDA 0.242764f
C1235 VD4.t17 GNDA 0.242764f
C1236 VD4.t36 GNDA 0.420453f
C1237 VD4.n30 GNDA 0.281683f
C1238 VD4.n31 GNDA 0.069509f
C1239 VD4.n32 GNDA 0.050655f
C1240 VD4.t35 GNDA 0.042516f
C1241 VD4.n33 GNDA 0.078578f
C1242 VD4.t37 GNDA 0.120449f
C1243 VDDA.t238 GNDA 0.020359f
C1244 VDDA.t223 GNDA 0.020359f
C1245 VDDA.n0 GNDA 0.084193f
C1246 VDDA.t73 GNDA 0.020359f
C1247 VDDA.t81 GNDA 0.020359f
C1248 VDDA.n1 GNDA 0.08387f
C1249 VDDA.n2 GNDA 0.116281f
C1250 VDDA.t80 GNDA 0.020359f
C1251 VDDA.t260 GNDA 0.020359f
C1252 VDDA.n3 GNDA 0.08387f
C1253 VDDA.n4 GNDA 0.060677f
C1254 VDDA.t101 GNDA 0.020359f
C1255 VDDA.t12 GNDA 0.020359f
C1256 VDDA.n5 GNDA 0.08387f
C1257 VDDA.n6 GNDA 0.060677f
C1258 VDDA.t90 GNDA 0.020359f
C1259 VDDA.t1 GNDA 0.020359f
C1260 VDDA.n7 GNDA 0.08387f
C1261 VDDA.n8 GNDA 0.060677f
C1262 VDDA.t222 GNDA 0.020359f
C1263 VDDA.t95 GNDA 0.020359f
C1264 VDDA.n9 GNDA 0.08387f
C1265 VDDA.n10 GNDA 0.175242f
C1266 VDDA.t112 GNDA 0.040718f
C1267 VDDA.t63 GNDA 0.040718f
C1268 VDDA.n11 GNDA 0.163354f
C1269 VDDA.n12 GNDA 0.082988f
C1270 VDDA.t173 GNDA 0.040562f
C1271 VDDA.n13 GNDA 0.054924f
C1272 VDDA.n14 GNDA 0.077525f
C1273 VDDA.t176 GNDA 0.045048f
C1274 VDDA.t174 GNDA 0.019727f
C1275 VDDA.n15 GNDA 0.071459f
C1276 VDDA.n16 GNDA 0.042068f
C1277 VDDA.t167 GNDA 0.045048f
C1278 VDDA.t165 GNDA 0.019727f
C1279 VDDA.n17 GNDA 0.071459f
C1280 VDDA.n18 GNDA 0.042068f
C1281 VDDA.n19 GNDA 0.044789f
C1282 VDDA.n20 GNDA 0.077525f
C1283 VDDA.n21 GNDA 0.224118f
C1284 VDDA.t166 GNDA 0.277564f
C1285 VDDA.t256 GNDA 0.160495f
C1286 VDDA.t40 GNDA 0.160495f
C1287 VDDA.t41 GNDA 0.160495f
C1288 VDDA.t21 GNDA 0.160495f
C1289 VDDA.t108 GNDA 0.120371f
C1290 VDDA.n22 GNDA 0.080247f
C1291 VDDA.t65 GNDA 0.120371f
C1292 VDDA.t27 GNDA 0.160495f
C1293 VDDA.t19 GNDA 0.160495f
C1294 VDDA.t28 GNDA 0.160495f
C1295 VDDA.t20 GNDA 0.160495f
C1296 VDDA.t175 GNDA 0.277564f
C1297 VDDA.n23 GNDA 0.224118f
C1298 VDDA.n24 GNDA 0.054924f
C1299 VDDA.n25 GNDA 0.103934f
C1300 VDDA.n26 GNDA 0.071129f
C1301 VDDA.n27 GNDA 0.105504f
C1302 VDDA.n28 GNDA 0.105504f
C1303 VDDA.n29 GNDA 0.104817f
C1304 VDDA.t161 GNDA 0.040562f
C1305 VDDA.t71 GNDA 0.040718f
C1306 VDDA.t30 GNDA 0.040718f
C1307 VDDA.n30 GNDA 0.163354f
C1308 VDDA.n31 GNDA 0.082988f
C1309 VDDA.t246 GNDA 0.040718f
C1310 VDDA.t14 GNDA 0.040718f
C1311 VDDA.n32 GNDA 0.163354f
C1312 VDDA.n33 GNDA 0.082988f
C1313 VDDA.t35 GNDA 0.040718f
C1314 VDDA.t26 GNDA 0.040718f
C1315 VDDA.n34 GNDA 0.163354f
C1316 VDDA.n35 GNDA 0.082988f
C1317 VDDA.t89 GNDA 0.040718f
C1318 VDDA.t235 GNDA 0.040718f
C1319 VDDA.n36 GNDA 0.163354f
C1320 VDDA.n37 GNDA 0.174387f
C1321 VDDA.n38 GNDA 0.131665f
C1322 VDDA.t159 GNDA 0.049215f
C1323 VDDA.n39 GNDA 0.094165f
C1324 VDDA.n40 GNDA 0.055014f
C1325 VDDA.n41 GNDA 0.082313f
C1326 VDDA.n42 GNDA 0.362312f
C1327 VDDA.t160 GNDA 0.559628f
C1328 VDDA.t88 GNDA 0.309793f
C1329 VDDA.t234 GNDA 0.309793f
C1330 VDDA.t34 GNDA 0.309793f
C1331 VDDA.t25 GNDA 0.309793f
C1332 VDDA.t245 GNDA 0.232345f
C1333 VDDA.n43 GNDA 0.154896f
C1334 VDDA.t13 GNDA 0.232345f
C1335 VDDA.t70 GNDA 0.309793f
C1336 VDDA.t29 GNDA 0.309793f
C1337 VDDA.t111 GNDA 0.309793f
C1338 VDDA.t62 GNDA 0.309793f
C1339 VDDA.t172 GNDA 0.559628f
C1340 VDDA.n44 GNDA 0.362312f
C1341 VDDA.n45 GNDA 0.082313f
C1342 VDDA.n46 GNDA 0.055014f
C1343 VDDA.t171 GNDA 0.049215f
C1344 VDDA.n47 GNDA 0.094165f
C1345 VDDA.n48 GNDA 0.131325f
C1346 VDDA.n49 GNDA 0.098525f
C1347 VDDA.t220 GNDA 0.020359f
C1348 VDDA.t109 GNDA 0.020359f
C1349 VDDA.n50 GNDA 0.084193f
C1350 VDDA.t110 GNDA 0.020359f
C1351 VDDA.t39 GNDA 0.020359f
C1352 VDDA.n51 GNDA 0.08387f
C1353 VDDA.n52 GNDA 0.116281f
C1354 VDDA.t33 GNDA 0.020359f
C1355 VDDA.t18 GNDA 0.020359f
C1356 VDDA.n53 GNDA 0.08387f
C1357 VDDA.n54 GNDA 0.060677f
C1358 VDDA.t42 GNDA 0.020359f
C1359 VDDA.t15 GNDA 0.020359f
C1360 VDDA.n55 GNDA 0.08387f
C1361 VDDA.n56 GNDA 0.060677f
C1362 VDDA.t64 GNDA 0.020359f
C1363 VDDA.t98 GNDA 0.020359f
C1364 VDDA.n57 GNDA 0.08387f
C1365 VDDA.n58 GNDA 0.060677f
C1366 VDDA.t259 GNDA 0.020359f
C1367 VDDA.t221 GNDA 0.020359f
C1368 VDDA.n59 GNDA 0.08387f
C1369 VDDA.n60 GNDA 0.209634f
C1370 VDDA.n61 GNDA 0.19375f
C1371 VDDA.t59 GNDA 0.023752f
C1372 VDDA.t87 GNDA 0.023752f
C1373 VDDA.n62 GNDA 0.082604f
C1374 VDDA.t255 GNDA 0.023752f
C1375 VDDA.t107 GNDA 0.023752f
C1376 VDDA.n63 GNDA 0.082311f
C1377 VDDA.n64 GNDA 0.155396f
C1378 VDDA.t48 GNDA 0.023752f
C1379 VDDA.t55 GNDA 0.023752f
C1380 VDDA.n65 GNDA 0.082604f
C1381 VDDA.t253 GNDA 0.023752f
C1382 VDDA.t242 GNDA 0.023752f
C1383 VDDA.n66 GNDA 0.082311f
C1384 VDDA.n67 GNDA 0.155396f
C1385 VDDA.n68 GNDA 0.021716f
C1386 VDDA.n69 GNDA 0.067619f
C1387 VDDA.n70 GNDA 0.091949f
C1388 VDDA.t179 GNDA 0.117173f
C1389 VDDA.t177 GNDA 0.04136f
C1390 VDDA.n71 GNDA 0.076441f
C1391 VDDA.n72 GNDA 0.049277f
C1392 VDDA.t130 GNDA 0.117173f
C1393 VDDA.t128 GNDA 0.04136f
C1394 VDDA.n73 GNDA 0.076441f
C1395 VDDA.n74 GNDA 0.049277f
C1396 VDDA.n75 GNDA 0.048861f
C1397 VDDA.n76 GNDA 0.091949f
C1398 VDDA.n77 GNDA 0.274023f
C1399 VDDA.t129 GNDA 0.409019f
C1400 VDDA.t58 GNDA 0.236162f
C1401 VDDA.t86 GNDA 0.236162f
C1402 VDDA.t254 GNDA 0.236162f
C1403 VDDA.t106 GNDA 0.236162f
C1404 VDDA.t16 GNDA 0.177121f
C1405 VDDA.n78 GNDA 0.118081f
C1406 VDDA.t250 GNDA 0.177121f
C1407 VDDA.t252 GNDA 0.236162f
C1408 VDDA.t241 GNDA 0.236162f
C1409 VDDA.t47 GNDA 0.236162f
C1410 VDDA.t54 GNDA 0.236162f
C1411 VDDA.t178 GNDA 0.409019f
C1412 VDDA.n79 GNDA 0.274023f
C1413 VDDA.n80 GNDA 0.067619f
C1414 VDDA.n81 GNDA 0.094663f
C1415 VDDA.t17 GNDA 0.023752f
C1416 VDDA.t251 GNDA 0.023752f
C1417 VDDA.n82 GNDA 0.077441f
C1418 VDDA.n83 GNDA 0.052855f
C1419 VDDA.n84 GNDA 0.029483f
C1420 VDDA.n85 GNDA 0.118458f
C1421 VDDA.t24 GNDA 0.023752f
C1422 VDDA.t248 GNDA 0.023752f
C1423 VDDA.n86 GNDA 0.082604f
C1424 VDDA.t44 GNDA 0.023752f
C1425 VDDA.t100 GNDA 0.023752f
C1426 VDDA.n87 GNDA 0.082311f
C1427 VDDA.n88 GNDA 0.155396f
C1428 VDDA.t52 GNDA 0.023752f
C1429 VDDA.t85 GNDA 0.023752f
C1430 VDDA.n89 GNDA 0.082604f
C1431 VDDA.t32 GNDA 0.023752f
C1432 VDDA.t244 GNDA 0.023752f
C1433 VDDA.n90 GNDA 0.082311f
C1434 VDDA.n91 GNDA 0.155396f
C1435 VDDA.n92 GNDA 0.021716f
C1436 VDDA.n93 GNDA 0.067619f
C1437 VDDA.n94 GNDA 0.091949f
C1438 VDDA.t155 GNDA 0.117173f
C1439 VDDA.t153 GNDA 0.04136f
C1440 VDDA.n95 GNDA 0.076441f
C1441 VDDA.n96 GNDA 0.049277f
C1442 VDDA.t133 GNDA 0.117173f
C1443 VDDA.t131 GNDA 0.04136f
C1444 VDDA.n97 GNDA 0.076441f
C1445 VDDA.n98 GNDA 0.049277f
C1446 VDDA.n99 GNDA 0.048861f
C1447 VDDA.n100 GNDA 0.091949f
C1448 VDDA.n101 GNDA 0.274023f
C1449 VDDA.t132 GNDA 0.409019f
C1450 VDDA.t23 GNDA 0.236162f
C1451 VDDA.t247 GNDA 0.236162f
C1452 VDDA.t43 GNDA 0.236162f
C1453 VDDA.t99 GNDA 0.236162f
C1454 VDDA.t7 GNDA 0.177121f
C1455 VDDA.n102 GNDA 0.118081f
C1456 VDDA.t82 GNDA 0.177121f
C1457 VDDA.t31 GNDA 0.236162f
C1458 VDDA.t243 GNDA 0.236162f
C1459 VDDA.t51 GNDA 0.236162f
C1460 VDDA.t84 GNDA 0.236162f
C1461 VDDA.t154 GNDA 0.409019f
C1462 VDDA.n103 GNDA 0.274023f
C1463 VDDA.n104 GNDA 0.067619f
C1464 VDDA.n105 GNDA 0.094663f
C1465 VDDA.t8 GNDA 0.023752f
C1466 VDDA.t83 GNDA 0.023752f
C1467 VDDA.n106 GNDA 0.077441f
C1468 VDDA.n107 GNDA 0.052855f
C1469 VDDA.n108 GNDA 0.029483f
C1470 VDDA.n109 GNDA 0.116422f
C1471 VDDA.t57 GNDA 0.040718f
C1472 VDDA.t3 GNDA 0.040718f
C1473 VDDA.n110 GNDA 0.163354f
C1474 VDDA.n111 GNDA 0.082988f
C1475 VDDA.t115 GNDA 0.040562f
C1476 VDDA.n112 GNDA 0.082313f
C1477 VDDA.n113 GNDA 0.054924f
C1478 VDDA.n114 GNDA 0.077525f
C1479 VDDA.t127 GNDA 0.045048f
C1480 VDDA.t125 GNDA 0.019727f
C1481 VDDA.n115 GNDA 0.071459f
C1482 VDDA.n116 GNDA 0.042068f
C1483 VDDA.t118 GNDA 0.045048f
C1484 VDDA.t116 GNDA 0.019727f
C1485 VDDA.n117 GNDA 0.071459f
C1486 VDDA.n118 GNDA 0.042068f
C1487 VDDA.n119 GNDA 0.044789f
C1488 VDDA.n120 GNDA 0.077525f
C1489 VDDA.n121 GNDA 0.224118f
C1490 VDDA.t117 GNDA 0.277564f
C1491 VDDA.t74 GNDA 0.160495f
C1492 VDDA.t4 GNDA 0.160495f
C1493 VDDA.t77 GNDA 0.160495f
C1494 VDDA.t236 GNDA 0.160495f
C1495 VDDA.t22 GNDA 0.120371f
C1496 VDDA.n122 GNDA 0.080247f
C1497 VDDA.t11 GNDA 0.120371f
C1498 VDDA.t239 GNDA 0.160495f
C1499 VDDA.t237 GNDA 0.160495f
C1500 VDDA.t0 GNDA 0.160495f
C1501 VDDA.t240 GNDA 0.160495f
C1502 VDDA.t126 GNDA 0.277564f
C1503 VDDA.n123 GNDA 0.224118f
C1504 VDDA.n124 GNDA 0.054924f
C1505 VDDA.n125 GNDA 0.103934f
C1506 VDDA.t121 GNDA 0.040562f
C1507 VDDA.t94 GNDA 0.040718f
C1508 VDDA.t10 GNDA 0.040718f
C1509 VDDA.n126 GNDA 0.163354f
C1510 VDDA.n127 GNDA 0.082988f
C1511 VDDA.t6 GNDA 0.040718f
C1512 VDDA.t76 GNDA 0.040718f
C1513 VDDA.n128 GNDA 0.163354f
C1514 VDDA.n129 GNDA 0.082988f
C1515 VDDA.t79 GNDA 0.040718f
C1516 VDDA.t46 GNDA 0.040718f
C1517 VDDA.n130 GNDA 0.163354f
C1518 VDDA.n131 GNDA 0.082988f
C1519 VDDA.t258 GNDA 0.040718f
C1520 VDDA.t97 GNDA 0.040718f
C1521 VDDA.n132 GNDA 0.163354f
C1522 VDDA.n133 GNDA 0.174387f
C1523 VDDA.n134 GNDA 0.131665f
C1524 VDDA.t119 GNDA 0.049215f
C1525 VDDA.n135 GNDA 0.094165f
C1526 VDDA.n136 GNDA 0.055014f
C1527 VDDA.n137 GNDA 0.362312f
C1528 VDDA.n138 GNDA 0.362312f
C1529 VDDA.t114 GNDA 0.559628f
C1530 VDDA.t56 GNDA 0.309793f
C1531 VDDA.t2 GNDA 0.309793f
C1532 VDDA.t93 GNDA 0.309793f
C1533 VDDA.t9 GNDA 0.309793f
C1534 VDDA.t5 GNDA 0.232345f
C1535 VDDA.n139 GNDA 0.082313f
C1536 VDDA.n140 GNDA 0.105504f
C1537 VDDA.n141 GNDA 0.105504f
C1538 VDDA.t120 GNDA 0.559628f
C1539 VDDA.t96 GNDA 0.309793f
C1540 VDDA.t257 GNDA 0.309793f
C1541 VDDA.t45 GNDA 0.309793f
C1542 VDDA.t78 GNDA 0.309793f
C1543 VDDA.t75 GNDA 0.232345f
C1544 VDDA.n142 GNDA 0.154896f
C1545 VDDA.n143 GNDA 0.104817f
C1546 VDDA.n144 GNDA 0.071129f
C1547 VDDA.n145 GNDA 0.055014f
C1548 VDDA.t113 GNDA 0.049215f
C1549 VDDA.n146 GNDA 0.094165f
C1550 VDDA.n147 GNDA 0.131325f
C1551 VDDA.n148 GNDA 0.100561f
C1552 VDDA.n149 GNDA 0.056326f
C1553 VDDA.n150 GNDA 0.190477f
C1554 VDDA.n151 GNDA 0.065742f
C1555 VDDA.n152 GNDA 0.175511f
C1556 VDDA.t145 GNDA 0.012787f
C1557 VDDA.n153 GNDA 0.027208f
C1558 VDDA.t139 GNDA 0.012787f
C1559 VDDA.n154 GNDA 0.027208f
C1560 VDDA.n155 GNDA 0.039506f
C1561 VDDA.n156 GNDA 0.066401f
C1562 VDDA.n157 GNDA 0.17696f
C1563 VDDA.t158 GNDA 0.012787f
C1564 VDDA.n158 GNDA 0.027208f
C1565 VDDA.t152 GNDA 0.012787f
C1566 VDDA.n159 GNDA 0.027208f
C1567 VDDA.n160 GNDA 0.036815f
C1568 VDDA.n161 GNDA 0.0457f
C1569 VDDA.n162 GNDA 0.17696f
C1570 VDDA.t151 GNDA 0.172148f
C1571 VDDA.t224 GNDA 0.106375f
C1572 VDDA.t68 GNDA 0.106375f
C1573 VDDA.t53 GNDA 0.106375f
C1574 VDDA.t230 GNDA 0.106375f
C1575 VDDA.t226 GNDA 0.079781f
C1576 VDDA.t157 GNDA 0.172148f
C1577 VDDA.t50 GNDA 0.106375f
C1578 VDDA.t231 GNDA 0.106375f
C1579 VDDA.t227 GNDA 0.106375f
C1580 VDDA.t69 GNDA 0.106375f
C1581 VDDA.t49 GNDA 0.079781f
C1582 VDDA.n163 GNDA 0.067059f
C1583 VDDA.n164 GNDA 0.053187f
C1584 VDDA.n165 GNDA 0.067059f
C1585 VDDA.n166 GNDA 0.044789f
C1586 VDDA.n167 GNDA 0.036239f
C1587 VDDA.n168 GNDA 0.08426f
C1588 VDDA.n169 GNDA 0.08426f
C1589 VDDA.n170 GNDA 0.175511f
C1590 VDDA.t138 GNDA 0.168677f
C1591 VDDA.t233 GNDA 0.104508f
C1592 VDDA.t38 GNDA 0.104508f
C1593 VDDA.t104 GNDA 0.104508f
C1594 VDDA.t228 GNDA 0.104508f
C1595 VDDA.t232 GNDA 0.078381f
C1596 VDDA.t144 GNDA 0.168677f
C1597 VDDA.t249 GNDA 0.104508f
C1598 VDDA.t229 GNDA 0.104508f
C1599 VDDA.t225 GNDA 0.104508f
C1600 VDDA.t105 GNDA 0.104508f
C1601 VDDA.t72 GNDA 0.078381f
C1602 VDDA.n171 GNDA 0.067059f
C1603 VDDA.n172 GNDA 0.052254f
C1604 VDDA.n173 GNDA 0.067059f
C1605 VDDA.n174 GNDA 0.044576f
C1606 VDDA.n175 GNDA 0.036239f
C1607 VDDA.n176 GNDA 0.070155f
C1608 VDDA.n177 GNDA 0.093844f
C1609 VDDA.n179 GNDA 0.051961f
C1610 VDDA.n180 GNDA 0.082114f
C1611 VDDA.n181 GNDA 0.104185f
C1612 VDDA.n182 GNDA 0.104185f
C1613 VDDA.n183 GNDA 0.104185f
C1614 VDDA.n185 GNDA 0.051961f
C1615 VDDA.n187 GNDA 0.051961f
C1616 VDDA.n189 GNDA 0.051961f
C1617 VDDA.n191 GNDA 0.051961f
C1618 VDDA.n193 GNDA 0.051961f
C1619 VDDA.n195 GNDA 0.051961f
C1620 VDDA.n197 GNDA 0.051961f
C1621 VDDA.n199 GNDA 0.051961f
C1622 VDDA.n201 GNDA 0.085029f
C1623 VDDA.t136 GNDA 0.012364f
C1624 VDDA.n202 GNDA 0.018358f
C1625 VDDA.n203 GNDA 0.016243f
C1626 VDDA.n204 GNDA 0.055478f
C1627 VDDA.n205 GNDA 0.064462f
C1628 VDDA.n206 GNDA 0.213035f
C1629 VDDA.t135 GNDA 0.168677f
C1630 VDDA.t214 GNDA 0.104508f
C1631 VDDA.t192 GNDA 0.104508f
C1632 VDDA.t208 GNDA 0.104508f
C1633 VDDA.t182 GNDA 0.104508f
C1634 VDDA.t196 GNDA 0.104508f
C1635 VDDA.t216 GNDA 0.104508f
C1636 VDDA.t194 GNDA 0.104508f
C1637 VDDA.t210 GNDA 0.104508f
C1638 VDDA.t206 GNDA 0.104508f
C1639 VDDA.t186 GNDA 0.078381f
C1640 VDDA.n207 GNDA 0.052254f
C1641 VDDA.t200 GNDA 0.078381f
C1642 VDDA.t180 GNDA 0.104508f
C1643 VDDA.t198 GNDA 0.104508f
C1644 VDDA.t218 GNDA 0.104508f
C1645 VDDA.t188 GNDA 0.104508f
C1646 VDDA.t204 GNDA 0.104508f
C1647 VDDA.t184 GNDA 0.104508f
C1648 VDDA.t212 GNDA 0.104508f
C1649 VDDA.t190 GNDA 0.104508f
C1650 VDDA.t202 GNDA 0.104508f
C1651 VDDA.t123 GNDA 0.168677f
C1652 VDDA.n208 GNDA 0.213035f
C1653 VDDA.n209 GNDA 0.064462f
C1654 VDDA.n210 GNDA 0.055478f
C1655 VDDA.n211 GNDA 0.016243f
C1656 VDDA.t124 GNDA 0.012364f
C1657 VDDA.n212 GNDA 0.01791f
C1658 VDDA.n213 GNDA 0.089101f
C1659 VDDA.n214 GNDA 0.082855f
C1660 VDDA.n215 GNDA 0.012309f
C1661 VDDA.n216 GNDA 0.058947f
C1662 VDDA.n217 GNDA 0.024431f
C1663 VDDA.t142 GNDA 0.016419f
C1664 VDDA.t140 GNDA 0.013308f
C1665 VDDA.n218 GNDA 0.030357f
C1666 VDDA.t149 GNDA 0.016419f
C1667 VDDA.t146 GNDA 0.013036f
C1668 VDDA.n219 GNDA 0.030357f
C1669 VDDA.n220 GNDA 0.067199f
C1670 VDDA.n221 GNDA 0.067199f
C1671 VDDA.n222 GNDA 0.065099f
C1672 VDDA.t170 GNDA 0.020451f
C1673 VDDA.n223 GNDA 0.015993f
C1674 VDDA.n224 GNDA 0.012309f
C1675 VDDA.n225 GNDA 0.081529f
C1676 VDDA.n226 GNDA 0.026199f
C1677 VDDA.t168 GNDA 0.023837f
C1678 VDDA.n227 GNDA 0.019088f
C1679 VDDA.n228 GNDA 0.037465f
C1680 VDDA.n229 GNDA 0.04765f
C1681 VDDA.n230 GNDA 0.189858f
C1682 VDDA.t169 GNDA 0.201075f
C1683 VDDA.t91 GNDA 0.12826f
C1684 VDDA.t36 GNDA 0.12826f
C1685 VDDA.t66 GNDA 0.12826f
C1686 VDDA.t60 GNDA 0.122916f
C1687 VDDA.n231 GNDA 0.06413f
C1688 VDDA.t163 GNDA 0.144293f
C1689 VDDA.t141 GNDA 0.203079f
C1690 VDDA.t102 GNDA 0.12826f
C1691 VDDA.t147 GNDA 0.201075f
C1692 VDDA.n232 GNDA 0.184374f
C1693 VDDA.n233 GNDA 0.044907f
C1694 VDDA.n234 GNDA 0.027625f
C1695 VDDA.n235 GNDA 0.019961f
C1696 VDDA.n236 GNDA 0.01012f
C1697 VDDA.t162 GNDA 0.014902f
C1698 VDDA.n237 GNDA 0.019088f
C1699 VDDA.t164 GNDA 0.020451f
C1700 VDDA.n238 GNDA 0.020929f
C1701 VDDA.n239 GNDA 0.045993f
C1702 VDDA.n241 GNDA 0.10512f
C1703 VDDA.n242 GNDA 0.630924f
C1704 V_err_gate.t30 GNDA 0.012427f
C1705 V_err_gate.t20 GNDA 0.012427f
C1706 V_err_gate.t28 GNDA 0.012427f
C1707 V_err_gate.t12 GNDA 0.012427f
C1708 V_err_gate.t22 GNDA 0.012427f
C1709 V_err_gate.t31 GNDA 0.012427f
C1710 V_err_gate.t21 GNDA 0.012427f
C1711 V_err_gate.t29 GNDA 0.012427f
C1712 V_err_gate.t19 GNDA 0.012427f
C1713 V_err_gate.t16 GNDA 0.012427f
C1714 V_err_gate.t24 GNDA 0.012427f
C1715 V_err_gate.t13 GNDA 0.012427f
C1716 V_err_gate.t23 GNDA 0.012427f
C1717 V_err_gate.t27 GNDA 0.012427f
C1718 V_err_gate.t17 GNDA 0.012427f
C1719 V_err_gate.t25 GNDA 0.012427f
C1720 V_err_gate.t14 GNDA 0.026925f
C1721 V_err_gate.n0 GNDA 0.041988f
C1722 V_err_gate.n1 GNDA 0.032762f
C1723 V_err_gate.n2 GNDA 0.032762f
C1724 V_err_gate.n3 GNDA 0.032762f
C1725 V_err_gate.n4 GNDA 0.032762f
C1726 V_err_gate.n5 GNDA 0.032762f
C1727 V_err_gate.n6 GNDA 0.032762f
C1728 V_err_gate.n7 GNDA 0.032762f
C1729 V_err_gate.n8 GNDA 0.032762f
C1730 V_err_gate.n9 GNDA 0.032762f
C1731 V_err_gate.n10 GNDA 0.032762f
C1732 V_err_gate.n11 GNDA 0.032762f
C1733 V_err_gate.n12 GNDA 0.032762f
C1734 V_err_gate.n13 GNDA 0.032762f
C1735 V_err_gate.n14 GNDA 0.032762f
C1736 V_err_gate.n15 GNDA 0.028035f
C1737 V_err_gate.t15 GNDA 0.012427f
C1738 V_err_gate.t26 GNDA 0.012427f
C1739 V_err_gate.t18 GNDA 0.026925f
C1740 V_err_gate.n16 GNDA 0.041988f
C1741 V_err_gate.n17 GNDA 0.028035f
C1742 V_err_gate.n18 GNDA 0.045175f
C1743 V_err_gate.t10 GNDA 0.015063f
C1744 V_err_gate.t8 GNDA 0.015063f
C1745 V_err_gate.n19 GNDA 0.034896f
C1746 V_err_gate.t0 GNDA 0.015063f
C1747 V_err_gate.t2 GNDA 0.015063f
C1748 V_err_gate.n20 GNDA 0.034933f
C1749 V_err_gate.n21 GNDA 0.530582f
C1750 V_err_gate.t11 GNDA 0.015063f
C1751 V_err_gate.t9 GNDA 0.015063f
C1752 V_err_gate.n22 GNDA 0.03516f
C1753 V_err_gate.t4 GNDA 0.015063f
C1754 V_err_gate.t6 GNDA 0.015063f
C1755 V_err_gate.n23 GNDA 0.034933f
C1756 V_err_gate.n24 GNDA 0.558034f
C1757 V_err_gate.t1 GNDA 0.015063f
C1758 V_err_gate.t3 GNDA 0.015063f
C1759 V_err_gate.n25 GNDA 0.034933f
C1760 V_err_gate.n26 GNDA 0.290428f
C1761 V_err_gate.n27 GNDA 0.223127f
C1762 V_err_gate.t5 GNDA 0.015063f
C1763 V_err_gate.t7 GNDA 0.015063f
C1764 V_err_gate.n28 GNDA 0.030126f
C1765 V_err_gate.n29 GNDA 0.089738f
C1766 V_err_amp_ref.t9 GNDA 0.040349f
C1767 V_err_amp_ref.t3 GNDA 0.012674f
C1768 V_err_amp_ref.t7 GNDA 0.023651f
C1769 V_err_amp_ref.n0 GNDA 0.056465f
C1770 V_err_amp_ref.n1 GNDA 0.353066f
C1771 V_err_amp_ref.t6 GNDA 0.012674f
C1772 V_err_amp_ref.t2 GNDA 0.023651f
C1773 V_err_amp_ref.n2 GNDA 0.056465f
C1774 V_err_amp_ref.n3 GNDA 0.32615f
C1775 V_err_amp_ref.t0 GNDA 0.039962f
C1776 V_err_amp_ref.n4 GNDA 0.317574f
C1777 V_err_amp_ref.t5 GNDA 0.012674f
C1778 V_err_amp_ref.t1 GNDA 0.023651f
C1779 V_err_amp_ref.n5 GNDA 0.056465f
C1780 V_err_amp_ref.n6 GNDA 0.197202f
C1781 V_err_amp_ref.t8 GNDA 0.012674f
C1782 V_err_amp_ref.t4 GNDA 0.023651f
C1783 V_err_amp_ref.n7 GNDA 0.056465f
C1784 V_err_amp_ref.n8 GNDA 0.306509f
C1785 V_p.t24 GNDA 0.024781f
C1786 V_p.n0 GNDA 0.049064f
C1787 V_p.t39 GNDA 0.014869f
C1788 V_p.t36 GNDA 0.014869f
C1789 V_p.n1 GNDA 0.050516f
C1790 V_p.t1 GNDA 0.014869f
C1791 V_p.t9 GNDA 0.014869f
C1792 V_p.n2 GNDA 0.053418f
C1793 V_p.t8 GNDA 0.014869f
C1794 V_p.t0 GNDA 0.014869f
C1795 V_p.n3 GNDA 0.053005f
C1796 V_p.n4 GNDA 0.179254f
C1797 V_p.t7 GNDA 0.014869f
C1798 V_p.t6 GNDA 0.014869f
C1799 V_p.n5 GNDA 0.053005f
C1800 V_p.n6 GNDA 0.093302f
C1801 V_p.t40 GNDA 0.014869f
C1802 V_p.t2 GNDA 0.014869f
C1803 V_p.n7 GNDA 0.053005f
C1804 V_p.n8 GNDA 0.092807f
C1805 V_p.t5 GNDA 0.014869f
C1806 V_p.t16 GNDA 0.014869f
C1807 V_p.n9 GNDA 0.053395f
C1808 V_p.t13 GNDA 0.014869f
C1809 V_p.t10 GNDA 0.014869f
C1810 V_p.n10 GNDA 0.053005f
C1811 V_p.n11 GNDA 0.177493f
C1812 V_p.t3 GNDA 0.014869f
C1813 V_p.t15 GNDA 0.014869f
C1814 V_p.n12 GNDA 0.053005f
C1815 V_p.n13 GNDA 0.093302f
C1816 V_p.t14 GNDA 0.014869f
C1817 V_p.t4 GNDA 0.014869f
C1818 V_p.n14 GNDA 0.053005f
C1819 V_p.n15 GNDA 0.093302f
C1820 V_p.t12 GNDA 0.014869f
C1821 V_p.t11 GNDA 0.014869f
C1822 V_p.n16 GNDA 0.053005f
C1823 V_p.n17 GNDA 0.142369f
C1824 V_p.n18 GNDA 0.078308f
C1825 V_p.n19 GNDA 0.0836f
C1826 V_p.t29 GNDA 0.024781f
C1827 V_p.t19 GNDA 0.024781f
C1828 V_p.n20 GNDA 0.095622f
C1829 V_p.n21 GNDA 0.079333f
C1830 V_p.n22 GNDA 0.16901f
C1831 V_p.t27 GNDA 0.024781f
C1832 V_p.t18 GNDA 0.024781f
C1833 V_p.n23 GNDA 0.098392f
C1834 V_p.n24 GNDA 0.087962f
C1835 V_p.t25 GNDA 0.024781f
C1836 V_p.t22 GNDA 0.024781f
C1837 V_p.n25 GNDA 0.098392f
C1838 V_p.n26 GNDA 0.087962f
C1839 V_p.t31 GNDA 0.024781f
C1840 V_p.t20 GNDA 0.024781f
C1841 V_p.n27 GNDA 0.098392f
C1842 V_p.n28 GNDA 0.087962f
C1843 V_p.t28 GNDA 0.024781f
C1844 V_p.t33 GNDA 0.024781f
C1845 V_p.n29 GNDA 0.098392f
C1846 V_p.n30 GNDA 0.087962f
C1847 V_p.t37 GNDA 0.086517f
C1848 V_p.t23 GNDA 0.024781f
C1849 V_p.t32 GNDA 0.024781f
C1850 V_p.n31 GNDA 0.095622f
C1851 V_p.n32 GNDA 0.572198f
C1852 V_p.n33 GNDA 0.029737f
C1853 V_p.t21 GNDA 0.024781f
C1854 V_p.t30 GNDA 0.024781f
C1855 V_p.n34 GNDA 0.098392f
C1856 V_p.n35 GNDA 0.087962f
C1857 V_p.t26 GNDA 0.024781f
C1858 V_p.t17 GNDA 0.024781f
C1859 V_p.n36 GNDA 0.098392f
C1860 V_p.n37 GNDA 0.168528f
C1861 V_p.n38 GNDA 0.098849f
C1862 V_p.t34 GNDA 0.024781f
C1863 cap_res_X.t8 GNDA 0.344645f
C1864 cap_res_X.t42 GNDA 0.167175f
C1865 cap_res_X.n0 GNDA 0.198327f
C1866 cap_res_X.t39 GNDA 0.344645f
C1867 cap_res_X.t82 GNDA 0.167175f
C1868 cap_res_X.n1 GNDA 0.216884f
C1869 cap_res_X.t79 GNDA 0.344645f
C1870 cap_res_X.t123 GNDA 0.167175f
C1871 cap_res_X.n2 GNDA 0.216884f
C1872 cap_res_X.t59 GNDA 0.344645f
C1873 cap_res_X.t102 GNDA 0.167175f
C1874 cap_res_X.n3 GNDA 0.216884f
C1875 cap_res_X.t101 GNDA 0.344645f
C1876 cap_res_X.t34 GNDA 0.345795f
C1877 cap_res_X.t1 GNDA 0.364353f
C1878 cap_res_X.t103 GNDA 0.364353f
C1879 cap_res_X.t134 GNDA 0.364353f
C1880 cap_res_X.t137 GNDA 0.185733f
C1881 cap_res_X.n4 GNDA 0.216884f
C1882 cap_res_X.t75 GNDA 0.344645f
C1883 cap_res_X.t135 GNDA 0.345795f
C1884 cap_res_X.t95 GNDA 0.364353f
C1885 cap_res_X.t54 GNDA 0.364353f
C1886 cap_res_X.t89 GNDA 0.364353f
C1887 cap_res_X.t120 GNDA 0.185733f
C1888 cap_res_X.n5 GNDA 0.216884f
C1889 cap_res_X.t126 GNDA 0.345795f
C1890 cap_res_X.t84 GNDA 0.347048f
C1891 cap_res_X.t83 GNDA 0.345795f
C1892 cap_res_X.t44 GNDA 0.348506f
C1893 cap_res_X.t14 GNDA 0.37905f
C1894 cap_res_X.t68 GNDA 0.345795f
C1895 cap_res_X.t107 GNDA 0.347048f
C1896 cap_res_X.t87 GNDA 0.345795f
C1897 cap_res_X.t48 GNDA 0.347048f
C1898 cap_res_X.t32 GNDA 0.345795f
C1899 cap_res_X.t70 GNDA 0.347048f
C1900 cap_res_X.t51 GNDA 0.345795f
C1901 cap_res_X.t20 GNDA 0.347048f
C1902 cap_res_X.t72 GNDA 0.345795f
C1903 cap_res_X.t116 GNDA 0.347048f
C1904 cap_res_X.t92 GNDA 0.345795f
C1905 cap_res_X.t58 GNDA 0.347048f
C1906 cap_res_X.t118 GNDA 0.345795f
C1907 cap_res_X.t15 GNDA 0.347048f
C1908 cap_res_X.t130 GNDA 0.345795f
C1909 cap_res_X.t99 GNDA 0.347048f
C1910 cap_res_X.t78 GNDA 0.345795f
C1911 cap_res_X.t119 GNDA 0.347048f
C1912 cap_res_X.t100 GNDA 0.345795f
C1913 cap_res_X.t64 GNDA 0.347048f
C1914 cap_res_X.t122 GNDA 0.345795f
C1915 cap_res_X.t17 GNDA 0.347048f
C1916 cap_res_X.t136 GNDA 0.345795f
C1917 cap_res_X.t105 GNDA 0.347048f
C1918 cap_res_X.t22 GNDA 0.345795f
C1919 cap_res_X.t55 GNDA 0.347048f
C1920 cap_res_X.t33 GNDA 0.345795f
C1921 cap_res_X.t5 GNDA 0.347048f
C1922 cap_res_X.t61 GNDA 0.345795f
C1923 cap_res_X.t97 GNDA 0.347048f
C1924 cap_res_X.t73 GNDA 0.345795f
C1925 cap_res_X.t37 GNDA 0.347048f
C1926 cap_res_X.t25 GNDA 0.345795f
C1927 cap_res_X.t62 GNDA 0.347048f
C1928 cap_res_X.t38 GNDA 0.345795f
C1929 cap_res_X.t13 GNDA 0.347048f
C1930 cap_res_X.t65 GNDA 0.345795f
C1931 cap_res_X.t104 GNDA 0.347048f
C1932 cap_res_X.t80 GNDA 0.345795f
C1933 cap_res_X.t45 GNDA 0.347048f
C1934 cap_res_X.t106 GNDA 0.345795f
C1935 cap_res_X.t4 GNDA 0.347048f
C1936 cap_res_X.t124 GNDA 0.345795f
C1937 cap_res_X.t86 GNDA 0.347048f
C1938 cap_res_X.t69 GNDA 0.345795f
C1939 cap_res_X.t109 GNDA 0.347048f
C1940 cap_res_X.t85 GNDA 0.345795f
C1941 cap_res_X.t49 GNDA 0.347048f
C1942 cap_res_X.t115 GNDA 0.345795f
C1943 cap_res_X.t11 GNDA 0.347048f
C1944 cap_res_X.t127 GNDA 0.345795f
C1945 cap_res_X.t91 GNDA 0.347048f
C1946 cap_res_X.t52 GNDA 0.345795f
C1947 cap_res_X.t6 GNDA 0.347048f
C1948 cap_res_X.t81 GNDA 0.345795f
C1949 cap_res_X.t132 GNDA 0.347048f
C1950 cap_res_X.t71 GNDA 0.345795f
C1951 cap_res_X.t128 GNDA 0.362749f
C1952 cap_res_X.t111 GNDA 0.345795f
C1953 cap_res_X.t76 GNDA 0.185733f
C1954 cap_res_X.n6 GNDA 0.198781f
C1955 cap_res_X.t7 GNDA 0.345795f
C1956 cap_res_X.t29 GNDA 0.185733f
C1957 cap_res_X.n7 GNDA 0.197177f
C1958 cap_res_X.t53 GNDA 0.345795f
C1959 cap_res_X.t21 GNDA 0.185733f
C1960 cap_res_X.n8 GNDA 0.197177f
C1961 cap_res_X.t88 GNDA 0.345795f
C1962 cap_res_X.t113 GNDA 0.185733f
C1963 cap_res_X.n9 GNDA 0.197177f
C1964 cap_res_X.t40 GNDA 0.345795f
C1965 cap_res_X.t112 GNDA 0.185733f
C1966 cap_res_X.n10 GNDA 0.197177f
C1967 cap_res_X.t94 GNDA 0.345795f
C1968 cap_res_X.t96 GNDA 0.185733f
C1969 cap_res_X.n11 GNDA 0.197177f
C1970 cap_res_X.t129 GNDA 0.345795f
C1971 cap_res_X.t46 GNDA 0.185733f
C1972 cap_res_X.n12 GNDA 0.197177f
C1973 cap_res_X.t24 GNDA 0.345795f
C1974 cap_res_X.t138 GNDA 0.185733f
C1975 cap_res_X.n13 GNDA 0.197177f
C1976 cap_res_X.t60 GNDA 0.345795f
C1977 cap_res_X.t90 GNDA 0.185733f
C1978 cap_res_X.n14 GNDA 0.197177f
C1979 cap_res_X.t121 GNDA 0.345795f
C1980 cap_res_X.t27 GNDA 0.347048f
C1981 cap_res_X.t36 GNDA 0.345795f
C1982 cap_res_X.t10 GNDA 0.347048f
C1983 cap_res_X.t114 GNDA 0.167175f
C1984 cap_res_X.n15 GNDA 0.215631f
C1985 cap_res_X.t74 GNDA 0.184584f
C1986 cap_res_X.n16 GNDA 0.234189f
C1987 cap_res_X.t41 GNDA 0.184584f
C1988 cap_res_X.n17 GNDA 0.251494f
C1989 cap_res_X.t57 GNDA 0.184584f
C1990 cap_res_X.n18 GNDA 0.251494f
C1991 cap_res_X.t19 GNDA 0.184584f
C1992 cap_res_X.n19 GNDA 0.251494f
C1993 cap_res_X.t50 GNDA 0.184584f
C1994 cap_res_X.n20 GNDA 0.251494f
C1995 cap_res_X.t16 GNDA 0.184584f
C1996 cap_res_X.n21 GNDA 0.251494f
C1997 cap_res_X.t117 GNDA 0.184584f
C1998 cap_res_X.n22 GNDA 0.251494f
C1999 cap_res_X.t12 GNDA 0.184584f
C2000 cap_res_X.n23 GNDA 0.251494f
C2001 cap_res_X.t110 GNDA 0.184584f
C2002 cap_res_X.n24 GNDA 0.251494f
C2003 cap_res_X.t66 GNDA 0.184584f
C2004 cap_res_X.n25 GNDA 0.251494f
C2005 cap_res_X.t26 GNDA 0.184584f
C2006 cap_res_X.n26 GNDA 0.251494f
C2007 cap_res_X.t63 GNDA 0.184584f
C2008 cap_res_X.n27 GNDA 0.251494f
C2009 cap_res_X.t23 GNDA 0.184584f
C2010 cap_res_X.n28 GNDA 0.251494f
C2011 cap_res_X.t125 GNDA 0.184584f
C2012 cap_res_X.n29 GNDA 0.251494f
C2013 cap_res_X.t18 GNDA 0.184584f
C2014 cap_res_X.n30 GNDA 0.251494f
C2015 cap_res_X.t47 GNDA 0.184584f
C2016 cap_res_X.n31 GNDA 0.234189f
C2017 cap_res_X.t28 GNDA 0.344645f
C2018 cap_res_X.t67 GNDA 0.167175f
C2019 cap_res_X.n32 GNDA 0.216884f
C2020 cap_res_X.t131 GNDA 0.344645f
C2021 cap_res_X.t30 GNDA 0.167175f
C2022 cap_res_X.n33 GNDA 0.216884f
C2023 cap_res_X.t93 GNDA 0.344645f
C2024 cap_res_X.t77 GNDA 0.345795f
C2025 cap_res_X.t35 GNDA 0.364353f
C2026 cap_res_X.t3 GNDA 0.364353f
C2027 cap_res_X.t31 GNDA 0.364353f
C2028 cap_res_X.t133 GNDA 0.185733f
C2029 cap_res_X.n34 GNDA 0.216884f
C2030 cap_res_X.t56 GNDA 0.344645f
C2031 cap_res_X.n35 GNDA 0.216884f
C2032 cap_res_X.t98 GNDA 0.185733f
C2033 cap_res_X.t2 GNDA 0.364353f
C2034 cap_res_X.t108 GNDA 0.364353f
C2035 cap_res_X.t9 GNDA 0.364353f
C2036 cap_res_X.t43 GNDA 0.337351f
C2037 cap_res_X.t0 GNDA 0.298183f
C2038 VOUT-.t9 GNDA 0.051003f
C2039 VOUT-.t8 GNDA 0.051003f
C2040 VOUT-.n0 GNDA 0.235943f
C2041 VOUT-.t7 GNDA 0.051003f
C2042 VOUT-.t4 GNDA 0.051003f
C2043 VOUT-.n1 GNDA 0.235153f
C2044 VOUT-.n2 GNDA 0.145313f
C2045 VOUT-.t3 GNDA 0.051003f
C2046 VOUT-.t17 GNDA 0.051003f
C2047 VOUT-.n3 GNDA 0.235153f
C2048 VOUT-.n4 GNDA 0.089445f
C2049 VOUT-.t15 GNDA 0.084326f
C2050 VOUT-.n5 GNDA 0.119504f
C2051 VOUT-.t13 GNDA 0.043717f
C2052 VOUT-.t6 GNDA 0.043717f
C2053 VOUT-.n6 GNDA 0.175711f
C2054 VOUT-.t16 GNDA 0.043717f
C2055 VOUT-.t12 GNDA 0.043717f
C2056 VOUT-.n7 GNDA 0.17571f
C2057 VOUT-.t5 GNDA 0.043717f
C2058 VOUT-.t18 GNDA 0.043717f
C2059 VOUT-.n8 GNDA 0.175387f
C2060 VOUT-.n9 GNDA 0.172777f
C2061 VOUT-.t10 GNDA 0.043717f
C2062 VOUT-.t11 GNDA 0.043717f
C2063 VOUT-.n10 GNDA 0.175387f
C2064 VOUT-.n11 GNDA 0.0891f
C2065 VOUT-.t2 GNDA 0.043717f
C2066 VOUT-.t1 GNDA 0.043717f
C2067 VOUT-.n12 GNDA 0.175387f
C2068 VOUT-.n13 GNDA 0.0891f
C2069 VOUT-.n14 GNDA 0.105535f
C2070 VOUT-.t0 GNDA 0.043717f
C2071 VOUT-.t14 GNDA 0.043717f
C2072 VOUT-.n15 GNDA 0.17324f
C2073 VOUT-.n16 GNDA 0.211953f
C2074 VOUT-.t43 GNDA 0.291446f
C2075 VOUT-.t121 GNDA 0.29641f
C2076 VOUT-.t147 GNDA 0.291446f
C2077 VOUT-.n17 GNDA 0.195405f
C2078 VOUT-.n18 GNDA 0.127508f
C2079 VOUT-.t97 GNDA 0.295788f
C2080 VOUT-.t133 GNDA 0.295788f
C2081 VOUT-.t28 GNDA 0.295788f
C2082 VOUT-.t63 GNDA 0.295788f
C2083 VOUT-.t117 GNDA 0.295788f
C2084 VOUT-.t69 GNDA 0.295788f
C2085 VOUT-.t104 GNDA 0.295788f
C2086 VOUT-.t150 GNDA 0.295788f
C2087 VOUT-.t46 GNDA 0.295788f
C2088 VOUT-.t86 GNDA 0.295788f
C2089 VOUT-.t29 GNDA 0.291446f
C2090 VOUT-.n19 GNDA 0.196026f
C2091 VOUT-.t81 GNDA 0.291446f
C2092 VOUT-.n20 GNDA 0.250673f
C2093 VOUT-.t128 GNDA 0.291446f
C2094 VOUT-.n21 GNDA 0.250673f
C2095 VOUT-.t136 GNDA 0.291446f
C2096 VOUT-.n22 GNDA 0.250673f
C2097 VOUT-.t44 GNDA 0.291446f
C2098 VOUT-.n23 GNDA 0.250673f
C2099 VOUT-.t45 GNDA 0.291446f
C2100 VOUT-.n24 GNDA 0.250673f
C2101 VOUT-.t61 GNDA 0.291446f
C2102 VOUT-.n25 GNDA 0.250673f
C2103 VOUT-.t111 GNDA 0.291446f
C2104 VOUT-.n26 GNDA 0.250673f
C2105 VOUT-.t19 GNDA 0.291446f
C2106 VOUT-.n27 GNDA 0.250673f
C2107 VOUT-.t67 GNDA 0.291446f
C2108 VOUT-.n28 GNDA 0.250673f
C2109 VOUT-.t83 GNDA 0.291446f
C2110 VOUT-.t36 GNDA 0.29641f
C2111 VOUT-.t130 GNDA 0.291446f
C2112 VOUT-.n29 GNDA 0.195405f
C2113 VOUT-.n30 GNDA 0.2368f
C2114 VOUT-.t105 GNDA 0.29641f
C2115 VOUT-.t151 GNDA 0.291446f
C2116 VOUT-.n31 GNDA 0.195405f
C2117 VOUT-.t116 GNDA 0.291446f
C2118 VOUT-.t76 GNDA 0.29641f
C2119 VOUT-.t25 GNDA 0.291446f
C2120 VOUT-.n32 GNDA 0.195405f
C2121 VOUT-.n33 GNDA 0.2368f
C2122 VOUT-.t42 GNDA 0.29641f
C2123 VOUT-.t146 GNDA 0.291446f
C2124 VOUT-.n34 GNDA 0.195405f
C2125 VOUT-.t100 GNDA 0.291446f
C2126 VOUT-.t30 GNDA 0.29641f
C2127 VOUT-.t66 GNDA 0.291446f
C2128 VOUT-.n35 GNDA 0.195405f
C2129 VOUT-.n36 GNDA 0.2368f
C2130 VOUT-.t88 GNDA 0.29641f
C2131 VOUT-.t48 GNDA 0.291446f
C2132 VOUT-.n37 GNDA 0.195405f
C2133 VOUT-.t138 GNDA 0.291446f
C2134 VOUT-.t72 GNDA 0.29641f
C2135 VOUT-.t108 GNDA 0.291446f
C2136 VOUT-.n38 GNDA 0.195405f
C2137 VOUT-.n39 GNDA 0.2368f
C2138 VOUT-.t51 GNDA 0.29641f
C2139 VOUT-.t153 GNDA 0.291446f
C2140 VOUT-.n40 GNDA 0.195405f
C2141 VOUT-.t107 GNDA 0.291446f
C2142 VOUT-.t33 GNDA 0.29641f
C2143 VOUT-.t71 GNDA 0.291446f
C2144 VOUT-.n41 GNDA 0.195405f
C2145 VOUT-.n42 GNDA 0.2368f
C2146 VOUT-.t92 GNDA 0.29641f
C2147 VOUT-.t53 GNDA 0.291446f
C2148 VOUT-.n43 GNDA 0.195405f
C2149 VOUT-.t141 GNDA 0.291446f
C2150 VOUT-.t77 GNDA 0.29641f
C2151 VOUT-.t112 GNDA 0.291446f
C2152 VOUT-.n44 GNDA 0.195405f
C2153 VOUT-.n45 GNDA 0.2368f
C2154 VOUT-.t143 GNDA 0.291446f
C2155 VOUT-.t74 GNDA 0.29641f
C2156 VOUT-.t113 GNDA 0.291446f
C2157 VOUT-.n46 GNDA 0.195405f
C2158 VOUT-.n47 GNDA 0.127508f
C2159 VOUT-.t129 GNDA 0.295788f
C2160 VOUT-.t26 GNDA 0.295788f
C2161 VOUT-.t80 GNDA 0.29641f
C2162 VOUT-.t122 GNDA 0.291446f
C2163 VOUT-.n48 GNDA 0.195405f
C2164 VOUT-.t154 GNDA 0.291446f
C2165 VOUT-.n49 GNDA 0.127508f
C2166 VOUT-.t126 GNDA 0.291446f
C2167 VOUT-.n50 GNDA 0.122954f
C2168 VOUT-.t64 GNDA 0.295788f
C2169 VOUT-.t114 GNDA 0.29641f
C2170 VOUT-.t148 GNDA 0.291446f
C2171 VOUT-.n51 GNDA 0.195405f
C2172 VOUT-.t49 GNDA 0.291446f
C2173 VOUT-.n52 GNDA 0.127508f
C2174 VOUT-.t155 GNDA 0.291446f
C2175 VOUT-.n53 GNDA 0.122954f
C2176 VOUT-.t101 GNDA 0.295788f
C2177 VOUT-.t22 GNDA 0.29641f
C2178 VOUT-.t62 GNDA 0.291446f
C2179 VOUT-.n54 GNDA 0.195405f
C2180 VOUT-.t103 GNDA 0.291446f
C2181 VOUT-.n55 GNDA 0.127508f
C2182 VOUT-.t68 GNDA 0.291446f
C2183 VOUT-.n56 GNDA 0.122954f
C2184 VOUT-.t82 GNDA 0.295788f
C2185 VOUT-.t123 GNDA 0.29641f
C2186 VOUT-.t156 GNDA 0.291446f
C2187 VOUT-.n57 GNDA 0.195405f
C2188 VOUT-.t54 GNDA 0.291446f
C2189 VOUT-.n58 GNDA 0.127508f
C2190 VOUT-.t23 GNDA 0.291446f
C2191 VOUT-.n59 GNDA 0.122954f
C2192 VOUT-.t56 GNDA 0.295788f
C2193 VOUT-.t98 GNDA 0.295788f
C2194 VOUT-.t78 GNDA 0.295788f
C2195 VOUT-.t118 GNDA 0.295788f
C2196 VOUT-.t149 GNDA 0.295788f
C2197 VOUT-.t115 GNDA 0.291446f
C2198 VOUT-.n60 GNDA 0.196026f
C2199 VOUT-.t75 GNDA 0.291446f
C2200 VOUT-.n61 GNDA 0.250673f
C2201 VOUT-.t34 GNDA 0.291446f
C2202 VOUT-.n62 GNDA 0.250673f
C2203 VOUT-.t55 GNDA 0.291446f
C2204 VOUT-.n63 GNDA 0.250673f
C2205 VOUT-.t20 GNDA 0.291446f
C2206 VOUT-.n64 GNDA 0.309872f
C2207 VOUT-.t37 GNDA 0.291446f
C2208 VOUT-.n65 GNDA 0.309872f
C2209 VOUT-.t59 GNDA 0.291446f
C2210 VOUT-.n66 GNDA 0.309872f
C2211 VOUT-.t24 GNDA 0.291446f
C2212 VOUT-.n67 GNDA 0.309872f
C2213 VOUT-.t127 GNDA 0.291446f
C2214 VOUT-.n68 GNDA 0.250673f
C2215 VOUT-.t90 GNDA 0.291446f
C2216 VOUT-.n69 GNDA 0.250673f
C2217 VOUT-.t110 GNDA 0.291446f
C2218 VOUT-.t31 GNDA 0.29641f
C2219 VOUT-.t73 GNDA 0.291446f
C2220 VOUT-.n70 GNDA 0.195405f
C2221 VOUT-.n71 GNDA 0.2368f
C2222 VOUT-.t89 GNDA 0.29641f
C2223 VOUT-.t50 GNDA 0.291446f
C2224 VOUT-.n72 GNDA 0.195405f
C2225 VOUT-.t139 GNDA 0.291446f
C2226 VOUT-.t70 GNDA 0.29641f
C2227 VOUT-.t109 GNDA 0.291446f
C2228 VOUT-.n73 GNDA 0.195405f
C2229 VOUT-.n74 GNDA 0.2368f
C2230 VOUT-.t125 GNDA 0.29641f
C2231 VOUT-.t87 GNDA 0.291446f
C2232 VOUT-.n75 GNDA 0.195405f
C2233 VOUT-.t32 GNDA 0.291446f
C2234 VOUT-.t106 GNDA 0.29641f
C2235 VOUT-.t137 GNDA 0.291446f
C2236 VOUT-.n76 GNDA 0.195405f
C2237 VOUT-.n77 GNDA 0.2368f
C2238 VOUT-.t85 GNDA 0.29641f
C2239 VOUT-.t41 GNDA 0.291446f
C2240 VOUT-.n78 GNDA 0.195405f
C2241 VOUT-.t134 GNDA 0.291446f
C2242 VOUT-.t65 GNDA 0.29641f
C2243 VOUT-.t99 GNDA 0.291446f
C2244 VOUT-.n79 GNDA 0.195405f
C2245 VOUT-.n80 GNDA 0.2368f
C2246 VOUT-.t39 GNDA 0.29641f
C2247 VOUT-.t142 GNDA 0.291446f
C2248 VOUT-.n81 GNDA 0.195405f
C2249 VOUT-.t94 GNDA 0.291446f
C2250 VOUT-.t27 GNDA 0.29641f
C2251 VOUT-.t58 GNDA 0.291446f
C2252 VOUT-.n82 GNDA 0.195405f
C2253 VOUT-.n83 GNDA 0.2368f
C2254 VOUT-.t79 GNDA 0.29641f
C2255 VOUT-.t38 GNDA 0.291446f
C2256 VOUT-.n84 GNDA 0.195405f
C2257 VOUT-.t131 GNDA 0.291446f
C2258 VOUT-.t57 GNDA 0.29641f
C2259 VOUT-.t93 GNDA 0.291446f
C2260 VOUT-.n85 GNDA 0.195405f
C2261 VOUT-.n86 GNDA 0.2368f
C2262 VOUT-.t35 GNDA 0.29641f
C2263 VOUT-.t140 GNDA 0.291446f
C2264 VOUT-.n87 GNDA 0.195405f
C2265 VOUT-.t91 GNDA 0.291446f
C2266 VOUT-.t21 GNDA 0.29641f
C2267 VOUT-.t52 GNDA 0.291446f
C2268 VOUT-.n88 GNDA 0.195405f
C2269 VOUT-.n89 GNDA 0.2368f
C2270 VOUT-.t135 GNDA 0.29641f
C2271 VOUT-.t102 GNDA 0.291446f
C2272 VOUT-.n90 GNDA 0.195405f
C2273 VOUT-.t47 GNDA 0.291446f
C2274 VOUT-.t124 GNDA 0.29641f
C2275 VOUT-.t152 GNDA 0.291446f
C2276 VOUT-.n91 GNDA 0.195405f
C2277 VOUT-.n92 GNDA 0.2368f
C2278 VOUT-.t96 GNDA 0.29641f
C2279 VOUT-.t60 GNDA 0.291446f
C2280 VOUT-.n93 GNDA 0.195405f
C2281 VOUT-.t145 GNDA 0.291446f
C2282 VOUT-.t84 GNDA 0.29641f
C2283 VOUT-.t120 GNDA 0.291446f
C2284 VOUT-.n94 GNDA 0.195405f
C2285 VOUT-.n95 GNDA 0.2368f
C2286 VOUT-.t119 GNDA 0.29641f
C2287 VOUT-.t144 GNDA 0.291446f
C2288 VOUT-.n96 GNDA 0.195405f
C2289 VOUT-.t40 GNDA 0.291446f
C2290 VOUT-.n97 GNDA 0.2368f
C2291 VOUT-.t95 GNDA 0.291446f
C2292 VOUT-.n98 GNDA 0.127508f
C2293 VOUT-.t132 GNDA 0.291446f
C2294 VOUT-.n99 GNDA 0.23878f
C2295 VOUT-.n100 GNDA 0.268998f
.ends

