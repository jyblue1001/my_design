* PEX produced on Wed Aug 20 07:39:19 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic_17.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic_17 VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 VDDA.t211 bgr_11_0.1st_Vout_2.t7 bgr_11_0.PFET_GATE_10uA.t9 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X1 VOUT-.t19 two_stage_opamp_dummy_magic_24_0.cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2 VOUT+.t19 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 VDDA.t362 two_stage_opamp_dummy_magic_24_0.Vb3.t8 two_stage_opamp_dummy_magic_24_0.VD4.t26 VDDA.t361 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X4 VOUT-.t20 two_stage_opamp_dummy_magic_24_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5 VDDA.t108 two_stage_opamp_dummy_magic_24_0.Vb3.t9 two_stage_opamp_dummy_magic_24_0.VD3.t31 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X6 two_stage_opamp_dummy_magic_24_0.VD2.t9 VIN+.t0 two_stage_opamp_dummy_magic_24_0.V_source.t9 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X7 GNDA.t160 GNDA.t158 two_stage_opamp_dummy_magic_24_0.Vb2.t3 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X8 two_stage_opamp_dummy_magic_24_0.VD3.t7 two_stage_opamp_dummy_magic_24_0.Vb2.t11 two_stage_opamp_dummy_magic_24_0.X.t14 two_stage_opamp_dummy_magic_24_0.VD3.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X9 VOUT-.t21 two_stage_opamp_dummy_magic_24_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 two_stage_opamp_dummy_magic_24_0.V_source.t28 two_stage_opamp_dummy_magic_24_0.Vb1.t12 two_stage_opamp_dummy_magic_24_0.Vb1_2.t4 GNDA.t229 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.6 ps=3.8 w=1.5 l=3
X11 VOUT+.t7 two_stage_opamp_dummy_magic_24_0.Y.t25 VDDA.t150 VDDA.t149 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X12 GNDA.t269 VDDA.t358 VDDA.t360 VDDA.t359 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X13 GNDA.t241 two_stage_opamp_dummy_magic_24_0.Y.t26 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t15 VDDA.t160 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X14 VOUT-.t22 two_stage_opamp_dummy_magic_24_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 VDDA.t385 bgr_11_0.V_TOP.t14 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t3 VDDA.t384 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X16 bgr_11_0.1st_Vout_1.t7 bgr_11_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 VDDA.t148 two_stage_opamp_dummy_magic_24_0.Y.t27 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t14 GNDA.t223 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X18 VOUT+.t20 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X19 VOUT-.t23 two_stage_opamp_dummy_magic_24_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 GNDA.t47 bgr_11_0.NFET_GATE_10uA.t5 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t1 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X21 two_stage_opamp_dummy_magic_24_0.VD2.t20 two_stage_opamp_dummy_magic_24_0.Vb1.t13 two_stage_opamp_dummy_magic_24_0.Y.t22 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X22 bgr_11_0.V_TOP.t15 VDDA.t386 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X23 two_stage_opamp_dummy_magic_24_0.Vb2.t2 GNDA.t155 GNDA.t157 GNDA.t156 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X24 VOUT-.t24 two_stage_opamp_dummy_magic_24_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 two_stage_opamp_dummy_magic_24_0.V_err_gate.t5 VDDA.t355 VDDA.t357 VDDA.t356 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X26 two_stage_opamp_dummy_magic_24_0.V_source.t18 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t12 GNDA.t52 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X27 bgr_11_0.START_UP_NFET1.t0 bgr_11_0.START_UP_NFET1 GNDA.t176 GNDA.t175 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X28 bgr_11_0.1st_Vout_1.t0 bgr_11_0.V_mir1.t13 VDDA.t11 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X29 two_stage_opamp_dummy_magic_24_0.V_err_p.t1 two_stage_opamp_dummy_magic_24_0.V_tot.t4 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t3 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X30 VDDA.t87 two_stage_opamp_dummy_magic_24_0.Vb3.t10 two_stage_opamp_dummy_magic_24_0.VD4.t25 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X31 VOUT-.t25 two_stage_opamp_dummy_magic_24_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 bgr_11_0.V_TOP.t16 VDDA.t392 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 GNDA.t285 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t13 two_stage_opamp_dummy_magic_24_0.V_source.t39 GNDA.t284 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X34 VOUT-.t2 two_stage_opamp_dummy_magic_24_0.X.t25 VDDA.t112 VDDA.t111 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X35 VOUT+.t21 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 two_stage_opamp_dummy_magic_24_0.VD3.t21 VDDA.t352 VDDA.t354 VDDA.t353 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X37 VOUT-.t14 two_stage_opamp_dummy_magic_24_0.X.t26 VDDA.t375 VDDA.t374 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X38 GNDA.t18 two_stage_opamp_dummy_magic_24_0.X.t27 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t9 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X39 a_6350_30238.t1 bgr_11_0.Vin+.t5 GNDA.t13 sky130_fd_pr__res_xhigh_po_0p35 l=6
X40 GNDA.t154 GNDA.t152 VDDA.t104 GNDA.t153 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X41 bgr_11_0.V_TOP.t17 VDDA.t393 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 two_stage_opamp_dummy_magic_24_0.V_err_gate.t3 bgr_11_0.NFET_GATE_10uA.t6 GNDA.t188 GNDA.t187 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X43 VOUT+.t22 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 VOUT-.t26 two_stage_opamp_dummy_magic_24_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 VOUT-.t27 two_stage_opamp_dummy_magic_24_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 VDDA.t159 a_6540_22450.t11 a_6540_22450.t12 VDDA.t158 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X47 VOUT-.t28 two_stage_opamp_dummy_magic_24_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X48 VOUT-.t29 two_stage_opamp_dummy_magic_24_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 VDDA.t81 two_stage_opamp_dummy_magic_24_0.Vb3.t11 two_stage_opamp_dummy_magic_24_0.VD4.t24 VDDA.t80 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X50 VDDA.t65 two_stage_opamp_dummy_magic_24_0.X.t28 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t9 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X51 VOUT-.t30 two_stage_opamp_dummy_magic_24_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 VDDA.t199 bgr_11_0.V_mir1.t11 bgr_11_0.V_mir1.t12 VDDA.t198 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X53 VOUT+.t23 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X54 VDDA.t351 VDDA.t349 two_stage_opamp_dummy_magic_24_0.V_err_gate.t4 VDDA.t350 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X55 VOUT+.t24 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X56 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t0 GNDA.t150 GNDA.t151 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X57 two_stage_opamp_dummy_magic_24_0.VD1.t21 VIN-.t0 two_stage_opamp_dummy_magic_24_0.V_source.t15 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X58 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t3 bgr_11_0.PFET_GATE_10uA.t10 VDDA.t249 VDDA.t248 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X59 VOUT+.t25 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X60 VDDA.t247 bgr_11_0.PFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t2 VDDA.t246 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X61 bgr_11_0.V_TOP.t18 VDDA.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X62 bgr_11_0.cap_res1.t20 bgr_11_0.V_TOP.t6 GNDA.t194 sky130_fd_pr__res_high_po_0p35 l=2.05
X63 VOUT+.t26 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X64 two_stage_opamp_dummy_magic_24_0.VD2.t12 GNDA.t148 GNDA.t149 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X65 two_stage_opamp_dummy_magic_24_0.Vb1.t5 two_stage_opamp_dummy_magic_24_0.Vb1.t4 two_stage_opamp_dummy_magic_24_0.Vb1_2.t3 GNDA.t307 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X66 two_stage_opamp_dummy_magic_24_0.VD3.t5 two_stage_opamp_dummy_magic_24_0.Vb2.t12 two_stage_opamp_dummy_magic_24_0.X.t13 two_stage_opamp_dummy_magic_24_0.VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X67 VOUT+.t27 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 VOUT+.t12 VDDA.t346 VDDA.t348 VDDA.t347 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X69 GNDA.t147 GNDA.t146 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t3 GNDA.t86 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X70 two_stage_opamp_dummy_magic_24_0.VD1.t20 VIN-.t1 two_stage_opamp_dummy_magic_24_0.V_source.t38 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X71 VOUT-.t31 two_stage_opamp_dummy_magic_24_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 VOUT+.t18 two_stage_opamp_dummy_magic_24_0.Y.t28 VDDA.t418 VDDA.t417 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X73 two_stage_opamp_dummy_magic_24_0.X.t12 two_stage_opamp_dummy_magic_24_0.Vb2.t13 two_stage_opamp_dummy_magic_24_0.VD3.t3 two_stage_opamp_dummy_magic_24_0.VD3.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X74 GNDA.t263 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t2 VOUT+.t10 GNDA.t262 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X75 GNDA.t295 two_stage_opamp_dummy_magic_24_0.Y.t29 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t14 VDDA.t404 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X76 VOUT-.t32 two_stage_opamp_dummy_magic_24_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X77 bgr_11_0.V_TOP.t19 VDDA.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X78 VOUT-.t33 two_stage_opamp_dummy_magic_24_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 VOUT-.t34 two_stage_opamp_dummy_magic_24_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X80 bgr_11_0.1st_Vout_2.t8 bgr_11_0.cap_res2.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X81 VOUT+.t28 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X82 GNDA.t62 GNDA.t145 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X83 two_stage_opamp_dummy_magic_24_0.VD4.t8 two_stage_opamp_dummy_magic_24_0.Vb2.t14 two_stage_opamp_dummy_magic_24_0.Y.t11 two_stage_opamp_dummy_magic_24_0.VD4.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X84 VDDA.t121 two_stage_opamp_dummy_magic_24_0.Vb3.t12 two_stage_opamp_dummy_magic_24_0.VD4.t23 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X85 VOUT+.t29 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X86 VOUT+.t30 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X87 VOUT+.t31 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 two_stage_opamp_dummy_magic_24_0.VD2.t11 two_stage_opamp_dummy_magic_24_0.Vb1.t14 two_stage_opamp_dummy_magic_24_0.Y.t21 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X89 two_stage_opamp_dummy_magic_24_0.Vb2_2.t8 two_stage_opamp_dummy_magic_24_0.Vb2_2.t6 two_stage_opamp_dummy_magic_24_0.Vb2_2.t8 two_stage_opamp_dummy_magic_24_0.Vb2_2.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X90 VDDA.t209 bgr_11_0.1st_Vout_2.t9 bgr_11_0.PFET_GATE_10uA.t8 VDDA.t208 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X91 VOUT-.t35 two_stage_opamp_dummy_magic_24_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X92 two_stage_opamp_dummy_magic_24_0.VD3.t30 two_stage_opamp_dummy_magic_24_0.Vb3.t13 VDDA.t369 VDDA.t368 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X93 bgr_11_0.1st_Vout_2.t10 bgr_11_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X94 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t11 bgr_11_0.PFET_GATE_10uA.t12 VDDA.t245 VDDA.t244 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X95 GNDA.t144 GNDA.t142 VOUT+.t8 GNDA.t143 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X96 VOUT+.t32 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 VOUT-.t36 two_stage_opamp_dummy_magic_24_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X98 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 bgr_11_0.Vin+.t4 GNDA.t165 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X99 VOUT-.t37 two_stage_opamp_dummy_magic_24_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 VOUT-.t38 two_stage_opamp_dummy_magic_24_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X101 VOUT+.t33 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X102 bgr_11_0.1st_Vout_1.t8 bgr_11_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X103 VDDA.t345 VDDA.t343 GNDA.t268 VDDA.t344 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X104 VOUT-.t39 two_stage_opamp_dummy_magic_24_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 VOUT-.t40 two_stage_opamp_dummy_magic_24_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X106 bgr_11_0.1st_Vout_2.t11 bgr_11_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 VOUT-.t3 two_stage_opamp_dummy_magic_24_0.X.t29 VDDA.t135 VDDA.t134 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X108 VOUT-.t41 two_stage_opamp_dummy_magic_24_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X109 bgr_11_0.V_TOP.t20 VDDA.t181 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X110 GNDA.t204 two_stage_opamp_dummy_magic_24_0.X.t30 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t8 VDDA.t127 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X111 VDDA.t243 bgr_11_0.PFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t14 VDDA.t242 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X112 VOUT+.t34 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 VOUT+.t35 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t16 VDDA.t340 VDDA.t342 VDDA.t341 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X115 two_stage_opamp_dummy_magic_24_0.V_source.t17 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t14 GNDA.t50 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X116 VDDA.t169 a_6540_22450.t13 bgr_11_0.1st_Vout_2.t5 VDDA.t168 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X117 VOUT+.t36 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X118 VOUT+.t37 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 VDDA.t183 bgr_11_0.V_TOP.t21 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t2 VDDA.t182 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X120 VDDA.t84 GNDA.t139 GNDA.t141 GNDA.t140 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X121 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.t3 two_stage_opamp_dummy_magic_24_0.V_err_gate.t6 VDDA.t119 VDDA.t118 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X122 VOUT+.t38 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 two_stage_opamp_dummy_magic_24_0.Y.t24 two_stage_opamp_dummy_magic_24_0.VD4.t30 two_stage_opamp_dummy_magic_24_0.VD4.t32 two_stage_opamp_dummy_magic_24_0.VD4.t31 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X124 two_stage_opamp_dummy_magic_24_0.VD1.t19 VIN-.t2 two_stage_opamp_dummy_magic_24_0.V_source.t37 GNDA.t205 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X125 GNDA.t6 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t15 two_stage_opamp_dummy_magic_24_0.V_source.t2 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X126 two_stage_opamp_dummy_magic_24_0.VD4.t22 two_stage_opamp_dummy_magic_24_0.Vb3.t14 VDDA.t75 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X127 VOUT-.t42 two_stage_opamp_dummy_magic_24_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 two_stage_opamp_dummy_magic_24_0.VD3.t29 two_stage_opamp_dummy_magic_24_0.Vb3.t15 VDDA.t77 VDDA.t76 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X129 VOUT+.t39 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 two_stage_opamp_dummy_magic_24_0.X.t11 two_stage_opamp_dummy_magic_24_0.Vb2.t15 two_stage_opamp_dummy_magic_24_0.VD3.t1 two_stage_opamp_dummy_magic_24_0.VD3.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X131 VOUT-.t43 two_stage_opamp_dummy_magic_24_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X132 VOUT+.t40 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t0 a_13940_n594.t0 GNDA.t167 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X134 VOUT+.t41 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X135 VOUT-.t44 two_stage_opamp_dummy_magic_24_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X136 GNDA.t162 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t16 two_stage_opamp_dummy_magic_24_0.V_p_mir.t1 GNDA.t161 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X137 VOUT-.t45 two_stage_opamp_dummy_magic_24_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 bgr_11_0.1st_Vout_2.t12 bgr_11_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 two_stage_opamp_dummy_magic_24_0.Vb1.t7 two_stage_opamp_dummy_magic_24_0.Vb1.t6 two_stage_opamp_dummy_magic_24_0.Vb1_2.t2 GNDA.t193 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X140 two_stage_opamp_dummy_magic_24_0.VD1.t18 VIN-.t3 two_stage_opamp_dummy_magic_24_0.V_source.t27 GNDA.t227 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X141 bgr_11_0.V_TOP.t22 VDDA.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X142 VOUT+.t17 two_stage_opamp_dummy_magic_24_0.Y.t30 VDDA.t416 VDDA.t415 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X143 VOUT+.t42 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 VOUT+.t43 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 VOUT-.t46 two_stage_opamp_dummy_magic_24_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X146 two_stage_opamp_dummy_magic_24_0.VD1.t11 two_stage_opamp_dummy_magic_24_0.Vb1.t15 two_stage_opamp_dummy_magic_24_0.X.t16 GNDA.t177 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X147 VOUT+.t44 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t6 VDDA.t337 VDDA.t339 VDDA.t338 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X149 two_stage_opamp_dummy_magic_24_0.V_source.t31 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t17 GNDA.t246 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X150 a_13840_3288.t1 two_stage_opamp_dummy_magic_24_0.V_tot.t0 GNDA.t230 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X151 GNDA.t198 bgr_11_0.NFET_GATE_10uA.t7 two_stage_opamp_dummy_magic_24_0.Vb3.t3 GNDA.t197 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X152 VOUT+.t45 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X153 two_stage_opamp_dummy_magic_24_0.VD2.t14 two_stage_opamp_dummy_magic_24_0.Vb1.t16 two_stage_opamp_dummy_magic_24_0.Y.t20 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X154 GNDA.t138 GNDA.t137 two_stage_opamp_dummy_magic_24_0.VD1.t1 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X155 GNDA.t171 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t18 two_stage_opamp_dummy_magic_24_0.V_source.t20 GNDA.t170 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X156 VDDA.t391 a_6540_22450.t9 a_6540_22450.t10 VDDA.t390 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X157 bgr_11_0.START_UP.t3 bgr_11_0.V_TOP.t23 VDDA.t57 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X158 two_stage_opamp_dummy_magic_24_0.VD1.t10 two_stage_opamp_dummy_magic_24_0.Vb1.t17 two_stage_opamp_dummy_magic_24_0.X.t15 GNDA.t172 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X159 VOUT-.t47 two_stage_opamp_dummy_magic_24_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X160 VOUT-.t48 two_stage_opamp_dummy_magic_24_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X161 VOUT-.t49 two_stage_opamp_dummy_magic_24_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 VOUT+.t46 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X163 VOUT+.t47 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 a_11420_30238.t1 bgr_11_0.Vin-.t7 GNDA.t309 sky130_fd_pr__res_xhigh_po_0p35 l=6
X165 bgr_11_0.V_TOP.t13 VDDA.t334 VDDA.t336 VDDA.t335 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.45 ps=2.9 w=1 l=0.15
X166 a_11300_30238.t1 a_11950_28880.t1 GNDA.t305 sky130_fd_pr__res_xhigh_po_0p35 l=4
X167 VOUT+.t48 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X168 GNDA.t136 GNDA.t135 two_stage_opamp_dummy_magic_24_0.VD2.t19 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X169 VOUT+.t49 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X170 bgr_11_0.V_TOP.t24 VDDA.t139 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 VDDA.t371 two_stage_opamp_dummy_magic_24_0.Vb3.t16 two_stage_opamp_dummy_magic_24_0.VD3.t28 VDDA.t370 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X172 VOUT-.t50 two_stage_opamp_dummy_magic_24_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X173 VDDA.t333 VDDA.t331 VOUT+.t11 VDDA.t332 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X174 VOUT+.t50 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 VOUT+.t3 GNDA.t132 GNDA.t134 GNDA.t133 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X176 VOUT+.t51 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 VOUT+.t52 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X178 bgr_11_0.Vin+.t3 bgr_11_0.V_TOP.t25 VDDA.t141 VDDA.t140 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X179 VOUT+.t53 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X180 VOUT+.t54 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 VOUT+.t55 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 VOUT-.t8 two_stage_opamp_dummy_magic_24_0.X.t31 VDDA.t172 VDDA.t171 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X183 VDDA.t197 bgr_11_0.V_mir1.t14 bgr_11_0.1st_Vout_1.t5 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X184 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t4 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0 ps=0 w=3.5 l=0.2
X185 two_stage_opamp_dummy_magic_24_0.Y.t10 two_stage_opamp_dummy_magic_24_0.Vb2.t16 two_stage_opamp_dummy_magic_24_0.VD4.t3 two_stage_opamp_dummy_magic_24_0.VD4.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X186 two_stage_opamp_dummy_magic_24_0.VD4.t21 two_stage_opamp_dummy_magic_24_0.Vb3.t17 VDDA.t4 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X187 GNDA.t267 VDDA.t328 VDDA.t330 VDDA.t329 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X188 VOUT-.t51 two_stage_opamp_dummy_magic_24_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 VOUT+.t56 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X190 VOUT-.t52 two_stage_opamp_dummy_magic_24_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 bgr_11_0.1st_Vout_2.t13 bgr_11_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 VDDA.t327 VDDA.t324 VDDA.t326 VDDA.t325 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.15
X193 VDDA.t323 VDDA.t320 VDDA.t322 VDDA.t321 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0 ps=0 w=1 l=0.15
X194 VOUT-.t53 two_stage_opamp_dummy_magic_24_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 VOUT-.t54 two_stage_opamp_dummy_magic_24_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 VDDA.t241 bgr_11_0.PFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t10 VDDA.t240 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X197 VOUT+.t57 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 VOUT-.t55 two_stage_opamp_dummy_magic_24_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 VOUT+.t9 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t3 GNDA.t257 GNDA.t256 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X200 GNDA.t252 bgr_11_0.NFET_GATE_10uA.t8 two_stage_opamp_dummy_magic_24_0.Vb2.t9 GNDA.t251 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X201 VOUT+.t58 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 two_stage_opamp_dummy_magic_24_0.X.t10 two_stage_opamp_dummy_magic_24_0.Vb2.t17 two_stage_opamp_dummy_magic_24_0.VD3.t37 two_stage_opamp_dummy_magic_24_0.VD3.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X203 VOUT-.t56 two_stage_opamp_dummy_magic_24_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X204 VOUT+.t59 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X205 two_stage_opamp_dummy_magic_24_0.Vb2.t6 bgr_11_0.NFET_GATE_10uA.t9 GNDA.t184 GNDA.t183 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X206 VDDA.t178 bgr_11_0.V_TOP.t26 bgr_11_0.Vin-.t3 VDDA.t177 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X207 VDDA.t319 VDDA.t317 bgr_11_0.V_TOP.t12 VDDA.t318 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X208 VOUT-.t57 two_stage_opamp_dummy_magic_24_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 two_stage_opamp_dummy_magic_24_0.V_source.t0 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t19 GNDA.t2 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X210 two_stage_opamp_dummy_magic_24_0.Vb1.t1 GNDA.t129 GNDA.t131 GNDA.t130 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X211 GNDA.t62 GNDA.t128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X212 VOUT+.t60 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 two_stage_opamp_dummy_magic_24_0.VD1.t0 GNDA.t126 GNDA.t127 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X214 two_stage_opamp_dummy_magic_24_0.Y.t9 two_stage_opamp_dummy_magic_24_0.Vb2.t18 two_stage_opamp_dummy_magic_24_0.VD4.t34 two_stage_opamp_dummy_magic_24_0.VD4.t33 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X215 two_stage_opamp_dummy_magic_24_0.VD4.t20 two_stage_opamp_dummy_magic_24_0.Vb3.t18 VDDA.t2 VDDA.t1 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X216 two_stage_opamp_dummy_magic_24_0.VD1.t9 two_stage_opamp_dummy_magic_24_0.Vb1.t18 two_stage_opamp_dummy_magic_24_0.X.t4 GNDA.t166 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X217 bgr_11_0.1st_Vout_1.t9 bgr_11_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X218 GNDA.t186 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t20 two_stage_opamp_dummy_magic_24_0.V_source.t22 GNDA.t185 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X219 GNDA.t101 GNDA.t118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X220 VDDA.t189 bgr_11_0.1st_Vout_1.t10 bgr_11_0.V_TOP.t8 VDDA.t188 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X221 VOUT-.t58 two_stage_opamp_dummy_magic_24_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 VOUT-.t59 two_stage_opamp_dummy_magic_24_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 VOUT-.t60 two_stage_opamp_dummy_magic_24_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X224 bgr_11_0.START_UP.t5 bgr_11_0.START_UP.t4 bgr_11_0.START_UP_NFET1.t0 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X225 GNDA.t125 GNDA.t123 VDDA.t124 GNDA.t124 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X226 VOUT-.t61 two_stage_opamp_dummy_magic_24_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X227 VDDA.t364 two_stage_opamp_dummy_magic_24_0.Vb3.t19 two_stage_opamp_dummy_magic_24_0.VD3.t27 VDDA.t363 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X228 VOUT-.t62 two_stage_opamp_dummy_magic_24_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 GNDA.t122 GNDA.t119 GNDA.t121 GNDA.t120 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X230 two_stage_opamp_dummy_magic_24_0.VD2.t17 two_stage_opamp_dummy_magic_24_0.Vb1.t19 two_stage_opamp_dummy_magic_24_0.Y.t19 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X231 a_3690_3288.t0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t3 GNDA.t207 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X232 VOUT+.t61 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X233 bgr_11_0.NFET_GATE_10uA.t2 bgr_11_0.NFET_GATE_10uA.t1 GNDA.t10 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X234 two_stage_opamp_dummy_magic_24_0.VD1.t8 two_stage_opamp_dummy_magic_24_0.Vb1.t20 two_stage_opamp_dummy_magic_24_0.X.t1 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X235 VOUT-.t63 two_stage_opamp_dummy_magic_24_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 a_13960_3288.t1 two_stage_opamp_dummy_magic_24_0.V_tot.t3 GNDA.t303 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X237 VDDA.t180 bgr_11_0.V_TOP.t27 bgr_11_0.Vin+.t2 VDDA.t179 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X238 bgr_11_0.1st_Vout_1.t11 bgr_11_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 VOUT+.t62 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 VOUT-.t64 two_stage_opamp_dummy_magic_24_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 two_stage_opamp_dummy_magic_24_0.V_source.t7 VIN+.t1 two_stage_opamp_dummy_magic_24_0.VD2.t8 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X242 bgr_11_0.V_TOP.t28 VDDA.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X243 GNDA.t62 GNDA.t117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X244 VDDA.t22 bgr_11_0.V_mir1.t9 bgr_11_0.V_mir1.t10 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X245 VDDA.t316 VDDA.t314 bgr_11_0.NFET_GATE_10uA.t4 VDDA.t315 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X246 VOUT-.t11 VDDA.t311 VDDA.t313 VDDA.t312 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X247 bgr_11_0.1st_Vout_1.t12 bgr_11_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X248 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t1 a_3830_n594.t1 GNDA.t190 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X249 VOUT+.t63 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t13 two_stage_opamp_dummy_magic_24_0.Y.t31 VDDA.t132 GNDA.t208 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X251 VDDA.t61 bgr_11_0.1st_Vout_1.t13 bgr_11_0.V_TOP.t5 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X252 two_stage_opamp_dummy_magic_24_0.X.t9 two_stage_opamp_dummy_magic_24_0.Vb2.t19 two_stage_opamp_dummy_magic_24_0.VD3.t33 two_stage_opamp_dummy_magic_24_0.VD3.t32 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X253 VOUT-.t65 two_stage_opamp_dummy_magic_24_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 two_stage_opamp_dummy_magic_24_0.VD4.t14 two_stage_opamp_dummy_magic_24_0.Vb2.t20 two_stage_opamp_dummy_magic_24_0.Y.t8 two_stage_opamp_dummy_magic_24_0.VD4.t13 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X255 VOUT-.t66 two_stage_opamp_dummy_magic_24_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 VOUT-.t67 two_stage_opamp_dummy_magic_24_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X257 VOUT+.t64 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 VOUT+.t65 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X259 VOUT+.t66 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X260 VDDA.t123 two_stage_opamp_dummy_magic_24_0.Vb3.t20 two_stage_opamp_dummy_magic_24_0.VD3.t26 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X261 VOUT+.t67 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 two_stage_opamp_dummy_magic_24_0.VD3.t17 two_stage_opamp_dummy_magic_24_0.VD3.t15 two_stage_opamp_dummy_magic_24_0.X.t22 two_stage_opamp_dummy_magic_24_0.VD3.t16 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X263 bgr_11_0.Vin+.t1 bgr_11_0.V_TOP.t29 VDDA.t54 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X264 two_stage_opamp_dummy_magic_24_0.err_amp_out.t2 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t5 GNDA.t36 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X265 VOUT+.t68 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 VOUT+.t69 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X267 bgr_11_0.V_TOP.t30 VDDA.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X268 bgr_11_0.PFET_GATE_10uA.t7 bgr_11_0.1st_Vout_2.t14 VDDA.t207 VDDA.t206 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X269 GNDA.t116 GNDA.t114 VOUT-.t17 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X270 two_stage_opamp_dummy_magic_24_0.Vb2.t7 bgr_11_0.NFET_GATE_10uA.t10 GNDA.t234 GNDA.t233 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X271 bgr_11_0.1st_Vout_1.t14 bgr_11_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X272 VDDA.t187 bgr_11_0.V_mir1.t7 bgr_11_0.V_mir1.t8 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X273 VOUT-.t68 two_stage_opamp_dummy_magic_24_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X274 bgr_11_0.V_TOP.t31 VDDA.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X275 VOUT+.t70 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X276 VOUT-.t69 two_stage_opamp_dummy_magic_24_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 VDDA.t310 VDDA.t308 GNDA.t266 VDDA.t309 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X278 VOUT-.t70 two_stage_opamp_dummy_magic_24_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X279 VDDA.t205 bgr_11_0.1st_Vout_2.t15 bgr_11_0.PFET_GATE_10uA.t6 VDDA.t204 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X280 VOUT+.t71 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X281 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t8 two_stage_opamp_dummy_magic_24_0.X.t32 VDDA.t153 GNDA.t226 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X282 VOUT+.t72 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X283 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t7 two_stage_opamp_dummy_magic_24_0.X.t33 VDDA.t14 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X284 a_11300_30238.t0 a_11300_28630.t0 GNDA.t181 sky130_fd_pr__res_xhigh_po_0p35 l=6
X285 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t4 bgr_11_0.NFET_GATE_10uA.t11 GNDA.t248 GNDA.t247 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X286 two_stage_opamp_dummy_magic_24_0.V_source.t4 two_stage_opamp_dummy_magic_24_0.err_amp_out.t4 GNDA.t12 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X287 two_stage_opamp_dummy_magic_24_0.V_source.t32 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t21 GNDA.t250 GNDA.t249 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X288 two_stage_opamp_dummy_magic_24_0.VD1.t7 two_stage_opamp_dummy_magic_24_0.Vb1.t21 two_stage_opamp_dummy_magic_24_0.X.t18 GNDA.t212 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X289 VOUT-.t71 two_stage_opamp_dummy_magic_24_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X290 bgr_11_0.1st_Vout_2.t16 bgr_11_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X291 bgr_11_0.V_TOP.t32 VDDA.t174 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 two_stage_opamp_dummy_magic_24_0.V_source.t5 VIN+.t2 two_stage_opamp_dummy_magic_24_0.VD2.t7 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X293 VOUT-.t72 two_stage_opamp_dummy_magic_24_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X294 GNDA.t42 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t22 two_stage_opamp_dummy_magic_24_0.V_source.t16 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X295 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t2 GNDA.t111 GNDA.t113 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X296 bgr_11_0.V_p_1.t1 bgr_11_0.Vin+.t6 bgr_11_0.1st_Vout_1.t2 GNDA.t209 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.2
X297 two_stage_opamp_dummy_magic_24_0.Vb3.t2 two_stage_opamp_dummy_magic_24_0.Vb2.t21 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X298 two_stage_opamp_dummy_magic_24_0.VD4.t1 two_stage_opamp_dummy_magic_24_0.Vb2.t22 two_stage_opamp_dummy_magic_24_0.Y.t7 two_stage_opamp_dummy_magic_24_0.VD4.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X299 VDDA.t24 a_6540_22450.t14 bgr_11_0.1st_Vout_2.t0 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X300 bgr_11_0.1st_Vout_1.t15 bgr_11_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t13 two_stage_opamp_dummy_magic_24_0.Y.t32 GNDA.t222 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X302 VOUT-.t73 two_stage_opamp_dummy_magic_24_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 two_stage_opamp_dummy_magic_24_0.cap_res_X.t0 two_stage_opamp_dummy_magic_24_0.X.t19 GNDA.t213 sky130_fd_pr__res_high_po_1p41 l=1.41
X304 VOUT+.t73 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X305 VOUT-.t74 two_stage_opamp_dummy_magic_24_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X306 two_stage_opamp_dummy_magic_24_0.X.t23 two_stage_opamp_dummy_magic_24_0.Vb1.t22 two_stage_opamp_dummy_magic_24_0.VD1.t6 GNDA.t239 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X307 VOUT+.t74 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X308 VOUT-.t75 two_stage_opamp_dummy_magic_24_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 VOUT+.t75 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 bgr_11_0.1st_Vout_2.t17 bgr_11_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X311 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t12 two_stage_opamp_dummy_magic_24_0.Y.t33 VDDA.t67 GNDA.t57 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X312 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t11 two_stage_opamp_dummy_magic_24_0.Y.t34 VDDA.t117 GNDA.t195 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X313 VOUT+.t76 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 VOUT+.t77 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 GNDA.t110 GNDA.t107 GNDA.t109 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0 ps=0 w=1 l=0.15
X316 two_stage_opamp_dummy_magic_24_0.VD3.t9 two_stage_opamp_dummy_magic_24_0.Vb2.t23 two_stage_opamp_dummy_magic_24_0.X.t8 two_stage_opamp_dummy_magic_24_0.VD3.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X317 two_stage_opamp_dummy_magic_24_0.Y.t18 two_stage_opamp_dummy_magic_24_0.Vb1.t23 two_stage_opamp_dummy_magic_24_0.VD2.t18 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X318 bgr_11_0.1st_Vout_1.t16 bgr_11_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 a_5700_30088.t0 a_5820_28824.t1 GNDA.t196 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X320 VOUT+.t78 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X321 bgr_11_0.1st_Vout_2.t18 bgr_11_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X322 VDDA.t239 bgr_11_0.PFET_GATE_10uA.t15 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t1 VDDA.t238 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X323 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t5 VDDA.t305 VDDA.t307 VDDA.t306 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X324 two_stage_opamp_dummy_magic_24_0.err_amp_out.t0 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t7 two_stage_opamp_dummy_magic_24_0.V_err_p.t0 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X325 VOUT+.t79 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X326 VOUT-.t76 two_stage_opamp_dummy_magic_24_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X327 a_6540_22450.t8 a_6540_22450.t7 VDDA.t50 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X328 bgr_11_0.1st_Vout_1.t17 bgr_11_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X329 two_stage_opamp_dummy_magic_24_0.VD4.t37 two_stage_opamp_dummy_magic_24_0.Vb2.t24 two_stage_opamp_dummy_magic_24_0.Y.t6 two_stage_opamp_dummy_magic_24_0.VD4.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X330 VOUT-.t77 two_stage_opamp_dummy_magic_24_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X331 bgr_11_0.1st_Vout_2.t19 bgr_11_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X332 VDDA.t409 a_5760_7230# two_stage_opamp_dummy_magic_24_0.VD4.t35 VDDA.t408 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X333 GNDA.t62 GNDA.t106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X334 VOUT+.t80 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X335 VOUT-.t78 two_stage_opamp_dummy_magic_24_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X336 VOUT-.t15 GNDA.t103 GNDA.t105 GNDA.t104 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X337 VDDA.t304 VDDA.t302 VOUT-.t10 VDDA.t303 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X338 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t7 two_stage_opamp_dummy_magic_24_0.X.t34 GNDA.t225 VDDA.t152 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X339 VOUT+.t81 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X340 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t6 two_stage_opamp_dummy_magic_24_0.X.t35 GNDA.t0 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X341 two_stage_opamp_dummy_magic_24_0.VD3.t25 two_stage_opamp_dummy_magic_24_0.Vb3.t21 VDDA.t89 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X342 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t6 two_stage_opamp_dummy_magic_24_0.X.t36 VDDA.t151 GNDA.t224 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X343 bgr_11_0.1st_Vout_2.t20 bgr_11_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X344 VOUT+.t82 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 VOUT-.t79 two_stage_opamp_dummy_magic_24_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X346 VOUT-.t80 two_stage_opamp_dummy_magic_24_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X347 VOUT-.t81 two_stage_opamp_dummy_magic_24_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X348 VOUT-.t82 two_stage_opamp_dummy_magic_24_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X349 VOUT+.t83 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 bgr_11_0.START_UP.t2 bgr_11_0.V_TOP.t33 VDDA.t176 VDDA.t175 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X351 VOUT+.t84 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X352 VDDA.t301 VDDA.t299 VDDA.t301 VDDA.t300 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0 ps=0 w=1 l=0.15
X353 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t9 VDDA.t296 VDDA.t298 VDDA.t297 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X354 VOUT-.t83 two_stage_opamp_dummy_magic_24_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X355 bgr_11_0.1st_Vout_1.t18 bgr_11_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X356 VOUT-.t12 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t4 GNDA.t283 GNDA.t282 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X357 VDDA.t406 bgr_11_0.V_mir1.t15 bgr_11_0.1st_Vout_1.t6 VDDA.t405 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X358 VDDA.t237 bgr_11_0.PFET_GATE_10uA.t16 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t9 VDDA.t236 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X359 bgr_11_0.cap_res2.t0 bgr_11_0.PFET_GATE_10uA.t3 GNDA.t41 sky130_fd_pr__res_high_po_0p35 l=2.05
X360 two_stage_opamp_dummy_magic_24_0.V_source.t10 VIN+.t3 two_stage_opamp_dummy_magic_24_0.VD2.t6 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X361 bgr_11_0.V_TOP.t34 VDDA.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X362 VOUT-.t84 two_stage_opamp_dummy_magic_24_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 VOUT-.t85 two_stage_opamp_dummy_magic_24_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 VOUT+.t2 a_3830_n594.t0 GNDA.t174 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X365 VDDA.t403 two_stage_opamp_dummy_magic_24_0.Y.t35 VOUT+.t16 VDDA.t402 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X366 VOUT+.t85 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X367 VOUT+.t86 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X368 VOUT+.t87 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X369 VOUT+.t88 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X370 GNDA.t62 GNDA.t102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X371 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t12 two_stage_opamp_dummy_magic_24_0.Y.t36 GNDA.t304 VDDA.t410 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X372 two_stage_opamp_dummy_magic_24_0.VD3.t35 two_stage_opamp_dummy_magic_24_0.Vb2.t25 two_stage_opamp_dummy_magic_24_0.X.t7 two_stage_opamp_dummy_magic_24_0.VD3.t34 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X373 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t11 two_stage_opamp_dummy_magic_24_0.Y.t37 GNDA.t191 VDDA.t101 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X374 VOUT+.t89 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t13 bgr_11_0.PFET_GATE_10uA.t17 VDDA.t235 VDDA.t234 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X376 two_stage_opamp_dummy_magic_24_0.VD3.t24 two_stage_opamp_dummy_magic_24_0.Vb3.t22 VDDA.t114 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X377 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t10 two_stage_opamp_dummy_magic_24_0.Y.t38 VDDA.t102 GNDA.t192 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X378 VOUT+.t90 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 a_6350_30238.t0 a_6470_28630.t1 GNDA.t13 sky130_fd_pr__res_xhigh_po_0p35 l=6
X380 two_stage_opamp_dummy_magic_24_0.Y.t17 two_stage_opamp_dummy_magic_24_0.Vb1.t24 two_stage_opamp_dummy_magic_24_0.VD2.t21 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X381 VOUT-.t86 two_stage_opamp_dummy_magic_24_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 VOUT-.t87 two_stage_opamp_dummy_magic_24_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 bgr_11_0.1st_Vout_2.t2 a_6540_22450.t15 VDDA.t44 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X384 VDDA.t155 bgr_11_0.1st_Vout_1.t19 bgr_11_0.V_TOP.t7 VDDA.t154 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X385 two_stage_opamp_dummy_magic_24_0.Y.t16 two_stage_opamp_dummy_magic_24_0.Vb1.t25 two_stage_opamp_dummy_magic_24_0.VD2.t15 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X386 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t8 two_stage_opamp_dummy_magic_24_0.V_err_gate.t0 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X387 VOUT+.t91 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 VOUT-.t88 two_stage_opamp_dummy_magic_24_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X389 two_stage_opamp_dummy_magic_24_0.V_source.t19 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t23 GNDA.t164 GNDA.t163 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X390 VDDA.t30 two_stage_opamp_dummy_magic_24_0.V_err_gate.t7 two_stage_opamp_dummy_magic_24_0.V_err_p.t3 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X391 VOUT+.t92 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X392 VDDA.t32 bgr_11_0.V_mir1.t16 bgr_11_0.1st_Vout_1.t1 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X393 VOUT+.t93 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 VOUT-.t89 two_stage_opamp_dummy_magic_24_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X395 VOUT-.t90 two_stage_opamp_dummy_magic_24_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X396 VOUT+.t94 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X397 VOUT+.t95 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X398 bgr_11_0.V_TOP.t35 VDDA.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 VDDA.t373 two_stage_opamp_dummy_magic_24_0.X.t37 VOUT-.t13 VDDA.t372 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X400 VOUT+.t96 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 VDDA.t64 two_stage_opamp_dummy_magic_24_0.X.t38 VOUT-.t0 VDDA.t63 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X402 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t5 two_stage_opamp_dummy_magic_24_0.X.t39 GNDA.t210 VDDA.t133 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X403 VOUT-.t91 two_stage_opamp_dummy_magic_24_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 GNDA.t101 GNDA.t100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X405 a_12070_30088.t1 a_11950_28880.t0 GNDA.t178 sky130_fd_pr__res_xhigh_po_0p35 l=4
X406 VOUT-.t92 two_stage_opamp_dummy_magic_24_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X407 VDDA.t165 bgr_11_0.V_TOP.t36 bgr_11_0.Vin+.t0 VDDA.t164 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X408 VOUT-.t93 two_stage_opamp_dummy_magic_24_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X409 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t5 two_stage_opamp_dummy_magic_24_0.X.t40 VDDA.t170 GNDA.t242 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X410 VOUT-.t94 two_stage_opamp_dummy_magic_24_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 GNDA.t99 GNDA.t97 two_stage_opamp_dummy_magic_24_0.Vb3.t6 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X412 GNDA.t290 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t1 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t2 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X413 VOUT+.t97 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 two_stage_opamp_dummy_magic_24_0.V_source.t21 VIN-.t4 two_stage_opamp_dummy_magic_24_0.VD1.t17 GNDA.t177 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X415 VOUT+.t98 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 bgr_11_0.V_TOP.t4 bgr_11_0.START_UP.t6 bgr_11_0.Vin-.t6 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X417 a_6540_22450.t6 a_6540_22450.t5 VDDA.t366 VDDA.t365 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X418 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t0 two_stage_opamp_dummy_magic_24_0.Vb3.t1 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t1 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X419 two_stage_opamp_dummy_magic_24_0.Y.t5 two_stage_opamp_dummy_magic_24_0.Vb2.t26 two_stage_opamp_dummy_magic_24_0.VD4.t5 two_stage_opamp_dummy_magic_24_0.VD4.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X420 bgr_11_0.1st_Vout_1.t20 bgr_11_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 VDDA.t295 VDDA.t293 bgr_11_0.V_TOP.t11 VDDA.t294 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X422 VOUT+.t99 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 VOUT-.t95 two_stage_opamp_dummy_magic_24_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X424 two_stage_opamp_dummy_magic_24_0.V_source.t11 VIN+.t4 two_stage_opamp_dummy_magic_24_0.VD2.t5 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X425 GNDA.t96 GNDA.t94 two_stage_opamp_dummy_magic_24_0.Vb1.t0 GNDA.t95 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X426 VOUT+.t100 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 VDDA.t116 two_stage_opamp_dummy_magic_24_0.Y.t39 VOUT+.t4 VDDA.t115 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X428 two_stage_opamp_dummy_magic_24_0.V_source.t26 VIN-.t5 two_stage_opamp_dummy_magic_24_0.VD1.t16 GNDA.t172 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X429 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t1 bgr_11_0.V_TOP.t37 VDDA.t167 VDDA.t166 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X430 VDDA.t381 two_stage_opamp_dummy_magic_24_0.Y.t40 VOUT+.t15 VDDA.t380 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X431 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t10 two_stage_opamp_dummy_magic_24_0.Y.t41 GNDA.t22 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X432 VOUT+.t101 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 VOUT-.t96 two_stage_opamp_dummy_magic_24_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 VOUT-.t97 two_stage_opamp_dummy_magic_24_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 VOUT-.t98 two_stage_opamp_dummy_magic_24_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t9 two_stage_opamp_dummy_magic_24_0.Y.t42 VDDA.t66 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X437 VOUT+.t102 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 VOUT-.t99 two_stage_opamp_dummy_magic_24_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 VOUT+.t103 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 VOUT-.t100 two_stage_opamp_dummy_magic_24_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 VDDA.t292 VDDA.t290 two_stage_opamp_dummy_magic_24_0.Vb1.t11 VDDA.t291 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X442 VDDA.t233 bgr_11_0.PFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t8 VDDA.t232 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X443 VOUT+.t104 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X444 two_stage_opamp_dummy_magic_24_0.Y.t15 two_stage_opamp_dummy_magic_24_0.Vb1.t26 two_stage_opamp_dummy_magic_24_0.VD2.t10 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X445 VOUT+.t105 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X446 VOUT+.t106 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X447 bgr_11_0.PFET_GATE_10uA.t5 bgr_11_0.1st_Vout_2.t21 VDDA.t203 VDDA.t202 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X448 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t7 bgr_11_0.PFET_GATE_10uA.t19 VDDA.t231 VDDA.t230 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X449 bgr_11_0.1st_Vout_1.t21 bgr_11_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X450 GNDA.t93 GNDA.t91 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t2 GNDA.t92 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X451 VOUT-.t101 two_stage_opamp_dummy_magic_24_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t4 VDDA.t287 VDDA.t289 VDDA.t288 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X453 VOUT+.t107 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X454 two_stage_opamp_dummy_magic_24_0.Y.t4 two_stage_opamp_dummy_magic_24_0.Vb2.t27 two_stage_opamp_dummy_magic_24_0.VD4.t12 two_stage_opamp_dummy_magic_24_0.VD4.t11 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X455 GNDA.t201 bgr_11_0.NFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t14 GNDA.t200 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X456 VDDA.t95 bgr_11_0.V_TOP.t38 bgr_11_0.START_UP.t1 VDDA.t94 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X457 VOUT+.t108 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X458 bgr_11_0.Vin-.t2 bgr_11_0.V_TOP.t39 VDDA.t97 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X459 VOUT+.t109 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 bgr_11_0.1st_Vout_1.t22 bgr_11_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 GNDA.t4 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t24 two_stage_opamp_dummy_magic_24_0.V_source.t1 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X462 VDDA.t399 two_stage_opamp_dummy_magic_24_0.X.t41 VOUT-.t16 VDDA.t398 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X463 VDDA.t7 two_stage_opamp_dummy_magic_24_0.Vb3.t23 two_stage_opamp_dummy_magic_24_0.VD3.t23 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X464 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t4 two_stage_opamp_dummy_magic_24_0.X.t42 GNDA.t306 VDDA.t413 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X465 VOUT-.t102 two_stage_opamp_dummy_magic_24_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X466 VOUT-.t103 two_stage_opamp_dummy_magic_24_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X467 VDDA.t136 two_stage_opamp_dummy_magic_24_0.Y.t43 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t8 GNDA.t214 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X468 VOUT+.t110 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X469 two_stage_opamp_dummy_magic_24_0.V_source.t40 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t25 GNDA.t299 GNDA.t298 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X470 VOUT-.t104 two_stage_opamp_dummy_magic_24_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X471 VOUT+.t111 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t4 two_stage_opamp_dummy_magic_24_0.X.t43 VDDA.t126 GNDA.t203 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X473 VOUT+.t14 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t5 GNDA.t280 GNDA.t279 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X474 GNDA.t275 VDDA.t419 bgr_11_0.V_TOP.t9 GNDA.t274 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X475 bgr_11_0.1st_Vout_1.t23 bgr_11_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X476 VDDA.t79 two_stage_opamp_dummy_magic_24_0.Vb3.t24 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t10 VDDA.t78 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X477 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_24_0.Y.t12 GNDA.t173 sky130_fd_pr__res_high_po_1p41 l=1.41
X478 two_stage_opamp_dummy_magic_24_0.V_err_gate.t1 two_stage_opamp_dummy_magic_24_0.V_tot.t5 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.t1 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X479 GNDA.t297 bgr_11_0.NFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_24_0.V_err_gate.t2 GNDA.t296 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X480 two_stage_opamp_dummy_magic_24_0.V_source.t33 VIN-.t6 two_stage_opamp_dummy_magic_24_0.VD1.t15 GNDA.t166 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X481 VOUT-.t105 two_stage_opamp_dummy_magic_24_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 VOUT+.t112 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 bgr_11_0.V_TOP.t40 VDDA.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X484 VOUT-.t106 two_stage_opamp_dummy_magic_24_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X485 bgr_11_0.1st_Vout_2.t3 a_6540_22450.t16 VDDA.t46 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X486 VOUT+.t113 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X487 a_3810_3288.t1 two_stage_opamp_dummy_magic_24_0.V_tot.t2 GNDA.t302 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X488 VOUT+.t114 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X489 a_13840_3288.t0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t10 GNDA.t48 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X490 two_stage_opamp_dummy_magic_24_0.Vb1_2.t1 two_stage_opamp_dummy_magic_24_0.Vb1.t2 two_stage_opamp_dummy_magic_24_0.Vb1.t3 GNDA.t206 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X491 bgr_11_0.V_p_1.t2 VDDA.t420 GNDA.t273 GNDA.t272 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X492 two_stage_opamp_dummy_magic_24_0.V_source.t13 VIN+.t5 two_stage_opamp_dummy_magic_24_0.VD2.t4 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X493 VOUT-.t107 two_stage_opamp_dummy_magic_24_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X494 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t1 VIN-.t7 two_stage_opamp_dummy_magic_24_0.V_p_mir.t3 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X495 two_stage_opamp_dummy_magic_24_0.V_source.t36 VIN-.t8 two_stage_opamp_dummy_magic_24_0.VD1.t14 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X496 VDDA.t131 two_stage_opamp_dummy_magic_24_0.Y.t44 VOUT+.t6 VDDA.t130 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X497 VOUT-.t108 two_stage_opamp_dummy_magic_24_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 VDDA.t286 VDDA.t284 two_stage_opamp_dummy_magic_24_0.VD3.t20 VDDA.t285 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X499 bgr_11_0.NFET_GATE_10uA.t3 bgr_11_0.PFET_GATE_10uA.t20 VDDA.t229 VDDA.t228 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X500 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t9 two_stage_opamp_dummy_magic_24_0.Y.t45 GNDA.t243 VDDA.t173 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X501 VOUT+.t115 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X502 VOUT-.t109 two_stage_opamp_dummy_magic_24_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X503 two_stage_opamp_dummy_magic_24_0.Vb3.t4 bgr_11_0.NFET_GATE_10uA.t14 GNDA.t236 GNDA.t235 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X504 VOUT-.t110 two_stage_opamp_dummy_magic_24_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X505 VOUT+.t116 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X506 bgr_11_0.1st_Vout_2.t22 bgr_11_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X507 bgr_11_0.V_mir1.t6 bgr_11_0.V_mir1.t5 VDDA.t71 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X508 VOUT+.t117 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X509 bgr_11_0.1st_Vout_2.t4 bgr_11_0.V_CUR_REF_REG.t3 bgr_11_0.V_p_2.t0 GNDA.t228 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.2
X510 two_stage_opamp_dummy_magic_24_0.Y.t14 two_stage_opamp_dummy_magic_24_0.Vb1.t27 two_stage_opamp_dummy_magic_24_0.VD2.t13 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X511 bgr_11_0.1st_Vout_1.t24 bgr_11_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X512 bgr_11_0.1st_Vout_2.t23 bgr_11_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X513 VOUT-.t7 a_13940_n594.t1 GNDA.t240 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X514 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t13 bgr_11_0.NFET_GATE_10uA.t15 GNDA.t216 GNDA.t215 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X515 GNDA.t62 GNDA.t61 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X516 GNDA.t169 bgr_11_0.NFET_GATE_10uA.t16 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t12 GNDA.t168 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X517 VOUT-.t111 two_stage_opamp_dummy_magic_24_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X518 VOUT+.t118 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X519 GNDA.t221 two_stage_opamp_dummy_magic_24_0.Y.t46 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t8 VDDA.t146 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X520 VOUT+.t119 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X521 bgr_11_0.1st_Vout_2.t24 bgr_11_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X522 VDDA.t143 two_stage_opamp_dummy_magic_24_0.X.t44 VOUT-.t4 VDDA.t142 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X523 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t3 two_stage_opamp_dummy_magic_24_0.X.t45 GNDA.t292 VDDA.t397 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X524 VOUT-.t112 two_stage_opamp_dummy_magic_24_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 bgr_11_0.1st_Vout_1.t25 bgr_11_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X526 two_stage_opamp_dummy_magic_24_0.Vb2.t0 bgr_11_0.NFET_GATE_10uA.t17 GNDA.t38 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X527 VOUT+.t120 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 bgr_11_0.1st_Vout_2.t25 bgr_11_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X529 GNDA.t254 bgr_11_0.NFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_24_0.Vb2.t10 GNDA.t253 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X530 bgr_11_0.PFET_GATE_10uA.t4 bgr_11_0.1st_Vout_2.t26 VDDA.t201 VDDA.t200 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X531 VDDA.t26 two_stage_opamp_dummy_magic_24_0.V_err_gate.t8 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.t2 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X532 two_stage_opamp_dummy_magic_24_0.VD4.t10 two_stage_opamp_dummy_magic_24_0.Vb2.t28 two_stage_opamp_dummy_magic_24_0.Y.t3 two_stage_opamp_dummy_magic_24_0.VD4.t9 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X533 VOUT-.t113 two_stage_opamp_dummy_magic_24_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X534 VOUT+.t121 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X535 GNDA.t259 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t26 two_stage_opamp_dummy_magic_24_0.V_source.t34 GNDA.t258 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X536 bgr_11_0.1st_Vout_1.t26 bgr_11_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X537 VOUT-.t114 two_stage_opamp_dummy_magic_24_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X538 VOUT-.t115 two_stage_opamp_dummy_magic_24_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X539 two_stage_opamp_dummy_magic_24_0.V_source.t25 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t27 GNDA.t218 GNDA.t217 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X540 VOUT-.t116 two_stage_opamp_dummy_magic_24_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X541 bgr_11_0.1st_Vout_2.t27 bgr_11_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X542 two_stage_opamp_dummy_magic_24_0.Vb1_2.t0 two_stage_opamp_dummy_magic_24_0.Vb1.t8 two_stage_opamp_dummy_magic_24_0.Vb1.t9 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X543 GNDA.t62 GNDA.t63 bgr_11_0.Vin-.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X544 VOUT-.t117 two_stage_opamp_dummy_magic_24_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X545 a_3690_3288.t1 two_stage_opamp_dummy_magic_24_0.V_tot.t1 GNDA.t289 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X546 VOUT+.t122 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 VOUT+.t123 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X548 VDDA.t17 two_stage_opamp_dummy_magic_24_0.Y.t47 VOUT+.t1 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X549 two_stage_opamp_dummy_magic_24_0.V_source.t30 VIN-.t9 two_stage_opamp_dummy_magic_24_0.VD1.t13 GNDA.t212 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X550 VOUT+.t124 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X551 VDDA.t91 two_stage_opamp_dummy_magic_24_0.Vb3.t25 two_stage_opamp_dummy_magic_24_0.VD4.t19 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X552 two_stage_opamp_dummy_magic_24_0.X.t24 two_stage_opamp_dummy_magic_24_0.Vb1.t28 two_stage_opamp_dummy_magic_24_0.VD1.t5 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X553 bgr_11_0.1st_Vout_2.t6 a_6540_22450.t17 VDDA.t383 VDDA.t382 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X554 bgr_11_0.1st_Vout_1.t27 bgr_11_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X555 two_stage_opamp_dummy_magic_24_0.V_p_mir.t0 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t28 GNDA.t287 GNDA.t286 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X556 bgr_11_0.V_TOP.t1 bgr_11_0.1st_Vout_1.t28 VDDA.t20 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X557 VOUT-.t118 two_stage_opamp_dummy_magic_24_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X558 GNDA.t278 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t6 VOUT+.t13 GNDA.t277 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X559 VOUT+.t125 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X560 VOUT-.t119 two_stage_opamp_dummy_magic_24_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 bgr_11_0.1st_Vout_1.t3 bgr_11_0.V_mir1.t17 VDDA.t185 VDDA.t184 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X562 VOUT-.t120 two_stage_opamp_dummy_magic_24_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X563 two_stage_opamp_dummy_magic_24_0.Y.t1 GNDA.t88 GNDA.t90 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X564 two_stage_opamp_dummy_magic_24_0.VD1.t12 VIN-.t10 two_stage_opamp_dummy_magic_24_0.V_source.t29 GNDA.t239 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X565 two_stage_opamp_dummy_magic_24_0.VD4.t29 two_stage_opamp_dummy_magic_24_0.VD4.t27 two_stage_opamp_dummy_magic_24_0.Y.t23 two_stage_opamp_dummy_magic_24_0.VD4.t28 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X566 GNDA.t276 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t29 two_stage_opamp_dummy_magic_24_0.V_source.t35 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X567 VDDA.t283 VDDA.t281 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t4 VDDA.t282 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X568 VOUT-.t121 two_stage_opamp_dummy_magic_24_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X569 VOUT-.t122 two_stage_opamp_dummy_magic_24_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 bgr_11_0.PFET_GATE_10uA.t0 VDDA.t421 GNDA.t271 GNDA.t270 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X571 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t0 bgr_11_0.PFET_GATE_10uA.t21 VDDA.t227 VDDA.t226 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X572 two_stage_opamp_dummy_magic_24_0.X.t0 two_stage_opamp_dummy_magic_24_0.Vb1.t29 two_stage_opamp_dummy_magic_24_0.VD1.t4 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X573 VOUT-.t123 two_stage_opamp_dummy_magic_24_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X574 VDDA.t280 VDDA.t277 VDDA.t279 VDDA.t278 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0 ps=0 w=1.8 l=0.2
X575 two_stage_opamp_dummy_magic_24_0.VD2.t3 VIN+.t6 two_stage_opamp_dummy_magic_24_0.V_source.t12 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X576 bgr_11_0.V_TOP.t41 VDDA.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X577 two_stage_opamp_dummy_magic_24_0.VD3.t22 two_stage_opamp_dummy_magic_24_0.Vb3.t26 VDDA.t93 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X578 VDDA.t276 VDDA.t274 bgr_11_0.PFET_GATE_10uA.t2 VDDA.t275 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X579 VDDA.t162 bgr_11_0.V_TOP.t42 bgr_11_0.START_UP.t0 VDDA.t161 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X580 VOUT+.t0 two_stage_opamp_dummy_magic_24_0.Y.t48 VDDA.t9 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X581 VDDA.t412 two_stage_opamp_dummy_magic_24_0.X.t46 VOUT-.t18 VDDA.t411 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X582 VDDA.t145 two_stage_opamp_dummy_magic_24_0.Y.t49 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t7 GNDA.t220 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X583 VOUT+.t126 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X584 VOUT-.t124 two_stage_opamp_dummy_magic_24_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X585 a_6540_22450.t4 a_6540_22450.t3 VDDA.t83 VDDA.t82 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X586 VDDA.t273 VDDA.t271 VDDA.t273 VDDA.t272 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X587 VOUT-.t125 two_stage_opamp_dummy_magic_24_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X588 bgr_11_0.V_TOP.t43 VDDA.t163 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X589 VOUT-.t126 two_stage_opamp_dummy_magic_24_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X590 two_stage_opamp_dummy_magic_24_0.X.t6 two_stage_opamp_dummy_magic_24_0.Vb2.t29 two_stage_opamp_dummy_magic_24_0.VD3.t11 two_stage_opamp_dummy_magic_24_0.VD3.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X591 a_11420_30238.t0 a_11300_28630.t1 GNDA.t182 sky130_fd_pr__res_xhigh_po_0p35 l=6
X592 a_3810_3288.t0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t16 GNDA.t301 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X593 GNDA.t87 GNDA.t85 two_stage_opamp_dummy_magic_24_0.err_amp_out.t1 GNDA.t86 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X594 VOUT+.t127 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X595 a_13960_3288.t0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t10 GNDA.t43 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X596 VOUT-.t127 two_stage_opamp_dummy_magic_24_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X597 VDDA.t225 bgr_11_0.PFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t6 VDDA.t224 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X598 VOUT+.t128 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X599 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t5 bgr_11_0.PFET_GATE_10uA.t23 VDDA.t223 VDDA.t222 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X600 bgr_11_0.V_TOP.t44 VDDA.t387 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X601 VOUT+.t129 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X602 VOUT+.t130 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X603 VOUT-.t128 two_stage_opamp_dummy_magic_24_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X604 two_stage_opamp_dummy_magic_24_0.Vb2.t1 two_stage_opamp_dummy_magic_24_0.Vb2_2.t3 two_stage_opamp_dummy_magic_24_0.Vb2_2.t5 two_stage_opamp_dummy_magic_24_0.Vb2_2.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X605 bgr_11_0.1st_Vout_1.t4 bgr_11_0.V_mir1.t18 VDDA.t195 VDDA.t194 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X606 VOUT+.t131 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X607 VOUT+.t132 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X608 bgr_11_0.V_mir1.t0 bgr_11_0.Vin-.t8 bgr_11_0.V_p_1.t0 GNDA.t255 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.2
X609 two_stage_opamp_dummy_magic_24_0.X.t17 two_stage_opamp_dummy_magic_24_0.Vb1.t30 two_stage_opamp_dummy_magic_24_0.VD1.t3 GNDA.t205 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X610 VOUT-.t129 two_stage_opamp_dummy_magic_24_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X611 GNDA.t84 GNDA.t82 two_stage_opamp_dummy_magic_24_0.V_source.t23 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X612 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t12 bgr_11_0.PFET_GATE_10uA.t24 VDDA.t221 VDDA.t220 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X613 GNDA.t8 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t30 two_stage_opamp_dummy_magic_24_0.V_source.t3 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X614 VDDA.t219 bgr_11_0.PFET_GATE_10uA.t25 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t11 VDDA.t218 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X615 VOUT-.t130 two_stage_opamp_dummy_magic_24_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X616 VOUT-.t131 two_stage_opamp_dummy_magic_24_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X617 VOUT-.t132 two_stage_opamp_dummy_magic_24_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X618 VDDA.t270 VDDA.t268 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t15 VDDA.t269 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X619 VOUT-.t133 two_stage_opamp_dummy_magic_24_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X620 VDDA.t125 two_stage_opamp_dummy_magic_24_0.X.t47 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t3 GNDA.t202 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X621 VOUT+.t133 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X622 VDDA.t267 VDDA.t265 two_stage_opamp_dummy_magic_24_0.Vb2_2.t9 VDDA.t266 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.36 ps=2.2 w=1.8 l=0.2
X623 VOUT+.t134 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X624 VOUT-.t9 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t7 GNDA.t261 GNDA.t260 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X625 two_stage_opamp_dummy_magic_24_0.V_source.t24 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t31 GNDA.t199 GNDA.t86 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X626 VOUT+.t135 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X627 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t0 bgr_11_0.V_TOP.t45 VDDA.t389 VDDA.t388 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X628 two_stage_opamp_dummy_magic_24_0.X.t20 two_stage_opamp_dummy_magic_24_0.Vb1.t31 two_stage_opamp_dummy_magic_24_0.VD1.t2 GNDA.t227 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X629 bgr_11_0.V_TOP.t46 VDDA.t394 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X630 GNDA.t180 a_5820_28824.t0 GNDA.t179 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X631 bgr_11_0.V_TOP.t3 bgr_11_0.1st_Vout_1.t29 VDDA.t48 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X632 two_stage_opamp_dummy_magic_24_0.VD2.t2 VIN+.t7 two_stage_opamp_dummy_magic_24_0.V_source.t8 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X633 VOUT+.t136 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X634 two_stage_opamp_dummy_magic_24_0.V_p_mir.t2 VIN+.t8 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t0 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X635 two_stage_opamp_dummy_magic_24_0.VD2.t1 VIN+.t9 two_stage_opamp_dummy_magic_24_0.V_source.t14 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X636 VOUT+.t137 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X637 two_stage_opamp_dummy_magic_24_0.VD4.t6 a_4440_7230# VDDA.t73 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X638 GNDA.t294 two_stage_opamp_dummy_magic_24_0.Y.t50 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t7 VDDA.t401 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X639 VOUT-.t134 two_stage_opamp_dummy_magic_24_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X640 GNDA.t81 GNDA.t79 two_stage_opamp_dummy_magic_24_0.X.t3 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X641 VOUT-.t135 two_stage_opamp_dummy_magic_24_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X642 VOUT-.t136 two_stage_opamp_dummy_magic_24_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X643 bgr_11_0.V_TOP.t2 bgr_11_0.1st_Vout_1.t30 VDDA.t34 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X644 VOUT-.t137 two_stage_opamp_dummy_magic_24_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X645 VOUT+.t138 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X646 VOUT-.t138 two_stage_opamp_dummy_magic_24_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X647 bgr_11_0.1st_Vout_2.t28 bgr_11_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X648 VDDA.t414 two_stage_opamp_dummy_magic_24_0.Y.t51 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t6 GNDA.t308 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X649 VOUT+.t139 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X650 VDDA.t264 VDDA.t262 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t5 VDDA.t263 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X651 two_stage_opamp_dummy_magic_24_0.Y.t2 two_stage_opamp_dummy_magic_24_0.Vb2.t30 two_stage_opamp_dummy_magic_24_0.VD4.t16 two_stage_opamp_dummy_magic_24_0.VD4.t15 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X652 VOUT+.t140 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X653 two_stage_opamp_dummy_magic_24_0.Vb3.t0 bgr_11_0.NFET_GATE_10uA.t19 GNDA.t40 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X654 GNDA.t78 GNDA.t76 two_stage_opamp_dummy_magic_24_0.Y.t0 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X655 VOUT-.t139 two_stage_opamp_dummy_magic_24_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X656 bgr_11_0.1st_Vout_1.t31 bgr_11_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X657 VDDA.t261 VDDA.t259 two_stage_opamp_dummy_magic_24_0.err_amp_out.t3 VDDA.t260 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X658 VOUT+.t141 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X659 VOUT-.t140 two_stage_opamp_dummy_magic_24_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X660 bgr_11_0.Vin-.t5 bgr_11_0.START_UP.t7 bgr_11_0.V_TOP.t0 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X661 VOUT-.t141 two_stage_opamp_dummy_magic_24_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X662 VOUT+.t142 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X663 VOUT+.t143 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X664 VOUT-.t142 two_stage_opamp_dummy_magic_24_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X665 bgr_11_0.V_mir1.t4 bgr_11_0.V_mir1.t3 VDDA.t191 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X666 two_stage_opamp_dummy_magic_24_0.VD4.t18 two_stage_opamp_dummy_magic_24_0.Vb3.t27 VDDA.t379 VDDA.t378 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X667 VOUT+.t144 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X668 bgr_11_0.V_p_2.t1 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t9 a_6540_22450.t0 GNDA.t281 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.2
X669 VOUT-.t143 two_stage_opamp_dummy_magic_24_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X670 VOUT-.t144 two_stage_opamp_dummy_magic_24_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X671 VOUT-.t145 two_stage_opamp_dummy_magic_24_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X672 bgr_11_0.V_TOP.t10 VDDA.t256 VDDA.t258 VDDA.t257 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X673 VOUT-.t146 two_stage_opamp_dummy_magic_24_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X674 VOUT+.t145 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X675 GNDA.t291 two_stage_opamp_dummy_magic_24_0.X.t48 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t2 VDDA.t396 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X676 bgr_11_0.V_TOP.t47 VDDA.t395 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X677 VDDA.t40 bgr_11_0.V_TOP.t48 bgr_11_0.Vin-.t1 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X678 VOUT+.t146 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X679 VDDA.t407 two_stage_opamp_dummy_magic_24_0.X.t49 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t2 GNDA.t300 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X680 VOUT+.t147 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X681 VOUT-.t147 two_stage_opamp_dummy_magic_24_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X682 two_stage_opamp_dummy_magic_24_0.Vb1.t10 bgr_11_0.PFET_GATE_10uA.t26 VDDA.t217 VDDA.t216 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X683 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t4 bgr_11_0.PFET_GATE_10uA.t27 VDDA.t215 VDDA.t214 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X684 VDDA.t100 two_stage_opamp_dummy_magic_24_0.X.t50 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t1 GNDA.t189 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X685 VOUT-.t148 two_stage_opamp_dummy_magic_24_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X686 GNDA.t14 a_6470_28630.t0 GNDA.t13 sky130_fd_pr__res_xhigh_po_0p35 l=6
X687 VOUT+.t148 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X688 VOUT-.t149 two_stage_opamp_dummy_magic_24_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X689 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t0 bgr_11_0.NFET_GATE_10uA.t20 GNDA.t45 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X690 two_stage_opamp_dummy_magic_24_0.Vb2_2.t2 two_stage_opamp_dummy_magic_24_0.Vb2.t31 VDDA.t28 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.36 ps=2.2 w=1.8 l=0.2
X691 two_stage_opamp_dummy_magic_24_0.X.t2 GNDA.t73 GNDA.t75 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X692 VDDA.t38 a_6540_22450.t18 bgr_11_0.1st_Vout_2.t1 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X693 bgr_11_0.1st_Vout_2.t29 bgr_11_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X694 GNDA.t245 bgr_11_0.NFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_24_0.Vb2.t8 GNDA.t244 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X695 two_stage_opamp_dummy_magic_24_0.VD2.t0 VIN+.t10 two_stage_opamp_dummy_magic_24_0.V_source.t6 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X696 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t11 GNDA.t70 GNDA.t72 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X697 GNDA.t265 VDDA.t422 bgr_11_0.V_p_2.t2 GNDA.t264 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X698 bgr_11_0.V_mir1.t2 bgr_11_0.V_mir1.t1 VDDA.t157 VDDA.t156 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X699 VOUT+.t5 two_stage_opamp_dummy_magic_24_0.Y.t52 VDDA.t129 VDDA.t128 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X700 VOUT+.t149 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X701 bgr_11_0.PFET_GATE_10uA.t1 VDDA.t253 VDDA.t255 VDDA.t254 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X702 two_stage_opamp_dummy_magic_24_0.X.t21 two_stage_opamp_dummy_magic_24_0.VD3.t12 two_stage_opamp_dummy_magic_24_0.VD3.t14 two_stage_opamp_dummy_magic_24_0.VD3.t13 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X703 GNDA.t219 two_stage_opamp_dummy_magic_24_0.Y.t53 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t6 VDDA.t144 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X704 VDDA.t85 GNDA.t67 GNDA.t69 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X705 two_stage_opamp_dummy_magic_24_0.VD3.t19 two_stage_opamp_dummy_magic_24_0.Vb2.t32 two_stage_opamp_dummy_magic_24_0.X.t5 two_stage_opamp_dummy_magic_24_0.VD3.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X706 VDDA.t400 two_stage_opamp_dummy_magic_24_0.Y.t54 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t5 GNDA.t293 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X707 a_12070_30088.t0 bgr_11_0.V_CUR_REF_REG.t0 GNDA.t19 sky130_fd_pr__res_xhigh_po_0p35 l=4
X708 GNDA.t232 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t8 VOUT-.t5 GNDA.t231 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X709 two_stage_opamp_dummy_magic_24_0.VD2.t16 two_stage_opamp_dummy_magic_24_0.Vb1.t32 two_stage_opamp_dummy_magic_24_0.Y.t13 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X710 two_stage_opamp_dummy_magic_24_0.VD4.t17 two_stage_opamp_dummy_magic_24_0.Vb3.t28 VDDA.t377 VDDA.t376 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X711 VOUT+.t150 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X712 bgr_11_0.1st_Vout_2.t30 bgr_11_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X713 GNDA.t66 GNDA.t64 bgr_11_0.NFET_GATE_10uA.t0 GNDA.t65 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X714 bgr_11_0.Vin-.t0 bgr_11_0.V_TOP.t49 VDDA.t42 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X715 VOUT-.t150 two_stage_opamp_dummy_magic_24_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X716 VOUT+.t151 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X717 two_stage_opamp_dummy_magic_24_0.V_err_p.t2 two_stage_opamp_dummy_magic_24_0.V_err_gate.t9 VDDA.t193 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X718 two_stage_opamp_dummy_magic_24_0.Vb2_2.t1 two_stage_opamp_dummy_magic_24_0.Vb2.t4 two_stage_opamp_dummy_magic_24_0.Vb2.t5 two_stage_opamp_dummy_magic_24_0.Vb2_2.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X719 VOUT-.t151 two_stage_opamp_dummy_magic_24_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X720 VOUT+.t152 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X721 VDDA.t106 a_6540_22450.t1 a_6540_22450.t2 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X722 VOUT-.t152 two_stage_opamp_dummy_magic_24_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X723 VOUT-.t153 two_stage_opamp_dummy_magic_24_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X724 VOUT+.t153 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X725 bgr_11_0.1st_Vout_2.t31 bgr_11_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X726 VOUT+.t154 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X727 bgr_11_0.V_CUR_REF_REG.t2 VDDA.t250 VDDA.t252 VDDA.t251 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X728 VOUT+.t155 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X729 two_stage_opamp_dummy_magic_24_0.Vb3.t5 GNDA.t58 GNDA.t60 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X730 VOUT-.t1 two_stage_opamp_dummy_magic_24_0.X.t51 VDDA.t110 VDDA.t109 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X731 VOUT+.t156 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X732 GNDA.t238 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t9 VOUT-.t6 GNDA.t237 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X733 VDDA.t213 bgr_11_0.PFET_GATE_10uA.t28 bgr_11_0.V_CUR_REF_REG.t1 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X734 GNDA.t288 two_stage_opamp_dummy_magic_24_0.X.t52 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t1 VDDA.t367 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X735 GNDA.t311 bgr_11_0.NFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_24_0.Vb3.t7 GNDA.t310 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X736 VOUT-.t154 two_stage_opamp_dummy_magic_24_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X737 bgr_11_0.1st_Vout_1.t32 bgr_11_0.cap_res1.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X738 GNDA.t16 two_stage_opamp_dummy_magic_24_0.X.t53 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t0 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X739 VDDA.t62 two_stage_opamp_dummy_magic_24_0.X.t54 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t0 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X740 a_5700_30088.t1 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t4 GNDA.t211 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X741 VOUT-.t155 two_stage_opamp_dummy_magic_24_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X742 bgr_11_0.1st_Vout_2.t32 bgr_11_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X743 VOUT-.t156 two_stage_opamp_dummy_magic_24_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 bgr_11_0.1st_Vout_2.n9 bgr_11_0.1st_Vout_2.t15 362.341
R1 bgr_11_0.1st_Vout_2.n7 bgr_11_0.1st_Vout_2.t14 355.094
R2 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.n10 302.183
R3 bgr_11_0.1st_Vout_2.n7 bgr_11_0.1st_Vout_2.n6 302.183
R4 bgr_11_0.1st_Vout_2.n12 bgr_11_0.1st_Vout_2.n5 297.683
R5 bgr_11_0.1st_Vout_2.n11 bgr_11_0.1st_Vout_2.t26 194.809
R6 bgr_11_0.1st_Vout_2.n11 bgr_11_0.1st_Vout_2.t9 194.809
R7 bgr_11_0.1st_Vout_2.n8 bgr_11_0.1st_Vout_2.t21 194.809
R8 bgr_11_0.1st_Vout_2.n8 bgr_11_0.1st_Vout_2.t7 194.809
R9 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.n11 166.03
R10 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.n8 166.03
R11 bgr_11_0.1st_Vout_2.t4 bgr_11_0.1st_Vout_2.n12 49.5021
R12 bgr_11_0.1st_Vout_2.n10 bgr_11_0.1st_Vout_2.t0 39.4005
R13 bgr_11_0.1st_Vout_2.n10 bgr_11_0.1st_Vout_2.t3 39.4005
R14 bgr_11_0.1st_Vout_2.n6 bgr_11_0.1st_Vout_2.t1 39.4005
R15 bgr_11_0.1st_Vout_2.n6 bgr_11_0.1st_Vout_2.t2 39.4005
R16 bgr_11_0.1st_Vout_2.n5 bgr_11_0.1st_Vout_2.t5 39.4005
R17 bgr_11_0.1st_Vout_2.n5 bgr_11_0.1st_Vout_2.t6 39.4005
R18 bgr_11_0.1st_Vout_2.n9 bgr_11_0.1st_Vout_2.n0 35.7185
R19 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t32 4.8295
R20 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t12 4.8295
R21 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t13 4.8295
R22 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t19 4.8295
R23 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t30 4.8295
R24 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t11 4.8295
R25 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t23 4.8295
R26 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t28 4.8295
R27 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t8 4.8295
R28 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t27 4.5005
R29 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t20 4.5005
R30 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t31 4.5005
R31 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t25 4.5005
R32 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t24 4.5005
R33 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t18 4.5005
R34 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t17 4.5005
R35 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t10 4.5005
R36 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t29 4.5005
R37 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t22 4.5005
R38 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t16 4.5005
R39 bgr_11_0.1st_Vout_2.n12 bgr_11_0.1st_Vout_2.n3 4.5005
R40 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.n9 2.90725
R41 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.n2 2.2095
R42 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.n4 1.1255
R43 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.n7 1.1255
R44 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.n1 0.8935
R45 bgr_11_0.PFET_GATE_10uA.n14 bgr_11_0.PFET_GATE_10uA.t26 758.64
R46 bgr_11_0.PFET_GATE_10uA.n4 bgr_11_0.PFET_GATE_10uA.n0 510.991
R47 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n25 509.226
R48 bgr_11_0.PFET_GATE_10uA.n22 bgr_11_0.PFET_GATE_10uA.t22 369.534
R49 bgr_11_0.PFET_GATE_10uA.n19 bgr_11_0.PFET_GATE_10uA.t27 369.534
R50 bgr_11_0.PFET_GATE_10uA.n16 bgr_11_0.PFET_GATE_10uA.t11 369.534
R51 bgr_11_0.PFET_GATE_10uA.n15 bgr_11_0.PFET_GATE_10uA.t10 369.534
R52 bgr_11_0.PFET_GATE_10uA.n2 bgr_11_0.PFET_GATE_10uA.t25 369.534
R53 bgr_11_0.PFET_GATE_10uA.n1 bgr_11_0.PFET_GATE_10uA.t24 369.534
R54 bgr_11_0.PFET_GATE_10uA.n12 bgr_11_0.PFET_GATE_10uA.n11 301.933
R55 bgr_11_0.PFET_GATE_10uA.n10 bgr_11_0.PFET_GATE_10uA.n9 301.933
R56 bgr_11_0.PFET_GATE_10uA.n8 bgr_11_0.PFET_GATE_10uA.n7 301.933
R57 bgr_11_0.PFET_GATE_10uA.n6 bgr_11_0.PFET_GATE_10uA.n5 301.933
R58 bgr_11_0.PFET_GATE_10uA.n0 bgr_11_0.PFET_GATE_10uA.t20 249.034
R59 bgr_11_0.PFET_GATE_10uA.n0 bgr_11_0.PFET_GATE_10uA.t28 249.034
R60 bgr_11_0.PFET_GATE_10uA.n22 bgr_11_0.PFET_GATE_10uA.t12 192.8
R61 bgr_11_0.PFET_GATE_10uA.n23 bgr_11_0.PFET_GATE_10uA.t16 192.8
R62 bgr_11_0.PFET_GATE_10uA.n24 bgr_11_0.PFET_GATE_10uA.t23 192.8
R63 bgr_11_0.PFET_GATE_10uA.n21 bgr_11_0.PFET_GATE_10uA.t14 192.8
R64 bgr_11_0.PFET_GATE_10uA.n20 bgr_11_0.PFET_GATE_10uA.t19 192.8
R65 bgr_11_0.PFET_GATE_10uA.n19 bgr_11_0.PFET_GATE_10uA.t18 192.8
R66 bgr_11_0.PFET_GATE_10uA.n16 bgr_11_0.PFET_GATE_10uA.t21 192.8
R67 bgr_11_0.PFET_GATE_10uA.n15 bgr_11_0.PFET_GATE_10uA.t15 192.8
R68 bgr_11_0.PFET_GATE_10uA.n2 bgr_11_0.PFET_GATE_10uA.t17 192.8
R69 bgr_11_0.PFET_GATE_10uA.n1 bgr_11_0.PFET_GATE_10uA.t13 192.8
R70 bgr_11_0.PFET_GATE_10uA.n21 bgr_11_0.PFET_GATE_10uA.n20 176.733
R71 bgr_11_0.PFET_GATE_10uA.n20 bgr_11_0.PFET_GATE_10uA.n19 176.733
R72 bgr_11_0.PFET_GATE_10uA.n23 bgr_11_0.PFET_GATE_10uA.n22 176.733
R73 bgr_11_0.PFET_GATE_10uA.n24 bgr_11_0.PFET_GATE_10uA.n23 176.733
R74 bgr_11_0.PFET_GATE_10uA.n18 bgr_11_0.PFET_GATE_10uA.n17 166.541
R75 bgr_11_0.PFET_GATE_10uA.n4 bgr_11_0.PFET_GATE_10uA.n3 166.343
R76 bgr_11_0.PFET_GATE_10uA.n13 bgr_11_0.PFET_GATE_10uA.t3 119.118
R77 bgr_11_0.PFET_GATE_10uA.n6 bgr_11_0.PFET_GATE_10uA.t0 104.474
R78 bgr_11_0.PFET_GATE_10uA.n17 bgr_11_0.PFET_GATE_10uA.n16 56.2338
R79 bgr_11_0.PFET_GATE_10uA.n17 bgr_11_0.PFET_GATE_10uA.n15 56.2338
R80 bgr_11_0.PFET_GATE_10uA.n3 bgr_11_0.PFET_GATE_10uA.n2 56.2338
R81 bgr_11_0.PFET_GATE_10uA.n3 bgr_11_0.PFET_GATE_10uA.n1 56.2338
R82 bgr_11_0.PFET_GATE_10uA.n25 bgr_11_0.PFET_GATE_10uA.n21 56.2338
R83 bgr_11_0.PFET_GATE_10uA.n25 bgr_11_0.PFET_GATE_10uA.n24 56.2338
R84 bgr_11_0.PFET_GATE_10uA.n11 bgr_11_0.PFET_GATE_10uA.t6 39.4005
R85 bgr_11_0.PFET_GATE_10uA.n11 bgr_11_0.PFET_GATE_10uA.t1 39.4005
R86 bgr_11_0.PFET_GATE_10uA.n9 bgr_11_0.PFET_GATE_10uA.t8 39.4005
R87 bgr_11_0.PFET_GATE_10uA.n9 bgr_11_0.PFET_GATE_10uA.t4 39.4005
R88 bgr_11_0.PFET_GATE_10uA.n7 bgr_11_0.PFET_GATE_10uA.t9 39.4005
R89 bgr_11_0.PFET_GATE_10uA.n7 bgr_11_0.PFET_GATE_10uA.t5 39.4005
R90 bgr_11_0.PFET_GATE_10uA.n5 bgr_11_0.PFET_GATE_10uA.t2 39.4005
R91 bgr_11_0.PFET_GATE_10uA.n5 bgr_11_0.PFET_GATE_10uA.t7 39.4005
R92 bgr_11_0.PFET_GATE_10uA.n18 bgr_11_0.PFET_GATE_10uA.n14 10.5161
R93 bgr_11_0.PFET_GATE_10uA.n13 bgr_11_0.PFET_GATE_10uA.n12 6.15675
R94 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n4 2.28175
R95 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n18 2.28175
R96 bgr_11_0.PFET_GATE_10uA.n14 bgr_11_0.PFET_GATE_10uA.n13 1.40675
R97 bgr_11_0.PFET_GATE_10uA.n8 bgr_11_0.PFET_GATE_10uA.n6 1.1255
R98 bgr_11_0.PFET_GATE_10uA.n10 bgr_11_0.PFET_GATE_10uA.n8 1.1255
R99 bgr_11_0.PFET_GATE_10uA.n12 bgr_11_0.PFET_GATE_10uA.n10 1.1255
R100 VDDA.n404 VDDA.t331 1231.74
R101 VDDA.n401 VDDA.t346 1231.74
R102 VDDA.n2301 VDDA.t302 1231.74
R103 VDDA.n2304 VDDA.t311 1231.74
R104 VDDA.n2360 VDDA.t259 826.801
R105 VDDA.n2392 VDDA.t355 826.801
R106 VDDA.n2366 VDDA.t349 826.801
R107 VDDA.n448 VDDA.t287 826.801
R108 VDDA.t276 VDDA.n1973 708.125
R109 VDDA.n1996 VDDA.t276 708.125
R110 VDDA.n1993 VDDA.t255 708.125
R111 VDDA.t255 VDDA.n1974 708.125
R112 VDDA.t319 VDDA.n1953 708.125
R113 VDDA.n2006 VDDA.t319 708.125
R114 VDDA.n2003 VDDA.t258 708.125
R115 VDDA.t258 VDDA.n1954 708.125
R116 VDDA.t335 VDDA.n2083 676.966
R117 VDDA.n380 VDDA.t271 661.375
R118 VDDA.n383 VDDA.t296 661.375
R119 VDDA.n1995 VDDA.t275 657.76
R120 VDDA.n2005 VDDA.t318 657.76
R121 VDDA.n2084 VDDA.t294 643.038
R122 VDDA.t282 VDDA.n2117 643.037
R123 VDDA.n2118 VDDA.t306 643.037
R124 VDDA.t269 VDDA.n2102 643.037
R125 VDDA.n2103 VDDA.t341 643.037
R126 VDDA.n2112 VDDA.t321 642.992
R127 VDDA.t300 VDDA.n2111 642.992
R128 VDDA.n2097 VDDA.t251 642.992
R129 VDDA.t315 VDDA.n2096 642.992
R130 VDDA.n1768 VDDA.t324 605.143
R131 VDDA.n1789 VDDA.t290 589.076
R132 VDDA.n2328 VDDA.t308 589.076
R133 VDDA.n2331 VDDA.t328 589.076
R134 VDDA.n435 VDDA.t343 589.076
R135 VDDA.n432 VDDA.t358 589.076
R136 VDDA.n2035 VDDA.n2033 587.407
R137 VDDA.n2039 VDDA.n2036 587.407
R138 VDDA.n2065 VDDA.n2064 587.407
R139 VDDA.n2060 VDDA.n2026 587.407
R140 VDDA.n2064 VDDA.n2063 585
R141 VDDA.n2062 VDDA.n2060 585
R142 VDDA.n2046 VDDA.n2035 585
R143 VDDA.n2043 VDDA.n2036 585
R144 VDDA.n2391 VDDA.n442 585
R145 VDDA.n2379 VDDA.n2378 585
R146 VDDA.n2376 VDDA.n2375 585
R147 VDDA.n2359 VDDA.n2358 585
R148 VDDA.t254 VDDA.n1994 540.818
R149 VDDA.t257 VDDA.n2004 540.818
R150 VDDA.n1779 VDDA.t292 464.281
R151 VDDA.t292 VDDA.n1395 464.281
R152 VDDA.n1774 VDDA.t327 464.281
R153 VDDA.t327 VDDA.n1773 464.281
R154 VDDA.n376 VDDA.t265 456.526
R155 VDDA.n373 VDDA.t277 456.526
R156 VDDA.n2105 VDDA.t299 441.2
R157 VDDA.n2113 VDDA.t320 441.2
R158 VDDA.n2094 VDDA.t314 441.2
R159 VDDA.n2098 VDDA.t250 441.2
R160 VDDA.n2085 VDDA.t293 413.084
R161 VDDA.n2082 VDDA.t334 413.084
R162 VDDA.n2114 VDDA.t281 409.067
R163 VDDA.n2119 VDDA.t305 409.067
R164 VDDA.t275 VDDA.t206 407.144
R165 VDDA.t206 VDDA.t37 407.144
R166 VDDA.t37 VDDA.t43 407.144
R167 VDDA.t43 VDDA.t158 407.144
R168 VDDA.t158 VDDA.t49 407.144
R169 VDDA.t49 VDDA.t210 407.144
R170 VDDA.t210 VDDA.t202 407.144
R171 VDDA.t202 VDDA.t168 407.144
R172 VDDA.t168 VDDA.t382 407.144
R173 VDDA.t382 VDDA.t105 407.144
R174 VDDA.t105 VDDA.t365 407.144
R175 VDDA.t365 VDDA.t208 407.144
R176 VDDA.t208 VDDA.t200 407.144
R177 VDDA.t200 VDDA.t23 407.144
R178 VDDA.t23 VDDA.t45 407.144
R179 VDDA.t45 VDDA.t390 407.144
R180 VDDA.t390 VDDA.t82 407.144
R181 VDDA.t82 VDDA.t204 407.144
R182 VDDA.t204 VDDA.t254 407.144
R183 VDDA.t318 VDDA.t47 407.144
R184 VDDA.t47 VDDA.t198 407.144
R185 VDDA.t198 VDDA.t70 407.144
R186 VDDA.t70 VDDA.t196 407.144
R187 VDDA.t196 VDDA.t194 407.144
R188 VDDA.t194 VDDA.t154 407.144
R189 VDDA.t154 VDDA.t19 407.144
R190 VDDA.t19 VDDA.t21 407.144
R191 VDDA.t21 VDDA.t190 407.144
R192 VDDA.t190 VDDA.t405 407.144
R193 VDDA.t405 VDDA.t10 407.144
R194 VDDA.t10 VDDA.t188 407.144
R195 VDDA.t188 VDDA.t33 407.144
R196 VDDA.t33 VDDA.t186 407.144
R197 VDDA.t186 VDDA.t156 407.144
R198 VDDA.t156 VDDA.t31 407.144
R199 VDDA.t31 VDDA.t184 407.144
R200 VDDA.t184 VDDA.t60 407.144
R201 VDDA.t60 VDDA.t257 407.144
R202 VDDA.n375 VDDA.t266 397.784
R203 VDDA.t278 VDDA.n374 397.784
R204 VDDA.n2099 VDDA.t268 390.322
R205 VDDA.n2104 VDDA.t340 390.322
R206 VDDA.t248 VDDA.t282 373.214
R207 VDDA.t238 VDDA.t248 373.214
R208 VDDA.t226 VDDA.t238 373.214
R209 VDDA.t246 VDDA.t226 373.214
R210 VDDA.t306 VDDA.t246 373.214
R211 VDDA.t224 VDDA.t300 373.214
R212 VDDA.t244 VDDA.t224 373.214
R213 VDDA.t236 VDDA.t244 373.214
R214 VDDA.t222 VDDA.t236 373.214
R215 VDDA.t240 VDDA.t222 373.214
R216 VDDA.t230 VDDA.t240 373.214
R217 VDDA.t232 VDDA.t230 373.214
R218 VDDA.t214 VDDA.t232 373.214
R219 VDDA.t321 VDDA.t214 373.214
R220 VDDA.t220 VDDA.t269 373.214
R221 VDDA.t242 VDDA.t220 373.214
R222 VDDA.t234 VDDA.t242 373.214
R223 VDDA.t218 VDDA.t234 373.214
R224 VDDA.t341 VDDA.t218 373.214
R225 VDDA.t228 VDDA.t315 373.214
R226 VDDA.t212 VDDA.t228 373.214
R227 VDDA.t251 VDDA.t212 373.214
R228 VDDA.t294 VDDA.t51 373.214
R229 VDDA.t51 VDDA.t0 373.214
R230 VDDA.t0 VDDA.t335 373.214
R231 VDDA.n1998 VDDA.t274 370.168
R232 VDDA.n1991 VDDA.t253 370.168
R233 VDDA.n2008 VDDA.t317 370.168
R234 VDDA.n2001 VDDA.t256 370.168
R235 VDDA.n2017 VDDA.t262 360.868
R236 VDDA.n2071 VDDA.t337 360.868
R237 VDDA.n2112 VDDA.t323 354.154
R238 VDDA.n2111 VDDA.t301 354.154
R239 VDDA.n2097 VDDA.t252 354.154
R240 VDDA.n2096 VDDA.t316 354.154
R241 VDDA.n2084 VDDA.t295 354.063
R242 VDDA.n2083 VDDA.t336 347.224
R243 VDDA.t309 VDDA.n2329 343.882
R244 VDDA.n2330 VDDA.t329 343.882
R245 VDDA.n434 VDDA.t344 343.882
R246 VDDA.t359 VDDA.n433 343.882
R247 VDDA.n2131 VDDA.n2101 342.197
R248 VDDA.n2132 VDDA.n2100 342.197
R249 VDDA.n2120 VDDA.n2116 341.769
R250 VDDA.n2121 VDDA.n2115 341.769
R251 VDDA.n2124 VDDA.n2110 336.341
R252 VDDA.n2125 VDDA.n2109 336.341
R253 VDDA.n2126 VDDA.n2108 336.341
R254 VDDA.n2127 VDDA.n2107 336.341
R255 VDDA.n2128 VDDA.n2106 336.341
R256 VDDA.n2135 VDDA.n2095 336.341
R257 VDDA.n2278 VDDA.t284 333.182
R258 VDDA.n2281 VDDA.t352 333.182
R259 VDDA.n2102 VDDA.t270 332.267
R260 VDDA.n2103 VDDA.t342 332.267
R261 VDDA.n2117 VDDA.t283 332.084
R262 VDDA.n2118 VDDA.t307 332.084
R263 VDDA.n1990 VDDA.n1989 299.231
R264 VDDA.n1988 VDDA.n1987 299.231
R265 VDDA.n1986 VDDA.n1985 299.231
R266 VDDA.n1984 VDDA.n1983 299.231
R267 VDDA.n1982 VDDA.n1981 299.231
R268 VDDA.n1980 VDDA.n1979 299.231
R269 VDDA.n1978 VDDA.n1977 299.231
R270 VDDA.n1976 VDDA.n1975 299.231
R271 VDDA.n1972 VDDA.n1971 299.231
R272 VDDA.n1970 VDDA.n1969 299.231
R273 VDDA.n1968 VDDA.n1967 299.231
R274 VDDA.n1966 VDDA.n1965 299.231
R275 VDDA.n1964 VDDA.n1963 299.231
R276 VDDA.n1962 VDDA.n1961 299.231
R277 VDDA.n1960 VDDA.n1959 299.231
R278 VDDA.n1958 VDDA.n1957 299.231
R279 VDDA.n1956 VDDA.n1955 299.231
R280 VDDA.n1952 VDDA.n1951 299.231
R281 VDDA.n2378 VDDA.n2370 291.053
R282 VDDA.n2378 VDDA.n2377 291.053
R283 VDDA.n2375 VDDA.n2368 291.053
R284 VDDA.n2375 VDDA.n2374 291.053
R285 VDDA.n2384 VDDA.n442 290.233
R286 VDDA.n2385 VDDA.n442 290.233
R287 VDDA.n2358 VDDA.n2348 290.233
R288 VDDA.n2358 VDDA.n2357 290.233
R289 VDDA.n1785 VDDA.t291 267.188
R290 VDDA.t325 VDDA.n1777 267.188
R291 VDDA.t266 VDDA.t27 259.091
R292 VDDA.t27 VDDA.t278 259.091
R293 VDDA.t166 VDDA.t263 251.471
R294 VDDA.t94 VDDA.t166 251.471
R295 VDDA.t56 VDDA.t94 251.471
R296 VDDA.t39 VDDA.t56 251.471
R297 VDDA.t96 VDDA.t39 251.471
R298 VDDA.t179 VDDA.t96 251.471
R299 VDDA.t53 VDDA.t179 251.471
R300 VDDA.t384 VDDA.t53 251.471
R301 VDDA.t388 VDDA.t384 251.471
R302 VDDA.t164 VDDA.t388 251.471
R303 VDDA.t140 VDDA.t164 251.471
R304 VDDA.t177 VDDA.t140 251.471
R305 VDDA.t41 VDDA.t177 251.471
R306 VDDA.t161 VDDA.t41 251.471
R307 VDDA.t175 VDDA.t161 251.471
R308 VDDA.t182 VDDA.t175 251.471
R309 VDDA.t338 VDDA.t182 251.471
R310 VDDA.n2385 VDDA.n2382 242.903
R311 VDDA.n2357 VDDA.n2356 242.903
R312 VDDA.n1776 VDDA.n1775 238.367
R313 VDDA.n1402 VDDA.n1398 238.367
R314 VDDA.n2067 VDDA.n2066 238.367
R315 VDDA.n1994 VDDA.n1993 238.367
R316 VDDA.n1994 VDDA.n1974 238.367
R317 VDDA.n2004 VDDA.n2003 238.367
R318 VDDA.n2004 VDDA.n1954 238.367
R319 VDDA.n2391 VDDA.n2390 238.367
R320 VDDA.n2380 VDDA.n2379 238.367
R321 VDDA.n2376 VDDA.n445 238.367
R322 VDDA.t263 VDDA.n2051 237.5
R323 VDDA.n2068 VDDA.t338 237.5
R324 VDDA.n2355 VDDA.t260 221.121
R325 VDDA.n2381 VDDA.t288 221.121
R326 VDDA.t350 VDDA.n2381 221.121
R327 VDDA.n2389 VDDA.t356 221.121
R328 VDDA.t291 VDDA.t216 217.708
R329 VDDA.t216 VDDA.t325 217.708
R330 VDDA.t396 VDDA.t309 217.708
R331 VDDA.t5 VDDA.t396 217.708
R332 VDDA.t13 VDDA.t5 217.708
R333 VDDA.t152 VDDA.t13 217.708
R334 VDDA.t367 VDDA.t152 217.708
R335 VDDA.t133 VDDA.t367 217.708
R336 VDDA.t15 VDDA.t133 217.708
R337 VDDA.t413 VDDA.t15 217.708
R338 VDDA.t127 VDDA.t413 217.708
R339 VDDA.t397 VDDA.t127 217.708
R340 VDDA.t329 VDDA.t397 217.708
R341 VDDA.t344 VDDA.t146 217.708
R342 VDDA.t146 VDDA.t101 217.708
R343 VDDA.t101 VDDA.t160 217.708
R344 VDDA.t160 VDDA.t18 217.708
R345 VDDA.t18 VDDA.t404 217.708
R346 VDDA.t404 VDDA.t173 217.708
R347 VDDA.t173 VDDA.t401 217.708
R348 VDDA.t401 VDDA.t147 217.708
R349 VDDA.t147 VDDA.t144 217.708
R350 VDDA.t144 VDDA.t410 217.708
R351 VDDA.t410 VDDA.t359 217.708
R352 VDDA.n441 VDDA.n440 216.677
R353 VDDA.n2363 VDDA.n2362 216.677
R354 VDDA.t272 VDDA.n381 213.131
R355 VDDA.n382 VDDA.t297 213.131
R356 VDDA.n2405 VDDA.t408 213.131
R357 VDDA.t72 VDDA.n367 213.131
R358 VDDA.t285 VDDA.n2279 213.131
R359 VDDA.n2280 VDDA.t353 213.131
R360 VDDA.n1401 VDDA.n1399 185
R361 VDDA.n1772 VDDA.n1771 185
R362 VDDA.n1784 VDDA.n1783 185
R363 VDDA.n1785 VDDA.n1784 185
R364 VDDA.n1781 VDDA.n1778 185
R365 VDDA.n1780 VDDA.n1396 185
R366 VDDA.n1787 VDDA.n1786 185
R367 VDDA.n1786 VDDA.n1785 185
R368 VDDA.n2056 VDDA.n2054 185
R369 VDDA.n2063 VDDA.n2053 185
R370 VDDA.n2068 VDDA.n2053 185
R371 VDDA.n2062 VDDA.n2061 185
R372 VDDA.n2059 VDDA.n2028 185
R373 VDDA.n2070 VDDA.n2069 185
R374 VDDA.n2069 VDDA.n2068 185
R375 VDDA.n2050 VDDA.n2049 185
R376 VDDA.n2051 VDDA.n2050 185
R377 VDDA.n2047 VDDA.n2032 185
R378 VDDA.n2046 VDDA.n2045 185
R379 VDDA.n2044 VDDA.n2043 185
R380 VDDA.n2038 VDDA.n2037 185
R381 VDDA.n2040 VDDA.n2031 185
R382 VDDA.n2051 VDDA.n2031 185
R383 VDDA.n2369 VDDA.n447 185
R384 VDDA.n2373 VDDA.n446 185
R385 VDDA.n2381 VDDA.n446 185
R386 VDDA.n2372 VDDA.n2371 185
R387 VDDA.n444 VDDA.n443 185
R388 VDDA.n2388 VDDA.n2387 185
R389 VDDA.n2389 VDDA.n2388 185
R390 VDDA.n2386 VDDA.n2383 185
R391 VDDA.n2359 VDDA.n2346 185
R392 VDDA.n2355 VDDA.n2346 185
R393 VDDA.n2351 VDDA.n2347 185
R394 VDDA.n2353 VDDA.n2352 185
R395 VDDA.n2350 VDDA.n2349 185
R396 VDDA.t260 VDDA.t12 180.173
R397 VDDA.t12 VDDA.t192 180.173
R398 VDDA.t192 VDDA.t29 180.173
R399 VDDA.t29 VDDA.t35 180.173
R400 VDDA.t35 VDDA.t288 180.173
R401 VDDA.t103 VDDA.t350 180.173
R402 VDDA.t118 VDDA.t103 180.173
R403 VDDA.t25 VDDA.t118 180.173
R404 VDDA.t36 VDDA.t25 180.173
R405 VDDA.t356 VDDA.t36 180.173
R406 VDDA.n375 VDDA.t267 168.139
R407 VDDA.n374 VDDA.t280 168.139
R408 VDDA.n372 VDDA.n371 150.643
R409 VDDA.n1771 VDDA.n1399 150
R410 VDDA.n1784 VDDA.n1778 150
R411 VDDA.n1786 VDDA.n1396 150
R412 VDDA.n2054 VDDA.n2053 150
R413 VDDA.n2061 VDDA.n2053 150
R414 VDDA.n2069 VDDA.n2028 150
R415 VDDA.n2050 VDDA.n2032 150
R416 VDDA.n2045 VDDA.n2044 150
R417 VDDA.n2037 VDDA.n2031 150
R418 VDDA.n2388 VDDA.n444 150
R419 VDDA.n2388 VDDA.n2383 150
R420 VDDA.n447 VDDA.n446 150
R421 VDDA.n2371 VDDA.n446 150
R422 VDDA.n2351 VDDA.n2346 150
R423 VDDA.n2353 VDDA.n2350 150
R424 VDDA.n1404 VDDA.n1403 149.112
R425 VDDA.t78 VDDA.t272 146.155
R426 VDDA.t297 VDDA.t78 146.155
R427 VDDA.t408 VDDA.t1 146.155
R428 VDDA.t1 VDDA.t120 146.155
R429 VDDA.t120 VDDA.t376 146.155
R430 VDDA.t376 VDDA.t86 146.155
R431 VDDA.t86 VDDA.t378 146.155
R432 VDDA.t378 VDDA.t90 146.155
R433 VDDA.t90 VDDA.t3 146.155
R434 VDDA.t3 VDDA.t80 146.155
R435 VDDA.t80 VDDA.t74 146.155
R436 VDDA.t74 VDDA.t361 146.155
R437 VDDA.t361 VDDA.t72 146.155
R438 VDDA.t113 VDDA.t285 146.155
R439 VDDA.t122 VDDA.t113 146.155
R440 VDDA.t76 VDDA.t122 146.155
R441 VDDA.t107 VDDA.t76 146.155
R442 VDDA.t92 VDDA.t107 146.155
R443 VDDA.t6 VDDA.t92 146.155
R444 VDDA.t88 VDDA.t6 146.155
R445 VDDA.t363 VDDA.t88 146.155
R446 VDDA.t368 VDDA.t363 146.155
R447 VDDA.t370 VDDA.t368 146.155
R448 VDDA.t353 VDDA.t370 146.155
R449 VDDA.n2072 VDDA.n2025 141.712
R450 VDDA.n2073 VDDA.n2024 141.712
R451 VDDA.n2074 VDDA.n2023 141.712
R452 VDDA.n2075 VDDA.n2022 141.712
R453 VDDA.n2076 VDDA.n2021 141.712
R454 VDDA.n2077 VDDA.n2020 141.712
R455 VDDA.n2078 VDDA.n2019 141.712
R456 VDDA.n2079 VDDA.n2018 141.712
R457 VDDA.n2329 VDDA.t310 136.701
R458 VDDA.n2330 VDDA.t330 136.701
R459 VDDA.n434 VDDA.t345 136.701
R460 VDDA.n433 VDDA.t360 136.701
R461 VDDA.t264 VDDA.n2035 123.126
R462 VDDA.n2036 VDDA.t264 123.126
R463 VDDA.n2064 VDDA.t339 123.126
R464 VDDA.n2060 VDDA.t339 123.126
R465 VDDA.n403 VDDA.t332 122.829
R466 VDDA.t347 VDDA.n402 122.829
R467 VDDA.t303 VDDA.n2302 122.829
R468 VDDA.n2303 VDDA.t312 122.829
R469 VDDA.t332 VDDA.t8 81.6411
R470 VDDA.t8 VDDA.t380 81.6411
R471 VDDA.t380 VDDA.t417 81.6411
R472 VDDA.t417 VDDA.t130 81.6411
R473 VDDA.t130 VDDA.t415 81.6411
R474 VDDA.t415 VDDA.t16 81.6411
R475 VDDA.t16 VDDA.t128 81.6411
R476 VDDA.t128 VDDA.t402 81.6411
R477 VDDA.t402 VDDA.t149 81.6411
R478 VDDA.t149 VDDA.t115 81.6411
R479 VDDA.t115 VDDA.t347 81.6411
R480 VDDA.t109 VDDA.t303 81.6411
R481 VDDA.t63 VDDA.t109 81.6411
R482 VDDA.t374 VDDA.t63 81.6411
R483 VDDA.t372 VDDA.t374 81.6411
R484 VDDA.t111 VDDA.t372 81.6411
R485 VDDA.t398 VDDA.t111 81.6411
R486 VDDA.t134 VDDA.t398 81.6411
R487 VDDA.t142 VDDA.t134 81.6411
R488 VDDA.t171 VDDA.t142 81.6411
R489 VDDA.t411 VDDA.t171 81.6411
R490 VDDA.t312 VDDA.t411 81.6411
R491 VDDA.n381 VDDA.t273 76.2576
R492 VDDA.n382 VDDA.t298 76.2576
R493 VDDA.n2405 VDDA.t409 76.2576
R494 VDDA.n367 VDDA.t73 76.2576
R495 VDDA.n2279 VDDA.t286 76.2576
R496 VDDA.n2280 VDDA.t354 76.2576
R497 VDDA.n2417 VDDA.n2416 71.388
R498 VDDA.n2415 VDDA.n2414 71.388
R499 VDDA.n2410 VDDA.n2409 71.388
R500 VDDA.n2408 VDDA.n2407 71.388
R501 VDDA.n2274 VDDA.n2273 71.388
R502 VDDA.n2276 VDDA.n2275 71.388
R503 VDDA.n455 VDDA.n454 71.388
R504 VDDA.n2269 VDDA.n2268 71.388
R505 VDDA.n379 VDDA.n378 68.4557
R506 VDDA.n2412 VDDA.n2411 66.888
R507 VDDA.n2271 VDDA.n2270 66.888
R508 VDDA.n1777 VDDA.n1776 65.8183
R509 VDDA.n1777 VDDA.n1398 65.8183
R510 VDDA.n1785 VDDA.n1397 65.8183
R511 VDDA.n2068 VDDA.n2067 65.8183
R512 VDDA.n2068 VDDA.n2052 65.8183
R513 VDDA.n2051 VDDA.n2029 65.8183
R514 VDDA.n2051 VDDA.n2030 65.8183
R515 VDDA.n2381 VDDA.n2380 65.8183
R516 VDDA.n2381 VDDA.n445 65.8183
R517 VDDA.n2390 VDDA.n2389 65.8183
R518 VDDA.n2389 VDDA.n2382 65.8183
R519 VDDA.n2355 VDDA.n2354 65.8183
R520 VDDA.n2356 VDDA.n2355 65.8183
R521 VDDA.n1942 VDDA.t419 58.8005
R522 VDDA.n1941 VDDA.t421 58.8005
R523 VDDA.n2392 VDDA.n2391 58.0576
R524 VDDA.n2360 VDDA.n2359 58.0576
R525 VDDA.n2367 VDDA.n2366 54.4005
R526 VDDA.n2367 VDDA.n448 54.4005
R527 VDDA.n1776 VDDA.n1399 53.3664
R528 VDDA.n1771 VDDA.n1398 53.3664
R529 VDDA.n1778 VDDA.n1397 53.3664
R530 VDDA.n1397 VDDA.n1396 53.3664
R531 VDDA.n2061 VDDA.n2052 53.3664
R532 VDDA.n2067 VDDA.n2054 53.3664
R533 VDDA.n2052 VDDA.n2028 53.3664
R534 VDDA.n2032 VDDA.n2029 53.3664
R535 VDDA.n2044 VDDA.n2030 53.3664
R536 VDDA.n2045 VDDA.n2029 53.3664
R537 VDDA.n2037 VDDA.n2030 53.3664
R538 VDDA.n2383 VDDA.n2382 53.3664
R539 VDDA.n2371 VDDA.n445 53.3664
R540 VDDA.n2380 VDDA.n447 53.3664
R541 VDDA.n2390 VDDA.n444 53.3664
R542 VDDA.n2354 VDDA.n2351 53.3664
R543 VDDA.n2356 VDDA.n2350 53.3664
R544 VDDA.n2354 VDDA.n2353 53.3664
R545 VDDA.n1941 VDDA.t422 49.1638
R546 VDDA.n1943 VDDA.t420 48.5162
R547 VDDA.n403 VDDA.t333 40.9789
R548 VDDA.n402 VDDA.t348 40.9789
R549 VDDA.n2302 VDDA.t304 40.9789
R550 VDDA.n2303 VDDA.t313 40.9789
R551 VDDA.n2116 VDDA.t227 39.4005
R552 VDDA.n2116 VDDA.t247 39.4005
R553 VDDA.n2115 VDDA.t249 39.4005
R554 VDDA.n2115 VDDA.t239 39.4005
R555 VDDA.n2110 VDDA.t215 39.4005
R556 VDDA.n2110 VDDA.t322 39.4005
R557 VDDA.n2109 VDDA.t231 39.4005
R558 VDDA.n2109 VDDA.t233 39.4005
R559 VDDA.n2108 VDDA.t223 39.4005
R560 VDDA.n2108 VDDA.t241 39.4005
R561 VDDA.n2107 VDDA.t245 39.4005
R562 VDDA.n2107 VDDA.t237 39.4005
R563 VDDA.t301 VDDA.n2106 39.4005
R564 VDDA.n2106 VDDA.t225 39.4005
R565 VDDA.n2101 VDDA.t235 39.4005
R566 VDDA.n2101 VDDA.t219 39.4005
R567 VDDA.n2100 VDDA.t221 39.4005
R568 VDDA.n2100 VDDA.t243 39.4005
R569 VDDA.n2095 VDDA.t229 39.4005
R570 VDDA.n2095 VDDA.t213 39.4005
R571 VDDA.n1989 VDDA.t83 39.4005
R572 VDDA.n1989 VDDA.t205 39.4005
R573 VDDA.n1987 VDDA.t46 39.4005
R574 VDDA.n1987 VDDA.t391 39.4005
R575 VDDA.n1985 VDDA.t201 39.4005
R576 VDDA.n1985 VDDA.t24 39.4005
R577 VDDA.n1983 VDDA.t366 39.4005
R578 VDDA.n1983 VDDA.t209 39.4005
R579 VDDA.n1981 VDDA.t383 39.4005
R580 VDDA.n1981 VDDA.t106 39.4005
R581 VDDA.n1979 VDDA.t203 39.4005
R582 VDDA.n1979 VDDA.t169 39.4005
R583 VDDA.n1977 VDDA.t50 39.4005
R584 VDDA.n1977 VDDA.t211 39.4005
R585 VDDA.n1975 VDDA.t44 39.4005
R586 VDDA.n1975 VDDA.t159 39.4005
R587 VDDA.n1971 VDDA.t207 39.4005
R588 VDDA.n1971 VDDA.t38 39.4005
R589 VDDA.n1969 VDDA.t185 39.4005
R590 VDDA.n1969 VDDA.t61 39.4005
R591 VDDA.n1967 VDDA.t157 39.4005
R592 VDDA.n1967 VDDA.t32 39.4005
R593 VDDA.n1965 VDDA.t34 39.4005
R594 VDDA.n1965 VDDA.t187 39.4005
R595 VDDA.n1963 VDDA.t11 39.4005
R596 VDDA.n1963 VDDA.t189 39.4005
R597 VDDA.n1961 VDDA.t191 39.4005
R598 VDDA.n1961 VDDA.t406 39.4005
R599 VDDA.n1959 VDDA.t20 39.4005
R600 VDDA.n1959 VDDA.t22 39.4005
R601 VDDA.n1957 VDDA.t195 39.4005
R602 VDDA.n1957 VDDA.t155 39.4005
R603 VDDA.n1955 VDDA.t71 39.4005
R604 VDDA.n1955 VDDA.t197 39.4005
R605 VDDA.n1951 VDDA.t48 39.4005
R606 VDDA.n1951 VDDA.t199 39.4005
R607 VDDA.n400 VDDA.n399 38.2279
R608 VDDA.n398 VDDA.n397 38.2279
R609 VDDA.n396 VDDA.n395 38.2279
R610 VDDA.n394 VDDA.n393 38.2279
R611 VDDA.n392 VDDA.n391 38.2279
R612 VDDA.n2292 VDDA.n2291 38.2279
R613 VDDA.n2294 VDDA.n2293 38.2279
R614 VDDA.n2296 VDDA.n2295 38.2279
R615 VDDA.n2298 VDDA.n2297 38.2279
R616 VDDA.n2300 VDDA.n2299 38.2279
R617 VDDA.n2119 VDDA.n2118 27.2462
R618 VDDA.n2117 VDDA.n2114 27.2462
R619 VDDA.n2104 VDDA.n2103 27.2462
R620 VDDA.n2102 VDDA.n2099 27.2462
R621 VDDA.n417 VDDA.n415 26.9096
R622 VDDA.n2314 VDDA.n2312 26.8887
R623 VDDA.n417 VDDA.n416 26.795
R624 VDDA.n419 VDDA.n418 26.795
R625 VDDA.n421 VDDA.n420 26.795
R626 VDDA.n423 VDDA.n422 26.795
R627 VDDA.n425 VDDA.n424 26.795
R628 VDDA.n2322 VDDA.n2321 26.7741
R629 VDDA.n2320 VDDA.n2319 26.7741
R630 VDDA.n2318 VDDA.n2317 26.7741
R631 VDDA.n2316 VDDA.n2315 26.7741
R632 VDDA.n2314 VDDA.n2313 26.7741
R633 VDDA.n2113 VDDA.n2112 24.9931
R634 VDDA.n2111 VDDA.n2105 24.9931
R635 VDDA.n2098 VDDA.n2097 24.9931
R636 VDDA.n2096 VDDA.n2094 24.9931
R637 VDDA.n1463 VDDA.t386 24.1029
R638 VDDA.n2085 VDDA.n2084 22.9536
R639 VDDA.n2071 VDDA.n2070 22.8576
R640 VDDA.n2040 VDDA.n2017 22.8576
R641 VDDA.n371 VDDA.t28 21.8894
R642 VDDA.n371 VDDA.t279 21.8894
R643 VDDA.n2083 VDDA.n2082 20.4312
R644 VDDA.n1403 VDDA.t217 19.7005
R645 VDDA.n1403 VDDA.t326 19.7005
R646 VDDA.n2358 VDDA.t261 15.7605
R647 VDDA.n442 VDDA.t357 15.7605
R648 VDDA.n2375 VDDA.t351 15.7605
R649 VDDA.n2378 VDDA.t289 15.7605
R650 VDDA.n440 VDDA.t119 15.7605
R651 VDDA.n440 VDDA.t26 15.7605
R652 VDDA.n2362 VDDA.t193 15.7605
R653 VDDA.n2362 VDDA.t30 15.7605
R654 VDDA.n2025 VDDA.t176 13.1338
R655 VDDA.n2025 VDDA.t183 13.1338
R656 VDDA.n2024 VDDA.t42 13.1338
R657 VDDA.n2024 VDDA.t162 13.1338
R658 VDDA.n2023 VDDA.t141 13.1338
R659 VDDA.n2023 VDDA.t178 13.1338
R660 VDDA.n2022 VDDA.t389 13.1338
R661 VDDA.n2022 VDDA.t165 13.1338
R662 VDDA.n2021 VDDA.t54 13.1338
R663 VDDA.n2021 VDDA.t385 13.1338
R664 VDDA.n2020 VDDA.t97 13.1338
R665 VDDA.n2020 VDDA.t180 13.1338
R666 VDDA.n2019 VDDA.t57 13.1338
R667 VDDA.n2019 VDDA.t40 13.1338
R668 VDDA.n2018 VDDA.t167 13.1338
R669 VDDA.n2018 VDDA.t95 13.1338
R670 VDDA.n2082 VDDA.n2081 11.37
R671 VDDA.n2086 VDDA.n2085 11.37
R672 VDDA.t273 VDDA.n379 11.2576
R673 VDDA.n379 VDDA.t79 11.2576
R674 VDDA.n2416 VDDA.t75 11.2576
R675 VDDA.n2416 VDDA.t362 11.2576
R676 VDDA.n2414 VDDA.t4 11.2576
R677 VDDA.n2414 VDDA.t81 11.2576
R678 VDDA.n2411 VDDA.t379 11.2576
R679 VDDA.n2411 VDDA.t91 11.2576
R680 VDDA.n2409 VDDA.t377 11.2576
R681 VDDA.n2409 VDDA.t87 11.2576
R682 VDDA.n2407 VDDA.t2 11.2576
R683 VDDA.n2407 VDDA.t121 11.2576
R684 VDDA.n2273 VDDA.t77 11.2576
R685 VDDA.n2273 VDDA.t108 11.2576
R686 VDDA.n2275 VDDA.t114 11.2576
R687 VDDA.n2275 VDDA.t123 11.2576
R688 VDDA.n454 VDDA.t369 11.2576
R689 VDDA.n454 VDDA.t371 11.2576
R690 VDDA.n2268 VDDA.t89 11.2576
R691 VDDA.n2268 VDDA.t364 11.2576
R692 VDDA.n2270 VDDA.t93 11.2576
R693 VDDA.n2270 VDDA.t7 11.2576
R694 VDDA.n2072 VDDA.n2071 11.0575
R695 VDDA.n2120 VDDA.n2119 10.9846
R696 VDDA.n2122 VDDA.n2114 10.87
R697 VDDA.n2129 VDDA.n2105 10.87
R698 VDDA.n2133 VDDA.n2099 10.87
R699 VDDA.n2136 VDDA.n2094 10.87
R700 VDDA.n2134 VDDA.n2098 10.87
R701 VDDA.n2130 VDDA.n2104 10.87
R702 VDDA.n2123 VDDA.n2113 10.87
R703 VDDA.n2080 VDDA.n2017 10.87
R704 VDDA.n2361 VDDA.n2360 10.8696
R705 VDDA.n2364 VDDA.n448 10.869
R706 VDDA.n2366 VDDA.n2365 10.869
R707 VDDA.n2393 VDDA.n2392 10.869
R708 VDDA.n1775 VDDA.n1400 9.50883
R709 VDDA.n1783 VDDA.n1782 9.50883
R710 VDDA.n2049 VDDA.n2048 9.50883
R711 VDDA.n2041 VDDA.n2040 9.50883
R712 VDDA.n2066 VDDA.n2055 9.50883
R713 VDDA.n2070 VDDA.n2027 9.50883
R714 VDDA.n1997 VDDA.n1973 9.50883
R715 VDDA.n2007 VDDA.n1953 9.50883
R716 VDDA.n1772 VDDA.n1770 9.3005
R717 VDDA.n1401 VDDA.n1400 9.3005
R718 VDDA.n1769 VDDA.n1402 9.3005
R719 VDDA.n1780 VDDA.n1394 9.3005
R720 VDDA.n1782 VDDA.n1781 9.3005
R721 VDDA.n1788 VDDA.n1787 9.3005
R722 VDDA.n2059 VDDA.n2027 9.3005
R723 VDDA.n2062 VDDA.n2058 9.3005
R724 VDDA.n2063 VDDA.n2057 9.3005
R725 VDDA.n2056 VDDA.n2055 9.3005
R726 VDDA.n2041 VDDA.n2038 9.3005
R727 VDDA.n2043 VDDA.n2042 9.3005
R728 VDDA.n2046 VDDA.n2034 9.3005
R729 VDDA.n2048 VDDA.n2047 9.3005
R730 VDDA.n1997 VDDA.n1996 9.3005
R731 VDDA.n2007 VDDA.n2006 9.3005
R732 VDDA.n1772 VDDA.n1401 9.14336
R733 VDDA.n1781 VDDA.n1780 9.14336
R734 VDDA.n2063 VDDA.n2056 9.14336
R735 VDDA.n2063 VDDA.n2062 9.14336
R736 VDDA.n2062 VDDA.n2059 9.14336
R737 VDDA.n2047 VDDA.n2046 9.14336
R738 VDDA.n2046 VDDA.n2043 9.14336
R739 VDDA.n2043 VDDA.n2038 9.14336
R740 VDDA.n2391 VDDA.n443 9.14336
R741 VDDA.n2387 VDDA.n2386 9.14336
R742 VDDA.n2359 VDDA.n2347 9.14336
R743 VDDA.n2352 VDDA.n2349 9.14336
R744 VDDA.n2321 VDDA.t126 8.0005
R745 VDDA.n2321 VDDA.t84 8.0005
R746 VDDA.n2319 VDDA.t170 8.0005
R747 VDDA.n2319 VDDA.t65 8.0005
R748 VDDA.n2317 VDDA.t151 8.0005
R749 VDDA.n2317 VDDA.t62 8.0005
R750 VDDA.n2315 VDDA.t153 8.0005
R751 VDDA.n2315 VDDA.t407 8.0005
R752 VDDA.n2313 VDDA.t14 8.0005
R753 VDDA.n2313 VDDA.t100 8.0005
R754 VDDA.n2312 VDDA.t124 8.0005
R755 VDDA.n2312 VDDA.t125 8.0005
R756 VDDA.n415 VDDA.t67 8.0005
R757 VDDA.n415 VDDA.t85 8.0005
R758 VDDA.n416 VDDA.t132 8.0005
R759 VDDA.n416 VDDA.t414 8.0005
R760 VDDA.n418 VDDA.t66 8.0005
R761 VDDA.n418 VDDA.t145 8.0005
R762 VDDA.n420 VDDA.t102 8.0005
R763 VDDA.n420 VDDA.t148 8.0005
R764 VDDA.n422 VDDA.t117 8.0005
R765 VDDA.n422 VDDA.t400 8.0005
R766 VDDA.n424 VDDA.t104 8.0005
R767 VDDA.n424 VDDA.t136 8.0005
R768 VDDA.n399 VDDA.t150 6.56717
R769 VDDA.n399 VDDA.t116 6.56717
R770 VDDA.n397 VDDA.t129 6.56717
R771 VDDA.n397 VDDA.t403 6.56717
R772 VDDA.n395 VDDA.t416 6.56717
R773 VDDA.n395 VDDA.t17 6.56717
R774 VDDA.n393 VDDA.t418 6.56717
R775 VDDA.n393 VDDA.t131 6.56717
R776 VDDA.n391 VDDA.t9 6.56717
R777 VDDA.n391 VDDA.t381 6.56717
R778 VDDA.n2291 VDDA.t172 6.56717
R779 VDDA.n2291 VDDA.t412 6.56717
R780 VDDA.n2293 VDDA.t135 6.56717
R781 VDDA.n2293 VDDA.t143 6.56717
R782 VDDA.n2295 VDDA.t112 6.56717
R783 VDDA.n2295 VDDA.t399 6.56717
R784 VDDA.n2297 VDDA.t375 6.56717
R785 VDDA.n2297 VDDA.t373 6.56717
R786 VDDA.n2299 VDDA.t110 6.56717
R787 VDDA.n2299 VDDA.t64 6.56717
R788 VDDA.n1775 VDDA.n1774 5.33286
R789 VDDA.n1773 VDDA.n1402 5.33286
R790 VDDA.n1783 VDDA.n1779 5.33286
R791 VDDA.n1787 VDDA.n1395 5.33286
R792 VDDA.n2066 VDDA.n2065 5.33286
R793 VDDA.n2070 VDDA.n2026 5.33286
R794 VDDA.n2049 VDDA.n2033 5.33286
R795 VDDA.n2040 VDDA.n2039 5.33286
R796 VDDA.n2408 VDDA.n2406 5.1255
R797 VDDA.n2418 VDDA.n2417 5.1255
R798 VDDA.n2282 VDDA.n455 5.1255
R799 VDDA.n2277 VDDA.n2276 5.1255
R800 VDDA.n2384 VDDA.n443 4.53698
R801 VDDA.n2386 VDDA.n2385 4.53698
R802 VDDA.n2387 VDDA.n2384 4.53698
R803 VDDA.n2348 VDDA.n2347 4.53698
R804 VDDA.n2357 VDDA.n2349 4.53698
R805 VDDA.n2352 VDDA.n2348 4.53698
R806 VDDA.n1792 VDDA.n1791 4.5005
R807 VDDA.n1795 VDDA.n1794 4.5005
R808 VDDA.n1796 VDDA.n1392 4.5005
R809 VDDA.n1800 VDDA.n1797 4.5005
R810 VDDA.n1801 VDDA.n1391 4.5005
R811 VDDA.n1805 VDDA.n1804 4.5005
R812 VDDA.n1806 VDDA.n1390 4.5005
R813 VDDA.n1810 VDDA.n1807 4.5005
R814 VDDA.n1811 VDDA.n1389 4.5005
R815 VDDA.n1815 VDDA.n1814 4.5005
R816 VDDA.n1816 VDDA.n1388 4.5005
R817 VDDA.n1820 VDDA.n1817 4.5005
R818 VDDA.n1821 VDDA.n1387 4.5005
R819 VDDA.n1825 VDDA.n1824 4.5005
R820 VDDA.n1826 VDDA.n1386 4.5005
R821 VDDA.n1830 VDDA.n1827 4.5005
R822 VDDA.n1831 VDDA.n1385 4.5005
R823 VDDA.n1835 VDDA.n1834 4.5005
R824 VDDA.n1836 VDDA.n1384 4.5005
R825 VDDA.n1840 VDDA.n1837 4.5005
R826 VDDA.n1841 VDDA.n1383 4.5005
R827 VDDA.n1845 VDDA.n1844 4.5005
R828 VDDA.n1846 VDDA.n1382 4.5005
R829 VDDA.n1850 VDDA.n1847 4.5005
R830 VDDA.n1851 VDDA.n1381 4.5005
R831 VDDA.n1855 VDDA.n1854 4.5005
R832 VDDA.n1856 VDDA.n1380 4.5005
R833 VDDA.n1860 VDDA.n1857 4.5005
R834 VDDA.n1861 VDDA.n1379 4.5005
R835 VDDA.n1865 VDDA.n1864 4.5005
R836 VDDA.n1866 VDDA.n1378 4.5005
R837 VDDA.n1870 VDDA.n1867 4.5005
R838 VDDA.n1871 VDDA.n1377 4.5005
R839 VDDA.n1875 VDDA.n1874 4.5005
R840 VDDA.n1876 VDDA.n1376 4.5005
R841 VDDA.n1880 VDDA.n1877 4.5005
R842 VDDA.n1881 VDDA.n1375 4.5005
R843 VDDA.n1885 VDDA.n1884 4.5005
R844 VDDA.n1886 VDDA.n1374 4.5005
R845 VDDA.n1890 VDDA.n1887 4.5005
R846 VDDA.n1891 VDDA.n1373 4.5005
R847 VDDA.n1895 VDDA.n1894 4.5005
R848 VDDA.n1896 VDDA.n1372 4.5005
R849 VDDA.n1900 VDDA.n1897 4.5005
R850 VDDA.n1901 VDDA.n1371 4.5005
R851 VDDA.n1905 VDDA.n1904 4.5005
R852 VDDA.n1464 VDDA.n1463 4.5005
R853 VDDA.n1467 VDDA.n1466 4.5005
R854 VDDA.n1468 VDDA.n1457 4.5005
R855 VDDA.n1472 VDDA.n1469 4.5005
R856 VDDA.n1473 VDDA.n1456 4.5005
R857 VDDA.n1477 VDDA.n1476 4.5005
R858 VDDA.n1478 VDDA.n1455 4.5005
R859 VDDA.n1482 VDDA.n1479 4.5005
R860 VDDA.n1483 VDDA.n1454 4.5005
R861 VDDA.n1487 VDDA.n1486 4.5005
R862 VDDA.n1488 VDDA.n1453 4.5005
R863 VDDA.n1492 VDDA.n1489 4.5005
R864 VDDA.n1493 VDDA.n1452 4.5005
R865 VDDA.n1497 VDDA.n1496 4.5005
R866 VDDA.n1498 VDDA.n1451 4.5005
R867 VDDA.n1502 VDDA.n1499 4.5005
R868 VDDA.n1503 VDDA.n1450 4.5005
R869 VDDA.n1507 VDDA.n1506 4.5005
R870 VDDA.n1508 VDDA.n1449 4.5005
R871 VDDA.n1512 VDDA.n1509 4.5005
R872 VDDA.n1513 VDDA.n1448 4.5005
R873 VDDA.n1517 VDDA.n1516 4.5005
R874 VDDA.n1518 VDDA.n1447 4.5005
R875 VDDA.n1522 VDDA.n1519 4.5005
R876 VDDA.n1523 VDDA.n1446 4.5005
R877 VDDA.n1527 VDDA.n1526 4.5005
R878 VDDA.n1528 VDDA.n1445 4.5005
R879 VDDA.n1532 VDDA.n1529 4.5005
R880 VDDA.n1533 VDDA.n1444 4.5005
R881 VDDA.n1537 VDDA.n1536 4.5005
R882 VDDA.n1538 VDDA.n1443 4.5005
R883 VDDA.n1542 VDDA.n1539 4.5005
R884 VDDA.n1543 VDDA.n1442 4.5005
R885 VDDA.n1547 VDDA.n1546 4.5005
R886 VDDA.n1548 VDDA.n1441 4.5005
R887 VDDA.n1552 VDDA.n1549 4.5005
R888 VDDA.n1553 VDDA.n1440 4.5005
R889 VDDA.n1557 VDDA.n1556 4.5005
R890 VDDA.n1558 VDDA.n1439 4.5005
R891 VDDA.n1562 VDDA.n1559 4.5005
R892 VDDA.n1563 VDDA.n1438 4.5005
R893 VDDA.n1567 VDDA.n1566 4.5005
R894 VDDA.n1568 VDDA.n1437 4.5005
R895 VDDA.n1572 VDDA.n1569 4.5005
R896 VDDA.n1573 VDDA.n1436 4.5005
R897 VDDA.n1577 VDDA.n1576 4.5005
R898 VDDA.n1947 VDDA.n1946 4.5005
R899 VDDA.n2013 VDDA.n2012 4.5005
R900 VDDA.n2090 VDDA.n2089 4.5005
R901 VDDA.n2140 VDDA.n2139 4.5005
R902 VDDA.n2144 VDDA.n2143 4.5005
R903 VDDA.n2145 VDDA.n1932 4.5005
R904 VDDA.n2149 VDDA.n2146 4.5005
R905 VDDA.n2150 VDDA.n1931 4.5005
R906 VDDA.n2154 VDDA.n2153 4.5005
R907 VDDA.n2155 VDDA.n1930 4.5005
R908 VDDA.n2159 VDDA.n2156 4.5005
R909 VDDA.n2160 VDDA.n1929 4.5005
R910 VDDA.n2164 VDDA.n2163 4.5005
R911 VDDA.n2165 VDDA.n1928 4.5005
R912 VDDA.n2169 VDDA.n2166 4.5005
R913 VDDA.n2170 VDDA.n1927 4.5005
R914 VDDA.n2174 VDDA.n2173 4.5005
R915 VDDA.n2175 VDDA.n1926 4.5005
R916 VDDA.n2179 VDDA.n2176 4.5005
R917 VDDA.n2180 VDDA.n1925 4.5005
R918 VDDA.n2184 VDDA.n2183 4.5005
R919 VDDA.n2185 VDDA.n1924 4.5005
R920 VDDA.n2189 VDDA.n2186 4.5005
R921 VDDA.n2190 VDDA.n1923 4.5005
R922 VDDA.n2194 VDDA.n2193 4.5005
R923 VDDA.n2195 VDDA.n1922 4.5005
R924 VDDA.n2199 VDDA.n2196 4.5005
R925 VDDA.n2200 VDDA.n1921 4.5005
R926 VDDA.n2204 VDDA.n2203 4.5005
R927 VDDA.n2205 VDDA.n1920 4.5005
R928 VDDA.n2209 VDDA.n2206 4.5005
R929 VDDA.n2210 VDDA.n1919 4.5005
R930 VDDA.n2214 VDDA.n2213 4.5005
R931 VDDA.n2215 VDDA.n1918 4.5005
R932 VDDA.n2219 VDDA.n2216 4.5005
R933 VDDA.n2220 VDDA.n1917 4.5005
R934 VDDA.n2224 VDDA.n2223 4.5005
R935 VDDA.n2225 VDDA.n1916 4.5005
R936 VDDA.n2229 VDDA.n2226 4.5005
R937 VDDA.n2230 VDDA.n1915 4.5005
R938 VDDA.n2234 VDDA.n2233 4.5005
R939 VDDA.n2235 VDDA.n1914 4.5005
R940 VDDA.n2239 VDDA.n2236 4.5005
R941 VDDA.n2240 VDDA.n1913 4.5005
R942 VDDA.n2244 VDDA.n2243 4.5005
R943 VDDA.n2245 VDDA.n1912 4.5005
R944 VDDA.n2249 VDDA.n2246 4.5005
R945 VDDA.n2250 VDDA.n1911 4.5005
R946 VDDA.n2254 VDDA.n2253 4.5005
R947 VDDA.n93 VDDA.n87 4.5005
R948 VDDA.n95 VDDA.n94 4.5005
R949 VDDA.n96 VDDA.n86 4.5005
R950 VDDA.n100 VDDA.n99 4.5005
R951 VDDA.n101 VDDA.n83 4.5005
R952 VDDA.n103 VDDA.n102 4.5005
R953 VDDA.n104 VDDA.n82 4.5005
R954 VDDA.n108 VDDA.n107 4.5005
R955 VDDA.n109 VDDA.n79 4.5005
R956 VDDA.n111 VDDA.n110 4.5005
R957 VDDA.n112 VDDA.n78 4.5005
R958 VDDA.n116 VDDA.n115 4.5005
R959 VDDA.n117 VDDA.n75 4.5005
R960 VDDA.n119 VDDA.n118 4.5005
R961 VDDA.n120 VDDA.n74 4.5005
R962 VDDA.n124 VDDA.n123 4.5005
R963 VDDA.n125 VDDA.n71 4.5005
R964 VDDA.n127 VDDA.n126 4.5005
R965 VDDA.n128 VDDA.n70 4.5005
R966 VDDA.n132 VDDA.n131 4.5005
R967 VDDA.n133 VDDA.n67 4.5005
R968 VDDA.n135 VDDA.n134 4.5005
R969 VDDA.n136 VDDA.n66 4.5005
R970 VDDA.n140 VDDA.n139 4.5005
R971 VDDA.n141 VDDA.n63 4.5005
R972 VDDA.n143 VDDA.n142 4.5005
R973 VDDA.n144 VDDA.n62 4.5005
R974 VDDA.n148 VDDA.n147 4.5005
R975 VDDA.n149 VDDA.n59 4.5005
R976 VDDA.n151 VDDA.n150 4.5005
R977 VDDA.n152 VDDA.n58 4.5005
R978 VDDA.n156 VDDA.n155 4.5005
R979 VDDA.n157 VDDA.n55 4.5005
R980 VDDA.n159 VDDA.n158 4.5005
R981 VDDA.n160 VDDA.n54 4.5005
R982 VDDA.n164 VDDA.n163 4.5005
R983 VDDA.n165 VDDA.n51 4.5005
R984 VDDA.n167 VDDA.n166 4.5005
R985 VDDA.n168 VDDA.n50 4.5005
R986 VDDA.n172 VDDA.n171 4.5005
R987 VDDA.n173 VDDA.n47 4.5005
R988 VDDA.n175 VDDA.n174 4.5005
R989 VDDA.n176 VDDA.n46 4.5005
R990 VDDA.n180 VDDA.n179 4.5005
R991 VDDA.n181 VDDA.n45 4.5005
R992 VDDA.n2945 VDDA.n2944 4.5005
R993 VDDA.n2814 VDDA.n2813 4.5005
R994 VDDA.n2824 VDDA.n2823 4.5005
R995 VDDA.n2825 VDDA.n2812 4.5005
R996 VDDA.n2827 VDDA.n2826 4.5005
R997 VDDA.n2810 VDDA.n2809 4.5005
R998 VDDA.n2834 VDDA.n2833 4.5005
R999 VDDA.n2835 VDDA.n2808 4.5005
R1000 VDDA.n2837 VDDA.n2836 4.5005
R1001 VDDA.n2806 VDDA.n2805 4.5005
R1002 VDDA.n2844 VDDA.n2843 4.5005
R1003 VDDA.n2845 VDDA.n2804 4.5005
R1004 VDDA.n2847 VDDA.n2846 4.5005
R1005 VDDA.n2802 VDDA.n2801 4.5005
R1006 VDDA.n2854 VDDA.n2853 4.5005
R1007 VDDA.n2855 VDDA.n2800 4.5005
R1008 VDDA.n2857 VDDA.n2856 4.5005
R1009 VDDA.n2798 VDDA.n2797 4.5005
R1010 VDDA.n2864 VDDA.n2863 4.5005
R1011 VDDA.n2865 VDDA.n2796 4.5005
R1012 VDDA.n2867 VDDA.n2866 4.5005
R1013 VDDA.n2794 VDDA.n2793 4.5005
R1014 VDDA.n2874 VDDA.n2873 4.5005
R1015 VDDA.n2875 VDDA.n2792 4.5005
R1016 VDDA.n2877 VDDA.n2876 4.5005
R1017 VDDA.n2790 VDDA.n2789 4.5005
R1018 VDDA.n2884 VDDA.n2883 4.5005
R1019 VDDA.n2885 VDDA.n2788 4.5005
R1020 VDDA.n2887 VDDA.n2886 4.5005
R1021 VDDA.n2786 VDDA.n2785 4.5005
R1022 VDDA.n2894 VDDA.n2893 4.5005
R1023 VDDA.n2895 VDDA.n2784 4.5005
R1024 VDDA.n2897 VDDA.n2896 4.5005
R1025 VDDA.n2782 VDDA.n2781 4.5005
R1026 VDDA.n2904 VDDA.n2903 4.5005
R1027 VDDA.n2905 VDDA.n2780 4.5005
R1028 VDDA.n2907 VDDA.n2906 4.5005
R1029 VDDA.n2778 VDDA.n2777 4.5005
R1030 VDDA.n2914 VDDA.n2913 4.5005
R1031 VDDA.n2915 VDDA.n2776 4.5005
R1032 VDDA.n2917 VDDA.n2916 4.5005
R1033 VDDA.n2774 VDDA.n2773 4.5005
R1034 VDDA.n2924 VDDA.n2923 4.5005
R1035 VDDA.n2925 VDDA.n2772 4.5005
R1036 VDDA.n2927 VDDA.n2926 4.5005
R1037 VDDA.n2770 VDDA.n2769 4.5005
R1038 VDDA.n2933 VDDA.n2932 4.5005
R1039 VDDA.n2669 VDDA.n2665 4.5005
R1040 VDDA.n2673 VDDA.n2672 4.5005
R1041 VDDA.n2674 VDDA.n2662 4.5005
R1042 VDDA.n2676 VDDA.n2675 4.5005
R1043 VDDA.n2677 VDDA.n2661 4.5005
R1044 VDDA.n2681 VDDA.n2680 4.5005
R1045 VDDA.n2682 VDDA.n2658 4.5005
R1046 VDDA.n2684 VDDA.n2683 4.5005
R1047 VDDA.n2685 VDDA.n2657 4.5005
R1048 VDDA.n2689 VDDA.n2688 4.5005
R1049 VDDA.n2690 VDDA.n2654 4.5005
R1050 VDDA.n2692 VDDA.n2691 4.5005
R1051 VDDA.n2693 VDDA.n2653 4.5005
R1052 VDDA.n2697 VDDA.n2696 4.5005
R1053 VDDA.n2698 VDDA.n2650 4.5005
R1054 VDDA.n2700 VDDA.n2699 4.5005
R1055 VDDA.n2701 VDDA.n2649 4.5005
R1056 VDDA.n2705 VDDA.n2704 4.5005
R1057 VDDA.n2706 VDDA.n2646 4.5005
R1058 VDDA.n2708 VDDA.n2707 4.5005
R1059 VDDA.n2709 VDDA.n2645 4.5005
R1060 VDDA.n2713 VDDA.n2712 4.5005
R1061 VDDA.n2714 VDDA.n2642 4.5005
R1062 VDDA.n2716 VDDA.n2715 4.5005
R1063 VDDA.n2717 VDDA.n2641 4.5005
R1064 VDDA.n2721 VDDA.n2720 4.5005
R1065 VDDA.n2722 VDDA.n2638 4.5005
R1066 VDDA.n2724 VDDA.n2723 4.5005
R1067 VDDA.n2725 VDDA.n2637 4.5005
R1068 VDDA.n2729 VDDA.n2728 4.5005
R1069 VDDA.n2730 VDDA.n2634 4.5005
R1070 VDDA.n2732 VDDA.n2731 4.5005
R1071 VDDA.n2733 VDDA.n2633 4.5005
R1072 VDDA.n2737 VDDA.n2736 4.5005
R1073 VDDA.n2738 VDDA.n2630 4.5005
R1074 VDDA.n2740 VDDA.n2739 4.5005
R1075 VDDA.n2741 VDDA.n2629 4.5005
R1076 VDDA.n2745 VDDA.n2744 4.5005
R1077 VDDA.n2746 VDDA.n2626 4.5005
R1078 VDDA.n2748 VDDA.n2747 4.5005
R1079 VDDA.n2749 VDDA.n2625 4.5005
R1080 VDDA.n2753 VDDA.n2752 4.5005
R1081 VDDA.n2754 VDDA.n2624 4.5005
R1082 VDDA.n2756 VDDA.n2755 4.5005
R1083 VDDA.n195 VDDA.n194 4.5005
R1084 VDDA.n2762 VDDA.n2761 4.5005
R1085 VDDA.n271 VDDA.n265 4.5005
R1086 VDDA.n273 VDDA.n272 4.5005
R1087 VDDA.n274 VDDA.n264 4.5005
R1088 VDDA.n278 VDDA.n277 4.5005
R1089 VDDA.n279 VDDA.n261 4.5005
R1090 VDDA.n281 VDDA.n280 4.5005
R1091 VDDA.n282 VDDA.n260 4.5005
R1092 VDDA.n286 VDDA.n285 4.5005
R1093 VDDA.n287 VDDA.n257 4.5005
R1094 VDDA.n289 VDDA.n288 4.5005
R1095 VDDA.n290 VDDA.n256 4.5005
R1096 VDDA.n294 VDDA.n293 4.5005
R1097 VDDA.n295 VDDA.n253 4.5005
R1098 VDDA.n297 VDDA.n296 4.5005
R1099 VDDA.n298 VDDA.n252 4.5005
R1100 VDDA.n302 VDDA.n301 4.5005
R1101 VDDA.n303 VDDA.n249 4.5005
R1102 VDDA.n305 VDDA.n304 4.5005
R1103 VDDA.n306 VDDA.n248 4.5005
R1104 VDDA.n310 VDDA.n309 4.5005
R1105 VDDA.n311 VDDA.n245 4.5005
R1106 VDDA.n313 VDDA.n312 4.5005
R1107 VDDA.n314 VDDA.n244 4.5005
R1108 VDDA.n318 VDDA.n317 4.5005
R1109 VDDA.n319 VDDA.n241 4.5005
R1110 VDDA.n321 VDDA.n320 4.5005
R1111 VDDA.n322 VDDA.n240 4.5005
R1112 VDDA.n326 VDDA.n325 4.5005
R1113 VDDA.n327 VDDA.n237 4.5005
R1114 VDDA.n329 VDDA.n328 4.5005
R1115 VDDA.n330 VDDA.n236 4.5005
R1116 VDDA.n334 VDDA.n333 4.5005
R1117 VDDA.n335 VDDA.n233 4.5005
R1118 VDDA.n337 VDDA.n336 4.5005
R1119 VDDA.n338 VDDA.n232 4.5005
R1120 VDDA.n342 VDDA.n341 4.5005
R1121 VDDA.n343 VDDA.n229 4.5005
R1122 VDDA.n345 VDDA.n344 4.5005
R1123 VDDA.n346 VDDA.n228 4.5005
R1124 VDDA.n350 VDDA.n349 4.5005
R1125 VDDA.n351 VDDA.n225 4.5005
R1126 VDDA.n353 VDDA.n352 4.5005
R1127 VDDA.n354 VDDA.n224 4.5005
R1128 VDDA.n358 VDDA.n357 4.5005
R1129 VDDA.n359 VDDA.n223 4.5005
R1130 VDDA.n2597 VDDA.n2596 4.5005
R1131 VDDA.n2466 VDDA.n2465 4.5005
R1132 VDDA.n2476 VDDA.n2475 4.5005
R1133 VDDA.n2477 VDDA.n2464 4.5005
R1134 VDDA.n2479 VDDA.n2478 4.5005
R1135 VDDA.n2462 VDDA.n2461 4.5005
R1136 VDDA.n2486 VDDA.n2485 4.5005
R1137 VDDA.n2487 VDDA.n2460 4.5005
R1138 VDDA.n2489 VDDA.n2488 4.5005
R1139 VDDA.n2458 VDDA.n2457 4.5005
R1140 VDDA.n2496 VDDA.n2495 4.5005
R1141 VDDA.n2497 VDDA.n2456 4.5005
R1142 VDDA.n2499 VDDA.n2498 4.5005
R1143 VDDA.n2454 VDDA.n2453 4.5005
R1144 VDDA.n2506 VDDA.n2505 4.5005
R1145 VDDA.n2507 VDDA.n2452 4.5005
R1146 VDDA.n2509 VDDA.n2508 4.5005
R1147 VDDA.n2450 VDDA.n2449 4.5005
R1148 VDDA.n2516 VDDA.n2515 4.5005
R1149 VDDA.n2517 VDDA.n2448 4.5005
R1150 VDDA.n2519 VDDA.n2518 4.5005
R1151 VDDA.n2446 VDDA.n2445 4.5005
R1152 VDDA.n2526 VDDA.n2525 4.5005
R1153 VDDA.n2527 VDDA.n2444 4.5005
R1154 VDDA.n2529 VDDA.n2528 4.5005
R1155 VDDA.n2442 VDDA.n2441 4.5005
R1156 VDDA.n2536 VDDA.n2535 4.5005
R1157 VDDA.n2537 VDDA.n2440 4.5005
R1158 VDDA.n2539 VDDA.n2538 4.5005
R1159 VDDA.n2438 VDDA.n2437 4.5005
R1160 VDDA.n2546 VDDA.n2545 4.5005
R1161 VDDA.n2547 VDDA.n2436 4.5005
R1162 VDDA.n2549 VDDA.n2548 4.5005
R1163 VDDA.n2434 VDDA.n2433 4.5005
R1164 VDDA.n2556 VDDA.n2555 4.5005
R1165 VDDA.n2557 VDDA.n2432 4.5005
R1166 VDDA.n2559 VDDA.n2558 4.5005
R1167 VDDA.n2430 VDDA.n2429 4.5005
R1168 VDDA.n2566 VDDA.n2565 4.5005
R1169 VDDA.n2567 VDDA.n2428 4.5005
R1170 VDDA.n2569 VDDA.n2568 4.5005
R1171 VDDA.n2426 VDDA.n2425 4.5005
R1172 VDDA.n2576 VDDA.n2575 4.5005
R1173 VDDA.n2577 VDDA.n2424 4.5005
R1174 VDDA.n2579 VDDA.n2578 4.5005
R1175 VDDA.n2422 VDDA.n2421 4.5005
R1176 VDDA.n2585 VDDA.n2584 4.5005
R1177 VDDA.n1231 VDDA.n1227 4.5005
R1178 VDDA.n1235 VDDA.n1234 4.5005
R1179 VDDA.n1236 VDDA.n1224 4.5005
R1180 VDDA.n1238 VDDA.n1237 4.5005
R1181 VDDA.n1239 VDDA.n1223 4.5005
R1182 VDDA.n1243 VDDA.n1242 4.5005
R1183 VDDA.n1244 VDDA.n1220 4.5005
R1184 VDDA.n1246 VDDA.n1245 4.5005
R1185 VDDA.n1247 VDDA.n1219 4.5005
R1186 VDDA.n1251 VDDA.n1250 4.5005
R1187 VDDA.n1252 VDDA.n1216 4.5005
R1188 VDDA.n1254 VDDA.n1253 4.5005
R1189 VDDA.n1255 VDDA.n1215 4.5005
R1190 VDDA.n1259 VDDA.n1258 4.5005
R1191 VDDA.n1260 VDDA.n1212 4.5005
R1192 VDDA.n1262 VDDA.n1261 4.5005
R1193 VDDA.n1263 VDDA.n1211 4.5005
R1194 VDDA.n1267 VDDA.n1266 4.5005
R1195 VDDA.n1268 VDDA.n1208 4.5005
R1196 VDDA.n1270 VDDA.n1269 4.5005
R1197 VDDA.n1271 VDDA.n1207 4.5005
R1198 VDDA.n1275 VDDA.n1274 4.5005
R1199 VDDA.n1276 VDDA.n1204 4.5005
R1200 VDDA.n1278 VDDA.n1277 4.5005
R1201 VDDA.n1279 VDDA.n1203 4.5005
R1202 VDDA.n1283 VDDA.n1282 4.5005
R1203 VDDA.n1284 VDDA.n1200 4.5005
R1204 VDDA.n1286 VDDA.n1285 4.5005
R1205 VDDA.n1287 VDDA.n1199 4.5005
R1206 VDDA.n1291 VDDA.n1290 4.5005
R1207 VDDA.n1292 VDDA.n1196 4.5005
R1208 VDDA.n1294 VDDA.n1293 4.5005
R1209 VDDA.n1295 VDDA.n1195 4.5005
R1210 VDDA.n1299 VDDA.n1298 4.5005
R1211 VDDA.n1300 VDDA.n1192 4.5005
R1212 VDDA.n1302 VDDA.n1301 4.5005
R1213 VDDA.n1303 VDDA.n1191 4.5005
R1214 VDDA.n1307 VDDA.n1306 4.5005
R1215 VDDA.n1308 VDDA.n1188 4.5005
R1216 VDDA.n1310 VDDA.n1309 4.5005
R1217 VDDA.n1311 VDDA.n1187 4.5005
R1218 VDDA.n1315 VDDA.n1314 4.5005
R1219 VDDA.n1316 VDDA.n1186 4.5005
R1220 VDDA.n1318 VDDA.n1317 4.5005
R1221 VDDA.n462 VDDA.n461 4.5005
R1222 VDDA.n2261 VDDA.n2260 4.5005
R1223 VDDA.n2413 VDDA.n2412 4.5005
R1224 VDDA.n409 VDDA.n408 4.5005
R1225 VDDA.n412 VDDA.n411 4.5005
R1226 VDDA.n2394 VDDA.n389 4.5005
R1227 VDDA.n2396 VDDA.n2395 4.5005
R1228 VDDA.n2395 VDDA.n2394 4.5005
R1229 VDDA.n2290 VDDA.n450 4.5005
R1230 VDDA.n2308 VDDA.n2307 4.5005
R1231 VDDA.n2311 VDDA.n2310 4.5005
R1232 VDDA.n2272 VDDA.n2271 4.5005
R1233 VDDA.n538 VDDA.n532 4.5005
R1234 VDDA.n540 VDDA.n539 4.5005
R1235 VDDA.n541 VDDA.n531 4.5005
R1236 VDDA.n545 VDDA.n544 4.5005
R1237 VDDA.n546 VDDA.n528 4.5005
R1238 VDDA.n548 VDDA.n547 4.5005
R1239 VDDA.n549 VDDA.n527 4.5005
R1240 VDDA.n553 VDDA.n552 4.5005
R1241 VDDA.n554 VDDA.n524 4.5005
R1242 VDDA.n556 VDDA.n555 4.5005
R1243 VDDA.n557 VDDA.n523 4.5005
R1244 VDDA.n561 VDDA.n560 4.5005
R1245 VDDA.n562 VDDA.n520 4.5005
R1246 VDDA.n564 VDDA.n563 4.5005
R1247 VDDA.n565 VDDA.n519 4.5005
R1248 VDDA.n569 VDDA.n568 4.5005
R1249 VDDA.n570 VDDA.n516 4.5005
R1250 VDDA.n572 VDDA.n571 4.5005
R1251 VDDA.n573 VDDA.n515 4.5005
R1252 VDDA.n577 VDDA.n576 4.5005
R1253 VDDA.n578 VDDA.n512 4.5005
R1254 VDDA.n580 VDDA.n579 4.5005
R1255 VDDA.n581 VDDA.n511 4.5005
R1256 VDDA.n585 VDDA.n584 4.5005
R1257 VDDA.n586 VDDA.n508 4.5005
R1258 VDDA.n588 VDDA.n587 4.5005
R1259 VDDA.n589 VDDA.n507 4.5005
R1260 VDDA.n593 VDDA.n592 4.5005
R1261 VDDA.n594 VDDA.n504 4.5005
R1262 VDDA.n596 VDDA.n595 4.5005
R1263 VDDA.n597 VDDA.n503 4.5005
R1264 VDDA.n601 VDDA.n600 4.5005
R1265 VDDA.n602 VDDA.n500 4.5005
R1266 VDDA.n604 VDDA.n603 4.5005
R1267 VDDA.n605 VDDA.n499 4.5005
R1268 VDDA.n609 VDDA.n608 4.5005
R1269 VDDA.n610 VDDA.n496 4.5005
R1270 VDDA.n612 VDDA.n611 4.5005
R1271 VDDA.n613 VDDA.n495 4.5005
R1272 VDDA.n617 VDDA.n616 4.5005
R1273 VDDA.n618 VDDA.n492 4.5005
R1274 VDDA.n620 VDDA.n619 4.5005
R1275 VDDA.n621 VDDA.n491 4.5005
R1276 VDDA.n625 VDDA.n624 4.5005
R1277 VDDA.n626 VDDA.n490 4.5005
R1278 VDDA.n1159 VDDA.n1158 4.5005
R1279 VDDA.n1028 VDDA.n1027 4.5005
R1280 VDDA.n1038 VDDA.n1037 4.5005
R1281 VDDA.n1039 VDDA.n1026 4.5005
R1282 VDDA.n1041 VDDA.n1040 4.5005
R1283 VDDA.n1024 VDDA.n1023 4.5005
R1284 VDDA.n1048 VDDA.n1047 4.5005
R1285 VDDA.n1049 VDDA.n1022 4.5005
R1286 VDDA.n1051 VDDA.n1050 4.5005
R1287 VDDA.n1020 VDDA.n1019 4.5005
R1288 VDDA.n1058 VDDA.n1057 4.5005
R1289 VDDA.n1059 VDDA.n1018 4.5005
R1290 VDDA.n1061 VDDA.n1060 4.5005
R1291 VDDA.n1016 VDDA.n1015 4.5005
R1292 VDDA.n1068 VDDA.n1067 4.5005
R1293 VDDA.n1069 VDDA.n1014 4.5005
R1294 VDDA.n1071 VDDA.n1070 4.5005
R1295 VDDA.n1012 VDDA.n1011 4.5005
R1296 VDDA.n1078 VDDA.n1077 4.5005
R1297 VDDA.n1079 VDDA.n1010 4.5005
R1298 VDDA.n1081 VDDA.n1080 4.5005
R1299 VDDA.n1008 VDDA.n1007 4.5005
R1300 VDDA.n1088 VDDA.n1087 4.5005
R1301 VDDA.n1089 VDDA.n1006 4.5005
R1302 VDDA.n1091 VDDA.n1090 4.5005
R1303 VDDA.n1004 VDDA.n1003 4.5005
R1304 VDDA.n1098 VDDA.n1097 4.5005
R1305 VDDA.n1099 VDDA.n1002 4.5005
R1306 VDDA.n1101 VDDA.n1100 4.5005
R1307 VDDA.n1000 VDDA.n999 4.5005
R1308 VDDA.n1108 VDDA.n1107 4.5005
R1309 VDDA.n1109 VDDA.n998 4.5005
R1310 VDDA.n1111 VDDA.n1110 4.5005
R1311 VDDA.n996 VDDA.n995 4.5005
R1312 VDDA.n1118 VDDA.n1117 4.5005
R1313 VDDA.n1119 VDDA.n994 4.5005
R1314 VDDA.n1121 VDDA.n1120 4.5005
R1315 VDDA.n992 VDDA.n991 4.5005
R1316 VDDA.n1128 VDDA.n1127 4.5005
R1317 VDDA.n1129 VDDA.n990 4.5005
R1318 VDDA.n1131 VDDA.n1130 4.5005
R1319 VDDA.n988 VDDA.n987 4.5005
R1320 VDDA.n1138 VDDA.n1137 4.5005
R1321 VDDA.n1139 VDDA.n986 4.5005
R1322 VDDA.n1141 VDDA.n1140 4.5005
R1323 VDDA.n984 VDDA.n983 4.5005
R1324 VDDA.n1147 VDDA.n1146 4.5005
R1325 VDDA.n883 VDDA.n879 4.5005
R1326 VDDA.n887 VDDA.n886 4.5005
R1327 VDDA.n888 VDDA.n876 4.5005
R1328 VDDA.n890 VDDA.n889 4.5005
R1329 VDDA.n891 VDDA.n875 4.5005
R1330 VDDA.n895 VDDA.n894 4.5005
R1331 VDDA.n896 VDDA.n872 4.5005
R1332 VDDA.n898 VDDA.n897 4.5005
R1333 VDDA.n899 VDDA.n871 4.5005
R1334 VDDA.n903 VDDA.n902 4.5005
R1335 VDDA.n904 VDDA.n868 4.5005
R1336 VDDA.n906 VDDA.n905 4.5005
R1337 VDDA.n907 VDDA.n867 4.5005
R1338 VDDA.n911 VDDA.n910 4.5005
R1339 VDDA.n912 VDDA.n864 4.5005
R1340 VDDA.n914 VDDA.n913 4.5005
R1341 VDDA.n915 VDDA.n863 4.5005
R1342 VDDA.n919 VDDA.n918 4.5005
R1343 VDDA.n920 VDDA.n860 4.5005
R1344 VDDA.n922 VDDA.n921 4.5005
R1345 VDDA.n923 VDDA.n859 4.5005
R1346 VDDA.n927 VDDA.n926 4.5005
R1347 VDDA.n928 VDDA.n856 4.5005
R1348 VDDA.n930 VDDA.n929 4.5005
R1349 VDDA.n931 VDDA.n855 4.5005
R1350 VDDA.n935 VDDA.n934 4.5005
R1351 VDDA.n936 VDDA.n852 4.5005
R1352 VDDA.n938 VDDA.n937 4.5005
R1353 VDDA.n939 VDDA.n851 4.5005
R1354 VDDA.n943 VDDA.n942 4.5005
R1355 VDDA.n944 VDDA.n848 4.5005
R1356 VDDA.n946 VDDA.n945 4.5005
R1357 VDDA.n947 VDDA.n847 4.5005
R1358 VDDA.n951 VDDA.n950 4.5005
R1359 VDDA.n952 VDDA.n844 4.5005
R1360 VDDA.n954 VDDA.n953 4.5005
R1361 VDDA.n955 VDDA.n843 4.5005
R1362 VDDA.n959 VDDA.n958 4.5005
R1363 VDDA.n960 VDDA.n840 4.5005
R1364 VDDA.n962 VDDA.n961 4.5005
R1365 VDDA.n963 VDDA.n839 4.5005
R1366 VDDA.n967 VDDA.n966 4.5005
R1367 VDDA.n968 VDDA.n838 4.5005
R1368 VDDA.n970 VDDA.n969 4.5005
R1369 VDDA.n639 VDDA.n638 4.5005
R1370 VDDA.n976 VDDA.n975 4.5005
R1371 VDDA.n979 VDDA.n637 4.5005
R1372 VDDA.n981 VDDA.n980 4.5005
R1373 VDDA.n980 VDDA.n979 4.5005
R1374 VDDA.n1150 VDDA.n982 4.5005
R1375 VDDA.n1152 VDDA.n1151 4.5005
R1376 VDDA.n1151 VDDA.n1150 4.5005
R1377 VDDA.n1155 VDDA.n1154 4.5005
R1378 VDDA.n1153 VDDA.n459 4.5005
R1379 VDDA.n1154 VDDA.n1153 4.5005
R1380 VDDA.n2288 VDDA.n2284 4.5005
R1381 VDDA.n2289 VDDA.n452 4.5005
R1382 VDDA.n2289 VDDA.n2288 4.5005
R1383 VDDA.n2403 VDDA.n2402 4.5005
R1384 VDDA.n2402 VDDA.n2401 4.5005
R1385 VDDA.n2401 VDDA.n387 4.5005
R1386 VDDA.n2264 VDDA.n460 4.5005
R1387 VDDA.n2266 VDDA.n2265 4.5005
R1388 VDDA.n2265 VDDA.n2264 4.5005
R1389 VDDA.n2588 VDDA.n2420 4.5005
R1390 VDDA.n2590 VDDA.n2589 4.5005
R1391 VDDA.n2589 VDDA.n2588 4.5005
R1392 VDDA.n2593 VDDA.n2592 4.5005
R1393 VDDA.n2591 VDDA.n192 4.5005
R1394 VDDA.n2592 VDDA.n2591 4.5005
R1395 VDDA.n2765 VDDA.n193 4.5005
R1396 VDDA.n2767 VDDA.n2766 4.5005
R1397 VDDA.n2766 VDDA.n2765 4.5005
R1398 VDDA.n2936 VDDA.n2768 4.5005
R1399 VDDA.n2938 VDDA.n2937 4.5005
R1400 VDDA.n2937 VDDA.n2936 4.5005
R1401 VDDA.n2939 VDDA.n183 4.5005
R1402 VDDA.n2941 VDDA.n2940 4.5005
R1403 VDDA.n2940 VDDA.n2939 4.5005
R1404 VDDA.n807 VDDA.n804 4.5005
R1405 VDDA.n692 VDDA.n688 4.5005
R1406 VDDA.n696 VDDA.n693 4.5005
R1407 VDDA.n697 VDDA.n687 4.5005
R1408 VDDA.n701 VDDA.n700 4.5005
R1409 VDDA.n702 VDDA.n686 4.5005
R1410 VDDA.n706 VDDA.n703 4.5005
R1411 VDDA.n707 VDDA.n685 4.5005
R1412 VDDA.n711 VDDA.n710 4.5005
R1413 VDDA.n712 VDDA.n684 4.5005
R1414 VDDA.n716 VDDA.n713 4.5005
R1415 VDDA.n717 VDDA.n683 4.5005
R1416 VDDA.n721 VDDA.n720 4.5005
R1417 VDDA.n722 VDDA.n682 4.5005
R1418 VDDA.n726 VDDA.n723 4.5005
R1419 VDDA.n727 VDDA.n681 4.5005
R1420 VDDA.n731 VDDA.n730 4.5005
R1421 VDDA.n732 VDDA.n680 4.5005
R1422 VDDA.n736 VDDA.n733 4.5005
R1423 VDDA.n737 VDDA.n679 4.5005
R1424 VDDA.n741 VDDA.n740 4.5005
R1425 VDDA.n742 VDDA.n678 4.5005
R1426 VDDA.n746 VDDA.n743 4.5005
R1427 VDDA.n747 VDDA.n677 4.5005
R1428 VDDA.n751 VDDA.n750 4.5005
R1429 VDDA.n752 VDDA.n676 4.5005
R1430 VDDA.n756 VDDA.n753 4.5005
R1431 VDDA.n757 VDDA.n675 4.5005
R1432 VDDA.n761 VDDA.n760 4.5005
R1433 VDDA.n762 VDDA.n674 4.5005
R1434 VDDA.n766 VDDA.n763 4.5005
R1435 VDDA.n767 VDDA.n673 4.5005
R1436 VDDA.n771 VDDA.n770 4.5005
R1437 VDDA.n772 VDDA.n672 4.5005
R1438 VDDA.n776 VDDA.n773 4.5005
R1439 VDDA.n777 VDDA.n671 4.5005
R1440 VDDA.n781 VDDA.n780 4.5005
R1441 VDDA.n782 VDDA.n670 4.5005
R1442 VDDA.n786 VDDA.n783 4.5005
R1443 VDDA.n787 VDDA.n669 4.5005
R1444 VDDA.n791 VDDA.n790 4.5005
R1445 VDDA.n792 VDDA.n668 4.5005
R1446 VDDA.n796 VDDA.n793 4.5005
R1447 VDDA.n797 VDDA.n667 4.5005
R1448 VDDA.n801 VDDA.n800 4.5005
R1449 VDDA.n802 VDDA.n666 4.5005
R1450 VDDA.n811 VDDA.n810 4.5005
R1451 VDDA.n1996 VDDA.n1995 4.48641
R1452 VDDA.n1995 VDDA.n1973 4.48641
R1453 VDDA.n2006 VDDA.n2005 4.48641
R1454 VDDA.n2005 VDDA.n1953 4.48641
R1455 VDDA.n1774 VDDA.n1401 3.75335
R1456 VDDA.n1773 VDDA.n1772 3.75335
R1457 VDDA.n1781 VDDA.n1779 3.75335
R1458 VDDA.n1780 VDDA.n1395 3.75335
R1459 VDDA.n2065 VDDA.n2056 3.75335
R1460 VDDA.n2059 VDDA.n2026 3.75335
R1461 VDDA.n2047 VDDA.n2033 3.75335
R1462 VDDA.n2039 VDDA.n2038 3.75335
R1463 VDDA.n1907 VDDA.n1906 3.48486
R1464 VDDA.n1579 VDDA.n1578 3.47821
R1465 VDDA.n2256 VDDA.n2255 3.47821
R1466 VDDA.n92 VDDA.n20 3.47821
R1467 VDDA.n2816 VDDA.n2815 3.47821
R1468 VDDA.n2666 VDDA.n2600 3.47821
R1469 VDDA.n270 VDDA.n198 3.47821
R1470 VDDA.n2468 VDDA.n2467 3.47821
R1471 VDDA.n1228 VDDA.n1162 3.47821
R1472 VDDA.n537 VDDA.n465 3.47821
R1473 VDDA.n1030 VDDA.n1029 3.47821
R1474 VDDA.n880 VDDA.n814 3.47821
R1475 VDDA.n691 VDDA.n641 3.47821
R1476 VDDA.n1992 VDDA.n1991 3.41464
R1477 VDDA.n2002 VDDA.n2001 3.41464
R1478 VDDA.n1370 VDDA.n1369 3.4105
R1479 VDDA.n1904 VDDA.n1903 3.4105
R1480 VDDA.n1902 VDDA.n1901 3.4105
R1481 VDDA.n1900 VDDA.n1899 3.4105
R1482 VDDA.n1898 VDDA.n1372 3.4105
R1483 VDDA.n1894 VDDA.n1893 3.4105
R1484 VDDA.n1892 VDDA.n1891 3.4105
R1485 VDDA.n1890 VDDA.n1889 3.4105
R1486 VDDA.n1888 VDDA.n1374 3.4105
R1487 VDDA.n1884 VDDA.n1883 3.4105
R1488 VDDA.n1882 VDDA.n1881 3.4105
R1489 VDDA.n1880 VDDA.n1879 3.4105
R1490 VDDA.n1878 VDDA.n1376 3.4105
R1491 VDDA.n1874 VDDA.n1873 3.4105
R1492 VDDA.n1872 VDDA.n1871 3.4105
R1493 VDDA.n1870 VDDA.n1869 3.4105
R1494 VDDA.n1868 VDDA.n1378 3.4105
R1495 VDDA.n1864 VDDA.n1863 3.4105
R1496 VDDA.n1862 VDDA.n1861 3.4105
R1497 VDDA.n1860 VDDA.n1859 3.4105
R1498 VDDA.n1858 VDDA.n1380 3.4105
R1499 VDDA.n1854 VDDA.n1853 3.4105
R1500 VDDA.n1852 VDDA.n1851 3.4105
R1501 VDDA.n1850 VDDA.n1849 3.4105
R1502 VDDA.n1848 VDDA.n1382 3.4105
R1503 VDDA.n1844 VDDA.n1843 3.4105
R1504 VDDA.n1842 VDDA.n1841 3.4105
R1505 VDDA.n1840 VDDA.n1839 3.4105
R1506 VDDA.n1838 VDDA.n1384 3.4105
R1507 VDDA.n1834 VDDA.n1833 3.4105
R1508 VDDA.n1832 VDDA.n1831 3.4105
R1509 VDDA.n1830 VDDA.n1829 3.4105
R1510 VDDA.n1828 VDDA.n1386 3.4105
R1511 VDDA.n1824 VDDA.n1823 3.4105
R1512 VDDA.n1822 VDDA.n1821 3.4105
R1513 VDDA.n1820 VDDA.n1819 3.4105
R1514 VDDA.n1818 VDDA.n1388 3.4105
R1515 VDDA.n1814 VDDA.n1813 3.4105
R1516 VDDA.n1812 VDDA.n1811 3.4105
R1517 VDDA.n1810 VDDA.n1809 3.4105
R1518 VDDA.n1808 VDDA.n1390 3.4105
R1519 VDDA.n1804 VDDA.n1803 3.4105
R1520 VDDA.n1802 VDDA.n1801 3.4105
R1521 VDDA.n1800 VDDA.n1799 3.4105
R1522 VDDA.n1798 VDDA.n1392 3.4105
R1523 VDDA.n1794 VDDA.n1793 3.4105
R1524 VDDA.n1792 VDDA.n1344 3.4105
R1525 VDDA.n1435 VDDA.n1434 3.4105
R1526 VDDA.n1576 VDDA.n1575 3.4105
R1527 VDDA.n1574 VDDA.n1573 3.4105
R1528 VDDA.n1572 VDDA.n1571 3.4105
R1529 VDDA.n1570 VDDA.n1437 3.4105
R1530 VDDA.n1566 VDDA.n1565 3.4105
R1531 VDDA.n1564 VDDA.n1563 3.4105
R1532 VDDA.n1562 VDDA.n1561 3.4105
R1533 VDDA.n1560 VDDA.n1439 3.4105
R1534 VDDA.n1556 VDDA.n1555 3.4105
R1535 VDDA.n1554 VDDA.n1553 3.4105
R1536 VDDA.n1552 VDDA.n1551 3.4105
R1537 VDDA.n1550 VDDA.n1441 3.4105
R1538 VDDA.n1546 VDDA.n1545 3.4105
R1539 VDDA.n1544 VDDA.n1543 3.4105
R1540 VDDA.n1542 VDDA.n1541 3.4105
R1541 VDDA.n1540 VDDA.n1443 3.4105
R1542 VDDA.n1536 VDDA.n1535 3.4105
R1543 VDDA.n1534 VDDA.n1533 3.4105
R1544 VDDA.n1532 VDDA.n1531 3.4105
R1545 VDDA.n1530 VDDA.n1445 3.4105
R1546 VDDA.n1526 VDDA.n1525 3.4105
R1547 VDDA.n1524 VDDA.n1523 3.4105
R1548 VDDA.n1522 VDDA.n1521 3.4105
R1549 VDDA.n1520 VDDA.n1447 3.4105
R1550 VDDA.n1516 VDDA.n1515 3.4105
R1551 VDDA.n1514 VDDA.n1513 3.4105
R1552 VDDA.n1512 VDDA.n1511 3.4105
R1553 VDDA.n1510 VDDA.n1449 3.4105
R1554 VDDA.n1506 VDDA.n1505 3.4105
R1555 VDDA.n1504 VDDA.n1503 3.4105
R1556 VDDA.n1502 VDDA.n1501 3.4105
R1557 VDDA.n1500 VDDA.n1451 3.4105
R1558 VDDA.n1496 VDDA.n1495 3.4105
R1559 VDDA.n1494 VDDA.n1493 3.4105
R1560 VDDA.n1492 VDDA.n1491 3.4105
R1561 VDDA.n1490 VDDA.n1453 3.4105
R1562 VDDA.n1486 VDDA.n1485 3.4105
R1563 VDDA.n1484 VDDA.n1483 3.4105
R1564 VDDA.n1482 VDDA.n1481 3.4105
R1565 VDDA.n1480 VDDA.n1455 3.4105
R1566 VDDA.n1476 VDDA.n1475 3.4105
R1567 VDDA.n1474 VDDA.n1473 3.4105
R1568 VDDA.n1472 VDDA.n1471 3.4105
R1569 VDDA.n1470 VDDA.n1457 3.4105
R1570 VDDA.n1466 VDDA.n1465 3.4105
R1571 VDDA.n1464 VDDA.n1410 3.4105
R1572 VDDA.n1910 VDDA.n1909 3.4105
R1573 VDDA.n2253 VDDA.n2252 3.4105
R1574 VDDA.n2251 VDDA.n2250 3.4105
R1575 VDDA.n2249 VDDA.n2248 3.4105
R1576 VDDA.n2247 VDDA.n1912 3.4105
R1577 VDDA.n2243 VDDA.n2242 3.4105
R1578 VDDA.n2241 VDDA.n2240 3.4105
R1579 VDDA.n2239 VDDA.n2238 3.4105
R1580 VDDA.n2237 VDDA.n1914 3.4105
R1581 VDDA.n2233 VDDA.n2232 3.4105
R1582 VDDA.n2231 VDDA.n2230 3.4105
R1583 VDDA.n2229 VDDA.n2228 3.4105
R1584 VDDA.n2227 VDDA.n1916 3.4105
R1585 VDDA.n2223 VDDA.n2222 3.4105
R1586 VDDA.n2221 VDDA.n2220 3.4105
R1587 VDDA.n2219 VDDA.n2218 3.4105
R1588 VDDA.n2217 VDDA.n1918 3.4105
R1589 VDDA.n2213 VDDA.n2212 3.4105
R1590 VDDA.n2211 VDDA.n2210 3.4105
R1591 VDDA.n2209 VDDA.n2208 3.4105
R1592 VDDA.n2207 VDDA.n1920 3.4105
R1593 VDDA.n2203 VDDA.n2202 3.4105
R1594 VDDA.n2201 VDDA.n2200 3.4105
R1595 VDDA.n2199 VDDA.n2198 3.4105
R1596 VDDA.n2197 VDDA.n1922 3.4105
R1597 VDDA.n2193 VDDA.n2192 3.4105
R1598 VDDA.n2191 VDDA.n2190 3.4105
R1599 VDDA.n2189 VDDA.n2188 3.4105
R1600 VDDA.n2187 VDDA.n1924 3.4105
R1601 VDDA.n2183 VDDA.n2182 3.4105
R1602 VDDA.n2181 VDDA.n2180 3.4105
R1603 VDDA.n2179 VDDA.n2178 3.4105
R1604 VDDA.n2177 VDDA.n1926 3.4105
R1605 VDDA.n2173 VDDA.n2172 3.4105
R1606 VDDA.n2171 VDDA.n2170 3.4105
R1607 VDDA.n2169 VDDA.n2168 3.4105
R1608 VDDA.n2167 VDDA.n1928 3.4105
R1609 VDDA.n2163 VDDA.n2162 3.4105
R1610 VDDA.n2161 VDDA.n2160 3.4105
R1611 VDDA.n2159 VDDA.n2158 3.4105
R1612 VDDA.n2157 VDDA.n1930 3.4105
R1613 VDDA.n2153 VDDA.n2152 3.4105
R1614 VDDA.n2151 VDDA.n2150 3.4105
R1615 VDDA.n2149 VDDA.n2148 3.4105
R1616 VDDA.n2147 VDDA.n1932 3.4105
R1617 VDDA.n45 VDDA.n44 3.4105
R1618 VDDA.n179 VDDA.n178 3.4105
R1619 VDDA.n177 VDDA.n176 3.4105
R1620 VDDA.n175 VDDA.n49 3.4105
R1621 VDDA.n48 VDDA.n47 3.4105
R1622 VDDA.n171 VDDA.n170 3.4105
R1623 VDDA.n169 VDDA.n168 3.4105
R1624 VDDA.n167 VDDA.n53 3.4105
R1625 VDDA.n52 VDDA.n51 3.4105
R1626 VDDA.n163 VDDA.n162 3.4105
R1627 VDDA.n161 VDDA.n160 3.4105
R1628 VDDA.n159 VDDA.n57 3.4105
R1629 VDDA.n56 VDDA.n55 3.4105
R1630 VDDA.n155 VDDA.n154 3.4105
R1631 VDDA.n153 VDDA.n152 3.4105
R1632 VDDA.n151 VDDA.n61 3.4105
R1633 VDDA.n60 VDDA.n59 3.4105
R1634 VDDA.n147 VDDA.n146 3.4105
R1635 VDDA.n145 VDDA.n144 3.4105
R1636 VDDA.n143 VDDA.n65 3.4105
R1637 VDDA.n64 VDDA.n63 3.4105
R1638 VDDA.n139 VDDA.n138 3.4105
R1639 VDDA.n137 VDDA.n136 3.4105
R1640 VDDA.n135 VDDA.n69 3.4105
R1641 VDDA.n68 VDDA.n67 3.4105
R1642 VDDA.n131 VDDA.n130 3.4105
R1643 VDDA.n129 VDDA.n128 3.4105
R1644 VDDA.n127 VDDA.n73 3.4105
R1645 VDDA.n72 VDDA.n71 3.4105
R1646 VDDA.n123 VDDA.n122 3.4105
R1647 VDDA.n121 VDDA.n120 3.4105
R1648 VDDA.n119 VDDA.n77 3.4105
R1649 VDDA.n76 VDDA.n75 3.4105
R1650 VDDA.n115 VDDA.n114 3.4105
R1651 VDDA.n113 VDDA.n112 3.4105
R1652 VDDA.n111 VDDA.n81 3.4105
R1653 VDDA.n80 VDDA.n79 3.4105
R1654 VDDA.n107 VDDA.n106 3.4105
R1655 VDDA.n105 VDDA.n104 3.4105
R1656 VDDA.n103 VDDA.n85 3.4105
R1657 VDDA.n84 VDDA.n83 3.4105
R1658 VDDA.n99 VDDA.n98 3.4105
R1659 VDDA.n97 VDDA.n96 3.4105
R1660 VDDA.n95 VDDA.n89 3.4105
R1661 VDDA.n88 VDDA.n87 3.4105
R1662 VDDA.n91 VDDA.n90 3.4105
R1663 VDDA.n2946 VDDA.n2945 3.4105
R1664 VDDA.n2930 VDDA.n2770 3.4105
R1665 VDDA.n2928 VDDA.n2927 3.4105
R1666 VDDA.n2772 VDDA.n2771 3.4105
R1667 VDDA.n2923 VDDA.n2922 3.4105
R1668 VDDA.n2920 VDDA.n2774 3.4105
R1669 VDDA.n2918 VDDA.n2917 3.4105
R1670 VDDA.n2776 VDDA.n2775 3.4105
R1671 VDDA.n2913 VDDA.n2912 3.4105
R1672 VDDA.n2910 VDDA.n2778 3.4105
R1673 VDDA.n2908 VDDA.n2907 3.4105
R1674 VDDA.n2780 VDDA.n2779 3.4105
R1675 VDDA.n2903 VDDA.n2902 3.4105
R1676 VDDA.n2900 VDDA.n2782 3.4105
R1677 VDDA.n2898 VDDA.n2897 3.4105
R1678 VDDA.n2784 VDDA.n2783 3.4105
R1679 VDDA.n2893 VDDA.n2892 3.4105
R1680 VDDA.n2890 VDDA.n2786 3.4105
R1681 VDDA.n2888 VDDA.n2887 3.4105
R1682 VDDA.n2788 VDDA.n2787 3.4105
R1683 VDDA.n2883 VDDA.n2882 3.4105
R1684 VDDA.n2880 VDDA.n2790 3.4105
R1685 VDDA.n2878 VDDA.n2877 3.4105
R1686 VDDA.n2792 VDDA.n2791 3.4105
R1687 VDDA.n2873 VDDA.n2872 3.4105
R1688 VDDA.n2870 VDDA.n2794 3.4105
R1689 VDDA.n2868 VDDA.n2867 3.4105
R1690 VDDA.n2796 VDDA.n2795 3.4105
R1691 VDDA.n2863 VDDA.n2862 3.4105
R1692 VDDA.n2860 VDDA.n2798 3.4105
R1693 VDDA.n2858 VDDA.n2857 3.4105
R1694 VDDA.n2800 VDDA.n2799 3.4105
R1695 VDDA.n2853 VDDA.n2852 3.4105
R1696 VDDA.n2850 VDDA.n2802 3.4105
R1697 VDDA.n2848 VDDA.n2847 3.4105
R1698 VDDA.n2804 VDDA.n2803 3.4105
R1699 VDDA.n2843 VDDA.n2842 3.4105
R1700 VDDA.n2840 VDDA.n2806 3.4105
R1701 VDDA.n2838 VDDA.n2837 3.4105
R1702 VDDA.n2808 VDDA.n2807 3.4105
R1703 VDDA.n2833 VDDA.n2832 3.4105
R1704 VDDA.n2830 VDDA.n2810 3.4105
R1705 VDDA.n2828 VDDA.n2827 3.4105
R1706 VDDA.n2812 VDDA.n2811 3.4105
R1707 VDDA.n2823 VDDA.n2822 3.4105
R1708 VDDA.n2820 VDDA.n2814 3.4105
R1709 VDDA.n2818 VDDA.n2817 3.4105
R1710 VDDA.n2932 VDDA.n2931 3.4105
R1711 VDDA.n196 VDDA.n195 3.4105
R1712 VDDA.n2757 VDDA.n2756 3.4105
R1713 VDDA.n2624 VDDA.n2623 3.4105
R1714 VDDA.n2752 VDDA.n2751 3.4105
R1715 VDDA.n2750 VDDA.n2749 3.4105
R1716 VDDA.n2748 VDDA.n2628 3.4105
R1717 VDDA.n2627 VDDA.n2626 3.4105
R1718 VDDA.n2744 VDDA.n2743 3.4105
R1719 VDDA.n2742 VDDA.n2741 3.4105
R1720 VDDA.n2740 VDDA.n2632 3.4105
R1721 VDDA.n2631 VDDA.n2630 3.4105
R1722 VDDA.n2736 VDDA.n2735 3.4105
R1723 VDDA.n2734 VDDA.n2733 3.4105
R1724 VDDA.n2732 VDDA.n2636 3.4105
R1725 VDDA.n2635 VDDA.n2634 3.4105
R1726 VDDA.n2728 VDDA.n2727 3.4105
R1727 VDDA.n2726 VDDA.n2725 3.4105
R1728 VDDA.n2724 VDDA.n2640 3.4105
R1729 VDDA.n2639 VDDA.n2638 3.4105
R1730 VDDA.n2720 VDDA.n2719 3.4105
R1731 VDDA.n2718 VDDA.n2717 3.4105
R1732 VDDA.n2716 VDDA.n2644 3.4105
R1733 VDDA.n2643 VDDA.n2642 3.4105
R1734 VDDA.n2712 VDDA.n2711 3.4105
R1735 VDDA.n2710 VDDA.n2709 3.4105
R1736 VDDA.n2708 VDDA.n2648 3.4105
R1737 VDDA.n2647 VDDA.n2646 3.4105
R1738 VDDA.n2704 VDDA.n2703 3.4105
R1739 VDDA.n2702 VDDA.n2701 3.4105
R1740 VDDA.n2700 VDDA.n2652 3.4105
R1741 VDDA.n2651 VDDA.n2650 3.4105
R1742 VDDA.n2696 VDDA.n2695 3.4105
R1743 VDDA.n2694 VDDA.n2693 3.4105
R1744 VDDA.n2692 VDDA.n2656 3.4105
R1745 VDDA.n2655 VDDA.n2654 3.4105
R1746 VDDA.n2688 VDDA.n2687 3.4105
R1747 VDDA.n2686 VDDA.n2685 3.4105
R1748 VDDA.n2684 VDDA.n2660 3.4105
R1749 VDDA.n2659 VDDA.n2658 3.4105
R1750 VDDA.n2680 VDDA.n2679 3.4105
R1751 VDDA.n2678 VDDA.n2677 3.4105
R1752 VDDA.n2676 VDDA.n2664 3.4105
R1753 VDDA.n2663 VDDA.n2662 3.4105
R1754 VDDA.n2672 VDDA.n2671 3.4105
R1755 VDDA.n2670 VDDA.n2669 3.4105
R1756 VDDA.n2668 VDDA.n2667 3.4105
R1757 VDDA.n2761 VDDA.n2760 3.4105
R1758 VDDA.n223 VDDA.n222 3.4105
R1759 VDDA.n357 VDDA.n356 3.4105
R1760 VDDA.n355 VDDA.n354 3.4105
R1761 VDDA.n353 VDDA.n227 3.4105
R1762 VDDA.n226 VDDA.n225 3.4105
R1763 VDDA.n349 VDDA.n348 3.4105
R1764 VDDA.n347 VDDA.n346 3.4105
R1765 VDDA.n345 VDDA.n231 3.4105
R1766 VDDA.n230 VDDA.n229 3.4105
R1767 VDDA.n341 VDDA.n340 3.4105
R1768 VDDA.n339 VDDA.n338 3.4105
R1769 VDDA.n337 VDDA.n235 3.4105
R1770 VDDA.n234 VDDA.n233 3.4105
R1771 VDDA.n333 VDDA.n332 3.4105
R1772 VDDA.n331 VDDA.n330 3.4105
R1773 VDDA.n329 VDDA.n239 3.4105
R1774 VDDA.n238 VDDA.n237 3.4105
R1775 VDDA.n325 VDDA.n324 3.4105
R1776 VDDA.n323 VDDA.n322 3.4105
R1777 VDDA.n321 VDDA.n243 3.4105
R1778 VDDA.n242 VDDA.n241 3.4105
R1779 VDDA.n317 VDDA.n316 3.4105
R1780 VDDA.n315 VDDA.n314 3.4105
R1781 VDDA.n313 VDDA.n247 3.4105
R1782 VDDA.n246 VDDA.n245 3.4105
R1783 VDDA.n309 VDDA.n308 3.4105
R1784 VDDA.n307 VDDA.n306 3.4105
R1785 VDDA.n305 VDDA.n251 3.4105
R1786 VDDA.n250 VDDA.n249 3.4105
R1787 VDDA.n301 VDDA.n300 3.4105
R1788 VDDA.n299 VDDA.n298 3.4105
R1789 VDDA.n297 VDDA.n255 3.4105
R1790 VDDA.n254 VDDA.n253 3.4105
R1791 VDDA.n293 VDDA.n292 3.4105
R1792 VDDA.n291 VDDA.n290 3.4105
R1793 VDDA.n289 VDDA.n259 3.4105
R1794 VDDA.n258 VDDA.n257 3.4105
R1795 VDDA.n285 VDDA.n284 3.4105
R1796 VDDA.n283 VDDA.n282 3.4105
R1797 VDDA.n281 VDDA.n263 3.4105
R1798 VDDA.n262 VDDA.n261 3.4105
R1799 VDDA.n277 VDDA.n276 3.4105
R1800 VDDA.n275 VDDA.n274 3.4105
R1801 VDDA.n273 VDDA.n267 3.4105
R1802 VDDA.n266 VDDA.n265 3.4105
R1803 VDDA.n269 VDDA.n268 3.4105
R1804 VDDA.n2598 VDDA.n2597 3.4105
R1805 VDDA.n2582 VDDA.n2422 3.4105
R1806 VDDA.n2580 VDDA.n2579 3.4105
R1807 VDDA.n2424 VDDA.n2423 3.4105
R1808 VDDA.n2575 VDDA.n2574 3.4105
R1809 VDDA.n2572 VDDA.n2426 3.4105
R1810 VDDA.n2570 VDDA.n2569 3.4105
R1811 VDDA.n2428 VDDA.n2427 3.4105
R1812 VDDA.n2565 VDDA.n2564 3.4105
R1813 VDDA.n2562 VDDA.n2430 3.4105
R1814 VDDA.n2560 VDDA.n2559 3.4105
R1815 VDDA.n2432 VDDA.n2431 3.4105
R1816 VDDA.n2555 VDDA.n2554 3.4105
R1817 VDDA.n2552 VDDA.n2434 3.4105
R1818 VDDA.n2550 VDDA.n2549 3.4105
R1819 VDDA.n2436 VDDA.n2435 3.4105
R1820 VDDA.n2545 VDDA.n2544 3.4105
R1821 VDDA.n2542 VDDA.n2438 3.4105
R1822 VDDA.n2540 VDDA.n2539 3.4105
R1823 VDDA.n2440 VDDA.n2439 3.4105
R1824 VDDA.n2535 VDDA.n2534 3.4105
R1825 VDDA.n2532 VDDA.n2442 3.4105
R1826 VDDA.n2530 VDDA.n2529 3.4105
R1827 VDDA.n2444 VDDA.n2443 3.4105
R1828 VDDA.n2525 VDDA.n2524 3.4105
R1829 VDDA.n2522 VDDA.n2446 3.4105
R1830 VDDA.n2520 VDDA.n2519 3.4105
R1831 VDDA.n2448 VDDA.n2447 3.4105
R1832 VDDA.n2515 VDDA.n2514 3.4105
R1833 VDDA.n2512 VDDA.n2450 3.4105
R1834 VDDA.n2510 VDDA.n2509 3.4105
R1835 VDDA.n2452 VDDA.n2451 3.4105
R1836 VDDA.n2505 VDDA.n2504 3.4105
R1837 VDDA.n2502 VDDA.n2454 3.4105
R1838 VDDA.n2500 VDDA.n2499 3.4105
R1839 VDDA.n2456 VDDA.n2455 3.4105
R1840 VDDA.n2495 VDDA.n2494 3.4105
R1841 VDDA.n2492 VDDA.n2458 3.4105
R1842 VDDA.n2490 VDDA.n2489 3.4105
R1843 VDDA.n2460 VDDA.n2459 3.4105
R1844 VDDA.n2485 VDDA.n2484 3.4105
R1845 VDDA.n2482 VDDA.n2462 3.4105
R1846 VDDA.n2480 VDDA.n2479 3.4105
R1847 VDDA.n2464 VDDA.n2463 3.4105
R1848 VDDA.n2475 VDDA.n2474 3.4105
R1849 VDDA.n2472 VDDA.n2466 3.4105
R1850 VDDA.n2470 VDDA.n2469 3.4105
R1851 VDDA.n2584 VDDA.n2583 3.4105
R1852 VDDA.n463 VDDA.n462 3.4105
R1853 VDDA.n1319 VDDA.n1318 3.4105
R1854 VDDA.n1186 VDDA.n1185 3.4105
R1855 VDDA.n1314 VDDA.n1313 3.4105
R1856 VDDA.n1312 VDDA.n1311 3.4105
R1857 VDDA.n1310 VDDA.n1190 3.4105
R1858 VDDA.n1189 VDDA.n1188 3.4105
R1859 VDDA.n1306 VDDA.n1305 3.4105
R1860 VDDA.n1304 VDDA.n1303 3.4105
R1861 VDDA.n1302 VDDA.n1194 3.4105
R1862 VDDA.n1193 VDDA.n1192 3.4105
R1863 VDDA.n1298 VDDA.n1297 3.4105
R1864 VDDA.n1296 VDDA.n1295 3.4105
R1865 VDDA.n1294 VDDA.n1198 3.4105
R1866 VDDA.n1197 VDDA.n1196 3.4105
R1867 VDDA.n1290 VDDA.n1289 3.4105
R1868 VDDA.n1288 VDDA.n1287 3.4105
R1869 VDDA.n1286 VDDA.n1202 3.4105
R1870 VDDA.n1201 VDDA.n1200 3.4105
R1871 VDDA.n1282 VDDA.n1281 3.4105
R1872 VDDA.n1280 VDDA.n1279 3.4105
R1873 VDDA.n1278 VDDA.n1206 3.4105
R1874 VDDA.n1205 VDDA.n1204 3.4105
R1875 VDDA.n1274 VDDA.n1273 3.4105
R1876 VDDA.n1272 VDDA.n1271 3.4105
R1877 VDDA.n1270 VDDA.n1210 3.4105
R1878 VDDA.n1209 VDDA.n1208 3.4105
R1879 VDDA.n1266 VDDA.n1265 3.4105
R1880 VDDA.n1264 VDDA.n1263 3.4105
R1881 VDDA.n1262 VDDA.n1214 3.4105
R1882 VDDA.n1213 VDDA.n1212 3.4105
R1883 VDDA.n1258 VDDA.n1257 3.4105
R1884 VDDA.n1256 VDDA.n1255 3.4105
R1885 VDDA.n1254 VDDA.n1218 3.4105
R1886 VDDA.n1217 VDDA.n1216 3.4105
R1887 VDDA.n1250 VDDA.n1249 3.4105
R1888 VDDA.n1248 VDDA.n1247 3.4105
R1889 VDDA.n1246 VDDA.n1222 3.4105
R1890 VDDA.n1221 VDDA.n1220 3.4105
R1891 VDDA.n1242 VDDA.n1241 3.4105
R1892 VDDA.n1240 VDDA.n1239 3.4105
R1893 VDDA.n1238 VDDA.n1226 3.4105
R1894 VDDA.n1225 VDDA.n1224 3.4105
R1895 VDDA.n1234 VDDA.n1233 3.4105
R1896 VDDA.n1232 VDDA.n1231 3.4105
R1897 VDDA.n1230 VDDA.n1229 3.4105
R1898 VDDA.n2260 VDDA.n2259 3.4105
R1899 VDDA.n490 VDDA.n489 3.4105
R1900 VDDA.n624 VDDA.n623 3.4105
R1901 VDDA.n622 VDDA.n621 3.4105
R1902 VDDA.n620 VDDA.n494 3.4105
R1903 VDDA.n493 VDDA.n492 3.4105
R1904 VDDA.n616 VDDA.n615 3.4105
R1905 VDDA.n614 VDDA.n613 3.4105
R1906 VDDA.n612 VDDA.n498 3.4105
R1907 VDDA.n497 VDDA.n496 3.4105
R1908 VDDA.n608 VDDA.n607 3.4105
R1909 VDDA.n606 VDDA.n605 3.4105
R1910 VDDA.n604 VDDA.n502 3.4105
R1911 VDDA.n501 VDDA.n500 3.4105
R1912 VDDA.n600 VDDA.n599 3.4105
R1913 VDDA.n598 VDDA.n597 3.4105
R1914 VDDA.n596 VDDA.n506 3.4105
R1915 VDDA.n505 VDDA.n504 3.4105
R1916 VDDA.n592 VDDA.n591 3.4105
R1917 VDDA.n590 VDDA.n589 3.4105
R1918 VDDA.n588 VDDA.n510 3.4105
R1919 VDDA.n509 VDDA.n508 3.4105
R1920 VDDA.n584 VDDA.n583 3.4105
R1921 VDDA.n582 VDDA.n581 3.4105
R1922 VDDA.n580 VDDA.n514 3.4105
R1923 VDDA.n513 VDDA.n512 3.4105
R1924 VDDA.n576 VDDA.n575 3.4105
R1925 VDDA.n574 VDDA.n573 3.4105
R1926 VDDA.n572 VDDA.n518 3.4105
R1927 VDDA.n517 VDDA.n516 3.4105
R1928 VDDA.n568 VDDA.n567 3.4105
R1929 VDDA.n566 VDDA.n565 3.4105
R1930 VDDA.n564 VDDA.n522 3.4105
R1931 VDDA.n521 VDDA.n520 3.4105
R1932 VDDA.n560 VDDA.n559 3.4105
R1933 VDDA.n558 VDDA.n557 3.4105
R1934 VDDA.n556 VDDA.n526 3.4105
R1935 VDDA.n525 VDDA.n524 3.4105
R1936 VDDA.n552 VDDA.n551 3.4105
R1937 VDDA.n550 VDDA.n549 3.4105
R1938 VDDA.n548 VDDA.n530 3.4105
R1939 VDDA.n529 VDDA.n528 3.4105
R1940 VDDA.n544 VDDA.n543 3.4105
R1941 VDDA.n542 VDDA.n541 3.4105
R1942 VDDA.n540 VDDA.n534 3.4105
R1943 VDDA.n533 VDDA.n532 3.4105
R1944 VDDA.n536 VDDA.n535 3.4105
R1945 VDDA.n1160 VDDA.n1159 3.4105
R1946 VDDA.n1144 VDDA.n984 3.4105
R1947 VDDA.n1142 VDDA.n1141 3.4105
R1948 VDDA.n986 VDDA.n985 3.4105
R1949 VDDA.n1137 VDDA.n1136 3.4105
R1950 VDDA.n1134 VDDA.n988 3.4105
R1951 VDDA.n1132 VDDA.n1131 3.4105
R1952 VDDA.n990 VDDA.n989 3.4105
R1953 VDDA.n1127 VDDA.n1126 3.4105
R1954 VDDA.n1124 VDDA.n992 3.4105
R1955 VDDA.n1122 VDDA.n1121 3.4105
R1956 VDDA.n994 VDDA.n993 3.4105
R1957 VDDA.n1117 VDDA.n1116 3.4105
R1958 VDDA.n1114 VDDA.n996 3.4105
R1959 VDDA.n1112 VDDA.n1111 3.4105
R1960 VDDA.n998 VDDA.n997 3.4105
R1961 VDDA.n1107 VDDA.n1106 3.4105
R1962 VDDA.n1104 VDDA.n1000 3.4105
R1963 VDDA.n1102 VDDA.n1101 3.4105
R1964 VDDA.n1002 VDDA.n1001 3.4105
R1965 VDDA.n1097 VDDA.n1096 3.4105
R1966 VDDA.n1094 VDDA.n1004 3.4105
R1967 VDDA.n1092 VDDA.n1091 3.4105
R1968 VDDA.n1006 VDDA.n1005 3.4105
R1969 VDDA.n1087 VDDA.n1086 3.4105
R1970 VDDA.n1084 VDDA.n1008 3.4105
R1971 VDDA.n1082 VDDA.n1081 3.4105
R1972 VDDA.n1010 VDDA.n1009 3.4105
R1973 VDDA.n1077 VDDA.n1076 3.4105
R1974 VDDA.n1074 VDDA.n1012 3.4105
R1975 VDDA.n1072 VDDA.n1071 3.4105
R1976 VDDA.n1014 VDDA.n1013 3.4105
R1977 VDDA.n1067 VDDA.n1066 3.4105
R1978 VDDA.n1064 VDDA.n1016 3.4105
R1979 VDDA.n1062 VDDA.n1061 3.4105
R1980 VDDA.n1018 VDDA.n1017 3.4105
R1981 VDDA.n1057 VDDA.n1056 3.4105
R1982 VDDA.n1054 VDDA.n1020 3.4105
R1983 VDDA.n1052 VDDA.n1051 3.4105
R1984 VDDA.n1022 VDDA.n1021 3.4105
R1985 VDDA.n1047 VDDA.n1046 3.4105
R1986 VDDA.n1044 VDDA.n1024 3.4105
R1987 VDDA.n1042 VDDA.n1041 3.4105
R1988 VDDA.n1026 VDDA.n1025 3.4105
R1989 VDDA.n1037 VDDA.n1036 3.4105
R1990 VDDA.n1034 VDDA.n1028 3.4105
R1991 VDDA.n1032 VDDA.n1031 3.4105
R1992 VDDA.n1146 VDDA.n1145 3.4105
R1993 VDDA.n640 VDDA.n639 3.4105
R1994 VDDA.n971 VDDA.n970 3.4105
R1995 VDDA.n838 VDDA.n837 3.4105
R1996 VDDA.n966 VDDA.n965 3.4105
R1997 VDDA.n964 VDDA.n963 3.4105
R1998 VDDA.n962 VDDA.n842 3.4105
R1999 VDDA.n841 VDDA.n840 3.4105
R2000 VDDA.n958 VDDA.n957 3.4105
R2001 VDDA.n956 VDDA.n955 3.4105
R2002 VDDA.n954 VDDA.n846 3.4105
R2003 VDDA.n845 VDDA.n844 3.4105
R2004 VDDA.n950 VDDA.n949 3.4105
R2005 VDDA.n948 VDDA.n947 3.4105
R2006 VDDA.n946 VDDA.n850 3.4105
R2007 VDDA.n849 VDDA.n848 3.4105
R2008 VDDA.n942 VDDA.n941 3.4105
R2009 VDDA.n940 VDDA.n939 3.4105
R2010 VDDA.n938 VDDA.n854 3.4105
R2011 VDDA.n853 VDDA.n852 3.4105
R2012 VDDA.n934 VDDA.n933 3.4105
R2013 VDDA.n932 VDDA.n931 3.4105
R2014 VDDA.n930 VDDA.n858 3.4105
R2015 VDDA.n857 VDDA.n856 3.4105
R2016 VDDA.n926 VDDA.n925 3.4105
R2017 VDDA.n924 VDDA.n923 3.4105
R2018 VDDA.n922 VDDA.n862 3.4105
R2019 VDDA.n861 VDDA.n860 3.4105
R2020 VDDA.n918 VDDA.n917 3.4105
R2021 VDDA.n916 VDDA.n915 3.4105
R2022 VDDA.n914 VDDA.n866 3.4105
R2023 VDDA.n865 VDDA.n864 3.4105
R2024 VDDA.n910 VDDA.n909 3.4105
R2025 VDDA.n908 VDDA.n907 3.4105
R2026 VDDA.n906 VDDA.n870 3.4105
R2027 VDDA.n869 VDDA.n868 3.4105
R2028 VDDA.n902 VDDA.n901 3.4105
R2029 VDDA.n900 VDDA.n899 3.4105
R2030 VDDA.n898 VDDA.n874 3.4105
R2031 VDDA.n873 VDDA.n872 3.4105
R2032 VDDA.n894 VDDA.n893 3.4105
R2033 VDDA.n892 VDDA.n891 3.4105
R2034 VDDA.n890 VDDA.n878 3.4105
R2035 VDDA.n877 VDDA.n876 3.4105
R2036 VDDA.n886 VDDA.n885 3.4105
R2037 VDDA.n884 VDDA.n883 3.4105
R2038 VDDA.n882 VDDA.n881 3.4105
R2039 VDDA.n975 VDDA.n974 3.4105
R2040 VDDA.n666 VDDA.n665 3.4105
R2041 VDDA.n800 VDDA.n799 3.4105
R2042 VDDA.n798 VDDA.n797 3.4105
R2043 VDDA.n796 VDDA.n795 3.4105
R2044 VDDA.n794 VDDA.n668 3.4105
R2045 VDDA.n790 VDDA.n789 3.4105
R2046 VDDA.n788 VDDA.n787 3.4105
R2047 VDDA.n786 VDDA.n785 3.4105
R2048 VDDA.n784 VDDA.n670 3.4105
R2049 VDDA.n780 VDDA.n779 3.4105
R2050 VDDA.n778 VDDA.n777 3.4105
R2051 VDDA.n776 VDDA.n775 3.4105
R2052 VDDA.n774 VDDA.n672 3.4105
R2053 VDDA.n770 VDDA.n769 3.4105
R2054 VDDA.n768 VDDA.n767 3.4105
R2055 VDDA.n766 VDDA.n765 3.4105
R2056 VDDA.n764 VDDA.n674 3.4105
R2057 VDDA.n760 VDDA.n759 3.4105
R2058 VDDA.n758 VDDA.n757 3.4105
R2059 VDDA.n756 VDDA.n755 3.4105
R2060 VDDA.n754 VDDA.n676 3.4105
R2061 VDDA.n750 VDDA.n749 3.4105
R2062 VDDA.n748 VDDA.n747 3.4105
R2063 VDDA.n746 VDDA.n745 3.4105
R2064 VDDA.n744 VDDA.n678 3.4105
R2065 VDDA.n740 VDDA.n739 3.4105
R2066 VDDA.n738 VDDA.n737 3.4105
R2067 VDDA.n736 VDDA.n735 3.4105
R2068 VDDA.n734 VDDA.n680 3.4105
R2069 VDDA.n730 VDDA.n729 3.4105
R2070 VDDA.n728 VDDA.n727 3.4105
R2071 VDDA.n726 VDDA.n725 3.4105
R2072 VDDA.n724 VDDA.n682 3.4105
R2073 VDDA.n720 VDDA.n719 3.4105
R2074 VDDA.n718 VDDA.n717 3.4105
R2075 VDDA.n716 VDDA.n715 3.4105
R2076 VDDA.n714 VDDA.n684 3.4105
R2077 VDDA.n710 VDDA.n709 3.4105
R2078 VDDA.n708 VDDA.n707 3.4105
R2079 VDDA.n706 VDDA.n705 3.4105
R2080 VDDA.n704 VDDA.n686 3.4105
R2081 VDDA.n700 VDDA.n699 3.4105
R2082 VDDA.n698 VDDA.n697 3.4105
R2083 VDDA.n696 VDDA.n695 3.4105
R2084 VDDA.n694 VDDA.n688 3.4105
R2085 VDDA.n690 VDDA.n689 3.4105
R2086 VDDA.n812 VDDA.n811 3.4105
R2087 VDDA.n813 VDDA.n641 3.4105
R2088 VDDA.n813 VDDA.n812 3.4105
R2089 VDDA.n973 VDDA.n814 3.4105
R2090 VDDA.n974 VDDA.n973 3.4105
R2091 VDDA.n1029 VDDA.n464 3.4105
R2092 VDDA.n1145 VDDA.n464 3.4105
R2093 VDDA.n1161 VDDA.n465 3.4105
R2094 VDDA.n1161 VDDA.n1160 3.4105
R2095 VDDA.n2258 VDDA.n1162 3.4105
R2096 VDDA.n2259 VDDA.n2258 3.4105
R2097 VDDA.n2257 VDDA.n2256 3.4105
R2098 VDDA.n2467 VDDA.n197 3.4105
R2099 VDDA.n2583 VDDA.n197 3.4105
R2100 VDDA.n2599 VDDA.n198 3.4105
R2101 VDDA.n2599 VDDA.n2598 3.4105
R2102 VDDA.n2759 VDDA.n2600 3.4105
R2103 VDDA.n2760 VDDA.n2759 3.4105
R2104 VDDA.n2815 VDDA.n19 3.4105
R2105 VDDA.n2931 VDDA.n19 3.4105
R2106 VDDA.n2947 VDDA.n20 3.4105
R2107 VDDA.n2947 VDDA.n2946 3.4105
R2108 VDDA.n1580 VDDA.n1410 3.4105
R2109 VDDA.n1580 VDDA.n1579 3.4105
R2110 VDDA.n1908 VDDA.n1344 3.4105
R2111 VDDA.n1908 VDDA.n1907 3.4105
R2112 VDDA.n1581 VDDA.n1409 3.4105
R2113 VDDA.n1646 VDDA.n1581 3.4105
R2114 VDDA.n3134 VDDA.n17 3.4105
R2115 VDDA.n3134 VDDA.n16 3.4105
R2116 VDDA.n3134 VDDA.n18 3.4105
R2117 VDDA.n3134 VDDA.n3133 3.4105
R2118 VDDA.n3133 VDDA.n2984 3.4105
R2119 VDDA.n2981 VDDA.n16 3.4105
R2120 VDDA.n3103 VDDA.n2981 3.4105
R2121 VDDA.n3100 VDDA.n2981 3.4105
R2122 VDDA.n3105 VDDA.n2981 3.4105
R2123 VDDA.n3099 VDDA.n2981 3.4105
R2124 VDDA.n3107 VDDA.n2981 3.4105
R2125 VDDA.n3098 VDDA.n2981 3.4105
R2126 VDDA.n3109 VDDA.n2981 3.4105
R2127 VDDA.n3097 VDDA.n2981 3.4105
R2128 VDDA.n3111 VDDA.n2981 3.4105
R2129 VDDA.n3096 VDDA.n2981 3.4105
R2130 VDDA.n3113 VDDA.n2981 3.4105
R2131 VDDA.n3095 VDDA.n2981 3.4105
R2132 VDDA.n3115 VDDA.n2981 3.4105
R2133 VDDA.n3094 VDDA.n2981 3.4105
R2134 VDDA.n3117 VDDA.n2981 3.4105
R2135 VDDA.n3093 VDDA.n2981 3.4105
R2136 VDDA.n3119 VDDA.n2981 3.4105
R2137 VDDA.n3092 VDDA.n2981 3.4105
R2138 VDDA.n3121 VDDA.n2981 3.4105
R2139 VDDA.n3091 VDDA.n2981 3.4105
R2140 VDDA.n3123 VDDA.n2981 3.4105
R2141 VDDA.n3090 VDDA.n2981 3.4105
R2142 VDDA.n3125 VDDA.n2981 3.4105
R2143 VDDA.n3089 VDDA.n2981 3.4105
R2144 VDDA.n3127 VDDA.n2981 3.4105
R2145 VDDA.n3088 VDDA.n2981 3.4105
R2146 VDDA.n3129 VDDA.n2981 3.4105
R2147 VDDA.n3087 VDDA.n2981 3.4105
R2148 VDDA.n3131 VDDA.n2981 3.4105
R2149 VDDA.n3086 VDDA.n2981 3.4105
R2150 VDDA.n2981 VDDA.n18 3.4105
R2151 VDDA.n3133 VDDA.n2981 3.4105
R2152 VDDA.n2987 VDDA.n16 3.4105
R2153 VDDA.n3103 VDDA.n2987 3.4105
R2154 VDDA.n3100 VDDA.n2987 3.4105
R2155 VDDA.n3105 VDDA.n2987 3.4105
R2156 VDDA.n3099 VDDA.n2987 3.4105
R2157 VDDA.n3107 VDDA.n2987 3.4105
R2158 VDDA.n3098 VDDA.n2987 3.4105
R2159 VDDA.n3109 VDDA.n2987 3.4105
R2160 VDDA.n3097 VDDA.n2987 3.4105
R2161 VDDA.n3111 VDDA.n2987 3.4105
R2162 VDDA.n3096 VDDA.n2987 3.4105
R2163 VDDA.n3113 VDDA.n2987 3.4105
R2164 VDDA.n3095 VDDA.n2987 3.4105
R2165 VDDA.n3115 VDDA.n2987 3.4105
R2166 VDDA.n3094 VDDA.n2987 3.4105
R2167 VDDA.n3117 VDDA.n2987 3.4105
R2168 VDDA.n3093 VDDA.n2987 3.4105
R2169 VDDA.n3119 VDDA.n2987 3.4105
R2170 VDDA.n3092 VDDA.n2987 3.4105
R2171 VDDA.n3121 VDDA.n2987 3.4105
R2172 VDDA.n3091 VDDA.n2987 3.4105
R2173 VDDA.n3123 VDDA.n2987 3.4105
R2174 VDDA.n3090 VDDA.n2987 3.4105
R2175 VDDA.n3125 VDDA.n2987 3.4105
R2176 VDDA.n3089 VDDA.n2987 3.4105
R2177 VDDA.n3127 VDDA.n2987 3.4105
R2178 VDDA.n3088 VDDA.n2987 3.4105
R2179 VDDA.n3129 VDDA.n2987 3.4105
R2180 VDDA.n3087 VDDA.n2987 3.4105
R2181 VDDA.n3131 VDDA.n2987 3.4105
R2182 VDDA.n3086 VDDA.n2987 3.4105
R2183 VDDA.n2987 VDDA.n18 3.4105
R2184 VDDA.n3133 VDDA.n2987 3.4105
R2185 VDDA.n2980 VDDA.n16 3.4105
R2186 VDDA.n3103 VDDA.n2980 3.4105
R2187 VDDA.n3100 VDDA.n2980 3.4105
R2188 VDDA.n3105 VDDA.n2980 3.4105
R2189 VDDA.n3099 VDDA.n2980 3.4105
R2190 VDDA.n3107 VDDA.n2980 3.4105
R2191 VDDA.n3098 VDDA.n2980 3.4105
R2192 VDDA.n3109 VDDA.n2980 3.4105
R2193 VDDA.n3097 VDDA.n2980 3.4105
R2194 VDDA.n3111 VDDA.n2980 3.4105
R2195 VDDA.n3096 VDDA.n2980 3.4105
R2196 VDDA.n3113 VDDA.n2980 3.4105
R2197 VDDA.n3095 VDDA.n2980 3.4105
R2198 VDDA.n3115 VDDA.n2980 3.4105
R2199 VDDA.n3094 VDDA.n2980 3.4105
R2200 VDDA.n3117 VDDA.n2980 3.4105
R2201 VDDA.n3093 VDDA.n2980 3.4105
R2202 VDDA.n3119 VDDA.n2980 3.4105
R2203 VDDA.n3092 VDDA.n2980 3.4105
R2204 VDDA.n3121 VDDA.n2980 3.4105
R2205 VDDA.n3091 VDDA.n2980 3.4105
R2206 VDDA.n3123 VDDA.n2980 3.4105
R2207 VDDA.n3090 VDDA.n2980 3.4105
R2208 VDDA.n3125 VDDA.n2980 3.4105
R2209 VDDA.n3089 VDDA.n2980 3.4105
R2210 VDDA.n3127 VDDA.n2980 3.4105
R2211 VDDA.n3088 VDDA.n2980 3.4105
R2212 VDDA.n3129 VDDA.n2980 3.4105
R2213 VDDA.n3087 VDDA.n2980 3.4105
R2214 VDDA.n3131 VDDA.n2980 3.4105
R2215 VDDA.n3086 VDDA.n2980 3.4105
R2216 VDDA.n2980 VDDA.n18 3.4105
R2217 VDDA.n3133 VDDA.n2980 3.4105
R2218 VDDA.n2990 VDDA.n16 3.4105
R2219 VDDA.n3103 VDDA.n2990 3.4105
R2220 VDDA.n3100 VDDA.n2990 3.4105
R2221 VDDA.n3105 VDDA.n2990 3.4105
R2222 VDDA.n3099 VDDA.n2990 3.4105
R2223 VDDA.n3107 VDDA.n2990 3.4105
R2224 VDDA.n3098 VDDA.n2990 3.4105
R2225 VDDA.n3109 VDDA.n2990 3.4105
R2226 VDDA.n3097 VDDA.n2990 3.4105
R2227 VDDA.n3111 VDDA.n2990 3.4105
R2228 VDDA.n3096 VDDA.n2990 3.4105
R2229 VDDA.n3113 VDDA.n2990 3.4105
R2230 VDDA.n3095 VDDA.n2990 3.4105
R2231 VDDA.n3115 VDDA.n2990 3.4105
R2232 VDDA.n3094 VDDA.n2990 3.4105
R2233 VDDA.n3117 VDDA.n2990 3.4105
R2234 VDDA.n3093 VDDA.n2990 3.4105
R2235 VDDA.n3119 VDDA.n2990 3.4105
R2236 VDDA.n3092 VDDA.n2990 3.4105
R2237 VDDA.n3121 VDDA.n2990 3.4105
R2238 VDDA.n3091 VDDA.n2990 3.4105
R2239 VDDA.n3123 VDDA.n2990 3.4105
R2240 VDDA.n3090 VDDA.n2990 3.4105
R2241 VDDA.n3125 VDDA.n2990 3.4105
R2242 VDDA.n3089 VDDA.n2990 3.4105
R2243 VDDA.n3127 VDDA.n2990 3.4105
R2244 VDDA.n3088 VDDA.n2990 3.4105
R2245 VDDA.n3129 VDDA.n2990 3.4105
R2246 VDDA.n3087 VDDA.n2990 3.4105
R2247 VDDA.n3131 VDDA.n2990 3.4105
R2248 VDDA.n3086 VDDA.n2990 3.4105
R2249 VDDA.n2990 VDDA.n18 3.4105
R2250 VDDA.n3133 VDDA.n2990 3.4105
R2251 VDDA.n2979 VDDA.n16 3.4105
R2252 VDDA.n3103 VDDA.n2979 3.4105
R2253 VDDA.n3100 VDDA.n2979 3.4105
R2254 VDDA.n3105 VDDA.n2979 3.4105
R2255 VDDA.n3099 VDDA.n2979 3.4105
R2256 VDDA.n3107 VDDA.n2979 3.4105
R2257 VDDA.n3098 VDDA.n2979 3.4105
R2258 VDDA.n3109 VDDA.n2979 3.4105
R2259 VDDA.n3097 VDDA.n2979 3.4105
R2260 VDDA.n3111 VDDA.n2979 3.4105
R2261 VDDA.n3096 VDDA.n2979 3.4105
R2262 VDDA.n3113 VDDA.n2979 3.4105
R2263 VDDA.n3095 VDDA.n2979 3.4105
R2264 VDDA.n3115 VDDA.n2979 3.4105
R2265 VDDA.n3094 VDDA.n2979 3.4105
R2266 VDDA.n3117 VDDA.n2979 3.4105
R2267 VDDA.n3093 VDDA.n2979 3.4105
R2268 VDDA.n3119 VDDA.n2979 3.4105
R2269 VDDA.n3092 VDDA.n2979 3.4105
R2270 VDDA.n3121 VDDA.n2979 3.4105
R2271 VDDA.n3091 VDDA.n2979 3.4105
R2272 VDDA.n3123 VDDA.n2979 3.4105
R2273 VDDA.n3090 VDDA.n2979 3.4105
R2274 VDDA.n3125 VDDA.n2979 3.4105
R2275 VDDA.n3089 VDDA.n2979 3.4105
R2276 VDDA.n3127 VDDA.n2979 3.4105
R2277 VDDA.n3088 VDDA.n2979 3.4105
R2278 VDDA.n3129 VDDA.n2979 3.4105
R2279 VDDA.n3087 VDDA.n2979 3.4105
R2280 VDDA.n3131 VDDA.n2979 3.4105
R2281 VDDA.n3086 VDDA.n2979 3.4105
R2282 VDDA.n2979 VDDA.n18 3.4105
R2283 VDDA.n3133 VDDA.n2979 3.4105
R2284 VDDA.n2993 VDDA.n16 3.4105
R2285 VDDA.n3103 VDDA.n2993 3.4105
R2286 VDDA.n3100 VDDA.n2993 3.4105
R2287 VDDA.n3105 VDDA.n2993 3.4105
R2288 VDDA.n3099 VDDA.n2993 3.4105
R2289 VDDA.n3107 VDDA.n2993 3.4105
R2290 VDDA.n3098 VDDA.n2993 3.4105
R2291 VDDA.n3109 VDDA.n2993 3.4105
R2292 VDDA.n3097 VDDA.n2993 3.4105
R2293 VDDA.n3111 VDDA.n2993 3.4105
R2294 VDDA.n3096 VDDA.n2993 3.4105
R2295 VDDA.n3113 VDDA.n2993 3.4105
R2296 VDDA.n3095 VDDA.n2993 3.4105
R2297 VDDA.n3115 VDDA.n2993 3.4105
R2298 VDDA.n3094 VDDA.n2993 3.4105
R2299 VDDA.n3117 VDDA.n2993 3.4105
R2300 VDDA.n3093 VDDA.n2993 3.4105
R2301 VDDA.n3119 VDDA.n2993 3.4105
R2302 VDDA.n3092 VDDA.n2993 3.4105
R2303 VDDA.n3121 VDDA.n2993 3.4105
R2304 VDDA.n3091 VDDA.n2993 3.4105
R2305 VDDA.n3123 VDDA.n2993 3.4105
R2306 VDDA.n3090 VDDA.n2993 3.4105
R2307 VDDA.n3125 VDDA.n2993 3.4105
R2308 VDDA.n3089 VDDA.n2993 3.4105
R2309 VDDA.n3127 VDDA.n2993 3.4105
R2310 VDDA.n3088 VDDA.n2993 3.4105
R2311 VDDA.n3129 VDDA.n2993 3.4105
R2312 VDDA.n3087 VDDA.n2993 3.4105
R2313 VDDA.n3131 VDDA.n2993 3.4105
R2314 VDDA.n3086 VDDA.n2993 3.4105
R2315 VDDA.n2993 VDDA.n18 3.4105
R2316 VDDA.n3133 VDDA.n2993 3.4105
R2317 VDDA.n2978 VDDA.n16 3.4105
R2318 VDDA.n3103 VDDA.n2978 3.4105
R2319 VDDA.n3100 VDDA.n2978 3.4105
R2320 VDDA.n3105 VDDA.n2978 3.4105
R2321 VDDA.n3099 VDDA.n2978 3.4105
R2322 VDDA.n3107 VDDA.n2978 3.4105
R2323 VDDA.n3098 VDDA.n2978 3.4105
R2324 VDDA.n3109 VDDA.n2978 3.4105
R2325 VDDA.n3097 VDDA.n2978 3.4105
R2326 VDDA.n3111 VDDA.n2978 3.4105
R2327 VDDA.n3096 VDDA.n2978 3.4105
R2328 VDDA.n3113 VDDA.n2978 3.4105
R2329 VDDA.n3095 VDDA.n2978 3.4105
R2330 VDDA.n3115 VDDA.n2978 3.4105
R2331 VDDA.n3094 VDDA.n2978 3.4105
R2332 VDDA.n3117 VDDA.n2978 3.4105
R2333 VDDA.n3093 VDDA.n2978 3.4105
R2334 VDDA.n3119 VDDA.n2978 3.4105
R2335 VDDA.n3092 VDDA.n2978 3.4105
R2336 VDDA.n3121 VDDA.n2978 3.4105
R2337 VDDA.n3091 VDDA.n2978 3.4105
R2338 VDDA.n3123 VDDA.n2978 3.4105
R2339 VDDA.n3090 VDDA.n2978 3.4105
R2340 VDDA.n3125 VDDA.n2978 3.4105
R2341 VDDA.n3089 VDDA.n2978 3.4105
R2342 VDDA.n3127 VDDA.n2978 3.4105
R2343 VDDA.n3088 VDDA.n2978 3.4105
R2344 VDDA.n3129 VDDA.n2978 3.4105
R2345 VDDA.n3087 VDDA.n2978 3.4105
R2346 VDDA.n3131 VDDA.n2978 3.4105
R2347 VDDA.n3086 VDDA.n2978 3.4105
R2348 VDDA.n2978 VDDA.n18 3.4105
R2349 VDDA.n3133 VDDA.n2978 3.4105
R2350 VDDA.n2996 VDDA.n16 3.4105
R2351 VDDA.n3103 VDDA.n2996 3.4105
R2352 VDDA.n3100 VDDA.n2996 3.4105
R2353 VDDA.n3105 VDDA.n2996 3.4105
R2354 VDDA.n3099 VDDA.n2996 3.4105
R2355 VDDA.n3107 VDDA.n2996 3.4105
R2356 VDDA.n3098 VDDA.n2996 3.4105
R2357 VDDA.n3109 VDDA.n2996 3.4105
R2358 VDDA.n3097 VDDA.n2996 3.4105
R2359 VDDA.n3111 VDDA.n2996 3.4105
R2360 VDDA.n3096 VDDA.n2996 3.4105
R2361 VDDA.n3113 VDDA.n2996 3.4105
R2362 VDDA.n3095 VDDA.n2996 3.4105
R2363 VDDA.n3115 VDDA.n2996 3.4105
R2364 VDDA.n3094 VDDA.n2996 3.4105
R2365 VDDA.n3117 VDDA.n2996 3.4105
R2366 VDDA.n3093 VDDA.n2996 3.4105
R2367 VDDA.n3119 VDDA.n2996 3.4105
R2368 VDDA.n3092 VDDA.n2996 3.4105
R2369 VDDA.n3121 VDDA.n2996 3.4105
R2370 VDDA.n3091 VDDA.n2996 3.4105
R2371 VDDA.n3123 VDDA.n2996 3.4105
R2372 VDDA.n3090 VDDA.n2996 3.4105
R2373 VDDA.n3125 VDDA.n2996 3.4105
R2374 VDDA.n3089 VDDA.n2996 3.4105
R2375 VDDA.n3127 VDDA.n2996 3.4105
R2376 VDDA.n3088 VDDA.n2996 3.4105
R2377 VDDA.n3129 VDDA.n2996 3.4105
R2378 VDDA.n3087 VDDA.n2996 3.4105
R2379 VDDA.n3131 VDDA.n2996 3.4105
R2380 VDDA.n3086 VDDA.n2996 3.4105
R2381 VDDA.n2996 VDDA.n18 3.4105
R2382 VDDA.n3133 VDDA.n2996 3.4105
R2383 VDDA.n2977 VDDA.n16 3.4105
R2384 VDDA.n3103 VDDA.n2977 3.4105
R2385 VDDA.n3100 VDDA.n2977 3.4105
R2386 VDDA.n3105 VDDA.n2977 3.4105
R2387 VDDA.n3099 VDDA.n2977 3.4105
R2388 VDDA.n3107 VDDA.n2977 3.4105
R2389 VDDA.n3098 VDDA.n2977 3.4105
R2390 VDDA.n3109 VDDA.n2977 3.4105
R2391 VDDA.n3097 VDDA.n2977 3.4105
R2392 VDDA.n3111 VDDA.n2977 3.4105
R2393 VDDA.n3096 VDDA.n2977 3.4105
R2394 VDDA.n3113 VDDA.n2977 3.4105
R2395 VDDA.n3095 VDDA.n2977 3.4105
R2396 VDDA.n3115 VDDA.n2977 3.4105
R2397 VDDA.n3094 VDDA.n2977 3.4105
R2398 VDDA.n3117 VDDA.n2977 3.4105
R2399 VDDA.n3093 VDDA.n2977 3.4105
R2400 VDDA.n3119 VDDA.n2977 3.4105
R2401 VDDA.n3092 VDDA.n2977 3.4105
R2402 VDDA.n3121 VDDA.n2977 3.4105
R2403 VDDA.n3091 VDDA.n2977 3.4105
R2404 VDDA.n3123 VDDA.n2977 3.4105
R2405 VDDA.n3090 VDDA.n2977 3.4105
R2406 VDDA.n3125 VDDA.n2977 3.4105
R2407 VDDA.n3089 VDDA.n2977 3.4105
R2408 VDDA.n3127 VDDA.n2977 3.4105
R2409 VDDA.n3088 VDDA.n2977 3.4105
R2410 VDDA.n3129 VDDA.n2977 3.4105
R2411 VDDA.n3087 VDDA.n2977 3.4105
R2412 VDDA.n3131 VDDA.n2977 3.4105
R2413 VDDA.n3086 VDDA.n2977 3.4105
R2414 VDDA.n2977 VDDA.n18 3.4105
R2415 VDDA.n3133 VDDA.n2977 3.4105
R2416 VDDA.n2999 VDDA.n16 3.4105
R2417 VDDA.n3103 VDDA.n2999 3.4105
R2418 VDDA.n3100 VDDA.n2999 3.4105
R2419 VDDA.n3105 VDDA.n2999 3.4105
R2420 VDDA.n3099 VDDA.n2999 3.4105
R2421 VDDA.n3107 VDDA.n2999 3.4105
R2422 VDDA.n3098 VDDA.n2999 3.4105
R2423 VDDA.n3109 VDDA.n2999 3.4105
R2424 VDDA.n3097 VDDA.n2999 3.4105
R2425 VDDA.n3111 VDDA.n2999 3.4105
R2426 VDDA.n3096 VDDA.n2999 3.4105
R2427 VDDA.n3113 VDDA.n2999 3.4105
R2428 VDDA.n3095 VDDA.n2999 3.4105
R2429 VDDA.n3115 VDDA.n2999 3.4105
R2430 VDDA.n3094 VDDA.n2999 3.4105
R2431 VDDA.n3117 VDDA.n2999 3.4105
R2432 VDDA.n3093 VDDA.n2999 3.4105
R2433 VDDA.n3119 VDDA.n2999 3.4105
R2434 VDDA.n3092 VDDA.n2999 3.4105
R2435 VDDA.n3121 VDDA.n2999 3.4105
R2436 VDDA.n3091 VDDA.n2999 3.4105
R2437 VDDA.n3123 VDDA.n2999 3.4105
R2438 VDDA.n3090 VDDA.n2999 3.4105
R2439 VDDA.n3125 VDDA.n2999 3.4105
R2440 VDDA.n3089 VDDA.n2999 3.4105
R2441 VDDA.n3127 VDDA.n2999 3.4105
R2442 VDDA.n3088 VDDA.n2999 3.4105
R2443 VDDA.n3129 VDDA.n2999 3.4105
R2444 VDDA.n3087 VDDA.n2999 3.4105
R2445 VDDA.n3131 VDDA.n2999 3.4105
R2446 VDDA.n3086 VDDA.n2999 3.4105
R2447 VDDA.n2999 VDDA.n18 3.4105
R2448 VDDA.n3133 VDDA.n2999 3.4105
R2449 VDDA.n2976 VDDA.n16 3.4105
R2450 VDDA.n3103 VDDA.n2976 3.4105
R2451 VDDA.n3100 VDDA.n2976 3.4105
R2452 VDDA.n3105 VDDA.n2976 3.4105
R2453 VDDA.n3099 VDDA.n2976 3.4105
R2454 VDDA.n3107 VDDA.n2976 3.4105
R2455 VDDA.n3098 VDDA.n2976 3.4105
R2456 VDDA.n3109 VDDA.n2976 3.4105
R2457 VDDA.n3097 VDDA.n2976 3.4105
R2458 VDDA.n3111 VDDA.n2976 3.4105
R2459 VDDA.n3096 VDDA.n2976 3.4105
R2460 VDDA.n3113 VDDA.n2976 3.4105
R2461 VDDA.n3095 VDDA.n2976 3.4105
R2462 VDDA.n3115 VDDA.n2976 3.4105
R2463 VDDA.n3094 VDDA.n2976 3.4105
R2464 VDDA.n3117 VDDA.n2976 3.4105
R2465 VDDA.n3093 VDDA.n2976 3.4105
R2466 VDDA.n3119 VDDA.n2976 3.4105
R2467 VDDA.n3092 VDDA.n2976 3.4105
R2468 VDDA.n3121 VDDA.n2976 3.4105
R2469 VDDA.n3091 VDDA.n2976 3.4105
R2470 VDDA.n3123 VDDA.n2976 3.4105
R2471 VDDA.n3090 VDDA.n2976 3.4105
R2472 VDDA.n3125 VDDA.n2976 3.4105
R2473 VDDA.n3089 VDDA.n2976 3.4105
R2474 VDDA.n3127 VDDA.n2976 3.4105
R2475 VDDA.n3088 VDDA.n2976 3.4105
R2476 VDDA.n3129 VDDA.n2976 3.4105
R2477 VDDA.n3087 VDDA.n2976 3.4105
R2478 VDDA.n3131 VDDA.n2976 3.4105
R2479 VDDA.n3086 VDDA.n2976 3.4105
R2480 VDDA.n2976 VDDA.n18 3.4105
R2481 VDDA.n3133 VDDA.n2976 3.4105
R2482 VDDA.n3002 VDDA.n16 3.4105
R2483 VDDA.n3103 VDDA.n3002 3.4105
R2484 VDDA.n3100 VDDA.n3002 3.4105
R2485 VDDA.n3105 VDDA.n3002 3.4105
R2486 VDDA.n3099 VDDA.n3002 3.4105
R2487 VDDA.n3107 VDDA.n3002 3.4105
R2488 VDDA.n3098 VDDA.n3002 3.4105
R2489 VDDA.n3109 VDDA.n3002 3.4105
R2490 VDDA.n3097 VDDA.n3002 3.4105
R2491 VDDA.n3111 VDDA.n3002 3.4105
R2492 VDDA.n3096 VDDA.n3002 3.4105
R2493 VDDA.n3113 VDDA.n3002 3.4105
R2494 VDDA.n3095 VDDA.n3002 3.4105
R2495 VDDA.n3115 VDDA.n3002 3.4105
R2496 VDDA.n3094 VDDA.n3002 3.4105
R2497 VDDA.n3117 VDDA.n3002 3.4105
R2498 VDDA.n3093 VDDA.n3002 3.4105
R2499 VDDA.n3119 VDDA.n3002 3.4105
R2500 VDDA.n3092 VDDA.n3002 3.4105
R2501 VDDA.n3121 VDDA.n3002 3.4105
R2502 VDDA.n3091 VDDA.n3002 3.4105
R2503 VDDA.n3123 VDDA.n3002 3.4105
R2504 VDDA.n3090 VDDA.n3002 3.4105
R2505 VDDA.n3125 VDDA.n3002 3.4105
R2506 VDDA.n3089 VDDA.n3002 3.4105
R2507 VDDA.n3127 VDDA.n3002 3.4105
R2508 VDDA.n3088 VDDA.n3002 3.4105
R2509 VDDA.n3129 VDDA.n3002 3.4105
R2510 VDDA.n3087 VDDA.n3002 3.4105
R2511 VDDA.n3131 VDDA.n3002 3.4105
R2512 VDDA.n3086 VDDA.n3002 3.4105
R2513 VDDA.n3002 VDDA.n18 3.4105
R2514 VDDA.n3133 VDDA.n3002 3.4105
R2515 VDDA.n2975 VDDA.n16 3.4105
R2516 VDDA.n3103 VDDA.n2975 3.4105
R2517 VDDA.n3100 VDDA.n2975 3.4105
R2518 VDDA.n3105 VDDA.n2975 3.4105
R2519 VDDA.n3099 VDDA.n2975 3.4105
R2520 VDDA.n3107 VDDA.n2975 3.4105
R2521 VDDA.n3098 VDDA.n2975 3.4105
R2522 VDDA.n3109 VDDA.n2975 3.4105
R2523 VDDA.n3097 VDDA.n2975 3.4105
R2524 VDDA.n3111 VDDA.n2975 3.4105
R2525 VDDA.n3096 VDDA.n2975 3.4105
R2526 VDDA.n3113 VDDA.n2975 3.4105
R2527 VDDA.n3095 VDDA.n2975 3.4105
R2528 VDDA.n3115 VDDA.n2975 3.4105
R2529 VDDA.n3094 VDDA.n2975 3.4105
R2530 VDDA.n3117 VDDA.n2975 3.4105
R2531 VDDA.n3093 VDDA.n2975 3.4105
R2532 VDDA.n3119 VDDA.n2975 3.4105
R2533 VDDA.n3092 VDDA.n2975 3.4105
R2534 VDDA.n3121 VDDA.n2975 3.4105
R2535 VDDA.n3091 VDDA.n2975 3.4105
R2536 VDDA.n3123 VDDA.n2975 3.4105
R2537 VDDA.n3090 VDDA.n2975 3.4105
R2538 VDDA.n3125 VDDA.n2975 3.4105
R2539 VDDA.n3089 VDDA.n2975 3.4105
R2540 VDDA.n3127 VDDA.n2975 3.4105
R2541 VDDA.n3088 VDDA.n2975 3.4105
R2542 VDDA.n3129 VDDA.n2975 3.4105
R2543 VDDA.n3087 VDDA.n2975 3.4105
R2544 VDDA.n3131 VDDA.n2975 3.4105
R2545 VDDA.n3086 VDDA.n2975 3.4105
R2546 VDDA.n2975 VDDA.n18 3.4105
R2547 VDDA.n3133 VDDA.n2975 3.4105
R2548 VDDA.n3005 VDDA.n16 3.4105
R2549 VDDA.n3103 VDDA.n3005 3.4105
R2550 VDDA.n3100 VDDA.n3005 3.4105
R2551 VDDA.n3105 VDDA.n3005 3.4105
R2552 VDDA.n3099 VDDA.n3005 3.4105
R2553 VDDA.n3107 VDDA.n3005 3.4105
R2554 VDDA.n3098 VDDA.n3005 3.4105
R2555 VDDA.n3109 VDDA.n3005 3.4105
R2556 VDDA.n3097 VDDA.n3005 3.4105
R2557 VDDA.n3111 VDDA.n3005 3.4105
R2558 VDDA.n3096 VDDA.n3005 3.4105
R2559 VDDA.n3113 VDDA.n3005 3.4105
R2560 VDDA.n3095 VDDA.n3005 3.4105
R2561 VDDA.n3115 VDDA.n3005 3.4105
R2562 VDDA.n3094 VDDA.n3005 3.4105
R2563 VDDA.n3117 VDDA.n3005 3.4105
R2564 VDDA.n3093 VDDA.n3005 3.4105
R2565 VDDA.n3119 VDDA.n3005 3.4105
R2566 VDDA.n3092 VDDA.n3005 3.4105
R2567 VDDA.n3121 VDDA.n3005 3.4105
R2568 VDDA.n3091 VDDA.n3005 3.4105
R2569 VDDA.n3123 VDDA.n3005 3.4105
R2570 VDDA.n3090 VDDA.n3005 3.4105
R2571 VDDA.n3125 VDDA.n3005 3.4105
R2572 VDDA.n3089 VDDA.n3005 3.4105
R2573 VDDA.n3127 VDDA.n3005 3.4105
R2574 VDDA.n3088 VDDA.n3005 3.4105
R2575 VDDA.n3129 VDDA.n3005 3.4105
R2576 VDDA.n3087 VDDA.n3005 3.4105
R2577 VDDA.n3131 VDDA.n3005 3.4105
R2578 VDDA.n3086 VDDA.n3005 3.4105
R2579 VDDA.n3005 VDDA.n18 3.4105
R2580 VDDA.n3133 VDDA.n3005 3.4105
R2581 VDDA.n2974 VDDA.n16 3.4105
R2582 VDDA.n3103 VDDA.n2974 3.4105
R2583 VDDA.n3100 VDDA.n2974 3.4105
R2584 VDDA.n3105 VDDA.n2974 3.4105
R2585 VDDA.n3099 VDDA.n2974 3.4105
R2586 VDDA.n3107 VDDA.n2974 3.4105
R2587 VDDA.n3098 VDDA.n2974 3.4105
R2588 VDDA.n3109 VDDA.n2974 3.4105
R2589 VDDA.n3097 VDDA.n2974 3.4105
R2590 VDDA.n3111 VDDA.n2974 3.4105
R2591 VDDA.n3096 VDDA.n2974 3.4105
R2592 VDDA.n3113 VDDA.n2974 3.4105
R2593 VDDA.n3095 VDDA.n2974 3.4105
R2594 VDDA.n3115 VDDA.n2974 3.4105
R2595 VDDA.n3094 VDDA.n2974 3.4105
R2596 VDDA.n3117 VDDA.n2974 3.4105
R2597 VDDA.n3093 VDDA.n2974 3.4105
R2598 VDDA.n3119 VDDA.n2974 3.4105
R2599 VDDA.n3092 VDDA.n2974 3.4105
R2600 VDDA.n3121 VDDA.n2974 3.4105
R2601 VDDA.n3091 VDDA.n2974 3.4105
R2602 VDDA.n3123 VDDA.n2974 3.4105
R2603 VDDA.n3090 VDDA.n2974 3.4105
R2604 VDDA.n3125 VDDA.n2974 3.4105
R2605 VDDA.n3089 VDDA.n2974 3.4105
R2606 VDDA.n3127 VDDA.n2974 3.4105
R2607 VDDA.n3088 VDDA.n2974 3.4105
R2608 VDDA.n3129 VDDA.n2974 3.4105
R2609 VDDA.n3087 VDDA.n2974 3.4105
R2610 VDDA.n3131 VDDA.n2974 3.4105
R2611 VDDA.n3086 VDDA.n2974 3.4105
R2612 VDDA.n2974 VDDA.n18 3.4105
R2613 VDDA.n3133 VDDA.n2974 3.4105
R2614 VDDA.n3008 VDDA.n16 3.4105
R2615 VDDA.n3103 VDDA.n3008 3.4105
R2616 VDDA.n3100 VDDA.n3008 3.4105
R2617 VDDA.n3105 VDDA.n3008 3.4105
R2618 VDDA.n3099 VDDA.n3008 3.4105
R2619 VDDA.n3107 VDDA.n3008 3.4105
R2620 VDDA.n3098 VDDA.n3008 3.4105
R2621 VDDA.n3109 VDDA.n3008 3.4105
R2622 VDDA.n3097 VDDA.n3008 3.4105
R2623 VDDA.n3111 VDDA.n3008 3.4105
R2624 VDDA.n3096 VDDA.n3008 3.4105
R2625 VDDA.n3113 VDDA.n3008 3.4105
R2626 VDDA.n3095 VDDA.n3008 3.4105
R2627 VDDA.n3115 VDDA.n3008 3.4105
R2628 VDDA.n3094 VDDA.n3008 3.4105
R2629 VDDA.n3117 VDDA.n3008 3.4105
R2630 VDDA.n3093 VDDA.n3008 3.4105
R2631 VDDA.n3119 VDDA.n3008 3.4105
R2632 VDDA.n3092 VDDA.n3008 3.4105
R2633 VDDA.n3121 VDDA.n3008 3.4105
R2634 VDDA.n3091 VDDA.n3008 3.4105
R2635 VDDA.n3123 VDDA.n3008 3.4105
R2636 VDDA.n3090 VDDA.n3008 3.4105
R2637 VDDA.n3125 VDDA.n3008 3.4105
R2638 VDDA.n3089 VDDA.n3008 3.4105
R2639 VDDA.n3127 VDDA.n3008 3.4105
R2640 VDDA.n3088 VDDA.n3008 3.4105
R2641 VDDA.n3129 VDDA.n3008 3.4105
R2642 VDDA.n3087 VDDA.n3008 3.4105
R2643 VDDA.n3131 VDDA.n3008 3.4105
R2644 VDDA.n3086 VDDA.n3008 3.4105
R2645 VDDA.n3008 VDDA.n18 3.4105
R2646 VDDA.n3133 VDDA.n3008 3.4105
R2647 VDDA.n2973 VDDA.n16 3.4105
R2648 VDDA.n3103 VDDA.n2973 3.4105
R2649 VDDA.n3100 VDDA.n2973 3.4105
R2650 VDDA.n3105 VDDA.n2973 3.4105
R2651 VDDA.n3099 VDDA.n2973 3.4105
R2652 VDDA.n3107 VDDA.n2973 3.4105
R2653 VDDA.n3098 VDDA.n2973 3.4105
R2654 VDDA.n3109 VDDA.n2973 3.4105
R2655 VDDA.n3097 VDDA.n2973 3.4105
R2656 VDDA.n3111 VDDA.n2973 3.4105
R2657 VDDA.n3096 VDDA.n2973 3.4105
R2658 VDDA.n3113 VDDA.n2973 3.4105
R2659 VDDA.n3095 VDDA.n2973 3.4105
R2660 VDDA.n3115 VDDA.n2973 3.4105
R2661 VDDA.n3094 VDDA.n2973 3.4105
R2662 VDDA.n3117 VDDA.n2973 3.4105
R2663 VDDA.n3093 VDDA.n2973 3.4105
R2664 VDDA.n3119 VDDA.n2973 3.4105
R2665 VDDA.n3092 VDDA.n2973 3.4105
R2666 VDDA.n3121 VDDA.n2973 3.4105
R2667 VDDA.n3091 VDDA.n2973 3.4105
R2668 VDDA.n3123 VDDA.n2973 3.4105
R2669 VDDA.n3090 VDDA.n2973 3.4105
R2670 VDDA.n3125 VDDA.n2973 3.4105
R2671 VDDA.n3089 VDDA.n2973 3.4105
R2672 VDDA.n3127 VDDA.n2973 3.4105
R2673 VDDA.n3088 VDDA.n2973 3.4105
R2674 VDDA.n3129 VDDA.n2973 3.4105
R2675 VDDA.n3087 VDDA.n2973 3.4105
R2676 VDDA.n3131 VDDA.n2973 3.4105
R2677 VDDA.n3086 VDDA.n2973 3.4105
R2678 VDDA.n2973 VDDA.n18 3.4105
R2679 VDDA.n3133 VDDA.n2973 3.4105
R2680 VDDA.n3011 VDDA.n16 3.4105
R2681 VDDA.n3103 VDDA.n3011 3.4105
R2682 VDDA.n3100 VDDA.n3011 3.4105
R2683 VDDA.n3105 VDDA.n3011 3.4105
R2684 VDDA.n3099 VDDA.n3011 3.4105
R2685 VDDA.n3107 VDDA.n3011 3.4105
R2686 VDDA.n3098 VDDA.n3011 3.4105
R2687 VDDA.n3109 VDDA.n3011 3.4105
R2688 VDDA.n3097 VDDA.n3011 3.4105
R2689 VDDA.n3111 VDDA.n3011 3.4105
R2690 VDDA.n3096 VDDA.n3011 3.4105
R2691 VDDA.n3113 VDDA.n3011 3.4105
R2692 VDDA.n3095 VDDA.n3011 3.4105
R2693 VDDA.n3115 VDDA.n3011 3.4105
R2694 VDDA.n3094 VDDA.n3011 3.4105
R2695 VDDA.n3117 VDDA.n3011 3.4105
R2696 VDDA.n3093 VDDA.n3011 3.4105
R2697 VDDA.n3119 VDDA.n3011 3.4105
R2698 VDDA.n3092 VDDA.n3011 3.4105
R2699 VDDA.n3121 VDDA.n3011 3.4105
R2700 VDDA.n3091 VDDA.n3011 3.4105
R2701 VDDA.n3123 VDDA.n3011 3.4105
R2702 VDDA.n3090 VDDA.n3011 3.4105
R2703 VDDA.n3125 VDDA.n3011 3.4105
R2704 VDDA.n3089 VDDA.n3011 3.4105
R2705 VDDA.n3127 VDDA.n3011 3.4105
R2706 VDDA.n3088 VDDA.n3011 3.4105
R2707 VDDA.n3129 VDDA.n3011 3.4105
R2708 VDDA.n3087 VDDA.n3011 3.4105
R2709 VDDA.n3131 VDDA.n3011 3.4105
R2710 VDDA.n3086 VDDA.n3011 3.4105
R2711 VDDA.n3011 VDDA.n18 3.4105
R2712 VDDA.n3133 VDDA.n3011 3.4105
R2713 VDDA.n2972 VDDA.n16 3.4105
R2714 VDDA.n3103 VDDA.n2972 3.4105
R2715 VDDA.n3100 VDDA.n2972 3.4105
R2716 VDDA.n3105 VDDA.n2972 3.4105
R2717 VDDA.n3099 VDDA.n2972 3.4105
R2718 VDDA.n3107 VDDA.n2972 3.4105
R2719 VDDA.n3098 VDDA.n2972 3.4105
R2720 VDDA.n3109 VDDA.n2972 3.4105
R2721 VDDA.n3097 VDDA.n2972 3.4105
R2722 VDDA.n3111 VDDA.n2972 3.4105
R2723 VDDA.n3096 VDDA.n2972 3.4105
R2724 VDDA.n3113 VDDA.n2972 3.4105
R2725 VDDA.n3095 VDDA.n2972 3.4105
R2726 VDDA.n3115 VDDA.n2972 3.4105
R2727 VDDA.n3094 VDDA.n2972 3.4105
R2728 VDDA.n3117 VDDA.n2972 3.4105
R2729 VDDA.n3093 VDDA.n2972 3.4105
R2730 VDDA.n3119 VDDA.n2972 3.4105
R2731 VDDA.n3092 VDDA.n2972 3.4105
R2732 VDDA.n3121 VDDA.n2972 3.4105
R2733 VDDA.n3091 VDDA.n2972 3.4105
R2734 VDDA.n3123 VDDA.n2972 3.4105
R2735 VDDA.n3090 VDDA.n2972 3.4105
R2736 VDDA.n3125 VDDA.n2972 3.4105
R2737 VDDA.n3089 VDDA.n2972 3.4105
R2738 VDDA.n3127 VDDA.n2972 3.4105
R2739 VDDA.n3088 VDDA.n2972 3.4105
R2740 VDDA.n3129 VDDA.n2972 3.4105
R2741 VDDA.n3087 VDDA.n2972 3.4105
R2742 VDDA.n3131 VDDA.n2972 3.4105
R2743 VDDA.n3086 VDDA.n2972 3.4105
R2744 VDDA.n2972 VDDA.n18 3.4105
R2745 VDDA.n3133 VDDA.n2972 3.4105
R2746 VDDA.n3014 VDDA.n16 3.4105
R2747 VDDA.n3103 VDDA.n3014 3.4105
R2748 VDDA.n3100 VDDA.n3014 3.4105
R2749 VDDA.n3105 VDDA.n3014 3.4105
R2750 VDDA.n3099 VDDA.n3014 3.4105
R2751 VDDA.n3107 VDDA.n3014 3.4105
R2752 VDDA.n3098 VDDA.n3014 3.4105
R2753 VDDA.n3109 VDDA.n3014 3.4105
R2754 VDDA.n3097 VDDA.n3014 3.4105
R2755 VDDA.n3111 VDDA.n3014 3.4105
R2756 VDDA.n3096 VDDA.n3014 3.4105
R2757 VDDA.n3113 VDDA.n3014 3.4105
R2758 VDDA.n3095 VDDA.n3014 3.4105
R2759 VDDA.n3115 VDDA.n3014 3.4105
R2760 VDDA.n3094 VDDA.n3014 3.4105
R2761 VDDA.n3117 VDDA.n3014 3.4105
R2762 VDDA.n3093 VDDA.n3014 3.4105
R2763 VDDA.n3119 VDDA.n3014 3.4105
R2764 VDDA.n3092 VDDA.n3014 3.4105
R2765 VDDA.n3121 VDDA.n3014 3.4105
R2766 VDDA.n3091 VDDA.n3014 3.4105
R2767 VDDA.n3123 VDDA.n3014 3.4105
R2768 VDDA.n3090 VDDA.n3014 3.4105
R2769 VDDA.n3125 VDDA.n3014 3.4105
R2770 VDDA.n3089 VDDA.n3014 3.4105
R2771 VDDA.n3127 VDDA.n3014 3.4105
R2772 VDDA.n3088 VDDA.n3014 3.4105
R2773 VDDA.n3129 VDDA.n3014 3.4105
R2774 VDDA.n3087 VDDA.n3014 3.4105
R2775 VDDA.n3131 VDDA.n3014 3.4105
R2776 VDDA.n3086 VDDA.n3014 3.4105
R2777 VDDA.n3014 VDDA.n18 3.4105
R2778 VDDA.n3133 VDDA.n3014 3.4105
R2779 VDDA.n2971 VDDA.n16 3.4105
R2780 VDDA.n3103 VDDA.n2971 3.4105
R2781 VDDA.n3100 VDDA.n2971 3.4105
R2782 VDDA.n3105 VDDA.n2971 3.4105
R2783 VDDA.n3099 VDDA.n2971 3.4105
R2784 VDDA.n3107 VDDA.n2971 3.4105
R2785 VDDA.n3098 VDDA.n2971 3.4105
R2786 VDDA.n3109 VDDA.n2971 3.4105
R2787 VDDA.n3097 VDDA.n2971 3.4105
R2788 VDDA.n3111 VDDA.n2971 3.4105
R2789 VDDA.n3096 VDDA.n2971 3.4105
R2790 VDDA.n3113 VDDA.n2971 3.4105
R2791 VDDA.n3095 VDDA.n2971 3.4105
R2792 VDDA.n3115 VDDA.n2971 3.4105
R2793 VDDA.n3094 VDDA.n2971 3.4105
R2794 VDDA.n3117 VDDA.n2971 3.4105
R2795 VDDA.n3093 VDDA.n2971 3.4105
R2796 VDDA.n3119 VDDA.n2971 3.4105
R2797 VDDA.n3092 VDDA.n2971 3.4105
R2798 VDDA.n3121 VDDA.n2971 3.4105
R2799 VDDA.n3091 VDDA.n2971 3.4105
R2800 VDDA.n3123 VDDA.n2971 3.4105
R2801 VDDA.n3090 VDDA.n2971 3.4105
R2802 VDDA.n3125 VDDA.n2971 3.4105
R2803 VDDA.n3089 VDDA.n2971 3.4105
R2804 VDDA.n3127 VDDA.n2971 3.4105
R2805 VDDA.n3088 VDDA.n2971 3.4105
R2806 VDDA.n3129 VDDA.n2971 3.4105
R2807 VDDA.n3087 VDDA.n2971 3.4105
R2808 VDDA.n3131 VDDA.n2971 3.4105
R2809 VDDA.n3086 VDDA.n2971 3.4105
R2810 VDDA.n2971 VDDA.n18 3.4105
R2811 VDDA.n3133 VDDA.n2971 3.4105
R2812 VDDA.n3017 VDDA.n16 3.4105
R2813 VDDA.n3103 VDDA.n3017 3.4105
R2814 VDDA.n3100 VDDA.n3017 3.4105
R2815 VDDA.n3105 VDDA.n3017 3.4105
R2816 VDDA.n3099 VDDA.n3017 3.4105
R2817 VDDA.n3107 VDDA.n3017 3.4105
R2818 VDDA.n3098 VDDA.n3017 3.4105
R2819 VDDA.n3109 VDDA.n3017 3.4105
R2820 VDDA.n3097 VDDA.n3017 3.4105
R2821 VDDA.n3111 VDDA.n3017 3.4105
R2822 VDDA.n3096 VDDA.n3017 3.4105
R2823 VDDA.n3113 VDDA.n3017 3.4105
R2824 VDDA.n3095 VDDA.n3017 3.4105
R2825 VDDA.n3115 VDDA.n3017 3.4105
R2826 VDDA.n3094 VDDA.n3017 3.4105
R2827 VDDA.n3117 VDDA.n3017 3.4105
R2828 VDDA.n3093 VDDA.n3017 3.4105
R2829 VDDA.n3119 VDDA.n3017 3.4105
R2830 VDDA.n3092 VDDA.n3017 3.4105
R2831 VDDA.n3121 VDDA.n3017 3.4105
R2832 VDDA.n3091 VDDA.n3017 3.4105
R2833 VDDA.n3123 VDDA.n3017 3.4105
R2834 VDDA.n3090 VDDA.n3017 3.4105
R2835 VDDA.n3125 VDDA.n3017 3.4105
R2836 VDDA.n3089 VDDA.n3017 3.4105
R2837 VDDA.n3127 VDDA.n3017 3.4105
R2838 VDDA.n3088 VDDA.n3017 3.4105
R2839 VDDA.n3129 VDDA.n3017 3.4105
R2840 VDDA.n3087 VDDA.n3017 3.4105
R2841 VDDA.n3131 VDDA.n3017 3.4105
R2842 VDDA.n3086 VDDA.n3017 3.4105
R2843 VDDA.n3017 VDDA.n18 3.4105
R2844 VDDA.n3133 VDDA.n3017 3.4105
R2845 VDDA.n2970 VDDA.n16 3.4105
R2846 VDDA.n3103 VDDA.n2970 3.4105
R2847 VDDA.n3100 VDDA.n2970 3.4105
R2848 VDDA.n3105 VDDA.n2970 3.4105
R2849 VDDA.n3099 VDDA.n2970 3.4105
R2850 VDDA.n3107 VDDA.n2970 3.4105
R2851 VDDA.n3098 VDDA.n2970 3.4105
R2852 VDDA.n3109 VDDA.n2970 3.4105
R2853 VDDA.n3097 VDDA.n2970 3.4105
R2854 VDDA.n3111 VDDA.n2970 3.4105
R2855 VDDA.n3096 VDDA.n2970 3.4105
R2856 VDDA.n3113 VDDA.n2970 3.4105
R2857 VDDA.n3095 VDDA.n2970 3.4105
R2858 VDDA.n3115 VDDA.n2970 3.4105
R2859 VDDA.n3094 VDDA.n2970 3.4105
R2860 VDDA.n3117 VDDA.n2970 3.4105
R2861 VDDA.n3093 VDDA.n2970 3.4105
R2862 VDDA.n3119 VDDA.n2970 3.4105
R2863 VDDA.n3092 VDDA.n2970 3.4105
R2864 VDDA.n3121 VDDA.n2970 3.4105
R2865 VDDA.n3091 VDDA.n2970 3.4105
R2866 VDDA.n3123 VDDA.n2970 3.4105
R2867 VDDA.n3090 VDDA.n2970 3.4105
R2868 VDDA.n3125 VDDA.n2970 3.4105
R2869 VDDA.n3089 VDDA.n2970 3.4105
R2870 VDDA.n3127 VDDA.n2970 3.4105
R2871 VDDA.n3088 VDDA.n2970 3.4105
R2872 VDDA.n3129 VDDA.n2970 3.4105
R2873 VDDA.n3087 VDDA.n2970 3.4105
R2874 VDDA.n3131 VDDA.n2970 3.4105
R2875 VDDA.n3086 VDDA.n2970 3.4105
R2876 VDDA.n2970 VDDA.n18 3.4105
R2877 VDDA.n3133 VDDA.n2970 3.4105
R2878 VDDA.n3020 VDDA.n16 3.4105
R2879 VDDA.n3103 VDDA.n3020 3.4105
R2880 VDDA.n3100 VDDA.n3020 3.4105
R2881 VDDA.n3105 VDDA.n3020 3.4105
R2882 VDDA.n3099 VDDA.n3020 3.4105
R2883 VDDA.n3107 VDDA.n3020 3.4105
R2884 VDDA.n3098 VDDA.n3020 3.4105
R2885 VDDA.n3109 VDDA.n3020 3.4105
R2886 VDDA.n3097 VDDA.n3020 3.4105
R2887 VDDA.n3111 VDDA.n3020 3.4105
R2888 VDDA.n3096 VDDA.n3020 3.4105
R2889 VDDA.n3113 VDDA.n3020 3.4105
R2890 VDDA.n3095 VDDA.n3020 3.4105
R2891 VDDA.n3115 VDDA.n3020 3.4105
R2892 VDDA.n3094 VDDA.n3020 3.4105
R2893 VDDA.n3117 VDDA.n3020 3.4105
R2894 VDDA.n3093 VDDA.n3020 3.4105
R2895 VDDA.n3119 VDDA.n3020 3.4105
R2896 VDDA.n3092 VDDA.n3020 3.4105
R2897 VDDA.n3121 VDDA.n3020 3.4105
R2898 VDDA.n3091 VDDA.n3020 3.4105
R2899 VDDA.n3123 VDDA.n3020 3.4105
R2900 VDDA.n3090 VDDA.n3020 3.4105
R2901 VDDA.n3125 VDDA.n3020 3.4105
R2902 VDDA.n3089 VDDA.n3020 3.4105
R2903 VDDA.n3127 VDDA.n3020 3.4105
R2904 VDDA.n3088 VDDA.n3020 3.4105
R2905 VDDA.n3129 VDDA.n3020 3.4105
R2906 VDDA.n3087 VDDA.n3020 3.4105
R2907 VDDA.n3131 VDDA.n3020 3.4105
R2908 VDDA.n3086 VDDA.n3020 3.4105
R2909 VDDA.n3020 VDDA.n18 3.4105
R2910 VDDA.n3133 VDDA.n3020 3.4105
R2911 VDDA.n2969 VDDA.n16 3.4105
R2912 VDDA.n3103 VDDA.n2969 3.4105
R2913 VDDA.n3100 VDDA.n2969 3.4105
R2914 VDDA.n3105 VDDA.n2969 3.4105
R2915 VDDA.n3099 VDDA.n2969 3.4105
R2916 VDDA.n3107 VDDA.n2969 3.4105
R2917 VDDA.n3098 VDDA.n2969 3.4105
R2918 VDDA.n3109 VDDA.n2969 3.4105
R2919 VDDA.n3097 VDDA.n2969 3.4105
R2920 VDDA.n3111 VDDA.n2969 3.4105
R2921 VDDA.n3096 VDDA.n2969 3.4105
R2922 VDDA.n3113 VDDA.n2969 3.4105
R2923 VDDA.n3095 VDDA.n2969 3.4105
R2924 VDDA.n3115 VDDA.n2969 3.4105
R2925 VDDA.n3094 VDDA.n2969 3.4105
R2926 VDDA.n3117 VDDA.n2969 3.4105
R2927 VDDA.n3093 VDDA.n2969 3.4105
R2928 VDDA.n3119 VDDA.n2969 3.4105
R2929 VDDA.n3092 VDDA.n2969 3.4105
R2930 VDDA.n3121 VDDA.n2969 3.4105
R2931 VDDA.n3091 VDDA.n2969 3.4105
R2932 VDDA.n3123 VDDA.n2969 3.4105
R2933 VDDA.n3090 VDDA.n2969 3.4105
R2934 VDDA.n3125 VDDA.n2969 3.4105
R2935 VDDA.n3089 VDDA.n2969 3.4105
R2936 VDDA.n3127 VDDA.n2969 3.4105
R2937 VDDA.n3088 VDDA.n2969 3.4105
R2938 VDDA.n3129 VDDA.n2969 3.4105
R2939 VDDA.n3087 VDDA.n2969 3.4105
R2940 VDDA.n3131 VDDA.n2969 3.4105
R2941 VDDA.n3086 VDDA.n2969 3.4105
R2942 VDDA.n2969 VDDA.n18 3.4105
R2943 VDDA.n3133 VDDA.n2969 3.4105
R2944 VDDA.n3023 VDDA.n16 3.4105
R2945 VDDA.n3103 VDDA.n3023 3.4105
R2946 VDDA.n3100 VDDA.n3023 3.4105
R2947 VDDA.n3105 VDDA.n3023 3.4105
R2948 VDDA.n3099 VDDA.n3023 3.4105
R2949 VDDA.n3107 VDDA.n3023 3.4105
R2950 VDDA.n3098 VDDA.n3023 3.4105
R2951 VDDA.n3109 VDDA.n3023 3.4105
R2952 VDDA.n3097 VDDA.n3023 3.4105
R2953 VDDA.n3111 VDDA.n3023 3.4105
R2954 VDDA.n3096 VDDA.n3023 3.4105
R2955 VDDA.n3113 VDDA.n3023 3.4105
R2956 VDDA.n3095 VDDA.n3023 3.4105
R2957 VDDA.n3115 VDDA.n3023 3.4105
R2958 VDDA.n3094 VDDA.n3023 3.4105
R2959 VDDA.n3117 VDDA.n3023 3.4105
R2960 VDDA.n3093 VDDA.n3023 3.4105
R2961 VDDA.n3119 VDDA.n3023 3.4105
R2962 VDDA.n3092 VDDA.n3023 3.4105
R2963 VDDA.n3121 VDDA.n3023 3.4105
R2964 VDDA.n3091 VDDA.n3023 3.4105
R2965 VDDA.n3123 VDDA.n3023 3.4105
R2966 VDDA.n3090 VDDA.n3023 3.4105
R2967 VDDA.n3125 VDDA.n3023 3.4105
R2968 VDDA.n3089 VDDA.n3023 3.4105
R2969 VDDA.n3127 VDDA.n3023 3.4105
R2970 VDDA.n3088 VDDA.n3023 3.4105
R2971 VDDA.n3129 VDDA.n3023 3.4105
R2972 VDDA.n3087 VDDA.n3023 3.4105
R2973 VDDA.n3131 VDDA.n3023 3.4105
R2974 VDDA.n3086 VDDA.n3023 3.4105
R2975 VDDA.n3023 VDDA.n18 3.4105
R2976 VDDA.n3133 VDDA.n3023 3.4105
R2977 VDDA.n2968 VDDA.n16 3.4105
R2978 VDDA.n3103 VDDA.n2968 3.4105
R2979 VDDA.n3100 VDDA.n2968 3.4105
R2980 VDDA.n3105 VDDA.n2968 3.4105
R2981 VDDA.n3099 VDDA.n2968 3.4105
R2982 VDDA.n3107 VDDA.n2968 3.4105
R2983 VDDA.n3098 VDDA.n2968 3.4105
R2984 VDDA.n3109 VDDA.n2968 3.4105
R2985 VDDA.n3097 VDDA.n2968 3.4105
R2986 VDDA.n3111 VDDA.n2968 3.4105
R2987 VDDA.n3096 VDDA.n2968 3.4105
R2988 VDDA.n3113 VDDA.n2968 3.4105
R2989 VDDA.n3095 VDDA.n2968 3.4105
R2990 VDDA.n3115 VDDA.n2968 3.4105
R2991 VDDA.n3094 VDDA.n2968 3.4105
R2992 VDDA.n3117 VDDA.n2968 3.4105
R2993 VDDA.n3093 VDDA.n2968 3.4105
R2994 VDDA.n3119 VDDA.n2968 3.4105
R2995 VDDA.n3092 VDDA.n2968 3.4105
R2996 VDDA.n3121 VDDA.n2968 3.4105
R2997 VDDA.n3091 VDDA.n2968 3.4105
R2998 VDDA.n3123 VDDA.n2968 3.4105
R2999 VDDA.n3090 VDDA.n2968 3.4105
R3000 VDDA.n3125 VDDA.n2968 3.4105
R3001 VDDA.n3089 VDDA.n2968 3.4105
R3002 VDDA.n3127 VDDA.n2968 3.4105
R3003 VDDA.n3088 VDDA.n2968 3.4105
R3004 VDDA.n3129 VDDA.n2968 3.4105
R3005 VDDA.n3087 VDDA.n2968 3.4105
R3006 VDDA.n3131 VDDA.n2968 3.4105
R3007 VDDA.n3086 VDDA.n2968 3.4105
R3008 VDDA.n2968 VDDA.n18 3.4105
R3009 VDDA.n3133 VDDA.n2968 3.4105
R3010 VDDA.n3026 VDDA.n16 3.4105
R3011 VDDA.n3103 VDDA.n3026 3.4105
R3012 VDDA.n3100 VDDA.n3026 3.4105
R3013 VDDA.n3105 VDDA.n3026 3.4105
R3014 VDDA.n3099 VDDA.n3026 3.4105
R3015 VDDA.n3107 VDDA.n3026 3.4105
R3016 VDDA.n3098 VDDA.n3026 3.4105
R3017 VDDA.n3109 VDDA.n3026 3.4105
R3018 VDDA.n3097 VDDA.n3026 3.4105
R3019 VDDA.n3111 VDDA.n3026 3.4105
R3020 VDDA.n3096 VDDA.n3026 3.4105
R3021 VDDA.n3113 VDDA.n3026 3.4105
R3022 VDDA.n3095 VDDA.n3026 3.4105
R3023 VDDA.n3115 VDDA.n3026 3.4105
R3024 VDDA.n3094 VDDA.n3026 3.4105
R3025 VDDA.n3117 VDDA.n3026 3.4105
R3026 VDDA.n3093 VDDA.n3026 3.4105
R3027 VDDA.n3119 VDDA.n3026 3.4105
R3028 VDDA.n3092 VDDA.n3026 3.4105
R3029 VDDA.n3121 VDDA.n3026 3.4105
R3030 VDDA.n3091 VDDA.n3026 3.4105
R3031 VDDA.n3123 VDDA.n3026 3.4105
R3032 VDDA.n3090 VDDA.n3026 3.4105
R3033 VDDA.n3125 VDDA.n3026 3.4105
R3034 VDDA.n3089 VDDA.n3026 3.4105
R3035 VDDA.n3127 VDDA.n3026 3.4105
R3036 VDDA.n3088 VDDA.n3026 3.4105
R3037 VDDA.n3129 VDDA.n3026 3.4105
R3038 VDDA.n3087 VDDA.n3026 3.4105
R3039 VDDA.n3131 VDDA.n3026 3.4105
R3040 VDDA.n3086 VDDA.n3026 3.4105
R3041 VDDA.n3026 VDDA.n18 3.4105
R3042 VDDA.n3133 VDDA.n3026 3.4105
R3043 VDDA.n2967 VDDA.n16 3.4105
R3044 VDDA.n3103 VDDA.n2967 3.4105
R3045 VDDA.n3100 VDDA.n2967 3.4105
R3046 VDDA.n3105 VDDA.n2967 3.4105
R3047 VDDA.n3099 VDDA.n2967 3.4105
R3048 VDDA.n3107 VDDA.n2967 3.4105
R3049 VDDA.n3098 VDDA.n2967 3.4105
R3050 VDDA.n3109 VDDA.n2967 3.4105
R3051 VDDA.n3097 VDDA.n2967 3.4105
R3052 VDDA.n3111 VDDA.n2967 3.4105
R3053 VDDA.n3096 VDDA.n2967 3.4105
R3054 VDDA.n3113 VDDA.n2967 3.4105
R3055 VDDA.n3095 VDDA.n2967 3.4105
R3056 VDDA.n3115 VDDA.n2967 3.4105
R3057 VDDA.n3094 VDDA.n2967 3.4105
R3058 VDDA.n3117 VDDA.n2967 3.4105
R3059 VDDA.n3093 VDDA.n2967 3.4105
R3060 VDDA.n3119 VDDA.n2967 3.4105
R3061 VDDA.n3092 VDDA.n2967 3.4105
R3062 VDDA.n3121 VDDA.n2967 3.4105
R3063 VDDA.n3091 VDDA.n2967 3.4105
R3064 VDDA.n3123 VDDA.n2967 3.4105
R3065 VDDA.n3090 VDDA.n2967 3.4105
R3066 VDDA.n3125 VDDA.n2967 3.4105
R3067 VDDA.n3089 VDDA.n2967 3.4105
R3068 VDDA.n3127 VDDA.n2967 3.4105
R3069 VDDA.n3088 VDDA.n2967 3.4105
R3070 VDDA.n3129 VDDA.n2967 3.4105
R3071 VDDA.n3087 VDDA.n2967 3.4105
R3072 VDDA.n3131 VDDA.n2967 3.4105
R3073 VDDA.n3086 VDDA.n2967 3.4105
R3074 VDDA.n2967 VDDA.n18 3.4105
R3075 VDDA.n3133 VDDA.n2967 3.4105
R3076 VDDA.n3029 VDDA.n16 3.4105
R3077 VDDA.n3103 VDDA.n3029 3.4105
R3078 VDDA.n3100 VDDA.n3029 3.4105
R3079 VDDA.n3105 VDDA.n3029 3.4105
R3080 VDDA.n3099 VDDA.n3029 3.4105
R3081 VDDA.n3107 VDDA.n3029 3.4105
R3082 VDDA.n3098 VDDA.n3029 3.4105
R3083 VDDA.n3109 VDDA.n3029 3.4105
R3084 VDDA.n3097 VDDA.n3029 3.4105
R3085 VDDA.n3111 VDDA.n3029 3.4105
R3086 VDDA.n3096 VDDA.n3029 3.4105
R3087 VDDA.n3113 VDDA.n3029 3.4105
R3088 VDDA.n3095 VDDA.n3029 3.4105
R3089 VDDA.n3115 VDDA.n3029 3.4105
R3090 VDDA.n3094 VDDA.n3029 3.4105
R3091 VDDA.n3117 VDDA.n3029 3.4105
R3092 VDDA.n3093 VDDA.n3029 3.4105
R3093 VDDA.n3119 VDDA.n3029 3.4105
R3094 VDDA.n3092 VDDA.n3029 3.4105
R3095 VDDA.n3121 VDDA.n3029 3.4105
R3096 VDDA.n3091 VDDA.n3029 3.4105
R3097 VDDA.n3123 VDDA.n3029 3.4105
R3098 VDDA.n3090 VDDA.n3029 3.4105
R3099 VDDA.n3125 VDDA.n3029 3.4105
R3100 VDDA.n3089 VDDA.n3029 3.4105
R3101 VDDA.n3127 VDDA.n3029 3.4105
R3102 VDDA.n3088 VDDA.n3029 3.4105
R3103 VDDA.n3129 VDDA.n3029 3.4105
R3104 VDDA.n3087 VDDA.n3029 3.4105
R3105 VDDA.n3131 VDDA.n3029 3.4105
R3106 VDDA.n3086 VDDA.n3029 3.4105
R3107 VDDA.n3029 VDDA.n18 3.4105
R3108 VDDA.n3133 VDDA.n3029 3.4105
R3109 VDDA.n2966 VDDA.n16 3.4105
R3110 VDDA.n3103 VDDA.n2966 3.4105
R3111 VDDA.n3100 VDDA.n2966 3.4105
R3112 VDDA.n3105 VDDA.n2966 3.4105
R3113 VDDA.n3099 VDDA.n2966 3.4105
R3114 VDDA.n3107 VDDA.n2966 3.4105
R3115 VDDA.n3098 VDDA.n2966 3.4105
R3116 VDDA.n3109 VDDA.n2966 3.4105
R3117 VDDA.n3097 VDDA.n2966 3.4105
R3118 VDDA.n3111 VDDA.n2966 3.4105
R3119 VDDA.n3096 VDDA.n2966 3.4105
R3120 VDDA.n3113 VDDA.n2966 3.4105
R3121 VDDA.n3095 VDDA.n2966 3.4105
R3122 VDDA.n3115 VDDA.n2966 3.4105
R3123 VDDA.n3094 VDDA.n2966 3.4105
R3124 VDDA.n3117 VDDA.n2966 3.4105
R3125 VDDA.n3093 VDDA.n2966 3.4105
R3126 VDDA.n3119 VDDA.n2966 3.4105
R3127 VDDA.n3092 VDDA.n2966 3.4105
R3128 VDDA.n3121 VDDA.n2966 3.4105
R3129 VDDA.n3091 VDDA.n2966 3.4105
R3130 VDDA.n3123 VDDA.n2966 3.4105
R3131 VDDA.n3090 VDDA.n2966 3.4105
R3132 VDDA.n3125 VDDA.n2966 3.4105
R3133 VDDA.n3089 VDDA.n2966 3.4105
R3134 VDDA.n3127 VDDA.n2966 3.4105
R3135 VDDA.n3088 VDDA.n2966 3.4105
R3136 VDDA.n3129 VDDA.n2966 3.4105
R3137 VDDA.n3087 VDDA.n2966 3.4105
R3138 VDDA.n3131 VDDA.n2966 3.4105
R3139 VDDA.n3086 VDDA.n2966 3.4105
R3140 VDDA.n2966 VDDA.n18 3.4105
R3141 VDDA.n3133 VDDA.n2966 3.4105
R3142 VDDA.n3032 VDDA.n16 3.4105
R3143 VDDA.n3103 VDDA.n3032 3.4105
R3144 VDDA.n3100 VDDA.n3032 3.4105
R3145 VDDA.n3105 VDDA.n3032 3.4105
R3146 VDDA.n3099 VDDA.n3032 3.4105
R3147 VDDA.n3107 VDDA.n3032 3.4105
R3148 VDDA.n3098 VDDA.n3032 3.4105
R3149 VDDA.n3109 VDDA.n3032 3.4105
R3150 VDDA.n3097 VDDA.n3032 3.4105
R3151 VDDA.n3111 VDDA.n3032 3.4105
R3152 VDDA.n3096 VDDA.n3032 3.4105
R3153 VDDA.n3113 VDDA.n3032 3.4105
R3154 VDDA.n3095 VDDA.n3032 3.4105
R3155 VDDA.n3115 VDDA.n3032 3.4105
R3156 VDDA.n3094 VDDA.n3032 3.4105
R3157 VDDA.n3117 VDDA.n3032 3.4105
R3158 VDDA.n3093 VDDA.n3032 3.4105
R3159 VDDA.n3119 VDDA.n3032 3.4105
R3160 VDDA.n3092 VDDA.n3032 3.4105
R3161 VDDA.n3121 VDDA.n3032 3.4105
R3162 VDDA.n3091 VDDA.n3032 3.4105
R3163 VDDA.n3123 VDDA.n3032 3.4105
R3164 VDDA.n3090 VDDA.n3032 3.4105
R3165 VDDA.n3125 VDDA.n3032 3.4105
R3166 VDDA.n3089 VDDA.n3032 3.4105
R3167 VDDA.n3127 VDDA.n3032 3.4105
R3168 VDDA.n3088 VDDA.n3032 3.4105
R3169 VDDA.n3129 VDDA.n3032 3.4105
R3170 VDDA.n3087 VDDA.n3032 3.4105
R3171 VDDA.n3131 VDDA.n3032 3.4105
R3172 VDDA.n3086 VDDA.n3032 3.4105
R3173 VDDA.n3032 VDDA.n18 3.4105
R3174 VDDA.n3133 VDDA.n3032 3.4105
R3175 VDDA.n2965 VDDA.n16 3.4105
R3176 VDDA.n3103 VDDA.n2965 3.4105
R3177 VDDA.n3100 VDDA.n2965 3.4105
R3178 VDDA.n3105 VDDA.n2965 3.4105
R3179 VDDA.n3099 VDDA.n2965 3.4105
R3180 VDDA.n3107 VDDA.n2965 3.4105
R3181 VDDA.n3098 VDDA.n2965 3.4105
R3182 VDDA.n3109 VDDA.n2965 3.4105
R3183 VDDA.n3097 VDDA.n2965 3.4105
R3184 VDDA.n3111 VDDA.n2965 3.4105
R3185 VDDA.n3096 VDDA.n2965 3.4105
R3186 VDDA.n3113 VDDA.n2965 3.4105
R3187 VDDA.n3095 VDDA.n2965 3.4105
R3188 VDDA.n3115 VDDA.n2965 3.4105
R3189 VDDA.n3094 VDDA.n2965 3.4105
R3190 VDDA.n3117 VDDA.n2965 3.4105
R3191 VDDA.n3093 VDDA.n2965 3.4105
R3192 VDDA.n3119 VDDA.n2965 3.4105
R3193 VDDA.n3092 VDDA.n2965 3.4105
R3194 VDDA.n3121 VDDA.n2965 3.4105
R3195 VDDA.n3091 VDDA.n2965 3.4105
R3196 VDDA.n3123 VDDA.n2965 3.4105
R3197 VDDA.n3090 VDDA.n2965 3.4105
R3198 VDDA.n3125 VDDA.n2965 3.4105
R3199 VDDA.n3089 VDDA.n2965 3.4105
R3200 VDDA.n3127 VDDA.n2965 3.4105
R3201 VDDA.n3088 VDDA.n2965 3.4105
R3202 VDDA.n3129 VDDA.n2965 3.4105
R3203 VDDA.n3087 VDDA.n2965 3.4105
R3204 VDDA.n3131 VDDA.n2965 3.4105
R3205 VDDA.n3086 VDDA.n2965 3.4105
R3206 VDDA.n2965 VDDA.n18 3.4105
R3207 VDDA.n3133 VDDA.n2965 3.4105
R3208 VDDA.n3035 VDDA.n16 3.4105
R3209 VDDA.n3103 VDDA.n3035 3.4105
R3210 VDDA.n3100 VDDA.n3035 3.4105
R3211 VDDA.n3105 VDDA.n3035 3.4105
R3212 VDDA.n3099 VDDA.n3035 3.4105
R3213 VDDA.n3107 VDDA.n3035 3.4105
R3214 VDDA.n3098 VDDA.n3035 3.4105
R3215 VDDA.n3109 VDDA.n3035 3.4105
R3216 VDDA.n3097 VDDA.n3035 3.4105
R3217 VDDA.n3111 VDDA.n3035 3.4105
R3218 VDDA.n3096 VDDA.n3035 3.4105
R3219 VDDA.n3113 VDDA.n3035 3.4105
R3220 VDDA.n3095 VDDA.n3035 3.4105
R3221 VDDA.n3115 VDDA.n3035 3.4105
R3222 VDDA.n3094 VDDA.n3035 3.4105
R3223 VDDA.n3117 VDDA.n3035 3.4105
R3224 VDDA.n3093 VDDA.n3035 3.4105
R3225 VDDA.n3119 VDDA.n3035 3.4105
R3226 VDDA.n3092 VDDA.n3035 3.4105
R3227 VDDA.n3121 VDDA.n3035 3.4105
R3228 VDDA.n3091 VDDA.n3035 3.4105
R3229 VDDA.n3123 VDDA.n3035 3.4105
R3230 VDDA.n3090 VDDA.n3035 3.4105
R3231 VDDA.n3125 VDDA.n3035 3.4105
R3232 VDDA.n3089 VDDA.n3035 3.4105
R3233 VDDA.n3127 VDDA.n3035 3.4105
R3234 VDDA.n3088 VDDA.n3035 3.4105
R3235 VDDA.n3129 VDDA.n3035 3.4105
R3236 VDDA.n3087 VDDA.n3035 3.4105
R3237 VDDA.n3131 VDDA.n3035 3.4105
R3238 VDDA.n3086 VDDA.n3035 3.4105
R3239 VDDA.n3035 VDDA.n18 3.4105
R3240 VDDA.n3133 VDDA.n3035 3.4105
R3241 VDDA.n2964 VDDA.n16 3.4105
R3242 VDDA.n3103 VDDA.n2964 3.4105
R3243 VDDA.n3100 VDDA.n2964 3.4105
R3244 VDDA.n3105 VDDA.n2964 3.4105
R3245 VDDA.n3099 VDDA.n2964 3.4105
R3246 VDDA.n3107 VDDA.n2964 3.4105
R3247 VDDA.n3098 VDDA.n2964 3.4105
R3248 VDDA.n3109 VDDA.n2964 3.4105
R3249 VDDA.n3097 VDDA.n2964 3.4105
R3250 VDDA.n3111 VDDA.n2964 3.4105
R3251 VDDA.n3096 VDDA.n2964 3.4105
R3252 VDDA.n3113 VDDA.n2964 3.4105
R3253 VDDA.n3095 VDDA.n2964 3.4105
R3254 VDDA.n3115 VDDA.n2964 3.4105
R3255 VDDA.n3094 VDDA.n2964 3.4105
R3256 VDDA.n3117 VDDA.n2964 3.4105
R3257 VDDA.n3093 VDDA.n2964 3.4105
R3258 VDDA.n3119 VDDA.n2964 3.4105
R3259 VDDA.n3092 VDDA.n2964 3.4105
R3260 VDDA.n3121 VDDA.n2964 3.4105
R3261 VDDA.n3091 VDDA.n2964 3.4105
R3262 VDDA.n3123 VDDA.n2964 3.4105
R3263 VDDA.n3090 VDDA.n2964 3.4105
R3264 VDDA.n3125 VDDA.n2964 3.4105
R3265 VDDA.n3089 VDDA.n2964 3.4105
R3266 VDDA.n3127 VDDA.n2964 3.4105
R3267 VDDA.n3088 VDDA.n2964 3.4105
R3268 VDDA.n3129 VDDA.n2964 3.4105
R3269 VDDA.n3087 VDDA.n2964 3.4105
R3270 VDDA.n3131 VDDA.n2964 3.4105
R3271 VDDA.n3086 VDDA.n2964 3.4105
R3272 VDDA.n2964 VDDA.n18 3.4105
R3273 VDDA.n3133 VDDA.n2964 3.4105
R3274 VDDA.n3038 VDDA.n16 3.4105
R3275 VDDA.n3103 VDDA.n3038 3.4105
R3276 VDDA.n3100 VDDA.n3038 3.4105
R3277 VDDA.n3105 VDDA.n3038 3.4105
R3278 VDDA.n3099 VDDA.n3038 3.4105
R3279 VDDA.n3107 VDDA.n3038 3.4105
R3280 VDDA.n3098 VDDA.n3038 3.4105
R3281 VDDA.n3109 VDDA.n3038 3.4105
R3282 VDDA.n3097 VDDA.n3038 3.4105
R3283 VDDA.n3111 VDDA.n3038 3.4105
R3284 VDDA.n3096 VDDA.n3038 3.4105
R3285 VDDA.n3113 VDDA.n3038 3.4105
R3286 VDDA.n3095 VDDA.n3038 3.4105
R3287 VDDA.n3115 VDDA.n3038 3.4105
R3288 VDDA.n3094 VDDA.n3038 3.4105
R3289 VDDA.n3117 VDDA.n3038 3.4105
R3290 VDDA.n3093 VDDA.n3038 3.4105
R3291 VDDA.n3119 VDDA.n3038 3.4105
R3292 VDDA.n3092 VDDA.n3038 3.4105
R3293 VDDA.n3121 VDDA.n3038 3.4105
R3294 VDDA.n3091 VDDA.n3038 3.4105
R3295 VDDA.n3123 VDDA.n3038 3.4105
R3296 VDDA.n3090 VDDA.n3038 3.4105
R3297 VDDA.n3125 VDDA.n3038 3.4105
R3298 VDDA.n3089 VDDA.n3038 3.4105
R3299 VDDA.n3127 VDDA.n3038 3.4105
R3300 VDDA.n3088 VDDA.n3038 3.4105
R3301 VDDA.n3129 VDDA.n3038 3.4105
R3302 VDDA.n3087 VDDA.n3038 3.4105
R3303 VDDA.n3131 VDDA.n3038 3.4105
R3304 VDDA.n3086 VDDA.n3038 3.4105
R3305 VDDA.n3038 VDDA.n18 3.4105
R3306 VDDA.n3133 VDDA.n3038 3.4105
R3307 VDDA.n2963 VDDA.n16 3.4105
R3308 VDDA.n3103 VDDA.n2963 3.4105
R3309 VDDA.n3100 VDDA.n2963 3.4105
R3310 VDDA.n3105 VDDA.n2963 3.4105
R3311 VDDA.n3099 VDDA.n2963 3.4105
R3312 VDDA.n3107 VDDA.n2963 3.4105
R3313 VDDA.n3098 VDDA.n2963 3.4105
R3314 VDDA.n3109 VDDA.n2963 3.4105
R3315 VDDA.n3097 VDDA.n2963 3.4105
R3316 VDDA.n3111 VDDA.n2963 3.4105
R3317 VDDA.n3096 VDDA.n2963 3.4105
R3318 VDDA.n3113 VDDA.n2963 3.4105
R3319 VDDA.n3095 VDDA.n2963 3.4105
R3320 VDDA.n3115 VDDA.n2963 3.4105
R3321 VDDA.n3094 VDDA.n2963 3.4105
R3322 VDDA.n3117 VDDA.n2963 3.4105
R3323 VDDA.n3093 VDDA.n2963 3.4105
R3324 VDDA.n3119 VDDA.n2963 3.4105
R3325 VDDA.n3092 VDDA.n2963 3.4105
R3326 VDDA.n3121 VDDA.n2963 3.4105
R3327 VDDA.n3091 VDDA.n2963 3.4105
R3328 VDDA.n3123 VDDA.n2963 3.4105
R3329 VDDA.n3090 VDDA.n2963 3.4105
R3330 VDDA.n3125 VDDA.n2963 3.4105
R3331 VDDA.n3089 VDDA.n2963 3.4105
R3332 VDDA.n3127 VDDA.n2963 3.4105
R3333 VDDA.n3088 VDDA.n2963 3.4105
R3334 VDDA.n3129 VDDA.n2963 3.4105
R3335 VDDA.n3087 VDDA.n2963 3.4105
R3336 VDDA.n3131 VDDA.n2963 3.4105
R3337 VDDA.n3086 VDDA.n2963 3.4105
R3338 VDDA.n2963 VDDA.n18 3.4105
R3339 VDDA.n3133 VDDA.n2963 3.4105
R3340 VDDA.n3041 VDDA.n16 3.4105
R3341 VDDA.n3103 VDDA.n3041 3.4105
R3342 VDDA.n3100 VDDA.n3041 3.4105
R3343 VDDA.n3105 VDDA.n3041 3.4105
R3344 VDDA.n3099 VDDA.n3041 3.4105
R3345 VDDA.n3107 VDDA.n3041 3.4105
R3346 VDDA.n3098 VDDA.n3041 3.4105
R3347 VDDA.n3109 VDDA.n3041 3.4105
R3348 VDDA.n3097 VDDA.n3041 3.4105
R3349 VDDA.n3111 VDDA.n3041 3.4105
R3350 VDDA.n3096 VDDA.n3041 3.4105
R3351 VDDA.n3113 VDDA.n3041 3.4105
R3352 VDDA.n3095 VDDA.n3041 3.4105
R3353 VDDA.n3115 VDDA.n3041 3.4105
R3354 VDDA.n3094 VDDA.n3041 3.4105
R3355 VDDA.n3117 VDDA.n3041 3.4105
R3356 VDDA.n3093 VDDA.n3041 3.4105
R3357 VDDA.n3119 VDDA.n3041 3.4105
R3358 VDDA.n3092 VDDA.n3041 3.4105
R3359 VDDA.n3121 VDDA.n3041 3.4105
R3360 VDDA.n3091 VDDA.n3041 3.4105
R3361 VDDA.n3123 VDDA.n3041 3.4105
R3362 VDDA.n3090 VDDA.n3041 3.4105
R3363 VDDA.n3125 VDDA.n3041 3.4105
R3364 VDDA.n3089 VDDA.n3041 3.4105
R3365 VDDA.n3127 VDDA.n3041 3.4105
R3366 VDDA.n3088 VDDA.n3041 3.4105
R3367 VDDA.n3129 VDDA.n3041 3.4105
R3368 VDDA.n3087 VDDA.n3041 3.4105
R3369 VDDA.n3131 VDDA.n3041 3.4105
R3370 VDDA.n3086 VDDA.n3041 3.4105
R3371 VDDA.n3041 VDDA.n18 3.4105
R3372 VDDA.n3133 VDDA.n3041 3.4105
R3373 VDDA.n2962 VDDA.n16 3.4105
R3374 VDDA.n3103 VDDA.n2962 3.4105
R3375 VDDA.n3100 VDDA.n2962 3.4105
R3376 VDDA.n3105 VDDA.n2962 3.4105
R3377 VDDA.n3099 VDDA.n2962 3.4105
R3378 VDDA.n3107 VDDA.n2962 3.4105
R3379 VDDA.n3098 VDDA.n2962 3.4105
R3380 VDDA.n3109 VDDA.n2962 3.4105
R3381 VDDA.n3097 VDDA.n2962 3.4105
R3382 VDDA.n3111 VDDA.n2962 3.4105
R3383 VDDA.n3096 VDDA.n2962 3.4105
R3384 VDDA.n3113 VDDA.n2962 3.4105
R3385 VDDA.n3095 VDDA.n2962 3.4105
R3386 VDDA.n3115 VDDA.n2962 3.4105
R3387 VDDA.n3094 VDDA.n2962 3.4105
R3388 VDDA.n3117 VDDA.n2962 3.4105
R3389 VDDA.n3093 VDDA.n2962 3.4105
R3390 VDDA.n3119 VDDA.n2962 3.4105
R3391 VDDA.n3092 VDDA.n2962 3.4105
R3392 VDDA.n3121 VDDA.n2962 3.4105
R3393 VDDA.n3091 VDDA.n2962 3.4105
R3394 VDDA.n3123 VDDA.n2962 3.4105
R3395 VDDA.n3090 VDDA.n2962 3.4105
R3396 VDDA.n3125 VDDA.n2962 3.4105
R3397 VDDA.n3089 VDDA.n2962 3.4105
R3398 VDDA.n3127 VDDA.n2962 3.4105
R3399 VDDA.n3088 VDDA.n2962 3.4105
R3400 VDDA.n3129 VDDA.n2962 3.4105
R3401 VDDA.n3087 VDDA.n2962 3.4105
R3402 VDDA.n3131 VDDA.n2962 3.4105
R3403 VDDA.n3086 VDDA.n2962 3.4105
R3404 VDDA.n2962 VDDA.n18 3.4105
R3405 VDDA.n3133 VDDA.n2962 3.4105
R3406 VDDA.n3044 VDDA.n16 3.4105
R3407 VDDA.n3103 VDDA.n3044 3.4105
R3408 VDDA.n3100 VDDA.n3044 3.4105
R3409 VDDA.n3105 VDDA.n3044 3.4105
R3410 VDDA.n3099 VDDA.n3044 3.4105
R3411 VDDA.n3107 VDDA.n3044 3.4105
R3412 VDDA.n3098 VDDA.n3044 3.4105
R3413 VDDA.n3109 VDDA.n3044 3.4105
R3414 VDDA.n3097 VDDA.n3044 3.4105
R3415 VDDA.n3111 VDDA.n3044 3.4105
R3416 VDDA.n3096 VDDA.n3044 3.4105
R3417 VDDA.n3113 VDDA.n3044 3.4105
R3418 VDDA.n3095 VDDA.n3044 3.4105
R3419 VDDA.n3115 VDDA.n3044 3.4105
R3420 VDDA.n3094 VDDA.n3044 3.4105
R3421 VDDA.n3117 VDDA.n3044 3.4105
R3422 VDDA.n3093 VDDA.n3044 3.4105
R3423 VDDA.n3119 VDDA.n3044 3.4105
R3424 VDDA.n3092 VDDA.n3044 3.4105
R3425 VDDA.n3121 VDDA.n3044 3.4105
R3426 VDDA.n3091 VDDA.n3044 3.4105
R3427 VDDA.n3123 VDDA.n3044 3.4105
R3428 VDDA.n3090 VDDA.n3044 3.4105
R3429 VDDA.n3125 VDDA.n3044 3.4105
R3430 VDDA.n3089 VDDA.n3044 3.4105
R3431 VDDA.n3127 VDDA.n3044 3.4105
R3432 VDDA.n3088 VDDA.n3044 3.4105
R3433 VDDA.n3129 VDDA.n3044 3.4105
R3434 VDDA.n3087 VDDA.n3044 3.4105
R3435 VDDA.n3131 VDDA.n3044 3.4105
R3436 VDDA.n3086 VDDA.n3044 3.4105
R3437 VDDA.n3044 VDDA.n18 3.4105
R3438 VDDA.n3133 VDDA.n3044 3.4105
R3439 VDDA.n2961 VDDA.n16 3.4105
R3440 VDDA.n3103 VDDA.n2961 3.4105
R3441 VDDA.n3100 VDDA.n2961 3.4105
R3442 VDDA.n3105 VDDA.n2961 3.4105
R3443 VDDA.n3099 VDDA.n2961 3.4105
R3444 VDDA.n3107 VDDA.n2961 3.4105
R3445 VDDA.n3098 VDDA.n2961 3.4105
R3446 VDDA.n3109 VDDA.n2961 3.4105
R3447 VDDA.n3097 VDDA.n2961 3.4105
R3448 VDDA.n3111 VDDA.n2961 3.4105
R3449 VDDA.n3096 VDDA.n2961 3.4105
R3450 VDDA.n3113 VDDA.n2961 3.4105
R3451 VDDA.n3095 VDDA.n2961 3.4105
R3452 VDDA.n3115 VDDA.n2961 3.4105
R3453 VDDA.n3094 VDDA.n2961 3.4105
R3454 VDDA.n3117 VDDA.n2961 3.4105
R3455 VDDA.n3093 VDDA.n2961 3.4105
R3456 VDDA.n3119 VDDA.n2961 3.4105
R3457 VDDA.n3092 VDDA.n2961 3.4105
R3458 VDDA.n3121 VDDA.n2961 3.4105
R3459 VDDA.n3091 VDDA.n2961 3.4105
R3460 VDDA.n3123 VDDA.n2961 3.4105
R3461 VDDA.n3090 VDDA.n2961 3.4105
R3462 VDDA.n3125 VDDA.n2961 3.4105
R3463 VDDA.n3089 VDDA.n2961 3.4105
R3464 VDDA.n3127 VDDA.n2961 3.4105
R3465 VDDA.n3088 VDDA.n2961 3.4105
R3466 VDDA.n3129 VDDA.n2961 3.4105
R3467 VDDA.n3087 VDDA.n2961 3.4105
R3468 VDDA.n3131 VDDA.n2961 3.4105
R3469 VDDA.n3086 VDDA.n2961 3.4105
R3470 VDDA.n2961 VDDA.n18 3.4105
R3471 VDDA.n3133 VDDA.n2961 3.4105
R3472 VDDA.n3047 VDDA.n16 3.4105
R3473 VDDA.n3103 VDDA.n3047 3.4105
R3474 VDDA.n3100 VDDA.n3047 3.4105
R3475 VDDA.n3105 VDDA.n3047 3.4105
R3476 VDDA.n3099 VDDA.n3047 3.4105
R3477 VDDA.n3107 VDDA.n3047 3.4105
R3478 VDDA.n3098 VDDA.n3047 3.4105
R3479 VDDA.n3109 VDDA.n3047 3.4105
R3480 VDDA.n3097 VDDA.n3047 3.4105
R3481 VDDA.n3111 VDDA.n3047 3.4105
R3482 VDDA.n3096 VDDA.n3047 3.4105
R3483 VDDA.n3113 VDDA.n3047 3.4105
R3484 VDDA.n3095 VDDA.n3047 3.4105
R3485 VDDA.n3115 VDDA.n3047 3.4105
R3486 VDDA.n3094 VDDA.n3047 3.4105
R3487 VDDA.n3117 VDDA.n3047 3.4105
R3488 VDDA.n3093 VDDA.n3047 3.4105
R3489 VDDA.n3119 VDDA.n3047 3.4105
R3490 VDDA.n3092 VDDA.n3047 3.4105
R3491 VDDA.n3121 VDDA.n3047 3.4105
R3492 VDDA.n3091 VDDA.n3047 3.4105
R3493 VDDA.n3123 VDDA.n3047 3.4105
R3494 VDDA.n3090 VDDA.n3047 3.4105
R3495 VDDA.n3125 VDDA.n3047 3.4105
R3496 VDDA.n3089 VDDA.n3047 3.4105
R3497 VDDA.n3127 VDDA.n3047 3.4105
R3498 VDDA.n3088 VDDA.n3047 3.4105
R3499 VDDA.n3129 VDDA.n3047 3.4105
R3500 VDDA.n3087 VDDA.n3047 3.4105
R3501 VDDA.n3131 VDDA.n3047 3.4105
R3502 VDDA.n3086 VDDA.n3047 3.4105
R3503 VDDA.n3047 VDDA.n18 3.4105
R3504 VDDA.n3133 VDDA.n3047 3.4105
R3505 VDDA.n2960 VDDA.n16 3.4105
R3506 VDDA.n3103 VDDA.n2960 3.4105
R3507 VDDA.n3100 VDDA.n2960 3.4105
R3508 VDDA.n3105 VDDA.n2960 3.4105
R3509 VDDA.n3099 VDDA.n2960 3.4105
R3510 VDDA.n3107 VDDA.n2960 3.4105
R3511 VDDA.n3098 VDDA.n2960 3.4105
R3512 VDDA.n3109 VDDA.n2960 3.4105
R3513 VDDA.n3097 VDDA.n2960 3.4105
R3514 VDDA.n3111 VDDA.n2960 3.4105
R3515 VDDA.n3096 VDDA.n2960 3.4105
R3516 VDDA.n3113 VDDA.n2960 3.4105
R3517 VDDA.n3095 VDDA.n2960 3.4105
R3518 VDDA.n3115 VDDA.n2960 3.4105
R3519 VDDA.n3094 VDDA.n2960 3.4105
R3520 VDDA.n3117 VDDA.n2960 3.4105
R3521 VDDA.n3093 VDDA.n2960 3.4105
R3522 VDDA.n3119 VDDA.n2960 3.4105
R3523 VDDA.n3092 VDDA.n2960 3.4105
R3524 VDDA.n3121 VDDA.n2960 3.4105
R3525 VDDA.n3091 VDDA.n2960 3.4105
R3526 VDDA.n3123 VDDA.n2960 3.4105
R3527 VDDA.n3090 VDDA.n2960 3.4105
R3528 VDDA.n3125 VDDA.n2960 3.4105
R3529 VDDA.n3089 VDDA.n2960 3.4105
R3530 VDDA.n3127 VDDA.n2960 3.4105
R3531 VDDA.n3088 VDDA.n2960 3.4105
R3532 VDDA.n3129 VDDA.n2960 3.4105
R3533 VDDA.n3087 VDDA.n2960 3.4105
R3534 VDDA.n3131 VDDA.n2960 3.4105
R3535 VDDA.n3086 VDDA.n2960 3.4105
R3536 VDDA.n2960 VDDA.n18 3.4105
R3537 VDDA.n3133 VDDA.n2960 3.4105
R3538 VDDA.n3050 VDDA.n16 3.4105
R3539 VDDA.n3103 VDDA.n3050 3.4105
R3540 VDDA.n3100 VDDA.n3050 3.4105
R3541 VDDA.n3105 VDDA.n3050 3.4105
R3542 VDDA.n3099 VDDA.n3050 3.4105
R3543 VDDA.n3107 VDDA.n3050 3.4105
R3544 VDDA.n3098 VDDA.n3050 3.4105
R3545 VDDA.n3109 VDDA.n3050 3.4105
R3546 VDDA.n3097 VDDA.n3050 3.4105
R3547 VDDA.n3111 VDDA.n3050 3.4105
R3548 VDDA.n3096 VDDA.n3050 3.4105
R3549 VDDA.n3113 VDDA.n3050 3.4105
R3550 VDDA.n3095 VDDA.n3050 3.4105
R3551 VDDA.n3115 VDDA.n3050 3.4105
R3552 VDDA.n3094 VDDA.n3050 3.4105
R3553 VDDA.n3117 VDDA.n3050 3.4105
R3554 VDDA.n3093 VDDA.n3050 3.4105
R3555 VDDA.n3119 VDDA.n3050 3.4105
R3556 VDDA.n3092 VDDA.n3050 3.4105
R3557 VDDA.n3121 VDDA.n3050 3.4105
R3558 VDDA.n3091 VDDA.n3050 3.4105
R3559 VDDA.n3123 VDDA.n3050 3.4105
R3560 VDDA.n3090 VDDA.n3050 3.4105
R3561 VDDA.n3125 VDDA.n3050 3.4105
R3562 VDDA.n3089 VDDA.n3050 3.4105
R3563 VDDA.n3127 VDDA.n3050 3.4105
R3564 VDDA.n3088 VDDA.n3050 3.4105
R3565 VDDA.n3129 VDDA.n3050 3.4105
R3566 VDDA.n3087 VDDA.n3050 3.4105
R3567 VDDA.n3131 VDDA.n3050 3.4105
R3568 VDDA.n3086 VDDA.n3050 3.4105
R3569 VDDA.n3050 VDDA.n18 3.4105
R3570 VDDA.n3133 VDDA.n3050 3.4105
R3571 VDDA.n2959 VDDA.n16 3.4105
R3572 VDDA.n3103 VDDA.n2959 3.4105
R3573 VDDA.n3100 VDDA.n2959 3.4105
R3574 VDDA.n3105 VDDA.n2959 3.4105
R3575 VDDA.n3099 VDDA.n2959 3.4105
R3576 VDDA.n3107 VDDA.n2959 3.4105
R3577 VDDA.n3098 VDDA.n2959 3.4105
R3578 VDDA.n3109 VDDA.n2959 3.4105
R3579 VDDA.n3097 VDDA.n2959 3.4105
R3580 VDDA.n3111 VDDA.n2959 3.4105
R3581 VDDA.n3096 VDDA.n2959 3.4105
R3582 VDDA.n3113 VDDA.n2959 3.4105
R3583 VDDA.n3095 VDDA.n2959 3.4105
R3584 VDDA.n3115 VDDA.n2959 3.4105
R3585 VDDA.n3094 VDDA.n2959 3.4105
R3586 VDDA.n3117 VDDA.n2959 3.4105
R3587 VDDA.n3093 VDDA.n2959 3.4105
R3588 VDDA.n3119 VDDA.n2959 3.4105
R3589 VDDA.n3092 VDDA.n2959 3.4105
R3590 VDDA.n3121 VDDA.n2959 3.4105
R3591 VDDA.n3091 VDDA.n2959 3.4105
R3592 VDDA.n3123 VDDA.n2959 3.4105
R3593 VDDA.n3090 VDDA.n2959 3.4105
R3594 VDDA.n3125 VDDA.n2959 3.4105
R3595 VDDA.n3089 VDDA.n2959 3.4105
R3596 VDDA.n3127 VDDA.n2959 3.4105
R3597 VDDA.n3088 VDDA.n2959 3.4105
R3598 VDDA.n3129 VDDA.n2959 3.4105
R3599 VDDA.n3087 VDDA.n2959 3.4105
R3600 VDDA.n3131 VDDA.n2959 3.4105
R3601 VDDA.n3086 VDDA.n2959 3.4105
R3602 VDDA.n2959 VDDA.n18 3.4105
R3603 VDDA.n3133 VDDA.n2959 3.4105
R3604 VDDA.n3053 VDDA.n16 3.4105
R3605 VDDA.n3103 VDDA.n3053 3.4105
R3606 VDDA.n3100 VDDA.n3053 3.4105
R3607 VDDA.n3105 VDDA.n3053 3.4105
R3608 VDDA.n3099 VDDA.n3053 3.4105
R3609 VDDA.n3107 VDDA.n3053 3.4105
R3610 VDDA.n3098 VDDA.n3053 3.4105
R3611 VDDA.n3109 VDDA.n3053 3.4105
R3612 VDDA.n3097 VDDA.n3053 3.4105
R3613 VDDA.n3111 VDDA.n3053 3.4105
R3614 VDDA.n3096 VDDA.n3053 3.4105
R3615 VDDA.n3113 VDDA.n3053 3.4105
R3616 VDDA.n3095 VDDA.n3053 3.4105
R3617 VDDA.n3115 VDDA.n3053 3.4105
R3618 VDDA.n3094 VDDA.n3053 3.4105
R3619 VDDA.n3117 VDDA.n3053 3.4105
R3620 VDDA.n3093 VDDA.n3053 3.4105
R3621 VDDA.n3119 VDDA.n3053 3.4105
R3622 VDDA.n3092 VDDA.n3053 3.4105
R3623 VDDA.n3121 VDDA.n3053 3.4105
R3624 VDDA.n3091 VDDA.n3053 3.4105
R3625 VDDA.n3123 VDDA.n3053 3.4105
R3626 VDDA.n3090 VDDA.n3053 3.4105
R3627 VDDA.n3125 VDDA.n3053 3.4105
R3628 VDDA.n3089 VDDA.n3053 3.4105
R3629 VDDA.n3127 VDDA.n3053 3.4105
R3630 VDDA.n3088 VDDA.n3053 3.4105
R3631 VDDA.n3129 VDDA.n3053 3.4105
R3632 VDDA.n3087 VDDA.n3053 3.4105
R3633 VDDA.n3131 VDDA.n3053 3.4105
R3634 VDDA.n3086 VDDA.n3053 3.4105
R3635 VDDA.n3053 VDDA.n18 3.4105
R3636 VDDA.n3133 VDDA.n3053 3.4105
R3637 VDDA.n2958 VDDA.n16 3.4105
R3638 VDDA.n3103 VDDA.n2958 3.4105
R3639 VDDA.n3100 VDDA.n2958 3.4105
R3640 VDDA.n3105 VDDA.n2958 3.4105
R3641 VDDA.n3099 VDDA.n2958 3.4105
R3642 VDDA.n3107 VDDA.n2958 3.4105
R3643 VDDA.n3098 VDDA.n2958 3.4105
R3644 VDDA.n3109 VDDA.n2958 3.4105
R3645 VDDA.n3097 VDDA.n2958 3.4105
R3646 VDDA.n3111 VDDA.n2958 3.4105
R3647 VDDA.n3096 VDDA.n2958 3.4105
R3648 VDDA.n3113 VDDA.n2958 3.4105
R3649 VDDA.n3095 VDDA.n2958 3.4105
R3650 VDDA.n3115 VDDA.n2958 3.4105
R3651 VDDA.n3094 VDDA.n2958 3.4105
R3652 VDDA.n3117 VDDA.n2958 3.4105
R3653 VDDA.n3093 VDDA.n2958 3.4105
R3654 VDDA.n3119 VDDA.n2958 3.4105
R3655 VDDA.n3092 VDDA.n2958 3.4105
R3656 VDDA.n3121 VDDA.n2958 3.4105
R3657 VDDA.n3091 VDDA.n2958 3.4105
R3658 VDDA.n3123 VDDA.n2958 3.4105
R3659 VDDA.n3090 VDDA.n2958 3.4105
R3660 VDDA.n3125 VDDA.n2958 3.4105
R3661 VDDA.n3089 VDDA.n2958 3.4105
R3662 VDDA.n3127 VDDA.n2958 3.4105
R3663 VDDA.n3088 VDDA.n2958 3.4105
R3664 VDDA.n3129 VDDA.n2958 3.4105
R3665 VDDA.n3087 VDDA.n2958 3.4105
R3666 VDDA.n3131 VDDA.n2958 3.4105
R3667 VDDA.n3086 VDDA.n2958 3.4105
R3668 VDDA.n2958 VDDA.n18 3.4105
R3669 VDDA.n3133 VDDA.n2958 3.4105
R3670 VDDA.n3056 VDDA.n16 3.4105
R3671 VDDA.n3103 VDDA.n3056 3.4105
R3672 VDDA.n3100 VDDA.n3056 3.4105
R3673 VDDA.n3105 VDDA.n3056 3.4105
R3674 VDDA.n3099 VDDA.n3056 3.4105
R3675 VDDA.n3107 VDDA.n3056 3.4105
R3676 VDDA.n3098 VDDA.n3056 3.4105
R3677 VDDA.n3109 VDDA.n3056 3.4105
R3678 VDDA.n3097 VDDA.n3056 3.4105
R3679 VDDA.n3111 VDDA.n3056 3.4105
R3680 VDDA.n3096 VDDA.n3056 3.4105
R3681 VDDA.n3113 VDDA.n3056 3.4105
R3682 VDDA.n3095 VDDA.n3056 3.4105
R3683 VDDA.n3115 VDDA.n3056 3.4105
R3684 VDDA.n3094 VDDA.n3056 3.4105
R3685 VDDA.n3117 VDDA.n3056 3.4105
R3686 VDDA.n3093 VDDA.n3056 3.4105
R3687 VDDA.n3119 VDDA.n3056 3.4105
R3688 VDDA.n3092 VDDA.n3056 3.4105
R3689 VDDA.n3121 VDDA.n3056 3.4105
R3690 VDDA.n3091 VDDA.n3056 3.4105
R3691 VDDA.n3123 VDDA.n3056 3.4105
R3692 VDDA.n3090 VDDA.n3056 3.4105
R3693 VDDA.n3125 VDDA.n3056 3.4105
R3694 VDDA.n3089 VDDA.n3056 3.4105
R3695 VDDA.n3127 VDDA.n3056 3.4105
R3696 VDDA.n3088 VDDA.n3056 3.4105
R3697 VDDA.n3129 VDDA.n3056 3.4105
R3698 VDDA.n3087 VDDA.n3056 3.4105
R3699 VDDA.n3131 VDDA.n3056 3.4105
R3700 VDDA.n3086 VDDA.n3056 3.4105
R3701 VDDA.n3056 VDDA.n18 3.4105
R3702 VDDA.n3133 VDDA.n3056 3.4105
R3703 VDDA.n2957 VDDA.n16 3.4105
R3704 VDDA.n3103 VDDA.n2957 3.4105
R3705 VDDA.n3100 VDDA.n2957 3.4105
R3706 VDDA.n3105 VDDA.n2957 3.4105
R3707 VDDA.n3099 VDDA.n2957 3.4105
R3708 VDDA.n3107 VDDA.n2957 3.4105
R3709 VDDA.n3098 VDDA.n2957 3.4105
R3710 VDDA.n3109 VDDA.n2957 3.4105
R3711 VDDA.n3097 VDDA.n2957 3.4105
R3712 VDDA.n3111 VDDA.n2957 3.4105
R3713 VDDA.n3096 VDDA.n2957 3.4105
R3714 VDDA.n3113 VDDA.n2957 3.4105
R3715 VDDA.n3095 VDDA.n2957 3.4105
R3716 VDDA.n3115 VDDA.n2957 3.4105
R3717 VDDA.n3094 VDDA.n2957 3.4105
R3718 VDDA.n3117 VDDA.n2957 3.4105
R3719 VDDA.n3093 VDDA.n2957 3.4105
R3720 VDDA.n3119 VDDA.n2957 3.4105
R3721 VDDA.n3092 VDDA.n2957 3.4105
R3722 VDDA.n3121 VDDA.n2957 3.4105
R3723 VDDA.n3091 VDDA.n2957 3.4105
R3724 VDDA.n3123 VDDA.n2957 3.4105
R3725 VDDA.n3090 VDDA.n2957 3.4105
R3726 VDDA.n3125 VDDA.n2957 3.4105
R3727 VDDA.n3089 VDDA.n2957 3.4105
R3728 VDDA.n3127 VDDA.n2957 3.4105
R3729 VDDA.n3088 VDDA.n2957 3.4105
R3730 VDDA.n3129 VDDA.n2957 3.4105
R3731 VDDA.n3087 VDDA.n2957 3.4105
R3732 VDDA.n3131 VDDA.n2957 3.4105
R3733 VDDA.n3086 VDDA.n2957 3.4105
R3734 VDDA.n2957 VDDA.n18 3.4105
R3735 VDDA.n3133 VDDA.n2957 3.4105
R3736 VDDA.n3059 VDDA.n16 3.4105
R3737 VDDA.n3103 VDDA.n3059 3.4105
R3738 VDDA.n3100 VDDA.n3059 3.4105
R3739 VDDA.n3105 VDDA.n3059 3.4105
R3740 VDDA.n3099 VDDA.n3059 3.4105
R3741 VDDA.n3107 VDDA.n3059 3.4105
R3742 VDDA.n3098 VDDA.n3059 3.4105
R3743 VDDA.n3109 VDDA.n3059 3.4105
R3744 VDDA.n3097 VDDA.n3059 3.4105
R3745 VDDA.n3111 VDDA.n3059 3.4105
R3746 VDDA.n3096 VDDA.n3059 3.4105
R3747 VDDA.n3113 VDDA.n3059 3.4105
R3748 VDDA.n3095 VDDA.n3059 3.4105
R3749 VDDA.n3115 VDDA.n3059 3.4105
R3750 VDDA.n3094 VDDA.n3059 3.4105
R3751 VDDA.n3117 VDDA.n3059 3.4105
R3752 VDDA.n3093 VDDA.n3059 3.4105
R3753 VDDA.n3119 VDDA.n3059 3.4105
R3754 VDDA.n3092 VDDA.n3059 3.4105
R3755 VDDA.n3121 VDDA.n3059 3.4105
R3756 VDDA.n3091 VDDA.n3059 3.4105
R3757 VDDA.n3123 VDDA.n3059 3.4105
R3758 VDDA.n3090 VDDA.n3059 3.4105
R3759 VDDA.n3125 VDDA.n3059 3.4105
R3760 VDDA.n3089 VDDA.n3059 3.4105
R3761 VDDA.n3127 VDDA.n3059 3.4105
R3762 VDDA.n3088 VDDA.n3059 3.4105
R3763 VDDA.n3129 VDDA.n3059 3.4105
R3764 VDDA.n3087 VDDA.n3059 3.4105
R3765 VDDA.n3131 VDDA.n3059 3.4105
R3766 VDDA.n3086 VDDA.n3059 3.4105
R3767 VDDA.n3059 VDDA.n18 3.4105
R3768 VDDA.n3133 VDDA.n3059 3.4105
R3769 VDDA.n2956 VDDA.n16 3.4105
R3770 VDDA.n3103 VDDA.n2956 3.4105
R3771 VDDA.n3100 VDDA.n2956 3.4105
R3772 VDDA.n3105 VDDA.n2956 3.4105
R3773 VDDA.n3099 VDDA.n2956 3.4105
R3774 VDDA.n3107 VDDA.n2956 3.4105
R3775 VDDA.n3098 VDDA.n2956 3.4105
R3776 VDDA.n3109 VDDA.n2956 3.4105
R3777 VDDA.n3097 VDDA.n2956 3.4105
R3778 VDDA.n3111 VDDA.n2956 3.4105
R3779 VDDA.n3096 VDDA.n2956 3.4105
R3780 VDDA.n3113 VDDA.n2956 3.4105
R3781 VDDA.n3095 VDDA.n2956 3.4105
R3782 VDDA.n3115 VDDA.n2956 3.4105
R3783 VDDA.n3094 VDDA.n2956 3.4105
R3784 VDDA.n3117 VDDA.n2956 3.4105
R3785 VDDA.n3093 VDDA.n2956 3.4105
R3786 VDDA.n3119 VDDA.n2956 3.4105
R3787 VDDA.n3092 VDDA.n2956 3.4105
R3788 VDDA.n3121 VDDA.n2956 3.4105
R3789 VDDA.n3091 VDDA.n2956 3.4105
R3790 VDDA.n3123 VDDA.n2956 3.4105
R3791 VDDA.n3090 VDDA.n2956 3.4105
R3792 VDDA.n3125 VDDA.n2956 3.4105
R3793 VDDA.n3089 VDDA.n2956 3.4105
R3794 VDDA.n3127 VDDA.n2956 3.4105
R3795 VDDA.n3088 VDDA.n2956 3.4105
R3796 VDDA.n3129 VDDA.n2956 3.4105
R3797 VDDA.n3087 VDDA.n2956 3.4105
R3798 VDDA.n3131 VDDA.n2956 3.4105
R3799 VDDA.n3086 VDDA.n2956 3.4105
R3800 VDDA.n2956 VDDA.n18 3.4105
R3801 VDDA.n3133 VDDA.n2956 3.4105
R3802 VDDA.n3062 VDDA.n16 3.4105
R3803 VDDA.n3103 VDDA.n3062 3.4105
R3804 VDDA.n3100 VDDA.n3062 3.4105
R3805 VDDA.n3105 VDDA.n3062 3.4105
R3806 VDDA.n3099 VDDA.n3062 3.4105
R3807 VDDA.n3107 VDDA.n3062 3.4105
R3808 VDDA.n3098 VDDA.n3062 3.4105
R3809 VDDA.n3109 VDDA.n3062 3.4105
R3810 VDDA.n3097 VDDA.n3062 3.4105
R3811 VDDA.n3111 VDDA.n3062 3.4105
R3812 VDDA.n3096 VDDA.n3062 3.4105
R3813 VDDA.n3113 VDDA.n3062 3.4105
R3814 VDDA.n3095 VDDA.n3062 3.4105
R3815 VDDA.n3115 VDDA.n3062 3.4105
R3816 VDDA.n3094 VDDA.n3062 3.4105
R3817 VDDA.n3117 VDDA.n3062 3.4105
R3818 VDDA.n3093 VDDA.n3062 3.4105
R3819 VDDA.n3119 VDDA.n3062 3.4105
R3820 VDDA.n3092 VDDA.n3062 3.4105
R3821 VDDA.n3121 VDDA.n3062 3.4105
R3822 VDDA.n3091 VDDA.n3062 3.4105
R3823 VDDA.n3123 VDDA.n3062 3.4105
R3824 VDDA.n3090 VDDA.n3062 3.4105
R3825 VDDA.n3125 VDDA.n3062 3.4105
R3826 VDDA.n3089 VDDA.n3062 3.4105
R3827 VDDA.n3127 VDDA.n3062 3.4105
R3828 VDDA.n3088 VDDA.n3062 3.4105
R3829 VDDA.n3129 VDDA.n3062 3.4105
R3830 VDDA.n3087 VDDA.n3062 3.4105
R3831 VDDA.n3131 VDDA.n3062 3.4105
R3832 VDDA.n3086 VDDA.n3062 3.4105
R3833 VDDA.n3062 VDDA.n18 3.4105
R3834 VDDA.n3133 VDDA.n3062 3.4105
R3835 VDDA.n2955 VDDA.n16 3.4105
R3836 VDDA.n3103 VDDA.n2955 3.4105
R3837 VDDA.n3100 VDDA.n2955 3.4105
R3838 VDDA.n3105 VDDA.n2955 3.4105
R3839 VDDA.n3099 VDDA.n2955 3.4105
R3840 VDDA.n3107 VDDA.n2955 3.4105
R3841 VDDA.n3098 VDDA.n2955 3.4105
R3842 VDDA.n3109 VDDA.n2955 3.4105
R3843 VDDA.n3097 VDDA.n2955 3.4105
R3844 VDDA.n3111 VDDA.n2955 3.4105
R3845 VDDA.n3096 VDDA.n2955 3.4105
R3846 VDDA.n3113 VDDA.n2955 3.4105
R3847 VDDA.n3095 VDDA.n2955 3.4105
R3848 VDDA.n3115 VDDA.n2955 3.4105
R3849 VDDA.n3094 VDDA.n2955 3.4105
R3850 VDDA.n3117 VDDA.n2955 3.4105
R3851 VDDA.n3093 VDDA.n2955 3.4105
R3852 VDDA.n3119 VDDA.n2955 3.4105
R3853 VDDA.n3092 VDDA.n2955 3.4105
R3854 VDDA.n3121 VDDA.n2955 3.4105
R3855 VDDA.n3091 VDDA.n2955 3.4105
R3856 VDDA.n3123 VDDA.n2955 3.4105
R3857 VDDA.n3090 VDDA.n2955 3.4105
R3858 VDDA.n3125 VDDA.n2955 3.4105
R3859 VDDA.n3089 VDDA.n2955 3.4105
R3860 VDDA.n3127 VDDA.n2955 3.4105
R3861 VDDA.n3088 VDDA.n2955 3.4105
R3862 VDDA.n3129 VDDA.n2955 3.4105
R3863 VDDA.n3087 VDDA.n2955 3.4105
R3864 VDDA.n3131 VDDA.n2955 3.4105
R3865 VDDA.n3086 VDDA.n2955 3.4105
R3866 VDDA.n2955 VDDA.n18 3.4105
R3867 VDDA.n3133 VDDA.n2955 3.4105
R3868 VDDA.n3065 VDDA.n16 3.4105
R3869 VDDA.n3103 VDDA.n3065 3.4105
R3870 VDDA.n3100 VDDA.n3065 3.4105
R3871 VDDA.n3105 VDDA.n3065 3.4105
R3872 VDDA.n3099 VDDA.n3065 3.4105
R3873 VDDA.n3107 VDDA.n3065 3.4105
R3874 VDDA.n3098 VDDA.n3065 3.4105
R3875 VDDA.n3109 VDDA.n3065 3.4105
R3876 VDDA.n3097 VDDA.n3065 3.4105
R3877 VDDA.n3111 VDDA.n3065 3.4105
R3878 VDDA.n3096 VDDA.n3065 3.4105
R3879 VDDA.n3113 VDDA.n3065 3.4105
R3880 VDDA.n3095 VDDA.n3065 3.4105
R3881 VDDA.n3115 VDDA.n3065 3.4105
R3882 VDDA.n3094 VDDA.n3065 3.4105
R3883 VDDA.n3117 VDDA.n3065 3.4105
R3884 VDDA.n3093 VDDA.n3065 3.4105
R3885 VDDA.n3119 VDDA.n3065 3.4105
R3886 VDDA.n3092 VDDA.n3065 3.4105
R3887 VDDA.n3121 VDDA.n3065 3.4105
R3888 VDDA.n3091 VDDA.n3065 3.4105
R3889 VDDA.n3123 VDDA.n3065 3.4105
R3890 VDDA.n3090 VDDA.n3065 3.4105
R3891 VDDA.n3125 VDDA.n3065 3.4105
R3892 VDDA.n3089 VDDA.n3065 3.4105
R3893 VDDA.n3127 VDDA.n3065 3.4105
R3894 VDDA.n3088 VDDA.n3065 3.4105
R3895 VDDA.n3129 VDDA.n3065 3.4105
R3896 VDDA.n3087 VDDA.n3065 3.4105
R3897 VDDA.n3131 VDDA.n3065 3.4105
R3898 VDDA.n3086 VDDA.n3065 3.4105
R3899 VDDA.n3065 VDDA.n18 3.4105
R3900 VDDA.n3133 VDDA.n3065 3.4105
R3901 VDDA.n2954 VDDA.n16 3.4105
R3902 VDDA.n3103 VDDA.n2954 3.4105
R3903 VDDA.n3100 VDDA.n2954 3.4105
R3904 VDDA.n3105 VDDA.n2954 3.4105
R3905 VDDA.n3099 VDDA.n2954 3.4105
R3906 VDDA.n3107 VDDA.n2954 3.4105
R3907 VDDA.n3098 VDDA.n2954 3.4105
R3908 VDDA.n3109 VDDA.n2954 3.4105
R3909 VDDA.n3097 VDDA.n2954 3.4105
R3910 VDDA.n3111 VDDA.n2954 3.4105
R3911 VDDA.n3096 VDDA.n2954 3.4105
R3912 VDDA.n3113 VDDA.n2954 3.4105
R3913 VDDA.n3095 VDDA.n2954 3.4105
R3914 VDDA.n3115 VDDA.n2954 3.4105
R3915 VDDA.n3094 VDDA.n2954 3.4105
R3916 VDDA.n3117 VDDA.n2954 3.4105
R3917 VDDA.n3093 VDDA.n2954 3.4105
R3918 VDDA.n3119 VDDA.n2954 3.4105
R3919 VDDA.n3092 VDDA.n2954 3.4105
R3920 VDDA.n3121 VDDA.n2954 3.4105
R3921 VDDA.n3091 VDDA.n2954 3.4105
R3922 VDDA.n3123 VDDA.n2954 3.4105
R3923 VDDA.n3090 VDDA.n2954 3.4105
R3924 VDDA.n3125 VDDA.n2954 3.4105
R3925 VDDA.n3089 VDDA.n2954 3.4105
R3926 VDDA.n3127 VDDA.n2954 3.4105
R3927 VDDA.n3088 VDDA.n2954 3.4105
R3928 VDDA.n3129 VDDA.n2954 3.4105
R3929 VDDA.n3087 VDDA.n2954 3.4105
R3930 VDDA.n3131 VDDA.n2954 3.4105
R3931 VDDA.n3086 VDDA.n2954 3.4105
R3932 VDDA.n2954 VDDA.n18 3.4105
R3933 VDDA.n3133 VDDA.n2954 3.4105
R3934 VDDA.n3068 VDDA.n16 3.4105
R3935 VDDA.n3103 VDDA.n3068 3.4105
R3936 VDDA.n3100 VDDA.n3068 3.4105
R3937 VDDA.n3105 VDDA.n3068 3.4105
R3938 VDDA.n3099 VDDA.n3068 3.4105
R3939 VDDA.n3107 VDDA.n3068 3.4105
R3940 VDDA.n3098 VDDA.n3068 3.4105
R3941 VDDA.n3109 VDDA.n3068 3.4105
R3942 VDDA.n3097 VDDA.n3068 3.4105
R3943 VDDA.n3111 VDDA.n3068 3.4105
R3944 VDDA.n3096 VDDA.n3068 3.4105
R3945 VDDA.n3113 VDDA.n3068 3.4105
R3946 VDDA.n3095 VDDA.n3068 3.4105
R3947 VDDA.n3115 VDDA.n3068 3.4105
R3948 VDDA.n3094 VDDA.n3068 3.4105
R3949 VDDA.n3117 VDDA.n3068 3.4105
R3950 VDDA.n3093 VDDA.n3068 3.4105
R3951 VDDA.n3119 VDDA.n3068 3.4105
R3952 VDDA.n3092 VDDA.n3068 3.4105
R3953 VDDA.n3121 VDDA.n3068 3.4105
R3954 VDDA.n3091 VDDA.n3068 3.4105
R3955 VDDA.n3123 VDDA.n3068 3.4105
R3956 VDDA.n3090 VDDA.n3068 3.4105
R3957 VDDA.n3125 VDDA.n3068 3.4105
R3958 VDDA.n3089 VDDA.n3068 3.4105
R3959 VDDA.n3127 VDDA.n3068 3.4105
R3960 VDDA.n3088 VDDA.n3068 3.4105
R3961 VDDA.n3129 VDDA.n3068 3.4105
R3962 VDDA.n3087 VDDA.n3068 3.4105
R3963 VDDA.n3131 VDDA.n3068 3.4105
R3964 VDDA.n3086 VDDA.n3068 3.4105
R3965 VDDA.n3068 VDDA.n18 3.4105
R3966 VDDA.n3133 VDDA.n3068 3.4105
R3967 VDDA.n2953 VDDA.n16 3.4105
R3968 VDDA.n3103 VDDA.n2953 3.4105
R3969 VDDA.n3100 VDDA.n2953 3.4105
R3970 VDDA.n3105 VDDA.n2953 3.4105
R3971 VDDA.n3099 VDDA.n2953 3.4105
R3972 VDDA.n3107 VDDA.n2953 3.4105
R3973 VDDA.n3098 VDDA.n2953 3.4105
R3974 VDDA.n3109 VDDA.n2953 3.4105
R3975 VDDA.n3097 VDDA.n2953 3.4105
R3976 VDDA.n3111 VDDA.n2953 3.4105
R3977 VDDA.n3096 VDDA.n2953 3.4105
R3978 VDDA.n3113 VDDA.n2953 3.4105
R3979 VDDA.n3095 VDDA.n2953 3.4105
R3980 VDDA.n3115 VDDA.n2953 3.4105
R3981 VDDA.n3094 VDDA.n2953 3.4105
R3982 VDDA.n3117 VDDA.n2953 3.4105
R3983 VDDA.n3093 VDDA.n2953 3.4105
R3984 VDDA.n3119 VDDA.n2953 3.4105
R3985 VDDA.n3092 VDDA.n2953 3.4105
R3986 VDDA.n3121 VDDA.n2953 3.4105
R3987 VDDA.n3091 VDDA.n2953 3.4105
R3988 VDDA.n3123 VDDA.n2953 3.4105
R3989 VDDA.n3090 VDDA.n2953 3.4105
R3990 VDDA.n3125 VDDA.n2953 3.4105
R3991 VDDA.n3089 VDDA.n2953 3.4105
R3992 VDDA.n3127 VDDA.n2953 3.4105
R3993 VDDA.n3088 VDDA.n2953 3.4105
R3994 VDDA.n3129 VDDA.n2953 3.4105
R3995 VDDA.n3087 VDDA.n2953 3.4105
R3996 VDDA.n3131 VDDA.n2953 3.4105
R3997 VDDA.n3086 VDDA.n2953 3.4105
R3998 VDDA.n2953 VDDA.n18 3.4105
R3999 VDDA.n3133 VDDA.n2953 3.4105
R4000 VDDA.n3071 VDDA.n16 3.4105
R4001 VDDA.n3103 VDDA.n3071 3.4105
R4002 VDDA.n3100 VDDA.n3071 3.4105
R4003 VDDA.n3105 VDDA.n3071 3.4105
R4004 VDDA.n3099 VDDA.n3071 3.4105
R4005 VDDA.n3107 VDDA.n3071 3.4105
R4006 VDDA.n3098 VDDA.n3071 3.4105
R4007 VDDA.n3109 VDDA.n3071 3.4105
R4008 VDDA.n3097 VDDA.n3071 3.4105
R4009 VDDA.n3111 VDDA.n3071 3.4105
R4010 VDDA.n3096 VDDA.n3071 3.4105
R4011 VDDA.n3113 VDDA.n3071 3.4105
R4012 VDDA.n3095 VDDA.n3071 3.4105
R4013 VDDA.n3115 VDDA.n3071 3.4105
R4014 VDDA.n3094 VDDA.n3071 3.4105
R4015 VDDA.n3117 VDDA.n3071 3.4105
R4016 VDDA.n3093 VDDA.n3071 3.4105
R4017 VDDA.n3119 VDDA.n3071 3.4105
R4018 VDDA.n3092 VDDA.n3071 3.4105
R4019 VDDA.n3121 VDDA.n3071 3.4105
R4020 VDDA.n3091 VDDA.n3071 3.4105
R4021 VDDA.n3123 VDDA.n3071 3.4105
R4022 VDDA.n3090 VDDA.n3071 3.4105
R4023 VDDA.n3125 VDDA.n3071 3.4105
R4024 VDDA.n3089 VDDA.n3071 3.4105
R4025 VDDA.n3127 VDDA.n3071 3.4105
R4026 VDDA.n3088 VDDA.n3071 3.4105
R4027 VDDA.n3129 VDDA.n3071 3.4105
R4028 VDDA.n3087 VDDA.n3071 3.4105
R4029 VDDA.n3131 VDDA.n3071 3.4105
R4030 VDDA.n3086 VDDA.n3071 3.4105
R4031 VDDA.n3071 VDDA.n18 3.4105
R4032 VDDA.n3133 VDDA.n3071 3.4105
R4033 VDDA.n2952 VDDA.n16 3.4105
R4034 VDDA.n3103 VDDA.n2952 3.4105
R4035 VDDA.n3100 VDDA.n2952 3.4105
R4036 VDDA.n3105 VDDA.n2952 3.4105
R4037 VDDA.n3099 VDDA.n2952 3.4105
R4038 VDDA.n3107 VDDA.n2952 3.4105
R4039 VDDA.n3098 VDDA.n2952 3.4105
R4040 VDDA.n3109 VDDA.n2952 3.4105
R4041 VDDA.n3097 VDDA.n2952 3.4105
R4042 VDDA.n3111 VDDA.n2952 3.4105
R4043 VDDA.n3096 VDDA.n2952 3.4105
R4044 VDDA.n3113 VDDA.n2952 3.4105
R4045 VDDA.n3095 VDDA.n2952 3.4105
R4046 VDDA.n3115 VDDA.n2952 3.4105
R4047 VDDA.n3094 VDDA.n2952 3.4105
R4048 VDDA.n3117 VDDA.n2952 3.4105
R4049 VDDA.n3093 VDDA.n2952 3.4105
R4050 VDDA.n3119 VDDA.n2952 3.4105
R4051 VDDA.n3092 VDDA.n2952 3.4105
R4052 VDDA.n3121 VDDA.n2952 3.4105
R4053 VDDA.n3091 VDDA.n2952 3.4105
R4054 VDDA.n3123 VDDA.n2952 3.4105
R4055 VDDA.n3090 VDDA.n2952 3.4105
R4056 VDDA.n3125 VDDA.n2952 3.4105
R4057 VDDA.n3089 VDDA.n2952 3.4105
R4058 VDDA.n3127 VDDA.n2952 3.4105
R4059 VDDA.n3088 VDDA.n2952 3.4105
R4060 VDDA.n3129 VDDA.n2952 3.4105
R4061 VDDA.n3087 VDDA.n2952 3.4105
R4062 VDDA.n3131 VDDA.n2952 3.4105
R4063 VDDA.n3086 VDDA.n2952 3.4105
R4064 VDDA.n2952 VDDA.n18 3.4105
R4065 VDDA.n3133 VDDA.n2952 3.4105
R4066 VDDA.n3074 VDDA.n16 3.4105
R4067 VDDA.n3103 VDDA.n3074 3.4105
R4068 VDDA.n3100 VDDA.n3074 3.4105
R4069 VDDA.n3105 VDDA.n3074 3.4105
R4070 VDDA.n3099 VDDA.n3074 3.4105
R4071 VDDA.n3107 VDDA.n3074 3.4105
R4072 VDDA.n3098 VDDA.n3074 3.4105
R4073 VDDA.n3109 VDDA.n3074 3.4105
R4074 VDDA.n3097 VDDA.n3074 3.4105
R4075 VDDA.n3111 VDDA.n3074 3.4105
R4076 VDDA.n3096 VDDA.n3074 3.4105
R4077 VDDA.n3113 VDDA.n3074 3.4105
R4078 VDDA.n3095 VDDA.n3074 3.4105
R4079 VDDA.n3115 VDDA.n3074 3.4105
R4080 VDDA.n3094 VDDA.n3074 3.4105
R4081 VDDA.n3117 VDDA.n3074 3.4105
R4082 VDDA.n3093 VDDA.n3074 3.4105
R4083 VDDA.n3119 VDDA.n3074 3.4105
R4084 VDDA.n3092 VDDA.n3074 3.4105
R4085 VDDA.n3121 VDDA.n3074 3.4105
R4086 VDDA.n3091 VDDA.n3074 3.4105
R4087 VDDA.n3123 VDDA.n3074 3.4105
R4088 VDDA.n3090 VDDA.n3074 3.4105
R4089 VDDA.n3125 VDDA.n3074 3.4105
R4090 VDDA.n3089 VDDA.n3074 3.4105
R4091 VDDA.n3127 VDDA.n3074 3.4105
R4092 VDDA.n3088 VDDA.n3074 3.4105
R4093 VDDA.n3129 VDDA.n3074 3.4105
R4094 VDDA.n3087 VDDA.n3074 3.4105
R4095 VDDA.n3131 VDDA.n3074 3.4105
R4096 VDDA.n3086 VDDA.n3074 3.4105
R4097 VDDA.n3074 VDDA.n18 3.4105
R4098 VDDA.n3133 VDDA.n3074 3.4105
R4099 VDDA.n2951 VDDA.n16 3.4105
R4100 VDDA.n3103 VDDA.n2951 3.4105
R4101 VDDA.n3100 VDDA.n2951 3.4105
R4102 VDDA.n3105 VDDA.n2951 3.4105
R4103 VDDA.n3099 VDDA.n2951 3.4105
R4104 VDDA.n3107 VDDA.n2951 3.4105
R4105 VDDA.n3098 VDDA.n2951 3.4105
R4106 VDDA.n3109 VDDA.n2951 3.4105
R4107 VDDA.n3097 VDDA.n2951 3.4105
R4108 VDDA.n3111 VDDA.n2951 3.4105
R4109 VDDA.n3096 VDDA.n2951 3.4105
R4110 VDDA.n3113 VDDA.n2951 3.4105
R4111 VDDA.n3095 VDDA.n2951 3.4105
R4112 VDDA.n3115 VDDA.n2951 3.4105
R4113 VDDA.n3094 VDDA.n2951 3.4105
R4114 VDDA.n3117 VDDA.n2951 3.4105
R4115 VDDA.n3093 VDDA.n2951 3.4105
R4116 VDDA.n3119 VDDA.n2951 3.4105
R4117 VDDA.n3092 VDDA.n2951 3.4105
R4118 VDDA.n3121 VDDA.n2951 3.4105
R4119 VDDA.n3091 VDDA.n2951 3.4105
R4120 VDDA.n3123 VDDA.n2951 3.4105
R4121 VDDA.n3090 VDDA.n2951 3.4105
R4122 VDDA.n3125 VDDA.n2951 3.4105
R4123 VDDA.n3089 VDDA.n2951 3.4105
R4124 VDDA.n3127 VDDA.n2951 3.4105
R4125 VDDA.n3088 VDDA.n2951 3.4105
R4126 VDDA.n3129 VDDA.n2951 3.4105
R4127 VDDA.n3087 VDDA.n2951 3.4105
R4128 VDDA.n3131 VDDA.n2951 3.4105
R4129 VDDA.n3086 VDDA.n2951 3.4105
R4130 VDDA.n2951 VDDA.n18 3.4105
R4131 VDDA.n3133 VDDA.n2951 3.4105
R4132 VDDA.n3077 VDDA.n16 3.4105
R4133 VDDA.n3103 VDDA.n3077 3.4105
R4134 VDDA.n3100 VDDA.n3077 3.4105
R4135 VDDA.n3105 VDDA.n3077 3.4105
R4136 VDDA.n3099 VDDA.n3077 3.4105
R4137 VDDA.n3107 VDDA.n3077 3.4105
R4138 VDDA.n3098 VDDA.n3077 3.4105
R4139 VDDA.n3109 VDDA.n3077 3.4105
R4140 VDDA.n3097 VDDA.n3077 3.4105
R4141 VDDA.n3111 VDDA.n3077 3.4105
R4142 VDDA.n3096 VDDA.n3077 3.4105
R4143 VDDA.n3113 VDDA.n3077 3.4105
R4144 VDDA.n3095 VDDA.n3077 3.4105
R4145 VDDA.n3115 VDDA.n3077 3.4105
R4146 VDDA.n3094 VDDA.n3077 3.4105
R4147 VDDA.n3117 VDDA.n3077 3.4105
R4148 VDDA.n3093 VDDA.n3077 3.4105
R4149 VDDA.n3119 VDDA.n3077 3.4105
R4150 VDDA.n3092 VDDA.n3077 3.4105
R4151 VDDA.n3121 VDDA.n3077 3.4105
R4152 VDDA.n3091 VDDA.n3077 3.4105
R4153 VDDA.n3123 VDDA.n3077 3.4105
R4154 VDDA.n3090 VDDA.n3077 3.4105
R4155 VDDA.n3125 VDDA.n3077 3.4105
R4156 VDDA.n3089 VDDA.n3077 3.4105
R4157 VDDA.n3127 VDDA.n3077 3.4105
R4158 VDDA.n3088 VDDA.n3077 3.4105
R4159 VDDA.n3129 VDDA.n3077 3.4105
R4160 VDDA.n3087 VDDA.n3077 3.4105
R4161 VDDA.n3131 VDDA.n3077 3.4105
R4162 VDDA.n3086 VDDA.n3077 3.4105
R4163 VDDA.n3077 VDDA.n18 3.4105
R4164 VDDA.n3133 VDDA.n3077 3.4105
R4165 VDDA.n2950 VDDA.n16 3.4105
R4166 VDDA.n3103 VDDA.n2950 3.4105
R4167 VDDA.n3100 VDDA.n2950 3.4105
R4168 VDDA.n3105 VDDA.n2950 3.4105
R4169 VDDA.n3099 VDDA.n2950 3.4105
R4170 VDDA.n3107 VDDA.n2950 3.4105
R4171 VDDA.n3098 VDDA.n2950 3.4105
R4172 VDDA.n3109 VDDA.n2950 3.4105
R4173 VDDA.n3097 VDDA.n2950 3.4105
R4174 VDDA.n3111 VDDA.n2950 3.4105
R4175 VDDA.n3096 VDDA.n2950 3.4105
R4176 VDDA.n3113 VDDA.n2950 3.4105
R4177 VDDA.n3095 VDDA.n2950 3.4105
R4178 VDDA.n3115 VDDA.n2950 3.4105
R4179 VDDA.n3094 VDDA.n2950 3.4105
R4180 VDDA.n3117 VDDA.n2950 3.4105
R4181 VDDA.n3093 VDDA.n2950 3.4105
R4182 VDDA.n3119 VDDA.n2950 3.4105
R4183 VDDA.n3092 VDDA.n2950 3.4105
R4184 VDDA.n3121 VDDA.n2950 3.4105
R4185 VDDA.n3091 VDDA.n2950 3.4105
R4186 VDDA.n3123 VDDA.n2950 3.4105
R4187 VDDA.n3090 VDDA.n2950 3.4105
R4188 VDDA.n3125 VDDA.n2950 3.4105
R4189 VDDA.n3089 VDDA.n2950 3.4105
R4190 VDDA.n3127 VDDA.n2950 3.4105
R4191 VDDA.n3088 VDDA.n2950 3.4105
R4192 VDDA.n3129 VDDA.n2950 3.4105
R4193 VDDA.n3087 VDDA.n2950 3.4105
R4194 VDDA.n3131 VDDA.n2950 3.4105
R4195 VDDA.n3086 VDDA.n2950 3.4105
R4196 VDDA.n2950 VDDA.n18 3.4105
R4197 VDDA.n3133 VDDA.n2950 3.4105
R4198 VDDA.n3080 VDDA.n16 3.4105
R4199 VDDA.n3103 VDDA.n3080 3.4105
R4200 VDDA.n3100 VDDA.n3080 3.4105
R4201 VDDA.n3105 VDDA.n3080 3.4105
R4202 VDDA.n3099 VDDA.n3080 3.4105
R4203 VDDA.n3107 VDDA.n3080 3.4105
R4204 VDDA.n3098 VDDA.n3080 3.4105
R4205 VDDA.n3109 VDDA.n3080 3.4105
R4206 VDDA.n3097 VDDA.n3080 3.4105
R4207 VDDA.n3111 VDDA.n3080 3.4105
R4208 VDDA.n3096 VDDA.n3080 3.4105
R4209 VDDA.n3113 VDDA.n3080 3.4105
R4210 VDDA.n3095 VDDA.n3080 3.4105
R4211 VDDA.n3115 VDDA.n3080 3.4105
R4212 VDDA.n3094 VDDA.n3080 3.4105
R4213 VDDA.n3117 VDDA.n3080 3.4105
R4214 VDDA.n3093 VDDA.n3080 3.4105
R4215 VDDA.n3119 VDDA.n3080 3.4105
R4216 VDDA.n3092 VDDA.n3080 3.4105
R4217 VDDA.n3121 VDDA.n3080 3.4105
R4218 VDDA.n3091 VDDA.n3080 3.4105
R4219 VDDA.n3123 VDDA.n3080 3.4105
R4220 VDDA.n3090 VDDA.n3080 3.4105
R4221 VDDA.n3125 VDDA.n3080 3.4105
R4222 VDDA.n3089 VDDA.n3080 3.4105
R4223 VDDA.n3127 VDDA.n3080 3.4105
R4224 VDDA.n3088 VDDA.n3080 3.4105
R4225 VDDA.n3129 VDDA.n3080 3.4105
R4226 VDDA.n3087 VDDA.n3080 3.4105
R4227 VDDA.n3131 VDDA.n3080 3.4105
R4228 VDDA.n3086 VDDA.n3080 3.4105
R4229 VDDA.n3080 VDDA.n18 3.4105
R4230 VDDA.n3133 VDDA.n3080 3.4105
R4231 VDDA.n2949 VDDA.n16 3.4105
R4232 VDDA.n3103 VDDA.n2949 3.4105
R4233 VDDA.n3100 VDDA.n2949 3.4105
R4234 VDDA.n3105 VDDA.n2949 3.4105
R4235 VDDA.n3099 VDDA.n2949 3.4105
R4236 VDDA.n3107 VDDA.n2949 3.4105
R4237 VDDA.n3098 VDDA.n2949 3.4105
R4238 VDDA.n3109 VDDA.n2949 3.4105
R4239 VDDA.n3097 VDDA.n2949 3.4105
R4240 VDDA.n3111 VDDA.n2949 3.4105
R4241 VDDA.n3096 VDDA.n2949 3.4105
R4242 VDDA.n3113 VDDA.n2949 3.4105
R4243 VDDA.n3095 VDDA.n2949 3.4105
R4244 VDDA.n3115 VDDA.n2949 3.4105
R4245 VDDA.n3094 VDDA.n2949 3.4105
R4246 VDDA.n3117 VDDA.n2949 3.4105
R4247 VDDA.n3093 VDDA.n2949 3.4105
R4248 VDDA.n3119 VDDA.n2949 3.4105
R4249 VDDA.n3092 VDDA.n2949 3.4105
R4250 VDDA.n3121 VDDA.n2949 3.4105
R4251 VDDA.n3091 VDDA.n2949 3.4105
R4252 VDDA.n3123 VDDA.n2949 3.4105
R4253 VDDA.n3090 VDDA.n2949 3.4105
R4254 VDDA.n3125 VDDA.n2949 3.4105
R4255 VDDA.n3089 VDDA.n2949 3.4105
R4256 VDDA.n3127 VDDA.n2949 3.4105
R4257 VDDA.n3088 VDDA.n2949 3.4105
R4258 VDDA.n3129 VDDA.n2949 3.4105
R4259 VDDA.n3087 VDDA.n2949 3.4105
R4260 VDDA.n3131 VDDA.n2949 3.4105
R4261 VDDA.n3086 VDDA.n2949 3.4105
R4262 VDDA.n2949 VDDA.n18 3.4105
R4263 VDDA.n3133 VDDA.n2949 3.4105
R4264 VDDA.n3083 VDDA.n16 3.4105
R4265 VDDA.n3103 VDDA.n3083 3.4105
R4266 VDDA.n3100 VDDA.n3083 3.4105
R4267 VDDA.n3105 VDDA.n3083 3.4105
R4268 VDDA.n3099 VDDA.n3083 3.4105
R4269 VDDA.n3107 VDDA.n3083 3.4105
R4270 VDDA.n3098 VDDA.n3083 3.4105
R4271 VDDA.n3109 VDDA.n3083 3.4105
R4272 VDDA.n3097 VDDA.n3083 3.4105
R4273 VDDA.n3111 VDDA.n3083 3.4105
R4274 VDDA.n3096 VDDA.n3083 3.4105
R4275 VDDA.n3113 VDDA.n3083 3.4105
R4276 VDDA.n3095 VDDA.n3083 3.4105
R4277 VDDA.n3115 VDDA.n3083 3.4105
R4278 VDDA.n3094 VDDA.n3083 3.4105
R4279 VDDA.n3117 VDDA.n3083 3.4105
R4280 VDDA.n3093 VDDA.n3083 3.4105
R4281 VDDA.n3119 VDDA.n3083 3.4105
R4282 VDDA.n3092 VDDA.n3083 3.4105
R4283 VDDA.n3121 VDDA.n3083 3.4105
R4284 VDDA.n3091 VDDA.n3083 3.4105
R4285 VDDA.n3123 VDDA.n3083 3.4105
R4286 VDDA.n3090 VDDA.n3083 3.4105
R4287 VDDA.n3125 VDDA.n3083 3.4105
R4288 VDDA.n3089 VDDA.n3083 3.4105
R4289 VDDA.n3127 VDDA.n3083 3.4105
R4290 VDDA.n3088 VDDA.n3083 3.4105
R4291 VDDA.n3129 VDDA.n3083 3.4105
R4292 VDDA.n3087 VDDA.n3083 3.4105
R4293 VDDA.n3131 VDDA.n3083 3.4105
R4294 VDDA.n3086 VDDA.n3083 3.4105
R4295 VDDA.n3083 VDDA.n18 3.4105
R4296 VDDA.n3133 VDDA.n3083 3.4105
R4297 VDDA.n2948 VDDA.n16 3.4105
R4298 VDDA.n3103 VDDA.n2948 3.4105
R4299 VDDA.n3100 VDDA.n2948 3.4105
R4300 VDDA.n3105 VDDA.n2948 3.4105
R4301 VDDA.n3099 VDDA.n2948 3.4105
R4302 VDDA.n3107 VDDA.n2948 3.4105
R4303 VDDA.n3098 VDDA.n2948 3.4105
R4304 VDDA.n3109 VDDA.n2948 3.4105
R4305 VDDA.n3097 VDDA.n2948 3.4105
R4306 VDDA.n3111 VDDA.n2948 3.4105
R4307 VDDA.n3096 VDDA.n2948 3.4105
R4308 VDDA.n3113 VDDA.n2948 3.4105
R4309 VDDA.n3095 VDDA.n2948 3.4105
R4310 VDDA.n3115 VDDA.n2948 3.4105
R4311 VDDA.n3094 VDDA.n2948 3.4105
R4312 VDDA.n3117 VDDA.n2948 3.4105
R4313 VDDA.n3093 VDDA.n2948 3.4105
R4314 VDDA.n3119 VDDA.n2948 3.4105
R4315 VDDA.n3092 VDDA.n2948 3.4105
R4316 VDDA.n3121 VDDA.n2948 3.4105
R4317 VDDA.n3091 VDDA.n2948 3.4105
R4318 VDDA.n3123 VDDA.n2948 3.4105
R4319 VDDA.n3090 VDDA.n2948 3.4105
R4320 VDDA.n3125 VDDA.n2948 3.4105
R4321 VDDA.n3089 VDDA.n2948 3.4105
R4322 VDDA.n3127 VDDA.n2948 3.4105
R4323 VDDA.n3088 VDDA.n2948 3.4105
R4324 VDDA.n3129 VDDA.n2948 3.4105
R4325 VDDA.n3087 VDDA.n2948 3.4105
R4326 VDDA.n3131 VDDA.n2948 3.4105
R4327 VDDA.n3086 VDDA.n2948 3.4105
R4328 VDDA.n2948 VDDA.n18 3.4105
R4329 VDDA.n3133 VDDA.n2948 3.4105
R4330 VDDA.n3132 VDDA.n3103 3.4105
R4331 VDDA.n3132 VDDA.n3100 3.4105
R4332 VDDA.n3132 VDDA.n3105 3.4105
R4333 VDDA.n3132 VDDA.n3099 3.4105
R4334 VDDA.n3132 VDDA.n3107 3.4105
R4335 VDDA.n3132 VDDA.n3098 3.4105
R4336 VDDA.n3132 VDDA.n3109 3.4105
R4337 VDDA.n3132 VDDA.n3097 3.4105
R4338 VDDA.n3132 VDDA.n3111 3.4105
R4339 VDDA.n3132 VDDA.n3096 3.4105
R4340 VDDA.n3132 VDDA.n3113 3.4105
R4341 VDDA.n3132 VDDA.n3095 3.4105
R4342 VDDA.n3132 VDDA.n3115 3.4105
R4343 VDDA.n3132 VDDA.n3094 3.4105
R4344 VDDA.n3132 VDDA.n3117 3.4105
R4345 VDDA.n3132 VDDA.n3093 3.4105
R4346 VDDA.n3132 VDDA.n3119 3.4105
R4347 VDDA.n3132 VDDA.n3092 3.4105
R4348 VDDA.n3132 VDDA.n3121 3.4105
R4349 VDDA.n3132 VDDA.n3091 3.4105
R4350 VDDA.n3132 VDDA.n3123 3.4105
R4351 VDDA.n3132 VDDA.n3090 3.4105
R4352 VDDA.n3132 VDDA.n3125 3.4105
R4353 VDDA.n3132 VDDA.n3089 3.4105
R4354 VDDA.n3132 VDDA.n3127 3.4105
R4355 VDDA.n3132 VDDA.n3088 3.4105
R4356 VDDA.n3132 VDDA.n3129 3.4105
R4357 VDDA.n3132 VDDA.n3087 3.4105
R4358 VDDA.n3132 VDDA.n3131 3.4105
R4359 VDDA.n3132 VDDA.n3086 3.4105
R4360 VDDA.n3132 VDDA.n18 3.4105
R4361 VDDA.n3133 VDDA.n3132 3.4105
R4362 VDDA.n1993 VDDA.n1992 3.11118
R4363 VDDA.n2003 VDDA.n2002 3.11118
R4364 VDDA.n386 VDDA.n385 3.06776
R4365 VDDA.n1992 VDDA.n1974 3.04304
R4366 VDDA.n2002 VDDA.n1954 3.04304
R4367 VDDA.n2332 VDDA.n2328 2.96402
R4368 VDDA.n436 VDDA.n432 2.96402
R4369 VDDA.n2369 VDDA.n2368 2.8957
R4370 VDDA.n2370 VDDA.n2369 2.8957
R4371 VDDA.n2374 VDDA.n2372 2.8957
R4372 VDDA.n2377 VDDA.n2372 2.8957
R4373 VDDA.n2373 VDDA.n2370 2.8957
R4374 VDDA.n2377 VDDA.n2376 2.8957
R4375 VDDA.n2379 VDDA.n2368 2.8957
R4376 VDDA.n2374 VDDA.n2373 2.8957
R4377 VDDA.n374 VDDA.n373 2.8255
R4378 VDDA.n376 VDDA.n375 2.8255
R4379 VDDA.n2283 VDDA.n2282 2.53872
R4380 VDDA.n2277 VDDA.n2267 2.53872
R4381 VDDA.n2412 VDDA.n366 2.53694
R4382 VDDA.n2419 VDDA.n2418 2.53694
R4383 VDDA.n2406 VDDA.n2404 2.53694
R4384 VDDA.n2271 VDDA.n453 2.53694
R4385 VDDA.n2331 VDDA.n2330 2.423
R4386 VDDA.n2329 VDDA.n2328 2.423
R4387 VDDA.n433 VDDA.n432 2.423
R4388 VDDA.n435 VDDA.n434 2.423
R4389 VDDA.n1906 VDDA.n1905 2.41009
R4390 VDDA.n1791 VDDA.n1790 2.36299
R4391 VDDA.n2379 VDDA.n2367 2.32777
R4392 VDDA.n93 VDDA.n92 2.30736
R4393 VDDA.n2816 VDDA.n2813 2.30736
R4394 VDDA.n2666 VDDA.n2665 2.30736
R4395 VDDA.n271 VDDA.n270 2.30736
R4396 VDDA.n2468 VDDA.n2465 2.30736
R4397 VDDA.n1228 VDDA.n1227 2.30736
R4398 VDDA.n538 VDDA.n537 2.30736
R4399 VDDA.n1030 VDDA.n1027 2.30736
R4400 VDDA.n880 VDDA.n879 2.30736
R4401 VDDA.n1578 VDDA.n1577 2.30736
R4402 VDDA.n2255 VDDA.n2254 2.30736
R4403 VDDA.n692 VDDA.n691 2.30736
R4404 VDDA.n1766 VDDA.n1404 2.2948
R4405 VDDA.n1767 VDDA.n1766 2.2948
R4406 VDDA.n2332 VDDA.n2331 2.27652
R4407 VDDA.n436 VDDA.n435 2.27652
R4408 VDDA.n1948 VDDA.n1940 2.26187
R4409 VDDA.n2014 VDDA.n1938 2.26187
R4410 VDDA.n2091 VDDA.n1936 2.26187
R4411 VDDA.n2141 VDDA.n1934 2.26187
R4412 VDDA.n429 VDDA.n407 2.26187
R4413 VDDA.n413 VDDA.n410 2.26187
R4414 VDDA.n414 VDDA.n413 2.26187
R4415 VDDA.n2325 VDDA.n2324 2.26187
R4416 VDDA.n806 VDDA.n803 2.26187
R4417 VDDA.n806 VDDA.n805 2.26187
R4418 VDDA.n1945 VDDA.n1940 2.26187
R4419 VDDA.n2326 VDDA.n2325 2.26187
R4420 VDDA.n2337 VDDA.n2336 2.26187
R4421 VDDA.n2287 VDDA.n2286 2.26187
R4422 VDDA.n1765 VDDA.n1405 2.2505
R4423 VDDA.n1764 VDDA.n1763 2.2505
R4424 VDDA.n1407 VDDA.n1406 2.2505
R4425 VDDA.n1585 VDDA.n1582 2.2505
R4426 VDDA.n1755 VDDA.n1754 2.2505
R4427 VDDA.n1753 VDDA.n1584 2.2505
R4428 VDDA.n1752 VDDA.n1751 2.2505
R4429 VDDA.n1587 VDDA.n1586 2.2505
R4430 VDDA.n1745 VDDA.n1744 2.2505
R4431 VDDA.n1743 VDDA.n1591 2.2505
R4432 VDDA.n1742 VDDA.n1741 2.2505
R4433 VDDA.n1593 VDDA.n1592 2.2505
R4434 VDDA.n1735 VDDA.n1734 2.2505
R4435 VDDA.n1733 VDDA.n1597 2.2505
R4436 VDDA.n1732 VDDA.n1731 2.2505
R4437 VDDA.n1599 VDDA.n1598 2.2505
R4438 VDDA.n1725 VDDA.n1724 2.2505
R4439 VDDA.n1723 VDDA.n1603 2.2505
R4440 VDDA.n1722 VDDA.n1721 2.2505
R4441 VDDA.n1605 VDDA.n1604 2.2505
R4442 VDDA.n1715 VDDA.n1714 2.2505
R4443 VDDA.n1713 VDDA.n1609 2.2505
R4444 VDDA.n1712 VDDA.n1711 2.2505
R4445 VDDA.n1611 VDDA.n1610 2.2505
R4446 VDDA.n1705 VDDA.n1704 2.2505
R4447 VDDA.n1703 VDDA.n1615 2.2505
R4448 VDDA.n1702 VDDA.n1701 2.2505
R4449 VDDA.n1617 VDDA.n1616 2.2505
R4450 VDDA.n1695 VDDA.n1694 2.2505
R4451 VDDA.n1693 VDDA.n1621 2.2505
R4452 VDDA.n1692 VDDA.n1691 2.2505
R4453 VDDA.n1623 VDDA.n1622 2.2505
R4454 VDDA.n1685 VDDA.n1684 2.2505
R4455 VDDA.n1683 VDDA.n1627 2.2505
R4456 VDDA.n1682 VDDA.n1681 2.2505
R4457 VDDA.n1629 VDDA.n1628 2.2505
R4458 VDDA.n1675 VDDA.n1674 2.2505
R4459 VDDA.n1673 VDDA.n1633 2.2505
R4460 VDDA.n1672 VDDA.n1671 2.2505
R4461 VDDA.n1635 VDDA.n1634 2.2505
R4462 VDDA.n1665 VDDA.n1664 2.2505
R4463 VDDA.n1663 VDDA.n1639 2.2505
R4464 VDDA.n1662 VDDA.n1661 2.2505
R4465 VDDA.n1641 VDDA.n1640 2.2505
R4466 VDDA.n1655 VDDA.n1654 2.2505
R4467 VDDA.n1653 VDDA.n1645 2.2505
R4468 VDDA.n1949 VDDA.n1939 2.24063
R4469 VDDA.n2015 VDDA.n1937 2.24063
R4470 VDDA.n2092 VDDA.n1935 2.24063
R4471 VDDA.n2142 VDDA.n1933 2.24063
R4472 VDDA.n431 VDDA.n430 2.24063
R4473 VDDA.n2397 VDDA.n2396 2.24063
R4474 VDDA.n406 VDDA.n390 2.24063
R4475 VDDA.n2341 VDDA.n2340 2.24063
R4476 VDDA.n2339 VDDA.n449 2.24063
R4477 VDDA.n2334 VDDA.n2333 2.24063
R4478 VDDA.n2336 VDDA.n2335 2.24063
R4479 VDDA.n2324 VDDA.n2323 2.24063
R4480 VDDA.n981 VDDA.n634 2.24063
R4481 VDDA.n635 VDDA.n633 2.24063
R4482 VDDA.n1152 VDDA.n631 2.24063
R4483 VDDA.n632 VDDA.n630 2.24063
R4484 VDDA.n1156 VDDA.n459 2.24063
R4485 VDDA.n629 VDDA.n628 2.24063
R4486 VDDA.n2286 VDDA.n452 2.24063
R4487 VDDA.n2285 VDDA.n451 2.24063
R4488 VDDA.n2403 VDDA.n369 2.24063
R4489 VDDA.n370 VDDA.n368 2.24063
R4490 VDDA.n2400 VDDA.n2399 2.24063
R4491 VDDA.n2266 VDDA.n457 2.24063
R4492 VDDA.n458 VDDA.n456 2.24063
R4493 VDDA.n2590 VDDA.n364 2.24063
R4494 VDDA.n365 VDDA.n363 2.24063
R4495 VDDA.n2594 VDDA.n192 2.24063
R4496 VDDA.n362 VDDA.n361 2.24063
R4497 VDDA.n2767 VDDA.n190 2.24063
R4498 VDDA.n191 VDDA.n189 2.24063
R4499 VDDA.n2938 VDDA.n187 2.24063
R4500 VDDA.n188 VDDA.n186 2.24063
R4501 VDDA.n2942 VDDA.n2941 2.24063
R4502 VDDA.n185 VDDA.n184 2.24063
R4503 VDDA.n1945 VDDA.n1944 2.24063
R4504 VDDA.n1950 VDDA.n1938 2.24063
R4505 VDDA.n2011 VDDA.n2010 2.24063
R4506 VDDA.n2016 VDDA.n1936 2.24063
R4507 VDDA.n2088 VDDA.n2087 2.24063
R4508 VDDA.n2093 VDDA.n1934 2.24063
R4509 VDDA.n2138 VDDA.n2137 2.24063
R4510 VDDA.n439 VDDA.n407 2.24063
R4511 VDDA.n438 VDDA.n437 2.24063
R4512 VDDA.n428 VDDA.n410 2.24063
R4513 VDDA.n427 VDDA.n426 2.24063
R4514 VDDA.n2398 VDDA.n388 2.24063
R4515 VDDA.n2343 VDDA.n2342 2.24063
R4516 VDDA.n2345 VDDA.n2344 2.24063
R4517 VDDA.n2338 VDDA.n2306 2.24063
R4518 VDDA.n2327 VDDA.n2309 2.24063
R4519 VDDA.n978 VDDA.n977 2.24063
R4520 VDDA.n1149 VDDA.n1148 2.24063
R4521 VDDA.n1157 VDDA.n627 2.24063
R4522 VDDA.n2263 VDDA.n2262 2.24063
R4523 VDDA.n2587 VDDA.n2586 2.24063
R4524 VDDA.n2595 VDDA.n360 2.24063
R4525 VDDA.n2764 VDDA.n2763 2.24063
R4526 VDDA.n2935 VDDA.n2934 2.24063
R4527 VDDA.n2943 VDDA.n182 2.24063
R4528 VDDA.n809 VDDA.n803 2.24063
R4529 VDDA.n808 VDDA.n636 2.24063
R4530 VDDA.n2944 VDDA.n2943 2.16196
R4531 VDDA.n2934 VDDA.n2933 2.16196
R4532 VDDA.n2763 VDDA.n2762 2.16196
R4533 VDDA.n2596 VDDA.n2595 2.16196
R4534 VDDA.n2586 VDDA.n2585 2.16196
R4535 VDDA.n2262 VDDA.n2261 2.16196
R4536 VDDA.n1158 VDDA.n1157 2.16196
R4537 VDDA.n1148 VDDA.n1147 2.16196
R4538 VDDA.n977 VDDA.n976 2.16196
R4539 VDDA.n810 VDDA.n809 2.16196
R4540 VDDA.n385 VDDA.n384 2.12369
R4541 VDDA.n402 VDDA.n401 1.97758
R4542 VDDA.n404 VDDA.n403 1.97758
R4543 VDDA.n2304 VDDA.n2303 1.97758
R4544 VDDA.n2302 VDDA.n2301 1.97758
R4545 VDDA.n401 VDDA.n400 1.95361
R4546 VDDA.n2301 VDDA.n2300 1.95361
R4547 VDDA.n1991 VDDA.n1990 1.90331
R4548 VDDA.n383 VDDA.n382 1.888
R4549 VDDA.n381 VDDA.n380 1.888
R4550 VDDA.n2418 VDDA.n367 1.888
R4551 VDDA.n2406 VDDA.n2405 1.888
R4552 VDDA.n405 VDDA.n404 1.83902
R4553 VDDA.n2305 VDDA.n2304 1.83902
R4554 VDDA.n1999 VDDA.n1998 1.77831
R4555 VDDA.n2001 VDDA.n2000 1.77831
R4556 VDDA.n2009 VDDA.n2008 1.77831
R4557 VDDA.n2143 VDDA.n1321 1.7622
R4558 VDDA.n1652 VDDA.n1646 1.74133
R4559 VDDA.n3134 VDDA.n15 1.70583
R4560 VDDA.n3134 VDDA.n14 1.70583
R4561 VDDA.n3134 VDDA.n13 1.70583
R4562 VDDA.n3134 VDDA.n12 1.70583
R4563 VDDA.n3134 VDDA.n11 1.70583
R4564 VDDA.n3134 VDDA.n10 1.70583
R4565 VDDA.n3134 VDDA.n9 1.70583
R4566 VDDA.n3134 VDDA.n8 1.70583
R4567 VDDA.n3134 VDDA.n7 1.70583
R4568 VDDA.n3134 VDDA.n6 1.70583
R4569 VDDA.n3134 VDDA.n5 1.70583
R4570 VDDA.n3134 VDDA.n4 1.70583
R4571 VDDA.n3134 VDDA.n3 1.70583
R4572 VDDA.n3134 VDDA.n2 1.70583
R4573 VDDA.n3134 VDDA.n1 1.70583
R4574 VDDA.n3102 VDDA.n2984 1.70583
R4575 VDDA.n3104 VDDA.n2984 1.70583
R4576 VDDA.n3106 VDDA.n2984 1.70583
R4577 VDDA.n3108 VDDA.n2984 1.70583
R4578 VDDA.n3110 VDDA.n2984 1.70583
R4579 VDDA.n3112 VDDA.n2984 1.70583
R4580 VDDA.n3114 VDDA.n2984 1.70583
R4581 VDDA.n3116 VDDA.n2984 1.70583
R4582 VDDA.n3118 VDDA.n2984 1.70583
R4583 VDDA.n3120 VDDA.n2984 1.70583
R4584 VDDA.n3122 VDDA.n2984 1.70583
R4585 VDDA.n3124 VDDA.n2984 1.70583
R4586 VDDA.n3126 VDDA.n2984 1.70583
R4587 VDDA.n3128 VDDA.n2984 1.70583
R4588 VDDA.n3130 VDDA.n2984 1.70583
R4589 VDDA.n3085 VDDA.n2984 1.70583
R4590 VDDA.n3132 VDDA.n3101 1.70583
R4591 VDDA.n2982 VDDA.n0 1.70567
R4592 VDDA.n2983 VDDA.n17 1.70567
R4593 VDDA.n2985 VDDA.n2982 1.70567
R4594 VDDA.n2986 VDDA.n17 1.70567
R4595 VDDA.n2988 VDDA.n2982 1.70567
R4596 VDDA.n2989 VDDA.n17 1.70567
R4597 VDDA.n2991 VDDA.n2982 1.70567
R4598 VDDA.n2992 VDDA.n17 1.70567
R4599 VDDA.n2994 VDDA.n2982 1.70567
R4600 VDDA.n2995 VDDA.n17 1.70567
R4601 VDDA.n2997 VDDA.n2982 1.70567
R4602 VDDA.n2998 VDDA.n17 1.70567
R4603 VDDA.n3000 VDDA.n2982 1.70567
R4604 VDDA.n3001 VDDA.n17 1.70567
R4605 VDDA.n3003 VDDA.n2982 1.70567
R4606 VDDA.n3004 VDDA.n17 1.70567
R4607 VDDA.n3006 VDDA.n2982 1.70567
R4608 VDDA.n3007 VDDA.n17 1.70567
R4609 VDDA.n3009 VDDA.n2982 1.70567
R4610 VDDA.n3010 VDDA.n17 1.70567
R4611 VDDA.n3012 VDDA.n2982 1.70567
R4612 VDDA.n3013 VDDA.n17 1.70567
R4613 VDDA.n3015 VDDA.n2982 1.70567
R4614 VDDA.n3016 VDDA.n17 1.70567
R4615 VDDA.n3018 VDDA.n2982 1.70567
R4616 VDDA.n3019 VDDA.n17 1.70567
R4617 VDDA.n3021 VDDA.n2982 1.70567
R4618 VDDA.n3022 VDDA.n17 1.70567
R4619 VDDA.n3024 VDDA.n2982 1.70567
R4620 VDDA.n3025 VDDA.n17 1.70567
R4621 VDDA.n3027 VDDA.n2982 1.70567
R4622 VDDA.n3028 VDDA.n17 1.70567
R4623 VDDA.n3030 VDDA.n2982 1.70567
R4624 VDDA.n3031 VDDA.n17 1.70567
R4625 VDDA.n3034 VDDA.n17 1.70567
R4626 VDDA.n3036 VDDA.n2982 1.70567
R4627 VDDA.n3037 VDDA.n17 1.70567
R4628 VDDA.n3039 VDDA.n2982 1.70567
R4629 VDDA.n3040 VDDA.n17 1.70567
R4630 VDDA.n3042 VDDA.n2982 1.70567
R4631 VDDA.n3043 VDDA.n17 1.70567
R4632 VDDA.n3045 VDDA.n2982 1.70567
R4633 VDDA.n3046 VDDA.n17 1.70567
R4634 VDDA.n3048 VDDA.n2982 1.70567
R4635 VDDA.n3049 VDDA.n17 1.70567
R4636 VDDA.n3051 VDDA.n2982 1.70567
R4637 VDDA.n3052 VDDA.n17 1.70567
R4638 VDDA.n3054 VDDA.n2982 1.70567
R4639 VDDA.n3055 VDDA.n17 1.70567
R4640 VDDA.n3057 VDDA.n2982 1.70567
R4641 VDDA.n3058 VDDA.n17 1.70567
R4642 VDDA.n3060 VDDA.n2982 1.70567
R4643 VDDA.n3061 VDDA.n17 1.70567
R4644 VDDA.n3063 VDDA.n2982 1.70567
R4645 VDDA.n3064 VDDA.n17 1.70567
R4646 VDDA.n3066 VDDA.n2982 1.70567
R4647 VDDA.n3067 VDDA.n17 1.70567
R4648 VDDA.n3069 VDDA.n2982 1.70567
R4649 VDDA.n3070 VDDA.n17 1.70567
R4650 VDDA.n3072 VDDA.n2982 1.70567
R4651 VDDA.n3073 VDDA.n17 1.70567
R4652 VDDA.n3075 VDDA.n2982 1.70567
R4653 VDDA.n3076 VDDA.n17 1.70567
R4654 VDDA.n3078 VDDA.n2982 1.70567
R4655 VDDA.n3079 VDDA.n17 1.70567
R4656 VDDA.n3081 VDDA.n2982 1.70567
R4657 VDDA.n3082 VDDA.n17 1.70567
R4658 VDDA.n3084 VDDA.n2982 1.70567
R4659 VDDA.n1651 VDDA.n1650 1.7055
R4660 VDDA.n1647 VDDA.n1645 1.7055
R4661 VDDA.n1656 VDDA.n1655 1.7055
R4662 VDDA.n1658 VDDA.n1641 1.7055
R4663 VDDA.n1661 VDDA.n1660 1.7055
R4664 VDDA.n1642 VDDA.n1639 1.7055
R4665 VDDA.n1666 VDDA.n1665 1.7055
R4666 VDDA.n1668 VDDA.n1635 1.7055
R4667 VDDA.n1671 VDDA.n1670 1.7055
R4668 VDDA.n1636 VDDA.n1633 1.7055
R4669 VDDA.n1676 VDDA.n1675 1.7055
R4670 VDDA.n1678 VDDA.n1629 1.7055
R4671 VDDA.n1681 VDDA.n1680 1.7055
R4672 VDDA.n1630 VDDA.n1627 1.7055
R4673 VDDA.n1686 VDDA.n1685 1.7055
R4674 VDDA.n1688 VDDA.n1623 1.7055
R4675 VDDA.n1691 VDDA.n1690 1.7055
R4676 VDDA.n1624 VDDA.n1621 1.7055
R4677 VDDA.n1696 VDDA.n1695 1.7055
R4678 VDDA.n1698 VDDA.n1617 1.7055
R4679 VDDA.n1701 VDDA.n1700 1.7055
R4680 VDDA.n1618 VDDA.n1615 1.7055
R4681 VDDA.n1706 VDDA.n1705 1.7055
R4682 VDDA.n1708 VDDA.n1611 1.7055
R4683 VDDA.n1711 VDDA.n1710 1.7055
R4684 VDDA.n1612 VDDA.n1609 1.7055
R4685 VDDA.n1716 VDDA.n1715 1.7055
R4686 VDDA.n1718 VDDA.n1605 1.7055
R4687 VDDA.n1721 VDDA.n1720 1.7055
R4688 VDDA.n1606 VDDA.n1603 1.7055
R4689 VDDA.n1726 VDDA.n1725 1.7055
R4690 VDDA.n1728 VDDA.n1599 1.7055
R4691 VDDA.n1731 VDDA.n1730 1.7055
R4692 VDDA.n1600 VDDA.n1597 1.7055
R4693 VDDA.n1736 VDDA.n1735 1.7055
R4694 VDDA.n1738 VDDA.n1593 1.7055
R4695 VDDA.n1741 VDDA.n1740 1.7055
R4696 VDDA.n1594 VDDA.n1591 1.7055
R4697 VDDA.n1746 VDDA.n1745 1.7055
R4698 VDDA.n1748 VDDA.n1587 1.7055
R4699 VDDA.n1751 VDDA.n1750 1.7055
R4700 VDDA.n1588 VDDA.n1584 1.7055
R4701 VDDA.n1756 VDDA.n1755 1.7055
R4702 VDDA.n1758 VDDA.n1582 1.7055
R4703 VDDA.n1760 VDDA.n1407 1.7055
R4704 VDDA.n1763 VDDA.n1762 1.7055
R4705 VDDA.n1409 VDDA.n1405 1.7055
R4706 VDDA.n3033 VDDA.n2982 1.70549
R4707 VDDA.n1643 VDDA.n1581 1.69989
R4708 VDDA.n1677 VDDA.n1581 1.69989
R4709 VDDA.n1625 VDDA.n1581 1.69989
R4710 VDDA.n1707 VDDA.n1581 1.69989
R4711 VDDA.n1607 VDDA.n1581 1.69989
R4712 VDDA.n1737 VDDA.n1581 1.69989
R4713 VDDA.n1589 VDDA.n1581 1.69989
R4714 VDDA.n1659 VDDA.n1368 1.69938
R4715 VDDA.n1638 VDDA.n1368 1.69938
R4716 VDDA.n1632 VDDA.n1368 1.69938
R4717 VDDA.n1679 VDDA.n1368 1.69938
R4718 VDDA.n1689 VDDA.n1368 1.69938
R4719 VDDA.n1620 VDDA.n1368 1.69938
R4720 VDDA.n1614 VDDA.n1368 1.69938
R4721 VDDA.n1709 VDDA.n1368 1.69938
R4722 VDDA.n1719 VDDA.n1368 1.69938
R4723 VDDA.n1602 VDDA.n1368 1.69938
R4724 VDDA.n1596 VDDA.n1368 1.69938
R4725 VDDA.n1739 VDDA.n1368 1.69938
R4726 VDDA.n1749 VDDA.n1368 1.69938
R4727 VDDA.n1583 VDDA.n1368 1.69938
R4728 VDDA.n1408 VDDA.n1368 1.69938
R4729 VDDA.n1649 VDDA.n1368 1.69938
R4730 VDDA.n1648 VDDA.n1581 1.69888
R4731 VDDA.n1644 VDDA.n1368 1.69888
R4732 VDDA.n1657 VDDA.n1581 1.69888
R4733 VDDA.n1667 VDDA.n1581 1.69888
R4734 VDDA.n1669 VDDA.n1368 1.69888
R4735 VDDA.n1637 VDDA.n1581 1.69888
R4736 VDDA.n1631 VDDA.n1581 1.69888
R4737 VDDA.n1626 VDDA.n1368 1.69888
R4738 VDDA.n1687 VDDA.n1581 1.69888
R4739 VDDA.n1697 VDDA.n1581 1.69888
R4740 VDDA.n1699 VDDA.n1368 1.69888
R4741 VDDA.n1619 VDDA.n1581 1.69888
R4742 VDDA.n1613 VDDA.n1581 1.69888
R4743 VDDA.n1608 VDDA.n1368 1.69888
R4744 VDDA.n1717 VDDA.n1581 1.69888
R4745 VDDA.n1727 VDDA.n1581 1.69888
R4746 VDDA.n1729 VDDA.n1368 1.69888
R4747 VDDA.n1601 VDDA.n1581 1.69888
R4748 VDDA.n1595 VDDA.n1581 1.69888
R4749 VDDA.n1590 VDDA.n1368 1.69888
R4750 VDDA.n1747 VDDA.n1581 1.69888
R4751 VDDA.n1757 VDDA.n1581 1.69888
R4752 VDDA.n1759 VDDA.n1368 1.69888
R4753 VDDA.n1761 VDDA.n1581 1.69888
R4754 VDDA.n813 VDDA.n662 1.69433
R4755 VDDA.n813 VDDA.n659 1.69433
R4756 VDDA.n813 VDDA.n656 1.69433
R4757 VDDA.n813 VDDA.n653 1.69433
R4758 VDDA.n813 VDDA.n650 1.69433
R4759 VDDA.n813 VDDA.n647 1.69433
R4760 VDDA.n813 VDDA.n644 1.69433
R4761 VDDA.n973 VDDA.n835 1.69433
R4762 VDDA.n973 VDDA.n832 1.69433
R4763 VDDA.n973 VDDA.n829 1.69433
R4764 VDDA.n973 VDDA.n826 1.69433
R4765 VDDA.n973 VDDA.n823 1.69433
R4766 VDDA.n973 VDDA.n820 1.69433
R4767 VDDA.n973 VDDA.n817 1.69433
R4768 VDDA.n1133 VDDA.n464 1.69433
R4769 VDDA.n1115 VDDA.n464 1.69433
R4770 VDDA.n1103 VDDA.n464 1.69433
R4771 VDDA.n1085 VDDA.n464 1.69433
R4772 VDDA.n1073 VDDA.n464 1.69433
R4773 VDDA.n1055 VDDA.n464 1.69433
R4774 VDDA.n1043 VDDA.n464 1.69433
R4775 VDDA.n1161 VDDA.n486 1.69433
R4776 VDDA.n1161 VDDA.n483 1.69433
R4777 VDDA.n1161 VDDA.n480 1.69433
R4778 VDDA.n1161 VDDA.n477 1.69433
R4779 VDDA.n1161 VDDA.n474 1.69433
R4780 VDDA.n1161 VDDA.n471 1.69433
R4781 VDDA.n1161 VDDA.n468 1.69433
R4782 VDDA.n2258 VDDA.n1183 1.69433
R4783 VDDA.n2258 VDDA.n1180 1.69433
R4784 VDDA.n2258 VDDA.n1177 1.69433
R4785 VDDA.n2258 VDDA.n1174 1.69433
R4786 VDDA.n2258 VDDA.n1171 1.69433
R4787 VDDA.n2258 VDDA.n1168 1.69433
R4788 VDDA.n2258 VDDA.n1165 1.69433
R4789 VDDA.n2257 VDDA.n1341 1.69433
R4790 VDDA.n2257 VDDA.n1338 1.69433
R4791 VDDA.n2257 VDDA.n1335 1.69433
R4792 VDDA.n2257 VDDA.n1332 1.69433
R4793 VDDA.n2257 VDDA.n1329 1.69433
R4794 VDDA.n2257 VDDA.n1326 1.69433
R4795 VDDA.n2257 VDDA.n1323 1.69433
R4796 VDDA.n2571 VDDA.n197 1.69433
R4797 VDDA.n2553 VDDA.n197 1.69433
R4798 VDDA.n2541 VDDA.n197 1.69433
R4799 VDDA.n2523 VDDA.n197 1.69433
R4800 VDDA.n2511 VDDA.n197 1.69433
R4801 VDDA.n2493 VDDA.n197 1.69433
R4802 VDDA.n2481 VDDA.n197 1.69433
R4803 VDDA.n2599 VDDA.n219 1.69433
R4804 VDDA.n2599 VDDA.n216 1.69433
R4805 VDDA.n2599 VDDA.n213 1.69433
R4806 VDDA.n2599 VDDA.n210 1.69433
R4807 VDDA.n2599 VDDA.n207 1.69433
R4808 VDDA.n2599 VDDA.n204 1.69433
R4809 VDDA.n2599 VDDA.n201 1.69433
R4810 VDDA.n2759 VDDA.n2621 1.69433
R4811 VDDA.n2759 VDDA.n2618 1.69433
R4812 VDDA.n2759 VDDA.n2615 1.69433
R4813 VDDA.n2759 VDDA.n2612 1.69433
R4814 VDDA.n2759 VDDA.n2609 1.69433
R4815 VDDA.n2759 VDDA.n2606 1.69433
R4816 VDDA.n2759 VDDA.n2603 1.69433
R4817 VDDA.n2919 VDDA.n19 1.69433
R4818 VDDA.n2901 VDDA.n19 1.69433
R4819 VDDA.n2889 VDDA.n19 1.69433
R4820 VDDA.n2871 VDDA.n19 1.69433
R4821 VDDA.n2859 VDDA.n19 1.69433
R4822 VDDA.n2841 VDDA.n19 1.69433
R4823 VDDA.n2829 VDDA.n19 1.69433
R4824 VDDA.n2947 VDDA.n41 1.69433
R4825 VDDA.n2947 VDDA.n38 1.69433
R4826 VDDA.n2947 VDDA.n35 1.69433
R4827 VDDA.n2947 VDDA.n32 1.69433
R4828 VDDA.n2947 VDDA.n29 1.69433
R4829 VDDA.n2947 VDDA.n26 1.69433
R4830 VDDA.n2947 VDDA.n23 1.69433
R4831 VDDA.n1580 VDDA.n1431 1.69433
R4832 VDDA.n1580 VDDA.n1428 1.69433
R4833 VDDA.n1580 VDDA.n1425 1.69433
R4834 VDDA.n1580 VDDA.n1422 1.69433
R4835 VDDA.n1580 VDDA.n1419 1.69433
R4836 VDDA.n1580 VDDA.n1416 1.69433
R4837 VDDA.n1580 VDDA.n1413 1.69433
R4838 VDDA.n1908 VDDA.n1365 1.69328
R4839 VDDA.n1908 VDDA.n1362 1.69328
R4840 VDDA.n1908 VDDA.n1359 1.69328
R4841 VDDA.n1908 VDDA.n1356 1.69328
R4842 VDDA.n1908 VDDA.n1353 1.69328
R4843 VDDA.n1908 VDDA.n1350 1.69328
R4844 VDDA.n1908 VDDA.n1347 1.69328
R4845 VDDA.n813 VDDA.n664 1.6924
R4846 VDDA.n813 VDDA.n663 1.6924
R4847 VDDA.n813 VDDA.n661 1.6924
R4848 VDDA.n813 VDDA.n660 1.6924
R4849 VDDA.n813 VDDA.n658 1.6924
R4850 VDDA.n813 VDDA.n657 1.6924
R4851 VDDA.n813 VDDA.n655 1.6924
R4852 VDDA.n813 VDDA.n654 1.6924
R4853 VDDA.n813 VDDA.n652 1.6924
R4854 VDDA.n813 VDDA.n651 1.6924
R4855 VDDA.n813 VDDA.n649 1.6924
R4856 VDDA.n813 VDDA.n648 1.6924
R4857 VDDA.n813 VDDA.n646 1.6924
R4858 VDDA.n813 VDDA.n645 1.6924
R4859 VDDA.n813 VDDA.n643 1.6924
R4860 VDDA.n813 VDDA.n642 1.6924
R4861 VDDA.n973 VDDA.n972 1.6924
R4862 VDDA.n973 VDDA.n836 1.6924
R4863 VDDA.n973 VDDA.n834 1.6924
R4864 VDDA.n973 VDDA.n833 1.6924
R4865 VDDA.n973 VDDA.n831 1.6924
R4866 VDDA.n973 VDDA.n830 1.6924
R4867 VDDA.n973 VDDA.n828 1.6924
R4868 VDDA.n973 VDDA.n827 1.6924
R4869 VDDA.n973 VDDA.n825 1.6924
R4870 VDDA.n973 VDDA.n824 1.6924
R4871 VDDA.n973 VDDA.n822 1.6924
R4872 VDDA.n973 VDDA.n821 1.6924
R4873 VDDA.n973 VDDA.n819 1.6924
R4874 VDDA.n973 VDDA.n818 1.6924
R4875 VDDA.n973 VDDA.n816 1.6924
R4876 VDDA.n973 VDDA.n815 1.6924
R4877 VDDA.n1143 VDDA.n464 1.6924
R4878 VDDA.n1135 VDDA.n464 1.6924
R4879 VDDA.n1125 VDDA.n464 1.6924
R4880 VDDA.n1123 VDDA.n464 1.6924
R4881 VDDA.n1113 VDDA.n464 1.6924
R4882 VDDA.n1105 VDDA.n464 1.6924
R4883 VDDA.n1095 VDDA.n464 1.6924
R4884 VDDA.n1093 VDDA.n464 1.6924
R4885 VDDA.n1083 VDDA.n464 1.6924
R4886 VDDA.n1075 VDDA.n464 1.6924
R4887 VDDA.n1065 VDDA.n464 1.6924
R4888 VDDA.n1063 VDDA.n464 1.6924
R4889 VDDA.n1053 VDDA.n464 1.6924
R4890 VDDA.n1045 VDDA.n464 1.6924
R4891 VDDA.n1035 VDDA.n464 1.6924
R4892 VDDA.n1033 VDDA.n464 1.6924
R4893 VDDA.n1161 VDDA.n488 1.6924
R4894 VDDA.n1161 VDDA.n487 1.6924
R4895 VDDA.n1161 VDDA.n485 1.6924
R4896 VDDA.n1161 VDDA.n484 1.6924
R4897 VDDA.n1161 VDDA.n482 1.6924
R4898 VDDA.n1161 VDDA.n481 1.6924
R4899 VDDA.n1161 VDDA.n479 1.6924
R4900 VDDA.n1161 VDDA.n478 1.6924
R4901 VDDA.n1161 VDDA.n476 1.6924
R4902 VDDA.n1161 VDDA.n475 1.6924
R4903 VDDA.n1161 VDDA.n473 1.6924
R4904 VDDA.n1161 VDDA.n472 1.6924
R4905 VDDA.n1161 VDDA.n470 1.6924
R4906 VDDA.n1161 VDDA.n469 1.6924
R4907 VDDA.n1161 VDDA.n467 1.6924
R4908 VDDA.n1161 VDDA.n466 1.6924
R4909 VDDA.n2258 VDDA.n1320 1.6924
R4910 VDDA.n2258 VDDA.n1184 1.6924
R4911 VDDA.n2258 VDDA.n1182 1.6924
R4912 VDDA.n2258 VDDA.n1181 1.6924
R4913 VDDA.n2258 VDDA.n1179 1.6924
R4914 VDDA.n2258 VDDA.n1178 1.6924
R4915 VDDA.n2258 VDDA.n1176 1.6924
R4916 VDDA.n2258 VDDA.n1175 1.6924
R4917 VDDA.n2258 VDDA.n1173 1.6924
R4918 VDDA.n2258 VDDA.n1172 1.6924
R4919 VDDA.n2258 VDDA.n1170 1.6924
R4920 VDDA.n2258 VDDA.n1169 1.6924
R4921 VDDA.n2258 VDDA.n1167 1.6924
R4922 VDDA.n2258 VDDA.n1166 1.6924
R4923 VDDA.n2258 VDDA.n1164 1.6924
R4924 VDDA.n2258 VDDA.n1163 1.6924
R4925 VDDA.n2257 VDDA.n1343 1.6924
R4926 VDDA.n2257 VDDA.n1342 1.6924
R4927 VDDA.n2257 VDDA.n1340 1.6924
R4928 VDDA.n2257 VDDA.n1339 1.6924
R4929 VDDA.n2257 VDDA.n1337 1.6924
R4930 VDDA.n2257 VDDA.n1336 1.6924
R4931 VDDA.n2257 VDDA.n1334 1.6924
R4932 VDDA.n2257 VDDA.n1333 1.6924
R4933 VDDA.n2257 VDDA.n1331 1.6924
R4934 VDDA.n2257 VDDA.n1330 1.6924
R4935 VDDA.n2257 VDDA.n1328 1.6924
R4936 VDDA.n2257 VDDA.n1327 1.6924
R4937 VDDA.n2257 VDDA.n1325 1.6924
R4938 VDDA.n2257 VDDA.n1324 1.6924
R4939 VDDA.n2257 VDDA.n1322 1.6924
R4940 VDDA.n2581 VDDA.n197 1.6924
R4941 VDDA.n2573 VDDA.n197 1.6924
R4942 VDDA.n2563 VDDA.n197 1.6924
R4943 VDDA.n2561 VDDA.n197 1.6924
R4944 VDDA.n2551 VDDA.n197 1.6924
R4945 VDDA.n2543 VDDA.n197 1.6924
R4946 VDDA.n2533 VDDA.n197 1.6924
R4947 VDDA.n2531 VDDA.n197 1.6924
R4948 VDDA.n2521 VDDA.n197 1.6924
R4949 VDDA.n2513 VDDA.n197 1.6924
R4950 VDDA.n2503 VDDA.n197 1.6924
R4951 VDDA.n2501 VDDA.n197 1.6924
R4952 VDDA.n2491 VDDA.n197 1.6924
R4953 VDDA.n2483 VDDA.n197 1.6924
R4954 VDDA.n2473 VDDA.n197 1.6924
R4955 VDDA.n2471 VDDA.n197 1.6924
R4956 VDDA.n2599 VDDA.n221 1.6924
R4957 VDDA.n2599 VDDA.n220 1.6924
R4958 VDDA.n2599 VDDA.n218 1.6924
R4959 VDDA.n2599 VDDA.n217 1.6924
R4960 VDDA.n2599 VDDA.n215 1.6924
R4961 VDDA.n2599 VDDA.n214 1.6924
R4962 VDDA.n2599 VDDA.n212 1.6924
R4963 VDDA.n2599 VDDA.n211 1.6924
R4964 VDDA.n2599 VDDA.n209 1.6924
R4965 VDDA.n2599 VDDA.n208 1.6924
R4966 VDDA.n2599 VDDA.n206 1.6924
R4967 VDDA.n2599 VDDA.n205 1.6924
R4968 VDDA.n2599 VDDA.n203 1.6924
R4969 VDDA.n2599 VDDA.n202 1.6924
R4970 VDDA.n2599 VDDA.n200 1.6924
R4971 VDDA.n2599 VDDA.n199 1.6924
R4972 VDDA.n2759 VDDA.n2758 1.6924
R4973 VDDA.n2759 VDDA.n2622 1.6924
R4974 VDDA.n2759 VDDA.n2620 1.6924
R4975 VDDA.n2759 VDDA.n2619 1.6924
R4976 VDDA.n2759 VDDA.n2617 1.6924
R4977 VDDA.n2759 VDDA.n2616 1.6924
R4978 VDDA.n2759 VDDA.n2614 1.6924
R4979 VDDA.n2759 VDDA.n2613 1.6924
R4980 VDDA.n2759 VDDA.n2611 1.6924
R4981 VDDA.n2759 VDDA.n2610 1.6924
R4982 VDDA.n2759 VDDA.n2608 1.6924
R4983 VDDA.n2759 VDDA.n2607 1.6924
R4984 VDDA.n2759 VDDA.n2605 1.6924
R4985 VDDA.n2759 VDDA.n2604 1.6924
R4986 VDDA.n2759 VDDA.n2602 1.6924
R4987 VDDA.n2759 VDDA.n2601 1.6924
R4988 VDDA.n2929 VDDA.n19 1.6924
R4989 VDDA.n2921 VDDA.n19 1.6924
R4990 VDDA.n2911 VDDA.n19 1.6924
R4991 VDDA.n2909 VDDA.n19 1.6924
R4992 VDDA.n2899 VDDA.n19 1.6924
R4993 VDDA.n2891 VDDA.n19 1.6924
R4994 VDDA.n2881 VDDA.n19 1.6924
R4995 VDDA.n2879 VDDA.n19 1.6924
R4996 VDDA.n2869 VDDA.n19 1.6924
R4997 VDDA.n2861 VDDA.n19 1.6924
R4998 VDDA.n2851 VDDA.n19 1.6924
R4999 VDDA.n2849 VDDA.n19 1.6924
R5000 VDDA.n2839 VDDA.n19 1.6924
R5001 VDDA.n2831 VDDA.n19 1.6924
R5002 VDDA.n2821 VDDA.n19 1.6924
R5003 VDDA.n2819 VDDA.n19 1.6924
R5004 VDDA.n2947 VDDA.n43 1.6924
R5005 VDDA.n2947 VDDA.n42 1.6924
R5006 VDDA.n2947 VDDA.n40 1.6924
R5007 VDDA.n2947 VDDA.n39 1.6924
R5008 VDDA.n2947 VDDA.n37 1.6924
R5009 VDDA.n2947 VDDA.n36 1.6924
R5010 VDDA.n2947 VDDA.n34 1.6924
R5011 VDDA.n2947 VDDA.n33 1.6924
R5012 VDDA.n2947 VDDA.n31 1.6924
R5013 VDDA.n2947 VDDA.n30 1.6924
R5014 VDDA.n2947 VDDA.n28 1.6924
R5015 VDDA.n2947 VDDA.n27 1.6924
R5016 VDDA.n2947 VDDA.n25 1.6924
R5017 VDDA.n2947 VDDA.n24 1.6924
R5018 VDDA.n2947 VDDA.n22 1.6924
R5019 VDDA.n2947 VDDA.n21 1.6924
R5020 VDDA.n1580 VDDA.n1433 1.6924
R5021 VDDA.n1580 VDDA.n1432 1.6924
R5022 VDDA.n1580 VDDA.n1430 1.6924
R5023 VDDA.n1580 VDDA.n1429 1.6924
R5024 VDDA.n1580 VDDA.n1427 1.6924
R5025 VDDA.n1580 VDDA.n1426 1.6924
R5026 VDDA.n1580 VDDA.n1424 1.6924
R5027 VDDA.n1580 VDDA.n1423 1.6924
R5028 VDDA.n1580 VDDA.n1421 1.6924
R5029 VDDA.n1580 VDDA.n1420 1.6924
R5030 VDDA.n1580 VDDA.n1418 1.6924
R5031 VDDA.n1580 VDDA.n1417 1.6924
R5032 VDDA.n1580 VDDA.n1415 1.6924
R5033 VDDA.n1580 VDDA.n1414 1.6924
R5034 VDDA.n1580 VDDA.n1412 1.6924
R5035 VDDA.n1580 VDDA.n1411 1.6924
R5036 VDDA.n1908 VDDA.n1367 1.69118
R5037 VDDA.n1908 VDDA.n1366 1.69118
R5038 VDDA.n1908 VDDA.n1364 1.69118
R5039 VDDA.n1908 VDDA.n1363 1.69118
R5040 VDDA.n1908 VDDA.n1361 1.69118
R5041 VDDA.n1908 VDDA.n1360 1.69118
R5042 VDDA.n1908 VDDA.n1358 1.69118
R5043 VDDA.n1908 VDDA.n1357 1.69118
R5044 VDDA.n1908 VDDA.n1355 1.69118
R5045 VDDA.n1908 VDDA.n1354 1.69118
R5046 VDDA.n1908 VDDA.n1352 1.69118
R5047 VDDA.n1908 VDDA.n1351 1.69118
R5048 VDDA.n1908 VDDA.n1349 1.69118
R5049 VDDA.n1908 VDDA.n1348 1.69118
R5050 VDDA.n1908 VDDA.n1346 1.69118
R5051 VDDA.n1908 VDDA.n1345 1.69118
R5052 VDDA.n373 VDDA.n372 1.63212
R5053 VDDA.n380 VDDA.n378 1.63212
R5054 VDDA.n385 VDDA.n377 1.59823
R5055 VDDA.n377 VDDA.n376 1.56962
R5056 VDDA.n384 VDDA.n383 1.56962
R5057 VDDA.n1790 VDDA.n1393 1.56177
R5058 VDDA.n1767 VDDA.n1393 1.50969
R5059 VDDA.n2279 VDDA.n2278 1.46464
R5060 VDDA.n2281 VDDA.n2280 1.46464
R5061 VDDA.n1404 VDDA.n1393 1.44719
R5062 VDDA.n452 VDDA.n386 1.31821
R5063 VDDA.n2401 VDDA.n386 1.31821
R5064 VDDA.n1944 VDDA.n1943 1.26222
R5065 VDDA.n1653 VDDA.n1652 1.20209
R5066 VDDA.n2395 VDDA.n439 1.13592
R5067 VDDA.n2339 VDDA.n2338 1.13592
R5068 VDDA.n2257 VDDA.n1321 1.12311
R5069 VDDA.n430 VDDA.n428 1.07342
R5070 VDDA.n2335 VDDA.n2327 1.06821
R5071 VDDA.n1950 VDDA.n1949 0.943208
R5072 VDDA.n2361 VDDA.n2345 0.932792
R5073 VDDA.n2394 VDDA.n2393 0.932792
R5074 VDDA.n2399 VDDA.n2398 0.922375
R5075 VDDA.n2343 VDDA.n2289 0.922375
R5076 VDDA.n2087 VDDA.n2086 0.880708
R5077 VDDA.n2010 VDDA.n2009 0.865083
R5078 VDDA.n2137 VDDA.n2136 0.807792
R5079 VDDA.n1942 VDDA.n1941 0.75233
R5080 VDDA.n2016 VDDA.n2015 0.672375
R5081 VDDA.n1943 VDDA.n1942 0.648711
R5082 VDDA.n2264 VDDA.n459 0.646333
R5083 VDDA.n2592 VDDA.n2590 0.646333
R5084 VDDA.n2410 VDDA.n2408 0.6255
R5085 VDDA.n2413 VDDA.n2410 0.6255
R5086 VDDA.n2415 VDDA.n2413 0.6255
R5087 VDDA.n2417 VDDA.n2415 0.6255
R5088 VDDA.n2272 VDDA.n2269 0.6255
R5089 VDDA.n2269 VDDA.n455 0.6255
R5090 VDDA.n2276 VDDA.n2274 0.6255
R5091 VDDA.n2274 VDDA.n2272 0.6255
R5092 VDDA.n3133 VDDA.n2947 0.546104
R5093 VDDA.n2267 VDDA.n2266 0.490083
R5094 VDDA.n2588 VDDA.n2419 0.490083
R5095 VDDA.n2144 VDDA.n2142 0.448417
R5096 VDDA.n2282 VDDA.n2281 0.424316
R5097 VDDA.n2278 VDDA.n2277 0.424316
R5098 VDDA.n2267 VDDA.n453 0.3755
R5099 VDDA.n2283 VDDA.n453 0.3755
R5100 VDDA.n2404 VDDA.n366 0.3755
R5101 VDDA.n2419 VDDA.n366 0.3755
R5102 VDDA.n2000 VDDA.n1999 0.333833
R5103 VDDA.n2081 VDDA.n2080 0.328625
R5104 VDDA.n2323 VDDA.n2322 0.323417
R5105 VDDA.n426 VDDA.n425 0.323417
R5106 VDDA.n2134 VDDA.n2133 0.292167
R5107 VDDA.n2130 VDDA.n2129 0.292167
R5108 VDDA.n2123 VDDA.n2122 0.292167
R5109 VDDA.n2093 VDDA.n2092 0.292167
R5110 VDDA.n979 VDDA.n636 0.28175
R5111 VDDA.n1150 VDDA.n981 0.28175
R5112 VDDA.n1154 VDDA.n1152 0.28175
R5113 VDDA.n2765 VDDA.n192 0.28175
R5114 VDDA.n2936 VDDA.n2767 0.28175
R5115 VDDA.n2939 VDDA.n2938 0.28175
R5116 VDDA.n2333 VDDA.n2332 0.266125
R5117 VDDA.n437 VDDA.n436 0.266125
R5118 VDDA.n2341 VDDA.n2305 0.266125
R5119 VDDA.n2396 VDDA.n405 0.266125
R5120 VDDA.n1998 VDDA.n1997 0.2505
R5121 VDDA.n2008 VDDA.n2007 0.2505
R5122 VDDA.n2288 VDDA.n2283 0.234875
R5123 VDDA.n2404 VDDA.n2403 0.234875
R5124 VDDA.n1769 VDDA.n1768 0.229667
R5125 VDDA.n1789 VDDA.n1788 0.229667
R5126 VDDA.n2086 VDDA.n2081 0.229667
R5127 VDDA.n1770 VDDA.n1400 0.208833
R5128 VDDA.n1770 VDDA.n1769 0.208833
R5129 VDDA.n1782 VDDA.n1394 0.208833
R5130 VDDA.n1788 VDDA.n1394 0.208833
R5131 VDDA.n2048 VDDA.n2034 0.208833
R5132 VDDA.n2042 VDDA.n2034 0.208833
R5133 VDDA.n2042 VDDA.n2041 0.208833
R5134 VDDA.n2057 VDDA.n2055 0.208833
R5135 VDDA.n2058 VDDA.n2057 0.208833
R5136 VDDA.n2058 VDDA.n2027 0.208833
R5137 VDDA.n2080 VDDA.n2079 0.188
R5138 VDDA.n2079 VDDA.n2078 0.188
R5139 VDDA.n2078 VDDA.n2077 0.188
R5140 VDDA.n2077 VDDA.n2076 0.188
R5141 VDDA.n2076 VDDA.n2075 0.188
R5142 VDDA.n2075 VDDA.n2074 0.188
R5143 VDDA.n2074 VDDA.n2073 0.188
R5144 VDDA.n2073 VDDA.n2072 0.188
R5145 VDDA.n2363 VDDA.n2361 0.172375
R5146 VDDA.n2364 VDDA.n2363 0.172375
R5147 VDDA.n2365 VDDA.n441 0.172375
R5148 VDDA.n2393 VDDA.n441 0.172375
R5149 VDDA.t52 VDDA.t181 0.1603
R5150 VDDA.t392 VDDA.t395 0.1603
R5151 VDDA.t137 VDDA.t55 0.1603
R5152 VDDA.t68 VDDA.t98 0.1603
R5153 VDDA.t174 VDDA.t139 0.1603
R5154 VDDA.n1796 VDDA.n1795 0.159591
R5155 VDDA.n1797 VDDA.n1796 0.159591
R5156 VDDA.n1797 VDDA.n1391 0.159591
R5157 VDDA.n1807 VDDA.n1389 0.159591
R5158 VDDA.n1815 VDDA.n1389 0.159591
R5159 VDDA.n1816 VDDA.n1815 0.159591
R5160 VDDA.n1826 VDDA.n1825 0.159591
R5161 VDDA.n1827 VDDA.n1826 0.159591
R5162 VDDA.n1827 VDDA.n1385 0.159591
R5163 VDDA.n1837 VDDA.n1383 0.159591
R5164 VDDA.n1845 VDDA.n1383 0.159591
R5165 VDDA.n1846 VDDA.n1845 0.159591
R5166 VDDA.n1856 VDDA.n1855 0.159591
R5167 VDDA.n1857 VDDA.n1856 0.159591
R5168 VDDA.n1857 VDDA.n1379 0.159591
R5169 VDDA.n1867 VDDA.n1377 0.159591
R5170 VDDA.n1875 VDDA.n1377 0.159591
R5171 VDDA.n1876 VDDA.n1875 0.159591
R5172 VDDA.n1886 VDDA.n1885 0.159591
R5173 VDDA.n1887 VDDA.n1886 0.159591
R5174 VDDA.n1887 VDDA.n1373 0.159591
R5175 VDDA.n1897 VDDA.n1371 0.159591
R5176 VDDA.n1905 VDDA.n1371 0.159591
R5177 VDDA.n1794 VDDA.n1392 0.159591
R5178 VDDA.n1800 VDDA.n1392 0.159591
R5179 VDDA.n1801 VDDA.n1800 0.159591
R5180 VDDA.n1811 VDDA.n1810 0.159591
R5181 VDDA.n1814 VDDA.n1811 0.159591
R5182 VDDA.n1814 VDDA.n1388 0.159591
R5183 VDDA.n1824 VDDA.n1386 0.159591
R5184 VDDA.n1830 VDDA.n1386 0.159591
R5185 VDDA.n1831 VDDA.n1830 0.159591
R5186 VDDA.n1841 VDDA.n1840 0.159591
R5187 VDDA.n1844 VDDA.n1841 0.159591
R5188 VDDA.n1844 VDDA.n1382 0.159591
R5189 VDDA.n1854 VDDA.n1380 0.159591
R5190 VDDA.n1860 VDDA.n1380 0.159591
R5191 VDDA.n1861 VDDA.n1860 0.159591
R5192 VDDA.n1871 VDDA.n1870 0.159591
R5193 VDDA.n1874 VDDA.n1871 0.159591
R5194 VDDA.n1874 VDDA.n1376 0.159591
R5195 VDDA.n1884 VDDA.n1374 0.159591
R5196 VDDA.n1890 VDDA.n1374 0.159591
R5197 VDDA.n1891 VDDA.n1890 0.159591
R5198 VDDA.n1901 VDDA.n1900 0.159591
R5199 VDDA.n1904 VDDA.n1901 0.159591
R5200 VDDA.n1904 VDDA.n1370 0.159591
R5201 VDDA.n1459 VDDA.t59 0.159278
R5202 VDDA.n1460 VDDA.t138 0.159278
R5203 VDDA.n1461 VDDA.t393 0.159278
R5204 VDDA.n1462 VDDA.t163 0.159278
R5205 VDDA.n1795 VDDA.n1791 0.148227
R5206 VDDA.n1805 VDDA.n1391 0.148227
R5207 VDDA.n1807 VDDA.n1806 0.148227
R5208 VDDA.n1817 VDDA.n1816 0.148227
R5209 VDDA.n1825 VDDA.n1387 0.148227
R5210 VDDA.n1835 VDDA.n1385 0.148227
R5211 VDDA.n1837 VDDA.n1836 0.148227
R5212 VDDA.n1847 VDDA.n1846 0.148227
R5213 VDDA.n1855 VDDA.n1381 0.148227
R5214 VDDA.n1865 VDDA.n1379 0.148227
R5215 VDDA.n1867 VDDA.n1866 0.148227
R5216 VDDA.n1877 VDDA.n1876 0.148227
R5217 VDDA.n1885 VDDA.n1375 0.148227
R5218 VDDA.n1895 VDDA.n1373 0.148227
R5219 VDDA.n1897 VDDA.n1896 0.148227
R5220 VDDA.n1794 VDDA.n1792 0.148227
R5221 VDDA.n1804 VDDA.n1801 0.148227
R5222 VDDA.n1810 VDDA.n1390 0.148227
R5223 VDDA.n1820 VDDA.n1388 0.148227
R5224 VDDA.n1824 VDDA.n1821 0.148227
R5225 VDDA.n1834 VDDA.n1831 0.148227
R5226 VDDA.n1840 VDDA.n1384 0.148227
R5227 VDDA.n1850 VDDA.n1382 0.148227
R5228 VDDA.n1854 VDDA.n1851 0.148227
R5229 VDDA.n1864 VDDA.n1861 0.148227
R5230 VDDA.n1870 VDDA.n1378 0.148227
R5231 VDDA.n1880 VDDA.n1376 0.148227
R5232 VDDA.n1884 VDDA.n1881 0.148227
R5233 VDDA.n1894 VDDA.n1891 0.148227
R5234 VDDA.n1900 VDDA.n1372 0.148227
R5235 VDDA.n1466 VDDA.n1457 0.146333
R5236 VDDA.n1472 VDDA.n1457 0.146333
R5237 VDDA.n1473 VDDA.n1472 0.146333
R5238 VDDA.n1483 VDDA.n1482 0.146333
R5239 VDDA.n1486 VDDA.n1483 0.146333
R5240 VDDA.n1486 VDDA.n1453 0.146333
R5241 VDDA.n1496 VDDA.n1451 0.146333
R5242 VDDA.n1502 VDDA.n1451 0.146333
R5243 VDDA.n1503 VDDA.n1502 0.146333
R5244 VDDA.n1513 VDDA.n1512 0.146333
R5245 VDDA.n1516 VDDA.n1513 0.146333
R5246 VDDA.n1516 VDDA.n1447 0.146333
R5247 VDDA.n1526 VDDA.n1445 0.146333
R5248 VDDA.n1532 VDDA.n1445 0.146333
R5249 VDDA.n1533 VDDA.n1532 0.146333
R5250 VDDA.n1543 VDDA.n1542 0.146333
R5251 VDDA.n1546 VDDA.n1543 0.146333
R5252 VDDA.n1546 VDDA.n1441 0.146333
R5253 VDDA.n1556 VDDA.n1439 0.146333
R5254 VDDA.n1562 VDDA.n1439 0.146333
R5255 VDDA.n1563 VDDA.n1562 0.146333
R5256 VDDA.n1573 VDDA.n1572 0.146333
R5257 VDDA.n1576 VDDA.n1573 0.146333
R5258 VDDA.n1576 VDDA.n1435 0.146333
R5259 VDDA.n2143 VDDA.n1932 0.146333
R5260 VDDA.n2149 VDDA.n1932 0.146333
R5261 VDDA.n2150 VDDA.n2149 0.146333
R5262 VDDA.n2160 VDDA.n2159 0.146333
R5263 VDDA.n2163 VDDA.n2160 0.146333
R5264 VDDA.n2163 VDDA.n1928 0.146333
R5265 VDDA.n2173 VDDA.n1926 0.146333
R5266 VDDA.n2179 VDDA.n1926 0.146333
R5267 VDDA.n2180 VDDA.n2179 0.146333
R5268 VDDA.n2190 VDDA.n2189 0.146333
R5269 VDDA.n2193 VDDA.n2190 0.146333
R5270 VDDA.n2193 VDDA.n1922 0.146333
R5271 VDDA.n2203 VDDA.n1920 0.146333
R5272 VDDA.n2209 VDDA.n1920 0.146333
R5273 VDDA.n2210 VDDA.n2209 0.146333
R5274 VDDA.n2220 VDDA.n2219 0.146333
R5275 VDDA.n2223 VDDA.n2220 0.146333
R5276 VDDA.n2223 VDDA.n1916 0.146333
R5277 VDDA.n2233 VDDA.n1914 0.146333
R5278 VDDA.n2239 VDDA.n1914 0.146333
R5279 VDDA.n2240 VDDA.n2239 0.146333
R5280 VDDA.n2250 VDDA.n2249 0.146333
R5281 VDDA.n2253 VDDA.n2250 0.146333
R5282 VDDA.n2253 VDDA.n1910 0.146333
R5283 VDDA.n91 VDDA.n87 0.146333
R5284 VDDA.n95 VDDA.n87 0.146333
R5285 VDDA.n96 VDDA.n95 0.146333
R5286 VDDA.n104 VDDA.n103 0.146333
R5287 VDDA.n107 VDDA.n104 0.146333
R5288 VDDA.n107 VDDA.n79 0.146333
R5289 VDDA.n115 VDDA.n75 0.146333
R5290 VDDA.n119 VDDA.n75 0.146333
R5291 VDDA.n120 VDDA.n119 0.146333
R5292 VDDA.n128 VDDA.n127 0.146333
R5293 VDDA.n131 VDDA.n128 0.146333
R5294 VDDA.n131 VDDA.n67 0.146333
R5295 VDDA.n139 VDDA.n63 0.146333
R5296 VDDA.n143 VDDA.n63 0.146333
R5297 VDDA.n144 VDDA.n143 0.146333
R5298 VDDA.n152 VDDA.n151 0.146333
R5299 VDDA.n155 VDDA.n152 0.146333
R5300 VDDA.n155 VDDA.n55 0.146333
R5301 VDDA.n163 VDDA.n51 0.146333
R5302 VDDA.n167 VDDA.n51 0.146333
R5303 VDDA.n168 VDDA.n167 0.146333
R5304 VDDA.n176 VDDA.n175 0.146333
R5305 VDDA.n179 VDDA.n176 0.146333
R5306 VDDA.n179 VDDA.n45 0.146333
R5307 VDDA.n2817 VDDA.n2814 0.146333
R5308 VDDA.n2823 VDDA.n2814 0.146333
R5309 VDDA.n2823 VDDA.n2812 0.146333
R5310 VDDA.n2833 VDDA.n2808 0.146333
R5311 VDDA.n2837 VDDA.n2808 0.146333
R5312 VDDA.n2837 VDDA.n2806 0.146333
R5313 VDDA.n2847 VDDA.n2802 0.146333
R5314 VDDA.n2853 VDDA.n2802 0.146333
R5315 VDDA.n2853 VDDA.n2800 0.146333
R5316 VDDA.n2863 VDDA.n2796 0.146333
R5317 VDDA.n2867 VDDA.n2796 0.146333
R5318 VDDA.n2867 VDDA.n2794 0.146333
R5319 VDDA.n2877 VDDA.n2790 0.146333
R5320 VDDA.n2883 VDDA.n2790 0.146333
R5321 VDDA.n2883 VDDA.n2788 0.146333
R5322 VDDA.n2893 VDDA.n2784 0.146333
R5323 VDDA.n2897 VDDA.n2784 0.146333
R5324 VDDA.n2897 VDDA.n2782 0.146333
R5325 VDDA.n2907 VDDA.n2778 0.146333
R5326 VDDA.n2913 VDDA.n2778 0.146333
R5327 VDDA.n2913 VDDA.n2776 0.146333
R5328 VDDA.n2923 VDDA.n2772 0.146333
R5329 VDDA.n2927 VDDA.n2772 0.146333
R5330 VDDA.n2927 VDDA.n2770 0.146333
R5331 VDDA.n2669 VDDA.n2668 0.146333
R5332 VDDA.n2672 VDDA.n2669 0.146333
R5333 VDDA.n2672 VDDA.n2662 0.146333
R5334 VDDA.n2680 VDDA.n2658 0.146333
R5335 VDDA.n2684 VDDA.n2658 0.146333
R5336 VDDA.n2685 VDDA.n2684 0.146333
R5337 VDDA.n2693 VDDA.n2692 0.146333
R5338 VDDA.n2696 VDDA.n2693 0.146333
R5339 VDDA.n2696 VDDA.n2650 0.146333
R5340 VDDA.n2704 VDDA.n2646 0.146333
R5341 VDDA.n2708 VDDA.n2646 0.146333
R5342 VDDA.n2709 VDDA.n2708 0.146333
R5343 VDDA.n2717 VDDA.n2716 0.146333
R5344 VDDA.n2720 VDDA.n2717 0.146333
R5345 VDDA.n2720 VDDA.n2638 0.146333
R5346 VDDA.n2728 VDDA.n2634 0.146333
R5347 VDDA.n2732 VDDA.n2634 0.146333
R5348 VDDA.n2733 VDDA.n2732 0.146333
R5349 VDDA.n2741 VDDA.n2740 0.146333
R5350 VDDA.n2744 VDDA.n2741 0.146333
R5351 VDDA.n2744 VDDA.n2626 0.146333
R5352 VDDA.n2752 VDDA.n2624 0.146333
R5353 VDDA.n2756 VDDA.n2624 0.146333
R5354 VDDA.n2756 VDDA.n195 0.146333
R5355 VDDA.n269 VDDA.n265 0.146333
R5356 VDDA.n273 VDDA.n265 0.146333
R5357 VDDA.n274 VDDA.n273 0.146333
R5358 VDDA.n282 VDDA.n281 0.146333
R5359 VDDA.n285 VDDA.n282 0.146333
R5360 VDDA.n285 VDDA.n257 0.146333
R5361 VDDA.n293 VDDA.n253 0.146333
R5362 VDDA.n297 VDDA.n253 0.146333
R5363 VDDA.n298 VDDA.n297 0.146333
R5364 VDDA.n306 VDDA.n305 0.146333
R5365 VDDA.n309 VDDA.n306 0.146333
R5366 VDDA.n309 VDDA.n245 0.146333
R5367 VDDA.n317 VDDA.n241 0.146333
R5368 VDDA.n321 VDDA.n241 0.146333
R5369 VDDA.n322 VDDA.n321 0.146333
R5370 VDDA.n330 VDDA.n329 0.146333
R5371 VDDA.n333 VDDA.n330 0.146333
R5372 VDDA.n333 VDDA.n233 0.146333
R5373 VDDA.n341 VDDA.n229 0.146333
R5374 VDDA.n345 VDDA.n229 0.146333
R5375 VDDA.n346 VDDA.n345 0.146333
R5376 VDDA.n354 VDDA.n353 0.146333
R5377 VDDA.n357 VDDA.n354 0.146333
R5378 VDDA.n357 VDDA.n223 0.146333
R5379 VDDA.n2469 VDDA.n2466 0.146333
R5380 VDDA.n2475 VDDA.n2466 0.146333
R5381 VDDA.n2475 VDDA.n2464 0.146333
R5382 VDDA.n2485 VDDA.n2460 0.146333
R5383 VDDA.n2489 VDDA.n2460 0.146333
R5384 VDDA.n2489 VDDA.n2458 0.146333
R5385 VDDA.n2499 VDDA.n2454 0.146333
R5386 VDDA.n2505 VDDA.n2454 0.146333
R5387 VDDA.n2505 VDDA.n2452 0.146333
R5388 VDDA.n2515 VDDA.n2448 0.146333
R5389 VDDA.n2519 VDDA.n2448 0.146333
R5390 VDDA.n2519 VDDA.n2446 0.146333
R5391 VDDA.n2529 VDDA.n2442 0.146333
R5392 VDDA.n2535 VDDA.n2442 0.146333
R5393 VDDA.n2535 VDDA.n2440 0.146333
R5394 VDDA.n2545 VDDA.n2436 0.146333
R5395 VDDA.n2549 VDDA.n2436 0.146333
R5396 VDDA.n2549 VDDA.n2434 0.146333
R5397 VDDA.n2559 VDDA.n2430 0.146333
R5398 VDDA.n2565 VDDA.n2430 0.146333
R5399 VDDA.n2565 VDDA.n2428 0.146333
R5400 VDDA.n2575 VDDA.n2424 0.146333
R5401 VDDA.n2579 VDDA.n2424 0.146333
R5402 VDDA.n2579 VDDA.n2422 0.146333
R5403 VDDA.n1231 VDDA.n1230 0.146333
R5404 VDDA.n1234 VDDA.n1231 0.146333
R5405 VDDA.n1234 VDDA.n1224 0.146333
R5406 VDDA.n1242 VDDA.n1220 0.146333
R5407 VDDA.n1246 VDDA.n1220 0.146333
R5408 VDDA.n1247 VDDA.n1246 0.146333
R5409 VDDA.n1255 VDDA.n1254 0.146333
R5410 VDDA.n1258 VDDA.n1255 0.146333
R5411 VDDA.n1258 VDDA.n1212 0.146333
R5412 VDDA.n1266 VDDA.n1208 0.146333
R5413 VDDA.n1270 VDDA.n1208 0.146333
R5414 VDDA.n1271 VDDA.n1270 0.146333
R5415 VDDA.n1279 VDDA.n1278 0.146333
R5416 VDDA.n1282 VDDA.n1279 0.146333
R5417 VDDA.n1282 VDDA.n1200 0.146333
R5418 VDDA.n1290 VDDA.n1196 0.146333
R5419 VDDA.n1294 VDDA.n1196 0.146333
R5420 VDDA.n1295 VDDA.n1294 0.146333
R5421 VDDA.n1303 VDDA.n1302 0.146333
R5422 VDDA.n1306 VDDA.n1303 0.146333
R5423 VDDA.n1306 VDDA.n1188 0.146333
R5424 VDDA.n1314 VDDA.n1186 0.146333
R5425 VDDA.n1318 VDDA.n1186 0.146333
R5426 VDDA.n1318 VDDA.n462 0.146333
R5427 VDDA.n536 VDDA.n532 0.146333
R5428 VDDA.n540 VDDA.n532 0.146333
R5429 VDDA.n541 VDDA.n540 0.146333
R5430 VDDA.n549 VDDA.n548 0.146333
R5431 VDDA.n552 VDDA.n549 0.146333
R5432 VDDA.n552 VDDA.n524 0.146333
R5433 VDDA.n560 VDDA.n520 0.146333
R5434 VDDA.n564 VDDA.n520 0.146333
R5435 VDDA.n565 VDDA.n564 0.146333
R5436 VDDA.n573 VDDA.n572 0.146333
R5437 VDDA.n576 VDDA.n573 0.146333
R5438 VDDA.n576 VDDA.n512 0.146333
R5439 VDDA.n584 VDDA.n508 0.146333
R5440 VDDA.n588 VDDA.n508 0.146333
R5441 VDDA.n589 VDDA.n588 0.146333
R5442 VDDA.n597 VDDA.n596 0.146333
R5443 VDDA.n600 VDDA.n597 0.146333
R5444 VDDA.n600 VDDA.n500 0.146333
R5445 VDDA.n608 VDDA.n496 0.146333
R5446 VDDA.n612 VDDA.n496 0.146333
R5447 VDDA.n613 VDDA.n612 0.146333
R5448 VDDA.n621 VDDA.n620 0.146333
R5449 VDDA.n624 VDDA.n621 0.146333
R5450 VDDA.n624 VDDA.n490 0.146333
R5451 VDDA.n1031 VDDA.n1028 0.146333
R5452 VDDA.n1037 VDDA.n1028 0.146333
R5453 VDDA.n1037 VDDA.n1026 0.146333
R5454 VDDA.n1047 VDDA.n1022 0.146333
R5455 VDDA.n1051 VDDA.n1022 0.146333
R5456 VDDA.n1051 VDDA.n1020 0.146333
R5457 VDDA.n1061 VDDA.n1016 0.146333
R5458 VDDA.n1067 VDDA.n1016 0.146333
R5459 VDDA.n1067 VDDA.n1014 0.146333
R5460 VDDA.n1077 VDDA.n1010 0.146333
R5461 VDDA.n1081 VDDA.n1010 0.146333
R5462 VDDA.n1081 VDDA.n1008 0.146333
R5463 VDDA.n1091 VDDA.n1004 0.146333
R5464 VDDA.n1097 VDDA.n1004 0.146333
R5465 VDDA.n1097 VDDA.n1002 0.146333
R5466 VDDA.n1107 VDDA.n998 0.146333
R5467 VDDA.n1111 VDDA.n998 0.146333
R5468 VDDA.n1111 VDDA.n996 0.146333
R5469 VDDA.n1121 VDDA.n992 0.146333
R5470 VDDA.n1127 VDDA.n992 0.146333
R5471 VDDA.n1127 VDDA.n990 0.146333
R5472 VDDA.n1137 VDDA.n986 0.146333
R5473 VDDA.n1141 VDDA.n986 0.146333
R5474 VDDA.n1141 VDDA.n984 0.146333
R5475 VDDA.n883 VDDA.n882 0.146333
R5476 VDDA.n886 VDDA.n883 0.146333
R5477 VDDA.n886 VDDA.n876 0.146333
R5478 VDDA.n894 VDDA.n872 0.146333
R5479 VDDA.n898 VDDA.n872 0.146333
R5480 VDDA.n899 VDDA.n898 0.146333
R5481 VDDA.n907 VDDA.n906 0.146333
R5482 VDDA.n910 VDDA.n907 0.146333
R5483 VDDA.n910 VDDA.n864 0.146333
R5484 VDDA.n918 VDDA.n860 0.146333
R5485 VDDA.n922 VDDA.n860 0.146333
R5486 VDDA.n923 VDDA.n922 0.146333
R5487 VDDA.n931 VDDA.n930 0.146333
R5488 VDDA.n934 VDDA.n931 0.146333
R5489 VDDA.n934 VDDA.n852 0.146333
R5490 VDDA.n942 VDDA.n848 0.146333
R5491 VDDA.n946 VDDA.n848 0.146333
R5492 VDDA.n947 VDDA.n946 0.146333
R5493 VDDA.n955 VDDA.n954 0.146333
R5494 VDDA.n958 VDDA.n955 0.146333
R5495 VDDA.n958 VDDA.n840 0.146333
R5496 VDDA.n966 VDDA.n838 0.146333
R5497 VDDA.n970 VDDA.n838 0.146333
R5498 VDDA.n970 VDDA.n639 0.146333
R5499 VDDA.n690 VDDA.n688 0.146333
R5500 VDDA.n696 VDDA.n688 0.146333
R5501 VDDA.n697 VDDA.n696 0.146333
R5502 VDDA.n707 VDDA.n706 0.146333
R5503 VDDA.n710 VDDA.n707 0.146333
R5504 VDDA.n710 VDDA.n684 0.146333
R5505 VDDA.n720 VDDA.n682 0.146333
R5506 VDDA.n726 VDDA.n682 0.146333
R5507 VDDA.n727 VDDA.n726 0.146333
R5508 VDDA.n737 VDDA.n736 0.146333
R5509 VDDA.n740 VDDA.n737 0.146333
R5510 VDDA.n740 VDDA.n678 0.146333
R5511 VDDA.n750 VDDA.n676 0.146333
R5512 VDDA.n756 VDDA.n676 0.146333
R5513 VDDA.n757 VDDA.n756 0.146333
R5514 VDDA.n767 VDDA.n766 0.146333
R5515 VDDA.n770 VDDA.n767 0.146333
R5516 VDDA.n770 VDDA.n672 0.146333
R5517 VDDA.n780 VDDA.n670 0.146333
R5518 VDDA.n786 VDDA.n670 0.146333
R5519 VDDA.n787 VDDA.n786 0.146333
R5520 VDDA.n797 VDDA.n796 0.146333
R5521 VDDA.n800 VDDA.n797 0.146333
R5522 VDDA.n800 VDDA.n666 0.146333
R5523 VDDA.n1806 VDDA.n1805 0.136864
R5524 VDDA.n1817 VDDA.n1387 0.136864
R5525 VDDA.n1836 VDDA.n1835 0.136864
R5526 VDDA.n1847 VDDA.n1381 0.136864
R5527 VDDA.n1866 VDDA.n1865 0.136864
R5528 VDDA.n1877 VDDA.n1375 0.136864
R5529 VDDA.n1896 VDDA.n1895 0.136864
R5530 VDDA.n1804 VDDA.n1390 0.136864
R5531 VDDA.n1821 VDDA.n1820 0.136864
R5532 VDDA.n1834 VDDA.n1384 0.136864
R5533 VDDA.n1851 VDDA.n1850 0.136864
R5534 VDDA.n1864 VDDA.n1378 0.136864
R5535 VDDA.n1881 VDDA.n1880 0.136864
R5536 VDDA.n1894 VDDA.n1372 0.136864
R5537 VDDA.n1462 VDDA.t69 0.1368
R5538 VDDA.n1462 VDDA.t52 0.1368
R5539 VDDA.n1461 VDDA.t99 0.1368
R5540 VDDA.n1461 VDDA.t392 0.1368
R5541 VDDA.n1460 VDDA.t387 0.1368
R5542 VDDA.n1460 VDDA.t137 0.1368
R5543 VDDA.n1459 VDDA.t58 0.1368
R5544 VDDA.n1459 VDDA.t68 0.1368
R5545 VDDA.n1458 VDDA.t394 0.1368
R5546 VDDA.n1458 VDDA.t174 0.1368
R5547 VDDA.n1466 VDDA.n1464 0.135917
R5548 VDDA.n1476 VDDA.n1473 0.135917
R5549 VDDA.n1482 VDDA.n1455 0.135917
R5550 VDDA.n1492 VDDA.n1453 0.135917
R5551 VDDA.n1496 VDDA.n1493 0.135917
R5552 VDDA.n1506 VDDA.n1503 0.135917
R5553 VDDA.n1512 VDDA.n1449 0.135917
R5554 VDDA.n1522 VDDA.n1447 0.135917
R5555 VDDA.n1526 VDDA.n1523 0.135917
R5556 VDDA.n1536 VDDA.n1533 0.135917
R5557 VDDA.n1542 VDDA.n1443 0.135917
R5558 VDDA.n1552 VDDA.n1441 0.135917
R5559 VDDA.n1556 VDDA.n1553 0.135917
R5560 VDDA.n1566 VDDA.n1563 0.135917
R5561 VDDA.n1572 VDDA.n1437 0.135917
R5562 VDDA.n2153 VDDA.n2150 0.135917
R5563 VDDA.n2159 VDDA.n1930 0.135917
R5564 VDDA.n2169 VDDA.n1928 0.135917
R5565 VDDA.n2173 VDDA.n2170 0.135917
R5566 VDDA.n2183 VDDA.n2180 0.135917
R5567 VDDA.n2189 VDDA.n1924 0.135917
R5568 VDDA.n2199 VDDA.n1922 0.135917
R5569 VDDA.n2203 VDDA.n2200 0.135917
R5570 VDDA.n2213 VDDA.n2210 0.135917
R5571 VDDA.n2219 VDDA.n1918 0.135917
R5572 VDDA.n2229 VDDA.n1916 0.135917
R5573 VDDA.n2233 VDDA.n2230 0.135917
R5574 VDDA.n2243 VDDA.n2240 0.135917
R5575 VDDA.n2249 VDDA.n1912 0.135917
R5576 VDDA.n99 VDDA.n96 0.135917
R5577 VDDA.n103 VDDA.n83 0.135917
R5578 VDDA.n111 VDDA.n79 0.135917
R5579 VDDA.n115 VDDA.n112 0.135917
R5580 VDDA.n123 VDDA.n120 0.135917
R5581 VDDA.n127 VDDA.n71 0.135917
R5582 VDDA.n135 VDDA.n67 0.135917
R5583 VDDA.n139 VDDA.n136 0.135917
R5584 VDDA.n147 VDDA.n144 0.135917
R5585 VDDA.n151 VDDA.n59 0.135917
R5586 VDDA.n159 VDDA.n55 0.135917
R5587 VDDA.n163 VDDA.n160 0.135917
R5588 VDDA.n171 VDDA.n168 0.135917
R5589 VDDA.n175 VDDA.n47 0.135917
R5590 VDDA.n2945 VDDA.n45 0.135917
R5591 VDDA.n2827 VDDA.n2812 0.135917
R5592 VDDA.n2833 VDDA.n2810 0.135917
R5593 VDDA.n2843 VDDA.n2806 0.135917
R5594 VDDA.n2847 VDDA.n2804 0.135917
R5595 VDDA.n2857 VDDA.n2800 0.135917
R5596 VDDA.n2863 VDDA.n2798 0.135917
R5597 VDDA.n2873 VDDA.n2794 0.135917
R5598 VDDA.n2877 VDDA.n2792 0.135917
R5599 VDDA.n2887 VDDA.n2788 0.135917
R5600 VDDA.n2893 VDDA.n2786 0.135917
R5601 VDDA.n2903 VDDA.n2782 0.135917
R5602 VDDA.n2907 VDDA.n2780 0.135917
R5603 VDDA.n2917 VDDA.n2776 0.135917
R5604 VDDA.n2923 VDDA.n2774 0.135917
R5605 VDDA.n2932 VDDA.n2770 0.135917
R5606 VDDA.n2676 VDDA.n2662 0.135917
R5607 VDDA.n2680 VDDA.n2677 0.135917
R5608 VDDA.n2688 VDDA.n2685 0.135917
R5609 VDDA.n2692 VDDA.n2654 0.135917
R5610 VDDA.n2700 VDDA.n2650 0.135917
R5611 VDDA.n2704 VDDA.n2701 0.135917
R5612 VDDA.n2712 VDDA.n2709 0.135917
R5613 VDDA.n2716 VDDA.n2642 0.135917
R5614 VDDA.n2724 VDDA.n2638 0.135917
R5615 VDDA.n2728 VDDA.n2725 0.135917
R5616 VDDA.n2736 VDDA.n2733 0.135917
R5617 VDDA.n2740 VDDA.n2630 0.135917
R5618 VDDA.n2748 VDDA.n2626 0.135917
R5619 VDDA.n2752 VDDA.n2749 0.135917
R5620 VDDA.n2761 VDDA.n195 0.135917
R5621 VDDA.n277 VDDA.n274 0.135917
R5622 VDDA.n281 VDDA.n261 0.135917
R5623 VDDA.n289 VDDA.n257 0.135917
R5624 VDDA.n293 VDDA.n290 0.135917
R5625 VDDA.n301 VDDA.n298 0.135917
R5626 VDDA.n305 VDDA.n249 0.135917
R5627 VDDA.n313 VDDA.n245 0.135917
R5628 VDDA.n317 VDDA.n314 0.135917
R5629 VDDA.n325 VDDA.n322 0.135917
R5630 VDDA.n329 VDDA.n237 0.135917
R5631 VDDA.n337 VDDA.n233 0.135917
R5632 VDDA.n341 VDDA.n338 0.135917
R5633 VDDA.n349 VDDA.n346 0.135917
R5634 VDDA.n353 VDDA.n225 0.135917
R5635 VDDA.n2597 VDDA.n223 0.135917
R5636 VDDA.n2479 VDDA.n2464 0.135917
R5637 VDDA.n2485 VDDA.n2462 0.135917
R5638 VDDA.n2495 VDDA.n2458 0.135917
R5639 VDDA.n2499 VDDA.n2456 0.135917
R5640 VDDA.n2509 VDDA.n2452 0.135917
R5641 VDDA.n2515 VDDA.n2450 0.135917
R5642 VDDA.n2525 VDDA.n2446 0.135917
R5643 VDDA.n2529 VDDA.n2444 0.135917
R5644 VDDA.n2539 VDDA.n2440 0.135917
R5645 VDDA.n2545 VDDA.n2438 0.135917
R5646 VDDA.n2555 VDDA.n2434 0.135917
R5647 VDDA.n2559 VDDA.n2432 0.135917
R5648 VDDA.n2569 VDDA.n2428 0.135917
R5649 VDDA.n2575 VDDA.n2426 0.135917
R5650 VDDA.n2584 VDDA.n2422 0.135917
R5651 VDDA.n1238 VDDA.n1224 0.135917
R5652 VDDA.n1242 VDDA.n1239 0.135917
R5653 VDDA.n1250 VDDA.n1247 0.135917
R5654 VDDA.n1254 VDDA.n1216 0.135917
R5655 VDDA.n1262 VDDA.n1212 0.135917
R5656 VDDA.n1266 VDDA.n1263 0.135917
R5657 VDDA.n1274 VDDA.n1271 0.135917
R5658 VDDA.n1278 VDDA.n1204 0.135917
R5659 VDDA.n1286 VDDA.n1200 0.135917
R5660 VDDA.n1290 VDDA.n1287 0.135917
R5661 VDDA.n1298 VDDA.n1295 0.135917
R5662 VDDA.n1302 VDDA.n1192 0.135917
R5663 VDDA.n1310 VDDA.n1188 0.135917
R5664 VDDA.n1314 VDDA.n1311 0.135917
R5665 VDDA.n2260 VDDA.n462 0.135917
R5666 VDDA.n544 VDDA.n541 0.135917
R5667 VDDA.n548 VDDA.n528 0.135917
R5668 VDDA.n556 VDDA.n524 0.135917
R5669 VDDA.n560 VDDA.n557 0.135917
R5670 VDDA.n568 VDDA.n565 0.135917
R5671 VDDA.n572 VDDA.n516 0.135917
R5672 VDDA.n580 VDDA.n512 0.135917
R5673 VDDA.n584 VDDA.n581 0.135917
R5674 VDDA.n592 VDDA.n589 0.135917
R5675 VDDA.n596 VDDA.n504 0.135917
R5676 VDDA.n604 VDDA.n500 0.135917
R5677 VDDA.n608 VDDA.n605 0.135917
R5678 VDDA.n616 VDDA.n613 0.135917
R5679 VDDA.n620 VDDA.n492 0.135917
R5680 VDDA.n1159 VDDA.n490 0.135917
R5681 VDDA.n1041 VDDA.n1026 0.135917
R5682 VDDA.n1047 VDDA.n1024 0.135917
R5683 VDDA.n1057 VDDA.n1020 0.135917
R5684 VDDA.n1061 VDDA.n1018 0.135917
R5685 VDDA.n1071 VDDA.n1014 0.135917
R5686 VDDA.n1077 VDDA.n1012 0.135917
R5687 VDDA.n1087 VDDA.n1008 0.135917
R5688 VDDA.n1091 VDDA.n1006 0.135917
R5689 VDDA.n1101 VDDA.n1002 0.135917
R5690 VDDA.n1107 VDDA.n1000 0.135917
R5691 VDDA.n1117 VDDA.n996 0.135917
R5692 VDDA.n1121 VDDA.n994 0.135917
R5693 VDDA.n1131 VDDA.n990 0.135917
R5694 VDDA.n1137 VDDA.n988 0.135917
R5695 VDDA.n1146 VDDA.n984 0.135917
R5696 VDDA.n890 VDDA.n876 0.135917
R5697 VDDA.n894 VDDA.n891 0.135917
R5698 VDDA.n902 VDDA.n899 0.135917
R5699 VDDA.n906 VDDA.n868 0.135917
R5700 VDDA.n914 VDDA.n864 0.135917
R5701 VDDA.n918 VDDA.n915 0.135917
R5702 VDDA.n926 VDDA.n923 0.135917
R5703 VDDA.n930 VDDA.n856 0.135917
R5704 VDDA.n938 VDDA.n852 0.135917
R5705 VDDA.n942 VDDA.n939 0.135917
R5706 VDDA.n950 VDDA.n947 0.135917
R5707 VDDA.n954 VDDA.n844 0.135917
R5708 VDDA.n962 VDDA.n840 0.135917
R5709 VDDA.n966 VDDA.n963 0.135917
R5710 VDDA.n975 VDDA.n639 0.135917
R5711 VDDA.n700 VDDA.n697 0.135917
R5712 VDDA.n706 VDDA.n686 0.135917
R5713 VDDA.n716 VDDA.n684 0.135917
R5714 VDDA.n720 VDDA.n717 0.135917
R5715 VDDA.n730 VDDA.n727 0.135917
R5716 VDDA.n736 VDDA.n680 0.135917
R5717 VDDA.n746 VDDA.n678 0.135917
R5718 VDDA.n750 VDDA.n747 0.135917
R5719 VDDA.n760 VDDA.n757 0.135917
R5720 VDDA.n766 VDDA.n674 0.135917
R5721 VDDA.n776 VDDA.n672 0.135917
R5722 VDDA.n780 VDDA.n777 0.135917
R5723 VDDA.n790 VDDA.n787 0.135917
R5724 VDDA.n796 VDDA.n668 0.135917
R5725 VDDA.n811 VDDA.n666 0.135917
R5726 VDDA.n1476 VDDA.n1455 0.1255
R5727 VDDA.n1493 VDDA.n1492 0.1255
R5728 VDDA.n1506 VDDA.n1449 0.1255
R5729 VDDA.n1523 VDDA.n1522 0.1255
R5730 VDDA.n1536 VDDA.n1443 0.1255
R5731 VDDA.n1553 VDDA.n1552 0.1255
R5732 VDDA.n1566 VDDA.n1437 0.1255
R5733 VDDA.n2136 VDDA.n2135 0.1255
R5734 VDDA.n2135 VDDA.n2134 0.1255
R5735 VDDA.n2009 VDDA.n1952 0.1255
R5736 VDDA.n1956 VDDA.n1952 0.1255
R5737 VDDA.n1958 VDDA.n1956 0.1255
R5738 VDDA.n1960 VDDA.n1958 0.1255
R5739 VDDA.n1962 VDDA.n1960 0.1255
R5740 VDDA.n1964 VDDA.n1962 0.1255
R5741 VDDA.n1966 VDDA.n1964 0.1255
R5742 VDDA.n1968 VDDA.n1966 0.1255
R5743 VDDA.n1970 VDDA.n1968 0.1255
R5744 VDDA.n2000 VDDA.n1970 0.1255
R5745 VDDA.n1999 VDDA.n1972 0.1255
R5746 VDDA.n1976 VDDA.n1972 0.1255
R5747 VDDA.n1978 VDDA.n1976 0.1255
R5748 VDDA.n1980 VDDA.n1978 0.1255
R5749 VDDA.n1982 VDDA.n1980 0.1255
R5750 VDDA.n1984 VDDA.n1982 0.1255
R5751 VDDA.n1986 VDDA.n1984 0.1255
R5752 VDDA.n1988 VDDA.n1986 0.1255
R5753 VDDA.n1990 VDDA.n1988 0.1255
R5754 VDDA.n2153 VDDA.n1930 0.1255
R5755 VDDA.n2170 VDDA.n2169 0.1255
R5756 VDDA.n2183 VDDA.n1924 0.1255
R5757 VDDA.n2200 VDDA.n2199 0.1255
R5758 VDDA.n2213 VDDA.n1918 0.1255
R5759 VDDA.n2230 VDDA.n2229 0.1255
R5760 VDDA.n2243 VDDA.n1912 0.1255
R5761 VDDA.n99 VDDA.n83 0.1255
R5762 VDDA.n112 VDDA.n111 0.1255
R5763 VDDA.n123 VDDA.n71 0.1255
R5764 VDDA.n136 VDDA.n135 0.1255
R5765 VDDA.n147 VDDA.n59 0.1255
R5766 VDDA.n160 VDDA.n159 0.1255
R5767 VDDA.n171 VDDA.n47 0.1255
R5768 VDDA.n2827 VDDA.n2810 0.1255
R5769 VDDA.n2843 VDDA.n2804 0.1255
R5770 VDDA.n2857 VDDA.n2798 0.1255
R5771 VDDA.n2873 VDDA.n2792 0.1255
R5772 VDDA.n2887 VDDA.n2786 0.1255
R5773 VDDA.n2903 VDDA.n2780 0.1255
R5774 VDDA.n2917 VDDA.n2774 0.1255
R5775 VDDA.n2677 VDDA.n2676 0.1255
R5776 VDDA.n2688 VDDA.n2654 0.1255
R5777 VDDA.n2701 VDDA.n2700 0.1255
R5778 VDDA.n2712 VDDA.n2642 0.1255
R5779 VDDA.n2725 VDDA.n2724 0.1255
R5780 VDDA.n2736 VDDA.n2630 0.1255
R5781 VDDA.n2749 VDDA.n2748 0.1255
R5782 VDDA.n277 VDDA.n261 0.1255
R5783 VDDA.n290 VDDA.n289 0.1255
R5784 VDDA.n301 VDDA.n249 0.1255
R5785 VDDA.n314 VDDA.n313 0.1255
R5786 VDDA.n325 VDDA.n237 0.1255
R5787 VDDA.n338 VDDA.n337 0.1255
R5788 VDDA.n349 VDDA.n225 0.1255
R5789 VDDA.n2479 VDDA.n2462 0.1255
R5790 VDDA.n2495 VDDA.n2456 0.1255
R5791 VDDA.n2509 VDDA.n2450 0.1255
R5792 VDDA.n2525 VDDA.n2444 0.1255
R5793 VDDA.n2539 VDDA.n2438 0.1255
R5794 VDDA.n2555 VDDA.n2432 0.1255
R5795 VDDA.n2569 VDDA.n2426 0.1255
R5796 VDDA.n1239 VDDA.n1238 0.1255
R5797 VDDA.n1250 VDDA.n1216 0.1255
R5798 VDDA.n1263 VDDA.n1262 0.1255
R5799 VDDA.n1274 VDDA.n1204 0.1255
R5800 VDDA.n1287 VDDA.n1286 0.1255
R5801 VDDA.n1298 VDDA.n1192 0.1255
R5802 VDDA.n1311 VDDA.n1310 0.1255
R5803 VDDA.n377 VDDA.n372 0.1255
R5804 VDDA.n384 VDDA.n378 0.1255
R5805 VDDA.n544 VDDA.n528 0.1255
R5806 VDDA.n557 VDDA.n556 0.1255
R5807 VDDA.n568 VDDA.n516 0.1255
R5808 VDDA.n581 VDDA.n580 0.1255
R5809 VDDA.n592 VDDA.n504 0.1255
R5810 VDDA.n605 VDDA.n604 0.1255
R5811 VDDA.n616 VDDA.n492 0.1255
R5812 VDDA.n1041 VDDA.n1024 0.1255
R5813 VDDA.n1057 VDDA.n1018 0.1255
R5814 VDDA.n1071 VDDA.n1012 0.1255
R5815 VDDA.n1087 VDDA.n1006 0.1255
R5816 VDDA.n1101 VDDA.n1000 0.1255
R5817 VDDA.n1117 VDDA.n994 0.1255
R5818 VDDA.n1131 VDDA.n988 0.1255
R5819 VDDA.n891 VDDA.n890 0.1255
R5820 VDDA.n902 VDDA.n868 0.1255
R5821 VDDA.n915 VDDA.n914 0.1255
R5822 VDDA.n926 VDDA.n856 0.1255
R5823 VDDA.n939 VDDA.n938 0.1255
R5824 VDDA.n950 VDDA.n844 0.1255
R5825 VDDA.n963 VDDA.n962 0.1255
R5826 VDDA.n700 VDDA.n686 0.1255
R5827 VDDA.n717 VDDA.n716 0.1255
R5828 VDDA.n730 VDDA.n680 0.1255
R5829 VDDA.n747 VDDA.n746 0.1255
R5830 VDDA.n760 VDDA.n674 0.1255
R5831 VDDA.n777 VDDA.n776 0.1255
R5832 VDDA.n790 VDDA.n668 0.1255
R5833 VDDA.n1768 VDDA.n1767 0.123287
R5834 VDDA.n1790 VDDA.n1789 0.123287
R5835 VDDA.n2133 VDDA.n2132 0.115083
R5836 VDDA.n2132 VDDA.n2131 0.115083
R5837 VDDA.n2131 VDDA.n2130 0.115083
R5838 VDDA.n2128 VDDA.n2127 0.115083
R5839 VDDA.n2127 VDDA.n2126 0.115083
R5840 VDDA.n2126 VDDA.n2125 0.115083
R5841 VDDA.n2125 VDDA.n2124 0.115083
R5842 VDDA.n2122 VDDA.n2121 0.115083
R5843 VDDA.n2121 VDDA.n2120 0.115083
R5844 VDDA.n2316 VDDA.n2314 0.115083
R5845 VDDA.n2318 VDDA.n2316 0.115083
R5846 VDDA.n2320 VDDA.n2318 0.115083
R5847 VDDA.n2322 VDDA.n2320 0.115083
R5848 VDDA.n425 VDDA.n423 0.115083
R5849 VDDA.n423 VDDA.n421 0.115083
R5850 VDDA.n421 VDDA.n419 0.115083
R5851 VDDA.n419 VDDA.n417 0.115083
R5852 VDDA.n2300 VDDA.n2298 0.115083
R5853 VDDA.n2298 VDDA.n2296 0.115083
R5854 VDDA.n2296 VDDA.n2294 0.115083
R5855 VDDA.n2294 VDDA.n2292 0.115083
R5856 VDDA.n2305 VDDA.n2292 0.115083
R5857 VDDA.n405 VDDA.n392 0.115083
R5858 VDDA.n394 VDDA.n392 0.115083
R5859 VDDA.n396 VDDA.n394 0.115083
R5860 VDDA.n398 VDDA.n396 0.115083
R5861 VDDA.n400 VDDA.n398 0.115083
R5862 VDDA.n2365 VDDA.n2364 0.0838333
R5863 VDDA.n1763 VDDA.n1407 0.076587
R5864 VDDA.n1582 VDDA.n1407 0.076587
R5865 VDDA.n1755 VDDA.n1582 0.076587
R5866 VDDA.n1745 VDDA.n1587 0.076587
R5867 VDDA.n1745 VDDA.n1591 0.076587
R5868 VDDA.n1741 VDDA.n1591 0.076587
R5869 VDDA.n1731 VDDA.n1597 0.076587
R5870 VDDA.n1731 VDDA.n1599 0.076587
R5871 VDDA.n1725 VDDA.n1599 0.076587
R5872 VDDA.n1715 VDDA.n1605 0.076587
R5873 VDDA.n1715 VDDA.n1609 0.076587
R5874 VDDA.n1711 VDDA.n1609 0.076587
R5875 VDDA.n1701 VDDA.n1615 0.076587
R5876 VDDA.n1701 VDDA.n1617 0.076587
R5877 VDDA.n1695 VDDA.n1617 0.076587
R5878 VDDA.n1685 VDDA.n1623 0.076587
R5879 VDDA.n1685 VDDA.n1627 0.076587
R5880 VDDA.n1681 VDDA.n1627 0.076587
R5881 VDDA.n1671 VDDA.n1633 0.076587
R5882 VDDA.n1671 VDDA.n1635 0.076587
R5883 VDDA.n1665 VDDA.n1635 0.076587
R5884 VDDA.n1655 VDDA.n1641 0.076587
R5885 VDDA.n1655 VDDA.n1645 0.076587
R5886 VDDA.n1651 VDDA.n1645 0.076587
R5887 VDDA.n1764 VDDA.n1406 0.076587
R5888 VDDA.n1585 VDDA.n1406 0.076587
R5889 VDDA.n1754 VDDA.n1585 0.076587
R5890 VDDA.n1744 VDDA.n1586 0.076587
R5891 VDDA.n1744 VDDA.n1743 0.076587
R5892 VDDA.n1743 VDDA.n1742 0.076587
R5893 VDDA.n1733 VDDA.n1732 0.076587
R5894 VDDA.n1732 VDDA.n1598 0.076587
R5895 VDDA.n1724 VDDA.n1598 0.076587
R5896 VDDA.n1714 VDDA.n1604 0.076587
R5897 VDDA.n1714 VDDA.n1713 0.076587
R5898 VDDA.n1713 VDDA.n1712 0.076587
R5899 VDDA.n1703 VDDA.n1702 0.076587
R5900 VDDA.n1702 VDDA.n1616 0.076587
R5901 VDDA.n1694 VDDA.n1616 0.076587
R5902 VDDA.n1684 VDDA.n1622 0.076587
R5903 VDDA.n1684 VDDA.n1683 0.076587
R5904 VDDA.n1683 VDDA.n1682 0.076587
R5905 VDDA.n1673 VDDA.n1672 0.076587
R5906 VDDA.n1672 VDDA.n1634 0.076587
R5907 VDDA.n1664 VDDA.n1634 0.076587
R5908 VDDA.n1654 VDDA.n1640 0.076587
R5909 VDDA.n1654 VDDA.n1653 0.076587
R5910 VDDA.n1468 VDDA.n1467 0.0734167
R5911 VDDA.n1469 VDDA.n1468 0.0734167
R5912 VDDA.n1469 VDDA.n1456 0.0734167
R5913 VDDA.n1479 VDDA.n1454 0.0734167
R5914 VDDA.n1487 VDDA.n1454 0.0734167
R5915 VDDA.n1488 VDDA.n1487 0.0734167
R5916 VDDA.n1498 VDDA.n1497 0.0734167
R5917 VDDA.n1499 VDDA.n1498 0.0734167
R5918 VDDA.n1499 VDDA.n1450 0.0734167
R5919 VDDA.n1509 VDDA.n1448 0.0734167
R5920 VDDA.n1517 VDDA.n1448 0.0734167
R5921 VDDA.n1518 VDDA.n1517 0.0734167
R5922 VDDA.n1528 VDDA.n1527 0.0734167
R5923 VDDA.n1529 VDDA.n1528 0.0734167
R5924 VDDA.n1529 VDDA.n1444 0.0734167
R5925 VDDA.n1539 VDDA.n1442 0.0734167
R5926 VDDA.n1547 VDDA.n1442 0.0734167
R5927 VDDA.n1548 VDDA.n1547 0.0734167
R5928 VDDA.n1558 VDDA.n1557 0.0734167
R5929 VDDA.n1559 VDDA.n1558 0.0734167
R5930 VDDA.n1559 VDDA.n1438 0.0734167
R5931 VDDA.n1569 VDDA.n1436 0.0734167
R5932 VDDA.n1577 VDDA.n1436 0.0734167
R5933 VDDA.n2145 VDDA.n2144 0.0734167
R5934 VDDA.n2146 VDDA.n2145 0.0734167
R5935 VDDA.n2146 VDDA.n1931 0.0734167
R5936 VDDA.n2156 VDDA.n1929 0.0734167
R5937 VDDA.n2164 VDDA.n1929 0.0734167
R5938 VDDA.n2165 VDDA.n2164 0.0734167
R5939 VDDA.n2175 VDDA.n2174 0.0734167
R5940 VDDA.n2176 VDDA.n2175 0.0734167
R5941 VDDA.n2176 VDDA.n1925 0.0734167
R5942 VDDA.n2186 VDDA.n1923 0.0734167
R5943 VDDA.n2194 VDDA.n1923 0.0734167
R5944 VDDA.n2195 VDDA.n2194 0.0734167
R5945 VDDA.n2205 VDDA.n2204 0.0734167
R5946 VDDA.n2206 VDDA.n2205 0.0734167
R5947 VDDA.n2206 VDDA.n1919 0.0734167
R5948 VDDA.n2216 VDDA.n1917 0.0734167
R5949 VDDA.n2224 VDDA.n1917 0.0734167
R5950 VDDA.n2225 VDDA.n2224 0.0734167
R5951 VDDA.n2235 VDDA.n2234 0.0734167
R5952 VDDA.n2236 VDDA.n2235 0.0734167
R5953 VDDA.n2236 VDDA.n1913 0.0734167
R5954 VDDA.n2246 VDDA.n1911 0.0734167
R5955 VDDA.n2254 VDDA.n1911 0.0734167
R5956 VDDA.n94 VDDA.n93 0.0734167
R5957 VDDA.n94 VDDA.n86 0.0734167
R5958 VDDA.n102 VDDA.n82 0.0734167
R5959 VDDA.n108 VDDA.n82 0.0734167
R5960 VDDA.n109 VDDA.n108 0.0734167
R5961 VDDA.n117 VDDA.n116 0.0734167
R5962 VDDA.n118 VDDA.n117 0.0734167
R5963 VDDA.n118 VDDA.n74 0.0734167
R5964 VDDA.n126 VDDA.n70 0.0734167
R5965 VDDA.n132 VDDA.n70 0.0734167
R5966 VDDA.n133 VDDA.n132 0.0734167
R5967 VDDA.n141 VDDA.n140 0.0734167
R5968 VDDA.n142 VDDA.n141 0.0734167
R5969 VDDA.n142 VDDA.n62 0.0734167
R5970 VDDA.n150 VDDA.n58 0.0734167
R5971 VDDA.n156 VDDA.n58 0.0734167
R5972 VDDA.n157 VDDA.n156 0.0734167
R5973 VDDA.n165 VDDA.n164 0.0734167
R5974 VDDA.n166 VDDA.n165 0.0734167
R5975 VDDA.n166 VDDA.n50 0.0734167
R5976 VDDA.n174 VDDA.n46 0.0734167
R5977 VDDA.n180 VDDA.n46 0.0734167
R5978 VDDA.n181 VDDA.n180 0.0734167
R5979 VDDA.n2824 VDDA.n2813 0.0734167
R5980 VDDA.n2825 VDDA.n2824 0.0734167
R5981 VDDA.n2835 VDDA.n2834 0.0734167
R5982 VDDA.n2836 VDDA.n2835 0.0734167
R5983 VDDA.n2836 VDDA.n2805 0.0734167
R5984 VDDA.n2846 VDDA.n2801 0.0734167
R5985 VDDA.n2854 VDDA.n2801 0.0734167
R5986 VDDA.n2855 VDDA.n2854 0.0734167
R5987 VDDA.n2865 VDDA.n2864 0.0734167
R5988 VDDA.n2866 VDDA.n2865 0.0734167
R5989 VDDA.n2866 VDDA.n2793 0.0734167
R5990 VDDA.n2876 VDDA.n2789 0.0734167
R5991 VDDA.n2884 VDDA.n2789 0.0734167
R5992 VDDA.n2885 VDDA.n2884 0.0734167
R5993 VDDA.n2895 VDDA.n2894 0.0734167
R5994 VDDA.n2896 VDDA.n2895 0.0734167
R5995 VDDA.n2896 VDDA.n2781 0.0734167
R5996 VDDA.n2906 VDDA.n2777 0.0734167
R5997 VDDA.n2914 VDDA.n2777 0.0734167
R5998 VDDA.n2915 VDDA.n2914 0.0734167
R5999 VDDA.n2925 VDDA.n2924 0.0734167
R6000 VDDA.n2926 VDDA.n2925 0.0734167
R6001 VDDA.n2926 VDDA.n2769 0.0734167
R6002 VDDA.n2673 VDDA.n2665 0.0734167
R6003 VDDA.n2674 VDDA.n2673 0.0734167
R6004 VDDA.n2682 VDDA.n2681 0.0734167
R6005 VDDA.n2683 VDDA.n2682 0.0734167
R6006 VDDA.n2683 VDDA.n2657 0.0734167
R6007 VDDA.n2691 VDDA.n2653 0.0734167
R6008 VDDA.n2697 VDDA.n2653 0.0734167
R6009 VDDA.n2698 VDDA.n2697 0.0734167
R6010 VDDA.n2706 VDDA.n2705 0.0734167
R6011 VDDA.n2707 VDDA.n2706 0.0734167
R6012 VDDA.n2707 VDDA.n2645 0.0734167
R6013 VDDA.n2715 VDDA.n2641 0.0734167
R6014 VDDA.n2721 VDDA.n2641 0.0734167
R6015 VDDA.n2722 VDDA.n2721 0.0734167
R6016 VDDA.n2730 VDDA.n2729 0.0734167
R6017 VDDA.n2731 VDDA.n2730 0.0734167
R6018 VDDA.n2731 VDDA.n2633 0.0734167
R6019 VDDA.n2739 VDDA.n2629 0.0734167
R6020 VDDA.n2745 VDDA.n2629 0.0734167
R6021 VDDA.n2746 VDDA.n2745 0.0734167
R6022 VDDA.n2754 VDDA.n2753 0.0734167
R6023 VDDA.n2755 VDDA.n2754 0.0734167
R6024 VDDA.n2755 VDDA.n194 0.0734167
R6025 VDDA.n272 VDDA.n271 0.0734167
R6026 VDDA.n272 VDDA.n264 0.0734167
R6027 VDDA.n280 VDDA.n260 0.0734167
R6028 VDDA.n286 VDDA.n260 0.0734167
R6029 VDDA.n287 VDDA.n286 0.0734167
R6030 VDDA.n295 VDDA.n294 0.0734167
R6031 VDDA.n296 VDDA.n295 0.0734167
R6032 VDDA.n296 VDDA.n252 0.0734167
R6033 VDDA.n304 VDDA.n248 0.0734167
R6034 VDDA.n310 VDDA.n248 0.0734167
R6035 VDDA.n311 VDDA.n310 0.0734167
R6036 VDDA.n319 VDDA.n318 0.0734167
R6037 VDDA.n320 VDDA.n319 0.0734167
R6038 VDDA.n320 VDDA.n240 0.0734167
R6039 VDDA.n328 VDDA.n236 0.0734167
R6040 VDDA.n334 VDDA.n236 0.0734167
R6041 VDDA.n335 VDDA.n334 0.0734167
R6042 VDDA.n343 VDDA.n342 0.0734167
R6043 VDDA.n344 VDDA.n343 0.0734167
R6044 VDDA.n344 VDDA.n228 0.0734167
R6045 VDDA.n352 VDDA.n224 0.0734167
R6046 VDDA.n358 VDDA.n224 0.0734167
R6047 VDDA.n359 VDDA.n358 0.0734167
R6048 VDDA.n2476 VDDA.n2465 0.0734167
R6049 VDDA.n2477 VDDA.n2476 0.0734167
R6050 VDDA.n2487 VDDA.n2486 0.0734167
R6051 VDDA.n2488 VDDA.n2487 0.0734167
R6052 VDDA.n2488 VDDA.n2457 0.0734167
R6053 VDDA.n2498 VDDA.n2453 0.0734167
R6054 VDDA.n2506 VDDA.n2453 0.0734167
R6055 VDDA.n2507 VDDA.n2506 0.0734167
R6056 VDDA.n2517 VDDA.n2516 0.0734167
R6057 VDDA.n2518 VDDA.n2517 0.0734167
R6058 VDDA.n2518 VDDA.n2445 0.0734167
R6059 VDDA.n2528 VDDA.n2441 0.0734167
R6060 VDDA.n2536 VDDA.n2441 0.0734167
R6061 VDDA.n2537 VDDA.n2536 0.0734167
R6062 VDDA.n2547 VDDA.n2546 0.0734167
R6063 VDDA.n2548 VDDA.n2547 0.0734167
R6064 VDDA.n2548 VDDA.n2433 0.0734167
R6065 VDDA.n2558 VDDA.n2429 0.0734167
R6066 VDDA.n2566 VDDA.n2429 0.0734167
R6067 VDDA.n2567 VDDA.n2566 0.0734167
R6068 VDDA.n2577 VDDA.n2576 0.0734167
R6069 VDDA.n2578 VDDA.n2577 0.0734167
R6070 VDDA.n2578 VDDA.n2421 0.0734167
R6071 VDDA.n1235 VDDA.n1227 0.0734167
R6072 VDDA.n1236 VDDA.n1235 0.0734167
R6073 VDDA.n1244 VDDA.n1243 0.0734167
R6074 VDDA.n1245 VDDA.n1244 0.0734167
R6075 VDDA.n1245 VDDA.n1219 0.0734167
R6076 VDDA.n1253 VDDA.n1215 0.0734167
R6077 VDDA.n1259 VDDA.n1215 0.0734167
R6078 VDDA.n1260 VDDA.n1259 0.0734167
R6079 VDDA.n1268 VDDA.n1267 0.0734167
R6080 VDDA.n1269 VDDA.n1268 0.0734167
R6081 VDDA.n1269 VDDA.n1207 0.0734167
R6082 VDDA.n1277 VDDA.n1203 0.0734167
R6083 VDDA.n1283 VDDA.n1203 0.0734167
R6084 VDDA.n1284 VDDA.n1283 0.0734167
R6085 VDDA.n1292 VDDA.n1291 0.0734167
R6086 VDDA.n1293 VDDA.n1292 0.0734167
R6087 VDDA.n1293 VDDA.n1195 0.0734167
R6088 VDDA.n1301 VDDA.n1191 0.0734167
R6089 VDDA.n1307 VDDA.n1191 0.0734167
R6090 VDDA.n1308 VDDA.n1307 0.0734167
R6091 VDDA.n1316 VDDA.n1315 0.0734167
R6092 VDDA.n1317 VDDA.n1316 0.0734167
R6093 VDDA.n1317 VDDA.n461 0.0734167
R6094 VDDA.n539 VDDA.n538 0.0734167
R6095 VDDA.n539 VDDA.n531 0.0734167
R6096 VDDA.n547 VDDA.n527 0.0734167
R6097 VDDA.n553 VDDA.n527 0.0734167
R6098 VDDA.n554 VDDA.n553 0.0734167
R6099 VDDA.n562 VDDA.n561 0.0734167
R6100 VDDA.n563 VDDA.n562 0.0734167
R6101 VDDA.n563 VDDA.n519 0.0734167
R6102 VDDA.n571 VDDA.n515 0.0734167
R6103 VDDA.n577 VDDA.n515 0.0734167
R6104 VDDA.n578 VDDA.n577 0.0734167
R6105 VDDA.n586 VDDA.n585 0.0734167
R6106 VDDA.n587 VDDA.n586 0.0734167
R6107 VDDA.n587 VDDA.n507 0.0734167
R6108 VDDA.n595 VDDA.n503 0.0734167
R6109 VDDA.n601 VDDA.n503 0.0734167
R6110 VDDA.n602 VDDA.n601 0.0734167
R6111 VDDA.n610 VDDA.n609 0.0734167
R6112 VDDA.n611 VDDA.n610 0.0734167
R6113 VDDA.n611 VDDA.n495 0.0734167
R6114 VDDA.n619 VDDA.n491 0.0734167
R6115 VDDA.n625 VDDA.n491 0.0734167
R6116 VDDA.n626 VDDA.n625 0.0734167
R6117 VDDA.n1038 VDDA.n1027 0.0734167
R6118 VDDA.n1039 VDDA.n1038 0.0734167
R6119 VDDA.n1049 VDDA.n1048 0.0734167
R6120 VDDA.n1050 VDDA.n1049 0.0734167
R6121 VDDA.n1050 VDDA.n1019 0.0734167
R6122 VDDA.n1060 VDDA.n1015 0.0734167
R6123 VDDA.n1068 VDDA.n1015 0.0734167
R6124 VDDA.n1069 VDDA.n1068 0.0734167
R6125 VDDA.n1079 VDDA.n1078 0.0734167
R6126 VDDA.n1080 VDDA.n1079 0.0734167
R6127 VDDA.n1080 VDDA.n1007 0.0734167
R6128 VDDA.n1090 VDDA.n1003 0.0734167
R6129 VDDA.n1098 VDDA.n1003 0.0734167
R6130 VDDA.n1099 VDDA.n1098 0.0734167
R6131 VDDA.n1109 VDDA.n1108 0.0734167
R6132 VDDA.n1110 VDDA.n1109 0.0734167
R6133 VDDA.n1110 VDDA.n995 0.0734167
R6134 VDDA.n1120 VDDA.n991 0.0734167
R6135 VDDA.n1128 VDDA.n991 0.0734167
R6136 VDDA.n1129 VDDA.n1128 0.0734167
R6137 VDDA.n1139 VDDA.n1138 0.0734167
R6138 VDDA.n1140 VDDA.n1139 0.0734167
R6139 VDDA.n1140 VDDA.n983 0.0734167
R6140 VDDA.n887 VDDA.n879 0.0734167
R6141 VDDA.n888 VDDA.n887 0.0734167
R6142 VDDA.n896 VDDA.n895 0.0734167
R6143 VDDA.n897 VDDA.n896 0.0734167
R6144 VDDA.n897 VDDA.n871 0.0734167
R6145 VDDA.n905 VDDA.n867 0.0734167
R6146 VDDA.n911 VDDA.n867 0.0734167
R6147 VDDA.n912 VDDA.n911 0.0734167
R6148 VDDA.n920 VDDA.n919 0.0734167
R6149 VDDA.n921 VDDA.n920 0.0734167
R6150 VDDA.n921 VDDA.n859 0.0734167
R6151 VDDA.n929 VDDA.n855 0.0734167
R6152 VDDA.n935 VDDA.n855 0.0734167
R6153 VDDA.n936 VDDA.n935 0.0734167
R6154 VDDA.n944 VDDA.n943 0.0734167
R6155 VDDA.n945 VDDA.n944 0.0734167
R6156 VDDA.n945 VDDA.n847 0.0734167
R6157 VDDA.n953 VDDA.n843 0.0734167
R6158 VDDA.n959 VDDA.n843 0.0734167
R6159 VDDA.n960 VDDA.n959 0.0734167
R6160 VDDA.n968 VDDA.n967 0.0734167
R6161 VDDA.n969 VDDA.n968 0.0734167
R6162 VDDA.n969 VDDA.n638 0.0734167
R6163 VDDA.n693 VDDA.n692 0.0734167
R6164 VDDA.n693 VDDA.n687 0.0734167
R6165 VDDA.n703 VDDA.n685 0.0734167
R6166 VDDA.n711 VDDA.n685 0.0734167
R6167 VDDA.n712 VDDA.n711 0.0734167
R6168 VDDA.n722 VDDA.n721 0.0734167
R6169 VDDA.n723 VDDA.n722 0.0734167
R6170 VDDA.n723 VDDA.n681 0.0734167
R6171 VDDA.n733 VDDA.n679 0.0734167
R6172 VDDA.n741 VDDA.n679 0.0734167
R6173 VDDA.n742 VDDA.n741 0.0734167
R6174 VDDA.n752 VDDA.n751 0.0734167
R6175 VDDA.n753 VDDA.n752 0.0734167
R6176 VDDA.n753 VDDA.n675 0.0734167
R6177 VDDA.n763 VDDA.n673 0.0734167
R6178 VDDA.n771 VDDA.n673 0.0734167
R6179 VDDA.n772 VDDA.n771 0.0734167
R6180 VDDA.n782 VDDA.n781 0.0734167
R6181 VDDA.n783 VDDA.n782 0.0734167
R6182 VDDA.n783 VDDA.n669 0.0734167
R6183 VDDA.n793 VDDA.n667 0.0734167
R6184 VDDA.n801 VDDA.n667 0.0734167
R6185 VDDA.n802 VDDA.n801 0.0734167
R6186 VDDA.n1906 VDDA.n1370 0.0725159
R6187 VDDA.n1763 VDDA.n1405 0.0711522
R6188 VDDA.n1755 VDDA.n1584 0.0711522
R6189 VDDA.n1751 VDDA.n1587 0.0711522
R6190 VDDA.n1741 VDDA.n1593 0.0711522
R6191 VDDA.n1735 VDDA.n1597 0.0711522
R6192 VDDA.n1725 VDDA.n1603 0.0711522
R6193 VDDA.n1721 VDDA.n1605 0.0711522
R6194 VDDA.n1711 VDDA.n1611 0.0711522
R6195 VDDA.n1705 VDDA.n1615 0.0711522
R6196 VDDA.n1695 VDDA.n1621 0.0711522
R6197 VDDA.n1691 VDDA.n1623 0.0711522
R6198 VDDA.n1681 VDDA.n1629 0.0711522
R6199 VDDA.n1675 VDDA.n1633 0.0711522
R6200 VDDA.n1665 VDDA.n1639 0.0711522
R6201 VDDA.n1661 VDDA.n1641 0.0711522
R6202 VDDA.n1765 VDDA.n1764 0.0711522
R6203 VDDA.n1754 VDDA.n1753 0.0711522
R6204 VDDA.n1752 VDDA.n1586 0.0711522
R6205 VDDA.n1742 VDDA.n1592 0.0711522
R6206 VDDA.n1734 VDDA.n1733 0.0711522
R6207 VDDA.n1724 VDDA.n1723 0.0711522
R6208 VDDA.n1722 VDDA.n1604 0.0711522
R6209 VDDA.n1712 VDDA.n1610 0.0711522
R6210 VDDA.n1704 VDDA.n1703 0.0711522
R6211 VDDA.n1694 VDDA.n1693 0.0711522
R6212 VDDA.n1692 VDDA.n1622 0.0711522
R6213 VDDA.n1682 VDDA.n1628 0.0711522
R6214 VDDA.n1674 VDDA.n1673 0.0711522
R6215 VDDA.n1664 VDDA.n1663 0.0711522
R6216 VDDA.n1662 VDDA.n1640 0.0711522
R6217 VDDA.n1467 VDDA.n1463 0.0682083
R6218 VDDA.n1477 VDDA.n1456 0.0682083
R6219 VDDA.n1479 VDDA.n1478 0.0682083
R6220 VDDA.n1489 VDDA.n1488 0.0682083
R6221 VDDA.n1497 VDDA.n1452 0.0682083
R6222 VDDA.n1507 VDDA.n1450 0.0682083
R6223 VDDA.n1509 VDDA.n1508 0.0682083
R6224 VDDA.n1519 VDDA.n1518 0.0682083
R6225 VDDA.n1527 VDDA.n1446 0.0682083
R6226 VDDA.n1537 VDDA.n1444 0.0682083
R6227 VDDA.n1539 VDDA.n1538 0.0682083
R6228 VDDA.n1549 VDDA.n1548 0.0682083
R6229 VDDA.n1557 VDDA.n1440 0.0682083
R6230 VDDA.n1567 VDDA.n1438 0.0682083
R6231 VDDA.n1569 VDDA.n1568 0.0682083
R6232 VDDA.n2129 VDDA.n2128 0.0682083
R6233 VDDA.n2124 VDDA.n2123 0.0682083
R6234 VDDA.n2154 VDDA.n1931 0.0682083
R6235 VDDA.n2156 VDDA.n2155 0.0682083
R6236 VDDA.n2166 VDDA.n2165 0.0682083
R6237 VDDA.n2174 VDDA.n1927 0.0682083
R6238 VDDA.n2184 VDDA.n1925 0.0682083
R6239 VDDA.n2186 VDDA.n2185 0.0682083
R6240 VDDA.n2196 VDDA.n2195 0.0682083
R6241 VDDA.n2204 VDDA.n1921 0.0682083
R6242 VDDA.n2214 VDDA.n1919 0.0682083
R6243 VDDA.n2216 VDDA.n2215 0.0682083
R6244 VDDA.n2226 VDDA.n2225 0.0682083
R6245 VDDA.n2234 VDDA.n1915 0.0682083
R6246 VDDA.n2244 VDDA.n1913 0.0682083
R6247 VDDA.n2246 VDDA.n2245 0.0682083
R6248 VDDA.n100 VDDA.n86 0.0682083
R6249 VDDA.n102 VDDA.n101 0.0682083
R6250 VDDA.n110 VDDA.n109 0.0682083
R6251 VDDA.n116 VDDA.n78 0.0682083
R6252 VDDA.n124 VDDA.n74 0.0682083
R6253 VDDA.n126 VDDA.n125 0.0682083
R6254 VDDA.n134 VDDA.n133 0.0682083
R6255 VDDA.n140 VDDA.n66 0.0682083
R6256 VDDA.n148 VDDA.n62 0.0682083
R6257 VDDA.n150 VDDA.n149 0.0682083
R6258 VDDA.n158 VDDA.n157 0.0682083
R6259 VDDA.n164 VDDA.n54 0.0682083
R6260 VDDA.n172 VDDA.n50 0.0682083
R6261 VDDA.n174 VDDA.n173 0.0682083
R6262 VDDA.n2944 VDDA.n181 0.0682083
R6263 VDDA.n2826 VDDA.n2825 0.0682083
R6264 VDDA.n2834 VDDA.n2809 0.0682083
R6265 VDDA.n2844 VDDA.n2805 0.0682083
R6266 VDDA.n2846 VDDA.n2845 0.0682083
R6267 VDDA.n2856 VDDA.n2855 0.0682083
R6268 VDDA.n2864 VDDA.n2797 0.0682083
R6269 VDDA.n2874 VDDA.n2793 0.0682083
R6270 VDDA.n2876 VDDA.n2875 0.0682083
R6271 VDDA.n2886 VDDA.n2885 0.0682083
R6272 VDDA.n2894 VDDA.n2785 0.0682083
R6273 VDDA.n2904 VDDA.n2781 0.0682083
R6274 VDDA.n2906 VDDA.n2905 0.0682083
R6275 VDDA.n2916 VDDA.n2915 0.0682083
R6276 VDDA.n2924 VDDA.n2773 0.0682083
R6277 VDDA.n2933 VDDA.n2769 0.0682083
R6278 VDDA.n2675 VDDA.n2674 0.0682083
R6279 VDDA.n2681 VDDA.n2661 0.0682083
R6280 VDDA.n2689 VDDA.n2657 0.0682083
R6281 VDDA.n2691 VDDA.n2690 0.0682083
R6282 VDDA.n2699 VDDA.n2698 0.0682083
R6283 VDDA.n2705 VDDA.n2649 0.0682083
R6284 VDDA.n2713 VDDA.n2645 0.0682083
R6285 VDDA.n2715 VDDA.n2714 0.0682083
R6286 VDDA.n2723 VDDA.n2722 0.0682083
R6287 VDDA.n2729 VDDA.n2637 0.0682083
R6288 VDDA.n2737 VDDA.n2633 0.0682083
R6289 VDDA.n2739 VDDA.n2738 0.0682083
R6290 VDDA.n2747 VDDA.n2746 0.0682083
R6291 VDDA.n2753 VDDA.n2625 0.0682083
R6292 VDDA.n2762 VDDA.n194 0.0682083
R6293 VDDA.n278 VDDA.n264 0.0682083
R6294 VDDA.n280 VDDA.n279 0.0682083
R6295 VDDA.n288 VDDA.n287 0.0682083
R6296 VDDA.n294 VDDA.n256 0.0682083
R6297 VDDA.n302 VDDA.n252 0.0682083
R6298 VDDA.n304 VDDA.n303 0.0682083
R6299 VDDA.n312 VDDA.n311 0.0682083
R6300 VDDA.n318 VDDA.n244 0.0682083
R6301 VDDA.n326 VDDA.n240 0.0682083
R6302 VDDA.n328 VDDA.n327 0.0682083
R6303 VDDA.n336 VDDA.n335 0.0682083
R6304 VDDA.n342 VDDA.n232 0.0682083
R6305 VDDA.n350 VDDA.n228 0.0682083
R6306 VDDA.n352 VDDA.n351 0.0682083
R6307 VDDA.n2596 VDDA.n359 0.0682083
R6308 VDDA.n2478 VDDA.n2477 0.0682083
R6309 VDDA.n2486 VDDA.n2461 0.0682083
R6310 VDDA.n2496 VDDA.n2457 0.0682083
R6311 VDDA.n2498 VDDA.n2497 0.0682083
R6312 VDDA.n2508 VDDA.n2507 0.0682083
R6313 VDDA.n2516 VDDA.n2449 0.0682083
R6314 VDDA.n2526 VDDA.n2445 0.0682083
R6315 VDDA.n2528 VDDA.n2527 0.0682083
R6316 VDDA.n2538 VDDA.n2537 0.0682083
R6317 VDDA.n2546 VDDA.n2437 0.0682083
R6318 VDDA.n2556 VDDA.n2433 0.0682083
R6319 VDDA.n2558 VDDA.n2557 0.0682083
R6320 VDDA.n2568 VDDA.n2567 0.0682083
R6321 VDDA.n2576 VDDA.n2425 0.0682083
R6322 VDDA.n2585 VDDA.n2421 0.0682083
R6323 VDDA.n1237 VDDA.n1236 0.0682083
R6324 VDDA.n1243 VDDA.n1223 0.0682083
R6325 VDDA.n1251 VDDA.n1219 0.0682083
R6326 VDDA.n1253 VDDA.n1252 0.0682083
R6327 VDDA.n1261 VDDA.n1260 0.0682083
R6328 VDDA.n1267 VDDA.n1211 0.0682083
R6329 VDDA.n1275 VDDA.n1207 0.0682083
R6330 VDDA.n1277 VDDA.n1276 0.0682083
R6331 VDDA.n1285 VDDA.n1284 0.0682083
R6332 VDDA.n1291 VDDA.n1199 0.0682083
R6333 VDDA.n1299 VDDA.n1195 0.0682083
R6334 VDDA.n1301 VDDA.n1300 0.0682083
R6335 VDDA.n1309 VDDA.n1308 0.0682083
R6336 VDDA.n1315 VDDA.n1187 0.0682083
R6337 VDDA.n2261 VDDA.n461 0.0682083
R6338 VDDA.n545 VDDA.n531 0.0682083
R6339 VDDA.n547 VDDA.n546 0.0682083
R6340 VDDA.n555 VDDA.n554 0.0682083
R6341 VDDA.n561 VDDA.n523 0.0682083
R6342 VDDA.n569 VDDA.n519 0.0682083
R6343 VDDA.n571 VDDA.n570 0.0682083
R6344 VDDA.n579 VDDA.n578 0.0682083
R6345 VDDA.n585 VDDA.n511 0.0682083
R6346 VDDA.n593 VDDA.n507 0.0682083
R6347 VDDA.n595 VDDA.n594 0.0682083
R6348 VDDA.n603 VDDA.n602 0.0682083
R6349 VDDA.n609 VDDA.n499 0.0682083
R6350 VDDA.n617 VDDA.n495 0.0682083
R6351 VDDA.n619 VDDA.n618 0.0682083
R6352 VDDA.n1158 VDDA.n626 0.0682083
R6353 VDDA.n1040 VDDA.n1039 0.0682083
R6354 VDDA.n1048 VDDA.n1023 0.0682083
R6355 VDDA.n1058 VDDA.n1019 0.0682083
R6356 VDDA.n1060 VDDA.n1059 0.0682083
R6357 VDDA.n1070 VDDA.n1069 0.0682083
R6358 VDDA.n1078 VDDA.n1011 0.0682083
R6359 VDDA.n1088 VDDA.n1007 0.0682083
R6360 VDDA.n1090 VDDA.n1089 0.0682083
R6361 VDDA.n1100 VDDA.n1099 0.0682083
R6362 VDDA.n1108 VDDA.n999 0.0682083
R6363 VDDA.n1118 VDDA.n995 0.0682083
R6364 VDDA.n1120 VDDA.n1119 0.0682083
R6365 VDDA.n1130 VDDA.n1129 0.0682083
R6366 VDDA.n1138 VDDA.n987 0.0682083
R6367 VDDA.n1147 VDDA.n983 0.0682083
R6368 VDDA.n889 VDDA.n888 0.0682083
R6369 VDDA.n895 VDDA.n875 0.0682083
R6370 VDDA.n903 VDDA.n871 0.0682083
R6371 VDDA.n905 VDDA.n904 0.0682083
R6372 VDDA.n913 VDDA.n912 0.0682083
R6373 VDDA.n919 VDDA.n863 0.0682083
R6374 VDDA.n927 VDDA.n859 0.0682083
R6375 VDDA.n929 VDDA.n928 0.0682083
R6376 VDDA.n937 VDDA.n936 0.0682083
R6377 VDDA.n943 VDDA.n851 0.0682083
R6378 VDDA.n951 VDDA.n847 0.0682083
R6379 VDDA.n953 VDDA.n952 0.0682083
R6380 VDDA.n961 VDDA.n960 0.0682083
R6381 VDDA.n967 VDDA.n839 0.0682083
R6382 VDDA.n976 VDDA.n638 0.0682083
R6383 VDDA.n701 VDDA.n687 0.0682083
R6384 VDDA.n703 VDDA.n702 0.0682083
R6385 VDDA.n713 VDDA.n712 0.0682083
R6386 VDDA.n721 VDDA.n683 0.0682083
R6387 VDDA.n731 VDDA.n681 0.0682083
R6388 VDDA.n733 VDDA.n732 0.0682083
R6389 VDDA.n743 VDDA.n742 0.0682083
R6390 VDDA.n751 VDDA.n677 0.0682083
R6391 VDDA.n761 VDDA.n675 0.0682083
R6392 VDDA.n763 VDDA.n762 0.0682083
R6393 VDDA.n773 VDDA.n772 0.0682083
R6394 VDDA.n781 VDDA.n671 0.0682083
R6395 VDDA.n791 VDDA.n669 0.0682083
R6396 VDDA.n793 VDDA.n792 0.0682083
R6397 VDDA.n810 VDDA.n802 0.0682083
R6398 VDDA.n92 VDDA.n91 0.0672139
R6399 VDDA.n2817 VDDA.n2816 0.0672139
R6400 VDDA.n2668 VDDA.n2666 0.0672139
R6401 VDDA.n270 VDDA.n269 0.0672139
R6402 VDDA.n2469 VDDA.n2468 0.0672139
R6403 VDDA.n1230 VDDA.n1228 0.0672139
R6404 VDDA.n537 VDDA.n536 0.0672139
R6405 VDDA.n1031 VDDA.n1030 0.0672139
R6406 VDDA.n882 VDDA.n880 0.0672139
R6407 VDDA.n1578 VDDA.n1435 0.0672139
R6408 VDDA.n2255 VDDA.n1910 0.0672139
R6409 VDDA.n691 VDDA.n690 0.0672139
R6410 VDDA.n1751 VDDA.n1584 0.0657174
R6411 VDDA.n1735 VDDA.n1593 0.0657174
R6412 VDDA.n1721 VDDA.n1603 0.0657174
R6413 VDDA.n1705 VDDA.n1611 0.0657174
R6414 VDDA.n1691 VDDA.n1621 0.0657174
R6415 VDDA.n1675 VDDA.n1629 0.0657174
R6416 VDDA.n1661 VDDA.n1639 0.0657174
R6417 VDDA.n1753 VDDA.n1752 0.0657174
R6418 VDDA.n1734 VDDA.n1592 0.0657174
R6419 VDDA.n1723 VDDA.n1722 0.0657174
R6420 VDDA.n1704 VDDA.n1610 0.0657174
R6421 VDDA.n1693 VDDA.n1692 0.0657174
R6422 VDDA.n1674 VDDA.n1628 0.0657174
R6423 VDDA.n1663 VDDA.n1662 0.0657174
R6424 VDDA.n1478 VDDA.n1477 0.063
R6425 VDDA.n1489 VDDA.n1452 0.063
R6426 VDDA.n1508 VDDA.n1507 0.063
R6427 VDDA.n1519 VDDA.n1446 0.063
R6428 VDDA.n1538 VDDA.n1537 0.063
R6429 VDDA.n1549 VDDA.n1440 0.063
R6430 VDDA.n1568 VDDA.n1567 0.063
R6431 VDDA.n2155 VDDA.n2154 0.063
R6432 VDDA.n2166 VDDA.n1927 0.063
R6433 VDDA.n2185 VDDA.n2184 0.063
R6434 VDDA.n2196 VDDA.n1921 0.063
R6435 VDDA.n2215 VDDA.n2214 0.063
R6436 VDDA.n2226 VDDA.n1915 0.063
R6437 VDDA.n2245 VDDA.n2244 0.063
R6438 VDDA.n101 VDDA.n100 0.063
R6439 VDDA.n110 VDDA.n78 0.063
R6440 VDDA.n125 VDDA.n124 0.063
R6441 VDDA.n134 VDDA.n66 0.063
R6442 VDDA.n149 VDDA.n148 0.063
R6443 VDDA.n158 VDDA.n54 0.063
R6444 VDDA.n173 VDDA.n172 0.063
R6445 VDDA.n2826 VDDA.n2809 0.063
R6446 VDDA.n2845 VDDA.n2844 0.063
R6447 VDDA.n2856 VDDA.n2797 0.063
R6448 VDDA.n2875 VDDA.n2874 0.063
R6449 VDDA.n2886 VDDA.n2785 0.063
R6450 VDDA.n2905 VDDA.n2904 0.063
R6451 VDDA.n2916 VDDA.n2773 0.063
R6452 VDDA.n2675 VDDA.n2661 0.063
R6453 VDDA.n2690 VDDA.n2689 0.063
R6454 VDDA.n2699 VDDA.n2649 0.063
R6455 VDDA.n2714 VDDA.n2713 0.063
R6456 VDDA.n2723 VDDA.n2637 0.063
R6457 VDDA.n2738 VDDA.n2737 0.063
R6458 VDDA.n2747 VDDA.n2625 0.063
R6459 VDDA.n279 VDDA.n278 0.063
R6460 VDDA.n288 VDDA.n256 0.063
R6461 VDDA.n303 VDDA.n302 0.063
R6462 VDDA.n312 VDDA.n244 0.063
R6463 VDDA.n327 VDDA.n326 0.063
R6464 VDDA.n336 VDDA.n232 0.063
R6465 VDDA.n351 VDDA.n350 0.063
R6466 VDDA.n2478 VDDA.n2461 0.063
R6467 VDDA.n2497 VDDA.n2496 0.063
R6468 VDDA.n2508 VDDA.n2449 0.063
R6469 VDDA.n2527 VDDA.n2526 0.063
R6470 VDDA.n2538 VDDA.n2437 0.063
R6471 VDDA.n2557 VDDA.n2556 0.063
R6472 VDDA.n2568 VDDA.n2425 0.063
R6473 VDDA.n1237 VDDA.n1223 0.063
R6474 VDDA.n1252 VDDA.n1251 0.063
R6475 VDDA.n1261 VDDA.n1211 0.063
R6476 VDDA.n1276 VDDA.n1275 0.063
R6477 VDDA.n1285 VDDA.n1199 0.063
R6478 VDDA.n1300 VDDA.n1299 0.063
R6479 VDDA.n1309 VDDA.n1187 0.063
R6480 VDDA.n546 VDDA.n545 0.063
R6481 VDDA.n555 VDDA.n523 0.063
R6482 VDDA.n570 VDDA.n569 0.063
R6483 VDDA.n579 VDDA.n511 0.063
R6484 VDDA.n594 VDDA.n593 0.063
R6485 VDDA.n603 VDDA.n499 0.063
R6486 VDDA.n618 VDDA.n617 0.063
R6487 VDDA.n1040 VDDA.n1023 0.063
R6488 VDDA.n1059 VDDA.n1058 0.063
R6489 VDDA.n1070 VDDA.n1011 0.063
R6490 VDDA.n1089 VDDA.n1088 0.063
R6491 VDDA.n1100 VDDA.n999 0.063
R6492 VDDA.n1119 VDDA.n1118 0.063
R6493 VDDA.n1130 VDDA.n987 0.063
R6494 VDDA.n889 VDDA.n875 0.063
R6495 VDDA.n904 VDDA.n903 0.063
R6496 VDDA.n913 VDDA.n863 0.063
R6497 VDDA.n928 VDDA.n927 0.063
R6498 VDDA.n937 VDDA.n851 0.063
R6499 VDDA.n952 VDDA.n951 0.063
R6500 VDDA.n961 VDDA.n839 0.063
R6501 VDDA.n702 VDDA.n701 0.063
R6502 VDDA.n713 VDDA.n683 0.063
R6503 VDDA.n732 VDDA.n731 0.063
R6504 VDDA.n743 VDDA.n677 0.063
R6505 VDDA.n762 VDDA.n761 0.063
R6506 VDDA.n773 VDDA.n671 0.063
R6507 VDDA.n792 VDDA.n791 0.063
R6508 VDDA.n1799 VDDA.n1798 0.0603182
R6509 VDDA.n1813 VDDA.n1812 0.0603182
R6510 VDDA.n1829 VDDA.n1828 0.0603182
R6511 VDDA.n1843 VDDA.n1842 0.0603182
R6512 VDDA.n1859 VDDA.n1858 0.0603182
R6513 VDDA.n1873 VDDA.n1872 0.0603182
R6514 VDDA.n1889 VDDA.n1888 0.0603182
R6515 VDDA.n1903 VDDA.n1902 0.0603182
R6516 VDDA.n1793 VDDA.n1344 0.0560455
R6517 VDDA.n1803 VDDA.n1802 0.0560455
R6518 VDDA.n1809 VDDA.n1808 0.0560455
R6519 VDDA.n1819 VDDA.n1818 0.0560455
R6520 VDDA.n1823 VDDA.n1822 0.0560455
R6521 VDDA.n1833 VDDA.n1832 0.0560455
R6522 VDDA.n1839 VDDA.n1838 0.0560455
R6523 VDDA.n1849 VDDA.n1848 0.0560455
R6524 VDDA.n1853 VDDA.n1852 0.0560455
R6525 VDDA.n1863 VDDA.n1862 0.0560455
R6526 VDDA.n1869 VDDA.n1868 0.0560455
R6527 VDDA.n1879 VDDA.n1878 0.0560455
R6528 VDDA.n1883 VDDA.n1882 0.0560455
R6529 VDDA.n1893 VDDA.n1892 0.0560455
R6530 VDDA.n1899 VDDA.n1898 0.0560455
R6531 VDDA.n1907 VDDA.n1369 0.0560455
R6532 VDDA.n1471 VDDA.n1470 0.0553333
R6533 VDDA.n1485 VDDA.n1484 0.0553333
R6534 VDDA.n1501 VDDA.n1500 0.0553333
R6535 VDDA.n1515 VDDA.n1514 0.0553333
R6536 VDDA.n1531 VDDA.n1530 0.0553333
R6537 VDDA.n1545 VDDA.n1544 0.0553333
R6538 VDDA.n1561 VDDA.n1560 0.0553333
R6539 VDDA.n1575 VDDA.n1574 0.0553333
R6540 VDDA.n2148 VDDA.n2147 0.0553333
R6541 VDDA.n2162 VDDA.n2161 0.0553333
R6542 VDDA.n2178 VDDA.n2177 0.0553333
R6543 VDDA.n2192 VDDA.n2191 0.0553333
R6544 VDDA.n2208 VDDA.n2207 0.0553333
R6545 VDDA.n2222 VDDA.n2221 0.0553333
R6546 VDDA.n2238 VDDA.n2237 0.0553333
R6547 VDDA.n2252 VDDA.n2251 0.0553333
R6548 VDDA.n89 VDDA.n88 0.0553333
R6549 VDDA.n106 VDDA.n105 0.0553333
R6550 VDDA.n77 VDDA.n76 0.0553333
R6551 VDDA.n130 VDDA.n129 0.0553333
R6552 VDDA.n65 VDDA.n64 0.0553333
R6553 VDDA.n154 VDDA.n153 0.0553333
R6554 VDDA.n53 VDDA.n52 0.0553333
R6555 VDDA.n178 VDDA.n177 0.0553333
R6556 VDDA.n2822 VDDA.n2820 0.0553333
R6557 VDDA.n2838 VDDA.n2807 0.0553333
R6558 VDDA.n2852 VDDA.n2850 0.0553333
R6559 VDDA.n2868 VDDA.n2795 0.0553333
R6560 VDDA.n2882 VDDA.n2880 0.0553333
R6561 VDDA.n2898 VDDA.n2783 0.0553333
R6562 VDDA.n2912 VDDA.n2910 0.0553333
R6563 VDDA.n2928 VDDA.n2771 0.0553333
R6564 VDDA.n2671 VDDA.n2670 0.0553333
R6565 VDDA.n2660 VDDA.n2659 0.0553333
R6566 VDDA.n2695 VDDA.n2694 0.0553333
R6567 VDDA.n2648 VDDA.n2647 0.0553333
R6568 VDDA.n2719 VDDA.n2718 0.0553333
R6569 VDDA.n2636 VDDA.n2635 0.0553333
R6570 VDDA.n2743 VDDA.n2742 0.0553333
R6571 VDDA.n2757 VDDA.n2623 0.0553333
R6572 VDDA.n267 VDDA.n266 0.0553333
R6573 VDDA.n284 VDDA.n283 0.0553333
R6574 VDDA.n255 VDDA.n254 0.0553333
R6575 VDDA.n308 VDDA.n307 0.0553333
R6576 VDDA.n243 VDDA.n242 0.0553333
R6577 VDDA.n332 VDDA.n331 0.0553333
R6578 VDDA.n231 VDDA.n230 0.0553333
R6579 VDDA.n356 VDDA.n355 0.0553333
R6580 VDDA.n2474 VDDA.n2472 0.0553333
R6581 VDDA.n2490 VDDA.n2459 0.0553333
R6582 VDDA.n2504 VDDA.n2502 0.0553333
R6583 VDDA.n2520 VDDA.n2447 0.0553333
R6584 VDDA.n2534 VDDA.n2532 0.0553333
R6585 VDDA.n2550 VDDA.n2435 0.0553333
R6586 VDDA.n2564 VDDA.n2562 0.0553333
R6587 VDDA.n2580 VDDA.n2423 0.0553333
R6588 VDDA.n1233 VDDA.n1232 0.0553333
R6589 VDDA.n1222 VDDA.n1221 0.0553333
R6590 VDDA.n1257 VDDA.n1256 0.0553333
R6591 VDDA.n1210 VDDA.n1209 0.0553333
R6592 VDDA.n1281 VDDA.n1280 0.0553333
R6593 VDDA.n1198 VDDA.n1197 0.0553333
R6594 VDDA.n1305 VDDA.n1304 0.0553333
R6595 VDDA.n1319 VDDA.n1185 0.0553333
R6596 VDDA.n534 VDDA.n533 0.0553333
R6597 VDDA.n551 VDDA.n550 0.0553333
R6598 VDDA.n522 VDDA.n521 0.0553333
R6599 VDDA.n575 VDDA.n574 0.0553333
R6600 VDDA.n510 VDDA.n509 0.0553333
R6601 VDDA.n599 VDDA.n598 0.0553333
R6602 VDDA.n498 VDDA.n497 0.0553333
R6603 VDDA.n623 VDDA.n622 0.0553333
R6604 VDDA.n1036 VDDA.n1034 0.0553333
R6605 VDDA.n1052 VDDA.n1021 0.0553333
R6606 VDDA.n1066 VDDA.n1064 0.0553333
R6607 VDDA.n1082 VDDA.n1009 0.0553333
R6608 VDDA.n1096 VDDA.n1094 0.0553333
R6609 VDDA.n1112 VDDA.n997 0.0553333
R6610 VDDA.n1126 VDDA.n1124 0.0553333
R6611 VDDA.n1142 VDDA.n985 0.0553333
R6612 VDDA.n885 VDDA.n884 0.0553333
R6613 VDDA.n874 VDDA.n873 0.0553333
R6614 VDDA.n909 VDDA.n908 0.0553333
R6615 VDDA.n862 VDDA.n861 0.0553333
R6616 VDDA.n933 VDDA.n932 0.0553333
R6617 VDDA.n850 VDDA.n849 0.0553333
R6618 VDDA.n957 VDDA.n956 0.0553333
R6619 VDDA.n971 VDDA.n837 0.0553333
R6620 VDDA.n695 VDDA.n694 0.0553333
R6621 VDDA.n709 VDDA.n708 0.0553333
R6622 VDDA.n725 VDDA.n724 0.0553333
R6623 VDDA.n739 VDDA.n738 0.0553333
R6624 VDDA.n755 VDDA.n754 0.0553333
R6625 VDDA.n769 VDDA.n768 0.0553333
R6626 VDDA.n785 VDDA.n784 0.0553333
R6627 VDDA.n799 VDDA.n798 0.0553333
R6628 VDDA.n1465 VDDA.n1410 0.0514167
R6629 VDDA.n1475 VDDA.n1474 0.0514167
R6630 VDDA.n1481 VDDA.n1480 0.0514167
R6631 VDDA.n1491 VDDA.n1490 0.0514167
R6632 VDDA.n1495 VDDA.n1494 0.0514167
R6633 VDDA.n1505 VDDA.n1504 0.0514167
R6634 VDDA.n1511 VDDA.n1510 0.0514167
R6635 VDDA.n1521 VDDA.n1520 0.0514167
R6636 VDDA.n1525 VDDA.n1524 0.0514167
R6637 VDDA.n1535 VDDA.n1534 0.0514167
R6638 VDDA.n1541 VDDA.n1540 0.0514167
R6639 VDDA.n1551 VDDA.n1550 0.0514167
R6640 VDDA.n1555 VDDA.n1554 0.0514167
R6641 VDDA.n1565 VDDA.n1564 0.0514167
R6642 VDDA.n1571 VDDA.n1570 0.0514167
R6643 VDDA.n1579 VDDA.n1434 0.0514167
R6644 VDDA.n2152 VDDA.n2151 0.0514167
R6645 VDDA.n2158 VDDA.n2157 0.0514167
R6646 VDDA.n2168 VDDA.n2167 0.0514167
R6647 VDDA.n2172 VDDA.n2171 0.0514167
R6648 VDDA.n2182 VDDA.n2181 0.0514167
R6649 VDDA.n2188 VDDA.n2187 0.0514167
R6650 VDDA.n2198 VDDA.n2197 0.0514167
R6651 VDDA.n2202 VDDA.n2201 0.0514167
R6652 VDDA.n2212 VDDA.n2211 0.0514167
R6653 VDDA.n2218 VDDA.n2217 0.0514167
R6654 VDDA.n2228 VDDA.n2227 0.0514167
R6655 VDDA.n2232 VDDA.n2231 0.0514167
R6656 VDDA.n2242 VDDA.n2241 0.0514167
R6657 VDDA.n2248 VDDA.n2247 0.0514167
R6658 VDDA.n2256 VDDA.n1909 0.0514167
R6659 VDDA.n90 VDDA.n20 0.0514167
R6660 VDDA.n98 VDDA.n97 0.0514167
R6661 VDDA.n85 VDDA.n84 0.0514167
R6662 VDDA.n81 VDDA.n80 0.0514167
R6663 VDDA.n114 VDDA.n113 0.0514167
R6664 VDDA.n122 VDDA.n121 0.0514167
R6665 VDDA.n73 VDDA.n72 0.0514167
R6666 VDDA.n69 VDDA.n68 0.0514167
R6667 VDDA.n138 VDDA.n137 0.0514167
R6668 VDDA.n146 VDDA.n145 0.0514167
R6669 VDDA.n61 VDDA.n60 0.0514167
R6670 VDDA.n57 VDDA.n56 0.0514167
R6671 VDDA.n162 VDDA.n161 0.0514167
R6672 VDDA.n170 VDDA.n169 0.0514167
R6673 VDDA.n49 VDDA.n48 0.0514167
R6674 VDDA.n2946 VDDA.n44 0.0514167
R6675 VDDA.n2818 VDDA.n2815 0.0514167
R6676 VDDA.n2828 VDDA.n2811 0.0514167
R6677 VDDA.n2832 VDDA.n2830 0.0514167
R6678 VDDA.n2842 VDDA.n2840 0.0514167
R6679 VDDA.n2848 VDDA.n2803 0.0514167
R6680 VDDA.n2858 VDDA.n2799 0.0514167
R6681 VDDA.n2862 VDDA.n2860 0.0514167
R6682 VDDA.n2872 VDDA.n2870 0.0514167
R6683 VDDA.n2878 VDDA.n2791 0.0514167
R6684 VDDA.n2888 VDDA.n2787 0.0514167
R6685 VDDA.n2892 VDDA.n2890 0.0514167
R6686 VDDA.n2902 VDDA.n2900 0.0514167
R6687 VDDA.n2908 VDDA.n2779 0.0514167
R6688 VDDA.n2918 VDDA.n2775 0.0514167
R6689 VDDA.n2922 VDDA.n2920 0.0514167
R6690 VDDA.n2931 VDDA.n2930 0.0514167
R6691 VDDA.n2667 VDDA.n2600 0.0514167
R6692 VDDA.n2664 VDDA.n2663 0.0514167
R6693 VDDA.n2679 VDDA.n2678 0.0514167
R6694 VDDA.n2687 VDDA.n2686 0.0514167
R6695 VDDA.n2656 VDDA.n2655 0.0514167
R6696 VDDA.n2652 VDDA.n2651 0.0514167
R6697 VDDA.n2703 VDDA.n2702 0.0514167
R6698 VDDA.n2711 VDDA.n2710 0.0514167
R6699 VDDA.n2644 VDDA.n2643 0.0514167
R6700 VDDA.n2640 VDDA.n2639 0.0514167
R6701 VDDA.n2727 VDDA.n2726 0.0514167
R6702 VDDA.n2735 VDDA.n2734 0.0514167
R6703 VDDA.n2632 VDDA.n2631 0.0514167
R6704 VDDA.n2628 VDDA.n2627 0.0514167
R6705 VDDA.n2751 VDDA.n2750 0.0514167
R6706 VDDA.n2760 VDDA.n196 0.0514167
R6707 VDDA.n268 VDDA.n198 0.0514167
R6708 VDDA.n276 VDDA.n275 0.0514167
R6709 VDDA.n263 VDDA.n262 0.0514167
R6710 VDDA.n259 VDDA.n258 0.0514167
R6711 VDDA.n292 VDDA.n291 0.0514167
R6712 VDDA.n300 VDDA.n299 0.0514167
R6713 VDDA.n251 VDDA.n250 0.0514167
R6714 VDDA.n247 VDDA.n246 0.0514167
R6715 VDDA.n316 VDDA.n315 0.0514167
R6716 VDDA.n324 VDDA.n323 0.0514167
R6717 VDDA.n239 VDDA.n238 0.0514167
R6718 VDDA.n235 VDDA.n234 0.0514167
R6719 VDDA.n340 VDDA.n339 0.0514167
R6720 VDDA.n348 VDDA.n347 0.0514167
R6721 VDDA.n227 VDDA.n226 0.0514167
R6722 VDDA.n2598 VDDA.n222 0.0514167
R6723 VDDA.n2470 VDDA.n2467 0.0514167
R6724 VDDA.n2480 VDDA.n2463 0.0514167
R6725 VDDA.n2484 VDDA.n2482 0.0514167
R6726 VDDA.n2494 VDDA.n2492 0.0514167
R6727 VDDA.n2500 VDDA.n2455 0.0514167
R6728 VDDA.n2510 VDDA.n2451 0.0514167
R6729 VDDA.n2514 VDDA.n2512 0.0514167
R6730 VDDA.n2524 VDDA.n2522 0.0514167
R6731 VDDA.n2530 VDDA.n2443 0.0514167
R6732 VDDA.n2540 VDDA.n2439 0.0514167
R6733 VDDA.n2544 VDDA.n2542 0.0514167
R6734 VDDA.n2554 VDDA.n2552 0.0514167
R6735 VDDA.n2560 VDDA.n2431 0.0514167
R6736 VDDA.n2570 VDDA.n2427 0.0514167
R6737 VDDA.n2574 VDDA.n2572 0.0514167
R6738 VDDA.n2583 VDDA.n2582 0.0514167
R6739 VDDA.n1229 VDDA.n1162 0.0514167
R6740 VDDA.n1226 VDDA.n1225 0.0514167
R6741 VDDA.n1241 VDDA.n1240 0.0514167
R6742 VDDA.n1249 VDDA.n1248 0.0514167
R6743 VDDA.n1218 VDDA.n1217 0.0514167
R6744 VDDA.n1214 VDDA.n1213 0.0514167
R6745 VDDA.n1265 VDDA.n1264 0.0514167
R6746 VDDA.n1273 VDDA.n1272 0.0514167
R6747 VDDA.n1206 VDDA.n1205 0.0514167
R6748 VDDA.n1202 VDDA.n1201 0.0514167
R6749 VDDA.n1289 VDDA.n1288 0.0514167
R6750 VDDA.n1297 VDDA.n1296 0.0514167
R6751 VDDA.n1194 VDDA.n1193 0.0514167
R6752 VDDA.n1190 VDDA.n1189 0.0514167
R6753 VDDA.n1313 VDDA.n1312 0.0514167
R6754 VDDA.n2259 VDDA.n463 0.0514167
R6755 VDDA.n535 VDDA.n465 0.0514167
R6756 VDDA.n543 VDDA.n542 0.0514167
R6757 VDDA.n530 VDDA.n529 0.0514167
R6758 VDDA.n526 VDDA.n525 0.0514167
R6759 VDDA.n559 VDDA.n558 0.0514167
R6760 VDDA.n567 VDDA.n566 0.0514167
R6761 VDDA.n518 VDDA.n517 0.0514167
R6762 VDDA.n514 VDDA.n513 0.0514167
R6763 VDDA.n583 VDDA.n582 0.0514167
R6764 VDDA.n591 VDDA.n590 0.0514167
R6765 VDDA.n506 VDDA.n505 0.0514167
R6766 VDDA.n502 VDDA.n501 0.0514167
R6767 VDDA.n607 VDDA.n606 0.0514167
R6768 VDDA.n615 VDDA.n614 0.0514167
R6769 VDDA.n494 VDDA.n493 0.0514167
R6770 VDDA.n1160 VDDA.n489 0.0514167
R6771 VDDA.n1032 VDDA.n1029 0.0514167
R6772 VDDA.n1042 VDDA.n1025 0.0514167
R6773 VDDA.n1046 VDDA.n1044 0.0514167
R6774 VDDA.n1056 VDDA.n1054 0.0514167
R6775 VDDA.n1062 VDDA.n1017 0.0514167
R6776 VDDA.n1072 VDDA.n1013 0.0514167
R6777 VDDA.n1076 VDDA.n1074 0.0514167
R6778 VDDA.n1086 VDDA.n1084 0.0514167
R6779 VDDA.n1092 VDDA.n1005 0.0514167
R6780 VDDA.n1102 VDDA.n1001 0.0514167
R6781 VDDA.n1106 VDDA.n1104 0.0514167
R6782 VDDA.n1116 VDDA.n1114 0.0514167
R6783 VDDA.n1122 VDDA.n993 0.0514167
R6784 VDDA.n1132 VDDA.n989 0.0514167
R6785 VDDA.n1136 VDDA.n1134 0.0514167
R6786 VDDA.n1145 VDDA.n1144 0.0514167
R6787 VDDA.n881 VDDA.n814 0.0514167
R6788 VDDA.n878 VDDA.n877 0.0514167
R6789 VDDA.n893 VDDA.n892 0.0514167
R6790 VDDA.n901 VDDA.n900 0.0514167
R6791 VDDA.n870 VDDA.n869 0.0514167
R6792 VDDA.n866 VDDA.n865 0.0514167
R6793 VDDA.n917 VDDA.n916 0.0514167
R6794 VDDA.n925 VDDA.n924 0.0514167
R6795 VDDA.n858 VDDA.n857 0.0514167
R6796 VDDA.n854 VDDA.n853 0.0514167
R6797 VDDA.n941 VDDA.n940 0.0514167
R6798 VDDA.n949 VDDA.n948 0.0514167
R6799 VDDA.n846 VDDA.n845 0.0514167
R6800 VDDA.n842 VDDA.n841 0.0514167
R6801 VDDA.n965 VDDA.n964 0.0514167
R6802 VDDA.n974 VDDA.n640 0.0514167
R6803 VDDA.n689 VDDA.n641 0.0514167
R6804 VDDA.n699 VDDA.n698 0.0514167
R6805 VDDA.n705 VDDA.n704 0.0514167
R6806 VDDA.n715 VDDA.n714 0.0514167
R6807 VDDA.n719 VDDA.n718 0.0514167
R6808 VDDA.n729 VDDA.n728 0.0514167
R6809 VDDA.n735 VDDA.n734 0.0514167
R6810 VDDA.n745 VDDA.n744 0.0514167
R6811 VDDA.n749 VDDA.n748 0.0514167
R6812 VDDA.n759 VDDA.n758 0.0514167
R6813 VDDA.n765 VDDA.n764 0.0514167
R6814 VDDA.n775 VDDA.n774 0.0514167
R6815 VDDA.n779 VDDA.n778 0.0514167
R6816 VDDA.n789 VDDA.n788 0.0514167
R6817 VDDA.n795 VDDA.n794 0.0514167
R6818 VDDA.n812 VDDA.n665 0.0514167
R6819 VDDA.n2257 VDDA.n1908 0.0497766
R6820 VDDA.n2147 VDDA.n1321 0.0459984
R6821 VDDA.n2396 VDDA.n390 0.0421667
R6822 VDDA.n981 VDDA.n633 0.0421667
R6823 VDDA.n1152 VDDA.n630 0.0421667
R6824 VDDA.n628 VDDA.n459 0.0421667
R6825 VDDA.n2266 VDDA.n456 0.0421667
R6826 VDDA.n2285 VDDA.n452 0.0421667
R6827 VDDA.n2403 VDDA.n368 0.0421667
R6828 VDDA.n2590 VDDA.n363 0.0421667
R6829 VDDA.n361 VDDA.n192 0.0421667
R6830 VDDA.n2767 VDDA.n189 0.0421667
R6831 VDDA.n2938 VDDA.n186 0.0421667
R6832 VDDA.n2941 VDDA.n184 0.0421667
R6833 VDDA.n1652 VDDA.n1651 0.0352506
R6834 VDDA.n1766 VDDA.n1765 0.0331087
R6835 VDDA.n1798 VDDA.n1345 0.030649
R6836 VDDA.n1802 VDDA.n1346 0.030649
R6837 VDDA.n1812 VDDA.n1348 0.030649
R6838 VDDA.n1818 VDDA.n1349 0.030649
R6839 VDDA.n1828 VDDA.n1351 0.030649
R6840 VDDA.n1832 VDDA.n1352 0.030649
R6841 VDDA.n1842 VDDA.n1354 0.030649
R6842 VDDA.n1848 VDDA.n1355 0.030649
R6843 VDDA.n1858 VDDA.n1357 0.030649
R6844 VDDA.n1862 VDDA.n1358 0.030649
R6845 VDDA.n1872 VDDA.n1360 0.030649
R6846 VDDA.n1878 VDDA.n1361 0.030649
R6847 VDDA.n1888 VDDA.n1363 0.030649
R6848 VDDA.n1892 VDDA.n1364 0.030649
R6849 VDDA.n1902 VDDA.n1366 0.030649
R6850 VDDA.n1369 VDDA.n1367 0.030649
R6851 VDDA.n1903 VDDA.n1367 0.030649
R6852 VDDA.n1899 VDDA.n1366 0.030649
R6853 VDDA.n1889 VDDA.n1364 0.030649
R6854 VDDA.n1883 VDDA.n1363 0.030649
R6855 VDDA.n1873 VDDA.n1361 0.030649
R6856 VDDA.n1869 VDDA.n1360 0.030649
R6857 VDDA.n1859 VDDA.n1358 0.030649
R6858 VDDA.n1853 VDDA.n1357 0.030649
R6859 VDDA.n1843 VDDA.n1355 0.030649
R6860 VDDA.n1839 VDDA.n1354 0.030649
R6861 VDDA.n1829 VDDA.n1352 0.030649
R6862 VDDA.n1823 VDDA.n1351 0.030649
R6863 VDDA.n1813 VDDA.n1349 0.030649
R6864 VDDA.n1809 VDDA.n1348 0.030649
R6865 VDDA.n1799 VDDA.n1346 0.030649
R6866 VDDA.n1793 VDDA.n1345 0.030649
R6867 VDDA.n1470 VDDA.n1411 0.028198
R6868 VDDA.n1474 VDDA.n1412 0.028198
R6869 VDDA.n1484 VDDA.n1414 0.028198
R6870 VDDA.n1490 VDDA.n1415 0.028198
R6871 VDDA.n1500 VDDA.n1417 0.028198
R6872 VDDA.n1504 VDDA.n1418 0.028198
R6873 VDDA.n1514 VDDA.n1420 0.028198
R6874 VDDA.n1520 VDDA.n1421 0.028198
R6875 VDDA.n1530 VDDA.n1423 0.028198
R6876 VDDA.n1534 VDDA.n1424 0.028198
R6877 VDDA.n1544 VDDA.n1426 0.028198
R6878 VDDA.n1550 VDDA.n1427 0.028198
R6879 VDDA.n1560 VDDA.n1429 0.028198
R6880 VDDA.n1564 VDDA.n1430 0.028198
R6881 VDDA.n1574 VDDA.n1432 0.028198
R6882 VDDA.n1434 VDDA.n1433 0.028198
R6883 VDDA.n2151 VDDA.n1322 0.028198
R6884 VDDA.n2161 VDDA.n1324 0.028198
R6885 VDDA.n2167 VDDA.n1325 0.028198
R6886 VDDA.n2177 VDDA.n1327 0.028198
R6887 VDDA.n2181 VDDA.n1328 0.028198
R6888 VDDA.n2191 VDDA.n1330 0.028198
R6889 VDDA.n2197 VDDA.n1331 0.028198
R6890 VDDA.n2207 VDDA.n1333 0.028198
R6891 VDDA.n2211 VDDA.n1334 0.028198
R6892 VDDA.n2221 VDDA.n1336 0.028198
R6893 VDDA.n2227 VDDA.n1337 0.028198
R6894 VDDA.n2237 VDDA.n1339 0.028198
R6895 VDDA.n2241 VDDA.n1340 0.028198
R6896 VDDA.n2251 VDDA.n1342 0.028198
R6897 VDDA.n1909 VDDA.n1343 0.028198
R6898 VDDA.n88 VDDA.n21 0.028198
R6899 VDDA.n97 VDDA.n22 0.028198
R6900 VDDA.n105 VDDA.n24 0.028198
R6901 VDDA.n80 VDDA.n25 0.028198
R6902 VDDA.n76 VDDA.n27 0.028198
R6903 VDDA.n121 VDDA.n28 0.028198
R6904 VDDA.n129 VDDA.n30 0.028198
R6905 VDDA.n68 VDDA.n31 0.028198
R6906 VDDA.n64 VDDA.n33 0.028198
R6907 VDDA.n145 VDDA.n34 0.028198
R6908 VDDA.n153 VDDA.n36 0.028198
R6909 VDDA.n56 VDDA.n37 0.028198
R6910 VDDA.n52 VDDA.n39 0.028198
R6911 VDDA.n169 VDDA.n40 0.028198
R6912 VDDA.n177 VDDA.n42 0.028198
R6913 VDDA.n44 VDDA.n43 0.028198
R6914 VDDA.n2820 VDDA.n2819 0.028198
R6915 VDDA.n2821 VDDA.n2811 0.028198
R6916 VDDA.n2831 VDDA.n2807 0.028198
R6917 VDDA.n2840 VDDA.n2839 0.028198
R6918 VDDA.n2850 VDDA.n2849 0.028198
R6919 VDDA.n2851 VDDA.n2799 0.028198
R6920 VDDA.n2861 VDDA.n2795 0.028198
R6921 VDDA.n2870 VDDA.n2869 0.028198
R6922 VDDA.n2880 VDDA.n2879 0.028198
R6923 VDDA.n2881 VDDA.n2787 0.028198
R6924 VDDA.n2891 VDDA.n2783 0.028198
R6925 VDDA.n2900 VDDA.n2899 0.028198
R6926 VDDA.n2910 VDDA.n2909 0.028198
R6927 VDDA.n2911 VDDA.n2775 0.028198
R6928 VDDA.n2921 VDDA.n2771 0.028198
R6929 VDDA.n2930 VDDA.n2929 0.028198
R6930 VDDA.n2670 VDDA.n2601 0.028198
R6931 VDDA.n2663 VDDA.n2602 0.028198
R6932 VDDA.n2659 VDDA.n2604 0.028198
R6933 VDDA.n2686 VDDA.n2605 0.028198
R6934 VDDA.n2694 VDDA.n2607 0.028198
R6935 VDDA.n2651 VDDA.n2608 0.028198
R6936 VDDA.n2647 VDDA.n2610 0.028198
R6937 VDDA.n2710 VDDA.n2611 0.028198
R6938 VDDA.n2718 VDDA.n2613 0.028198
R6939 VDDA.n2639 VDDA.n2614 0.028198
R6940 VDDA.n2635 VDDA.n2616 0.028198
R6941 VDDA.n2734 VDDA.n2617 0.028198
R6942 VDDA.n2742 VDDA.n2619 0.028198
R6943 VDDA.n2627 VDDA.n2620 0.028198
R6944 VDDA.n2623 VDDA.n2622 0.028198
R6945 VDDA.n2758 VDDA.n196 0.028198
R6946 VDDA.n266 VDDA.n199 0.028198
R6947 VDDA.n275 VDDA.n200 0.028198
R6948 VDDA.n283 VDDA.n202 0.028198
R6949 VDDA.n258 VDDA.n203 0.028198
R6950 VDDA.n254 VDDA.n205 0.028198
R6951 VDDA.n299 VDDA.n206 0.028198
R6952 VDDA.n307 VDDA.n208 0.028198
R6953 VDDA.n246 VDDA.n209 0.028198
R6954 VDDA.n242 VDDA.n211 0.028198
R6955 VDDA.n323 VDDA.n212 0.028198
R6956 VDDA.n331 VDDA.n214 0.028198
R6957 VDDA.n234 VDDA.n215 0.028198
R6958 VDDA.n230 VDDA.n217 0.028198
R6959 VDDA.n347 VDDA.n218 0.028198
R6960 VDDA.n355 VDDA.n220 0.028198
R6961 VDDA.n222 VDDA.n221 0.028198
R6962 VDDA.n2472 VDDA.n2471 0.028198
R6963 VDDA.n2473 VDDA.n2463 0.028198
R6964 VDDA.n2483 VDDA.n2459 0.028198
R6965 VDDA.n2492 VDDA.n2491 0.028198
R6966 VDDA.n2502 VDDA.n2501 0.028198
R6967 VDDA.n2503 VDDA.n2451 0.028198
R6968 VDDA.n2513 VDDA.n2447 0.028198
R6969 VDDA.n2522 VDDA.n2521 0.028198
R6970 VDDA.n2532 VDDA.n2531 0.028198
R6971 VDDA.n2533 VDDA.n2439 0.028198
R6972 VDDA.n2543 VDDA.n2435 0.028198
R6973 VDDA.n2552 VDDA.n2551 0.028198
R6974 VDDA.n2562 VDDA.n2561 0.028198
R6975 VDDA.n2563 VDDA.n2427 0.028198
R6976 VDDA.n2573 VDDA.n2423 0.028198
R6977 VDDA.n2582 VDDA.n2581 0.028198
R6978 VDDA.n1232 VDDA.n1163 0.028198
R6979 VDDA.n1225 VDDA.n1164 0.028198
R6980 VDDA.n1221 VDDA.n1166 0.028198
R6981 VDDA.n1248 VDDA.n1167 0.028198
R6982 VDDA.n1256 VDDA.n1169 0.028198
R6983 VDDA.n1213 VDDA.n1170 0.028198
R6984 VDDA.n1209 VDDA.n1172 0.028198
R6985 VDDA.n1272 VDDA.n1173 0.028198
R6986 VDDA.n1280 VDDA.n1175 0.028198
R6987 VDDA.n1201 VDDA.n1176 0.028198
R6988 VDDA.n1197 VDDA.n1178 0.028198
R6989 VDDA.n1296 VDDA.n1179 0.028198
R6990 VDDA.n1304 VDDA.n1181 0.028198
R6991 VDDA.n1189 VDDA.n1182 0.028198
R6992 VDDA.n1185 VDDA.n1184 0.028198
R6993 VDDA.n1320 VDDA.n463 0.028198
R6994 VDDA.n533 VDDA.n466 0.028198
R6995 VDDA.n542 VDDA.n467 0.028198
R6996 VDDA.n550 VDDA.n469 0.028198
R6997 VDDA.n525 VDDA.n470 0.028198
R6998 VDDA.n521 VDDA.n472 0.028198
R6999 VDDA.n566 VDDA.n473 0.028198
R7000 VDDA.n574 VDDA.n475 0.028198
R7001 VDDA.n513 VDDA.n476 0.028198
R7002 VDDA.n509 VDDA.n478 0.028198
R7003 VDDA.n590 VDDA.n479 0.028198
R7004 VDDA.n598 VDDA.n481 0.028198
R7005 VDDA.n501 VDDA.n482 0.028198
R7006 VDDA.n497 VDDA.n484 0.028198
R7007 VDDA.n614 VDDA.n485 0.028198
R7008 VDDA.n622 VDDA.n487 0.028198
R7009 VDDA.n489 VDDA.n488 0.028198
R7010 VDDA.n1034 VDDA.n1033 0.028198
R7011 VDDA.n1035 VDDA.n1025 0.028198
R7012 VDDA.n1045 VDDA.n1021 0.028198
R7013 VDDA.n1054 VDDA.n1053 0.028198
R7014 VDDA.n1064 VDDA.n1063 0.028198
R7015 VDDA.n1065 VDDA.n1013 0.028198
R7016 VDDA.n1075 VDDA.n1009 0.028198
R7017 VDDA.n1084 VDDA.n1083 0.028198
R7018 VDDA.n1094 VDDA.n1093 0.028198
R7019 VDDA.n1095 VDDA.n1001 0.028198
R7020 VDDA.n1105 VDDA.n997 0.028198
R7021 VDDA.n1114 VDDA.n1113 0.028198
R7022 VDDA.n1124 VDDA.n1123 0.028198
R7023 VDDA.n1125 VDDA.n989 0.028198
R7024 VDDA.n1135 VDDA.n985 0.028198
R7025 VDDA.n1144 VDDA.n1143 0.028198
R7026 VDDA.n884 VDDA.n815 0.028198
R7027 VDDA.n877 VDDA.n816 0.028198
R7028 VDDA.n873 VDDA.n818 0.028198
R7029 VDDA.n900 VDDA.n819 0.028198
R7030 VDDA.n908 VDDA.n821 0.028198
R7031 VDDA.n865 VDDA.n822 0.028198
R7032 VDDA.n861 VDDA.n824 0.028198
R7033 VDDA.n924 VDDA.n825 0.028198
R7034 VDDA.n932 VDDA.n827 0.028198
R7035 VDDA.n853 VDDA.n828 0.028198
R7036 VDDA.n849 VDDA.n830 0.028198
R7037 VDDA.n948 VDDA.n831 0.028198
R7038 VDDA.n956 VDDA.n833 0.028198
R7039 VDDA.n841 VDDA.n834 0.028198
R7040 VDDA.n837 VDDA.n836 0.028198
R7041 VDDA.n972 VDDA.n640 0.028198
R7042 VDDA.n694 VDDA.n642 0.028198
R7043 VDDA.n698 VDDA.n643 0.028198
R7044 VDDA.n708 VDDA.n645 0.028198
R7045 VDDA.n714 VDDA.n646 0.028198
R7046 VDDA.n724 VDDA.n648 0.028198
R7047 VDDA.n728 VDDA.n649 0.028198
R7048 VDDA.n738 VDDA.n651 0.028198
R7049 VDDA.n744 VDDA.n652 0.028198
R7050 VDDA.n754 VDDA.n654 0.028198
R7051 VDDA.n758 VDDA.n655 0.028198
R7052 VDDA.n768 VDDA.n657 0.028198
R7053 VDDA.n774 VDDA.n658 0.028198
R7054 VDDA.n784 VDDA.n660 0.028198
R7055 VDDA.n788 VDDA.n661 0.028198
R7056 VDDA.n798 VDDA.n663 0.028198
R7057 VDDA.n665 VDDA.n664 0.028198
R7058 VDDA.n799 VDDA.n664 0.028198
R7059 VDDA.n795 VDDA.n663 0.028198
R7060 VDDA.n785 VDDA.n661 0.028198
R7061 VDDA.n779 VDDA.n660 0.028198
R7062 VDDA.n769 VDDA.n658 0.028198
R7063 VDDA.n765 VDDA.n657 0.028198
R7064 VDDA.n755 VDDA.n655 0.028198
R7065 VDDA.n749 VDDA.n654 0.028198
R7066 VDDA.n739 VDDA.n652 0.028198
R7067 VDDA.n735 VDDA.n651 0.028198
R7068 VDDA.n725 VDDA.n649 0.028198
R7069 VDDA.n719 VDDA.n648 0.028198
R7070 VDDA.n709 VDDA.n646 0.028198
R7071 VDDA.n705 VDDA.n645 0.028198
R7072 VDDA.n695 VDDA.n643 0.028198
R7073 VDDA.n689 VDDA.n642 0.028198
R7074 VDDA.n972 VDDA.n971 0.028198
R7075 VDDA.n965 VDDA.n836 0.028198
R7076 VDDA.n957 VDDA.n834 0.028198
R7077 VDDA.n846 VDDA.n833 0.028198
R7078 VDDA.n850 VDDA.n831 0.028198
R7079 VDDA.n941 VDDA.n830 0.028198
R7080 VDDA.n933 VDDA.n828 0.028198
R7081 VDDA.n858 VDDA.n827 0.028198
R7082 VDDA.n862 VDDA.n825 0.028198
R7083 VDDA.n917 VDDA.n824 0.028198
R7084 VDDA.n909 VDDA.n822 0.028198
R7085 VDDA.n870 VDDA.n821 0.028198
R7086 VDDA.n874 VDDA.n819 0.028198
R7087 VDDA.n893 VDDA.n818 0.028198
R7088 VDDA.n885 VDDA.n816 0.028198
R7089 VDDA.n881 VDDA.n815 0.028198
R7090 VDDA.n1143 VDDA.n1142 0.028198
R7091 VDDA.n1136 VDDA.n1135 0.028198
R7092 VDDA.n1126 VDDA.n1125 0.028198
R7093 VDDA.n1123 VDDA.n1122 0.028198
R7094 VDDA.n1113 VDDA.n1112 0.028198
R7095 VDDA.n1106 VDDA.n1105 0.028198
R7096 VDDA.n1096 VDDA.n1095 0.028198
R7097 VDDA.n1093 VDDA.n1092 0.028198
R7098 VDDA.n1083 VDDA.n1082 0.028198
R7099 VDDA.n1076 VDDA.n1075 0.028198
R7100 VDDA.n1066 VDDA.n1065 0.028198
R7101 VDDA.n1063 VDDA.n1062 0.028198
R7102 VDDA.n1053 VDDA.n1052 0.028198
R7103 VDDA.n1046 VDDA.n1045 0.028198
R7104 VDDA.n1036 VDDA.n1035 0.028198
R7105 VDDA.n1033 VDDA.n1032 0.028198
R7106 VDDA.n623 VDDA.n488 0.028198
R7107 VDDA.n494 VDDA.n487 0.028198
R7108 VDDA.n498 VDDA.n485 0.028198
R7109 VDDA.n607 VDDA.n484 0.028198
R7110 VDDA.n599 VDDA.n482 0.028198
R7111 VDDA.n506 VDDA.n481 0.028198
R7112 VDDA.n510 VDDA.n479 0.028198
R7113 VDDA.n583 VDDA.n478 0.028198
R7114 VDDA.n575 VDDA.n476 0.028198
R7115 VDDA.n518 VDDA.n475 0.028198
R7116 VDDA.n522 VDDA.n473 0.028198
R7117 VDDA.n559 VDDA.n472 0.028198
R7118 VDDA.n551 VDDA.n470 0.028198
R7119 VDDA.n530 VDDA.n469 0.028198
R7120 VDDA.n534 VDDA.n467 0.028198
R7121 VDDA.n535 VDDA.n466 0.028198
R7122 VDDA.n1320 VDDA.n1319 0.028198
R7123 VDDA.n1313 VDDA.n1184 0.028198
R7124 VDDA.n1305 VDDA.n1182 0.028198
R7125 VDDA.n1194 VDDA.n1181 0.028198
R7126 VDDA.n1198 VDDA.n1179 0.028198
R7127 VDDA.n1289 VDDA.n1178 0.028198
R7128 VDDA.n1281 VDDA.n1176 0.028198
R7129 VDDA.n1206 VDDA.n1175 0.028198
R7130 VDDA.n1210 VDDA.n1173 0.028198
R7131 VDDA.n1265 VDDA.n1172 0.028198
R7132 VDDA.n1257 VDDA.n1170 0.028198
R7133 VDDA.n1218 VDDA.n1169 0.028198
R7134 VDDA.n1222 VDDA.n1167 0.028198
R7135 VDDA.n1241 VDDA.n1166 0.028198
R7136 VDDA.n1233 VDDA.n1164 0.028198
R7137 VDDA.n1229 VDDA.n1163 0.028198
R7138 VDDA.n2252 VDDA.n1343 0.028198
R7139 VDDA.n2248 VDDA.n1342 0.028198
R7140 VDDA.n2238 VDDA.n1340 0.028198
R7141 VDDA.n2232 VDDA.n1339 0.028198
R7142 VDDA.n2222 VDDA.n1337 0.028198
R7143 VDDA.n2218 VDDA.n1336 0.028198
R7144 VDDA.n2208 VDDA.n1334 0.028198
R7145 VDDA.n2202 VDDA.n1333 0.028198
R7146 VDDA.n2192 VDDA.n1331 0.028198
R7147 VDDA.n2188 VDDA.n1330 0.028198
R7148 VDDA.n2178 VDDA.n1328 0.028198
R7149 VDDA.n2172 VDDA.n1327 0.028198
R7150 VDDA.n2162 VDDA.n1325 0.028198
R7151 VDDA.n2158 VDDA.n1324 0.028198
R7152 VDDA.n2148 VDDA.n1322 0.028198
R7153 VDDA.n2581 VDDA.n2580 0.028198
R7154 VDDA.n2574 VDDA.n2573 0.028198
R7155 VDDA.n2564 VDDA.n2563 0.028198
R7156 VDDA.n2561 VDDA.n2560 0.028198
R7157 VDDA.n2551 VDDA.n2550 0.028198
R7158 VDDA.n2544 VDDA.n2543 0.028198
R7159 VDDA.n2534 VDDA.n2533 0.028198
R7160 VDDA.n2531 VDDA.n2530 0.028198
R7161 VDDA.n2521 VDDA.n2520 0.028198
R7162 VDDA.n2514 VDDA.n2513 0.028198
R7163 VDDA.n2504 VDDA.n2503 0.028198
R7164 VDDA.n2501 VDDA.n2500 0.028198
R7165 VDDA.n2491 VDDA.n2490 0.028198
R7166 VDDA.n2484 VDDA.n2483 0.028198
R7167 VDDA.n2474 VDDA.n2473 0.028198
R7168 VDDA.n2471 VDDA.n2470 0.028198
R7169 VDDA.n356 VDDA.n221 0.028198
R7170 VDDA.n227 VDDA.n220 0.028198
R7171 VDDA.n231 VDDA.n218 0.028198
R7172 VDDA.n340 VDDA.n217 0.028198
R7173 VDDA.n332 VDDA.n215 0.028198
R7174 VDDA.n239 VDDA.n214 0.028198
R7175 VDDA.n243 VDDA.n212 0.028198
R7176 VDDA.n316 VDDA.n211 0.028198
R7177 VDDA.n308 VDDA.n209 0.028198
R7178 VDDA.n251 VDDA.n208 0.028198
R7179 VDDA.n255 VDDA.n206 0.028198
R7180 VDDA.n292 VDDA.n205 0.028198
R7181 VDDA.n284 VDDA.n203 0.028198
R7182 VDDA.n263 VDDA.n202 0.028198
R7183 VDDA.n267 VDDA.n200 0.028198
R7184 VDDA.n268 VDDA.n199 0.028198
R7185 VDDA.n2758 VDDA.n2757 0.028198
R7186 VDDA.n2751 VDDA.n2622 0.028198
R7187 VDDA.n2743 VDDA.n2620 0.028198
R7188 VDDA.n2632 VDDA.n2619 0.028198
R7189 VDDA.n2636 VDDA.n2617 0.028198
R7190 VDDA.n2727 VDDA.n2616 0.028198
R7191 VDDA.n2719 VDDA.n2614 0.028198
R7192 VDDA.n2644 VDDA.n2613 0.028198
R7193 VDDA.n2648 VDDA.n2611 0.028198
R7194 VDDA.n2703 VDDA.n2610 0.028198
R7195 VDDA.n2695 VDDA.n2608 0.028198
R7196 VDDA.n2656 VDDA.n2607 0.028198
R7197 VDDA.n2660 VDDA.n2605 0.028198
R7198 VDDA.n2679 VDDA.n2604 0.028198
R7199 VDDA.n2671 VDDA.n2602 0.028198
R7200 VDDA.n2667 VDDA.n2601 0.028198
R7201 VDDA.n2929 VDDA.n2928 0.028198
R7202 VDDA.n2922 VDDA.n2921 0.028198
R7203 VDDA.n2912 VDDA.n2911 0.028198
R7204 VDDA.n2909 VDDA.n2908 0.028198
R7205 VDDA.n2899 VDDA.n2898 0.028198
R7206 VDDA.n2892 VDDA.n2891 0.028198
R7207 VDDA.n2882 VDDA.n2881 0.028198
R7208 VDDA.n2879 VDDA.n2878 0.028198
R7209 VDDA.n2869 VDDA.n2868 0.028198
R7210 VDDA.n2862 VDDA.n2861 0.028198
R7211 VDDA.n2852 VDDA.n2851 0.028198
R7212 VDDA.n2849 VDDA.n2848 0.028198
R7213 VDDA.n2839 VDDA.n2838 0.028198
R7214 VDDA.n2832 VDDA.n2831 0.028198
R7215 VDDA.n2822 VDDA.n2821 0.028198
R7216 VDDA.n2819 VDDA.n2818 0.028198
R7217 VDDA.n178 VDDA.n43 0.028198
R7218 VDDA.n49 VDDA.n42 0.028198
R7219 VDDA.n53 VDDA.n40 0.028198
R7220 VDDA.n162 VDDA.n39 0.028198
R7221 VDDA.n154 VDDA.n37 0.028198
R7222 VDDA.n61 VDDA.n36 0.028198
R7223 VDDA.n65 VDDA.n34 0.028198
R7224 VDDA.n138 VDDA.n33 0.028198
R7225 VDDA.n130 VDDA.n31 0.028198
R7226 VDDA.n73 VDDA.n30 0.028198
R7227 VDDA.n77 VDDA.n28 0.028198
R7228 VDDA.n114 VDDA.n27 0.028198
R7229 VDDA.n106 VDDA.n25 0.028198
R7230 VDDA.n85 VDDA.n24 0.028198
R7231 VDDA.n89 VDDA.n22 0.028198
R7232 VDDA.n90 VDDA.n21 0.028198
R7233 VDDA.n1575 VDDA.n1433 0.028198
R7234 VDDA.n1571 VDDA.n1432 0.028198
R7235 VDDA.n1561 VDDA.n1430 0.028198
R7236 VDDA.n1555 VDDA.n1429 0.028198
R7237 VDDA.n1545 VDDA.n1427 0.028198
R7238 VDDA.n1541 VDDA.n1426 0.028198
R7239 VDDA.n1531 VDDA.n1424 0.028198
R7240 VDDA.n1525 VDDA.n1423 0.028198
R7241 VDDA.n1515 VDDA.n1421 0.028198
R7242 VDDA.n1511 VDDA.n1420 0.028198
R7243 VDDA.n1501 VDDA.n1418 0.028198
R7244 VDDA.n1495 VDDA.n1417 0.028198
R7245 VDDA.n1485 VDDA.n1415 0.028198
R7246 VDDA.n1481 VDDA.n1414 0.028198
R7247 VDDA.n1471 VDDA.n1412 0.028198
R7248 VDDA.n1465 VDDA.n1411 0.028198
R7249 VDDA.n1808 VDDA.n1347 0.0264451
R7250 VDDA.n1822 VDDA.n1350 0.0264451
R7251 VDDA.n1838 VDDA.n1353 0.0264451
R7252 VDDA.n1852 VDDA.n1356 0.0264451
R7253 VDDA.n1868 VDDA.n1359 0.0264451
R7254 VDDA.n1882 VDDA.n1362 0.0264451
R7255 VDDA.n1898 VDDA.n1365 0.0264451
R7256 VDDA.n1893 VDDA.n1365 0.0264451
R7257 VDDA.n1879 VDDA.n1362 0.0264451
R7258 VDDA.n1863 VDDA.n1359 0.0264451
R7259 VDDA.n1849 VDDA.n1356 0.0264451
R7260 VDDA.n1833 VDDA.n1353 0.0264451
R7261 VDDA.n1819 VDDA.n1350 0.0264451
R7262 VDDA.n1803 VDDA.n1347 0.0264451
R7263 VDDA.n1480 VDDA.n1413 0.0243392
R7264 VDDA.n1494 VDDA.n1416 0.0243392
R7265 VDDA.n1510 VDDA.n1419 0.0243392
R7266 VDDA.n1524 VDDA.n1422 0.0243392
R7267 VDDA.n1540 VDDA.n1425 0.0243392
R7268 VDDA.n1554 VDDA.n1428 0.0243392
R7269 VDDA.n1570 VDDA.n1431 0.0243392
R7270 VDDA.n2157 VDDA.n1323 0.0243392
R7271 VDDA.n2171 VDDA.n1326 0.0243392
R7272 VDDA.n2187 VDDA.n1329 0.0243392
R7273 VDDA.n2201 VDDA.n1332 0.0243392
R7274 VDDA.n2217 VDDA.n1335 0.0243392
R7275 VDDA.n2231 VDDA.n1338 0.0243392
R7276 VDDA.n2247 VDDA.n1341 0.0243392
R7277 VDDA.n84 VDDA.n23 0.0243392
R7278 VDDA.n113 VDDA.n26 0.0243392
R7279 VDDA.n72 VDDA.n29 0.0243392
R7280 VDDA.n137 VDDA.n32 0.0243392
R7281 VDDA.n60 VDDA.n35 0.0243392
R7282 VDDA.n161 VDDA.n38 0.0243392
R7283 VDDA.n48 VDDA.n41 0.0243392
R7284 VDDA.n2830 VDDA.n2829 0.0243392
R7285 VDDA.n2841 VDDA.n2803 0.0243392
R7286 VDDA.n2860 VDDA.n2859 0.0243392
R7287 VDDA.n2871 VDDA.n2791 0.0243392
R7288 VDDA.n2890 VDDA.n2889 0.0243392
R7289 VDDA.n2901 VDDA.n2779 0.0243392
R7290 VDDA.n2920 VDDA.n2919 0.0243392
R7291 VDDA.n2678 VDDA.n2603 0.0243392
R7292 VDDA.n2655 VDDA.n2606 0.0243392
R7293 VDDA.n2702 VDDA.n2609 0.0243392
R7294 VDDA.n2643 VDDA.n2612 0.0243392
R7295 VDDA.n2726 VDDA.n2615 0.0243392
R7296 VDDA.n2631 VDDA.n2618 0.0243392
R7297 VDDA.n2750 VDDA.n2621 0.0243392
R7298 VDDA.n262 VDDA.n201 0.0243392
R7299 VDDA.n291 VDDA.n204 0.0243392
R7300 VDDA.n250 VDDA.n207 0.0243392
R7301 VDDA.n315 VDDA.n210 0.0243392
R7302 VDDA.n238 VDDA.n213 0.0243392
R7303 VDDA.n339 VDDA.n216 0.0243392
R7304 VDDA.n226 VDDA.n219 0.0243392
R7305 VDDA.n2482 VDDA.n2481 0.0243392
R7306 VDDA.n2493 VDDA.n2455 0.0243392
R7307 VDDA.n2512 VDDA.n2511 0.0243392
R7308 VDDA.n2523 VDDA.n2443 0.0243392
R7309 VDDA.n2542 VDDA.n2541 0.0243392
R7310 VDDA.n2553 VDDA.n2431 0.0243392
R7311 VDDA.n2572 VDDA.n2571 0.0243392
R7312 VDDA.n1240 VDDA.n1165 0.0243392
R7313 VDDA.n1217 VDDA.n1168 0.0243392
R7314 VDDA.n1264 VDDA.n1171 0.0243392
R7315 VDDA.n1205 VDDA.n1174 0.0243392
R7316 VDDA.n1288 VDDA.n1177 0.0243392
R7317 VDDA.n1193 VDDA.n1180 0.0243392
R7318 VDDA.n1312 VDDA.n1183 0.0243392
R7319 VDDA.n529 VDDA.n468 0.0243392
R7320 VDDA.n558 VDDA.n471 0.0243392
R7321 VDDA.n517 VDDA.n474 0.0243392
R7322 VDDA.n582 VDDA.n477 0.0243392
R7323 VDDA.n505 VDDA.n480 0.0243392
R7324 VDDA.n606 VDDA.n483 0.0243392
R7325 VDDA.n493 VDDA.n486 0.0243392
R7326 VDDA.n1044 VDDA.n1043 0.0243392
R7327 VDDA.n1055 VDDA.n1017 0.0243392
R7328 VDDA.n1074 VDDA.n1073 0.0243392
R7329 VDDA.n1085 VDDA.n1005 0.0243392
R7330 VDDA.n1104 VDDA.n1103 0.0243392
R7331 VDDA.n1115 VDDA.n993 0.0243392
R7332 VDDA.n1134 VDDA.n1133 0.0243392
R7333 VDDA.n892 VDDA.n817 0.0243392
R7334 VDDA.n869 VDDA.n820 0.0243392
R7335 VDDA.n916 VDDA.n823 0.0243392
R7336 VDDA.n857 VDDA.n826 0.0243392
R7337 VDDA.n940 VDDA.n829 0.0243392
R7338 VDDA.n845 VDDA.n832 0.0243392
R7339 VDDA.n964 VDDA.n835 0.0243392
R7340 VDDA.n704 VDDA.n644 0.0243392
R7341 VDDA.n718 VDDA.n647 0.0243392
R7342 VDDA.n734 VDDA.n650 0.0243392
R7343 VDDA.n748 VDDA.n653 0.0243392
R7344 VDDA.n764 VDDA.n656 0.0243392
R7345 VDDA.n778 VDDA.n659 0.0243392
R7346 VDDA.n794 VDDA.n662 0.0243392
R7347 VDDA.n789 VDDA.n662 0.0243392
R7348 VDDA.n775 VDDA.n659 0.0243392
R7349 VDDA.n759 VDDA.n656 0.0243392
R7350 VDDA.n745 VDDA.n653 0.0243392
R7351 VDDA.n729 VDDA.n650 0.0243392
R7352 VDDA.n715 VDDA.n647 0.0243392
R7353 VDDA.n699 VDDA.n644 0.0243392
R7354 VDDA.n842 VDDA.n835 0.0243392
R7355 VDDA.n949 VDDA.n832 0.0243392
R7356 VDDA.n854 VDDA.n829 0.0243392
R7357 VDDA.n925 VDDA.n826 0.0243392
R7358 VDDA.n866 VDDA.n823 0.0243392
R7359 VDDA.n901 VDDA.n820 0.0243392
R7360 VDDA.n878 VDDA.n817 0.0243392
R7361 VDDA.n1133 VDDA.n1132 0.0243392
R7362 VDDA.n1116 VDDA.n1115 0.0243392
R7363 VDDA.n1103 VDDA.n1102 0.0243392
R7364 VDDA.n1086 VDDA.n1085 0.0243392
R7365 VDDA.n1073 VDDA.n1072 0.0243392
R7366 VDDA.n1056 VDDA.n1055 0.0243392
R7367 VDDA.n1043 VDDA.n1042 0.0243392
R7368 VDDA.n615 VDDA.n486 0.0243392
R7369 VDDA.n502 VDDA.n483 0.0243392
R7370 VDDA.n591 VDDA.n480 0.0243392
R7371 VDDA.n514 VDDA.n477 0.0243392
R7372 VDDA.n567 VDDA.n474 0.0243392
R7373 VDDA.n526 VDDA.n471 0.0243392
R7374 VDDA.n543 VDDA.n468 0.0243392
R7375 VDDA.n1190 VDDA.n1183 0.0243392
R7376 VDDA.n1297 VDDA.n1180 0.0243392
R7377 VDDA.n1202 VDDA.n1177 0.0243392
R7378 VDDA.n1273 VDDA.n1174 0.0243392
R7379 VDDA.n1214 VDDA.n1171 0.0243392
R7380 VDDA.n1249 VDDA.n1168 0.0243392
R7381 VDDA.n1226 VDDA.n1165 0.0243392
R7382 VDDA.n2242 VDDA.n1341 0.0243392
R7383 VDDA.n2228 VDDA.n1338 0.0243392
R7384 VDDA.n2212 VDDA.n1335 0.0243392
R7385 VDDA.n2198 VDDA.n1332 0.0243392
R7386 VDDA.n2182 VDDA.n1329 0.0243392
R7387 VDDA.n2168 VDDA.n1326 0.0243392
R7388 VDDA.n2152 VDDA.n1323 0.0243392
R7389 VDDA.n2571 VDDA.n2570 0.0243392
R7390 VDDA.n2554 VDDA.n2553 0.0243392
R7391 VDDA.n2541 VDDA.n2540 0.0243392
R7392 VDDA.n2524 VDDA.n2523 0.0243392
R7393 VDDA.n2511 VDDA.n2510 0.0243392
R7394 VDDA.n2494 VDDA.n2493 0.0243392
R7395 VDDA.n2481 VDDA.n2480 0.0243392
R7396 VDDA.n348 VDDA.n219 0.0243392
R7397 VDDA.n235 VDDA.n216 0.0243392
R7398 VDDA.n324 VDDA.n213 0.0243392
R7399 VDDA.n247 VDDA.n210 0.0243392
R7400 VDDA.n300 VDDA.n207 0.0243392
R7401 VDDA.n259 VDDA.n204 0.0243392
R7402 VDDA.n276 VDDA.n201 0.0243392
R7403 VDDA.n2628 VDDA.n2621 0.0243392
R7404 VDDA.n2735 VDDA.n2618 0.0243392
R7405 VDDA.n2640 VDDA.n2615 0.0243392
R7406 VDDA.n2711 VDDA.n2612 0.0243392
R7407 VDDA.n2652 VDDA.n2609 0.0243392
R7408 VDDA.n2687 VDDA.n2606 0.0243392
R7409 VDDA.n2664 VDDA.n2603 0.0243392
R7410 VDDA.n2919 VDDA.n2918 0.0243392
R7411 VDDA.n2902 VDDA.n2901 0.0243392
R7412 VDDA.n2889 VDDA.n2888 0.0243392
R7413 VDDA.n2872 VDDA.n2871 0.0243392
R7414 VDDA.n2859 VDDA.n2858 0.0243392
R7415 VDDA.n2842 VDDA.n2841 0.0243392
R7416 VDDA.n2829 VDDA.n2828 0.0243392
R7417 VDDA.n170 VDDA.n41 0.0243392
R7418 VDDA.n57 VDDA.n38 0.0243392
R7419 VDDA.n146 VDDA.n35 0.0243392
R7420 VDDA.n69 VDDA.n32 0.0243392
R7421 VDDA.n122 VDDA.n29 0.0243392
R7422 VDDA.n81 VDDA.n26 0.0243392
R7423 VDDA.n98 VDDA.n23 0.0243392
R7424 VDDA.n1565 VDDA.n1431 0.0243392
R7425 VDDA.n1551 VDDA.n1428 0.0243392
R7426 VDDA.n1535 VDDA.n1425 0.0243392
R7427 VDDA.n1521 VDDA.n1422 0.0243392
R7428 VDDA.n1505 VDDA.n1419 0.0243392
R7429 VDDA.n1491 VDDA.n1416 0.0243392
R7430 VDDA.n1475 VDDA.n1413 0.0243392
R7431 VDDA.n2137 VDDA.n1933 0.0217373
R7432 VDDA.n2087 VDDA.n1935 0.0217373
R7433 VDDA.n2010 VDDA.n1937 0.0217373
R7434 VDDA.n1944 VDDA.n1939 0.0217373
R7435 VDDA.n1948 VDDA.n1947 0.0217373
R7436 VDDA.n2014 VDDA.n2013 0.0217373
R7437 VDDA.n2091 VDDA.n2090 0.0217373
R7438 VDDA.n2141 VDDA.n2140 0.0217373
R7439 VDDA.n1946 VDDA.n1939 0.0217373
R7440 VDDA.n1949 VDDA.n1948 0.0217373
R7441 VDDA.n2012 VDDA.n1937 0.0217373
R7442 VDDA.n2015 VDDA.n2014 0.0217373
R7443 VDDA.n2089 VDDA.n1935 0.0217373
R7444 VDDA.n2092 VDDA.n2091 0.0217373
R7445 VDDA.n2139 VDDA.n1933 0.0217373
R7446 VDDA.n2142 VDDA.n2141 0.0217373
R7447 VDDA.n2943 VDDA.n2942 0.0217373
R7448 VDDA.n2940 VDDA.n185 0.0217373
R7449 VDDA.n2934 VDDA.n187 0.0217373
R7450 VDDA.n2937 VDDA.n188 0.0217373
R7451 VDDA.n2763 VDDA.n190 0.0217373
R7452 VDDA.n2766 VDDA.n191 0.0217373
R7453 VDDA.n2595 VDDA.n2594 0.0217373
R7454 VDDA.n2591 VDDA.n362 0.0217373
R7455 VDDA.n2586 VDDA.n364 0.0217373
R7456 VDDA.n2589 VDDA.n365 0.0217373
R7457 VDDA.n2262 VDDA.n457 0.0217373
R7458 VDDA.n2265 VDDA.n458 0.0217373
R7459 VDDA.n426 VDDA.n414 0.0217373
R7460 VDDA.n437 VDDA.n431 0.0217373
R7461 VDDA.n387 VDDA.n370 0.0217373
R7462 VDDA.n387 VDDA.n369 0.0217373
R7463 VDDA.n2398 VDDA.n2397 0.0217373
R7464 VDDA.n2395 VDDA.n406 0.0217373
R7465 VDDA.n429 VDDA.n408 0.0217373
R7466 VDDA.n413 VDDA.n411 0.0217373
R7467 VDDA.n431 VDDA.n409 0.0217373
R7468 VDDA.n430 VDDA.n429 0.0217373
R7469 VDDA.n414 VDDA.n412 0.0217373
R7470 VDDA.n2345 VDDA.n449 0.0217373
R7471 VDDA.n2397 VDDA.n389 0.0217373
R7472 VDDA.n406 VDDA.n389 0.0217373
R7473 VDDA.n2289 VDDA.n451 0.0217373
R7474 VDDA.n2340 VDDA.n450 0.0217373
R7475 VDDA.n2334 VDDA.n2307 0.0217373
R7476 VDDA.n2324 VDDA.n2310 0.0217373
R7477 VDDA.n2290 VDDA.n449 0.0217373
R7478 VDDA.n2340 VDDA.n2339 0.0217373
R7479 VDDA.n2336 VDDA.n2308 0.0217373
R7480 VDDA.n2335 VDDA.n2334 0.0217373
R7481 VDDA.n2325 VDDA.n2311 0.0217373
R7482 VDDA.n1157 VDDA.n1156 0.0217373
R7483 VDDA.n1153 VDDA.n629 0.0217373
R7484 VDDA.n1148 VDDA.n631 0.0217373
R7485 VDDA.n1151 VDDA.n632 0.0217373
R7486 VDDA.n977 VDDA.n634 0.0217373
R7487 VDDA.n980 VDDA.n635 0.0217373
R7488 VDDA.n805 VDDA.n636 0.0217373
R7489 VDDA.n2400 VDDA.n368 0.0217373
R7490 VDDA.n637 VDDA.n634 0.0217373
R7491 VDDA.n637 VDDA.n635 0.0217373
R7492 VDDA.n982 VDDA.n631 0.0217373
R7493 VDDA.n982 VDDA.n632 0.0217373
R7494 VDDA.n1156 VDDA.n1155 0.0217373
R7495 VDDA.n1155 VDDA.n629 0.0217373
R7496 VDDA.n2286 VDDA.n2284 0.0217373
R7497 VDDA.n2284 VDDA.n451 0.0217373
R7498 VDDA.n2402 VDDA.n370 0.0217373
R7499 VDDA.n2399 VDDA.n369 0.0217373
R7500 VDDA.n2401 VDDA.n2400 0.0217373
R7501 VDDA.n460 VDDA.n457 0.0217373
R7502 VDDA.n460 VDDA.n458 0.0217373
R7503 VDDA.n2420 VDDA.n364 0.0217373
R7504 VDDA.n2420 VDDA.n365 0.0217373
R7505 VDDA.n2594 VDDA.n2593 0.0217373
R7506 VDDA.n2593 VDDA.n362 0.0217373
R7507 VDDA.n193 VDDA.n190 0.0217373
R7508 VDDA.n193 VDDA.n191 0.0217373
R7509 VDDA.n2768 VDDA.n187 0.0217373
R7510 VDDA.n2768 VDDA.n188 0.0217373
R7511 VDDA.n2942 VDDA.n183 0.0217373
R7512 VDDA.n185 VDDA.n183 0.0217373
R7513 VDDA.n807 VDDA.n806 0.0217373
R7514 VDDA.n805 VDDA.n804 0.0217373
R7515 VDDA.n2139 VDDA.n1934 0.0217373
R7516 VDDA.n2089 VDDA.n1936 0.0217373
R7517 VDDA.n2012 VDDA.n1938 0.0217373
R7518 VDDA.n1946 VDDA.n1940 0.0217373
R7519 VDDA.n1947 VDDA.n1945 0.0217373
R7520 VDDA.n2013 VDDA.n2011 0.0217373
R7521 VDDA.n2090 VDDA.n2088 0.0217373
R7522 VDDA.n2140 VDDA.n2138 0.0217373
R7523 VDDA.n2011 VDDA.n1950 0.0217373
R7524 VDDA.n2088 VDDA.n2016 0.0217373
R7525 VDDA.n2138 VDDA.n2093 0.0217373
R7526 VDDA.n2311 VDDA.n2309 0.0217373
R7527 VDDA.n2308 VDDA.n2306 0.0217373
R7528 VDDA.n412 VDDA.n410 0.0217373
R7529 VDDA.n409 VDDA.n407 0.0217373
R7530 VDDA.n438 VDDA.n408 0.0217373
R7531 VDDA.n427 VDDA.n411 0.0217373
R7532 VDDA.n439 VDDA.n438 0.0217373
R7533 VDDA.n428 VDDA.n427 0.0217373
R7534 VDDA.n2342 VDDA.n2290 0.0217373
R7535 VDDA.n2394 VDDA.n388 0.0217373
R7536 VDDA.n390 VDDA.n388 0.0217373
R7537 VDDA.n2344 VDDA.n450 0.0217373
R7538 VDDA.n2337 VDDA.n2307 0.0217373
R7539 VDDA.n2326 VDDA.n2310 0.0217373
R7540 VDDA.n2344 VDDA.n2343 0.0217373
R7541 VDDA.n2342 VDDA.n2341 0.0217373
R7542 VDDA.n2338 VDDA.n2337 0.0217373
R7543 VDDA.n2333 VDDA.n2306 0.0217373
R7544 VDDA.n2327 VDDA.n2326 0.0217373
R7545 VDDA.n2323 VDDA.n2309 0.0217373
R7546 VDDA.n804 VDDA.n803 0.0217373
R7547 VDDA.n979 VDDA.n978 0.0217373
R7548 VDDA.n1150 VDDA.n1149 0.0217373
R7549 VDDA.n1154 VDDA.n627 0.0217373
R7550 VDDA.n2264 VDDA.n2263 0.0217373
R7551 VDDA.n2288 VDDA.n2287 0.0217373
R7552 VDDA.n2588 VDDA.n2587 0.0217373
R7553 VDDA.n2592 VDDA.n360 0.0217373
R7554 VDDA.n2765 VDDA.n2764 0.0217373
R7555 VDDA.n2936 VDDA.n2935 0.0217373
R7556 VDDA.n2939 VDDA.n182 0.0217373
R7557 VDDA.n978 VDDA.n633 0.0217373
R7558 VDDA.n1149 VDDA.n630 0.0217373
R7559 VDDA.n628 VDDA.n627 0.0217373
R7560 VDDA.n2287 VDDA.n2285 0.0217373
R7561 VDDA.n2263 VDDA.n456 0.0217373
R7562 VDDA.n2587 VDDA.n363 0.0217373
R7563 VDDA.n361 VDDA.n360 0.0217373
R7564 VDDA.n2764 VDDA.n189 0.0217373
R7565 VDDA.n2935 VDDA.n186 0.0217373
R7566 VDDA.n184 VDDA.n182 0.0217373
R7567 VDDA.n808 VDDA.n807 0.0217373
R7568 VDDA.n809 VDDA.n808 0.0217373
R7569 VDDA VDDA.n3134 0.0164359
R7570 VDDA.n1761 VDDA.n1760 0.0152446
R7571 VDDA.n1759 VDDA.n1758 0.0152446
R7572 VDDA.n1757 VDDA.n1756 0.0152446
R7573 VDDA.n1747 VDDA.n1746 0.0152446
R7574 VDDA.n1594 VDDA.n1590 0.0152446
R7575 VDDA.n1740 VDDA.n1595 0.0152446
R7576 VDDA.n1730 VDDA.n1601 0.0152446
R7577 VDDA.n1729 VDDA.n1728 0.0152446
R7578 VDDA.n1727 VDDA.n1726 0.0152446
R7579 VDDA.n1717 VDDA.n1716 0.0152446
R7580 VDDA.n1612 VDDA.n1608 0.0152446
R7581 VDDA.n1710 VDDA.n1613 0.0152446
R7582 VDDA.n1700 VDDA.n1619 0.0152446
R7583 VDDA.n1699 VDDA.n1698 0.0152446
R7584 VDDA.n1697 VDDA.n1696 0.0152446
R7585 VDDA.n1687 VDDA.n1686 0.0152446
R7586 VDDA.n1630 VDDA.n1626 0.0152446
R7587 VDDA.n1680 VDDA.n1631 0.0152446
R7588 VDDA.n1670 VDDA.n1637 0.0152446
R7589 VDDA.n1669 VDDA.n1668 0.0152446
R7590 VDDA.n1667 VDDA.n1666 0.0152446
R7591 VDDA.n1657 VDDA.n1656 0.0152446
R7592 VDDA.n1647 VDDA.n1644 0.0152446
R7593 VDDA.n1650 VDDA.n1648 0.0152446
R7594 VDDA.n1648 VDDA.n1647 0.0152446
R7595 VDDA.n1656 VDDA.n1644 0.0152446
R7596 VDDA.n1658 VDDA.n1657 0.0152446
R7597 VDDA.n1668 VDDA.n1667 0.0152446
R7598 VDDA.n1670 VDDA.n1669 0.0152446
R7599 VDDA.n1637 VDDA.n1636 0.0152446
R7600 VDDA.n1631 VDDA.n1630 0.0152446
R7601 VDDA.n1686 VDDA.n1626 0.0152446
R7602 VDDA.n1688 VDDA.n1687 0.0152446
R7603 VDDA.n1698 VDDA.n1697 0.0152446
R7604 VDDA.n1700 VDDA.n1699 0.0152446
R7605 VDDA.n1619 VDDA.n1618 0.0152446
R7606 VDDA.n1613 VDDA.n1612 0.0152446
R7607 VDDA.n1716 VDDA.n1608 0.0152446
R7608 VDDA.n1718 VDDA.n1717 0.0152446
R7609 VDDA.n1728 VDDA.n1727 0.0152446
R7610 VDDA.n1730 VDDA.n1729 0.0152446
R7611 VDDA.n1601 VDDA.n1600 0.0152446
R7612 VDDA.n1595 VDDA.n1594 0.0152446
R7613 VDDA.n1746 VDDA.n1590 0.0152446
R7614 VDDA.n1748 VDDA.n1747 0.0152446
R7615 VDDA.n1758 VDDA.n1757 0.0152446
R7616 VDDA.n1760 VDDA.n1759 0.0152446
R7617 VDDA.n1762 VDDA.n1761 0.0152446
R7618 VDDA.n1762 VDDA.n1408 0.0142311
R7619 VDDA.n1588 VDDA.n1583 0.0142311
R7620 VDDA.n1749 VDDA.n1748 0.0142311
R7621 VDDA.n1739 VDDA.n1738 0.0142311
R7622 VDDA.n1600 VDDA.n1596 0.0142311
R7623 VDDA.n1606 VDDA.n1602 0.0142311
R7624 VDDA.n1719 VDDA.n1718 0.0142311
R7625 VDDA.n1709 VDDA.n1708 0.0142311
R7626 VDDA.n1618 VDDA.n1614 0.0142311
R7627 VDDA.n1624 VDDA.n1620 0.0142311
R7628 VDDA.n1689 VDDA.n1688 0.0142311
R7629 VDDA.n1679 VDDA.n1678 0.0142311
R7630 VDDA.n1636 VDDA.n1632 0.0142311
R7631 VDDA.n1642 VDDA.n1638 0.0142311
R7632 VDDA.n1659 VDDA.n1658 0.0142311
R7633 VDDA.n1649 VDDA.n1646 0.0142311
R7634 VDDA.n1650 VDDA.n1649 0.0142311
R7635 VDDA.n1660 VDDA.n1659 0.0142311
R7636 VDDA.n1666 VDDA.n1638 0.0142311
R7637 VDDA.n1676 VDDA.n1632 0.0142311
R7638 VDDA.n1680 VDDA.n1679 0.0142311
R7639 VDDA.n1690 VDDA.n1689 0.0142311
R7640 VDDA.n1696 VDDA.n1620 0.0142311
R7641 VDDA.n1706 VDDA.n1614 0.0142311
R7642 VDDA.n1710 VDDA.n1709 0.0142311
R7643 VDDA.n1720 VDDA.n1719 0.0142311
R7644 VDDA.n1726 VDDA.n1602 0.0142311
R7645 VDDA.n1736 VDDA.n1596 0.0142311
R7646 VDDA.n1740 VDDA.n1739 0.0142311
R7647 VDDA.n1750 VDDA.n1749 0.0142311
R7648 VDDA.n1756 VDDA.n1583 0.0142311
R7649 VDDA.n1409 VDDA.n1408 0.0142311
R7650 VDDA.n1581 VDDA.n1580 0.0141594
R7651 VDDA.n1750 VDDA.n1589 0.0132169
R7652 VDDA.n1737 VDDA.n1736 0.0132169
R7653 VDDA.n1720 VDDA.n1607 0.0132169
R7654 VDDA.n1707 VDDA.n1706 0.0132169
R7655 VDDA.n1690 VDDA.n1625 0.0132169
R7656 VDDA.n1677 VDDA.n1676 0.0132169
R7657 VDDA.n1660 VDDA.n1643 0.0132169
R7658 VDDA.n1643 VDDA.n1642 0.0132169
R7659 VDDA.n1678 VDDA.n1677 0.0132169
R7660 VDDA.n1625 VDDA.n1624 0.0132169
R7661 VDDA.n1708 VDDA.n1707 0.0132169
R7662 VDDA.n1607 VDDA.n1606 0.0132169
R7663 VDDA.n1738 VDDA.n1737 0.0132169
R7664 VDDA.n1589 VDDA.n1588 0.0132169
R7665 VDDA.n2258 VDDA.n1161 0.0107812
R7666 VDDA.n2599 VDDA.n197 0.0107812
R7667 VDDA.n1580 VDDA.n197 0.00894531
R7668 VDDA.n2258 VDDA.n2257 0.00887187
R7669 VDDA.n973 VDDA.n813 0.00564062
R7670 VDDA.n973 VDDA.n464 0.00564062
R7671 VDDA.n1161 VDDA.n464 0.00564062
R7672 VDDA.n2759 VDDA.n2599 0.00564062
R7673 VDDA.n2759 VDDA.n19 0.00564062
R7674 VDDA.n2947 VDDA.n19 0.00564062
R7675 VDDA.n1908 VDDA.n1368 0.00211562
R7676 VDDA.n3035 VDDA.n3033 0.00202782
R7677 VDDA.n3033 VDDA.n2965 0.00202782
R7678 VDDA.n2984 VDDA.n0 0.00166081
R7679 VDDA.n2983 VDDA.n2981 0.00166081
R7680 VDDA.n2987 VDDA.n2985 0.00166081
R7681 VDDA.n2986 VDDA.n2980 0.00166081
R7682 VDDA.n2990 VDDA.n2988 0.00166081
R7683 VDDA.n2989 VDDA.n2979 0.00166081
R7684 VDDA.n2993 VDDA.n2991 0.00166081
R7685 VDDA.n2992 VDDA.n2978 0.00166081
R7686 VDDA.n2996 VDDA.n2994 0.00166081
R7687 VDDA.n2995 VDDA.n2977 0.00166081
R7688 VDDA.n2999 VDDA.n2997 0.00166081
R7689 VDDA.n2998 VDDA.n2976 0.00166081
R7690 VDDA.n3002 VDDA.n3000 0.00166081
R7691 VDDA.n3001 VDDA.n2975 0.00166081
R7692 VDDA.n3005 VDDA.n3003 0.00166081
R7693 VDDA.n3004 VDDA.n2974 0.00166081
R7694 VDDA.n3008 VDDA.n3006 0.00166081
R7695 VDDA.n3007 VDDA.n2973 0.00166081
R7696 VDDA.n3011 VDDA.n3009 0.00166081
R7697 VDDA.n3010 VDDA.n2972 0.00166081
R7698 VDDA.n3014 VDDA.n3012 0.00166081
R7699 VDDA.n3013 VDDA.n2971 0.00166081
R7700 VDDA.n3017 VDDA.n3015 0.00166081
R7701 VDDA.n3016 VDDA.n2970 0.00166081
R7702 VDDA.n3020 VDDA.n3018 0.00166081
R7703 VDDA.n3019 VDDA.n2969 0.00166081
R7704 VDDA.n3023 VDDA.n3021 0.00166081
R7705 VDDA.n3022 VDDA.n2968 0.00166081
R7706 VDDA.n3026 VDDA.n3024 0.00166081
R7707 VDDA.n3025 VDDA.n2967 0.00166081
R7708 VDDA.n3029 VDDA.n3027 0.00166081
R7709 VDDA.n3028 VDDA.n2966 0.00166081
R7710 VDDA.n3032 VDDA.n3030 0.00166081
R7711 VDDA.n3031 VDDA.n2965 0.00166081
R7712 VDDA.n3034 VDDA.n2964 0.00166081
R7713 VDDA.n3038 VDDA.n3036 0.00166081
R7714 VDDA.n3037 VDDA.n2963 0.00166081
R7715 VDDA.n3041 VDDA.n3039 0.00166081
R7716 VDDA.n3040 VDDA.n2962 0.00166081
R7717 VDDA.n3044 VDDA.n3042 0.00166081
R7718 VDDA.n3043 VDDA.n2961 0.00166081
R7719 VDDA.n3047 VDDA.n3045 0.00166081
R7720 VDDA.n3046 VDDA.n2960 0.00166081
R7721 VDDA.n3050 VDDA.n3048 0.00166081
R7722 VDDA.n3049 VDDA.n2959 0.00166081
R7723 VDDA.n3053 VDDA.n3051 0.00166081
R7724 VDDA.n3052 VDDA.n2958 0.00166081
R7725 VDDA.n3056 VDDA.n3054 0.00166081
R7726 VDDA.n3055 VDDA.n2957 0.00166081
R7727 VDDA.n3059 VDDA.n3057 0.00166081
R7728 VDDA.n3058 VDDA.n2956 0.00166081
R7729 VDDA.n3062 VDDA.n3060 0.00166081
R7730 VDDA.n3061 VDDA.n2955 0.00166081
R7731 VDDA.n3065 VDDA.n3063 0.00166081
R7732 VDDA.n3064 VDDA.n2954 0.00166081
R7733 VDDA.n3068 VDDA.n3066 0.00166081
R7734 VDDA.n3067 VDDA.n2953 0.00166081
R7735 VDDA.n3071 VDDA.n3069 0.00166081
R7736 VDDA.n3070 VDDA.n2952 0.00166081
R7737 VDDA.n3074 VDDA.n3072 0.00166081
R7738 VDDA.n3073 VDDA.n2951 0.00166081
R7739 VDDA.n3077 VDDA.n3075 0.00166081
R7740 VDDA.n3076 VDDA.n2950 0.00166081
R7741 VDDA.n3080 VDDA.n3078 0.00166081
R7742 VDDA.n3079 VDDA.n2949 0.00166081
R7743 VDDA.n3083 VDDA.n3081 0.00166081
R7744 VDDA.n3082 VDDA.n2948 0.00166081
R7745 VDDA.n3132 VDDA.n3084 0.00166081
R7746 VDDA.n3134 VDDA.n0 0.00166081
R7747 VDDA.n2984 VDDA.n2983 0.00166081
R7748 VDDA.n2985 VDDA.n2981 0.00166081
R7749 VDDA.n2987 VDDA.n2986 0.00166081
R7750 VDDA.n2988 VDDA.n2980 0.00166081
R7751 VDDA.n2990 VDDA.n2989 0.00166081
R7752 VDDA.n2991 VDDA.n2979 0.00166081
R7753 VDDA.n2993 VDDA.n2992 0.00166081
R7754 VDDA.n2994 VDDA.n2978 0.00166081
R7755 VDDA.n2996 VDDA.n2995 0.00166081
R7756 VDDA.n2997 VDDA.n2977 0.00166081
R7757 VDDA.n2999 VDDA.n2998 0.00166081
R7758 VDDA.n3000 VDDA.n2976 0.00166081
R7759 VDDA.n3002 VDDA.n3001 0.00166081
R7760 VDDA.n3003 VDDA.n2975 0.00166081
R7761 VDDA.n3005 VDDA.n3004 0.00166081
R7762 VDDA.n3006 VDDA.n2974 0.00166081
R7763 VDDA.n3008 VDDA.n3007 0.00166081
R7764 VDDA.n3009 VDDA.n2973 0.00166081
R7765 VDDA.n3011 VDDA.n3010 0.00166081
R7766 VDDA.n3012 VDDA.n2972 0.00166081
R7767 VDDA.n3014 VDDA.n3013 0.00166081
R7768 VDDA.n3015 VDDA.n2971 0.00166081
R7769 VDDA.n3017 VDDA.n3016 0.00166081
R7770 VDDA.n3018 VDDA.n2970 0.00166081
R7771 VDDA.n3020 VDDA.n3019 0.00166081
R7772 VDDA.n3021 VDDA.n2969 0.00166081
R7773 VDDA.n3023 VDDA.n3022 0.00166081
R7774 VDDA.n3024 VDDA.n2968 0.00166081
R7775 VDDA.n3026 VDDA.n3025 0.00166081
R7776 VDDA.n3027 VDDA.n2967 0.00166081
R7777 VDDA.n3029 VDDA.n3028 0.00166081
R7778 VDDA.n3030 VDDA.n2966 0.00166081
R7779 VDDA.n3032 VDDA.n3031 0.00166081
R7780 VDDA.n3035 VDDA.n3034 0.00166081
R7781 VDDA.n3036 VDDA.n2964 0.00166081
R7782 VDDA.n3038 VDDA.n3037 0.00166081
R7783 VDDA.n3039 VDDA.n2963 0.00166081
R7784 VDDA.n3041 VDDA.n3040 0.00166081
R7785 VDDA.n3042 VDDA.n2962 0.00166081
R7786 VDDA.n3044 VDDA.n3043 0.00166081
R7787 VDDA.n3045 VDDA.n2961 0.00166081
R7788 VDDA.n3047 VDDA.n3046 0.00166081
R7789 VDDA.n3048 VDDA.n2960 0.00166081
R7790 VDDA.n3050 VDDA.n3049 0.00166081
R7791 VDDA.n3051 VDDA.n2959 0.00166081
R7792 VDDA.n3053 VDDA.n3052 0.00166081
R7793 VDDA.n3054 VDDA.n2958 0.00166081
R7794 VDDA.n3056 VDDA.n3055 0.00166081
R7795 VDDA.n3057 VDDA.n2957 0.00166081
R7796 VDDA.n3059 VDDA.n3058 0.00166081
R7797 VDDA.n3060 VDDA.n2956 0.00166081
R7798 VDDA.n3062 VDDA.n3061 0.00166081
R7799 VDDA.n3063 VDDA.n2955 0.00166081
R7800 VDDA.n3065 VDDA.n3064 0.00166081
R7801 VDDA.n3066 VDDA.n2954 0.00166081
R7802 VDDA.n3068 VDDA.n3067 0.00166081
R7803 VDDA.n3069 VDDA.n2953 0.00166081
R7804 VDDA.n3071 VDDA.n3070 0.00166081
R7805 VDDA.n3072 VDDA.n2952 0.00166081
R7806 VDDA.n3074 VDDA.n3073 0.00166081
R7807 VDDA.n3075 VDDA.n2951 0.00166081
R7808 VDDA.n3077 VDDA.n3076 0.00166081
R7809 VDDA.n3078 VDDA.n2950 0.00166081
R7810 VDDA.n3080 VDDA.n3079 0.00166081
R7811 VDDA.n3081 VDDA.n2949 0.00166081
R7812 VDDA.n3083 VDDA.n3082 0.00166081
R7813 VDDA.n3084 VDDA.n2948 0.00166081
R7814 VDDA.t59 VDDA.n1458 0.00152174
R7815 VDDA.t138 VDDA.n1459 0.00152174
R7816 VDDA.t393 VDDA.n1460 0.00152174
R7817 VDDA.t163 VDDA.n1461 0.00152174
R7818 VDDA.t386 VDDA.n1462 0.00152174
R7819 VDDA.n1581 VDDA.n1368 0.00138125
R7820 VDDA.n3086 VDDA.n3085 0.00133044
R7821 VDDA.n3086 VDDA.n1 0.00133044
R7822 VDDA.n3130 VDDA.n3087 0.00133044
R7823 VDDA.n3087 VDDA.n2 0.00133044
R7824 VDDA.n3128 VDDA.n3088 0.00133044
R7825 VDDA.n3088 VDDA.n3 0.00133044
R7826 VDDA.n3126 VDDA.n3089 0.00133044
R7827 VDDA.n3089 VDDA.n4 0.00133044
R7828 VDDA.n3124 VDDA.n3090 0.00133044
R7829 VDDA.n3090 VDDA.n5 0.00133044
R7830 VDDA.n3122 VDDA.n3091 0.00133044
R7831 VDDA.n3091 VDDA.n6 0.00133044
R7832 VDDA.n3120 VDDA.n3092 0.00133044
R7833 VDDA.n3092 VDDA.n7 0.00133044
R7834 VDDA.n3118 VDDA.n3093 0.00133044
R7835 VDDA.n3093 VDDA.n8 0.00133044
R7836 VDDA.n3116 VDDA.n3094 0.00133044
R7837 VDDA.n3094 VDDA.n9 0.00133044
R7838 VDDA.n3114 VDDA.n3095 0.00133044
R7839 VDDA.n3095 VDDA.n10 0.00133044
R7840 VDDA.n3112 VDDA.n3096 0.00133044
R7841 VDDA.n3096 VDDA.n11 0.00133044
R7842 VDDA.n3110 VDDA.n3097 0.00133044
R7843 VDDA.n3097 VDDA.n12 0.00133044
R7844 VDDA.n3108 VDDA.n3098 0.00133044
R7845 VDDA.n3098 VDDA.n13 0.00133044
R7846 VDDA.n3106 VDDA.n3099 0.00133044
R7847 VDDA.n3099 VDDA.n14 0.00133044
R7848 VDDA.n3104 VDDA.n3100 0.00133044
R7849 VDDA.n3100 VDDA.n15 0.00133044
R7850 VDDA.n3102 VDDA.n16 0.00133044
R7851 VDDA.n3101 VDDA.n17 0.00133044
R7852 VDDA.n3103 VDDA.n15 0.00133044
R7853 VDDA.n3105 VDDA.n14 0.00133044
R7854 VDDA.n3107 VDDA.n13 0.00133044
R7855 VDDA.n3109 VDDA.n12 0.00133044
R7856 VDDA.n3111 VDDA.n11 0.00133044
R7857 VDDA.n3113 VDDA.n10 0.00133044
R7858 VDDA.n3115 VDDA.n9 0.00133044
R7859 VDDA.n3117 VDDA.n8 0.00133044
R7860 VDDA.n3119 VDDA.n7 0.00133044
R7861 VDDA.n3121 VDDA.n6 0.00133044
R7862 VDDA.n3123 VDDA.n5 0.00133044
R7863 VDDA.n3125 VDDA.n4 0.00133044
R7864 VDDA.n3127 VDDA.n3 0.00133044
R7865 VDDA.n3129 VDDA.n2 0.00133044
R7866 VDDA.n3131 VDDA.n1 0.00133044
R7867 VDDA.n3103 VDDA.n3102 0.00133044
R7868 VDDA.n3105 VDDA.n3104 0.00133044
R7869 VDDA.n3107 VDDA.n3106 0.00133044
R7870 VDDA.n3109 VDDA.n3108 0.00133044
R7871 VDDA.n3111 VDDA.n3110 0.00133044
R7872 VDDA.n3113 VDDA.n3112 0.00133044
R7873 VDDA.n3115 VDDA.n3114 0.00133044
R7874 VDDA.n3117 VDDA.n3116 0.00133044
R7875 VDDA.n3119 VDDA.n3118 0.00133044
R7876 VDDA.n3121 VDDA.n3120 0.00133044
R7877 VDDA.n3123 VDDA.n3122 0.00133044
R7878 VDDA.n3125 VDDA.n3124 0.00133044
R7879 VDDA.n3127 VDDA.n3126 0.00133044
R7880 VDDA.n3129 VDDA.n3128 0.00133044
R7881 VDDA.n3131 VDDA.n3130 0.00133044
R7882 VDDA.n3085 VDDA.n18 0.00133044
R7883 VDDA.n3101 VDDA.n16 0.00133044
R7884 VDDA.n3133 VDDA.n2982 0.00116094
R7885 VDDA.n2982 VDDA.n18 0.00116094
R7886 VOUT-.n178 VOUT-.t7 110.386
R7887 VOUT-.n39 VOUT-.n38 34.9935
R7888 VOUT-.n28 VOUT-.n27 34.9935
R7889 VOUT-.n30 VOUT-.n29 34.9935
R7890 VOUT-.n33 VOUT-.n32 34.9935
R7891 VOUT-.n36 VOUT-.n35 34.9935
R7892 VOUT-.n42 VOUT-.n41 34.9935
R7893 VOUT-.n185 VOUT-.n184 9.73997
R7894 VOUT-.n181 VOUT-.n180 9.73997
R7895 VOUT-.n188 VOUT-.n187 9.73997
R7896 VOUT-.n186 VOUT-.n181 6.64633
R7897 VOUT-.n186 VOUT-.n185 6.64633
R7898 VOUT-.n38 VOUT-.t18 6.56717
R7899 VOUT-.n38 VOUT-.t11 6.56717
R7900 VOUT-.n27 VOUT-.t10 6.56717
R7901 VOUT-.n27 VOUT-.t1 6.56717
R7902 VOUT-.n29 VOUT-.t0 6.56717
R7903 VOUT-.n29 VOUT-.t14 6.56717
R7904 VOUT-.n32 VOUT-.t13 6.56717
R7905 VOUT-.n32 VOUT-.t2 6.56717
R7906 VOUT-.n35 VOUT-.t16 6.56717
R7907 VOUT-.n35 VOUT-.t3 6.56717
R7908 VOUT-.n41 VOUT-.t4 6.56717
R7909 VOUT-.n41 VOUT-.t8 6.56717
R7910 VOUT-.n31 VOUT-.n28 6.3755
R7911 VOUT-.n40 VOUT-.n39 6.3755
R7912 VOUT-.n188 VOUT-.n186 6.02133
R7913 VOUT-.n31 VOUT-.n30 5.813
R7914 VOUT-.n34 VOUT-.n33 5.813
R7915 VOUT-.n37 VOUT-.n36 5.813
R7916 VOUT-.n42 VOUT-.n40 5.813
R7917 VOUT-.n46 VOUT-.n26 5.063
R7918 VOUT-.n43 VOUT-.n19 5.063
R7919 VOUT-.n109 VOUT-.t35 4.8295
R7920 VOUT-.n108 VOUT-.t71 4.8295
R7921 VOUT-.n107 VOUT-.t106 4.8295
R7922 VOUT-.n106 VOUT-.t141 4.8295
R7923 VOUT-.n105 VOUT-.t54 4.8295
R7924 VOUT-.n104 VOUT-.t100 4.8295
R7925 VOUT-.n110 VOUT-.t147 4.8295
R7926 VOUT-.n121 VOUT-.t132 4.8295
R7927 VOUT-.n122 VOUT-.t42 4.8295
R7928 VOUT-.n124 VOUT-.t103 4.8295
R7929 VOUT-.n125 VOUT-.t86 4.8295
R7930 VOUT-.n127 VOUT-.t67 4.8295
R7931 VOUT-.n128 VOUT-.t48 4.8295
R7932 VOUT-.n130 VOUT-.t98 4.8295
R7933 VOUT-.n131 VOUT-.t80 4.8295
R7934 VOUT-.n133 VOUT-.t61 4.8295
R7935 VOUT-.n134 VOUT-.t43 4.8295
R7936 VOUT-.n136 VOUT-.t19 4.8295
R7937 VOUT-.n137 VOUT-.t142 4.8295
R7938 VOUT-.n139 VOUT-.t55 4.8295
R7939 VOUT-.n140 VOUT-.t36 4.8295
R7940 VOUT-.n142 VOUT-.t151 4.8295
R7941 VOUT-.n143 VOUT-.t134 4.8295
R7942 VOUT-.n145 VOUT-.t111 4.8295
R7943 VOUT-.n146 VOUT-.t97 4.8295
R7944 VOUT-.n148 VOUT-.t74 4.8295
R7945 VOUT-.n149 VOUT-.t59 4.8295
R7946 VOUT-.n71 VOUT-.t96 4.8295
R7947 VOUT-.n73 VOUT-.t58 4.8295
R7948 VOUT-.n86 VOUT-.t117 4.8295
R7949 VOUT-.n87 VOUT-.t102 4.8295
R7950 VOUT-.n89 VOUT-.t153 4.8295
R7951 VOUT-.n90 VOUT-.t136 4.8295
R7952 VOUT-.n92 VOUT-.t62 4.8295
R7953 VOUT-.n93 VOUT-.t30 4.8295
R7954 VOUT-.n95 VOUT-.t66 4.8295
R7955 VOUT-.n96 VOUT-.t47 4.8295
R7956 VOUT-.n98 VOUT-.t29 4.8295
R7957 VOUT-.n99 VOUT-.t150 4.8295
R7958 VOUT-.n101 VOUT-.t70 4.8295
R7959 VOUT-.n102 VOUT-.t53 4.8295
R7960 VOUT-.n151 VOUT-.t108 4.8295
R7961 VOUT-.n112 VOUT-.t75 4.8154
R7962 VOUT-.n74 VOUT-.t146 4.806
R7963 VOUT-.n75 VOUT-.t119 4.806
R7964 VOUT-.n76 VOUT-.t139 4.806
R7965 VOUT-.n77 VOUT-.t38 4.806
R7966 VOUT-.n78 VOUT-.t154 4.806
R7967 VOUT-.n79 VOUT-.t56 4.806
R7968 VOUT-.n80 VOUT-.t91 4.806
R7969 VOUT-.n81 VOUT-.t127 4.806
R7970 VOUT-.n82 VOUT-.t107 4.806
R7971 VOUT-.n83 VOUT-.t148 4.806
R7972 VOUT-.n84 VOUT-.t45 4.806
R7973 VOUT-.n109 VOUT-.t52 4.5005
R7974 VOUT-.n108 VOUT-.t90 4.5005
R7975 VOUT-.n107 VOUT-.t125 4.5005
R7976 VOUT-.n106 VOUT-.t25 4.5005
R7977 VOUT-.n105 VOUT-.t145 4.5005
R7978 VOUT-.n104 VOUT-.t64 4.5005
R7979 VOUT-.n120 VOUT-.t23 4.5005
R7980 VOUT-.n119 VOUT-.t46 4.5005
R7981 VOUT-.n118 VOUT-.t149 4.5005
R7982 VOUT-.n117 VOUT-.t109 4.5005
R7983 VOUT-.n116 VOUT-.t128 4.5005
R7984 VOUT-.n115 VOUT-.t94 4.5005
R7985 VOUT-.n114 VOUT-.t57 4.5005
R7986 VOUT-.n113 VOUT-.t155 4.5005
R7987 VOUT-.n112 VOUT-.t41 4.5005
R7988 VOUT-.n111 VOUT-.t140 4.5005
R7989 VOUT-.n110 VOUT-.t122 4.5005
R7990 VOUT-.n121 VOUT-.t95 4.5005
R7991 VOUT-.n123 VOUT-.t60 4.5005
R7992 VOUT-.n122 VOUT-.t78 4.5005
R7993 VOUT-.n124 VOUT-.t69 4.5005
R7994 VOUT-.n126 VOUT-.t32 4.5005
R7995 VOUT-.n125 VOUT-.t120 4.5005
R7996 VOUT-.n127 VOUT-.t27 4.5005
R7997 VOUT-.n129 VOUT-.t131 4.5005
R7998 VOUT-.n128 VOUT-.t82 4.5005
R7999 VOUT-.n130 VOUT-.t65 4.5005
R8000 VOUT-.n132 VOUT-.t26 4.5005
R8001 VOUT-.n131 VOUT-.t113 4.5005
R8002 VOUT-.n133 VOUT-.t24 4.5005
R8003 VOUT-.n135 VOUT-.t126 4.5005
R8004 VOUT-.n134 VOUT-.t76 4.5005
R8005 VOUT-.n136 VOUT-.t123 4.5005
R8006 VOUT-.n138 VOUT-.t88 4.5005
R8007 VOUT-.n137 VOUT-.t37 4.5005
R8008 VOUT-.n139 VOUT-.t156 4.5005
R8009 VOUT-.n141 VOUT-.t121 4.5005
R8010 VOUT-.n140 VOUT-.t72 4.5005
R8011 VOUT-.n142 VOUT-.t115 4.5005
R8012 VOUT-.n144 VOUT-.t83 4.5005
R8013 VOUT-.n143 VOUT-.t31 4.5005
R8014 VOUT-.n145 VOUT-.t77 4.5005
R8015 VOUT-.n147 VOUT-.t44 4.5005
R8016 VOUT-.n146 VOUT-.t129 4.5005
R8017 VOUT-.n148 VOUT-.t40 4.5005
R8018 VOUT-.n150 VOUT-.t143 4.5005
R8019 VOUT-.n149 VOUT-.t93 4.5005
R8020 VOUT-.n71 VOUT-.t63 4.5005
R8021 VOUT-.n72 VOUT-.t22 4.5005
R8022 VOUT-.n73 VOUT-.t20 4.5005
R8023 VOUT-.n85 VOUT-.t118 4.5005
R8024 VOUT-.n84 VOUT-.t144 4.5005
R8025 VOUT-.n83 VOUT-.t105 4.5005
R8026 VOUT-.n82 VOUT-.t68 4.5005
R8027 VOUT-.n81 VOUT-.t89 4.5005
R8028 VOUT-.n80 VOUT-.t51 4.5005
R8029 VOUT-.n79 VOUT-.t152 4.5005
R8030 VOUT-.n78 VOUT-.t112 4.5005
R8031 VOUT-.n77 VOUT-.t135 4.5005
R8032 VOUT-.n76 VOUT-.t101 4.5005
R8033 VOUT-.n75 VOUT-.t79 4.5005
R8034 VOUT-.n74 VOUT-.t104 4.5005
R8035 VOUT-.n86 VOUT-.t85 4.5005
R8036 VOUT-.n88 VOUT-.t50 4.5005
R8037 VOUT-.n87 VOUT-.t137 4.5005
R8038 VOUT-.n89 VOUT-.t116 4.5005
R8039 VOUT-.n91 VOUT-.t84 4.5005
R8040 VOUT-.n90 VOUT-.t33 4.5005
R8041 VOUT-.n92 VOUT-.t110 4.5005
R8042 VOUT-.n94 VOUT-.t21 4.5005
R8043 VOUT-.n93 VOUT-.t114 4.5005
R8044 VOUT-.n95 VOUT-.t28 4.5005
R8045 VOUT-.n97 VOUT-.t130 4.5005
R8046 VOUT-.n96 VOUT-.t81 4.5005
R8047 VOUT-.n98 VOUT-.t133 4.5005
R8048 VOUT-.n100 VOUT-.t99 4.5005
R8049 VOUT-.n99 VOUT-.t49 4.5005
R8050 VOUT-.n101 VOUT-.t34 4.5005
R8051 VOUT-.n103 VOUT-.t138 4.5005
R8052 VOUT-.n102 VOUT-.t87 4.5005
R8053 VOUT-.n151 VOUT-.t73 4.5005
R8054 VOUT-.n152 VOUT-.t39 4.5005
R8055 VOUT-.n153 VOUT-.t124 4.5005
R8056 VOUT-.n154 VOUT-.t92 4.5005
R8057 VOUT-.n47 VOUT-.n46 4.5005
R8058 VOUT-.n45 VOUT-.n24 4.5005
R8059 VOUT-.n44 VOUT-.n23 4.5005
R8060 VOUT-.n43 VOUT-.n20 4.5005
R8061 VOUT-.n65 VOUT-.n64 4.5005
R8062 VOUT-.n16 VOUT-.n13 4.5005
R8063 VOUT-.n65 VOUT-.n13 4.5005
R8064 VOUT-.n66 VOUT-.n9 4.5005
R8065 VOUT-.n66 VOUT-.n11 4.5005
R8066 VOUT-.n66 VOUT-.n65 4.5005
R8067 VOUT-.n163 VOUT-.n69 4.5005
R8068 VOUT-.n164 VOUT-.n163 4.5005
R8069 VOUT-.n164 VOUT-.n5 4.5005
R8070 VOUT-.n165 VOUT-.n4 4.5005
R8071 VOUT-.n165 VOUT-.n164 4.5005
R8072 VOUT-.n177 VOUT-.n176 4.5005
R8073 VOUT-.n177 VOUT-.n1 4.5005
R8074 VOUT-.n173 VOUT-.n1 4.5005
R8075 VOUT-.n170 VOUT-.n1 4.5005
R8076 VOUT-.n171 VOUT-.n1 4.5005
R8077 VOUT-.n173 VOUT-.n172 4.5005
R8078 VOUT-.n172 VOUT-.n170 4.5005
R8079 VOUT-.n172 VOUT-.n171 4.5005
R8080 VOUT-.n184 VOUT-.t5 3.42907
R8081 VOUT-.n184 VOUT-.t15 3.42907
R8082 VOUT-.n180 VOUT-.t17 3.42907
R8083 VOUT-.n180 VOUT-.t9 3.42907
R8084 VOUT-.n187 VOUT-.t6 3.42907
R8085 VOUT-.n187 VOUT-.t12 3.42907
R8086 VOUT-.n63 VOUT-.n62 2.24601
R8087 VOUT-.n14 VOUT-.n8 2.24601
R8088 VOUT-.n175 VOUT-.n174 2.24601
R8089 VOUT-.n169 VOUT-.n168 2.24601
R8090 VOUT-.n162 VOUT-.n161 2.24477
R8091 VOUT-.n7 VOUT-.n2 2.24477
R8092 VOUT-.n66 VOUT-.n10 2.24063
R8093 VOUT-.n165 VOUT-.n3 2.24063
R8094 VOUT-.n172 VOUT-.n0 2.24063
R8095 VOUT-.n13 VOUT-.n12 2.24063
R8096 VOUT-.n163 VOUT-.n67 2.24063
R8097 VOUT-.n68 VOUT-.n5 2.24063
R8098 VOUT-.n176 VOUT-.n167 2.24063
R8099 VOUT-.n176 VOUT-.n166 2.24063
R8100 VOUT-.n64 VOUT-.n17 2.23934
R8101 VOUT-.n64 VOUT-.n15 2.23934
R8102 VOUT-.n185 VOUT-.n183 1.83719
R8103 VOUT-.n196 VOUT-.n181 1.72967
R8104 VOUT-.n189 VOUT-.n188 1.72967
R8105 VOUT-.n50 VOUT-.n25 1.5005
R8106 VOUT-.n52 VOUT-.n51 1.5005
R8107 VOUT-.n53 VOUT-.n22 1.5005
R8108 VOUT-.n55 VOUT-.n54 1.5005
R8109 VOUT-.n56 VOUT-.n21 1.5005
R8110 VOUT-.n58 VOUT-.n57 1.5005
R8111 VOUT-.n59 VOUT-.n18 1.5005
R8112 VOUT-.n61 VOUT-.n60 1.5005
R8113 VOUT-.n191 VOUT-.n190 1.5005
R8114 VOUT-.n192 VOUT-.n182 1.5005
R8115 VOUT-.n194 VOUT-.n193 1.5005
R8116 VOUT-.n195 VOUT-.n179 1.5005
R8117 VOUT-.n197 VOUT-.n196 1.5005
R8118 VOUT-.n30 VOUT-.n20 1.313
R8119 VOUT-.n33 VOUT-.n23 1.313
R8120 VOUT-.n36 VOUT-.n24 1.313
R8121 VOUT-.n47 VOUT-.n42 1.313
R8122 VOUT-.n28 VOUT-.n19 1.313
R8123 VOUT-.n39 VOUT-.n26 1.313
R8124 VOUT-.n161 VOUT-.n160 1.1455
R8125 VOUT-.n155 VOUT-.n6 1.13717
R8126 VOUT-.n157 VOUT-.n156 1.13717
R8127 VOUT-.n159 VOUT-.n158 1.13717
R8128 VOUT-.n164 VOUT-.n6 1.13717
R8129 VOUT-.n157 VOUT-.n7 1.13717
R8130 VOUT-.n158 VOUT-.n4 1.13717
R8131 VOUT-.n70 VOUT-.n69 1.13717
R8132 VOUT-.n49 VOUT-.n26 0.715216
R8133 VOUT-.n58 VOUT-.n20 0.65675
R8134 VOUT-.n54 VOUT-.n23 0.65675
R8135 VOUT-.n52 VOUT-.n24 0.65675
R8136 VOUT-.n48 VOUT-.n47 0.65675
R8137 VOUT-.n60 VOUT-.n19 0.65675
R8138 VOUT-.n160 VOUT-.n159 0.585
R8139 VOUT-.n50 VOUT-.n49 0.564601
R8140 VOUT-.n46 VOUT-.n45 0.563
R8141 VOUT-.n45 VOUT-.n44 0.563
R8142 VOUT-.n44 VOUT-.n43 0.563
R8143 VOUT-.n34 VOUT-.n31 0.563
R8144 VOUT-.n37 VOUT-.n34 0.563
R8145 VOUT-.n40 VOUT-.n37 0.563
R8146 VOUT-.n176 VOUT-.n165 0.5455
R8147 VOUT-.n62 VOUT-.n61 0.495292
R8148 VOUT-.n120 VOUT-.n104 0.3295
R8149 VOUT-.n120 VOUT-.n119 0.3295
R8150 VOUT-.n119 VOUT-.n118 0.3295
R8151 VOUT-.n118 VOUT-.n117 0.3295
R8152 VOUT-.n117 VOUT-.n116 0.3295
R8153 VOUT-.n116 VOUT-.n115 0.3295
R8154 VOUT-.n115 VOUT-.n114 0.3295
R8155 VOUT-.n114 VOUT-.n113 0.3295
R8156 VOUT-.n113 VOUT-.n112 0.3295
R8157 VOUT-.n112 VOUT-.n111 0.3295
R8158 VOUT-.n111 VOUT-.n110 0.3295
R8159 VOUT-.n123 VOUT-.n121 0.3295
R8160 VOUT-.n123 VOUT-.n122 0.3295
R8161 VOUT-.n126 VOUT-.n124 0.3295
R8162 VOUT-.n126 VOUT-.n125 0.3295
R8163 VOUT-.n129 VOUT-.n127 0.3295
R8164 VOUT-.n129 VOUT-.n128 0.3295
R8165 VOUT-.n132 VOUT-.n130 0.3295
R8166 VOUT-.n132 VOUT-.n131 0.3295
R8167 VOUT-.n135 VOUT-.n133 0.3295
R8168 VOUT-.n135 VOUT-.n134 0.3295
R8169 VOUT-.n138 VOUT-.n136 0.3295
R8170 VOUT-.n138 VOUT-.n137 0.3295
R8171 VOUT-.n141 VOUT-.n139 0.3295
R8172 VOUT-.n141 VOUT-.n140 0.3295
R8173 VOUT-.n144 VOUT-.n142 0.3295
R8174 VOUT-.n144 VOUT-.n143 0.3295
R8175 VOUT-.n147 VOUT-.n145 0.3295
R8176 VOUT-.n147 VOUT-.n146 0.3295
R8177 VOUT-.n150 VOUT-.n148 0.3295
R8178 VOUT-.n150 VOUT-.n149 0.3295
R8179 VOUT-.n72 VOUT-.n71 0.3295
R8180 VOUT-.n85 VOUT-.n73 0.3295
R8181 VOUT-.n85 VOUT-.n84 0.3295
R8182 VOUT-.n84 VOUT-.n83 0.3295
R8183 VOUT-.n83 VOUT-.n82 0.3295
R8184 VOUT-.n82 VOUT-.n81 0.3295
R8185 VOUT-.n81 VOUT-.n80 0.3295
R8186 VOUT-.n80 VOUT-.n79 0.3295
R8187 VOUT-.n79 VOUT-.n78 0.3295
R8188 VOUT-.n78 VOUT-.n77 0.3295
R8189 VOUT-.n77 VOUT-.n76 0.3295
R8190 VOUT-.n76 VOUT-.n75 0.3295
R8191 VOUT-.n75 VOUT-.n74 0.3295
R8192 VOUT-.n88 VOUT-.n86 0.3295
R8193 VOUT-.n88 VOUT-.n87 0.3295
R8194 VOUT-.n91 VOUT-.n89 0.3295
R8195 VOUT-.n91 VOUT-.n90 0.3295
R8196 VOUT-.n94 VOUT-.n92 0.3295
R8197 VOUT-.n94 VOUT-.n93 0.3295
R8198 VOUT-.n97 VOUT-.n95 0.3295
R8199 VOUT-.n97 VOUT-.n96 0.3295
R8200 VOUT-.n100 VOUT-.n98 0.3295
R8201 VOUT-.n100 VOUT-.n99 0.3295
R8202 VOUT-.n103 VOUT-.n101 0.3295
R8203 VOUT-.n103 VOUT-.n102 0.3295
R8204 VOUT-.n152 VOUT-.n151 0.3295
R8205 VOUT-.n153 VOUT-.n152 0.3295
R8206 VOUT-.n113 VOUT-.n109 0.3154
R8207 VOUT-.n191 VOUT-.n183 0.314966
R8208 VOUT-.n154 VOUT-.n153 0.3107
R8209 VOUT-.n114 VOUT-.n108 0.306
R8210 VOUT-.n115 VOUT-.n107 0.306
R8211 VOUT-.n116 VOUT-.n106 0.306
R8212 VOUT-.n117 VOUT-.n105 0.306
R8213 VOUT-.n123 VOUT-.n120 0.2825
R8214 VOUT-.n126 VOUT-.n123 0.2825
R8215 VOUT-.n129 VOUT-.n126 0.2825
R8216 VOUT-.n132 VOUT-.n129 0.2825
R8217 VOUT-.n135 VOUT-.n132 0.2825
R8218 VOUT-.n138 VOUT-.n135 0.2825
R8219 VOUT-.n141 VOUT-.n138 0.2825
R8220 VOUT-.n144 VOUT-.n141 0.2825
R8221 VOUT-.n147 VOUT-.n144 0.2825
R8222 VOUT-.n150 VOUT-.n147 0.2825
R8223 VOUT-.n85 VOUT-.n72 0.2825
R8224 VOUT-.n88 VOUT-.n85 0.2825
R8225 VOUT-.n91 VOUT-.n88 0.2825
R8226 VOUT-.n94 VOUT-.n91 0.2825
R8227 VOUT-.n97 VOUT-.n94 0.2825
R8228 VOUT-.n100 VOUT-.n97 0.2825
R8229 VOUT-.n103 VOUT-.n100 0.2825
R8230 VOUT-.n152 VOUT-.n103 0.2825
R8231 VOUT-.n152 VOUT-.n150 0.2825
R8232 VOUT-.n163 VOUT-.n66 0.2655
R8233 VOUT- VOUT-.n178 0.198417
R8234 VOUT-.n178 VOUT-.n177 0.193208
R8235 VOUT- VOUT-.n197 0.182792
R8236 VOUT-.n155 VOUT-.n154 0.138367
R8237 VOUT-.n189 VOUT-.n183 0.0891864
R8238 VOUT-.n60 VOUT-.n59 0.0577917
R8239 VOUT-.n59 VOUT-.n58 0.0577917
R8240 VOUT-.n58 VOUT-.n21 0.0577917
R8241 VOUT-.n54 VOUT-.n21 0.0577917
R8242 VOUT-.n54 VOUT-.n53 0.0577917
R8243 VOUT-.n53 VOUT-.n52 0.0577917
R8244 VOUT-.n52 VOUT-.n25 0.0577917
R8245 VOUT-.n48 VOUT-.n25 0.0577917
R8246 VOUT-.n61 VOUT-.n18 0.0577917
R8247 VOUT-.n57 VOUT-.n18 0.0577917
R8248 VOUT-.n57 VOUT-.n56 0.0577917
R8249 VOUT-.n56 VOUT-.n55 0.0577917
R8250 VOUT-.n55 VOUT-.n22 0.0577917
R8251 VOUT-.n51 VOUT-.n22 0.0577917
R8252 VOUT-.n51 VOUT-.n50 0.0577917
R8253 VOUT-.n49 VOUT-.n48 0.054517
R8254 VOUT-.n170 VOUT-.n169 0.047375
R8255 VOUT-.n174 VOUT-.n173 0.047375
R8256 VOUT-.n164 VOUT-.n7 0.0421667
R8257 VOUT-.n65 VOUT-.n14 0.0421667
R8258 VOUT-.n196 VOUT-.n195 0.0421667
R8259 VOUT-.n195 VOUT-.n194 0.0421667
R8260 VOUT-.n194 VOUT-.n182 0.0421667
R8261 VOUT-.n190 VOUT-.n182 0.0421667
R8262 VOUT-.n190 VOUT-.n189 0.0421667
R8263 VOUT-.n197 VOUT-.n179 0.0421667
R8264 VOUT-.n193 VOUT-.n179 0.0421667
R8265 VOUT-.n193 VOUT-.n192 0.0421667
R8266 VOUT-.n192 VOUT-.n191 0.0421667
R8267 VOUT-.n15 VOUT-.n14 0.0243161
R8268 VOUT-.n17 VOUT-.n9 0.0243161
R8269 VOUT-.n17 VOUT-.n16 0.0243161
R8270 VOUT-.n15 VOUT-.n11 0.0243161
R8271 VOUT-.n161 VOUT-.n3 0.0217373
R8272 VOUT-.n62 VOUT-.n10 0.0217373
R8273 VOUT-.n16 VOUT-.n10 0.0217373
R8274 VOUT-.n69 VOUT-.n3 0.0217373
R8275 VOUT-.n177 VOUT-.n0 0.0217373
R8276 VOUT-.n174 VOUT-.n0 0.0217373
R8277 VOUT-.n67 VOUT-.n7 0.0217373
R8278 VOUT-.n69 VOUT-.n68 0.0217373
R8279 VOUT-.n12 VOUT-.n9 0.0217373
R8280 VOUT-.n12 VOUT-.n11 0.0217373
R8281 VOUT-.n67 VOUT-.n4 0.0217373
R8282 VOUT-.n68 VOUT-.n4 0.0217373
R8283 VOUT-.n171 VOUT-.n166 0.0217373
R8284 VOUT-.n170 VOUT-.n167 0.0217373
R8285 VOUT-.n173 VOUT-.n167 0.0217373
R8286 VOUT-.n169 VOUT-.n166 0.0217373
R8287 VOUT-.n156 VOUT-.n155 0.0161667
R8288 VOUT-.n159 VOUT-.n156 0.0161667
R8289 VOUT-.n157 VOUT-.n6 0.0161667
R8290 VOUT-.n158 VOUT-.n157 0.0161667
R8291 VOUT-.n158 VOUT-.n70 0.0161667
R8292 VOUT-.n162 VOUT-.n5 0.0134654
R8293 VOUT-.n165 VOUT-.n2 0.0134654
R8294 VOUT-.n163 VOUT-.n162 0.0134654
R8295 VOUT-.n5 VOUT-.n2 0.0134654
R8296 VOUT-.n63 VOUT-.n13 0.0109778
R8297 VOUT-.n66 VOUT-.n8 0.0109778
R8298 VOUT-.n175 VOUT-.n1 0.0109778
R8299 VOUT-.n172 VOUT-.n168 0.0109778
R8300 VOUT-.n64 VOUT-.n63 0.0109778
R8301 VOUT-.n13 VOUT-.n8 0.0109778
R8302 VOUT-.n176 VOUT-.n175 0.0109778
R8303 VOUT-.n168 VOUT-.n1 0.0109778
R8304 VOUT-.n160 VOUT-.n70 0.00872683
R8305 two_stage_opamp_dummy_magic_24_0.cap_res_X two_stage_opamp_dummy_magic_24_0.cap_res_X.t0 49.4254
R8306 two_stage_opamp_dummy_magic_24_0.cap_res_X two_stage_opamp_dummy_magic_24_0.cap_res_X.t16 1.481
R8307 two_stage_opamp_dummy_magic_24_0.cap_res_X.t35 two_stage_opamp_dummy_magic_24_0.cap_res_X.t10 0.1603
R8308 two_stage_opamp_dummy_magic_24_0.cap_res_X.t17 two_stage_opamp_dummy_magic_24_0.cap_res_X.t35 0.1603
R8309 two_stage_opamp_dummy_magic_24_0.cap_res_X.t116 two_stage_opamp_dummy_magic_24_0.cap_res_X.t82 0.1603
R8310 two_stage_opamp_dummy_magic_24_0.cap_res_X.t105 two_stage_opamp_dummy_magic_24_0.cap_res_X.t122 0.1603
R8311 two_stage_opamp_dummy_magic_24_0.cap_res_X.t2 two_stage_opamp_dummy_magic_24_0.cap_res_X.t105 0.1603
R8312 two_stage_opamp_dummy_magic_24_0.cap_res_X.t67 two_stage_opamp_dummy_magic_24_0.cap_res_X.t86 0.1603
R8313 two_stage_opamp_dummy_magic_24_0.cap_res_X.t100 two_stage_opamp_dummy_magic_24_0.cap_res_X.t67 0.1603
R8314 two_stage_opamp_dummy_magic_24_0.cap_res_X.t32 two_stage_opamp_dummy_magic_24_0.cap_res_X.t51 0.1603
R8315 two_stage_opamp_dummy_magic_24_0.cap_res_X.t63 two_stage_opamp_dummy_magic_24_0.cap_res_X.t32 0.1603
R8316 two_stage_opamp_dummy_magic_24_0.cap_res_X.t93 two_stage_opamp_dummy_magic_24_0.cap_res_X.t57 0.1603
R8317 two_stage_opamp_dummy_magic_24_0.cap_res_X.t79 two_stage_opamp_dummy_magic_24_0.cap_res_X.t115 0.1603
R8318 two_stage_opamp_dummy_magic_24_0.cap_res_X.t62 two_stage_opamp_dummy_magic_24_0.cap_res_X.t25 0.1603
R8319 two_stage_opamp_dummy_magic_24_0.cap_res_X.t37 two_stage_opamp_dummy_magic_24_0.cap_res_X.t71 0.1603
R8320 two_stage_opamp_dummy_magic_24_0.cap_res_X.t88 two_stage_opamp_dummy_magic_24_0.cap_res_X.t54 0.1603
R8321 two_stage_opamp_dummy_magic_24_0.cap_res_X.t75 two_stage_opamp_dummy_magic_24_0.cap_res_X.t109 0.1603
R8322 two_stage_opamp_dummy_magic_24_0.cap_res_X.t130 two_stage_opamp_dummy_magic_24_0.cap_res_X.t90 0.1603
R8323 two_stage_opamp_dummy_magic_24_0.cap_res_X.t44 two_stage_opamp_dummy_magic_24_0.cap_res_X.t77 0.1603
R8324 two_stage_opamp_dummy_magic_24_0.cap_res_X.t92 two_stage_opamp_dummy_magic_24_0.cap_res_X.t59 0.1603
R8325 two_stage_opamp_dummy_magic_24_0.cap_res_X.t81 two_stage_opamp_dummy_magic_24_0.cap_res_X.t114 0.1603
R8326 two_stage_opamp_dummy_magic_24_0.cap_res_X.t133 two_stage_opamp_dummy_magic_24_0.cap_res_X.t96 0.1603
R8327 two_stage_opamp_dummy_magic_24_0.cap_res_X.t120 two_stage_opamp_dummy_magic_24_0.cap_res_X.t15 0.1603
R8328 two_stage_opamp_dummy_magic_24_0.cap_res_X.t34 two_stage_opamp_dummy_magic_24_0.cap_res_X.t138 0.1603
R8329 two_stage_opamp_dummy_magic_24_0.cap_res_X.t85 two_stage_opamp_dummy_magic_24_0.cap_res_X.t121 0.1603
R8330 two_stage_opamp_dummy_magic_24_0.cap_res_X.t1 two_stage_opamp_dummy_magic_24_0.cap_res_X.t102 0.1603
R8331 two_stage_opamp_dummy_magic_24_0.cap_res_X.t126 two_stage_opamp_dummy_magic_24_0.cap_res_X.t23 0.1603
R8332 two_stage_opamp_dummy_magic_24_0.cap_res_X.t42 two_stage_opamp_dummy_magic_24_0.cap_res_X.t6 0.1603
R8333 two_stage_opamp_dummy_magic_24_0.cap_res_X.t28 two_stage_opamp_dummy_magic_24_0.cap_res_X.t60 0.1603
R8334 two_stage_opamp_dummy_magic_24_0.cap_res_X.t80 two_stage_opamp_dummy_magic_24_0.cap_res_X.t46 0.1603
R8335 two_stage_opamp_dummy_magic_24_0.cap_res_X.t64 two_stage_opamp_dummy_magic_24_0.cap_res_X.t98 0.1603
R8336 two_stage_opamp_dummy_magic_24_0.cap_res_X.t117 two_stage_opamp_dummy_magic_24_0.cap_res_X.t83 0.1603
R8337 two_stage_opamp_dummy_magic_24_0.cap_res_X.t33 two_stage_opamp_dummy_magic_24_0.cap_res_X.t65 0.1603
R8338 two_stage_opamp_dummy_magic_24_0.cap_res_X.t84 two_stage_opamp_dummy_magic_24_0.cap_res_X.t49 0.1603
R8339 two_stage_opamp_dummy_magic_24_0.cap_res_X.t70 two_stage_opamp_dummy_magic_24_0.cap_res_X.t104 0.1603
R8340 two_stage_opamp_dummy_magic_24_0.cap_res_X.t123 two_stage_opamp_dummy_magic_24_0.cap_res_X.t87 0.1603
R8341 two_stage_opamp_dummy_magic_24_0.cap_res_X.t108 two_stage_opamp_dummy_magic_24_0.cap_res_X.t7 0.1603
R8342 two_stage_opamp_dummy_magic_24_0.cap_res_X.t24 two_stage_opamp_dummy_magic_24_0.cap_res_X.t128 0.1603
R8343 two_stage_opamp_dummy_magic_24_0.cap_res_X.t76 two_stage_opamp_dummy_magic_24_0.cap_res_X.t110 0.1603
R8344 two_stage_opamp_dummy_magic_24_0.cap_res_X.t129 two_stage_opamp_dummy_magic_24_0.cap_res_X.t91 0.1603
R8345 two_stage_opamp_dummy_magic_24_0.cap_res_X.t43 two_stage_opamp_dummy_magic_24_0.cap_res_X.t127 0.1603
R8346 two_stage_opamp_dummy_magic_24_0.cap_res_X.t47 two_stage_opamp_dummy_magic_24_0.cap_res_X.t95 0.1603
R8347 two_stage_opamp_dummy_magic_24_0.cap_res_X.t124 two_stage_opamp_dummy_magic_24_0.cap_res_X.t21 0.1603
R8348 two_stage_opamp_dummy_magic_24_0.cap_res_X.t41 two_stage_opamp_dummy_magic_24_0.cap_res_X.t4 0.1603
R8349 two_stage_opamp_dummy_magic_24_0.cap_res_X.t20 two_stage_opamp_dummy_magic_24_0.cap_res_X.t55 0.1603
R8350 two_stage_opamp_dummy_magic_24_0.cap_res_X.t72 two_stage_opamp_dummy_magic_24_0.cap_res_X.t40 0.1603
R8351 two_stage_opamp_dummy_magic_24_0.cap_res_X.t53 two_stage_opamp_dummy_magic_24_0.cap_res_X.t11 0.1603
R8352 two_stage_opamp_dummy_magic_24_0.cap_res_X.t78 two_stage_opamp_dummy_magic_24_0.cap_res_X.t38 0.1603
R8353 two_stage_opamp_dummy_magic_24_0.cap_res_X.t56 two_stage_opamp_dummy_magic_24_0.cap_res_X.t18 0.1603
R8354 two_stage_opamp_dummy_magic_24_0.cap_res_X.t22 two_stage_opamp_dummy_magic_24_0.cap_res_X.t119 0.1603
R8355 two_stage_opamp_dummy_magic_24_0.cap_res_X.t45 two_stage_opamp_dummy_magic_24_0.cap_res_X.t3 0.1603
R8356 two_stage_opamp_dummy_magic_24_0.cap_res_X.t5 two_stage_opamp_dummy_magic_24_0.cap_res_X.t101 0.1603
R8357 two_stage_opamp_dummy_magic_24_0.cap_res_X.t106 two_stage_opamp_dummy_magic_24_0.cap_res_X.t66 0.1603
R8358 two_stage_opamp_dummy_magic_24_0.cap_res_X.t68 two_stage_opamp_dummy_magic_24_0.cap_res_X.t30 0.1603
R8359 two_stage_opamp_dummy_magic_24_0.cap_res_X.t89 two_stage_opamp_dummy_magic_24_0.cap_res_X.t50 0.1603
R8360 two_stage_opamp_dummy_magic_24_0.cap_res_X.t52 two_stage_opamp_dummy_magic_24_0.cap_res_X.t9 0.1603
R8361 two_stage_opamp_dummy_magic_24_0.cap_res_X.t13 two_stage_opamp_dummy_magic_24_0.cap_res_X.t112 0.1603
R8362 two_stage_opamp_dummy_magic_24_0.cap_res_X.t137 two_stage_opamp_dummy_magic_24_0.cap_res_X.t99 0.1603
R8363 two_stage_opamp_dummy_magic_24_0.cap_res_X.t94 two_stage_opamp_dummy_magic_24_0.cap_res_X.t61 0.1603
R8364 two_stage_opamp_dummy_magic_24_0.cap_res_X.t8 two_stage_opamp_dummy_magic_24_0.cap_res_X.t111 0.1603
R8365 two_stage_opamp_dummy_magic_24_0.cap_res_X.t12 two_stage_opamp_dummy_magic_24_0.cap_res_X.t103 0.1603
R8366 two_stage_opamp_dummy_magic_24_0.cap_res_X.t48 two_stage_opamp_dummy_magic_24_0.cap_res_X.t12 0.1603
R8367 two_stage_opamp_dummy_magic_24_0.cap_res_X.t132 two_stage_opamp_dummy_magic_24_0.cap_res_X.t29 0.1603
R8368 two_stage_opamp_dummy_magic_24_0.cap_res_X.t16 two_stage_opamp_dummy_magic_24_0.cap_res_X.t132 0.1603
R8369 two_stage_opamp_dummy_magic_24_0.cap_res_X.t39 two_stage_opamp_dummy_magic_24_0.cap_res_X.n10 0.159278
R8370 two_stage_opamp_dummy_magic_24_0.cap_res_X.t107 two_stage_opamp_dummy_magic_24_0.cap_res_X.n11 0.159278
R8371 two_stage_opamp_dummy_magic_24_0.cap_res_X.t73 two_stage_opamp_dummy_magic_24_0.cap_res_X.n12 0.159278
R8372 two_stage_opamp_dummy_magic_24_0.cap_res_X.t136 two_stage_opamp_dummy_magic_24_0.cap_res_X.n13 0.159278
R8373 two_stage_opamp_dummy_magic_24_0.cap_res_X.t27 two_stage_opamp_dummy_magic_24_0.cap_res_X.n14 0.159278
R8374 two_stage_opamp_dummy_magic_24_0.cap_res_X.t58 two_stage_opamp_dummy_magic_24_0.cap_res_X.n15 0.159278
R8375 two_stage_opamp_dummy_magic_24_0.cap_res_X.t19 two_stage_opamp_dummy_magic_24_0.cap_res_X.n16 0.159278
R8376 two_stage_opamp_dummy_magic_24_0.cap_res_X.t118 two_stage_opamp_dummy_magic_24_0.cap_res_X.n17 0.159278
R8377 two_stage_opamp_dummy_magic_24_0.cap_res_X.t14 two_stage_opamp_dummy_magic_24_0.cap_res_X.n18 0.159278
R8378 two_stage_opamp_dummy_magic_24_0.cap_res_X.t113 two_stage_opamp_dummy_magic_24_0.cap_res_X.n19 0.159278
R8379 two_stage_opamp_dummy_magic_24_0.cap_res_X.t74 two_stage_opamp_dummy_magic_24_0.cap_res_X.n20 0.159278
R8380 two_stage_opamp_dummy_magic_24_0.cap_res_X.t36 two_stage_opamp_dummy_magic_24_0.cap_res_X.n21 0.159278
R8381 two_stage_opamp_dummy_magic_24_0.cap_res_X.t69 two_stage_opamp_dummy_magic_24_0.cap_res_X.n22 0.159278
R8382 two_stage_opamp_dummy_magic_24_0.cap_res_X.t31 two_stage_opamp_dummy_magic_24_0.cap_res_X.n23 0.159278
R8383 two_stage_opamp_dummy_magic_24_0.cap_res_X.t131 two_stage_opamp_dummy_magic_24_0.cap_res_X.n24 0.159278
R8384 two_stage_opamp_dummy_magic_24_0.cap_res_X.t26 two_stage_opamp_dummy_magic_24_0.cap_res_X.n25 0.159278
R8385 two_stage_opamp_dummy_magic_24_0.cap_res_X.t125 two_stage_opamp_dummy_magic_24_0.cap_res_X.n26 0.159278
R8386 two_stage_opamp_dummy_magic_24_0.cap_res_X.t97 two_stage_opamp_dummy_magic_24_0.cap_res_X.n27 0.159278
R8387 two_stage_opamp_dummy_magic_24_0.cap_res_X.t134 two_stage_opamp_dummy_magic_24_0.cap_res_X.n28 0.159278
R8388 two_stage_opamp_dummy_magic_24_0.cap_res_X.n31 two_stage_opamp_dummy_magic_24_0.cap_res_X.t17 0.1368
R8389 two_stage_opamp_dummy_magic_24_0.cap_res_X.n29 two_stage_opamp_dummy_magic_24_0.cap_res_X.t93 0.1368
R8390 two_stage_opamp_dummy_magic_24_0.cap_res_X.n28 two_stage_opamp_dummy_magic_24_0.cap_res_X.t79 0.1368
R8391 two_stage_opamp_dummy_magic_24_0.cap_res_X.n28 two_stage_opamp_dummy_magic_24_0.cap_res_X.t62 0.1368
R8392 two_stage_opamp_dummy_magic_24_0.cap_res_X.n27 two_stage_opamp_dummy_magic_24_0.cap_res_X.t37 0.1368
R8393 two_stage_opamp_dummy_magic_24_0.cap_res_X.n27 two_stage_opamp_dummy_magic_24_0.cap_res_X.t88 0.1368
R8394 two_stage_opamp_dummy_magic_24_0.cap_res_X.n26 two_stage_opamp_dummy_magic_24_0.cap_res_X.t75 0.1368
R8395 two_stage_opamp_dummy_magic_24_0.cap_res_X.n26 two_stage_opamp_dummy_magic_24_0.cap_res_X.t130 0.1368
R8396 two_stage_opamp_dummy_magic_24_0.cap_res_X.n25 two_stage_opamp_dummy_magic_24_0.cap_res_X.t44 0.1368
R8397 two_stage_opamp_dummy_magic_24_0.cap_res_X.n25 two_stage_opamp_dummy_magic_24_0.cap_res_X.t92 0.1368
R8398 two_stage_opamp_dummy_magic_24_0.cap_res_X.n24 two_stage_opamp_dummy_magic_24_0.cap_res_X.t81 0.1368
R8399 two_stage_opamp_dummy_magic_24_0.cap_res_X.n24 two_stage_opamp_dummy_magic_24_0.cap_res_X.t133 0.1368
R8400 two_stage_opamp_dummy_magic_24_0.cap_res_X.n23 two_stage_opamp_dummy_magic_24_0.cap_res_X.t120 0.1368
R8401 two_stage_opamp_dummy_magic_24_0.cap_res_X.n23 two_stage_opamp_dummy_magic_24_0.cap_res_X.t34 0.1368
R8402 two_stage_opamp_dummy_magic_24_0.cap_res_X.n22 two_stage_opamp_dummy_magic_24_0.cap_res_X.t85 0.1368
R8403 two_stage_opamp_dummy_magic_24_0.cap_res_X.n22 two_stage_opamp_dummy_magic_24_0.cap_res_X.t1 0.1368
R8404 two_stage_opamp_dummy_magic_24_0.cap_res_X.n21 two_stage_opamp_dummy_magic_24_0.cap_res_X.t126 0.1368
R8405 two_stage_opamp_dummy_magic_24_0.cap_res_X.n21 two_stage_opamp_dummy_magic_24_0.cap_res_X.t42 0.1368
R8406 two_stage_opamp_dummy_magic_24_0.cap_res_X.n20 two_stage_opamp_dummy_magic_24_0.cap_res_X.t28 0.1368
R8407 two_stage_opamp_dummy_magic_24_0.cap_res_X.n20 two_stage_opamp_dummy_magic_24_0.cap_res_X.t80 0.1368
R8408 two_stage_opamp_dummy_magic_24_0.cap_res_X.n19 two_stage_opamp_dummy_magic_24_0.cap_res_X.t64 0.1368
R8409 two_stage_opamp_dummy_magic_24_0.cap_res_X.n19 two_stage_opamp_dummy_magic_24_0.cap_res_X.t117 0.1368
R8410 two_stage_opamp_dummy_magic_24_0.cap_res_X.n18 two_stage_opamp_dummy_magic_24_0.cap_res_X.t33 0.1368
R8411 two_stage_opamp_dummy_magic_24_0.cap_res_X.n18 two_stage_opamp_dummy_magic_24_0.cap_res_X.t84 0.1368
R8412 two_stage_opamp_dummy_magic_24_0.cap_res_X.n17 two_stage_opamp_dummy_magic_24_0.cap_res_X.t70 0.1368
R8413 two_stage_opamp_dummy_magic_24_0.cap_res_X.n17 two_stage_opamp_dummy_magic_24_0.cap_res_X.t123 0.1368
R8414 two_stage_opamp_dummy_magic_24_0.cap_res_X.n16 two_stage_opamp_dummy_magic_24_0.cap_res_X.t108 0.1368
R8415 two_stage_opamp_dummy_magic_24_0.cap_res_X.n16 two_stage_opamp_dummy_magic_24_0.cap_res_X.t24 0.1368
R8416 two_stage_opamp_dummy_magic_24_0.cap_res_X.n15 two_stage_opamp_dummy_magic_24_0.cap_res_X.t76 0.1368
R8417 two_stage_opamp_dummy_magic_24_0.cap_res_X.n15 two_stage_opamp_dummy_magic_24_0.cap_res_X.t129 0.1368
R8418 two_stage_opamp_dummy_magic_24_0.cap_res_X.n14 two_stage_opamp_dummy_magic_24_0.cap_res_X.t43 0.1368
R8419 two_stage_opamp_dummy_magic_24_0.cap_res_X.n14 two_stage_opamp_dummy_magic_24_0.cap_res_X.t47 0.1368
R8420 two_stage_opamp_dummy_magic_24_0.cap_res_X.n13 two_stage_opamp_dummy_magic_24_0.cap_res_X.t124 0.1368
R8421 two_stage_opamp_dummy_magic_24_0.cap_res_X.n13 two_stage_opamp_dummy_magic_24_0.cap_res_X.t41 0.1368
R8422 two_stage_opamp_dummy_magic_24_0.cap_res_X.n12 two_stage_opamp_dummy_magic_24_0.cap_res_X.t20 0.1368
R8423 two_stage_opamp_dummy_magic_24_0.cap_res_X.n12 two_stage_opamp_dummy_magic_24_0.cap_res_X.t72 0.1368
R8424 two_stage_opamp_dummy_magic_24_0.cap_res_X.n11 two_stage_opamp_dummy_magic_24_0.cap_res_X.t137 0.1368
R8425 two_stage_opamp_dummy_magic_24_0.cap_res_X.n10 two_stage_opamp_dummy_magic_24_0.cap_res_X.t94 0.1368
R8426 two_stage_opamp_dummy_magic_24_0.cap_res_X.t111 two_stage_opamp_dummy_magic_24_0.cap_res_X.n29 0.1368
R8427 two_stage_opamp_dummy_magic_24_0.cap_res_X.n30 two_stage_opamp_dummy_magic_24_0.cap_res_X.t8 0.1368
R8428 two_stage_opamp_dummy_magic_24_0.cap_res_X.n0 two_stage_opamp_dummy_magic_24_0.cap_res_X.t53 0.114322
R8429 two_stage_opamp_dummy_magic_24_0.cap_res_X.n32 two_stage_opamp_dummy_magic_24_0.cap_res_X.n31 0.1133
R8430 two_stage_opamp_dummy_magic_24_0.cap_res_X.n33 two_stage_opamp_dummy_magic_24_0.cap_res_X.n32 0.1133
R8431 two_stage_opamp_dummy_magic_24_0.cap_res_X.n34 two_stage_opamp_dummy_magic_24_0.cap_res_X.n33 0.1133
R8432 two_stage_opamp_dummy_magic_24_0.cap_res_X.n1 two_stage_opamp_dummy_magic_24_0.cap_res_X.n0 0.1133
R8433 two_stage_opamp_dummy_magic_24_0.cap_res_X.n2 two_stage_opamp_dummy_magic_24_0.cap_res_X.n1 0.1133
R8434 two_stage_opamp_dummy_magic_24_0.cap_res_X.n3 two_stage_opamp_dummy_magic_24_0.cap_res_X.n2 0.1133
R8435 two_stage_opamp_dummy_magic_24_0.cap_res_X.n4 two_stage_opamp_dummy_magic_24_0.cap_res_X.n3 0.1133
R8436 two_stage_opamp_dummy_magic_24_0.cap_res_X.n5 two_stage_opamp_dummy_magic_24_0.cap_res_X.n4 0.1133
R8437 two_stage_opamp_dummy_magic_24_0.cap_res_X.n6 two_stage_opamp_dummy_magic_24_0.cap_res_X.n5 0.1133
R8438 two_stage_opamp_dummy_magic_24_0.cap_res_X.n7 two_stage_opamp_dummy_magic_24_0.cap_res_X.n6 0.1133
R8439 two_stage_opamp_dummy_magic_24_0.cap_res_X.n8 two_stage_opamp_dummy_magic_24_0.cap_res_X.n7 0.1133
R8440 two_stage_opamp_dummy_magic_24_0.cap_res_X.n9 two_stage_opamp_dummy_magic_24_0.cap_res_X.n8 0.1133
R8441 two_stage_opamp_dummy_magic_24_0.cap_res_X.n11 two_stage_opamp_dummy_magic_24_0.cap_res_X.n9 0.1133
R8442 two_stage_opamp_dummy_magic_24_0.cap_res_X.n35 two_stage_opamp_dummy_magic_24_0.cap_res_X.n30 0.1133
R8443 two_stage_opamp_dummy_magic_24_0.cap_res_X.n35 two_stage_opamp_dummy_magic_24_0.cap_res_X.n34 0.1133
R8444 two_stage_opamp_dummy_magic_24_0.cap_res_X.n31 two_stage_opamp_dummy_magic_24_0.cap_res_X.t116 0.00152174
R8445 two_stage_opamp_dummy_magic_24_0.cap_res_X.n32 two_stage_opamp_dummy_magic_24_0.cap_res_X.t2 0.00152174
R8446 two_stage_opamp_dummy_magic_24_0.cap_res_X.n33 two_stage_opamp_dummy_magic_24_0.cap_res_X.t100 0.00152174
R8447 two_stage_opamp_dummy_magic_24_0.cap_res_X.n34 two_stage_opamp_dummy_magic_24_0.cap_res_X.t63 0.00152174
R8448 two_stage_opamp_dummy_magic_24_0.cap_res_X.n0 two_stage_opamp_dummy_magic_24_0.cap_res_X.t78 0.00152174
R8449 two_stage_opamp_dummy_magic_24_0.cap_res_X.n1 two_stage_opamp_dummy_magic_24_0.cap_res_X.t56 0.00152174
R8450 two_stage_opamp_dummy_magic_24_0.cap_res_X.n2 two_stage_opamp_dummy_magic_24_0.cap_res_X.t22 0.00152174
R8451 two_stage_opamp_dummy_magic_24_0.cap_res_X.n3 two_stage_opamp_dummy_magic_24_0.cap_res_X.t45 0.00152174
R8452 two_stage_opamp_dummy_magic_24_0.cap_res_X.n4 two_stage_opamp_dummy_magic_24_0.cap_res_X.t5 0.00152174
R8453 two_stage_opamp_dummy_magic_24_0.cap_res_X.n5 two_stage_opamp_dummy_magic_24_0.cap_res_X.t106 0.00152174
R8454 two_stage_opamp_dummy_magic_24_0.cap_res_X.n6 two_stage_opamp_dummy_magic_24_0.cap_res_X.t68 0.00152174
R8455 two_stage_opamp_dummy_magic_24_0.cap_res_X.n7 two_stage_opamp_dummy_magic_24_0.cap_res_X.t89 0.00152174
R8456 two_stage_opamp_dummy_magic_24_0.cap_res_X.n8 two_stage_opamp_dummy_magic_24_0.cap_res_X.t52 0.00152174
R8457 two_stage_opamp_dummy_magic_24_0.cap_res_X.n9 two_stage_opamp_dummy_magic_24_0.cap_res_X.t13 0.00152174
R8458 two_stage_opamp_dummy_magic_24_0.cap_res_X.n10 two_stage_opamp_dummy_magic_24_0.cap_res_X.t135 0.00152174
R8459 two_stage_opamp_dummy_magic_24_0.cap_res_X.n11 two_stage_opamp_dummy_magic_24_0.cap_res_X.t39 0.00152174
R8460 two_stage_opamp_dummy_magic_24_0.cap_res_X.n12 two_stage_opamp_dummy_magic_24_0.cap_res_X.t107 0.00152174
R8461 two_stage_opamp_dummy_magic_24_0.cap_res_X.n13 two_stage_opamp_dummy_magic_24_0.cap_res_X.t73 0.00152174
R8462 two_stage_opamp_dummy_magic_24_0.cap_res_X.n14 two_stage_opamp_dummy_magic_24_0.cap_res_X.t136 0.00152174
R8463 two_stage_opamp_dummy_magic_24_0.cap_res_X.n15 two_stage_opamp_dummy_magic_24_0.cap_res_X.t27 0.00152174
R8464 two_stage_opamp_dummy_magic_24_0.cap_res_X.n16 two_stage_opamp_dummy_magic_24_0.cap_res_X.t58 0.00152174
R8465 two_stage_opamp_dummy_magic_24_0.cap_res_X.n17 two_stage_opamp_dummy_magic_24_0.cap_res_X.t19 0.00152174
R8466 two_stage_opamp_dummy_magic_24_0.cap_res_X.n18 two_stage_opamp_dummy_magic_24_0.cap_res_X.t118 0.00152174
R8467 two_stage_opamp_dummy_magic_24_0.cap_res_X.n19 two_stage_opamp_dummy_magic_24_0.cap_res_X.t14 0.00152174
R8468 two_stage_opamp_dummy_magic_24_0.cap_res_X.n20 two_stage_opamp_dummy_magic_24_0.cap_res_X.t113 0.00152174
R8469 two_stage_opamp_dummy_magic_24_0.cap_res_X.n21 two_stage_opamp_dummy_magic_24_0.cap_res_X.t74 0.00152174
R8470 two_stage_opamp_dummy_magic_24_0.cap_res_X.n22 two_stage_opamp_dummy_magic_24_0.cap_res_X.t36 0.00152174
R8471 two_stage_opamp_dummy_magic_24_0.cap_res_X.n23 two_stage_opamp_dummy_magic_24_0.cap_res_X.t69 0.00152174
R8472 two_stage_opamp_dummy_magic_24_0.cap_res_X.n24 two_stage_opamp_dummy_magic_24_0.cap_res_X.t31 0.00152174
R8473 two_stage_opamp_dummy_magic_24_0.cap_res_X.n25 two_stage_opamp_dummy_magic_24_0.cap_res_X.t131 0.00152174
R8474 two_stage_opamp_dummy_magic_24_0.cap_res_X.n26 two_stage_opamp_dummy_magic_24_0.cap_res_X.t26 0.00152174
R8475 two_stage_opamp_dummy_magic_24_0.cap_res_X.n27 two_stage_opamp_dummy_magic_24_0.cap_res_X.t125 0.00152174
R8476 two_stage_opamp_dummy_magic_24_0.cap_res_X.n28 two_stage_opamp_dummy_magic_24_0.cap_res_X.t97 0.00152174
R8477 two_stage_opamp_dummy_magic_24_0.cap_res_X.n29 two_stage_opamp_dummy_magic_24_0.cap_res_X.t134 0.00152174
R8478 two_stage_opamp_dummy_magic_24_0.cap_res_X.n30 two_stage_opamp_dummy_magic_24_0.cap_res_X.t48 0.00152174
R8479 two_stage_opamp_dummy_magic_24_0.cap_res_X.t29 two_stage_opamp_dummy_magic_24_0.cap_res_X.n35 0.00152174
R8480 VOUT+.n196 VOUT+.t2 110.386
R8481 VOUT+.n47 VOUT+.n46 34.9935
R8482 VOUT+.n45 VOUT+.n44 34.9935
R8483 VOUT+.n59 VOUT+.n58 34.9935
R8484 VOUT+.n55 VOUT+.n54 34.9935
R8485 VOUT+.n52 VOUT+.n51 34.9935
R8486 VOUT+.n49 VOUT+.n48 34.9935
R8487 VOUT+.n2 VOUT+.n1 9.73997
R8488 VOUT+.n6 VOUT+.n5 9.73997
R8489 VOUT+.n9 VOUT+.n8 9.73997
R8490 VOUT+.n7 VOUT+.n6 6.64633
R8491 VOUT+.n7 VOUT+.n2 6.64633
R8492 VOUT+.n46 VOUT+.t4 6.56717
R8493 VOUT+.n46 VOUT+.t12 6.56717
R8494 VOUT+.n44 VOUT+.t11 6.56717
R8495 VOUT+.n44 VOUT+.t0 6.56717
R8496 VOUT+.n58 VOUT+.t15 6.56717
R8497 VOUT+.n58 VOUT+.t18 6.56717
R8498 VOUT+.n54 VOUT+.t6 6.56717
R8499 VOUT+.n54 VOUT+.t17 6.56717
R8500 VOUT+.n51 VOUT+.t1 6.56717
R8501 VOUT+.n51 VOUT+.t5 6.56717
R8502 VOUT+.n48 VOUT+.t16 6.56717
R8503 VOUT+.n48 VOUT+.t7 6.56717
R8504 VOUT+.n57 VOUT+.n45 6.3755
R8505 VOUT+.n50 VOUT+.n47 6.3755
R8506 VOUT+.n9 VOUT+.n7 6.02133
R8507 VOUT+.n59 VOUT+.n57 5.813
R8508 VOUT+.n56 VOUT+.n55 5.813
R8509 VOUT+.n53 VOUT+.n52 5.813
R8510 VOUT+.n50 VOUT+.n49 5.813
R8511 VOUT+.n60 VOUT+.n36 5.063
R8512 VOUT+.n63 VOUT+.n43 5.063
R8513 VOUT+.n130 VOUT+.t52 4.8295
R8514 VOUT+.n131 VOUT+.t88 4.8295
R8515 VOUT+.n132 VOUT+.t123 4.8295
R8516 VOUT+.n133 VOUT+.t26 4.8295
R8517 VOUT+.n134 VOUT+.t68 4.8295
R8518 VOUT+.n135 VOUT+.t114 4.8295
R8519 VOUT+.n145 VOUT+.t144 4.8295
R8520 VOUT+.n147 VOUT+.t124 4.8295
R8521 VOUT+.n148 VOUT+.t33 4.8295
R8522 VOUT+.n150 VOUT+.t139 4.8295
R8523 VOUT+.n151 VOUT+.t27 4.8295
R8524 VOUT+.n153 VOUT+.t106 4.8295
R8525 VOUT+.n154 VOUT+.t132 4.8295
R8526 VOUT+.n156 VOUT+.t133 4.8295
R8527 VOUT+.n157 VOUT+.t21 4.8295
R8528 VOUT+.n159 VOUT+.t98 4.8295
R8529 VOUT+.n160 VOUT+.t126 4.8295
R8530 VOUT+.n162 VOUT+.t59 4.8295
R8531 VOUT+.n163 VOUT+.t90 4.8295
R8532 VOUT+.n165 VOUT+.t92 4.8295
R8533 VOUT+.n166 VOUT+.t125 4.8295
R8534 VOUT+.n168 VOUT+.t49 4.8295
R8535 VOUT+.n169 VOUT+.t82 4.8295
R8536 VOUT+.n171 VOUT+.t149 4.8295
R8537 VOUT+.n172 VOUT+.t39 4.8295
R8538 VOUT+.n174 VOUT+.t116 4.8295
R8539 VOUT+.n175 VOUT+.t143 4.8295
R8540 VOUT+.n97 VOUT+.t142 4.8295
R8541 VOUT+.n110 VOUT+.t109 4.8295
R8542 VOUT+.n112 VOUT+.t155 4.8295
R8543 VOUT+.n113 VOUT+.t47 4.8295
R8544 VOUT+.n115 VOUT+.t51 4.8295
R8545 VOUT+.n116 VOUT+.t84 4.8295
R8546 VOUT+.n118 VOUT+.t41 4.8295
R8547 VOUT+.n119 VOUT+.t48 4.8295
R8548 VOUT+.n121 VOUT+.t105 4.8295
R8549 VOUT+.n122 VOUT+.t131 4.8295
R8550 VOUT+.n124 VOUT+.t67 4.8295
R8551 VOUT+.n125 VOUT+.t101 4.8295
R8552 VOUT+.n127 VOUT+.t111 4.8295
R8553 VOUT+.n128 VOUT+.t137 4.8295
R8554 VOUT+.n177 VOUT+.t32 4.8295
R8555 VOUT+.n137 VOUT+.t91 4.8154
R8556 VOUT+.n109 VOUT+.t45 4.806
R8557 VOUT+.n108 VOUT+.t85 4.806
R8558 VOUT+.n107 VOUT+.t63 4.806
R8559 VOUT+.n106 VOUT+.t107 4.806
R8560 VOUT+.n105 VOUT+.t138 4.806
R8561 VOUT+.n104 VOUT+.t120 4.806
R8562 VOUT+.n103 VOUT+.t153 4.806
R8563 VOUT+.n102 VOUT+.t56 4.806
R8564 VOUT+.n101 VOUT+.t94 4.806
R8565 VOUT+.n100 VOUT+.t70 4.806
R8566 VOUT+.n99 VOUT+.t112 4.806
R8567 VOUT+.n130 VOUT+.t103 4.5005
R8568 VOUT+.n131 VOUT+.t136 4.5005
R8569 VOUT+.n132 VOUT+.t29 4.5005
R8570 VOUT+.n133 VOUT+.t151 4.5005
R8571 VOUT+.n134 VOUT+.t55 4.5005
R8572 VOUT+.n135 VOUT+.t72 4.5005
R8573 VOUT+.n136 VOUT+.t96 4.5005
R8574 VOUT+.n137 VOUT+.t57 4.5005
R8575 VOUT+.n138 VOUT+.t156 4.5005
R8576 VOUT+.n139 VOUT+.t121 4.5005
R8577 VOUT+.n140 VOUT+.t140 4.5005
R8578 VOUT+.n141 VOUT+.t108 4.5005
R8579 VOUT+.n142 VOUT+.t64 4.5005
R8580 VOUT+.n143 VOUT+.t89 4.5005
R8581 VOUT+.n144 VOUT+.t46 4.5005
R8582 VOUT+.n146 VOUT+.t40 4.5005
R8583 VOUT+.n145 VOUT+.t77 4.5005
R8584 VOUT+.n147 VOUT+.t83 4.5005
R8585 VOUT+.n149 VOUT+.t79 4.5005
R8586 VOUT+.n148 VOUT+.t117 4.5005
R8587 VOUT+.n150 VOUT+.t110 4.5005
R8588 VOUT+.n152 VOUT+.t80 4.5005
R8589 VOUT+.n151 VOUT+.t81 4.5005
R8590 VOUT+.n153 VOUT+.t66 4.5005
R8591 VOUT+.n155 VOUT+.t35 4.5005
R8592 VOUT+.n154 VOUT+.t37 4.5005
R8593 VOUT+.n156 VOUT+.t104 4.5005
R8594 VOUT+.n158 VOUT+.t75 4.5005
R8595 VOUT+.n157 VOUT+.t76 4.5005
R8596 VOUT+.n159 VOUT+.t61 4.5005
R8597 VOUT+.n161 VOUT+.t30 4.5005
R8598 VOUT+.n160 VOUT+.t31 4.5005
R8599 VOUT+.n162 VOUT+.t19 4.5005
R8600 VOUT+.n164 VOUT+.t134 4.5005
R8601 VOUT+.n163 VOUT+.t135 4.5005
R8602 VOUT+.n165 VOUT+.t58 4.5005
R8603 VOUT+.n167 VOUT+.t24 4.5005
R8604 VOUT+.n166 VOUT+.t25 4.5005
R8605 VOUT+.n168 VOUT+.t152 4.5005
R8606 VOUT+.n170 VOUT+.t127 4.5005
R8607 VOUT+.n169 VOUT+.t128 4.5005
R8608 VOUT+.n171 VOUT+.t118 4.5005
R8609 VOUT+.n173 VOUT+.t93 4.5005
R8610 VOUT+.n172 VOUT+.t95 4.5005
R8611 VOUT+.n174 VOUT+.t74 4.5005
R8612 VOUT+.n176 VOUT+.t50 4.5005
R8613 VOUT+.n175 VOUT+.t54 4.5005
R8614 VOUT+.n98 VOUT+.t38 4.5005
R8615 VOUT+.n97 VOUT+.t73 4.5005
R8616 VOUT+.n99 VOUT+.t69 4.5005
R8617 VOUT+.n100 VOUT+.t22 4.5005
R8618 VOUT+.n101 VOUT+.t53 4.5005
R8619 VOUT+.n102 VOUT+.t150 4.5005
R8620 VOUT+.n103 VOUT+.t119 4.5005
R8621 VOUT+.n104 VOUT+.t78 4.5005
R8622 VOUT+.n105 VOUT+.t102 4.5005
R8623 VOUT+.n106 VOUT+.t62 4.5005
R8624 VOUT+.n107 VOUT+.t20 4.5005
R8625 VOUT+.n108 VOUT+.t42 4.5005
R8626 VOUT+.n109 VOUT+.t148 4.5005
R8627 VOUT+.n111 VOUT+.t141 4.5005
R8628 VOUT+.n110 VOUT+.t28 4.5005
R8629 VOUT+.n112 VOUT+.t122 4.5005
R8630 VOUT+.n114 VOUT+.t99 4.5005
R8631 VOUT+.n113 VOUT+.t100 4.5005
R8632 VOUT+.n115 VOUT+.t154 4.5005
R8633 VOUT+.n117 VOUT+.t129 4.5005
R8634 VOUT+.n116 VOUT+.t130 4.5005
R8635 VOUT+.n118 VOUT+.t97 4.5005
R8636 VOUT+.n120 VOUT+.t60 4.5005
R8637 VOUT+.n119 VOUT+.t113 4.5005
R8638 VOUT+.n121 VOUT+.t65 4.5005
R8639 VOUT+.n123 VOUT+.t34 4.5005
R8640 VOUT+.n122 VOUT+.t36 4.5005
R8641 VOUT+.n124 VOUT+.t23 4.5005
R8642 VOUT+.n126 VOUT+.t146 4.5005
R8643 VOUT+.n125 VOUT+.t147 4.5005
R8644 VOUT+.n127 VOUT+.t71 4.5005
R8645 VOUT+.n129 VOUT+.t43 4.5005
R8646 VOUT+.n128 VOUT+.t44 4.5005
R8647 VOUT+.n179 VOUT+.t115 4.5005
R8648 VOUT+.n178 VOUT+.t86 4.5005
R8649 VOUT+.n177 VOUT+.t87 4.5005
R8650 VOUT+.n180 VOUT+.t145 4.5005
R8651 VOUT+.n60 VOUT+.n37 4.5005
R8652 VOUT+.n61 VOUT+.n40 4.5005
R8653 VOUT+.n62 VOUT+.n41 4.5005
R8654 VOUT+.n64 VOUT+.n63 4.5005
R8655 VOUT+.n87 VOUT+.n86 4.5005
R8656 VOUT+.n83 VOUT+.n80 4.5005
R8657 VOUT+.n87 VOUT+.n80 4.5005
R8658 VOUT+.n88 VOUT+.n32 4.5005
R8659 VOUT+.n88 VOUT+.n34 4.5005
R8660 VOUT+.n88 VOUT+.n87 4.5005
R8661 VOUT+.n185 VOUT+.n91 4.5005
R8662 VOUT+.n186 VOUT+.n185 4.5005
R8663 VOUT+.n186 VOUT+.n28 4.5005
R8664 VOUT+.n187 VOUT+.n27 4.5005
R8665 VOUT+.n187 VOUT+.n186 4.5005
R8666 VOUT+.n191 VOUT+.n190 4.5005
R8667 VOUT+.n190 VOUT+.n19 4.5005
R8668 VOUT+.n22 VOUT+.n19 4.5005
R8669 VOUT+.n193 VOUT+.n19 4.5005
R8670 VOUT+.n195 VOUT+.n19 4.5005
R8671 VOUT+.n194 VOUT+.n22 4.5005
R8672 VOUT+.n194 VOUT+.n193 4.5005
R8673 VOUT+.n195 VOUT+.n194 4.5005
R8674 VOUT+.n1 VOUT+.t13 3.42907
R8675 VOUT+.n1 VOUT+.t3 3.42907
R8676 VOUT+.n5 VOUT+.t8 3.42907
R8677 VOUT+.n5 VOUT+.t14 3.42907
R8678 VOUT+.n8 VOUT+.t10 3.42907
R8679 VOUT+.n8 VOUT+.t9 3.42907
R8680 VOUT+.n85 VOUT+.n33 2.26725
R8681 VOUT+.n81 VOUT+.n31 2.24601
R8682 VOUT+.n189 VOUT+.n188 2.24601
R8683 VOUT+.n24 VOUT+.n21 2.24601
R8684 VOUT+.n184 VOUT+.n183 2.24477
R8685 VOUT+.n30 VOUT+.n25 2.24477
R8686 VOUT+.n88 VOUT+.n33 2.24063
R8687 VOUT+.n187 VOUT+.n26 2.24063
R8688 VOUT+.n194 VOUT+.n23 2.24063
R8689 VOUT+.n80 VOUT+.n79 2.24063
R8690 VOUT+.n185 VOUT+.n89 2.24063
R8691 VOUT+.n90 VOUT+.n28 2.24063
R8692 VOUT+.n192 VOUT+.n191 2.24063
R8693 VOUT+.n191 VOUT+.n20 2.24063
R8694 VOUT+.n86 VOUT+.n84 2.23934
R8695 VOUT+.n86 VOUT+.n82 2.23934
R8696 VOUT+.n6 VOUT+.n4 1.83719
R8697 VOUT+.n10 VOUT+.n9 1.72967
R8698 VOUT+.n17 VOUT+.n2 1.72967
R8699 VOUT+.n78 VOUT+.n77 1.5005
R8700 VOUT+.n76 VOUT+.n35 1.5005
R8701 VOUT+.n75 VOUT+.n74 1.5005
R8702 VOUT+.n73 VOUT+.n38 1.5005
R8703 VOUT+.n72 VOUT+.n71 1.5005
R8704 VOUT+.n70 VOUT+.n39 1.5005
R8705 VOUT+.n69 VOUT+.n68 1.5005
R8706 VOUT+.n67 VOUT+.n42 1.5005
R8707 VOUT+.n18 VOUT+.n17 1.5005
R8708 VOUT+.n16 VOUT+.n0 1.5005
R8709 VOUT+.n15 VOUT+.n14 1.5005
R8710 VOUT+.n13 VOUT+.n3 1.5005
R8711 VOUT+.n12 VOUT+.n11 1.5005
R8712 VOUT+.n64 VOUT+.n59 1.313
R8713 VOUT+.n55 VOUT+.n41 1.313
R8714 VOUT+.n52 VOUT+.n40 1.313
R8715 VOUT+.n49 VOUT+.n37 1.313
R8716 VOUT+.n45 VOUT+.n43 1.313
R8717 VOUT+.n47 VOUT+.n36 1.313
R8718 VOUT+.n186 VOUT+.n29 1.1455
R8719 VOUT+.n95 VOUT+.n94 1.13717
R8720 VOUT+.n96 VOUT+.n92 1.13717
R8721 VOUT+.n182 VOUT+.n181 1.13717
R8722 VOUT+.n93 VOUT+.n30 1.13717
R8723 VOUT+.n94 VOUT+.n27 1.13717
R8724 VOUT+.n92 VOUT+.n91 1.13717
R8725 VOUT+.n183 VOUT+.n182 1.13717
R8726 VOUT+.n66 VOUT+.n43 0.715216
R8727 VOUT+.n65 VOUT+.n64 0.65675
R8728 VOUT+.n69 VOUT+.n41 0.65675
R8729 VOUT+.n71 VOUT+.n40 0.65675
R8730 VOUT+.n75 VOUT+.n37 0.65675
R8731 VOUT+.n77 VOUT+.n36 0.65675
R8732 VOUT+.n95 VOUT+.n29 0.585
R8733 VOUT+.n67 VOUT+.n66 0.564601
R8734 VOUT+.n61 VOUT+.n60 0.563
R8735 VOUT+.n62 VOUT+.n61 0.563
R8736 VOUT+.n63 VOUT+.n62 0.563
R8737 VOUT+.n57 VOUT+.n56 0.563
R8738 VOUT+.n56 VOUT+.n53 0.563
R8739 VOUT+.n53 VOUT+.n50 0.563
R8740 VOUT+.n191 VOUT+.n187 0.5455
R8741 VOUT+.n87 VOUT+.n78 0.495292
R8742 VOUT+.n136 VOUT+.n135 0.3295
R8743 VOUT+.n137 VOUT+.n136 0.3295
R8744 VOUT+.n138 VOUT+.n137 0.3295
R8745 VOUT+.n139 VOUT+.n138 0.3295
R8746 VOUT+.n140 VOUT+.n139 0.3295
R8747 VOUT+.n141 VOUT+.n140 0.3295
R8748 VOUT+.n142 VOUT+.n141 0.3295
R8749 VOUT+.n143 VOUT+.n142 0.3295
R8750 VOUT+.n144 VOUT+.n143 0.3295
R8751 VOUT+.n146 VOUT+.n144 0.3295
R8752 VOUT+.n146 VOUT+.n145 0.3295
R8753 VOUT+.n149 VOUT+.n147 0.3295
R8754 VOUT+.n149 VOUT+.n148 0.3295
R8755 VOUT+.n152 VOUT+.n150 0.3295
R8756 VOUT+.n152 VOUT+.n151 0.3295
R8757 VOUT+.n155 VOUT+.n153 0.3295
R8758 VOUT+.n155 VOUT+.n154 0.3295
R8759 VOUT+.n158 VOUT+.n156 0.3295
R8760 VOUT+.n158 VOUT+.n157 0.3295
R8761 VOUT+.n161 VOUT+.n159 0.3295
R8762 VOUT+.n161 VOUT+.n160 0.3295
R8763 VOUT+.n164 VOUT+.n162 0.3295
R8764 VOUT+.n164 VOUT+.n163 0.3295
R8765 VOUT+.n167 VOUT+.n165 0.3295
R8766 VOUT+.n167 VOUT+.n166 0.3295
R8767 VOUT+.n170 VOUT+.n168 0.3295
R8768 VOUT+.n170 VOUT+.n169 0.3295
R8769 VOUT+.n173 VOUT+.n171 0.3295
R8770 VOUT+.n173 VOUT+.n172 0.3295
R8771 VOUT+.n176 VOUT+.n174 0.3295
R8772 VOUT+.n176 VOUT+.n175 0.3295
R8773 VOUT+.n98 VOUT+.n97 0.3295
R8774 VOUT+.n100 VOUT+.n99 0.3295
R8775 VOUT+.n101 VOUT+.n100 0.3295
R8776 VOUT+.n102 VOUT+.n101 0.3295
R8777 VOUT+.n103 VOUT+.n102 0.3295
R8778 VOUT+.n104 VOUT+.n103 0.3295
R8779 VOUT+.n105 VOUT+.n104 0.3295
R8780 VOUT+.n106 VOUT+.n105 0.3295
R8781 VOUT+.n107 VOUT+.n106 0.3295
R8782 VOUT+.n108 VOUT+.n107 0.3295
R8783 VOUT+.n109 VOUT+.n108 0.3295
R8784 VOUT+.n111 VOUT+.n109 0.3295
R8785 VOUT+.n111 VOUT+.n110 0.3295
R8786 VOUT+.n114 VOUT+.n112 0.3295
R8787 VOUT+.n114 VOUT+.n113 0.3295
R8788 VOUT+.n117 VOUT+.n115 0.3295
R8789 VOUT+.n117 VOUT+.n116 0.3295
R8790 VOUT+.n120 VOUT+.n118 0.3295
R8791 VOUT+.n120 VOUT+.n119 0.3295
R8792 VOUT+.n123 VOUT+.n121 0.3295
R8793 VOUT+.n123 VOUT+.n122 0.3295
R8794 VOUT+.n126 VOUT+.n124 0.3295
R8795 VOUT+.n126 VOUT+.n125 0.3295
R8796 VOUT+.n129 VOUT+.n127 0.3295
R8797 VOUT+.n129 VOUT+.n128 0.3295
R8798 VOUT+.n179 VOUT+.n178 0.3295
R8799 VOUT+.n178 VOUT+.n177 0.3295
R8800 VOUT+.n138 VOUT+.n134 0.3154
R8801 VOUT+.n12 VOUT+.n4 0.314966
R8802 VOUT+.n180 VOUT+.n179 0.313833
R8803 VOUT+.n142 VOUT+.n130 0.306
R8804 VOUT+.n141 VOUT+.n131 0.306
R8805 VOUT+.n140 VOUT+.n132 0.306
R8806 VOUT+.n139 VOUT+.n133 0.306
R8807 VOUT+.n149 VOUT+.n146 0.2825
R8808 VOUT+.n152 VOUT+.n149 0.2825
R8809 VOUT+.n155 VOUT+.n152 0.2825
R8810 VOUT+.n158 VOUT+.n155 0.2825
R8811 VOUT+.n161 VOUT+.n158 0.2825
R8812 VOUT+.n164 VOUT+.n161 0.2825
R8813 VOUT+.n167 VOUT+.n164 0.2825
R8814 VOUT+.n170 VOUT+.n167 0.2825
R8815 VOUT+.n173 VOUT+.n170 0.2825
R8816 VOUT+.n176 VOUT+.n173 0.2825
R8817 VOUT+.n111 VOUT+.n98 0.2825
R8818 VOUT+.n114 VOUT+.n111 0.2825
R8819 VOUT+.n117 VOUT+.n114 0.2825
R8820 VOUT+.n120 VOUT+.n117 0.2825
R8821 VOUT+.n123 VOUT+.n120 0.2825
R8822 VOUT+.n126 VOUT+.n123 0.2825
R8823 VOUT+.n129 VOUT+.n126 0.2825
R8824 VOUT+.n178 VOUT+.n129 0.2825
R8825 VOUT+.n178 VOUT+.n176 0.2825
R8826 VOUT+.n185 VOUT+.n88 0.2655
R8827 VOUT+ VOUT+.n196 0.198417
R8828 VOUT+.n196 VOUT+.n195 0.193208
R8829 VOUT+ VOUT+.n18 0.182792
R8830 VOUT+.n181 VOUT+.n180 0.138367
R8831 VOUT+.n10 VOUT+.n4 0.0891864
R8832 VOUT+.n65 VOUT+.n42 0.0577917
R8833 VOUT+.n69 VOUT+.n42 0.0577917
R8834 VOUT+.n70 VOUT+.n69 0.0577917
R8835 VOUT+.n71 VOUT+.n70 0.0577917
R8836 VOUT+.n71 VOUT+.n38 0.0577917
R8837 VOUT+.n75 VOUT+.n38 0.0577917
R8838 VOUT+.n76 VOUT+.n75 0.0577917
R8839 VOUT+.n77 VOUT+.n76 0.0577917
R8840 VOUT+.n68 VOUT+.n67 0.0577917
R8841 VOUT+.n68 VOUT+.n39 0.0577917
R8842 VOUT+.n72 VOUT+.n39 0.0577917
R8843 VOUT+.n73 VOUT+.n72 0.0577917
R8844 VOUT+.n74 VOUT+.n73 0.0577917
R8845 VOUT+.n74 VOUT+.n35 0.0577917
R8846 VOUT+.n78 VOUT+.n35 0.0577917
R8847 VOUT+.n66 VOUT+.n65 0.054517
R8848 VOUT+.n193 VOUT+.n24 0.047375
R8849 VOUT+.n188 VOUT+.n22 0.047375
R8850 VOUT+.n186 VOUT+.n30 0.0421667
R8851 VOUT+.n87 VOUT+.n81 0.0421667
R8852 VOUT+.n11 VOUT+.n10 0.0421667
R8853 VOUT+.n11 VOUT+.n3 0.0421667
R8854 VOUT+.n15 VOUT+.n3 0.0421667
R8855 VOUT+.n16 VOUT+.n15 0.0421667
R8856 VOUT+.n17 VOUT+.n16 0.0421667
R8857 VOUT+.n13 VOUT+.n12 0.0421667
R8858 VOUT+.n14 VOUT+.n13 0.0421667
R8859 VOUT+.n14 VOUT+.n0 0.0421667
R8860 VOUT+.n18 VOUT+.n0 0.0421667
R8861 VOUT+.n82 VOUT+.n81 0.0243161
R8862 VOUT+.n84 VOUT+.n32 0.0243161
R8863 VOUT+.n84 VOUT+.n83 0.0243161
R8864 VOUT+.n82 VOUT+.n34 0.0243161
R8865 VOUT+.n183 VOUT+.n26 0.0217373
R8866 VOUT+.n83 VOUT+.n33 0.0217373
R8867 VOUT+.n91 VOUT+.n26 0.0217373
R8868 VOUT+.n190 VOUT+.n23 0.0217373
R8869 VOUT+.n188 VOUT+.n23 0.0217373
R8870 VOUT+.n89 VOUT+.n30 0.0217373
R8871 VOUT+.n91 VOUT+.n90 0.0217373
R8872 VOUT+.n79 VOUT+.n32 0.0217373
R8873 VOUT+.n79 VOUT+.n34 0.0217373
R8874 VOUT+.n89 VOUT+.n27 0.0217373
R8875 VOUT+.n90 VOUT+.n27 0.0217373
R8876 VOUT+.n195 VOUT+.n20 0.0217373
R8877 VOUT+.n193 VOUT+.n192 0.0217373
R8878 VOUT+.n192 VOUT+.n22 0.0217373
R8879 VOUT+.n24 VOUT+.n20 0.0217373
R8880 VOUT+.n96 VOUT+.n95 0.0161667
R8881 VOUT+.n181 VOUT+.n96 0.0161667
R8882 VOUT+.n94 VOUT+.n93 0.0161667
R8883 VOUT+.n94 VOUT+.n92 0.0161667
R8884 VOUT+.n182 VOUT+.n92 0.0161667
R8885 VOUT+.n184 VOUT+.n28 0.0134654
R8886 VOUT+.n187 VOUT+.n25 0.0134654
R8887 VOUT+.n185 VOUT+.n184 0.0134654
R8888 VOUT+.n28 VOUT+.n25 0.0134654
R8889 VOUT+.n85 VOUT+.n80 0.0109778
R8890 VOUT+.n88 VOUT+.n31 0.0109778
R8891 VOUT+.n189 VOUT+.n19 0.0109778
R8892 VOUT+.n194 VOUT+.n21 0.0109778
R8893 VOUT+.n86 VOUT+.n85 0.0109778
R8894 VOUT+.n80 VOUT+.n31 0.0109778
R8895 VOUT+.n191 VOUT+.n189 0.0109778
R8896 VOUT+.n21 VOUT+.n19 0.0109778
R8897 VOUT+.n93 VOUT+.n29 0.00872683
R8898 two_stage_opamp_dummy_magic_24_0.cap_res_Y two_stage_opamp_dummy_magic_24_0.cap_res_Y.t138 49.4263
R8899 two_stage_opamp_dummy_magic_24_0.cap_res_Y two_stage_opamp_dummy_magic_24_0.cap_res_Y.t68 1.481
R8900 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t79 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t12 0.1603
R8901 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t39 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t123 0.1603
R8902 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t73 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t32 0.1603
R8903 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t75 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t129 0.1603
R8904 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t46 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t17 0.1603
R8905 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t119 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t24 0.1603
R8906 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t90 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t50 0.1603
R8907 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t80 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t135 0.1603
R8908 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t52 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t23 0.1603
R8909 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t125 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t30 0.1603
R8910 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t95 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t58 0.1603
R8911 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t21 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t66 0.1603
R8912 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t137 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t97 0.1603
R8913 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t131 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t31 0.1603
R8914 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t98 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t64 0.1603
R8915 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t28 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t74 0.1603
R8916 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t4 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t107 0.1603
R8917 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t61 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t117 0.1603
R8918 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t38 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t7 0.1603
R8919 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t102 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t13 0.1603
R8920 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t82 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t40 0.1603
R8921 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t69 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t124 0.1603
R8922 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t41 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t11 0.1603
R8923 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t112 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t19 0.1603
R8924 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t85 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t45 0.1603
R8925 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t9 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t55 0.1603
R8926 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t133 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t89 0.1603
R8927 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t120 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t25 0.1603
R8928 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t91 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t51 0.1603
R8929 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t43 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t108 0.1603
R8930 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t115 0.1603
R8931 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t26 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t72 0.1603
R8932 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t2 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t105 0.1603
R8933 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t56 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t109 0.1603
R8934 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t34 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t1 0.1603
R8935 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t128 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t47 0.1603
R8936 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t87 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t44 0.1603
R8937 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t134 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t86 0.1603
R8938 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t103 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t62 0.1603
R8939 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t6 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t100 0.1603
R8940 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t37 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t3 0.1603
R8941 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t78 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t36 0.1603
R8942 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t54 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t18 0.1603
R8943 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t94 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t49 0.1603
R8944 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t136 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t93 0.1603
R8945 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t114 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t71 0.1603
R8946 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t8 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t111 0.1603
R8947 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t83 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t14 0.1603
R8948 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t67 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t110 0.1603
R8949 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t53 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t104 0.1603
R8950 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t92 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t53 0.1603
R8951 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t84 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t42 0.1603
R8952 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t60 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t84 0.1603
R8953 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t99 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t65 0.1603
R8954 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t101 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t88 0.1603
R8955 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t101 0.1603
R8956 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t5 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t130 0.1603
R8957 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t35 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t5 0.1603
R8958 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t127 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t33 0.1603
R8959 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t127 0.1603
R8960 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t20 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t48 0.1603
R8961 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t68 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t20 0.1603
R8962 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t15 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n14 0.159278
R8963 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t57 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n15 0.159278
R8964 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t27 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n16 0.159278
R8965 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t96 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n17 0.159278
R8966 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t122 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n18 0.159278
R8967 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t10 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n19 0.159278
R8968 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t113 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n20 0.159278
R8969 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t70 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n21 0.159278
R8970 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t106 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n22 0.159278
R8971 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t63 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n23 0.159278
R8972 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t29 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n24 0.159278
R8973 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t132 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n25 0.159278
R8974 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t22 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n26 0.159278
R8975 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t126 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n27 0.159278
R8976 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t81 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n28 0.159278
R8977 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t121 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n29 0.159278
R8978 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t76 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n30 0.159278
R8979 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t77 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n31 0.159278
R8980 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t116 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n32 0.159278
R8981 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t79 0.1368
R8982 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t39 0.1368
R8983 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t73 0.1368
R8984 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t75 0.1368
R8985 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t46 0.1368
R8986 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t119 0.1368
R8987 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t90 0.1368
R8988 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t80 0.1368
R8989 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t52 0.1368
R8990 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t125 0.1368
R8991 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t95 0.1368
R8992 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t21 0.1368
R8993 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t137 0.1368
R8994 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t131 0.1368
R8995 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t98 0.1368
R8996 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t28 0.1368
R8997 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t4 0.1368
R8998 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t61 0.1368
R8999 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t38 0.1368
R9000 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t102 0.1368
R9001 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t82 0.1368
R9002 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t69 0.1368
R9003 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t41 0.1368
R9004 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t112 0.1368
R9005 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t85 0.1368
R9006 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t9 0.1368
R9007 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t133 0.1368
R9008 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t120 0.1368
R9009 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t91 0.1368
R9010 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t43 0.1368
R9011 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t59 0.1368
R9012 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t26 0.1368
R9013 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t2 0.1368
R9014 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t56 0.1368
R9015 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t34 0.1368
R9016 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t128 0.1368
R9017 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t83 0.1368
R9018 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t110 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n33 0.1368
R9019 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t67 0.1368
R9020 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t60 0.1368
R9021 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t87 0.114322
R9022 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n4 0.1133
R9023 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n5 0.1133
R9024 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n6 0.1133
R9025 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n7 0.1133
R9026 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n8 0.1133
R9027 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n9 0.1133
R9028 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n10 0.1133
R9029 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n11 0.1133
R9030 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n12 0.1133
R9031 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n13 0.1133
R9032 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n0 0.1133
R9033 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n1 0.1133
R9034 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n2 0.1133
R9035 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n3 0.1133
R9036 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n34 0.1133
R9037 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t134 0.00152174
R9038 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t103 0.00152174
R9039 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t6 0.00152174
R9040 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t37 0.00152174
R9041 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t78 0.00152174
R9042 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t54 0.00152174
R9043 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t94 0.00152174
R9044 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t136 0.00152174
R9045 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t114 0.00152174
R9046 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t8 0.00152174
R9047 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t118 0.00152174
R9048 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t15 0.00152174
R9049 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t57 0.00152174
R9050 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t27 0.00152174
R9051 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t96 0.00152174
R9052 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t122 0.00152174
R9053 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t10 0.00152174
R9054 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t113 0.00152174
R9055 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t70 0.00152174
R9056 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t106 0.00152174
R9057 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t63 0.00152174
R9058 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t29 0.00152174
R9059 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t132 0.00152174
R9060 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t22 0.00152174
R9061 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t126 0.00152174
R9062 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t81 0.00152174
R9063 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t121 0.00152174
R9064 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t76 0.00152174
R9065 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t77 0.00152174
R9066 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t116 0.00152174
R9067 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t92 0.00152174
R9068 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t99 0.00152174
R9069 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t0 0.00152174
R9070 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t35 0.00152174
R9071 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t16 0.00152174
R9072 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t48 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n35 0.00152174
R9073 two_stage_opamp_dummy_magic_24_0.Vb3.n13 two_stage_opamp_dummy_magic_24_0.Vb3.t24 768.551
R9074 two_stage_opamp_dummy_magic_24_0.Vb3.n3 two_stage_opamp_dummy_magic_24_0.Vb3.t8 752.422
R9075 two_stage_opamp_dummy_magic_24_0.Vb3.n2 two_stage_opamp_dummy_magic_24_0.Vb3.t18 752.422
R9076 two_stage_opamp_dummy_magic_24_0.Vb3.n1 two_stage_opamp_dummy_magic_24_0.Vb3.t16 752.422
R9077 two_stage_opamp_dummy_magic_24_0.Vb3.n0 two_stage_opamp_dummy_magic_24_0.Vb3.t22 752.422
R9078 two_stage_opamp_dummy_magic_24_0.Vb3.n3 two_stage_opamp_dummy_magic_24_0.Vb3.t14 752.234
R9079 two_stage_opamp_dummy_magic_24_0.Vb3.n3 two_stage_opamp_dummy_magic_24_0.Vb3.t11 752.234
R9080 two_stage_opamp_dummy_magic_24_0.Vb3.n3 two_stage_opamp_dummy_magic_24_0.Vb3.t17 752.234
R9081 two_stage_opamp_dummy_magic_24_0.Vb3.n2 two_stage_opamp_dummy_magic_24_0.Vb3.t10 752.234
R9082 two_stage_opamp_dummy_magic_24_0.Vb3.n2 two_stage_opamp_dummy_magic_24_0.Vb3.t28 752.234
R9083 two_stage_opamp_dummy_magic_24_0.Vb3.n2 two_stage_opamp_dummy_magic_24_0.Vb3.t12 752.234
R9084 two_stage_opamp_dummy_magic_24_0.Vb3.n1 two_stage_opamp_dummy_magic_24_0.Vb3.t13 752.234
R9085 two_stage_opamp_dummy_magic_24_0.Vb3.n1 two_stage_opamp_dummy_magic_24_0.Vb3.t19 752.234
R9086 two_stage_opamp_dummy_magic_24_0.Vb3.n1 two_stage_opamp_dummy_magic_24_0.Vb3.t21 752.234
R9087 two_stage_opamp_dummy_magic_24_0.Vb3.n0 two_stage_opamp_dummy_magic_24_0.Vb3.t9 752.234
R9088 two_stage_opamp_dummy_magic_24_0.Vb3.n0 two_stage_opamp_dummy_magic_24_0.Vb3.t15 752.234
R9089 two_stage_opamp_dummy_magic_24_0.Vb3.n0 two_stage_opamp_dummy_magic_24_0.Vb3.t20 752.234
R9090 two_stage_opamp_dummy_magic_24_0.Vb3.n4 two_stage_opamp_dummy_magic_24_0.Vb3.t25 747.734
R9091 two_stage_opamp_dummy_magic_24_0.Vb3.n4 two_stage_opamp_dummy_magic_24_0.Vb3.t27 747.734
R9092 two_stage_opamp_dummy_magic_24_0.Vb3.n5 two_stage_opamp_dummy_magic_24_0.Vb3.t23 747.734
R9093 two_stage_opamp_dummy_magic_24_0.Vb3.n5 two_stage_opamp_dummy_magic_24_0.Vb3.t26 747.734
R9094 two_stage_opamp_dummy_magic_24_0.Vb3.n9 two_stage_opamp_dummy_magic_24_0.Vb3.n7 139.639
R9095 two_stage_opamp_dummy_magic_24_0.Vb3.n9 two_stage_opamp_dummy_magic_24_0.Vb3.n8 139.638
R9096 two_stage_opamp_dummy_magic_24_0.Vb3.n11 two_stage_opamp_dummy_magic_24_0.Vb3.n10 134.577
R9097 two_stage_opamp_dummy_magic_24_0.Vb3.n12 two_stage_opamp_dummy_magic_24_0.Vb3.n6 73.3081
R9098 two_stage_opamp_dummy_magic_24_0.Vb3.n12 two_stage_opamp_dummy_magic_24_0.Vb3 68.6255
R9099 two_stage_opamp_dummy_magic_24_0.Vb3 two_stage_opamp_dummy_magic_24_0.Vb3.n11 43.0317
R9100 two_stage_opamp_dummy_magic_24_0.Vb3.n10 two_stage_opamp_dummy_magic_24_0.Vb3.t3 24.0005
R9101 two_stage_opamp_dummy_magic_24_0.Vb3.n10 two_stage_opamp_dummy_magic_24_0.Vb3.t4 24.0005
R9102 two_stage_opamp_dummy_magic_24_0.Vb3.n8 two_stage_opamp_dummy_magic_24_0.Vb3.t7 24.0005
R9103 two_stage_opamp_dummy_magic_24_0.Vb3.n8 two_stage_opamp_dummy_magic_24_0.Vb3.t5 24.0005
R9104 two_stage_opamp_dummy_magic_24_0.Vb3.n7 two_stage_opamp_dummy_magic_24_0.Vb3.t6 24.0005
R9105 two_stage_opamp_dummy_magic_24_0.Vb3.n7 two_stage_opamp_dummy_magic_24_0.Vb3.t0 24.0005
R9106 two_stage_opamp_dummy_magic_24_0.Vb3 two_stage_opamp_dummy_magic_24_0.Vb3.n13 16.3443
R9107 two_stage_opamp_dummy_magic_24_0.Vb3.n6 two_stage_opamp_dummy_magic_24_0.Vb3.t1 11.2576
R9108 two_stage_opamp_dummy_magic_24_0.Vb3.n6 two_stage_opamp_dummy_magic_24_0.Vb3.t2 11.2576
R9109 two_stage_opamp_dummy_magic_24_0.Vb3 two_stage_opamp_dummy_magic_24_0.Vb3.n4 10.7974
R9110 two_stage_opamp_dummy_magic_24_0.Vb3 two_stage_opamp_dummy_magic_24_0.Vb3.n5 10.5161
R9111 two_stage_opamp_dummy_magic_24_0.Vb3.n11 two_stage_opamp_dummy_magic_24_0.Vb3.n9 4.5005
R9112 two_stage_opamp_dummy_magic_24_0.Vb3.n3 two_stage_opamp_dummy_magic_24_0.Vb3.n4 2.251
R9113 two_stage_opamp_dummy_magic_24_0.Vb3.n1 two_stage_opamp_dummy_magic_24_0.Vb3.n5 2.251
R9114 two_stage_opamp_dummy_magic_24_0.Vb3.n3 two_stage_opamp_dummy_magic_24_0.Vb3.n2 1.31025
R9115 two_stage_opamp_dummy_magic_24_0.Vb3.n1 two_stage_opamp_dummy_magic_24_0.Vb3.n0 1.31025
R9116 two_stage_opamp_dummy_magic_24_0.Vb3.n13 two_stage_opamp_dummy_magic_24_0.Vb3.n12 1.21231
R9117 two_stage_opamp_dummy_magic_24_0.VD4.n12 two_stage_opamp_dummy_magic_24_0.VD4.t27 671.418
R9118 two_stage_opamp_dummy_magic_24_0.VD4.n15 two_stage_opamp_dummy_magic_24_0.VD4.t30 671.418
R9119 two_stage_opamp_dummy_magic_24_0.VD4.t28 two_stage_opamp_dummy_magic_24_0.VD4.n13 213.131
R9120 two_stage_opamp_dummy_magic_24_0.VD4.n14 two_stage_opamp_dummy_magic_24_0.VD4.t31 213.131
R9121 two_stage_opamp_dummy_magic_24_0.VD4.t11 two_stage_opamp_dummy_magic_24_0.VD4.t28 146.155
R9122 two_stage_opamp_dummy_magic_24_0.VD4.t36 two_stage_opamp_dummy_magic_24_0.VD4.t11 146.155
R9123 two_stage_opamp_dummy_magic_24_0.VD4.t33 two_stage_opamp_dummy_magic_24_0.VD4.t36 146.155
R9124 two_stage_opamp_dummy_magic_24_0.VD4.t7 two_stage_opamp_dummy_magic_24_0.VD4.t33 146.155
R9125 two_stage_opamp_dummy_magic_24_0.VD4.t15 two_stage_opamp_dummy_magic_24_0.VD4.t7 146.155
R9126 two_stage_opamp_dummy_magic_24_0.VD4.t9 two_stage_opamp_dummy_magic_24_0.VD4.t15 146.155
R9127 two_stage_opamp_dummy_magic_24_0.VD4.t4 two_stage_opamp_dummy_magic_24_0.VD4.t9 146.155
R9128 two_stage_opamp_dummy_magic_24_0.VD4.t0 two_stage_opamp_dummy_magic_24_0.VD4.t4 146.155
R9129 two_stage_opamp_dummy_magic_24_0.VD4.t2 two_stage_opamp_dummy_magic_24_0.VD4.t0 146.155
R9130 two_stage_opamp_dummy_magic_24_0.VD4.t13 two_stage_opamp_dummy_magic_24_0.VD4.t2 146.155
R9131 two_stage_opamp_dummy_magic_24_0.VD4.t31 two_stage_opamp_dummy_magic_24_0.VD4.t13 146.155
R9132 two_stage_opamp_dummy_magic_24_0.VD4.n13 two_stage_opamp_dummy_magic_24_0.VD4.t29 76.2576
R9133 two_stage_opamp_dummy_magic_24_0.VD4.n14 two_stage_opamp_dummy_magic_24_0.VD4.t32 76.2576
R9134 two_stage_opamp_dummy_magic_24_0.VD4.n3 two_stage_opamp_dummy_magic_24_0.VD4.n2 68.0435
R9135 two_stage_opamp_dummy_magic_24_0.VD4.n5 two_stage_opamp_dummy_magic_24_0.VD4.n4 68.0435
R9136 two_stage_opamp_dummy_magic_24_0.VD4.n7 two_stage_opamp_dummy_magic_24_0.VD4.n6 68.0435
R9137 two_stage_opamp_dummy_magic_24_0.VD4.n9 two_stage_opamp_dummy_magic_24_0.VD4.n8 68.0435
R9138 two_stage_opamp_dummy_magic_24_0.VD4.n11 two_stage_opamp_dummy_magic_24_0.VD4.n10 68.0435
R9139 two_stage_opamp_dummy_magic_24_0.VD4.n19 two_stage_opamp_dummy_magic_24_0.VD4.n18 66.0338
R9140 two_stage_opamp_dummy_magic_24_0.VD4.n32 two_stage_opamp_dummy_magic_24_0.VD4.n31 66.0338
R9141 two_stage_opamp_dummy_magic_24_0.VD4.n29 two_stage_opamp_dummy_magic_24_0.VD4.n28 66.0338
R9142 two_stage_opamp_dummy_magic_24_0.VD4.n25 two_stage_opamp_dummy_magic_24_0.VD4.n24 66.0338
R9143 two_stage_opamp_dummy_magic_24_0.VD4.n22 two_stage_opamp_dummy_magic_24_0.VD4.n21 66.0338
R9144 two_stage_opamp_dummy_magic_24_0.VD4.n35 two_stage_opamp_dummy_magic_24_0.VD4.n34 66.0338
R9145 two_stage_opamp_dummy_magic_24_0.VD4.n18 two_stage_opamp_dummy_magic_24_0.VD4.t35 11.2576
R9146 two_stage_opamp_dummy_magic_24_0.VD4.n18 two_stage_opamp_dummy_magic_24_0.VD4.t20 11.2576
R9147 two_stage_opamp_dummy_magic_24_0.VD4.n31 two_stage_opamp_dummy_magic_24_0.VD4.t24 11.2576
R9148 two_stage_opamp_dummy_magic_24_0.VD4.n31 two_stage_opamp_dummy_magic_24_0.VD4.t22 11.2576
R9149 two_stage_opamp_dummy_magic_24_0.VD4.n28 two_stage_opamp_dummy_magic_24_0.VD4.t19 11.2576
R9150 two_stage_opamp_dummy_magic_24_0.VD4.n28 two_stage_opamp_dummy_magic_24_0.VD4.t21 11.2576
R9151 two_stage_opamp_dummy_magic_24_0.VD4.n24 two_stage_opamp_dummy_magic_24_0.VD4.t25 11.2576
R9152 two_stage_opamp_dummy_magic_24_0.VD4.n24 two_stage_opamp_dummy_magic_24_0.VD4.t18 11.2576
R9153 two_stage_opamp_dummy_magic_24_0.VD4.n21 two_stage_opamp_dummy_magic_24_0.VD4.t23 11.2576
R9154 two_stage_opamp_dummy_magic_24_0.VD4.n21 two_stage_opamp_dummy_magic_24_0.VD4.t17 11.2576
R9155 two_stage_opamp_dummy_magic_24_0.VD4.n2 two_stage_opamp_dummy_magic_24_0.VD4.t3 11.2576
R9156 two_stage_opamp_dummy_magic_24_0.VD4.n2 two_stage_opamp_dummy_magic_24_0.VD4.t14 11.2576
R9157 two_stage_opamp_dummy_magic_24_0.VD4.n4 two_stage_opamp_dummy_magic_24_0.VD4.t5 11.2576
R9158 two_stage_opamp_dummy_magic_24_0.VD4.n4 two_stage_opamp_dummy_magic_24_0.VD4.t1 11.2576
R9159 two_stage_opamp_dummy_magic_24_0.VD4.n6 two_stage_opamp_dummy_magic_24_0.VD4.t16 11.2576
R9160 two_stage_opamp_dummy_magic_24_0.VD4.n6 two_stage_opamp_dummy_magic_24_0.VD4.t10 11.2576
R9161 two_stage_opamp_dummy_magic_24_0.VD4.n8 two_stage_opamp_dummy_magic_24_0.VD4.t34 11.2576
R9162 two_stage_opamp_dummy_magic_24_0.VD4.n8 two_stage_opamp_dummy_magic_24_0.VD4.t8 11.2576
R9163 two_stage_opamp_dummy_magic_24_0.VD4.n10 two_stage_opamp_dummy_magic_24_0.VD4.t12 11.2576
R9164 two_stage_opamp_dummy_magic_24_0.VD4.n10 two_stage_opamp_dummy_magic_24_0.VD4.t37 11.2576
R9165 two_stage_opamp_dummy_magic_24_0.VD4.t26 two_stage_opamp_dummy_magic_24_0.VD4.n35 11.2576
R9166 two_stage_opamp_dummy_magic_24_0.VD4.n35 two_stage_opamp_dummy_magic_24_0.VD4.t6 11.2576
R9167 two_stage_opamp_dummy_magic_24_0.VD4.n20 two_stage_opamp_dummy_magic_24_0.VD4.n19 5.91717
R9168 two_stage_opamp_dummy_magic_24_0.VD4.n34 two_stage_opamp_dummy_magic_24_0.VD4.n33 5.91717
R9169 two_stage_opamp_dummy_magic_24_0.VD4.n33 two_stage_opamp_dummy_magic_24_0.VD4.n32 5.29217
R9170 two_stage_opamp_dummy_magic_24_0.VD4.n30 two_stage_opamp_dummy_magic_24_0.VD4.n29 5.29217
R9171 two_stage_opamp_dummy_magic_24_0.VD4.n25 two_stage_opamp_dummy_magic_24_0.VD4.n1 5.29217
R9172 two_stage_opamp_dummy_magic_24_0.VD4.n22 two_stage_opamp_dummy_magic_24_0.VD4.n20 5.29217
R9173 two_stage_opamp_dummy_magic_24_0.VD4.n34 two_stage_opamp_dummy_magic_24_0.VD4.n0 2.07265
R9174 two_stage_opamp_dummy_magic_24_0.VD4.n19 two_stage_opamp_dummy_magic_24_0.VD4.n17 2.01265
R9175 two_stage_opamp_dummy_magic_24_0.VD4.n32 two_stage_opamp_dummy_magic_24_0.VD4.n0 2.01015
R9176 two_stage_opamp_dummy_magic_24_0.VD4.n29 two_stage_opamp_dummy_magic_24_0.VD4.n27 2.01015
R9177 two_stage_opamp_dummy_magic_24_0.VD4.n26 two_stage_opamp_dummy_magic_24_0.VD4.n25 2.01015
R9178 two_stage_opamp_dummy_magic_24_0.VD4.n23 two_stage_opamp_dummy_magic_24_0.VD4.n22 2.01015
R9179 two_stage_opamp_dummy_magic_24_0.VD4.n15 two_stage_opamp_dummy_magic_24_0.VD4.n14 1.90883
R9180 two_stage_opamp_dummy_magic_24_0.VD4.n13 two_stage_opamp_dummy_magic_24_0.VD4.n12 1.90883
R9181 two_stage_opamp_dummy_magic_24_0.VD4.n12 two_stage_opamp_dummy_magic_24_0.VD4.n11 1.19765
R9182 two_stage_opamp_dummy_magic_24_0.VD4.n16 two_stage_opamp_dummy_magic_24_0.VD4.n15 1.13515
R9183 two_stage_opamp_dummy_magic_24_0.VD4.n20 two_stage_opamp_dummy_magic_24_0.VD4.n1 0.6255
R9184 two_stage_opamp_dummy_magic_24_0.VD4.n30 two_stage_opamp_dummy_magic_24_0.VD4.n1 0.6255
R9185 two_stage_opamp_dummy_magic_24_0.VD4.n33 two_stage_opamp_dummy_magic_24_0.VD4.n30 0.6255
R9186 two_stage_opamp_dummy_magic_24_0.VD4.n17 two_stage_opamp_dummy_magic_24_0.VD4.n16 0.393729
R9187 two_stage_opamp_dummy_magic_24_0.VD4.n11 two_stage_opamp_dummy_magic_24_0.VD4.n9 0.063
R9188 two_stage_opamp_dummy_magic_24_0.VD4.n9 two_stage_opamp_dummy_magic_24_0.VD4.n7 0.063
R9189 two_stage_opamp_dummy_magic_24_0.VD4.n7 two_stage_opamp_dummy_magic_24_0.VD4.n5 0.063
R9190 two_stage_opamp_dummy_magic_24_0.VD4.n5 two_stage_opamp_dummy_magic_24_0.VD4.n3 0.063
R9191 two_stage_opamp_dummy_magic_24_0.VD4.n16 two_stage_opamp_dummy_magic_24_0.VD4.n3 0.063
R9192 two_stage_opamp_dummy_magic_24_0.VD4.n23 two_stage_opamp_dummy_magic_24_0.VD4.n17 0.063
R9193 two_stage_opamp_dummy_magic_24_0.VD4.n26 two_stage_opamp_dummy_magic_24_0.VD4.n23 0.063
R9194 two_stage_opamp_dummy_magic_24_0.VD4.n27 two_stage_opamp_dummy_magic_24_0.VD4.n26 0.063
R9195 two_stage_opamp_dummy_magic_24_0.VD4.n27 two_stage_opamp_dummy_magic_24_0.VD4.n0 0.063
R9196 two_stage_opamp_dummy_magic_24_0.VD3.n21 two_stage_opamp_dummy_magic_24_0.VD3.t15 671.418
R9197 two_stage_opamp_dummy_magic_24_0.VD3.n18 two_stage_opamp_dummy_magic_24_0.VD3.t12 671.418
R9198 two_stage_opamp_dummy_magic_24_0.VD3.n20 two_stage_opamp_dummy_magic_24_0.VD3.t16 213.131
R9199 two_stage_opamp_dummy_magic_24_0.VD3.t13 two_stage_opamp_dummy_magic_24_0.VD3.n19 213.131
R9200 two_stage_opamp_dummy_magic_24_0.VD3.t16 two_stage_opamp_dummy_magic_24_0.VD3.t0 146.155
R9201 two_stage_opamp_dummy_magic_24_0.VD3.t0 two_stage_opamp_dummy_magic_24_0.VD3.t6 146.155
R9202 two_stage_opamp_dummy_magic_24_0.VD3.t6 two_stage_opamp_dummy_magic_24_0.VD3.t2 146.155
R9203 two_stage_opamp_dummy_magic_24_0.VD3.t2 two_stage_opamp_dummy_magic_24_0.VD3.t18 146.155
R9204 two_stage_opamp_dummy_magic_24_0.VD3.t18 two_stage_opamp_dummy_magic_24_0.VD3.t10 146.155
R9205 two_stage_opamp_dummy_magic_24_0.VD3.t10 two_stage_opamp_dummy_magic_24_0.VD3.t34 146.155
R9206 two_stage_opamp_dummy_magic_24_0.VD3.t34 two_stage_opamp_dummy_magic_24_0.VD3.t32 146.155
R9207 two_stage_opamp_dummy_magic_24_0.VD3.t32 two_stage_opamp_dummy_magic_24_0.VD3.t8 146.155
R9208 two_stage_opamp_dummy_magic_24_0.VD3.t8 two_stage_opamp_dummy_magic_24_0.VD3.t36 146.155
R9209 two_stage_opamp_dummy_magic_24_0.VD3.t36 two_stage_opamp_dummy_magic_24_0.VD3.t4 146.155
R9210 two_stage_opamp_dummy_magic_24_0.VD3.t4 two_stage_opamp_dummy_magic_24_0.VD3.t13 146.155
R9211 two_stage_opamp_dummy_magic_24_0.VD3.n20 two_stage_opamp_dummy_magic_24_0.VD3.t17 76.2576
R9212 two_stage_opamp_dummy_magic_24_0.VD3.n19 two_stage_opamp_dummy_magic_24_0.VD3.t14 76.2576
R9213 two_stage_opamp_dummy_magic_24_0.VD3.n17 two_stage_opamp_dummy_magic_24_0.VD3.n16 68.0435
R9214 two_stage_opamp_dummy_magic_24_0.VD3.n15 two_stage_opamp_dummy_magic_24_0.VD3.n14 68.0435
R9215 two_stage_opamp_dummy_magic_24_0.VD3.n13 two_stage_opamp_dummy_magic_24_0.VD3.n12 68.0435
R9216 two_stage_opamp_dummy_magic_24_0.VD3.n11 two_stage_opamp_dummy_magic_24_0.VD3.n10 68.0435
R9217 two_stage_opamp_dummy_magic_24_0.VD3.n9 two_stage_opamp_dummy_magic_24_0.VD3.n8 68.0435
R9218 two_stage_opamp_dummy_magic_24_0.VD3.n2 two_stage_opamp_dummy_magic_24_0.VD3.n1 66.0338
R9219 two_stage_opamp_dummy_magic_24_0.VD3.n31 two_stage_opamp_dummy_magic_24_0.VD3.n30 66.0338
R9220 two_stage_opamp_dummy_magic_24_0.VD3.n27 two_stage_opamp_dummy_magic_24_0.VD3.n26 66.0338
R9221 two_stage_opamp_dummy_magic_24_0.VD3.n24 two_stage_opamp_dummy_magic_24_0.VD3.n23 66.0338
R9222 two_stage_opamp_dummy_magic_24_0.VD3.n5 two_stage_opamp_dummy_magic_24_0.VD3.n4 66.0338
R9223 two_stage_opamp_dummy_magic_24_0.VD3.n35 two_stage_opamp_dummy_magic_24_0.VD3.n34 66.0338
R9224 two_stage_opamp_dummy_magic_24_0.VD3.n1 two_stage_opamp_dummy_magic_24_0.VD3.t20 11.2576
R9225 two_stage_opamp_dummy_magic_24_0.VD3.n1 two_stage_opamp_dummy_magic_24_0.VD3.t24 11.2576
R9226 two_stage_opamp_dummy_magic_24_0.VD3.n16 two_stage_opamp_dummy_magic_24_0.VD3.t37 11.2576
R9227 two_stage_opamp_dummy_magic_24_0.VD3.n16 two_stage_opamp_dummy_magic_24_0.VD3.t5 11.2576
R9228 two_stage_opamp_dummy_magic_24_0.VD3.n14 two_stage_opamp_dummy_magic_24_0.VD3.t33 11.2576
R9229 two_stage_opamp_dummy_magic_24_0.VD3.n14 two_stage_opamp_dummy_magic_24_0.VD3.t9 11.2576
R9230 two_stage_opamp_dummy_magic_24_0.VD3.n12 two_stage_opamp_dummy_magic_24_0.VD3.t11 11.2576
R9231 two_stage_opamp_dummy_magic_24_0.VD3.n12 two_stage_opamp_dummy_magic_24_0.VD3.t35 11.2576
R9232 two_stage_opamp_dummy_magic_24_0.VD3.n10 two_stage_opamp_dummy_magic_24_0.VD3.t3 11.2576
R9233 two_stage_opamp_dummy_magic_24_0.VD3.n10 two_stage_opamp_dummy_magic_24_0.VD3.t19 11.2576
R9234 two_stage_opamp_dummy_magic_24_0.VD3.n8 two_stage_opamp_dummy_magic_24_0.VD3.t1 11.2576
R9235 two_stage_opamp_dummy_magic_24_0.VD3.n8 two_stage_opamp_dummy_magic_24_0.VD3.t7 11.2576
R9236 two_stage_opamp_dummy_magic_24_0.VD3.n30 two_stage_opamp_dummy_magic_24_0.VD3.t23 11.2576
R9237 two_stage_opamp_dummy_magic_24_0.VD3.n30 two_stage_opamp_dummy_magic_24_0.VD3.t25 11.2576
R9238 two_stage_opamp_dummy_magic_24_0.VD3.n26 two_stage_opamp_dummy_magic_24_0.VD3.t27 11.2576
R9239 two_stage_opamp_dummy_magic_24_0.VD3.n26 two_stage_opamp_dummy_magic_24_0.VD3.t30 11.2576
R9240 two_stage_opamp_dummy_magic_24_0.VD3.n23 two_stage_opamp_dummy_magic_24_0.VD3.t28 11.2576
R9241 two_stage_opamp_dummy_magic_24_0.VD3.n23 two_stage_opamp_dummy_magic_24_0.VD3.t21 11.2576
R9242 two_stage_opamp_dummy_magic_24_0.VD3.n4 two_stage_opamp_dummy_magic_24_0.VD3.t26 11.2576
R9243 two_stage_opamp_dummy_magic_24_0.VD3.n4 two_stage_opamp_dummy_magic_24_0.VD3.t29 11.2576
R9244 two_stage_opamp_dummy_magic_24_0.VD3.t31 two_stage_opamp_dummy_magic_24_0.VD3.n35 11.2576
R9245 two_stage_opamp_dummy_magic_24_0.VD3.n35 two_stage_opamp_dummy_magic_24_0.VD3.t22 11.2576
R9246 two_stage_opamp_dummy_magic_24_0.VD3.n24 two_stage_opamp_dummy_magic_24_0.VD3.n7 5.91717
R9247 two_stage_opamp_dummy_magic_24_0.VD3.n6 two_stage_opamp_dummy_magic_24_0.VD3.n2 5.91717
R9248 two_stage_opamp_dummy_magic_24_0.VD3.n27 two_stage_opamp_dummy_magic_24_0.VD3.n7 5.29217
R9249 two_stage_opamp_dummy_magic_24_0.VD3.n32 two_stage_opamp_dummy_magic_24_0.VD3.n31 5.29217
R9250 two_stage_opamp_dummy_magic_24_0.VD3.n6 two_stage_opamp_dummy_magic_24_0.VD3.n5 5.29217
R9251 two_stage_opamp_dummy_magic_24_0.VD3.n34 two_stage_opamp_dummy_magic_24_0.VD3.n33 5.29217
R9252 two_stage_opamp_dummy_magic_24_0.VD3.n3 two_stage_opamp_dummy_magic_24_0.VD3.n2 2.07515
R9253 two_stage_opamp_dummy_magic_24_0.VD3.n28 two_stage_opamp_dummy_magic_24_0.VD3.n27 2.01015
R9254 two_stage_opamp_dummy_magic_24_0.VD3.n25 two_stage_opamp_dummy_magic_24_0.VD3.n24 2.01015
R9255 two_stage_opamp_dummy_magic_24_0.VD3.n31 two_stage_opamp_dummy_magic_24_0.VD3.n29 2.01015
R9256 two_stage_opamp_dummy_magic_24_0.VD3.n34 two_stage_opamp_dummy_magic_24_0.VD3.n0 2.01015
R9257 two_stage_opamp_dummy_magic_24_0.VD3.n5 two_stage_opamp_dummy_magic_24_0.VD3.n3 2.01015
R9258 two_stage_opamp_dummy_magic_24_0.VD3.n19 two_stage_opamp_dummy_magic_24_0.VD3.n18 1.90883
R9259 two_stage_opamp_dummy_magic_24_0.VD3.n21 two_stage_opamp_dummy_magic_24_0.VD3.n20 1.90883
R9260 two_stage_opamp_dummy_magic_24_0.VD3.n18 two_stage_opamp_dummy_magic_24_0.VD3.n17 1.19765
R9261 two_stage_opamp_dummy_magic_24_0.VD3.n22 two_stage_opamp_dummy_magic_24_0.VD3.n21 1.13515
R9262 two_stage_opamp_dummy_magic_24_0.VD3.n32 two_stage_opamp_dummy_magic_24_0.VD3.n7 0.6255
R9263 two_stage_opamp_dummy_magic_24_0.VD3.n33 two_stage_opamp_dummy_magic_24_0.VD3.n32 0.6255
R9264 two_stage_opamp_dummy_magic_24_0.VD3.n33 two_stage_opamp_dummy_magic_24_0.VD3.n6 0.6255
R9265 two_stage_opamp_dummy_magic_24_0.VD3.n25 two_stage_opamp_dummy_magic_24_0.VD3.n22 0.393729
R9266 two_stage_opamp_dummy_magic_24_0.VD3.n3 two_stage_opamp_dummy_magic_24_0.VD3.n0 0.063
R9267 two_stage_opamp_dummy_magic_24_0.VD3.n29 two_stage_opamp_dummy_magic_24_0.VD3.n0 0.063
R9268 two_stage_opamp_dummy_magic_24_0.VD3.n29 two_stage_opamp_dummy_magic_24_0.VD3.n28 0.063
R9269 two_stage_opamp_dummy_magic_24_0.VD3.n28 two_stage_opamp_dummy_magic_24_0.VD3.n25 0.063
R9270 two_stage_opamp_dummy_magic_24_0.VD3.n22 two_stage_opamp_dummy_magic_24_0.VD3.n9 0.063
R9271 two_stage_opamp_dummy_magic_24_0.VD3.n11 two_stage_opamp_dummy_magic_24_0.VD3.n9 0.063
R9272 two_stage_opamp_dummy_magic_24_0.VD3.n13 two_stage_opamp_dummy_magic_24_0.VD3.n11 0.063
R9273 two_stage_opamp_dummy_magic_24_0.VD3.n15 two_stage_opamp_dummy_magic_24_0.VD3.n13 0.063
R9274 two_stage_opamp_dummy_magic_24_0.VD3.n17 two_stage_opamp_dummy_magic_24_0.VD3.n15 0.063
R9275 VIN+.n0 VIN+.t8 1097.62
R9276 VIN+ VIN+.n9 433.019
R9277 VIN+.n9 VIN+.t4 273.134
R9278 VIN+.n0 VIN+.t6 273.134
R9279 VIN+.n8 VIN+.t0 273.134
R9280 VIN+.n7 VIN+.t3 273.134
R9281 VIN+.n6 VIN+.t10 273.134
R9282 VIN+.n5 VIN+.t2 273.134
R9283 VIN+.n4 VIN+.t7 273.134
R9284 VIN+.n3 VIN+.t5 273.134
R9285 VIN+.n2 VIN+.t9 273.134
R9286 VIN+.n1 VIN+.t1 273.134
R9287 VIN+.n1 VIN+.n0 176.733
R9288 VIN+.n2 VIN+.n1 176.733
R9289 VIN+.n3 VIN+.n2 176.733
R9290 VIN+.n4 VIN+.n3 176.733
R9291 VIN+.n5 VIN+.n4 176.733
R9292 VIN+.n6 VIN+.n5 176.733
R9293 VIN+.n7 VIN+.n6 176.733
R9294 VIN+.n8 VIN+.n7 176.733
R9295 VIN+.n9 VIN+.n8 176.733
R9296 two_stage_opamp_dummy_magic_24_0.V_source.n29 two_stage_opamp_dummy_magic_24_0.V_source.n28 49.3505
R9297 two_stage_opamp_dummy_magic_24_0.V_source.n27 two_stage_opamp_dummy_magic_24_0.V_source.n26 49.3505
R9298 two_stage_opamp_dummy_magic_24_0.V_source.n19 two_stage_opamp_dummy_magic_24_0.V_source.n18 49.3505
R9299 two_stage_opamp_dummy_magic_24_0.V_source.n35 two_stage_opamp_dummy_magic_24_0.V_source.n34 49.3505
R9300 two_stage_opamp_dummy_magic_24_0.V_source.n32 two_stage_opamp_dummy_magic_24_0.V_source.n31 49.3505
R9301 two_stage_opamp_dummy_magic_24_0.V_source.n44 two_stage_opamp_dummy_magic_24_0.V_source.n43 49.3505
R9302 two_stage_opamp_dummy_magic_24_0.V_source.n40 two_stage_opamp_dummy_magic_24_0.V_source.n39 49.3505
R9303 two_stage_opamp_dummy_magic_24_0.V_source.n38 two_stage_opamp_dummy_magic_24_0.V_source.n37 49.3505
R9304 two_stage_opamp_dummy_magic_24_0.V_source.n23 two_stage_opamp_dummy_magic_24_0.V_source.n22 49.3505
R9305 two_stage_opamp_dummy_magic_24_0.V_source.n21 two_stage_opamp_dummy_magic_24_0.V_source.n20 49.3505
R9306 two_stage_opamp_dummy_magic_24_0.V_source.n47 two_stage_opamp_dummy_magic_24_0.V_source.n46 32.3838
R9307 two_stage_opamp_dummy_magic_24_0.V_source.n9 two_stage_opamp_dummy_magic_24_0.V_source.n48 32.3838
R9308 two_stage_opamp_dummy_magic_24_0.V_source.n8 two_stage_opamp_dummy_magic_24_0.V_source.n10 32.3838
R9309 two_stage_opamp_dummy_magic_24_0.V_source.n14 two_stage_opamp_dummy_magic_24_0.V_source.n13 32.3838
R9310 two_stage_opamp_dummy_magic_24_0.V_source.n12 two_stage_opamp_dummy_magic_24_0.V_source.n11 32.3838
R9311 two_stage_opamp_dummy_magic_24_0.V_source.n16 two_stage_opamp_dummy_magic_24_0.V_source.n15 32.3838
R9312 two_stage_opamp_dummy_magic_24_0.V_source.n52 two_stage_opamp_dummy_magic_24_0.V_source.n51 32.3838
R9313 two_stage_opamp_dummy_magic_24_0.V_source.n54 two_stage_opamp_dummy_magic_24_0.V_source.n53 32.3838
R9314 two_stage_opamp_dummy_magic_24_0.V_source.n56 two_stage_opamp_dummy_magic_24_0.V_source.n55 32.3838
R9315 two_stage_opamp_dummy_magic_24_0.V_source.n50 two_stage_opamp_dummy_magic_24_0.V_source.n49 32.3838
R9316 two_stage_opamp_dummy_magic_24_0.V_source.n28 two_stage_opamp_dummy_magic_24_0.V_source.t27 16.0005
R9317 two_stage_opamp_dummy_magic_24_0.V_source.n28 two_stage_opamp_dummy_magic_24_0.V_source.t30 16.0005
R9318 two_stage_opamp_dummy_magic_24_0.V_source.n26 two_stage_opamp_dummy_magic_24_0.V_source.t38 16.0005
R9319 two_stage_opamp_dummy_magic_24_0.V_source.n26 two_stage_opamp_dummy_magic_24_0.V_source.t36 16.0005
R9320 two_stage_opamp_dummy_magic_24_0.V_source.n18 two_stage_opamp_dummy_magic_24_0.V_source.t29 16.0005
R9321 two_stage_opamp_dummy_magic_24_0.V_source.n18 two_stage_opamp_dummy_magic_24_0.V_source.t21 16.0005
R9322 two_stage_opamp_dummy_magic_24_0.V_source.n34 two_stage_opamp_dummy_magic_24_0.V_source.t14 16.0005
R9323 two_stage_opamp_dummy_magic_24_0.V_source.n34 two_stage_opamp_dummy_magic_24_0.V_source.t13 16.0005
R9324 two_stage_opamp_dummy_magic_24_0.V_source.n31 two_stage_opamp_dummy_magic_24_0.V_source.t12 16.0005
R9325 two_stage_opamp_dummy_magic_24_0.V_source.n31 two_stage_opamp_dummy_magic_24_0.V_source.t7 16.0005
R9326 two_stage_opamp_dummy_magic_24_0.V_source.n43 two_stage_opamp_dummy_magic_24_0.V_source.t8 16.0005
R9327 two_stage_opamp_dummy_magic_24_0.V_source.n43 two_stage_opamp_dummy_magic_24_0.V_source.t5 16.0005
R9328 two_stage_opamp_dummy_magic_24_0.V_source.n39 two_stage_opamp_dummy_magic_24_0.V_source.t6 16.0005
R9329 two_stage_opamp_dummy_magic_24_0.V_source.n39 two_stage_opamp_dummy_magic_24_0.V_source.t10 16.0005
R9330 two_stage_opamp_dummy_magic_24_0.V_source.n37 two_stage_opamp_dummy_magic_24_0.V_source.t9 16.0005
R9331 two_stage_opamp_dummy_magic_24_0.V_source.n37 two_stage_opamp_dummy_magic_24_0.V_source.t11 16.0005
R9332 two_stage_opamp_dummy_magic_24_0.V_source.n22 two_stage_opamp_dummy_magic_24_0.V_source.t37 16.0005
R9333 two_stage_opamp_dummy_magic_24_0.V_source.n22 two_stage_opamp_dummy_magic_24_0.V_source.t26 16.0005
R9334 two_stage_opamp_dummy_magic_24_0.V_source.n20 two_stage_opamp_dummy_magic_24_0.V_source.t15 16.0005
R9335 two_stage_opamp_dummy_magic_24_0.V_source.n20 two_stage_opamp_dummy_magic_24_0.V_source.t33 16.0005
R9336 two_stage_opamp_dummy_magic_24_0.V_source.n46 two_stage_opamp_dummy_magic_24_0.V_source.t1 9.6005
R9337 two_stage_opamp_dummy_magic_24_0.V_source.n46 two_stage_opamp_dummy_magic_24_0.V_source.t17 9.6005
R9338 two_stage_opamp_dummy_magic_24_0.V_source.n48 two_stage_opamp_dummy_magic_24_0.V_source.t3 9.6005
R9339 two_stage_opamp_dummy_magic_24_0.V_source.n48 two_stage_opamp_dummy_magic_24_0.V_source.t32 9.6005
R9340 two_stage_opamp_dummy_magic_24_0.V_source.n10 two_stage_opamp_dummy_magic_24_0.V_source.t23 9.6005
R9341 two_stage_opamp_dummy_magic_24_0.V_source.n10 two_stage_opamp_dummy_magic_24_0.V_source.t4 9.6005
R9342 two_stage_opamp_dummy_magic_24_0.V_source.n13 two_stage_opamp_dummy_magic_24_0.V_source.t39 9.6005
R9343 two_stage_opamp_dummy_magic_24_0.V_source.n13 two_stage_opamp_dummy_magic_24_0.V_source.t40 9.6005
R9344 two_stage_opamp_dummy_magic_24_0.V_source.n11 two_stage_opamp_dummy_magic_24_0.V_source.t20 9.6005
R9345 two_stage_opamp_dummy_magic_24_0.V_source.n11 two_stage_opamp_dummy_magic_24_0.V_source.t19 9.6005
R9346 two_stage_opamp_dummy_magic_24_0.V_source.n15 two_stage_opamp_dummy_magic_24_0.V_source.t2 9.6005
R9347 two_stage_opamp_dummy_magic_24_0.V_source.n15 two_stage_opamp_dummy_magic_24_0.V_source.t25 9.6005
R9348 two_stage_opamp_dummy_magic_24_0.V_source.n51 two_stage_opamp_dummy_magic_24_0.V_source.t35 9.6005
R9349 two_stage_opamp_dummy_magic_24_0.V_source.n51 two_stage_opamp_dummy_magic_24_0.V_source.t18 9.6005
R9350 two_stage_opamp_dummy_magic_24_0.V_source.n53 two_stage_opamp_dummy_magic_24_0.V_source.t16 9.6005
R9351 two_stage_opamp_dummy_magic_24_0.V_source.n53 two_stage_opamp_dummy_magic_24_0.V_source.t31 9.6005
R9352 two_stage_opamp_dummy_magic_24_0.V_source.n55 two_stage_opamp_dummy_magic_24_0.V_source.t22 9.6005
R9353 two_stage_opamp_dummy_magic_24_0.V_source.n55 two_stage_opamp_dummy_magic_24_0.V_source.t24 9.6005
R9354 two_stage_opamp_dummy_magic_24_0.V_source.n49 two_stage_opamp_dummy_magic_24_0.V_source.t34 9.6005
R9355 two_stage_opamp_dummy_magic_24_0.V_source.n49 two_stage_opamp_dummy_magic_24_0.V_source.t0 9.6005
R9356 two_stage_opamp_dummy_magic_24_0.V_source.n58 two_stage_opamp_dummy_magic_24_0.V_source.n8 5.85227
R9357 two_stage_opamp_dummy_magic_24_0.V_source.n38 two_stage_opamp_dummy_magic_24_0.V_source.n4 5.51092
R9358 two_stage_opamp_dummy_magic_24_0.V_source.n3 two_stage_opamp_dummy_magic_24_0.V_source.n19 5.51092
R9359 two_stage_opamp_dummy_magic_24_0.V_source.n41 two_stage_opamp_dummy_magic_24_0.V_source.n38 5.45883
R9360 two_stage_opamp_dummy_magic_24_0.V_source.n19 two_stage_opamp_dummy_magic_24_0.V_source.n17 5.45883
R9361 two_stage_opamp_dummy_magic_24_0.V_source.n52 two_stage_opamp_dummy_magic_24_0.V_source.n5 5.188
R9362 two_stage_opamp_dummy_magic_24_0.V_source.n54 two_stage_opamp_dummy_magic_24_0.V_source.n5 5.188
R9363 two_stage_opamp_dummy_magic_24_0.V_source.n57 two_stage_opamp_dummy_magic_24_0.V_source.n56 5.188
R9364 two_stage_opamp_dummy_magic_24_0.V_source.n4 two_stage_opamp_dummy_magic_24_0.V_source.n44 5.16717
R9365 two_stage_opamp_dummy_magic_24_0.V_source.n40 two_stage_opamp_dummy_magic_24_0.V_source.n4 5.16717
R9366 two_stage_opamp_dummy_magic_24_0.V_source.n23 two_stage_opamp_dummy_magic_24_0.V_source.n3 5.16717
R9367 two_stage_opamp_dummy_magic_24_0.V_source.n3 two_stage_opamp_dummy_magic_24_0.V_source.n21 5.16717
R9368 two_stage_opamp_dummy_magic_24_0.V_source.n36 two_stage_opamp_dummy_magic_24_0.V_source.n35 4.89633
R9369 two_stage_opamp_dummy_magic_24_0.V_source.n44 two_stage_opamp_dummy_magic_24_0.V_source.n42 4.89633
R9370 two_stage_opamp_dummy_magic_24_0.V_source.n41 two_stage_opamp_dummy_magic_24_0.V_source.n40 4.89633
R9371 two_stage_opamp_dummy_magic_24_0.V_source.n30 two_stage_opamp_dummy_magic_24_0.V_source.n29 4.89633
R9372 two_stage_opamp_dummy_magic_24_0.V_source.n33 two_stage_opamp_dummy_magic_24_0.V_source.n32 4.89633
R9373 two_stage_opamp_dummy_magic_24_0.V_source.n24 two_stage_opamp_dummy_magic_24_0.V_source.n23 4.89633
R9374 two_stage_opamp_dummy_magic_24_0.V_source.n21 two_stage_opamp_dummy_magic_24_0.V_source.n17 4.89633
R9375 two_stage_opamp_dummy_magic_24_0.V_source.n27 two_stage_opamp_dummy_magic_24_0.V_source.n25 4.89633
R9376 two_stage_opamp_dummy_magic_24_0.V_source.n33 two_stage_opamp_dummy_magic_24_0.V_source.n30 3.6255
R9377 two_stage_opamp_dummy_magic_24_0.V_source.n1 two_stage_opamp_dummy_magic_24_0.V_source.n9 2.55956
R9378 two_stage_opamp_dummy_magic_24_0.V_source.n47 two_stage_opamp_dummy_magic_24_0.V_source.n1 2.44497
R9379 two_stage_opamp_dummy_magic_24_0.V_source.n0 two_stage_opamp_dummy_magic_24_0.V_source.n14 2.44497
R9380 two_stage_opamp_dummy_magic_24_0.V_source.n0 two_stage_opamp_dummy_magic_24_0.V_source.n12 2.44497
R9381 two_stage_opamp_dummy_magic_24_0.V_source.n1 two_stage_opamp_dummy_magic_24_0.V_source.n16 2.44497
R9382 two_stage_opamp_dummy_magic_24_0.V_source.n1 two_stage_opamp_dummy_magic_24_0.V_source.n52 2.44497
R9383 two_stage_opamp_dummy_magic_24_0.V_source.n1 two_stage_opamp_dummy_magic_24_0.V_source.n54 2.44497
R9384 two_stage_opamp_dummy_magic_24_0.V_source.n56 two_stage_opamp_dummy_magic_24_0.V_source.n1 2.44497
R9385 two_stage_opamp_dummy_magic_24_0.V_source.n0 two_stage_opamp_dummy_magic_24_0.V_source.n8 2.44497
R9386 two_stage_opamp_dummy_magic_24_0.V_source.n50 two_stage_opamp_dummy_magic_24_0.V_source.n1 2.44462
R9387 two_stage_opamp_dummy_magic_24_0.V_source.n45 two_stage_opamp_dummy_magic_24_0.V_source.n2 2.2076
R9388 two_stage_opamp_dummy_magic_24_0.V_source.n7 two_stage_opamp_dummy_magic_24_0.V_source.n45 2.16822
R9389 two_stage_opamp_dummy_magic_24_0.V_source.n2 two_stage_opamp_dummy_magic_24_0.V_source.n6 2.16822
R9390 two_stage_opamp_dummy_magic_24_0.V_source.n5 two_stage_opamp_dummy_magic_24_0.V_source.n7 2.02255
R9391 two_stage_opamp_dummy_magic_24_0.V_source.n6 two_stage_opamp_dummy_magic_24_0.V_source.n58 1.36007
R9392 two_stage_opamp_dummy_magic_24_0.V_source.n58 two_stage_opamp_dummy_magic_24_0.V_source.n57 0.664374
R9393 two_stage_opamp_dummy_magic_24_0.V_source.n7 two_stage_opamp_dummy_magic_24_0.V_source.n47 0.6255
R9394 two_stage_opamp_dummy_magic_24_0.V_source.n7 two_stage_opamp_dummy_magic_24_0.V_source.n9 0.6255
R9395 two_stage_opamp_dummy_magic_24_0.V_source.n16 two_stage_opamp_dummy_magic_24_0.V_source.n6 0.6255
R9396 two_stage_opamp_dummy_magic_24_0.V_source.n12 two_stage_opamp_dummy_magic_24_0.V_source.n6 0.6255
R9397 two_stage_opamp_dummy_magic_24_0.V_source.n14 two_stage_opamp_dummy_magic_24_0.V_source.n6 0.6255
R9398 two_stage_opamp_dummy_magic_24_0.V_source.n7 two_stage_opamp_dummy_magic_24_0.V_source.n50 0.6255
R9399 two_stage_opamp_dummy_magic_24_0.V_source.n32 two_stage_opamp_dummy_magic_24_0.V_source.n7 0.604667
R9400 two_stage_opamp_dummy_magic_24_0.V_source.n6 two_stage_opamp_dummy_magic_24_0.V_source.n27 0.604667
R9401 two_stage_opamp_dummy_magic_24_0.V_source.n42 two_stage_opamp_dummy_magic_24_0.V_source.n41 0.563
R9402 two_stage_opamp_dummy_magic_24_0.V_source.n42 two_stage_opamp_dummy_magic_24_0.V_source.n36 0.563
R9403 two_stage_opamp_dummy_magic_24_0.V_source.n36 two_stage_opamp_dummy_magic_24_0.V_source.n33 0.563
R9404 two_stage_opamp_dummy_magic_24_0.V_source.n30 two_stage_opamp_dummy_magic_24_0.V_source.n25 0.563
R9405 two_stage_opamp_dummy_magic_24_0.V_source.n24 two_stage_opamp_dummy_magic_24_0.V_source.n17 0.563
R9406 two_stage_opamp_dummy_magic_24_0.V_source.n25 two_stage_opamp_dummy_magic_24_0.V_source.n24 0.563
R9407 two_stage_opamp_dummy_magic_24_0.V_source.n0 two_stage_opamp_dummy_magic_24_0.V_source.t28 84.5617
R9408 two_stage_opamp_dummy_magic_24_0.V_source.n1 two_stage_opamp_dummy_magic_24_0.V_source.n0 0.917167
R9409 two_stage_opamp_dummy_magic_24_0.V_source.n35 two_stage_opamp_dummy_magic_24_0.V_source.n7 0.854667
R9410 two_stage_opamp_dummy_magic_24_0.V_source.n29 two_stage_opamp_dummy_magic_24_0.V_source.n6 0.854667
R9411 two_stage_opamp_dummy_magic_24_0.V_source.n45 two_stage_opamp_dummy_magic_24_0.V_source.n4 0.854052
R9412 two_stage_opamp_dummy_magic_24_0.V_source.n3 two_stage_opamp_dummy_magic_24_0.V_source.n2 0.854052
R9413 two_stage_opamp_dummy_magic_24_0.V_source.n57 two_stage_opamp_dummy_magic_24_0.V_source.n5 0.688
R9414 two_stage_opamp_dummy_magic_24_0.VD2.n25 two_stage_opamp_dummy_magic_24_0.VD2.n24 49.7255
R9415 two_stage_opamp_dummy_magic_24_0.VD2.n1 two_stage_opamp_dummy_magic_24_0.VD2.n0 49.7255
R9416 two_stage_opamp_dummy_magic_24_0.VD2.n21 two_stage_opamp_dummy_magic_24_0.VD2.n12 49.7255
R9417 two_stage_opamp_dummy_magic_24_0.VD2.n11 two_stage_opamp_dummy_magic_24_0.VD2.n10 49.7255
R9418 two_stage_opamp_dummy_magic_24_0.VD2.n27 two_stage_opamp_dummy_magic_24_0.VD2.n9 49.7255
R9419 two_stage_opamp_dummy_magic_24_0.VD2.n15 two_stage_opamp_dummy_magic_24_0.VD2.n14 49.3505
R9420 two_stage_opamp_dummy_magic_24_0.VD2.n18 two_stage_opamp_dummy_magic_24_0.VD2.n17 49.3505
R9421 two_stage_opamp_dummy_magic_24_0.VD2.n5 two_stage_opamp_dummy_magic_24_0.VD2.n4 49.3505
R9422 two_stage_opamp_dummy_magic_24_0.VD2.n35 two_stage_opamp_dummy_magic_24_0.VD2.n34 49.3505
R9423 two_stage_opamp_dummy_magic_24_0.VD2.n8 two_stage_opamp_dummy_magic_24_0.VD2.n7 49.3505
R9424 two_stage_opamp_dummy_magic_24_0.VD2.n31 two_stage_opamp_dummy_magic_24_0.VD2.n30 49.3505
R9425 two_stage_opamp_dummy_magic_24_0.VD2.n14 two_stage_opamp_dummy_magic_24_0.VD2.t19 16.0005
R9426 two_stage_opamp_dummy_magic_24_0.VD2.n14 two_stage_opamp_dummy_magic_24_0.VD2.t3 16.0005
R9427 two_stage_opamp_dummy_magic_24_0.VD2.n17 two_stage_opamp_dummy_magic_24_0.VD2.t8 16.0005
R9428 two_stage_opamp_dummy_magic_24_0.VD2.n17 two_stage_opamp_dummy_magic_24_0.VD2.t1 16.0005
R9429 two_stage_opamp_dummy_magic_24_0.VD2.n4 two_stage_opamp_dummy_magic_24_0.VD2.t4 16.0005
R9430 two_stage_opamp_dummy_magic_24_0.VD2.n4 two_stage_opamp_dummy_magic_24_0.VD2.t2 16.0005
R9431 two_stage_opamp_dummy_magic_24_0.VD2.n34 two_stage_opamp_dummy_magic_24_0.VD2.t7 16.0005
R9432 two_stage_opamp_dummy_magic_24_0.VD2.n34 two_stage_opamp_dummy_magic_24_0.VD2.t0 16.0005
R9433 two_stage_opamp_dummy_magic_24_0.VD2.n24 two_stage_opamp_dummy_magic_24_0.VD2.t10 16.0005
R9434 two_stage_opamp_dummy_magic_24_0.VD2.n24 two_stage_opamp_dummy_magic_24_0.VD2.t11 16.0005
R9435 two_stage_opamp_dummy_magic_24_0.VD2.n0 two_stage_opamp_dummy_magic_24_0.VD2.t21 16.0005
R9436 two_stage_opamp_dummy_magic_24_0.VD2.n0 two_stage_opamp_dummy_magic_24_0.VD2.t20 16.0005
R9437 two_stage_opamp_dummy_magic_24_0.VD2.n12 two_stage_opamp_dummy_magic_24_0.VD2.t15 16.0005
R9438 two_stage_opamp_dummy_magic_24_0.VD2.n12 two_stage_opamp_dummy_magic_24_0.VD2.t17 16.0005
R9439 two_stage_opamp_dummy_magic_24_0.VD2.n10 two_stage_opamp_dummy_magic_24_0.VD2.t18 16.0005
R9440 two_stage_opamp_dummy_magic_24_0.VD2.n10 two_stage_opamp_dummy_magic_24_0.VD2.t16 16.0005
R9441 two_stage_opamp_dummy_magic_24_0.VD2.n9 two_stage_opamp_dummy_magic_24_0.VD2.t13 16.0005
R9442 two_stage_opamp_dummy_magic_24_0.VD2.n9 two_stage_opamp_dummy_magic_24_0.VD2.t14 16.0005
R9443 two_stage_opamp_dummy_magic_24_0.VD2.n7 two_stage_opamp_dummy_magic_24_0.VD2.t5 16.0005
R9444 two_stage_opamp_dummy_magic_24_0.VD2.n7 two_stage_opamp_dummy_magic_24_0.VD2.t12 16.0005
R9445 two_stage_opamp_dummy_magic_24_0.VD2.n30 two_stage_opamp_dummy_magic_24_0.VD2.t6 16.0005
R9446 two_stage_opamp_dummy_magic_24_0.VD2.n30 two_stage_opamp_dummy_magic_24_0.VD2.t9 16.0005
R9447 two_stage_opamp_dummy_magic_24_0.VD2.n25 two_stage_opamp_dummy_magic_24_0.VD2.n3 6.29217
R9448 two_stage_opamp_dummy_magic_24_0.VD2.n21 two_stage_opamp_dummy_magic_24_0.VD2.n20 6.29217
R9449 two_stage_opamp_dummy_magic_24_0.VD2.n13 two_stage_opamp_dummy_magic_24_0.VD2.n11 6.29217
R9450 two_stage_opamp_dummy_magic_24_0.VD2.n28 two_stage_opamp_dummy_magic_24_0.VD2.n27 6.29217
R9451 two_stage_opamp_dummy_magic_24_0.VD2.n32 two_stage_opamp_dummy_magic_24_0.VD2.n8 5.438
R9452 two_stage_opamp_dummy_magic_24_0.VD2.n16 two_stage_opamp_dummy_magic_24_0.VD2.n15 5.438
R9453 two_stage_opamp_dummy_magic_24_0.VD2.n28 two_stage_opamp_dummy_magic_24_0.VD2.n8 5.31821
R9454 two_stage_opamp_dummy_magic_24_0.VD2.n15 two_stage_opamp_dummy_magic_24_0.VD2.n13 5.31821
R9455 two_stage_opamp_dummy_magic_24_0.VD2.n19 two_stage_opamp_dummy_magic_24_0.VD2.n18 5.08383
R9456 two_stage_opamp_dummy_magic_24_0.VD2.n5 two_stage_opamp_dummy_magic_24_0.VD2.n2 5.08383
R9457 two_stage_opamp_dummy_magic_24_0.VD2.n36 two_stage_opamp_dummy_magic_24_0.VD2.n35 5.08383
R9458 two_stage_opamp_dummy_magic_24_0.VD2.n31 two_stage_opamp_dummy_magic_24_0.VD2.n29 5.08383
R9459 two_stage_opamp_dummy_magic_24_0.VD2.n22 two_stage_opamp_dummy_magic_24_0.VD2.n11 5.063
R9460 two_stage_opamp_dummy_magic_24_0.VD2.n27 two_stage_opamp_dummy_magic_24_0.VD2.n26 5.063
R9461 two_stage_opamp_dummy_magic_24_0.VD2.n18 two_stage_opamp_dummy_magic_24_0.VD2.n16 4.8755
R9462 two_stage_opamp_dummy_magic_24_0.VD2.n6 two_stage_opamp_dummy_magic_24_0.VD2.n5 4.8755
R9463 two_stage_opamp_dummy_magic_24_0.VD2.n35 two_stage_opamp_dummy_magic_24_0.VD2.n33 4.8755
R9464 two_stage_opamp_dummy_magic_24_0.VD2.n32 two_stage_opamp_dummy_magic_24_0.VD2.n31 4.8755
R9465 two_stage_opamp_dummy_magic_24_0.VD2 two_stage_opamp_dummy_magic_24_0.VD2.n37 4.60467
R9466 two_stage_opamp_dummy_magic_24_0.VD2.n22 two_stage_opamp_dummy_magic_24_0.VD2.n21 4.5005
R9467 two_stage_opamp_dummy_magic_24_0.VD2.n23 two_stage_opamp_dummy_magic_24_0.VD2.n1 4.5005
R9468 two_stage_opamp_dummy_magic_24_0.VD2.n26 two_stage_opamp_dummy_magic_24_0.VD2.n25 4.5005
R9469 two_stage_opamp_dummy_magic_24_0.VD2 two_stage_opamp_dummy_magic_24_0.VD2.n1 1.688
R9470 two_stage_opamp_dummy_magic_24_0.VD2.n23 two_stage_opamp_dummy_magic_24_0.VD2.n22 0.563
R9471 two_stage_opamp_dummy_magic_24_0.VD2.n26 two_stage_opamp_dummy_magic_24_0.VD2.n23 0.563
R9472 two_stage_opamp_dummy_magic_24_0.VD2.n16 two_stage_opamp_dummy_magic_24_0.VD2.n6 0.563
R9473 two_stage_opamp_dummy_magic_24_0.VD2.n33 two_stage_opamp_dummy_magic_24_0.VD2.n6 0.563
R9474 two_stage_opamp_dummy_magic_24_0.VD2.n33 two_stage_opamp_dummy_magic_24_0.VD2.n32 0.563
R9475 two_stage_opamp_dummy_magic_24_0.VD2.n29 two_stage_opamp_dummy_magic_24_0.VD2.n28 0.234875
R9476 two_stage_opamp_dummy_magic_24_0.VD2.n29 two_stage_opamp_dummy_magic_24_0.VD2.n3 0.234875
R9477 two_stage_opamp_dummy_magic_24_0.VD2.n36 two_stage_opamp_dummy_magic_24_0.VD2.n3 0.234875
R9478 two_stage_opamp_dummy_magic_24_0.VD2.n37 two_stage_opamp_dummy_magic_24_0.VD2.n36 0.234875
R9479 two_stage_opamp_dummy_magic_24_0.VD2.n37 two_stage_opamp_dummy_magic_24_0.VD2.n2 0.234875
R9480 two_stage_opamp_dummy_magic_24_0.VD2.n20 two_stage_opamp_dummy_magic_24_0.VD2.n2 0.234875
R9481 two_stage_opamp_dummy_magic_24_0.VD2.n20 two_stage_opamp_dummy_magic_24_0.VD2.n19 0.234875
R9482 two_stage_opamp_dummy_magic_24_0.VD2.n19 two_stage_opamp_dummy_magic_24_0.VD2.n13 0.234875
R9483 GNDA.n3318 GNDA.n3317 396244
R9484 GNDA.n1466 GNDA.n1464 287100
R9485 GNDA.n3324 GNDA.n3323 284429
R9486 GNDA.n4623 GNDA.n4622 280024
R9487 GNDA.n4627 GNDA.n428 212953
R9488 GNDA.n3321 GNDA.n3320 192657
R9489 GNDA.n3321 GNDA.n1464 175770
R9490 GNDA.n3320 GNDA.n3319 171600
R9491 GNDA.n4622 GNDA.n4621 147745
R9492 GNDA.n4622 GNDA.t173 138700
R9493 GNDA.n1466 GNDA.n742 135705
R9494 GNDA.n3323 GNDA.n3322 124143
R9495 GNDA.n3317 GNDA.n3316 105027
R9496 GNDA.n3324 GNDA.n746 77980.7
R9497 GNDA.n3317 GNDA.n3304 71214.8
R9498 GNDA.n3318 GNDA.t309 55812.1
R9499 GNDA.n3306 GNDA.n3305 44241
R9500 GNDA.n3313 GNDA.n3312 37118.9
R9501 GNDA.n3609 GNDA.n571 36266
R9502 GNDA.n3311 GNDA.n3310 34786.4
R9503 GNDA.n431 GNDA.n430 30642.9
R9504 GNDA.n3316 GNDA.n1467 23059.8
R9505 GNDA.n3312 GNDA.n1467 22000
R9506 GNDA.n430 GNDA.n429 20900
R9507 GNDA.n3312 GNDA.n3311 20388.3
R9508 GNDA.n3318 GNDA.n1465 19727.9
R9509 GNDA.n4622 GNDA.t289 19113.8
R9510 GNDA.n4623 GNDA.n431 17600
R9511 GNDA.n3322 GNDA.n3321 17285.7
R9512 GNDA.n4625 GNDA.n4624 17160
R9513 GNDA.n4641 GNDA.n4640 17109.1
R9514 GNDA.n4626 GNDA.n4625 16010.8
R9515 GNDA.n3314 GNDA.n3313 13613.1
R9516 GNDA.n3310 GNDA.n3307 13528.5
R9517 GNDA.n3315 GNDA.n3314 13460.8
R9518 GNDA.n4621 GNDA.n431 12238.2
R9519 GNDA.n4621 GNDA.n4620 11720.7
R9520 GNDA.n3303 GNDA.n428 11693.7
R9521 GNDA.n3309 GNDA.n1463 11440
R9522 GNDA.n3325 GNDA.n1463 9920.29
R9523 GNDA.n3311 GNDA.n3306 9541.89
R9524 GNDA.n3304 GNDA.n3303 9511.11
R9525 GNDA.n3313 GNDA.n428 8875.99
R9526 GNDA.n3213 GNDA.n3212 7286.54
R9527 GNDA.n3314 GNDA.n1467 7240.76
R9528 GNDA.n3307 GNDA.n1467 6386.29
R9529 GNDA.n4622 GNDA.t41 6264.76
R9530 GNDA.n3305 GNDA.n1463 6187.5
R9531 GNDA.n3308 GNDA.n3307 5929.09
R9532 GNDA.n3323 GNDA.n1464 5689.59
R9533 GNDA.n571 GNDA.n429 5235.44
R9534 GNDA.n3308 GNDA.n1465 4407.11
R9535 GNDA.n3315 GNDA.n3304 4106.67
R9536 GNDA.n3303 GNDA.t62 4106.67
R9537 GNDA.n3320 GNDA.n1465 3818.87
R9538 GNDA.n3318 GNDA.n1467 3606.56
R9539 GNDA.n3310 GNDA.n3309 3390.16
R9540 GNDA.t33 GNDA.n571 2556.19
R9541 GNDA.n3322 GNDA.n1462 1911.48
R9542 GNDA.n4625 GNDA.n429 1885.71
R9543 GNDA.n3325 GNDA.n1462 1821.31
R9544 GNDA.n3223 GNDA.n3222 1684.55
R9545 GNDA.n3320 GNDA.n1462 1618.87
R9546 GNDA.n3309 GNDA.n3308 1522.77
R9547 GNDA.n3305 GNDA.n571 1215.24
R9548 GNDA.n3316 GNDA.n3315 1031.25
R9549 GNDA.n740 GNDA.t123 749.742
R9550 GNDA.n4618 GNDA.t152 747.734
R9551 GNDA.n4615 GNDA.t67 747.734
R9552 GNDA.n744 GNDA.t139 747.734
R9553 GNDA.t62 GNDA.n102 741.376
R9554 GNDA.n3247 GNDA.n3246 686.717
R9555 GNDA.n2826 GNDA.n2825 686.717
R9556 GNDA.n2818 GNDA.n2692 686.717
R9557 GNDA.n3243 GNDA.n1521 686.717
R9558 GNDA.n1738 GNDA.t13 671.187
R9559 GNDA.n2804 GNDA.n2803 669.307
R9560 GNDA.n2707 GNDA.n2706 669.307
R9561 GNDA.n568 GNDA.t119 659.367
R9562 GNDA.n3365 GNDA.t82 659.367
R9563 GNDA.n3586 GNDA.t150 659.367
R9564 GNDA.n3569 GNDA.t85 659.367
R9565 GNDA.n4682 GNDA.n357 654.447
R9566 GNDA.n2657 GNDA.n2656 585.003
R9567 GNDA.n2931 GNDA.n2930 585.001
R9568 GNDA.n2919 GNDA.n2918 585.001
R9569 GNDA.n2736 GNDA.n2735 585.001
R9570 GNDA.n3277 GNDA.n3276 585.001
R9571 GNDA.n2801 GNDA.n2800 585.001
R9572 GNDA.n1829 GNDA.n1828 585.001
R9573 GNDA.n3265 GNDA.n3264 585.001
R9574 GNDA.n4697 GNDA.n4696 585
R9575 GNDA.n4698 GNDA.n4697 585
R9576 GNDA.n299 GNDA.n298 585
R9577 GNDA.n4699 GNDA.n299 585
R9578 GNDA.n4702 GNDA.n4701 585
R9579 GNDA.n4701 GNDA.n4700 585
R9580 GNDA.n4703 GNDA.n297 585
R9581 GNDA.n297 GNDA.n296 585
R9582 GNDA.n4705 GNDA.n4704 585
R9583 GNDA.n4706 GNDA.n4705 585
R9584 GNDA.n295 GNDA.n294 585
R9585 GNDA.n4707 GNDA.n295 585
R9586 GNDA.n4710 GNDA.n4709 585
R9587 GNDA.n4709 GNDA.n4708 585
R9588 GNDA.n4711 GNDA.n293 585
R9589 GNDA.n293 GNDA.n292 585
R9590 GNDA.n4713 GNDA.n4712 585
R9591 GNDA.n4714 GNDA.n4713 585
R9592 GNDA.n291 GNDA.n290 585
R9593 GNDA.n4715 GNDA.n291 585
R9594 GNDA.n4718 GNDA.n4717 585
R9595 GNDA.n4717 GNDA.n4716 585
R9596 GNDA.n4719 GNDA.n289 585
R9597 GNDA.n289 GNDA.n99 585
R9598 GNDA.n4681 GNDA.n4680 585
R9599 GNDA.n4679 GNDA.n355 585
R9600 GNDA.t62 GNDA.n355 585
R9601 GNDA.n5078 GNDA.n5077 585
R9602 GNDA.n131 GNDA.n129 585
R9603 GNDA.n242 GNDA.n241 585
R9604 GNDA.n244 GNDA.n243 585
R9605 GNDA.n246 GNDA.n245 585
R9606 GNDA.n248 GNDA.n247 585
R9607 GNDA.n250 GNDA.n249 585
R9608 GNDA.n252 GNDA.n251 585
R9609 GNDA.n254 GNDA.n253 585
R9610 GNDA.n256 GNDA.n255 585
R9611 GNDA.n258 GNDA.n257 585
R9612 GNDA.n260 GNDA.n259 585
R9613 GNDA.n1587 GNDA.n1586 585
R9614 GNDA.n1584 GNDA.n1583 585
R9615 GNDA.n1582 GNDA.n1581 585
R9616 GNDA.n1580 GNDA.n1579 585
R9617 GNDA.n1578 GNDA.n1577 585
R9618 GNDA.n1576 GNDA.n1575 585
R9619 GNDA.n1574 GNDA.n1573 585
R9620 GNDA.n1572 GNDA.n1571 585
R9621 GNDA.n1570 GNDA.n1569 585
R9622 GNDA.n1568 GNDA.n1567 585
R9623 GNDA.n1566 GNDA.n1565 585
R9624 GNDA.n135 GNDA.n132 585
R9625 GNDA.n1741 GNDA.n1740 585
R9626 GNDA.n1743 GNDA.n1742 585
R9627 GNDA.n1745 GNDA.n1744 585
R9628 GNDA.n1747 GNDA.n1746 585
R9629 GNDA.n1749 GNDA.n1748 585
R9630 GNDA.n1751 GNDA.n1750 585
R9631 GNDA.n1753 GNDA.n1752 585
R9632 GNDA.n1755 GNDA.n1754 585
R9633 GNDA.n1757 GNDA.n1756 585
R9634 GNDA.n1759 GNDA.n1758 585
R9635 GNDA.n1761 GNDA.n1760 585
R9636 GNDA.n1763 GNDA.n1762 585
R9637 GNDA.n5258 GNDA.n5257 585
R9638 GNDA.n5255 GNDA.n54 585
R9639 GNDA.n59 GNDA.n58 585
R9640 GNDA.n5250 GNDA.n5249 585
R9641 GNDA.n5248 GNDA.n5247 585
R9642 GNDA.n5174 GNDA.n63 585
R9643 GNDA.n5176 GNDA.n5175 585
R9644 GNDA.n5181 GNDA.n5180 585
R9645 GNDA.n5179 GNDA.n5172 585
R9646 GNDA.n5187 GNDA.n5186 585
R9647 GNDA.n5189 GNDA.n5188 585
R9648 GNDA.n5170 GNDA.n5169 585
R9649 GNDA.n4835 GNDA.n4834 585
R9650 GNDA.n4832 GNDA.n4831 585
R9651 GNDA.n4830 GNDA.n4829 585
R9652 GNDA.n4746 GNDA.n4722 585
R9653 GNDA.n4748 GNDA.n4747 585
R9654 GNDA.n4752 GNDA.n4751 585
R9655 GNDA.n4754 GNDA.n4753 585
R9656 GNDA.n4761 GNDA.n4760 585
R9657 GNDA.n4759 GNDA.n4744 585
R9658 GNDA.n4767 GNDA.n4766 585
R9659 GNDA.n4769 GNDA.n4768 585
R9660 GNDA.n4742 GNDA.n4741 585
R9661 GNDA.n328 GNDA.n325 585
R9662 GNDA.n329 GNDA.n323 585
R9663 GNDA.n330 GNDA.n322 585
R9664 GNDA.n320 GNDA.n318 585
R9665 GNDA.n336 GNDA.n317 585
R9666 GNDA.n337 GNDA.n315 585
R9667 GNDA.n338 GNDA.n314 585
R9668 GNDA.n312 GNDA.n310 585
R9669 GNDA.n344 GNDA.n309 585
R9670 GNDA.n345 GNDA.n307 585
R9671 GNDA.n346 GNDA.n306 585
R9672 GNDA.n302 GNDA.n301 585
R9673 GNDA.n133 GNDA.n85 585
R9674 GNDA.n5167 GNDA.n85 585
R9675 GNDA.n349 GNDA.n302 585
R9676 GNDA.n347 GNDA.n346 585
R9677 GNDA.n345 GNDA.n304 585
R9678 GNDA.n344 GNDA.n343 585
R9679 GNDA.n341 GNDA.n310 585
R9680 GNDA.n339 GNDA.n338 585
R9681 GNDA.n337 GNDA.n311 585
R9682 GNDA.n336 GNDA.n335 585
R9683 GNDA.n333 GNDA.n318 585
R9684 GNDA.n331 GNDA.n330 585
R9685 GNDA.n329 GNDA.n319 585
R9686 GNDA.n328 GNDA.n327 585
R9687 GNDA.n133 GNDA.n55 585
R9688 GNDA.n5167 GNDA.n55 585
R9689 GNDA.n5053 GNDA.n159 585
R9690 GNDA.n5054 GNDA.n150 585
R9691 GNDA.n5057 GNDA.n149 585
R9692 GNDA.n5058 GNDA.n148 585
R9693 GNDA.n5061 GNDA.n147 585
R9694 GNDA.n5062 GNDA.n146 585
R9695 GNDA.n5065 GNDA.n145 585
R9696 GNDA.n5067 GNDA.n144 585
R9697 GNDA.n5068 GNDA.n143 585
R9698 GNDA.n5069 GNDA.n142 585
R9699 GNDA.n151 GNDA.n134 585
R9700 GNDA.n5075 GNDA.n130 585
R9701 GNDA.n5075 GNDA.n5074 585
R9702 GNDA.n136 GNDA.n134 585
R9703 GNDA.n5070 GNDA.n5069 585
R9704 GNDA.n5068 GNDA.n141 585
R9705 GNDA.n5067 GNDA.n5066 585
R9706 GNDA.n5065 GNDA.n5064 585
R9707 GNDA.n5063 GNDA.n5062 585
R9708 GNDA.n5061 GNDA.n5060 585
R9709 GNDA.n5059 GNDA.n5058 585
R9710 GNDA.n5057 GNDA.n5056 585
R9711 GNDA.n5055 GNDA.n5054 585
R9712 GNDA.n5053 GNDA.n5052 585
R9713 GNDA.n3043 GNDA.n1833 585
R9714 GNDA.n3041 GNDA.n3040 585
R9715 GNDA.n1835 GNDA.n1834 585
R9716 GNDA.n1841 GNDA.n1837 585
R9717 GNDA.n3033 GNDA.n3032 585
R9718 GNDA.n3030 GNDA.n1839 585
R9719 GNDA.n3029 GNDA.n1842 585
R9720 GNDA.n3027 GNDA.n3026 585
R9721 GNDA.n1844 GNDA.n1843 585
R9722 GNDA.n3021 GNDA.n3020 585
R9723 GNDA.n3018 GNDA.n1848 585
R9724 GNDA.n3016 GNDA.n3015 585
R9725 GNDA.n3015 GNDA.n3014 585
R9726 GNDA.n1848 GNDA.n1847 585
R9727 GNDA.n3022 GNDA.n3021 585
R9728 GNDA.n3022 GNDA.n1468 585
R9729 GNDA.n3023 GNDA.n1844 585
R9730 GNDA.n3026 GNDA.n3025 585
R9731 GNDA.n1846 GNDA.n1842 585
R9732 GNDA.n1839 GNDA.n1838 585
R9733 GNDA.n3034 GNDA.n3033 585
R9734 GNDA.n3036 GNDA.n1837 585
R9735 GNDA.n3037 GNDA.n1835 585
R9736 GNDA.n3040 GNDA.n3039 585
R9737 GNDA.n1836 GNDA.n1833 585
R9738 GNDA.n1836 GNDA.n1468 585
R9739 GNDA.n2981 GNDA.n1849 585
R9740 GNDA.n2980 GNDA.n2979 585
R9741 GNDA.n2977 GNDA.n1850 585
R9742 GNDA.n2975 GNDA.n2974 585
R9743 GNDA.n2973 GNDA.n1851 585
R9744 GNDA.n2972 GNDA.n2971 585
R9745 GNDA.n2969 GNDA.n1852 585
R9746 GNDA.n2967 GNDA.n2966 585
R9747 GNDA.n2965 GNDA.n1853 585
R9748 GNDA.n2964 GNDA.n2963 585
R9749 GNDA.n2961 GNDA.n1854 585
R9750 GNDA.n2959 GNDA.n2958 585
R9751 GNDA.n2993 GNDA.n2992 585
R9752 GNDA.n2994 GNDA.n2990 585
R9753 GNDA.n2996 GNDA.n2995 585
R9754 GNDA.n2998 GNDA.n2988 585
R9755 GNDA.n3000 GNDA.n2999 585
R9756 GNDA.n3001 GNDA.n2987 585
R9757 GNDA.n3003 GNDA.n3002 585
R9758 GNDA.n3005 GNDA.n2985 585
R9759 GNDA.n3007 GNDA.n3006 585
R9760 GNDA.n3008 GNDA.n2984 585
R9761 GNDA.n3010 GNDA.n3009 585
R9762 GNDA.n3012 GNDA.n2983 585
R9763 GNDA.n3193 GNDA.n1543 585
R9764 GNDA.n3191 GNDA.n3190 585
R9765 GNDA.n3189 GNDA.n1544 585
R9766 GNDA.n3188 GNDA.n3187 585
R9767 GNDA.n3185 GNDA.n1545 585
R9768 GNDA.n3183 GNDA.n3182 585
R9769 GNDA.n3181 GNDA.n1546 585
R9770 GNDA.n3180 GNDA.n3179 585
R9771 GNDA.n3177 GNDA.n1547 585
R9772 GNDA.n3175 GNDA.n3174 585
R9773 GNDA.n3173 GNDA.n1548 585
R9774 GNDA.n3172 GNDA.n3171 585
R9775 GNDA.n4889 GNDA.n162 585
R9776 GNDA.n4889 GNDA.n161 585
R9777 GNDA.n4979 GNDA.n4978 585
R9778 GNDA.n4976 GNDA.n226 585
R9779 GNDA.n4866 GNDA.n4865 585
R9780 GNDA.n4971 GNDA.n4970 585
R9781 GNDA.n4969 GNDA.n4968 585
R9782 GNDA.n4895 GNDA.n4870 585
R9783 GNDA.n4897 GNDA.n4896 585
R9784 GNDA.n4902 GNDA.n4901 585
R9785 GNDA.n4900 GNDA.n4893 585
R9786 GNDA.n4908 GNDA.n4907 585
R9787 GNDA.n4910 GNDA.n4909 585
R9788 GNDA.n4891 GNDA.n4890 585
R9789 GNDA.n5051 GNDA.n162 585
R9790 GNDA.n5051 GNDA.n161 585
R9791 GNDA.n5050 GNDA.n5049 585
R9792 GNDA.n5047 GNDA.n5046 585
R9793 GNDA.n5045 GNDA.n5044 585
R9794 GNDA.n199 GNDA.n167 585
R9795 GNDA.n219 GNDA.n218 585
R9796 GNDA.n215 GNDA.n198 585
R9797 GNDA.n202 GNDA.n201 585
R9798 GNDA.n210 GNDA.n209 585
R9799 GNDA.n208 GNDA.n207 585
R9800 GNDA.n188 GNDA.n187 585
R9801 GNDA.n4984 GNDA.n4983 585
R9802 GNDA.n1549 GNDA.n189 585
R9803 GNDA.n1676 GNDA.n1552 585
R9804 GNDA.n1700 GNDA.n1678 585
R9805 GNDA.n1702 GNDA.n1701 585
R9806 GNDA.n1698 GNDA.n1697 585
R9807 GNDA.n1696 GNDA.n1695 585
R9808 GNDA.n1691 GNDA.n1690 585
R9809 GNDA.n1689 GNDA.n1688 585
R9810 GNDA.n1684 GNDA.n1683 585
R9811 GNDA.n1682 GNDA.n1603 585
R9812 GNDA.n1710 GNDA.n1709 585
R9813 GNDA.n1712 GNDA.n1711 585
R9814 GNDA.n1715 GNDA.n1714 585
R9815 GNDA.n1529 GNDA.n1528 585
R9816 GNDA.n3212 GNDA.n1529 585
R9817 GNDA.n3225 GNDA.n3224 585
R9818 GNDA.n3224 GNDA.n3223 585
R9819 GNDA.n3214 GNDA.n1535 585
R9820 GNDA.n3217 GNDA.n3216 585
R9821 GNDA.n3216 GNDA.n3215 585
R9822 GNDA.n1534 GNDA.n1533 585
R9823 GNDA.n3211 GNDA.n1534 585
R9824 GNDA.n3209 GNDA.n3208 585
R9825 GNDA.n3210 GNDA.n3209 585
R9826 GNDA.n3207 GNDA.n1537 585
R9827 GNDA.n1537 GNDA.n1536 585
R9828 GNDA.n3206 GNDA.n3205 585
R9829 GNDA.n3205 GNDA.n1518 585
R9830 GNDA.n3204 GNDA.n1538 585
R9831 GNDA.n3204 GNDA.n1517 585
R9832 GNDA.n3203 GNDA.n1540 585
R9833 GNDA.n3203 GNDA.n3202 585
R9834 GNDA.n3197 GNDA.n1539 585
R9835 GNDA.n3201 GNDA.n1539 585
R9836 GNDA.n3199 GNDA.n3198 585
R9837 GNDA.n3200 GNDA.n3199 585
R9838 GNDA.n3196 GNDA.n1542 585
R9839 GNDA.n1542 GNDA.n1541 585
R9840 GNDA.n3195 GNDA.n3194 585
R9841 GNDA.n3194 GNDA.n102 585
R9842 GNDA.n3213 GNDA.n1530 585
R9843 GNDA.n1600 GNDA.n1599 585
R9844 GNDA.n1720 GNDA.n1719 585
R9845 GNDA.n1721 GNDA.n1720 585
R9846 GNDA.n1597 GNDA.n1596 585
R9847 GNDA.n1722 GNDA.n1597 585
R9848 GNDA.n1725 GNDA.n1724 585
R9849 GNDA.n1724 GNDA.n1723 585
R9850 GNDA.n1726 GNDA.n1595 585
R9851 GNDA.n1598 GNDA.n1595 585
R9852 GNDA.n1728 GNDA.n1727 585
R9853 GNDA.n1728 GNDA.n108 585
R9854 GNDA.n1729 GNDA.n1594 585
R9855 GNDA.n1729 GNDA.n109 585
R9856 GNDA.n1732 GNDA.n1731 585
R9857 GNDA.n1731 GNDA.n1730 585
R9858 GNDA.n1733 GNDA.n1592 585
R9859 GNDA.n1592 GNDA.n1591 585
R9860 GNDA.n1735 GNDA.n1734 585
R9861 GNDA.n1736 GNDA.n1735 585
R9862 GNDA.n1593 GNDA.n1590 585
R9863 GNDA.n1737 GNDA.n1590 585
R9864 GNDA.n1739 GNDA.n1589 585
R9865 GNDA.n1739 GNDA.n1738 585
R9866 GNDA.n1716 GNDA.n103 585
R9867 GNDA.n5092 GNDA.n5091 585
R9868 GNDA.n5094 GNDA.n88 585
R9869 GNDA.n5165 GNDA.n5164 585
R9870 GNDA.n24 GNDA.n22 585
R9871 GNDA.n5263 GNDA.n5262 585
R9872 GNDA.n32 GNDA.n25 585
R9873 GNDA.n40 GNDA.n39 585
R9874 GNDA.n35 GNDA.n31 585
R9875 GNDA.n30 GNDA.n0 585
R9876 GNDA.n5099 GNDA.n1 585
R9877 GNDA.n5101 GNDA.n5100 585
R9878 GNDA.n5105 GNDA.n5104 585
R9879 GNDA.n5107 GNDA.n5106 585
R9880 GNDA.n5096 GNDA.n5095 585
R9881 GNDA.n5086 GNDA.n89 585
R9882 GNDA.n5090 GNDA.n89 585
R9883 GNDA.n5088 GNDA.n5087 585
R9884 GNDA.n5089 GNDA.n5088 585
R9885 GNDA.n5085 GNDA.n91 585
R9886 GNDA.n91 GNDA.n90 585
R9887 GNDA.n5084 GNDA.n5083 585
R9888 GNDA.n5083 GNDA.n5082 585
R9889 GNDA.n93 GNDA.n92 585
R9890 GNDA.n5081 GNDA.n93 585
R9891 GNDA.n4629 GNDA.n4628 585
R9892 GNDA.n4628 GNDA.n110 585
R9893 GNDA.n4631 GNDA.n4630 585
R9894 GNDA.n4632 GNDA.n4631 585
R9895 GNDA.n427 GNDA.n426 585
R9896 GNDA.n4633 GNDA.n427 585
R9897 GNDA.n4636 GNDA.n4635 585
R9898 GNDA.n4635 GNDA.n4634 585
R9899 GNDA.n4637 GNDA.n425 585
R9900 GNDA.n425 GNDA.n424 585
R9901 GNDA.n4639 GNDA.n4638 585
R9902 GNDA.n4640 GNDA.n4639 585
R9903 GNDA.n423 GNDA.n422 585
R9904 GNDA.n4641 GNDA.n423 585
R9905 GNDA.n4644 GNDA.n4643 585
R9906 GNDA.n4643 GNDA.n4642 585
R9907 GNDA.n4645 GNDA.n421 585
R9908 GNDA.n421 GNDA.n420 585
R9909 GNDA.n4647 GNDA.n4646 585
R9910 GNDA.n4648 GNDA.n4647 585
R9911 GNDA.n419 GNDA.n418 585
R9912 GNDA.n4649 GNDA.n419 585
R9913 GNDA.n4652 GNDA.n4651 585
R9914 GNDA.n4651 GNDA.n4650 585
R9915 GNDA.n4653 GNDA.n417 585
R9916 GNDA.n417 GNDA.n416 585
R9917 GNDA.n4655 GNDA.n4654 585
R9918 GNDA.n4656 GNDA.n4655 585
R9919 GNDA.n415 GNDA.n414 585
R9920 GNDA.n4657 GNDA.n415 585
R9921 GNDA.n4660 GNDA.n4659 585
R9922 GNDA.n4659 GNDA.n4658 585
R9923 GNDA.n4661 GNDA.n413 585
R9924 GNDA.n413 GNDA.n367 585
R9925 GNDA.n4663 GNDA.n4662 585
R9926 GNDA.n4664 GNDA.n4663 585
R9927 GNDA.n4668 GNDA.n4667 585
R9928 GNDA.n4667 GNDA.n4666 585
R9929 GNDA.n4669 GNDA.n363 585
R9930 GNDA.n363 GNDA.n362 585
R9931 GNDA.n4671 GNDA.n4670 585
R9932 GNDA.n4672 GNDA.n4671 585
R9933 GNDA.n364 GNDA.n361 585
R9934 GNDA.n4673 GNDA.n361 585
R9935 GNDA.n4675 GNDA.n360 585
R9936 GNDA.n4675 GNDA.n4674 585
R9937 GNDA.n4677 GNDA.n4676 585
R9938 GNDA.n4676 GNDA.n356 585
R9939 GNDA.n354 GNDA.n353 585
R9940 GNDA.n4683 GNDA.n354 585
R9941 GNDA.n4686 GNDA.n4685 585
R9942 GNDA.n4685 GNDA.n4684 585
R9943 GNDA.n4687 GNDA.n352 585
R9944 GNDA.n352 GNDA.n351 585
R9945 GNDA.n4689 GNDA.n4688 585
R9946 GNDA.n4690 GNDA.n4689 585
R9947 GNDA.n350 GNDA.n303 585
R9948 GNDA.n4691 GNDA.n350 585
R9949 GNDA.n4694 GNDA.n4693 585
R9950 GNDA.n4693 GNDA.n4692 585
R9951 GNDA.n389 GNDA.n83 585
R9952 GNDA.n390 GNDA.n388 585
R9953 GNDA.n395 GNDA.n386 585
R9954 GNDA.n396 GNDA.n384 585
R9955 GNDA.n397 GNDA.n383 585
R9956 GNDA.n381 GNDA.n379 585
R9957 GNDA.n403 GNDA.n378 585
R9958 GNDA.n404 GNDA.n376 585
R9959 GNDA.n405 GNDA.n375 585
R9960 GNDA.n373 GNDA.n371 585
R9961 GNDA.n410 GNDA.n370 585
R9962 GNDA.n411 GNDA.n366 585
R9963 GNDA.n5168 GNDA.n84 585
R9964 GNDA.n5168 GNDA.n5167 585
R9965 GNDA.n412 GNDA.n411 585
R9966 GNDA.n410 GNDA.n409 585
R9967 GNDA.n408 GNDA.n371 585
R9968 GNDA.n406 GNDA.n405 585
R9969 GNDA.n404 GNDA.n372 585
R9970 GNDA.n403 GNDA.n402 585
R9971 GNDA.n400 GNDA.n379 585
R9972 GNDA.n398 GNDA.n397 585
R9973 GNDA.n396 GNDA.n380 585
R9974 GNDA.n395 GNDA.n394 585
R9975 GNDA.n392 GNDA.n390 585
R9976 GNDA.n389 GNDA.n86 585
R9977 GNDA.n5166 GNDA.n84 585
R9978 GNDA.n5167 GNDA.n5166 585
R9979 GNDA.n1796 GNDA.n1795 585
R9980 GNDA.n1793 GNDA.n1554 585
R9981 GNDA.n1792 GNDA.n1791 585
R9982 GNDA.n1783 GNDA.n1556 585
R9983 GNDA.n1785 GNDA.n1784 585
R9984 GNDA.n1781 GNDA.n1558 585
R9985 GNDA.n1780 GNDA.n1779 585
R9986 GNDA.n1771 GNDA.n1560 585
R9987 GNDA.n1773 GNDA.n1772 585
R9988 GNDA.n1769 GNDA.n1562 585
R9989 GNDA.n1768 GNDA.n1767 585
R9990 GNDA.n1585 GNDA.n1564 585
R9991 GNDA.n1799 GNDA.n1551 585
R9992 GNDA.n1551 GNDA.n161 585
R9993 GNDA.n1764 GNDA.n1564 585
R9994 GNDA.n1767 GNDA.n1766 585
R9995 GNDA.n1562 GNDA.n1561 585
R9996 GNDA.n1561 GNDA.n111 585
R9997 GNDA.n1774 GNDA.n1773 585
R9998 GNDA.n1776 GNDA.n1560 585
R9999 GNDA.n1779 GNDA.n1778 585
R10000 GNDA.n1558 GNDA.n1557 585
R10001 GNDA.n1786 GNDA.n1785 585
R10002 GNDA.n1788 GNDA.n1556 585
R10003 GNDA.n1791 GNDA.n1790 585
R10004 GNDA.n1554 GNDA.n1553 585
R10005 GNDA.n1797 GNDA.n1796 585
R10006 GNDA.n1797 GNDA.n111 585
R10007 GNDA.n1799 GNDA.n1798 585
R10008 GNDA.n1798 GNDA.n161 585
R10009 GNDA.n3148 GNDA.n3147 585
R10010 GNDA.n3149 GNDA.n1823 585
R10011 GNDA.n1822 GNDA.n1819 585
R10012 GNDA.n3155 GNDA.n1818 585
R10013 GNDA.n3156 GNDA.n1817 585
R10014 GNDA.n3157 GNDA.n1815 585
R10015 GNDA.n1814 GNDA.n1811 585
R10016 GNDA.n3162 GNDA.n1810 585
R10017 GNDA.n3163 GNDA.n1809 585
R10018 GNDA.n1807 GNDA.n1805 585
R10019 GNDA.n3167 GNDA.n1804 585
R10020 GNDA.n3168 GNDA.n1802 585
R10021 GNDA.n3169 GNDA.n3168 585
R10022 GNDA.n3167 GNDA.n3166 585
R10023 GNDA.n3165 GNDA.n1805 585
R10024 GNDA.n3165 GNDA.n1519 585
R10025 GNDA.n3164 GNDA.n3163 585
R10026 GNDA.n3162 GNDA.n3161 585
R10027 GNDA.n3160 GNDA.n1811 585
R10028 GNDA.n3158 GNDA.n3157 585
R10029 GNDA.n3156 GNDA.n1812 585
R10030 GNDA.n3155 GNDA.n3154 585
R10031 GNDA.n3152 GNDA.n1819 585
R10032 GNDA.n3150 GNDA.n3149 585
R10033 GNDA.n3148 GNDA.n1820 585
R10034 GNDA.n1820 GNDA.n1519 585
R10035 GNDA.n2708 GNDA.n2705 585
R10036 GNDA.n2710 GNDA.n2709 585
R10037 GNDA.n2709 GNDA.n1497 585
R10038 GNDA.n2719 GNDA.n2718 585
R10039 GNDA.n2807 GNDA.n2806 585
R10040 GNDA.n2806 GNDA.n2805 585
R10041 GNDA.n2816 GNDA.n2694 585
R10042 GNDA.n2823 GNDA.n2693 585
R10043 GNDA.n2827 GNDA.n2693 585
R10044 GNDA.n2821 GNDA.n2820 585
R10045 GNDA.n3236 GNDA.n1523 585
R10046 GNDA.n3240 GNDA.n1522 585
R10047 GNDA.n3248 GNDA.n1522 585
R10048 GNDA.n3239 GNDA.n3238 585
R10049 GNDA.n3044 GNDA.n1832 585
R10050 GNDA.n3045 GNDA.n3044 585
R10051 GNDA.n2935 GNDA.n2934 585
R10052 GNDA.n2934 GNDA.n2933 585
R10053 GNDA.n2907 GNDA.n1858 585
R10054 GNDA.n2932 GNDA.n1858 585
R10055 GNDA.n2908 GNDA.n2664 585
R10056 GNDA.n2664 GNDA.n1859 585
R10057 GNDA.n2916 GNDA.n2915 585
R10058 GNDA.n2917 GNDA.n2916 585
R10059 GNDA.n2668 GNDA.n2666 585
R10060 GNDA.n2666 GNDA.n2665 585
R10061 GNDA.n2832 GNDA.n2831 585
R10062 GNDA.n2831 GNDA.n106 585
R10063 GNDA.n2833 GNDA.n2829 585
R10064 GNDA.n2829 GNDA.n2828 585
R10065 GNDA.n2842 GNDA.n2841 585
R10066 GNDA.n2843 GNDA.n2842 585
R10067 GNDA.n2689 GNDA.n2688 585
R10068 GNDA.n2844 GNDA.n2689 585
R10069 GNDA.n2849 GNDA.n2848 585
R10070 GNDA.n2848 GNDA.n2847 585
R10071 GNDA.n2691 GNDA.n2690 585
R10072 GNDA.n2846 GNDA.n2691 585
R10073 GNDA.n2731 GNDA.n1831 585
R10074 GNDA.n2845 GNDA.n1831 585
R10075 GNDA.n3146 GNDA.n1827 585
R10076 GNDA.n3146 GNDA.n3145 585
R10077 GNDA.n2733 GNDA.n1832 585
R10078 GNDA.n2733 GNDA.n1830 585
R10079 GNDA.n2739 GNDA.n2738 585
R10080 GNDA.n2738 GNDA.n2737 585
R10081 GNDA.n1495 GNDA.n1493 585
R10082 GNDA.n3278 GNDA.n1495 585
R10083 GNDA.n3293 GNDA.n3292 585
R10084 GNDA.n3292 GNDA.n3291 585
R10085 GNDA.n3280 GNDA.n1496 585
R10086 GNDA.n3290 GNDA.n1496 585
R10087 GNDA.n3288 GNDA.n3287 585
R10088 GNDA.n3289 GNDA.n3288 585
R10089 GNDA.n3283 GNDA.n1470 585
R10090 GNDA.n3279 GNDA.n1470 585
R10091 GNDA.n3301 GNDA.n3300 585
R10092 GNDA.n3302 GNDA.n3301 585
R10093 GNDA.n1472 GNDA.n1471 585
R10094 GNDA.n2723 GNDA.n1471 585
R10095 GNDA.n2726 GNDA.n2725 585
R10096 GNDA.n2725 GNDA.n2724 585
R10097 GNDA.n2729 GNDA.n2721 585
R10098 GNDA.n2721 GNDA.n2720 585
R10099 GNDA.n2798 GNDA.n2797 585
R10100 GNDA.n2799 GNDA.n2798 585
R10101 GNDA.n2795 GNDA.n1826 585
R10102 GNDA.n2802 GNDA.n1826 585
R10103 GNDA.n3143 GNDA.n1827 585
R10104 GNDA.n3144 GNDA.n3143 585
R10105 GNDA.n3142 GNDA.n3139 585
R10106 GNDA.n3142 GNDA.n3141 585
R10107 GNDA.n3137 GNDA.n3046 585
R10108 GNDA.n3140 GNDA.n3046 585
R10109 GNDA.n3117 GNDA.n3048 585
R10110 GNDA.n3128 GNDA.n3117 585
R10111 GNDA.n3132 GNDA.n3131 585
R10112 GNDA.n3131 GNDA.n3130 585
R10113 GNDA.n3127 GNDA.n3126 585
R10114 GNDA.n3129 GNDA.n3127 585
R10115 GNDA.n3121 GNDA.n3118 585
R10116 GNDA.n3118 GNDA.n1520 585
R10117 GNDA.n3119 GNDA.n1516 585
R10118 GNDA.n3249 GNDA.n1516 585
R10119 GNDA.n3252 GNDA.n3251 585
R10120 GNDA.n3251 GNDA.n3250 585
R10121 GNDA.n1513 GNDA.n1508 585
R10122 GNDA.n1508 GNDA.n1506 585
R10123 GNDA.n3262 GNDA.n3261 585
R10124 GNDA.n3263 GNDA.n3262 585
R10125 GNDA.n1511 GNDA.n1509 585
R10126 GNDA.n1509 GNDA.n1507 585
R10127 GNDA.n3220 GNDA.n3219 585
R10128 GNDA.n3221 GNDA.n3220 585
R10129 GNDA.n2957 GNDA.n1855 585
R10130 GNDA.n2956 GNDA.n2955 585
R10131 GNDA.n2954 GNDA.n2953 585
R10132 GNDA.n2952 GNDA.n2951 585
R10133 GNDA.n2950 GNDA.n2949 585
R10134 GNDA.n2948 GNDA.n2947 585
R10135 GNDA.n2946 GNDA.n2945 585
R10136 GNDA.n2944 GNDA.n2943 585
R10137 GNDA.n2942 GNDA.n2941 585
R10138 GNDA.n2940 GNDA.n2939 585
R10139 GNDA.n2938 GNDA.n2937 585
R10140 GNDA.n4860 GNDA.n280 585
R10141 GNDA.n262 GNDA.n261 585
R10142 GNDA.n264 GNDA.n263 585
R10143 GNDA.n266 GNDA.n265 585
R10144 GNDA.n268 GNDA.n267 585
R10145 GNDA.n270 GNDA.n269 585
R10146 GNDA.n272 GNDA.n271 585
R10147 GNDA.n274 GNDA.n273 585
R10148 GNDA.n275 GNDA.n240 585
R10149 GNDA.n278 GNDA.n277 585
R10150 GNDA.n276 GNDA.n239 585
R10151 GNDA.n229 GNDA.n228 585
R10152 GNDA.n4860 GNDA.n229 585
R10153 GNDA.n4863 GNDA.n4862 585
R10154 GNDA.n4863 GNDA.n227 585
R10155 GNDA.n4858 GNDA.n4857 585
R10156 GNDA.n4856 GNDA.n288 585
R10157 GNDA.n4855 GNDA.n287 585
R10158 GNDA.n4860 GNDA.n287 585
R10159 GNDA.n4854 GNDA.n4853 585
R10160 GNDA.n4852 GNDA.n4851 585
R10161 GNDA.n4850 GNDA.n4849 585
R10162 GNDA.n4848 GNDA.n4847 585
R10163 GNDA.n4846 GNDA.n4845 585
R10164 GNDA.n4844 GNDA.n4843 585
R10165 GNDA.n4842 GNDA.n4841 585
R10166 GNDA.n4840 GNDA.n4839 585
R10167 GNDA.n4838 GNDA.n4837 585
R10168 GNDA.n4837 GNDA.n4836 585
R10169 GNDA.n3385 GNDA.t114 524.808
R10170 GNDA.n3380 GNDA.t103 524.808
R10171 GNDA.n4610 GNDA.t132 524.808
R10172 GNDA.n3851 GNDA.t142 524.808
R10173 GNDA.n3614 GNDA.t129 508.743
R10174 GNDA.n1452 GNDA.t94 508.743
R10175 GNDA.n583 GNDA.t76 508.743
R10176 GNDA.n3335 GNDA.t73 508.743
R10177 GNDA.n3607 GNDA.t88 499.442
R10178 GNDA.n3338 GNDA.t79 499.442
R10179 GNDA.n572 GNDA.t148 499.442
R10180 GNDA.n3326 GNDA.t137 499.442
R10181 GNDA.t62 GNDA.n88 486.94
R10182 GNDA.t62 GNDA.n103 486.94
R10183 GNDA.n3579 GNDA.t135 475.976
R10184 GNDA.n3579 GNDA.t111 475.976
R10185 GNDA.n3575 GNDA.t146 475.976
R10186 GNDA.n3575 GNDA.t126 475.976
R10187 GNDA.n2929 GNDA.t107 425.134
R10188 GNDA.n2658 GNDA.t64 409.067
R10189 GNDA.n3266 GNDA.t155 409.067
R10190 GNDA.n1502 GNDA.t91 409.067
R10191 GNDA.n1501 GNDA.t58 409.067
R10192 GNDA.n3275 GNDA.t97 409.067
R10193 GNDA.n2734 GNDA.t70 409.067
R10194 GNDA.n2920 GNDA.t158 409.067
R10195 GNDA.n4640 GNDA.n424 394.817
R10196 GNDA.n4634 GNDA.n4633 394.817
R10197 GNDA.n4633 GNDA.n4632 394.817
R10198 GNDA.n4632 GNDA.n110 394.817
R10199 GNDA.n5082 GNDA.n5081 394.817
R10200 GNDA.n5082 GNDA.n90 394.817
R10201 GNDA.n5089 GNDA.n90 394.817
R10202 GNDA.n5090 GNDA.n5089 394.817
R10203 GNDA.n5091 GNDA.n5090 394.817
R10204 GNDA.n5091 GNDA.n88 394.817
R10205 GNDA.n1738 GNDA.n1737 394.817
R10206 GNDA.n1737 GNDA.n1736 394.817
R10207 GNDA.n1736 GNDA.n1591 394.817
R10208 GNDA.n1730 GNDA.n1591 394.817
R10209 GNDA.n1730 GNDA.n109 394.817
R10210 GNDA.n1598 GNDA.n108 394.817
R10211 GNDA.n1723 GNDA.n1598 394.817
R10212 GNDA.n1723 GNDA.n1722 394.817
R10213 GNDA.n1722 GNDA.n1721 394.817
R10214 GNDA.n1721 GNDA.n1599 394.817
R10215 GNDA.n1599 GNDA.n103 394.817
R10216 GNDA.n1541 GNDA.n102 394.817
R10217 GNDA.n3200 GNDA.n1541 394.817
R10218 GNDA.n3201 GNDA.n3200 394.817
R10219 GNDA.n3202 GNDA.n3201 394.817
R10220 GNDA.n3202 GNDA.n1517 394.817
R10221 GNDA.n1536 GNDA.n1518 394.817
R10222 GNDA.n3210 GNDA.n1536 394.817
R10223 GNDA.n3211 GNDA.n3210 394.817
R10224 GNDA.n3215 GNDA.n3211 394.817
R10225 GNDA.n3215 GNDA.n3214 394.817
R10226 GNDA.n3214 GNDA.n3213 394.817
R10227 GNDA.n3325 GNDA.n3324 386.587
R10228 GNDA.n4627 GNDA.n424 377.269
R10229 GNDA.n300 GNDA.n96 370.214
R10230 GNDA.n4665 GNDA.n98 370.214
R10231 GNDA.n300 GNDA.n95 365.957
R10232 GNDA.n4665 GNDA.n97 365.957
R10233 GNDA.n3306 GNDA.n429 334.178
R10234 GNDA.n4624 GNDA.n430 328.358
R10235 GNDA.t62 GNDA.n94 172.876
R10236 GNDA.t62 GNDA.n95 327.661
R10237 GNDA.t62 GNDA.n97 327.661
R10238 GNDA.t62 GNDA.n1469 172.876
R10239 GNDA.t62 GNDA.n1468 172.615
R10240 GNDA.t62 GNDA.n96 323.404
R10241 GNDA.t62 GNDA.n98 323.404
R10242 GNDA.t62 GNDA.n1519 172.615
R10243 GNDA.n3613 GNDA.n3612 296.158
R10244 GNDA.n1451 GNDA.n1450 296.158
R10245 GNDA.n3584 GNDA.n584 296.158
R10246 GNDA.n3571 GNDA.n588 296.158
R10247 GNDA.n3340 GNDA.n3327 292.5
R10248 GNDA.n3572 GNDA.n3571 292.5
R10249 GNDA.n3584 GNDA.n3583 292.5
R10250 GNDA.n3609 GNDA.n573 292.5
R10251 GNDA.n3340 GNDA.n3339 292.5
R10252 GNDA.n3609 GNDA.n3608 292.5
R10253 GNDA.t62 GNDA.n110 267.598
R10254 GNDA.t62 GNDA.n109 267.598
R10255 GNDA.t62 GNDA.n1517 267.598
R10256 GNDA.n3218 GNDA.n1532 264.301
R10257 GNDA.n1718 GNDA.n1717 264.301
R10258 GNDA.n5093 GNDA.n87 264.301
R10259 GNDA.n2936 GNDA.n1856 264.301
R10260 GNDA.n4861 GNDA.n4860 264.301
R10261 GNDA.n4860 GNDA.n234 264.301
R10262 GNDA.t176 GNDA.n1528 260
R10263 GNDA.n3225 GNDA.t176 260
R10264 GNDA.n3194 GNDA.n3193 259.416
R10265 GNDA.n2992 GNDA.n1802 259.416
R10266 GNDA.n3016 GNDA.n1849 259.416
R10267 GNDA.n4667 GNDA.n366 259.416
R10268 GNDA.n1740 GNDA.n1739 259.416
R10269 GNDA.n1586 GNDA.n1585 259.416
R10270 GNDA.n5078 GNDA.n130 259.416
R10271 GNDA.n4697 GNDA.n301 259.416
R10272 GNDA.n4639 GNDA.n423 259.416
R10273 GNDA.n3098 GNDA.n3096 258.334
R10274 GNDA.n2758 GNDA.n2757 258.334
R10275 GNDA.n5023 GNDA.n5022 258.334
R10276 GNDA.n4808 GNDA.n4807 258.334
R10277 GNDA.n1659 GNDA.n1658 258.334
R10278 GNDA.n4947 GNDA.n4887 258.334
R10279 GNDA.n5226 GNDA.n80 258.334
R10280 GNDA.n2889 GNDA.n2674 258.334
R10281 GNDA.n5146 GNDA.n5145 258.334
R10282 GNDA.t62 GNDA.n4682 257.779
R10283 GNDA.n5080 GNDA.n5079 254.34
R10284 GNDA.n5080 GNDA.n128 254.34
R10285 GNDA.n5080 GNDA.n127 254.34
R10286 GNDA.n5080 GNDA.n126 254.34
R10287 GNDA.n5080 GNDA.n125 254.34
R10288 GNDA.n5080 GNDA.n124 254.34
R10289 GNDA.n5080 GNDA.n123 254.34
R10290 GNDA.n5080 GNDA.n122 254.34
R10291 GNDA.n5080 GNDA.n121 254.34
R10292 GNDA.n5080 GNDA.n120 254.34
R10293 GNDA.n5080 GNDA.n119 254.34
R10294 GNDA.n5080 GNDA.n118 254.34
R10295 GNDA.n5080 GNDA.n117 254.34
R10296 GNDA.n5080 GNDA.n116 254.34
R10297 GNDA.n5080 GNDA.n115 254.34
R10298 GNDA.n5080 GNDA.n114 254.34
R10299 GNDA.n5080 GNDA.n113 254.34
R10300 GNDA.n5080 GNDA.n112 254.34
R10301 GNDA.n5260 GNDA.n5259 254.34
R10302 GNDA.n5260 GNDA.n53 254.34
R10303 GNDA.n5260 GNDA.n52 254.34
R10304 GNDA.n5260 GNDA.n51 254.34
R10305 GNDA.n5260 GNDA.n50 254.34
R10306 GNDA.n5260 GNDA.n49 254.34
R10307 GNDA.n5260 GNDA.n48 254.34
R10308 GNDA.n5260 GNDA.n47 254.34
R10309 GNDA.n5260 GNDA.n46 254.34
R10310 GNDA.n5260 GNDA.n45 254.34
R10311 GNDA.n5260 GNDA.n44 254.34
R10312 GNDA.n5260 GNDA.n43 254.34
R10313 GNDA.n324 GNDA.n95 254.34
R10314 GNDA.n321 GNDA.n95 254.34
R10315 GNDA.n316 GNDA.n95 254.34
R10316 GNDA.n313 GNDA.n95 254.34
R10317 GNDA.n308 GNDA.n95 254.34
R10318 GNDA.n305 GNDA.n95 254.34
R10319 GNDA.n348 GNDA.n96 254.34
R10320 GNDA.n342 GNDA.n96 254.34
R10321 GNDA.n340 GNDA.n96 254.34
R10322 GNDA.n334 GNDA.n96 254.34
R10323 GNDA.n332 GNDA.n96 254.34
R10324 GNDA.n326 GNDA.n96 254.34
R10325 GNDA.n158 GNDA.n157 254.34
R10326 GNDA.n157 GNDA.n156 254.34
R10327 GNDA.n157 GNDA.n155 254.34
R10328 GNDA.n157 GNDA.n154 254.34
R10329 GNDA.n157 GNDA.n153 254.34
R10330 GNDA.n157 GNDA.n152 254.34
R10331 GNDA.n5073 GNDA.n5072 254.34
R10332 GNDA.n5072 GNDA.n5071 254.34
R10333 GNDA.n5072 GNDA.n140 254.34
R10334 GNDA.n5072 GNDA.n139 254.34
R10335 GNDA.n5072 GNDA.n138 254.34
R10336 GNDA.n5072 GNDA.n137 254.34
R10337 GNDA.n3042 GNDA.n94 254.34
R10338 GNDA.n1840 GNDA.n94 254.34
R10339 GNDA.n3031 GNDA.n94 254.34
R10340 GNDA.n3028 GNDA.n94 254.34
R10341 GNDA.n3019 GNDA.n94 254.34
R10342 GNDA.n3017 GNDA.n94 254.34
R10343 GNDA.n3013 GNDA.n1468 254.34
R10344 GNDA.n3024 GNDA.n1468 254.34
R10345 GNDA.n1845 GNDA.n1468 254.34
R10346 GNDA.n3035 GNDA.n1468 254.34
R10347 GNDA.n3038 GNDA.n1468 254.34
R10348 GNDA.n2978 GNDA.n104 254.34
R10349 GNDA.n2976 GNDA.n104 254.34
R10350 GNDA.n2970 GNDA.n104 254.34
R10351 GNDA.n2968 GNDA.n104 254.34
R10352 GNDA.n2962 GNDA.n104 254.34
R10353 GNDA.n2960 GNDA.n104 254.34
R10354 GNDA.n2991 GNDA.n104 254.34
R10355 GNDA.n2997 GNDA.n104 254.34
R10356 GNDA.n2989 GNDA.n104 254.34
R10357 GNDA.n3004 GNDA.n104 254.34
R10358 GNDA.n2986 GNDA.n104 254.34
R10359 GNDA.n3011 GNDA.n104 254.34
R10360 GNDA.n3192 GNDA.n104 254.34
R10361 GNDA.n3186 GNDA.n104 254.34
R10362 GNDA.n3184 GNDA.n104 254.34
R10363 GNDA.n3178 GNDA.n104 254.34
R10364 GNDA.n3176 GNDA.n104 254.34
R10365 GNDA.n3170 GNDA.n104 254.34
R10366 GNDA.n4981 GNDA.n4980 254.34
R10367 GNDA.n4981 GNDA.n225 254.34
R10368 GNDA.n4981 GNDA.n224 254.34
R10369 GNDA.n4981 GNDA.n223 254.34
R10370 GNDA.n4981 GNDA.n222 254.34
R10371 GNDA.n4981 GNDA.n221 254.34
R10372 GNDA.n4981 GNDA.n163 254.34
R10373 GNDA.n4981 GNDA.n166 254.34
R10374 GNDA.n4981 GNDA.n220 254.34
R10375 GNDA.n4981 GNDA.n197 254.34
R10376 GNDA.n4981 GNDA.n196 254.34
R10377 GNDA.n4982 GNDA.n4981 254.34
R10378 GNDA.n4981 GNDA.n195 254.34
R10379 GNDA.n4981 GNDA.n194 254.34
R10380 GNDA.n4981 GNDA.n193 254.34
R10381 GNDA.n4981 GNDA.n192 254.34
R10382 GNDA.n4981 GNDA.n191 254.34
R10383 GNDA.n4981 GNDA.n190 254.34
R10384 GNDA.n5260 GNDA.n42 254.34
R10385 GNDA.n5261 GNDA.n5260 254.34
R10386 GNDA.n5260 GNDA.n41 254.34
R10387 GNDA.n5260 GNDA.n29 254.34
R10388 GNDA.n5260 GNDA.n28 254.34
R10389 GNDA.n5260 GNDA.n27 254.34
R10390 GNDA.n387 GNDA.n97 254.34
R10391 GNDA.n385 GNDA.n97 254.34
R10392 GNDA.n382 GNDA.n97 254.34
R10393 GNDA.n377 GNDA.n97 254.34
R10394 GNDA.n374 GNDA.n97 254.34
R10395 GNDA.n369 GNDA.n97 254.34
R10396 GNDA.n368 GNDA.n98 254.34
R10397 GNDA.n407 GNDA.n98 254.34
R10398 GNDA.n401 GNDA.n98 254.34
R10399 GNDA.n399 GNDA.n98 254.34
R10400 GNDA.n393 GNDA.n98 254.34
R10401 GNDA.n391 GNDA.n98 254.34
R10402 GNDA.n1794 GNDA.n101 254.34
R10403 GNDA.n1555 GNDA.n101 254.34
R10404 GNDA.n1782 GNDA.n101 254.34
R10405 GNDA.n1559 GNDA.n101 254.34
R10406 GNDA.n1770 GNDA.n101 254.34
R10407 GNDA.n1563 GNDA.n101 254.34
R10408 GNDA.n1765 GNDA.n111 254.34
R10409 GNDA.n1775 GNDA.n111 254.34
R10410 GNDA.n1777 GNDA.n111 254.34
R10411 GNDA.n1787 GNDA.n111 254.34
R10412 GNDA.n1789 GNDA.n111 254.34
R10413 GNDA.n1825 GNDA.n1469 254.34
R10414 GNDA.n1821 GNDA.n1469 254.34
R10415 GNDA.n1816 GNDA.n1469 254.34
R10416 GNDA.n1813 GNDA.n1469 254.34
R10417 GNDA.n1808 GNDA.n1469 254.34
R10418 GNDA.n1803 GNDA.n1469 254.34
R10419 GNDA.n1801 GNDA.n1519 254.34
R10420 GNDA.n1806 GNDA.n1519 254.34
R10421 GNDA.n3159 GNDA.n1519 254.34
R10422 GNDA.n3153 GNDA.n1519 254.34
R10423 GNDA.n3151 GNDA.n1519 254.34
R10424 GNDA.n4860 GNDA.n286 254.34
R10425 GNDA.n4860 GNDA.n285 254.34
R10426 GNDA.n4860 GNDA.n284 254.34
R10427 GNDA.n4860 GNDA.n283 254.34
R10428 GNDA.n4860 GNDA.n282 254.34
R10429 GNDA.n4860 GNDA.n281 254.34
R10430 GNDA.n4860 GNDA.n235 254.34
R10431 GNDA.n4860 GNDA.n236 254.34
R10432 GNDA.n4860 GNDA.n237 254.34
R10433 GNDA.n4860 GNDA.n238 254.34
R10434 GNDA.n4860 GNDA.n279 254.34
R10435 GNDA.n4860 GNDA.n4859 254.34
R10436 GNDA.n4860 GNDA.n230 254.34
R10437 GNDA.n4860 GNDA.n231 254.34
R10438 GNDA.n4860 GNDA.n232 254.34
R10439 GNDA.n4860 GNDA.n233 254.34
R10440 GNDA.n2707 GNDA.n1497 250.349
R10441 GNDA.n2805 GNDA.n2804 250.349
R10442 GNDA.n3171 GNDA.n3169 249.663
R10443 GNDA.n3014 GNDA.n3012 249.663
R10444 GNDA.n2959 GNDA.n1855 249.663
R10445 GNDA.n4693 GNDA.n349 249.663
R10446 GNDA.n1764 GNDA.n1763 249.663
R10447 GNDA.n5074 GNDA.n135 249.663
R10448 GNDA.n261 GNDA.n260 249.663
R10449 GNDA.n4858 GNDA.n289 249.663
R10450 GNDA.n4663 GNDA.n412 249.663
R10451 GNDA.n1523 GNDA.n1522 246.25
R10452 GNDA.n3238 GNDA.n1522 246.25
R10453 GNDA.n2694 GNDA.n2693 246.25
R10454 GNDA.n2820 GNDA.n2693 246.25
R10455 GNDA.n3224 GNDA.n1529 246.25
R10456 GNDA.n2827 GNDA.n2826 241.643
R10457 GNDA.n2827 GNDA.n2692 241.643
R10458 GNDA.n3248 GNDA.n3247 241.643
R10459 GNDA.n3248 GNDA.n1521 241.643
R10460 GNDA.t15 GNDA.t108 227.873
R10461 GNDA.n3212 GNDA.t175 219.343
R10462 GNDA.n3223 GNDA.t175 219.343
R10463 GNDA.n3342 GNDA.n3341 197.133
R10464 GNDA.n3585 GNDA.n3584 197.133
R10465 GNDA.n3571 GNDA.n3570 197.133
R10466 GNDA.n3611 GNDA.n3610 197.133
R10467 GNDA.n4624 GNDA.n4623 197.016
R10468 GNDA.n2806 GNDA.n2719 197
R10469 GNDA.n2709 GNDA.n2708 197
R10470 GNDA.n3220 GNDA.n1530 197
R10471 GNDA.n3146 GNDA.n1826 197
R10472 GNDA.n3044 GNDA.n1831 197
R10473 GNDA.n1716 GNDA.n1715 197
R10474 GNDA.n1551 GNDA.n189 197
R10475 GNDA.n4890 GNDA.n4889 197
R10476 GNDA.n4741 GNDA.n85 197
R10477 GNDA.n5169 GNDA.n5168 197
R10478 GNDA.n5095 GNDA.n5094 197
R10479 GNDA.n3143 GNDA.n3142 187.249
R10480 GNDA.n2738 GNDA.n2733 187.249
R10481 GNDA.n2934 GNDA.n280 187.249
R10482 GNDA.n1798 GNDA.n1552 187.249
R10483 GNDA.n5051 GNDA.n5050 187.249
R10484 GNDA.n4979 GNDA.n227 187.249
R10485 GNDA.n4836 GNDA.n4835 187.249
R10486 GNDA.n5258 GNDA.n55 187.249
R10487 GNDA.n5166 GNDA.n5165 187.249
R10488 GNDA.n3099 GNDA.n3098 185
R10489 GNDA.n3100 GNDA.n3052 185
R10490 GNDA.n3102 GNDA.n3101 185
R10491 GNDA.n3104 GNDA.n3051 185
R10492 GNDA.n3107 GNDA.n3106 185
R10493 GNDA.n3108 GNDA.n3050 185
R10494 GNDA.n3110 GNDA.n3109 185
R10495 GNDA.n3112 GNDA.n3049 185
R10496 GNDA.n3113 GNDA.n3047 185
R10497 GNDA.n3080 GNDA.n3057 185
R10498 GNDA.n3083 GNDA.n3082 185
R10499 GNDA.n3084 GNDA.n3056 185
R10500 GNDA.n3086 GNDA.n3085 185
R10501 GNDA.n3088 GNDA.n3055 185
R10502 GNDA.n3091 GNDA.n3090 185
R10503 GNDA.n3092 GNDA.n3054 185
R10504 GNDA.n3094 GNDA.n3093 185
R10505 GNDA.n3096 GNDA.n3053 185
R10506 GNDA.n3062 GNDA.n1512 185
R10507 GNDA.n3066 GNDA.n3063 185
R10508 GNDA.n3068 GNDA.n3067 185
R10509 GNDA.n3069 GNDA.n3061 185
R10510 GNDA.n3071 GNDA.n3070 185
R10511 GNDA.n3073 GNDA.n3059 185
R10512 GNDA.n3075 GNDA.n3074 185
R10513 GNDA.n3076 GNDA.n3058 185
R10514 GNDA.n3078 GNDA.n3077 185
R10515 GNDA.n3260 GNDA.n3259 185
R10516 GNDA.n3257 GNDA.n1510 185
R10517 GNDA.n3256 GNDA.n1514 185
R10518 GNDA.n3254 GNDA.n3253 185
R10519 GNDA.n3120 GNDA.n1515 185
R10520 GNDA.n3125 GNDA.n3124 185
R10521 GNDA.n3122 GNDA.n3116 185
R10522 GNDA.n3134 GNDA.n3133 185
R10523 GNDA.n3136 GNDA.n3135 185
R10524 GNDA.n2757 GNDA.n2756 185
R10525 GNDA.n2755 GNDA.n2754 185
R10526 GNDA.n2753 GNDA.n2752 185
R10527 GNDA.n2751 GNDA.n2750 185
R10528 GNDA.n2749 GNDA.n2748 185
R10529 GNDA.n2747 GNDA.n2746 185
R10530 GNDA.n2745 GNDA.n2744 185
R10531 GNDA.n2743 GNDA.n2742 185
R10532 GNDA.n2741 GNDA.n1491 185
R10533 GNDA.n2775 GNDA.n2774 185
R10534 GNDA.n2773 GNDA.n2772 185
R10535 GNDA.n2771 GNDA.n2770 185
R10536 GNDA.n2769 GNDA.n2768 185
R10537 GNDA.n2767 GNDA.n2766 185
R10538 GNDA.n2765 GNDA.n2764 185
R10539 GNDA.n2763 GNDA.n2762 185
R10540 GNDA.n2761 GNDA.n2760 185
R10541 GNDA.n2759 GNDA.n2758 185
R10542 GNDA.n2794 GNDA.n2793 185
R10543 GNDA.n2791 GNDA.n2790 185
R10544 GNDA.n2789 GNDA.n2788 185
R10545 GNDA.n2787 GNDA.n2786 185
R10546 GNDA.n2785 GNDA.n2784 185
R10547 GNDA.n2783 GNDA.n2782 185
R10548 GNDA.n2781 GNDA.n2780 185
R10549 GNDA.n2779 GNDA.n2778 185
R10550 GNDA.n2777 GNDA.n2776 185
R10551 GNDA.n2792 GNDA.n2730 185
R10552 GNDA.n2728 GNDA.n2727 185
R10553 GNDA.n2722 GNDA.n1474 185
R10554 GNDA.n3299 GNDA.n3298 185
R10555 GNDA.n3282 GNDA.n1473 185
R10556 GNDA.n3286 GNDA.n3285 185
R10557 GNDA.n3284 GNDA.n3281 185
R10558 GNDA.n1494 GNDA.n1492 185
R10559 GNDA.n3295 GNDA.n3294 185
R10560 GNDA.n5024 GNDA.n5023 185
R10561 GNDA.n5026 GNDA.n5025 185
R10562 GNDA.n5028 GNDA.n5027 185
R10563 GNDA.n5030 GNDA.n5029 185
R10564 GNDA.n5032 GNDA.n5031 185
R10565 GNDA.n5034 GNDA.n5033 185
R10566 GNDA.n5036 GNDA.n5035 185
R10567 GNDA.n5038 GNDA.n5037 185
R10568 GNDA.n5039 GNDA.n164 185
R10569 GNDA.n5006 GNDA.n5005 185
R10570 GNDA.n5008 GNDA.n5007 185
R10571 GNDA.n5010 GNDA.n5009 185
R10572 GNDA.n5012 GNDA.n5011 185
R10573 GNDA.n5014 GNDA.n5013 185
R10574 GNDA.n5016 GNDA.n5015 185
R10575 GNDA.n5018 GNDA.n5017 185
R10576 GNDA.n5020 GNDA.n5019 185
R10577 GNDA.n5022 GNDA.n5021 185
R10578 GNDA.n4988 GNDA.n4987 185
R10579 GNDA.n4990 GNDA.n4989 185
R10580 GNDA.n4992 GNDA.n4991 185
R10581 GNDA.n4994 GNDA.n4993 185
R10582 GNDA.n4996 GNDA.n4995 185
R10583 GNDA.n4998 GNDA.n4997 185
R10584 GNDA.n5000 GNDA.n4999 185
R10585 GNDA.n5002 GNDA.n5001 185
R10586 GNDA.n5004 GNDA.n5003 185
R10587 GNDA.n4986 GNDA.n4985 185
R10588 GNDA.n206 GNDA.n205 185
R10589 GNDA.n204 GNDA.n203 185
R10590 GNDA.n212 GNDA.n211 185
R10591 GNDA.n214 GNDA.n213 185
R10592 GNDA.n217 GNDA.n216 185
R10593 GNDA.n200 GNDA.n169 185
R10594 GNDA.n5043 GNDA.n5042 185
R10595 GNDA.n168 GNDA.n165 185
R10596 GNDA.n4809 GNDA.n4808 185
R10597 GNDA.n4811 GNDA.n4810 185
R10598 GNDA.n4813 GNDA.n4812 185
R10599 GNDA.n4815 GNDA.n4814 185
R10600 GNDA.n4817 GNDA.n4816 185
R10601 GNDA.n4819 GNDA.n4818 185
R10602 GNDA.n4821 GNDA.n4820 185
R10603 GNDA.n4823 GNDA.n4822 185
R10604 GNDA.n4824 GNDA.n4720 185
R10605 GNDA.n4791 GNDA.n4790 185
R10606 GNDA.n4793 GNDA.n4792 185
R10607 GNDA.n4795 GNDA.n4794 185
R10608 GNDA.n4797 GNDA.n4796 185
R10609 GNDA.n4799 GNDA.n4798 185
R10610 GNDA.n4801 GNDA.n4800 185
R10611 GNDA.n4803 GNDA.n4802 185
R10612 GNDA.n4805 GNDA.n4804 185
R10613 GNDA.n4807 GNDA.n4806 185
R10614 GNDA.n4773 GNDA.n4772 185
R10615 GNDA.n4775 GNDA.n4774 185
R10616 GNDA.n4777 GNDA.n4776 185
R10617 GNDA.n4779 GNDA.n4778 185
R10618 GNDA.n4781 GNDA.n4780 185
R10619 GNDA.n4783 GNDA.n4782 185
R10620 GNDA.n4785 GNDA.n4784 185
R10621 GNDA.n4787 GNDA.n4786 185
R10622 GNDA.n4789 GNDA.n4788 185
R10623 GNDA.n1660 GNDA.n1659 185
R10624 GNDA.n1662 GNDA.n1661 185
R10625 GNDA.n1664 GNDA.n1663 185
R10626 GNDA.n1666 GNDA.n1665 185
R10627 GNDA.n1668 GNDA.n1667 185
R10628 GNDA.n1670 GNDA.n1669 185
R10629 GNDA.n1672 GNDA.n1671 185
R10630 GNDA.n1674 GNDA.n1673 185
R10631 GNDA.n1675 GNDA.n1623 185
R10632 GNDA.n1642 GNDA.n1641 185
R10633 GNDA.n1644 GNDA.n1643 185
R10634 GNDA.n1646 GNDA.n1645 185
R10635 GNDA.n1648 GNDA.n1647 185
R10636 GNDA.n1650 GNDA.n1649 185
R10637 GNDA.n1652 GNDA.n1651 185
R10638 GNDA.n1654 GNDA.n1653 185
R10639 GNDA.n1656 GNDA.n1655 185
R10640 GNDA.n1658 GNDA.n1657 185
R10641 GNDA.n1615 GNDA.n1601 185
R10642 GNDA.n1626 GNDA.n1625 185
R10643 GNDA.n1628 GNDA.n1627 185
R10644 GNDA.n1630 GNDA.n1629 185
R10645 GNDA.n1632 GNDA.n1631 185
R10646 GNDA.n1634 GNDA.n1633 185
R10647 GNDA.n1636 GNDA.n1635 185
R10648 GNDA.n1638 GNDA.n1637 185
R10649 GNDA.n1640 GNDA.n1639 185
R10650 GNDA.n1605 GNDA.n1602 185
R10651 GNDA.n1708 GNDA.n1707 185
R10652 GNDA.n1681 GNDA.n1604 185
R10653 GNDA.n1687 GNDA.n1686 185
R10654 GNDA.n1685 GNDA.n1680 185
R10655 GNDA.n1694 GNDA.n1693 185
R10656 GNDA.n1692 GNDA.n1679 185
R10657 GNDA.n1699 GNDA.n1624 185
R10658 GNDA.n1704 GNDA.n1703 185
R10659 GNDA.n4949 GNDA.n4887 185
R10660 GNDA.n4963 GNDA.n4962 185
R10661 GNDA.n4961 GNDA.n4888 185
R10662 GNDA.n4960 GNDA.n4959 185
R10663 GNDA.n4958 GNDA.n4957 185
R10664 GNDA.n4956 GNDA.n4955 185
R10665 GNDA.n4954 GNDA.n4953 185
R10666 GNDA.n4952 GNDA.n4951 185
R10667 GNDA.n4950 GNDA.n4864 185
R10668 GNDA.n4932 GNDA.n4931 185
R10669 GNDA.n4934 GNDA.n4933 185
R10670 GNDA.n4936 GNDA.n4935 185
R10671 GNDA.n4938 GNDA.n4937 185
R10672 GNDA.n4940 GNDA.n4939 185
R10673 GNDA.n4942 GNDA.n4941 185
R10674 GNDA.n4944 GNDA.n4943 185
R10675 GNDA.n4946 GNDA.n4945 185
R10676 GNDA.n4948 GNDA.n4947 185
R10677 GNDA.n4914 GNDA.n4913 185
R10678 GNDA.n4916 GNDA.n4915 185
R10679 GNDA.n4918 GNDA.n4917 185
R10680 GNDA.n4920 GNDA.n4919 185
R10681 GNDA.n4922 GNDA.n4921 185
R10682 GNDA.n4924 GNDA.n4923 185
R10683 GNDA.n4926 GNDA.n4925 185
R10684 GNDA.n4928 GNDA.n4927 185
R10685 GNDA.n4930 GNDA.n4929 185
R10686 GNDA.n4912 GNDA.n4911 185
R10687 GNDA.n4906 GNDA.n4905 185
R10688 GNDA.n4904 GNDA.n4903 185
R10689 GNDA.n4899 GNDA.n4898 185
R10690 GNDA.n4894 GNDA.n4872 185
R10691 GNDA.n4967 GNDA.n4966 185
R10692 GNDA.n4871 GNDA.n4869 185
R10693 GNDA.n4973 GNDA.n4972 185
R10694 GNDA.n4975 GNDA.n4974 185
R10695 GNDA.n3246 GNDA.n3245 185
R10696 GNDA.n3243 GNDA.n3242 185
R10697 GNDA.n2825 GNDA.n2824 185
R10698 GNDA.n2824 GNDA.n2823 185
R10699 GNDA.n2825 GNDA.n2815 185
R10700 GNDA.n2818 GNDA.n2815 185
R10701 GNDA.n5228 GNDA.n80 185
R10702 GNDA.n5242 GNDA.n5241 185
R10703 GNDA.n5240 GNDA.n81 185
R10704 GNDA.n5239 GNDA.n5238 185
R10705 GNDA.n5237 GNDA.n5236 185
R10706 GNDA.n5235 GNDA.n5234 185
R10707 GNDA.n5233 GNDA.n5232 185
R10708 GNDA.n5231 GNDA.n5230 185
R10709 GNDA.n5229 GNDA.n57 185
R10710 GNDA.n5211 GNDA.n5210 185
R10711 GNDA.n5213 GNDA.n5212 185
R10712 GNDA.n5215 GNDA.n5214 185
R10713 GNDA.n5217 GNDA.n5216 185
R10714 GNDA.n5219 GNDA.n5218 185
R10715 GNDA.n5221 GNDA.n5220 185
R10716 GNDA.n5223 GNDA.n5222 185
R10717 GNDA.n5225 GNDA.n5224 185
R10718 GNDA.n5227 GNDA.n5226 185
R10719 GNDA.n5193 GNDA.n5192 185
R10720 GNDA.n5195 GNDA.n5194 185
R10721 GNDA.n5197 GNDA.n5196 185
R10722 GNDA.n5199 GNDA.n5198 185
R10723 GNDA.n5201 GNDA.n5200 185
R10724 GNDA.n5203 GNDA.n5202 185
R10725 GNDA.n5205 GNDA.n5204 185
R10726 GNDA.n5207 GNDA.n5206 185
R10727 GNDA.n5209 GNDA.n5208 185
R10728 GNDA.n5191 GNDA.n5190 185
R10729 GNDA.n5185 GNDA.n5184 185
R10730 GNDA.n5183 GNDA.n5182 185
R10731 GNDA.n5178 GNDA.n5177 185
R10732 GNDA.n5173 GNDA.n65 185
R10733 GNDA.n5246 GNDA.n5245 185
R10734 GNDA.n64 GNDA.n62 185
R10735 GNDA.n5252 GNDA.n5251 185
R10736 GNDA.n5254 GNDA.n5253 185
R10737 GNDA.n4771 GNDA.n4770 185
R10738 GNDA.n4765 GNDA.n4764 185
R10739 GNDA.n4763 GNDA.n4762 185
R10740 GNDA.n4758 GNDA.n4757 185
R10741 GNDA.n4756 GNDA.n4755 185
R10742 GNDA.n4750 GNDA.n4749 185
R10743 GNDA.n4745 GNDA.n4724 185
R10744 GNDA.n4828 GNDA.n4827 185
R10745 GNDA.n4723 GNDA.n4721 185
R10746 GNDA.n2889 GNDA.n2888 185
R10747 GNDA.n2891 GNDA.n2673 185
R10748 GNDA.n2894 GNDA.n2893 185
R10749 GNDA.n2895 GNDA.n2672 185
R10750 GNDA.n2897 GNDA.n2896 185
R10751 GNDA.n2899 GNDA.n2671 185
R10752 GNDA.n2902 GNDA.n2901 185
R10753 GNDA.n2903 GNDA.n2670 185
R10754 GNDA.n2905 GNDA.n2904 185
R10755 GNDA.n2871 GNDA.n2678 185
R10756 GNDA.n2873 GNDA.n2872 185
R10757 GNDA.n2875 GNDA.n2677 185
R10758 GNDA.n2878 GNDA.n2877 185
R10759 GNDA.n2879 GNDA.n2676 185
R10760 GNDA.n2881 GNDA.n2880 185
R10761 GNDA.n2883 GNDA.n2675 185
R10762 GNDA.n2886 GNDA.n2885 185
R10763 GNDA.n2887 GNDA.n2674 185
R10764 GNDA.n2855 GNDA.n2854 185
R10765 GNDA.n2856 GNDA.n2683 185
R10766 GNDA.n2858 GNDA.n2857 185
R10767 GNDA.n2860 GNDA.n2681 185
R10768 GNDA.n2862 GNDA.n2861 185
R10769 GNDA.n2863 GNDA.n2680 185
R10770 GNDA.n2865 GNDA.n2864 185
R10771 GNDA.n2867 GNDA.n2679 185
R10772 GNDA.n2870 GNDA.n2869 185
R10773 GNDA.n2853 GNDA.n2686 185
R10774 GNDA.n2851 GNDA.n2850 185
R10775 GNDA.n2840 GNDA.n2687 185
R10776 GNDA.n2839 GNDA.n2838 185
R10777 GNDA.n2836 GNDA.n2834 185
R10778 GNDA.n2830 GNDA.n2669 185
R10779 GNDA.n2914 GNDA.n2913 185
R10780 GNDA.n2911 GNDA.n2667 185
R10781 GNDA.n2910 GNDA.n2909 185
R10782 GNDA.n5147 GNDA.n5146 185
R10783 GNDA.n5149 GNDA.n5148 185
R10784 GNDA.n5151 GNDA.n5150 185
R10785 GNDA.n5153 GNDA.n5152 185
R10786 GNDA.n5155 GNDA.n5154 185
R10787 GNDA.n5157 GNDA.n5156 185
R10788 GNDA.n5159 GNDA.n5158 185
R10789 GNDA.n5161 GNDA.n5160 185
R10790 GNDA.n5162 GNDA.n20 185
R10791 GNDA.n5129 GNDA.n5128 185
R10792 GNDA.n5131 GNDA.n5130 185
R10793 GNDA.n5133 GNDA.n5132 185
R10794 GNDA.n5135 GNDA.n5134 185
R10795 GNDA.n5137 GNDA.n5136 185
R10796 GNDA.n5139 GNDA.n5138 185
R10797 GNDA.n5141 GNDA.n5140 185
R10798 GNDA.n5143 GNDA.n5142 185
R10799 GNDA.n5145 GNDA.n5144 185
R10800 GNDA.n5111 GNDA.n5110 185
R10801 GNDA.n5113 GNDA.n5112 185
R10802 GNDA.n5115 GNDA.n5114 185
R10803 GNDA.n5117 GNDA.n5116 185
R10804 GNDA.n5119 GNDA.n5118 185
R10805 GNDA.n5121 GNDA.n5120 185
R10806 GNDA.n5123 GNDA.n5122 185
R10807 GNDA.n5125 GNDA.n5124 185
R10808 GNDA.n5127 GNDA.n5126 185
R10809 GNDA.n5109 GNDA.n5108 185
R10810 GNDA.n5103 GNDA.n5102 185
R10811 GNDA.n5098 GNDA.n3 185
R10812 GNDA.n5269 GNDA.n5268 185
R10813 GNDA.n34 GNDA.n2 185
R10814 GNDA.n38 GNDA.n37 185
R10815 GNDA.n36 GNDA.n33 185
R10816 GNDA.n23 GNDA.n21 185
R10817 GNDA.n5265 GNDA.n5264 185
R10818 GNDA.n3194 GNDA.n1542 175.546
R10819 GNDA.n3199 GNDA.n1542 175.546
R10820 GNDA.n3199 GNDA.n1539 175.546
R10821 GNDA.n3203 GNDA.n1539 175.546
R10822 GNDA.n3204 GNDA.n3203 175.546
R10823 GNDA.n3205 GNDA.n3204 175.546
R10824 GNDA.n3205 GNDA.n1537 175.546
R10825 GNDA.n3209 GNDA.n1537 175.546
R10826 GNDA.n3209 GNDA.n1534 175.546
R10827 GNDA.n3216 GNDA.n1534 175.546
R10828 GNDA.n3216 GNDA.n1535 175.546
R10829 GNDA.n3142 GNDA.n3046 175.546
R10830 GNDA.n3117 GNDA.n3046 175.546
R10831 GNDA.n3131 GNDA.n3117 175.546
R10832 GNDA.n3131 GNDA.n3127 175.546
R10833 GNDA.n3127 GNDA.n3118 175.546
R10834 GNDA.n3118 GNDA.n1516 175.546
R10835 GNDA.n3251 GNDA.n1516 175.546
R10836 GNDA.n3251 GNDA.n1508 175.546
R10837 GNDA.n3262 GNDA.n1508 175.546
R10838 GNDA.n3262 GNDA.n1509 175.546
R10839 GNDA.n3220 GNDA.n1509 175.546
R10840 GNDA.n3166 GNDA.n3165 175.546
R10841 GNDA.n3165 GNDA.n3164 175.546
R10842 GNDA.n3161 GNDA.n3160 175.546
R10843 GNDA.n3158 GNDA.n1812 175.546
R10844 GNDA.n3154 GNDA.n3152 175.546
R10845 GNDA.n3150 GNDA.n1820 175.546
R10846 GNDA.n3175 GNDA.n1548 175.546
R10847 GNDA.n3179 GNDA.n3177 175.546
R10848 GNDA.n3183 GNDA.n1546 175.546
R10849 GNDA.n3187 GNDA.n3185 175.546
R10850 GNDA.n3191 GNDA.n1544 175.546
R10851 GNDA.n1807 GNDA.n1804 175.546
R10852 GNDA.n1810 GNDA.n1809 175.546
R10853 GNDA.n1815 GNDA.n1814 175.546
R10854 GNDA.n1818 GNDA.n1817 175.546
R10855 GNDA.n1823 GNDA.n1822 175.546
R10856 GNDA.n3010 GNDA.n2984 175.546
R10857 GNDA.n3006 GNDA.n3005 175.546
R10858 GNDA.n3003 GNDA.n2987 175.546
R10859 GNDA.n2999 GNDA.n2998 175.546
R10860 GNDA.n2996 GNDA.n2990 175.546
R10861 GNDA.n2738 GNDA.n1495 175.546
R10862 GNDA.n3292 GNDA.n1495 175.546
R10863 GNDA.n3292 GNDA.n1496 175.546
R10864 GNDA.n3288 GNDA.n1496 175.546
R10865 GNDA.n3288 GNDA.n1470 175.546
R10866 GNDA.n3301 GNDA.n1470 175.546
R10867 GNDA.n3301 GNDA.n1471 175.546
R10868 GNDA.n2725 GNDA.n1471 175.546
R10869 GNDA.n2725 GNDA.n2721 175.546
R10870 GNDA.n2798 GNDA.n2721 175.546
R10871 GNDA.n2798 GNDA.n1826 175.546
R10872 GNDA.n3022 GNDA.n1847 175.546
R10873 GNDA.n3023 GNDA.n3022 175.546
R10874 GNDA.n3025 GNDA.n1846 175.546
R10875 GNDA.n3034 GNDA.n1838 175.546
R10876 GNDA.n3037 GNDA.n3036 175.546
R10877 GNDA.n3039 GNDA.n1836 175.546
R10878 GNDA.n2955 GNDA.n2954 175.546
R10879 GNDA.n2951 GNDA.n2950 175.546
R10880 GNDA.n2947 GNDA.n2946 175.546
R10881 GNDA.n2943 GNDA.n2942 175.546
R10882 GNDA.n2939 GNDA.n2938 175.546
R10883 GNDA.n2963 GNDA.n2961 175.546
R10884 GNDA.n2967 GNDA.n1853 175.546
R10885 GNDA.n2971 GNDA.n2969 175.546
R10886 GNDA.n2975 GNDA.n1851 175.546
R10887 GNDA.n2979 GNDA.n2977 175.546
R10888 GNDA.n2934 GNDA.n1858 175.546
R10889 GNDA.n2664 GNDA.n1858 175.546
R10890 GNDA.n2916 GNDA.n2664 175.546
R10891 GNDA.n2916 GNDA.n2666 175.546
R10892 GNDA.n2831 GNDA.n2666 175.546
R10893 GNDA.n2831 GNDA.n2829 175.546
R10894 GNDA.n2842 GNDA.n2829 175.546
R10895 GNDA.n2842 GNDA.n2689 175.546
R10896 GNDA.n2848 GNDA.n2689 175.546
R10897 GNDA.n2848 GNDA.n2691 175.546
R10898 GNDA.n2691 GNDA.n1831 175.546
R10899 GNDA.n3020 GNDA.n3018 175.546
R10900 GNDA.n3027 GNDA.n1843 175.546
R10901 GNDA.n3030 GNDA.n3029 175.546
R10902 GNDA.n3032 GNDA.n1841 175.546
R10903 GNDA.n3041 GNDA.n1834 175.546
R10904 GNDA.n373 GNDA.n370 175.546
R10905 GNDA.n376 GNDA.n375 175.546
R10906 GNDA.n381 GNDA.n378 175.546
R10907 GNDA.n384 GNDA.n383 175.546
R10908 GNDA.n388 GNDA.n386 175.546
R10909 GNDA.n4693 GNDA.n350 175.546
R10910 GNDA.n4689 GNDA.n350 175.546
R10911 GNDA.n4689 GNDA.n352 175.546
R10912 GNDA.n4685 GNDA.n352 175.546
R10913 GNDA.n4685 GNDA.n354 175.546
R10914 GNDA.n4676 GNDA.n354 175.546
R10915 GNDA.n4676 GNDA.n4675 175.546
R10916 GNDA.n4675 GNDA.n361 175.546
R10917 GNDA.n4671 GNDA.n361 175.546
R10918 GNDA.n4671 GNDA.n363 175.546
R10919 GNDA.n4667 GNDA.n363 175.546
R10920 GNDA.n347 GNDA.n304 175.546
R10921 GNDA.n343 GNDA.n341 175.546
R10922 GNDA.n339 GNDA.n311 175.546
R10923 GNDA.n335 GNDA.n333 175.546
R10924 GNDA.n331 GNDA.n319 175.546
R10925 GNDA.n1739 GNDA.n1590 175.546
R10926 GNDA.n1735 GNDA.n1590 175.546
R10927 GNDA.n1735 GNDA.n1592 175.546
R10928 GNDA.n1731 GNDA.n1592 175.546
R10929 GNDA.n1731 GNDA.n1729 175.546
R10930 GNDA.n1729 GNDA.n1728 175.546
R10931 GNDA.n1728 GNDA.n1595 175.546
R10932 GNDA.n1724 GNDA.n1595 175.546
R10933 GNDA.n1724 GNDA.n1597 175.546
R10934 GNDA.n1720 GNDA.n1597 175.546
R10935 GNDA.n1720 GNDA.n1600 175.546
R10936 GNDA.n1701 GNDA.n1700 175.546
R10937 GNDA.n1697 GNDA.n1696 175.546
R10938 GNDA.n1690 GNDA.n1689 175.546
R10939 GNDA.n1683 GNDA.n1682 175.546
R10940 GNDA.n1711 GNDA.n1710 175.546
R10941 GNDA.n1766 GNDA.n1561 175.546
R10942 GNDA.n1774 GNDA.n1561 175.546
R10943 GNDA.n1778 GNDA.n1776 175.546
R10944 GNDA.n1786 GNDA.n1557 175.546
R10945 GNDA.n1790 GNDA.n1788 175.546
R10946 GNDA.n1797 GNDA.n1553 175.546
R10947 GNDA.n1760 GNDA.n1759 175.546
R10948 GNDA.n1756 GNDA.n1755 175.546
R10949 GNDA.n1752 GNDA.n1751 175.546
R10950 GNDA.n1748 GNDA.n1747 175.546
R10951 GNDA.n1744 GNDA.n1743 175.546
R10952 GNDA.n1769 GNDA.n1768 175.546
R10953 GNDA.n1772 GNDA.n1771 175.546
R10954 GNDA.n1781 GNDA.n1780 175.546
R10955 GNDA.n1784 GNDA.n1783 175.546
R10956 GNDA.n1793 GNDA.n1792 175.546
R10957 GNDA.n5046 GNDA.n5045 175.546
R10958 GNDA.n219 GNDA.n199 175.546
R10959 GNDA.n201 GNDA.n198 175.546
R10960 GNDA.n209 GNDA.n208 175.546
R10961 GNDA.n4983 GNDA.n188 175.546
R10962 GNDA.n5070 GNDA.n136 175.546
R10963 GNDA.n5066 GNDA.n141 175.546
R10964 GNDA.n5064 GNDA.n5063 175.546
R10965 GNDA.n5060 GNDA.n5059 175.546
R10966 GNDA.n5056 GNDA.n5055 175.546
R10967 GNDA.n1567 GNDA.n1566 175.546
R10968 GNDA.n1571 GNDA.n1570 175.546
R10969 GNDA.n1575 GNDA.n1574 175.546
R10970 GNDA.n1579 GNDA.n1578 175.546
R10971 GNDA.n1583 GNDA.n1582 175.546
R10972 GNDA.n151 GNDA.n142 175.546
R10973 GNDA.n144 GNDA.n143 175.546
R10974 GNDA.n146 GNDA.n145 175.546
R10975 GNDA.n148 GNDA.n147 175.546
R10976 GNDA.n150 GNDA.n149 175.546
R10977 GNDA.n4865 GNDA.n226 175.546
R10978 GNDA.n4970 GNDA.n4969 175.546
R10979 GNDA.n4896 GNDA.n4895 175.546
R10980 GNDA.n4901 GNDA.n4900 175.546
R10981 GNDA.n4909 GNDA.n4908 175.546
R10982 GNDA.n265 GNDA.n264 175.546
R10983 GNDA.n269 GNDA.n268 175.546
R10984 GNDA.n273 GNDA.n272 175.546
R10985 GNDA.n278 GNDA.n240 175.546
R10986 GNDA.n239 GNDA.n229 175.546
R10987 GNDA.n4862 GNDA.n229 175.546
R10988 GNDA.n257 GNDA.n256 175.546
R10989 GNDA.n253 GNDA.n252 175.546
R10990 GNDA.n249 GNDA.n248 175.546
R10991 GNDA.n245 GNDA.n244 175.546
R10992 GNDA.n241 GNDA.n129 175.546
R10993 GNDA.n307 GNDA.n306 175.546
R10994 GNDA.n312 GNDA.n309 175.546
R10995 GNDA.n315 GNDA.n314 175.546
R10996 GNDA.n320 GNDA.n317 175.546
R10997 GNDA.n323 GNDA.n322 175.546
R10998 GNDA.n4831 GNDA.n4830 175.546
R10999 GNDA.n4747 GNDA.n4746 175.546
R11000 GNDA.n4753 GNDA.n4752 175.546
R11001 GNDA.n4760 GNDA.n4759 175.546
R11002 GNDA.n4768 GNDA.n4767 175.546
R11003 GNDA.n288 GNDA.n287 175.546
R11004 GNDA.n4853 GNDA.n287 175.546
R11005 GNDA.n4851 GNDA.n4850 175.546
R11006 GNDA.n4847 GNDA.n4846 175.546
R11007 GNDA.n4843 GNDA.n4842 175.546
R11008 GNDA.n4839 GNDA.n4838 175.546
R11009 GNDA.n4717 GNDA.n289 175.546
R11010 GNDA.n4717 GNDA.n291 175.546
R11011 GNDA.n4713 GNDA.n291 175.546
R11012 GNDA.n4713 GNDA.n293 175.546
R11013 GNDA.n4709 GNDA.n293 175.546
R11014 GNDA.n4709 GNDA.n295 175.546
R11015 GNDA.n4705 GNDA.n295 175.546
R11016 GNDA.n4705 GNDA.n297 175.546
R11017 GNDA.n4701 GNDA.n297 175.546
R11018 GNDA.n4701 GNDA.n299 175.546
R11019 GNDA.n4697 GNDA.n299 175.546
R11020 GNDA.n58 GNDA.n54 175.546
R11021 GNDA.n5249 GNDA.n5248 175.546
R11022 GNDA.n5175 GNDA.n5174 175.546
R11023 GNDA.n5180 GNDA.n5179 175.546
R11024 GNDA.n5188 GNDA.n5187 175.546
R11025 GNDA.n409 GNDA.n408 175.546
R11026 GNDA.n406 GNDA.n372 175.546
R11027 GNDA.n402 GNDA.n400 175.546
R11028 GNDA.n398 GNDA.n380 175.546
R11029 GNDA.n394 GNDA.n392 175.546
R11030 GNDA.n4663 GNDA.n413 175.546
R11031 GNDA.n4659 GNDA.n413 175.546
R11032 GNDA.n4659 GNDA.n415 175.546
R11033 GNDA.n4655 GNDA.n415 175.546
R11034 GNDA.n4655 GNDA.n417 175.546
R11035 GNDA.n4651 GNDA.n417 175.546
R11036 GNDA.n4651 GNDA.n419 175.546
R11037 GNDA.n4647 GNDA.n419 175.546
R11038 GNDA.n4647 GNDA.n421 175.546
R11039 GNDA.n4643 GNDA.n421 175.546
R11040 GNDA.n4643 GNDA.n423 175.546
R11041 GNDA.n5262 GNDA.n24 175.546
R11042 GNDA.n40 GNDA.n25 175.546
R11043 GNDA.n31 GNDA.n30 175.546
R11044 GNDA.n5100 GNDA.n5099 175.546
R11045 GNDA.n5106 GNDA.n5105 175.546
R11046 GNDA.n4639 GNDA.n425 175.546
R11047 GNDA.n4635 GNDA.n425 175.546
R11048 GNDA.n4635 GNDA.n427 175.546
R11049 GNDA.n4631 GNDA.n427 175.546
R11050 GNDA.n4631 GNDA.n4628 175.546
R11051 GNDA.n4628 GNDA.n93 175.546
R11052 GNDA.n5083 GNDA.n93 175.546
R11053 GNDA.n5083 GNDA.n91 175.546
R11054 GNDA.n5088 GNDA.n91 175.546
R11055 GNDA.n5088 GNDA.n89 175.546
R11056 GNDA.n5092 GNDA.n89 175.546
R11057 GNDA.n157 GNDA.n100 173.881
R11058 GNDA.t62 GNDA.n101 172.876
R11059 GNDA.t62 GNDA.n111 172.615
R11060 GNDA.n5072 GNDA.n100 171.624
R11061 GNDA.n3259 GNDA.n1512 163.333
R11062 GNDA.n2793 GNDA.n2792 163.333
R11063 GNDA.n4987 GNDA.n4986 163.333
R11064 GNDA.n4772 GNDA.n4771 163.333
R11065 GNDA.n1615 GNDA.n1605 163.333
R11066 GNDA.n4913 GNDA.n4912 163.333
R11067 GNDA.n5192 GNDA.n5191 163.333
R11068 GNDA.n2854 GNDA.n2853 163.333
R11069 GNDA.n5110 GNDA.n5109 163.333
R11070 GNDA.n3580 GNDA.n3579 161.3
R11071 GNDA.n3576 GNDA.n3575 161.3
R11072 GNDA.n4681 GNDA.n355 157.601
R11073 GNDA.t194 GNDA.n1466 154.323
R11074 GNDA.n3094 GNDA.n3054 150
R11075 GNDA.n3090 GNDA.n3088 150
R11076 GNDA.n3086 GNDA.n3056 150
R11077 GNDA.n3082 GNDA.n3080 150
R11078 GNDA.n3078 GNDA.n3058 150
R11079 GNDA.n3074 GNDA.n3073 150
R11080 GNDA.n3071 GNDA.n3061 150
R11081 GNDA.n3067 GNDA.n3066 150
R11082 GNDA.n3135 GNDA.n3134 150
R11083 GNDA.n3124 GNDA.n3122 150
R11084 GNDA.n3254 GNDA.n1515 150
R11085 GNDA.n3257 GNDA.n3256 150
R11086 GNDA.n3102 GNDA.n3052 150
R11087 GNDA.n3106 GNDA.n3104 150
R11088 GNDA.n3110 GNDA.n3050 150
R11089 GNDA.n3113 GNDA.n3112 150
R11090 GNDA.n2762 GNDA.n2761 150
R11091 GNDA.n2766 GNDA.n2765 150
R11092 GNDA.n2770 GNDA.n2769 150
R11093 GNDA.n2774 GNDA.n2773 150
R11094 GNDA.n2778 GNDA.n2777 150
R11095 GNDA.n2782 GNDA.n2781 150
R11096 GNDA.n2786 GNDA.n2785 150
R11097 GNDA.n2790 GNDA.n2789 150
R11098 GNDA.n3295 GNDA.n1492 150
R11099 GNDA.n3285 GNDA.n3284 150
R11100 GNDA.n3298 GNDA.n1473 150
R11101 GNDA.n2727 GNDA.n1474 150
R11102 GNDA.n2754 GNDA.n2753 150
R11103 GNDA.n2750 GNDA.n2749 150
R11104 GNDA.n2746 GNDA.n2745 150
R11105 GNDA.n2742 GNDA.n1491 150
R11106 GNDA.n5019 GNDA.n5018 150
R11107 GNDA.n5015 GNDA.n5014 150
R11108 GNDA.n5011 GNDA.n5010 150
R11109 GNDA.n5007 GNDA.n5006 150
R11110 GNDA.n5003 GNDA.n5002 150
R11111 GNDA.n4999 GNDA.n4998 150
R11112 GNDA.n4995 GNDA.n4994 150
R11113 GNDA.n4991 GNDA.n4990 150
R11114 GNDA.n5042 GNDA.n168 150
R11115 GNDA.n216 GNDA.n169 150
R11116 GNDA.n213 GNDA.n212 150
R11117 GNDA.n205 GNDA.n204 150
R11118 GNDA.n5027 GNDA.n5026 150
R11119 GNDA.n5031 GNDA.n5030 150
R11120 GNDA.n5035 GNDA.n5034 150
R11121 GNDA.n5039 GNDA.n5038 150
R11122 GNDA.n4804 GNDA.n4803 150
R11123 GNDA.n4800 GNDA.n4799 150
R11124 GNDA.n4796 GNDA.n4795 150
R11125 GNDA.n4792 GNDA.n4791 150
R11126 GNDA.n4788 GNDA.n4787 150
R11127 GNDA.n4784 GNDA.n4783 150
R11128 GNDA.n4780 GNDA.n4779 150
R11129 GNDA.n4776 GNDA.n4775 150
R11130 GNDA.n4827 GNDA.n4723 150
R11131 GNDA.n4749 GNDA.n4724 150
R11132 GNDA.n4757 GNDA.n4756 150
R11133 GNDA.n4764 GNDA.n4763 150
R11134 GNDA.n4812 GNDA.n4811 150
R11135 GNDA.n4816 GNDA.n4815 150
R11136 GNDA.n4820 GNDA.n4819 150
R11137 GNDA.n4824 GNDA.n4823 150
R11138 GNDA.n1655 GNDA.n1654 150
R11139 GNDA.n1651 GNDA.n1650 150
R11140 GNDA.n1647 GNDA.n1646 150
R11141 GNDA.n1643 GNDA.n1642 150
R11142 GNDA.n1639 GNDA.n1638 150
R11143 GNDA.n1635 GNDA.n1634 150
R11144 GNDA.n1631 GNDA.n1630 150
R11145 GNDA.n1627 GNDA.n1626 150
R11146 GNDA.n1704 GNDA.n1624 150
R11147 GNDA.n1693 GNDA.n1692 150
R11148 GNDA.n1686 GNDA.n1685 150
R11149 GNDA.n1707 GNDA.n1604 150
R11150 GNDA.n1663 GNDA.n1662 150
R11151 GNDA.n1667 GNDA.n1666 150
R11152 GNDA.n1671 GNDA.n1670 150
R11153 GNDA.n1673 GNDA.n1623 150
R11154 GNDA.n4945 GNDA.n4944 150
R11155 GNDA.n4941 GNDA.n4940 150
R11156 GNDA.n4937 GNDA.n4936 150
R11157 GNDA.n4933 GNDA.n4932 150
R11158 GNDA.n4929 GNDA.n4928 150
R11159 GNDA.n4925 GNDA.n4924 150
R11160 GNDA.n4921 GNDA.n4920 150
R11161 GNDA.n4917 GNDA.n4916 150
R11162 GNDA.n4974 GNDA.n4973 150
R11163 GNDA.n4966 GNDA.n4871 150
R11164 GNDA.n4898 GNDA.n4872 150
R11165 GNDA.n4905 GNDA.n4904 150
R11166 GNDA.n4963 GNDA.n4888 150
R11167 GNDA.n4959 GNDA.n4958 150
R11168 GNDA.n4955 GNDA.n4954 150
R11169 GNDA.n4951 GNDA.n4950 150
R11170 GNDA.n5224 GNDA.n5223 150
R11171 GNDA.n5220 GNDA.n5219 150
R11172 GNDA.n5216 GNDA.n5215 150
R11173 GNDA.n5212 GNDA.n5211 150
R11174 GNDA.n5208 GNDA.n5207 150
R11175 GNDA.n5204 GNDA.n5203 150
R11176 GNDA.n5200 GNDA.n5199 150
R11177 GNDA.n5196 GNDA.n5195 150
R11178 GNDA.n5253 GNDA.n5252 150
R11179 GNDA.n5245 GNDA.n64 150
R11180 GNDA.n5177 GNDA.n65 150
R11181 GNDA.n5184 GNDA.n5183 150
R11182 GNDA.n5242 GNDA.n81 150
R11183 GNDA.n5238 GNDA.n5237 150
R11184 GNDA.n5234 GNDA.n5233 150
R11185 GNDA.n5230 GNDA.n5229 150
R11186 GNDA.n2885 GNDA.n2883 150
R11187 GNDA.n2881 GNDA.n2676 150
R11188 GNDA.n2877 GNDA.n2875 150
R11189 GNDA.n2873 GNDA.n2678 150
R11190 GNDA.n2869 GNDA.n2867 150
R11191 GNDA.n2865 GNDA.n2680 150
R11192 GNDA.n2861 GNDA.n2860 150
R11193 GNDA.n2858 GNDA.n2683 150
R11194 GNDA.n2911 GNDA.n2910 150
R11195 GNDA.n2913 GNDA.n2669 150
R11196 GNDA.n2838 GNDA.n2836 150
R11197 GNDA.n2851 GNDA.n2687 150
R11198 GNDA.n2893 GNDA.n2891 150
R11199 GNDA.n2897 GNDA.n2672 150
R11200 GNDA.n2901 GNDA.n2899 150
R11201 GNDA.n2905 GNDA.n2670 150
R11202 GNDA.n5142 GNDA.n5141 150
R11203 GNDA.n5138 GNDA.n5137 150
R11204 GNDA.n5134 GNDA.n5133 150
R11205 GNDA.n5130 GNDA.n5129 150
R11206 GNDA.n5126 GNDA.n5125 150
R11207 GNDA.n5122 GNDA.n5121 150
R11208 GNDA.n5118 GNDA.n5117 150
R11209 GNDA.n5114 GNDA.n5113 150
R11210 GNDA.n5265 GNDA.n21 150
R11211 GNDA.n37 GNDA.n36 150
R11212 GNDA.n5268 GNDA.n2 150
R11213 GNDA.n5102 GNDA.n3 150
R11214 GNDA.n5150 GNDA.n5149 150
R11215 GNDA.n5154 GNDA.n5153 150
R11216 GNDA.n5158 GNDA.n5157 150
R11217 GNDA.n5160 GNDA.n20 150
R11218 GNDA.n4614 GNDA.n4613 148.017
R11219 GNDA.n746 GNDA.n745 148.017
R11220 GNDA.n742 GNDA.n741 148.017
R11221 GNDA.n4620 GNDA.n4619 148.017
R11222 GNDA.n4613 GNDA.t207 139.571
R11223 GNDA.n3267 GNDA.n1505 136.145
R11224 GNDA.n3268 GNDA.n1504 136.145
R11225 GNDA.n3269 GNDA.n1503 136.145
R11226 GNDA.n3272 GNDA.n1500 136.145
R11227 GNDA.n3273 GNDA.n1499 136.145
R11228 GNDA.n2924 GNDA.n2923 136.145
R11229 GNDA.n2925 GNDA.n2922 136.145
R11230 GNDA.n2926 GNDA.n2921 136.145
R11231 GNDA.n2663 GNDA.n2662 136.145
R11232 GNDA.n2661 GNDA.n2660 136.145
R11233 GNDA.n2824 GNDA.n2817 134.268
R11234 GNDA.n2817 GNDA.n2815 134.268
R11235 GNDA.n1856 GNDA.n281 132.721
R11236 GNDA.n3265 GNDA.t157 130.001
R11237 GNDA.n1828 GNDA.t93 130.001
R11238 GNDA.n2800 GNDA.t60 130.001
R11239 GNDA.n3276 GNDA.t99 130.001
R11240 GNDA.n2735 GNDA.t72 130.001
R11241 GNDA.n2919 GNDA.t160 130.001
R11242 GNDA.n2930 GNDA.t110 130.001
R11243 GNDA.n2657 GNDA.t66 130
R11244 GNDA.n5081 GNDA.t62 127.219
R11245 GNDA.t62 GNDA.n108 127.219
R11246 GNDA.t62 GNDA.n1518 127.219
R11247 GNDA.n3143 GNDA.n1820 124.832
R11248 GNDA.n3147 GNDA.n3146 124.832
R11249 GNDA.n2733 GNDA.n1836 124.832
R11250 GNDA.n3044 GNDA.n3043 124.832
R11251 GNDA.n5168 GNDA.n83 124.832
R11252 GNDA.n327 GNDA.n55 124.832
R11253 GNDA.n1798 GNDA.n1797 124.832
R11254 GNDA.n1795 GNDA.n1551 124.832
R11255 GNDA.n5052 GNDA.n5051 124.832
R11256 GNDA.n4889 GNDA.n159 124.832
R11257 GNDA.n325 GNDA.n85 124.832
R11258 GNDA.n5166 GNDA.n86 124.832
R11259 GNDA.n453 GNDA.n451 121.251
R11260 GNDA.n461 GNDA.n460 121.136
R11261 GNDA.n459 GNDA.n458 121.136
R11262 GNDA.n457 GNDA.n456 121.136
R11263 GNDA.n455 GNDA.n454 121.136
R11264 GNDA.n453 GNDA.n452 121.136
R11265 GNDA.n3557 GNDA.n3556 121.136
R11266 GNDA.n3555 GNDA.n3554 121.136
R11267 GNDA.n3553 GNDA.n3552 121.136
R11268 GNDA.n3551 GNDA.n3550 121.136
R11269 GNDA.n3549 GNDA.n3548 121.136
R11270 GNDA.n3547 GNDA.n3546 121.136
R11271 GNDA.n2628 GNDA.t180 111.799
R11272 GNDA.n2627 GNDA.t14 111.331
R11273 GNDA.n4698 GNDA.n300 105.719
R11274 GNDA.n4666 GNDA.n4665 105.719
R11275 GNDA.n4692 GNDA.n300 103.457
R11276 GNDA.n4665 GNDA.n4664 103.457
R11277 GNDA.n3238 GNDA.n1521 101.718
R11278 GNDA.n2820 GNDA.n2692 101.718
R11279 GNDA.n2826 GNDA.n2694 101.718
R11280 GNDA.n3247 GNDA.n1523 101.718
R11281 GNDA.t62 GNDA.n104 47.6748
R11282 GNDA.n3245 GNDA.n3237 91.069
R11283 GNDA.n3245 GNDA.n3244 91.069
R11284 GNDA.n3242 GNDA.n3235 91.069
R11285 GNDA.n3242 GNDA.n3241 91.069
R11286 GNDA.n2824 GNDA.n2819 91.069
R11287 GNDA.n2822 GNDA.n2815 91.069
R11288 GNDA.n2933 GNDA.n2932 90.1439
R11289 GNDA.n2844 GNDA.n2843 90.1439
R11290 GNDA.n3291 GNDA.n3278 90.1439
R11291 GNDA.n2799 GNDA.n2720 90.1439
R11292 GNDA.n3130 GNDA.n3129 90.1439
R11293 GNDA.n3263 GNDA.n1507 90.1439
R11294 GNDA.n3221 GNDA.n1507 90.1439
R11295 GNDA.n2918 GNDA.n1859 87.1391
R11296 GNDA.t62 GNDA.n1830 87.1391
R11297 GNDA.n3250 GNDA.t281 87.1391
R11298 GNDA.n3145 GNDA.t62 86.1375
R11299 GNDA.n2708 GNDA.n2707 84.306
R11300 GNDA.n2804 GNDA.n2719 84.306
R11301 GNDA.n2665 GNDA.t255 83.1328
R11302 GNDA.n3264 GNDA.n3263 83.1328
R11303 GNDA.n2828 GNDA.t168 82.1312
R11304 GNDA.n3289 GNDA.t197 82.1312
R11305 GNDA.t46 GNDA.n3128 82.1312
R11306 GNDA.n3222 GNDA.t264 78.5658
R11307 GNDA.n2847 GNDA.t215 78.1248
R11308 GNDA.n2723 GNDA.t235 78.1248
R11309 GNDA.t247 GNDA.n1520 78.1248
R11310 GNDA.t62 GNDA.n100 76.3879
R11311 GNDA.n3169 GNDA.n1801 76.3222
R11312 GNDA.n3164 GNDA.n1806 76.3222
R11313 GNDA.n3160 GNDA.n3159 76.3222
R11314 GNDA.n3153 GNDA.n1812 76.3222
R11315 GNDA.n3152 GNDA.n3151 76.3222
R11316 GNDA.n3170 GNDA.n1548 76.3222
R11317 GNDA.n3177 GNDA.n3176 76.3222
R11318 GNDA.n3178 GNDA.n1546 76.3222
R11319 GNDA.n3185 GNDA.n3184 76.3222
R11320 GNDA.n3186 GNDA.n1544 76.3222
R11321 GNDA.n3193 GNDA.n3192 76.3222
R11322 GNDA.n1804 GNDA.n1803 76.3222
R11323 GNDA.n1809 GNDA.n1808 76.3222
R11324 GNDA.n1814 GNDA.n1813 76.3222
R11325 GNDA.n1817 GNDA.n1816 76.3222
R11326 GNDA.n1822 GNDA.n1821 76.3222
R11327 GNDA.n3147 GNDA.n1825 76.3222
R11328 GNDA.n3011 GNDA.n3010 76.3222
R11329 GNDA.n3006 GNDA.n2986 76.3222
R11330 GNDA.n3004 GNDA.n3003 76.3222
R11331 GNDA.n2999 GNDA.n2989 76.3222
R11332 GNDA.n2997 GNDA.n2996 76.3222
R11333 GNDA.n2992 GNDA.n2991 76.3222
R11334 GNDA.n3014 GNDA.n3013 76.3222
R11335 GNDA.n3024 GNDA.n3023 76.3222
R11336 GNDA.n1846 GNDA.n1845 76.3222
R11337 GNDA.n3035 GNDA.n3034 76.3222
R11338 GNDA.n3038 GNDA.n3037 76.3222
R11339 GNDA.n1855 GNDA.n286 76.3222
R11340 GNDA.n2954 GNDA.n285 76.3222
R11341 GNDA.n2950 GNDA.n284 76.3222
R11342 GNDA.n2946 GNDA.n283 76.3222
R11343 GNDA.n2942 GNDA.n282 76.3222
R11344 GNDA.n2938 GNDA.n281 76.3222
R11345 GNDA.n2961 GNDA.n2960 76.3222
R11346 GNDA.n2962 GNDA.n1853 76.3222
R11347 GNDA.n2969 GNDA.n2968 76.3222
R11348 GNDA.n2970 GNDA.n1851 76.3222
R11349 GNDA.n2977 GNDA.n2976 76.3222
R11350 GNDA.n2978 GNDA.n1849 76.3222
R11351 GNDA.n3017 GNDA.n3016 76.3222
R11352 GNDA.n3020 GNDA.n3019 76.3222
R11353 GNDA.n3028 GNDA.n3027 76.3222
R11354 GNDA.n3031 GNDA.n3030 76.3222
R11355 GNDA.n1841 GNDA.n1840 76.3222
R11356 GNDA.n3042 GNDA.n3041 76.3222
R11357 GNDA.n370 GNDA.n369 76.3222
R11358 GNDA.n375 GNDA.n374 76.3222
R11359 GNDA.n378 GNDA.n377 76.3222
R11360 GNDA.n383 GNDA.n382 76.3222
R11361 GNDA.n386 GNDA.n385 76.3222
R11362 GNDA.n387 GNDA.n83 76.3222
R11363 GNDA.n349 GNDA.n348 76.3222
R11364 GNDA.n342 GNDA.n304 76.3222
R11365 GNDA.n341 GNDA.n340 76.3222
R11366 GNDA.n334 GNDA.n311 76.3222
R11367 GNDA.n333 GNDA.n332 76.3222
R11368 GNDA.n326 GNDA.n319 76.3222
R11369 GNDA.n1552 GNDA.n195 76.3222
R11370 GNDA.n1701 GNDA.n194 76.3222
R11371 GNDA.n1696 GNDA.n193 76.3222
R11372 GNDA.n1689 GNDA.n192 76.3222
R11373 GNDA.n1682 GNDA.n191 76.3222
R11374 GNDA.n1711 GNDA.n190 76.3222
R11375 GNDA.n1765 GNDA.n1764 76.3222
R11376 GNDA.n1775 GNDA.n1774 76.3222
R11377 GNDA.n1778 GNDA.n1777 76.3222
R11378 GNDA.n1787 GNDA.n1786 76.3222
R11379 GNDA.n1790 GNDA.n1789 76.3222
R11380 GNDA.n1760 GNDA.n112 76.3222
R11381 GNDA.n1756 GNDA.n113 76.3222
R11382 GNDA.n1752 GNDA.n114 76.3222
R11383 GNDA.n1748 GNDA.n115 76.3222
R11384 GNDA.n1744 GNDA.n116 76.3222
R11385 GNDA.n1740 GNDA.n117 76.3222
R11386 GNDA.n1768 GNDA.n1563 76.3222
R11387 GNDA.n1772 GNDA.n1770 76.3222
R11388 GNDA.n1780 GNDA.n1559 76.3222
R11389 GNDA.n1784 GNDA.n1782 76.3222
R11390 GNDA.n1792 GNDA.n1555 76.3222
R11391 GNDA.n1795 GNDA.n1794 76.3222
R11392 GNDA.n5050 GNDA.n163 76.3222
R11393 GNDA.n5045 GNDA.n166 76.3222
R11394 GNDA.n220 GNDA.n219 76.3222
R11395 GNDA.n201 GNDA.n197 76.3222
R11396 GNDA.n208 GNDA.n196 76.3222
R11397 GNDA.n4983 GNDA.n4982 76.3222
R11398 GNDA.n5074 GNDA.n5073 76.3222
R11399 GNDA.n5071 GNDA.n5070 76.3222
R11400 GNDA.n5066 GNDA.n140 76.3222
R11401 GNDA.n5063 GNDA.n139 76.3222
R11402 GNDA.n5059 GNDA.n138 76.3222
R11403 GNDA.n5055 GNDA.n137 76.3222
R11404 GNDA.n1566 GNDA.n118 76.3222
R11405 GNDA.n1570 GNDA.n119 76.3222
R11406 GNDA.n1574 GNDA.n120 76.3222
R11407 GNDA.n1578 GNDA.n121 76.3222
R11408 GNDA.n1582 GNDA.n122 76.3222
R11409 GNDA.n1586 GNDA.n123 76.3222
R11410 GNDA.n152 GNDA.n151 76.3222
R11411 GNDA.n153 GNDA.n143 76.3222
R11412 GNDA.n154 GNDA.n145 76.3222
R11413 GNDA.n155 GNDA.n147 76.3222
R11414 GNDA.n156 GNDA.n149 76.3222
R11415 GNDA.n159 GNDA.n158 76.3222
R11416 GNDA.n4980 GNDA.n4979 76.3222
R11417 GNDA.n4865 GNDA.n225 76.3222
R11418 GNDA.n4969 GNDA.n224 76.3222
R11419 GNDA.n4896 GNDA.n223 76.3222
R11420 GNDA.n4900 GNDA.n222 76.3222
R11421 GNDA.n4909 GNDA.n221 76.3222
R11422 GNDA.n261 GNDA.n235 76.3222
R11423 GNDA.n265 GNDA.n236 76.3222
R11424 GNDA.n269 GNDA.n237 76.3222
R11425 GNDA.n273 GNDA.n238 76.3222
R11426 GNDA.n279 GNDA.n278 76.3222
R11427 GNDA.n257 GNDA.n124 76.3222
R11428 GNDA.n253 GNDA.n125 76.3222
R11429 GNDA.n249 GNDA.n126 76.3222
R11430 GNDA.n245 GNDA.n127 76.3222
R11431 GNDA.n241 GNDA.n128 76.3222
R11432 GNDA.n5079 GNDA.n5078 76.3222
R11433 GNDA.n306 GNDA.n305 76.3222
R11434 GNDA.n309 GNDA.n308 76.3222
R11435 GNDA.n314 GNDA.n313 76.3222
R11436 GNDA.n317 GNDA.n316 76.3222
R11437 GNDA.n322 GNDA.n321 76.3222
R11438 GNDA.n325 GNDA.n324 76.3222
R11439 GNDA.n4831 GNDA.n48 76.3222
R11440 GNDA.n4746 GNDA.n47 76.3222
R11441 GNDA.n4752 GNDA.n46 76.3222
R11442 GNDA.n4760 GNDA.n45 76.3222
R11443 GNDA.n4767 GNDA.n44 76.3222
R11444 GNDA.n4741 GNDA.n43 76.3222
R11445 GNDA.n4859 GNDA.n4858 76.3222
R11446 GNDA.n4853 GNDA.n230 76.3222
R11447 GNDA.n4850 GNDA.n231 76.3222
R11448 GNDA.n4846 GNDA.n232 76.3222
R11449 GNDA.n4842 GNDA.n233 76.3222
R11450 GNDA.n5079 GNDA.n129 76.3222
R11451 GNDA.n244 GNDA.n128 76.3222
R11452 GNDA.n248 GNDA.n127 76.3222
R11453 GNDA.n252 GNDA.n126 76.3222
R11454 GNDA.n256 GNDA.n125 76.3222
R11455 GNDA.n260 GNDA.n124 76.3222
R11456 GNDA.n1583 GNDA.n123 76.3222
R11457 GNDA.n1579 GNDA.n122 76.3222
R11458 GNDA.n1575 GNDA.n121 76.3222
R11459 GNDA.n1571 GNDA.n120 76.3222
R11460 GNDA.n1567 GNDA.n119 76.3222
R11461 GNDA.n135 GNDA.n118 76.3222
R11462 GNDA.n1743 GNDA.n117 76.3222
R11463 GNDA.n1747 GNDA.n116 76.3222
R11464 GNDA.n1751 GNDA.n115 76.3222
R11465 GNDA.n1755 GNDA.n114 76.3222
R11466 GNDA.n1759 GNDA.n113 76.3222
R11467 GNDA.n1763 GNDA.n112 76.3222
R11468 GNDA.n5259 GNDA.n54 76.3222
R11469 GNDA.n5249 GNDA.n53 76.3222
R11470 GNDA.n5174 GNDA.n52 76.3222
R11471 GNDA.n5180 GNDA.n51 76.3222
R11472 GNDA.n5187 GNDA.n50 76.3222
R11473 GNDA.n5169 GNDA.n49 76.3222
R11474 GNDA.n5259 GNDA.n5258 76.3222
R11475 GNDA.n58 GNDA.n53 76.3222
R11476 GNDA.n5248 GNDA.n52 76.3222
R11477 GNDA.n5175 GNDA.n51 76.3222
R11478 GNDA.n5179 GNDA.n50 76.3222
R11479 GNDA.n5188 GNDA.n49 76.3222
R11480 GNDA.n4835 GNDA.n48 76.3222
R11481 GNDA.n4830 GNDA.n47 76.3222
R11482 GNDA.n4747 GNDA.n46 76.3222
R11483 GNDA.n4753 GNDA.n45 76.3222
R11484 GNDA.n4759 GNDA.n44 76.3222
R11485 GNDA.n4768 GNDA.n43 76.3222
R11486 GNDA.n324 GNDA.n323 76.3222
R11487 GNDA.n321 GNDA.n320 76.3222
R11488 GNDA.n316 GNDA.n315 76.3222
R11489 GNDA.n313 GNDA.n312 76.3222
R11490 GNDA.n308 GNDA.n307 76.3222
R11491 GNDA.n305 GNDA.n301 76.3222
R11492 GNDA.n348 GNDA.n347 76.3222
R11493 GNDA.n343 GNDA.n342 76.3222
R11494 GNDA.n340 GNDA.n339 76.3222
R11495 GNDA.n335 GNDA.n334 76.3222
R11496 GNDA.n332 GNDA.n331 76.3222
R11497 GNDA.n327 GNDA.n326 76.3222
R11498 GNDA.n158 GNDA.n150 76.3222
R11499 GNDA.n156 GNDA.n148 76.3222
R11500 GNDA.n155 GNDA.n146 76.3222
R11501 GNDA.n154 GNDA.n144 76.3222
R11502 GNDA.n153 GNDA.n142 76.3222
R11503 GNDA.n152 GNDA.n130 76.3222
R11504 GNDA.n5073 GNDA.n136 76.3222
R11505 GNDA.n5071 GNDA.n141 76.3222
R11506 GNDA.n5064 GNDA.n140 76.3222
R11507 GNDA.n5060 GNDA.n139 76.3222
R11508 GNDA.n5056 GNDA.n138 76.3222
R11509 GNDA.n5052 GNDA.n137 76.3222
R11510 GNDA.n3043 GNDA.n3042 76.3222
R11511 GNDA.n1840 GNDA.n1834 76.3222
R11512 GNDA.n3032 GNDA.n3031 76.3222
R11513 GNDA.n3029 GNDA.n3028 76.3222
R11514 GNDA.n3019 GNDA.n1843 76.3222
R11515 GNDA.n3018 GNDA.n3017 76.3222
R11516 GNDA.n3013 GNDA.n1847 76.3222
R11517 GNDA.n3025 GNDA.n3024 76.3222
R11518 GNDA.n1845 GNDA.n1838 76.3222
R11519 GNDA.n3036 GNDA.n3035 76.3222
R11520 GNDA.n3039 GNDA.n3038 76.3222
R11521 GNDA.n2979 GNDA.n2978 76.3222
R11522 GNDA.n2976 GNDA.n2975 76.3222
R11523 GNDA.n2971 GNDA.n2970 76.3222
R11524 GNDA.n2968 GNDA.n2967 76.3222
R11525 GNDA.n2963 GNDA.n2962 76.3222
R11526 GNDA.n2960 GNDA.n2959 76.3222
R11527 GNDA.n2991 GNDA.n2990 76.3222
R11528 GNDA.n2998 GNDA.n2997 76.3222
R11529 GNDA.n2989 GNDA.n2987 76.3222
R11530 GNDA.n3005 GNDA.n3004 76.3222
R11531 GNDA.n2986 GNDA.n2984 76.3222
R11532 GNDA.n3012 GNDA.n3011 76.3222
R11533 GNDA.n3192 GNDA.n3191 76.3222
R11534 GNDA.n3187 GNDA.n3186 76.3222
R11535 GNDA.n3184 GNDA.n3183 76.3222
R11536 GNDA.n3179 GNDA.n3178 76.3222
R11537 GNDA.n3176 GNDA.n3175 76.3222
R11538 GNDA.n3171 GNDA.n3170 76.3222
R11539 GNDA.n4980 GNDA.n226 76.3222
R11540 GNDA.n4970 GNDA.n225 76.3222
R11541 GNDA.n4895 GNDA.n224 76.3222
R11542 GNDA.n4901 GNDA.n223 76.3222
R11543 GNDA.n4908 GNDA.n222 76.3222
R11544 GNDA.n4890 GNDA.n221 76.3222
R11545 GNDA.n5046 GNDA.n163 76.3222
R11546 GNDA.n199 GNDA.n166 76.3222
R11547 GNDA.n220 GNDA.n198 76.3222
R11548 GNDA.n209 GNDA.n197 76.3222
R11549 GNDA.n196 GNDA.n188 76.3222
R11550 GNDA.n4982 GNDA.n189 76.3222
R11551 GNDA.n1700 GNDA.n195 76.3222
R11552 GNDA.n1697 GNDA.n194 76.3222
R11553 GNDA.n1690 GNDA.n193 76.3222
R11554 GNDA.n1683 GNDA.n192 76.3222
R11555 GNDA.n1710 GNDA.n191 76.3222
R11556 GNDA.n1715 GNDA.n190 76.3222
R11557 GNDA.n412 GNDA.n368 76.3222
R11558 GNDA.n408 GNDA.n407 76.3222
R11559 GNDA.n401 GNDA.n372 76.3222
R11560 GNDA.n400 GNDA.n399 76.3222
R11561 GNDA.n393 GNDA.n380 76.3222
R11562 GNDA.n392 GNDA.n391 76.3222
R11563 GNDA.n42 GNDA.n24 76.3222
R11564 GNDA.n5261 GNDA.n25 76.3222
R11565 GNDA.n41 GNDA.n31 76.3222
R11566 GNDA.n5099 GNDA.n29 76.3222
R11567 GNDA.n5105 GNDA.n28 76.3222
R11568 GNDA.n5095 GNDA.n27 76.3222
R11569 GNDA.n5165 GNDA.n42 76.3222
R11570 GNDA.n5262 GNDA.n5261 76.3222
R11571 GNDA.n41 GNDA.n40 76.3222
R11572 GNDA.n30 GNDA.n29 76.3222
R11573 GNDA.n5100 GNDA.n28 76.3222
R11574 GNDA.n5106 GNDA.n27 76.3222
R11575 GNDA.n388 GNDA.n387 76.3222
R11576 GNDA.n385 GNDA.n384 76.3222
R11577 GNDA.n382 GNDA.n381 76.3222
R11578 GNDA.n377 GNDA.n376 76.3222
R11579 GNDA.n374 GNDA.n373 76.3222
R11580 GNDA.n369 GNDA.n366 76.3222
R11581 GNDA.n409 GNDA.n368 76.3222
R11582 GNDA.n407 GNDA.n406 76.3222
R11583 GNDA.n402 GNDA.n401 76.3222
R11584 GNDA.n399 GNDA.n398 76.3222
R11585 GNDA.n394 GNDA.n393 76.3222
R11586 GNDA.n391 GNDA.n86 76.3222
R11587 GNDA.n1794 GNDA.n1793 76.3222
R11588 GNDA.n1783 GNDA.n1555 76.3222
R11589 GNDA.n1782 GNDA.n1781 76.3222
R11590 GNDA.n1771 GNDA.n1559 76.3222
R11591 GNDA.n1770 GNDA.n1769 76.3222
R11592 GNDA.n1585 GNDA.n1563 76.3222
R11593 GNDA.n1766 GNDA.n1765 76.3222
R11594 GNDA.n1776 GNDA.n1775 76.3222
R11595 GNDA.n1777 GNDA.n1557 76.3222
R11596 GNDA.n1788 GNDA.n1787 76.3222
R11597 GNDA.n1789 GNDA.n1553 76.3222
R11598 GNDA.n1825 GNDA.n1823 76.3222
R11599 GNDA.n1821 GNDA.n1818 76.3222
R11600 GNDA.n1816 GNDA.n1815 76.3222
R11601 GNDA.n1813 GNDA.n1810 76.3222
R11602 GNDA.n1808 GNDA.n1807 76.3222
R11603 GNDA.n1803 GNDA.n1802 76.3222
R11604 GNDA.n3166 GNDA.n1801 76.3222
R11605 GNDA.n3161 GNDA.n1806 76.3222
R11606 GNDA.n3159 GNDA.n3158 76.3222
R11607 GNDA.n3154 GNDA.n3153 76.3222
R11608 GNDA.n3151 GNDA.n3150 76.3222
R11609 GNDA.n2955 GNDA.n286 76.3222
R11610 GNDA.n2951 GNDA.n285 76.3222
R11611 GNDA.n2947 GNDA.n284 76.3222
R11612 GNDA.n2943 GNDA.n283 76.3222
R11613 GNDA.n2939 GNDA.n282 76.3222
R11614 GNDA.n264 GNDA.n235 76.3222
R11615 GNDA.n268 GNDA.n236 76.3222
R11616 GNDA.n272 GNDA.n237 76.3222
R11617 GNDA.n240 GNDA.n238 76.3222
R11618 GNDA.n279 GNDA.n239 76.3222
R11619 GNDA.n4859 GNDA.n288 76.3222
R11620 GNDA.n4851 GNDA.n230 76.3222
R11621 GNDA.n4847 GNDA.n231 76.3222
R11622 GNDA.n4843 GNDA.n232 76.3222
R11623 GNDA.n4839 GNDA.n233 76.3222
R11624 GNDA.n3080 GNDA.n3079 74.5978
R11625 GNDA.n3079 GNDA.n3078 74.5978
R11626 GNDA.n2774 GNDA.n1480 74.5978
R11627 GNDA.n2777 GNDA.n1480 74.5978
R11628 GNDA.n5006 GNDA.n175 74.5978
R11629 GNDA.n5003 GNDA.n175 74.5978
R11630 GNDA.n4791 GNDA.n4730 74.5978
R11631 GNDA.n4788 GNDA.n4730 74.5978
R11632 GNDA.n1642 GNDA.n1611 74.5978
R11633 GNDA.n1639 GNDA.n1611 74.5978
R11634 GNDA.n4932 GNDA.n4877 74.5978
R11635 GNDA.n4929 GNDA.n4877 74.5978
R11636 GNDA.n5211 GNDA.n70 74.5978
R11637 GNDA.n5208 GNDA.n70 74.5978
R11638 GNDA.n2868 GNDA.n2678 74.5978
R11639 GNDA.n2869 GNDA.n2868 74.5978
R11640 GNDA.n5129 GNDA.n9 74.5978
R11641 GNDA.n5126 GNDA.n9 74.5978
R11642 GNDA.n2845 GNDA.t200 72.1152
R11643 GNDA.t62 GNDA.t13 70.1899
R11644 GNDA.n4682 GNDA.n4681 69.4466
R11645 GNDA.n3135 GNDA.n3114 69.3109
R11646 GNDA.n3114 GNDA.n3113 69.3109
R11647 GNDA.n3296 GNDA.n3295 69.3109
R11648 GNDA.n3296 GNDA.n1491 69.3109
R11649 GNDA.n5040 GNDA.n168 69.3109
R11650 GNDA.n5040 GNDA.n5039 69.3109
R11651 GNDA.n4825 GNDA.n4723 69.3109
R11652 GNDA.n4825 GNDA.n4824 69.3109
R11653 GNDA.n1705 GNDA.n1704 69.3109
R11654 GNDA.n1705 GNDA.n1623 69.3109
R11655 GNDA.n4974 GNDA.n4867 69.3109
R11656 GNDA.n4950 GNDA.n4867 69.3109
R11657 GNDA.n5253 GNDA.n60 69.3109
R11658 GNDA.n5229 GNDA.n60 69.3109
R11659 GNDA.n2910 GNDA.n2906 69.3109
R11660 GNDA.n2906 GNDA.n2905 69.3109
R11661 GNDA.n5266 GNDA.n5265 69.3109
R11662 GNDA.n5266 GNDA.n20 69.3109
R11663 GNDA.n3141 GNDA.t44 68.1089
R11664 GNDA.n3097 GNDA.t118 65.8183
R11665 GNDA.n3103 GNDA.t118 65.8183
R11666 GNDA.n3105 GNDA.t118 65.8183
R11667 GNDA.n3111 GNDA.t118 65.8183
R11668 GNDA.n3081 GNDA.t118 65.8183
R11669 GNDA.n3087 GNDA.t118 65.8183
R11670 GNDA.n3089 GNDA.t118 65.8183
R11671 GNDA.n3095 GNDA.t118 65.8183
R11672 GNDA.n3065 GNDA.t118 65.8183
R11673 GNDA.n3064 GNDA.t118 65.8183
R11674 GNDA.n3072 GNDA.t118 65.8183
R11675 GNDA.n3060 GNDA.t118 65.8183
R11676 GNDA.n3258 GNDA.t118 65.8183
R11677 GNDA.n3255 GNDA.t118 65.8183
R11678 GNDA.n3123 GNDA.t118 65.8183
R11679 GNDA.n3115 GNDA.t118 65.8183
R11680 GNDA.t100 GNDA.n1490 65.8183
R11681 GNDA.t100 GNDA.n1489 65.8183
R11682 GNDA.t100 GNDA.n1488 65.8183
R11683 GNDA.t100 GNDA.n1487 65.8183
R11684 GNDA.t100 GNDA.n1478 65.8183
R11685 GNDA.t100 GNDA.n1485 65.8183
R11686 GNDA.t100 GNDA.n1476 65.8183
R11687 GNDA.t100 GNDA.n1486 65.8183
R11688 GNDA.t100 GNDA.n1484 65.8183
R11689 GNDA.t100 GNDA.n1483 65.8183
R11690 GNDA.t100 GNDA.n1482 65.8183
R11691 GNDA.t100 GNDA.n1481 65.8183
R11692 GNDA.t100 GNDA.n1479 65.8183
R11693 GNDA.n3297 GNDA.t100 65.8183
R11694 GNDA.t100 GNDA.n1477 65.8183
R11695 GNDA.t100 GNDA.n1475 65.8183
R11696 GNDA.t63 GNDA.n185 65.8183
R11697 GNDA.t63 GNDA.n184 65.8183
R11698 GNDA.t63 GNDA.n183 65.8183
R11699 GNDA.t63 GNDA.n182 65.8183
R11700 GNDA.t63 GNDA.n173 65.8183
R11701 GNDA.t63 GNDA.n180 65.8183
R11702 GNDA.t63 GNDA.n170 65.8183
R11703 GNDA.t63 GNDA.n181 65.8183
R11704 GNDA.t63 GNDA.n179 65.8183
R11705 GNDA.t63 GNDA.n178 65.8183
R11706 GNDA.t63 GNDA.n177 65.8183
R11707 GNDA.t63 GNDA.n176 65.8183
R11708 GNDA.t63 GNDA.n174 65.8183
R11709 GNDA.t63 GNDA.n172 65.8183
R11710 GNDA.t63 GNDA.n171 65.8183
R11711 GNDA.n5041 GNDA.t63 65.8183
R11712 GNDA.t128 GNDA.n4740 65.8183
R11713 GNDA.t128 GNDA.n4739 65.8183
R11714 GNDA.t128 GNDA.n4738 65.8183
R11715 GNDA.t128 GNDA.n4737 65.8183
R11716 GNDA.t128 GNDA.n4728 65.8183
R11717 GNDA.t128 GNDA.n4735 65.8183
R11718 GNDA.t128 GNDA.n4725 65.8183
R11719 GNDA.t128 GNDA.n4736 65.8183
R11720 GNDA.t128 GNDA.n4734 65.8183
R11721 GNDA.t128 GNDA.n4733 65.8183
R11722 GNDA.t128 GNDA.n4732 65.8183
R11723 GNDA.t128 GNDA.n4731 65.8183
R11724 GNDA.t102 GNDA.n1622 65.8183
R11725 GNDA.t102 GNDA.n1621 65.8183
R11726 GNDA.t102 GNDA.n1620 65.8183
R11727 GNDA.t102 GNDA.n1619 65.8183
R11728 GNDA.t102 GNDA.n1610 65.8183
R11729 GNDA.t102 GNDA.n1617 65.8183
R11730 GNDA.t102 GNDA.n1607 65.8183
R11731 GNDA.t102 GNDA.n1618 65.8183
R11732 GNDA.t102 GNDA.n1616 65.8183
R11733 GNDA.t102 GNDA.n1614 65.8183
R11734 GNDA.t102 GNDA.n1613 65.8183
R11735 GNDA.t102 GNDA.n1612 65.8183
R11736 GNDA.n1706 GNDA.t102 65.8183
R11737 GNDA.t102 GNDA.n1609 65.8183
R11738 GNDA.t102 GNDA.n1608 65.8183
R11739 GNDA.t102 GNDA.n1606 65.8183
R11740 GNDA.t117 GNDA.n4964 65.8183
R11741 GNDA.t117 GNDA.n4886 65.8183
R11742 GNDA.t117 GNDA.n4885 65.8183
R11743 GNDA.t117 GNDA.n4884 65.8183
R11744 GNDA.t117 GNDA.n4875 65.8183
R11745 GNDA.t117 GNDA.n4882 65.8183
R11746 GNDA.t117 GNDA.n4873 65.8183
R11747 GNDA.t117 GNDA.n4883 65.8183
R11748 GNDA.t117 GNDA.n4881 65.8183
R11749 GNDA.t117 GNDA.n4880 65.8183
R11750 GNDA.t117 GNDA.n4879 65.8183
R11751 GNDA.t117 GNDA.n4878 65.8183
R11752 GNDA.t117 GNDA.n4876 65.8183
R11753 GNDA.t117 GNDA.n4874 65.8183
R11754 GNDA.n4965 GNDA.t117 65.8183
R11755 GNDA.t117 GNDA.n4868 65.8183
R11756 GNDA.t61 GNDA.n5243 65.8183
R11757 GNDA.t61 GNDA.n79 65.8183
R11758 GNDA.t61 GNDA.n78 65.8183
R11759 GNDA.t61 GNDA.n77 65.8183
R11760 GNDA.t61 GNDA.n68 65.8183
R11761 GNDA.t61 GNDA.n75 65.8183
R11762 GNDA.t61 GNDA.n66 65.8183
R11763 GNDA.t61 GNDA.n76 65.8183
R11764 GNDA.t61 GNDA.n74 65.8183
R11765 GNDA.t61 GNDA.n73 65.8183
R11766 GNDA.t61 GNDA.n72 65.8183
R11767 GNDA.t61 GNDA.n71 65.8183
R11768 GNDA.t61 GNDA.n69 65.8183
R11769 GNDA.t61 GNDA.n67 65.8183
R11770 GNDA.n5244 GNDA.t61 65.8183
R11771 GNDA.t61 GNDA.n61 65.8183
R11772 GNDA.t128 GNDA.n4729 65.8183
R11773 GNDA.t128 GNDA.n4727 65.8183
R11774 GNDA.t128 GNDA.n4726 65.8183
R11775 GNDA.n4826 GNDA.t128 65.8183
R11776 GNDA.n2890 GNDA.t145 65.8183
R11777 GNDA.n2892 GNDA.t145 65.8183
R11778 GNDA.n2898 GNDA.t145 65.8183
R11779 GNDA.n2900 GNDA.t145 65.8183
R11780 GNDA.n2874 GNDA.t145 65.8183
R11781 GNDA.n2876 GNDA.t145 65.8183
R11782 GNDA.n2882 GNDA.t145 65.8183
R11783 GNDA.n2884 GNDA.t145 65.8183
R11784 GNDA.n2685 GNDA.t145 65.8183
R11785 GNDA.n2859 GNDA.t145 65.8183
R11786 GNDA.n2682 GNDA.t145 65.8183
R11787 GNDA.n2866 GNDA.t145 65.8183
R11788 GNDA.n2852 GNDA.t145 65.8183
R11789 GNDA.n2837 GNDA.t145 65.8183
R11790 GNDA.n2835 GNDA.t145 65.8183
R11791 GNDA.n2912 GNDA.t145 65.8183
R11792 GNDA.t106 GNDA.n19 65.8183
R11793 GNDA.t106 GNDA.n18 65.8183
R11794 GNDA.t106 GNDA.n17 65.8183
R11795 GNDA.t106 GNDA.n16 65.8183
R11796 GNDA.t106 GNDA.n7 65.8183
R11797 GNDA.t106 GNDA.n14 65.8183
R11798 GNDA.t106 GNDA.n5 65.8183
R11799 GNDA.t106 GNDA.n15 65.8183
R11800 GNDA.t106 GNDA.n13 65.8183
R11801 GNDA.t106 GNDA.n12 65.8183
R11802 GNDA.t106 GNDA.n11 65.8183
R11803 GNDA.t106 GNDA.n10 65.8183
R11804 GNDA.t106 GNDA.n8 65.8183
R11805 GNDA.n5267 GNDA.t106 65.8183
R11806 GNDA.t106 GNDA.n6 65.8183
R11807 GNDA.t106 GNDA.n4 65.8183
R11808 GNDA.n3613 GNDA.t131 62.2505
R11809 GNDA.n1451 GNDA.t96 62.2505
R11810 GNDA.n584 GNDA.t78 62.2505
R11811 GNDA.n588 GNDA.t75 62.2505
R11812 GNDA.n3608 GNDA.t90 62.2505
R11813 GNDA.n3339 GNDA.t81 62.2505
R11814 GNDA.n3582 GNDA.t136 62.2505
R11815 GNDA.n585 GNDA.t113 62.2505
R11816 GNDA.n3573 GNDA.t147 62.2505
R11817 GNDA.n587 GNDA.t127 62.2505
R11818 GNDA.n573 GNDA.t149 62.2505
R11819 GNDA.n3327 GNDA.t138 62.2505
R11820 GNDA.n3290 GNDA.t39 62.0993
R11821 GNDA.n3140 GNDA.t37 62.0993
R11822 GNDA.t19 GNDA.t194 60.2941
R11823 GNDA.n3382 GNDA.n3381 59.2425
R11824 GNDA.n4612 GNDA.n4611 59.2425
R11825 GNDA.n3850 GNDA.n432 59.2425
R11826 GNDA.n3384 GNDA.n3383 59.2425
R11827 GNDA.t41 GNDA.t211 58.8586
R11828 GNDA.t244 GNDA.n2846 58.0929
R11829 GNDA.n2724 GNDA.t310 58.0929
R11830 GNDA.n3340 GNDA.n3325 57.8952
R11831 GNDA.n3114 GNDA.t118 57.8461
R11832 GNDA.t100 GNDA.n3296 57.8461
R11833 GNDA.t63 GNDA.n5040 57.8461
R11834 GNDA.t102 GNDA.n1705 57.8461
R11835 GNDA.t117 GNDA.n4867 57.8461
R11836 GNDA.t61 GNDA.n60 57.8461
R11837 GNDA.t128 GNDA.n4825 57.8461
R11838 GNDA.n2906 GNDA.t145 57.8461
R11839 GNDA.t106 GNDA.n5266 57.8461
R11840 GNDA.n2737 GNDA.n1497 57.0913
R11841 GNDA.n2802 GNDA.n1829 57.0913
R11842 GNDA.t302 GNDA.t289 56.7747
R11843 GNDA.n1535 GNDA.n1532 56.3995
R11844 GNDA.n1717 GNDA.n1600 56.3995
R11845 GNDA.n4862 GNDA.n4861 56.3995
R11846 GNDA.n4838 GNDA.n234 56.3995
R11847 GNDA.n1532 GNDA.n1530 56.3995
R11848 GNDA.n1717 GNDA.n1716 56.3995
R11849 GNDA.n5093 GNDA.n5092 56.3995
R11850 GNDA.n5094 GNDA.n5093 56.3995
R11851 GNDA.n1856 GNDA.n280 56.3995
R11852 GNDA.n4861 GNDA.n227 56.3995
R11853 GNDA.n4836 GNDA.n234 56.3995
R11854 GNDA.n3079 GNDA.t118 55.2026
R11855 GNDA.t100 GNDA.n1480 55.2026
R11856 GNDA.t63 GNDA.n175 55.2026
R11857 GNDA.t128 GNDA.n4730 55.2026
R11858 GNDA.t102 GNDA.n1611 55.2026
R11859 GNDA.t117 GNDA.n4877 55.2026
R11860 GNDA.t61 GNDA.n70 55.2026
R11861 GNDA.n2868 GNDA.t145 55.2026
R11862 GNDA.t106 GNDA.n9 55.2026
R11863 GNDA.n3096 GNDA.n3095 53.3664
R11864 GNDA.n3089 GNDA.n3054 53.3664
R11865 GNDA.n3088 GNDA.n3087 53.3664
R11866 GNDA.n3081 GNDA.n3056 53.3664
R11867 GNDA.n3074 GNDA.n3060 53.3664
R11868 GNDA.n3072 GNDA.n3071 53.3664
R11869 GNDA.n3067 GNDA.n3064 53.3664
R11870 GNDA.n3065 GNDA.n1512 53.3664
R11871 GNDA.n3134 GNDA.n3115 53.3664
R11872 GNDA.n3124 GNDA.n3123 53.3664
R11873 GNDA.n3255 GNDA.n3254 53.3664
R11874 GNDA.n3258 GNDA.n3257 53.3664
R11875 GNDA.n3097 GNDA.n3052 53.3664
R11876 GNDA.n3103 GNDA.n3102 53.3664
R11877 GNDA.n3106 GNDA.n3105 53.3664
R11878 GNDA.n3111 GNDA.n3110 53.3664
R11879 GNDA.n3098 GNDA.n3097 53.3664
R11880 GNDA.n3104 GNDA.n3103 53.3664
R11881 GNDA.n3105 GNDA.n3050 53.3664
R11882 GNDA.n3112 GNDA.n3111 53.3664
R11883 GNDA.n3082 GNDA.n3081 53.3664
R11884 GNDA.n3087 GNDA.n3086 53.3664
R11885 GNDA.n3090 GNDA.n3089 53.3664
R11886 GNDA.n3095 GNDA.n3094 53.3664
R11887 GNDA.n3066 GNDA.n3065 53.3664
R11888 GNDA.n3064 GNDA.n3061 53.3664
R11889 GNDA.n3073 GNDA.n3072 53.3664
R11890 GNDA.n3060 GNDA.n3058 53.3664
R11891 GNDA.n3259 GNDA.n3258 53.3664
R11892 GNDA.n3256 GNDA.n3255 53.3664
R11893 GNDA.n3123 GNDA.n1515 53.3664
R11894 GNDA.n3122 GNDA.n3115 53.3664
R11895 GNDA.n2758 GNDA.n1486 53.3664
R11896 GNDA.n2762 GNDA.n1476 53.3664
R11897 GNDA.n2766 GNDA.n1485 53.3664
R11898 GNDA.n2770 GNDA.n1478 53.3664
R11899 GNDA.n2781 GNDA.n1481 53.3664
R11900 GNDA.n2785 GNDA.n1482 53.3664
R11901 GNDA.n2789 GNDA.n1483 53.3664
R11902 GNDA.n2793 GNDA.n1484 53.3664
R11903 GNDA.n1492 GNDA.n1475 53.3664
R11904 GNDA.n3285 GNDA.n1477 53.3664
R11905 GNDA.n3298 GNDA.n3297 53.3664
R11906 GNDA.n2727 GNDA.n1479 53.3664
R11907 GNDA.n2754 GNDA.n1490 53.3664
R11908 GNDA.n2753 GNDA.n1489 53.3664
R11909 GNDA.n2749 GNDA.n1488 53.3664
R11910 GNDA.n2745 GNDA.n1487 53.3664
R11911 GNDA.n2757 GNDA.n1490 53.3664
R11912 GNDA.n2750 GNDA.n1489 53.3664
R11913 GNDA.n2746 GNDA.n1488 53.3664
R11914 GNDA.n2742 GNDA.n1487 53.3664
R11915 GNDA.n2773 GNDA.n1478 53.3664
R11916 GNDA.n2769 GNDA.n1485 53.3664
R11917 GNDA.n2765 GNDA.n1476 53.3664
R11918 GNDA.n2761 GNDA.n1486 53.3664
R11919 GNDA.n2790 GNDA.n1484 53.3664
R11920 GNDA.n2786 GNDA.n1483 53.3664
R11921 GNDA.n2782 GNDA.n1482 53.3664
R11922 GNDA.n2778 GNDA.n1481 53.3664
R11923 GNDA.n2792 GNDA.n1479 53.3664
R11924 GNDA.n3297 GNDA.n1474 53.3664
R11925 GNDA.n1477 GNDA.n1473 53.3664
R11926 GNDA.n3284 GNDA.n1475 53.3664
R11927 GNDA.n5022 GNDA.n181 53.3664
R11928 GNDA.n5018 GNDA.n170 53.3664
R11929 GNDA.n5014 GNDA.n180 53.3664
R11930 GNDA.n5010 GNDA.n173 53.3664
R11931 GNDA.n4999 GNDA.n176 53.3664
R11932 GNDA.n4995 GNDA.n177 53.3664
R11933 GNDA.n4991 GNDA.n178 53.3664
R11934 GNDA.n4987 GNDA.n179 53.3664
R11935 GNDA.n5042 GNDA.n5041 53.3664
R11936 GNDA.n216 GNDA.n171 53.3664
R11937 GNDA.n212 GNDA.n172 53.3664
R11938 GNDA.n205 GNDA.n174 53.3664
R11939 GNDA.n5026 GNDA.n185 53.3664
R11940 GNDA.n5027 GNDA.n184 53.3664
R11941 GNDA.n5031 GNDA.n183 53.3664
R11942 GNDA.n5035 GNDA.n182 53.3664
R11943 GNDA.n5023 GNDA.n185 53.3664
R11944 GNDA.n5030 GNDA.n184 53.3664
R11945 GNDA.n5034 GNDA.n183 53.3664
R11946 GNDA.n5038 GNDA.n182 53.3664
R11947 GNDA.n5007 GNDA.n173 53.3664
R11948 GNDA.n5011 GNDA.n180 53.3664
R11949 GNDA.n5015 GNDA.n170 53.3664
R11950 GNDA.n5019 GNDA.n181 53.3664
R11951 GNDA.n4990 GNDA.n179 53.3664
R11952 GNDA.n4994 GNDA.n178 53.3664
R11953 GNDA.n4998 GNDA.n177 53.3664
R11954 GNDA.n5002 GNDA.n176 53.3664
R11955 GNDA.n4986 GNDA.n174 53.3664
R11956 GNDA.n204 GNDA.n172 53.3664
R11957 GNDA.n213 GNDA.n171 53.3664
R11958 GNDA.n5041 GNDA.n169 53.3664
R11959 GNDA.n4807 GNDA.n4736 53.3664
R11960 GNDA.n4803 GNDA.n4725 53.3664
R11961 GNDA.n4799 GNDA.n4735 53.3664
R11962 GNDA.n4795 GNDA.n4728 53.3664
R11963 GNDA.n4784 GNDA.n4731 53.3664
R11964 GNDA.n4780 GNDA.n4732 53.3664
R11965 GNDA.n4776 GNDA.n4733 53.3664
R11966 GNDA.n4772 GNDA.n4734 53.3664
R11967 GNDA.n4827 GNDA.n4826 53.3664
R11968 GNDA.n4749 GNDA.n4726 53.3664
R11969 GNDA.n4757 GNDA.n4727 53.3664
R11970 GNDA.n4764 GNDA.n4729 53.3664
R11971 GNDA.n4811 GNDA.n4740 53.3664
R11972 GNDA.n4812 GNDA.n4739 53.3664
R11973 GNDA.n4816 GNDA.n4738 53.3664
R11974 GNDA.n4820 GNDA.n4737 53.3664
R11975 GNDA.n4808 GNDA.n4740 53.3664
R11976 GNDA.n4815 GNDA.n4739 53.3664
R11977 GNDA.n4819 GNDA.n4738 53.3664
R11978 GNDA.n4823 GNDA.n4737 53.3664
R11979 GNDA.n4792 GNDA.n4728 53.3664
R11980 GNDA.n4796 GNDA.n4735 53.3664
R11981 GNDA.n4800 GNDA.n4725 53.3664
R11982 GNDA.n4804 GNDA.n4736 53.3664
R11983 GNDA.n4775 GNDA.n4734 53.3664
R11984 GNDA.n4779 GNDA.n4733 53.3664
R11985 GNDA.n4783 GNDA.n4732 53.3664
R11986 GNDA.n4787 GNDA.n4731 53.3664
R11987 GNDA.n1658 GNDA.n1618 53.3664
R11988 GNDA.n1654 GNDA.n1607 53.3664
R11989 GNDA.n1650 GNDA.n1617 53.3664
R11990 GNDA.n1646 GNDA.n1610 53.3664
R11991 GNDA.n1635 GNDA.n1612 53.3664
R11992 GNDA.n1631 GNDA.n1613 53.3664
R11993 GNDA.n1627 GNDA.n1614 53.3664
R11994 GNDA.n1616 GNDA.n1615 53.3664
R11995 GNDA.n1624 GNDA.n1606 53.3664
R11996 GNDA.n1693 GNDA.n1608 53.3664
R11997 GNDA.n1686 GNDA.n1609 53.3664
R11998 GNDA.n1707 GNDA.n1706 53.3664
R11999 GNDA.n1662 GNDA.n1622 53.3664
R12000 GNDA.n1663 GNDA.n1621 53.3664
R12001 GNDA.n1667 GNDA.n1620 53.3664
R12002 GNDA.n1671 GNDA.n1619 53.3664
R12003 GNDA.n1659 GNDA.n1622 53.3664
R12004 GNDA.n1666 GNDA.n1621 53.3664
R12005 GNDA.n1670 GNDA.n1620 53.3664
R12006 GNDA.n1673 GNDA.n1619 53.3664
R12007 GNDA.n1643 GNDA.n1610 53.3664
R12008 GNDA.n1647 GNDA.n1617 53.3664
R12009 GNDA.n1651 GNDA.n1607 53.3664
R12010 GNDA.n1655 GNDA.n1618 53.3664
R12011 GNDA.n1626 GNDA.n1616 53.3664
R12012 GNDA.n1630 GNDA.n1614 53.3664
R12013 GNDA.n1634 GNDA.n1613 53.3664
R12014 GNDA.n1638 GNDA.n1612 53.3664
R12015 GNDA.n1706 GNDA.n1605 53.3664
R12016 GNDA.n1609 GNDA.n1604 53.3664
R12017 GNDA.n1685 GNDA.n1608 53.3664
R12018 GNDA.n1692 GNDA.n1606 53.3664
R12019 GNDA.n4947 GNDA.n4883 53.3664
R12020 GNDA.n4944 GNDA.n4873 53.3664
R12021 GNDA.n4940 GNDA.n4882 53.3664
R12022 GNDA.n4936 GNDA.n4875 53.3664
R12023 GNDA.n4925 GNDA.n4878 53.3664
R12024 GNDA.n4921 GNDA.n4879 53.3664
R12025 GNDA.n4917 GNDA.n4880 53.3664
R12026 GNDA.n4913 GNDA.n4881 53.3664
R12027 GNDA.n4973 GNDA.n4868 53.3664
R12028 GNDA.n4966 GNDA.n4965 53.3664
R12029 GNDA.n4898 GNDA.n4874 53.3664
R12030 GNDA.n4905 GNDA.n4876 53.3664
R12031 GNDA.n4964 GNDA.n4963 53.3664
R12032 GNDA.n4888 GNDA.n4886 53.3664
R12033 GNDA.n4958 GNDA.n4885 53.3664
R12034 GNDA.n4954 GNDA.n4884 53.3664
R12035 GNDA.n4964 GNDA.n4887 53.3664
R12036 GNDA.n4959 GNDA.n4886 53.3664
R12037 GNDA.n4955 GNDA.n4885 53.3664
R12038 GNDA.n4951 GNDA.n4884 53.3664
R12039 GNDA.n4933 GNDA.n4875 53.3664
R12040 GNDA.n4937 GNDA.n4882 53.3664
R12041 GNDA.n4941 GNDA.n4873 53.3664
R12042 GNDA.n4945 GNDA.n4883 53.3664
R12043 GNDA.n4916 GNDA.n4881 53.3664
R12044 GNDA.n4920 GNDA.n4880 53.3664
R12045 GNDA.n4924 GNDA.n4879 53.3664
R12046 GNDA.n4928 GNDA.n4878 53.3664
R12047 GNDA.n4912 GNDA.n4876 53.3664
R12048 GNDA.n4904 GNDA.n4874 53.3664
R12049 GNDA.n4965 GNDA.n4872 53.3664
R12050 GNDA.n4871 GNDA.n4868 53.3664
R12051 GNDA.n5226 GNDA.n76 53.3664
R12052 GNDA.n5223 GNDA.n66 53.3664
R12053 GNDA.n5219 GNDA.n75 53.3664
R12054 GNDA.n5215 GNDA.n68 53.3664
R12055 GNDA.n5204 GNDA.n71 53.3664
R12056 GNDA.n5200 GNDA.n72 53.3664
R12057 GNDA.n5196 GNDA.n73 53.3664
R12058 GNDA.n5192 GNDA.n74 53.3664
R12059 GNDA.n5252 GNDA.n61 53.3664
R12060 GNDA.n5245 GNDA.n5244 53.3664
R12061 GNDA.n5177 GNDA.n67 53.3664
R12062 GNDA.n5184 GNDA.n69 53.3664
R12063 GNDA.n5243 GNDA.n5242 53.3664
R12064 GNDA.n81 GNDA.n79 53.3664
R12065 GNDA.n5237 GNDA.n78 53.3664
R12066 GNDA.n5233 GNDA.n77 53.3664
R12067 GNDA.n5243 GNDA.n80 53.3664
R12068 GNDA.n5238 GNDA.n79 53.3664
R12069 GNDA.n5234 GNDA.n78 53.3664
R12070 GNDA.n5230 GNDA.n77 53.3664
R12071 GNDA.n5212 GNDA.n68 53.3664
R12072 GNDA.n5216 GNDA.n75 53.3664
R12073 GNDA.n5220 GNDA.n66 53.3664
R12074 GNDA.n5224 GNDA.n76 53.3664
R12075 GNDA.n5195 GNDA.n74 53.3664
R12076 GNDA.n5199 GNDA.n73 53.3664
R12077 GNDA.n5203 GNDA.n72 53.3664
R12078 GNDA.n5207 GNDA.n71 53.3664
R12079 GNDA.n5191 GNDA.n69 53.3664
R12080 GNDA.n5183 GNDA.n67 53.3664
R12081 GNDA.n5244 GNDA.n65 53.3664
R12082 GNDA.n64 GNDA.n61 53.3664
R12083 GNDA.n4771 GNDA.n4729 53.3664
R12084 GNDA.n4763 GNDA.n4727 53.3664
R12085 GNDA.n4756 GNDA.n4726 53.3664
R12086 GNDA.n4826 GNDA.n4724 53.3664
R12087 GNDA.n2884 GNDA.n2674 53.3664
R12088 GNDA.n2883 GNDA.n2882 53.3664
R12089 GNDA.n2876 GNDA.n2676 53.3664
R12090 GNDA.n2875 GNDA.n2874 53.3664
R12091 GNDA.n2866 GNDA.n2865 53.3664
R12092 GNDA.n2861 GNDA.n2682 53.3664
R12093 GNDA.n2859 GNDA.n2858 53.3664
R12094 GNDA.n2854 GNDA.n2685 53.3664
R12095 GNDA.n2912 GNDA.n2911 53.3664
R12096 GNDA.n2835 GNDA.n2669 53.3664
R12097 GNDA.n2838 GNDA.n2837 53.3664
R12098 GNDA.n2852 GNDA.n2851 53.3664
R12099 GNDA.n2891 GNDA.n2890 53.3664
R12100 GNDA.n2893 GNDA.n2892 53.3664
R12101 GNDA.n2898 GNDA.n2897 53.3664
R12102 GNDA.n2901 GNDA.n2900 53.3664
R12103 GNDA.n2890 GNDA.n2889 53.3664
R12104 GNDA.n2892 GNDA.n2672 53.3664
R12105 GNDA.n2899 GNDA.n2898 53.3664
R12106 GNDA.n2900 GNDA.n2670 53.3664
R12107 GNDA.n2874 GNDA.n2873 53.3664
R12108 GNDA.n2877 GNDA.n2876 53.3664
R12109 GNDA.n2882 GNDA.n2881 53.3664
R12110 GNDA.n2885 GNDA.n2884 53.3664
R12111 GNDA.n2685 GNDA.n2683 53.3664
R12112 GNDA.n2860 GNDA.n2859 53.3664
R12113 GNDA.n2682 GNDA.n2680 53.3664
R12114 GNDA.n2867 GNDA.n2866 53.3664
R12115 GNDA.n2853 GNDA.n2852 53.3664
R12116 GNDA.n2837 GNDA.n2687 53.3664
R12117 GNDA.n2836 GNDA.n2835 53.3664
R12118 GNDA.n2913 GNDA.n2912 53.3664
R12119 GNDA.n5145 GNDA.n15 53.3664
R12120 GNDA.n5141 GNDA.n5 53.3664
R12121 GNDA.n5137 GNDA.n14 53.3664
R12122 GNDA.n5133 GNDA.n7 53.3664
R12123 GNDA.n5122 GNDA.n10 53.3664
R12124 GNDA.n5118 GNDA.n11 53.3664
R12125 GNDA.n5114 GNDA.n12 53.3664
R12126 GNDA.n5110 GNDA.n13 53.3664
R12127 GNDA.n21 GNDA.n4 53.3664
R12128 GNDA.n37 GNDA.n6 53.3664
R12129 GNDA.n5268 GNDA.n5267 53.3664
R12130 GNDA.n5102 GNDA.n8 53.3664
R12131 GNDA.n5149 GNDA.n19 53.3664
R12132 GNDA.n5150 GNDA.n18 53.3664
R12133 GNDA.n5154 GNDA.n17 53.3664
R12134 GNDA.n5158 GNDA.n16 53.3664
R12135 GNDA.n5146 GNDA.n19 53.3664
R12136 GNDA.n5153 GNDA.n18 53.3664
R12137 GNDA.n5157 GNDA.n17 53.3664
R12138 GNDA.n5160 GNDA.n16 53.3664
R12139 GNDA.n5130 GNDA.n7 53.3664
R12140 GNDA.n5134 GNDA.n14 53.3664
R12141 GNDA.n5138 GNDA.n5 53.3664
R12142 GNDA.n5142 GNDA.n15 53.3664
R12143 GNDA.n5113 GNDA.n13 53.3664
R12144 GNDA.n5117 GNDA.n12 53.3664
R12145 GNDA.n5121 GNDA.n11 53.3664
R12146 GNDA.n5125 GNDA.n10 53.3664
R12147 GNDA.n5109 GNDA.n8 53.3664
R12148 GNDA.n5267 GNDA.n3 53.3664
R12149 GNDA.n6 GNDA.n2 53.3664
R12150 GNDA.n36 GNDA.n4 53.3664
R12151 GNDA.n2931 GNDA.n1859 53.085
R12152 GNDA.n2737 GNDA.n2736 53.085
R12153 GNDA.n2805 GNDA.n2802 53.085
R12154 GNDA.n2846 GNDA.t183 52.0834
R12155 GNDA.n2724 GNDA.t59 52.0834
R12156 GNDA.t156 GNDA.n3249 52.0834
R12157 GNDA.t195 GNDA.t214 52.0435
R12158 GNDA.t192 GNDA.t293 52.0435
R12159 GNDA.t56 GNDA.t223 52.0435
R12160 GNDA.t208 GNDA.t220 52.0435
R12161 GNDA.t57 GNDA.t308 52.0435
R12162 GNDA.t202 GNDA.t17 52.0435
R12163 GNDA.t189 GNDA.t226 52.0435
R12164 GNDA.t300 GNDA.t224 52.0435
R12165 GNDA.t53 GNDA.t242 52.0435
R12166 GNDA.t54 GNDA.t203 52.0435
R12167 GNDA.n4716 GNDA.n99 50.8806
R12168 GNDA.n4716 GNDA.n4715 50.8806
R12169 GNDA.n4715 GNDA.n4714 50.8806
R12170 GNDA.n4714 GNDA.n292 50.8806
R12171 GNDA.n4708 GNDA.n292 50.8806
R12172 GNDA.n4707 GNDA.n4706 50.8806
R12173 GNDA.n4706 GNDA.n296 50.8806
R12174 GNDA.n4700 GNDA.n296 50.8806
R12175 GNDA.n4700 GNDA.n4699 50.8806
R12176 GNDA.n4699 GNDA.n4698 50.8806
R12177 GNDA.n4692 GNDA.n4691 50.8806
R12178 GNDA.n4691 GNDA.n4690 50.8806
R12179 GNDA.n4690 GNDA.n351 50.8806
R12180 GNDA.n4684 GNDA.n351 50.8806
R12181 GNDA.n4684 GNDA.n4683 50.8806
R12182 GNDA.n4674 GNDA.n356 50.8806
R12183 GNDA.n4674 GNDA.n4673 50.8806
R12184 GNDA.n4673 GNDA.n4672 50.8806
R12185 GNDA.n4672 GNDA.n362 50.8806
R12186 GNDA.n4666 GNDA.n362 50.8806
R12187 GNDA.n4664 GNDA.n367 50.8806
R12188 GNDA.n4658 GNDA.n367 50.8806
R12189 GNDA.n4658 GNDA.n4657 50.8806
R12190 GNDA.n4657 GNDA.n4656 50.8806
R12191 GNDA.n4656 GNDA.n416 50.8806
R12192 GNDA.n4650 GNDA.n4649 50.8806
R12193 GNDA.n4649 GNDA.n4648 50.8806
R12194 GNDA.n4648 GNDA.n420 50.8806
R12195 GNDA.n4642 GNDA.n420 50.8806
R12196 GNDA.n4642 GNDA.n4641 50.8806
R12197 GNDA.t80 GNDA.n3340 50.4249
R12198 GNDA.t89 GNDA.n3609 50.4249
R12199 GNDA.t143 GNDA.t153 49.6779
R12200 GNDA.t68 GNDA.t133 49.6779
R12201 GNDA.t124 GNDA.t115 49.6779
R12202 GNDA.t104 GNDA.t140 49.6779
R12203 GNDA.t159 GNDA.n106 48.077
R12204 GNDA.t98 GNDA.n3290 48.077
R12205 GNDA.t251 GNDA.n3140 48.077
R12206 GNDA.t62 GNDA.n5080 47.6748
R12207 GNDA.t207 GNDA.t174 47.3123
R12208 GNDA.t301 GNDA.t190 47.3123
R12209 GNDA.t62 GNDA.n106 47.0754
R12210 GNDA.t270 GNDA.n3144 47.0754
R12211 GNDA.t274 GNDA.n3045 46.0738
R12212 GNDA.n3145 GNDA.n1829 44.0706
R12213 GNDA.n2736 GNDA.n1830 43.069
R12214 GNDA.t62 GNDA.n3302 43.069
R12215 GNDA.n3249 GNDA.t62 43.069
R12216 GNDA.n3291 GNDA.t98 42.0674
R12217 GNDA.n3141 GNDA.t251 42.0674
R12218 GNDA.t239 GNDA.t80 41.0871
R12219 GNDA.t177 GNDA.t239 41.0871
R12220 GNDA.t34 GNDA.t177 41.0871
R12221 GNDA.t86 GNDA.t185 41.0871
R12222 GNDA.t35 GNDA.t86 41.0871
R12223 GNDA.t25 GNDA.t35 41.0871
R12224 GNDA.t112 GNDA.t51 41.0871
R12225 GNDA.t33 GNDA.t29 41.0871
R12226 GNDA.t29 GNDA.t89 41.0871
R12227 GNDA.n3279 GNDA.t165 41.0658
R12228 GNDA.n3342 GNDA.t84 40.4338
R12229 GNDA.n3585 GNDA.t151 40.4338
R12230 GNDA.n3570 GNDA.t87 40.4338
R12231 GNDA.n3610 GNDA.t122 40.4338
R12232 GNDA.t279 GNDA.t195 40.2156
R12233 GNDA.t308 GNDA.t277 40.2156
R12234 GNDA.t17 GNDA.t260 40.2156
R12235 GNDA.t231 GNDA.t54 40.2156
R12236 GNDA.n1450 GNDA.t25 39.2195
R12237 GNDA.t183 GNDA.n2845 38.0611
R12238 GNDA.t59 GNDA.n2720 38.0611
R12239 GNDA.n3364 GNDA.n3363 37.5297
R12240 GNDA.n3362 GNDA.n3361 37.5297
R12241 GNDA.n3360 GNDA.n3359 37.5297
R12242 GNDA.n3358 GNDA.n3357 37.5297
R12243 GNDA.n3356 GNDA.n3355 37.5297
R12244 GNDA.n3354 GNDA.n3353 37.5297
R12245 GNDA.n3352 GNDA.n3351 37.5297
R12246 GNDA.n3350 GNDA.n3349 37.5297
R12247 GNDA.n3348 GNDA.n3347 37.5297
R12248 GNDA.n3346 GNDA.n3345 37.5297
R12249 GNDA.n3344 GNDA.n3343 37.5297
R12250 GNDA.n2932 GNDA.n2931 37.0595
R12251 GNDA.n2665 GNDA.t209 37.0595
R12252 GNDA.t153 GNDA.n432 35.4844
R12253 GNDA.n4612 GNDA.t68 35.4844
R12254 GNDA.n3383 GNDA.t124 35.4844
R12255 GNDA.t140 GNDA.n3382 35.4844
R12256 GNDA.t71 GNDA.t274 35.0563
R12257 GNDA.t92 GNDA.t270 35.0563
R12258 GNDA.n582 GNDA.n581 34.5991
R12259 GNDA.t182 GNDA.t309 33.1455
R12260 GNDA.n2825 GNDA.n2814 33.0531
R12261 GNDA.n3250 GNDA.t228 33.0531
R12262 GNDA.t62 GNDA.n26 32.9056
R12263 GNDA.t62 GNDA.n107 32.9056
R12264 GNDA.n3246 GNDA.n3234 32.3969
R12265 GNDA.t310 GNDA.n2723 32.0515
R12266 GNDA.n3341 GNDA.t166 31.7492
R12267 GNDA.n3584 GNDA.t3 31.7492
R12268 GNDA.t30 GNDA.n3611 31.7492
R12269 GNDA.n573 GNDA.n572 31.5738
R12270 GNDA.n4679 GNDA.n4678 31.3605
R12271 GNDA.n4619 GNDA.t154 31.1255
R12272 GNDA.n4614 GNDA.t69 31.1255
R12273 GNDA.n745 GNDA.t141 31.1255
R12274 GNDA.n741 GNDA.t125 31.1255
R12275 GNDA.t262 GNDA.t192 30.7532
R12276 GNDA.t220 GNDA.t256 30.7532
R12277 GNDA.t226 GNDA.t237 30.7532
R12278 GNDA.t282 GNDA.t53 30.7532
R12279 GNDA.t65 GNDA.t9 30.3834
R12280 GNDA.t9 GNDA.t296 30.3834
R12281 GNDA.t296 GNDA.t187 30.3834
R12282 GNDA.n3277 GNDA.n1497 30.0483
R12283 GNDA.n2805 GNDA.n2801 30.0483
R12284 GNDA.n3608 GNDA.n3607 29.8672
R12285 GNDA.n3339 GNDA.n3338 29.8672
R12286 GNDA.n3327 GNDA.n3326 29.8672
R12287 GNDA.n3045 GNDA.t200 29.0467
R12288 GNDA.n4620 GNDA.n432 28.3876
R12289 GNDA.n4613 GNDA.n4612 28.3876
R12290 GNDA.n3383 GNDA.n742 28.3876
R12291 GNDA.n3382 GNDA.n746 28.3876
R12292 GNDA.t39 GNDA.n3289 28.0451
R12293 GNDA.n3144 GNDA.t44 28.0451
R12294 GNDA.n3099 GNDA.n3053 27.5561
R12295 GNDA.n2759 GNDA.n2756 27.5561
R12296 GNDA.n5024 GNDA.n5021 27.5561
R12297 GNDA.n4809 GNDA.n4806 27.5561
R12298 GNDA.n1660 GNDA.n1657 27.5561
R12299 GNDA.n4949 GNDA.n4948 27.5561
R12300 GNDA.n5228 GNDA.n5227 27.5561
R12301 GNDA.n2888 GNDA.n2887 27.5561
R12302 GNDA.n5147 GNDA.n5144 27.5561
R12303 GNDA.n3248 GNDA.n1520 27.0435
R12304 GNDA.n3077 GNDA.n3057 26.6672
R12305 GNDA.n2776 GNDA.n2775 26.6672
R12306 GNDA.n5005 GNDA.n5004 26.6672
R12307 GNDA.n4790 GNDA.n4789 26.6672
R12308 GNDA.n1641 GNDA.n1640 26.6672
R12309 GNDA.n4931 GNDA.n4930 26.6672
R12310 GNDA.n5210 GNDA.n5209 26.6672
R12311 GNDA.n2871 GNDA.n2870 26.6672
R12312 GNDA.n5128 GNDA.n5127 26.6672
R12313 GNDA.n4708 GNDA.t62 26.5712
R12314 GNDA.n4683 GNDA.t62 26.5712
R12315 GNDA.t62 GNDA.n416 26.5712
R12316 GNDA.n2817 GNDA.n2816 25.3679
R12317 GNDA.t15 GNDA.t244 25.0403
R12318 GNDA.t37 GNDA.t175 25.0403
R12319 GNDA.t62 GNDA.n4707 24.3099
R12320 GNDA.t62 GNDA.n356 24.3099
R12321 GNDA.n4650 GNDA.t62 24.3099
R12322 GNDA.t217 GNDA.t229 24.2789
R12323 GNDA.n3222 GNDA.n3221 24.0387
R12324 GNDA.n1505 GNDA.t248 24.0005
R12325 GNDA.n1505 GNDA.t254 24.0005
R12326 GNDA.n1504 GNDA.t38 24.0005
R12327 GNDA.n1504 GNDA.t47 24.0005
R12328 GNDA.n1503 GNDA.t45 24.0005
R12329 GNDA.n1503 GNDA.t252 24.0005
R12330 GNDA.n1500 GNDA.t236 24.0005
R12331 GNDA.n1500 GNDA.t311 24.0005
R12332 GNDA.n1499 GNDA.t40 24.0005
R12333 GNDA.n1499 GNDA.t198 24.0005
R12334 GNDA.n2923 GNDA.t184 24.0005
R12335 GNDA.n2923 GNDA.t201 24.0005
R12336 GNDA.n2922 GNDA.t216 24.0005
R12337 GNDA.n2922 GNDA.t245 24.0005
R12338 GNDA.n2921 GNDA.t234 24.0005
R12339 GNDA.n2921 GNDA.t169 24.0005
R12340 GNDA.n2662 GNDA.t188 24.0005
R12341 GNDA.n2662 GNDA.t109 24.0005
R12342 GNDA.n2660 GNDA.t10 24.0005
R12343 GNDA.n2660 GNDA.t297 24.0005
R12344 GNDA.n2656 GNDA.t181 23.4782
R12345 GNDA.n2828 GNDA.n2827 23.0371
R12346 GNDA.t83 GNDA.t205 22.4114
R12347 GNDA.t11 GNDA.t172 22.4114
R12348 GNDA.t170 GNDA.t20 22.4114
R12349 GNDA.t163 GNDA.t55 22.4114
R12350 GNDA.t284 GNDA.t227 22.4114
R12351 GNDA.t298 GNDA.t212 22.4114
R12352 GNDA.t5 GNDA.t74 22.4114
R12353 GNDA.t77 GNDA.t49 22.4114
R12354 GNDA.t27 GNDA.t258 22.4114
R12355 GNDA.t32 GNDA.t1 22.4114
R12356 GNDA.t24 GNDA.t7 22.4114
R12357 GNDA.t28 GNDA.t249 22.4114
R12358 GNDA.t26 GNDA.t161 22.4114
R12359 GNDA.t31 GNDA.t286 22.4114
R12360 GNDA.t23 GNDA.t120 22.4114
R12361 GNDA.t223 GNDA.t262 21.2908
R12362 GNDA.t256 GNDA.t56 21.2908
R12363 GNDA.t237 GNDA.t300 21.2908
R12364 GNDA.t224 GNDA.t282 21.2908
R12365 GNDA.n3266 GNDA.n3265 20.8233
R12366 GNDA.n1828 GNDA.n1502 20.8233
R12367 GNDA.n2800 GNDA.n1501 20.8233
R12368 GNDA.n3276 GNDA.n3275 20.8233
R12369 GNDA.n2735 GNDA.n2734 20.8233
R12370 GNDA.n2920 GNDA.n2919 20.8233
R12371 GNDA.n2930 GNDA.n2929 20.8233
R12372 GNDA.n2658 GNDA.n2657 20.8233
R12373 GNDA.n460 GNDA.t304 19.7005
R12374 GNDA.n460 GNDA.t269 19.7005
R12375 GNDA.n458 GNDA.t222 19.7005
R12376 GNDA.n458 GNDA.t219 19.7005
R12377 GNDA.n456 GNDA.t243 19.7005
R12378 GNDA.n456 GNDA.t294 19.7005
R12379 GNDA.n454 GNDA.t22 19.7005
R12380 GNDA.n454 GNDA.t295 19.7005
R12381 GNDA.n452 GNDA.t191 19.7005
R12382 GNDA.n452 GNDA.t241 19.7005
R12383 GNDA.n451 GNDA.t268 19.7005
R12384 GNDA.n451 GNDA.t221 19.7005
R12385 GNDA.n3556 GNDA.t292 19.7005
R12386 GNDA.n3556 GNDA.t267 19.7005
R12387 GNDA.n3554 GNDA.t306 19.7005
R12388 GNDA.n3554 GNDA.t204 19.7005
R12389 GNDA.n3552 GNDA.t210 19.7005
R12390 GNDA.n3552 GNDA.t18 19.7005
R12391 GNDA.n3550 GNDA.t225 19.7005
R12392 GNDA.n3550 GNDA.t288 19.7005
R12393 GNDA.n3548 GNDA.t0 19.7005
R12394 GNDA.n3548 GNDA.t16 19.7005
R12395 GNDA.n3546 GNDA.t266 19.7005
R12396 GNDA.n3546 GNDA.t291 19.7005
R12397 GNDA.t166 GNDA.t83 18.6762
R12398 GNDA.t205 GNDA.t11 18.6762
R12399 GNDA.t172 GNDA.t170 18.6762
R12400 GNDA.t20 GNDA.t163 18.6762
R12401 GNDA.t55 GNDA.t284 18.6762
R12402 GNDA.t227 GNDA.t298 18.6762
R12403 GNDA.t212 GNDA.t5 18.6762
R12404 GNDA.t74 GNDA.t217 18.6762
R12405 GNDA.t161 GNDA.t31 18.6762
R12406 GNDA.t286 GNDA.t23 18.6762
R12407 GNDA.t120 GNDA.t30 18.6762
R12408 GNDA.n3195 GNDA.n1543 17.5843
R12409 GNDA.n1741 GNDA.n1589 17.5843
R12410 GNDA.n4638 GNDA.n422 17.5843
R12411 GNDA.n4634 GNDA.n4627 17.5479
R12412 GNDA.t196 GNDA.t179 17.2273
R12413 GNDA.t211 GNDA.t196 17.2273
R12414 GNDA.t178 GNDA.t19 17.2273
R12415 GNDA.t305 GNDA.t178 17.2273
R12416 GNDA.n262 GNDA.n259 16.9379
R12417 GNDA.n4857 GNDA.n4719 16.9379
R12418 GNDA.n2958 GNDA.n2957 16.9379
R12419 GNDA.n3612 GNDA.t249 16.8086
R12420 GNDA.n5076 GNDA.n133 16.7709
R12421 GNDA.n2982 GNDA.n162 16.7709
R12422 GNDA.n1588 GNDA.n84 16.7709
R12423 GNDA.n1800 GNDA.n1799 16.7709
R12424 GNDA.t62 GNDA.n105 16.4553
R12425 GNDA.n3100 GNDA.n3099 16.0005
R12426 GNDA.n3101 GNDA.n3100 16.0005
R12427 GNDA.n3101 GNDA.n3051 16.0005
R12428 GNDA.n3107 GNDA.n3051 16.0005
R12429 GNDA.n3108 GNDA.n3107 16.0005
R12430 GNDA.n3109 GNDA.n3108 16.0005
R12431 GNDA.n3109 GNDA.n3049 16.0005
R12432 GNDA.n3049 GNDA.n3047 16.0005
R12433 GNDA.n3093 GNDA.n3053 16.0005
R12434 GNDA.n3093 GNDA.n3092 16.0005
R12435 GNDA.n3092 GNDA.n3091 16.0005
R12436 GNDA.n3091 GNDA.n3055 16.0005
R12437 GNDA.n3085 GNDA.n3055 16.0005
R12438 GNDA.n3085 GNDA.n3084 16.0005
R12439 GNDA.n3084 GNDA.n3083 16.0005
R12440 GNDA.n3083 GNDA.n3057 16.0005
R12441 GNDA.n3077 GNDA.n3076 16.0005
R12442 GNDA.n3076 GNDA.n3075 16.0005
R12443 GNDA.n3075 GNDA.n3059 16.0005
R12444 GNDA.n3070 GNDA.n3059 16.0005
R12445 GNDA.n3070 GNDA.n3069 16.0005
R12446 GNDA.n3069 GNDA.n3068 16.0005
R12447 GNDA.n3068 GNDA.n3063 16.0005
R12448 GNDA.n3063 GNDA.n3062 16.0005
R12449 GNDA.n2756 GNDA.n2755 16.0005
R12450 GNDA.n2755 GNDA.n2752 16.0005
R12451 GNDA.n2752 GNDA.n2751 16.0005
R12452 GNDA.n2751 GNDA.n2748 16.0005
R12453 GNDA.n2748 GNDA.n2747 16.0005
R12454 GNDA.n2747 GNDA.n2744 16.0005
R12455 GNDA.n2744 GNDA.n2743 16.0005
R12456 GNDA.n2743 GNDA.n2741 16.0005
R12457 GNDA.n2760 GNDA.n2759 16.0005
R12458 GNDA.n2763 GNDA.n2760 16.0005
R12459 GNDA.n2764 GNDA.n2763 16.0005
R12460 GNDA.n2767 GNDA.n2764 16.0005
R12461 GNDA.n2768 GNDA.n2767 16.0005
R12462 GNDA.n2771 GNDA.n2768 16.0005
R12463 GNDA.n2772 GNDA.n2771 16.0005
R12464 GNDA.n2775 GNDA.n2772 16.0005
R12465 GNDA.n2779 GNDA.n2776 16.0005
R12466 GNDA.n2780 GNDA.n2779 16.0005
R12467 GNDA.n2783 GNDA.n2780 16.0005
R12468 GNDA.n2784 GNDA.n2783 16.0005
R12469 GNDA.n2787 GNDA.n2784 16.0005
R12470 GNDA.n2788 GNDA.n2787 16.0005
R12471 GNDA.n2791 GNDA.n2788 16.0005
R12472 GNDA.n2794 GNDA.n2791 16.0005
R12473 GNDA.n5025 GNDA.n5024 16.0005
R12474 GNDA.n5028 GNDA.n5025 16.0005
R12475 GNDA.n5029 GNDA.n5028 16.0005
R12476 GNDA.n5032 GNDA.n5029 16.0005
R12477 GNDA.n5033 GNDA.n5032 16.0005
R12478 GNDA.n5036 GNDA.n5033 16.0005
R12479 GNDA.n5037 GNDA.n5036 16.0005
R12480 GNDA.n5037 GNDA.n164 16.0005
R12481 GNDA.n5021 GNDA.n5020 16.0005
R12482 GNDA.n5020 GNDA.n5017 16.0005
R12483 GNDA.n5017 GNDA.n5016 16.0005
R12484 GNDA.n5016 GNDA.n5013 16.0005
R12485 GNDA.n5013 GNDA.n5012 16.0005
R12486 GNDA.n5012 GNDA.n5009 16.0005
R12487 GNDA.n5009 GNDA.n5008 16.0005
R12488 GNDA.n5008 GNDA.n5005 16.0005
R12489 GNDA.n5004 GNDA.n5001 16.0005
R12490 GNDA.n5001 GNDA.n5000 16.0005
R12491 GNDA.n5000 GNDA.n4997 16.0005
R12492 GNDA.n4997 GNDA.n4996 16.0005
R12493 GNDA.n4996 GNDA.n4993 16.0005
R12494 GNDA.n4993 GNDA.n4992 16.0005
R12495 GNDA.n4992 GNDA.n4989 16.0005
R12496 GNDA.n4989 GNDA.n4988 16.0005
R12497 GNDA.n4810 GNDA.n4809 16.0005
R12498 GNDA.n4813 GNDA.n4810 16.0005
R12499 GNDA.n4814 GNDA.n4813 16.0005
R12500 GNDA.n4817 GNDA.n4814 16.0005
R12501 GNDA.n4818 GNDA.n4817 16.0005
R12502 GNDA.n4821 GNDA.n4818 16.0005
R12503 GNDA.n4822 GNDA.n4821 16.0005
R12504 GNDA.n4822 GNDA.n4720 16.0005
R12505 GNDA.n4806 GNDA.n4805 16.0005
R12506 GNDA.n4805 GNDA.n4802 16.0005
R12507 GNDA.n4802 GNDA.n4801 16.0005
R12508 GNDA.n4801 GNDA.n4798 16.0005
R12509 GNDA.n4798 GNDA.n4797 16.0005
R12510 GNDA.n4797 GNDA.n4794 16.0005
R12511 GNDA.n4794 GNDA.n4793 16.0005
R12512 GNDA.n4793 GNDA.n4790 16.0005
R12513 GNDA.n4789 GNDA.n4786 16.0005
R12514 GNDA.n4786 GNDA.n4785 16.0005
R12515 GNDA.n4785 GNDA.n4782 16.0005
R12516 GNDA.n4782 GNDA.n4781 16.0005
R12517 GNDA.n4781 GNDA.n4778 16.0005
R12518 GNDA.n4778 GNDA.n4777 16.0005
R12519 GNDA.n4777 GNDA.n4774 16.0005
R12520 GNDA.n4774 GNDA.n4773 16.0005
R12521 GNDA.n1661 GNDA.n1660 16.0005
R12522 GNDA.n1664 GNDA.n1661 16.0005
R12523 GNDA.n1665 GNDA.n1664 16.0005
R12524 GNDA.n1668 GNDA.n1665 16.0005
R12525 GNDA.n1669 GNDA.n1668 16.0005
R12526 GNDA.n1672 GNDA.n1669 16.0005
R12527 GNDA.n1674 GNDA.n1672 16.0005
R12528 GNDA.n1675 GNDA.n1674 16.0005
R12529 GNDA.n1657 GNDA.n1656 16.0005
R12530 GNDA.n1656 GNDA.n1653 16.0005
R12531 GNDA.n1653 GNDA.n1652 16.0005
R12532 GNDA.n1652 GNDA.n1649 16.0005
R12533 GNDA.n1649 GNDA.n1648 16.0005
R12534 GNDA.n1648 GNDA.n1645 16.0005
R12535 GNDA.n1645 GNDA.n1644 16.0005
R12536 GNDA.n1644 GNDA.n1641 16.0005
R12537 GNDA.n1640 GNDA.n1637 16.0005
R12538 GNDA.n1637 GNDA.n1636 16.0005
R12539 GNDA.n1636 GNDA.n1633 16.0005
R12540 GNDA.n1633 GNDA.n1632 16.0005
R12541 GNDA.n1632 GNDA.n1629 16.0005
R12542 GNDA.n1629 GNDA.n1628 16.0005
R12543 GNDA.n1628 GNDA.n1625 16.0005
R12544 GNDA.n1625 GNDA.n1601 16.0005
R12545 GNDA.n4962 GNDA.n4949 16.0005
R12546 GNDA.n4962 GNDA.n4961 16.0005
R12547 GNDA.n4961 GNDA.n4960 16.0005
R12548 GNDA.n4960 GNDA.n4957 16.0005
R12549 GNDA.n4957 GNDA.n4956 16.0005
R12550 GNDA.n4956 GNDA.n4953 16.0005
R12551 GNDA.n4953 GNDA.n4952 16.0005
R12552 GNDA.n4952 GNDA.n4864 16.0005
R12553 GNDA.n4948 GNDA.n4946 16.0005
R12554 GNDA.n4946 GNDA.n4943 16.0005
R12555 GNDA.n4943 GNDA.n4942 16.0005
R12556 GNDA.n4942 GNDA.n4939 16.0005
R12557 GNDA.n4939 GNDA.n4938 16.0005
R12558 GNDA.n4938 GNDA.n4935 16.0005
R12559 GNDA.n4935 GNDA.n4934 16.0005
R12560 GNDA.n4934 GNDA.n4931 16.0005
R12561 GNDA.n4930 GNDA.n4927 16.0005
R12562 GNDA.n4927 GNDA.n4926 16.0005
R12563 GNDA.n4926 GNDA.n4923 16.0005
R12564 GNDA.n4923 GNDA.n4922 16.0005
R12565 GNDA.n4922 GNDA.n4919 16.0005
R12566 GNDA.n4919 GNDA.n4918 16.0005
R12567 GNDA.n4918 GNDA.n4915 16.0005
R12568 GNDA.n4915 GNDA.n4914 16.0005
R12569 GNDA.n5241 GNDA.n5228 16.0005
R12570 GNDA.n5241 GNDA.n5240 16.0005
R12571 GNDA.n5240 GNDA.n5239 16.0005
R12572 GNDA.n5239 GNDA.n5236 16.0005
R12573 GNDA.n5236 GNDA.n5235 16.0005
R12574 GNDA.n5235 GNDA.n5232 16.0005
R12575 GNDA.n5232 GNDA.n5231 16.0005
R12576 GNDA.n5231 GNDA.n57 16.0005
R12577 GNDA.n5227 GNDA.n5225 16.0005
R12578 GNDA.n5225 GNDA.n5222 16.0005
R12579 GNDA.n5222 GNDA.n5221 16.0005
R12580 GNDA.n5221 GNDA.n5218 16.0005
R12581 GNDA.n5218 GNDA.n5217 16.0005
R12582 GNDA.n5217 GNDA.n5214 16.0005
R12583 GNDA.n5214 GNDA.n5213 16.0005
R12584 GNDA.n5213 GNDA.n5210 16.0005
R12585 GNDA.n5209 GNDA.n5206 16.0005
R12586 GNDA.n5206 GNDA.n5205 16.0005
R12587 GNDA.n5205 GNDA.n5202 16.0005
R12588 GNDA.n5202 GNDA.n5201 16.0005
R12589 GNDA.n5201 GNDA.n5198 16.0005
R12590 GNDA.n5198 GNDA.n5197 16.0005
R12591 GNDA.n5197 GNDA.n5194 16.0005
R12592 GNDA.n5194 GNDA.n5193 16.0005
R12593 GNDA.n2888 GNDA.n2673 16.0005
R12594 GNDA.n2894 GNDA.n2673 16.0005
R12595 GNDA.n2895 GNDA.n2894 16.0005
R12596 GNDA.n2896 GNDA.n2895 16.0005
R12597 GNDA.n2896 GNDA.n2671 16.0005
R12598 GNDA.n2902 GNDA.n2671 16.0005
R12599 GNDA.n2903 GNDA.n2902 16.0005
R12600 GNDA.n2904 GNDA.n2903 16.0005
R12601 GNDA.n2887 GNDA.n2886 16.0005
R12602 GNDA.n2886 GNDA.n2675 16.0005
R12603 GNDA.n2880 GNDA.n2675 16.0005
R12604 GNDA.n2880 GNDA.n2879 16.0005
R12605 GNDA.n2879 GNDA.n2878 16.0005
R12606 GNDA.n2878 GNDA.n2677 16.0005
R12607 GNDA.n2872 GNDA.n2677 16.0005
R12608 GNDA.n2872 GNDA.n2871 16.0005
R12609 GNDA.n2870 GNDA.n2679 16.0005
R12610 GNDA.n2864 GNDA.n2679 16.0005
R12611 GNDA.n2864 GNDA.n2863 16.0005
R12612 GNDA.n2863 GNDA.n2862 16.0005
R12613 GNDA.n2862 GNDA.n2681 16.0005
R12614 GNDA.n2857 GNDA.n2681 16.0005
R12615 GNDA.n2857 GNDA.n2856 16.0005
R12616 GNDA.n2856 GNDA.n2855 16.0005
R12617 GNDA.n5148 GNDA.n5147 16.0005
R12618 GNDA.n5151 GNDA.n5148 16.0005
R12619 GNDA.n5152 GNDA.n5151 16.0005
R12620 GNDA.n5155 GNDA.n5152 16.0005
R12621 GNDA.n5156 GNDA.n5155 16.0005
R12622 GNDA.n5159 GNDA.n5156 16.0005
R12623 GNDA.n5161 GNDA.n5159 16.0005
R12624 GNDA.n5162 GNDA.n5161 16.0005
R12625 GNDA.n5144 GNDA.n5143 16.0005
R12626 GNDA.n5143 GNDA.n5140 16.0005
R12627 GNDA.n5140 GNDA.n5139 16.0005
R12628 GNDA.n5139 GNDA.n5136 16.0005
R12629 GNDA.n5136 GNDA.n5135 16.0005
R12630 GNDA.n5135 GNDA.n5132 16.0005
R12631 GNDA.n5132 GNDA.n5131 16.0005
R12632 GNDA.n5131 GNDA.n5128 16.0005
R12633 GNDA.n5127 GNDA.n5124 16.0005
R12634 GNDA.n5124 GNDA.n5123 16.0005
R12635 GNDA.n5123 GNDA.n5120 16.0005
R12636 GNDA.n5120 GNDA.n5119 16.0005
R12637 GNDA.n5119 GNDA.n5116 16.0005
R12638 GNDA.n5116 GNDA.n5115 16.0005
R12639 GNDA.n5115 GNDA.n5112 16.0005
R12640 GNDA.n5112 GNDA.n5111 16.0005
R12641 GNDA.n1466 GNDA.t48 15.3505
R12642 GNDA.t62 GNDA.t233 15.0244
R12643 GNDA.t62 GNDA.t253 15.0244
R12644 GNDA.n5260 GNDA.n26 14.555
R12645 GNDA.n4981 GNDA.n107 14.555
R12646 GNDA.t181 GNDA.t65 13.8109
R12647 GNDA.n2803 GNDA.n2718 12.8005
R12648 GNDA.n2807 GNDA.n2718 12.8005
R12649 GNDA.n2706 GNDA.n2705 12.8005
R12650 GNDA.n2710 GNDA.n2705 12.8005
R12651 GNDA.n4680 GNDA.n357 12.8005
R12652 GNDA.n4680 GNDA.n4679 12.8005
R12653 GNDA.n3384 GNDA.t116 12.6791
R12654 GNDA.n3381 GNDA.t105 12.6791
R12655 GNDA.n4611 GNDA.t134 12.6791
R12656 GNDA.n3850 GNDA.t144 12.6791
R12657 GNDA.n3937 GNDA.n3936 12.1358
R12658 GNDA.n895 GNDA.n803 12.1358
R12659 GNDA.n3940 GNDA.n3939 12.1114
R12660 GNDA.n892 GNDA.n889 12.1114
R12661 GNDA.t215 GNDA.n2844 12.0196
R12662 GNDA.n3302 GNDA.t235 12.0196
R12663 GNDA.n3129 GNDA.t247 12.0196
R12664 GNDA.t293 GNDA.t279 11.8285
R12665 GNDA.t277 GNDA.t208 11.8285
R12666 GNDA.t260 GNDA.t189 11.8285
R12667 GNDA.t242 GNDA.t231 11.8285
R12668 GNDA.n3196 GNDA.n3195 11.6369
R12669 GNDA.n3198 GNDA.n3196 11.6369
R12670 GNDA.n3198 GNDA.n3197 11.6369
R12671 GNDA.n3197 GNDA.n1540 11.6369
R12672 GNDA.n1540 GNDA.n1538 11.6369
R12673 GNDA.n3206 GNDA.n1538 11.6369
R12674 GNDA.n3207 GNDA.n3206 11.6369
R12675 GNDA.n3208 GNDA.n3207 11.6369
R12676 GNDA.n3208 GNDA.n1533 11.6369
R12677 GNDA.n3217 GNDA.n1533 11.6369
R12678 GNDA.n3173 GNDA.n3172 11.6369
R12679 GNDA.n3174 GNDA.n3173 11.6369
R12680 GNDA.n3174 GNDA.n1547 11.6369
R12681 GNDA.n3180 GNDA.n1547 11.6369
R12682 GNDA.n3181 GNDA.n3180 11.6369
R12683 GNDA.n3182 GNDA.n3181 11.6369
R12684 GNDA.n3182 GNDA.n1545 11.6369
R12685 GNDA.n3188 GNDA.n1545 11.6369
R12686 GNDA.n3189 GNDA.n3188 11.6369
R12687 GNDA.n3190 GNDA.n3189 11.6369
R12688 GNDA.n3190 GNDA.n1543 11.6369
R12689 GNDA.n3009 GNDA.n2983 11.6369
R12690 GNDA.n3009 GNDA.n3008 11.6369
R12691 GNDA.n3008 GNDA.n3007 11.6369
R12692 GNDA.n3007 GNDA.n2985 11.6369
R12693 GNDA.n3002 GNDA.n2985 11.6369
R12694 GNDA.n3002 GNDA.n3001 11.6369
R12695 GNDA.n3001 GNDA.n3000 11.6369
R12696 GNDA.n3000 GNDA.n2988 11.6369
R12697 GNDA.n2995 GNDA.n2988 11.6369
R12698 GNDA.n2995 GNDA.n2994 11.6369
R12699 GNDA.n2994 GNDA.n2993 11.6369
R12700 GNDA.n1593 GNDA.n1589 11.6369
R12701 GNDA.n1734 GNDA.n1593 11.6369
R12702 GNDA.n1734 GNDA.n1733 11.6369
R12703 GNDA.n1733 GNDA.n1732 11.6369
R12704 GNDA.n1732 GNDA.n1594 11.6369
R12705 GNDA.n1727 GNDA.n1594 11.6369
R12706 GNDA.n1727 GNDA.n1726 11.6369
R12707 GNDA.n1726 GNDA.n1725 11.6369
R12708 GNDA.n1725 GNDA.n1596 11.6369
R12709 GNDA.n1719 GNDA.n1596 11.6369
R12710 GNDA.n1762 GNDA.n1761 11.6369
R12711 GNDA.n1761 GNDA.n1758 11.6369
R12712 GNDA.n1758 GNDA.n1757 11.6369
R12713 GNDA.n1757 GNDA.n1754 11.6369
R12714 GNDA.n1754 GNDA.n1753 11.6369
R12715 GNDA.n1753 GNDA.n1750 11.6369
R12716 GNDA.n1750 GNDA.n1749 11.6369
R12717 GNDA.n1749 GNDA.n1746 11.6369
R12718 GNDA.n1746 GNDA.n1745 11.6369
R12719 GNDA.n1745 GNDA.n1742 11.6369
R12720 GNDA.n1742 GNDA.n1741 11.6369
R12721 GNDA.n1565 GNDA.n132 11.6369
R12722 GNDA.n1568 GNDA.n1565 11.6369
R12723 GNDA.n1569 GNDA.n1568 11.6369
R12724 GNDA.n1572 GNDA.n1569 11.6369
R12725 GNDA.n1573 GNDA.n1572 11.6369
R12726 GNDA.n1576 GNDA.n1573 11.6369
R12727 GNDA.n1577 GNDA.n1576 11.6369
R12728 GNDA.n1580 GNDA.n1577 11.6369
R12729 GNDA.n1581 GNDA.n1580 11.6369
R12730 GNDA.n1584 GNDA.n1581 11.6369
R12731 GNDA.n1587 GNDA.n1584 11.6369
R12732 GNDA.n263 GNDA.n262 11.6369
R12733 GNDA.n266 GNDA.n263 11.6369
R12734 GNDA.n267 GNDA.n266 11.6369
R12735 GNDA.n270 GNDA.n267 11.6369
R12736 GNDA.n271 GNDA.n270 11.6369
R12737 GNDA.n274 GNDA.n271 11.6369
R12738 GNDA.n275 GNDA.n274 11.6369
R12739 GNDA.n277 GNDA.n275 11.6369
R12740 GNDA.n277 GNDA.n276 11.6369
R12741 GNDA.n276 GNDA.n228 11.6369
R12742 GNDA.n259 GNDA.n258 11.6369
R12743 GNDA.n258 GNDA.n255 11.6369
R12744 GNDA.n255 GNDA.n254 11.6369
R12745 GNDA.n254 GNDA.n251 11.6369
R12746 GNDA.n251 GNDA.n250 11.6369
R12747 GNDA.n250 GNDA.n247 11.6369
R12748 GNDA.n247 GNDA.n246 11.6369
R12749 GNDA.n246 GNDA.n243 11.6369
R12750 GNDA.n243 GNDA.n242 11.6369
R12751 GNDA.n242 GNDA.n131 11.6369
R12752 GNDA.n5077 GNDA.n131 11.6369
R12753 GNDA.n4857 GNDA.n4856 11.6369
R12754 GNDA.n4856 GNDA.n4855 11.6369
R12755 GNDA.n4855 GNDA.n4854 11.6369
R12756 GNDA.n4854 GNDA.n4852 11.6369
R12757 GNDA.n4852 GNDA.n4849 11.6369
R12758 GNDA.n4849 GNDA.n4848 11.6369
R12759 GNDA.n4848 GNDA.n4845 11.6369
R12760 GNDA.n4845 GNDA.n4844 11.6369
R12761 GNDA.n4844 GNDA.n4841 11.6369
R12762 GNDA.n4841 GNDA.n4840 11.6369
R12763 GNDA.n4719 GNDA.n4718 11.6369
R12764 GNDA.n4718 GNDA.n290 11.6369
R12765 GNDA.n4712 GNDA.n290 11.6369
R12766 GNDA.n4712 GNDA.n4711 11.6369
R12767 GNDA.n4711 GNDA.n4710 11.6369
R12768 GNDA.n4710 GNDA.n294 11.6369
R12769 GNDA.n4704 GNDA.n294 11.6369
R12770 GNDA.n4704 GNDA.n4703 11.6369
R12771 GNDA.n4703 GNDA.n4702 11.6369
R12772 GNDA.n4702 GNDA.n298 11.6369
R12773 GNDA.n4696 GNDA.n298 11.6369
R12774 GNDA.n2957 GNDA.n2956 11.6369
R12775 GNDA.n2956 GNDA.n2953 11.6369
R12776 GNDA.n2953 GNDA.n2952 11.6369
R12777 GNDA.n2952 GNDA.n2949 11.6369
R12778 GNDA.n2949 GNDA.n2948 11.6369
R12779 GNDA.n2948 GNDA.n2945 11.6369
R12780 GNDA.n2945 GNDA.n2944 11.6369
R12781 GNDA.n2944 GNDA.n2941 11.6369
R12782 GNDA.n2941 GNDA.n2940 11.6369
R12783 GNDA.n2940 GNDA.n2937 11.6369
R12784 GNDA.n2958 GNDA.n1854 11.6369
R12785 GNDA.n2964 GNDA.n1854 11.6369
R12786 GNDA.n2965 GNDA.n2964 11.6369
R12787 GNDA.n2966 GNDA.n2965 11.6369
R12788 GNDA.n2966 GNDA.n1852 11.6369
R12789 GNDA.n2972 GNDA.n1852 11.6369
R12790 GNDA.n2973 GNDA.n2972 11.6369
R12791 GNDA.n2974 GNDA.n2973 11.6369
R12792 GNDA.n2974 GNDA.n1850 11.6369
R12793 GNDA.n2980 GNDA.n1850 11.6369
R12794 GNDA.n2981 GNDA.n2980 11.6369
R12795 GNDA.n4638 GNDA.n4637 11.6369
R12796 GNDA.n4637 GNDA.n4636 11.6369
R12797 GNDA.n4636 GNDA.n426 11.6369
R12798 GNDA.n4630 GNDA.n426 11.6369
R12799 GNDA.n4630 GNDA.n4629 11.6369
R12800 GNDA.n4629 GNDA.n92 11.6369
R12801 GNDA.n5084 GNDA.n92 11.6369
R12802 GNDA.n5085 GNDA.n5084 11.6369
R12803 GNDA.n5087 GNDA.n5085 11.6369
R12804 GNDA.n5087 GNDA.n5086 11.6369
R12805 GNDA.n4662 GNDA.n4661 11.6369
R12806 GNDA.n4661 GNDA.n4660 11.6369
R12807 GNDA.n4660 GNDA.n414 11.6369
R12808 GNDA.n4654 GNDA.n414 11.6369
R12809 GNDA.n4654 GNDA.n4653 11.6369
R12810 GNDA.n4653 GNDA.n4652 11.6369
R12811 GNDA.n4652 GNDA.n418 11.6369
R12812 GNDA.n4646 GNDA.n418 11.6369
R12813 GNDA.n4646 GNDA.n4645 11.6369
R12814 GNDA.n4645 GNDA.n4644 11.6369
R12815 GNDA.n4644 GNDA.n422 11.6369
R12816 GNDA.n4694 GNDA.n303 11.6369
R12817 GNDA.n4688 GNDA.n303 11.6369
R12818 GNDA.n4688 GNDA.n4687 11.6369
R12819 GNDA.n4687 GNDA.n4686 11.6369
R12820 GNDA.n4686 GNDA.n353 11.6369
R12821 GNDA.n4677 GNDA.n360 11.6369
R12822 GNDA.n364 GNDA.n360 11.6369
R12823 GNDA.n4670 GNDA.n364 11.6369
R12824 GNDA.n4670 GNDA.n4669 11.6369
R12825 GNDA.n4669 GNDA.n4668 11.6369
R12826 GNDA.t303 GNDA.t213 11.4882
R12827 GNDA.n572 GNDA.n433 11.4533
R12828 GNDA.n3326 GNDA.n586 11.4533
R12829 GNDA.t62 GNDA.n99 11.3072
R12830 GNDA.n4626 GNDA.t179 11.2482
R12831 GNDA.n3607 GNDA.n3606 11.245
R12832 GNDA.n3338 GNDA.n3337 11.245
R12833 GNDA.t307 GNDA.t77 11.2059
R12834 GNDA.t206 GNDA.t27 11.2059
R12835 GNDA.t193 GNDA.t32 11.2059
R12836 GNDA.t21 GNDA.t24 11.2059
R12837 GNDA.t130 GNDA.t28 11.2059
R12838 GNDA.n3267 GNDA.n3266 10.9846
R12839 GNDA.n2659 GNDA.n2658 10.87
R12840 GNDA.n2929 GNDA.n2928 10.87
R12841 GNDA.n2927 GNDA.n2920 10.87
R12842 GNDA.n2734 GNDA.n1498 10.87
R12843 GNDA.n3275 GNDA.n3274 10.87
R12844 GNDA.n3271 GNDA.n1501 10.87
R12845 GNDA.n3270 GNDA.n1502 10.87
R12846 GNDA.t43 GNDA.t167 9.90372
R12847 GNDA.t48 GNDA.t240 9.90372
R12848 GNDA.n2656 GNDA.t182 9.66779
R12849 GNDA.n3363 GNDA.t12 9.6005
R12850 GNDA.n3363 GNDA.t171 9.6005
R12851 GNDA.n3361 GNDA.t164 9.6005
R12852 GNDA.n3361 GNDA.t285 9.6005
R12853 GNDA.n3359 GNDA.t299 9.6005
R12854 GNDA.n3359 GNDA.t6 9.6005
R12855 GNDA.n3357 GNDA.t218 9.6005
R12856 GNDA.n3357 GNDA.t186 9.6005
R12857 GNDA.n3355 GNDA.t199 9.6005
R12858 GNDA.n3355 GNDA.t42 9.6005
R12859 GNDA.n3353 GNDA.t246 9.6005
R12860 GNDA.n3353 GNDA.t276 9.6005
R12861 GNDA.n3351 GNDA.t52 9.6005
R12862 GNDA.n3351 GNDA.t4 9.6005
R12863 GNDA.n3349 GNDA.t50 9.6005
R12864 GNDA.n3349 GNDA.t259 9.6005
R12865 GNDA.n3347 GNDA.t2 9.6005
R12866 GNDA.n3347 GNDA.t8 9.6005
R12867 GNDA.n3345 GNDA.t250 9.6005
R12868 GNDA.n3345 GNDA.t162 9.6005
R12869 GNDA.n3343 GNDA.t287 9.6005
R12870 GNDA.n3343 GNDA.t121 9.6005
R12871 GNDA.n581 GNDA.t36 9.6005
R12872 GNDA.n581 GNDA.t290 9.6005
R12873 GNDA.n3242 GNDA.t265 9.6005
R12874 GNDA.n3245 GNDA.t271 9.6005
R12875 GNDA.n2815 GNDA.t273 9.6005
R12876 GNDA.n2824 GNDA.t275 9.6005
R12877 GNDA.t174 GNDA.t301 9.46287
R12878 GNDA.t190 GNDA.t302 9.46287
R12879 GNDA.n2803 GNDA.n2716 9.36264
R12880 GNDA.n2706 GNDA.n2703 9.36264
R12881 GNDA.n2625 GNDA.n357 9.36264
R12882 GNDA.n3341 GNDA.t34 9.33836
R12883 GNDA.n3571 GNDA.t185 9.33836
R12884 GNDA.n3611 GNDA.t33 9.33836
R12885 GNDA.n2718 GNDA.n2717 9.3005
R12886 GNDA.n2808 GNDA.n2807 9.3005
R12887 GNDA.n2705 GNDA.n2704 9.3005
R12888 GNDA.n2711 GNDA.n2710 9.3005
R12889 GNDA.n4680 GNDA.n358 9.3005
R12890 GNDA.n4679 GNDA.n359 9.3005
R12891 GNDA.n3227 GNDA.n3226 8.62751
R12892 GNDA.n5167 GNDA.n26 8.60107
R12893 GNDA.n161 GNDA.n107 8.60107
R12894 GNDA.n2933 GNDA.t108 8.01325
R12895 GNDA.n2843 GNDA.t168 8.01325
R12896 GNDA.t197 GNDA.n3279 8.01325
R12897 GNDA.n3130 GNDA.t46 8.01325
R12898 GNDA.n3571 GNDA.t229 7.47079
R12899 GNDA.t51 GNDA.t95 7.47079
R12900 GNDA.t3 GNDA.t307 7.47079
R12901 GNDA.t49 GNDA.t206 7.47079
R12902 GNDA.t258 GNDA.t193 7.47079
R12903 GNDA.t1 GNDA.t21 7.47079
R12904 GNDA.t7 GNDA.t130 7.47079
R12905 GNDA.n2917 GNDA.t255 7.01165
R12906 GNDA.n2847 GNDA.t15 7.01165
R12907 GNDA.n2801 GNDA.n2799 7.01165
R12908 GNDA.n3264 GNDA.n1506 7.01165
R12909 GNDA.n2993 GNDA.n1800 6.72373
R12910 GNDA.n1588 GNDA.n1587 6.72373
R12911 GNDA.n5077 GNDA.n5076 6.72373
R12912 GNDA.n4696 GNDA.n4695 6.72373
R12913 GNDA.n2982 GNDA.n2981 6.72373
R12914 GNDA.n4668 GNDA.n365 6.72373
R12915 GNDA.n4627 GNDA.n4626 6.69811
R12916 GNDA.n3172 GNDA.n1800 6.20656
R12917 GNDA.n2983 GNDA.n2982 6.20656
R12918 GNDA.n1762 GNDA.n1588 6.20656
R12919 GNDA.n5076 GNDA.n132 6.20656
R12920 GNDA.n4662 GNDA.n365 6.20656
R12921 GNDA.n4695 GNDA.n4694 6.20656
R12922 GNDA.n4678 GNDA.n353 6.07727
R12923 GNDA.t62 GNDA.t165 6.01006
R12924 GNDA.n2825 GNDA.n2816 5.81868
R12925 GNDA.n2823 GNDA.n2816 5.81868
R12926 GNDA.n4678 GNDA.n4677 5.5601
R12927 GNDA.n3062 GNDA.n1531 5.51161
R12928 GNDA.n2796 GNDA.n2794 5.51161
R12929 GNDA.n4988 GNDA.n186 5.51161
R12930 GNDA.n4773 GNDA.n4743 5.51161
R12931 GNDA.n1713 GNDA.n1601 5.51161
R12932 GNDA.n4914 GNDA.n4892 5.51161
R12933 GNDA.n5193 GNDA.n5171 5.51161
R12934 GNDA.n2855 GNDA.n2684 5.51161
R12935 GNDA.n5111 GNDA.n5097 5.51161
R12936 GNDA.n3219 GNDA.n3218 5.1717
R12937 GNDA.n1718 GNDA.n1714 5.1717
R12938 GNDA.n5096 GNDA.n87 5.1717
R12939 GNDA.n3365 GNDA.n3364 5.063
R12940 GNDA.t209 GNDA.t159 5.00847
R12941 GNDA.n2827 GNDA.t233 5.00847
R12942 GNDA.t62 GNDA.t71 5.00847
R12943 GNDA.t62 GNDA.t92 5.00847
R12944 GNDA.t253 GNDA.n3248 5.00847
R12945 GNDA.t228 GNDA.t156 5.00847
R12946 GNDA.n4978 GNDA.n4863 4.9157
R12947 GNDA.n4837 GNDA.n4834 4.9157
R12948 GNDA.n2936 GNDA.n2935 4.9157
R12949 GNDA.n3344 GNDA.n568 4.71925
R12950 GNDA.n466 GNDA.n465 4.5005
R12951 GNDA.n3597 GNDA.n3596 4.5005
R12952 GNDA.n3600 GNDA.n576 4.5005
R12953 GNDA.n3592 GNDA.n3588 4.5005
R12954 GNDA.n3593 GNDA.n580 4.5005
R12955 GNDA.n3593 GNDA.n3592 4.5005
R12956 GNDA.n591 GNDA.n590 4.5005
R12957 GNDA.n3334 GNDA.n596 4.5005
R12958 GNDA.n3331 GNDA.n596 4.5005
R12959 GNDA.n3332 GNDA.n3331 4.5005
R12960 GNDA.n3558 GNDA.n593 4.5005
R12961 GNDA.n3560 GNDA.n3559 4.5005
R12962 GNDA.n3559 GNDA.n3558 4.5005
R12963 GNDA.n599 GNDA.n598 4.5005
R12964 GNDA.n3536 GNDA.n601 4.5005
R12965 GNDA.n3538 GNDA.n3537 4.5005
R12966 GNDA.n3537 GNDA.n3536 4.5005
R12967 GNDA.n449 GNDA.n434 4.5005
R12968 GNDA.n473 GNDA.n472 4.5005
R12969 GNDA.n473 GNDA.n434 4.5005
R12970 GNDA.n2712 GNDA.n2711 4.5005
R12971 GNDA.n2809 GNDA.n2808 4.5005
R12972 GNDA.n2702 GNDA.n2701 4.5005
R12973 GNDA.n2814 GNDA.n2695 4.5005
R12974 GNDA.n2813 GNDA.n1524 4.5005
R12975 GNDA.n2814 GNDA.n2813 4.5005
R12976 GNDA.n2583 GNDA.n2577 4.5005
R12977 GNDA.n2585 GNDA.n2584 4.5005
R12978 GNDA.n2586 GNDA.n2576 4.5005
R12979 GNDA.n2590 GNDA.n2589 4.5005
R12980 GNDA.n2591 GNDA.n2573 4.5005
R12981 GNDA.n2593 GNDA.n2592 4.5005
R12982 GNDA.n2594 GNDA.n2572 4.5005
R12983 GNDA.n2598 GNDA.n2597 4.5005
R12984 GNDA.n2599 GNDA.n2569 4.5005
R12985 GNDA.n2601 GNDA.n2600 4.5005
R12986 GNDA.n2602 GNDA.n2568 4.5005
R12987 GNDA.n2606 GNDA.n2605 4.5005
R12988 GNDA.n2607 GNDA.n2565 4.5005
R12989 GNDA.n2609 GNDA.n2608 4.5005
R12990 GNDA.n2610 GNDA.n2564 4.5005
R12991 GNDA.n2614 GNDA.n2613 4.5005
R12992 GNDA.n2615 GNDA.n2561 4.5005
R12993 GNDA.n2617 GNDA.n2616 4.5005
R12994 GNDA.n2618 GNDA.n2560 4.5005
R12995 GNDA.n2622 GNDA.n2621 4.5005
R12996 GNDA.n2623 GNDA.n2559 4.5005
R12997 GNDA.n2637 GNDA.n2636 4.5005
R12998 GNDA.n3228 GNDA.n1526 4.5005
R12999 GNDA.n2630 GNDA.n2629 4.5005
R13000 GNDA.n2633 GNDA.n1527 4.5005
R13001 GNDA.n2629 GNDA.n1527 4.5005
R13002 GNDA.n2626 GNDA.n359 4.5005
R13003 GNDA.n3697 GNDA.n3696 4.5005
R13004 GNDA.n3618 GNDA.n3617 4.5005
R13005 GNDA.n3640 GNDA.n3619 4.5005
R13006 GNDA.n3641 GNDA.n3620 4.5005
R13007 GNDA.n3642 GNDA.n3621 4.5005
R13008 GNDA.n3643 GNDA.n3622 4.5005
R13009 GNDA.n3644 GNDA.n3623 4.5005
R13010 GNDA.n3645 GNDA.n3624 4.5005
R13011 GNDA.n3646 GNDA.n3625 4.5005
R13012 GNDA.n3647 GNDA.n3626 4.5005
R13013 GNDA.n3648 GNDA.n3627 4.5005
R13014 GNDA.n3649 GNDA.n3628 4.5005
R13015 GNDA.n3650 GNDA.n3629 4.5005
R13016 GNDA.n3651 GNDA.n3630 4.5005
R13017 GNDA.n3652 GNDA.n3631 4.5005
R13018 GNDA.n3653 GNDA.n3632 4.5005
R13019 GNDA.n3654 GNDA.n3633 4.5005
R13020 GNDA.n3655 GNDA.n3634 4.5005
R13021 GNDA.n3656 GNDA.n3635 4.5005
R13022 GNDA.n3657 GNDA.n3636 4.5005
R13023 GNDA.n3658 GNDA.n3637 4.5005
R13024 GNDA.n3659 GNDA.n3638 4.5005
R13025 GNDA.n4573 GNDA.n4572 4.5005
R13026 GNDA.n500 GNDA.n499 4.5005
R13027 GNDA.n4518 GNDA.n4517 4.5005
R13028 GNDA.n4522 GNDA.n4519 4.5005
R13029 GNDA.n4523 GNDA.n4516 4.5005
R13030 GNDA.n4527 GNDA.n4526 4.5005
R13031 GNDA.n4528 GNDA.n4515 4.5005
R13032 GNDA.n4532 GNDA.n4529 4.5005
R13033 GNDA.n4533 GNDA.n4514 4.5005
R13034 GNDA.n4537 GNDA.n4536 4.5005
R13035 GNDA.n4538 GNDA.n4513 4.5005
R13036 GNDA.n4542 GNDA.n4539 4.5005
R13037 GNDA.n4543 GNDA.n4512 4.5005
R13038 GNDA.n4547 GNDA.n4546 4.5005
R13039 GNDA.n4548 GNDA.n4511 4.5005
R13040 GNDA.n4552 GNDA.n4549 4.5005
R13041 GNDA.n4553 GNDA.n4510 4.5005
R13042 GNDA.n4557 GNDA.n4556 4.5005
R13043 GNDA.n4558 GNDA.n4509 4.5005
R13044 GNDA.n4562 GNDA.n4559 4.5005
R13045 GNDA.n4563 GNDA.n4508 4.5005
R13046 GNDA.n4567 GNDA.n4566 4.5005
R13047 GNDA.n4438 GNDA.n4437 4.5005
R13048 GNDA.n4441 GNDA.n4440 4.5005
R13049 GNDA.n4442 GNDA.n4436 4.5005
R13050 GNDA.n4446 GNDA.n4443 4.5005
R13051 GNDA.n4447 GNDA.n4435 4.5005
R13052 GNDA.n4451 GNDA.n4450 4.5005
R13053 GNDA.n4452 GNDA.n4434 4.5005
R13054 GNDA.n4456 GNDA.n4453 4.5005
R13055 GNDA.n4457 GNDA.n4433 4.5005
R13056 GNDA.n4461 GNDA.n4460 4.5005
R13057 GNDA.n4462 GNDA.n4432 4.5005
R13058 GNDA.n4466 GNDA.n4463 4.5005
R13059 GNDA.n4467 GNDA.n4431 4.5005
R13060 GNDA.n4471 GNDA.n4470 4.5005
R13061 GNDA.n4472 GNDA.n4430 4.5005
R13062 GNDA.n4476 GNDA.n4473 4.5005
R13063 GNDA.n4477 GNDA.n4429 4.5005
R13064 GNDA.n4481 GNDA.n4480 4.5005
R13065 GNDA.n4482 GNDA.n4428 4.5005
R13066 GNDA.n4486 GNDA.n4483 4.5005
R13067 GNDA.n4487 GNDA.n4427 4.5005
R13068 GNDA.n4491 GNDA.n4490 4.5005
R13069 GNDA.n4356 GNDA.n4355 4.5005
R13070 GNDA.n4359 GNDA.n4358 4.5005
R13071 GNDA.n4360 GNDA.n4354 4.5005
R13072 GNDA.n4364 GNDA.n4361 4.5005
R13073 GNDA.n4365 GNDA.n4353 4.5005
R13074 GNDA.n4369 GNDA.n4368 4.5005
R13075 GNDA.n4370 GNDA.n4352 4.5005
R13076 GNDA.n4374 GNDA.n4371 4.5005
R13077 GNDA.n4375 GNDA.n4351 4.5005
R13078 GNDA.n4379 GNDA.n4378 4.5005
R13079 GNDA.n4380 GNDA.n4350 4.5005
R13080 GNDA.n4384 GNDA.n4381 4.5005
R13081 GNDA.n4385 GNDA.n4349 4.5005
R13082 GNDA.n4389 GNDA.n4388 4.5005
R13083 GNDA.n4390 GNDA.n4348 4.5005
R13084 GNDA.n4394 GNDA.n4391 4.5005
R13085 GNDA.n4395 GNDA.n4347 4.5005
R13086 GNDA.n4399 GNDA.n4398 4.5005
R13087 GNDA.n4400 GNDA.n4346 4.5005
R13088 GNDA.n4404 GNDA.n4401 4.5005
R13089 GNDA.n4405 GNDA.n4345 4.5005
R13090 GNDA.n4409 GNDA.n4408 4.5005
R13091 GNDA.n4274 GNDA.n4273 4.5005
R13092 GNDA.n4277 GNDA.n4276 4.5005
R13093 GNDA.n4278 GNDA.n4272 4.5005
R13094 GNDA.n4282 GNDA.n4279 4.5005
R13095 GNDA.n4283 GNDA.n4271 4.5005
R13096 GNDA.n4287 GNDA.n4286 4.5005
R13097 GNDA.n4288 GNDA.n4270 4.5005
R13098 GNDA.n4292 GNDA.n4289 4.5005
R13099 GNDA.n4293 GNDA.n4269 4.5005
R13100 GNDA.n4297 GNDA.n4296 4.5005
R13101 GNDA.n4298 GNDA.n4268 4.5005
R13102 GNDA.n4302 GNDA.n4299 4.5005
R13103 GNDA.n4303 GNDA.n4267 4.5005
R13104 GNDA.n4307 GNDA.n4306 4.5005
R13105 GNDA.n4308 GNDA.n4266 4.5005
R13106 GNDA.n4312 GNDA.n4309 4.5005
R13107 GNDA.n4313 GNDA.n4265 4.5005
R13108 GNDA.n4317 GNDA.n4316 4.5005
R13109 GNDA.n4318 GNDA.n4264 4.5005
R13110 GNDA.n4322 GNDA.n4319 4.5005
R13111 GNDA.n4323 GNDA.n4263 4.5005
R13112 GNDA.n4327 GNDA.n4326 4.5005
R13113 GNDA.n4192 GNDA.n4191 4.5005
R13114 GNDA.n4195 GNDA.n4194 4.5005
R13115 GNDA.n4196 GNDA.n4190 4.5005
R13116 GNDA.n4200 GNDA.n4197 4.5005
R13117 GNDA.n4201 GNDA.n4189 4.5005
R13118 GNDA.n4205 GNDA.n4204 4.5005
R13119 GNDA.n4206 GNDA.n4188 4.5005
R13120 GNDA.n4210 GNDA.n4207 4.5005
R13121 GNDA.n4211 GNDA.n4187 4.5005
R13122 GNDA.n4215 GNDA.n4214 4.5005
R13123 GNDA.n4216 GNDA.n4186 4.5005
R13124 GNDA.n4220 GNDA.n4217 4.5005
R13125 GNDA.n4221 GNDA.n4185 4.5005
R13126 GNDA.n4225 GNDA.n4224 4.5005
R13127 GNDA.n4226 GNDA.n4184 4.5005
R13128 GNDA.n4230 GNDA.n4227 4.5005
R13129 GNDA.n4231 GNDA.n4183 4.5005
R13130 GNDA.n4235 GNDA.n4234 4.5005
R13131 GNDA.n4236 GNDA.n4182 4.5005
R13132 GNDA.n4240 GNDA.n4237 4.5005
R13133 GNDA.n4241 GNDA.n4181 4.5005
R13134 GNDA.n4245 GNDA.n4244 4.5005
R13135 GNDA.n3946 GNDA.n3945 4.5005
R13136 GNDA.n3949 GNDA.n3948 4.5005
R13137 GNDA.n3950 GNDA.n526 4.5005
R13138 GNDA.n3954 GNDA.n3951 4.5005
R13139 GNDA.n3955 GNDA.n525 4.5005
R13140 GNDA.n3959 GNDA.n3958 4.5005
R13141 GNDA.n3960 GNDA.n524 4.5005
R13142 GNDA.n3964 GNDA.n3961 4.5005
R13143 GNDA.n3965 GNDA.n523 4.5005
R13144 GNDA.n3969 GNDA.n3968 4.5005
R13145 GNDA.n3970 GNDA.n522 4.5005
R13146 GNDA.n3974 GNDA.n3971 4.5005
R13147 GNDA.n3975 GNDA.n521 4.5005
R13148 GNDA.n3979 GNDA.n3978 4.5005
R13149 GNDA.n3980 GNDA.n520 4.5005
R13150 GNDA.n3984 GNDA.n3981 4.5005
R13151 GNDA.n3985 GNDA.n519 4.5005
R13152 GNDA.n3989 GNDA.n3988 4.5005
R13153 GNDA.n3990 GNDA.n518 4.5005
R13154 GNDA.n3994 GNDA.n3991 4.5005
R13155 GNDA.n3995 GNDA.n517 4.5005
R13156 GNDA.n3999 GNDA.n3998 4.5005
R13157 GNDA.n4110 GNDA.n4109 4.5005
R13158 GNDA.n4113 GNDA.n4112 4.5005
R13159 GNDA.n4114 GNDA.n4108 4.5005
R13160 GNDA.n4118 GNDA.n4115 4.5005
R13161 GNDA.n4119 GNDA.n4107 4.5005
R13162 GNDA.n4123 GNDA.n4122 4.5005
R13163 GNDA.n4124 GNDA.n4106 4.5005
R13164 GNDA.n4128 GNDA.n4125 4.5005
R13165 GNDA.n4129 GNDA.n4105 4.5005
R13166 GNDA.n4133 GNDA.n4132 4.5005
R13167 GNDA.n4134 GNDA.n4104 4.5005
R13168 GNDA.n4138 GNDA.n4135 4.5005
R13169 GNDA.n4139 GNDA.n4103 4.5005
R13170 GNDA.n4143 GNDA.n4142 4.5005
R13171 GNDA.n4144 GNDA.n4102 4.5005
R13172 GNDA.n4148 GNDA.n4145 4.5005
R13173 GNDA.n4149 GNDA.n4101 4.5005
R13174 GNDA.n4153 GNDA.n4152 4.5005
R13175 GNDA.n4154 GNDA.n4100 4.5005
R13176 GNDA.n4158 GNDA.n4155 4.5005
R13177 GNDA.n4159 GNDA.n4099 4.5005
R13178 GNDA.n4163 GNDA.n4162 4.5005
R13179 GNDA.n4028 GNDA.n4027 4.5005
R13180 GNDA.n4031 GNDA.n4030 4.5005
R13181 GNDA.n4032 GNDA.n4026 4.5005
R13182 GNDA.n4036 GNDA.n4033 4.5005
R13183 GNDA.n4037 GNDA.n4025 4.5005
R13184 GNDA.n4041 GNDA.n4040 4.5005
R13185 GNDA.n4042 GNDA.n4024 4.5005
R13186 GNDA.n4046 GNDA.n4043 4.5005
R13187 GNDA.n4047 GNDA.n4023 4.5005
R13188 GNDA.n4051 GNDA.n4050 4.5005
R13189 GNDA.n4052 GNDA.n4022 4.5005
R13190 GNDA.n4056 GNDA.n4053 4.5005
R13191 GNDA.n4057 GNDA.n4021 4.5005
R13192 GNDA.n4061 GNDA.n4060 4.5005
R13193 GNDA.n4062 GNDA.n4020 4.5005
R13194 GNDA.n4066 GNDA.n4063 4.5005
R13195 GNDA.n4067 GNDA.n4019 4.5005
R13196 GNDA.n4071 GNDA.n4070 4.5005
R13197 GNDA.n4072 GNDA.n4018 4.5005
R13198 GNDA.n4076 GNDA.n4073 4.5005
R13199 GNDA.n4077 GNDA.n4017 4.5005
R13200 GNDA.n4081 GNDA.n4080 4.5005
R13201 GNDA.n3934 GNDA.n3933 4.5005
R13202 GNDA.n3855 GNDA.n3854 4.5005
R13203 GNDA.n3877 GNDA.n3856 4.5005
R13204 GNDA.n3878 GNDA.n3857 4.5005
R13205 GNDA.n3879 GNDA.n3858 4.5005
R13206 GNDA.n3880 GNDA.n3859 4.5005
R13207 GNDA.n3881 GNDA.n3860 4.5005
R13208 GNDA.n3882 GNDA.n3861 4.5005
R13209 GNDA.n3883 GNDA.n3862 4.5005
R13210 GNDA.n3884 GNDA.n3863 4.5005
R13211 GNDA.n3885 GNDA.n3864 4.5005
R13212 GNDA.n3886 GNDA.n3865 4.5005
R13213 GNDA.n3887 GNDA.n3866 4.5005
R13214 GNDA.n3888 GNDA.n3867 4.5005
R13215 GNDA.n3889 GNDA.n3868 4.5005
R13216 GNDA.n3890 GNDA.n3869 4.5005
R13217 GNDA.n3891 GNDA.n3870 4.5005
R13218 GNDA.n3892 GNDA.n3871 4.5005
R13219 GNDA.n3893 GNDA.n3872 4.5005
R13220 GNDA.n3894 GNDA.n3873 4.5005
R13221 GNDA.n3895 GNDA.n3874 4.5005
R13222 GNDA.n3896 GNDA.n3875 4.5005
R13223 GNDA.n3844 GNDA.n3843 4.5005
R13224 GNDA.n536 GNDA.n535 4.5005
R13225 GNDA.n3789 GNDA.n3788 4.5005
R13226 GNDA.n3793 GNDA.n3790 4.5005
R13227 GNDA.n3794 GNDA.n3787 4.5005
R13228 GNDA.n3798 GNDA.n3797 4.5005
R13229 GNDA.n3799 GNDA.n3786 4.5005
R13230 GNDA.n3803 GNDA.n3800 4.5005
R13231 GNDA.n3804 GNDA.n3785 4.5005
R13232 GNDA.n3808 GNDA.n3807 4.5005
R13233 GNDA.n3809 GNDA.n3784 4.5005
R13234 GNDA.n3813 GNDA.n3810 4.5005
R13235 GNDA.n3814 GNDA.n3783 4.5005
R13236 GNDA.n3818 GNDA.n3817 4.5005
R13237 GNDA.n3819 GNDA.n3782 4.5005
R13238 GNDA.n3823 GNDA.n3820 4.5005
R13239 GNDA.n3824 GNDA.n3781 4.5005
R13240 GNDA.n3828 GNDA.n3827 4.5005
R13241 GNDA.n3829 GNDA.n3780 4.5005
R13242 GNDA.n3833 GNDA.n3830 4.5005
R13243 GNDA.n3834 GNDA.n3779 4.5005
R13244 GNDA.n3838 GNDA.n3837 4.5005
R13245 GNDA.n3709 GNDA.n3708 4.5005
R13246 GNDA.n3712 GNDA.n3711 4.5005
R13247 GNDA.n3713 GNDA.n562 4.5005
R13248 GNDA.n3717 GNDA.n3714 4.5005
R13249 GNDA.n3718 GNDA.n561 4.5005
R13250 GNDA.n3722 GNDA.n3721 4.5005
R13251 GNDA.n3723 GNDA.n560 4.5005
R13252 GNDA.n3727 GNDA.n3724 4.5005
R13253 GNDA.n3728 GNDA.n559 4.5005
R13254 GNDA.n3732 GNDA.n3731 4.5005
R13255 GNDA.n3733 GNDA.n558 4.5005
R13256 GNDA.n3737 GNDA.n3734 4.5005
R13257 GNDA.n3738 GNDA.n557 4.5005
R13258 GNDA.n3742 GNDA.n3741 4.5005
R13259 GNDA.n3743 GNDA.n556 4.5005
R13260 GNDA.n3747 GNDA.n3744 4.5005
R13261 GNDA.n3748 GNDA.n555 4.5005
R13262 GNDA.n3752 GNDA.n3751 4.5005
R13263 GNDA.n3753 GNDA.n554 4.5005
R13264 GNDA.n3757 GNDA.n3754 4.5005
R13265 GNDA.n3758 GNDA.n553 4.5005
R13266 GNDA.n3762 GNDA.n3761 4.5005
R13267 GNDA.n1443 GNDA.n1442 4.5005
R13268 GNDA.n776 GNDA.n775 4.5005
R13269 GNDA.n1388 GNDA.n1387 4.5005
R13270 GNDA.n1392 GNDA.n1389 4.5005
R13271 GNDA.n1393 GNDA.n1386 4.5005
R13272 GNDA.n1397 GNDA.n1396 4.5005
R13273 GNDA.n1398 GNDA.n1385 4.5005
R13274 GNDA.n1402 GNDA.n1399 4.5005
R13275 GNDA.n1403 GNDA.n1384 4.5005
R13276 GNDA.n1407 GNDA.n1406 4.5005
R13277 GNDA.n1408 GNDA.n1383 4.5005
R13278 GNDA.n1412 GNDA.n1409 4.5005
R13279 GNDA.n1413 GNDA.n1382 4.5005
R13280 GNDA.n1417 GNDA.n1416 4.5005
R13281 GNDA.n1418 GNDA.n1381 4.5005
R13282 GNDA.n1422 GNDA.n1419 4.5005
R13283 GNDA.n1423 GNDA.n1380 4.5005
R13284 GNDA.n1427 GNDA.n1426 4.5005
R13285 GNDA.n1428 GNDA.n1379 4.5005
R13286 GNDA.n1432 GNDA.n1429 4.5005
R13287 GNDA.n1433 GNDA.n1378 4.5005
R13288 GNDA.n1437 GNDA.n1436 4.5005
R13289 GNDA.n1308 GNDA.n1307 4.5005
R13290 GNDA.n1311 GNDA.n1310 4.5005
R13291 GNDA.n1312 GNDA.n1306 4.5005
R13292 GNDA.n1316 GNDA.n1313 4.5005
R13293 GNDA.n1317 GNDA.n1305 4.5005
R13294 GNDA.n1321 GNDA.n1320 4.5005
R13295 GNDA.n1322 GNDA.n1304 4.5005
R13296 GNDA.n1326 GNDA.n1323 4.5005
R13297 GNDA.n1327 GNDA.n1303 4.5005
R13298 GNDA.n1331 GNDA.n1330 4.5005
R13299 GNDA.n1332 GNDA.n1302 4.5005
R13300 GNDA.n1336 GNDA.n1333 4.5005
R13301 GNDA.n1337 GNDA.n1301 4.5005
R13302 GNDA.n1341 GNDA.n1340 4.5005
R13303 GNDA.n1342 GNDA.n1300 4.5005
R13304 GNDA.n1346 GNDA.n1343 4.5005
R13305 GNDA.n1347 GNDA.n1299 4.5005
R13306 GNDA.n1351 GNDA.n1350 4.5005
R13307 GNDA.n1352 GNDA.n1298 4.5005
R13308 GNDA.n1356 GNDA.n1353 4.5005
R13309 GNDA.n1357 GNDA.n1297 4.5005
R13310 GNDA.n1361 GNDA.n1360 4.5005
R13311 GNDA.n1226 GNDA.n1225 4.5005
R13312 GNDA.n1229 GNDA.n1228 4.5005
R13313 GNDA.n1230 GNDA.n1224 4.5005
R13314 GNDA.n1234 GNDA.n1231 4.5005
R13315 GNDA.n1235 GNDA.n1223 4.5005
R13316 GNDA.n1239 GNDA.n1238 4.5005
R13317 GNDA.n1240 GNDA.n1222 4.5005
R13318 GNDA.n1244 GNDA.n1241 4.5005
R13319 GNDA.n1245 GNDA.n1221 4.5005
R13320 GNDA.n1249 GNDA.n1248 4.5005
R13321 GNDA.n1250 GNDA.n1220 4.5005
R13322 GNDA.n1254 GNDA.n1251 4.5005
R13323 GNDA.n1255 GNDA.n1219 4.5005
R13324 GNDA.n1259 GNDA.n1258 4.5005
R13325 GNDA.n1260 GNDA.n1218 4.5005
R13326 GNDA.n1264 GNDA.n1261 4.5005
R13327 GNDA.n1265 GNDA.n1217 4.5005
R13328 GNDA.n1269 GNDA.n1268 4.5005
R13329 GNDA.n1270 GNDA.n1216 4.5005
R13330 GNDA.n1274 GNDA.n1271 4.5005
R13331 GNDA.n1275 GNDA.n1215 4.5005
R13332 GNDA.n1279 GNDA.n1278 4.5005
R13333 GNDA.n898 GNDA.n897 4.5005
R13334 GNDA.n901 GNDA.n900 4.5005
R13335 GNDA.n902 GNDA.n802 4.5005
R13336 GNDA.n906 GNDA.n903 4.5005
R13337 GNDA.n907 GNDA.n801 4.5005
R13338 GNDA.n911 GNDA.n910 4.5005
R13339 GNDA.n912 GNDA.n800 4.5005
R13340 GNDA.n916 GNDA.n913 4.5005
R13341 GNDA.n917 GNDA.n799 4.5005
R13342 GNDA.n921 GNDA.n920 4.5005
R13343 GNDA.n922 GNDA.n798 4.5005
R13344 GNDA.n926 GNDA.n923 4.5005
R13345 GNDA.n927 GNDA.n797 4.5005
R13346 GNDA.n931 GNDA.n930 4.5005
R13347 GNDA.n932 GNDA.n796 4.5005
R13348 GNDA.n936 GNDA.n933 4.5005
R13349 GNDA.n937 GNDA.n795 4.5005
R13350 GNDA.n941 GNDA.n940 4.5005
R13351 GNDA.n942 GNDA.n794 4.5005
R13352 GNDA.n946 GNDA.n943 4.5005
R13353 GNDA.n947 GNDA.n793 4.5005
R13354 GNDA.n951 GNDA.n950 4.5005
R13355 GNDA.n1144 GNDA.n1143 4.5005
R13356 GNDA.n1147 GNDA.n1146 4.5005
R13357 GNDA.n1148 GNDA.n1142 4.5005
R13358 GNDA.n1152 GNDA.n1149 4.5005
R13359 GNDA.n1153 GNDA.n1141 4.5005
R13360 GNDA.n1157 GNDA.n1156 4.5005
R13361 GNDA.n1158 GNDA.n1140 4.5005
R13362 GNDA.n1162 GNDA.n1159 4.5005
R13363 GNDA.n1163 GNDA.n1139 4.5005
R13364 GNDA.n1167 GNDA.n1166 4.5005
R13365 GNDA.n1168 GNDA.n1138 4.5005
R13366 GNDA.n1172 GNDA.n1169 4.5005
R13367 GNDA.n1173 GNDA.n1137 4.5005
R13368 GNDA.n1177 GNDA.n1176 4.5005
R13369 GNDA.n1178 GNDA.n1136 4.5005
R13370 GNDA.n1182 GNDA.n1179 4.5005
R13371 GNDA.n1183 GNDA.n1135 4.5005
R13372 GNDA.n1187 GNDA.n1186 4.5005
R13373 GNDA.n1188 GNDA.n1134 4.5005
R13374 GNDA.n1192 GNDA.n1189 4.5005
R13375 GNDA.n1193 GNDA.n1133 4.5005
R13376 GNDA.n1197 GNDA.n1196 4.5005
R13377 GNDA.n1062 GNDA.n1061 4.5005
R13378 GNDA.n1065 GNDA.n1064 4.5005
R13379 GNDA.n1066 GNDA.n1060 4.5005
R13380 GNDA.n1070 GNDA.n1067 4.5005
R13381 GNDA.n1071 GNDA.n1059 4.5005
R13382 GNDA.n1075 GNDA.n1074 4.5005
R13383 GNDA.n1076 GNDA.n1058 4.5005
R13384 GNDA.n1080 GNDA.n1077 4.5005
R13385 GNDA.n1081 GNDA.n1057 4.5005
R13386 GNDA.n1085 GNDA.n1084 4.5005
R13387 GNDA.n1086 GNDA.n1056 4.5005
R13388 GNDA.n1090 GNDA.n1087 4.5005
R13389 GNDA.n1091 GNDA.n1055 4.5005
R13390 GNDA.n1095 GNDA.n1094 4.5005
R13391 GNDA.n1096 GNDA.n1054 4.5005
R13392 GNDA.n1100 GNDA.n1097 4.5005
R13393 GNDA.n1101 GNDA.n1053 4.5005
R13394 GNDA.n1105 GNDA.n1104 4.5005
R13395 GNDA.n1106 GNDA.n1052 4.5005
R13396 GNDA.n1110 GNDA.n1107 4.5005
R13397 GNDA.n1111 GNDA.n1051 4.5005
R13398 GNDA.n1115 GNDA.n1114 4.5005
R13399 GNDA.n980 GNDA.n979 4.5005
R13400 GNDA.n983 GNDA.n982 4.5005
R13401 GNDA.n984 GNDA.n978 4.5005
R13402 GNDA.n988 GNDA.n985 4.5005
R13403 GNDA.n989 GNDA.n977 4.5005
R13404 GNDA.n993 GNDA.n992 4.5005
R13405 GNDA.n994 GNDA.n976 4.5005
R13406 GNDA.n998 GNDA.n995 4.5005
R13407 GNDA.n999 GNDA.n975 4.5005
R13408 GNDA.n1003 GNDA.n1002 4.5005
R13409 GNDA.n1004 GNDA.n974 4.5005
R13410 GNDA.n1008 GNDA.n1005 4.5005
R13411 GNDA.n1009 GNDA.n973 4.5005
R13412 GNDA.n1013 GNDA.n1012 4.5005
R13413 GNDA.n1014 GNDA.n972 4.5005
R13414 GNDA.n1018 GNDA.n1015 4.5005
R13415 GNDA.n1019 GNDA.n971 4.5005
R13416 GNDA.n1023 GNDA.n1022 4.5005
R13417 GNDA.n1024 GNDA.n970 4.5005
R13418 GNDA.n1028 GNDA.n1025 4.5005
R13419 GNDA.n1029 GNDA.n969 4.5005
R13420 GNDA.n1033 GNDA.n1032 4.5005
R13421 GNDA.n886 GNDA.n885 4.5005
R13422 GNDA.n807 GNDA.n806 4.5005
R13423 GNDA.n829 GNDA.n808 4.5005
R13424 GNDA.n830 GNDA.n809 4.5005
R13425 GNDA.n831 GNDA.n810 4.5005
R13426 GNDA.n832 GNDA.n811 4.5005
R13427 GNDA.n833 GNDA.n812 4.5005
R13428 GNDA.n834 GNDA.n813 4.5005
R13429 GNDA.n835 GNDA.n814 4.5005
R13430 GNDA.n836 GNDA.n815 4.5005
R13431 GNDA.n837 GNDA.n816 4.5005
R13432 GNDA.n838 GNDA.n817 4.5005
R13433 GNDA.n839 GNDA.n818 4.5005
R13434 GNDA.n840 GNDA.n819 4.5005
R13435 GNDA.n841 GNDA.n820 4.5005
R13436 GNDA.n842 GNDA.n821 4.5005
R13437 GNDA.n843 GNDA.n822 4.5005
R13438 GNDA.n844 GNDA.n823 4.5005
R13439 GNDA.n845 GNDA.n824 4.5005
R13440 GNDA.n846 GNDA.n825 4.5005
R13441 GNDA.n847 GNDA.n826 4.5005
R13442 GNDA.n848 GNDA.n827 4.5005
R13443 GNDA.n735 GNDA.n734 4.5005
R13444 GNDA.n656 GNDA.n655 4.5005
R13445 GNDA.n678 GNDA.n657 4.5005
R13446 GNDA.n679 GNDA.n658 4.5005
R13447 GNDA.n680 GNDA.n659 4.5005
R13448 GNDA.n681 GNDA.n660 4.5005
R13449 GNDA.n682 GNDA.n661 4.5005
R13450 GNDA.n683 GNDA.n662 4.5005
R13451 GNDA.n684 GNDA.n663 4.5005
R13452 GNDA.n685 GNDA.n664 4.5005
R13453 GNDA.n686 GNDA.n665 4.5005
R13454 GNDA.n687 GNDA.n666 4.5005
R13455 GNDA.n688 GNDA.n667 4.5005
R13456 GNDA.n689 GNDA.n668 4.5005
R13457 GNDA.n690 GNDA.n669 4.5005
R13458 GNDA.n691 GNDA.n670 4.5005
R13459 GNDA.n692 GNDA.n671 4.5005
R13460 GNDA.n693 GNDA.n672 4.5005
R13461 GNDA.n694 GNDA.n673 4.5005
R13462 GNDA.n695 GNDA.n674 4.5005
R13463 GNDA.n696 GNDA.n675 4.5005
R13464 GNDA.n697 GNDA.n676 4.5005
R13465 GNDA.n3400 GNDA.n3399 4.5005
R13466 GNDA.n3403 GNDA.n3402 4.5005
R13467 GNDA.n3404 GNDA.n651 4.5005
R13468 GNDA.n3408 GNDA.n3405 4.5005
R13469 GNDA.n3409 GNDA.n650 4.5005
R13470 GNDA.n3413 GNDA.n3412 4.5005
R13471 GNDA.n3414 GNDA.n649 4.5005
R13472 GNDA.n3418 GNDA.n3415 4.5005
R13473 GNDA.n3419 GNDA.n648 4.5005
R13474 GNDA.n3423 GNDA.n3422 4.5005
R13475 GNDA.n3424 GNDA.n647 4.5005
R13476 GNDA.n3428 GNDA.n3425 4.5005
R13477 GNDA.n3429 GNDA.n646 4.5005
R13478 GNDA.n3433 GNDA.n3432 4.5005
R13479 GNDA.n3434 GNDA.n645 4.5005
R13480 GNDA.n3438 GNDA.n3435 4.5005
R13481 GNDA.n3439 GNDA.n644 4.5005
R13482 GNDA.n3443 GNDA.n3442 4.5005
R13483 GNDA.n3444 GNDA.n643 4.5005
R13484 GNDA.n3448 GNDA.n3445 4.5005
R13485 GNDA.n3449 GNDA.n642 4.5005
R13486 GNDA.n3453 GNDA.n3452 4.5005
R13487 GNDA.n3524 GNDA.n3523 4.5005
R13488 GNDA.n613 GNDA.n612 4.5005
R13489 GNDA.n3469 GNDA.n3468 4.5005
R13490 GNDA.n3473 GNDA.n3470 4.5005
R13491 GNDA.n3474 GNDA.n3467 4.5005
R13492 GNDA.n3478 GNDA.n3477 4.5005
R13493 GNDA.n3479 GNDA.n3466 4.5005
R13494 GNDA.n3483 GNDA.n3480 4.5005
R13495 GNDA.n3484 GNDA.n3465 4.5005
R13496 GNDA.n3488 GNDA.n3487 4.5005
R13497 GNDA.n3489 GNDA.n3464 4.5005
R13498 GNDA.n3493 GNDA.n3490 4.5005
R13499 GNDA.n3494 GNDA.n3463 4.5005
R13500 GNDA.n3498 GNDA.n3497 4.5005
R13501 GNDA.n3499 GNDA.n3462 4.5005
R13502 GNDA.n3503 GNDA.n3500 4.5005
R13503 GNDA.n3504 GNDA.n3461 4.5005
R13504 GNDA.n3508 GNDA.n3507 4.5005
R13505 GNDA.n3509 GNDA.n3460 4.5005
R13506 GNDA.n3513 GNDA.n3510 4.5005
R13507 GNDA.n3514 GNDA.n3459 4.5005
R13508 GNDA.n3518 GNDA.n3517 4.5005
R13509 GNDA.n2258 GNDA.n2257 4.5005
R13510 GNDA.n2179 GNDA.n2178 4.5005
R13511 GNDA.n2201 GNDA.n2180 4.5005
R13512 GNDA.n2202 GNDA.n2181 4.5005
R13513 GNDA.n2203 GNDA.n2182 4.5005
R13514 GNDA.n2204 GNDA.n2183 4.5005
R13515 GNDA.n2205 GNDA.n2184 4.5005
R13516 GNDA.n2206 GNDA.n2185 4.5005
R13517 GNDA.n2207 GNDA.n2186 4.5005
R13518 GNDA.n2208 GNDA.n2187 4.5005
R13519 GNDA.n2209 GNDA.n2188 4.5005
R13520 GNDA.n2210 GNDA.n2189 4.5005
R13521 GNDA.n2211 GNDA.n2190 4.5005
R13522 GNDA.n2212 GNDA.n2191 4.5005
R13523 GNDA.n2213 GNDA.n2192 4.5005
R13524 GNDA.n2214 GNDA.n2193 4.5005
R13525 GNDA.n2215 GNDA.n2194 4.5005
R13526 GNDA.n2216 GNDA.n2195 4.5005
R13527 GNDA.n2217 GNDA.n2196 4.5005
R13528 GNDA.n2218 GNDA.n2197 4.5005
R13529 GNDA.n2219 GNDA.n2198 4.5005
R13530 GNDA.n2220 GNDA.n2199 4.5005
R13531 GNDA.n2288 GNDA.n2174 4.5005
R13532 GNDA.n2290 GNDA.n2289 4.5005
R13533 GNDA.n2293 GNDA.n2173 4.5005
R13534 GNDA.n2297 GNDA.n2296 4.5005
R13535 GNDA.n2298 GNDA.n2172 4.5005
R13536 GNDA.n2300 GNDA.n2299 4.5005
R13537 GNDA.n2303 GNDA.n2171 4.5005
R13538 GNDA.n2307 GNDA.n2306 4.5005
R13539 GNDA.n2308 GNDA.n2170 4.5005
R13540 GNDA.n2310 GNDA.n2309 4.5005
R13541 GNDA.n2313 GNDA.n2169 4.5005
R13542 GNDA.n2317 GNDA.n2316 4.5005
R13543 GNDA.n2318 GNDA.n2168 4.5005
R13544 GNDA.n2320 GNDA.n2319 4.5005
R13545 GNDA.n2323 GNDA.n2167 4.5005
R13546 GNDA.n2327 GNDA.n2326 4.5005
R13547 GNDA.n2328 GNDA.n2166 4.5005
R13548 GNDA.n2330 GNDA.n2329 4.5005
R13549 GNDA.n2333 GNDA.n2165 4.5005
R13550 GNDA.n2336 GNDA.n2335 4.5005
R13551 GNDA.n2337 GNDA.n2163 4.5005
R13552 GNDA.n2340 GNDA.n2339 4.5005
R13553 GNDA.n2274 GNDA.n2272 4.5005
R13554 GNDA.n2276 GNDA.n2275 4.5005
R13555 GNDA.n2275 GNDA.n2274 4.5005
R13556 GNDA.n2279 GNDA.n2277 4.5005
R13557 GNDA.n2281 GNDA.n2280 4.5005
R13558 GNDA.n2280 GNDA.n2279 4.5005
R13559 GNDA.n2286 GNDA.n2282 4.5005
R13560 GNDA.n2287 GNDA.n2265 4.5005
R13561 GNDA.n2287 GNDA.n2286 4.5005
R13562 GNDA.n2177 GNDA.n610 4.5005
R13563 GNDA.n2264 GNDA.n2177 4.5005
R13564 GNDA.n2264 GNDA.n2176 4.5005
R13565 GNDA.n3529 GNDA.n3528 4.5005
R13566 GNDA.n3528 GNDA.n3527 4.5005
R13567 GNDA.n3527 GNDA.n611 4.5005
R13568 GNDA.n3394 GNDA.n3391 4.5005
R13569 GNDA.n3395 GNDA.n3394 4.5005
R13570 GNDA.n3396 GNDA.n3395 4.5005
R13571 GNDA.n3387 GNDA.n654 4.5005
R13572 GNDA.n3390 GNDA.n654 4.5005
R13573 GNDA.n3390 GNDA.n653 4.5005
R13574 GNDA.n893 GNDA.n892 4.5005
R13575 GNDA.n892 GNDA.n739 4.5005
R13576 GNDA.n890 GNDA.n739 4.5005
R13577 GNDA.n3375 GNDA.n749 4.5005
R13578 GNDA.n3378 GNDA.n749 4.5005
R13579 GNDA.n3378 GNDA.n748 4.5005
R13580 GNDA.n3371 GNDA.n754 4.5005
R13581 GNDA.n3374 GNDA.n754 4.5005
R13582 GNDA.n3374 GNDA.n753 4.5005
R13583 GNDA.n3367 GNDA.n759 4.5005
R13584 GNDA.n3370 GNDA.n759 4.5005
R13585 GNDA.n3370 GNDA.n758 4.5005
R13586 GNDA.n1458 GNDA.n764 4.5005
R13587 GNDA.n1461 GNDA.n764 4.5005
R13588 GNDA.n1461 GNDA.n763 4.5005
R13589 GNDA.n1454 GNDA.n769 4.5005
R13590 GNDA.n1457 GNDA.n769 4.5005
R13591 GNDA.n1457 GNDA.n768 4.5005
R13592 GNDA.n774 GNDA.n570 4.5005
R13593 GNDA.n1449 GNDA.n774 4.5005
R13594 GNDA.n1449 GNDA.n773 4.5005
R13595 GNDA.n3703 GNDA.n533 4.5005
R13596 GNDA.n3704 GNDA.n3703 4.5005
R13597 GNDA.n3705 GNDA.n3704 4.5005
R13598 GNDA.n3849 GNDA.n3848 4.5005
R13599 GNDA.n3848 GNDA.n3847 4.5005
R13600 GNDA.n3847 GNDA.n534 4.5005
R13601 GNDA.n4605 GNDA.n437 4.5005
R13602 GNDA.n4608 GNDA.n437 4.5005
R13603 GNDA.n4608 GNDA.n436 4.5005
R13604 GNDA.n4601 GNDA.n442 4.5005
R13605 GNDA.n4604 GNDA.n442 4.5005
R13606 GNDA.n4604 GNDA.n441 4.5005
R13607 GNDA.n3940 GNDA.n435 4.5005
R13608 GNDA.n3941 GNDA.n3940 4.5005
R13609 GNDA.n3942 GNDA.n3941 4.5005
R13610 GNDA.n4593 GNDA.n478 4.5005
R13611 GNDA.n4596 GNDA.n478 4.5005
R13612 GNDA.n4596 GNDA.n477 4.5005
R13613 GNDA.n4589 GNDA.n483 4.5005
R13614 GNDA.n4592 GNDA.n483 4.5005
R13615 GNDA.n4592 GNDA.n482 4.5005
R13616 GNDA.n4585 GNDA.n488 4.5005
R13617 GNDA.n4588 GNDA.n488 4.5005
R13618 GNDA.n4588 GNDA.n487 4.5005
R13619 GNDA.n4581 GNDA.n493 4.5005
R13620 GNDA.n4584 GNDA.n493 4.5005
R13621 GNDA.n4584 GNDA.n492 4.5005
R13622 GNDA.n4577 GNDA.n498 4.5005
R13623 GNDA.n4580 GNDA.n498 4.5005
R13624 GNDA.n4580 GNDA.n497 4.5005
R13625 GNDA.n3535 GNDA.n606 4.5005
R13626 GNDA.n3535 GNDA.n3534 4.5005
R13627 GNDA.n3534 GNDA.n3530 4.5005
R13628 GNDA.n4597 GNDA.n474 4.5005
R13629 GNDA.n4600 GNDA.n474 4.5005
R13630 GNDA.n4600 GNDA.n446 4.5005
R13631 GNDA.n3702 GNDA.n3701 4.5005
R13632 GNDA.n3701 GNDA.n3700 4.5005
R13633 GNDA.n3700 GNDA.n3616 4.5005
R13634 GNDA.n2647 GNDA.n2646 4.5005
R13635 GNDA.n2650 GNDA.n1861 4.5005
R13636 GNDA.n2496 GNDA.n2492 4.5005
R13637 GNDA.n2500 GNDA.n2499 4.5005
R13638 GNDA.n2501 GNDA.n2491 4.5005
R13639 GNDA.n2505 GNDA.n2502 4.5005
R13640 GNDA.n2506 GNDA.n2490 4.5005
R13641 GNDA.n2510 GNDA.n2509 4.5005
R13642 GNDA.n2511 GNDA.n2489 4.5005
R13643 GNDA.n2515 GNDA.n2512 4.5005
R13644 GNDA.n2516 GNDA.n2488 4.5005
R13645 GNDA.n2520 GNDA.n2519 4.5005
R13646 GNDA.n2521 GNDA.n2487 4.5005
R13647 GNDA.n2525 GNDA.n2522 4.5005
R13648 GNDA.n2526 GNDA.n2486 4.5005
R13649 GNDA.n2530 GNDA.n2529 4.5005
R13650 GNDA.n2531 GNDA.n2485 4.5005
R13651 GNDA.n2535 GNDA.n2532 4.5005
R13652 GNDA.n2536 GNDA.n2484 4.5005
R13653 GNDA.n2540 GNDA.n2539 4.5005
R13654 GNDA.n2541 GNDA.n2483 4.5005
R13655 GNDA.n2543 GNDA.n2542 4.5005
R13656 GNDA.n1865 GNDA.n1864 4.5005
R13657 GNDA.n2643 GNDA.n2642 4.5005
R13658 GNDA.n3319 GNDA.t305 4.30719
R13659 GNDA.n346 GNDA.n302 4.26717
R13660 GNDA.n346 GNDA.n345 4.26717
R13661 GNDA.n345 GNDA.n344 4.26717
R13662 GNDA.n344 GNDA.n310 4.26717
R13663 GNDA.n338 GNDA.n310 4.26717
R13664 GNDA.n338 GNDA.n337 4.26717
R13665 GNDA.n337 GNDA.n336 4.26717
R13666 GNDA.n336 GNDA.n318 4.26717
R13667 GNDA.n330 GNDA.n318 4.26717
R13668 GNDA.n330 GNDA.n329 4.26717
R13669 GNDA.n329 GNDA.n328 4.26717
R13670 GNDA.n5075 GNDA.n134 4.26717
R13671 GNDA.n5069 GNDA.n134 4.26717
R13672 GNDA.n5069 GNDA.n5068 4.26717
R13673 GNDA.n5068 GNDA.n5067 4.26717
R13674 GNDA.n5067 GNDA.n5065 4.26717
R13675 GNDA.n5065 GNDA.n5062 4.26717
R13676 GNDA.n5062 GNDA.n5061 4.26717
R13677 GNDA.n5061 GNDA.n5058 4.26717
R13678 GNDA.n5058 GNDA.n5057 4.26717
R13679 GNDA.n5057 GNDA.n5054 4.26717
R13680 GNDA.n5054 GNDA.n5053 4.26717
R13681 GNDA.n3015 GNDA.n1848 4.26717
R13682 GNDA.n3021 GNDA.n1848 4.26717
R13683 GNDA.n3021 GNDA.n1844 4.26717
R13684 GNDA.n3026 GNDA.n1844 4.26717
R13685 GNDA.n3026 GNDA.n1842 4.26717
R13686 GNDA.n1842 GNDA.n1839 4.26717
R13687 GNDA.n3033 GNDA.n1839 4.26717
R13688 GNDA.n3033 GNDA.n1837 4.26717
R13689 GNDA.n1837 GNDA.n1835 4.26717
R13690 GNDA.n3040 GNDA.n1835 4.26717
R13691 GNDA.n3040 GNDA.n1833 4.26717
R13692 GNDA.n411 GNDA.n410 4.26717
R13693 GNDA.n410 GNDA.n371 4.26717
R13694 GNDA.n405 GNDA.n371 4.26717
R13695 GNDA.n405 GNDA.n404 4.26717
R13696 GNDA.n404 GNDA.n403 4.26717
R13697 GNDA.n403 GNDA.n379 4.26717
R13698 GNDA.n397 GNDA.n379 4.26717
R13699 GNDA.n397 GNDA.n396 4.26717
R13700 GNDA.n396 GNDA.n395 4.26717
R13701 GNDA.n395 GNDA.n390 4.26717
R13702 GNDA.n390 GNDA.n389 4.26717
R13703 GNDA.n1767 GNDA.n1564 4.26717
R13704 GNDA.n1767 GNDA.n1562 4.26717
R13705 GNDA.n1773 GNDA.n1562 4.26717
R13706 GNDA.n1773 GNDA.n1560 4.26717
R13707 GNDA.n1779 GNDA.n1560 4.26717
R13708 GNDA.n1779 GNDA.n1558 4.26717
R13709 GNDA.n1785 GNDA.n1558 4.26717
R13710 GNDA.n1785 GNDA.n1556 4.26717
R13711 GNDA.n1791 GNDA.n1556 4.26717
R13712 GNDA.n1791 GNDA.n1554 4.26717
R13713 GNDA.n1796 GNDA.n1554 4.26717
R13714 GNDA.n3168 GNDA.n3167 4.26717
R13715 GNDA.n3167 GNDA.n1805 4.26717
R13716 GNDA.n3163 GNDA.n1805 4.26717
R13717 GNDA.n3163 GNDA.n3162 4.26717
R13718 GNDA.n3162 GNDA.n1811 4.26717
R13719 GNDA.n3157 GNDA.n1811 4.26717
R13720 GNDA.n3157 GNDA.n3156 4.26717
R13721 GNDA.n3156 GNDA.n3155 4.26717
R13722 GNDA.n3155 GNDA.n1819 4.26717
R13723 GNDA.n3149 GNDA.n1819 4.26717
R13724 GNDA.n3149 GNDA.n3148 4.26717
R13725 GNDA.t187 GNDA.t272 4.14363
R13726 GNDA.n3366 GNDA.n3365 3.9606
R13727 GNDA.n4695 GNDA.n302 3.93531
R13728 GNDA.n5076 GNDA.n5075 3.93531
R13729 GNDA.n3015 GNDA.n2982 3.93531
R13730 GNDA.n411 GNDA.n365 3.93531
R13731 GNDA.n1588 GNDA.n1564 3.93531
R13732 GNDA.n3168 GNDA.n1800 3.93531
R13733 GNDA.n3137 GNDA.n3136 3.7893
R13734 GNDA.n3133 GNDA.n3048 3.7893
R13735 GNDA.n3132 GNDA.n3116 3.7893
R13736 GNDA.n3126 GNDA.n3125 3.7893
R13737 GNDA.n3121 GNDA.n3120 3.7893
R13738 GNDA.n3252 GNDA.n1514 3.7893
R13739 GNDA.n1513 GNDA.n1510 3.7893
R13740 GNDA.n3261 GNDA.n3260 3.7893
R13741 GNDA.n3294 GNDA.n1493 3.7893
R13742 GNDA.n3293 GNDA.n1494 3.7893
R13743 GNDA.n3281 GNDA.n3280 3.7893
R13744 GNDA.n3287 GNDA.n3286 3.7893
R13745 GNDA.n3283 GNDA.n3282 3.7893
R13746 GNDA.n2722 GNDA.n1472 3.7893
R13747 GNDA.n2728 GNDA.n2726 3.7893
R13748 GNDA.n2730 GNDA.n2729 3.7893
R13749 GNDA.n5047 GNDA.n165 3.7893
R13750 GNDA.n5044 GNDA.n5043 3.7893
R13751 GNDA.n200 GNDA.n167 3.7893
R13752 GNDA.n218 GNDA.n217 3.7893
R13753 GNDA.n215 GNDA.n214 3.7893
R13754 GNDA.n210 GNDA.n203 3.7893
R13755 GNDA.n207 GNDA.n206 3.7893
R13756 GNDA.n4985 GNDA.n187 3.7893
R13757 GNDA.n1703 GNDA.n1678 3.7893
R13758 GNDA.n1702 GNDA.n1699 3.7893
R13759 GNDA.n1698 GNDA.n1679 3.7893
R13760 GNDA.n1695 GNDA.n1694 3.7893
R13761 GNDA.n1691 GNDA.n1680 3.7893
R13762 GNDA.n1684 GNDA.n1681 3.7893
R13763 GNDA.n1708 GNDA.n1603 3.7893
R13764 GNDA.n1709 GNDA.n1602 3.7893
R13765 GNDA.n4976 GNDA.n4975 3.7893
R13766 GNDA.n4972 GNDA.n4866 3.7893
R13767 GNDA.n4971 GNDA.n4869 3.7893
R13768 GNDA.n4968 GNDA.n4967 3.7893
R13769 GNDA.n4894 GNDA.n4870 3.7893
R13770 GNDA.n4903 GNDA.n4902 3.7893
R13771 GNDA.n4906 GNDA.n4893 3.7893
R13772 GNDA.n4911 GNDA.n4907 3.7893
R13773 GNDA.n5255 GNDA.n5254 3.7893
R13774 GNDA.n5251 GNDA.n59 3.7893
R13775 GNDA.n5250 GNDA.n62 3.7893
R13776 GNDA.n5247 GNDA.n5246 3.7893
R13777 GNDA.n5173 GNDA.n63 3.7893
R13778 GNDA.n5182 GNDA.n5181 3.7893
R13779 GNDA.n5185 GNDA.n5172 3.7893
R13780 GNDA.n5190 GNDA.n5186 3.7893
R13781 GNDA.n4832 GNDA.n4721 3.7893
R13782 GNDA.n4829 GNDA.n4828 3.7893
R13783 GNDA.n4745 GNDA.n4722 3.7893
R13784 GNDA.n4750 GNDA.n4748 3.7893
R13785 GNDA.n4755 GNDA.n4751 3.7893
R13786 GNDA.n4762 GNDA.n4761 3.7893
R13787 GNDA.n4765 GNDA.n4744 3.7893
R13788 GNDA.n4770 GNDA.n4766 3.7893
R13789 GNDA.n2909 GNDA.n2907 3.7893
R13790 GNDA.n2908 GNDA.n2667 3.7893
R13791 GNDA.n2915 GNDA.n2914 3.7893
R13792 GNDA.n2830 GNDA.n2668 3.7893
R13793 GNDA.n2834 GNDA.n2832 3.7893
R13794 GNDA.n2841 GNDA.n2840 3.7893
R13795 GNDA.n2850 GNDA.n2688 3.7893
R13796 GNDA.n2849 GNDA.n2686 3.7893
R13797 GNDA.n5264 GNDA.n22 3.7893
R13798 GNDA.n5263 GNDA.n23 3.7893
R13799 GNDA.n33 GNDA.n32 3.7893
R13800 GNDA.n39 GNDA.n38 3.7893
R13801 GNDA.n35 GNDA.n34 3.7893
R13802 GNDA.n5098 GNDA.n1 3.7893
R13803 GNDA.n5103 GNDA.n5101 3.7893
R13804 GNDA.n5108 GNDA.n5104 3.7893
R13805 GNDA.n3253 GNDA 3.7381
R13806 GNDA GNDA.n3299 3.7381
R13807 GNDA.n211 GNDA 3.7381
R13808 GNDA GNDA.n1687 3.7381
R13809 GNDA.n4899 GNDA 3.7381
R13810 GNDA.n5178 GNDA 3.7381
R13811 GNDA.n4758 GNDA 3.7381
R13812 GNDA.n2839 GNDA 3.7381
R13813 GNDA GNDA.n5269 3.7381
R13814 GNDA.n3583 GNDA.n585 3.65764
R13815 GNDA.n3583 GNDA.n3582 3.65764
R13816 GNDA.n3572 GNDA.n587 3.65764
R13817 GNDA.n3573 GNDA.n3572 3.65764
R13818 GNDA.n2338 GNDA.n2150 3.50398
R13819 GNDA.n2493 GNDA.n2471 3.47871
R13820 GNDA.n2582 GNDA.n2546 3.47821
R13821 GNDA.n3661 GNDA.n3660 3.47821
R13822 GNDA.n4569 GNDA.n4568 3.47821
R13823 GNDA.n4493 GNDA.n4492 3.47821
R13824 GNDA.n4411 GNDA.n4410 3.47821
R13825 GNDA.n4329 GNDA.n4328 3.47821
R13826 GNDA.n4247 GNDA.n4246 3.47821
R13827 GNDA.n4001 GNDA.n4000 3.47821
R13828 GNDA.n4165 GNDA.n4164 3.47821
R13829 GNDA.n4083 GNDA.n4082 3.47821
R13830 GNDA.n3898 GNDA.n3897 3.47821
R13831 GNDA.n3840 GNDA.n3839 3.47821
R13832 GNDA.n3764 GNDA.n3763 3.47821
R13833 GNDA.n1439 GNDA.n1438 3.47821
R13834 GNDA.n1363 GNDA.n1362 3.47821
R13835 GNDA.n1281 GNDA.n1280 3.47821
R13836 GNDA.n953 GNDA.n952 3.47821
R13837 GNDA.n1199 GNDA.n1198 3.47821
R13838 GNDA.n1117 GNDA.n1116 3.47821
R13839 GNDA.n1035 GNDA.n1034 3.47821
R13840 GNDA.n850 GNDA.n849 3.47821
R13841 GNDA.n699 GNDA.n698 3.47821
R13842 GNDA.n3455 GNDA.n3454 3.47821
R13843 GNDA.n3520 GNDA.n3519 3.47821
R13844 GNDA.n2222 GNDA.n2221 3.47821
R13845 GNDA.n2174 GNDA.n2151 3.43627
R13846 GNDA.n3939 GNDA.t257 3.42907
R13847 GNDA.n3939 GNDA.t278 3.42907
R13848 GNDA.n3936 GNDA.t280 3.42907
R13849 GNDA.n3936 GNDA.t263 3.42907
R13850 GNDA.n803 GNDA.t283 3.42907
R13851 GNDA.n803 GNDA.t232 3.42907
R13852 GNDA.n889 GNDA.t261 3.42907
R13853 GNDA.n889 GNDA.t238 3.42907
R13854 GNDA.n2559 GNDA.n2558 3.4105
R13855 GNDA.n2621 GNDA.n2620 3.4105
R13856 GNDA.n2619 GNDA.n2618 3.4105
R13857 GNDA.n2617 GNDA.n2563 3.4105
R13858 GNDA.n2562 GNDA.n2561 3.4105
R13859 GNDA.n2613 GNDA.n2612 3.4105
R13860 GNDA.n2611 GNDA.n2610 3.4105
R13861 GNDA.n2609 GNDA.n2567 3.4105
R13862 GNDA.n2566 GNDA.n2565 3.4105
R13863 GNDA.n2605 GNDA.n2604 3.4105
R13864 GNDA.n2603 GNDA.n2602 3.4105
R13865 GNDA.n2601 GNDA.n2571 3.4105
R13866 GNDA.n2570 GNDA.n2569 3.4105
R13867 GNDA.n2597 GNDA.n2596 3.4105
R13868 GNDA.n2595 GNDA.n2594 3.4105
R13869 GNDA.n2593 GNDA.n2575 3.4105
R13870 GNDA.n2574 GNDA.n2573 3.4105
R13871 GNDA.n2589 GNDA.n2588 3.4105
R13872 GNDA.n2587 GNDA.n2586 3.4105
R13873 GNDA.n2585 GNDA.n2579 3.4105
R13874 GNDA.n2578 GNDA.n2577 3.4105
R13875 GNDA.n2581 GNDA.n2580 3.4105
R13876 GNDA.n2638 GNDA.n2637 3.4105
R13877 GNDA.n3662 GNDA.n3639 3.4105
R13878 GNDA.n3664 GNDA.n3638 3.4105
R13879 GNDA.n3665 GNDA.n3637 3.4105
R13880 GNDA.n3667 GNDA.n3636 3.4105
R13881 GNDA.n3668 GNDA.n3635 3.4105
R13882 GNDA.n3670 GNDA.n3634 3.4105
R13883 GNDA.n3671 GNDA.n3633 3.4105
R13884 GNDA.n3673 GNDA.n3632 3.4105
R13885 GNDA.n3674 GNDA.n3631 3.4105
R13886 GNDA.n3676 GNDA.n3630 3.4105
R13887 GNDA.n3677 GNDA.n3629 3.4105
R13888 GNDA.n3679 GNDA.n3628 3.4105
R13889 GNDA.n3680 GNDA.n3627 3.4105
R13890 GNDA.n3682 GNDA.n3626 3.4105
R13891 GNDA.n3683 GNDA.n3625 3.4105
R13892 GNDA.n3685 GNDA.n3624 3.4105
R13893 GNDA.n3686 GNDA.n3623 3.4105
R13894 GNDA.n3688 GNDA.n3622 3.4105
R13895 GNDA.n3689 GNDA.n3621 3.4105
R13896 GNDA.n3691 GNDA.n3620 3.4105
R13897 GNDA.n3692 GNDA.n3619 3.4105
R13898 GNDA.n3694 GNDA.n3618 3.4105
R13899 GNDA.n3696 GNDA.n3695 3.4105
R13900 GNDA.n4507 GNDA.n4506 3.4105
R13901 GNDA.n4566 GNDA.n4565 3.4105
R13902 GNDA.n4564 GNDA.n4563 3.4105
R13903 GNDA.n4562 GNDA.n4561 3.4105
R13904 GNDA.n4560 GNDA.n4509 3.4105
R13905 GNDA.n4556 GNDA.n4555 3.4105
R13906 GNDA.n4554 GNDA.n4553 3.4105
R13907 GNDA.n4552 GNDA.n4551 3.4105
R13908 GNDA.n4550 GNDA.n4511 3.4105
R13909 GNDA.n4546 GNDA.n4545 3.4105
R13910 GNDA.n4544 GNDA.n4543 3.4105
R13911 GNDA.n4542 GNDA.n4541 3.4105
R13912 GNDA.n4540 GNDA.n4513 3.4105
R13913 GNDA.n4536 GNDA.n4535 3.4105
R13914 GNDA.n4534 GNDA.n4533 3.4105
R13915 GNDA.n4532 GNDA.n4531 3.4105
R13916 GNDA.n4530 GNDA.n4515 3.4105
R13917 GNDA.n4526 GNDA.n4525 3.4105
R13918 GNDA.n4524 GNDA.n4523 3.4105
R13919 GNDA.n4522 GNDA.n4521 3.4105
R13920 GNDA.n4520 GNDA.n4517 3.4105
R13921 GNDA.n501 GNDA.n500 3.4105
R13922 GNDA.n4572 GNDA.n4571 3.4105
R13923 GNDA.n4426 GNDA.n4425 3.4105
R13924 GNDA.n4490 GNDA.n4489 3.4105
R13925 GNDA.n4488 GNDA.n4487 3.4105
R13926 GNDA.n4486 GNDA.n4485 3.4105
R13927 GNDA.n4484 GNDA.n4428 3.4105
R13928 GNDA.n4480 GNDA.n4479 3.4105
R13929 GNDA.n4478 GNDA.n4477 3.4105
R13930 GNDA.n4476 GNDA.n4475 3.4105
R13931 GNDA.n4474 GNDA.n4430 3.4105
R13932 GNDA.n4470 GNDA.n4469 3.4105
R13933 GNDA.n4468 GNDA.n4467 3.4105
R13934 GNDA.n4466 GNDA.n4465 3.4105
R13935 GNDA.n4464 GNDA.n4432 3.4105
R13936 GNDA.n4460 GNDA.n4459 3.4105
R13937 GNDA.n4458 GNDA.n4457 3.4105
R13938 GNDA.n4456 GNDA.n4455 3.4105
R13939 GNDA.n4454 GNDA.n4434 3.4105
R13940 GNDA.n4450 GNDA.n4449 3.4105
R13941 GNDA.n4448 GNDA.n4447 3.4105
R13942 GNDA.n4446 GNDA.n4445 3.4105
R13943 GNDA.n4444 GNDA.n4436 3.4105
R13944 GNDA.n4440 GNDA.n4439 3.4105
R13945 GNDA.n4438 GNDA.n4413 3.4105
R13946 GNDA.n4344 GNDA.n4343 3.4105
R13947 GNDA.n4408 GNDA.n4407 3.4105
R13948 GNDA.n4406 GNDA.n4405 3.4105
R13949 GNDA.n4404 GNDA.n4403 3.4105
R13950 GNDA.n4402 GNDA.n4346 3.4105
R13951 GNDA.n4398 GNDA.n4397 3.4105
R13952 GNDA.n4396 GNDA.n4395 3.4105
R13953 GNDA.n4394 GNDA.n4393 3.4105
R13954 GNDA.n4392 GNDA.n4348 3.4105
R13955 GNDA.n4388 GNDA.n4387 3.4105
R13956 GNDA.n4386 GNDA.n4385 3.4105
R13957 GNDA.n4384 GNDA.n4383 3.4105
R13958 GNDA.n4382 GNDA.n4350 3.4105
R13959 GNDA.n4378 GNDA.n4377 3.4105
R13960 GNDA.n4376 GNDA.n4375 3.4105
R13961 GNDA.n4374 GNDA.n4373 3.4105
R13962 GNDA.n4372 GNDA.n4352 3.4105
R13963 GNDA.n4368 GNDA.n4367 3.4105
R13964 GNDA.n4366 GNDA.n4365 3.4105
R13965 GNDA.n4364 GNDA.n4363 3.4105
R13966 GNDA.n4362 GNDA.n4354 3.4105
R13967 GNDA.n4358 GNDA.n4357 3.4105
R13968 GNDA.n4356 GNDA.n4331 3.4105
R13969 GNDA.n4262 GNDA.n4261 3.4105
R13970 GNDA.n4326 GNDA.n4325 3.4105
R13971 GNDA.n4324 GNDA.n4323 3.4105
R13972 GNDA.n4322 GNDA.n4321 3.4105
R13973 GNDA.n4320 GNDA.n4264 3.4105
R13974 GNDA.n4316 GNDA.n4315 3.4105
R13975 GNDA.n4314 GNDA.n4313 3.4105
R13976 GNDA.n4312 GNDA.n4311 3.4105
R13977 GNDA.n4310 GNDA.n4266 3.4105
R13978 GNDA.n4306 GNDA.n4305 3.4105
R13979 GNDA.n4304 GNDA.n4303 3.4105
R13980 GNDA.n4302 GNDA.n4301 3.4105
R13981 GNDA.n4300 GNDA.n4268 3.4105
R13982 GNDA.n4296 GNDA.n4295 3.4105
R13983 GNDA.n4294 GNDA.n4293 3.4105
R13984 GNDA.n4292 GNDA.n4291 3.4105
R13985 GNDA.n4290 GNDA.n4270 3.4105
R13986 GNDA.n4286 GNDA.n4285 3.4105
R13987 GNDA.n4284 GNDA.n4283 3.4105
R13988 GNDA.n4282 GNDA.n4281 3.4105
R13989 GNDA.n4280 GNDA.n4272 3.4105
R13990 GNDA.n4276 GNDA.n4275 3.4105
R13991 GNDA.n4274 GNDA.n4249 3.4105
R13992 GNDA.n4180 GNDA.n4179 3.4105
R13993 GNDA.n4244 GNDA.n4243 3.4105
R13994 GNDA.n4242 GNDA.n4241 3.4105
R13995 GNDA.n4240 GNDA.n4239 3.4105
R13996 GNDA.n4238 GNDA.n4182 3.4105
R13997 GNDA.n4234 GNDA.n4233 3.4105
R13998 GNDA.n4232 GNDA.n4231 3.4105
R13999 GNDA.n4230 GNDA.n4229 3.4105
R14000 GNDA.n4228 GNDA.n4184 3.4105
R14001 GNDA.n4224 GNDA.n4223 3.4105
R14002 GNDA.n4222 GNDA.n4221 3.4105
R14003 GNDA.n4220 GNDA.n4219 3.4105
R14004 GNDA.n4218 GNDA.n4186 3.4105
R14005 GNDA.n4214 GNDA.n4213 3.4105
R14006 GNDA.n4212 GNDA.n4211 3.4105
R14007 GNDA.n4210 GNDA.n4209 3.4105
R14008 GNDA.n4208 GNDA.n4188 3.4105
R14009 GNDA.n4204 GNDA.n4203 3.4105
R14010 GNDA.n4202 GNDA.n4201 3.4105
R14011 GNDA.n4200 GNDA.n4199 3.4105
R14012 GNDA.n4198 GNDA.n4190 3.4105
R14013 GNDA.n4194 GNDA.n4193 3.4105
R14014 GNDA.n4192 GNDA.n4167 3.4105
R14015 GNDA.n516 GNDA.n515 3.4105
R14016 GNDA.n3998 GNDA.n3997 3.4105
R14017 GNDA.n3996 GNDA.n3995 3.4105
R14018 GNDA.n3994 GNDA.n3993 3.4105
R14019 GNDA.n3992 GNDA.n518 3.4105
R14020 GNDA.n3988 GNDA.n3987 3.4105
R14021 GNDA.n3986 GNDA.n3985 3.4105
R14022 GNDA.n3984 GNDA.n3983 3.4105
R14023 GNDA.n3982 GNDA.n520 3.4105
R14024 GNDA.n3978 GNDA.n3977 3.4105
R14025 GNDA.n3976 GNDA.n3975 3.4105
R14026 GNDA.n3974 GNDA.n3973 3.4105
R14027 GNDA.n3972 GNDA.n522 3.4105
R14028 GNDA.n3968 GNDA.n3967 3.4105
R14029 GNDA.n3966 GNDA.n3965 3.4105
R14030 GNDA.n3964 GNDA.n3963 3.4105
R14031 GNDA.n3962 GNDA.n524 3.4105
R14032 GNDA.n3958 GNDA.n3957 3.4105
R14033 GNDA.n3956 GNDA.n3955 3.4105
R14034 GNDA.n3954 GNDA.n3953 3.4105
R14035 GNDA.n3952 GNDA.n526 3.4105
R14036 GNDA.n3948 GNDA.n3947 3.4105
R14037 GNDA.n3946 GNDA.n503 3.4105
R14038 GNDA.n4098 GNDA.n4097 3.4105
R14039 GNDA.n4162 GNDA.n4161 3.4105
R14040 GNDA.n4160 GNDA.n4159 3.4105
R14041 GNDA.n4158 GNDA.n4157 3.4105
R14042 GNDA.n4156 GNDA.n4100 3.4105
R14043 GNDA.n4152 GNDA.n4151 3.4105
R14044 GNDA.n4150 GNDA.n4149 3.4105
R14045 GNDA.n4148 GNDA.n4147 3.4105
R14046 GNDA.n4146 GNDA.n4102 3.4105
R14047 GNDA.n4142 GNDA.n4141 3.4105
R14048 GNDA.n4140 GNDA.n4139 3.4105
R14049 GNDA.n4138 GNDA.n4137 3.4105
R14050 GNDA.n4136 GNDA.n4104 3.4105
R14051 GNDA.n4132 GNDA.n4131 3.4105
R14052 GNDA.n4130 GNDA.n4129 3.4105
R14053 GNDA.n4128 GNDA.n4127 3.4105
R14054 GNDA.n4126 GNDA.n4106 3.4105
R14055 GNDA.n4122 GNDA.n4121 3.4105
R14056 GNDA.n4120 GNDA.n4119 3.4105
R14057 GNDA.n4118 GNDA.n4117 3.4105
R14058 GNDA.n4116 GNDA.n4108 3.4105
R14059 GNDA.n4112 GNDA.n4111 3.4105
R14060 GNDA.n4110 GNDA.n4085 3.4105
R14061 GNDA.n4016 GNDA.n4015 3.4105
R14062 GNDA.n4080 GNDA.n4079 3.4105
R14063 GNDA.n4078 GNDA.n4077 3.4105
R14064 GNDA.n4076 GNDA.n4075 3.4105
R14065 GNDA.n4074 GNDA.n4018 3.4105
R14066 GNDA.n4070 GNDA.n4069 3.4105
R14067 GNDA.n4068 GNDA.n4067 3.4105
R14068 GNDA.n4066 GNDA.n4065 3.4105
R14069 GNDA.n4064 GNDA.n4020 3.4105
R14070 GNDA.n4060 GNDA.n4059 3.4105
R14071 GNDA.n4058 GNDA.n4057 3.4105
R14072 GNDA.n4056 GNDA.n4055 3.4105
R14073 GNDA.n4054 GNDA.n4022 3.4105
R14074 GNDA.n4050 GNDA.n4049 3.4105
R14075 GNDA.n4048 GNDA.n4047 3.4105
R14076 GNDA.n4046 GNDA.n4045 3.4105
R14077 GNDA.n4044 GNDA.n4024 3.4105
R14078 GNDA.n4040 GNDA.n4039 3.4105
R14079 GNDA.n4038 GNDA.n4037 3.4105
R14080 GNDA.n4036 GNDA.n4035 3.4105
R14081 GNDA.n4034 GNDA.n4026 3.4105
R14082 GNDA.n4030 GNDA.n4029 3.4105
R14083 GNDA.n4028 GNDA.n4003 3.4105
R14084 GNDA.n3899 GNDA.n3876 3.4105
R14085 GNDA.n3901 GNDA.n3875 3.4105
R14086 GNDA.n3902 GNDA.n3874 3.4105
R14087 GNDA.n3904 GNDA.n3873 3.4105
R14088 GNDA.n3905 GNDA.n3872 3.4105
R14089 GNDA.n3907 GNDA.n3871 3.4105
R14090 GNDA.n3908 GNDA.n3870 3.4105
R14091 GNDA.n3910 GNDA.n3869 3.4105
R14092 GNDA.n3911 GNDA.n3868 3.4105
R14093 GNDA.n3913 GNDA.n3867 3.4105
R14094 GNDA.n3914 GNDA.n3866 3.4105
R14095 GNDA.n3916 GNDA.n3865 3.4105
R14096 GNDA.n3917 GNDA.n3864 3.4105
R14097 GNDA.n3919 GNDA.n3863 3.4105
R14098 GNDA.n3920 GNDA.n3862 3.4105
R14099 GNDA.n3922 GNDA.n3861 3.4105
R14100 GNDA.n3923 GNDA.n3860 3.4105
R14101 GNDA.n3925 GNDA.n3859 3.4105
R14102 GNDA.n3926 GNDA.n3858 3.4105
R14103 GNDA.n3928 GNDA.n3857 3.4105
R14104 GNDA.n3929 GNDA.n3856 3.4105
R14105 GNDA.n3931 GNDA.n3855 3.4105
R14106 GNDA.n3933 GNDA.n3932 3.4105
R14107 GNDA.n3778 GNDA.n3777 3.4105
R14108 GNDA.n3837 GNDA.n3836 3.4105
R14109 GNDA.n3835 GNDA.n3834 3.4105
R14110 GNDA.n3833 GNDA.n3832 3.4105
R14111 GNDA.n3831 GNDA.n3780 3.4105
R14112 GNDA.n3827 GNDA.n3826 3.4105
R14113 GNDA.n3825 GNDA.n3824 3.4105
R14114 GNDA.n3823 GNDA.n3822 3.4105
R14115 GNDA.n3821 GNDA.n3782 3.4105
R14116 GNDA.n3817 GNDA.n3816 3.4105
R14117 GNDA.n3815 GNDA.n3814 3.4105
R14118 GNDA.n3813 GNDA.n3812 3.4105
R14119 GNDA.n3811 GNDA.n3784 3.4105
R14120 GNDA.n3807 GNDA.n3806 3.4105
R14121 GNDA.n3805 GNDA.n3804 3.4105
R14122 GNDA.n3803 GNDA.n3802 3.4105
R14123 GNDA.n3801 GNDA.n3786 3.4105
R14124 GNDA.n3797 GNDA.n3796 3.4105
R14125 GNDA.n3795 GNDA.n3794 3.4105
R14126 GNDA.n3793 GNDA.n3792 3.4105
R14127 GNDA.n3791 GNDA.n3788 3.4105
R14128 GNDA.n537 GNDA.n536 3.4105
R14129 GNDA.n3843 GNDA.n3842 3.4105
R14130 GNDA.n552 GNDA.n551 3.4105
R14131 GNDA.n3761 GNDA.n3760 3.4105
R14132 GNDA.n3759 GNDA.n3758 3.4105
R14133 GNDA.n3757 GNDA.n3756 3.4105
R14134 GNDA.n3755 GNDA.n554 3.4105
R14135 GNDA.n3751 GNDA.n3750 3.4105
R14136 GNDA.n3749 GNDA.n3748 3.4105
R14137 GNDA.n3747 GNDA.n3746 3.4105
R14138 GNDA.n3745 GNDA.n556 3.4105
R14139 GNDA.n3741 GNDA.n3740 3.4105
R14140 GNDA.n3739 GNDA.n3738 3.4105
R14141 GNDA.n3737 GNDA.n3736 3.4105
R14142 GNDA.n3735 GNDA.n558 3.4105
R14143 GNDA.n3731 GNDA.n3730 3.4105
R14144 GNDA.n3729 GNDA.n3728 3.4105
R14145 GNDA.n3727 GNDA.n3726 3.4105
R14146 GNDA.n3725 GNDA.n560 3.4105
R14147 GNDA.n3721 GNDA.n3720 3.4105
R14148 GNDA.n3719 GNDA.n3718 3.4105
R14149 GNDA.n3717 GNDA.n3716 3.4105
R14150 GNDA.n3715 GNDA.n562 3.4105
R14151 GNDA.n3711 GNDA.n3710 3.4105
R14152 GNDA.n3709 GNDA.n539 3.4105
R14153 GNDA.n1377 GNDA.n1376 3.4105
R14154 GNDA.n1436 GNDA.n1435 3.4105
R14155 GNDA.n1434 GNDA.n1433 3.4105
R14156 GNDA.n1432 GNDA.n1431 3.4105
R14157 GNDA.n1430 GNDA.n1379 3.4105
R14158 GNDA.n1426 GNDA.n1425 3.4105
R14159 GNDA.n1424 GNDA.n1423 3.4105
R14160 GNDA.n1422 GNDA.n1421 3.4105
R14161 GNDA.n1420 GNDA.n1381 3.4105
R14162 GNDA.n1416 GNDA.n1415 3.4105
R14163 GNDA.n1414 GNDA.n1413 3.4105
R14164 GNDA.n1412 GNDA.n1411 3.4105
R14165 GNDA.n1410 GNDA.n1383 3.4105
R14166 GNDA.n1406 GNDA.n1405 3.4105
R14167 GNDA.n1404 GNDA.n1403 3.4105
R14168 GNDA.n1402 GNDA.n1401 3.4105
R14169 GNDA.n1400 GNDA.n1385 3.4105
R14170 GNDA.n1396 GNDA.n1395 3.4105
R14171 GNDA.n1394 GNDA.n1393 3.4105
R14172 GNDA.n1392 GNDA.n1391 3.4105
R14173 GNDA.n1390 GNDA.n1387 3.4105
R14174 GNDA.n777 GNDA.n776 3.4105
R14175 GNDA.n1442 GNDA.n1441 3.4105
R14176 GNDA.n1296 GNDA.n1295 3.4105
R14177 GNDA.n1360 GNDA.n1359 3.4105
R14178 GNDA.n1358 GNDA.n1357 3.4105
R14179 GNDA.n1356 GNDA.n1355 3.4105
R14180 GNDA.n1354 GNDA.n1298 3.4105
R14181 GNDA.n1350 GNDA.n1349 3.4105
R14182 GNDA.n1348 GNDA.n1347 3.4105
R14183 GNDA.n1346 GNDA.n1345 3.4105
R14184 GNDA.n1344 GNDA.n1300 3.4105
R14185 GNDA.n1340 GNDA.n1339 3.4105
R14186 GNDA.n1338 GNDA.n1337 3.4105
R14187 GNDA.n1336 GNDA.n1335 3.4105
R14188 GNDA.n1334 GNDA.n1302 3.4105
R14189 GNDA.n1330 GNDA.n1329 3.4105
R14190 GNDA.n1328 GNDA.n1327 3.4105
R14191 GNDA.n1326 GNDA.n1325 3.4105
R14192 GNDA.n1324 GNDA.n1304 3.4105
R14193 GNDA.n1320 GNDA.n1319 3.4105
R14194 GNDA.n1318 GNDA.n1317 3.4105
R14195 GNDA.n1316 GNDA.n1315 3.4105
R14196 GNDA.n1314 GNDA.n1306 3.4105
R14197 GNDA.n1310 GNDA.n1309 3.4105
R14198 GNDA.n1308 GNDA.n1283 3.4105
R14199 GNDA.n1214 GNDA.n1213 3.4105
R14200 GNDA.n1278 GNDA.n1277 3.4105
R14201 GNDA.n1276 GNDA.n1275 3.4105
R14202 GNDA.n1274 GNDA.n1273 3.4105
R14203 GNDA.n1272 GNDA.n1216 3.4105
R14204 GNDA.n1268 GNDA.n1267 3.4105
R14205 GNDA.n1266 GNDA.n1265 3.4105
R14206 GNDA.n1264 GNDA.n1263 3.4105
R14207 GNDA.n1262 GNDA.n1218 3.4105
R14208 GNDA.n1258 GNDA.n1257 3.4105
R14209 GNDA.n1256 GNDA.n1255 3.4105
R14210 GNDA.n1254 GNDA.n1253 3.4105
R14211 GNDA.n1252 GNDA.n1220 3.4105
R14212 GNDA.n1248 GNDA.n1247 3.4105
R14213 GNDA.n1246 GNDA.n1245 3.4105
R14214 GNDA.n1244 GNDA.n1243 3.4105
R14215 GNDA.n1242 GNDA.n1222 3.4105
R14216 GNDA.n1238 GNDA.n1237 3.4105
R14217 GNDA.n1236 GNDA.n1235 3.4105
R14218 GNDA.n1234 GNDA.n1233 3.4105
R14219 GNDA.n1232 GNDA.n1224 3.4105
R14220 GNDA.n1228 GNDA.n1227 3.4105
R14221 GNDA.n1226 GNDA.n1201 3.4105
R14222 GNDA.n792 GNDA.n791 3.4105
R14223 GNDA.n950 GNDA.n949 3.4105
R14224 GNDA.n948 GNDA.n947 3.4105
R14225 GNDA.n946 GNDA.n945 3.4105
R14226 GNDA.n944 GNDA.n794 3.4105
R14227 GNDA.n940 GNDA.n939 3.4105
R14228 GNDA.n938 GNDA.n937 3.4105
R14229 GNDA.n936 GNDA.n935 3.4105
R14230 GNDA.n934 GNDA.n796 3.4105
R14231 GNDA.n930 GNDA.n929 3.4105
R14232 GNDA.n928 GNDA.n927 3.4105
R14233 GNDA.n926 GNDA.n925 3.4105
R14234 GNDA.n924 GNDA.n798 3.4105
R14235 GNDA.n920 GNDA.n919 3.4105
R14236 GNDA.n918 GNDA.n917 3.4105
R14237 GNDA.n916 GNDA.n915 3.4105
R14238 GNDA.n914 GNDA.n800 3.4105
R14239 GNDA.n910 GNDA.n909 3.4105
R14240 GNDA.n908 GNDA.n907 3.4105
R14241 GNDA.n906 GNDA.n905 3.4105
R14242 GNDA.n904 GNDA.n802 3.4105
R14243 GNDA.n900 GNDA.n899 3.4105
R14244 GNDA.n898 GNDA.n779 3.4105
R14245 GNDA.n1132 GNDA.n1131 3.4105
R14246 GNDA.n1196 GNDA.n1195 3.4105
R14247 GNDA.n1194 GNDA.n1193 3.4105
R14248 GNDA.n1192 GNDA.n1191 3.4105
R14249 GNDA.n1190 GNDA.n1134 3.4105
R14250 GNDA.n1186 GNDA.n1185 3.4105
R14251 GNDA.n1184 GNDA.n1183 3.4105
R14252 GNDA.n1182 GNDA.n1181 3.4105
R14253 GNDA.n1180 GNDA.n1136 3.4105
R14254 GNDA.n1176 GNDA.n1175 3.4105
R14255 GNDA.n1174 GNDA.n1173 3.4105
R14256 GNDA.n1172 GNDA.n1171 3.4105
R14257 GNDA.n1170 GNDA.n1138 3.4105
R14258 GNDA.n1166 GNDA.n1165 3.4105
R14259 GNDA.n1164 GNDA.n1163 3.4105
R14260 GNDA.n1162 GNDA.n1161 3.4105
R14261 GNDA.n1160 GNDA.n1140 3.4105
R14262 GNDA.n1156 GNDA.n1155 3.4105
R14263 GNDA.n1154 GNDA.n1153 3.4105
R14264 GNDA.n1152 GNDA.n1151 3.4105
R14265 GNDA.n1150 GNDA.n1142 3.4105
R14266 GNDA.n1146 GNDA.n1145 3.4105
R14267 GNDA.n1144 GNDA.n1119 3.4105
R14268 GNDA.n1050 GNDA.n1049 3.4105
R14269 GNDA.n1114 GNDA.n1113 3.4105
R14270 GNDA.n1112 GNDA.n1111 3.4105
R14271 GNDA.n1110 GNDA.n1109 3.4105
R14272 GNDA.n1108 GNDA.n1052 3.4105
R14273 GNDA.n1104 GNDA.n1103 3.4105
R14274 GNDA.n1102 GNDA.n1101 3.4105
R14275 GNDA.n1100 GNDA.n1099 3.4105
R14276 GNDA.n1098 GNDA.n1054 3.4105
R14277 GNDA.n1094 GNDA.n1093 3.4105
R14278 GNDA.n1092 GNDA.n1091 3.4105
R14279 GNDA.n1090 GNDA.n1089 3.4105
R14280 GNDA.n1088 GNDA.n1056 3.4105
R14281 GNDA.n1084 GNDA.n1083 3.4105
R14282 GNDA.n1082 GNDA.n1081 3.4105
R14283 GNDA.n1080 GNDA.n1079 3.4105
R14284 GNDA.n1078 GNDA.n1058 3.4105
R14285 GNDA.n1074 GNDA.n1073 3.4105
R14286 GNDA.n1072 GNDA.n1071 3.4105
R14287 GNDA.n1070 GNDA.n1069 3.4105
R14288 GNDA.n1068 GNDA.n1060 3.4105
R14289 GNDA.n1064 GNDA.n1063 3.4105
R14290 GNDA.n1062 GNDA.n1037 3.4105
R14291 GNDA.n968 GNDA.n967 3.4105
R14292 GNDA.n1032 GNDA.n1031 3.4105
R14293 GNDA.n1030 GNDA.n1029 3.4105
R14294 GNDA.n1028 GNDA.n1027 3.4105
R14295 GNDA.n1026 GNDA.n970 3.4105
R14296 GNDA.n1022 GNDA.n1021 3.4105
R14297 GNDA.n1020 GNDA.n1019 3.4105
R14298 GNDA.n1018 GNDA.n1017 3.4105
R14299 GNDA.n1016 GNDA.n972 3.4105
R14300 GNDA.n1012 GNDA.n1011 3.4105
R14301 GNDA.n1010 GNDA.n1009 3.4105
R14302 GNDA.n1008 GNDA.n1007 3.4105
R14303 GNDA.n1006 GNDA.n974 3.4105
R14304 GNDA.n1002 GNDA.n1001 3.4105
R14305 GNDA.n1000 GNDA.n999 3.4105
R14306 GNDA.n998 GNDA.n997 3.4105
R14307 GNDA.n996 GNDA.n976 3.4105
R14308 GNDA.n992 GNDA.n991 3.4105
R14309 GNDA.n990 GNDA.n989 3.4105
R14310 GNDA.n988 GNDA.n987 3.4105
R14311 GNDA.n986 GNDA.n978 3.4105
R14312 GNDA.n982 GNDA.n981 3.4105
R14313 GNDA.n980 GNDA.n955 3.4105
R14314 GNDA.n851 GNDA.n828 3.4105
R14315 GNDA.n853 GNDA.n827 3.4105
R14316 GNDA.n854 GNDA.n826 3.4105
R14317 GNDA.n856 GNDA.n825 3.4105
R14318 GNDA.n857 GNDA.n824 3.4105
R14319 GNDA.n859 GNDA.n823 3.4105
R14320 GNDA.n860 GNDA.n822 3.4105
R14321 GNDA.n862 GNDA.n821 3.4105
R14322 GNDA.n863 GNDA.n820 3.4105
R14323 GNDA.n865 GNDA.n819 3.4105
R14324 GNDA.n866 GNDA.n818 3.4105
R14325 GNDA.n868 GNDA.n817 3.4105
R14326 GNDA.n869 GNDA.n816 3.4105
R14327 GNDA.n871 GNDA.n815 3.4105
R14328 GNDA.n872 GNDA.n814 3.4105
R14329 GNDA.n874 GNDA.n813 3.4105
R14330 GNDA.n875 GNDA.n812 3.4105
R14331 GNDA.n877 GNDA.n811 3.4105
R14332 GNDA.n878 GNDA.n810 3.4105
R14333 GNDA.n880 GNDA.n809 3.4105
R14334 GNDA.n881 GNDA.n808 3.4105
R14335 GNDA.n883 GNDA.n807 3.4105
R14336 GNDA.n885 GNDA.n884 3.4105
R14337 GNDA.n700 GNDA.n677 3.4105
R14338 GNDA.n702 GNDA.n676 3.4105
R14339 GNDA.n703 GNDA.n675 3.4105
R14340 GNDA.n705 GNDA.n674 3.4105
R14341 GNDA.n706 GNDA.n673 3.4105
R14342 GNDA.n708 GNDA.n672 3.4105
R14343 GNDA.n709 GNDA.n671 3.4105
R14344 GNDA.n711 GNDA.n670 3.4105
R14345 GNDA.n712 GNDA.n669 3.4105
R14346 GNDA.n714 GNDA.n668 3.4105
R14347 GNDA.n715 GNDA.n667 3.4105
R14348 GNDA.n717 GNDA.n666 3.4105
R14349 GNDA.n718 GNDA.n665 3.4105
R14350 GNDA.n720 GNDA.n664 3.4105
R14351 GNDA.n721 GNDA.n663 3.4105
R14352 GNDA.n723 GNDA.n662 3.4105
R14353 GNDA.n724 GNDA.n661 3.4105
R14354 GNDA.n726 GNDA.n660 3.4105
R14355 GNDA.n727 GNDA.n659 3.4105
R14356 GNDA.n729 GNDA.n658 3.4105
R14357 GNDA.n730 GNDA.n657 3.4105
R14358 GNDA.n732 GNDA.n656 3.4105
R14359 GNDA.n734 GNDA.n733 3.4105
R14360 GNDA.n641 GNDA.n640 3.4105
R14361 GNDA.n3452 GNDA.n3451 3.4105
R14362 GNDA.n3450 GNDA.n3449 3.4105
R14363 GNDA.n3448 GNDA.n3447 3.4105
R14364 GNDA.n3446 GNDA.n643 3.4105
R14365 GNDA.n3442 GNDA.n3441 3.4105
R14366 GNDA.n3440 GNDA.n3439 3.4105
R14367 GNDA.n3438 GNDA.n3437 3.4105
R14368 GNDA.n3436 GNDA.n645 3.4105
R14369 GNDA.n3432 GNDA.n3431 3.4105
R14370 GNDA.n3430 GNDA.n3429 3.4105
R14371 GNDA.n3428 GNDA.n3427 3.4105
R14372 GNDA.n3426 GNDA.n647 3.4105
R14373 GNDA.n3422 GNDA.n3421 3.4105
R14374 GNDA.n3420 GNDA.n3419 3.4105
R14375 GNDA.n3418 GNDA.n3417 3.4105
R14376 GNDA.n3416 GNDA.n649 3.4105
R14377 GNDA.n3412 GNDA.n3411 3.4105
R14378 GNDA.n3410 GNDA.n3409 3.4105
R14379 GNDA.n3408 GNDA.n3407 3.4105
R14380 GNDA.n3406 GNDA.n651 3.4105
R14381 GNDA.n3402 GNDA.n3401 3.4105
R14382 GNDA.n3400 GNDA.n627 3.4105
R14383 GNDA.n3458 GNDA.n3457 3.4105
R14384 GNDA.n3517 GNDA.n3516 3.4105
R14385 GNDA.n3515 GNDA.n3514 3.4105
R14386 GNDA.n3513 GNDA.n3512 3.4105
R14387 GNDA.n3511 GNDA.n3460 3.4105
R14388 GNDA.n3507 GNDA.n3506 3.4105
R14389 GNDA.n3505 GNDA.n3504 3.4105
R14390 GNDA.n3503 GNDA.n3502 3.4105
R14391 GNDA.n3501 GNDA.n3462 3.4105
R14392 GNDA.n3497 GNDA.n3496 3.4105
R14393 GNDA.n3495 GNDA.n3494 3.4105
R14394 GNDA.n3493 GNDA.n3492 3.4105
R14395 GNDA.n3491 GNDA.n3464 3.4105
R14396 GNDA.n3487 GNDA.n3486 3.4105
R14397 GNDA.n3485 GNDA.n3484 3.4105
R14398 GNDA.n3483 GNDA.n3482 3.4105
R14399 GNDA.n3481 GNDA.n3466 3.4105
R14400 GNDA.n3477 GNDA.n3476 3.4105
R14401 GNDA.n3475 GNDA.n3474 3.4105
R14402 GNDA.n3473 GNDA.n3472 3.4105
R14403 GNDA.n3471 GNDA.n3468 3.4105
R14404 GNDA.n614 GNDA.n613 3.4105
R14405 GNDA.n3523 GNDA.n3522 3.4105
R14406 GNDA.n2223 GNDA.n2200 3.4105
R14407 GNDA.n2225 GNDA.n2199 3.4105
R14408 GNDA.n2226 GNDA.n2198 3.4105
R14409 GNDA.n2228 GNDA.n2197 3.4105
R14410 GNDA.n2229 GNDA.n2196 3.4105
R14411 GNDA.n2231 GNDA.n2195 3.4105
R14412 GNDA.n2232 GNDA.n2194 3.4105
R14413 GNDA.n2234 GNDA.n2193 3.4105
R14414 GNDA.n2235 GNDA.n2192 3.4105
R14415 GNDA.n2237 GNDA.n2191 3.4105
R14416 GNDA.n2238 GNDA.n2190 3.4105
R14417 GNDA.n2240 GNDA.n2189 3.4105
R14418 GNDA.n2241 GNDA.n2188 3.4105
R14419 GNDA.n2243 GNDA.n2187 3.4105
R14420 GNDA.n2244 GNDA.n2186 3.4105
R14421 GNDA.n2246 GNDA.n2185 3.4105
R14422 GNDA.n2247 GNDA.n2184 3.4105
R14423 GNDA.n2249 GNDA.n2183 3.4105
R14424 GNDA.n2250 GNDA.n2182 3.4105
R14425 GNDA.n2252 GNDA.n2181 3.4105
R14426 GNDA.n2253 GNDA.n2180 3.4105
R14427 GNDA.n2255 GNDA.n2179 3.4105
R14428 GNDA.n2257 GNDA.n2256 3.4105
R14429 GNDA.n2256 GNDA.n615 3.4105
R14430 GNDA.n2222 GNDA.n615 3.4105
R14431 GNDA.n3522 GNDA.n3521 3.4105
R14432 GNDA.n3521 GNDA.n3520 3.4105
R14433 GNDA.n3456 GNDA.n627 3.4105
R14434 GNDA.n3456 GNDA.n3455 3.4105
R14435 GNDA.n733 GNDA.n639 3.4105
R14436 GNDA.n699 GNDA.n639 3.4105
R14437 GNDA.n884 GNDA.n778 3.4105
R14438 GNDA.n850 GNDA.n778 3.4105
R14439 GNDA.n1036 GNDA.n955 3.4105
R14440 GNDA.n1036 GNDA.n1035 3.4105
R14441 GNDA.n1118 GNDA.n1037 3.4105
R14442 GNDA.n1118 GNDA.n1117 3.4105
R14443 GNDA.n1200 GNDA.n1119 3.4105
R14444 GNDA.n1200 GNDA.n1199 3.4105
R14445 GNDA.n954 GNDA.n779 3.4105
R14446 GNDA.n954 GNDA.n953 3.4105
R14447 GNDA.n1282 GNDA.n1201 3.4105
R14448 GNDA.n1282 GNDA.n1281 3.4105
R14449 GNDA.n1364 GNDA.n1283 3.4105
R14450 GNDA.n1364 GNDA.n1363 3.4105
R14451 GNDA.n1441 GNDA.n1440 3.4105
R14452 GNDA.n1440 GNDA.n1439 3.4105
R14453 GNDA.n3765 GNDA.n539 3.4105
R14454 GNDA.n3765 GNDA.n3764 3.4105
R14455 GNDA.n3842 GNDA.n3841 3.4105
R14456 GNDA.n3841 GNDA.n3840 3.4105
R14457 GNDA.n3932 GNDA.n502 3.4105
R14458 GNDA.n3898 GNDA.n502 3.4105
R14459 GNDA.n4084 GNDA.n4003 3.4105
R14460 GNDA.n4084 GNDA.n4083 3.4105
R14461 GNDA.n4166 GNDA.n4085 3.4105
R14462 GNDA.n4166 GNDA.n4165 3.4105
R14463 GNDA.n4002 GNDA.n503 3.4105
R14464 GNDA.n4002 GNDA.n4001 3.4105
R14465 GNDA.n4248 GNDA.n4167 3.4105
R14466 GNDA.n4248 GNDA.n4247 3.4105
R14467 GNDA.n4330 GNDA.n4249 3.4105
R14468 GNDA.n4330 GNDA.n4329 3.4105
R14469 GNDA.n4412 GNDA.n4331 3.4105
R14470 GNDA.n4412 GNDA.n4411 3.4105
R14471 GNDA.n4494 GNDA.n4413 3.4105
R14472 GNDA.n4494 GNDA.n4493 3.4105
R14473 GNDA.n4571 GNDA.n4570 3.4105
R14474 GNDA.n4570 GNDA.n4569 3.4105
R14475 GNDA.n3695 GNDA.n538 3.4105
R14476 GNDA.n3661 GNDA.n538 3.4105
R14477 GNDA.n2164 GNDA.n2162 3.4105
R14478 GNDA.n2341 GNDA.n2340 3.4105
R14479 GNDA.n2163 GNDA.n2161 3.4105
R14480 GNDA.n2335 GNDA.n2334 3.4105
R14481 GNDA.n2333 GNDA.n2332 3.4105
R14482 GNDA.n2331 GNDA.n2330 3.4105
R14483 GNDA.n2324 GNDA.n2166 3.4105
R14484 GNDA.n2326 GNDA.n2325 3.4105
R14485 GNDA.n2323 GNDA.n2322 3.4105
R14486 GNDA.n2321 GNDA.n2320 3.4105
R14487 GNDA.n2314 GNDA.n2168 3.4105
R14488 GNDA.n2316 GNDA.n2315 3.4105
R14489 GNDA.n2313 GNDA.n2312 3.4105
R14490 GNDA.n2311 GNDA.n2310 3.4105
R14491 GNDA.n2304 GNDA.n2170 3.4105
R14492 GNDA.n2306 GNDA.n2305 3.4105
R14493 GNDA.n2303 GNDA.n2302 3.4105
R14494 GNDA.n2301 GNDA.n2300 3.4105
R14495 GNDA.n2294 GNDA.n2172 3.4105
R14496 GNDA.n2296 GNDA.n2295 3.4105
R14497 GNDA.n2293 GNDA.n2292 3.4105
R14498 GNDA.n2291 GNDA.n2290 3.4105
R14499 GNDA.n1866 GNDA.n1865 3.4105
R14500 GNDA.n2544 GNDA.n2543 3.4105
R14501 GNDA.n2483 GNDA.n2482 3.4105
R14502 GNDA.n2539 GNDA.n2538 3.4105
R14503 GNDA.n2537 GNDA.n2536 3.4105
R14504 GNDA.n2535 GNDA.n2534 3.4105
R14505 GNDA.n2533 GNDA.n2485 3.4105
R14506 GNDA.n2529 GNDA.n2528 3.4105
R14507 GNDA.n2527 GNDA.n2526 3.4105
R14508 GNDA.n2525 GNDA.n2524 3.4105
R14509 GNDA.n2523 GNDA.n2487 3.4105
R14510 GNDA.n2519 GNDA.n2518 3.4105
R14511 GNDA.n2517 GNDA.n2516 3.4105
R14512 GNDA.n2515 GNDA.n2514 3.4105
R14513 GNDA.n2513 GNDA.n2489 3.4105
R14514 GNDA.n2509 GNDA.n2508 3.4105
R14515 GNDA.n2507 GNDA.n2506 3.4105
R14516 GNDA.n2505 GNDA.n2504 3.4105
R14517 GNDA.n2503 GNDA.n2491 3.4105
R14518 GNDA.n2499 GNDA.n2498 3.4105
R14519 GNDA.n2497 GNDA.n2496 3.4105
R14520 GNDA.n2495 GNDA.n2494 3.4105
R14521 GNDA.n2642 GNDA.n2641 3.4105
R14522 GNDA.n2640 GNDA.n2471 3.4105
R14523 GNDA.n2641 GNDA.n2640 3.4105
R14524 GNDA.n2639 GNDA.n2546 3.4105
R14525 GNDA.n2639 GNDA.n2638 3.4105
R14526 GNDA.n2468 GNDA.n1901 3.4105
R14527 GNDA.n2468 GNDA.n2467 3.4105
R14528 GNDA.n2467 GNDA.n1884 3.4105
R14529 GNDA.n1920 GNDA.n1901 3.4105
R14530 GNDA.n2435 GNDA.n1920 3.4105
R14531 GNDA.n1966 GNDA.n1920 3.4105
R14532 GNDA.n2437 GNDA.n1920 3.4105
R14533 GNDA.n1965 GNDA.n1920 3.4105
R14534 GNDA.n2439 GNDA.n1920 3.4105
R14535 GNDA.n1964 GNDA.n1920 3.4105
R14536 GNDA.n2441 GNDA.n1920 3.4105
R14537 GNDA.n1963 GNDA.n1920 3.4105
R14538 GNDA.n2443 GNDA.n1920 3.4105
R14539 GNDA.n1962 GNDA.n1920 3.4105
R14540 GNDA.n2445 GNDA.n1920 3.4105
R14541 GNDA.n1961 GNDA.n1920 3.4105
R14542 GNDA.n2447 GNDA.n1920 3.4105
R14543 GNDA.n1960 GNDA.n1920 3.4105
R14544 GNDA.n2449 GNDA.n1920 3.4105
R14545 GNDA.n1959 GNDA.n1920 3.4105
R14546 GNDA.n2451 GNDA.n1920 3.4105
R14547 GNDA.n1958 GNDA.n1920 3.4105
R14548 GNDA.n2453 GNDA.n1920 3.4105
R14549 GNDA.n1957 GNDA.n1920 3.4105
R14550 GNDA.n2455 GNDA.n1920 3.4105
R14551 GNDA.n1956 GNDA.n1920 3.4105
R14552 GNDA.n2457 GNDA.n1920 3.4105
R14553 GNDA.n1955 GNDA.n1920 3.4105
R14554 GNDA.n2459 GNDA.n1920 3.4105
R14555 GNDA.n1954 GNDA.n1920 3.4105
R14556 GNDA.n2461 GNDA.n1920 3.4105
R14557 GNDA.n1953 GNDA.n1920 3.4105
R14558 GNDA.n2463 GNDA.n1920 3.4105
R14559 GNDA.n1952 GNDA.n1920 3.4105
R14560 GNDA.n2465 GNDA.n1920 3.4105
R14561 GNDA.n2467 GNDA.n1920 3.4105
R14562 GNDA.n1917 GNDA.n1901 3.4105
R14563 GNDA.n2435 GNDA.n1917 3.4105
R14564 GNDA.n1966 GNDA.n1917 3.4105
R14565 GNDA.n2437 GNDA.n1917 3.4105
R14566 GNDA.n1965 GNDA.n1917 3.4105
R14567 GNDA.n2439 GNDA.n1917 3.4105
R14568 GNDA.n1964 GNDA.n1917 3.4105
R14569 GNDA.n2441 GNDA.n1917 3.4105
R14570 GNDA.n1963 GNDA.n1917 3.4105
R14571 GNDA.n2443 GNDA.n1917 3.4105
R14572 GNDA.n1962 GNDA.n1917 3.4105
R14573 GNDA.n2445 GNDA.n1917 3.4105
R14574 GNDA.n1961 GNDA.n1917 3.4105
R14575 GNDA.n2447 GNDA.n1917 3.4105
R14576 GNDA.n1960 GNDA.n1917 3.4105
R14577 GNDA.n2449 GNDA.n1917 3.4105
R14578 GNDA.n1959 GNDA.n1917 3.4105
R14579 GNDA.n2451 GNDA.n1917 3.4105
R14580 GNDA.n1958 GNDA.n1917 3.4105
R14581 GNDA.n2453 GNDA.n1917 3.4105
R14582 GNDA.n1957 GNDA.n1917 3.4105
R14583 GNDA.n2455 GNDA.n1917 3.4105
R14584 GNDA.n1956 GNDA.n1917 3.4105
R14585 GNDA.n2457 GNDA.n1917 3.4105
R14586 GNDA.n1955 GNDA.n1917 3.4105
R14587 GNDA.n2459 GNDA.n1917 3.4105
R14588 GNDA.n1954 GNDA.n1917 3.4105
R14589 GNDA.n2461 GNDA.n1917 3.4105
R14590 GNDA.n1953 GNDA.n1917 3.4105
R14591 GNDA.n2463 GNDA.n1917 3.4105
R14592 GNDA.n1952 GNDA.n1917 3.4105
R14593 GNDA.n2465 GNDA.n1917 3.4105
R14594 GNDA.n2467 GNDA.n1917 3.4105
R14595 GNDA.n1922 GNDA.n1901 3.4105
R14596 GNDA.n2435 GNDA.n1922 3.4105
R14597 GNDA.n1966 GNDA.n1922 3.4105
R14598 GNDA.n2437 GNDA.n1922 3.4105
R14599 GNDA.n1965 GNDA.n1922 3.4105
R14600 GNDA.n2439 GNDA.n1922 3.4105
R14601 GNDA.n1964 GNDA.n1922 3.4105
R14602 GNDA.n2441 GNDA.n1922 3.4105
R14603 GNDA.n1963 GNDA.n1922 3.4105
R14604 GNDA.n2443 GNDA.n1922 3.4105
R14605 GNDA.n1962 GNDA.n1922 3.4105
R14606 GNDA.n2445 GNDA.n1922 3.4105
R14607 GNDA.n1961 GNDA.n1922 3.4105
R14608 GNDA.n2447 GNDA.n1922 3.4105
R14609 GNDA.n1960 GNDA.n1922 3.4105
R14610 GNDA.n2449 GNDA.n1922 3.4105
R14611 GNDA.n1959 GNDA.n1922 3.4105
R14612 GNDA.n2451 GNDA.n1922 3.4105
R14613 GNDA.n1958 GNDA.n1922 3.4105
R14614 GNDA.n2453 GNDA.n1922 3.4105
R14615 GNDA.n1957 GNDA.n1922 3.4105
R14616 GNDA.n2455 GNDA.n1922 3.4105
R14617 GNDA.n1956 GNDA.n1922 3.4105
R14618 GNDA.n2457 GNDA.n1922 3.4105
R14619 GNDA.n1955 GNDA.n1922 3.4105
R14620 GNDA.n2459 GNDA.n1922 3.4105
R14621 GNDA.n1954 GNDA.n1922 3.4105
R14622 GNDA.n2461 GNDA.n1922 3.4105
R14623 GNDA.n1953 GNDA.n1922 3.4105
R14624 GNDA.n2463 GNDA.n1922 3.4105
R14625 GNDA.n1952 GNDA.n1922 3.4105
R14626 GNDA.n2465 GNDA.n1922 3.4105
R14627 GNDA.n2467 GNDA.n1922 3.4105
R14628 GNDA.n1916 GNDA.n1901 3.4105
R14629 GNDA.n2435 GNDA.n1916 3.4105
R14630 GNDA.n1966 GNDA.n1916 3.4105
R14631 GNDA.n2437 GNDA.n1916 3.4105
R14632 GNDA.n1965 GNDA.n1916 3.4105
R14633 GNDA.n2439 GNDA.n1916 3.4105
R14634 GNDA.n1964 GNDA.n1916 3.4105
R14635 GNDA.n2441 GNDA.n1916 3.4105
R14636 GNDA.n1963 GNDA.n1916 3.4105
R14637 GNDA.n2443 GNDA.n1916 3.4105
R14638 GNDA.n1962 GNDA.n1916 3.4105
R14639 GNDA.n2445 GNDA.n1916 3.4105
R14640 GNDA.n1961 GNDA.n1916 3.4105
R14641 GNDA.n2447 GNDA.n1916 3.4105
R14642 GNDA.n1960 GNDA.n1916 3.4105
R14643 GNDA.n2449 GNDA.n1916 3.4105
R14644 GNDA.n1959 GNDA.n1916 3.4105
R14645 GNDA.n2451 GNDA.n1916 3.4105
R14646 GNDA.n1958 GNDA.n1916 3.4105
R14647 GNDA.n2453 GNDA.n1916 3.4105
R14648 GNDA.n1957 GNDA.n1916 3.4105
R14649 GNDA.n2455 GNDA.n1916 3.4105
R14650 GNDA.n1956 GNDA.n1916 3.4105
R14651 GNDA.n2457 GNDA.n1916 3.4105
R14652 GNDA.n1955 GNDA.n1916 3.4105
R14653 GNDA.n2459 GNDA.n1916 3.4105
R14654 GNDA.n1954 GNDA.n1916 3.4105
R14655 GNDA.n2461 GNDA.n1916 3.4105
R14656 GNDA.n1953 GNDA.n1916 3.4105
R14657 GNDA.n2463 GNDA.n1916 3.4105
R14658 GNDA.n1952 GNDA.n1916 3.4105
R14659 GNDA.n2465 GNDA.n1916 3.4105
R14660 GNDA.n2467 GNDA.n1916 3.4105
R14661 GNDA.n1924 GNDA.n1901 3.4105
R14662 GNDA.n2435 GNDA.n1924 3.4105
R14663 GNDA.n1966 GNDA.n1924 3.4105
R14664 GNDA.n2437 GNDA.n1924 3.4105
R14665 GNDA.n1965 GNDA.n1924 3.4105
R14666 GNDA.n2439 GNDA.n1924 3.4105
R14667 GNDA.n1964 GNDA.n1924 3.4105
R14668 GNDA.n2441 GNDA.n1924 3.4105
R14669 GNDA.n1963 GNDA.n1924 3.4105
R14670 GNDA.n2443 GNDA.n1924 3.4105
R14671 GNDA.n1962 GNDA.n1924 3.4105
R14672 GNDA.n2445 GNDA.n1924 3.4105
R14673 GNDA.n1961 GNDA.n1924 3.4105
R14674 GNDA.n2447 GNDA.n1924 3.4105
R14675 GNDA.n1960 GNDA.n1924 3.4105
R14676 GNDA.n2449 GNDA.n1924 3.4105
R14677 GNDA.n1959 GNDA.n1924 3.4105
R14678 GNDA.n2451 GNDA.n1924 3.4105
R14679 GNDA.n1958 GNDA.n1924 3.4105
R14680 GNDA.n2453 GNDA.n1924 3.4105
R14681 GNDA.n1957 GNDA.n1924 3.4105
R14682 GNDA.n2455 GNDA.n1924 3.4105
R14683 GNDA.n1956 GNDA.n1924 3.4105
R14684 GNDA.n2457 GNDA.n1924 3.4105
R14685 GNDA.n1955 GNDA.n1924 3.4105
R14686 GNDA.n2459 GNDA.n1924 3.4105
R14687 GNDA.n1954 GNDA.n1924 3.4105
R14688 GNDA.n2461 GNDA.n1924 3.4105
R14689 GNDA.n1953 GNDA.n1924 3.4105
R14690 GNDA.n2463 GNDA.n1924 3.4105
R14691 GNDA.n1952 GNDA.n1924 3.4105
R14692 GNDA.n2465 GNDA.n1924 3.4105
R14693 GNDA.n2467 GNDA.n1924 3.4105
R14694 GNDA.n1915 GNDA.n1901 3.4105
R14695 GNDA.n2435 GNDA.n1915 3.4105
R14696 GNDA.n1966 GNDA.n1915 3.4105
R14697 GNDA.n2437 GNDA.n1915 3.4105
R14698 GNDA.n1965 GNDA.n1915 3.4105
R14699 GNDA.n2439 GNDA.n1915 3.4105
R14700 GNDA.n1964 GNDA.n1915 3.4105
R14701 GNDA.n2441 GNDA.n1915 3.4105
R14702 GNDA.n1963 GNDA.n1915 3.4105
R14703 GNDA.n2443 GNDA.n1915 3.4105
R14704 GNDA.n1962 GNDA.n1915 3.4105
R14705 GNDA.n2445 GNDA.n1915 3.4105
R14706 GNDA.n1961 GNDA.n1915 3.4105
R14707 GNDA.n2447 GNDA.n1915 3.4105
R14708 GNDA.n1960 GNDA.n1915 3.4105
R14709 GNDA.n2449 GNDA.n1915 3.4105
R14710 GNDA.n1959 GNDA.n1915 3.4105
R14711 GNDA.n2451 GNDA.n1915 3.4105
R14712 GNDA.n1958 GNDA.n1915 3.4105
R14713 GNDA.n2453 GNDA.n1915 3.4105
R14714 GNDA.n1957 GNDA.n1915 3.4105
R14715 GNDA.n2455 GNDA.n1915 3.4105
R14716 GNDA.n1956 GNDA.n1915 3.4105
R14717 GNDA.n2457 GNDA.n1915 3.4105
R14718 GNDA.n1955 GNDA.n1915 3.4105
R14719 GNDA.n2459 GNDA.n1915 3.4105
R14720 GNDA.n1954 GNDA.n1915 3.4105
R14721 GNDA.n2461 GNDA.n1915 3.4105
R14722 GNDA.n1953 GNDA.n1915 3.4105
R14723 GNDA.n2463 GNDA.n1915 3.4105
R14724 GNDA.n1952 GNDA.n1915 3.4105
R14725 GNDA.n2465 GNDA.n1915 3.4105
R14726 GNDA.n2467 GNDA.n1915 3.4105
R14727 GNDA.n1926 GNDA.n1901 3.4105
R14728 GNDA.n2435 GNDA.n1926 3.4105
R14729 GNDA.n1966 GNDA.n1926 3.4105
R14730 GNDA.n2437 GNDA.n1926 3.4105
R14731 GNDA.n1965 GNDA.n1926 3.4105
R14732 GNDA.n2439 GNDA.n1926 3.4105
R14733 GNDA.n1964 GNDA.n1926 3.4105
R14734 GNDA.n2441 GNDA.n1926 3.4105
R14735 GNDA.n1963 GNDA.n1926 3.4105
R14736 GNDA.n2443 GNDA.n1926 3.4105
R14737 GNDA.n1962 GNDA.n1926 3.4105
R14738 GNDA.n2445 GNDA.n1926 3.4105
R14739 GNDA.n1961 GNDA.n1926 3.4105
R14740 GNDA.n2447 GNDA.n1926 3.4105
R14741 GNDA.n1960 GNDA.n1926 3.4105
R14742 GNDA.n2449 GNDA.n1926 3.4105
R14743 GNDA.n1959 GNDA.n1926 3.4105
R14744 GNDA.n2451 GNDA.n1926 3.4105
R14745 GNDA.n1958 GNDA.n1926 3.4105
R14746 GNDA.n2453 GNDA.n1926 3.4105
R14747 GNDA.n1957 GNDA.n1926 3.4105
R14748 GNDA.n2455 GNDA.n1926 3.4105
R14749 GNDA.n1956 GNDA.n1926 3.4105
R14750 GNDA.n2457 GNDA.n1926 3.4105
R14751 GNDA.n1955 GNDA.n1926 3.4105
R14752 GNDA.n2459 GNDA.n1926 3.4105
R14753 GNDA.n1954 GNDA.n1926 3.4105
R14754 GNDA.n2461 GNDA.n1926 3.4105
R14755 GNDA.n1953 GNDA.n1926 3.4105
R14756 GNDA.n2463 GNDA.n1926 3.4105
R14757 GNDA.n1952 GNDA.n1926 3.4105
R14758 GNDA.n2465 GNDA.n1926 3.4105
R14759 GNDA.n2467 GNDA.n1926 3.4105
R14760 GNDA.n1914 GNDA.n1901 3.4105
R14761 GNDA.n2435 GNDA.n1914 3.4105
R14762 GNDA.n1966 GNDA.n1914 3.4105
R14763 GNDA.n2437 GNDA.n1914 3.4105
R14764 GNDA.n1965 GNDA.n1914 3.4105
R14765 GNDA.n2439 GNDA.n1914 3.4105
R14766 GNDA.n1964 GNDA.n1914 3.4105
R14767 GNDA.n2441 GNDA.n1914 3.4105
R14768 GNDA.n1963 GNDA.n1914 3.4105
R14769 GNDA.n2443 GNDA.n1914 3.4105
R14770 GNDA.n1962 GNDA.n1914 3.4105
R14771 GNDA.n2445 GNDA.n1914 3.4105
R14772 GNDA.n1961 GNDA.n1914 3.4105
R14773 GNDA.n2447 GNDA.n1914 3.4105
R14774 GNDA.n1960 GNDA.n1914 3.4105
R14775 GNDA.n2449 GNDA.n1914 3.4105
R14776 GNDA.n1959 GNDA.n1914 3.4105
R14777 GNDA.n2451 GNDA.n1914 3.4105
R14778 GNDA.n1958 GNDA.n1914 3.4105
R14779 GNDA.n2453 GNDA.n1914 3.4105
R14780 GNDA.n1957 GNDA.n1914 3.4105
R14781 GNDA.n2455 GNDA.n1914 3.4105
R14782 GNDA.n1956 GNDA.n1914 3.4105
R14783 GNDA.n2457 GNDA.n1914 3.4105
R14784 GNDA.n1955 GNDA.n1914 3.4105
R14785 GNDA.n2459 GNDA.n1914 3.4105
R14786 GNDA.n1954 GNDA.n1914 3.4105
R14787 GNDA.n2461 GNDA.n1914 3.4105
R14788 GNDA.n1953 GNDA.n1914 3.4105
R14789 GNDA.n2463 GNDA.n1914 3.4105
R14790 GNDA.n1952 GNDA.n1914 3.4105
R14791 GNDA.n2465 GNDA.n1914 3.4105
R14792 GNDA.n2467 GNDA.n1914 3.4105
R14793 GNDA.n1928 GNDA.n1901 3.4105
R14794 GNDA.n2435 GNDA.n1928 3.4105
R14795 GNDA.n1966 GNDA.n1928 3.4105
R14796 GNDA.n2437 GNDA.n1928 3.4105
R14797 GNDA.n1965 GNDA.n1928 3.4105
R14798 GNDA.n2439 GNDA.n1928 3.4105
R14799 GNDA.n1964 GNDA.n1928 3.4105
R14800 GNDA.n2441 GNDA.n1928 3.4105
R14801 GNDA.n1963 GNDA.n1928 3.4105
R14802 GNDA.n2443 GNDA.n1928 3.4105
R14803 GNDA.n1962 GNDA.n1928 3.4105
R14804 GNDA.n2445 GNDA.n1928 3.4105
R14805 GNDA.n1961 GNDA.n1928 3.4105
R14806 GNDA.n2447 GNDA.n1928 3.4105
R14807 GNDA.n1960 GNDA.n1928 3.4105
R14808 GNDA.n2449 GNDA.n1928 3.4105
R14809 GNDA.n1959 GNDA.n1928 3.4105
R14810 GNDA.n2451 GNDA.n1928 3.4105
R14811 GNDA.n1958 GNDA.n1928 3.4105
R14812 GNDA.n2453 GNDA.n1928 3.4105
R14813 GNDA.n1957 GNDA.n1928 3.4105
R14814 GNDA.n2455 GNDA.n1928 3.4105
R14815 GNDA.n1956 GNDA.n1928 3.4105
R14816 GNDA.n2457 GNDA.n1928 3.4105
R14817 GNDA.n1955 GNDA.n1928 3.4105
R14818 GNDA.n2459 GNDA.n1928 3.4105
R14819 GNDA.n1954 GNDA.n1928 3.4105
R14820 GNDA.n2461 GNDA.n1928 3.4105
R14821 GNDA.n1953 GNDA.n1928 3.4105
R14822 GNDA.n2463 GNDA.n1928 3.4105
R14823 GNDA.n1952 GNDA.n1928 3.4105
R14824 GNDA.n2465 GNDA.n1928 3.4105
R14825 GNDA.n2467 GNDA.n1928 3.4105
R14826 GNDA.n1913 GNDA.n1901 3.4105
R14827 GNDA.n2435 GNDA.n1913 3.4105
R14828 GNDA.n1966 GNDA.n1913 3.4105
R14829 GNDA.n2437 GNDA.n1913 3.4105
R14830 GNDA.n1965 GNDA.n1913 3.4105
R14831 GNDA.n2439 GNDA.n1913 3.4105
R14832 GNDA.n1964 GNDA.n1913 3.4105
R14833 GNDA.n2441 GNDA.n1913 3.4105
R14834 GNDA.n1963 GNDA.n1913 3.4105
R14835 GNDA.n2443 GNDA.n1913 3.4105
R14836 GNDA.n1962 GNDA.n1913 3.4105
R14837 GNDA.n2445 GNDA.n1913 3.4105
R14838 GNDA.n1961 GNDA.n1913 3.4105
R14839 GNDA.n2447 GNDA.n1913 3.4105
R14840 GNDA.n1960 GNDA.n1913 3.4105
R14841 GNDA.n2449 GNDA.n1913 3.4105
R14842 GNDA.n1959 GNDA.n1913 3.4105
R14843 GNDA.n2451 GNDA.n1913 3.4105
R14844 GNDA.n1958 GNDA.n1913 3.4105
R14845 GNDA.n2453 GNDA.n1913 3.4105
R14846 GNDA.n1957 GNDA.n1913 3.4105
R14847 GNDA.n2455 GNDA.n1913 3.4105
R14848 GNDA.n1956 GNDA.n1913 3.4105
R14849 GNDA.n2457 GNDA.n1913 3.4105
R14850 GNDA.n1955 GNDA.n1913 3.4105
R14851 GNDA.n2459 GNDA.n1913 3.4105
R14852 GNDA.n1954 GNDA.n1913 3.4105
R14853 GNDA.n2461 GNDA.n1913 3.4105
R14854 GNDA.n1953 GNDA.n1913 3.4105
R14855 GNDA.n2463 GNDA.n1913 3.4105
R14856 GNDA.n1952 GNDA.n1913 3.4105
R14857 GNDA.n2465 GNDA.n1913 3.4105
R14858 GNDA.n2467 GNDA.n1913 3.4105
R14859 GNDA.n1930 GNDA.n1901 3.4105
R14860 GNDA.n2435 GNDA.n1930 3.4105
R14861 GNDA.n1966 GNDA.n1930 3.4105
R14862 GNDA.n2437 GNDA.n1930 3.4105
R14863 GNDA.n1965 GNDA.n1930 3.4105
R14864 GNDA.n2439 GNDA.n1930 3.4105
R14865 GNDA.n1964 GNDA.n1930 3.4105
R14866 GNDA.n2441 GNDA.n1930 3.4105
R14867 GNDA.n1963 GNDA.n1930 3.4105
R14868 GNDA.n2443 GNDA.n1930 3.4105
R14869 GNDA.n1962 GNDA.n1930 3.4105
R14870 GNDA.n2445 GNDA.n1930 3.4105
R14871 GNDA.n1961 GNDA.n1930 3.4105
R14872 GNDA.n2447 GNDA.n1930 3.4105
R14873 GNDA.n1960 GNDA.n1930 3.4105
R14874 GNDA.n2449 GNDA.n1930 3.4105
R14875 GNDA.n1959 GNDA.n1930 3.4105
R14876 GNDA.n2451 GNDA.n1930 3.4105
R14877 GNDA.n1958 GNDA.n1930 3.4105
R14878 GNDA.n2453 GNDA.n1930 3.4105
R14879 GNDA.n1957 GNDA.n1930 3.4105
R14880 GNDA.n2455 GNDA.n1930 3.4105
R14881 GNDA.n1956 GNDA.n1930 3.4105
R14882 GNDA.n2457 GNDA.n1930 3.4105
R14883 GNDA.n1955 GNDA.n1930 3.4105
R14884 GNDA.n2459 GNDA.n1930 3.4105
R14885 GNDA.n1954 GNDA.n1930 3.4105
R14886 GNDA.n2461 GNDA.n1930 3.4105
R14887 GNDA.n1953 GNDA.n1930 3.4105
R14888 GNDA.n2463 GNDA.n1930 3.4105
R14889 GNDA.n1952 GNDA.n1930 3.4105
R14890 GNDA.n2465 GNDA.n1930 3.4105
R14891 GNDA.n2467 GNDA.n1930 3.4105
R14892 GNDA.n1912 GNDA.n1901 3.4105
R14893 GNDA.n2435 GNDA.n1912 3.4105
R14894 GNDA.n1966 GNDA.n1912 3.4105
R14895 GNDA.n2437 GNDA.n1912 3.4105
R14896 GNDA.n1965 GNDA.n1912 3.4105
R14897 GNDA.n2439 GNDA.n1912 3.4105
R14898 GNDA.n1964 GNDA.n1912 3.4105
R14899 GNDA.n2441 GNDA.n1912 3.4105
R14900 GNDA.n1963 GNDA.n1912 3.4105
R14901 GNDA.n2443 GNDA.n1912 3.4105
R14902 GNDA.n1962 GNDA.n1912 3.4105
R14903 GNDA.n2445 GNDA.n1912 3.4105
R14904 GNDA.n1961 GNDA.n1912 3.4105
R14905 GNDA.n2447 GNDA.n1912 3.4105
R14906 GNDA.n1960 GNDA.n1912 3.4105
R14907 GNDA.n2449 GNDA.n1912 3.4105
R14908 GNDA.n1959 GNDA.n1912 3.4105
R14909 GNDA.n2451 GNDA.n1912 3.4105
R14910 GNDA.n1958 GNDA.n1912 3.4105
R14911 GNDA.n2453 GNDA.n1912 3.4105
R14912 GNDA.n1957 GNDA.n1912 3.4105
R14913 GNDA.n2455 GNDA.n1912 3.4105
R14914 GNDA.n1956 GNDA.n1912 3.4105
R14915 GNDA.n2457 GNDA.n1912 3.4105
R14916 GNDA.n1955 GNDA.n1912 3.4105
R14917 GNDA.n2459 GNDA.n1912 3.4105
R14918 GNDA.n1954 GNDA.n1912 3.4105
R14919 GNDA.n2461 GNDA.n1912 3.4105
R14920 GNDA.n1953 GNDA.n1912 3.4105
R14921 GNDA.n2463 GNDA.n1912 3.4105
R14922 GNDA.n1952 GNDA.n1912 3.4105
R14923 GNDA.n2465 GNDA.n1912 3.4105
R14924 GNDA.n2467 GNDA.n1912 3.4105
R14925 GNDA.n1932 GNDA.n1901 3.4105
R14926 GNDA.n2435 GNDA.n1932 3.4105
R14927 GNDA.n1966 GNDA.n1932 3.4105
R14928 GNDA.n2437 GNDA.n1932 3.4105
R14929 GNDA.n1965 GNDA.n1932 3.4105
R14930 GNDA.n2439 GNDA.n1932 3.4105
R14931 GNDA.n1964 GNDA.n1932 3.4105
R14932 GNDA.n2441 GNDA.n1932 3.4105
R14933 GNDA.n1963 GNDA.n1932 3.4105
R14934 GNDA.n2443 GNDA.n1932 3.4105
R14935 GNDA.n1962 GNDA.n1932 3.4105
R14936 GNDA.n2445 GNDA.n1932 3.4105
R14937 GNDA.n1961 GNDA.n1932 3.4105
R14938 GNDA.n2447 GNDA.n1932 3.4105
R14939 GNDA.n1960 GNDA.n1932 3.4105
R14940 GNDA.n2449 GNDA.n1932 3.4105
R14941 GNDA.n1959 GNDA.n1932 3.4105
R14942 GNDA.n2451 GNDA.n1932 3.4105
R14943 GNDA.n1958 GNDA.n1932 3.4105
R14944 GNDA.n2453 GNDA.n1932 3.4105
R14945 GNDA.n1957 GNDA.n1932 3.4105
R14946 GNDA.n2455 GNDA.n1932 3.4105
R14947 GNDA.n1956 GNDA.n1932 3.4105
R14948 GNDA.n2457 GNDA.n1932 3.4105
R14949 GNDA.n1955 GNDA.n1932 3.4105
R14950 GNDA.n2459 GNDA.n1932 3.4105
R14951 GNDA.n1954 GNDA.n1932 3.4105
R14952 GNDA.n2461 GNDA.n1932 3.4105
R14953 GNDA.n1953 GNDA.n1932 3.4105
R14954 GNDA.n2463 GNDA.n1932 3.4105
R14955 GNDA.n1952 GNDA.n1932 3.4105
R14956 GNDA.n2465 GNDA.n1932 3.4105
R14957 GNDA.n2467 GNDA.n1932 3.4105
R14958 GNDA.n1911 GNDA.n1901 3.4105
R14959 GNDA.n2435 GNDA.n1911 3.4105
R14960 GNDA.n1966 GNDA.n1911 3.4105
R14961 GNDA.n2437 GNDA.n1911 3.4105
R14962 GNDA.n1965 GNDA.n1911 3.4105
R14963 GNDA.n2439 GNDA.n1911 3.4105
R14964 GNDA.n1964 GNDA.n1911 3.4105
R14965 GNDA.n2441 GNDA.n1911 3.4105
R14966 GNDA.n1963 GNDA.n1911 3.4105
R14967 GNDA.n2443 GNDA.n1911 3.4105
R14968 GNDA.n1962 GNDA.n1911 3.4105
R14969 GNDA.n2445 GNDA.n1911 3.4105
R14970 GNDA.n1961 GNDA.n1911 3.4105
R14971 GNDA.n2447 GNDA.n1911 3.4105
R14972 GNDA.n1960 GNDA.n1911 3.4105
R14973 GNDA.n2449 GNDA.n1911 3.4105
R14974 GNDA.n1959 GNDA.n1911 3.4105
R14975 GNDA.n2451 GNDA.n1911 3.4105
R14976 GNDA.n1958 GNDA.n1911 3.4105
R14977 GNDA.n2453 GNDA.n1911 3.4105
R14978 GNDA.n1957 GNDA.n1911 3.4105
R14979 GNDA.n2455 GNDA.n1911 3.4105
R14980 GNDA.n1956 GNDA.n1911 3.4105
R14981 GNDA.n2457 GNDA.n1911 3.4105
R14982 GNDA.n1955 GNDA.n1911 3.4105
R14983 GNDA.n2459 GNDA.n1911 3.4105
R14984 GNDA.n1954 GNDA.n1911 3.4105
R14985 GNDA.n2461 GNDA.n1911 3.4105
R14986 GNDA.n1953 GNDA.n1911 3.4105
R14987 GNDA.n2463 GNDA.n1911 3.4105
R14988 GNDA.n1952 GNDA.n1911 3.4105
R14989 GNDA.n2465 GNDA.n1911 3.4105
R14990 GNDA.n2467 GNDA.n1911 3.4105
R14991 GNDA.n1934 GNDA.n1901 3.4105
R14992 GNDA.n2435 GNDA.n1934 3.4105
R14993 GNDA.n1966 GNDA.n1934 3.4105
R14994 GNDA.n2437 GNDA.n1934 3.4105
R14995 GNDA.n1965 GNDA.n1934 3.4105
R14996 GNDA.n2439 GNDA.n1934 3.4105
R14997 GNDA.n1964 GNDA.n1934 3.4105
R14998 GNDA.n2441 GNDA.n1934 3.4105
R14999 GNDA.n1963 GNDA.n1934 3.4105
R15000 GNDA.n2443 GNDA.n1934 3.4105
R15001 GNDA.n1962 GNDA.n1934 3.4105
R15002 GNDA.n2445 GNDA.n1934 3.4105
R15003 GNDA.n1961 GNDA.n1934 3.4105
R15004 GNDA.n2447 GNDA.n1934 3.4105
R15005 GNDA.n1960 GNDA.n1934 3.4105
R15006 GNDA.n2449 GNDA.n1934 3.4105
R15007 GNDA.n1959 GNDA.n1934 3.4105
R15008 GNDA.n2451 GNDA.n1934 3.4105
R15009 GNDA.n1958 GNDA.n1934 3.4105
R15010 GNDA.n2453 GNDA.n1934 3.4105
R15011 GNDA.n1957 GNDA.n1934 3.4105
R15012 GNDA.n2455 GNDA.n1934 3.4105
R15013 GNDA.n1956 GNDA.n1934 3.4105
R15014 GNDA.n2457 GNDA.n1934 3.4105
R15015 GNDA.n1955 GNDA.n1934 3.4105
R15016 GNDA.n2459 GNDA.n1934 3.4105
R15017 GNDA.n1954 GNDA.n1934 3.4105
R15018 GNDA.n2461 GNDA.n1934 3.4105
R15019 GNDA.n1953 GNDA.n1934 3.4105
R15020 GNDA.n2463 GNDA.n1934 3.4105
R15021 GNDA.n1952 GNDA.n1934 3.4105
R15022 GNDA.n2465 GNDA.n1934 3.4105
R15023 GNDA.n2467 GNDA.n1934 3.4105
R15024 GNDA.n1910 GNDA.n1901 3.4105
R15025 GNDA.n2435 GNDA.n1910 3.4105
R15026 GNDA.n1966 GNDA.n1910 3.4105
R15027 GNDA.n2437 GNDA.n1910 3.4105
R15028 GNDA.n1965 GNDA.n1910 3.4105
R15029 GNDA.n2439 GNDA.n1910 3.4105
R15030 GNDA.n1964 GNDA.n1910 3.4105
R15031 GNDA.n2441 GNDA.n1910 3.4105
R15032 GNDA.n1963 GNDA.n1910 3.4105
R15033 GNDA.n2443 GNDA.n1910 3.4105
R15034 GNDA.n1962 GNDA.n1910 3.4105
R15035 GNDA.n2445 GNDA.n1910 3.4105
R15036 GNDA.n1961 GNDA.n1910 3.4105
R15037 GNDA.n2447 GNDA.n1910 3.4105
R15038 GNDA.n1960 GNDA.n1910 3.4105
R15039 GNDA.n2449 GNDA.n1910 3.4105
R15040 GNDA.n1959 GNDA.n1910 3.4105
R15041 GNDA.n2451 GNDA.n1910 3.4105
R15042 GNDA.n1958 GNDA.n1910 3.4105
R15043 GNDA.n2453 GNDA.n1910 3.4105
R15044 GNDA.n1957 GNDA.n1910 3.4105
R15045 GNDA.n2455 GNDA.n1910 3.4105
R15046 GNDA.n1956 GNDA.n1910 3.4105
R15047 GNDA.n2457 GNDA.n1910 3.4105
R15048 GNDA.n1955 GNDA.n1910 3.4105
R15049 GNDA.n2459 GNDA.n1910 3.4105
R15050 GNDA.n1954 GNDA.n1910 3.4105
R15051 GNDA.n2461 GNDA.n1910 3.4105
R15052 GNDA.n1953 GNDA.n1910 3.4105
R15053 GNDA.n2463 GNDA.n1910 3.4105
R15054 GNDA.n1952 GNDA.n1910 3.4105
R15055 GNDA.n2465 GNDA.n1910 3.4105
R15056 GNDA.n2467 GNDA.n1910 3.4105
R15057 GNDA.n1936 GNDA.n1901 3.4105
R15058 GNDA.n2435 GNDA.n1936 3.4105
R15059 GNDA.n1966 GNDA.n1936 3.4105
R15060 GNDA.n2437 GNDA.n1936 3.4105
R15061 GNDA.n1965 GNDA.n1936 3.4105
R15062 GNDA.n2439 GNDA.n1936 3.4105
R15063 GNDA.n1964 GNDA.n1936 3.4105
R15064 GNDA.n2441 GNDA.n1936 3.4105
R15065 GNDA.n1963 GNDA.n1936 3.4105
R15066 GNDA.n2443 GNDA.n1936 3.4105
R15067 GNDA.n1962 GNDA.n1936 3.4105
R15068 GNDA.n2445 GNDA.n1936 3.4105
R15069 GNDA.n1961 GNDA.n1936 3.4105
R15070 GNDA.n2447 GNDA.n1936 3.4105
R15071 GNDA.n1960 GNDA.n1936 3.4105
R15072 GNDA.n2449 GNDA.n1936 3.4105
R15073 GNDA.n1959 GNDA.n1936 3.4105
R15074 GNDA.n2451 GNDA.n1936 3.4105
R15075 GNDA.n1958 GNDA.n1936 3.4105
R15076 GNDA.n2453 GNDA.n1936 3.4105
R15077 GNDA.n1957 GNDA.n1936 3.4105
R15078 GNDA.n2455 GNDA.n1936 3.4105
R15079 GNDA.n1956 GNDA.n1936 3.4105
R15080 GNDA.n2457 GNDA.n1936 3.4105
R15081 GNDA.n1955 GNDA.n1936 3.4105
R15082 GNDA.n2459 GNDA.n1936 3.4105
R15083 GNDA.n1954 GNDA.n1936 3.4105
R15084 GNDA.n2461 GNDA.n1936 3.4105
R15085 GNDA.n1953 GNDA.n1936 3.4105
R15086 GNDA.n2463 GNDA.n1936 3.4105
R15087 GNDA.n1952 GNDA.n1936 3.4105
R15088 GNDA.n2465 GNDA.n1936 3.4105
R15089 GNDA.n2467 GNDA.n1936 3.4105
R15090 GNDA.n1909 GNDA.n1901 3.4105
R15091 GNDA.n2435 GNDA.n1909 3.4105
R15092 GNDA.n1966 GNDA.n1909 3.4105
R15093 GNDA.n2437 GNDA.n1909 3.4105
R15094 GNDA.n1965 GNDA.n1909 3.4105
R15095 GNDA.n2439 GNDA.n1909 3.4105
R15096 GNDA.n1964 GNDA.n1909 3.4105
R15097 GNDA.n2441 GNDA.n1909 3.4105
R15098 GNDA.n1963 GNDA.n1909 3.4105
R15099 GNDA.n2443 GNDA.n1909 3.4105
R15100 GNDA.n1962 GNDA.n1909 3.4105
R15101 GNDA.n2445 GNDA.n1909 3.4105
R15102 GNDA.n1961 GNDA.n1909 3.4105
R15103 GNDA.n2447 GNDA.n1909 3.4105
R15104 GNDA.n1960 GNDA.n1909 3.4105
R15105 GNDA.n2449 GNDA.n1909 3.4105
R15106 GNDA.n1959 GNDA.n1909 3.4105
R15107 GNDA.n2451 GNDA.n1909 3.4105
R15108 GNDA.n1958 GNDA.n1909 3.4105
R15109 GNDA.n2453 GNDA.n1909 3.4105
R15110 GNDA.n1957 GNDA.n1909 3.4105
R15111 GNDA.n2455 GNDA.n1909 3.4105
R15112 GNDA.n1956 GNDA.n1909 3.4105
R15113 GNDA.n2457 GNDA.n1909 3.4105
R15114 GNDA.n1955 GNDA.n1909 3.4105
R15115 GNDA.n2459 GNDA.n1909 3.4105
R15116 GNDA.n1954 GNDA.n1909 3.4105
R15117 GNDA.n2461 GNDA.n1909 3.4105
R15118 GNDA.n1953 GNDA.n1909 3.4105
R15119 GNDA.n2463 GNDA.n1909 3.4105
R15120 GNDA.n1952 GNDA.n1909 3.4105
R15121 GNDA.n2465 GNDA.n1909 3.4105
R15122 GNDA.n2467 GNDA.n1909 3.4105
R15123 GNDA.n1938 GNDA.n1901 3.4105
R15124 GNDA.n2435 GNDA.n1938 3.4105
R15125 GNDA.n1966 GNDA.n1938 3.4105
R15126 GNDA.n2437 GNDA.n1938 3.4105
R15127 GNDA.n1965 GNDA.n1938 3.4105
R15128 GNDA.n2439 GNDA.n1938 3.4105
R15129 GNDA.n1964 GNDA.n1938 3.4105
R15130 GNDA.n2441 GNDA.n1938 3.4105
R15131 GNDA.n1963 GNDA.n1938 3.4105
R15132 GNDA.n2443 GNDA.n1938 3.4105
R15133 GNDA.n1962 GNDA.n1938 3.4105
R15134 GNDA.n2445 GNDA.n1938 3.4105
R15135 GNDA.n1961 GNDA.n1938 3.4105
R15136 GNDA.n2447 GNDA.n1938 3.4105
R15137 GNDA.n1960 GNDA.n1938 3.4105
R15138 GNDA.n2449 GNDA.n1938 3.4105
R15139 GNDA.n1959 GNDA.n1938 3.4105
R15140 GNDA.n2451 GNDA.n1938 3.4105
R15141 GNDA.n1958 GNDA.n1938 3.4105
R15142 GNDA.n2453 GNDA.n1938 3.4105
R15143 GNDA.n1957 GNDA.n1938 3.4105
R15144 GNDA.n2455 GNDA.n1938 3.4105
R15145 GNDA.n1956 GNDA.n1938 3.4105
R15146 GNDA.n2457 GNDA.n1938 3.4105
R15147 GNDA.n1955 GNDA.n1938 3.4105
R15148 GNDA.n2459 GNDA.n1938 3.4105
R15149 GNDA.n1954 GNDA.n1938 3.4105
R15150 GNDA.n2461 GNDA.n1938 3.4105
R15151 GNDA.n1953 GNDA.n1938 3.4105
R15152 GNDA.n2463 GNDA.n1938 3.4105
R15153 GNDA.n1952 GNDA.n1938 3.4105
R15154 GNDA.n2465 GNDA.n1938 3.4105
R15155 GNDA.n2467 GNDA.n1938 3.4105
R15156 GNDA.n1908 GNDA.n1901 3.4105
R15157 GNDA.n2435 GNDA.n1908 3.4105
R15158 GNDA.n1966 GNDA.n1908 3.4105
R15159 GNDA.n2437 GNDA.n1908 3.4105
R15160 GNDA.n1965 GNDA.n1908 3.4105
R15161 GNDA.n2439 GNDA.n1908 3.4105
R15162 GNDA.n1964 GNDA.n1908 3.4105
R15163 GNDA.n2441 GNDA.n1908 3.4105
R15164 GNDA.n1963 GNDA.n1908 3.4105
R15165 GNDA.n2443 GNDA.n1908 3.4105
R15166 GNDA.n1962 GNDA.n1908 3.4105
R15167 GNDA.n2445 GNDA.n1908 3.4105
R15168 GNDA.n1961 GNDA.n1908 3.4105
R15169 GNDA.n2447 GNDA.n1908 3.4105
R15170 GNDA.n1960 GNDA.n1908 3.4105
R15171 GNDA.n2449 GNDA.n1908 3.4105
R15172 GNDA.n1959 GNDA.n1908 3.4105
R15173 GNDA.n2451 GNDA.n1908 3.4105
R15174 GNDA.n1958 GNDA.n1908 3.4105
R15175 GNDA.n2453 GNDA.n1908 3.4105
R15176 GNDA.n1957 GNDA.n1908 3.4105
R15177 GNDA.n2455 GNDA.n1908 3.4105
R15178 GNDA.n1956 GNDA.n1908 3.4105
R15179 GNDA.n2457 GNDA.n1908 3.4105
R15180 GNDA.n1955 GNDA.n1908 3.4105
R15181 GNDA.n2459 GNDA.n1908 3.4105
R15182 GNDA.n1954 GNDA.n1908 3.4105
R15183 GNDA.n2461 GNDA.n1908 3.4105
R15184 GNDA.n1953 GNDA.n1908 3.4105
R15185 GNDA.n2463 GNDA.n1908 3.4105
R15186 GNDA.n1952 GNDA.n1908 3.4105
R15187 GNDA.n2465 GNDA.n1908 3.4105
R15188 GNDA.n2467 GNDA.n1908 3.4105
R15189 GNDA.n1940 GNDA.n1901 3.4105
R15190 GNDA.n2435 GNDA.n1940 3.4105
R15191 GNDA.n1966 GNDA.n1940 3.4105
R15192 GNDA.n2437 GNDA.n1940 3.4105
R15193 GNDA.n1965 GNDA.n1940 3.4105
R15194 GNDA.n2439 GNDA.n1940 3.4105
R15195 GNDA.n1964 GNDA.n1940 3.4105
R15196 GNDA.n2441 GNDA.n1940 3.4105
R15197 GNDA.n1963 GNDA.n1940 3.4105
R15198 GNDA.n2443 GNDA.n1940 3.4105
R15199 GNDA.n1962 GNDA.n1940 3.4105
R15200 GNDA.n2445 GNDA.n1940 3.4105
R15201 GNDA.n1961 GNDA.n1940 3.4105
R15202 GNDA.n2447 GNDA.n1940 3.4105
R15203 GNDA.n1960 GNDA.n1940 3.4105
R15204 GNDA.n2449 GNDA.n1940 3.4105
R15205 GNDA.n1959 GNDA.n1940 3.4105
R15206 GNDA.n2451 GNDA.n1940 3.4105
R15207 GNDA.n1958 GNDA.n1940 3.4105
R15208 GNDA.n2453 GNDA.n1940 3.4105
R15209 GNDA.n1957 GNDA.n1940 3.4105
R15210 GNDA.n2455 GNDA.n1940 3.4105
R15211 GNDA.n1956 GNDA.n1940 3.4105
R15212 GNDA.n2457 GNDA.n1940 3.4105
R15213 GNDA.n1955 GNDA.n1940 3.4105
R15214 GNDA.n2459 GNDA.n1940 3.4105
R15215 GNDA.n1954 GNDA.n1940 3.4105
R15216 GNDA.n2461 GNDA.n1940 3.4105
R15217 GNDA.n1953 GNDA.n1940 3.4105
R15218 GNDA.n2463 GNDA.n1940 3.4105
R15219 GNDA.n1952 GNDA.n1940 3.4105
R15220 GNDA.n2465 GNDA.n1940 3.4105
R15221 GNDA.n2467 GNDA.n1940 3.4105
R15222 GNDA.n1907 GNDA.n1901 3.4105
R15223 GNDA.n2435 GNDA.n1907 3.4105
R15224 GNDA.n1966 GNDA.n1907 3.4105
R15225 GNDA.n2437 GNDA.n1907 3.4105
R15226 GNDA.n1965 GNDA.n1907 3.4105
R15227 GNDA.n2439 GNDA.n1907 3.4105
R15228 GNDA.n1964 GNDA.n1907 3.4105
R15229 GNDA.n2441 GNDA.n1907 3.4105
R15230 GNDA.n1963 GNDA.n1907 3.4105
R15231 GNDA.n2443 GNDA.n1907 3.4105
R15232 GNDA.n1962 GNDA.n1907 3.4105
R15233 GNDA.n2445 GNDA.n1907 3.4105
R15234 GNDA.n1961 GNDA.n1907 3.4105
R15235 GNDA.n2447 GNDA.n1907 3.4105
R15236 GNDA.n1960 GNDA.n1907 3.4105
R15237 GNDA.n2449 GNDA.n1907 3.4105
R15238 GNDA.n1959 GNDA.n1907 3.4105
R15239 GNDA.n2451 GNDA.n1907 3.4105
R15240 GNDA.n1958 GNDA.n1907 3.4105
R15241 GNDA.n2453 GNDA.n1907 3.4105
R15242 GNDA.n1957 GNDA.n1907 3.4105
R15243 GNDA.n2455 GNDA.n1907 3.4105
R15244 GNDA.n1956 GNDA.n1907 3.4105
R15245 GNDA.n2457 GNDA.n1907 3.4105
R15246 GNDA.n1955 GNDA.n1907 3.4105
R15247 GNDA.n2459 GNDA.n1907 3.4105
R15248 GNDA.n1954 GNDA.n1907 3.4105
R15249 GNDA.n2461 GNDA.n1907 3.4105
R15250 GNDA.n1953 GNDA.n1907 3.4105
R15251 GNDA.n2463 GNDA.n1907 3.4105
R15252 GNDA.n1952 GNDA.n1907 3.4105
R15253 GNDA.n2465 GNDA.n1907 3.4105
R15254 GNDA.n2467 GNDA.n1907 3.4105
R15255 GNDA.n1942 GNDA.n1901 3.4105
R15256 GNDA.n2435 GNDA.n1942 3.4105
R15257 GNDA.n1966 GNDA.n1942 3.4105
R15258 GNDA.n2437 GNDA.n1942 3.4105
R15259 GNDA.n1965 GNDA.n1942 3.4105
R15260 GNDA.n2439 GNDA.n1942 3.4105
R15261 GNDA.n1964 GNDA.n1942 3.4105
R15262 GNDA.n2441 GNDA.n1942 3.4105
R15263 GNDA.n1963 GNDA.n1942 3.4105
R15264 GNDA.n2443 GNDA.n1942 3.4105
R15265 GNDA.n1962 GNDA.n1942 3.4105
R15266 GNDA.n2445 GNDA.n1942 3.4105
R15267 GNDA.n1961 GNDA.n1942 3.4105
R15268 GNDA.n2447 GNDA.n1942 3.4105
R15269 GNDA.n1960 GNDA.n1942 3.4105
R15270 GNDA.n2449 GNDA.n1942 3.4105
R15271 GNDA.n1959 GNDA.n1942 3.4105
R15272 GNDA.n2451 GNDA.n1942 3.4105
R15273 GNDA.n1958 GNDA.n1942 3.4105
R15274 GNDA.n2453 GNDA.n1942 3.4105
R15275 GNDA.n1957 GNDA.n1942 3.4105
R15276 GNDA.n2455 GNDA.n1942 3.4105
R15277 GNDA.n1956 GNDA.n1942 3.4105
R15278 GNDA.n2457 GNDA.n1942 3.4105
R15279 GNDA.n1955 GNDA.n1942 3.4105
R15280 GNDA.n2459 GNDA.n1942 3.4105
R15281 GNDA.n1954 GNDA.n1942 3.4105
R15282 GNDA.n2461 GNDA.n1942 3.4105
R15283 GNDA.n1953 GNDA.n1942 3.4105
R15284 GNDA.n2463 GNDA.n1942 3.4105
R15285 GNDA.n1952 GNDA.n1942 3.4105
R15286 GNDA.n2465 GNDA.n1942 3.4105
R15287 GNDA.n2467 GNDA.n1942 3.4105
R15288 GNDA.n1906 GNDA.n1901 3.4105
R15289 GNDA.n2435 GNDA.n1906 3.4105
R15290 GNDA.n1966 GNDA.n1906 3.4105
R15291 GNDA.n2437 GNDA.n1906 3.4105
R15292 GNDA.n1965 GNDA.n1906 3.4105
R15293 GNDA.n2439 GNDA.n1906 3.4105
R15294 GNDA.n1964 GNDA.n1906 3.4105
R15295 GNDA.n2441 GNDA.n1906 3.4105
R15296 GNDA.n1963 GNDA.n1906 3.4105
R15297 GNDA.n2443 GNDA.n1906 3.4105
R15298 GNDA.n1962 GNDA.n1906 3.4105
R15299 GNDA.n2445 GNDA.n1906 3.4105
R15300 GNDA.n1961 GNDA.n1906 3.4105
R15301 GNDA.n2447 GNDA.n1906 3.4105
R15302 GNDA.n1960 GNDA.n1906 3.4105
R15303 GNDA.n2449 GNDA.n1906 3.4105
R15304 GNDA.n1959 GNDA.n1906 3.4105
R15305 GNDA.n2451 GNDA.n1906 3.4105
R15306 GNDA.n1958 GNDA.n1906 3.4105
R15307 GNDA.n2453 GNDA.n1906 3.4105
R15308 GNDA.n1957 GNDA.n1906 3.4105
R15309 GNDA.n2455 GNDA.n1906 3.4105
R15310 GNDA.n1956 GNDA.n1906 3.4105
R15311 GNDA.n2457 GNDA.n1906 3.4105
R15312 GNDA.n1955 GNDA.n1906 3.4105
R15313 GNDA.n2459 GNDA.n1906 3.4105
R15314 GNDA.n1954 GNDA.n1906 3.4105
R15315 GNDA.n2461 GNDA.n1906 3.4105
R15316 GNDA.n1953 GNDA.n1906 3.4105
R15317 GNDA.n2463 GNDA.n1906 3.4105
R15318 GNDA.n1952 GNDA.n1906 3.4105
R15319 GNDA.n2465 GNDA.n1906 3.4105
R15320 GNDA.n2467 GNDA.n1906 3.4105
R15321 GNDA.n1944 GNDA.n1901 3.4105
R15322 GNDA.n2435 GNDA.n1944 3.4105
R15323 GNDA.n1966 GNDA.n1944 3.4105
R15324 GNDA.n2437 GNDA.n1944 3.4105
R15325 GNDA.n1965 GNDA.n1944 3.4105
R15326 GNDA.n2439 GNDA.n1944 3.4105
R15327 GNDA.n1964 GNDA.n1944 3.4105
R15328 GNDA.n2441 GNDA.n1944 3.4105
R15329 GNDA.n1963 GNDA.n1944 3.4105
R15330 GNDA.n2443 GNDA.n1944 3.4105
R15331 GNDA.n1962 GNDA.n1944 3.4105
R15332 GNDA.n2445 GNDA.n1944 3.4105
R15333 GNDA.n1961 GNDA.n1944 3.4105
R15334 GNDA.n2447 GNDA.n1944 3.4105
R15335 GNDA.n1960 GNDA.n1944 3.4105
R15336 GNDA.n2449 GNDA.n1944 3.4105
R15337 GNDA.n1959 GNDA.n1944 3.4105
R15338 GNDA.n2451 GNDA.n1944 3.4105
R15339 GNDA.n1958 GNDA.n1944 3.4105
R15340 GNDA.n2453 GNDA.n1944 3.4105
R15341 GNDA.n1957 GNDA.n1944 3.4105
R15342 GNDA.n2455 GNDA.n1944 3.4105
R15343 GNDA.n1956 GNDA.n1944 3.4105
R15344 GNDA.n2457 GNDA.n1944 3.4105
R15345 GNDA.n1955 GNDA.n1944 3.4105
R15346 GNDA.n2459 GNDA.n1944 3.4105
R15347 GNDA.n1954 GNDA.n1944 3.4105
R15348 GNDA.n2461 GNDA.n1944 3.4105
R15349 GNDA.n1953 GNDA.n1944 3.4105
R15350 GNDA.n2463 GNDA.n1944 3.4105
R15351 GNDA.n1952 GNDA.n1944 3.4105
R15352 GNDA.n2465 GNDA.n1944 3.4105
R15353 GNDA.n2467 GNDA.n1944 3.4105
R15354 GNDA.n1905 GNDA.n1901 3.4105
R15355 GNDA.n2435 GNDA.n1905 3.4105
R15356 GNDA.n1966 GNDA.n1905 3.4105
R15357 GNDA.n2437 GNDA.n1905 3.4105
R15358 GNDA.n1965 GNDA.n1905 3.4105
R15359 GNDA.n2439 GNDA.n1905 3.4105
R15360 GNDA.n1964 GNDA.n1905 3.4105
R15361 GNDA.n2441 GNDA.n1905 3.4105
R15362 GNDA.n1963 GNDA.n1905 3.4105
R15363 GNDA.n2443 GNDA.n1905 3.4105
R15364 GNDA.n1962 GNDA.n1905 3.4105
R15365 GNDA.n2445 GNDA.n1905 3.4105
R15366 GNDA.n1961 GNDA.n1905 3.4105
R15367 GNDA.n2447 GNDA.n1905 3.4105
R15368 GNDA.n1960 GNDA.n1905 3.4105
R15369 GNDA.n2449 GNDA.n1905 3.4105
R15370 GNDA.n1959 GNDA.n1905 3.4105
R15371 GNDA.n2451 GNDA.n1905 3.4105
R15372 GNDA.n1958 GNDA.n1905 3.4105
R15373 GNDA.n2453 GNDA.n1905 3.4105
R15374 GNDA.n1957 GNDA.n1905 3.4105
R15375 GNDA.n2455 GNDA.n1905 3.4105
R15376 GNDA.n1956 GNDA.n1905 3.4105
R15377 GNDA.n2457 GNDA.n1905 3.4105
R15378 GNDA.n1955 GNDA.n1905 3.4105
R15379 GNDA.n2459 GNDA.n1905 3.4105
R15380 GNDA.n1954 GNDA.n1905 3.4105
R15381 GNDA.n2461 GNDA.n1905 3.4105
R15382 GNDA.n1953 GNDA.n1905 3.4105
R15383 GNDA.n2463 GNDA.n1905 3.4105
R15384 GNDA.n1952 GNDA.n1905 3.4105
R15385 GNDA.n2465 GNDA.n1905 3.4105
R15386 GNDA.n2467 GNDA.n1905 3.4105
R15387 GNDA.n1946 GNDA.n1901 3.4105
R15388 GNDA.n2435 GNDA.n1946 3.4105
R15389 GNDA.n1966 GNDA.n1946 3.4105
R15390 GNDA.n2437 GNDA.n1946 3.4105
R15391 GNDA.n1965 GNDA.n1946 3.4105
R15392 GNDA.n2439 GNDA.n1946 3.4105
R15393 GNDA.n1964 GNDA.n1946 3.4105
R15394 GNDA.n2441 GNDA.n1946 3.4105
R15395 GNDA.n1963 GNDA.n1946 3.4105
R15396 GNDA.n2443 GNDA.n1946 3.4105
R15397 GNDA.n1962 GNDA.n1946 3.4105
R15398 GNDA.n2445 GNDA.n1946 3.4105
R15399 GNDA.n1961 GNDA.n1946 3.4105
R15400 GNDA.n2447 GNDA.n1946 3.4105
R15401 GNDA.n1960 GNDA.n1946 3.4105
R15402 GNDA.n2449 GNDA.n1946 3.4105
R15403 GNDA.n1959 GNDA.n1946 3.4105
R15404 GNDA.n2451 GNDA.n1946 3.4105
R15405 GNDA.n1958 GNDA.n1946 3.4105
R15406 GNDA.n2453 GNDA.n1946 3.4105
R15407 GNDA.n1957 GNDA.n1946 3.4105
R15408 GNDA.n2455 GNDA.n1946 3.4105
R15409 GNDA.n1956 GNDA.n1946 3.4105
R15410 GNDA.n2457 GNDA.n1946 3.4105
R15411 GNDA.n1955 GNDA.n1946 3.4105
R15412 GNDA.n2459 GNDA.n1946 3.4105
R15413 GNDA.n1954 GNDA.n1946 3.4105
R15414 GNDA.n2461 GNDA.n1946 3.4105
R15415 GNDA.n1953 GNDA.n1946 3.4105
R15416 GNDA.n2463 GNDA.n1946 3.4105
R15417 GNDA.n1952 GNDA.n1946 3.4105
R15418 GNDA.n2465 GNDA.n1946 3.4105
R15419 GNDA.n2467 GNDA.n1946 3.4105
R15420 GNDA.n1904 GNDA.n1901 3.4105
R15421 GNDA.n2435 GNDA.n1904 3.4105
R15422 GNDA.n1966 GNDA.n1904 3.4105
R15423 GNDA.n2437 GNDA.n1904 3.4105
R15424 GNDA.n1965 GNDA.n1904 3.4105
R15425 GNDA.n2439 GNDA.n1904 3.4105
R15426 GNDA.n1964 GNDA.n1904 3.4105
R15427 GNDA.n2441 GNDA.n1904 3.4105
R15428 GNDA.n1963 GNDA.n1904 3.4105
R15429 GNDA.n2443 GNDA.n1904 3.4105
R15430 GNDA.n1962 GNDA.n1904 3.4105
R15431 GNDA.n2445 GNDA.n1904 3.4105
R15432 GNDA.n1961 GNDA.n1904 3.4105
R15433 GNDA.n2447 GNDA.n1904 3.4105
R15434 GNDA.n1960 GNDA.n1904 3.4105
R15435 GNDA.n2449 GNDA.n1904 3.4105
R15436 GNDA.n1959 GNDA.n1904 3.4105
R15437 GNDA.n2451 GNDA.n1904 3.4105
R15438 GNDA.n1958 GNDA.n1904 3.4105
R15439 GNDA.n2453 GNDA.n1904 3.4105
R15440 GNDA.n1957 GNDA.n1904 3.4105
R15441 GNDA.n2455 GNDA.n1904 3.4105
R15442 GNDA.n1956 GNDA.n1904 3.4105
R15443 GNDA.n2457 GNDA.n1904 3.4105
R15444 GNDA.n1955 GNDA.n1904 3.4105
R15445 GNDA.n2459 GNDA.n1904 3.4105
R15446 GNDA.n1954 GNDA.n1904 3.4105
R15447 GNDA.n2461 GNDA.n1904 3.4105
R15448 GNDA.n1953 GNDA.n1904 3.4105
R15449 GNDA.n2463 GNDA.n1904 3.4105
R15450 GNDA.n1952 GNDA.n1904 3.4105
R15451 GNDA.n2465 GNDA.n1904 3.4105
R15452 GNDA.n2467 GNDA.n1904 3.4105
R15453 GNDA.n1948 GNDA.n1901 3.4105
R15454 GNDA.n2435 GNDA.n1948 3.4105
R15455 GNDA.n1966 GNDA.n1948 3.4105
R15456 GNDA.n2437 GNDA.n1948 3.4105
R15457 GNDA.n1965 GNDA.n1948 3.4105
R15458 GNDA.n2439 GNDA.n1948 3.4105
R15459 GNDA.n1964 GNDA.n1948 3.4105
R15460 GNDA.n2441 GNDA.n1948 3.4105
R15461 GNDA.n1963 GNDA.n1948 3.4105
R15462 GNDA.n2443 GNDA.n1948 3.4105
R15463 GNDA.n1962 GNDA.n1948 3.4105
R15464 GNDA.n2445 GNDA.n1948 3.4105
R15465 GNDA.n1961 GNDA.n1948 3.4105
R15466 GNDA.n2447 GNDA.n1948 3.4105
R15467 GNDA.n1960 GNDA.n1948 3.4105
R15468 GNDA.n2449 GNDA.n1948 3.4105
R15469 GNDA.n1959 GNDA.n1948 3.4105
R15470 GNDA.n2451 GNDA.n1948 3.4105
R15471 GNDA.n1958 GNDA.n1948 3.4105
R15472 GNDA.n2453 GNDA.n1948 3.4105
R15473 GNDA.n1957 GNDA.n1948 3.4105
R15474 GNDA.n2455 GNDA.n1948 3.4105
R15475 GNDA.n1956 GNDA.n1948 3.4105
R15476 GNDA.n2457 GNDA.n1948 3.4105
R15477 GNDA.n1955 GNDA.n1948 3.4105
R15478 GNDA.n2459 GNDA.n1948 3.4105
R15479 GNDA.n1954 GNDA.n1948 3.4105
R15480 GNDA.n2461 GNDA.n1948 3.4105
R15481 GNDA.n1953 GNDA.n1948 3.4105
R15482 GNDA.n2463 GNDA.n1948 3.4105
R15483 GNDA.n1952 GNDA.n1948 3.4105
R15484 GNDA.n2465 GNDA.n1948 3.4105
R15485 GNDA.n2467 GNDA.n1948 3.4105
R15486 GNDA.n1903 GNDA.n1901 3.4105
R15487 GNDA.n2435 GNDA.n1903 3.4105
R15488 GNDA.n1966 GNDA.n1903 3.4105
R15489 GNDA.n2437 GNDA.n1903 3.4105
R15490 GNDA.n1965 GNDA.n1903 3.4105
R15491 GNDA.n2439 GNDA.n1903 3.4105
R15492 GNDA.n1964 GNDA.n1903 3.4105
R15493 GNDA.n2441 GNDA.n1903 3.4105
R15494 GNDA.n1963 GNDA.n1903 3.4105
R15495 GNDA.n2443 GNDA.n1903 3.4105
R15496 GNDA.n1962 GNDA.n1903 3.4105
R15497 GNDA.n2445 GNDA.n1903 3.4105
R15498 GNDA.n1961 GNDA.n1903 3.4105
R15499 GNDA.n2447 GNDA.n1903 3.4105
R15500 GNDA.n1960 GNDA.n1903 3.4105
R15501 GNDA.n2449 GNDA.n1903 3.4105
R15502 GNDA.n1959 GNDA.n1903 3.4105
R15503 GNDA.n2451 GNDA.n1903 3.4105
R15504 GNDA.n1958 GNDA.n1903 3.4105
R15505 GNDA.n2453 GNDA.n1903 3.4105
R15506 GNDA.n1957 GNDA.n1903 3.4105
R15507 GNDA.n2455 GNDA.n1903 3.4105
R15508 GNDA.n1956 GNDA.n1903 3.4105
R15509 GNDA.n2457 GNDA.n1903 3.4105
R15510 GNDA.n1955 GNDA.n1903 3.4105
R15511 GNDA.n2459 GNDA.n1903 3.4105
R15512 GNDA.n1954 GNDA.n1903 3.4105
R15513 GNDA.n2461 GNDA.n1903 3.4105
R15514 GNDA.n1953 GNDA.n1903 3.4105
R15515 GNDA.n2463 GNDA.n1903 3.4105
R15516 GNDA.n1952 GNDA.n1903 3.4105
R15517 GNDA.n2465 GNDA.n1903 3.4105
R15518 GNDA.n2467 GNDA.n1903 3.4105
R15519 GNDA.n1950 GNDA.n1901 3.4105
R15520 GNDA.n2435 GNDA.n1950 3.4105
R15521 GNDA.n1966 GNDA.n1950 3.4105
R15522 GNDA.n2437 GNDA.n1950 3.4105
R15523 GNDA.n1965 GNDA.n1950 3.4105
R15524 GNDA.n2439 GNDA.n1950 3.4105
R15525 GNDA.n1964 GNDA.n1950 3.4105
R15526 GNDA.n2441 GNDA.n1950 3.4105
R15527 GNDA.n1963 GNDA.n1950 3.4105
R15528 GNDA.n2443 GNDA.n1950 3.4105
R15529 GNDA.n1962 GNDA.n1950 3.4105
R15530 GNDA.n2445 GNDA.n1950 3.4105
R15531 GNDA.n1961 GNDA.n1950 3.4105
R15532 GNDA.n2447 GNDA.n1950 3.4105
R15533 GNDA.n1960 GNDA.n1950 3.4105
R15534 GNDA.n2449 GNDA.n1950 3.4105
R15535 GNDA.n1959 GNDA.n1950 3.4105
R15536 GNDA.n2451 GNDA.n1950 3.4105
R15537 GNDA.n1958 GNDA.n1950 3.4105
R15538 GNDA.n2453 GNDA.n1950 3.4105
R15539 GNDA.n1957 GNDA.n1950 3.4105
R15540 GNDA.n2455 GNDA.n1950 3.4105
R15541 GNDA.n1956 GNDA.n1950 3.4105
R15542 GNDA.n2457 GNDA.n1950 3.4105
R15543 GNDA.n1955 GNDA.n1950 3.4105
R15544 GNDA.n2459 GNDA.n1950 3.4105
R15545 GNDA.n1954 GNDA.n1950 3.4105
R15546 GNDA.n2461 GNDA.n1950 3.4105
R15547 GNDA.n1953 GNDA.n1950 3.4105
R15548 GNDA.n2463 GNDA.n1950 3.4105
R15549 GNDA.n1952 GNDA.n1950 3.4105
R15550 GNDA.n2465 GNDA.n1950 3.4105
R15551 GNDA.n2467 GNDA.n1950 3.4105
R15552 GNDA.n1902 GNDA.n1901 3.4105
R15553 GNDA.n2435 GNDA.n1902 3.4105
R15554 GNDA.n1966 GNDA.n1902 3.4105
R15555 GNDA.n2437 GNDA.n1902 3.4105
R15556 GNDA.n1965 GNDA.n1902 3.4105
R15557 GNDA.n2439 GNDA.n1902 3.4105
R15558 GNDA.n1964 GNDA.n1902 3.4105
R15559 GNDA.n2441 GNDA.n1902 3.4105
R15560 GNDA.n1963 GNDA.n1902 3.4105
R15561 GNDA.n2443 GNDA.n1902 3.4105
R15562 GNDA.n1962 GNDA.n1902 3.4105
R15563 GNDA.n2445 GNDA.n1902 3.4105
R15564 GNDA.n1961 GNDA.n1902 3.4105
R15565 GNDA.n2447 GNDA.n1902 3.4105
R15566 GNDA.n1960 GNDA.n1902 3.4105
R15567 GNDA.n2449 GNDA.n1902 3.4105
R15568 GNDA.n1959 GNDA.n1902 3.4105
R15569 GNDA.n2451 GNDA.n1902 3.4105
R15570 GNDA.n1958 GNDA.n1902 3.4105
R15571 GNDA.n2453 GNDA.n1902 3.4105
R15572 GNDA.n1957 GNDA.n1902 3.4105
R15573 GNDA.n2455 GNDA.n1902 3.4105
R15574 GNDA.n1956 GNDA.n1902 3.4105
R15575 GNDA.n2457 GNDA.n1902 3.4105
R15576 GNDA.n1955 GNDA.n1902 3.4105
R15577 GNDA.n2459 GNDA.n1902 3.4105
R15578 GNDA.n1954 GNDA.n1902 3.4105
R15579 GNDA.n2461 GNDA.n1902 3.4105
R15580 GNDA.n1953 GNDA.n1902 3.4105
R15581 GNDA.n2463 GNDA.n1902 3.4105
R15582 GNDA.n1952 GNDA.n1902 3.4105
R15583 GNDA.n2465 GNDA.n1902 3.4105
R15584 GNDA.n2467 GNDA.n1902 3.4105
R15585 GNDA.n2466 GNDA.n2435 3.4105
R15586 GNDA.n2466 GNDA.n1966 3.4105
R15587 GNDA.n2466 GNDA.n2437 3.4105
R15588 GNDA.n2466 GNDA.n1965 3.4105
R15589 GNDA.n2466 GNDA.n2439 3.4105
R15590 GNDA.n2466 GNDA.n1964 3.4105
R15591 GNDA.n2466 GNDA.n2441 3.4105
R15592 GNDA.n2466 GNDA.n1963 3.4105
R15593 GNDA.n2466 GNDA.n2443 3.4105
R15594 GNDA.n2466 GNDA.n1962 3.4105
R15595 GNDA.n2466 GNDA.n2445 3.4105
R15596 GNDA.n2466 GNDA.n1961 3.4105
R15597 GNDA.n2466 GNDA.n2447 3.4105
R15598 GNDA.n2466 GNDA.n1960 3.4105
R15599 GNDA.n2466 GNDA.n2449 3.4105
R15600 GNDA.n2466 GNDA.n1959 3.4105
R15601 GNDA.n2466 GNDA.n2451 3.4105
R15602 GNDA.n2466 GNDA.n1958 3.4105
R15603 GNDA.n2466 GNDA.n2453 3.4105
R15604 GNDA.n2466 GNDA.n1957 3.4105
R15605 GNDA.n2466 GNDA.n2455 3.4105
R15606 GNDA.n2466 GNDA.n1956 3.4105
R15607 GNDA.n2466 GNDA.n2457 3.4105
R15608 GNDA.n2466 GNDA.n1955 3.4105
R15609 GNDA.n2466 GNDA.n2459 3.4105
R15610 GNDA.n2466 GNDA.n1954 3.4105
R15611 GNDA.n2466 GNDA.n2461 3.4105
R15612 GNDA.n2466 GNDA.n1953 3.4105
R15613 GNDA.n2466 GNDA.n2463 3.4105
R15614 GNDA.n2466 GNDA.n1952 3.4105
R15615 GNDA.n2466 GNDA.n2465 3.4105
R15616 GNDA.n2467 GNDA.n2466 3.4105
R15617 GNDA.n2378 GNDA.n2066 3.4105
R15618 GNDA.n2378 GNDA.n2377 3.4105
R15619 GNDA.n2344 GNDA.n2083 3.4105
R15620 GNDA.n2083 GNDA.n2066 3.4105
R15621 GNDA.n2377 GNDA.n2083 3.4105
R15622 GNDA.n2344 GNDA.n2086 3.4105
R15623 GNDA.n2149 GNDA.n2086 3.4105
R15624 GNDA.n2346 GNDA.n2086 3.4105
R15625 GNDA.n2148 GNDA.n2086 3.4105
R15626 GNDA.n2348 GNDA.n2086 3.4105
R15627 GNDA.n2147 GNDA.n2086 3.4105
R15628 GNDA.n2350 GNDA.n2086 3.4105
R15629 GNDA.n2146 GNDA.n2086 3.4105
R15630 GNDA.n2352 GNDA.n2086 3.4105
R15631 GNDA.n2145 GNDA.n2086 3.4105
R15632 GNDA.n2354 GNDA.n2086 3.4105
R15633 GNDA.n2144 GNDA.n2086 3.4105
R15634 GNDA.n2356 GNDA.n2086 3.4105
R15635 GNDA.n2143 GNDA.n2086 3.4105
R15636 GNDA.n2358 GNDA.n2086 3.4105
R15637 GNDA.n2142 GNDA.n2086 3.4105
R15638 GNDA.n2360 GNDA.n2086 3.4105
R15639 GNDA.n2141 GNDA.n2086 3.4105
R15640 GNDA.n2362 GNDA.n2086 3.4105
R15641 GNDA.n2140 GNDA.n2086 3.4105
R15642 GNDA.n2364 GNDA.n2086 3.4105
R15643 GNDA.n2139 GNDA.n2086 3.4105
R15644 GNDA.n2366 GNDA.n2086 3.4105
R15645 GNDA.n2138 GNDA.n2086 3.4105
R15646 GNDA.n2368 GNDA.n2086 3.4105
R15647 GNDA.n2137 GNDA.n2086 3.4105
R15648 GNDA.n2370 GNDA.n2086 3.4105
R15649 GNDA.n2136 GNDA.n2086 3.4105
R15650 GNDA.n2372 GNDA.n2086 3.4105
R15651 GNDA.n2135 GNDA.n2086 3.4105
R15652 GNDA.n2374 GNDA.n2086 3.4105
R15653 GNDA.n2086 GNDA.n2066 3.4105
R15654 GNDA.n2377 GNDA.n2086 3.4105
R15655 GNDA.n2344 GNDA.n2082 3.4105
R15656 GNDA.n2149 GNDA.n2082 3.4105
R15657 GNDA.n2346 GNDA.n2082 3.4105
R15658 GNDA.n2148 GNDA.n2082 3.4105
R15659 GNDA.n2348 GNDA.n2082 3.4105
R15660 GNDA.n2147 GNDA.n2082 3.4105
R15661 GNDA.n2350 GNDA.n2082 3.4105
R15662 GNDA.n2146 GNDA.n2082 3.4105
R15663 GNDA.n2352 GNDA.n2082 3.4105
R15664 GNDA.n2145 GNDA.n2082 3.4105
R15665 GNDA.n2354 GNDA.n2082 3.4105
R15666 GNDA.n2144 GNDA.n2082 3.4105
R15667 GNDA.n2356 GNDA.n2082 3.4105
R15668 GNDA.n2143 GNDA.n2082 3.4105
R15669 GNDA.n2358 GNDA.n2082 3.4105
R15670 GNDA.n2142 GNDA.n2082 3.4105
R15671 GNDA.n2360 GNDA.n2082 3.4105
R15672 GNDA.n2141 GNDA.n2082 3.4105
R15673 GNDA.n2362 GNDA.n2082 3.4105
R15674 GNDA.n2140 GNDA.n2082 3.4105
R15675 GNDA.n2364 GNDA.n2082 3.4105
R15676 GNDA.n2139 GNDA.n2082 3.4105
R15677 GNDA.n2366 GNDA.n2082 3.4105
R15678 GNDA.n2138 GNDA.n2082 3.4105
R15679 GNDA.n2368 GNDA.n2082 3.4105
R15680 GNDA.n2137 GNDA.n2082 3.4105
R15681 GNDA.n2370 GNDA.n2082 3.4105
R15682 GNDA.n2136 GNDA.n2082 3.4105
R15683 GNDA.n2372 GNDA.n2082 3.4105
R15684 GNDA.n2135 GNDA.n2082 3.4105
R15685 GNDA.n2374 GNDA.n2082 3.4105
R15686 GNDA.n2082 GNDA.n2066 3.4105
R15687 GNDA.n2377 GNDA.n2082 3.4105
R15688 GNDA.n2344 GNDA.n2088 3.4105
R15689 GNDA.n2149 GNDA.n2088 3.4105
R15690 GNDA.n2346 GNDA.n2088 3.4105
R15691 GNDA.n2148 GNDA.n2088 3.4105
R15692 GNDA.n2348 GNDA.n2088 3.4105
R15693 GNDA.n2147 GNDA.n2088 3.4105
R15694 GNDA.n2350 GNDA.n2088 3.4105
R15695 GNDA.n2146 GNDA.n2088 3.4105
R15696 GNDA.n2352 GNDA.n2088 3.4105
R15697 GNDA.n2145 GNDA.n2088 3.4105
R15698 GNDA.n2354 GNDA.n2088 3.4105
R15699 GNDA.n2144 GNDA.n2088 3.4105
R15700 GNDA.n2356 GNDA.n2088 3.4105
R15701 GNDA.n2143 GNDA.n2088 3.4105
R15702 GNDA.n2358 GNDA.n2088 3.4105
R15703 GNDA.n2142 GNDA.n2088 3.4105
R15704 GNDA.n2360 GNDA.n2088 3.4105
R15705 GNDA.n2141 GNDA.n2088 3.4105
R15706 GNDA.n2362 GNDA.n2088 3.4105
R15707 GNDA.n2140 GNDA.n2088 3.4105
R15708 GNDA.n2364 GNDA.n2088 3.4105
R15709 GNDA.n2139 GNDA.n2088 3.4105
R15710 GNDA.n2366 GNDA.n2088 3.4105
R15711 GNDA.n2138 GNDA.n2088 3.4105
R15712 GNDA.n2368 GNDA.n2088 3.4105
R15713 GNDA.n2137 GNDA.n2088 3.4105
R15714 GNDA.n2370 GNDA.n2088 3.4105
R15715 GNDA.n2136 GNDA.n2088 3.4105
R15716 GNDA.n2372 GNDA.n2088 3.4105
R15717 GNDA.n2135 GNDA.n2088 3.4105
R15718 GNDA.n2374 GNDA.n2088 3.4105
R15719 GNDA.n2088 GNDA.n2066 3.4105
R15720 GNDA.n2377 GNDA.n2088 3.4105
R15721 GNDA.n2344 GNDA.n2081 3.4105
R15722 GNDA.n2149 GNDA.n2081 3.4105
R15723 GNDA.n2346 GNDA.n2081 3.4105
R15724 GNDA.n2148 GNDA.n2081 3.4105
R15725 GNDA.n2348 GNDA.n2081 3.4105
R15726 GNDA.n2147 GNDA.n2081 3.4105
R15727 GNDA.n2350 GNDA.n2081 3.4105
R15728 GNDA.n2146 GNDA.n2081 3.4105
R15729 GNDA.n2352 GNDA.n2081 3.4105
R15730 GNDA.n2145 GNDA.n2081 3.4105
R15731 GNDA.n2354 GNDA.n2081 3.4105
R15732 GNDA.n2144 GNDA.n2081 3.4105
R15733 GNDA.n2356 GNDA.n2081 3.4105
R15734 GNDA.n2143 GNDA.n2081 3.4105
R15735 GNDA.n2358 GNDA.n2081 3.4105
R15736 GNDA.n2142 GNDA.n2081 3.4105
R15737 GNDA.n2360 GNDA.n2081 3.4105
R15738 GNDA.n2141 GNDA.n2081 3.4105
R15739 GNDA.n2362 GNDA.n2081 3.4105
R15740 GNDA.n2140 GNDA.n2081 3.4105
R15741 GNDA.n2364 GNDA.n2081 3.4105
R15742 GNDA.n2139 GNDA.n2081 3.4105
R15743 GNDA.n2366 GNDA.n2081 3.4105
R15744 GNDA.n2138 GNDA.n2081 3.4105
R15745 GNDA.n2368 GNDA.n2081 3.4105
R15746 GNDA.n2137 GNDA.n2081 3.4105
R15747 GNDA.n2370 GNDA.n2081 3.4105
R15748 GNDA.n2136 GNDA.n2081 3.4105
R15749 GNDA.n2372 GNDA.n2081 3.4105
R15750 GNDA.n2135 GNDA.n2081 3.4105
R15751 GNDA.n2374 GNDA.n2081 3.4105
R15752 GNDA.n2081 GNDA.n2066 3.4105
R15753 GNDA.n2377 GNDA.n2081 3.4105
R15754 GNDA.n2344 GNDA.n2090 3.4105
R15755 GNDA.n2149 GNDA.n2090 3.4105
R15756 GNDA.n2346 GNDA.n2090 3.4105
R15757 GNDA.n2148 GNDA.n2090 3.4105
R15758 GNDA.n2348 GNDA.n2090 3.4105
R15759 GNDA.n2147 GNDA.n2090 3.4105
R15760 GNDA.n2350 GNDA.n2090 3.4105
R15761 GNDA.n2146 GNDA.n2090 3.4105
R15762 GNDA.n2352 GNDA.n2090 3.4105
R15763 GNDA.n2145 GNDA.n2090 3.4105
R15764 GNDA.n2354 GNDA.n2090 3.4105
R15765 GNDA.n2144 GNDA.n2090 3.4105
R15766 GNDA.n2356 GNDA.n2090 3.4105
R15767 GNDA.n2143 GNDA.n2090 3.4105
R15768 GNDA.n2358 GNDA.n2090 3.4105
R15769 GNDA.n2142 GNDA.n2090 3.4105
R15770 GNDA.n2360 GNDA.n2090 3.4105
R15771 GNDA.n2141 GNDA.n2090 3.4105
R15772 GNDA.n2362 GNDA.n2090 3.4105
R15773 GNDA.n2140 GNDA.n2090 3.4105
R15774 GNDA.n2364 GNDA.n2090 3.4105
R15775 GNDA.n2139 GNDA.n2090 3.4105
R15776 GNDA.n2366 GNDA.n2090 3.4105
R15777 GNDA.n2138 GNDA.n2090 3.4105
R15778 GNDA.n2368 GNDA.n2090 3.4105
R15779 GNDA.n2137 GNDA.n2090 3.4105
R15780 GNDA.n2370 GNDA.n2090 3.4105
R15781 GNDA.n2136 GNDA.n2090 3.4105
R15782 GNDA.n2372 GNDA.n2090 3.4105
R15783 GNDA.n2135 GNDA.n2090 3.4105
R15784 GNDA.n2374 GNDA.n2090 3.4105
R15785 GNDA.n2090 GNDA.n2066 3.4105
R15786 GNDA.n2377 GNDA.n2090 3.4105
R15787 GNDA.n2344 GNDA.n2080 3.4105
R15788 GNDA.n2149 GNDA.n2080 3.4105
R15789 GNDA.n2346 GNDA.n2080 3.4105
R15790 GNDA.n2148 GNDA.n2080 3.4105
R15791 GNDA.n2348 GNDA.n2080 3.4105
R15792 GNDA.n2147 GNDA.n2080 3.4105
R15793 GNDA.n2350 GNDA.n2080 3.4105
R15794 GNDA.n2146 GNDA.n2080 3.4105
R15795 GNDA.n2352 GNDA.n2080 3.4105
R15796 GNDA.n2145 GNDA.n2080 3.4105
R15797 GNDA.n2354 GNDA.n2080 3.4105
R15798 GNDA.n2144 GNDA.n2080 3.4105
R15799 GNDA.n2356 GNDA.n2080 3.4105
R15800 GNDA.n2143 GNDA.n2080 3.4105
R15801 GNDA.n2358 GNDA.n2080 3.4105
R15802 GNDA.n2142 GNDA.n2080 3.4105
R15803 GNDA.n2360 GNDA.n2080 3.4105
R15804 GNDA.n2141 GNDA.n2080 3.4105
R15805 GNDA.n2362 GNDA.n2080 3.4105
R15806 GNDA.n2140 GNDA.n2080 3.4105
R15807 GNDA.n2364 GNDA.n2080 3.4105
R15808 GNDA.n2139 GNDA.n2080 3.4105
R15809 GNDA.n2366 GNDA.n2080 3.4105
R15810 GNDA.n2138 GNDA.n2080 3.4105
R15811 GNDA.n2368 GNDA.n2080 3.4105
R15812 GNDA.n2137 GNDA.n2080 3.4105
R15813 GNDA.n2370 GNDA.n2080 3.4105
R15814 GNDA.n2136 GNDA.n2080 3.4105
R15815 GNDA.n2372 GNDA.n2080 3.4105
R15816 GNDA.n2135 GNDA.n2080 3.4105
R15817 GNDA.n2374 GNDA.n2080 3.4105
R15818 GNDA.n2080 GNDA.n2066 3.4105
R15819 GNDA.n2377 GNDA.n2080 3.4105
R15820 GNDA.n2344 GNDA.n2092 3.4105
R15821 GNDA.n2149 GNDA.n2092 3.4105
R15822 GNDA.n2346 GNDA.n2092 3.4105
R15823 GNDA.n2148 GNDA.n2092 3.4105
R15824 GNDA.n2348 GNDA.n2092 3.4105
R15825 GNDA.n2147 GNDA.n2092 3.4105
R15826 GNDA.n2350 GNDA.n2092 3.4105
R15827 GNDA.n2146 GNDA.n2092 3.4105
R15828 GNDA.n2352 GNDA.n2092 3.4105
R15829 GNDA.n2145 GNDA.n2092 3.4105
R15830 GNDA.n2354 GNDA.n2092 3.4105
R15831 GNDA.n2144 GNDA.n2092 3.4105
R15832 GNDA.n2356 GNDA.n2092 3.4105
R15833 GNDA.n2143 GNDA.n2092 3.4105
R15834 GNDA.n2358 GNDA.n2092 3.4105
R15835 GNDA.n2142 GNDA.n2092 3.4105
R15836 GNDA.n2360 GNDA.n2092 3.4105
R15837 GNDA.n2141 GNDA.n2092 3.4105
R15838 GNDA.n2362 GNDA.n2092 3.4105
R15839 GNDA.n2140 GNDA.n2092 3.4105
R15840 GNDA.n2364 GNDA.n2092 3.4105
R15841 GNDA.n2139 GNDA.n2092 3.4105
R15842 GNDA.n2366 GNDA.n2092 3.4105
R15843 GNDA.n2138 GNDA.n2092 3.4105
R15844 GNDA.n2368 GNDA.n2092 3.4105
R15845 GNDA.n2137 GNDA.n2092 3.4105
R15846 GNDA.n2370 GNDA.n2092 3.4105
R15847 GNDA.n2136 GNDA.n2092 3.4105
R15848 GNDA.n2372 GNDA.n2092 3.4105
R15849 GNDA.n2135 GNDA.n2092 3.4105
R15850 GNDA.n2374 GNDA.n2092 3.4105
R15851 GNDA.n2092 GNDA.n2066 3.4105
R15852 GNDA.n2377 GNDA.n2092 3.4105
R15853 GNDA.n2344 GNDA.n2079 3.4105
R15854 GNDA.n2149 GNDA.n2079 3.4105
R15855 GNDA.n2346 GNDA.n2079 3.4105
R15856 GNDA.n2148 GNDA.n2079 3.4105
R15857 GNDA.n2348 GNDA.n2079 3.4105
R15858 GNDA.n2147 GNDA.n2079 3.4105
R15859 GNDA.n2350 GNDA.n2079 3.4105
R15860 GNDA.n2146 GNDA.n2079 3.4105
R15861 GNDA.n2352 GNDA.n2079 3.4105
R15862 GNDA.n2145 GNDA.n2079 3.4105
R15863 GNDA.n2354 GNDA.n2079 3.4105
R15864 GNDA.n2144 GNDA.n2079 3.4105
R15865 GNDA.n2356 GNDA.n2079 3.4105
R15866 GNDA.n2143 GNDA.n2079 3.4105
R15867 GNDA.n2358 GNDA.n2079 3.4105
R15868 GNDA.n2142 GNDA.n2079 3.4105
R15869 GNDA.n2360 GNDA.n2079 3.4105
R15870 GNDA.n2141 GNDA.n2079 3.4105
R15871 GNDA.n2362 GNDA.n2079 3.4105
R15872 GNDA.n2140 GNDA.n2079 3.4105
R15873 GNDA.n2364 GNDA.n2079 3.4105
R15874 GNDA.n2139 GNDA.n2079 3.4105
R15875 GNDA.n2366 GNDA.n2079 3.4105
R15876 GNDA.n2138 GNDA.n2079 3.4105
R15877 GNDA.n2368 GNDA.n2079 3.4105
R15878 GNDA.n2137 GNDA.n2079 3.4105
R15879 GNDA.n2370 GNDA.n2079 3.4105
R15880 GNDA.n2136 GNDA.n2079 3.4105
R15881 GNDA.n2372 GNDA.n2079 3.4105
R15882 GNDA.n2135 GNDA.n2079 3.4105
R15883 GNDA.n2374 GNDA.n2079 3.4105
R15884 GNDA.n2079 GNDA.n2066 3.4105
R15885 GNDA.n2377 GNDA.n2079 3.4105
R15886 GNDA.n2344 GNDA.n2094 3.4105
R15887 GNDA.n2149 GNDA.n2094 3.4105
R15888 GNDA.n2346 GNDA.n2094 3.4105
R15889 GNDA.n2148 GNDA.n2094 3.4105
R15890 GNDA.n2348 GNDA.n2094 3.4105
R15891 GNDA.n2147 GNDA.n2094 3.4105
R15892 GNDA.n2350 GNDA.n2094 3.4105
R15893 GNDA.n2146 GNDA.n2094 3.4105
R15894 GNDA.n2352 GNDA.n2094 3.4105
R15895 GNDA.n2145 GNDA.n2094 3.4105
R15896 GNDA.n2354 GNDA.n2094 3.4105
R15897 GNDA.n2144 GNDA.n2094 3.4105
R15898 GNDA.n2356 GNDA.n2094 3.4105
R15899 GNDA.n2143 GNDA.n2094 3.4105
R15900 GNDA.n2358 GNDA.n2094 3.4105
R15901 GNDA.n2142 GNDA.n2094 3.4105
R15902 GNDA.n2360 GNDA.n2094 3.4105
R15903 GNDA.n2141 GNDA.n2094 3.4105
R15904 GNDA.n2362 GNDA.n2094 3.4105
R15905 GNDA.n2140 GNDA.n2094 3.4105
R15906 GNDA.n2364 GNDA.n2094 3.4105
R15907 GNDA.n2139 GNDA.n2094 3.4105
R15908 GNDA.n2366 GNDA.n2094 3.4105
R15909 GNDA.n2138 GNDA.n2094 3.4105
R15910 GNDA.n2368 GNDA.n2094 3.4105
R15911 GNDA.n2137 GNDA.n2094 3.4105
R15912 GNDA.n2370 GNDA.n2094 3.4105
R15913 GNDA.n2136 GNDA.n2094 3.4105
R15914 GNDA.n2372 GNDA.n2094 3.4105
R15915 GNDA.n2135 GNDA.n2094 3.4105
R15916 GNDA.n2374 GNDA.n2094 3.4105
R15917 GNDA.n2094 GNDA.n2066 3.4105
R15918 GNDA.n2377 GNDA.n2094 3.4105
R15919 GNDA.n2344 GNDA.n2078 3.4105
R15920 GNDA.n2149 GNDA.n2078 3.4105
R15921 GNDA.n2346 GNDA.n2078 3.4105
R15922 GNDA.n2148 GNDA.n2078 3.4105
R15923 GNDA.n2348 GNDA.n2078 3.4105
R15924 GNDA.n2147 GNDA.n2078 3.4105
R15925 GNDA.n2350 GNDA.n2078 3.4105
R15926 GNDA.n2146 GNDA.n2078 3.4105
R15927 GNDA.n2352 GNDA.n2078 3.4105
R15928 GNDA.n2145 GNDA.n2078 3.4105
R15929 GNDA.n2354 GNDA.n2078 3.4105
R15930 GNDA.n2144 GNDA.n2078 3.4105
R15931 GNDA.n2356 GNDA.n2078 3.4105
R15932 GNDA.n2143 GNDA.n2078 3.4105
R15933 GNDA.n2358 GNDA.n2078 3.4105
R15934 GNDA.n2142 GNDA.n2078 3.4105
R15935 GNDA.n2360 GNDA.n2078 3.4105
R15936 GNDA.n2141 GNDA.n2078 3.4105
R15937 GNDA.n2362 GNDA.n2078 3.4105
R15938 GNDA.n2140 GNDA.n2078 3.4105
R15939 GNDA.n2364 GNDA.n2078 3.4105
R15940 GNDA.n2139 GNDA.n2078 3.4105
R15941 GNDA.n2366 GNDA.n2078 3.4105
R15942 GNDA.n2138 GNDA.n2078 3.4105
R15943 GNDA.n2368 GNDA.n2078 3.4105
R15944 GNDA.n2137 GNDA.n2078 3.4105
R15945 GNDA.n2370 GNDA.n2078 3.4105
R15946 GNDA.n2136 GNDA.n2078 3.4105
R15947 GNDA.n2372 GNDA.n2078 3.4105
R15948 GNDA.n2135 GNDA.n2078 3.4105
R15949 GNDA.n2374 GNDA.n2078 3.4105
R15950 GNDA.n2078 GNDA.n2066 3.4105
R15951 GNDA.n2377 GNDA.n2078 3.4105
R15952 GNDA.n2344 GNDA.n2096 3.4105
R15953 GNDA.n2149 GNDA.n2096 3.4105
R15954 GNDA.n2346 GNDA.n2096 3.4105
R15955 GNDA.n2148 GNDA.n2096 3.4105
R15956 GNDA.n2348 GNDA.n2096 3.4105
R15957 GNDA.n2147 GNDA.n2096 3.4105
R15958 GNDA.n2350 GNDA.n2096 3.4105
R15959 GNDA.n2146 GNDA.n2096 3.4105
R15960 GNDA.n2352 GNDA.n2096 3.4105
R15961 GNDA.n2145 GNDA.n2096 3.4105
R15962 GNDA.n2354 GNDA.n2096 3.4105
R15963 GNDA.n2144 GNDA.n2096 3.4105
R15964 GNDA.n2356 GNDA.n2096 3.4105
R15965 GNDA.n2143 GNDA.n2096 3.4105
R15966 GNDA.n2358 GNDA.n2096 3.4105
R15967 GNDA.n2142 GNDA.n2096 3.4105
R15968 GNDA.n2360 GNDA.n2096 3.4105
R15969 GNDA.n2141 GNDA.n2096 3.4105
R15970 GNDA.n2362 GNDA.n2096 3.4105
R15971 GNDA.n2140 GNDA.n2096 3.4105
R15972 GNDA.n2364 GNDA.n2096 3.4105
R15973 GNDA.n2139 GNDA.n2096 3.4105
R15974 GNDA.n2366 GNDA.n2096 3.4105
R15975 GNDA.n2138 GNDA.n2096 3.4105
R15976 GNDA.n2368 GNDA.n2096 3.4105
R15977 GNDA.n2137 GNDA.n2096 3.4105
R15978 GNDA.n2370 GNDA.n2096 3.4105
R15979 GNDA.n2136 GNDA.n2096 3.4105
R15980 GNDA.n2372 GNDA.n2096 3.4105
R15981 GNDA.n2135 GNDA.n2096 3.4105
R15982 GNDA.n2374 GNDA.n2096 3.4105
R15983 GNDA.n2096 GNDA.n2066 3.4105
R15984 GNDA.n2377 GNDA.n2096 3.4105
R15985 GNDA.n2344 GNDA.n2077 3.4105
R15986 GNDA.n2149 GNDA.n2077 3.4105
R15987 GNDA.n2346 GNDA.n2077 3.4105
R15988 GNDA.n2148 GNDA.n2077 3.4105
R15989 GNDA.n2348 GNDA.n2077 3.4105
R15990 GNDA.n2147 GNDA.n2077 3.4105
R15991 GNDA.n2350 GNDA.n2077 3.4105
R15992 GNDA.n2146 GNDA.n2077 3.4105
R15993 GNDA.n2352 GNDA.n2077 3.4105
R15994 GNDA.n2145 GNDA.n2077 3.4105
R15995 GNDA.n2354 GNDA.n2077 3.4105
R15996 GNDA.n2144 GNDA.n2077 3.4105
R15997 GNDA.n2356 GNDA.n2077 3.4105
R15998 GNDA.n2143 GNDA.n2077 3.4105
R15999 GNDA.n2358 GNDA.n2077 3.4105
R16000 GNDA.n2142 GNDA.n2077 3.4105
R16001 GNDA.n2360 GNDA.n2077 3.4105
R16002 GNDA.n2141 GNDA.n2077 3.4105
R16003 GNDA.n2362 GNDA.n2077 3.4105
R16004 GNDA.n2140 GNDA.n2077 3.4105
R16005 GNDA.n2364 GNDA.n2077 3.4105
R16006 GNDA.n2139 GNDA.n2077 3.4105
R16007 GNDA.n2366 GNDA.n2077 3.4105
R16008 GNDA.n2138 GNDA.n2077 3.4105
R16009 GNDA.n2368 GNDA.n2077 3.4105
R16010 GNDA.n2137 GNDA.n2077 3.4105
R16011 GNDA.n2370 GNDA.n2077 3.4105
R16012 GNDA.n2136 GNDA.n2077 3.4105
R16013 GNDA.n2372 GNDA.n2077 3.4105
R16014 GNDA.n2135 GNDA.n2077 3.4105
R16015 GNDA.n2374 GNDA.n2077 3.4105
R16016 GNDA.n2077 GNDA.n2066 3.4105
R16017 GNDA.n2377 GNDA.n2077 3.4105
R16018 GNDA.n2344 GNDA.n2098 3.4105
R16019 GNDA.n2149 GNDA.n2098 3.4105
R16020 GNDA.n2346 GNDA.n2098 3.4105
R16021 GNDA.n2148 GNDA.n2098 3.4105
R16022 GNDA.n2348 GNDA.n2098 3.4105
R16023 GNDA.n2147 GNDA.n2098 3.4105
R16024 GNDA.n2350 GNDA.n2098 3.4105
R16025 GNDA.n2146 GNDA.n2098 3.4105
R16026 GNDA.n2352 GNDA.n2098 3.4105
R16027 GNDA.n2145 GNDA.n2098 3.4105
R16028 GNDA.n2354 GNDA.n2098 3.4105
R16029 GNDA.n2144 GNDA.n2098 3.4105
R16030 GNDA.n2356 GNDA.n2098 3.4105
R16031 GNDA.n2143 GNDA.n2098 3.4105
R16032 GNDA.n2358 GNDA.n2098 3.4105
R16033 GNDA.n2142 GNDA.n2098 3.4105
R16034 GNDA.n2360 GNDA.n2098 3.4105
R16035 GNDA.n2141 GNDA.n2098 3.4105
R16036 GNDA.n2362 GNDA.n2098 3.4105
R16037 GNDA.n2140 GNDA.n2098 3.4105
R16038 GNDA.n2364 GNDA.n2098 3.4105
R16039 GNDA.n2139 GNDA.n2098 3.4105
R16040 GNDA.n2366 GNDA.n2098 3.4105
R16041 GNDA.n2138 GNDA.n2098 3.4105
R16042 GNDA.n2368 GNDA.n2098 3.4105
R16043 GNDA.n2137 GNDA.n2098 3.4105
R16044 GNDA.n2370 GNDA.n2098 3.4105
R16045 GNDA.n2136 GNDA.n2098 3.4105
R16046 GNDA.n2372 GNDA.n2098 3.4105
R16047 GNDA.n2135 GNDA.n2098 3.4105
R16048 GNDA.n2374 GNDA.n2098 3.4105
R16049 GNDA.n2098 GNDA.n2066 3.4105
R16050 GNDA.n2377 GNDA.n2098 3.4105
R16051 GNDA.n2344 GNDA.n2076 3.4105
R16052 GNDA.n2149 GNDA.n2076 3.4105
R16053 GNDA.n2346 GNDA.n2076 3.4105
R16054 GNDA.n2148 GNDA.n2076 3.4105
R16055 GNDA.n2348 GNDA.n2076 3.4105
R16056 GNDA.n2147 GNDA.n2076 3.4105
R16057 GNDA.n2350 GNDA.n2076 3.4105
R16058 GNDA.n2146 GNDA.n2076 3.4105
R16059 GNDA.n2352 GNDA.n2076 3.4105
R16060 GNDA.n2145 GNDA.n2076 3.4105
R16061 GNDA.n2354 GNDA.n2076 3.4105
R16062 GNDA.n2144 GNDA.n2076 3.4105
R16063 GNDA.n2356 GNDA.n2076 3.4105
R16064 GNDA.n2143 GNDA.n2076 3.4105
R16065 GNDA.n2358 GNDA.n2076 3.4105
R16066 GNDA.n2142 GNDA.n2076 3.4105
R16067 GNDA.n2360 GNDA.n2076 3.4105
R16068 GNDA.n2141 GNDA.n2076 3.4105
R16069 GNDA.n2362 GNDA.n2076 3.4105
R16070 GNDA.n2140 GNDA.n2076 3.4105
R16071 GNDA.n2364 GNDA.n2076 3.4105
R16072 GNDA.n2139 GNDA.n2076 3.4105
R16073 GNDA.n2366 GNDA.n2076 3.4105
R16074 GNDA.n2138 GNDA.n2076 3.4105
R16075 GNDA.n2368 GNDA.n2076 3.4105
R16076 GNDA.n2137 GNDA.n2076 3.4105
R16077 GNDA.n2370 GNDA.n2076 3.4105
R16078 GNDA.n2136 GNDA.n2076 3.4105
R16079 GNDA.n2372 GNDA.n2076 3.4105
R16080 GNDA.n2135 GNDA.n2076 3.4105
R16081 GNDA.n2374 GNDA.n2076 3.4105
R16082 GNDA.n2076 GNDA.n2066 3.4105
R16083 GNDA.n2377 GNDA.n2076 3.4105
R16084 GNDA.n2344 GNDA.n2100 3.4105
R16085 GNDA.n2149 GNDA.n2100 3.4105
R16086 GNDA.n2346 GNDA.n2100 3.4105
R16087 GNDA.n2148 GNDA.n2100 3.4105
R16088 GNDA.n2348 GNDA.n2100 3.4105
R16089 GNDA.n2147 GNDA.n2100 3.4105
R16090 GNDA.n2350 GNDA.n2100 3.4105
R16091 GNDA.n2146 GNDA.n2100 3.4105
R16092 GNDA.n2352 GNDA.n2100 3.4105
R16093 GNDA.n2145 GNDA.n2100 3.4105
R16094 GNDA.n2354 GNDA.n2100 3.4105
R16095 GNDA.n2144 GNDA.n2100 3.4105
R16096 GNDA.n2356 GNDA.n2100 3.4105
R16097 GNDA.n2143 GNDA.n2100 3.4105
R16098 GNDA.n2358 GNDA.n2100 3.4105
R16099 GNDA.n2142 GNDA.n2100 3.4105
R16100 GNDA.n2360 GNDA.n2100 3.4105
R16101 GNDA.n2141 GNDA.n2100 3.4105
R16102 GNDA.n2362 GNDA.n2100 3.4105
R16103 GNDA.n2140 GNDA.n2100 3.4105
R16104 GNDA.n2364 GNDA.n2100 3.4105
R16105 GNDA.n2139 GNDA.n2100 3.4105
R16106 GNDA.n2366 GNDA.n2100 3.4105
R16107 GNDA.n2138 GNDA.n2100 3.4105
R16108 GNDA.n2368 GNDA.n2100 3.4105
R16109 GNDA.n2137 GNDA.n2100 3.4105
R16110 GNDA.n2370 GNDA.n2100 3.4105
R16111 GNDA.n2136 GNDA.n2100 3.4105
R16112 GNDA.n2372 GNDA.n2100 3.4105
R16113 GNDA.n2135 GNDA.n2100 3.4105
R16114 GNDA.n2374 GNDA.n2100 3.4105
R16115 GNDA.n2100 GNDA.n2066 3.4105
R16116 GNDA.n2377 GNDA.n2100 3.4105
R16117 GNDA.n2344 GNDA.n2075 3.4105
R16118 GNDA.n2149 GNDA.n2075 3.4105
R16119 GNDA.n2346 GNDA.n2075 3.4105
R16120 GNDA.n2148 GNDA.n2075 3.4105
R16121 GNDA.n2348 GNDA.n2075 3.4105
R16122 GNDA.n2147 GNDA.n2075 3.4105
R16123 GNDA.n2350 GNDA.n2075 3.4105
R16124 GNDA.n2146 GNDA.n2075 3.4105
R16125 GNDA.n2352 GNDA.n2075 3.4105
R16126 GNDA.n2145 GNDA.n2075 3.4105
R16127 GNDA.n2354 GNDA.n2075 3.4105
R16128 GNDA.n2144 GNDA.n2075 3.4105
R16129 GNDA.n2356 GNDA.n2075 3.4105
R16130 GNDA.n2143 GNDA.n2075 3.4105
R16131 GNDA.n2358 GNDA.n2075 3.4105
R16132 GNDA.n2142 GNDA.n2075 3.4105
R16133 GNDA.n2360 GNDA.n2075 3.4105
R16134 GNDA.n2141 GNDA.n2075 3.4105
R16135 GNDA.n2362 GNDA.n2075 3.4105
R16136 GNDA.n2140 GNDA.n2075 3.4105
R16137 GNDA.n2364 GNDA.n2075 3.4105
R16138 GNDA.n2139 GNDA.n2075 3.4105
R16139 GNDA.n2366 GNDA.n2075 3.4105
R16140 GNDA.n2138 GNDA.n2075 3.4105
R16141 GNDA.n2368 GNDA.n2075 3.4105
R16142 GNDA.n2137 GNDA.n2075 3.4105
R16143 GNDA.n2370 GNDA.n2075 3.4105
R16144 GNDA.n2136 GNDA.n2075 3.4105
R16145 GNDA.n2372 GNDA.n2075 3.4105
R16146 GNDA.n2135 GNDA.n2075 3.4105
R16147 GNDA.n2374 GNDA.n2075 3.4105
R16148 GNDA.n2075 GNDA.n2066 3.4105
R16149 GNDA.n2377 GNDA.n2075 3.4105
R16150 GNDA.n2344 GNDA.n2102 3.4105
R16151 GNDA.n2149 GNDA.n2102 3.4105
R16152 GNDA.n2346 GNDA.n2102 3.4105
R16153 GNDA.n2148 GNDA.n2102 3.4105
R16154 GNDA.n2348 GNDA.n2102 3.4105
R16155 GNDA.n2147 GNDA.n2102 3.4105
R16156 GNDA.n2350 GNDA.n2102 3.4105
R16157 GNDA.n2146 GNDA.n2102 3.4105
R16158 GNDA.n2352 GNDA.n2102 3.4105
R16159 GNDA.n2145 GNDA.n2102 3.4105
R16160 GNDA.n2354 GNDA.n2102 3.4105
R16161 GNDA.n2144 GNDA.n2102 3.4105
R16162 GNDA.n2356 GNDA.n2102 3.4105
R16163 GNDA.n2143 GNDA.n2102 3.4105
R16164 GNDA.n2358 GNDA.n2102 3.4105
R16165 GNDA.n2142 GNDA.n2102 3.4105
R16166 GNDA.n2360 GNDA.n2102 3.4105
R16167 GNDA.n2141 GNDA.n2102 3.4105
R16168 GNDA.n2362 GNDA.n2102 3.4105
R16169 GNDA.n2140 GNDA.n2102 3.4105
R16170 GNDA.n2364 GNDA.n2102 3.4105
R16171 GNDA.n2139 GNDA.n2102 3.4105
R16172 GNDA.n2366 GNDA.n2102 3.4105
R16173 GNDA.n2138 GNDA.n2102 3.4105
R16174 GNDA.n2368 GNDA.n2102 3.4105
R16175 GNDA.n2137 GNDA.n2102 3.4105
R16176 GNDA.n2370 GNDA.n2102 3.4105
R16177 GNDA.n2136 GNDA.n2102 3.4105
R16178 GNDA.n2372 GNDA.n2102 3.4105
R16179 GNDA.n2135 GNDA.n2102 3.4105
R16180 GNDA.n2374 GNDA.n2102 3.4105
R16181 GNDA.n2102 GNDA.n2066 3.4105
R16182 GNDA.n2377 GNDA.n2102 3.4105
R16183 GNDA.n2344 GNDA.n2074 3.4105
R16184 GNDA.n2149 GNDA.n2074 3.4105
R16185 GNDA.n2346 GNDA.n2074 3.4105
R16186 GNDA.n2148 GNDA.n2074 3.4105
R16187 GNDA.n2348 GNDA.n2074 3.4105
R16188 GNDA.n2147 GNDA.n2074 3.4105
R16189 GNDA.n2350 GNDA.n2074 3.4105
R16190 GNDA.n2146 GNDA.n2074 3.4105
R16191 GNDA.n2352 GNDA.n2074 3.4105
R16192 GNDA.n2145 GNDA.n2074 3.4105
R16193 GNDA.n2354 GNDA.n2074 3.4105
R16194 GNDA.n2144 GNDA.n2074 3.4105
R16195 GNDA.n2356 GNDA.n2074 3.4105
R16196 GNDA.n2143 GNDA.n2074 3.4105
R16197 GNDA.n2358 GNDA.n2074 3.4105
R16198 GNDA.n2142 GNDA.n2074 3.4105
R16199 GNDA.n2360 GNDA.n2074 3.4105
R16200 GNDA.n2141 GNDA.n2074 3.4105
R16201 GNDA.n2362 GNDA.n2074 3.4105
R16202 GNDA.n2140 GNDA.n2074 3.4105
R16203 GNDA.n2364 GNDA.n2074 3.4105
R16204 GNDA.n2139 GNDA.n2074 3.4105
R16205 GNDA.n2366 GNDA.n2074 3.4105
R16206 GNDA.n2138 GNDA.n2074 3.4105
R16207 GNDA.n2368 GNDA.n2074 3.4105
R16208 GNDA.n2137 GNDA.n2074 3.4105
R16209 GNDA.n2370 GNDA.n2074 3.4105
R16210 GNDA.n2136 GNDA.n2074 3.4105
R16211 GNDA.n2372 GNDA.n2074 3.4105
R16212 GNDA.n2135 GNDA.n2074 3.4105
R16213 GNDA.n2374 GNDA.n2074 3.4105
R16214 GNDA.n2074 GNDA.n2066 3.4105
R16215 GNDA.n2377 GNDA.n2074 3.4105
R16216 GNDA.n2344 GNDA.n2104 3.4105
R16217 GNDA.n2149 GNDA.n2104 3.4105
R16218 GNDA.n2346 GNDA.n2104 3.4105
R16219 GNDA.n2148 GNDA.n2104 3.4105
R16220 GNDA.n2348 GNDA.n2104 3.4105
R16221 GNDA.n2147 GNDA.n2104 3.4105
R16222 GNDA.n2350 GNDA.n2104 3.4105
R16223 GNDA.n2146 GNDA.n2104 3.4105
R16224 GNDA.n2352 GNDA.n2104 3.4105
R16225 GNDA.n2145 GNDA.n2104 3.4105
R16226 GNDA.n2354 GNDA.n2104 3.4105
R16227 GNDA.n2144 GNDA.n2104 3.4105
R16228 GNDA.n2356 GNDA.n2104 3.4105
R16229 GNDA.n2143 GNDA.n2104 3.4105
R16230 GNDA.n2358 GNDA.n2104 3.4105
R16231 GNDA.n2142 GNDA.n2104 3.4105
R16232 GNDA.n2360 GNDA.n2104 3.4105
R16233 GNDA.n2141 GNDA.n2104 3.4105
R16234 GNDA.n2362 GNDA.n2104 3.4105
R16235 GNDA.n2140 GNDA.n2104 3.4105
R16236 GNDA.n2364 GNDA.n2104 3.4105
R16237 GNDA.n2139 GNDA.n2104 3.4105
R16238 GNDA.n2366 GNDA.n2104 3.4105
R16239 GNDA.n2138 GNDA.n2104 3.4105
R16240 GNDA.n2368 GNDA.n2104 3.4105
R16241 GNDA.n2137 GNDA.n2104 3.4105
R16242 GNDA.n2370 GNDA.n2104 3.4105
R16243 GNDA.n2136 GNDA.n2104 3.4105
R16244 GNDA.n2372 GNDA.n2104 3.4105
R16245 GNDA.n2135 GNDA.n2104 3.4105
R16246 GNDA.n2374 GNDA.n2104 3.4105
R16247 GNDA.n2104 GNDA.n2066 3.4105
R16248 GNDA.n2377 GNDA.n2104 3.4105
R16249 GNDA.n2344 GNDA.n2073 3.4105
R16250 GNDA.n2149 GNDA.n2073 3.4105
R16251 GNDA.n2346 GNDA.n2073 3.4105
R16252 GNDA.n2148 GNDA.n2073 3.4105
R16253 GNDA.n2348 GNDA.n2073 3.4105
R16254 GNDA.n2147 GNDA.n2073 3.4105
R16255 GNDA.n2350 GNDA.n2073 3.4105
R16256 GNDA.n2146 GNDA.n2073 3.4105
R16257 GNDA.n2352 GNDA.n2073 3.4105
R16258 GNDA.n2145 GNDA.n2073 3.4105
R16259 GNDA.n2354 GNDA.n2073 3.4105
R16260 GNDA.n2144 GNDA.n2073 3.4105
R16261 GNDA.n2356 GNDA.n2073 3.4105
R16262 GNDA.n2143 GNDA.n2073 3.4105
R16263 GNDA.n2358 GNDA.n2073 3.4105
R16264 GNDA.n2142 GNDA.n2073 3.4105
R16265 GNDA.n2360 GNDA.n2073 3.4105
R16266 GNDA.n2141 GNDA.n2073 3.4105
R16267 GNDA.n2362 GNDA.n2073 3.4105
R16268 GNDA.n2140 GNDA.n2073 3.4105
R16269 GNDA.n2364 GNDA.n2073 3.4105
R16270 GNDA.n2139 GNDA.n2073 3.4105
R16271 GNDA.n2366 GNDA.n2073 3.4105
R16272 GNDA.n2138 GNDA.n2073 3.4105
R16273 GNDA.n2368 GNDA.n2073 3.4105
R16274 GNDA.n2137 GNDA.n2073 3.4105
R16275 GNDA.n2370 GNDA.n2073 3.4105
R16276 GNDA.n2136 GNDA.n2073 3.4105
R16277 GNDA.n2372 GNDA.n2073 3.4105
R16278 GNDA.n2135 GNDA.n2073 3.4105
R16279 GNDA.n2374 GNDA.n2073 3.4105
R16280 GNDA.n2073 GNDA.n2066 3.4105
R16281 GNDA.n2377 GNDA.n2073 3.4105
R16282 GNDA.n2344 GNDA.n2106 3.4105
R16283 GNDA.n2149 GNDA.n2106 3.4105
R16284 GNDA.n2346 GNDA.n2106 3.4105
R16285 GNDA.n2148 GNDA.n2106 3.4105
R16286 GNDA.n2348 GNDA.n2106 3.4105
R16287 GNDA.n2147 GNDA.n2106 3.4105
R16288 GNDA.n2350 GNDA.n2106 3.4105
R16289 GNDA.n2146 GNDA.n2106 3.4105
R16290 GNDA.n2352 GNDA.n2106 3.4105
R16291 GNDA.n2145 GNDA.n2106 3.4105
R16292 GNDA.n2354 GNDA.n2106 3.4105
R16293 GNDA.n2144 GNDA.n2106 3.4105
R16294 GNDA.n2356 GNDA.n2106 3.4105
R16295 GNDA.n2143 GNDA.n2106 3.4105
R16296 GNDA.n2358 GNDA.n2106 3.4105
R16297 GNDA.n2142 GNDA.n2106 3.4105
R16298 GNDA.n2360 GNDA.n2106 3.4105
R16299 GNDA.n2141 GNDA.n2106 3.4105
R16300 GNDA.n2362 GNDA.n2106 3.4105
R16301 GNDA.n2140 GNDA.n2106 3.4105
R16302 GNDA.n2364 GNDA.n2106 3.4105
R16303 GNDA.n2139 GNDA.n2106 3.4105
R16304 GNDA.n2366 GNDA.n2106 3.4105
R16305 GNDA.n2138 GNDA.n2106 3.4105
R16306 GNDA.n2368 GNDA.n2106 3.4105
R16307 GNDA.n2137 GNDA.n2106 3.4105
R16308 GNDA.n2370 GNDA.n2106 3.4105
R16309 GNDA.n2136 GNDA.n2106 3.4105
R16310 GNDA.n2372 GNDA.n2106 3.4105
R16311 GNDA.n2135 GNDA.n2106 3.4105
R16312 GNDA.n2374 GNDA.n2106 3.4105
R16313 GNDA.n2106 GNDA.n2066 3.4105
R16314 GNDA.n2377 GNDA.n2106 3.4105
R16315 GNDA.n2344 GNDA.n2072 3.4105
R16316 GNDA.n2149 GNDA.n2072 3.4105
R16317 GNDA.n2346 GNDA.n2072 3.4105
R16318 GNDA.n2148 GNDA.n2072 3.4105
R16319 GNDA.n2348 GNDA.n2072 3.4105
R16320 GNDA.n2147 GNDA.n2072 3.4105
R16321 GNDA.n2350 GNDA.n2072 3.4105
R16322 GNDA.n2146 GNDA.n2072 3.4105
R16323 GNDA.n2352 GNDA.n2072 3.4105
R16324 GNDA.n2145 GNDA.n2072 3.4105
R16325 GNDA.n2354 GNDA.n2072 3.4105
R16326 GNDA.n2144 GNDA.n2072 3.4105
R16327 GNDA.n2356 GNDA.n2072 3.4105
R16328 GNDA.n2143 GNDA.n2072 3.4105
R16329 GNDA.n2358 GNDA.n2072 3.4105
R16330 GNDA.n2142 GNDA.n2072 3.4105
R16331 GNDA.n2360 GNDA.n2072 3.4105
R16332 GNDA.n2141 GNDA.n2072 3.4105
R16333 GNDA.n2362 GNDA.n2072 3.4105
R16334 GNDA.n2140 GNDA.n2072 3.4105
R16335 GNDA.n2364 GNDA.n2072 3.4105
R16336 GNDA.n2139 GNDA.n2072 3.4105
R16337 GNDA.n2366 GNDA.n2072 3.4105
R16338 GNDA.n2138 GNDA.n2072 3.4105
R16339 GNDA.n2368 GNDA.n2072 3.4105
R16340 GNDA.n2137 GNDA.n2072 3.4105
R16341 GNDA.n2370 GNDA.n2072 3.4105
R16342 GNDA.n2136 GNDA.n2072 3.4105
R16343 GNDA.n2372 GNDA.n2072 3.4105
R16344 GNDA.n2135 GNDA.n2072 3.4105
R16345 GNDA.n2374 GNDA.n2072 3.4105
R16346 GNDA.n2072 GNDA.n2066 3.4105
R16347 GNDA.n2377 GNDA.n2072 3.4105
R16348 GNDA.n2344 GNDA.n2108 3.4105
R16349 GNDA.n2149 GNDA.n2108 3.4105
R16350 GNDA.n2346 GNDA.n2108 3.4105
R16351 GNDA.n2148 GNDA.n2108 3.4105
R16352 GNDA.n2348 GNDA.n2108 3.4105
R16353 GNDA.n2147 GNDA.n2108 3.4105
R16354 GNDA.n2350 GNDA.n2108 3.4105
R16355 GNDA.n2146 GNDA.n2108 3.4105
R16356 GNDA.n2352 GNDA.n2108 3.4105
R16357 GNDA.n2145 GNDA.n2108 3.4105
R16358 GNDA.n2354 GNDA.n2108 3.4105
R16359 GNDA.n2144 GNDA.n2108 3.4105
R16360 GNDA.n2356 GNDA.n2108 3.4105
R16361 GNDA.n2143 GNDA.n2108 3.4105
R16362 GNDA.n2358 GNDA.n2108 3.4105
R16363 GNDA.n2142 GNDA.n2108 3.4105
R16364 GNDA.n2360 GNDA.n2108 3.4105
R16365 GNDA.n2141 GNDA.n2108 3.4105
R16366 GNDA.n2362 GNDA.n2108 3.4105
R16367 GNDA.n2140 GNDA.n2108 3.4105
R16368 GNDA.n2364 GNDA.n2108 3.4105
R16369 GNDA.n2139 GNDA.n2108 3.4105
R16370 GNDA.n2366 GNDA.n2108 3.4105
R16371 GNDA.n2138 GNDA.n2108 3.4105
R16372 GNDA.n2368 GNDA.n2108 3.4105
R16373 GNDA.n2137 GNDA.n2108 3.4105
R16374 GNDA.n2370 GNDA.n2108 3.4105
R16375 GNDA.n2136 GNDA.n2108 3.4105
R16376 GNDA.n2372 GNDA.n2108 3.4105
R16377 GNDA.n2135 GNDA.n2108 3.4105
R16378 GNDA.n2374 GNDA.n2108 3.4105
R16379 GNDA.n2108 GNDA.n2066 3.4105
R16380 GNDA.n2377 GNDA.n2108 3.4105
R16381 GNDA.n2344 GNDA.n2071 3.4105
R16382 GNDA.n2149 GNDA.n2071 3.4105
R16383 GNDA.n2346 GNDA.n2071 3.4105
R16384 GNDA.n2148 GNDA.n2071 3.4105
R16385 GNDA.n2348 GNDA.n2071 3.4105
R16386 GNDA.n2147 GNDA.n2071 3.4105
R16387 GNDA.n2350 GNDA.n2071 3.4105
R16388 GNDA.n2146 GNDA.n2071 3.4105
R16389 GNDA.n2352 GNDA.n2071 3.4105
R16390 GNDA.n2145 GNDA.n2071 3.4105
R16391 GNDA.n2354 GNDA.n2071 3.4105
R16392 GNDA.n2144 GNDA.n2071 3.4105
R16393 GNDA.n2356 GNDA.n2071 3.4105
R16394 GNDA.n2143 GNDA.n2071 3.4105
R16395 GNDA.n2358 GNDA.n2071 3.4105
R16396 GNDA.n2142 GNDA.n2071 3.4105
R16397 GNDA.n2360 GNDA.n2071 3.4105
R16398 GNDA.n2141 GNDA.n2071 3.4105
R16399 GNDA.n2362 GNDA.n2071 3.4105
R16400 GNDA.n2140 GNDA.n2071 3.4105
R16401 GNDA.n2364 GNDA.n2071 3.4105
R16402 GNDA.n2139 GNDA.n2071 3.4105
R16403 GNDA.n2366 GNDA.n2071 3.4105
R16404 GNDA.n2138 GNDA.n2071 3.4105
R16405 GNDA.n2368 GNDA.n2071 3.4105
R16406 GNDA.n2137 GNDA.n2071 3.4105
R16407 GNDA.n2370 GNDA.n2071 3.4105
R16408 GNDA.n2136 GNDA.n2071 3.4105
R16409 GNDA.n2372 GNDA.n2071 3.4105
R16410 GNDA.n2135 GNDA.n2071 3.4105
R16411 GNDA.n2374 GNDA.n2071 3.4105
R16412 GNDA.n2071 GNDA.n2066 3.4105
R16413 GNDA.n2377 GNDA.n2071 3.4105
R16414 GNDA.n2344 GNDA.n2110 3.4105
R16415 GNDA.n2149 GNDA.n2110 3.4105
R16416 GNDA.n2346 GNDA.n2110 3.4105
R16417 GNDA.n2148 GNDA.n2110 3.4105
R16418 GNDA.n2348 GNDA.n2110 3.4105
R16419 GNDA.n2147 GNDA.n2110 3.4105
R16420 GNDA.n2350 GNDA.n2110 3.4105
R16421 GNDA.n2146 GNDA.n2110 3.4105
R16422 GNDA.n2352 GNDA.n2110 3.4105
R16423 GNDA.n2145 GNDA.n2110 3.4105
R16424 GNDA.n2354 GNDA.n2110 3.4105
R16425 GNDA.n2144 GNDA.n2110 3.4105
R16426 GNDA.n2356 GNDA.n2110 3.4105
R16427 GNDA.n2143 GNDA.n2110 3.4105
R16428 GNDA.n2358 GNDA.n2110 3.4105
R16429 GNDA.n2142 GNDA.n2110 3.4105
R16430 GNDA.n2360 GNDA.n2110 3.4105
R16431 GNDA.n2141 GNDA.n2110 3.4105
R16432 GNDA.n2362 GNDA.n2110 3.4105
R16433 GNDA.n2140 GNDA.n2110 3.4105
R16434 GNDA.n2364 GNDA.n2110 3.4105
R16435 GNDA.n2139 GNDA.n2110 3.4105
R16436 GNDA.n2366 GNDA.n2110 3.4105
R16437 GNDA.n2138 GNDA.n2110 3.4105
R16438 GNDA.n2368 GNDA.n2110 3.4105
R16439 GNDA.n2137 GNDA.n2110 3.4105
R16440 GNDA.n2370 GNDA.n2110 3.4105
R16441 GNDA.n2136 GNDA.n2110 3.4105
R16442 GNDA.n2372 GNDA.n2110 3.4105
R16443 GNDA.n2135 GNDA.n2110 3.4105
R16444 GNDA.n2374 GNDA.n2110 3.4105
R16445 GNDA.n2110 GNDA.n2066 3.4105
R16446 GNDA.n2377 GNDA.n2110 3.4105
R16447 GNDA.n2344 GNDA.n2070 3.4105
R16448 GNDA.n2149 GNDA.n2070 3.4105
R16449 GNDA.n2346 GNDA.n2070 3.4105
R16450 GNDA.n2148 GNDA.n2070 3.4105
R16451 GNDA.n2348 GNDA.n2070 3.4105
R16452 GNDA.n2147 GNDA.n2070 3.4105
R16453 GNDA.n2350 GNDA.n2070 3.4105
R16454 GNDA.n2146 GNDA.n2070 3.4105
R16455 GNDA.n2352 GNDA.n2070 3.4105
R16456 GNDA.n2145 GNDA.n2070 3.4105
R16457 GNDA.n2354 GNDA.n2070 3.4105
R16458 GNDA.n2144 GNDA.n2070 3.4105
R16459 GNDA.n2356 GNDA.n2070 3.4105
R16460 GNDA.n2143 GNDA.n2070 3.4105
R16461 GNDA.n2358 GNDA.n2070 3.4105
R16462 GNDA.n2142 GNDA.n2070 3.4105
R16463 GNDA.n2360 GNDA.n2070 3.4105
R16464 GNDA.n2141 GNDA.n2070 3.4105
R16465 GNDA.n2362 GNDA.n2070 3.4105
R16466 GNDA.n2140 GNDA.n2070 3.4105
R16467 GNDA.n2364 GNDA.n2070 3.4105
R16468 GNDA.n2139 GNDA.n2070 3.4105
R16469 GNDA.n2366 GNDA.n2070 3.4105
R16470 GNDA.n2138 GNDA.n2070 3.4105
R16471 GNDA.n2368 GNDA.n2070 3.4105
R16472 GNDA.n2137 GNDA.n2070 3.4105
R16473 GNDA.n2370 GNDA.n2070 3.4105
R16474 GNDA.n2136 GNDA.n2070 3.4105
R16475 GNDA.n2372 GNDA.n2070 3.4105
R16476 GNDA.n2135 GNDA.n2070 3.4105
R16477 GNDA.n2374 GNDA.n2070 3.4105
R16478 GNDA.n2070 GNDA.n2066 3.4105
R16479 GNDA.n2377 GNDA.n2070 3.4105
R16480 GNDA.n2344 GNDA.n2112 3.4105
R16481 GNDA.n2149 GNDA.n2112 3.4105
R16482 GNDA.n2346 GNDA.n2112 3.4105
R16483 GNDA.n2148 GNDA.n2112 3.4105
R16484 GNDA.n2348 GNDA.n2112 3.4105
R16485 GNDA.n2147 GNDA.n2112 3.4105
R16486 GNDA.n2350 GNDA.n2112 3.4105
R16487 GNDA.n2146 GNDA.n2112 3.4105
R16488 GNDA.n2352 GNDA.n2112 3.4105
R16489 GNDA.n2145 GNDA.n2112 3.4105
R16490 GNDA.n2354 GNDA.n2112 3.4105
R16491 GNDA.n2144 GNDA.n2112 3.4105
R16492 GNDA.n2356 GNDA.n2112 3.4105
R16493 GNDA.n2143 GNDA.n2112 3.4105
R16494 GNDA.n2358 GNDA.n2112 3.4105
R16495 GNDA.n2142 GNDA.n2112 3.4105
R16496 GNDA.n2360 GNDA.n2112 3.4105
R16497 GNDA.n2141 GNDA.n2112 3.4105
R16498 GNDA.n2362 GNDA.n2112 3.4105
R16499 GNDA.n2140 GNDA.n2112 3.4105
R16500 GNDA.n2364 GNDA.n2112 3.4105
R16501 GNDA.n2139 GNDA.n2112 3.4105
R16502 GNDA.n2366 GNDA.n2112 3.4105
R16503 GNDA.n2138 GNDA.n2112 3.4105
R16504 GNDA.n2368 GNDA.n2112 3.4105
R16505 GNDA.n2137 GNDA.n2112 3.4105
R16506 GNDA.n2370 GNDA.n2112 3.4105
R16507 GNDA.n2136 GNDA.n2112 3.4105
R16508 GNDA.n2372 GNDA.n2112 3.4105
R16509 GNDA.n2135 GNDA.n2112 3.4105
R16510 GNDA.n2374 GNDA.n2112 3.4105
R16511 GNDA.n2112 GNDA.n2066 3.4105
R16512 GNDA.n2377 GNDA.n2112 3.4105
R16513 GNDA.n2344 GNDA.n2069 3.4105
R16514 GNDA.n2149 GNDA.n2069 3.4105
R16515 GNDA.n2346 GNDA.n2069 3.4105
R16516 GNDA.n2148 GNDA.n2069 3.4105
R16517 GNDA.n2348 GNDA.n2069 3.4105
R16518 GNDA.n2147 GNDA.n2069 3.4105
R16519 GNDA.n2350 GNDA.n2069 3.4105
R16520 GNDA.n2146 GNDA.n2069 3.4105
R16521 GNDA.n2352 GNDA.n2069 3.4105
R16522 GNDA.n2145 GNDA.n2069 3.4105
R16523 GNDA.n2354 GNDA.n2069 3.4105
R16524 GNDA.n2144 GNDA.n2069 3.4105
R16525 GNDA.n2356 GNDA.n2069 3.4105
R16526 GNDA.n2143 GNDA.n2069 3.4105
R16527 GNDA.n2358 GNDA.n2069 3.4105
R16528 GNDA.n2142 GNDA.n2069 3.4105
R16529 GNDA.n2360 GNDA.n2069 3.4105
R16530 GNDA.n2141 GNDA.n2069 3.4105
R16531 GNDA.n2362 GNDA.n2069 3.4105
R16532 GNDA.n2140 GNDA.n2069 3.4105
R16533 GNDA.n2364 GNDA.n2069 3.4105
R16534 GNDA.n2139 GNDA.n2069 3.4105
R16535 GNDA.n2366 GNDA.n2069 3.4105
R16536 GNDA.n2138 GNDA.n2069 3.4105
R16537 GNDA.n2368 GNDA.n2069 3.4105
R16538 GNDA.n2137 GNDA.n2069 3.4105
R16539 GNDA.n2370 GNDA.n2069 3.4105
R16540 GNDA.n2136 GNDA.n2069 3.4105
R16541 GNDA.n2372 GNDA.n2069 3.4105
R16542 GNDA.n2135 GNDA.n2069 3.4105
R16543 GNDA.n2374 GNDA.n2069 3.4105
R16544 GNDA.n2069 GNDA.n2066 3.4105
R16545 GNDA.n2377 GNDA.n2069 3.4105
R16546 GNDA.n2344 GNDA.n2114 3.4105
R16547 GNDA.n2149 GNDA.n2114 3.4105
R16548 GNDA.n2346 GNDA.n2114 3.4105
R16549 GNDA.n2148 GNDA.n2114 3.4105
R16550 GNDA.n2348 GNDA.n2114 3.4105
R16551 GNDA.n2147 GNDA.n2114 3.4105
R16552 GNDA.n2350 GNDA.n2114 3.4105
R16553 GNDA.n2146 GNDA.n2114 3.4105
R16554 GNDA.n2352 GNDA.n2114 3.4105
R16555 GNDA.n2145 GNDA.n2114 3.4105
R16556 GNDA.n2354 GNDA.n2114 3.4105
R16557 GNDA.n2144 GNDA.n2114 3.4105
R16558 GNDA.n2356 GNDA.n2114 3.4105
R16559 GNDA.n2143 GNDA.n2114 3.4105
R16560 GNDA.n2358 GNDA.n2114 3.4105
R16561 GNDA.n2142 GNDA.n2114 3.4105
R16562 GNDA.n2360 GNDA.n2114 3.4105
R16563 GNDA.n2141 GNDA.n2114 3.4105
R16564 GNDA.n2362 GNDA.n2114 3.4105
R16565 GNDA.n2140 GNDA.n2114 3.4105
R16566 GNDA.n2364 GNDA.n2114 3.4105
R16567 GNDA.n2139 GNDA.n2114 3.4105
R16568 GNDA.n2366 GNDA.n2114 3.4105
R16569 GNDA.n2138 GNDA.n2114 3.4105
R16570 GNDA.n2368 GNDA.n2114 3.4105
R16571 GNDA.n2137 GNDA.n2114 3.4105
R16572 GNDA.n2370 GNDA.n2114 3.4105
R16573 GNDA.n2136 GNDA.n2114 3.4105
R16574 GNDA.n2372 GNDA.n2114 3.4105
R16575 GNDA.n2135 GNDA.n2114 3.4105
R16576 GNDA.n2374 GNDA.n2114 3.4105
R16577 GNDA.n2114 GNDA.n2066 3.4105
R16578 GNDA.n2377 GNDA.n2114 3.4105
R16579 GNDA.n2344 GNDA.n2068 3.4105
R16580 GNDA.n2149 GNDA.n2068 3.4105
R16581 GNDA.n2346 GNDA.n2068 3.4105
R16582 GNDA.n2148 GNDA.n2068 3.4105
R16583 GNDA.n2348 GNDA.n2068 3.4105
R16584 GNDA.n2147 GNDA.n2068 3.4105
R16585 GNDA.n2350 GNDA.n2068 3.4105
R16586 GNDA.n2146 GNDA.n2068 3.4105
R16587 GNDA.n2352 GNDA.n2068 3.4105
R16588 GNDA.n2145 GNDA.n2068 3.4105
R16589 GNDA.n2354 GNDA.n2068 3.4105
R16590 GNDA.n2144 GNDA.n2068 3.4105
R16591 GNDA.n2356 GNDA.n2068 3.4105
R16592 GNDA.n2143 GNDA.n2068 3.4105
R16593 GNDA.n2358 GNDA.n2068 3.4105
R16594 GNDA.n2142 GNDA.n2068 3.4105
R16595 GNDA.n2360 GNDA.n2068 3.4105
R16596 GNDA.n2141 GNDA.n2068 3.4105
R16597 GNDA.n2362 GNDA.n2068 3.4105
R16598 GNDA.n2140 GNDA.n2068 3.4105
R16599 GNDA.n2364 GNDA.n2068 3.4105
R16600 GNDA.n2139 GNDA.n2068 3.4105
R16601 GNDA.n2366 GNDA.n2068 3.4105
R16602 GNDA.n2138 GNDA.n2068 3.4105
R16603 GNDA.n2368 GNDA.n2068 3.4105
R16604 GNDA.n2137 GNDA.n2068 3.4105
R16605 GNDA.n2370 GNDA.n2068 3.4105
R16606 GNDA.n2136 GNDA.n2068 3.4105
R16607 GNDA.n2372 GNDA.n2068 3.4105
R16608 GNDA.n2135 GNDA.n2068 3.4105
R16609 GNDA.n2374 GNDA.n2068 3.4105
R16610 GNDA.n2068 GNDA.n2066 3.4105
R16611 GNDA.n2377 GNDA.n2068 3.4105
R16612 GNDA.n2344 GNDA.n2116 3.4105
R16613 GNDA.n2149 GNDA.n2116 3.4105
R16614 GNDA.n2346 GNDA.n2116 3.4105
R16615 GNDA.n2148 GNDA.n2116 3.4105
R16616 GNDA.n2348 GNDA.n2116 3.4105
R16617 GNDA.n2147 GNDA.n2116 3.4105
R16618 GNDA.n2350 GNDA.n2116 3.4105
R16619 GNDA.n2146 GNDA.n2116 3.4105
R16620 GNDA.n2352 GNDA.n2116 3.4105
R16621 GNDA.n2145 GNDA.n2116 3.4105
R16622 GNDA.n2354 GNDA.n2116 3.4105
R16623 GNDA.n2144 GNDA.n2116 3.4105
R16624 GNDA.n2356 GNDA.n2116 3.4105
R16625 GNDA.n2143 GNDA.n2116 3.4105
R16626 GNDA.n2358 GNDA.n2116 3.4105
R16627 GNDA.n2142 GNDA.n2116 3.4105
R16628 GNDA.n2360 GNDA.n2116 3.4105
R16629 GNDA.n2141 GNDA.n2116 3.4105
R16630 GNDA.n2362 GNDA.n2116 3.4105
R16631 GNDA.n2140 GNDA.n2116 3.4105
R16632 GNDA.n2364 GNDA.n2116 3.4105
R16633 GNDA.n2139 GNDA.n2116 3.4105
R16634 GNDA.n2366 GNDA.n2116 3.4105
R16635 GNDA.n2138 GNDA.n2116 3.4105
R16636 GNDA.n2368 GNDA.n2116 3.4105
R16637 GNDA.n2137 GNDA.n2116 3.4105
R16638 GNDA.n2370 GNDA.n2116 3.4105
R16639 GNDA.n2136 GNDA.n2116 3.4105
R16640 GNDA.n2372 GNDA.n2116 3.4105
R16641 GNDA.n2135 GNDA.n2116 3.4105
R16642 GNDA.n2374 GNDA.n2116 3.4105
R16643 GNDA.n2116 GNDA.n2066 3.4105
R16644 GNDA.n2377 GNDA.n2116 3.4105
R16645 GNDA.n2344 GNDA.n2067 3.4105
R16646 GNDA.n2149 GNDA.n2067 3.4105
R16647 GNDA.n2346 GNDA.n2067 3.4105
R16648 GNDA.n2148 GNDA.n2067 3.4105
R16649 GNDA.n2348 GNDA.n2067 3.4105
R16650 GNDA.n2147 GNDA.n2067 3.4105
R16651 GNDA.n2350 GNDA.n2067 3.4105
R16652 GNDA.n2146 GNDA.n2067 3.4105
R16653 GNDA.n2352 GNDA.n2067 3.4105
R16654 GNDA.n2145 GNDA.n2067 3.4105
R16655 GNDA.n2354 GNDA.n2067 3.4105
R16656 GNDA.n2144 GNDA.n2067 3.4105
R16657 GNDA.n2356 GNDA.n2067 3.4105
R16658 GNDA.n2143 GNDA.n2067 3.4105
R16659 GNDA.n2358 GNDA.n2067 3.4105
R16660 GNDA.n2142 GNDA.n2067 3.4105
R16661 GNDA.n2360 GNDA.n2067 3.4105
R16662 GNDA.n2141 GNDA.n2067 3.4105
R16663 GNDA.n2362 GNDA.n2067 3.4105
R16664 GNDA.n2140 GNDA.n2067 3.4105
R16665 GNDA.n2364 GNDA.n2067 3.4105
R16666 GNDA.n2139 GNDA.n2067 3.4105
R16667 GNDA.n2366 GNDA.n2067 3.4105
R16668 GNDA.n2138 GNDA.n2067 3.4105
R16669 GNDA.n2368 GNDA.n2067 3.4105
R16670 GNDA.n2137 GNDA.n2067 3.4105
R16671 GNDA.n2370 GNDA.n2067 3.4105
R16672 GNDA.n2136 GNDA.n2067 3.4105
R16673 GNDA.n2372 GNDA.n2067 3.4105
R16674 GNDA.n2135 GNDA.n2067 3.4105
R16675 GNDA.n2374 GNDA.n2067 3.4105
R16676 GNDA.n2067 GNDA.n2066 3.4105
R16677 GNDA.n2377 GNDA.n2067 3.4105
R16678 GNDA.n2376 GNDA.n2344 3.4105
R16679 GNDA.n2376 GNDA.n2149 3.4105
R16680 GNDA.n2376 GNDA.n2346 3.4105
R16681 GNDA.n2376 GNDA.n2148 3.4105
R16682 GNDA.n2376 GNDA.n2348 3.4105
R16683 GNDA.n2376 GNDA.n2147 3.4105
R16684 GNDA.n2376 GNDA.n2350 3.4105
R16685 GNDA.n2376 GNDA.n2146 3.4105
R16686 GNDA.n2376 GNDA.n2352 3.4105
R16687 GNDA.n2376 GNDA.n2145 3.4105
R16688 GNDA.n2376 GNDA.n2354 3.4105
R16689 GNDA.n2376 GNDA.n2144 3.4105
R16690 GNDA.n2376 GNDA.n2356 3.4105
R16691 GNDA.n2376 GNDA.n2143 3.4105
R16692 GNDA.n2376 GNDA.n2358 3.4105
R16693 GNDA.n2376 GNDA.n2142 3.4105
R16694 GNDA.n2376 GNDA.n2360 3.4105
R16695 GNDA.n2376 GNDA.n2141 3.4105
R16696 GNDA.n2376 GNDA.n2362 3.4105
R16697 GNDA.n2376 GNDA.n2140 3.4105
R16698 GNDA.n2376 GNDA.n2364 3.4105
R16699 GNDA.n2376 GNDA.n2139 3.4105
R16700 GNDA.n2376 GNDA.n2366 3.4105
R16701 GNDA.n2376 GNDA.n2138 3.4105
R16702 GNDA.n2376 GNDA.n2368 3.4105
R16703 GNDA.n2376 GNDA.n2137 3.4105
R16704 GNDA.n2376 GNDA.n2370 3.4105
R16705 GNDA.n2376 GNDA.n2136 3.4105
R16706 GNDA.n2376 GNDA.n2372 3.4105
R16707 GNDA.n2376 GNDA.n2135 3.4105
R16708 GNDA.n2376 GNDA.n2374 3.4105
R16709 GNDA.n2377 GNDA.n2376 3.4105
R16710 GNDA.n2048 GNDA.n1984 3.4105
R16711 GNDA.n2409 GNDA.n1984 3.4105
R16712 GNDA.n2429 GNDA.n1984 3.4105
R16713 GNDA.n2428 GNDA.n2380 3.4105
R16714 GNDA.n2428 GNDA.n2047 3.4105
R16715 GNDA.n2428 GNDA.n2382 3.4105
R16716 GNDA.n2428 GNDA.n2046 3.4105
R16717 GNDA.n2428 GNDA.n2384 3.4105
R16718 GNDA.n2428 GNDA.n2045 3.4105
R16719 GNDA.n2428 GNDA.n2386 3.4105
R16720 GNDA.n2428 GNDA.n2044 3.4105
R16721 GNDA.n2428 GNDA.n2388 3.4105
R16722 GNDA.n2428 GNDA.n2043 3.4105
R16723 GNDA.n2428 GNDA.n2390 3.4105
R16724 GNDA.n2428 GNDA.n2042 3.4105
R16725 GNDA.n2428 GNDA.n2392 3.4105
R16726 GNDA.n2428 GNDA.n2041 3.4105
R16727 GNDA.n2428 GNDA.n2394 3.4105
R16728 GNDA.n2428 GNDA.n2040 3.4105
R16729 GNDA.n2428 GNDA.n2396 3.4105
R16730 GNDA.n2428 GNDA.n2039 3.4105
R16731 GNDA.n2428 GNDA.n2398 3.4105
R16732 GNDA.n2428 GNDA.n2038 3.4105
R16733 GNDA.n2428 GNDA.n2400 3.4105
R16734 GNDA.n2428 GNDA.n2037 3.4105
R16735 GNDA.n2428 GNDA.n2402 3.4105
R16736 GNDA.n2428 GNDA.n2036 3.4105
R16737 GNDA.n2428 GNDA.n2404 3.4105
R16738 GNDA.n2428 GNDA.n2035 3.4105
R16739 GNDA.n2428 GNDA.n2406 3.4105
R16740 GNDA.n2428 GNDA.n2034 3.4105
R16741 GNDA.n2428 GNDA.n2408 3.4105
R16742 GNDA.n2428 GNDA.n2409 3.4105
R16743 GNDA.n2429 GNDA.n2428 3.4105
R16744 GNDA.n2431 GNDA.n2000 3.4105
R16745 GNDA.n2048 GNDA.n2000 3.4105
R16746 GNDA.n2380 GNDA.n2000 3.4105
R16747 GNDA.n2047 GNDA.n2000 3.4105
R16748 GNDA.n2382 GNDA.n2000 3.4105
R16749 GNDA.n2046 GNDA.n2000 3.4105
R16750 GNDA.n2384 GNDA.n2000 3.4105
R16751 GNDA.n2045 GNDA.n2000 3.4105
R16752 GNDA.n2386 GNDA.n2000 3.4105
R16753 GNDA.n2044 GNDA.n2000 3.4105
R16754 GNDA.n2388 GNDA.n2000 3.4105
R16755 GNDA.n2043 GNDA.n2000 3.4105
R16756 GNDA.n2390 GNDA.n2000 3.4105
R16757 GNDA.n2042 GNDA.n2000 3.4105
R16758 GNDA.n2392 GNDA.n2000 3.4105
R16759 GNDA.n2041 GNDA.n2000 3.4105
R16760 GNDA.n2394 GNDA.n2000 3.4105
R16761 GNDA.n2040 GNDA.n2000 3.4105
R16762 GNDA.n2396 GNDA.n2000 3.4105
R16763 GNDA.n2039 GNDA.n2000 3.4105
R16764 GNDA.n2398 GNDA.n2000 3.4105
R16765 GNDA.n2038 GNDA.n2000 3.4105
R16766 GNDA.n2400 GNDA.n2000 3.4105
R16767 GNDA.n2037 GNDA.n2000 3.4105
R16768 GNDA.n2402 GNDA.n2000 3.4105
R16769 GNDA.n2036 GNDA.n2000 3.4105
R16770 GNDA.n2404 GNDA.n2000 3.4105
R16771 GNDA.n2035 GNDA.n2000 3.4105
R16772 GNDA.n2406 GNDA.n2000 3.4105
R16773 GNDA.n2034 GNDA.n2000 3.4105
R16774 GNDA.n2408 GNDA.n2000 3.4105
R16775 GNDA.n2409 GNDA.n2000 3.4105
R16776 GNDA.n2429 GNDA.n2000 3.4105
R16777 GNDA.n2431 GNDA.n2002 3.4105
R16778 GNDA.n2048 GNDA.n2002 3.4105
R16779 GNDA.n2380 GNDA.n2002 3.4105
R16780 GNDA.n2047 GNDA.n2002 3.4105
R16781 GNDA.n2382 GNDA.n2002 3.4105
R16782 GNDA.n2046 GNDA.n2002 3.4105
R16783 GNDA.n2384 GNDA.n2002 3.4105
R16784 GNDA.n2045 GNDA.n2002 3.4105
R16785 GNDA.n2386 GNDA.n2002 3.4105
R16786 GNDA.n2044 GNDA.n2002 3.4105
R16787 GNDA.n2388 GNDA.n2002 3.4105
R16788 GNDA.n2043 GNDA.n2002 3.4105
R16789 GNDA.n2390 GNDA.n2002 3.4105
R16790 GNDA.n2042 GNDA.n2002 3.4105
R16791 GNDA.n2392 GNDA.n2002 3.4105
R16792 GNDA.n2041 GNDA.n2002 3.4105
R16793 GNDA.n2394 GNDA.n2002 3.4105
R16794 GNDA.n2040 GNDA.n2002 3.4105
R16795 GNDA.n2396 GNDA.n2002 3.4105
R16796 GNDA.n2039 GNDA.n2002 3.4105
R16797 GNDA.n2398 GNDA.n2002 3.4105
R16798 GNDA.n2038 GNDA.n2002 3.4105
R16799 GNDA.n2400 GNDA.n2002 3.4105
R16800 GNDA.n2037 GNDA.n2002 3.4105
R16801 GNDA.n2402 GNDA.n2002 3.4105
R16802 GNDA.n2036 GNDA.n2002 3.4105
R16803 GNDA.n2404 GNDA.n2002 3.4105
R16804 GNDA.n2035 GNDA.n2002 3.4105
R16805 GNDA.n2406 GNDA.n2002 3.4105
R16806 GNDA.n2034 GNDA.n2002 3.4105
R16807 GNDA.n2408 GNDA.n2002 3.4105
R16808 GNDA.n2409 GNDA.n2002 3.4105
R16809 GNDA.n2429 GNDA.n2002 3.4105
R16810 GNDA.n2431 GNDA.n1999 3.4105
R16811 GNDA.n2048 GNDA.n1999 3.4105
R16812 GNDA.n2380 GNDA.n1999 3.4105
R16813 GNDA.n2047 GNDA.n1999 3.4105
R16814 GNDA.n2382 GNDA.n1999 3.4105
R16815 GNDA.n2046 GNDA.n1999 3.4105
R16816 GNDA.n2384 GNDA.n1999 3.4105
R16817 GNDA.n2045 GNDA.n1999 3.4105
R16818 GNDA.n2386 GNDA.n1999 3.4105
R16819 GNDA.n2044 GNDA.n1999 3.4105
R16820 GNDA.n2388 GNDA.n1999 3.4105
R16821 GNDA.n2043 GNDA.n1999 3.4105
R16822 GNDA.n2390 GNDA.n1999 3.4105
R16823 GNDA.n2042 GNDA.n1999 3.4105
R16824 GNDA.n2392 GNDA.n1999 3.4105
R16825 GNDA.n2041 GNDA.n1999 3.4105
R16826 GNDA.n2394 GNDA.n1999 3.4105
R16827 GNDA.n2040 GNDA.n1999 3.4105
R16828 GNDA.n2396 GNDA.n1999 3.4105
R16829 GNDA.n2039 GNDA.n1999 3.4105
R16830 GNDA.n2398 GNDA.n1999 3.4105
R16831 GNDA.n2038 GNDA.n1999 3.4105
R16832 GNDA.n2400 GNDA.n1999 3.4105
R16833 GNDA.n2037 GNDA.n1999 3.4105
R16834 GNDA.n2402 GNDA.n1999 3.4105
R16835 GNDA.n2036 GNDA.n1999 3.4105
R16836 GNDA.n2404 GNDA.n1999 3.4105
R16837 GNDA.n2035 GNDA.n1999 3.4105
R16838 GNDA.n2406 GNDA.n1999 3.4105
R16839 GNDA.n2034 GNDA.n1999 3.4105
R16840 GNDA.n2408 GNDA.n1999 3.4105
R16841 GNDA.n2409 GNDA.n1999 3.4105
R16842 GNDA.n2429 GNDA.n1999 3.4105
R16843 GNDA.n2431 GNDA.n2003 3.4105
R16844 GNDA.n2048 GNDA.n2003 3.4105
R16845 GNDA.n2380 GNDA.n2003 3.4105
R16846 GNDA.n2047 GNDA.n2003 3.4105
R16847 GNDA.n2382 GNDA.n2003 3.4105
R16848 GNDA.n2046 GNDA.n2003 3.4105
R16849 GNDA.n2384 GNDA.n2003 3.4105
R16850 GNDA.n2045 GNDA.n2003 3.4105
R16851 GNDA.n2386 GNDA.n2003 3.4105
R16852 GNDA.n2044 GNDA.n2003 3.4105
R16853 GNDA.n2388 GNDA.n2003 3.4105
R16854 GNDA.n2043 GNDA.n2003 3.4105
R16855 GNDA.n2390 GNDA.n2003 3.4105
R16856 GNDA.n2042 GNDA.n2003 3.4105
R16857 GNDA.n2392 GNDA.n2003 3.4105
R16858 GNDA.n2041 GNDA.n2003 3.4105
R16859 GNDA.n2394 GNDA.n2003 3.4105
R16860 GNDA.n2040 GNDA.n2003 3.4105
R16861 GNDA.n2396 GNDA.n2003 3.4105
R16862 GNDA.n2039 GNDA.n2003 3.4105
R16863 GNDA.n2398 GNDA.n2003 3.4105
R16864 GNDA.n2038 GNDA.n2003 3.4105
R16865 GNDA.n2400 GNDA.n2003 3.4105
R16866 GNDA.n2037 GNDA.n2003 3.4105
R16867 GNDA.n2402 GNDA.n2003 3.4105
R16868 GNDA.n2036 GNDA.n2003 3.4105
R16869 GNDA.n2404 GNDA.n2003 3.4105
R16870 GNDA.n2035 GNDA.n2003 3.4105
R16871 GNDA.n2406 GNDA.n2003 3.4105
R16872 GNDA.n2034 GNDA.n2003 3.4105
R16873 GNDA.n2408 GNDA.n2003 3.4105
R16874 GNDA.n2409 GNDA.n2003 3.4105
R16875 GNDA.n2429 GNDA.n2003 3.4105
R16876 GNDA.n2431 GNDA.n1998 3.4105
R16877 GNDA.n2048 GNDA.n1998 3.4105
R16878 GNDA.n2380 GNDA.n1998 3.4105
R16879 GNDA.n2047 GNDA.n1998 3.4105
R16880 GNDA.n2382 GNDA.n1998 3.4105
R16881 GNDA.n2046 GNDA.n1998 3.4105
R16882 GNDA.n2384 GNDA.n1998 3.4105
R16883 GNDA.n2045 GNDA.n1998 3.4105
R16884 GNDA.n2386 GNDA.n1998 3.4105
R16885 GNDA.n2044 GNDA.n1998 3.4105
R16886 GNDA.n2388 GNDA.n1998 3.4105
R16887 GNDA.n2043 GNDA.n1998 3.4105
R16888 GNDA.n2390 GNDA.n1998 3.4105
R16889 GNDA.n2042 GNDA.n1998 3.4105
R16890 GNDA.n2392 GNDA.n1998 3.4105
R16891 GNDA.n2041 GNDA.n1998 3.4105
R16892 GNDA.n2394 GNDA.n1998 3.4105
R16893 GNDA.n2040 GNDA.n1998 3.4105
R16894 GNDA.n2396 GNDA.n1998 3.4105
R16895 GNDA.n2039 GNDA.n1998 3.4105
R16896 GNDA.n2398 GNDA.n1998 3.4105
R16897 GNDA.n2038 GNDA.n1998 3.4105
R16898 GNDA.n2400 GNDA.n1998 3.4105
R16899 GNDA.n2037 GNDA.n1998 3.4105
R16900 GNDA.n2402 GNDA.n1998 3.4105
R16901 GNDA.n2036 GNDA.n1998 3.4105
R16902 GNDA.n2404 GNDA.n1998 3.4105
R16903 GNDA.n2035 GNDA.n1998 3.4105
R16904 GNDA.n2406 GNDA.n1998 3.4105
R16905 GNDA.n2034 GNDA.n1998 3.4105
R16906 GNDA.n2408 GNDA.n1998 3.4105
R16907 GNDA.n2409 GNDA.n1998 3.4105
R16908 GNDA.n2429 GNDA.n1998 3.4105
R16909 GNDA.n2431 GNDA.n2004 3.4105
R16910 GNDA.n2048 GNDA.n2004 3.4105
R16911 GNDA.n2380 GNDA.n2004 3.4105
R16912 GNDA.n2047 GNDA.n2004 3.4105
R16913 GNDA.n2382 GNDA.n2004 3.4105
R16914 GNDA.n2046 GNDA.n2004 3.4105
R16915 GNDA.n2384 GNDA.n2004 3.4105
R16916 GNDA.n2045 GNDA.n2004 3.4105
R16917 GNDA.n2386 GNDA.n2004 3.4105
R16918 GNDA.n2044 GNDA.n2004 3.4105
R16919 GNDA.n2388 GNDA.n2004 3.4105
R16920 GNDA.n2043 GNDA.n2004 3.4105
R16921 GNDA.n2390 GNDA.n2004 3.4105
R16922 GNDA.n2042 GNDA.n2004 3.4105
R16923 GNDA.n2392 GNDA.n2004 3.4105
R16924 GNDA.n2041 GNDA.n2004 3.4105
R16925 GNDA.n2394 GNDA.n2004 3.4105
R16926 GNDA.n2040 GNDA.n2004 3.4105
R16927 GNDA.n2396 GNDA.n2004 3.4105
R16928 GNDA.n2039 GNDA.n2004 3.4105
R16929 GNDA.n2398 GNDA.n2004 3.4105
R16930 GNDA.n2038 GNDA.n2004 3.4105
R16931 GNDA.n2400 GNDA.n2004 3.4105
R16932 GNDA.n2037 GNDA.n2004 3.4105
R16933 GNDA.n2402 GNDA.n2004 3.4105
R16934 GNDA.n2036 GNDA.n2004 3.4105
R16935 GNDA.n2404 GNDA.n2004 3.4105
R16936 GNDA.n2035 GNDA.n2004 3.4105
R16937 GNDA.n2406 GNDA.n2004 3.4105
R16938 GNDA.n2034 GNDA.n2004 3.4105
R16939 GNDA.n2408 GNDA.n2004 3.4105
R16940 GNDA.n2409 GNDA.n2004 3.4105
R16941 GNDA.n2429 GNDA.n2004 3.4105
R16942 GNDA.n2431 GNDA.n1997 3.4105
R16943 GNDA.n2048 GNDA.n1997 3.4105
R16944 GNDA.n2380 GNDA.n1997 3.4105
R16945 GNDA.n2047 GNDA.n1997 3.4105
R16946 GNDA.n2382 GNDA.n1997 3.4105
R16947 GNDA.n2046 GNDA.n1997 3.4105
R16948 GNDA.n2384 GNDA.n1997 3.4105
R16949 GNDA.n2045 GNDA.n1997 3.4105
R16950 GNDA.n2386 GNDA.n1997 3.4105
R16951 GNDA.n2044 GNDA.n1997 3.4105
R16952 GNDA.n2388 GNDA.n1997 3.4105
R16953 GNDA.n2043 GNDA.n1997 3.4105
R16954 GNDA.n2390 GNDA.n1997 3.4105
R16955 GNDA.n2042 GNDA.n1997 3.4105
R16956 GNDA.n2392 GNDA.n1997 3.4105
R16957 GNDA.n2041 GNDA.n1997 3.4105
R16958 GNDA.n2394 GNDA.n1997 3.4105
R16959 GNDA.n2040 GNDA.n1997 3.4105
R16960 GNDA.n2396 GNDA.n1997 3.4105
R16961 GNDA.n2039 GNDA.n1997 3.4105
R16962 GNDA.n2398 GNDA.n1997 3.4105
R16963 GNDA.n2038 GNDA.n1997 3.4105
R16964 GNDA.n2400 GNDA.n1997 3.4105
R16965 GNDA.n2037 GNDA.n1997 3.4105
R16966 GNDA.n2402 GNDA.n1997 3.4105
R16967 GNDA.n2036 GNDA.n1997 3.4105
R16968 GNDA.n2404 GNDA.n1997 3.4105
R16969 GNDA.n2035 GNDA.n1997 3.4105
R16970 GNDA.n2406 GNDA.n1997 3.4105
R16971 GNDA.n2034 GNDA.n1997 3.4105
R16972 GNDA.n2408 GNDA.n1997 3.4105
R16973 GNDA.n2409 GNDA.n1997 3.4105
R16974 GNDA.n2429 GNDA.n1997 3.4105
R16975 GNDA.n2431 GNDA.n2005 3.4105
R16976 GNDA.n2048 GNDA.n2005 3.4105
R16977 GNDA.n2380 GNDA.n2005 3.4105
R16978 GNDA.n2047 GNDA.n2005 3.4105
R16979 GNDA.n2382 GNDA.n2005 3.4105
R16980 GNDA.n2046 GNDA.n2005 3.4105
R16981 GNDA.n2384 GNDA.n2005 3.4105
R16982 GNDA.n2045 GNDA.n2005 3.4105
R16983 GNDA.n2386 GNDA.n2005 3.4105
R16984 GNDA.n2044 GNDA.n2005 3.4105
R16985 GNDA.n2388 GNDA.n2005 3.4105
R16986 GNDA.n2043 GNDA.n2005 3.4105
R16987 GNDA.n2390 GNDA.n2005 3.4105
R16988 GNDA.n2042 GNDA.n2005 3.4105
R16989 GNDA.n2392 GNDA.n2005 3.4105
R16990 GNDA.n2041 GNDA.n2005 3.4105
R16991 GNDA.n2394 GNDA.n2005 3.4105
R16992 GNDA.n2040 GNDA.n2005 3.4105
R16993 GNDA.n2396 GNDA.n2005 3.4105
R16994 GNDA.n2039 GNDA.n2005 3.4105
R16995 GNDA.n2398 GNDA.n2005 3.4105
R16996 GNDA.n2038 GNDA.n2005 3.4105
R16997 GNDA.n2400 GNDA.n2005 3.4105
R16998 GNDA.n2037 GNDA.n2005 3.4105
R16999 GNDA.n2402 GNDA.n2005 3.4105
R17000 GNDA.n2036 GNDA.n2005 3.4105
R17001 GNDA.n2404 GNDA.n2005 3.4105
R17002 GNDA.n2035 GNDA.n2005 3.4105
R17003 GNDA.n2406 GNDA.n2005 3.4105
R17004 GNDA.n2034 GNDA.n2005 3.4105
R17005 GNDA.n2408 GNDA.n2005 3.4105
R17006 GNDA.n2409 GNDA.n2005 3.4105
R17007 GNDA.n2429 GNDA.n2005 3.4105
R17008 GNDA.n2431 GNDA.n1996 3.4105
R17009 GNDA.n2048 GNDA.n1996 3.4105
R17010 GNDA.n2380 GNDA.n1996 3.4105
R17011 GNDA.n2047 GNDA.n1996 3.4105
R17012 GNDA.n2382 GNDA.n1996 3.4105
R17013 GNDA.n2046 GNDA.n1996 3.4105
R17014 GNDA.n2384 GNDA.n1996 3.4105
R17015 GNDA.n2045 GNDA.n1996 3.4105
R17016 GNDA.n2386 GNDA.n1996 3.4105
R17017 GNDA.n2044 GNDA.n1996 3.4105
R17018 GNDA.n2388 GNDA.n1996 3.4105
R17019 GNDA.n2043 GNDA.n1996 3.4105
R17020 GNDA.n2390 GNDA.n1996 3.4105
R17021 GNDA.n2042 GNDA.n1996 3.4105
R17022 GNDA.n2392 GNDA.n1996 3.4105
R17023 GNDA.n2041 GNDA.n1996 3.4105
R17024 GNDA.n2394 GNDA.n1996 3.4105
R17025 GNDA.n2040 GNDA.n1996 3.4105
R17026 GNDA.n2396 GNDA.n1996 3.4105
R17027 GNDA.n2039 GNDA.n1996 3.4105
R17028 GNDA.n2398 GNDA.n1996 3.4105
R17029 GNDA.n2038 GNDA.n1996 3.4105
R17030 GNDA.n2400 GNDA.n1996 3.4105
R17031 GNDA.n2037 GNDA.n1996 3.4105
R17032 GNDA.n2402 GNDA.n1996 3.4105
R17033 GNDA.n2036 GNDA.n1996 3.4105
R17034 GNDA.n2404 GNDA.n1996 3.4105
R17035 GNDA.n2035 GNDA.n1996 3.4105
R17036 GNDA.n2406 GNDA.n1996 3.4105
R17037 GNDA.n2034 GNDA.n1996 3.4105
R17038 GNDA.n2408 GNDA.n1996 3.4105
R17039 GNDA.n2409 GNDA.n1996 3.4105
R17040 GNDA.n2429 GNDA.n1996 3.4105
R17041 GNDA.n2431 GNDA.n2006 3.4105
R17042 GNDA.n2048 GNDA.n2006 3.4105
R17043 GNDA.n2380 GNDA.n2006 3.4105
R17044 GNDA.n2047 GNDA.n2006 3.4105
R17045 GNDA.n2382 GNDA.n2006 3.4105
R17046 GNDA.n2046 GNDA.n2006 3.4105
R17047 GNDA.n2384 GNDA.n2006 3.4105
R17048 GNDA.n2045 GNDA.n2006 3.4105
R17049 GNDA.n2386 GNDA.n2006 3.4105
R17050 GNDA.n2044 GNDA.n2006 3.4105
R17051 GNDA.n2388 GNDA.n2006 3.4105
R17052 GNDA.n2043 GNDA.n2006 3.4105
R17053 GNDA.n2390 GNDA.n2006 3.4105
R17054 GNDA.n2042 GNDA.n2006 3.4105
R17055 GNDA.n2392 GNDA.n2006 3.4105
R17056 GNDA.n2041 GNDA.n2006 3.4105
R17057 GNDA.n2394 GNDA.n2006 3.4105
R17058 GNDA.n2040 GNDA.n2006 3.4105
R17059 GNDA.n2396 GNDA.n2006 3.4105
R17060 GNDA.n2039 GNDA.n2006 3.4105
R17061 GNDA.n2398 GNDA.n2006 3.4105
R17062 GNDA.n2038 GNDA.n2006 3.4105
R17063 GNDA.n2400 GNDA.n2006 3.4105
R17064 GNDA.n2037 GNDA.n2006 3.4105
R17065 GNDA.n2402 GNDA.n2006 3.4105
R17066 GNDA.n2036 GNDA.n2006 3.4105
R17067 GNDA.n2404 GNDA.n2006 3.4105
R17068 GNDA.n2035 GNDA.n2006 3.4105
R17069 GNDA.n2406 GNDA.n2006 3.4105
R17070 GNDA.n2034 GNDA.n2006 3.4105
R17071 GNDA.n2408 GNDA.n2006 3.4105
R17072 GNDA.n2409 GNDA.n2006 3.4105
R17073 GNDA.n2429 GNDA.n2006 3.4105
R17074 GNDA.n2431 GNDA.n1995 3.4105
R17075 GNDA.n2048 GNDA.n1995 3.4105
R17076 GNDA.n2380 GNDA.n1995 3.4105
R17077 GNDA.n2047 GNDA.n1995 3.4105
R17078 GNDA.n2382 GNDA.n1995 3.4105
R17079 GNDA.n2046 GNDA.n1995 3.4105
R17080 GNDA.n2384 GNDA.n1995 3.4105
R17081 GNDA.n2045 GNDA.n1995 3.4105
R17082 GNDA.n2386 GNDA.n1995 3.4105
R17083 GNDA.n2044 GNDA.n1995 3.4105
R17084 GNDA.n2388 GNDA.n1995 3.4105
R17085 GNDA.n2043 GNDA.n1995 3.4105
R17086 GNDA.n2390 GNDA.n1995 3.4105
R17087 GNDA.n2042 GNDA.n1995 3.4105
R17088 GNDA.n2392 GNDA.n1995 3.4105
R17089 GNDA.n2041 GNDA.n1995 3.4105
R17090 GNDA.n2394 GNDA.n1995 3.4105
R17091 GNDA.n2040 GNDA.n1995 3.4105
R17092 GNDA.n2396 GNDA.n1995 3.4105
R17093 GNDA.n2039 GNDA.n1995 3.4105
R17094 GNDA.n2398 GNDA.n1995 3.4105
R17095 GNDA.n2038 GNDA.n1995 3.4105
R17096 GNDA.n2400 GNDA.n1995 3.4105
R17097 GNDA.n2037 GNDA.n1995 3.4105
R17098 GNDA.n2402 GNDA.n1995 3.4105
R17099 GNDA.n2036 GNDA.n1995 3.4105
R17100 GNDA.n2404 GNDA.n1995 3.4105
R17101 GNDA.n2035 GNDA.n1995 3.4105
R17102 GNDA.n2406 GNDA.n1995 3.4105
R17103 GNDA.n2034 GNDA.n1995 3.4105
R17104 GNDA.n2408 GNDA.n1995 3.4105
R17105 GNDA.n2409 GNDA.n1995 3.4105
R17106 GNDA.n2429 GNDA.n1995 3.4105
R17107 GNDA.n2431 GNDA.n2007 3.4105
R17108 GNDA.n2048 GNDA.n2007 3.4105
R17109 GNDA.n2380 GNDA.n2007 3.4105
R17110 GNDA.n2047 GNDA.n2007 3.4105
R17111 GNDA.n2382 GNDA.n2007 3.4105
R17112 GNDA.n2046 GNDA.n2007 3.4105
R17113 GNDA.n2384 GNDA.n2007 3.4105
R17114 GNDA.n2045 GNDA.n2007 3.4105
R17115 GNDA.n2386 GNDA.n2007 3.4105
R17116 GNDA.n2044 GNDA.n2007 3.4105
R17117 GNDA.n2388 GNDA.n2007 3.4105
R17118 GNDA.n2043 GNDA.n2007 3.4105
R17119 GNDA.n2390 GNDA.n2007 3.4105
R17120 GNDA.n2042 GNDA.n2007 3.4105
R17121 GNDA.n2392 GNDA.n2007 3.4105
R17122 GNDA.n2041 GNDA.n2007 3.4105
R17123 GNDA.n2394 GNDA.n2007 3.4105
R17124 GNDA.n2040 GNDA.n2007 3.4105
R17125 GNDA.n2396 GNDA.n2007 3.4105
R17126 GNDA.n2039 GNDA.n2007 3.4105
R17127 GNDA.n2398 GNDA.n2007 3.4105
R17128 GNDA.n2038 GNDA.n2007 3.4105
R17129 GNDA.n2400 GNDA.n2007 3.4105
R17130 GNDA.n2037 GNDA.n2007 3.4105
R17131 GNDA.n2402 GNDA.n2007 3.4105
R17132 GNDA.n2036 GNDA.n2007 3.4105
R17133 GNDA.n2404 GNDA.n2007 3.4105
R17134 GNDA.n2035 GNDA.n2007 3.4105
R17135 GNDA.n2406 GNDA.n2007 3.4105
R17136 GNDA.n2034 GNDA.n2007 3.4105
R17137 GNDA.n2408 GNDA.n2007 3.4105
R17138 GNDA.n2409 GNDA.n2007 3.4105
R17139 GNDA.n2429 GNDA.n2007 3.4105
R17140 GNDA.n2431 GNDA.n1994 3.4105
R17141 GNDA.n2048 GNDA.n1994 3.4105
R17142 GNDA.n2380 GNDA.n1994 3.4105
R17143 GNDA.n2047 GNDA.n1994 3.4105
R17144 GNDA.n2382 GNDA.n1994 3.4105
R17145 GNDA.n2046 GNDA.n1994 3.4105
R17146 GNDA.n2384 GNDA.n1994 3.4105
R17147 GNDA.n2045 GNDA.n1994 3.4105
R17148 GNDA.n2386 GNDA.n1994 3.4105
R17149 GNDA.n2044 GNDA.n1994 3.4105
R17150 GNDA.n2388 GNDA.n1994 3.4105
R17151 GNDA.n2043 GNDA.n1994 3.4105
R17152 GNDA.n2390 GNDA.n1994 3.4105
R17153 GNDA.n2042 GNDA.n1994 3.4105
R17154 GNDA.n2392 GNDA.n1994 3.4105
R17155 GNDA.n2041 GNDA.n1994 3.4105
R17156 GNDA.n2394 GNDA.n1994 3.4105
R17157 GNDA.n2040 GNDA.n1994 3.4105
R17158 GNDA.n2396 GNDA.n1994 3.4105
R17159 GNDA.n2039 GNDA.n1994 3.4105
R17160 GNDA.n2398 GNDA.n1994 3.4105
R17161 GNDA.n2038 GNDA.n1994 3.4105
R17162 GNDA.n2400 GNDA.n1994 3.4105
R17163 GNDA.n2037 GNDA.n1994 3.4105
R17164 GNDA.n2402 GNDA.n1994 3.4105
R17165 GNDA.n2036 GNDA.n1994 3.4105
R17166 GNDA.n2404 GNDA.n1994 3.4105
R17167 GNDA.n2035 GNDA.n1994 3.4105
R17168 GNDA.n2406 GNDA.n1994 3.4105
R17169 GNDA.n2034 GNDA.n1994 3.4105
R17170 GNDA.n2408 GNDA.n1994 3.4105
R17171 GNDA.n2409 GNDA.n1994 3.4105
R17172 GNDA.n2429 GNDA.n1994 3.4105
R17173 GNDA.n2431 GNDA.n2008 3.4105
R17174 GNDA.n2048 GNDA.n2008 3.4105
R17175 GNDA.n2380 GNDA.n2008 3.4105
R17176 GNDA.n2047 GNDA.n2008 3.4105
R17177 GNDA.n2382 GNDA.n2008 3.4105
R17178 GNDA.n2046 GNDA.n2008 3.4105
R17179 GNDA.n2384 GNDA.n2008 3.4105
R17180 GNDA.n2045 GNDA.n2008 3.4105
R17181 GNDA.n2386 GNDA.n2008 3.4105
R17182 GNDA.n2044 GNDA.n2008 3.4105
R17183 GNDA.n2388 GNDA.n2008 3.4105
R17184 GNDA.n2043 GNDA.n2008 3.4105
R17185 GNDA.n2390 GNDA.n2008 3.4105
R17186 GNDA.n2042 GNDA.n2008 3.4105
R17187 GNDA.n2392 GNDA.n2008 3.4105
R17188 GNDA.n2041 GNDA.n2008 3.4105
R17189 GNDA.n2394 GNDA.n2008 3.4105
R17190 GNDA.n2040 GNDA.n2008 3.4105
R17191 GNDA.n2396 GNDA.n2008 3.4105
R17192 GNDA.n2039 GNDA.n2008 3.4105
R17193 GNDA.n2398 GNDA.n2008 3.4105
R17194 GNDA.n2038 GNDA.n2008 3.4105
R17195 GNDA.n2400 GNDA.n2008 3.4105
R17196 GNDA.n2037 GNDA.n2008 3.4105
R17197 GNDA.n2402 GNDA.n2008 3.4105
R17198 GNDA.n2036 GNDA.n2008 3.4105
R17199 GNDA.n2404 GNDA.n2008 3.4105
R17200 GNDA.n2035 GNDA.n2008 3.4105
R17201 GNDA.n2406 GNDA.n2008 3.4105
R17202 GNDA.n2034 GNDA.n2008 3.4105
R17203 GNDA.n2408 GNDA.n2008 3.4105
R17204 GNDA.n2409 GNDA.n2008 3.4105
R17205 GNDA.n2429 GNDA.n2008 3.4105
R17206 GNDA.n2431 GNDA.n1993 3.4105
R17207 GNDA.n2048 GNDA.n1993 3.4105
R17208 GNDA.n2380 GNDA.n1993 3.4105
R17209 GNDA.n2047 GNDA.n1993 3.4105
R17210 GNDA.n2382 GNDA.n1993 3.4105
R17211 GNDA.n2046 GNDA.n1993 3.4105
R17212 GNDA.n2384 GNDA.n1993 3.4105
R17213 GNDA.n2045 GNDA.n1993 3.4105
R17214 GNDA.n2386 GNDA.n1993 3.4105
R17215 GNDA.n2044 GNDA.n1993 3.4105
R17216 GNDA.n2388 GNDA.n1993 3.4105
R17217 GNDA.n2043 GNDA.n1993 3.4105
R17218 GNDA.n2390 GNDA.n1993 3.4105
R17219 GNDA.n2042 GNDA.n1993 3.4105
R17220 GNDA.n2392 GNDA.n1993 3.4105
R17221 GNDA.n2041 GNDA.n1993 3.4105
R17222 GNDA.n2394 GNDA.n1993 3.4105
R17223 GNDA.n2040 GNDA.n1993 3.4105
R17224 GNDA.n2396 GNDA.n1993 3.4105
R17225 GNDA.n2039 GNDA.n1993 3.4105
R17226 GNDA.n2398 GNDA.n1993 3.4105
R17227 GNDA.n2038 GNDA.n1993 3.4105
R17228 GNDA.n2400 GNDA.n1993 3.4105
R17229 GNDA.n2037 GNDA.n1993 3.4105
R17230 GNDA.n2402 GNDA.n1993 3.4105
R17231 GNDA.n2036 GNDA.n1993 3.4105
R17232 GNDA.n2404 GNDA.n1993 3.4105
R17233 GNDA.n2035 GNDA.n1993 3.4105
R17234 GNDA.n2406 GNDA.n1993 3.4105
R17235 GNDA.n2034 GNDA.n1993 3.4105
R17236 GNDA.n2408 GNDA.n1993 3.4105
R17237 GNDA.n2409 GNDA.n1993 3.4105
R17238 GNDA.n2429 GNDA.n1993 3.4105
R17239 GNDA.n2431 GNDA.n2009 3.4105
R17240 GNDA.n2048 GNDA.n2009 3.4105
R17241 GNDA.n2380 GNDA.n2009 3.4105
R17242 GNDA.n2047 GNDA.n2009 3.4105
R17243 GNDA.n2382 GNDA.n2009 3.4105
R17244 GNDA.n2046 GNDA.n2009 3.4105
R17245 GNDA.n2384 GNDA.n2009 3.4105
R17246 GNDA.n2045 GNDA.n2009 3.4105
R17247 GNDA.n2386 GNDA.n2009 3.4105
R17248 GNDA.n2044 GNDA.n2009 3.4105
R17249 GNDA.n2388 GNDA.n2009 3.4105
R17250 GNDA.n2043 GNDA.n2009 3.4105
R17251 GNDA.n2390 GNDA.n2009 3.4105
R17252 GNDA.n2042 GNDA.n2009 3.4105
R17253 GNDA.n2392 GNDA.n2009 3.4105
R17254 GNDA.n2041 GNDA.n2009 3.4105
R17255 GNDA.n2394 GNDA.n2009 3.4105
R17256 GNDA.n2040 GNDA.n2009 3.4105
R17257 GNDA.n2396 GNDA.n2009 3.4105
R17258 GNDA.n2039 GNDA.n2009 3.4105
R17259 GNDA.n2398 GNDA.n2009 3.4105
R17260 GNDA.n2038 GNDA.n2009 3.4105
R17261 GNDA.n2400 GNDA.n2009 3.4105
R17262 GNDA.n2037 GNDA.n2009 3.4105
R17263 GNDA.n2402 GNDA.n2009 3.4105
R17264 GNDA.n2036 GNDA.n2009 3.4105
R17265 GNDA.n2404 GNDA.n2009 3.4105
R17266 GNDA.n2035 GNDA.n2009 3.4105
R17267 GNDA.n2406 GNDA.n2009 3.4105
R17268 GNDA.n2034 GNDA.n2009 3.4105
R17269 GNDA.n2408 GNDA.n2009 3.4105
R17270 GNDA.n2409 GNDA.n2009 3.4105
R17271 GNDA.n2429 GNDA.n2009 3.4105
R17272 GNDA.n2431 GNDA.n1992 3.4105
R17273 GNDA.n2048 GNDA.n1992 3.4105
R17274 GNDA.n2380 GNDA.n1992 3.4105
R17275 GNDA.n2047 GNDA.n1992 3.4105
R17276 GNDA.n2382 GNDA.n1992 3.4105
R17277 GNDA.n2046 GNDA.n1992 3.4105
R17278 GNDA.n2384 GNDA.n1992 3.4105
R17279 GNDA.n2045 GNDA.n1992 3.4105
R17280 GNDA.n2386 GNDA.n1992 3.4105
R17281 GNDA.n2044 GNDA.n1992 3.4105
R17282 GNDA.n2388 GNDA.n1992 3.4105
R17283 GNDA.n2043 GNDA.n1992 3.4105
R17284 GNDA.n2390 GNDA.n1992 3.4105
R17285 GNDA.n2042 GNDA.n1992 3.4105
R17286 GNDA.n2392 GNDA.n1992 3.4105
R17287 GNDA.n2041 GNDA.n1992 3.4105
R17288 GNDA.n2394 GNDA.n1992 3.4105
R17289 GNDA.n2040 GNDA.n1992 3.4105
R17290 GNDA.n2396 GNDA.n1992 3.4105
R17291 GNDA.n2039 GNDA.n1992 3.4105
R17292 GNDA.n2398 GNDA.n1992 3.4105
R17293 GNDA.n2038 GNDA.n1992 3.4105
R17294 GNDA.n2400 GNDA.n1992 3.4105
R17295 GNDA.n2037 GNDA.n1992 3.4105
R17296 GNDA.n2402 GNDA.n1992 3.4105
R17297 GNDA.n2036 GNDA.n1992 3.4105
R17298 GNDA.n2404 GNDA.n1992 3.4105
R17299 GNDA.n2035 GNDA.n1992 3.4105
R17300 GNDA.n2406 GNDA.n1992 3.4105
R17301 GNDA.n2034 GNDA.n1992 3.4105
R17302 GNDA.n2408 GNDA.n1992 3.4105
R17303 GNDA.n2409 GNDA.n1992 3.4105
R17304 GNDA.n2429 GNDA.n1992 3.4105
R17305 GNDA.n2431 GNDA.n2010 3.4105
R17306 GNDA.n2048 GNDA.n2010 3.4105
R17307 GNDA.n2380 GNDA.n2010 3.4105
R17308 GNDA.n2047 GNDA.n2010 3.4105
R17309 GNDA.n2382 GNDA.n2010 3.4105
R17310 GNDA.n2046 GNDA.n2010 3.4105
R17311 GNDA.n2384 GNDA.n2010 3.4105
R17312 GNDA.n2045 GNDA.n2010 3.4105
R17313 GNDA.n2386 GNDA.n2010 3.4105
R17314 GNDA.n2044 GNDA.n2010 3.4105
R17315 GNDA.n2388 GNDA.n2010 3.4105
R17316 GNDA.n2043 GNDA.n2010 3.4105
R17317 GNDA.n2390 GNDA.n2010 3.4105
R17318 GNDA.n2042 GNDA.n2010 3.4105
R17319 GNDA.n2392 GNDA.n2010 3.4105
R17320 GNDA.n2041 GNDA.n2010 3.4105
R17321 GNDA.n2394 GNDA.n2010 3.4105
R17322 GNDA.n2040 GNDA.n2010 3.4105
R17323 GNDA.n2396 GNDA.n2010 3.4105
R17324 GNDA.n2039 GNDA.n2010 3.4105
R17325 GNDA.n2398 GNDA.n2010 3.4105
R17326 GNDA.n2038 GNDA.n2010 3.4105
R17327 GNDA.n2400 GNDA.n2010 3.4105
R17328 GNDA.n2037 GNDA.n2010 3.4105
R17329 GNDA.n2402 GNDA.n2010 3.4105
R17330 GNDA.n2036 GNDA.n2010 3.4105
R17331 GNDA.n2404 GNDA.n2010 3.4105
R17332 GNDA.n2035 GNDA.n2010 3.4105
R17333 GNDA.n2406 GNDA.n2010 3.4105
R17334 GNDA.n2034 GNDA.n2010 3.4105
R17335 GNDA.n2408 GNDA.n2010 3.4105
R17336 GNDA.n2409 GNDA.n2010 3.4105
R17337 GNDA.n2429 GNDA.n2010 3.4105
R17338 GNDA.n2431 GNDA.n1991 3.4105
R17339 GNDA.n2048 GNDA.n1991 3.4105
R17340 GNDA.n2380 GNDA.n1991 3.4105
R17341 GNDA.n2047 GNDA.n1991 3.4105
R17342 GNDA.n2382 GNDA.n1991 3.4105
R17343 GNDA.n2046 GNDA.n1991 3.4105
R17344 GNDA.n2384 GNDA.n1991 3.4105
R17345 GNDA.n2045 GNDA.n1991 3.4105
R17346 GNDA.n2386 GNDA.n1991 3.4105
R17347 GNDA.n2044 GNDA.n1991 3.4105
R17348 GNDA.n2388 GNDA.n1991 3.4105
R17349 GNDA.n2043 GNDA.n1991 3.4105
R17350 GNDA.n2390 GNDA.n1991 3.4105
R17351 GNDA.n2042 GNDA.n1991 3.4105
R17352 GNDA.n2392 GNDA.n1991 3.4105
R17353 GNDA.n2041 GNDA.n1991 3.4105
R17354 GNDA.n2394 GNDA.n1991 3.4105
R17355 GNDA.n2040 GNDA.n1991 3.4105
R17356 GNDA.n2396 GNDA.n1991 3.4105
R17357 GNDA.n2039 GNDA.n1991 3.4105
R17358 GNDA.n2398 GNDA.n1991 3.4105
R17359 GNDA.n2038 GNDA.n1991 3.4105
R17360 GNDA.n2400 GNDA.n1991 3.4105
R17361 GNDA.n2037 GNDA.n1991 3.4105
R17362 GNDA.n2402 GNDA.n1991 3.4105
R17363 GNDA.n2036 GNDA.n1991 3.4105
R17364 GNDA.n2404 GNDA.n1991 3.4105
R17365 GNDA.n2035 GNDA.n1991 3.4105
R17366 GNDA.n2406 GNDA.n1991 3.4105
R17367 GNDA.n2034 GNDA.n1991 3.4105
R17368 GNDA.n2408 GNDA.n1991 3.4105
R17369 GNDA.n2409 GNDA.n1991 3.4105
R17370 GNDA.n2429 GNDA.n1991 3.4105
R17371 GNDA.n2431 GNDA.n2011 3.4105
R17372 GNDA.n2048 GNDA.n2011 3.4105
R17373 GNDA.n2380 GNDA.n2011 3.4105
R17374 GNDA.n2047 GNDA.n2011 3.4105
R17375 GNDA.n2382 GNDA.n2011 3.4105
R17376 GNDA.n2046 GNDA.n2011 3.4105
R17377 GNDA.n2384 GNDA.n2011 3.4105
R17378 GNDA.n2045 GNDA.n2011 3.4105
R17379 GNDA.n2386 GNDA.n2011 3.4105
R17380 GNDA.n2044 GNDA.n2011 3.4105
R17381 GNDA.n2388 GNDA.n2011 3.4105
R17382 GNDA.n2043 GNDA.n2011 3.4105
R17383 GNDA.n2390 GNDA.n2011 3.4105
R17384 GNDA.n2042 GNDA.n2011 3.4105
R17385 GNDA.n2392 GNDA.n2011 3.4105
R17386 GNDA.n2041 GNDA.n2011 3.4105
R17387 GNDA.n2394 GNDA.n2011 3.4105
R17388 GNDA.n2040 GNDA.n2011 3.4105
R17389 GNDA.n2396 GNDA.n2011 3.4105
R17390 GNDA.n2039 GNDA.n2011 3.4105
R17391 GNDA.n2398 GNDA.n2011 3.4105
R17392 GNDA.n2038 GNDA.n2011 3.4105
R17393 GNDA.n2400 GNDA.n2011 3.4105
R17394 GNDA.n2037 GNDA.n2011 3.4105
R17395 GNDA.n2402 GNDA.n2011 3.4105
R17396 GNDA.n2036 GNDA.n2011 3.4105
R17397 GNDA.n2404 GNDA.n2011 3.4105
R17398 GNDA.n2035 GNDA.n2011 3.4105
R17399 GNDA.n2406 GNDA.n2011 3.4105
R17400 GNDA.n2034 GNDA.n2011 3.4105
R17401 GNDA.n2408 GNDA.n2011 3.4105
R17402 GNDA.n2409 GNDA.n2011 3.4105
R17403 GNDA.n2429 GNDA.n2011 3.4105
R17404 GNDA.n2431 GNDA.n1990 3.4105
R17405 GNDA.n2048 GNDA.n1990 3.4105
R17406 GNDA.n2380 GNDA.n1990 3.4105
R17407 GNDA.n2047 GNDA.n1990 3.4105
R17408 GNDA.n2382 GNDA.n1990 3.4105
R17409 GNDA.n2046 GNDA.n1990 3.4105
R17410 GNDA.n2384 GNDA.n1990 3.4105
R17411 GNDA.n2045 GNDA.n1990 3.4105
R17412 GNDA.n2386 GNDA.n1990 3.4105
R17413 GNDA.n2044 GNDA.n1990 3.4105
R17414 GNDA.n2388 GNDA.n1990 3.4105
R17415 GNDA.n2043 GNDA.n1990 3.4105
R17416 GNDA.n2390 GNDA.n1990 3.4105
R17417 GNDA.n2042 GNDA.n1990 3.4105
R17418 GNDA.n2392 GNDA.n1990 3.4105
R17419 GNDA.n2041 GNDA.n1990 3.4105
R17420 GNDA.n2394 GNDA.n1990 3.4105
R17421 GNDA.n2040 GNDA.n1990 3.4105
R17422 GNDA.n2396 GNDA.n1990 3.4105
R17423 GNDA.n2039 GNDA.n1990 3.4105
R17424 GNDA.n2398 GNDA.n1990 3.4105
R17425 GNDA.n2038 GNDA.n1990 3.4105
R17426 GNDA.n2400 GNDA.n1990 3.4105
R17427 GNDA.n2037 GNDA.n1990 3.4105
R17428 GNDA.n2402 GNDA.n1990 3.4105
R17429 GNDA.n2036 GNDA.n1990 3.4105
R17430 GNDA.n2404 GNDA.n1990 3.4105
R17431 GNDA.n2035 GNDA.n1990 3.4105
R17432 GNDA.n2406 GNDA.n1990 3.4105
R17433 GNDA.n2034 GNDA.n1990 3.4105
R17434 GNDA.n2408 GNDA.n1990 3.4105
R17435 GNDA.n2409 GNDA.n1990 3.4105
R17436 GNDA.n2429 GNDA.n1990 3.4105
R17437 GNDA.n2431 GNDA.n2012 3.4105
R17438 GNDA.n2048 GNDA.n2012 3.4105
R17439 GNDA.n2380 GNDA.n2012 3.4105
R17440 GNDA.n2047 GNDA.n2012 3.4105
R17441 GNDA.n2382 GNDA.n2012 3.4105
R17442 GNDA.n2046 GNDA.n2012 3.4105
R17443 GNDA.n2384 GNDA.n2012 3.4105
R17444 GNDA.n2045 GNDA.n2012 3.4105
R17445 GNDA.n2386 GNDA.n2012 3.4105
R17446 GNDA.n2044 GNDA.n2012 3.4105
R17447 GNDA.n2388 GNDA.n2012 3.4105
R17448 GNDA.n2043 GNDA.n2012 3.4105
R17449 GNDA.n2390 GNDA.n2012 3.4105
R17450 GNDA.n2042 GNDA.n2012 3.4105
R17451 GNDA.n2392 GNDA.n2012 3.4105
R17452 GNDA.n2041 GNDA.n2012 3.4105
R17453 GNDA.n2394 GNDA.n2012 3.4105
R17454 GNDA.n2040 GNDA.n2012 3.4105
R17455 GNDA.n2396 GNDA.n2012 3.4105
R17456 GNDA.n2039 GNDA.n2012 3.4105
R17457 GNDA.n2398 GNDA.n2012 3.4105
R17458 GNDA.n2038 GNDA.n2012 3.4105
R17459 GNDA.n2400 GNDA.n2012 3.4105
R17460 GNDA.n2037 GNDA.n2012 3.4105
R17461 GNDA.n2402 GNDA.n2012 3.4105
R17462 GNDA.n2036 GNDA.n2012 3.4105
R17463 GNDA.n2404 GNDA.n2012 3.4105
R17464 GNDA.n2035 GNDA.n2012 3.4105
R17465 GNDA.n2406 GNDA.n2012 3.4105
R17466 GNDA.n2034 GNDA.n2012 3.4105
R17467 GNDA.n2408 GNDA.n2012 3.4105
R17468 GNDA.n2409 GNDA.n2012 3.4105
R17469 GNDA.n2429 GNDA.n2012 3.4105
R17470 GNDA.n2431 GNDA.n1989 3.4105
R17471 GNDA.n2048 GNDA.n1989 3.4105
R17472 GNDA.n2380 GNDA.n1989 3.4105
R17473 GNDA.n2047 GNDA.n1989 3.4105
R17474 GNDA.n2382 GNDA.n1989 3.4105
R17475 GNDA.n2046 GNDA.n1989 3.4105
R17476 GNDA.n2384 GNDA.n1989 3.4105
R17477 GNDA.n2045 GNDA.n1989 3.4105
R17478 GNDA.n2386 GNDA.n1989 3.4105
R17479 GNDA.n2044 GNDA.n1989 3.4105
R17480 GNDA.n2388 GNDA.n1989 3.4105
R17481 GNDA.n2043 GNDA.n1989 3.4105
R17482 GNDA.n2390 GNDA.n1989 3.4105
R17483 GNDA.n2042 GNDA.n1989 3.4105
R17484 GNDA.n2392 GNDA.n1989 3.4105
R17485 GNDA.n2041 GNDA.n1989 3.4105
R17486 GNDA.n2394 GNDA.n1989 3.4105
R17487 GNDA.n2040 GNDA.n1989 3.4105
R17488 GNDA.n2396 GNDA.n1989 3.4105
R17489 GNDA.n2039 GNDA.n1989 3.4105
R17490 GNDA.n2398 GNDA.n1989 3.4105
R17491 GNDA.n2038 GNDA.n1989 3.4105
R17492 GNDA.n2400 GNDA.n1989 3.4105
R17493 GNDA.n2037 GNDA.n1989 3.4105
R17494 GNDA.n2402 GNDA.n1989 3.4105
R17495 GNDA.n2036 GNDA.n1989 3.4105
R17496 GNDA.n2404 GNDA.n1989 3.4105
R17497 GNDA.n2035 GNDA.n1989 3.4105
R17498 GNDA.n2406 GNDA.n1989 3.4105
R17499 GNDA.n2034 GNDA.n1989 3.4105
R17500 GNDA.n2408 GNDA.n1989 3.4105
R17501 GNDA.n2409 GNDA.n1989 3.4105
R17502 GNDA.n2429 GNDA.n1989 3.4105
R17503 GNDA.n2431 GNDA.n2013 3.4105
R17504 GNDA.n2048 GNDA.n2013 3.4105
R17505 GNDA.n2380 GNDA.n2013 3.4105
R17506 GNDA.n2047 GNDA.n2013 3.4105
R17507 GNDA.n2382 GNDA.n2013 3.4105
R17508 GNDA.n2046 GNDA.n2013 3.4105
R17509 GNDA.n2384 GNDA.n2013 3.4105
R17510 GNDA.n2045 GNDA.n2013 3.4105
R17511 GNDA.n2386 GNDA.n2013 3.4105
R17512 GNDA.n2044 GNDA.n2013 3.4105
R17513 GNDA.n2388 GNDA.n2013 3.4105
R17514 GNDA.n2043 GNDA.n2013 3.4105
R17515 GNDA.n2390 GNDA.n2013 3.4105
R17516 GNDA.n2042 GNDA.n2013 3.4105
R17517 GNDA.n2392 GNDA.n2013 3.4105
R17518 GNDA.n2041 GNDA.n2013 3.4105
R17519 GNDA.n2394 GNDA.n2013 3.4105
R17520 GNDA.n2040 GNDA.n2013 3.4105
R17521 GNDA.n2396 GNDA.n2013 3.4105
R17522 GNDA.n2039 GNDA.n2013 3.4105
R17523 GNDA.n2398 GNDA.n2013 3.4105
R17524 GNDA.n2038 GNDA.n2013 3.4105
R17525 GNDA.n2400 GNDA.n2013 3.4105
R17526 GNDA.n2037 GNDA.n2013 3.4105
R17527 GNDA.n2402 GNDA.n2013 3.4105
R17528 GNDA.n2036 GNDA.n2013 3.4105
R17529 GNDA.n2404 GNDA.n2013 3.4105
R17530 GNDA.n2035 GNDA.n2013 3.4105
R17531 GNDA.n2406 GNDA.n2013 3.4105
R17532 GNDA.n2034 GNDA.n2013 3.4105
R17533 GNDA.n2408 GNDA.n2013 3.4105
R17534 GNDA.n2409 GNDA.n2013 3.4105
R17535 GNDA.n2429 GNDA.n2013 3.4105
R17536 GNDA.n2431 GNDA.n1988 3.4105
R17537 GNDA.n2048 GNDA.n1988 3.4105
R17538 GNDA.n2380 GNDA.n1988 3.4105
R17539 GNDA.n2047 GNDA.n1988 3.4105
R17540 GNDA.n2382 GNDA.n1988 3.4105
R17541 GNDA.n2046 GNDA.n1988 3.4105
R17542 GNDA.n2384 GNDA.n1988 3.4105
R17543 GNDA.n2045 GNDA.n1988 3.4105
R17544 GNDA.n2386 GNDA.n1988 3.4105
R17545 GNDA.n2044 GNDA.n1988 3.4105
R17546 GNDA.n2388 GNDA.n1988 3.4105
R17547 GNDA.n2043 GNDA.n1988 3.4105
R17548 GNDA.n2390 GNDA.n1988 3.4105
R17549 GNDA.n2042 GNDA.n1988 3.4105
R17550 GNDA.n2392 GNDA.n1988 3.4105
R17551 GNDA.n2041 GNDA.n1988 3.4105
R17552 GNDA.n2394 GNDA.n1988 3.4105
R17553 GNDA.n2040 GNDA.n1988 3.4105
R17554 GNDA.n2396 GNDA.n1988 3.4105
R17555 GNDA.n2039 GNDA.n1988 3.4105
R17556 GNDA.n2398 GNDA.n1988 3.4105
R17557 GNDA.n2038 GNDA.n1988 3.4105
R17558 GNDA.n2400 GNDA.n1988 3.4105
R17559 GNDA.n2037 GNDA.n1988 3.4105
R17560 GNDA.n2402 GNDA.n1988 3.4105
R17561 GNDA.n2036 GNDA.n1988 3.4105
R17562 GNDA.n2404 GNDA.n1988 3.4105
R17563 GNDA.n2035 GNDA.n1988 3.4105
R17564 GNDA.n2406 GNDA.n1988 3.4105
R17565 GNDA.n2034 GNDA.n1988 3.4105
R17566 GNDA.n2408 GNDA.n1988 3.4105
R17567 GNDA.n2409 GNDA.n1988 3.4105
R17568 GNDA.n2429 GNDA.n1988 3.4105
R17569 GNDA.n2431 GNDA.n2014 3.4105
R17570 GNDA.n2048 GNDA.n2014 3.4105
R17571 GNDA.n2380 GNDA.n2014 3.4105
R17572 GNDA.n2047 GNDA.n2014 3.4105
R17573 GNDA.n2382 GNDA.n2014 3.4105
R17574 GNDA.n2046 GNDA.n2014 3.4105
R17575 GNDA.n2384 GNDA.n2014 3.4105
R17576 GNDA.n2045 GNDA.n2014 3.4105
R17577 GNDA.n2386 GNDA.n2014 3.4105
R17578 GNDA.n2044 GNDA.n2014 3.4105
R17579 GNDA.n2388 GNDA.n2014 3.4105
R17580 GNDA.n2043 GNDA.n2014 3.4105
R17581 GNDA.n2390 GNDA.n2014 3.4105
R17582 GNDA.n2042 GNDA.n2014 3.4105
R17583 GNDA.n2392 GNDA.n2014 3.4105
R17584 GNDA.n2041 GNDA.n2014 3.4105
R17585 GNDA.n2394 GNDA.n2014 3.4105
R17586 GNDA.n2040 GNDA.n2014 3.4105
R17587 GNDA.n2396 GNDA.n2014 3.4105
R17588 GNDA.n2039 GNDA.n2014 3.4105
R17589 GNDA.n2398 GNDA.n2014 3.4105
R17590 GNDA.n2038 GNDA.n2014 3.4105
R17591 GNDA.n2400 GNDA.n2014 3.4105
R17592 GNDA.n2037 GNDA.n2014 3.4105
R17593 GNDA.n2402 GNDA.n2014 3.4105
R17594 GNDA.n2036 GNDA.n2014 3.4105
R17595 GNDA.n2404 GNDA.n2014 3.4105
R17596 GNDA.n2035 GNDA.n2014 3.4105
R17597 GNDA.n2406 GNDA.n2014 3.4105
R17598 GNDA.n2034 GNDA.n2014 3.4105
R17599 GNDA.n2408 GNDA.n2014 3.4105
R17600 GNDA.n2409 GNDA.n2014 3.4105
R17601 GNDA.n2429 GNDA.n2014 3.4105
R17602 GNDA.n2431 GNDA.n1987 3.4105
R17603 GNDA.n2048 GNDA.n1987 3.4105
R17604 GNDA.n2380 GNDA.n1987 3.4105
R17605 GNDA.n2047 GNDA.n1987 3.4105
R17606 GNDA.n2382 GNDA.n1987 3.4105
R17607 GNDA.n2046 GNDA.n1987 3.4105
R17608 GNDA.n2384 GNDA.n1987 3.4105
R17609 GNDA.n2045 GNDA.n1987 3.4105
R17610 GNDA.n2386 GNDA.n1987 3.4105
R17611 GNDA.n2044 GNDA.n1987 3.4105
R17612 GNDA.n2388 GNDA.n1987 3.4105
R17613 GNDA.n2043 GNDA.n1987 3.4105
R17614 GNDA.n2390 GNDA.n1987 3.4105
R17615 GNDA.n2042 GNDA.n1987 3.4105
R17616 GNDA.n2392 GNDA.n1987 3.4105
R17617 GNDA.n2041 GNDA.n1987 3.4105
R17618 GNDA.n2394 GNDA.n1987 3.4105
R17619 GNDA.n2040 GNDA.n1987 3.4105
R17620 GNDA.n2396 GNDA.n1987 3.4105
R17621 GNDA.n2039 GNDA.n1987 3.4105
R17622 GNDA.n2398 GNDA.n1987 3.4105
R17623 GNDA.n2038 GNDA.n1987 3.4105
R17624 GNDA.n2400 GNDA.n1987 3.4105
R17625 GNDA.n2037 GNDA.n1987 3.4105
R17626 GNDA.n2402 GNDA.n1987 3.4105
R17627 GNDA.n2036 GNDA.n1987 3.4105
R17628 GNDA.n2404 GNDA.n1987 3.4105
R17629 GNDA.n2035 GNDA.n1987 3.4105
R17630 GNDA.n2406 GNDA.n1987 3.4105
R17631 GNDA.n2034 GNDA.n1987 3.4105
R17632 GNDA.n2408 GNDA.n1987 3.4105
R17633 GNDA.n2409 GNDA.n1987 3.4105
R17634 GNDA.n2429 GNDA.n1987 3.4105
R17635 GNDA.n2431 GNDA.n2015 3.4105
R17636 GNDA.n2048 GNDA.n2015 3.4105
R17637 GNDA.n2380 GNDA.n2015 3.4105
R17638 GNDA.n2047 GNDA.n2015 3.4105
R17639 GNDA.n2382 GNDA.n2015 3.4105
R17640 GNDA.n2046 GNDA.n2015 3.4105
R17641 GNDA.n2384 GNDA.n2015 3.4105
R17642 GNDA.n2045 GNDA.n2015 3.4105
R17643 GNDA.n2386 GNDA.n2015 3.4105
R17644 GNDA.n2044 GNDA.n2015 3.4105
R17645 GNDA.n2388 GNDA.n2015 3.4105
R17646 GNDA.n2043 GNDA.n2015 3.4105
R17647 GNDA.n2390 GNDA.n2015 3.4105
R17648 GNDA.n2042 GNDA.n2015 3.4105
R17649 GNDA.n2392 GNDA.n2015 3.4105
R17650 GNDA.n2041 GNDA.n2015 3.4105
R17651 GNDA.n2394 GNDA.n2015 3.4105
R17652 GNDA.n2040 GNDA.n2015 3.4105
R17653 GNDA.n2396 GNDA.n2015 3.4105
R17654 GNDA.n2039 GNDA.n2015 3.4105
R17655 GNDA.n2398 GNDA.n2015 3.4105
R17656 GNDA.n2038 GNDA.n2015 3.4105
R17657 GNDA.n2400 GNDA.n2015 3.4105
R17658 GNDA.n2037 GNDA.n2015 3.4105
R17659 GNDA.n2402 GNDA.n2015 3.4105
R17660 GNDA.n2036 GNDA.n2015 3.4105
R17661 GNDA.n2404 GNDA.n2015 3.4105
R17662 GNDA.n2035 GNDA.n2015 3.4105
R17663 GNDA.n2406 GNDA.n2015 3.4105
R17664 GNDA.n2034 GNDA.n2015 3.4105
R17665 GNDA.n2408 GNDA.n2015 3.4105
R17666 GNDA.n2409 GNDA.n2015 3.4105
R17667 GNDA.n2429 GNDA.n2015 3.4105
R17668 GNDA.n2431 GNDA.n1986 3.4105
R17669 GNDA.n2048 GNDA.n1986 3.4105
R17670 GNDA.n2380 GNDA.n1986 3.4105
R17671 GNDA.n2047 GNDA.n1986 3.4105
R17672 GNDA.n2382 GNDA.n1986 3.4105
R17673 GNDA.n2046 GNDA.n1986 3.4105
R17674 GNDA.n2384 GNDA.n1986 3.4105
R17675 GNDA.n2045 GNDA.n1986 3.4105
R17676 GNDA.n2386 GNDA.n1986 3.4105
R17677 GNDA.n2044 GNDA.n1986 3.4105
R17678 GNDA.n2388 GNDA.n1986 3.4105
R17679 GNDA.n2043 GNDA.n1986 3.4105
R17680 GNDA.n2390 GNDA.n1986 3.4105
R17681 GNDA.n2042 GNDA.n1986 3.4105
R17682 GNDA.n2392 GNDA.n1986 3.4105
R17683 GNDA.n2041 GNDA.n1986 3.4105
R17684 GNDA.n2394 GNDA.n1986 3.4105
R17685 GNDA.n2040 GNDA.n1986 3.4105
R17686 GNDA.n2396 GNDA.n1986 3.4105
R17687 GNDA.n2039 GNDA.n1986 3.4105
R17688 GNDA.n2398 GNDA.n1986 3.4105
R17689 GNDA.n2038 GNDA.n1986 3.4105
R17690 GNDA.n2400 GNDA.n1986 3.4105
R17691 GNDA.n2037 GNDA.n1986 3.4105
R17692 GNDA.n2402 GNDA.n1986 3.4105
R17693 GNDA.n2036 GNDA.n1986 3.4105
R17694 GNDA.n2404 GNDA.n1986 3.4105
R17695 GNDA.n2035 GNDA.n1986 3.4105
R17696 GNDA.n2406 GNDA.n1986 3.4105
R17697 GNDA.n2034 GNDA.n1986 3.4105
R17698 GNDA.n2408 GNDA.n1986 3.4105
R17699 GNDA.n2409 GNDA.n1986 3.4105
R17700 GNDA.n2429 GNDA.n1986 3.4105
R17701 GNDA.n2431 GNDA.n2016 3.4105
R17702 GNDA.n2048 GNDA.n2016 3.4105
R17703 GNDA.n2380 GNDA.n2016 3.4105
R17704 GNDA.n2047 GNDA.n2016 3.4105
R17705 GNDA.n2382 GNDA.n2016 3.4105
R17706 GNDA.n2046 GNDA.n2016 3.4105
R17707 GNDA.n2384 GNDA.n2016 3.4105
R17708 GNDA.n2045 GNDA.n2016 3.4105
R17709 GNDA.n2386 GNDA.n2016 3.4105
R17710 GNDA.n2044 GNDA.n2016 3.4105
R17711 GNDA.n2388 GNDA.n2016 3.4105
R17712 GNDA.n2043 GNDA.n2016 3.4105
R17713 GNDA.n2390 GNDA.n2016 3.4105
R17714 GNDA.n2042 GNDA.n2016 3.4105
R17715 GNDA.n2392 GNDA.n2016 3.4105
R17716 GNDA.n2041 GNDA.n2016 3.4105
R17717 GNDA.n2394 GNDA.n2016 3.4105
R17718 GNDA.n2040 GNDA.n2016 3.4105
R17719 GNDA.n2396 GNDA.n2016 3.4105
R17720 GNDA.n2039 GNDA.n2016 3.4105
R17721 GNDA.n2398 GNDA.n2016 3.4105
R17722 GNDA.n2038 GNDA.n2016 3.4105
R17723 GNDA.n2400 GNDA.n2016 3.4105
R17724 GNDA.n2037 GNDA.n2016 3.4105
R17725 GNDA.n2402 GNDA.n2016 3.4105
R17726 GNDA.n2036 GNDA.n2016 3.4105
R17727 GNDA.n2404 GNDA.n2016 3.4105
R17728 GNDA.n2035 GNDA.n2016 3.4105
R17729 GNDA.n2406 GNDA.n2016 3.4105
R17730 GNDA.n2034 GNDA.n2016 3.4105
R17731 GNDA.n2408 GNDA.n2016 3.4105
R17732 GNDA.n2409 GNDA.n2016 3.4105
R17733 GNDA.n2429 GNDA.n2016 3.4105
R17734 GNDA.n2431 GNDA.n1985 3.4105
R17735 GNDA.n2048 GNDA.n1985 3.4105
R17736 GNDA.n2380 GNDA.n1985 3.4105
R17737 GNDA.n2047 GNDA.n1985 3.4105
R17738 GNDA.n2382 GNDA.n1985 3.4105
R17739 GNDA.n2046 GNDA.n1985 3.4105
R17740 GNDA.n2384 GNDA.n1985 3.4105
R17741 GNDA.n2045 GNDA.n1985 3.4105
R17742 GNDA.n2386 GNDA.n1985 3.4105
R17743 GNDA.n2044 GNDA.n1985 3.4105
R17744 GNDA.n2388 GNDA.n1985 3.4105
R17745 GNDA.n2043 GNDA.n1985 3.4105
R17746 GNDA.n2390 GNDA.n1985 3.4105
R17747 GNDA.n2042 GNDA.n1985 3.4105
R17748 GNDA.n2392 GNDA.n1985 3.4105
R17749 GNDA.n2041 GNDA.n1985 3.4105
R17750 GNDA.n2394 GNDA.n1985 3.4105
R17751 GNDA.n2040 GNDA.n1985 3.4105
R17752 GNDA.n2396 GNDA.n1985 3.4105
R17753 GNDA.n2039 GNDA.n1985 3.4105
R17754 GNDA.n2398 GNDA.n1985 3.4105
R17755 GNDA.n2038 GNDA.n1985 3.4105
R17756 GNDA.n2400 GNDA.n1985 3.4105
R17757 GNDA.n2037 GNDA.n1985 3.4105
R17758 GNDA.n2402 GNDA.n1985 3.4105
R17759 GNDA.n2036 GNDA.n1985 3.4105
R17760 GNDA.n2404 GNDA.n1985 3.4105
R17761 GNDA.n2035 GNDA.n1985 3.4105
R17762 GNDA.n2406 GNDA.n1985 3.4105
R17763 GNDA.n2034 GNDA.n1985 3.4105
R17764 GNDA.n2408 GNDA.n1985 3.4105
R17765 GNDA.n2409 GNDA.n1985 3.4105
R17766 GNDA.n2429 GNDA.n1985 3.4105
R17767 GNDA.n2431 GNDA.n2430 3.4105
R17768 GNDA.n2430 GNDA.n2048 3.4105
R17769 GNDA.n2430 GNDA.n2380 3.4105
R17770 GNDA.n2430 GNDA.n2047 3.4105
R17771 GNDA.n2430 GNDA.n2382 3.4105
R17772 GNDA.n2430 GNDA.n2046 3.4105
R17773 GNDA.n2430 GNDA.n2384 3.4105
R17774 GNDA.n2430 GNDA.n2045 3.4105
R17775 GNDA.n2430 GNDA.n2386 3.4105
R17776 GNDA.n2430 GNDA.n2044 3.4105
R17777 GNDA.n2430 GNDA.n2388 3.4105
R17778 GNDA.n2430 GNDA.n2043 3.4105
R17779 GNDA.n2430 GNDA.n2390 3.4105
R17780 GNDA.n2430 GNDA.n2042 3.4105
R17781 GNDA.n2430 GNDA.n2392 3.4105
R17782 GNDA.n2430 GNDA.n2041 3.4105
R17783 GNDA.n2430 GNDA.n2394 3.4105
R17784 GNDA.n2430 GNDA.n2040 3.4105
R17785 GNDA.n2430 GNDA.n2396 3.4105
R17786 GNDA.n2430 GNDA.n2039 3.4105
R17787 GNDA.n2430 GNDA.n2398 3.4105
R17788 GNDA.n2430 GNDA.n2038 3.4105
R17789 GNDA.n2430 GNDA.n2400 3.4105
R17790 GNDA.n2430 GNDA.n2037 3.4105
R17791 GNDA.n2430 GNDA.n2402 3.4105
R17792 GNDA.n2430 GNDA.n2036 3.4105
R17793 GNDA.n2430 GNDA.n2404 3.4105
R17794 GNDA.n2430 GNDA.n2035 3.4105
R17795 GNDA.n2430 GNDA.n2406 3.4105
R17796 GNDA.n2430 GNDA.n2034 3.4105
R17797 GNDA.n2430 GNDA.n2408 3.4105
R17798 GNDA.n2430 GNDA.n2033 3.4105
R17799 GNDA.n2430 GNDA.n2409 3.4105
R17800 GNDA.n2430 GNDA.n2429 3.4105
R17801 GNDA.n3614 GNDA.n3613 3.39217
R17802 GNDA.n1452 GNDA.n1451 3.39217
R17803 GNDA.n584 GNDA.n583 3.39217
R17804 GNDA.n3335 GNDA.n588 3.39217
R17805 GNDA.n3581 GNDA.n585 3.13621
R17806 GNDA.n3582 GNDA.n3581 3.13621
R17807 GNDA.n3574 GNDA.n587 3.13621
R17808 GNDA.n3574 GNDA.n3573 3.13621
R17809 GNDA.n3227 GNDA.n1527 3.04346
R17810 GNDA.n2918 GNDA.n2917 3.00528
R17811 GNDA.n3278 GNDA.n3277 3.00528
R17812 GNDA.n3128 GNDA.t175 3.00528
R17813 GNDA.t281 GNDA.n1506 3.00528
R17814 GNDA.n3236 GNDA.n3235 2.86505
R17815 GNDA.n3237 GNDA.n3236 2.86505
R17816 GNDA.n3241 GNDA.n3239 2.86505
R17817 GNDA.n3244 GNDA.n3239 2.86505
R17818 GNDA.n3240 GNDA.n3237 2.86505
R17819 GNDA.n3244 GNDA.n3243 2.86505
R17820 GNDA.n3246 GNDA.n3235 2.86505
R17821 GNDA.n3241 GNDA.n3240 2.86505
R17822 GNDA.n2822 GNDA.n2821 2.86505
R17823 GNDA.n2821 GNDA.n2819 2.86505
R17824 GNDA.n2819 GNDA.n2818 2.86505
R17825 GNDA.n2823 GNDA.n2822 2.86505
R17826 GNDA.n3139 GNDA.n3138 2.6629
R17827 GNDA.n2740 GNDA.n2739 2.6629
R17828 GNDA.n2795 GNDA.n1824 2.6629
R17829 GNDA.n5049 GNDA.n5048 2.6629
R17830 GNDA.n1550 GNDA.n1549 2.6629
R17831 GNDA.n1677 GNDA.n1676 2.6629
R17832 GNDA.n4978 GNDA.n4977 2.6629
R17833 GNDA.n4891 GNDA.n160 2.6629
R17834 GNDA.n5257 GNDA.n5256 2.6629
R17835 GNDA.n5170 GNDA.n82 2.6629
R17836 GNDA.n4834 GNDA.n4833 2.6629
R17837 GNDA.n4742 GNDA.n56 2.6629
R17838 GNDA.n2935 GNDA.n1857 2.6629
R17839 GNDA.n2732 GNDA.n2731 2.6629
R17840 GNDA.n5164 GNDA.n5163 2.6629
R17841 GNDA.t62 GNDA.t108 2.59854
R17842 GNDA.n2644 GNDA.n2643 2.56821
R17843 GNDA.n3139 GNDA.n1824 2.4581
R17844 GNDA.n3219 GNDA.n1531 2.4581
R17845 GNDA.n2739 GNDA.n2732 2.4581
R17846 GNDA.n2796 GNDA.n2795 2.4581
R17847 GNDA.n5049 GNDA.n160 2.4581
R17848 GNDA.n1549 GNDA.n186 2.4581
R17849 GNDA.n1676 GNDA.n1550 2.4581
R17850 GNDA.n1714 GNDA.n1713 2.4581
R17851 GNDA.n4892 GNDA.n4891 2.4581
R17852 GNDA.n5257 GNDA.n56 2.4581
R17853 GNDA.n5171 GNDA.n5170 2.4581
R17854 GNDA.n4743 GNDA.n4742 2.4581
R17855 GNDA.n2731 GNDA.n2684 2.4581
R17856 GNDA.n5164 GNDA.n82 2.4581
R17857 GNDA.n5097 GNDA.n5096 2.4581
R17858 GNDA.n3226 GNDA.n1528 2.44675
R17859 GNDA.n3226 GNDA.n3225 2.44675
R17860 GNDA.n2653 GNDA.n2649 2.42758
R17861 GNDA.n2493 GNDA.n2492 2.39683
R17862 GNDA.n3380 GNDA.n3379 2.38247
R17863 GNDA.n4610 GNDA.n4609 2.38247
R17864 GNDA.n3852 GNDA.n3851 2.38247
R17865 GNDA.n3386 GNDA.n3385 2.38212
R17866 GNDA.t214 GNDA.t143 2.36609
R17867 GNDA.t133 GNDA.t57 2.36609
R17868 GNDA.t115 GNDA.t202 2.36609
R17869 GNDA.t203 GNDA.t104 2.36609
R17870 GNDA.n3701 GNDA.n568 2.34946
R17871 GNDA.n2583 GNDA.n2582 2.30736
R17872 GNDA.n3660 GNDA.n3659 2.30736
R17873 GNDA.n4568 GNDA.n4567 2.30736
R17874 GNDA.n4492 GNDA.n4491 2.30736
R17875 GNDA.n4410 GNDA.n4409 2.30736
R17876 GNDA.n4328 GNDA.n4327 2.30736
R17877 GNDA.n4246 GNDA.n4245 2.30736
R17878 GNDA.n4000 GNDA.n3999 2.30736
R17879 GNDA.n4164 GNDA.n4163 2.30736
R17880 GNDA.n4082 GNDA.n4081 2.30736
R17881 GNDA.n3897 GNDA.n3896 2.30736
R17882 GNDA.n3839 GNDA.n3838 2.30736
R17883 GNDA.n3763 GNDA.n3762 2.30736
R17884 GNDA.n1438 GNDA.n1437 2.30736
R17885 GNDA.n1362 GNDA.n1361 2.30736
R17886 GNDA.n1280 GNDA.n1279 2.30736
R17887 GNDA.n952 GNDA.n951 2.30736
R17888 GNDA.n1198 GNDA.n1197 2.30736
R17889 GNDA.n1116 GNDA.n1115 2.30736
R17890 GNDA.n1034 GNDA.n1033 2.30736
R17891 GNDA.n849 GNDA.n848 2.30736
R17892 GNDA.n698 GNDA.n697 2.30736
R17893 GNDA.n3454 GNDA.n3453 2.30736
R17894 GNDA.n3519 GNDA.n3518 2.30736
R17895 GNDA.n2221 GNDA.n2220 2.30736
R17896 GNDA.n2339 GNDA.n2338 2.30736
R17897 GNDA.n4616 GNDA.n4615 2.29914
R17898 GNDA.n744 GNDA.n743 2.29914
R17899 GNDA.n740 GNDA.n603 2.29914
R17900 GNDA.n4618 GNDA.n4617 2.29878
R17901 GNDA.n3598 GNDA.n578 2.26187
R17902 GNDA.n3601 GNDA.n575 2.26187
R17903 GNDA.n3565 GNDA.n3564 2.26187
R17904 GNDA.n3333 GNDA.n3329 2.26187
R17905 GNDA.n3543 GNDA.n3542 2.26187
R17906 GNDA.n2715 GNDA.n2714 2.26187
R17907 GNDA.n3229 GNDA.n1525 2.26187
R17908 GNDA.n3533 GNDA.n3531 2.26187
R17909 GNDA.n4599 GNDA.n475 2.26187
R17910 GNDA.n2648 GNDA.n1863 2.26187
R17911 GNDA.n2652 GNDA.n2651 2.26187
R17912 GNDA.n2651 GNDA.n1860 2.26187
R17913 GNDA.n463 GNDA.n450 2.26187
R17914 GNDA.n464 GNDA.n463 2.26187
R17915 GNDA.n3602 GNDA.n3601 2.26187
R17916 GNDA.n3595 GNDA.n577 2.26187
R17917 GNDA.n3591 GNDA.n3590 2.26187
R17918 GNDA.n3566 GNDA.n3565 2.26187
R17919 GNDA.n3544 GNDA.n3543 2.26187
R17920 GNDA.n3230 GNDA.n3229 2.26187
R17921 GNDA.n2697 GNDA.n2696 2.26187
R17922 GNDA.n2273 GNDA.n2270 2.26187
R17923 GNDA.n2278 GNDA.n2267 2.26187
R17924 GNDA.n2285 GNDA.n2284 2.26187
R17925 GNDA.n2645 GNDA.n1862 2.26187
R17926 GNDA.n893 GNDA.n888 2.24241
R17927 GNDA.n891 GNDA.n804 2.24241
R17928 GNDA.n3943 GNDA.n435 2.24241
R17929 GNDA.n529 GNDA.n528 2.24241
R17930 GNDA.n467 GNDA.n462 2.24063
R17931 GNDA.n468 GNDA.n450 2.24063
R17932 GNDA.n3599 GNDA.n577 2.24063
R17933 GNDA.n3605 GNDA.n575 2.24063
R17934 GNDA.n3590 GNDA.n580 2.24063
R17935 GNDA.n3589 GNDA.n579 2.24063
R17936 GNDA.n3563 GNDA.n589 2.24063
R17937 GNDA.n3334 GNDA.n3333 2.24063
R17938 GNDA.n3330 GNDA.n3328 2.24063
R17939 GNDA.n3561 GNDA.n3560 2.24063
R17940 GNDA.n595 GNDA.n594 2.24063
R17941 GNDA.n3541 GNDA.n597 2.24063
R17942 GNDA.n3539 GNDA.n3538 2.24063
R17943 GNDA.n604 GNDA.n602 2.24063
R17944 GNDA.n472 GNDA.n471 2.24063
R17945 GNDA.n448 GNDA.n447 2.24063
R17946 GNDA.n2714 GNDA.n2713 2.24063
R17947 GNDA.n2696 GNDA.n1524 2.24063
R17948 GNDA.n2699 GNDA.n2698 2.24063
R17949 GNDA.n3233 GNDA.n1525 2.24063
R17950 GNDA.n2634 GNDA.n2633 2.24063
R17951 GNDA.n2632 GNDA.n2631 2.24063
R17952 GNDA.n2276 GNDA.n2270 2.24063
R17953 GNDA.n2271 GNDA.n2269 2.24063
R17954 GNDA.n2281 GNDA.n2267 2.24063
R17955 GNDA.n2268 GNDA.n2266 2.24063
R17956 GNDA.n2284 GNDA.n2265 2.24063
R17957 GNDA.n2283 GNDA.n2175 2.24063
R17958 GNDA.n2259 GNDA.n610 2.24063
R17959 GNDA.n2262 GNDA.n2261 2.24063
R17960 GNDA.n2263 GNDA.n2260 2.24063
R17961 GNDA.n3529 GNDA.n608 2.24063
R17962 GNDA.n609 GNDA.n607 2.24063
R17963 GNDA.n3526 GNDA.n3525 2.24063
R17964 GNDA.n3397 GNDA.n3391 2.24063
R17965 GNDA.n3393 GNDA.n3392 2.24063
R17966 GNDA.n3398 GNDA.n652 2.24063
R17967 GNDA.n3387 GNDA.n738 2.24063
R17968 GNDA.n3388 GNDA.n737 2.24063
R17969 GNDA.n3389 GNDA.n736 2.24063
R17970 GNDA.n887 GNDA.n805 2.24063
R17971 GNDA.n3375 GNDA.n752 2.24063
R17972 GNDA.n3376 GNDA.n751 2.24063
R17973 GNDA.n3377 GNDA.n750 2.24063
R17974 GNDA.n3371 GNDA.n757 2.24063
R17975 GNDA.n3372 GNDA.n756 2.24063
R17976 GNDA.n3373 GNDA.n755 2.24063
R17977 GNDA.n3367 GNDA.n762 2.24063
R17978 GNDA.n3368 GNDA.n761 2.24063
R17979 GNDA.n3369 GNDA.n760 2.24063
R17980 GNDA.n1458 GNDA.n767 2.24063
R17981 GNDA.n1459 GNDA.n766 2.24063
R17982 GNDA.n1460 GNDA.n765 2.24063
R17983 GNDA.n1454 GNDA.n772 2.24063
R17984 GNDA.n1455 GNDA.n771 2.24063
R17985 GNDA.n1456 GNDA.n770 2.24063
R17986 GNDA.n1444 GNDA.n570 2.24063
R17987 GNDA.n1447 GNDA.n1446 2.24063
R17988 GNDA.n1448 GNDA.n1445 2.24063
R17989 GNDA.n3706 GNDA.n533 2.24063
R17990 GNDA.n565 GNDA.n564 2.24063
R17991 GNDA.n3707 GNDA.n563 2.24063
R17992 GNDA.n3849 GNDA.n531 2.24063
R17993 GNDA.n532 GNDA.n530 2.24063
R17994 GNDA.n3846 GNDA.n3845 2.24063
R17995 GNDA.n4605 GNDA.n440 2.24063
R17996 GNDA.n4606 GNDA.n439 2.24063
R17997 GNDA.n4607 GNDA.n438 2.24063
R17998 GNDA.n4601 GNDA.n445 2.24063
R17999 GNDA.n4602 GNDA.n444 2.24063
R18000 GNDA.n4603 GNDA.n443 2.24063
R18001 GNDA.n3944 GNDA.n527 2.24063
R18002 GNDA.n4593 GNDA.n481 2.24063
R18003 GNDA.n4594 GNDA.n480 2.24063
R18004 GNDA.n4595 GNDA.n479 2.24063
R18005 GNDA.n4589 GNDA.n486 2.24063
R18006 GNDA.n4590 GNDA.n485 2.24063
R18007 GNDA.n4591 GNDA.n484 2.24063
R18008 GNDA.n4585 GNDA.n491 2.24063
R18009 GNDA.n4586 GNDA.n490 2.24063
R18010 GNDA.n4587 GNDA.n489 2.24063
R18011 GNDA.n4581 GNDA.n496 2.24063
R18012 GNDA.n4582 GNDA.n495 2.24063
R18013 GNDA.n4583 GNDA.n494 2.24063
R18014 GNDA.n4577 GNDA.n4576 2.24063
R18015 GNDA.n4578 GNDA.n4575 2.24063
R18016 GNDA.n4579 GNDA.n4574 2.24063
R18017 GNDA.n3531 GNDA.n606 2.24063
R18018 GNDA.n3532 GNDA.n605 2.24063
R18019 GNDA.n4597 GNDA.n475 2.24063
R18020 GNDA.n4598 GNDA.n476 2.24063
R18021 GNDA.n3702 GNDA.n567 2.24063
R18022 GNDA.n569 GNDA.n566 2.24063
R18023 GNDA.n3699 GNDA.n3698 2.24063
R18024 GNDA.n2649 GNDA.n1862 2.24063
R18025 GNDA.n3594 GNDA.n578 2.24063
R18026 GNDA.n3604 GNDA.n3603 2.24063
R18027 GNDA.n3567 GNDA.n3566 2.24063
R18028 GNDA.n3562 GNDA.n592 2.24063
R18029 GNDA.n3545 GNDA.n3544 2.24063
R18030 GNDA.n3540 GNDA.n600 2.24063
R18031 GNDA.n470 GNDA.n469 2.24063
R18032 GNDA.n2812 GNDA.n2700 2.24063
R18033 GNDA.n2811 GNDA.n2810 2.24063
R18034 GNDA.n3232 GNDA.n3231 2.24063
R18035 GNDA.n2635 GNDA.n2624 2.24063
R18036 GNDA.n2644 GNDA.n1863 2.24063
R18037 GNDA.n2653 GNDA.n2652 2.24063
R18038 GNDA.n2655 GNDA.n2654 2.24063
R18039 GNDA.n2712 GNDA.n2703 2.22018
R18040 GNDA.n2809 GNDA.n2716 2.22018
R18041 GNDA.n2626 GNDA.n2625 2.22018
R18042 GNDA.n3365 GNDA.n3342 2.19633
R18043 GNDA.n3586 GNDA.n3585 2.19633
R18044 GNDA.n3570 GNDA.n3569 2.19633
R18045 GNDA.n328 GNDA.n56 2.18124
R18046 GNDA.n5053 GNDA.n160 2.18124
R18047 GNDA.n2732 GNDA.n1833 2.18124
R18048 GNDA.n389 GNDA.n82 2.18124
R18049 GNDA.n1796 GNDA.n1550 2.18124
R18050 GNDA.n3148 GNDA.n1824 2.18124
R18051 GNDA.n2636 GNDA.n2635 2.16717
R18052 GNDA.n3580 GNDA.n3578 2.15331
R18053 GNDA.n3577 GNDA.n3576 2.15331
R18054 GNDA.n1531 GNDA.n1511 2.1509
R18055 GNDA.n2797 GNDA.n2796 2.1509
R18056 GNDA.n4984 GNDA.n186 2.1509
R18057 GNDA.n1713 GNDA.n1712 2.1509
R18058 GNDA.n4910 GNDA.n4892 2.1509
R18059 GNDA.n5189 GNDA.n5171 2.1509
R18060 GNDA.n4769 GNDA.n4743 2.1509
R18061 GNDA.n2690 GNDA.n2684 2.1509
R18062 GNDA.n5107 GNDA.n5097 2.1509
R18063 GNDA.n3138 GNDA.n3047 2.13383
R18064 GNDA.n2741 GNDA.n2740 2.13383
R18065 GNDA.n5048 GNDA.n164 2.13383
R18066 GNDA.n4833 GNDA.n4720 2.13383
R18067 GNDA.n1677 GNDA.n1675 2.13383
R18068 GNDA.n4977 GNDA.n4864 2.13383
R18069 GNDA.n5256 GNDA.n57 2.13383
R18070 GNDA.n2904 GNDA.n1857 2.13383
R18071 GNDA.n5163 GNDA.n5162 2.13383
R18072 GNDA.n3381 GNDA.n3380 2.09414
R18073 GNDA.n4611 GNDA.n4610 2.09414
R18074 GNDA.n3851 GNDA.n3850 2.09414
R18075 GNDA.n3385 GNDA.n3384 2.09414
R18076 GNDA.n133 GNDA.n56 2.08643
R18077 GNDA.n162 GNDA.n160 2.08643
R18078 GNDA.n2732 GNDA.n1832 2.08643
R18079 GNDA.n84 GNDA.n82 2.08643
R18080 GNDA.n1799 GNDA.n1550 2.08643
R18081 GNDA.n1827 GNDA.n1824 2.08643
R18082 GNDA.n3615 GNDA.n3614 2.00747
R18083 GNDA.n1453 GNDA.n1452 2.00747
R18084 GNDA.t167 GNDA.t303 1.98114
R18085 GNDA.t240 GNDA.t43 1.98114
R18086 GNDA.n3138 GNDA.n3137 1.9461
R18087 GNDA.n2740 GNDA.n1493 1.9461
R18088 GNDA.n5048 GNDA.n5047 1.9461
R18089 GNDA.n1678 GNDA.n1677 1.9461
R18090 GNDA.n4977 GNDA.n4976 1.9461
R18091 GNDA.n5256 GNDA.n5255 1.9461
R18092 GNDA.n4833 GNDA.n4832 1.9461
R18093 GNDA.n2907 GNDA.n1857 1.9461
R18094 GNDA.n5163 GNDA.n22 1.9461
R18095 GNDA.n583 GNDA.n574 1.94497
R18096 GNDA.n3336 GNDA.n3335 1.94497
R18097 GNDA.n4615 GNDA.n4614 1.93383
R18098 GNDA.n745 GNDA.n744 1.93383
R18099 GNDA.n741 GNDA.n740 1.93383
R18100 GNDA.n4619 GNDA.n4618 1.93383
R18101 GNDA.n3610 GNDA.n568 1.91062
R18102 GNDA.n1450 GNDA.t112 1.86807
R18103 GNDA.n3584 GNDA.t95 1.86807
R18104 GNDA.n3612 GNDA.t26 1.86807
R18105 GNDA.n3234 GNDA.n3233 1.71925
R18106 GNDA.n2468 GNDA.n1900 1.70567
R18107 GNDA.n2468 GNDA.n1899 1.70567
R18108 GNDA.n2468 GNDA.n1898 1.70567
R18109 GNDA.n2468 GNDA.n1897 1.70567
R18110 GNDA.n2468 GNDA.n1896 1.70567
R18111 GNDA.n2468 GNDA.n1895 1.70567
R18112 GNDA.n2468 GNDA.n1894 1.70567
R18113 GNDA.n2468 GNDA.n1893 1.70567
R18114 GNDA.n2468 GNDA.n1892 1.70567
R18115 GNDA.n2468 GNDA.n1891 1.70567
R18116 GNDA.n2468 GNDA.n1890 1.70567
R18117 GNDA.n2468 GNDA.n1889 1.70567
R18118 GNDA.n2468 GNDA.n1888 1.70567
R18119 GNDA.n2468 GNDA.n1887 1.70567
R18120 GNDA.n2468 GNDA.n1886 1.70567
R18121 GNDA.n2468 GNDA.n1885 1.70567
R18122 GNDA.n2470 GNDA.n2469 1.70567
R18123 GNDA.n2434 GNDA.n1884 1.70567
R18124 GNDA.n2436 GNDA.n1884 1.70567
R18125 GNDA.n2438 GNDA.n1884 1.70567
R18126 GNDA.n2440 GNDA.n1884 1.70567
R18127 GNDA.n2442 GNDA.n1884 1.70567
R18128 GNDA.n2444 GNDA.n1884 1.70567
R18129 GNDA.n2446 GNDA.n1884 1.70567
R18130 GNDA.n2448 GNDA.n1884 1.70567
R18131 GNDA.n2450 GNDA.n1884 1.70567
R18132 GNDA.n2452 GNDA.n1884 1.70567
R18133 GNDA.n2454 GNDA.n1884 1.70567
R18134 GNDA.n2456 GNDA.n1884 1.70567
R18135 GNDA.n2458 GNDA.n1884 1.70567
R18136 GNDA.n2460 GNDA.n1884 1.70567
R18137 GNDA.n2462 GNDA.n1884 1.70567
R18138 GNDA.n2464 GNDA.n1884 1.70567
R18139 GNDA.n1919 GNDA.n1918 1.70567
R18140 GNDA.n2470 GNDA.n1883 1.70567
R18141 GNDA.n1921 GNDA.n1918 1.70567
R18142 GNDA.n2470 GNDA.n1882 1.70567
R18143 GNDA.n1923 GNDA.n1918 1.70567
R18144 GNDA.n2470 GNDA.n1881 1.70567
R18145 GNDA.n1925 GNDA.n1918 1.70567
R18146 GNDA.n2470 GNDA.n1880 1.70567
R18147 GNDA.n1927 GNDA.n1918 1.70567
R18148 GNDA.n2470 GNDA.n1879 1.70567
R18149 GNDA.n1929 GNDA.n1918 1.70567
R18150 GNDA.n2470 GNDA.n1878 1.70567
R18151 GNDA.n1931 GNDA.n1918 1.70567
R18152 GNDA.n2470 GNDA.n1877 1.70567
R18153 GNDA.n1933 GNDA.n1918 1.70567
R18154 GNDA.n2470 GNDA.n1876 1.70567
R18155 GNDA.n1935 GNDA.n1918 1.70567
R18156 GNDA.n2470 GNDA.n1875 1.70567
R18157 GNDA.n1937 GNDA.n1918 1.70567
R18158 GNDA.n2470 GNDA.n1874 1.70567
R18159 GNDA.n1939 GNDA.n1918 1.70567
R18160 GNDA.n2470 GNDA.n1873 1.70567
R18161 GNDA.n1941 GNDA.n1918 1.70567
R18162 GNDA.n2470 GNDA.n1872 1.70567
R18163 GNDA.n1943 GNDA.n1918 1.70567
R18164 GNDA.n2470 GNDA.n1871 1.70567
R18165 GNDA.n1945 GNDA.n1918 1.70567
R18166 GNDA.n2470 GNDA.n1870 1.70567
R18167 GNDA.n1947 GNDA.n1918 1.70567
R18168 GNDA.n2470 GNDA.n1869 1.70567
R18169 GNDA.n1949 GNDA.n1918 1.70567
R18170 GNDA.n2470 GNDA.n1868 1.70567
R18171 GNDA.n2466 GNDA.n1867 1.70567
R18172 GNDA.n1951 GNDA.n1918 1.70567
R18173 GNDA.n2378 GNDA.n2065 1.70567
R18174 GNDA.n2378 GNDA.n2064 1.70567
R18175 GNDA.n2378 GNDA.n2063 1.70567
R18176 GNDA.n2378 GNDA.n2062 1.70567
R18177 GNDA.n2378 GNDA.n2061 1.70567
R18178 GNDA.n2378 GNDA.n2060 1.70567
R18179 GNDA.n2378 GNDA.n2059 1.70567
R18180 GNDA.n2378 GNDA.n2058 1.70567
R18181 GNDA.n2378 GNDA.n2057 1.70567
R18182 GNDA.n2378 GNDA.n2056 1.70567
R18183 GNDA.n2378 GNDA.n2055 1.70567
R18184 GNDA.n2378 GNDA.n2054 1.70567
R18185 GNDA.n2378 GNDA.n2053 1.70567
R18186 GNDA.n2378 GNDA.n2052 1.70567
R18187 GNDA.n2378 GNDA.n2051 1.70567
R18188 GNDA.n2378 GNDA.n2050 1.70567
R18189 GNDA.n2345 GNDA.n2083 1.70567
R18190 GNDA.n2347 GNDA.n2083 1.70567
R18191 GNDA.n2349 GNDA.n2083 1.70567
R18192 GNDA.n2351 GNDA.n2083 1.70567
R18193 GNDA.n2353 GNDA.n2083 1.70567
R18194 GNDA.n2355 GNDA.n2083 1.70567
R18195 GNDA.n2357 GNDA.n2083 1.70567
R18196 GNDA.n2359 GNDA.n2083 1.70567
R18197 GNDA.n2361 GNDA.n2083 1.70567
R18198 GNDA.n2363 GNDA.n2083 1.70567
R18199 GNDA.n2365 GNDA.n2083 1.70567
R18200 GNDA.n2367 GNDA.n2083 1.70567
R18201 GNDA.n2369 GNDA.n2083 1.70567
R18202 GNDA.n2371 GNDA.n2083 1.70567
R18203 GNDA.n2373 GNDA.n2083 1.70567
R18204 GNDA.n2084 GNDA.n2049 1.70567
R18205 GNDA.n2133 GNDA.n2117 1.70567
R18206 GNDA.n2085 GNDA.n2084 1.70567
R18207 GNDA.n2133 GNDA.n2118 1.70567
R18208 GNDA.n2087 GNDA.n2084 1.70567
R18209 GNDA.n2133 GNDA.n2119 1.70567
R18210 GNDA.n2089 GNDA.n2084 1.70567
R18211 GNDA.n2133 GNDA.n2120 1.70567
R18212 GNDA.n2091 GNDA.n2084 1.70567
R18213 GNDA.n2133 GNDA.n2121 1.70567
R18214 GNDA.n2093 GNDA.n2084 1.70567
R18215 GNDA.n2133 GNDA.n2122 1.70567
R18216 GNDA.n2095 GNDA.n2084 1.70567
R18217 GNDA.n2133 GNDA.n2123 1.70567
R18218 GNDA.n2097 GNDA.n2084 1.70567
R18219 GNDA.n2133 GNDA.n2124 1.70567
R18220 GNDA.n2099 GNDA.n2084 1.70567
R18221 GNDA.n2133 GNDA.n2125 1.70567
R18222 GNDA.n2101 GNDA.n2084 1.70567
R18223 GNDA.n2133 GNDA.n2126 1.70567
R18224 GNDA.n2103 GNDA.n2084 1.70567
R18225 GNDA.n2133 GNDA.n2127 1.70567
R18226 GNDA.n2105 GNDA.n2084 1.70567
R18227 GNDA.n2133 GNDA.n2128 1.70567
R18228 GNDA.n2107 GNDA.n2084 1.70567
R18229 GNDA.n2133 GNDA.n2129 1.70567
R18230 GNDA.n2109 GNDA.n2084 1.70567
R18231 GNDA.n2133 GNDA.n2130 1.70567
R18232 GNDA.n2111 GNDA.n2084 1.70567
R18233 GNDA.n2133 GNDA.n2131 1.70567
R18234 GNDA.n2113 GNDA.n2084 1.70567
R18235 GNDA.n2133 GNDA.n2132 1.70567
R18236 GNDA.n2115 GNDA.n2084 1.70567
R18237 GNDA.n2134 GNDA.n2133 1.70567
R18238 GNDA.n2376 GNDA.n2375 1.70567
R18239 GNDA.n2432 GNDA.n2431 1.70567
R18240 GNDA.n2433 GNDA.n1983 1.70567
R18241 GNDA.n2433 GNDA.n1982 1.70567
R18242 GNDA.n2433 GNDA.n1981 1.70567
R18243 GNDA.n2433 GNDA.n1980 1.70567
R18244 GNDA.n2433 GNDA.n1979 1.70567
R18245 GNDA.n2433 GNDA.n1978 1.70567
R18246 GNDA.n2433 GNDA.n1977 1.70567
R18247 GNDA.n2433 GNDA.n1976 1.70567
R18248 GNDA.n2433 GNDA.n1975 1.70567
R18249 GNDA.n2433 GNDA.n1974 1.70567
R18250 GNDA.n2433 GNDA.n1973 1.70567
R18251 GNDA.n2433 GNDA.n1972 1.70567
R18252 GNDA.n2433 GNDA.n1971 1.70567
R18253 GNDA.n2433 GNDA.n1970 1.70567
R18254 GNDA.n2433 GNDA.n1969 1.70567
R18255 GNDA.n2433 GNDA.n1968 1.70567
R18256 GNDA.n2433 GNDA.n1967 1.70567
R18257 GNDA.n2379 GNDA.n1984 1.70567
R18258 GNDA.n2381 GNDA.n1984 1.70567
R18259 GNDA.n2383 GNDA.n1984 1.70567
R18260 GNDA.n2385 GNDA.n1984 1.70567
R18261 GNDA.n2387 GNDA.n1984 1.70567
R18262 GNDA.n2389 GNDA.n1984 1.70567
R18263 GNDA.n2391 GNDA.n1984 1.70567
R18264 GNDA.n2393 GNDA.n1984 1.70567
R18265 GNDA.n2395 GNDA.n1984 1.70567
R18266 GNDA.n2397 GNDA.n1984 1.70567
R18267 GNDA.n2399 GNDA.n1984 1.70567
R18268 GNDA.n2401 GNDA.n1984 1.70567
R18269 GNDA.n2403 GNDA.n1984 1.70567
R18270 GNDA.n2405 GNDA.n1984 1.70567
R18271 GNDA.n2407 GNDA.n1984 1.70567
R18272 GNDA.n2428 GNDA.n2001 1.70567
R18273 GNDA.n2426 GNDA.n2425 1.70567
R18274 GNDA.n2427 GNDA.n2033 1.70567
R18275 GNDA.n2425 GNDA.n2410 1.70567
R18276 GNDA.n2033 GNDA.n2032 1.70567
R18277 GNDA.n2425 GNDA.n2411 1.70567
R18278 GNDA.n2033 GNDA.n2031 1.70567
R18279 GNDA.n2425 GNDA.n2412 1.70567
R18280 GNDA.n2033 GNDA.n2030 1.70567
R18281 GNDA.n2425 GNDA.n2413 1.70567
R18282 GNDA.n2033 GNDA.n2029 1.70567
R18283 GNDA.n2425 GNDA.n2414 1.70567
R18284 GNDA.n2033 GNDA.n2028 1.70567
R18285 GNDA.n2425 GNDA.n2415 1.70567
R18286 GNDA.n2033 GNDA.n2027 1.70567
R18287 GNDA.n2425 GNDA.n2416 1.70567
R18288 GNDA.n2033 GNDA.n2026 1.70567
R18289 GNDA.n2425 GNDA.n2417 1.70567
R18290 GNDA.n2033 GNDA.n2025 1.70567
R18291 GNDA.n2425 GNDA.n2418 1.70567
R18292 GNDA.n2033 GNDA.n2024 1.70567
R18293 GNDA.n2425 GNDA.n2419 1.70567
R18294 GNDA.n2033 GNDA.n2023 1.70567
R18295 GNDA.n2425 GNDA.n2420 1.70567
R18296 GNDA.n2033 GNDA.n2022 1.70567
R18297 GNDA.n2425 GNDA.n2421 1.70567
R18298 GNDA.n2033 GNDA.n2021 1.70567
R18299 GNDA.n2425 GNDA.n2422 1.70567
R18300 GNDA.n2033 GNDA.n2020 1.70567
R18301 GNDA.n2425 GNDA.n2423 1.70567
R18302 GNDA.n2033 GNDA.n2019 1.70567
R18303 GNDA.n2425 GNDA.n2424 1.70567
R18304 GNDA.n2033 GNDA.n2018 1.70567
R18305 GNDA.n2425 GNDA.n2017 1.70567
R18306 GNDA.n2230 GNDA.n615 1.69433
R18307 GNDA.n2239 GNDA.n615 1.69433
R18308 GNDA.n2248 GNDA.n615 1.69433
R18309 GNDA.n3521 GNDA.n624 1.69433
R18310 GNDA.n3521 GNDA.n621 1.69433
R18311 GNDA.n3521 GNDA.n618 1.69433
R18312 GNDA.n3456 GNDA.n636 1.69433
R18313 GNDA.n3456 GNDA.n633 1.69433
R18314 GNDA.n3456 GNDA.n630 1.69433
R18315 GNDA.n707 GNDA.n639 1.69433
R18316 GNDA.n716 GNDA.n639 1.69433
R18317 GNDA.n725 GNDA.n639 1.69433
R18318 GNDA.n858 GNDA.n778 1.69433
R18319 GNDA.n867 GNDA.n778 1.69433
R18320 GNDA.n876 GNDA.n778 1.69433
R18321 GNDA.n1036 GNDA.n964 1.69433
R18322 GNDA.n1036 GNDA.n961 1.69433
R18323 GNDA.n1036 GNDA.n958 1.69433
R18324 GNDA.n1118 GNDA.n1046 1.69433
R18325 GNDA.n1118 GNDA.n1043 1.69433
R18326 GNDA.n1118 GNDA.n1040 1.69433
R18327 GNDA.n1200 GNDA.n1128 1.69433
R18328 GNDA.n1200 GNDA.n1125 1.69433
R18329 GNDA.n1200 GNDA.n1122 1.69433
R18330 GNDA.n954 GNDA.n788 1.69433
R18331 GNDA.n954 GNDA.n785 1.69433
R18332 GNDA.n954 GNDA.n782 1.69433
R18333 GNDA.n1282 GNDA.n1210 1.69433
R18334 GNDA.n1282 GNDA.n1207 1.69433
R18335 GNDA.n1282 GNDA.n1204 1.69433
R18336 GNDA.n1364 GNDA.n1292 1.69433
R18337 GNDA.n1364 GNDA.n1289 1.69433
R18338 GNDA.n1364 GNDA.n1286 1.69433
R18339 GNDA.n1440 GNDA.n1373 1.69433
R18340 GNDA.n1440 GNDA.n1370 1.69433
R18341 GNDA.n1440 GNDA.n1367 1.69433
R18342 GNDA.n3765 GNDA.n548 1.69433
R18343 GNDA.n3765 GNDA.n545 1.69433
R18344 GNDA.n3765 GNDA.n542 1.69433
R18345 GNDA.n3841 GNDA.n3774 1.69433
R18346 GNDA.n3841 GNDA.n3771 1.69433
R18347 GNDA.n3841 GNDA.n3768 1.69433
R18348 GNDA.n3906 GNDA.n502 1.69433
R18349 GNDA.n3915 GNDA.n502 1.69433
R18350 GNDA.n3924 GNDA.n502 1.69433
R18351 GNDA.n4084 GNDA.n4012 1.69433
R18352 GNDA.n4084 GNDA.n4009 1.69433
R18353 GNDA.n4084 GNDA.n4006 1.69433
R18354 GNDA.n4166 GNDA.n4094 1.69433
R18355 GNDA.n4166 GNDA.n4091 1.69433
R18356 GNDA.n4166 GNDA.n4088 1.69433
R18357 GNDA.n4002 GNDA.n512 1.69433
R18358 GNDA.n4002 GNDA.n509 1.69433
R18359 GNDA.n4002 GNDA.n506 1.69433
R18360 GNDA.n4248 GNDA.n4176 1.69433
R18361 GNDA.n4248 GNDA.n4173 1.69433
R18362 GNDA.n4248 GNDA.n4170 1.69433
R18363 GNDA.n4330 GNDA.n4258 1.69433
R18364 GNDA.n4330 GNDA.n4255 1.69433
R18365 GNDA.n4330 GNDA.n4252 1.69433
R18366 GNDA.n4412 GNDA.n4340 1.69433
R18367 GNDA.n4412 GNDA.n4337 1.69433
R18368 GNDA.n4412 GNDA.n4334 1.69433
R18369 GNDA.n4494 GNDA.n4422 1.69433
R18370 GNDA.n4494 GNDA.n4419 1.69433
R18371 GNDA.n4494 GNDA.n4416 1.69433
R18372 GNDA.n4570 GNDA.n4503 1.69433
R18373 GNDA.n4570 GNDA.n4500 1.69433
R18374 GNDA.n4570 GNDA.n4497 1.69433
R18375 GNDA.n3669 GNDA.n538 1.69433
R18376 GNDA.n3678 GNDA.n538 1.69433
R18377 GNDA.n3687 GNDA.n538 1.69433
R18378 GNDA.n2640 GNDA.n2480 1.69433
R18379 GNDA.n2640 GNDA.n2477 1.69433
R18380 GNDA.n2640 GNDA.n2474 1.69433
R18381 GNDA.n2639 GNDA.n2555 1.69433
R18382 GNDA.n2639 GNDA.n2552 1.69433
R18383 GNDA.n2639 GNDA.n2549 1.69433
R18384 GNDA.n2343 GNDA.n2160 1.69337
R18385 GNDA.n2343 GNDA.n2159 1.69337
R18386 GNDA.n2343 GNDA.n2157 1.69337
R18387 GNDA.n2343 GNDA.n2156 1.69337
R18388 GNDA.n2343 GNDA.n2154 1.69337
R18389 GNDA.n2343 GNDA.n2153 1.69337
R18390 GNDA.n2343 GNDA.n2151 1.69337
R18391 GNDA.n2343 GNDA.n2150 1.69337
R18392 GNDA.n2224 GNDA.n615 1.6924
R18393 GNDA.n2227 GNDA.n615 1.6924
R18394 GNDA.n2233 GNDA.n615 1.6924
R18395 GNDA.n2236 GNDA.n615 1.6924
R18396 GNDA.n2242 GNDA.n615 1.6924
R18397 GNDA.n2245 GNDA.n615 1.6924
R18398 GNDA.n2251 GNDA.n615 1.6924
R18399 GNDA.n2254 GNDA.n615 1.6924
R18400 GNDA.n3521 GNDA.n626 1.6924
R18401 GNDA.n3521 GNDA.n625 1.6924
R18402 GNDA.n3521 GNDA.n623 1.6924
R18403 GNDA.n3521 GNDA.n622 1.6924
R18404 GNDA.n3521 GNDA.n620 1.6924
R18405 GNDA.n3521 GNDA.n619 1.6924
R18406 GNDA.n3521 GNDA.n617 1.6924
R18407 GNDA.n3521 GNDA.n616 1.6924
R18408 GNDA.n3456 GNDA.n638 1.6924
R18409 GNDA.n3456 GNDA.n637 1.6924
R18410 GNDA.n3456 GNDA.n635 1.6924
R18411 GNDA.n3456 GNDA.n634 1.6924
R18412 GNDA.n3456 GNDA.n632 1.6924
R18413 GNDA.n3456 GNDA.n631 1.6924
R18414 GNDA.n3456 GNDA.n629 1.6924
R18415 GNDA.n3456 GNDA.n628 1.6924
R18416 GNDA.n701 GNDA.n639 1.6924
R18417 GNDA.n704 GNDA.n639 1.6924
R18418 GNDA.n710 GNDA.n639 1.6924
R18419 GNDA.n713 GNDA.n639 1.6924
R18420 GNDA.n719 GNDA.n639 1.6924
R18421 GNDA.n722 GNDA.n639 1.6924
R18422 GNDA.n728 GNDA.n639 1.6924
R18423 GNDA.n731 GNDA.n639 1.6924
R18424 GNDA.n852 GNDA.n778 1.6924
R18425 GNDA.n855 GNDA.n778 1.6924
R18426 GNDA.n861 GNDA.n778 1.6924
R18427 GNDA.n864 GNDA.n778 1.6924
R18428 GNDA.n870 GNDA.n778 1.6924
R18429 GNDA.n873 GNDA.n778 1.6924
R18430 GNDA.n879 GNDA.n778 1.6924
R18431 GNDA.n882 GNDA.n778 1.6924
R18432 GNDA.n1036 GNDA.n966 1.6924
R18433 GNDA.n1036 GNDA.n965 1.6924
R18434 GNDA.n1036 GNDA.n963 1.6924
R18435 GNDA.n1036 GNDA.n962 1.6924
R18436 GNDA.n1036 GNDA.n960 1.6924
R18437 GNDA.n1036 GNDA.n959 1.6924
R18438 GNDA.n1036 GNDA.n957 1.6924
R18439 GNDA.n1036 GNDA.n956 1.6924
R18440 GNDA.n1118 GNDA.n1048 1.6924
R18441 GNDA.n1118 GNDA.n1047 1.6924
R18442 GNDA.n1118 GNDA.n1045 1.6924
R18443 GNDA.n1118 GNDA.n1044 1.6924
R18444 GNDA.n1118 GNDA.n1042 1.6924
R18445 GNDA.n1118 GNDA.n1041 1.6924
R18446 GNDA.n1118 GNDA.n1039 1.6924
R18447 GNDA.n1118 GNDA.n1038 1.6924
R18448 GNDA.n1200 GNDA.n1130 1.6924
R18449 GNDA.n1200 GNDA.n1129 1.6924
R18450 GNDA.n1200 GNDA.n1127 1.6924
R18451 GNDA.n1200 GNDA.n1126 1.6924
R18452 GNDA.n1200 GNDA.n1124 1.6924
R18453 GNDA.n1200 GNDA.n1123 1.6924
R18454 GNDA.n1200 GNDA.n1121 1.6924
R18455 GNDA.n1200 GNDA.n1120 1.6924
R18456 GNDA.n954 GNDA.n790 1.6924
R18457 GNDA.n954 GNDA.n789 1.6924
R18458 GNDA.n954 GNDA.n787 1.6924
R18459 GNDA.n954 GNDA.n786 1.6924
R18460 GNDA.n954 GNDA.n784 1.6924
R18461 GNDA.n954 GNDA.n783 1.6924
R18462 GNDA.n954 GNDA.n781 1.6924
R18463 GNDA.n954 GNDA.n780 1.6924
R18464 GNDA.n1282 GNDA.n1212 1.6924
R18465 GNDA.n1282 GNDA.n1211 1.6924
R18466 GNDA.n1282 GNDA.n1209 1.6924
R18467 GNDA.n1282 GNDA.n1208 1.6924
R18468 GNDA.n1282 GNDA.n1206 1.6924
R18469 GNDA.n1282 GNDA.n1205 1.6924
R18470 GNDA.n1282 GNDA.n1203 1.6924
R18471 GNDA.n1282 GNDA.n1202 1.6924
R18472 GNDA.n1364 GNDA.n1294 1.6924
R18473 GNDA.n1364 GNDA.n1293 1.6924
R18474 GNDA.n1364 GNDA.n1291 1.6924
R18475 GNDA.n1364 GNDA.n1290 1.6924
R18476 GNDA.n1364 GNDA.n1288 1.6924
R18477 GNDA.n1364 GNDA.n1287 1.6924
R18478 GNDA.n1364 GNDA.n1285 1.6924
R18479 GNDA.n1364 GNDA.n1284 1.6924
R18480 GNDA.n1440 GNDA.n1375 1.6924
R18481 GNDA.n1440 GNDA.n1374 1.6924
R18482 GNDA.n1440 GNDA.n1372 1.6924
R18483 GNDA.n1440 GNDA.n1371 1.6924
R18484 GNDA.n1440 GNDA.n1369 1.6924
R18485 GNDA.n1440 GNDA.n1368 1.6924
R18486 GNDA.n1440 GNDA.n1366 1.6924
R18487 GNDA.n1440 GNDA.n1365 1.6924
R18488 GNDA.n3765 GNDA.n550 1.6924
R18489 GNDA.n3765 GNDA.n549 1.6924
R18490 GNDA.n3765 GNDA.n547 1.6924
R18491 GNDA.n3765 GNDA.n546 1.6924
R18492 GNDA.n3765 GNDA.n544 1.6924
R18493 GNDA.n3765 GNDA.n543 1.6924
R18494 GNDA.n3765 GNDA.n541 1.6924
R18495 GNDA.n3765 GNDA.n540 1.6924
R18496 GNDA.n3841 GNDA.n3776 1.6924
R18497 GNDA.n3841 GNDA.n3775 1.6924
R18498 GNDA.n3841 GNDA.n3773 1.6924
R18499 GNDA.n3841 GNDA.n3772 1.6924
R18500 GNDA.n3841 GNDA.n3770 1.6924
R18501 GNDA.n3841 GNDA.n3769 1.6924
R18502 GNDA.n3841 GNDA.n3767 1.6924
R18503 GNDA.n3841 GNDA.n3766 1.6924
R18504 GNDA.n3900 GNDA.n502 1.6924
R18505 GNDA.n3903 GNDA.n502 1.6924
R18506 GNDA.n3909 GNDA.n502 1.6924
R18507 GNDA.n3912 GNDA.n502 1.6924
R18508 GNDA.n3918 GNDA.n502 1.6924
R18509 GNDA.n3921 GNDA.n502 1.6924
R18510 GNDA.n3927 GNDA.n502 1.6924
R18511 GNDA.n3930 GNDA.n502 1.6924
R18512 GNDA.n4084 GNDA.n4014 1.6924
R18513 GNDA.n4084 GNDA.n4013 1.6924
R18514 GNDA.n4084 GNDA.n4011 1.6924
R18515 GNDA.n4084 GNDA.n4010 1.6924
R18516 GNDA.n4084 GNDA.n4008 1.6924
R18517 GNDA.n4084 GNDA.n4007 1.6924
R18518 GNDA.n4084 GNDA.n4005 1.6924
R18519 GNDA.n4084 GNDA.n4004 1.6924
R18520 GNDA.n4166 GNDA.n4096 1.6924
R18521 GNDA.n4166 GNDA.n4095 1.6924
R18522 GNDA.n4166 GNDA.n4093 1.6924
R18523 GNDA.n4166 GNDA.n4092 1.6924
R18524 GNDA.n4166 GNDA.n4090 1.6924
R18525 GNDA.n4166 GNDA.n4089 1.6924
R18526 GNDA.n4166 GNDA.n4087 1.6924
R18527 GNDA.n4166 GNDA.n4086 1.6924
R18528 GNDA.n4002 GNDA.n514 1.6924
R18529 GNDA.n4002 GNDA.n513 1.6924
R18530 GNDA.n4002 GNDA.n511 1.6924
R18531 GNDA.n4002 GNDA.n510 1.6924
R18532 GNDA.n4002 GNDA.n508 1.6924
R18533 GNDA.n4002 GNDA.n507 1.6924
R18534 GNDA.n4002 GNDA.n505 1.6924
R18535 GNDA.n4002 GNDA.n504 1.6924
R18536 GNDA.n4248 GNDA.n4178 1.6924
R18537 GNDA.n4248 GNDA.n4177 1.6924
R18538 GNDA.n4248 GNDA.n4175 1.6924
R18539 GNDA.n4248 GNDA.n4174 1.6924
R18540 GNDA.n4248 GNDA.n4172 1.6924
R18541 GNDA.n4248 GNDA.n4171 1.6924
R18542 GNDA.n4248 GNDA.n4169 1.6924
R18543 GNDA.n4248 GNDA.n4168 1.6924
R18544 GNDA.n4330 GNDA.n4260 1.6924
R18545 GNDA.n4330 GNDA.n4259 1.6924
R18546 GNDA.n4330 GNDA.n4257 1.6924
R18547 GNDA.n4330 GNDA.n4256 1.6924
R18548 GNDA.n4330 GNDA.n4254 1.6924
R18549 GNDA.n4330 GNDA.n4253 1.6924
R18550 GNDA.n4330 GNDA.n4251 1.6924
R18551 GNDA.n4330 GNDA.n4250 1.6924
R18552 GNDA.n4412 GNDA.n4342 1.6924
R18553 GNDA.n4412 GNDA.n4341 1.6924
R18554 GNDA.n4412 GNDA.n4339 1.6924
R18555 GNDA.n4412 GNDA.n4338 1.6924
R18556 GNDA.n4412 GNDA.n4336 1.6924
R18557 GNDA.n4412 GNDA.n4335 1.6924
R18558 GNDA.n4412 GNDA.n4333 1.6924
R18559 GNDA.n4412 GNDA.n4332 1.6924
R18560 GNDA.n4494 GNDA.n4424 1.6924
R18561 GNDA.n4494 GNDA.n4423 1.6924
R18562 GNDA.n4494 GNDA.n4421 1.6924
R18563 GNDA.n4494 GNDA.n4420 1.6924
R18564 GNDA.n4494 GNDA.n4418 1.6924
R18565 GNDA.n4494 GNDA.n4417 1.6924
R18566 GNDA.n4494 GNDA.n4415 1.6924
R18567 GNDA.n4494 GNDA.n4414 1.6924
R18568 GNDA.n4570 GNDA.n4505 1.6924
R18569 GNDA.n4570 GNDA.n4504 1.6924
R18570 GNDA.n4570 GNDA.n4502 1.6924
R18571 GNDA.n4570 GNDA.n4501 1.6924
R18572 GNDA.n4570 GNDA.n4499 1.6924
R18573 GNDA.n4570 GNDA.n4498 1.6924
R18574 GNDA.n4570 GNDA.n4496 1.6924
R18575 GNDA.n4570 GNDA.n4495 1.6924
R18576 GNDA.n3663 GNDA.n538 1.6924
R18577 GNDA.n3666 GNDA.n538 1.6924
R18578 GNDA.n3672 GNDA.n538 1.6924
R18579 GNDA.n3675 GNDA.n538 1.6924
R18580 GNDA.n3681 GNDA.n538 1.6924
R18581 GNDA.n3684 GNDA.n538 1.6924
R18582 GNDA.n3690 GNDA.n538 1.6924
R18583 GNDA.n3693 GNDA.n538 1.6924
R18584 GNDA.n2640 GNDA.n2545 1.6924
R18585 GNDA.n2640 GNDA.n2481 1.6924
R18586 GNDA.n2640 GNDA.n2479 1.6924
R18587 GNDA.n2640 GNDA.n2478 1.6924
R18588 GNDA.n2640 GNDA.n2476 1.6924
R18589 GNDA.n2640 GNDA.n2475 1.6924
R18590 GNDA.n2640 GNDA.n2473 1.6924
R18591 GNDA.n2640 GNDA.n2472 1.6924
R18592 GNDA.n2639 GNDA.n2557 1.6924
R18593 GNDA.n2639 GNDA.n2556 1.6924
R18594 GNDA.n2639 GNDA.n2554 1.6924
R18595 GNDA.n2639 GNDA.n2553 1.6924
R18596 GNDA.n2639 GNDA.n2551 1.6924
R18597 GNDA.n2639 GNDA.n2550 1.6924
R18598 GNDA.n2639 GNDA.n2548 1.6924
R18599 GNDA.n2639 GNDA.n2547 1.6924
R18600 GNDA.n2343 GNDA.n2342 1.6924
R18601 GNDA.n2343 GNDA.n2158 1.6924
R18602 GNDA.n2343 GNDA.n2155 1.6924
R18603 GNDA.n2343 GNDA.n2152 1.6924
R18604 GNDA.n3569 GNDA.n3568 1.56997
R18605 GNDA.n3587 GNDA.n3586 1.56997
R18606 GNDA.t272 GNDA.n105 1.51652
R18607 GNDA.n474 GNDA.n473 1.5005
R18608 GNDA.n3537 GNDA.n3535 1.5005
R18609 GNDA.n895 GNDA.n894 1.5005
R18610 GNDA.n3938 GNDA.n3937 1.5005
R18611 GNDA.n3218 GNDA.n3217 1.47392
R18612 GNDA.n1719 GNDA.n1718 1.47392
R18613 GNDA.n4863 GNDA.n228 1.47392
R18614 GNDA.n4840 GNDA.n4837 1.47392
R18615 GNDA.n2937 GNDA.n2936 1.47392
R18616 GNDA.n5086 GNDA.n87 1.47392
R18617 GNDA.n2627 GNDA.n2626 1.22446
R18618 GNDA.n470 GNDA.n468 1.07342
R18619 GNDA.n3541 GNDA.n3540 1.07342
R18620 GNDA.n3568 GNDA.n3567 1.063
R18621 GNDA.n3592 GNDA.n3587 1.063
R18622 GNDA.n2659 GNDA.n2655 1.05258
R18623 GNDA.n2629 GNDA.n2628 0.854667
R18624 GNDA.n3136 GNDA.n3048 0.8197
R18625 GNDA.n3133 GNDA.n3132 0.8197
R18626 GNDA.n3126 GNDA.n3116 0.8197
R18627 GNDA.n3125 GNDA.n3121 0.8197
R18628 GNDA.n3253 GNDA.n3252 0.8197
R18629 GNDA.n1514 GNDA.n1513 0.8197
R18630 GNDA.n3261 GNDA.n1510 0.8197
R18631 GNDA.n3260 GNDA.n1511 0.8197
R18632 GNDA.n3294 GNDA.n3293 0.8197
R18633 GNDA.n3280 GNDA.n1494 0.8197
R18634 GNDA.n3287 GNDA.n3281 0.8197
R18635 GNDA.n3286 GNDA.n3283 0.8197
R18636 GNDA.n3299 GNDA.n1472 0.8197
R18637 GNDA.n2726 GNDA.n2722 0.8197
R18638 GNDA.n2729 GNDA.n2728 0.8197
R18639 GNDA.n2797 GNDA.n2730 0.8197
R18640 GNDA.n5044 GNDA.n165 0.8197
R18641 GNDA.n5043 GNDA.n167 0.8197
R18642 GNDA.n218 GNDA.n200 0.8197
R18643 GNDA.n217 GNDA.n215 0.8197
R18644 GNDA.n211 GNDA.n210 0.8197
R18645 GNDA.n207 GNDA.n203 0.8197
R18646 GNDA.n206 GNDA.n187 0.8197
R18647 GNDA.n4985 GNDA.n4984 0.8197
R18648 GNDA.n1703 GNDA.n1702 0.8197
R18649 GNDA.n1699 GNDA.n1698 0.8197
R18650 GNDA.n1695 GNDA.n1679 0.8197
R18651 GNDA.n1694 GNDA.n1691 0.8197
R18652 GNDA.n1687 GNDA.n1684 0.8197
R18653 GNDA.n1681 GNDA.n1603 0.8197
R18654 GNDA.n1709 GNDA.n1708 0.8197
R18655 GNDA.n1712 GNDA.n1602 0.8197
R18656 GNDA.n4975 GNDA.n4866 0.8197
R18657 GNDA.n4972 GNDA.n4971 0.8197
R18658 GNDA.n4968 GNDA.n4869 0.8197
R18659 GNDA.n4967 GNDA.n4870 0.8197
R18660 GNDA.n4902 GNDA.n4899 0.8197
R18661 GNDA.n4903 GNDA.n4893 0.8197
R18662 GNDA.n4907 GNDA.n4906 0.8197
R18663 GNDA.n4911 GNDA.n4910 0.8197
R18664 GNDA.n5254 GNDA.n59 0.8197
R18665 GNDA.n5251 GNDA.n5250 0.8197
R18666 GNDA.n5247 GNDA.n62 0.8197
R18667 GNDA.n5246 GNDA.n63 0.8197
R18668 GNDA.n5181 GNDA.n5178 0.8197
R18669 GNDA.n5182 GNDA.n5172 0.8197
R18670 GNDA.n5186 GNDA.n5185 0.8197
R18671 GNDA.n5190 GNDA.n5189 0.8197
R18672 GNDA.n4829 GNDA.n4721 0.8197
R18673 GNDA.n4828 GNDA.n4722 0.8197
R18674 GNDA.n4748 GNDA.n4745 0.8197
R18675 GNDA.n4751 GNDA.n4750 0.8197
R18676 GNDA.n4761 GNDA.n4758 0.8197
R18677 GNDA.n4762 GNDA.n4744 0.8197
R18678 GNDA.n4766 GNDA.n4765 0.8197
R18679 GNDA.n4770 GNDA.n4769 0.8197
R18680 GNDA.n2909 GNDA.n2908 0.8197
R18681 GNDA.n2915 GNDA.n2667 0.8197
R18682 GNDA.n2914 GNDA.n2668 0.8197
R18683 GNDA.n2832 GNDA.n2830 0.8197
R18684 GNDA.n2841 GNDA.n2839 0.8197
R18685 GNDA.n2840 GNDA.n2688 0.8197
R18686 GNDA.n2850 GNDA.n2849 0.8197
R18687 GNDA.n2690 GNDA.n2686 0.8197
R18688 GNDA.n5264 GNDA.n5263 0.8197
R18689 GNDA.n32 GNDA.n23 0.8197
R18690 GNDA.n39 GNDA.n33 0.8197
R18691 GNDA.n38 GNDA.n35 0.8197
R18692 GNDA.n5269 GNDA.n1 0.8197
R18693 GNDA.n5101 GNDA.n5098 0.8197
R18694 GNDA.n5104 GNDA.n5103 0.8197
R18695 GNDA.n5108 GNDA.n5107 0.8197
R18696 GNDA.n462 GNDA.n461 0.786958
R18697 GNDA.n3547 GNDA.n3545 0.786958
R18698 GNDA.n743 GNDA.n586 0.78175
R18699 GNDA.n4617 GNDA.n433 0.78175
R18700 GNDA.n2813 GNDA.n2812 0.776542
R18701 GNDA.n3698 GNDA.n3697 0.776542
R18702 GNDA.n4574 GNDA.n4573 0.776542
R18703 GNDA.n4437 GNDA.n494 0.776542
R18704 GNDA.n4355 GNDA.n489 0.776542
R18705 GNDA.n4273 GNDA.n484 0.776542
R18706 GNDA.n4191 GNDA.n479 0.776542
R18707 GNDA.n4109 GNDA.n443 0.776542
R18708 GNDA.n4027 GNDA.n438 0.776542
R18709 GNDA.n3845 GNDA.n3844 0.776542
R18710 GNDA.n3708 GNDA.n3707 0.776542
R18711 GNDA.n1445 GNDA.n1443 0.776542
R18712 GNDA.n1307 GNDA.n770 0.776542
R18713 GNDA.n1225 GNDA.n765 0.776542
R18714 GNDA.n1143 GNDA.n760 0.776542
R18715 GNDA.n1061 GNDA.n755 0.776542
R18716 GNDA.n979 GNDA.n750 0.776542
R18717 GNDA.n3399 GNDA.n3398 0.776542
R18718 GNDA.n3525 GNDA.n3524 0.776542
R18719 GNDA.n2260 GNDA.n2258 0.776542
R18720 GNDA.n2288 GNDA.n2287 0.776542
R18721 GNDA.n736 GNDA.n735 0.776542
R18722 GNDA.n3945 GNDA.n3944 0.77295
R18723 GNDA.n887 GNDA.n886 0.77295
R18724 GNDA.n3935 GNDA.n3934 0.755708
R18725 GNDA.n897 GNDA.n896 0.755708
R18726 GNDA.n3935 GNDA.n3853 0.751
R18727 GNDA.n896 GNDA.n747 0.751
R18728 GNDA.n3538 GNDA.n603 0.729667
R18729 GNDA.n3577 GNDA.n586 0.729667
R18730 GNDA.n3578 GNDA.n433 0.729667
R18731 GNDA.n4616 GNDA.n434 0.729667
R18732 GNDA.n2640 GNDA.n2470 0.723198
R18733 GNDA.n3319 GNDA.n3318 0.718281
R18734 GNDA.n3337 GNDA.n3336 0.688
R18735 GNDA.n3606 GNDA.n574 0.688
R18736 GNDA.n743 GNDA.n603 0.688
R18737 GNDA.n4617 GNDA.n4616 0.688
R18738 GNDA.n2344 GNDA.n2343 0.675611
R18739 GNDA.n3234 GNDA.n1524 0.65675
R18740 GNDA.n3120 GNDA 0.5637
R18741 GNDA.n3282 GNDA 0.5637
R18742 GNDA.n214 GNDA 0.5637
R18743 GNDA GNDA.n1680 0.5637
R18744 GNDA GNDA.n4894 0.5637
R18745 GNDA GNDA.n5173 0.5637
R18746 GNDA.n4755 GNDA 0.5637
R18747 GNDA.n2834 GNDA 0.5637
R18748 GNDA.n34 GNDA 0.5637
R18749 GNDA.n3346 GNDA.n3344 0.563
R18750 GNDA.n3348 GNDA.n3346 0.563
R18751 GNDA.n3350 GNDA.n3348 0.563
R18752 GNDA.n3352 GNDA.n3350 0.563
R18753 GNDA.n3354 GNDA.n3352 0.563
R18754 GNDA.n3356 GNDA.n3354 0.563
R18755 GNDA.n3358 GNDA.n3356 0.563
R18756 GNDA.n3360 GNDA.n3358 0.563
R18757 GNDA.n3362 GNDA.n3360 0.563
R18758 GNDA.n3364 GNDA.n3362 0.563
R18759 GNDA.n3558 GNDA.n3557 0.464042
R18760 GNDA.t213 GNDA.t230 0.396629
R18761 GNDA.n3336 GNDA.n574 0.396333
R18762 GNDA.n4860 GNDA.n105 0.383687
R18763 GNDA.n3603 GNDA.n3599 0.34425
R18764 GNDA.n3559 GNDA.n596 0.34425
R18765 GNDA.n2628 GNDA.n2627 0.339042
R18766 GNDA.n3578 GNDA.n3577 0.313
R18767 GNDA.n3337 GNDA.n3334 0.292167
R18768 GNDA.n3606 GNDA.n3605 0.292167
R18769 GNDA.n2466 GNDA.n2433 0.286759
R18770 GNDA.n2279 GNDA.n2276 0.28175
R18771 GNDA.n2286 GNDA.n2281 0.28175
R18772 GNDA.n2265 GNDA.n2264 0.28175
R18773 GNDA.n3527 GNDA.n610 0.28175
R18774 GNDA.n894 GNDA.n893 0.28175
R18775 GNDA.n3375 GNDA.n3374 0.28175
R18776 GNDA.n3371 GNDA.n3370 0.28175
R18777 GNDA.n1458 GNDA.n1457 0.28175
R18778 GNDA.n3704 GNDA.n3702 0.28175
R18779 GNDA.n3847 GNDA.n533 0.28175
R18780 GNDA.n3941 GNDA.n3938 0.28175
R18781 GNDA.n4605 GNDA.n4604 0.28175
R18782 GNDA.n4593 GNDA.n4592 0.28175
R18783 GNDA.n4589 GNDA.n4588 0.28175
R18784 GNDA.n4585 GNDA.n4584 0.28175
R18785 GNDA.n4581 GNDA.n4580 0.28175
R18786 GNDA.n3387 GNDA.n3386 0.271333
R18787 GNDA GNDA.n3119 0.2565
R18788 GNDA.n3300 GNDA 0.2565
R18789 GNDA.n202 GNDA 0.2565
R18790 GNDA.n1688 GNDA 0.2565
R18791 GNDA.n4897 GNDA 0.2565
R18792 GNDA.n5176 GNDA 0.2565
R18793 GNDA GNDA.n4754 0.2565
R18794 GNDA GNDA.n2833 0.2565
R18795 GNDA GNDA.n0 0.2565
R18796 GNDA.n2430 GNDA.n2378 0.229919
R18797 GNDA.n3366 GNDA.n1461 0.224458
R18798 GNDA.n3700 GNDA.n3615 0.21925
R18799 GNDA.n3581 GNDA.n3580 0.208833
R18800 GNDA.n3576 GNDA.n3574 0.208833
R18801 GNDA.n3391 GNDA.n3390 0.198417
R18802 GNDA.n3379 GNDA.n3378 0.198417
R18803 GNDA.n1453 GNDA.n1449 0.198417
R18804 GNDA.n3852 GNDA.n3849 0.198417
R18805 GNDA.n2713 GNDA.n2712 0.188
R18806 GNDA.n2810 GNDA.n2809 0.188
R18807 GNDA.n4609 GNDA.n4608 0.188
R18808 GNDA.n3594 GNDA.n3593 0.172375
R18809 GNDA.n3563 GNDA.n3562 0.172375
R18810 GNDA.n3274 GNDA.n1498 0.15675
R18811 GNDA.n3271 GNDA.n3270 0.15675
R18812 GNDA.n2928 GNDA.n2927 0.151542
R18813 GNDA.n3231 GNDA.n3227 0.147453
R18814 GNDA.n2581 GNDA.n2577 0.146333
R18815 GNDA.n2585 GNDA.n2577 0.146333
R18816 GNDA.n2586 GNDA.n2585 0.146333
R18817 GNDA.n2594 GNDA.n2593 0.146333
R18818 GNDA.n2597 GNDA.n2594 0.146333
R18819 GNDA.n2597 GNDA.n2569 0.146333
R18820 GNDA.n2605 GNDA.n2565 0.146333
R18821 GNDA.n2609 GNDA.n2565 0.146333
R18822 GNDA.n2610 GNDA.n2609 0.146333
R18823 GNDA.n2618 GNDA.n2617 0.146333
R18824 GNDA.n2621 GNDA.n2618 0.146333
R18825 GNDA.n2621 GNDA.n2559 0.146333
R18826 GNDA.n3619 GNDA.n3618 0.146333
R18827 GNDA.n3620 GNDA.n3619 0.146333
R18828 GNDA.n3621 GNDA.n3620 0.146333
R18829 GNDA.n3625 GNDA.n3624 0.146333
R18830 GNDA.n3626 GNDA.n3625 0.146333
R18831 GNDA.n3627 GNDA.n3626 0.146333
R18832 GNDA.n3631 GNDA.n3630 0.146333
R18833 GNDA.n3632 GNDA.n3631 0.146333
R18834 GNDA.n3633 GNDA.n3632 0.146333
R18835 GNDA.n3637 GNDA.n3636 0.146333
R18836 GNDA.n3638 GNDA.n3637 0.146333
R18837 GNDA.n3639 GNDA.n3638 0.146333
R18838 GNDA.n4517 GNDA.n500 0.146333
R18839 GNDA.n4522 GNDA.n4517 0.146333
R18840 GNDA.n4523 GNDA.n4522 0.146333
R18841 GNDA.n4533 GNDA.n4532 0.146333
R18842 GNDA.n4536 GNDA.n4533 0.146333
R18843 GNDA.n4536 GNDA.n4513 0.146333
R18844 GNDA.n4546 GNDA.n4511 0.146333
R18845 GNDA.n4552 GNDA.n4511 0.146333
R18846 GNDA.n4553 GNDA.n4552 0.146333
R18847 GNDA.n4563 GNDA.n4562 0.146333
R18848 GNDA.n4566 GNDA.n4563 0.146333
R18849 GNDA.n4566 GNDA.n4507 0.146333
R18850 GNDA.n4440 GNDA.n4436 0.146333
R18851 GNDA.n4446 GNDA.n4436 0.146333
R18852 GNDA.n4447 GNDA.n4446 0.146333
R18853 GNDA.n4457 GNDA.n4456 0.146333
R18854 GNDA.n4460 GNDA.n4457 0.146333
R18855 GNDA.n4460 GNDA.n4432 0.146333
R18856 GNDA.n4470 GNDA.n4430 0.146333
R18857 GNDA.n4476 GNDA.n4430 0.146333
R18858 GNDA.n4477 GNDA.n4476 0.146333
R18859 GNDA.n4487 GNDA.n4486 0.146333
R18860 GNDA.n4490 GNDA.n4487 0.146333
R18861 GNDA.n4490 GNDA.n4426 0.146333
R18862 GNDA.n4358 GNDA.n4354 0.146333
R18863 GNDA.n4364 GNDA.n4354 0.146333
R18864 GNDA.n4365 GNDA.n4364 0.146333
R18865 GNDA.n4375 GNDA.n4374 0.146333
R18866 GNDA.n4378 GNDA.n4375 0.146333
R18867 GNDA.n4378 GNDA.n4350 0.146333
R18868 GNDA.n4388 GNDA.n4348 0.146333
R18869 GNDA.n4394 GNDA.n4348 0.146333
R18870 GNDA.n4395 GNDA.n4394 0.146333
R18871 GNDA.n4405 GNDA.n4404 0.146333
R18872 GNDA.n4408 GNDA.n4405 0.146333
R18873 GNDA.n4408 GNDA.n4344 0.146333
R18874 GNDA.n4276 GNDA.n4272 0.146333
R18875 GNDA.n4282 GNDA.n4272 0.146333
R18876 GNDA.n4283 GNDA.n4282 0.146333
R18877 GNDA.n4293 GNDA.n4292 0.146333
R18878 GNDA.n4296 GNDA.n4293 0.146333
R18879 GNDA.n4296 GNDA.n4268 0.146333
R18880 GNDA.n4306 GNDA.n4266 0.146333
R18881 GNDA.n4312 GNDA.n4266 0.146333
R18882 GNDA.n4313 GNDA.n4312 0.146333
R18883 GNDA.n4323 GNDA.n4322 0.146333
R18884 GNDA.n4326 GNDA.n4323 0.146333
R18885 GNDA.n4326 GNDA.n4262 0.146333
R18886 GNDA.n4194 GNDA.n4190 0.146333
R18887 GNDA.n4200 GNDA.n4190 0.146333
R18888 GNDA.n4201 GNDA.n4200 0.146333
R18889 GNDA.n4211 GNDA.n4210 0.146333
R18890 GNDA.n4214 GNDA.n4211 0.146333
R18891 GNDA.n4214 GNDA.n4186 0.146333
R18892 GNDA.n4224 GNDA.n4184 0.146333
R18893 GNDA.n4230 GNDA.n4184 0.146333
R18894 GNDA.n4231 GNDA.n4230 0.146333
R18895 GNDA.n4241 GNDA.n4240 0.146333
R18896 GNDA.n4244 GNDA.n4241 0.146333
R18897 GNDA.n4244 GNDA.n4180 0.146333
R18898 GNDA.n3948 GNDA.n526 0.146333
R18899 GNDA.n3954 GNDA.n526 0.146333
R18900 GNDA.n3955 GNDA.n3954 0.146333
R18901 GNDA.n3965 GNDA.n3964 0.146333
R18902 GNDA.n3968 GNDA.n3965 0.146333
R18903 GNDA.n3968 GNDA.n522 0.146333
R18904 GNDA.n3978 GNDA.n520 0.146333
R18905 GNDA.n3984 GNDA.n520 0.146333
R18906 GNDA.n3985 GNDA.n3984 0.146333
R18907 GNDA.n3995 GNDA.n3994 0.146333
R18908 GNDA.n3998 GNDA.n3995 0.146333
R18909 GNDA.n3998 GNDA.n516 0.146333
R18910 GNDA.n4112 GNDA.n4108 0.146333
R18911 GNDA.n4118 GNDA.n4108 0.146333
R18912 GNDA.n4119 GNDA.n4118 0.146333
R18913 GNDA.n4129 GNDA.n4128 0.146333
R18914 GNDA.n4132 GNDA.n4129 0.146333
R18915 GNDA.n4132 GNDA.n4104 0.146333
R18916 GNDA.n4142 GNDA.n4102 0.146333
R18917 GNDA.n4148 GNDA.n4102 0.146333
R18918 GNDA.n4149 GNDA.n4148 0.146333
R18919 GNDA.n4159 GNDA.n4158 0.146333
R18920 GNDA.n4162 GNDA.n4159 0.146333
R18921 GNDA.n4162 GNDA.n4098 0.146333
R18922 GNDA.n4030 GNDA.n4026 0.146333
R18923 GNDA.n4036 GNDA.n4026 0.146333
R18924 GNDA.n4037 GNDA.n4036 0.146333
R18925 GNDA.n4047 GNDA.n4046 0.146333
R18926 GNDA.n4050 GNDA.n4047 0.146333
R18927 GNDA.n4050 GNDA.n4022 0.146333
R18928 GNDA.n4060 GNDA.n4020 0.146333
R18929 GNDA.n4066 GNDA.n4020 0.146333
R18930 GNDA.n4067 GNDA.n4066 0.146333
R18931 GNDA.n4077 GNDA.n4076 0.146333
R18932 GNDA.n4080 GNDA.n4077 0.146333
R18933 GNDA.n4080 GNDA.n4016 0.146333
R18934 GNDA.n3856 GNDA.n3855 0.146333
R18935 GNDA.n3857 GNDA.n3856 0.146333
R18936 GNDA.n3858 GNDA.n3857 0.146333
R18937 GNDA.n3862 GNDA.n3861 0.146333
R18938 GNDA.n3863 GNDA.n3862 0.146333
R18939 GNDA.n3864 GNDA.n3863 0.146333
R18940 GNDA.n3868 GNDA.n3867 0.146333
R18941 GNDA.n3869 GNDA.n3868 0.146333
R18942 GNDA.n3870 GNDA.n3869 0.146333
R18943 GNDA.n3874 GNDA.n3873 0.146333
R18944 GNDA.n3875 GNDA.n3874 0.146333
R18945 GNDA.n3876 GNDA.n3875 0.146333
R18946 GNDA.n3788 GNDA.n536 0.146333
R18947 GNDA.n3793 GNDA.n3788 0.146333
R18948 GNDA.n3794 GNDA.n3793 0.146333
R18949 GNDA.n3804 GNDA.n3803 0.146333
R18950 GNDA.n3807 GNDA.n3804 0.146333
R18951 GNDA.n3807 GNDA.n3784 0.146333
R18952 GNDA.n3817 GNDA.n3782 0.146333
R18953 GNDA.n3823 GNDA.n3782 0.146333
R18954 GNDA.n3824 GNDA.n3823 0.146333
R18955 GNDA.n3834 GNDA.n3833 0.146333
R18956 GNDA.n3837 GNDA.n3834 0.146333
R18957 GNDA.n3837 GNDA.n3778 0.146333
R18958 GNDA.n3711 GNDA.n562 0.146333
R18959 GNDA.n3717 GNDA.n562 0.146333
R18960 GNDA.n3718 GNDA.n3717 0.146333
R18961 GNDA.n3728 GNDA.n3727 0.146333
R18962 GNDA.n3731 GNDA.n3728 0.146333
R18963 GNDA.n3731 GNDA.n558 0.146333
R18964 GNDA.n3741 GNDA.n556 0.146333
R18965 GNDA.n3747 GNDA.n556 0.146333
R18966 GNDA.n3748 GNDA.n3747 0.146333
R18967 GNDA.n3758 GNDA.n3757 0.146333
R18968 GNDA.n3761 GNDA.n3758 0.146333
R18969 GNDA.n3761 GNDA.n552 0.146333
R18970 GNDA.n1387 GNDA.n776 0.146333
R18971 GNDA.n1392 GNDA.n1387 0.146333
R18972 GNDA.n1393 GNDA.n1392 0.146333
R18973 GNDA.n1403 GNDA.n1402 0.146333
R18974 GNDA.n1406 GNDA.n1403 0.146333
R18975 GNDA.n1406 GNDA.n1383 0.146333
R18976 GNDA.n1416 GNDA.n1381 0.146333
R18977 GNDA.n1422 GNDA.n1381 0.146333
R18978 GNDA.n1423 GNDA.n1422 0.146333
R18979 GNDA.n1433 GNDA.n1432 0.146333
R18980 GNDA.n1436 GNDA.n1433 0.146333
R18981 GNDA.n1436 GNDA.n1377 0.146333
R18982 GNDA.n1310 GNDA.n1306 0.146333
R18983 GNDA.n1316 GNDA.n1306 0.146333
R18984 GNDA.n1317 GNDA.n1316 0.146333
R18985 GNDA.n1327 GNDA.n1326 0.146333
R18986 GNDA.n1330 GNDA.n1327 0.146333
R18987 GNDA.n1330 GNDA.n1302 0.146333
R18988 GNDA.n1340 GNDA.n1300 0.146333
R18989 GNDA.n1346 GNDA.n1300 0.146333
R18990 GNDA.n1347 GNDA.n1346 0.146333
R18991 GNDA.n1357 GNDA.n1356 0.146333
R18992 GNDA.n1360 GNDA.n1357 0.146333
R18993 GNDA.n1360 GNDA.n1296 0.146333
R18994 GNDA.n1228 GNDA.n1224 0.146333
R18995 GNDA.n1234 GNDA.n1224 0.146333
R18996 GNDA.n1235 GNDA.n1234 0.146333
R18997 GNDA.n1245 GNDA.n1244 0.146333
R18998 GNDA.n1248 GNDA.n1245 0.146333
R18999 GNDA.n1248 GNDA.n1220 0.146333
R19000 GNDA.n1258 GNDA.n1218 0.146333
R19001 GNDA.n1264 GNDA.n1218 0.146333
R19002 GNDA.n1265 GNDA.n1264 0.146333
R19003 GNDA.n1275 GNDA.n1274 0.146333
R19004 GNDA.n1278 GNDA.n1275 0.146333
R19005 GNDA.n1278 GNDA.n1214 0.146333
R19006 GNDA.n900 GNDA.n802 0.146333
R19007 GNDA.n906 GNDA.n802 0.146333
R19008 GNDA.n907 GNDA.n906 0.146333
R19009 GNDA.n917 GNDA.n916 0.146333
R19010 GNDA.n920 GNDA.n917 0.146333
R19011 GNDA.n920 GNDA.n798 0.146333
R19012 GNDA.n930 GNDA.n796 0.146333
R19013 GNDA.n936 GNDA.n796 0.146333
R19014 GNDA.n937 GNDA.n936 0.146333
R19015 GNDA.n947 GNDA.n946 0.146333
R19016 GNDA.n950 GNDA.n947 0.146333
R19017 GNDA.n950 GNDA.n792 0.146333
R19018 GNDA.n1146 GNDA.n1142 0.146333
R19019 GNDA.n1152 GNDA.n1142 0.146333
R19020 GNDA.n1153 GNDA.n1152 0.146333
R19021 GNDA.n1163 GNDA.n1162 0.146333
R19022 GNDA.n1166 GNDA.n1163 0.146333
R19023 GNDA.n1166 GNDA.n1138 0.146333
R19024 GNDA.n1176 GNDA.n1136 0.146333
R19025 GNDA.n1182 GNDA.n1136 0.146333
R19026 GNDA.n1183 GNDA.n1182 0.146333
R19027 GNDA.n1193 GNDA.n1192 0.146333
R19028 GNDA.n1196 GNDA.n1193 0.146333
R19029 GNDA.n1196 GNDA.n1132 0.146333
R19030 GNDA.n1064 GNDA.n1060 0.146333
R19031 GNDA.n1070 GNDA.n1060 0.146333
R19032 GNDA.n1071 GNDA.n1070 0.146333
R19033 GNDA.n1081 GNDA.n1080 0.146333
R19034 GNDA.n1084 GNDA.n1081 0.146333
R19035 GNDA.n1084 GNDA.n1056 0.146333
R19036 GNDA.n1094 GNDA.n1054 0.146333
R19037 GNDA.n1100 GNDA.n1054 0.146333
R19038 GNDA.n1101 GNDA.n1100 0.146333
R19039 GNDA.n1111 GNDA.n1110 0.146333
R19040 GNDA.n1114 GNDA.n1111 0.146333
R19041 GNDA.n1114 GNDA.n1050 0.146333
R19042 GNDA.n982 GNDA.n978 0.146333
R19043 GNDA.n988 GNDA.n978 0.146333
R19044 GNDA.n989 GNDA.n988 0.146333
R19045 GNDA.n999 GNDA.n998 0.146333
R19046 GNDA.n1002 GNDA.n999 0.146333
R19047 GNDA.n1002 GNDA.n974 0.146333
R19048 GNDA.n1012 GNDA.n972 0.146333
R19049 GNDA.n1018 GNDA.n972 0.146333
R19050 GNDA.n1019 GNDA.n1018 0.146333
R19051 GNDA.n1029 GNDA.n1028 0.146333
R19052 GNDA.n1032 GNDA.n1029 0.146333
R19053 GNDA.n1032 GNDA.n968 0.146333
R19054 GNDA.n808 GNDA.n807 0.146333
R19055 GNDA.n809 GNDA.n808 0.146333
R19056 GNDA.n810 GNDA.n809 0.146333
R19057 GNDA.n814 GNDA.n813 0.146333
R19058 GNDA.n815 GNDA.n814 0.146333
R19059 GNDA.n816 GNDA.n815 0.146333
R19060 GNDA.n820 GNDA.n819 0.146333
R19061 GNDA.n821 GNDA.n820 0.146333
R19062 GNDA.n822 GNDA.n821 0.146333
R19063 GNDA.n826 GNDA.n825 0.146333
R19064 GNDA.n827 GNDA.n826 0.146333
R19065 GNDA.n828 GNDA.n827 0.146333
R19066 GNDA.n657 GNDA.n656 0.146333
R19067 GNDA.n658 GNDA.n657 0.146333
R19068 GNDA.n659 GNDA.n658 0.146333
R19069 GNDA.n663 GNDA.n662 0.146333
R19070 GNDA.n664 GNDA.n663 0.146333
R19071 GNDA.n665 GNDA.n664 0.146333
R19072 GNDA.n669 GNDA.n668 0.146333
R19073 GNDA.n670 GNDA.n669 0.146333
R19074 GNDA.n671 GNDA.n670 0.146333
R19075 GNDA.n675 GNDA.n674 0.146333
R19076 GNDA.n676 GNDA.n675 0.146333
R19077 GNDA.n677 GNDA.n676 0.146333
R19078 GNDA.n3402 GNDA.n651 0.146333
R19079 GNDA.n3408 GNDA.n651 0.146333
R19080 GNDA.n3409 GNDA.n3408 0.146333
R19081 GNDA.n3419 GNDA.n3418 0.146333
R19082 GNDA.n3422 GNDA.n3419 0.146333
R19083 GNDA.n3422 GNDA.n647 0.146333
R19084 GNDA.n3432 GNDA.n645 0.146333
R19085 GNDA.n3438 GNDA.n645 0.146333
R19086 GNDA.n3439 GNDA.n3438 0.146333
R19087 GNDA.n3449 GNDA.n3448 0.146333
R19088 GNDA.n3452 GNDA.n3449 0.146333
R19089 GNDA.n3452 GNDA.n641 0.146333
R19090 GNDA.n3468 GNDA.n613 0.146333
R19091 GNDA.n3473 GNDA.n3468 0.146333
R19092 GNDA.n3474 GNDA.n3473 0.146333
R19093 GNDA.n3484 GNDA.n3483 0.146333
R19094 GNDA.n3487 GNDA.n3484 0.146333
R19095 GNDA.n3487 GNDA.n3464 0.146333
R19096 GNDA.n3497 GNDA.n3462 0.146333
R19097 GNDA.n3503 GNDA.n3462 0.146333
R19098 GNDA.n3504 GNDA.n3503 0.146333
R19099 GNDA.n3514 GNDA.n3513 0.146333
R19100 GNDA.n3517 GNDA.n3514 0.146333
R19101 GNDA.n3517 GNDA.n3458 0.146333
R19102 GNDA.n2180 GNDA.n2179 0.146333
R19103 GNDA.n2181 GNDA.n2180 0.146333
R19104 GNDA.n2182 GNDA.n2181 0.146333
R19105 GNDA.n2186 GNDA.n2185 0.146333
R19106 GNDA.n2187 GNDA.n2186 0.146333
R19107 GNDA.n2188 GNDA.n2187 0.146333
R19108 GNDA.n2192 GNDA.n2191 0.146333
R19109 GNDA.n2193 GNDA.n2192 0.146333
R19110 GNDA.n2194 GNDA.n2193 0.146333
R19111 GNDA.n2198 GNDA.n2197 0.146333
R19112 GNDA.n2199 GNDA.n2198 0.146333
R19113 GNDA.n2200 GNDA.n2199 0.146333
R19114 GNDA.n2293 GNDA.n2290 0.146333
R19115 GNDA.n2296 GNDA.n2293 0.146333
R19116 GNDA.n2296 GNDA.n2172 0.146333
R19117 GNDA.n2306 GNDA.n2170 0.146333
R19118 GNDA.n2310 GNDA.n2170 0.146333
R19119 GNDA.n2313 GNDA.n2310 0.146333
R19120 GNDA.n2323 GNDA.n2320 0.146333
R19121 GNDA.n2326 GNDA.n2323 0.146333
R19122 GNDA.n2326 GNDA.n2166 0.146333
R19123 GNDA.n2335 GNDA.n2163 0.146333
R19124 GNDA.n2340 GNDA.n2163 0.146333
R19125 GNDA.n2340 GNDA.n2164 0.146333
R19126 GNDA.n2500 GNDA.n2492 0.146333
R19127 GNDA.n2501 GNDA.n2500 0.146333
R19128 GNDA.n2511 GNDA.n2510 0.146333
R19129 GNDA.n2512 GNDA.n2511 0.146333
R19130 GNDA.n2512 GNDA.n2488 0.146333
R19131 GNDA.n2522 GNDA.n2486 0.146333
R19132 GNDA.n2530 GNDA.n2486 0.146333
R19133 GNDA.n2531 GNDA.n2530 0.146333
R19134 GNDA.n2541 GNDA.n2540 0.146333
R19135 GNDA.n2542 GNDA.n2541 0.146333
R19136 GNDA.n2542 GNDA.n1864 0.146333
R19137 GNDA.n2496 GNDA.n2495 0.146333
R19138 GNDA.n2499 GNDA.n2496 0.146333
R19139 GNDA.n2499 GNDA.n2491 0.146333
R19140 GNDA.n2509 GNDA.n2489 0.146333
R19141 GNDA.n2515 GNDA.n2489 0.146333
R19142 GNDA.n2516 GNDA.n2515 0.146333
R19143 GNDA.n2526 GNDA.n2525 0.146333
R19144 GNDA.n2529 GNDA.n2526 0.146333
R19145 GNDA.n2529 GNDA.n2485 0.146333
R19146 GNDA.n2539 GNDA.n2483 0.146333
R19147 GNDA.n2543 GNDA.n2483 0.146333
R19148 GNDA.n2543 GNDA.n1865 0.146333
R19149 GNDA.n2589 GNDA.n2586 0.135917
R19150 GNDA.n2593 GNDA.n2573 0.135917
R19151 GNDA.n2601 GNDA.n2569 0.135917
R19152 GNDA.n2605 GNDA.n2602 0.135917
R19153 GNDA.n2613 GNDA.n2610 0.135917
R19154 GNDA.n2617 GNDA.n2561 0.135917
R19155 GNDA.n2637 GNDA.n2559 0.135917
R19156 GNDA.n3696 GNDA.n3618 0.135917
R19157 GNDA.n3622 GNDA.n3621 0.135917
R19158 GNDA.n3624 GNDA.n3623 0.135917
R19159 GNDA.n3628 GNDA.n3627 0.135917
R19160 GNDA.n3630 GNDA.n3629 0.135917
R19161 GNDA.n3634 GNDA.n3633 0.135917
R19162 GNDA.n3636 GNDA.n3635 0.135917
R19163 GNDA.n4572 GNDA.n500 0.135917
R19164 GNDA.n4526 GNDA.n4523 0.135917
R19165 GNDA.n4532 GNDA.n4515 0.135917
R19166 GNDA.n4542 GNDA.n4513 0.135917
R19167 GNDA.n4546 GNDA.n4543 0.135917
R19168 GNDA.n4556 GNDA.n4553 0.135917
R19169 GNDA.n4562 GNDA.n4509 0.135917
R19170 GNDA.n4440 GNDA.n4438 0.135917
R19171 GNDA.n4450 GNDA.n4447 0.135917
R19172 GNDA.n4456 GNDA.n4434 0.135917
R19173 GNDA.n4466 GNDA.n4432 0.135917
R19174 GNDA.n4470 GNDA.n4467 0.135917
R19175 GNDA.n4480 GNDA.n4477 0.135917
R19176 GNDA.n4486 GNDA.n4428 0.135917
R19177 GNDA.n4358 GNDA.n4356 0.135917
R19178 GNDA.n4368 GNDA.n4365 0.135917
R19179 GNDA.n4374 GNDA.n4352 0.135917
R19180 GNDA.n4384 GNDA.n4350 0.135917
R19181 GNDA.n4388 GNDA.n4385 0.135917
R19182 GNDA.n4398 GNDA.n4395 0.135917
R19183 GNDA.n4404 GNDA.n4346 0.135917
R19184 GNDA.n4276 GNDA.n4274 0.135917
R19185 GNDA.n4286 GNDA.n4283 0.135917
R19186 GNDA.n4292 GNDA.n4270 0.135917
R19187 GNDA.n4302 GNDA.n4268 0.135917
R19188 GNDA.n4306 GNDA.n4303 0.135917
R19189 GNDA.n4316 GNDA.n4313 0.135917
R19190 GNDA.n4322 GNDA.n4264 0.135917
R19191 GNDA.n4194 GNDA.n4192 0.135917
R19192 GNDA.n4204 GNDA.n4201 0.135917
R19193 GNDA.n4210 GNDA.n4188 0.135917
R19194 GNDA.n4220 GNDA.n4186 0.135917
R19195 GNDA.n4224 GNDA.n4221 0.135917
R19196 GNDA.n4234 GNDA.n4231 0.135917
R19197 GNDA.n4240 GNDA.n4182 0.135917
R19198 GNDA.n3948 GNDA.n3946 0.135917
R19199 GNDA.n3958 GNDA.n3955 0.135917
R19200 GNDA.n3964 GNDA.n524 0.135917
R19201 GNDA.n3974 GNDA.n522 0.135917
R19202 GNDA.n3978 GNDA.n3975 0.135917
R19203 GNDA.n3988 GNDA.n3985 0.135917
R19204 GNDA.n3994 GNDA.n518 0.135917
R19205 GNDA.n4112 GNDA.n4110 0.135917
R19206 GNDA.n4122 GNDA.n4119 0.135917
R19207 GNDA.n4128 GNDA.n4106 0.135917
R19208 GNDA.n4138 GNDA.n4104 0.135917
R19209 GNDA.n4142 GNDA.n4139 0.135917
R19210 GNDA.n4152 GNDA.n4149 0.135917
R19211 GNDA.n4158 GNDA.n4100 0.135917
R19212 GNDA.n4030 GNDA.n4028 0.135917
R19213 GNDA.n4040 GNDA.n4037 0.135917
R19214 GNDA.n4046 GNDA.n4024 0.135917
R19215 GNDA.n4056 GNDA.n4022 0.135917
R19216 GNDA.n4060 GNDA.n4057 0.135917
R19217 GNDA.n4070 GNDA.n4067 0.135917
R19218 GNDA.n4076 GNDA.n4018 0.135917
R19219 GNDA.n3933 GNDA.n3855 0.135917
R19220 GNDA.n3859 GNDA.n3858 0.135917
R19221 GNDA.n3861 GNDA.n3860 0.135917
R19222 GNDA.n3865 GNDA.n3864 0.135917
R19223 GNDA.n3867 GNDA.n3866 0.135917
R19224 GNDA.n3871 GNDA.n3870 0.135917
R19225 GNDA.n3873 GNDA.n3872 0.135917
R19226 GNDA.n3843 GNDA.n536 0.135917
R19227 GNDA.n3797 GNDA.n3794 0.135917
R19228 GNDA.n3803 GNDA.n3786 0.135917
R19229 GNDA.n3813 GNDA.n3784 0.135917
R19230 GNDA.n3817 GNDA.n3814 0.135917
R19231 GNDA.n3827 GNDA.n3824 0.135917
R19232 GNDA.n3833 GNDA.n3780 0.135917
R19233 GNDA.n3711 GNDA.n3709 0.135917
R19234 GNDA.n3721 GNDA.n3718 0.135917
R19235 GNDA.n3727 GNDA.n560 0.135917
R19236 GNDA.n3737 GNDA.n558 0.135917
R19237 GNDA.n3741 GNDA.n3738 0.135917
R19238 GNDA.n3751 GNDA.n3748 0.135917
R19239 GNDA.n3757 GNDA.n554 0.135917
R19240 GNDA.n1442 GNDA.n776 0.135917
R19241 GNDA.n1396 GNDA.n1393 0.135917
R19242 GNDA.n1402 GNDA.n1385 0.135917
R19243 GNDA.n1412 GNDA.n1383 0.135917
R19244 GNDA.n1416 GNDA.n1413 0.135917
R19245 GNDA.n1426 GNDA.n1423 0.135917
R19246 GNDA.n1432 GNDA.n1379 0.135917
R19247 GNDA.n1310 GNDA.n1308 0.135917
R19248 GNDA.n1320 GNDA.n1317 0.135917
R19249 GNDA.n1326 GNDA.n1304 0.135917
R19250 GNDA.n1336 GNDA.n1302 0.135917
R19251 GNDA.n1340 GNDA.n1337 0.135917
R19252 GNDA.n1350 GNDA.n1347 0.135917
R19253 GNDA.n1356 GNDA.n1298 0.135917
R19254 GNDA.n1228 GNDA.n1226 0.135917
R19255 GNDA.n1238 GNDA.n1235 0.135917
R19256 GNDA.n1244 GNDA.n1222 0.135917
R19257 GNDA.n1254 GNDA.n1220 0.135917
R19258 GNDA.n1258 GNDA.n1255 0.135917
R19259 GNDA.n1268 GNDA.n1265 0.135917
R19260 GNDA.n1274 GNDA.n1216 0.135917
R19261 GNDA.n900 GNDA.n898 0.135917
R19262 GNDA.n910 GNDA.n907 0.135917
R19263 GNDA.n916 GNDA.n800 0.135917
R19264 GNDA.n926 GNDA.n798 0.135917
R19265 GNDA.n930 GNDA.n927 0.135917
R19266 GNDA.n940 GNDA.n937 0.135917
R19267 GNDA.n946 GNDA.n794 0.135917
R19268 GNDA.n1146 GNDA.n1144 0.135917
R19269 GNDA.n1156 GNDA.n1153 0.135917
R19270 GNDA.n1162 GNDA.n1140 0.135917
R19271 GNDA.n1172 GNDA.n1138 0.135917
R19272 GNDA.n1176 GNDA.n1173 0.135917
R19273 GNDA.n1186 GNDA.n1183 0.135917
R19274 GNDA.n1192 GNDA.n1134 0.135917
R19275 GNDA.n1064 GNDA.n1062 0.135917
R19276 GNDA.n1074 GNDA.n1071 0.135917
R19277 GNDA.n1080 GNDA.n1058 0.135917
R19278 GNDA.n1090 GNDA.n1056 0.135917
R19279 GNDA.n1094 GNDA.n1091 0.135917
R19280 GNDA.n1104 GNDA.n1101 0.135917
R19281 GNDA.n1110 GNDA.n1052 0.135917
R19282 GNDA.n982 GNDA.n980 0.135917
R19283 GNDA.n992 GNDA.n989 0.135917
R19284 GNDA.n998 GNDA.n976 0.135917
R19285 GNDA.n1008 GNDA.n974 0.135917
R19286 GNDA.n1012 GNDA.n1009 0.135917
R19287 GNDA.n1022 GNDA.n1019 0.135917
R19288 GNDA.n1028 GNDA.n970 0.135917
R19289 GNDA.n885 GNDA.n807 0.135917
R19290 GNDA.n811 GNDA.n810 0.135917
R19291 GNDA.n813 GNDA.n812 0.135917
R19292 GNDA.n817 GNDA.n816 0.135917
R19293 GNDA.n819 GNDA.n818 0.135917
R19294 GNDA.n823 GNDA.n822 0.135917
R19295 GNDA.n825 GNDA.n824 0.135917
R19296 GNDA.n734 GNDA.n656 0.135917
R19297 GNDA.n660 GNDA.n659 0.135917
R19298 GNDA.n662 GNDA.n661 0.135917
R19299 GNDA.n666 GNDA.n665 0.135917
R19300 GNDA.n668 GNDA.n667 0.135917
R19301 GNDA.n672 GNDA.n671 0.135917
R19302 GNDA.n674 GNDA.n673 0.135917
R19303 GNDA.n3402 GNDA.n3400 0.135917
R19304 GNDA.n3412 GNDA.n3409 0.135917
R19305 GNDA.n3418 GNDA.n649 0.135917
R19306 GNDA.n3428 GNDA.n647 0.135917
R19307 GNDA.n3432 GNDA.n3429 0.135917
R19308 GNDA.n3442 GNDA.n3439 0.135917
R19309 GNDA.n3448 GNDA.n643 0.135917
R19310 GNDA.n3523 GNDA.n613 0.135917
R19311 GNDA.n3477 GNDA.n3474 0.135917
R19312 GNDA.n3483 GNDA.n3466 0.135917
R19313 GNDA.n3493 GNDA.n3464 0.135917
R19314 GNDA.n3497 GNDA.n3494 0.135917
R19315 GNDA.n3507 GNDA.n3504 0.135917
R19316 GNDA.n3513 GNDA.n3460 0.135917
R19317 GNDA.n2257 GNDA.n2179 0.135917
R19318 GNDA.n2183 GNDA.n2182 0.135917
R19319 GNDA.n2185 GNDA.n2184 0.135917
R19320 GNDA.n2189 GNDA.n2188 0.135917
R19321 GNDA.n2191 GNDA.n2190 0.135917
R19322 GNDA.n2195 GNDA.n2194 0.135917
R19323 GNDA.n2197 GNDA.n2196 0.135917
R19324 GNDA.n2290 GNDA.n2174 0.135917
R19325 GNDA.n2300 GNDA.n2172 0.135917
R19326 GNDA.n2306 GNDA.n2303 0.135917
R19327 GNDA.n2316 GNDA.n2313 0.135917
R19328 GNDA.n2320 GNDA.n2168 0.135917
R19329 GNDA.n2330 GNDA.n2166 0.135917
R19330 GNDA.n2335 GNDA.n2333 0.135917
R19331 GNDA.n2502 GNDA.n2501 0.135917
R19332 GNDA.n2510 GNDA.n2490 0.135917
R19333 GNDA.n2520 GNDA.n2488 0.135917
R19334 GNDA.n2522 GNDA.n2521 0.135917
R19335 GNDA.n2532 GNDA.n2531 0.135917
R19336 GNDA.n2540 GNDA.n2484 0.135917
R19337 GNDA.n2643 GNDA.n1864 0.135917
R19338 GNDA.n2505 GNDA.n2491 0.135917
R19339 GNDA.n2509 GNDA.n2506 0.135917
R19340 GNDA.n2519 GNDA.n2516 0.135917
R19341 GNDA.n2525 GNDA.n2487 0.135917
R19342 GNDA.n2535 GNDA.n2485 0.135917
R19343 GNDA.n2539 GNDA.n2536 0.135917
R19344 GNDA.n2642 GNDA.n1865 0.135917
R19345 GNDA.n2640 GNDA.n2639 0.135331
R19346 GNDA.n2808 GNDA.n2717 0.1255
R19347 GNDA.n2711 GNDA.n2704 0.1255
R19348 GNDA.n2589 GNDA.n2573 0.1255
R19349 GNDA.n2602 GNDA.n2601 0.1255
R19350 GNDA.n2613 GNDA.n2561 0.1255
R19351 GNDA.n359 GNDA.n358 0.1255
R19352 GNDA.n3623 GNDA.n3622 0.1255
R19353 GNDA.n3629 GNDA.n3628 0.1255
R19354 GNDA.n3635 GNDA.n3634 0.1255
R19355 GNDA.n4526 GNDA.n4515 0.1255
R19356 GNDA.n4543 GNDA.n4542 0.1255
R19357 GNDA.n4556 GNDA.n4509 0.1255
R19358 GNDA.n4450 GNDA.n4434 0.1255
R19359 GNDA.n4467 GNDA.n4466 0.1255
R19360 GNDA.n4480 GNDA.n4428 0.1255
R19361 GNDA.n4368 GNDA.n4352 0.1255
R19362 GNDA.n4385 GNDA.n4384 0.1255
R19363 GNDA.n4398 GNDA.n4346 0.1255
R19364 GNDA.n4286 GNDA.n4270 0.1255
R19365 GNDA.n4303 GNDA.n4302 0.1255
R19366 GNDA.n4316 GNDA.n4264 0.1255
R19367 GNDA.n4204 GNDA.n4188 0.1255
R19368 GNDA.n4221 GNDA.n4220 0.1255
R19369 GNDA.n4234 GNDA.n4182 0.1255
R19370 GNDA.n3958 GNDA.n524 0.1255
R19371 GNDA.n3975 GNDA.n3974 0.1255
R19372 GNDA.n3988 GNDA.n518 0.1255
R19373 GNDA.n4122 GNDA.n4106 0.1255
R19374 GNDA.n4139 GNDA.n4138 0.1255
R19375 GNDA.n4152 GNDA.n4100 0.1255
R19376 GNDA.n4040 GNDA.n4024 0.1255
R19377 GNDA.n4057 GNDA.n4056 0.1255
R19378 GNDA.n4070 GNDA.n4018 0.1255
R19379 GNDA.n3860 GNDA.n3859 0.1255
R19380 GNDA.n3866 GNDA.n3865 0.1255
R19381 GNDA.n3872 GNDA.n3871 0.1255
R19382 GNDA.n3797 GNDA.n3786 0.1255
R19383 GNDA.n3814 GNDA.n3813 0.1255
R19384 GNDA.n3827 GNDA.n3780 0.1255
R19385 GNDA.n3721 GNDA.n560 0.1255
R19386 GNDA.n3738 GNDA.n3737 0.1255
R19387 GNDA.n3751 GNDA.n554 0.1255
R19388 GNDA.n1396 GNDA.n1385 0.1255
R19389 GNDA.n1413 GNDA.n1412 0.1255
R19390 GNDA.n1426 GNDA.n1379 0.1255
R19391 GNDA.n1320 GNDA.n1304 0.1255
R19392 GNDA.n1337 GNDA.n1336 0.1255
R19393 GNDA.n1350 GNDA.n1298 0.1255
R19394 GNDA.n1238 GNDA.n1222 0.1255
R19395 GNDA.n1255 GNDA.n1254 0.1255
R19396 GNDA.n1268 GNDA.n1216 0.1255
R19397 GNDA.n910 GNDA.n800 0.1255
R19398 GNDA.n927 GNDA.n926 0.1255
R19399 GNDA.n940 GNDA.n794 0.1255
R19400 GNDA.n1156 GNDA.n1140 0.1255
R19401 GNDA.n1173 GNDA.n1172 0.1255
R19402 GNDA.n1186 GNDA.n1134 0.1255
R19403 GNDA.n1074 GNDA.n1058 0.1255
R19404 GNDA.n1091 GNDA.n1090 0.1255
R19405 GNDA.n1104 GNDA.n1052 0.1255
R19406 GNDA.n992 GNDA.n976 0.1255
R19407 GNDA.n1009 GNDA.n1008 0.1255
R19408 GNDA.n1022 GNDA.n970 0.1255
R19409 GNDA.n812 GNDA.n811 0.1255
R19410 GNDA.n818 GNDA.n817 0.1255
R19411 GNDA.n824 GNDA.n823 0.1255
R19412 GNDA.n661 GNDA.n660 0.1255
R19413 GNDA.n667 GNDA.n666 0.1255
R19414 GNDA.n673 GNDA.n672 0.1255
R19415 GNDA.n3412 GNDA.n649 0.1255
R19416 GNDA.n3429 GNDA.n3428 0.1255
R19417 GNDA.n3442 GNDA.n643 0.1255
R19418 GNDA.n3477 GNDA.n3466 0.1255
R19419 GNDA.n3494 GNDA.n3493 0.1255
R19420 GNDA.n3507 GNDA.n3460 0.1255
R19421 GNDA.n2184 GNDA.n2183 0.1255
R19422 GNDA.n2190 GNDA.n2189 0.1255
R19423 GNDA.n2196 GNDA.n2195 0.1255
R19424 GNDA.n2303 GNDA.n2300 0.1255
R19425 GNDA.n2316 GNDA.n2168 0.1255
R19426 GNDA.n2333 GNDA.n2330 0.1255
R19427 GNDA.n3395 GNDA.n606 0.1255
R19428 GNDA.n4601 GNDA.n4600 0.1255
R19429 GNDA.n2502 GNDA.n2490 0.1255
R19430 GNDA.n2521 GNDA.n2520 0.1255
R19431 GNDA.n2532 GNDA.n2484 0.1255
R19432 GNDA.n2506 GNDA.n2505 0.1255
R19433 GNDA.n2519 GNDA.n2487 0.1255
R19434 GNDA.n2536 GNDA.n2535 0.1255
R19435 GNDA.n455 GNDA.n453 0.115083
R19436 GNDA.n457 GNDA.n455 0.115083
R19437 GNDA.n459 GNDA.n457 0.115083
R19438 GNDA.n461 GNDA.n459 0.115083
R19439 GNDA.n3568 GNDA.n582 0.115083
R19440 GNDA.n3587 GNDA.n582 0.115083
R19441 GNDA.n3549 GNDA.n3547 0.115083
R19442 GNDA.n3551 GNDA.n3549 0.115083
R19443 GNDA.n3553 GNDA.n3551 0.115083
R19444 GNDA.n3555 GNDA.n3553 0.115083
R19445 GNDA.n3557 GNDA.n3555 0.115083
R19446 GNDA.n2661 GNDA.n2659 0.115083
R19447 GNDA.n2663 GNDA.n2661 0.115083
R19448 GNDA.n2927 GNDA.n2926 0.115083
R19449 GNDA.n2926 GNDA.n2925 0.115083
R19450 GNDA.n2925 GNDA.n2924 0.115083
R19451 GNDA.n2924 GNDA.n1498 0.115083
R19452 GNDA.n3274 GNDA.n3273 0.115083
R19453 GNDA.n3273 GNDA.n3272 0.115083
R19454 GNDA.n3272 GNDA.n3271 0.115083
R19455 GNDA.n3270 GNDA.n3269 0.115083
R19456 GNDA.n3269 GNDA.n3268 0.115083
R19457 GNDA.n3268 GNDA.n3267 0.115083
R19458 GNDA.n3379 GNDA.n747 0.105167
R19459 GNDA.n3853 GNDA.n3852 0.105167
R19460 GNDA.n3386 GNDA.n739 0.09425
R19461 GNDA.n4609 GNDA.n435 0.09425
R19462 GNDA.n1454 GNDA.n1453 0.0838333
R19463 GNDA.n2429 GNDA 0.0817953
R19464 GNDA.n2584 GNDA.n2583 0.0734167
R19465 GNDA.n2584 GNDA.n2576 0.0734167
R19466 GNDA.n2592 GNDA.n2572 0.0734167
R19467 GNDA.n2598 GNDA.n2572 0.0734167
R19468 GNDA.n2599 GNDA.n2598 0.0734167
R19469 GNDA.n2607 GNDA.n2606 0.0734167
R19470 GNDA.n2608 GNDA.n2607 0.0734167
R19471 GNDA.n2608 GNDA.n2564 0.0734167
R19472 GNDA.n2616 GNDA.n2560 0.0734167
R19473 GNDA.n2622 GNDA.n2560 0.0734167
R19474 GNDA.n2623 GNDA.n2622 0.0734167
R19475 GNDA.n3640 GNDA.n3617 0.0734167
R19476 GNDA.n3641 GNDA.n3640 0.0734167
R19477 GNDA.n3642 GNDA.n3641 0.0734167
R19478 GNDA.n3646 GNDA.n3645 0.0734167
R19479 GNDA.n3647 GNDA.n3646 0.0734167
R19480 GNDA.n3648 GNDA.n3647 0.0734167
R19481 GNDA.n3652 GNDA.n3651 0.0734167
R19482 GNDA.n3653 GNDA.n3652 0.0734167
R19483 GNDA.n3654 GNDA.n3653 0.0734167
R19484 GNDA.n3658 GNDA.n3657 0.0734167
R19485 GNDA.n3659 GNDA.n3658 0.0734167
R19486 GNDA.n4518 GNDA.n499 0.0734167
R19487 GNDA.n4519 GNDA.n4518 0.0734167
R19488 GNDA.n4519 GNDA.n4516 0.0734167
R19489 GNDA.n4529 GNDA.n4514 0.0734167
R19490 GNDA.n4537 GNDA.n4514 0.0734167
R19491 GNDA.n4538 GNDA.n4537 0.0734167
R19492 GNDA.n4548 GNDA.n4547 0.0734167
R19493 GNDA.n4549 GNDA.n4548 0.0734167
R19494 GNDA.n4549 GNDA.n4510 0.0734167
R19495 GNDA.n4559 GNDA.n4508 0.0734167
R19496 GNDA.n4567 GNDA.n4508 0.0734167
R19497 GNDA.n4442 GNDA.n4441 0.0734167
R19498 GNDA.n4443 GNDA.n4442 0.0734167
R19499 GNDA.n4443 GNDA.n4435 0.0734167
R19500 GNDA.n4453 GNDA.n4433 0.0734167
R19501 GNDA.n4461 GNDA.n4433 0.0734167
R19502 GNDA.n4462 GNDA.n4461 0.0734167
R19503 GNDA.n4472 GNDA.n4471 0.0734167
R19504 GNDA.n4473 GNDA.n4472 0.0734167
R19505 GNDA.n4473 GNDA.n4429 0.0734167
R19506 GNDA.n4483 GNDA.n4427 0.0734167
R19507 GNDA.n4491 GNDA.n4427 0.0734167
R19508 GNDA.n4360 GNDA.n4359 0.0734167
R19509 GNDA.n4361 GNDA.n4360 0.0734167
R19510 GNDA.n4361 GNDA.n4353 0.0734167
R19511 GNDA.n4371 GNDA.n4351 0.0734167
R19512 GNDA.n4379 GNDA.n4351 0.0734167
R19513 GNDA.n4380 GNDA.n4379 0.0734167
R19514 GNDA.n4390 GNDA.n4389 0.0734167
R19515 GNDA.n4391 GNDA.n4390 0.0734167
R19516 GNDA.n4391 GNDA.n4347 0.0734167
R19517 GNDA.n4401 GNDA.n4345 0.0734167
R19518 GNDA.n4409 GNDA.n4345 0.0734167
R19519 GNDA.n4278 GNDA.n4277 0.0734167
R19520 GNDA.n4279 GNDA.n4278 0.0734167
R19521 GNDA.n4279 GNDA.n4271 0.0734167
R19522 GNDA.n4289 GNDA.n4269 0.0734167
R19523 GNDA.n4297 GNDA.n4269 0.0734167
R19524 GNDA.n4298 GNDA.n4297 0.0734167
R19525 GNDA.n4308 GNDA.n4307 0.0734167
R19526 GNDA.n4309 GNDA.n4308 0.0734167
R19527 GNDA.n4309 GNDA.n4265 0.0734167
R19528 GNDA.n4319 GNDA.n4263 0.0734167
R19529 GNDA.n4327 GNDA.n4263 0.0734167
R19530 GNDA.n4196 GNDA.n4195 0.0734167
R19531 GNDA.n4197 GNDA.n4196 0.0734167
R19532 GNDA.n4197 GNDA.n4189 0.0734167
R19533 GNDA.n4207 GNDA.n4187 0.0734167
R19534 GNDA.n4215 GNDA.n4187 0.0734167
R19535 GNDA.n4216 GNDA.n4215 0.0734167
R19536 GNDA.n4226 GNDA.n4225 0.0734167
R19537 GNDA.n4227 GNDA.n4226 0.0734167
R19538 GNDA.n4227 GNDA.n4183 0.0734167
R19539 GNDA.n4237 GNDA.n4181 0.0734167
R19540 GNDA.n4245 GNDA.n4181 0.0734167
R19541 GNDA.n3950 GNDA.n3949 0.0734167
R19542 GNDA.n3951 GNDA.n3950 0.0734167
R19543 GNDA.n3951 GNDA.n525 0.0734167
R19544 GNDA.n3961 GNDA.n523 0.0734167
R19545 GNDA.n3969 GNDA.n523 0.0734167
R19546 GNDA.n3970 GNDA.n3969 0.0734167
R19547 GNDA.n3980 GNDA.n3979 0.0734167
R19548 GNDA.n3981 GNDA.n3980 0.0734167
R19549 GNDA.n3981 GNDA.n519 0.0734167
R19550 GNDA.n3991 GNDA.n517 0.0734167
R19551 GNDA.n3999 GNDA.n517 0.0734167
R19552 GNDA.n4114 GNDA.n4113 0.0734167
R19553 GNDA.n4115 GNDA.n4114 0.0734167
R19554 GNDA.n4115 GNDA.n4107 0.0734167
R19555 GNDA.n4125 GNDA.n4105 0.0734167
R19556 GNDA.n4133 GNDA.n4105 0.0734167
R19557 GNDA.n4134 GNDA.n4133 0.0734167
R19558 GNDA.n4144 GNDA.n4143 0.0734167
R19559 GNDA.n4145 GNDA.n4144 0.0734167
R19560 GNDA.n4145 GNDA.n4101 0.0734167
R19561 GNDA.n4155 GNDA.n4099 0.0734167
R19562 GNDA.n4163 GNDA.n4099 0.0734167
R19563 GNDA.n4032 GNDA.n4031 0.0734167
R19564 GNDA.n4033 GNDA.n4032 0.0734167
R19565 GNDA.n4033 GNDA.n4025 0.0734167
R19566 GNDA.n4043 GNDA.n4023 0.0734167
R19567 GNDA.n4051 GNDA.n4023 0.0734167
R19568 GNDA.n4052 GNDA.n4051 0.0734167
R19569 GNDA.n4062 GNDA.n4061 0.0734167
R19570 GNDA.n4063 GNDA.n4062 0.0734167
R19571 GNDA.n4063 GNDA.n4019 0.0734167
R19572 GNDA.n4073 GNDA.n4017 0.0734167
R19573 GNDA.n4081 GNDA.n4017 0.0734167
R19574 GNDA.n3877 GNDA.n3854 0.0734167
R19575 GNDA.n3878 GNDA.n3877 0.0734167
R19576 GNDA.n3879 GNDA.n3878 0.0734167
R19577 GNDA.n3883 GNDA.n3882 0.0734167
R19578 GNDA.n3884 GNDA.n3883 0.0734167
R19579 GNDA.n3885 GNDA.n3884 0.0734167
R19580 GNDA.n3889 GNDA.n3888 0.0734167
R19581 GNDA.n3890 GNDA.n3889 0.0734167
R19582 GNDA.n3891 GNDA.n3890 0.0734167
R19583 GNDA.n3895 GNDA.n3894 0.0734167
R19584 GNDA.n3896 GNDA.n3895 0.0734167
R19585 GNDA.n3789 GNDA.n535 0.0734167
R19586 GNDA.n3790 GNDA.n3789 0.0734167
R19587 GNDA.n3790 GNDA.n3787 0.0734167
R19588 GNDA.n3800 GNDA.n3785 0.0734167
R19589 GNDA.n3808 GNDA.n3785 0.0734167
R19590 GNDA.n3809 GNDA.n3808 0.0734167
R19591 GNDA.n3819 GNDA.n3818 0.0734167
R19592 GNDA.n3820 GNDA.n3819 0.0734167
R19593 GNDA.n3820 GNDA.n3781 0.0734167
R19594 GNDA.n3830 GNDA.n3779 0.0734167
R19595 GNDA.n3838 GNDA.n3779 0.0734167
R19596 GNDA.n3713 GNDA.n3712 0.0734167
R19597 GNDA.n3714 GNDA.n3713 0.0734167
R19598 GNDA.n3714 GNDA.n561 0.0734167
R19599 GNDA.n3724 GNDA.n559 0.0734167
R19600 GNDA.n3732 GNDA.n559 0.0734167
R19601 GNDA.n3733 GNDA.n3732 0.0734167
R19602 GNDA.n3743 GNDA.n3742 0.0734167
R19603 GNDA.n3744 GNDA.n3743 0.0734167
R19604 GNDA.n3744 GNDA.n555 0.0734167
R19605 GNDA.n3754 GNDA.n553 0.0734167
R19606 GNDA.n3762 GNDA.n553 0.0734167
R19607 GNDA.n1388 GNDA.n775 0.0734167
R19608 GNDA.n1389 GNDA.n1388 0.0734167
R19609 GNDA.n1389 GNDA.n1386 0.0734167
R19610 GNDA.n1399 GNDA.n1384 0.0734167
R19611 GNDA.n1407 GNDA.n1384 0.0734167
R19612 GNDA.n1408 GNDA.n1407 0.0734167
R19613 GNDA.n1418 GNDA.n1417 0.0734167
R19614 GNDA.n1419 GNDA.n1418 0.0734167
R19615 GNDA.n1419 GNDA.n1380 0.0734167
R19616 GNDA.n1429 GNDA.n1378 0.0734167
R19617 GNDA.n1437 GNDA.n1378 0.0734167
R19618 GNDA.n1312 GNDA.n1311 0.0734167
R19619 GNDA.n1313 GNDA.n1312 0.0734167
R19620 GNDA.n1313 GNDA.n1305 0.0734167
R19621 GNDA.n1323 GNDA.n1303 0.0734167
R19622 GNDA.n1331 GNDA.n1303 0.0734167
R19623 GNDA.n1332 GNDA.n1331 0.0734167
R19624 GNDA.n1342 GNDA.n1341 0.0734167
R19625 GNDA.n1343 GNDA.n1342 0.0734167
R19626 GNDA.n1343 GNDA.n1299 0.0734167
R19627 GNDA.n1353 GNDA.n1297 0.0734167
R19628 GNDA.n1361 GNDA.n1297 0.0734167
R19629 GNDA.n1230 GNDA.n1229 0.0734167
R19630 GNDA.n1231 GNDA.n1230 0.0734167
R19631 GNDA.n1231 GNDA.n1223 0.0734167
R19632 GNDA.n1241 GNDA.n1221 0.0734167
R19633 GNDA.n1249 GNDA.n1221 0.0734167
R19634 GNDA.n1250 GNDA.n1249 0.0734167
R19635 GNDA.n1260 GNDA.n1259 0.0734167
R19636 GNDA.n1261 GNDA.n1260 0.0734167
R19637 GNDA.n1261 GNDA.n1217 0.0734167
R19638 GNDA.n1271 GNDA.n1215 0.0734167
R19639 GNDA.n1279 GNDA.n1215 0.0734167
R19640 GNDA.n902 GNDA.n901 0.0734167
R19641 GNDA.n903 GNDA.n902 0.0734167
R19642 GNDA.n903 GNDA.n801 0.0734167
R19643 GNDA.n913 GNDA.n799 0.0734167
R19644 GNDA.n921 GNDA.n799 0.0734167
R19645 GNDA.n922 GNDA.n921 0.0734167
R19646 GNDA.n932 GNDA.n931 0.0734167
R19647 GNDA.n933 GNDA.n932 0.0734167
R19648 GNDA.n933 GNDA.n795 0.0734167
R19649 GNDA.n943 GNDA.n793 0.0734167
R19650 GNDA.n951 GNDA.n793 0.0734167
R19651 GNDA.n1148 GNDA.n1147 0.0734167
R19652 GNDA.n1149 GNDA.n1148 0.0734167
R19653 GNDA.n1149 GNDA.n1141 0.0734167
R19654 GNDA.n1159 GNDA.n1139 0.0734167
R19655 GNDA.n1167 GNDA.n1139 0.0734167
R19656 GNDA.n1168 GNDA.n1167 0.0734167
R19657 GNDA.n1178 GNDA.n1177 0.0734167
R19658 GNDA.n1179 GNDA.n1178 0.0734167
R19659 GNDA.n1179 GNDA.n1135 0.0734167
R19660 GNDA.n1189 GNDA.n1133 0.0734167
R19661 GNDA.n1197 GNDA.n1133 0.0734167
R19662 GNDA.n1066 GNDA.n1065 0.0734167
R19663 GNDA.n1067 GNDA.n1066 0.0734167
R19664 GNDA.n1067 GNDA.n1059 0.0734167
R19665 GNDA.n1077 GNDA.n1057 0.0734167
R19666 GNDA.n1085 GNDA.n1057 0.0734167
R19667 GNDA.n1086 GNDA.n1085 0.0734167
R19668 GNDA.n1096 GNDA.n1095 0.0734167
R19669 GNDA.n1097 GNDA.n1096 0.0734167
R19670 GNDA.n1097 GNDA.n1053 0.0734167
R19671 GNDA.n1107 GNDA.n1051 0.0734167
R19672 GNDA.n1115 GNDA.n1051 0.0734167
R19673 GNDA.n984 GNDA.n983 0.0734167
R19674 GNDA.n985 GNDA.n984 0.0734167
R19675 GNDA.n985 GNDA.n977 0.0734167
R19676 GNDA.n995 GNDA.n975 0.0734167
R19677 GNDA.n1003 GNDA.n975 0.0734167
R19678 GNDA.n1004 GNDA.n1003 0.0734167
R19679 GNDA.n1014 GNDA.n1013 0.0734167
R19680 GNDA.n1015 GNDA.n1014 0.0734167
R19681 GNDA.n1015 GNDA.n971 0.0734167
R19682 GNDA.n1025 GNDA.n969 0.0734167
R19683 GNDA.n1033 GNDA.n969 0.0734167
R19684 GNDA.n829 GNDA.n806 0.0734167
R19685 GNDA.n830 GNDA.n829 0.0734167
R19686 GNDA.n831 GNDA.n830 0.0734167
R19687 GNDA.n835 GNDA.n834 0.0734167
R19688 GNDA.n836 GNDA.n835 0.0734167
R19689 GNDA.n837 GNDA.n836 0.0734167
R19690 GNDA.n841 GNDA.n840 0.0734167
R19691 GNDA.n842 GNDA.n841 0.0734167
R19692 GNDA.n843 GNDA.n842 0.0734167
R19693 GNDA.n847 GNDA.n846 0.0734167
R19694 GNDA.n848 GNDA.n847 0.0734167
R19695 GNDA.n678 GNDA.n655 0.0734167
R19696 GNDA.n679 GNDA.n678 0.0734167
R19697 GNDA.n680 GNDA.n679 0.0734167
R19698 GNDA.n684 GNDA.n683 0.0734167
R19699 GNDA.n685 GNDA.n684 0.0734167
R19700 GNDA.n686 GNDA.n685 0.0734167
R19701 GNDA.n690 GNDA.n689 0.0734167
R19702 GNDA.n691 GNDA.n690 0.0734167
R19703 GNDA.n692 GNDA.n691 0.0734167
R19704 GNDA.n696 GNDA.n695 0.0734167
R19705 GNDA.n697 GNDA.n696 0.0734167
R19706 GNDA.n3404 GNDA.n3403 0.0734167
R19707 GNDA.n3405 GNDA.n3404 0.0734167
R19708 GNDA.n3405 GNDA.n650 0.0734167
R19709 GNDA.n3415 GNDA.n648 0.0734167
R19710 GNDA.n3423 GNDA.n648 0.0734167
R19711 GNDA.n3424 GNDA.n3423 0.0734167
R19712 GNDA.n3434 GNDA.n3433 0.0734167
R19713 GNDA.n3435 GNDA.n3434 0.0734167
R19714 GNDA.n3435 GNDA.n644 0.0734167
R19715 GNDA.n3445 GNDA.n642 0.0734167
R19716 GNDA.n3453 GNDA.n642 0.0734167
R19717 GNDA.n3469 GNDA.n612 0.0734167
R19718 GNDA.n3470 GNDA.n3469 0.0734167
R19719 GNDA.n3470 GNDA.n3467 0.0734167
R19720 GNDA.n3480 GNDA.n3465 0.0734167
R19721 GNDA.n3488 GNDA.n3465 0.0734167
R19722 GNDA.n3489 GNDA.n3488 0.0734167
R19723 GNDA.n3499 GNDA.n3498 0.0734167
R19724 GNDA.n3500 GNDA.n3499 0.0734167
R19725 GNDA.n3500 GNDA.n3461 0.0734167
R19726 GNDA.n3510 GNDA.n3459 0.0734167
R19727 GNDA.n3518 GNDA.n3459 0.0734167
R19728 GNDA.n2201 GNDA.n2178 0.0734167
R19729 GNDA.n2202 GNDA.n2201 0.0734167
R19730 GNDA.n2203 GNDA.n2202 0.0734167
R19731 GNDA.n2207 GNDA.n2206 0.0734167
R19732 GNDA.n2208 GNDA.n2207 0.0734167
R19733 GNDA.n2209 GNDA.n2208 0.0734167
R19734 GNDA.n2213 GNDA.n2212 0.0734167
R19735 GNDA.n2214 GNDA.n2213 0.0734167
R19736 GNDA.n2215 GNDA.n2214 0.0734167
R19737 GNDA.n2219 GNDA.n2218 0.0734167
R19738 GNDA.n2220 GNDA.n2219 0.0734167
R19739 GNDA.n2289 GNDA.n2173 0.0734167
R19740 GNDA.n2297 GNDA.n2173 0.0734167
R19741 GNDA.n2298 GNDA.n2297 0.0734167
R19742 GNDA.n2308 GNDA.n2307 0.0734167
R19743 GNDA.n2309 GNDA.n2308 0.0734167
R19744 GNDA.n2309 GNDA.n2169 0.0734167
R19745 GNDA.n2319 GNDA.n2167 0.0734167
R19746 GNDA.n2327 GNDA.n2167 0.0734167
R19747 GNDA.n2328 GNDA.n2327 0.0734167
R19748 GNDA.n2337 GNDA.n2336 0.0734167
R19749 GNDA.n2339 GNDA.n2337 0.0734167
R19750 GNDA.n3534 GNDA.n3529 0.0734167
R19751 GNDA.n4597 GNDA.n4596 0.0734167
R19752 GNDA.n2590 GNDA.n2576 0.0682083
R19753 GNDA.n2592 GNDA.n2591 0.0682083
R19754 GNDA.n2600 GNDA.n2599 0.0682083
R19755 GNDA.n2606 GNDA.n2568 0.0682083
R19756 GNDA.n2614 GNDA.n2564 0.0682083
R19757 GNDA.n2616 GNDA.n2615 0.0682083
R19758 GNDA.n2636 GNDA.n2623 0.0682083
R19759 GNDA.n3697 GNDA.n3617 0.0682083
R19760 GNDA.n3643 GNDA.n3642 0.0682083
R19761 GNDA.n3645 GNDA.n3644 0.0682083
R19762 GNDA.n3649 GNDA.n3648 0.0682083
R19763 GNDA.n3651 GNDA.n3650 0.0682083
R19764 GNDA.n3655 GNDA.n3654 0.0682083
R19765 GNDA.n3657 GNDA.n3656 0.0682083
R19766 GNDA.n4573 GNDA.n499 0.0682083
R19767 GNDA.n4527 GNDA.n4516 0.0682083
R19768 GNDA.n4529 GNDA.n4528 0.0682083
R19769 GNDA.n4539 GNDA.n4538 0.0682083
R19770 GNDA.n4547 GNDA.n4512 0.0682083
R19771 GNDA.n4557 GNDA.n4510 0.0682083
R19772 GNDA.n4559 GNDA.n4558 0.0682083
R19773 GNDA.n4441 GNDA.n4437 0.0682083
R19774 GNDA.n4451 GNDA.n4435 0.0682083
R19775 GNDA.n4453 GNDA.n4452 0.0682083
R19776 GNDA.n4463 GNDA.n4462 0.0682083
R19777 GNDA.n4471 GNDA.n4431 0.0682083
R19778 GNDA.n4481 GNDA.n4429 0.0682083
R19779 GNDA.n4483 GNDA.n4482 0.0682083
R19780 GNDA.n4359 GNDA.n4355 0.0682083
R19781 GNDA.n4369 GNDA.n4353 0.0682083
R19782 GNDA.n4371 GNDA.n4370 0.0682083
R19783 GNDA.n4381 GNDA.n4380 0.0682083
R19784 GNDA.n4389 GNDA.n4349 0.0682083
R19785 GNDA.n4399 GNDA.n4347 0.0682083
R19786 GNDA.n4401 GNDA.n4400 0.0682083
R19787 GNDA.n4277 GNDA.n4273 0.0682083
R19788 GNDA.n4287 GNDA.n4271 0.0682083
R19789 GNDA.n4289 GNDA.n4288 0.0682083
R19790 GNDA.n4299 GNDA.n4298 0.0682083
R19791 GNDA.n4307 GNDA.n4267 0.0682083
R19792 GNDA.n4317 GNDA.n4265 0.0682083
R19793 GNDA.n4319 GNDA.n4318 0.0682083
R19794 GNDA.n4195 GNDA.n4191 0.0682083
R19795 GNDA.n4205 GNDA.n4189 0.0682083
R19796 GNDA.n4207 GNDA.n4206 0.0682083
R19797 GNDA.n4217 GNDA.n4216 0.0682083
R19798 GNDA.n4225 GNDA.n4185 0.0682083
R19799 GNDA.n4235 GNDA.n4183 0.0682083
R19800 GNDA.n4237 GNDA.n4236 0.0682083
R19801 GNDA.n3949 GNDA.n3945 0.0682083
R19802 GNDA.n3959 GNDA.n525 0.0682083
R19803 GNDA.n3961 GNDA.n3960 0.0682083
R19804 GNDA.n3971 GNDA.n3970 0.0682083
R19805 GNDA.n3979 GNDA.n521 0.0682083
R19806 GNDA.n3989 GNDA.n519 0.0682083
R19807 GNDA.n3991 GNDA.n3990 0.0682083
R19808 GNDA.n4113 GNDA.n4109 0.0682083
R19809 GNDA.n4123 GNDA.n4107 0.0682083
R19810 GNDA.n4125 GNDA.n4124 0.0682083
R19811 GNDA.n4135 GNDA.n4134 0.0682083
R19812 GNDA.n4143 GNDA.n4103 0.0682083
R19813 GNDA.n4153 GNDA.n4101 0.0682083
R19814 GNDA.n4155 GNDA.n4154 0.0682083
R19815 GNDA.n4031 GNDA.n4027 0.0682083
R19816 GNDA.n4041 GNDA.n4025 0.0682083
R19817 GNDA.n4043 GNDA.n4042 0.0682083
R19818 GNDA.n4053 GNDA.n4052 0.0682083
R19819 GNDA.n4061 GNDA.n4021 0.0682083
R19820 GNDA.n4071 GNDA.n4019 0.0682083
R19821 GNDA.n4073 GNDA.n4072 0.0682083
R19822 GNDA.n3934 GNDA.n3854 0.0682083
R19823 GNDA.n3880 GNDA.n3879 0.0682083
R19824 GNDA.n3882 GNDA.n3881 0.0682083
R19825 GNDA.n3886 GNDA.n3885 0.0682083
R19826 GNDA.n3888 GNDA.n3887 0.0682083
R19827 GNDA.n3892 GNDA.n3891 0.0682083
R19828 GNDA.n3894 GNDA.n3893 0.0682083
R19829 GNDA.n3844 GNDA.n535 0.0682083
R19830 GNDA.n3798 GNDA.n3787 0.0682083
R19831 GNDA.n3800 GNDA.n3799 0.0682083
R19832 GNDA.n3810 GNDA.n3809 0.0682083
R19833 GNDA.n3818 GNDA.n3783 0.0682083
R19834 GNDA.n3828 GNDA.n3781 0.0682083
R19835 GNDA.n3830 GNDA.n3829 0.0682083
R19836 GNDA.n3712 GNDA.n3708 0.0682083
R19837 GNDA.n3722 GNDA.n561 0.0682083
R19838 GNDA.n3724 GNDA.n3723 0.0682083
R19839 GNDA.n3734 GNDA.n3733 0.0682083
R19840 GNDA.n3742 GNDA.n557 0.0682083
R19841 GNDA.n3752 GNDA.n555 0.0682083
R19842 GNDA.n3754 GNDA.n3753 0.0682083
R19843 GNDA.n1443 GNDA.n775 0.0682083
R19844 GNDA.n1397 GNDA.n1386 0.0682083
R19845 GNDA.n1399 GNDA.n1398 0.0682083
R19846 GNDA.n1409 GNDA.n1408 0.0682083
R19847 GNDA.n1417 GNDA.n1382 0.0682083
R19848 GNDA.n1427 GNDA.n1380 0.0682083
R19849 GNDA.n1429 GNDA.n1428 0.0682083
R19850 GNDA.n1311 GNDA.n1307 0.0682083
R19851 GNDA.n1321 GNDA.n1305 0.0682083
R19852 GNDA.n1323 GNDA.n1322 0.0682083
R19853 GNDA.n1333 GNDA.n1332 0.0682083
R19854 GNDA.n1341 GNDA.n1301 0.0682083
R19855 GNDA.n1351 GNDA.n1299 0.0682083
R19856 GNDA.n1353 GNDA.n1352 0.0682083
R19857 GNDA.n1229 GNDA.n1225 0.0682083
R19858 GNDA.n1239 GNDA.n1223 0.0682083
R19859 GNDA.n1241 GNDA.n1240 0.0682083
R19860 GNDA.n1251 GNDA.n1250 0.0682083
R19861 GNDA.n1259 GNDA.n1219 0.0682083
R19862 GNDA.n1269 GNDA.n1217 0.0682083
R19863 GNDA.n1271 GNDA.n1270 0.0682083
R19864 GNDA.n901 GNDA.n897 0.0682083
R19865 GNDA.n911 GNDA.n801 0.0682083
R19866 GNDA.n913 GNDA.n912 0.0682083
R19867 GNDA.n923 GNDA.n922 0.0682083
R19868 GNDA.n931 GNDA.n797 0.0682083
R19869 GNDA.n941 GNDA.n795 0.0682083
R19870 GNDA.n943 GNDA.n942 0.0682083
R19871 GNDA.n1147 GNDA.n1143 0.0682083
R19872 GNDA.n1157 GNDA.n1141 0.0682083
R19873 GNDA.n1159 GNDA.n1158 0.0682083
R19874 GNDA.n1169 GNDA.n1168 0.0682083
R19875 GNDA.n1177 GNDA.n1137 0.0682083
R19876 GNDA.n1187 GNDA.n1135 0.0682083
R19877 GNDA.n1189 GNDA.n1188 0.0682083
R19878 GNDA.n1065 GNDA.n1061 0.0682083
R19879 GNDA.n1075 GNDA.n1059 0.0682083
R19880 GNDA.n1077 GNDA.n1076 0.0682083
R19881 GNDA.n1087 GNDA.n1086 0.0682083
R19882 GNDA.n1095 GNDA.n1055 0.0682083
R19883 GNDA.n1105 GNDA.n1053 0.0682083
R19884 GNDA.n1107 GNDA.n1106 0.0682083
R19885 GNDA.n983 GNDA.n979 0.0682083
R19886 GNDA.n993 GNDA.n977 0.0682083
R19887 GNDA.n995 GNDA.n994 0.0682083
R19888 GNDA.n1005 GNDA.n1004 0.0682083
R19889 GNDA.n1013 GNDA.n973 0.0682083
R19890 GNDA.n1023 GNDA.n971 0.0682083
R19891 GNDA.n1025 GNDA.n1024 0.0682083
R19892 GNDA.n886 GNDA.n806 0.0682083
R19893 GNDA.n832 GNDA.n831 0.0682083
R19894 GNDA.n834 GNDA.n833 0.0682083
R19895 GNDA.n838 GNDA.n837 0.0682083
R19896 GNDA.n840 GNDA.n839 0.0682083
R19897 GNDA.n844 GNDA.n843 0.0682083
R19898 GNDA.n846 GNDA.n845 0.0682083
R19899 GNDA.n735 GNDA.n655 0.0682083
R19900 GNDA.n681 GNDA.n680 0.0682083
R19901 GNDA.n683 GNDA.n682 0.0682083
R19902 GNDA.n687 GNDA.n686 0.0682083
R19903 GNDA.n689 GNDA.n688 0.0682083
R19904 GNDA.n693 GNDA.n692 0.0682083
R19905 GNDA.n695 GNDA.n694 0.0682083
R19906 GNDA.n3403 GNDA.n3399 0.0682083
R19907 GNDA.n3413 GNDA.n650 0.0682083
R19908 GNDA.n3415 GNDA.n3414 0.0682083
R19909 GNDA.n3425 GNDA.n3424 0.0682083
R19910 GNDA.n3433 GNDA.n646 0.0682083
R19911 GNDA.n3443 GNDA.n644 0.0682083
R19912 GNDA.n3445 GNDA.n3444 0.0682083
R19913 GNDA.n3524 GNDA.n612 0.0682083
R19914 GNDA.n3478 GNDA.n3467 0.0682083
R19915 GNDA.n3480 GNDA.n3479 0.0682083
R19916 GNDA.n3490 GNDA.n3489 0.0682083
R19917 GNDA.n3498 GNDA.n3463 0.0682083
R19918 GNDA.n3508 GNDA.n3461 0.0682083
R19919 GNDA.n3510 GNDA.n3509 0.0682083
R19920 GNDA.n2258 GNDA.n2178 0.0682083
R19921 GNDA.n2204 GNDA.n2203 0.0682083
R19922 GNDA.n2206 GNDA.n2205 0.0682083
R19923 GNDA.n2210 GNDA.n2209 0.0682083
R19924 GNDA.n2212 GNDA.n2211 0.0682083
R19925 GNDA.n2216 GNDA.n2215 0.0682083
R19926 GNDA.n2218 GNDA.n2217 0.0682083
R19927 GNDA.n2289 GNDA.n2288 0.0682083
R19928 GNDA.n2299 GNDA.n2298 0.0682083
R19929 GNDA.n2307 GNDA.n2171 0.0682083
R19930 GNDA.n2317 GNDA.n2169 0.0682083
R19931 GNDA.n2319 GNDA.n2318 0.0682083
R19932 GNDA.n2329 GNDA.n2328 0.0682083
R19933 GNDA.n2336 GNDA.n2165 0.0682083
R19934 GNDA.n2582 GNDA.n2581 0.0672139
R19935 GNDA.n3660 GNDA.n3639 0.0672139
R19936 GNDA.n4568 GNDA.n4507 0.0672139
R19937 GNDA.n4492 GNDA.n4426 0.0672139
R19938 GNDA.n4410 GNDA.n4344 0.0672139
R19939 GNDA.n4328 GNDA.n4262 0.0672139
R19940 GNDA.n4246 GNDA.n4180 0.0672139
R19941 GNDA.n4000 GNDA.n516 0.0672139
R19942 GNDA.n4164 GNDA.n4098 0.0672139
R19943 GNDA.n4082 GNDA.n4016 0.0672139
R19944 GNDA.n3897 GNDA.n3876 0.0672139
R19945 GNDA.n3839 GNDA.n3778 0.0672139
R19946 GNDA.n3763 GNDA.n552 0.0672139
R19947 GNDA.n1438 GNDA.n1377 0.0672139
R19948 GNDA.n1362 GNDA.n1296 0.0672139
R19949 GNDA.n1280 GNDA.n1214 0.0672139
R19950 GNDA.n952 GNDA.n792 0.0672139
R19951 GNDA.n1198 GNDA.n1132 0.0672139
R19952 GNDA.n1116 GNDA.n1050 0.0672139
R19953 GNDA.n1034 GNDA.n968 0.0672139
R19954 GNDA.n849 GNDA.n828 0.0672139
R19955 GNDA.n698 GNDA.n677 0.0672139
R19956 GNDA.n3454 GNDA.n641 0.0672139
R19957 GNDA.n3519 GNDA.n3458 0.0672139
R19958 GNDA.n2221 GNDA.n2200 0.0672139
R19959 GNDA.n2338 GNDA.n2164 0.0672139
R19960 GNDA.n2495 GNDA.n2493 0.0667303
R19961 GNDA.n2591 GNDA.n2590 0.063
R19962 GNDA.n2600 GNDA.n2568 0.063
R19963 GNDA.n2615 GNDA.n2614 0.063
R19964 GNDA.n3644 GNDA.n3643 0.063
R19965 GNDA.n3650 GNDA.n3649 0.063
R19966 GNDA.n3656 GNDA.n3655 0.063
R19967 GNDA.n4528 GNDA.n4527 0.063
R19968 GNDA.n4539 GNDA.n4512 0.063
R19969 GNDA.n4558 GNDA.n4557 0.063
R19970 GNDA.n4452 GNDA.n4451 0.063
R19971 GNDA.n4463 GNDA.n4431 0.063
R19972 GNDA.n4482 GNDA.n4481 0.063
R19973 GNDA.n4370 GNDA.n4369 0.063
R19974 GNDA.n4381 GNDA.n4349 0.063
R19975 GNDA.n4400 GNDA.n4399 0.063
R19976 GNDA.n4288 GNDA.n4287 0.063
R19977 GNDA.n4299 GNDA.n4267 0.063
R19978 GNDA.n4318 GNDA.n4317 0.063
R19979 GNDA.n4206 GNDA.n4205 0.063
R19980 GNDA.n4217 GNDA.n4185 0.063
R19981 GNDA.n4236 GNDA.n4235 0.063
R19982 GNDA.n3960 GNDA.n3959 0.063
R19983 GNDA.n3971 GNDA.n521 0.063
R19984 GNDA.n3990 GNDA.n3989 0.063
R19985 GNDA.n4124 GNDA.n4123 0.063
R19986 GNDA.n4135 GNDA.n4103 0.063
R19987 GNDA.n4154 GNDA.n4153 0.063
R19988 GNDA.n4042 GNDA.n4041 0.063
R19989 GNDA.n4053 GNDA.n4021 0.063
R19990 GNDA.n4072 GNDA.n4071 0.063
R19991 GNDA.n3881 GNDA.n3880 0.063
R19992 GNDA.n3887 GNDA.n3886 0.063
R19993 GNDA.n3893 GNDA.n3892 0.063
R19994 GNDA.n3799 GNDA.n3798 0.063
R19995 GNDA.n3810 GNDA.n3783 0.063
R19996 GNDA.n3829 GNDA.n3828 0.063
R19997 GNDA.n3723 GNDA.n3722 0.063
R19998 GNDA.n3734 GNDA.n557 0.063
R19999 GNDA.n3753 GNDA.n3752 0.063
R20000 GNDA.n1398 GNDA.n1397 0.063
R20001 GNDA.n1409 GNDA.n1382 0.063
R20002 GNDA.n1428 GNDA.n1427 0.063
R20003 GNDA.n1322 GNDA.n1321 0.063
R20004 GNDA.n1333 GNDA.n1301 0.063
R20005 GNDA.n1352 GNDA.n1351 0.063
R20006 GNDA.n1240 GNDA.n1239 0.063
R20007 GNDA.n1251 GNDA.n1219 0.063
R20008 GNDA.n1270 GNDA.n1269 0.063
R20009 GNDA.n912 GNDA.n911 0.063
R20010 GNDA.n923 GNDA.n797 0.063
R20011 GNDA.n942 GNDA.n941 0.063
R20012 GNDA.n1158 GNDA.n1157 0.063
R20013 GNDA.n1169 GNDA.n1137 0.063
R20014 GNDA.n1188 GNDA.n1187 0.063
R20015 GNDA.n1076 GNDA.n1075 0.063
R20016 GNDA.n1087 GNDA.n1055 0.063
R20017 GNDA.n1106 GNDA.n1105 0.063
R20018 GNDA.n994 GNDA.n993 0.063
R20019 GNDA.n1005 GNDA.n973 0.063
R20020 GNDA.n1024 GNDA.n1023 0.063
R20021 GNDA.n833 GNDA.n832 0.063
R20022 GNDA.n839 GNDA.n838 0.063
R20023 GNDA.n845 GNDA.n844 0.063
R20024 GNDA.n682 GNDA.n681 0.063
R20025 GNDA.n688 GNDA.n687 0.063
R20026 GNDA.n694 GNDA.n693 0.063
R20027 GNDA.n3414 GNDA.n3413 0.063
R20028 GNDA.n3425 GNDA.n646 0.063
R20029 GNDA.n3444 GNDA.n3443 0.063
R20030 GNDA.n3479 GNDA.n3478 0.063
R20031 GNDA.n3490 GNDA.n3463 0.063
R20032 GNDA.n3509 GNDA.n3508 0.063
R20033 GNDA.n2205 GNDA.n2204 0.063
R20034 GNDA.n2211 GNDA.n2210 0.063
R20035 GNDA.n2217 GNDA.n2216 0.063
R20036 GNDA.n2299 GNDA.n2171 0.063
R20037 GNDA.n2318 GNDA.n2317 0.063
R20038 GNDA.n2329 GNDA.n2165 0.063
R20039 GNDA.n3615 GNDA.n570 0.063
R20040 GNDA.n2928 GNDA.n2663 0.063
R20041 GNDA.n894 GNDA.n747 0.0629369
R20042 GNDA.n3938 GNDA.n3853 0.0629369
R20043 GNDA.n2717 GNDA.n2716 0.0626438
R20044 GNDA.n2704 GNDA.n2703 0.0626438
R20045 GNDA.n2625 GNDA.n358 0.0626438
R20046 GNDA.n3367 GNDA.n3366 0.0577917
R20047 GNDA.n2579 GNDA.n2578 0.0553333
R20048 GNDA.n2596 GNDA.n2595 0.0553333
R20049 GNDA.n2567 GNDA.n2566 0.0553333
R20050 GNDA.n2620 GNDA.n2619 0.0553333
R20051 GNDA.n3692 GNDA.n3691 0.0553333
R20052 GNDA.n3683 GNDA.n3682 0.0553333
R20053 GNDA.n3674 GNDA.n3673 0.0553333
R20054 GNDA.n3665 GNDA.n3664 0.0553333
R20055 GNDA.n4521 GNDA.n4520 0.0553333
R20056 GNDA.n4535 GNDA.n4534 0.0553333
R20057 GNDA.n4551 GNDA.n4550 0.0553333
R20058 GNDA.n4565 GNDA.n4564 0.0553333
R20059 GNDA.n4445 GNDA.n4444 0.0553333
R20060 GNDA.n4459 GNDA.n4458 0.0553333
R20061 GNDA.n4475 GNDA.n4474 0.0553333
R20062 GNDA.n4489 GNDA.n4488 0.0553333
R20063 GNDA.n4363 GNDA.n4362 0.0553333
R20064 GNDA.n4377 GNDA.n4376 0.0553333
R20065 GNDA.n4393 GNDA.n4392 0.0553333
R20066 GNDA.n4407 GNDA.n4406 0.0553333
R20067 GNDA.n4281 GNDA.n4280 0.0553333
R20068 GNDA.n4295 GNDA.n4294 0.0553333
R20069 GNDA.n4311 GNDA.n4310 0.0553333
R20070 GNDA.n4325 GNDA.n4324 0.0553333
R20071 GNDA.n4199 GNDA.n4198 0.0553333
R20072 GNDA.n4213 GNDA.n4212 0.0553333
R20073 GNDA.n4229 GNDA.n4228 0.0553333
R20074 GNDA.n4243 GNDA.n4242 0.0553333
R20075 GNDA.n3953 GNDA.n3952 0.0553333
R20076 GNDA.n3967 GNDA.n3966 0.0553333
R20077 GNDA.n3983 GNDA.n3982 0.0553333
R20078 GNDA.n3997 GNDA.n3996 0.0553333
R20079 GNDA.n4117 GNDA.n4116 0.0553333
R20080 GNDA.n4131 GNDA.n4130 0.0553333
R20081 GNDA.n4147 GNDA.n4146 0.0553333
R20082 GNDA.n4161 GNDA.n4160 0.0553333
R20083 GNDA.n4035 GNDA.n4034 0.0553333
R20084 GNDA.n4049 GNDA.n4048 0.0553333
R20085 GNDA.n4065 GNDA.n4064 0.0553333
R20086 GNDA.n4079 GNDA.n4078 0.0553333
R20087 GNDA.n3929 GNDA.n3928 0.0553333
R20088 GNDA.n3920 GNDA.n3919 0.0553333
R20089 GNDA.n3911 GNDA.n3910 0.0553333
R20090 GNDA.n3902 GNDA.n3901 0.0553333
R20091 GNDA.n3792 GNDA.n3791 0.0553333
R20092 GNDA.n3806 GNDA.n3805 0.0553333
R20093 GNDA.n3822 GNDA.n3821 0.0553333
R20094 GNDA.n3836 GNDA.n3835 0.0553333
R20095 GNDA.n3716 GNDA.n3715 0.0553333
R20096 GNDA.n3730 GNDA.n3729 0.0553333
R20097 GNDA.n3746 GNDA.n3745 0.0553333
R20098 GNDA.n3760 GNDA.n3759 0.0553333
R20099 GNDA.n1391 GNDA.n1390 0.0553333
R20100 GNDA.n1405 GNDA.n1404 0.0553333
R20101 GNDA.n1421 GNDA.n1420 0.0553333
R20102 GNDA.n1435 GNDA.n1434 0.0553333
R20103 GNDA.n1315 GNDA.n1314 0.0553333
R20104 GNDA.n1329 GNDA.n1328 0.0553333
R20105 GNDA.n1345 GNDA.n1344 0.0553333
R20106 GNDA.n1359 GNDA.n1358 0.0553333
R20107 GNDA.n1233 GNDA.n1232 0.0553333
R20108 GNDA.n1247 GNDA.n1246 0.0553333
R20109 GNDA.n1263 GNDA.n1262 0.0553333
R20110 GNDA.n1277 GNDA.n1276 0.0553333
R20111 GNDA.n905 GNDA.n904 0.0553333
R20112 GNDA.n919 GNDA.n918 0.0553333
R20113 GNDA.n935 GNDA.n934 0.0553333
R20114 GNDA.n949 GNDA.n948 0.0553333
R20115 GNDA.n1151 GNDA.n1150 0.0553333
R20116 GNDA.n1165 GNDA.n1164 0.0553333
R20117 GNDA.n1181 GNDA.n1180 0.0553333
R20118 GNDA.n1195 GNDA.n1194 0.0553333
R20119 GNDA.n1069 GNDA.n1068 0.0553333
R20120 GNDA.n1083 GNDA.n1082 0.0553333
R20121 GNDA.n1099 GNDA.n1098 0.0553333
R20122 GNDA.n1113 GNDA.n1112 0.0553333
R20123 GNDA.n987 GNDA.n986 0.0553333
R20124 GNDA.n1001 GNDA.n1000 0.0553333
R20125 GNDA.n1017 GNDA.n1016 0.0553333
R20126 GNDA.n1031 GNDA.n1030 0.0553333
R20127 GNDA.n881 GNDA.n880 0.0553333
R20128 GNDA.n872 GNDA.n871 0.0553333
R20129 GNDA.n863 GNDA.n862 0.0553333
R20130 GNDA.n854 GNDA.n853 0.0553333
R20131 GNDA.n730 GNDA.n729 0.0553333
R20132 GNDA.n721 GNDA.n720 0.0553333
R20133 GNDA.n712 GNDA.n711 0.0553333
R20134 GNDA.n703 GNDA.n702 0.0553333
R20135 GNDA.n3407 GNDA.n3406 0.0553333
R20136 GNDA.n3421 GNDA.n3420 0.0553333
R20137 GNDA.n3437 GNDA.n3436 0.0553333
R20138 GNDA.n3451 GNDA.n3450 0.0553333
R20139 GNDA.n3472 GNDA.n3471 0.0553333
R20140 GNDA.n3486 GNDA.n3485 0.0553333
R20141 GNDA.n3502 GNDA.n3501 0.0553333
R20142 GNDA.n3516 GNDA.n3515 0.0553333
R20143 GNDA.n2253 GNDA.n2252 0.0553333
R20144 GNDA.n2244 GNDA.n2243 0.0553333
R20145 GNDA.n2235 GNDA.n2234 0.0553333
R20146 GNDA.n2226 GNDA.n2225 0.0553333
R20147 GNDA.n2292 GNDA.n2291 0.0553333
R20148 GNDA.n2295 GNDA.n2294 0.0553333
R20149 GNDA.n2305 GNDA.n2304 0.0553333
R20150 GNDA.n2312 GNDA.n2311 0.0553333
R20151 GNDA.n2322 GNDA.n2321 0.0553333
R20152 GNDA.n2325 GNDA.n2324 0.0553333
R20153 GNDA.n2334 GNDA.n2161 0.0553333
R20154 GNDA.n2341 GNDA.n2162 0.0553333
R20155 GNDA.n2498 GNDA.n2497 0.0553333
R20156 GNDA.n2514 GNDA.n2513 0.0553333
R20157 GNDA.n2528 GNDA.n2527 0.0553333
R20158 GNDA.n2544 GNDA.n2482 0.0553333
R20159 GNDA.n3119 GNDA 0.0517
R20160 GNDA.n3300 GNDA 0.0517
R20161 GNDA GNDA.n202 0.0517
R20162 GNDA.n1688 GNDA 0.0517
R20163 GNDA GNDA.n4897 0.0517
R20164 GNDA GNDA.n5176 0.0517
R20165 GNDA.n4754 GNDA 0.0517
R20166 GNDA.n2833 GNDA 0.0517
R20167 GNDA GNDA.n0 0.0517
R20168 GNDA.n2580 GNDA.n2546 0.0514167
R20169 GNDA.n2588 GNDA.n2587 0.0514167
R20170 GNDA.n2575 GNDA.n2574 0.0514167
R20171 GNDA.n2571 GNDA.n2570 0.0514167
R20172 GNDA.n2604 GNDA.n2603 0.0514167
R20173 GNDA.n2612 GNDA.n2611 0.0514167
R20174 GNDA.n2563 GNDA.n2562 0.0514167
R20175 GNDA.n2638 GNDA.n2558 0.0514167
R20176 GNDA.n3695 GNDA.n3694 0.0514167
R20177 GNDA.n3689 GNDA.n3688 0.0514167
R20178 GNDA.n3686 GNDA.n3685 0.0514167
R20179 GNDA.n3680 GNDA.n3679 0.0514167
R20180 GNDA.n3677 GNDA.n3676 0.0514167
R20181 GNDA.n3671 GNDA.n3670 0.0514167
R20182 GNDA.n3668 GNDA.n3667 0.0514167
R20183 GNDA.n3662 GNDA.n3661 0.0514167
R20184 GNDA.n4571 GNDA.n501 0.0514167
R20185 GNDA.n4525 GNDA.n4524 0.0514167
R20186 GNDA.n4531 GNDA.n4530 0.0514167
R20187 GNDA.n4541 GNDA.n4540 0.0514167
R20188 GNDA.n4545 GNDA.n4544 0.0514167
R20189 GNDA.n4555 GNDA.n4554 0.0514167
R20190 GNDA.n4561 GNDA.n4560 0.0514167
R20191 GNDA.n4569 GNDA.n4506 0.0514167
R20192 GNDA.n4439 GNDA.n4413 0.0514167
R20193 GNDA.n4449 GNDA.n4448 0.0514167
R20194 GNDA.n4455 GNDA.n4454 0.0514167
R20195 GNDA.n4465 GNDA.n4464 0.0514167
R20196 GNDA.n4469 GNDA.n4468 0.0514167
R20197 GNDA.n4479 GNDA.n4478 0.0514167
R20198 GNDA.n4485 GNDA.n4484 0.0514167
R20199 GNDA.n4493 GNDA.n4425 0.0514167
R20200 GNDA.n4357 GNDA.n4331 0.0514167
R20201 GNDA.n4367 GNDA.n4366 0.0514167
R20202 GNDA.n4373 GNDA.n4372 0.0514167
R20203 GNDA.n4383 GNDA.n4382 0.0514167
R20204 GNDA.n4387 GNDA.n4386 0.0514167
R20205 GNDA.n4397 GNDA.n4396 0.0514167
R20206 GNDA.n4403 GNDA.n4402 0.0514167
R20207 GNDA.n4411 GNDA.n4343 0.0514167
R20208 GNDA.n4275 GNDA.n4249 0.0514167
R20209 GNDA.n4285 GNDA.n4284 0.0514167
R20210 GNDA.n4291 GNDA.n4290 0.0514167
R20211 GNDA.n4301 GNDA.n4300 0.0514167
R20212 GNDA.n4305 GNDA.n4304 0.0514167
R20213 GNDA.n4315 GNDA.n4314 0.0514167
R20214 GNDA.n4321 GNDA.n4320 0.0514167
R20215 GNDA.n4329 GNDA.n4261 0.0514167
R20216 GNDA.n4193 GNDA.n4167 0.0514167
R20217 GNDA.n4203 GNDA.n4202 0.0514167
R20218 GNDA.n4209 GNDA.n4208 0.0514167
R20219 GNDA.n4219 GNDA.n4218 0.0514167
R20220 GNDA.n4223 GNDA.n4222 0.0514167
R20221 GNDA.n4233 GNDA.n4232 0.0514167
R20222 GNDA.n4239 GNDA.n4238 0.0514167
R20223 GNDA.n4247 GNDA.n4179 0.0514167
R20224 GNDA.n3947 GNDA.n503 0.0514167
R20225 GNDA.n3957 GNDA.n3956 0.0514167
R20226 GNDA.n3963 GNDA.n3962 0.0514167
R20227 GNDA.n3973 GNDA.n3972 0.0514167
R20228 GNDA.n3977 GNDA.n3976 0.0514167
R20229 GNDA.n3987 GNDA.n3986 0.0514167
R20230 GNDA.n3993 GNDA.n3992 0.0514167
R20231 GNDA.n4001 GNDA.n515 0.0514167
R20232 GNDA.n4111 GNDA.n4085 0.0514167
R20233 GNDA.n4121 GNDA.n4120 0.0514167
R20234 GNDA.n4127 GNDA.n4126 0.0514167
R20235 GNDA.n4137 GNDA.n4136 0.0514167
R20236 GNDA.n4141 GNDA.n4140 0.0514167
R20237 GNDA.n4151 GNDA.n4150 0.0514167
R20238 GNDA.n4157 GNDA.n4156 0.0514167
R20239 GNDA.n4165 GNDA.n4097 0.0514167
R20240 GNDA.n4029 GNDA.n4003 0.0514167
R20241 GNDA.n4039 GNDA.n4038 0.0514167
R20242 GNDA.n4045 GNDA.n4044 0.0514167
R20243 GNDA.n4055 GNDA.n4054 0.0514167
R20244 GNDA.n4059 GNDA.n4058 0.0514167
R20245 GNDA.n4069 GNDA.n4068 0.0514167
R20246 GNDA.n4075 GNDA.n4074 0.0514167
R20247 GNDA.n4083 GNDA.n4015 0.0514167
R20248 GNDA.n3932 GNDA.n3931 0.0514167
R20249 GNDA.n3926 GNDA.n3925 0.0514167
R20250 GNDA.n3923 GNDA.n3922 0.0514167
R20251 GNDA.n3917 GNDA.n3916 0.0514167
R20252 GNDA.n3914 GNDA.n3913 0.0514167
R20253 GNDA.n3908 GNDA.n3907 0.0514167
R20254 GNDA.n3905 GNDA.n3904 0.0514167
R20255 GNDA.n3899 GNDA.n3898 0.0514167
R20256 GNDA.n3842 GNDA.n537 0.0514167
R20257 GNDA.n3796 GNDA.n3795 0.0514167
R20258 GNDA.n3802 GNDA.n3801 0.0514167
R20259 GNDA.n3812 GNDA.n3811 0.0514167
R20260 GNDA.n3816 GNDA.n3815 0.0514167
R20261 GNDA.n3826 GNDA.n3825 0.0514167
R20262 GNDA.n3832 GNDA.n3831 0.0514167
R20263 GNDA.n3840 GNDA.n3777 0.0514167
R20264 GNDA.n3710 GNDA.n539 0.0514167
R20265 GNDA.n3720 GNDA.n3719 0.0514167
R20266 GNDA.n3726 GNDA.n3725 0.0514167
R20267 GNDA.n3736 GNDA.n3735 0.0514167
R20268 GNDA.n3740 GNDA.n3739 0.0514167
R20269 GNDA.n3750 GNDA.n3749 0.0514167
R20270 GNDA.n3756 GNDA.n3755 0.0514167
R20271 GNDA.n3764 GNDA.n551 0.0514167
R20272 GNDA.n1441 GNDA.n777 0.0514167
R20273 GNDA.n1395 GNDA.n1394 0.0514167
R20274 GNDA.n1401 GNDA.n1400 0.0514167
R20275 GNDA.n1411 GNDA.n1410 0.0514167
R20276 GNDA.n1415 GNDA.n1414 0.0514167
R20277 GNDA.n1425 GNDA.n1424 0.0514167
R20278 GNDA.n1431 GNDA.n1430 0.0514167
R20279 GNDA.n1439 GNDA.n1376 0.0514167
R20280 GNDA.n1309 GNDA.n1283 0.0514167
R20281 GNDA.n1319 GNDA.n1318 0.0514167
R20282 GNDA.n1325 GNDA.n1324 0.0514167
R20283 GNDA.n1335 GNDA.n1334 0.0514167
R20284 GNDA.n1339 GNDA.n1338 0.0514167
R20285 GNDA.n1349 GNDA.n1348 0.0514167
R20286 GNDA.n1355 GNDA.n1354 0.0514167
R20287 GNDA.n1363 GNDA.n1295 0.0514167
R20288 GNDA.n1227 GNDA.n1201 0.0514167
R20289 GNDA.n1237 GNDA.n1236 0.0514167
R20290 GNDA.n1243 GNDA.n1242 0.0514167
R20291 GNDA.n1253 GNDA.n1252 0.0514167
R20292 GNDA.n1257 GNDA.n1256 0.0514167
R20293 GNDA.n1267 GNDA.n1266 0.0514167
R20294 GNDA.n1273 GNDA.n1272 0.0514167
R20295 GNDA.n1281 GNDA.n1213 0.0514167
R20296 GNDA.n899 GNDA.n779 0.0514167
R20297 GNDA.n909 GNDA.n908 0.0514167
R20298 GNDA.n915 GNDA.n914 0.0514167
R20299 GNDA.n925 GNDA.n924 0.0514167
R20300 GNDA.n929 GNDA.n928 0.0514167
R20301 GNDA.n939 GNDA.n938 0.0514167
R20302 GNDA.n945 GNDA.n944 0.0514167
R20303 GNDA.n953 GNDA.n791 0.0514167
R20304 GNDA.n1145 GNDA.n1119 0.0514167
R20305 GNDA.n1155 GNDA.n1154 0.0514167
R20306 GNDA.n1161 GNDA.n1160 0.0514167
R20307 GNDA.n1171 GNDA.n1170 0.0514167
R20308 GNDA.n1175 GNDA.n1174 0.0514167
R20309 GNDA.n1185 GNDA.n1184 0.0514167
R20310 GNDA.n1191 GNDA.n1190 0.0514167
R20311 GNDA.n1199 GNDA.n1131 0.0514167
R20312 GNDA.n1063 GNDA.n1037 0.0514167
R20313 GNDA.n1073 GNDA.n1072 0.0514167
R20314 GNDA.n1079 GNDA.n1078 0.0514167
R20315 GNDA.n1089 GNDA.n1088 0.0514167
R20316 GNDA.n1093 GNDA.n1092 0.0514167
R20317 GNDA.n1103 GNDA.n1102 0.0514167
R20318 GNDA.n1109 GNDA.n1108 0.0514167
R20319 GNDA.n1117 GNDA.n1049 0.0514167
R20320 GNDA.n981 GNDA.n955 0.0514167
R20321 GNDA.n991 GNDA.n990 0.0514167
R20322 GNDA.n997 GNDA.n996 0.0514167
R20323 GNDA.n1007 GNDA.n1006 0.0514167
R20324 GNDA.n1011 GNDA.n1010 0.0514167
R20325 GNDA.n1021 GNDA.n1020 0.0514167
R20326 GNDA.n1027 GNDA.n1026 0.0514167
R20327 GNDA.n1035 GNDA.n967 0.0514167
R20328 GNDA.n884 GNDA.n883 0.0514167
R20329 GNDA.n878 GNDA.n877 0.0514167
R20330 GNDA.n875 GNDA.n874 0.0514167
R20331 GNDA.n869 GNDA.n868 0.0514167
R20332 GNDA.n866 GNDA.n865 0.0514167
R20333 GNDA.n860 GNDA.n859 0.0514167
R20334 GNDA.n857 GNDA.n856 0.0514167
R20335 GNDA.n851 GNDA.n850 0.0514167
R20336 GNDA.n733 GNDA.n732 0.0514167
R20337 GNDA.n727 GNDA.n726 0.0514167
R20338 GNDA.n724 GNDA.n723 0.0514167
R20339 GNDA.n718 GNDA.n717 0.0514167
R20340 GNDA.n715 GNDA.n714 0.0514167
R20341 GNDA.n709 GNDA.n708 0.0514167
R20342 GNDA.n706 GNDA.n705 0.0514167
R20343 GNDA.n700 GNDA.n699 0.0514167
R20344 GNDA.n3401 GNDA.n627 0.0514167
R20345 GNDA.n3411 GNDA.n3410 0.0514167
R20346 GNDA.n3417 GNDA.n3416 0.0514167
R20347 GNDA.n3427 GNDA.n3426 0.0514167
R20348 GNDA.n3431 GNDA.n3430 0.0514167
R20349 GNDA.n3441 GNDA.n3440 0.0514167
R20350 GNDA.n3447 GNDA.n3446 0.0514167
R20351 GNDA.n3455 GNDA.n640 0.0514167
R20352 GNDA.n3522 GNDA.n614 0.0514167
R20353 GNDA.n3476 GNDA.n3475 0.0514167
R20354 GNDA.n3482 GNDA.n3481 0.0514167
R20355 GNDA.n3492 GNDA.n3491 0.0514167
R20356 GNDA.n3496 GNDA.n3495 0.0514167
R20357 GNDA.n3506 GNDA.n3505 0.0514167
R20358 GNDA.n3512 GNDA.n3511 0.0514167
R20359 GNDA.n3520 GNDA.n3457 0.0514167
R20360 GNDA.n2256 GNDA.n2255 0.0514167
R20361 GNDA.n2250 GNDA.n2249 0.0514167
R20362 GNDA.n2247 GNDA.n2246 0.0514167
R20363 GNDA.n2241 GNDA.n2240 0.0514167
R20364 GNDA.n2238 GNDA.n2237 0.0514167
R20365 GNDA.n2232 GNDA.n2231 0.0514167
R20366 GNDA.n2229 GNDA.n2228 0.0514167
R20367 GNDA.n2223 GNDA.n2222 0.0514167
R20368 GNDA.n2494 GNDA.n2471 0.0514167
R20369 GNDA.n2504 GNDA.n2503 0.0514167
R20370 GNDA.n2508 GNDA.n2507 0.0514167
R20371 GNDA.n2518 GNDA.n2517 0.0514167
R20372 GNDA.n2524 GNDA.n2523 0.0514167
R20373 GNDA.n2534 GNDA.n2533 0.0514167
R20374 GNDA.n2538 GNDA.n2537 0.0514167
R20375 GNDA.n2641 GNDA.n1866 0.0514167
R20376 GNDA.n2302 GNDA.n2301 0.0475
R20377 GNDA.n2315 GNDA.n2314 0.0475
R20378 GNDA.n2332 GNDA.n2331 0.0475
R20379 GNDA.n3334 GNDA.n3328 0.0421667
R20380 GNDA.n3589 GNDA.n580 0.0421667
R20381 GNDA.n3560 GNDA.n594 0.0421667
R20382 GNDA.n3538 GNDA.n602 0.0421667
R20383 GNDA.n472 GNDA.n448 0.0421667
R20384 GNDA.n2698 GNDA.n1524 0.0421667
R20385 GNDA.n2633 GNDA.n2632 0.0421667
R20386 GNDA.n3937 GNDA.n3935 0.0421667
R20387 GNDA.n896 GNDA.n895 0.0421667
R20388 GNDA.n2276 GNDA.n2269 0.0421667
R20389 GNDA.n2281 GNDA.n2266 0.0421667
R20390 GNDA.n2283 GNDA.n2265 0.0421667
R20391 GNDA.n2262 GNDA.n610 0.0421667
R20392 GNDA.n3529 GNDA.n607 0.0421667
R20393 GNDA.n3532 GNDA.n606 0.0421667
R20394 GNDA.n3392 GNDA.n3391 0.0421667
R20395 GNDA.n3388 GNDA.n3387 0.0421667
R20396 GNDA.n893 GNDA.n804 0.0421667
R20397 GNDA.n3376 GNDA.n3375 0.0421667
R20398 GNDA.n3372 GNDA.n3371 0.0421667
R20399 GNDA.n3368 GNDA.n3367 0.0421667
R20400 GNDA.n1459 GNDA.n1458 0.0421667
R20401 GNDA.n1455 GNDA.n1454 0.0421667
R20402 GNDA.n1447 GNDA.n570 0.0421667
R20403 GNDA.n3702 GNDA.n566 0.0421667
R20404 GNDA.n564 GNDA.n533 0.0421667
R20405 GNDA.n3849 GNDA.n530 0.0421667
R20406 GNDA.n528 GNDA.n435 0.0421667
R20407 GNDA.n4606 GNDA.n4605 0.0421667
R20408 GNDA.n4602 GNDA.n4601 0.0421667
R20409 GNDA.n4598 GNDA.n4597 0.0421667
R20410 GNDA.n4594 GNDA.n4593 0.0421667
R20411 GNDA.n4590 GNDA.n4589 0.0421667
R20412 GNDA.n4586 GNDA.n4585 0.0421667
R20413 GNDA.n4582 GNDA.n4581 0.0421667
R20414 GNDA.n4578 GNDA.n4577 0.0421667
R20415 GNDA.n2578 GNDA.n2547 0.028198
R20416 GNDA.n2587 GNDA.n2548 0.028198
R20417 GNDA.n2595 GNDA.n2550 0.028198
R20418 GNDA.n2570 GNDA.n2551 0.028198
R20419 GNDA.n2566 GNDA.n2553 0.028198
R20420 GNDA.n2611 GNDA.n2554 0.028198
R20421 GNDA.n2619 GNDA.n2556 0.028198
R20422 GNDA.n2558 GNDA.n2557 0.028198
R20423 GNDA.n3693 GNDA.n3692 0.028198
R20424 GNDA.n3690 GNDA.n3689 0.028198
R20425 GNDA.n3684 GNDA.n3683 0.028198
R20426 GNDA.n3681 GNDA.n3680 0.028198
R20427 GNDA.n3675 GNDA.n3674 0.028198
R20428 GNDA.n3672 GNDA.n3671 0.028198
R20429 GNDA.n3666 GNDA.n3665 0.028198
R20430 GNDA.n3663 GNDA.n3662 0.028198
R20431 GNDA.n4520 GNDA.n4495 0.028198
R20432 GNDA.n4524 GNDA.n4496 0.028198
R20433 GNDA.n4534 GNDA.n4498 0.028198
R20434 GNDA.n4540 GNDA.n4499 0.028198
R20435 GNDA.n4550 GNDA.n4501 0.028198
R20436 GNDA.n4554 GNDA.n4502 0.028198
R20437 GNDA.n4564 GNDA.n4504 0.028198
R20438 GNDA.n4506 GNDA.n4505 0.028198
R20439 GNDA.n4444 GNDA.n4414 0.028198
R20440 GNDA.n4448 GNDA.n4415 0.028198
R20441 GNDA.n4458 GNDA.n4417 0.028198
R20442 GNDA.n4464 GNDA.n4418 0.028198
R20443 GNDA.n4474 GNDA.n4420 0.028198
R20444 GNDA.n4478 GNDA.n4421 0.028198
R20445 GNDA.n4488 GNDA.n4423 0.028198
R20446 GNDA.n4425 GNDA.n4424 0.028198
R20447 GNDA.n4362 GNDA.n4332 0.028198
R20448 GNDA.n4366 GNDA.n4333 0.028198
R20449 GNDA.n4376 GNDA.n4335 0.028198
R20450 GNDA.n4382 GNDA.n4336 0.028198
R20451 GNDA.n4392 GNDA.n4338 0.028198
R20452 GNDA.n4396 GNDA.n4339 0.028198
R20453 GNDA.n4406 GNDA.n4341 0.028198
R20454 GNDA.n4343 GNDA.n4342 0.028198
R20455 GNDA.n4280 GNDA.n4250 0.028198
R20456 GNDA.n4284 GNDA.n4251 0.028198
R20457 GNDA.n4294 GNDA.n4253 0.028198
R20458 GNDA.n4300 GNDA.n4254 0.028198
R20459 GNDA.n4310 GNDA.n4256 0.028198
R20460 GNDA.n4314 GNDA.n4257 0.028198
R20461 GNDA.n4324 GNDA.n4259 0.028198
R20462 GNDA.n4261 GNDA.n4260 0.028198
R20463 GNDA.n4198 GNDA.n4168 0.028198
R20464 GNDA.n4202 GNDA.n4169 0.028198
R20465 GNDA.n4212 GNDA.n4171 0.028198
R20466 GNDA.n4218 GNDA.n4172 0.028198
R20467 GNDA.n4228 GNDA.n4174 0.028198
R20468 GNDA.n4232 GNDA.n4175 0.028198
R20469 GNDA.n4242 GNDA.n4177 0.028198
R20470 GNDA.n4179 GNDA.n4178 0.028198
R20471 GNDA.n3952 GNDA.n504 0.028198
R20472 GNDA.n3956 GNDA.n505 0.028198
R20473 GNDA.n3966 GNDA.n507 0.028198
R20474 GNDA.n3972 GNDA.n508 0.028198
R20475 GNDA.n3982 GNDA.n510 0.028198
R20476 GNDA.n3986 GNDA.n511 0.028198
R20477 GNDA.n3996 GNDA.n513 0.028198
R20478 GNDA.n515 GNDA.n514 0.028198
R20479 GNDA.n4116 GNDA.n4086 0.028198
R20480 GNDA.n4120 GNDA.n4087 0.028198
R20481 GNDA.n4130 GNDA.n4089 0.028198
R20482 GNDA.n4136 GNDA.n4090 0.028198
R20483 GNDA.n4146 GNDA.n4092 0.028198
R20484 GNDA.n4150 GNDA.n4093 0.028198
R20485 GNDA.n4160 GNDA.n4095 0.028198
R20486 GNDA.n4097 GNDA.n4096 0.028198
R20487 GNDA.n4034 GNDA.n4004 0.028198
R20488 GNDA.n4038 GNDA.n4005 0.028198
R20489 GNDA.n4048 GNDA.n4007 0.028198
R20490 GNDA.n4054 GNDA.n4008 0.028198
R20491 GNDA.n4064 GNDA.n4010 0.028198
R20492 GNDA.n4068 GNDA.n4011 0.028198
R20493 GNDA.n4078 GNDA.n4013 0.028198
R20494 GNDA.n4015 GNDA.n4014 0.028198
R20495 GNDA.n3930 GNDA.n3929 0.028198
R20496 GNDA.n3927 GNDA.n3926 0.028198
R20497 GNDA.n3921 GNDA.n3920 0.028198
R20498 GNDA.n3918 GNDA.n3917 0.028198
R20499 GNDA.n3912 GNDA.n3911 0.028198
R20500 GNDA.n3909 GNDA.n3908 0.028198
R20501 GNDA.n3903 GNDA.n3902 0.028198
R20502 GNDA.n3900 GNDA.n3899 0.028198
R20503 GNDA.n3791 GNDA.n3766 0.028198
R20504 GNDA.n3795 GNDA.n3767 0.028198
R20505 GNDA.n3805 GNDA.n3769 0.028198
R20506 GNDA.n3811 GNDA.n3770 0.028198
R20507 GNDA.n3821 GNDA.n3772 0.028198
R20508 GNDA.n3825 GNDA.n3773 0.028198
R20509 GNDA.n3835 GNDA.n3775 0.028198
R20510 GNDA.n3777 GNDA.n3776 0.028198
R20511 GNDA.n3715 GNDA.n540 0.028198
R20512 GNDA.n3719 GNDA.n541 0.028198
R20513 GNDA.n3729 GNDA.n543 0.028198
R20514 GNDA.n3735 GNDA.n544 0.028198
R20515 GNDA.n3745 GNDA.n546 0.028198
R20516 GNDA.n3749 GNDA.n547 0.028198
R20517 GNDA.n3759 GNDA.n549 0.028198
R20518 GNDA.n551 GNDA.n550 0.028198
R20519 GNDA.n1390 GNDA.n1365 0.028198
R20520 GNDA.n1394 GNDA.n1366 0.028198
R20521 GNDA.n1404 GNDA.n1368 0.028198
R20522 GNDA.n1410 GNDA.n1369 0.028198
R20523 GNDA.n1420 GNDA.n1371 0.028198
R20524 GNDA.n1424 GNDA.n1372 0.028198
R20525 GNDA.n1434 GNDA.n1374 0.028198
R20526 GNDA.n1376 GNDA.n1375 0.028198
R20527 GNDA.n1314 GNDA.n1284 0.028198
R20528 GNDA.n1318 GNDA.n1285 0.028198
R20529 GNDA.n1328 GNDA.n1287 0.028198
R20530 GNDA.n1334 GNDA.n1288 0.028198
R20531 GNDA.n1344 GNDA.n1290 0.028198
R20532 GNDA.n1348 GNDA.n1291 0.028198
R20533 GNDA.n1358 GNDA.n1293 0.028198
R20534 GNDA.n1295 GNDA.n1294 0.028198
R20535 GNDA.n1232 GNDA.n1202 0.028198
R20536 GNDA.n1236 GNDA.n1203 0.028198
R20537 GNDA.n1246 GNDA.n1205 0.028198
R20538 GNDA.n1252 GNDA.n1206 0.028198
R20539 GNDA.n1262 GNDA.n1208 0.028198
R20540 GNDA.n1266 GNDA.n1209 0.028198
R20541 GNDA.n1276 GNDA.n1211 0.028198
R20542 GNDA.n1213 GNDA.n1212 0.028198
R20543 GNDA.n904 GNDA.n780 0.028198
R20544 GNDA.n908 GNDA.n781 0.028198
R20545 GNDA.n918 GNDA.n783 0.028198
R20546 GNDA.n924 GNDA.n784 0.028198
R20547 GNDA.n934 GNDA.n786 0.028198
R20548 GNDA.n938 GNDA.n787 0.028198
R20549 GNDA.n948 GNDA.n789 0.028198
R20550 GNDA.n791 GNDA.n790 0.028198
R20551 GNDA.n1150 GNDA.n1120 0.028198
R20552 GNDA.n1154 GNDA.n1121 0.028198
R20553 GNDA.n1164 GNDA.n1123 0.028198
R20554 GNDA.n1170 GNDA.n1124 0.028198
R20555 GNDA.n1180 GNDA.n1126 0.028198
R20556 GNDA.n1184 GNDA.n1127 0.028198
R20557 GNDA.n1194 GNDA.n1129 0.028198
R20558 GNDA.n1131 GNDA.n1130 0.028198
R20559 GNDA.n1068 GNDA.n1038 0.028198
R20560 GNDA.n1072 GNDA.n1039 0.028198
R20561 GNDA.n1082 GNDA.n1041 0.028198
R20562 GNDA.n1088 GNDA.n1042 0.028198
R20563 GNDA.n1098 GNDA.n1044 0.028198
R20564 GNDA.n1102 GNDA.n1045 0.028198
R20565 GNDA.n1112 GNDA.n1047 0.028198
R20566 GNDA.n1049 GNDA.n1048 0.028198
R20567 GNDA.n986 GNDA.n956 0.028198
R20568 GNDA.n990 GNDA.n957 0.028198
R20569 GNDA.n1000 GNDA.n959 0.028198
R20570 GNDA.n1006 GNDA.n960 0.028198
R20571 GNDA.n1016 GNDA.n962 0.028198
R20572 GNDA.n1020 GNDA.n963 0.028198
R20573 GNDA.n1030 GNDA.n965 0.028198
R20574 GNDA.n967 GNDA.n966 0.028198
R20575 GNDA.n882 GNDA.n881 0.028198
R20576 GNDA.n879 GNDA.n878 0.028198
R20577 GNDA.n873 GNDA.n872 0.028198
R20578 GNDA.n870 GNDA.n869 0.028198
R20579 GNDA.n864 GNDA.n863 0.028198
R20580 GNDA.n861 GNDA.n860 0.028198
R20581 GNDA.n855 GNDA.n854 0.028198
R20582 GNDA.n852 GNDA.n851 0.028198
R20583 GNDA.n731 GNDA.n730 0.028198
R20584 GNDA.n728 GNDA.n727 0.028198
R20585 GNDA.n722 GNDA.n721 0.028198
R20586 GNDA.n719 GNDA.n718 0.028198
R20587 GNDA.n713 GNDA.n712 0.028198
R20588 GNDA.n710 GNDA.n709 0.028198
R20589 GNDA.n704 GNDA.n703 0.028198
R20590 GNDA.n701 GNDA.n700 0.028198
R20591 GNDA.n3406 GNDA.n628 0.028198
R20592 GNDA.n3410 GNDA.n629 0.028198
R20593 GNDA.n3420 GNDA.n631 0.028198
R20594 GNDA.n3426 GNDA.n632 0.028198
R20595 GNDA.n3436 GNDA.n634 0.028198
R20596 GNDA.n3440 GNDA.n635 0.028198
R20597 GNDA.n3450 GNDA.n637 0.028198
R20598 GNDA.n640 GNDA.n638 0.028198
R20599 GNDA.n3471 GNDA.n616 0.028198
R20600 GNDA.n3475 GNDA.n617 0.028198
R20601 GNDA.n3485 GNDA.n619 0.028198
R20602 GNDA.n3491 GNDA.n620 0.028198
R20603 GNDA.n3501 GNDA.n622 0.028198
R20604 GNDA.n3505 GNDA.n623 0.028198
R20605 GNDA.n3515 GNDA.n625 0.028198
R20606 GNDA.n3457 GNDA.n626 0.028198
R20607 GNDA.n2254 GNDA.n2253 0.028198
R20608 GNDA.n2251 GNDA.n2250 0.028198
R20609 GNDA.n2245 GNDA.n2244 0.028198
R20610 GNDA.n2242 GNDA.n2241 0.028198
R20611 GNDA.n2236 GNDA.n2235 0.028198
R20612 GNDA.n2233 GNDA.n2232 0.028198
R20613 GNDA.n2227 GNDA.n2226 0.028198
R20614 GNDA.n2224 GNDA.n2223 0.028198
R20615 GNDA.n2225 GNDA.n2224 0.028198
R20616 GNDA.n2228 GNDA.n2227 0.028198
R20617 GNDA.n2234 GNDA.n2233 0.028198
R20618 GNDA.n2237 GNDA.n2236 0.028198
R20619 GNDA.n2243 GNDA.n2242 0.028198
R20620 GNDA.n2246 GNDA.n2245 0.028198
R20621 GNDA.n2252 GNDA.n2251 0.028198
R20622 GNDA.n2255 GNDA.n2254 0.028198
R20623 GNDA.n3516 GNDA.n626 0.028198
R20624 GNDA.n3512 GNDA.n625 0.028198
R20625 GNDA.n3502 GNDA.n623 0.028198
R20626 GNDA.n3496 GNDA.n622 0.028198
R20627 GNDA.n3486 GNDA.n620 0.028198
R20628 GNDA.n3482 GNDA.n619 0.028198
R20629 GNDA.n3472 GNDA.n617 0.028198
R20630 GNDA.n616 GNDA.n614 0.028198
R20631 GNDA.n3451 GNDA.n638 0.028198
R20632 GNDA.n3447 GNDA.n637 0.028198
R20633 GNDA.n3437 GNDA.n635 0.028198
R20634 GNDA.n3431 GNDA.n634 0.028198
R20635 GNDA.n3421 GNDA.n632 0.028198
R20636 GNDA.n3417 GNDA.n631 0.028198
R20637 GNDA.n3407 GNDA.n629 0.028198
R20638 GNDA.n3401 GNDA.n628 0.028198
R20639 GNDA.n702 GNDA.n701 0.028198
R20640 GNDA.n705 GNDA.n704 0.028198
R20641 GNDA.n711 GNDA.n710 0.028198
R20642 GNDA.n714 GNDA.n713 0.028198
R20643 GNDA.n720 GNDA.n719 0.028198
R20644 GNDA.n723 GNDA.n722 0.028198
R20645 GNDA.n729 GNDA.n728 0.028198
R20646 GNDA.n732 GNDA.n731 0.028198
R20647 GNDA.n853 GNDA.n852 0.028198
R20648 GNDA.n856 GNDA.n855 0.028198
R20649 GNDA.n862 GNDA.n861 0.028198
R20650 GNDA.n865 GNDA.n864 0.028198
R20651 GNDA.n871 GNDA.n870 0.028198
R20652 GNDA.n874 GNDA.n873 0.028198
R20653 GNDA.n880 GNDA.n879 0.028198
R20654 GNDA.n883 GNDA.n882 0.028198
R20655 GNDA.n1031 GNDA.n966 0.028198
R20656 GNDA.n1027 GNDA.n965 0.028198
R20657 GNDA.n1017 GNDA.n963 0.028198
R20658 GNDA.n1011 GNDA.n962 0.028198
R20659 GNDA.n1001 GNDA.n960 0.028198
R20660 GNDA.n997 GNDA.n959 0.028198
R20661 GNDA.n987 GNDA.n957 0.028198
R20662 GNDA.n981 GNDA.n956 0.028198
R20663 GNDA.n1113 GNDA.n1048 0.028198
R20664 GNDA.n1109 GNDA.n1047 0.028198
R20665 GNDA.n1099 GNDA.n1045 0.028198
R20666 GNDA.n1093 GNDA.n1044 0.028198
R20667 GNDA.n1083 GNDA.n1042 0.028198
R20668 GNDA.n1079 GNDA.n1041 0.028198
R20669 GNDA.n1069 GNDA.n1039 0.028198
R20670 GNDA.n1063 GNDA.n1038 0.028198
R20671 GNDA.n1195 GNDA.n1130 0.028198
R20672 GNDA.n1191 GNDA.n1129 0.028198
R20673 GNDA.n1181 GNDA.n1127 0.028198
R20674 GNDA.n1175 GNDA.n1126 0.028198
R20675 GNDA.n1165 GNDA.n1124 0.028198
R20676 GNDA.n1161 GNDA.n1123 0.028198
R20677 GNDA.n1151 GNDA.n1121 0.028198
R20678 GNDA.n1145 GNDA.n1120 0.028198
R20679 GNDA.n949 GNDA.n790 0.028198
R20680 GNDA.n945 GNDA.n789 0.028198
R20681 GNDA.n935 GNDA.n787 0.028198
R20682 GNDA.n929 GNDA.n786 0.028198
R20683 GNDA.n919 GNDA.n784 0.028198
R20684 GNDA.n915 GNDA.n783 0.028198
R20685 GNDA.n905 GNDA.n781 0.028198
R20686 GNDA.n899 GNDA.n780 0.028198
R20687 GNDA.n1277 GNDA.n1212 0.028198
R20688 GNDA.n1273 GNDA.n1211 0.028198
R20689 GNDA.n1263 GNDA.n1209 0.028198
R20690 GNDA.n1257 GNDA.n1208 0.028198
R20691 GNDA.n1247 GNDA.n1206 0.028198
R20692 GNDA.n1243 GNDA.n1205 0.028198
R20693 GNDA.n1233 GNDA.n1203 0.028198
R20694 GNDA.n1227 GNDA.n1202 0.028198
R20695 GNDA.n1359 GNDA.n1294 0.028198
R20696 GNDA.n1355 GNDA.n1293 0.028198
R20697 GNDA.n1345 GNDA.n1291 0.028198
R20698 GNDA.n1339 GNDA.n1290 0.028198
R20699 GNDA.n1329 GNDA.n1288 0.028198
R20700 GNDA.n1325 GNDA.n1287 0.028198
R20701 GNDA.n1315 GNDA.n1285 0.028198
R20702 GNDA.n1309 GNDA.n1284 0.028198
R20703 GNDA.n1435 GNDA.n1375 0.028198
R20704 GNDA.n1431 GNDA.n1374 0.028198
R20705 GNDA.n1421 GNDA.n1372 0.028198
R20706 GNDA.n1415 GNDA.n1371 0.028198
R20707 GNDA.n1405 GNDA.n1369 0.028198
R20708 GNDA.n1401 GNDA.n1368 0.028198
R20709 GNDA.n1391 GNDA.n1366 0.028198
R20710 GNDA.n1365 GNDA.n777 0.028198
R20711 GNDA.n3760 GNDA.n550 0.028198
R20712 GNDA.n3756 GNDA.n549 0.028198
R20713 GNDA.n3746 GNDA.n547 0.028198
R20714 GNDA.n3740 GNDA.n546 0.028198
R20715 GNDA.n3730 GNDA.n544 0.028198
R20716 GNDA.n3726 GNDA.n543 0.028198
R20717 GNDA.n3716 GNDA.n541 0.028198
R20718 GNDA.n3710 GNDA.n540 0.028198
R20719 GNDA.n3836 GNDA.n3776 0.028198
R20720 GNDA.n3832 GNDA.n3775 0.028198
R20721 GNDA.n3822 GNDA.n3773 0.028198
R20722 GNDA.n3816 GNDA.n3772 0.028198
R20723 GNDA.n3806 GNDA.n3770 0.028198
R20724 GNDA.n3802 GNDA.n3769 0.028198
R20725 GNDA.n3792 GNDA.n3767 0.028198
R20726 GNDA.n3766 GNDA.n537 0.028198
R20727 GNDA.n3901 GNDA.n3900 0.028198
R20728 GNDA.n3904 GNDA.n3903 0.028198
R20729 GNDA.n3910 GNDA.n3909 0.028198
R20730 GNDA.n3913 GNDA.n3912 0.028198
R20731 GNDA.n3919 GNDA.n3918 0.028198
R20732 GNDA.n3922 GNDA.n3921 0.028198
R20733 GNDA.n3928 GNDA.n3927 0.028198
R20734 GNDA.n3931 GNDA.n3930 0.028198
R20735 GNDA.n4079 GNDA.n4014 0.028198
R20736 GNDA.n4075 GNDA.n4013 0.028198
R20737 GNDA.n4065 GNDA.n4011 0.028198
R20738 GNDA.n4059 GNDA.n4010 0.028198
R20739 GNDA.n4049 GNDA.n4008 0.028198
R20740 GNDA.n4045 GNDA.n4007 0.028198
R20741 GNDA.n4035 GNDA.n4005 0.028198
R20742 GNDA.n4029 GNDA.n4004 0.028198
R20743 GNDA.n4161 GNDA.n4096 0.028198
R20744 GNDA.n4157 GNDA.n4095 0.028198
R20745 GNDA.n4147 GNDA.n4093 0.028198
R20746 GNDA.n4141 GNDA.n4092 0.028198
R20747 GNDA.n4131 GNDA.n4090 0.028198
R20748 GNDA.n4127 GNDA.n4089 0.028198
R20749 GNDA.n4117 GNDA.n4087 0.028198
R20750 GNDA.n4111 GNDA.n4086 0.028198
R20751 GNDA.n3997 GNDA.n514 0.028198
R20752 GNDA.n3993 GNDA.n513 0.028198
R20753 GNDA.n3983 GNDA.n511 0.028198
R20754 GNDA.n3977 GNDA.n510 0.028198
R20755 GNDA.n3967 GNDA.n508 0.028198
R20756 GNDA.n3963 GNDA.n507 0.028198
R20757 GNDA.n3953 GNDA.n505 0.028198
R20758 GNDA.n3947 GNDA.n504 0.028198
R20759 GNDA.n4243 GNDA.n4178 0.028198
R20760 GNDA.n4239 GNDA.n4177 0.028198
R20761 GNDA.n4229 GNDA.n4175 0.028198
R20762 GNDA.n4223 GNDA.n4174 0.028198
R20763 GNDA.n4213 GNDA.n4172 0.028198
R20764 GNDA.n4209 GNDA.n4171 0.028198
R20765 GNDA.n4199 GNDA.n4169 0.028198
R20766 GNDA.n4193 GNDA.n4168 0.028198
R20767 GNDA.n4325 GNDA.n4260 0.028198
R20768 GNDA.n4321 GNDA.n4259 0.028198
R20769 GNDA.n4311 GNDA.n4257 0.028198
R20770 GNDA.n4305 GNDA.n4256 0.028198
R20771 GNDA.n4295 GNDA.n4254 0.028198
R20772 GNDA.n4291 GNDA.n4253 0.028198
R20773 GNDA.n4281 GNDA.n4251 0.028198
R20774 GNDA.n4275 GNDA.n4250 0.028198
R20775 GNDA.n4407 GNDA.n4342 0.028198
R20776 GNDA.n4403 GNDA.n4341 0.028198
R20777 GNDA.n4393 GNDA.n4339 0.028198
R20778 GNDA.n4387 GNDA.n4338 0.028198
R20779 GNDA.n4377 GNDA.n4336 0.028198
R20780 GNDA.n4373 GNDA.n4335 0.028198
R20781 GNDA.n4363 GNDA.n4333 0.028198
R20782 GNDA.n4357 GNDA.n4332 0.028198
R20783 GNDA.n4489 GNDA.n4424 0.028198
R20784 GNDA.n4485 GNDA.n4423 0.028198
R20785 GNDA.n4475 GNDA.n4421 0.028198
R20786 GNDA.n4469 GNDA.n4420 0.028198
R20787 GNDA.n4459 GNDA.n4418 0.028198
R20788 GNDA.n4455 GNDA.n4417 0.028198
R20789 GNDA.n4445 GNDA.n4415 0.028198
R20790 GNDA.n4439 GNDA.n4414 0.028198
R20791 GNDA.n4565 GNDA.n4505 0.028198
R20792 GNDA.n4561 GNDA.n4504 0.028198
R20793 GNDA.n4551 GNDA.n4502 0.028198
R20794 GNDA.n4545 GNDA.n4501 0.028198
R20795 GNDA.n4535 GNDA.n4499 0.028198
R20796 GNDA.n4531 GNDA.n4498 0.028198
R20797 GNDA.n4521 GNDA.n4496 0.028198
R20798 GNDA.n4495 GNDA.n501 0.028198
R20799 GNDA.n3664 GNDA.n3663 0.028198
R20800 GNDA.n3667 GNDA.n3666 0.028198
R20801 GNDA.n3673 GNDA.n3672 0.028198
R20802 GNDA.n3676 GNDA.n3675 0.028198
R20803 GNDA.n3682 GNDA.n3681 0.028198
R20804 GNDA.n3685 GNDA.n3684 0.028198
R20805 GNDA.n3691 GNDA.n3690 0.028198
R20806 GNDA.n3694 GNDA.n3693 0.028198
R20807 GNDA.n2497 GNDA.n2472 0.028198
R20808 GNDA.n2503 GNDA.n2473 0.028198
R20809 GNDA.n2513 GNDA.n2475 0.028198
R20810 GNDA.n2517 GNDA.n2476 0.028198
R20811 GNDA.n2527 GNDA.n2478 0.028198
R20812 GNDA.n2533 GNDA.n2479 0.028198
R20813 GNDA.n2482 GNDA.n2481 0.028198
R20814 GNDA.n2545 GNDA.n1866 0.028198
R20815 GNDA.n2545 GNDA.n2544 0.028198
R20816 GNDA.n2538 GNDA.n2481 0.028198
R20817 GNDA.n2528 GNDA.n2479 0.028198
R20818 GNDA.n2524 GNDA.n2478 0.028198
R20819 GNDA.n2514 GNDA.n2476 0.028198
R20820 GNDA.n2508 GNDA.n2475 0.028198
R20821 GNDA.n2498 GNDA.n2473 0.028198
R20822 GNDA.n2494 GNDA.n2472 0.028198
R20823 GNDA.n2620 GNDA.n2557 0.028198
R20824 GNDA.n2563 GNDA.n2556 0.028198
R20825 GNDA.n2567 GNDA.n2554 0.028198
R20826 GNDA.n2604 GNDA.n2553 0.028198
R20827 GNDA.n2596 GNDA.n2551 0.028198
R20828 GNDA.n2575 GNDA.n2550 0.028198
R20829 GNDA.n2579 GNDA.n2548 0.028198
R20830 GNDA.n2580 GNDA.n2547 0.028198
R20831 GNDA.n2292 GNDA.n2152 0.028198
R20832 GNDA.n2304 GNDA.n2155 0.028198
R20833 GNDA.n2322 GNDA.n2158 0.028198
R20834 GNDA.n2342 GNDA.n2161 0.028198
R20835 GNDA.n2342 GNDA.n2341 0.028198
R20836 GNDA.n2325 GNDA.n2158 0.028198
R20837 GNDA.n2311 GNDA.n2155 0.028198
R20838 GNDA.n2295 GNDA.n2152 0.028198
R20839 GNDA.n2294 GNDA.n2153 0.0262697
R20840 GNDA.n2302 GNDA.n2154 0.0262697
R20841 GNDA.n2312 GNDA.n2156 0.0262697
R20842 GNDA.n2314 GNDA.n2157 0.0262697
R20843 GNDA.n2324 GNDA.n2159 0.0262697
R20844 GNDA.n2332 GNDA.n2160 0.0262697
R20845 GNDA.n2162 GNDA.n2150 0.0262697
R20846 GNDA.n2334 GNDA.n2160 0.0262697
R20847 GNDA.n2331 GNDA.n2159 0.0262697
R20848 GNDA.n2321 GNDA.n2157 0.0262697
R20849 GNDA.n2315 GNDA.n2156 0.0262697
R20850 GNDA.n2305 GNDA.n2154 0.0262697
R20851 GNDA.n2301 GNDA.n2153 0.0262697
R20852 GNDA.n2291 GNDA.n2151 0.0262697
R20853 GNDA.n2574 GNDA.n2549 0.0243392
R20854 GNDA.n2603 GNDA.n2552 0.0243392
R20855 GNDA.n2562 GNDA.n2555 0.0243392
R20856 GNDA.n3687 GNDA.n3686 0.0243392
R20857 GNDA.n3678 GNDA.n3677 0.0243392
R20858 GNDA.n3669 GNDA.n3668 0.0243392
R20859 GNDA.n4530 GNDA.n4497 0.0243392
R20860 GNDA.n4544 GNDA.n4500 0.0243392
R20861 GNDA.n4560 GNDA.n4503 0.0243392
R20862 GNDA.n4454 GNDA.n4416 0.0243392
R20863 GNDA.n4468 GNDA.n4419 0.0243392
R20864 GNDA.n4484 GNDA.n4422 0.0243392
R20865 GNDA.n4372 GNDA.n4334 0.0243392
R20866 GNDA.n4386 GNDA.n4337 0.0243392
R20867 GNDA.n4402 GNDA.n4340 0.0243392
R20868 GNDA.n4290 GNDA.n4252 0.0243392
R20869 GNDA.n4304 GNDA.n4255 0.0243392
R20870 GNDA.n4320 GNDA.n4258 0.0243392
R20871 GNDA.n4208 GNDA.n4170 0.0243392
R20872 GNDA.n4222 GNDA.n4173 0.0243392
R20873 GNDA.n4238 GNDA.n4176 0.0243392
R20874 GNDA.n3962 GNDA.n506 0.0243392
R20875 GNDA.n3976 GNDA.n509 0.0243392
R20876 GNDA.n3992 GNDA.n512 0.0243392
R20877 GNDA.n4126 GNDA.n4088 0.0243392
R20878 GNDA.n4140 GNDA.n4091 0.0243392
R20879 GNDA.n4156 GNDA.n4094 0.0243392
R20880 GNDA.n4044 GNDA.n4006 0.0243392
R20881 GNDA.n4058 GNDA.n4009 0.0243392
R20882 GNDA.n4074 GNDA.n4012 0.0243392
R20883 GNDA.n3924 GNDA.n3923 0.0243392
R20884 GNDA.n3915 GNDA.n3914 0.0243392
R20885 GNDA.n3906 GNDA.n3905 0.0243392
R20886 GNDA.n3801 GNDA.n3768 0.0243392
R20887 GNDA.n3815 GNDA.n3771 0.0243392
R20888 GNDA.n3831 GNDA.n3774 0.0243392
R20889 GNDA.n3725 GNDA.n542 0.0243392
R20890 GNDA.n3739 GNDA.n545 0.0243392
R20891 GNDA.n3755 GNDA.n548 0.0243392
R20892 GNDA.n1400 GNDA.n1367 0.0243392
R20893 GNDA.n1414 GNDA.n1370 0.0243392
R20894 GNDA.n1430 GNDA.n1373 0.0243392
R20895 GNDA.n1324 GNDA.n1286 0.0243392
R20896 GNDA.n1338 GNDA.n1289 0.0243392
R20897 GNDA.n1354 GNDA.n1292 0.0243392
R20898 GNDA.n1242 GNDA.n1204 0.0243392
R20899 GNDA.n1256 GNDA.n1207 0.0243392
R20900 GNDA.n1272 GNDA.n1210 0.0243392
R20901 GNDA.n914 GNDA.n782 0.0243392
R20902 GNDA.n928 GNDA.n785 0.0243392
R20903 GNDA.n944 GNDA.n788 0.0243392
R20904 GNDA.n1160 GNDA.n1122 0.0243392
R20905 GNDA.n1174 GNDA.n1125 0.0243392
R20906 GNDA.n1190 GNDA.n1128 0.0243392
R20907 GNDA.n1078 GNDA.n1040 0.0243392
R20908 GNDA.n1092 GNDA.n1043 0.0243392
R20909 GNDA.n1108 GNDA.n1046 0.0243392
R20910 GNDA.n996 GNDA.n958 0.0243392
R20911 GNDA.n1010 GNDA.n961 0.0243392
R20912 GNDA.n1026 GNDA.n964 0.0243392
R20913 GNDA.n876 GNDA.n875 0.0243392
R20914 GNDA.n867 GNDA.n866 0.0243392
R20915 GNDA.n858 GNDA.n857 0.0243392
R20916 GNDA.n725 GNDA.n724 0.0243392
R20917 GNDA.n716 GNDA.n715 0.0243392
R20918 GNDA.n707 GNDA.n706 0.0243392
R20919 GNDA.n3416 GNDA.n630 0.0243392
R20920 GNDA.n3430 GNDA.n633 0.0243392
R20921 GNDA.n3446 GNDA.n636 0.0243392
R20922 GNDA.n3481 GNDA.n618 0.0243392
R20923 GNDA.n3495 GNDA.n621 0.0243392
R20924 GNDA.n3511 GNDA.n624 0.0243392
R20925 GNDA.n2248 GNDA.n2247 0.0243392
R20926 GNDA.n2239 GNDA.n2238 0.0243392
R20927 GNDA.n2230 GNDA.n2229 0.0243392
R20928 GNDA.n2231 GNDA.n2230 0.0243392
R20929 GNDA.n2240 GNDA.n2239 0.0243392
R20930 GNDA.n2249 GNDA.n2248 0.0243392
R20931 GNDA.n3506 GNDA.n624 0.0243392
R20932 GNDA.n3492 GNDA.n621 0.0243392
R20933 GNDA.n3476 GNDA.n618 0.0243392
R20934 GNDA.n3441 GNDA.n636 0.0243392
R20935 GNDA.n3427 GNDA.n633 0.0243392
R20936 GNDA.n3411 GNDA.n630 0.0243392
R20937 GNDA.n708 GNDA.n707 0.0243392
R20938 GNDA.n717 GNDA.n716 0.0243392
R20939 GNDA.n726 GNDA.n725 0.0243392
R20940 GNDA.n859 GNDA.n858 0.0243392
R20941 GNDA.n868 GNDA.n867 0.0243392
R20942 GNDA.n877 GNDA.n876 0.0243392
R20943 GNDA.n1021 GNDA.n964 0.0243392
R20944 GNDA.n1007 GNDA.n961 0.0243392
R20945 GNDA.n991 GNDA.n958 0.0243392
R20946 GNDA.n1103 GNDA.n1046 0.0243392
R20947 GNDA.n1089 GNDA.n1043 0.0243392
R20948 GNDA.n1073 GNDA.n1040 0.0243392
R20949 GNDA.n1185 GNDA.n1128 0.0243392
R20950 GNDA.n1171 GNDA.n1125 0.0243392
R20951 GNDA.n1155 GNDA.n1122 0.0243392
R20952 GNDA.n939 GNDA.n788 0.0243392
R20953 GNDA.n925 GNDA.n785 0.0243392
R20954 GNDA.n909 GNDA.n782 0.0243392
R20955 GNDA.n1267 GNDA.n1210 0.0243392
R20956 GNDA.n1253 GNDA.n1207 0.0243392
R20957 GNDA.n1237 GNDA.n1204 0.0243392
R20958 GNDA.n1349 GNDA.n1292 0.0243392
R20959 GNDA.n1335 GNDA.n1289 0.0243392
R20960 GNDA.n1319 GNDA.n1286 0.0243392
R20961 GNDA.n1425 GNDA.n1373 0.0243392
R20962 GNDA.n1411 GNDA.n1370 0.0243392
R20963 GNDA.n1395 GNDA.n1367 0.0243392
R20964 GNDA.n3750 GNDA.n548 0.0243392
R20965 GNDA.n3736 GNDA.n545 0.0243392
R20966 GNDA.n3720 GNDA.n542 0.0243392
R20967 GNDA.n3826 GNDA.n3774 0.0243392
R20968 GNDA.n3812 GNDA.n3771 0.0243392
R20969 GNDA.n3796 GNDA.n3768 0.0243392
R20970 GNDA.n3907 GNDA.n3906 0.0243392
R20971 GNDA.n3916 GNDA.n3915 0.0243392
R20972 GNDA.n3925 GNDA.n3924 0.0243392
R20973 GNDA.n4069 GNDA.n4012 0.0243392
R20974 GNDA.n4055 GNDA.n4009 0.0243392
R20975 GNDA.n4039 GNDA.n4006 0.0243392
R20976 GNDA.n4151 GNDA.n4094 0.0243392
R20977 GNDA.n4137 GNDA.n4091 0.0243392
R20978 GNDA.n4121 GNDA.n4088 0.0243392
R20979 GNDA.n3987 GNDA.n512 0.0243392
R20980 GNDA.n3973 GNDA.n509 0.0243392
R20981 GNDA.n3957 GNDA.n506 0.0243392
R20982 GNDA.n4233 GNDA.n4176 0.0243392
R20983 GNDA.n4219 GNDA.n4173 0.0243392
R20984 GNDA.n4203 GNDA.n4170 0.0243392
R20985 GNDA.n4315 GNDA.n4258 0.0243392
R20986 GNDA.n4301 GNDA.n4255 0.0243392
R20987 GNDA.n4285 GNDA.n4252 0.0243392
R20988 GNDA.n4397 GNDA.n4340 0.0243392
R20989 GNDA.n4383 GNDA.n4337 0.0243392
R20990 GNDA.n4367 GNDA.n4334 0.0243392
R20991 GNDA.n4479 GNDA.n4422 0.0243392
R20992 GNDA.n4465 GNDA.n4419 0.0243392
R20993 GNDA.n4449 GNDA.n4416 0.0243392
R20994 GNDA.n4555 GNDA.n4503 0.0243392
R20995 GNDA.n4541 GNDA.n4500 0.0243392
R20996 GNDA.n4525 GNDA.n4497 0.0243392
R20997 GNDA.n3670 GNDA.n3669 0.0243392
R20998 GNDA.n3679 GNDA.n3678 0.0243392
R20999 GNDA.n3688 GNDA.n3687 0.0243392
R21000 GNDA.n2507 GNDA.n2474 0.0243392
R21001 GNDA.n2523 GNDA.n2477 0.0243392
R21002 GNDA.n2537 GNDA.n2480 0.0243392
R21003 GNDA.n2534 GNDA.n2480 0.0243392
R21004 GNDA.n2518 GNDA.n2477 0.0243392
R21005 GNDA.n2504 GNDA.n2474 0.0243392
R21006 GNDA.n2612 GNDA.n2555 0.0243392
R21007 GNDA.n2571 GNDA.n2552 0.0243392
R21008 GNDA.n2588 GNDA.n2549 0.0243392
R21009 GNDA.n467 GNDA.n466 0.0217373
R21010 GNDA.n471 GNDA.n470 0.0217373
R21011 GNDA.n473 GNDA.n447 0.0217373
R21012 GNDA.n476 GNDA.n446 0.0217373
R21013 GNDA.n475 GNDA.n446 0.0217373
R21014 GNDA.n465 GNDA.n450 0.0217373
R21015 GNDA.n468 GNDA.n467 0.0217373
R21016 GNDA.n3329 GNDA.n3328 0.0217373
R21017 GNDA.n3593 GNDA.n579 0.0217373
R21018 GNDA.n3598 GNDA.n3597 0.0217373
R21019 GNDA.n3600 GNDA.n575 0.0217373
R21020 GNDA.n3596 GNDA.n577 0.0217373
R21021 GNDA.n3599 GNDA.n3598 0.0217373
R21022 GNDA.n3601 GNDA.n576 0.0217373
R21023 GNDA.n3567 GNDA.n589 0.0217373
R21024 GNDA.n3590 GNDA.n3588 0.0217373
R21025 GNDA.n3588 GNDA.n579 0.0217373
R21026 GNDA.n3564 GNDA.n590 0.0217373
R21027 GNDA.n3562 GNDA.n3561 0.0217373
R21028 GNDA.n3559 GNDA.n595 0.0217373
R21029 GNDA.n3332 GNDA.n3330 0.0217373
R21030 GNDA.n3333 GNDA.n3332 0.0217373
R21031 GNDA.n591 GNDA.n589 0.0217373
R21032 GNDA.n3564 GNDA.n3563 0.0217373
R21033 GNDA.n3330 GNDA.n596 0.0217373
R21034 GNDA.n3331 GNDA.n3329 0.0217373
R21035 GNDA.n3545 GNDA.n597 0.0217373
R21036 GNDA.n3561 GNDA.n593 0.0217373
R21037 GNDA.n595 GNDA.n593 0.0217373
R21038 GNDA.n3542 GNDA.n598 0.0217373
R21039 GNDA.n3540 GNDA.n3539 0.0217373
R21040 GNDA.n3537 GNDA.n604 0.0217373
R21041 GNDA.n3530 GNDA.n605 0.0217373
R21042 GNDA.n3531 GNDA.n3530 0.0217373
R21043 GNDA.n599 GNDA.n597 0.0217373
R21044 GNDA.n3542 GNDA.n3541 0.0217373
R21045 GNDA.n3539 GNDA.n601 0.0217373
R21046 GNDA.n604 GNDA.n601 0.0217373
R21047 GNDA.n471 GNDA.n449 0.0217373
R21048 GNDA.n449 GNDA.n447 0.0217373
R21049 GNDA.n2810 GNDA.n2715 0.0217373
R21050 GNDA.n2813 GNDA.n2699 0.0217373
R21051 GNDA.n2714 GNDA.n2701 0.0217373
R21052 GNDA.n2715 GNDA.n2702 0.0217373
R21053 GNDA.n2696 GNDA.n2695 0.0217373
R21054 GNDA.n2699 GNDA.n2695 0.0217373
R21055 GNDA.n2635 GNDA.n2634 0.0217373
R21056 GNDA.n2631 GNDA.n1527 0.0217373
R21057 GNDA.n3228 GNDA.n1525 0.0217373
R21058 GNDA.n3229 GNDA.n1526 0.0217373
R21059 GNDA.n2634 GNDA.n2630 0.0217373
R21060 GNDA.n2631 GNDA.n2630 0.0217373
R21061 GNDA.n3616 GNDA.n569 0.0217373
R21062 GNDA.n3616 GNDA.n567 0.0217373
R21063 GNDA.n4575 GNDA.n497 0.0217373
R21064 GNDA.n4576 GNDA.n497 0.0217373
R21065 GNDA.n495 GNDA.n492 0.0217373
R21066 GNDA.n496 GNDA.n492 0.0217373
R21067 GNDA.n490 GNDA.n487 0.0217373
R21068 GNDA.n491 GNDA.n487 0.0217373
R21069 GNDA.n485 GNDA.n482 0.0217373
R21070 GNDA.n486 GNDA.n482 0.0217373
R21071 GNDA.n480 GNDA.n477 0.0217373
R21072 GNDA.n481 GNDA.n477 0.0217373
R21073 GNDA.n444 GNDA.n441 0.0217373
R21074 GNDA.n445 GNDA.n441 0.0217373
R21075 GNDA.n439 GNDA.n436 0.0217373
R21076 GNDA.n440 GNDA.n436 0.0217373
R21077 GNDA.n534 GNDA.n532 0.0217373
R21078 GNDA.n534 GNDA.n531 0.0217373
R21079 GNDA.n3705 GNDA.n565 0.0217373
R21080 GNDA.n3706 GNDA.n3705 0.0217373
R21081 GNDA.n1446 GNDA.n773 0.0217373
R21082 GNDA.n1444 GNDA.n773 0.0217373
R21083 GNDA.n771 GNDA.n768 0.0217373
R21084 GNDA.n772 GNDA.n768 0.0217373
R21085 GNDA.n766 GNDA.n763 0.0217373
R21086 GNDA.n767 GNDA.n763 0.0217373
R21087 GNDA.n761 GNDA.n758 0.0217373
R21088 GNDA.n762 GNDA.n758 0.0217373
R21089 GNDA.n756 GNDA.n753 0.0217373
R21090 GNDA.n757 GNDA.n753 0.0217373
R21091 GNDA.n751 GNDA.n748 0.0217373
R21092 GNDA.n752 GNDA.n748 0.0217373
R21093 GNDA.n737 GNDA.n653 0.0217373
R21094 GNDA.n738 GNDA.n653 0.0217373
R21095 GNDA.n3396 GNDA.n3393 0.0217373
R21096 GNDA.n3397 GNDA.n3396 0.0217373
R21097 GNDA.n611 GNDA.n609 0.0217373
R21098 GNDA.n611 GNDA.n608 0.0217373
R21099 GNDA.n2261 GNDA.n2176 0.0217373
R21100 GNDA.n2259 GNDA.n2176 0.0217373
R21101 GNDA.n2287 GNDA.n2175 0.0217373
R21102 GNDA.n2280 GNDA.n2268 0.0217373
R21103 GNDA.n2275 GNDA.n2271 0.0217373
R21104 GNDA.n2263 GNDA.n2262 0.0217373
R21105 GNDA.n3526 GNDA.n607 0.0217373
R21106 GNDA.n3533 GNDA.n3532 0.0217373
R21107 GNDA.n3392 GNDA.n652 0.0217373
R21108 GNDA.n3389 GNDA.n3388 0.0217373
R21109 GNDA.n805 GNDA.n804 0.0217373
R21110 GNDA.n3377 GNDA.n3376 0.0217373
R21111 GNDA.n3373 GNDA.n3372 0.0217373
R21112 GNDA.n3369 GNDA.n3368 0.0217373
R21113 GNDA.n1460 GNDA.n1459 0.0217373
R21114 GNDA.n1456 GNDA.n1455 0.0217373
R21115 GNDA.n1448 GNDA.n1447 0.0217373
R21116 GNDA.n3699 GNDA.n566 0.0217373
R21117 GNDA.n564 GNDA.n563 0.0217373
R21118 GNDA.n3846 GNDA.n530 0.0217373
R21119 GNDA.n528 GNDA.n527 0.0217373
R21120 GNDA.n4607 GNDA.n4606 0.0217373
R21121 GNDA.n4603 GNDA.n4602 0.0217373
R21122 GNDA.n4599 GNDA.n4598 0.0217373
R21123 GNDA.n4595 GNDA.n4594 0.0217373
R21124 GNDA.n4591 GNDA.n4590 0.0217373
R21125 GNDA.n4587 GNDA.n4586 0.0217373
R21126 GNDA.n4583 GNDA.n4582 0.0217373
R21127 GNDA.n4579 GNDA.n4578 0.0217373
R21128 GNDA.n2272 GNDA.n2270 0.0217373
R21129 GNDA.n2272 GNDA.n2271 0.0217373
R21130 GNDA.n2277 GNDA.n2267 0.0217373
R21131 GNDA.n2277 GNDA.n2268 0.0217373
R21132 GNDA.n2284 GNDA.n2282 0.0217373
R21133 GNDA.n2282 GNDA.n2175 0.0217373
R21134 GNDA.n2261 GNDA.n2177 0.0217373
R21135 GNDA.n2260 GNDA.n2259 0.0217373
R21136 GNDA.n2264 GNDA.n2263 0.0217373
R21137 GNDA.n3528 GNDA.n609 0.0217373
R21138 GNDA.n3525 GNDA.n608 0.0217373
R21139 GNDA.n3527 GNDA.n3526 0.0217373
R21140 GNDA.n3394 GNDA.n3393 0.0217373
R21141 GNDA.n3398 GNDA.n3397 0.0217373
R21142 GNDA.n3395 GNDA.n652 0.0217373
R21143 GNDA.n737 GNDA.n654 0.0217373
R21144 GNDA.n738 GNDA.n736 0.0217373
R21145 GNDA.n3390 GNDA.n3389 0.0217373
R21146 GNDA.n805 GNDA.n739 0.0217373
R21147 GNDA.n751 GNDA.n749 0.0217373
R21148 GNDA.n752 GNDA.n750 0.0217373
R21149 GNDA.n3378 GNDA.n3377 0.0217373
R21150 GNDA.n756 GNDA.n754 0.0217373
R21151 GNDA.n757 GNDA.n755 0.0217373
R21152 GNDA.n3374 GNDA.n3373 0.0217373
R21153 GNDA.n761 GNDA.n759 0.0217373
R21154 GNDA.n762 GNDA.n760 0.0217373
R21155 GNDA.n3370 GNDA.n3369 0.0217373
R21156 GNDA.n766 GNDA.n764 0.0217373
R21157 GNDA.n767 GNDA.n765 0.0217373
R21158 GNDA.n1461 GNDA.n1460 0.0217373
R21159 GNDA.n771 GNDA.n769 0.0217373
R21160 GNDA.n772 GNDA.n770 0.0217373
R21161 GNDA.n1457 GNDA.n1456 0.0217373
R21162 GNDA.n1446 GNDA.n774 0.0217373
R21163 GNDA.n1445 GNDA.n1444 0.0217373
R21164 GNDA.n1449 GNDA.n1448 0.0217373
R21165 GNDA.n3703 GNDA.n565 0.0217373
R21166 GNDA.n3707 GNDA.n3706 0.0217373
R21167 GNDA.n3704 GNDA.n563 0.0217373
R21168 GNDA.n3848 GNDA.n532 0.0217373
R21169 GNDA.n3845 GNDA.n531 0.0217373
R21170 GNDA.n3847 GNDA.n3846 0.0217373
R21171 GNDA.n439 GNDA.n437 0.0217373
R21172 GNDA.n440 GNDA.n438 0.0217373
R21173 GNDA.n4608 GNDA.n4607 0.0217373
R21174 GNDA.n444 GNDA.n442 0.0217373
R21175 GNDA.n445 GNDA.n443 0.0217373
R21176 GNDA.n4604 GNDA.n4603 0.0217373
R21177 GNDA.n3941 GNDA.n527 0.0217373
R21178 GNDA.n480 GNDA.n478 0.0217373
R21179 GNDA.n481 GNDA.n479 0.0217373
R21180 GNDA.n4596 GNDA.n4595 0.0217373
R21181 GNDA.n485 GNDA.n483 0.0217373
R21182 GNDA.n486 GNDA.n484 0.0217373
R21183 GNDA.n4592 GNDA.n4591 0.0217373
R21184 GNDA.n490 GNDA.n488 0.0217373
R21185 GNDA.n491 GNDA.n489 0.0217373
R21186 GNDA.n4588 GNDA.n4587 0.0217373
R21187 GNDA.n495 GNDA.n493 0.0217373
R21188 GNDA.n496 GNDA.n494 0.0217373
R21189 GNDA.n4584 GNDA.n4583 0.0217373
R21190 GNDA.n4575 GNDA.n498 0.0217373
R21191 GNDA.n4576 GNDA.n4574 0.0217373
R21192 GNDA.n4580 GNDA.n4579 0.0217373
R21193 GNDA.n3535 GNDA.n605 0.0217373
R21194 GNDA.n3534 GNDA.n3533 0.0217373
R21195 GNDA.n476 GNDA.n474 0.0217373
R21196 GNDA.n4600 GNDA.n4599 0.0217373
R21197 GNDA.n3701 GNDA.n569 0.0217373
R21198 GNDA.n3698 GNDA.n567 0.0217373
R21199 GNDA.n3700 GNDA.n3699 0.0217373
R21200 GNDA.n2655 GNDA.n1860 0.0217373
R21201 GNDA.n2648 GNDA.n2647 0.0217373
R21202 GNDA.n2651 GNDA.n1861 0.0217373
R21203 GNDA.n2646 GNDA.n1862 0.0217373
R21204 GNDA.n2649 GNDA.n2648 0.0217373
R21205 GNDA.n2650 GNDA.n1860 0.0217373
R21206 GNDA.n465 GNDA.n464 0.0217373
R21207 GNDA.n466 GNDA.n463 0.0217373
R21208 GNDA.n464 GNDA.n462 0.0217373
R21209 GNDA.n3604 GNDA.n576 0.0217373
R21210 GNDA.n3596 GNDA.n578 0.0217373
R21211 GNDA.n3597 GNDA.n3595 0.0217373
R21212 GNDA.n3602 GNDA.n3600 0.0217373
R21213 GNDA.n3595 GNDA.n3594 0.0217373
R21214 GNDA.n3603 GNDA.n3602 0.0217373
R21215 GNDA.n3605 GNDA.n3604 0.0217373
R21216 GNDA.n3565 GNDA.n591 0.0217373
R21217 GNDA.n3592 GNDA.n3591 0.0217373
R21218 GNDA.n3591 GNDA.n3589 0.0217373
R21219 GNDA.n3566 GNDA.n590 0.0217373
R21220 GNDA.n3543 GNDA.n599 0.0217373
R21221 GNDA.n3558 GNDA.n592 0.0217373
R21222 GNDA.n594 GNDA.n592 0.0217373
R21223 GNDA.n3544 GNDA.n598 0.0217373
R21224 GNDA.n3536 GNDA.n600 0.0217373
R21225 GNDA.n469 GNDA.n434 0.0217373
R21226 GNDA.n602 GNDA.n600 0.0217373
R21227 GNDA.n469 GNDA.n448 0.0217373
R21228 GNDA.n2702 GNDA.n2700 0.0217373
R21229 GNDA.n2811 GNDA.n2701 0.0217373
R21230 GNDA.n2812 GNDA.n2811 0.0217373
R21231 GNDA.n2713 GNDA.n2700 0.0217373
R21232 GNDA.n2814 GNDA.n2697 0.0217373
R21233 GNDA.n3232 GNDA.n1526 0.0217373
R21234 GNDA.n2698 GNDA.n2697 0.0217373
R21235 GNDA.n3230 GNDA.n3228 0.0217373
R21236 GNDA.n3231 GNDA.n3230 0.0217373
R21237 GNDA.n3233 GNDA.n3232 0.0217373
R21238 GNDA.n2629 GNDA.n2624 0.0217373
R21239 GNDA.n2632 GNDA.n2624 0.0217373
R21240 GNDA.n2274 GNDA.n2273 0.0217373
R21241 GNDA.n2279 GNDA.n2278 0.0217373
R21242 GNDA.n2286 GNDA.n2285 0.0217373
R21243 GNDA.n2273 GNDA.n2269 0.0217373
R21244 GNDA.n2278 GNDA.n2266 0.0217373
R21245 GNDA.n2285 GNDA.n2283 0.0217373
R21246 GNDA.n2652 GNDA.n2650 0.0217373
R21247 GNDA.n2646 GNDA.n1863 0.0217373
R21248 GNDA.n2647 GNDA.n2645 0.0217373
R21249 GNDA.n2654 GNDA.n1861 0.0217373
R21250 GNDA.n2645 GNDA.n2644 0.0217373
R21251 GNDA.n2654 GNDA.n2653 0.0217373
R21252 GNDA.n3942 GNDA.n529 0.0181756
R21253 GNDA.n3943 GNDA.n3942 0.0181756
R21254 GNDA.n891 GNDA.n890 0.0181756
R21255 GNDA.n890 GNDA.n888 0.0181756
R21256 GNDA.n892 GNDA.n891 0.0181756
R21257 GNDA.n888 GNDA.n887 0.0181756
R21258 GNDA.n3940 GNDA.n529 0.0181756
R21259 GNDA.n3944 GNDA.n3943 0.0181756
R21260 GNDA.n2343 GNDA.n615 0.0107812
R21261 GNDA.n3521 GNDA.n615 0.0107812
R21262 GNDA.n3521 GNDA.n3456 0.0107812
R21263 GNDA.n3456 GNDA.n639 0.0107812
R21264 GNDA.n778 GNDA.n639 0.0107812
R21265 GNDA.n954 GNDA.n778 0.0107812
R21266 GNDA.n1036 GNDA.n954 0.0107812
R21267 GNDA.n1118 GNDA.n1036 0.0107812
R21268 GNDA.n1200 GNDA.n1118 0.0107812
R21269 GNDA.n1282 GNDA.n1200 0.0107812
R21270 GNDA.n1364 GNDA.n1282 0.0107812
R21271 GNDA.n1440 GNDA.n1364 0.0107812
R21272 GNDA.n1440 GNDA.n538 0.0107812
R21273 GNDA.n3765 GNDA.n538 0.0107812
R21274 GNDA.n3841 GNDA.n3765 0.0107812
R21275 GNDA.n3841 GNDA.n502 0.0107812
R21276 GNDA.n4002 GNDA.n502 0.0107812
R21277 GNDA.n4084 GNDA.n4002 0.0107812
R21278 GNDA.n4166 GNDA.n4084 0.0107812
R21279 GNDA.n4248 GNDA.n4166 0.0107812
R21280 GNDA.n4330 GNDA.n4248 0.0107812
R21281 GNDA.n4412 GNDA.n4330 0.0107812
R21282 GNDA.n4494 GNDA.n4412 0.0107812
R21283 GNDA.n4570 GNDA.n4494 0.0107812
R21284 GNDA.n2377 GNDA.n2084 0.00182188
R21285 GNDA.n2133 GNDA.n2066 0.00182188
R21286 GNDA.n2467 GNDA.n1918 0.00182188
R21287 GNDA.n2425 GNDA.n2409 0.00182188
R21288 GNDA.n2375 GNDA.n2066 0.00166081
R21289 GNDA.n2133 GNDA.n2050 0.00166081
R21290 GNDA.n2373 GNDA.n2135 0.00166081
R21291 GNDA.n2135 GNDA.n2051 0.00166081
R21292 GNDA.n2371 GNDA.n2136 0.00166081
R21293 GNDA.n2136 GNDA.n2052 0.00166081
R21294 GNDA.n2369 GNDA.n2137 0.00166081
R21295 GNDA.n2137 GNDA.n2053 0.00166081
R21296 GNDA.n2367 GNDA.n2138 0.00166081
R21297 GNDA.n2138 GNDA.n2054 0.00166081
R21298 GNDA.n2365 GNDA.n2139 0.00166081
R21299 GNDA.n2139 GNDA.n2055 0.00166081
R21300 GNDA.n2363 GNDA.n2140 0.00166081
R21301 GNDA.n2140 GNDA.n2056 0.00166081
R21302 GNDA.n2361 GNDA.n2141 0.00166081
R21303 GNDA.n2141 GNDA.n2057 0.00166081
R21304 GNDA.n2359 GNDA.n2142 0.00166081
R21305 GNDA.n2142 GNDA.n2058 0.00166081
R21306 GNDA.n2357 GNDA.n2143 0.00166081
R21307 GNDA.n2143 GNDA.n2059 0.00166081
R21308 GNDA.n2355 GNDA.n2144 0.00166081
R21309 GNDA.n2144 GNDA.n2060 0.00166081
R21310 GNDA.n2353 GNDA.n2145 0.00166081
R21311 GNDA.n2145 GNDA.n2061 0.00166081
R21312 GNDA.n2351 GNDA.n2146 0.00166081
R21313 GNDA.n2146 GNDA.n2062 0.00166081
R21314 GNDA.n2349 GNDA.n2147 0.00166081
R21315 GNDA.n2147 GNDA.n2063 0.00166081
R21316 GNDA.n2347 GNDA.n2148 0.00166081
R21317 GNDA.n2148 GNDA.n2064 0.00166081
R21318 GNDA.n2345 GNDA.n2149 0.00166081
R21319 GNDA.n2149 GNDA.n2065 0.00166081
R21320 GNDA.n1918 GNDA.n1885 0.00166081
R21321 GNDA.n2464 GNDA.n1952 0.00166081
R21322 GNDA.n1952 GNDA.n1886 0.00166081
R21323 GNDA.n2462 GNDA.n1953 0.00166081
R21324 GNDA.n1953 GNDA.n1887 0.00166081
R21325 GNDA.n2460 GNDA.n1954 0.00166081
R21326 GNDA.n1954 GNDA.n1888 0.00166081
R21327 GNDA.n2458 GNDA.n1955 0.00166081
R21328 GNDA.n1955 GNDA.n1889 0.00166081
R21329 GNDA.n2456 GNDA.n1956 0.00166081
R21330 GNDA.n1956 GNDA.n1890 0.00166081
R21331 GNDA.n2454 GNDA.n1957 0.00166081
R21332 GNDA.n1957 GNDA.n1891 0.00166081
R21333 GNDA.n2452 GNDA.n1958 0.00166081
R21334 GNDA.n1958 GNDA.n1892 0.00166081
R21335 GNDA.n2450 GNDA.n1959 0.00166081
R21336 GNDA.n1959 GNDA.n1893 0.00166081
R21337 GNDA.n2448 GNDA.n1960 0.00166081
R21338 GNDA.n1960 GNDA.n1894 0.00166081
R21339 GNDA.n2446 GNDA.n1961 0.00166081
R21340 GNDA.n1961 GNDA.n1895 0.00166081
R21341 GNDA.n2444 GNDA.n1962 0.00166081
R21342 GNDA.n1962 GNDA.n1896 0.00166081
R21343 GNDA.n2442 GNDA.n1963 0.00166081
R21344 GNDA.n1963 GNDA.n1897 0.00166081
R21345 GNDA.n2440 GNDA.n1964 0.00166081
R21346 GNDA.n1964 GNDA.n1898 0.00166081
R21347 GNDA.n2438 GNDA.n1965 0.00166081
R21348 GNDA.n1965 GNDA.n1899 0.00166081
R21349 GNDA.n2436 GNDA.n1966 0.00166081
R21350 GNDA.n1966 GNDA.n1900 0.00166081
R21351 GNDA.n2434 GNDA.n1901 0.00166081
R21352 GNDA.n2470 GNDA.n1867 0.00166081
R21353 GNDA.n2469 GNDA.n1884 0.00166081
R21354 GNDA.n1920 GNDA.n1919 0.00166081
R21355 GNDA.n1917 GNDA.n1883 0.00166081
R21356 GNDA.n1922 GNDA.n1921 0.00166081
R21357 GNDA.n1916 GNDA.n1882 0.00166081
R21358 GNDA.n1924 GNDA.n1923 0.00166081
R21359 GNDA.n1915 GNDA.n1881 0.00166081
R21360 GNDA.n1926 GNDA.n1925 0.00166081
R21361 GNDA.n1914 GNDA.n1880 0.00166081
R21362 GNDA.n1928 GNDA.n1927 0.00166081
R21363 GNDA.n1913 GNDA.n1879 0.00166081
R21364 GNDA.n1930 GNDA.n1929 0.00166081
R21365 GNDA.n1912 GNDA.n1878 0.00166081
R21366 GNDA.n1932 GNDA.n1931 0.00166081
R21367 GNDA.n1911 GNDA.n1877 0.00166081
R21368 GNDA.n1934 GNDA.n1933 0.00166081
R21369 GNDA.n1910 GNDA.n1876 0.00166081
R21370 GNDA.n1936 GNDA.n1935 0.00166081
R21371 GNDA.n1909 GNDA.n1875 0.00166081
R21372 GNDA.n1938 GNDA.n1937 0.00166081
R21373 GNDA.n1908 GNDA.n1874 0.00166081
R21374 GNDA.n1940 GNDA.n1939 0.00166081
R21375 GNDA.n1907 GNDA.n1873 0.00166081
R21376 GNDA.n1942 GNDA.n1941 0.00166081
R21377 GNDA.n1906 GNDA.n1872 0.00166081
R21378 GNDA.n1944 GNDA.n1943 0.00166081
R21379 GNDA.n1905 GNDA.n1871 0.00166081
R21380 GNDA.n1946 GNDA.n1945 0.00166081
R21381 GNDA.n1904 GNDA.n1870 0.00166081
R21382 GNDA.n1948 GNDA.n1947 0.00166081
R21383 GNDA.n1903 GNDA.n1869 0.00166081
R21384 GNDA.n1950 GNDA.n1949 0.00166081
R21385 GNDA.n1902 GNDA.n1868 0.00166081
R21386 GNDA.n2466 GNDA.n1951 0.00166081
R21387 GNDA.n2433 GNDA.n2432 0.00166081
R21388 GNDA.n2428 GNDA.n2426 0.00166081
R21389 GNDA.n2427 GNDA.n2000 0.00166081
R21390 GNDA.n2410 GNDA.n2002 0.00166081
R21391 GNDA.n2032 GNDA.n1999 0.00166081
R21392 GNDA.n2411 GNDA.n2003 0.00166081
R21393 GNDA.n2031 GNDA.n1998 0.00166081
R21394 GNDA.n2412 GNDA.n2004 0.00166081
R21395 GNDA.n2030 GNDA.n1997 0.00166081
R21396 GNDA.n2413 GNDA.n2005 0.00166081
R21397 GNDA.n2029 GNDA.n1996 0.00166081
R21398 GNDA.n2414 GNDA.n2006 0.00166081
R21399 GNDA.n2028 GNDA.n1995 0.00166081
R21400 GNDA.n2415 GNDA.n2007 0.00166081
R21401 GNDA.n2027 GNDA.n1994 0.00166081
R21402 GNDA.n2416 GNDA.n2008 0.00166081
R21403 GNDA.n2026 GNDA.n1993 0.00166081
R21404 GNDA.n2417 GNDA.n2009 0.00166081
R21405 GNDA.n2025 GNDA.n1992 0.00166081
R21406 GNDA.n2418 GNDA.n2010 0.00166081
R21407 GNDA.n2024 GNDA.n1991 0.00166081
R21408 GNDA.n2419 GNDA.n2011 0.00166081
R21409 GNDA.n2023 GNDA.n1990 0.00166081
R21410 GNDA.n2420 GNDA.n2012 0.00166081
R21411 GNDA.n2022 GNDA.n1989 0.00166081
R21412 GNDA.n2421 GNDA.n2013 0.00166081
R21413 GNDA.n2021 GNDA.n1988 0.00166081
R21414 GNDA.n2422 GNDA.n2014 0.00166081
R21415 GNDA.n2020 GNDA.n1987 0.00166081
R21416 GNDA.n2423 GNDA.n2015 0.00166081
R21417 GNDA.n2019 GNDA.n1986 0.00166081
R21418 GNDA.n2424 GNDA.n2016 0.00166081
R21419 GNDA.n2018 GNDA.n1985 0.00166081
R21420 GNDA.n2430 GNDA.n2017 0.00166081
R21421 GNDA.n2083 GNDA.n2049 0.00166081
R21422 GNDA.n2117 GNDA.n2086 0.00166081
R21423 GNDA.n2085 GNDA.n2082 0.00166081
R21424 GNDA.n2118 GNDA.n2088 0.00166081
R21425 GNDA.n2087 GNDA.n2081 0.00166081
R21426 GNDA.n2119 GNDA.n2090 0.00166081
R21427 GNDA.n2089 GNDA.n2080 0.00166081
R21428 GNDA.n2120 GNDA.n2092 0.00166081
R21429 GNDA.n2091 GNDA.n2079 0.00166081
R21430 GNDA.n2121 GNDA.n2094 0.00166081
R21431 GNDA.n2093 GNDA.n2078 0.00166081
R21432 GNDA.n2122 GNDA.n2096 0.00166081
R21433 GNDA.n2095 GNDA.n2077 0.00166081
R21434 GNDA.n2123 GNDA.n2098 0.00166081
R21435 GNDA.n2097 GNDA.n2076 0.00166081
R21436 GNDA.n2124 GNDA.n2100 0.00166081
R21437 GNDA.n2099 GNDA.n2075 0.00166081
R21438 GNDA.n2125 GNDA.n2102 0.00166081
R21439 GNDA.n2101 GNDA.n2074 0.00166081
R21440 GNDA.n2126 GNDA.n2104 0.00166081
R21441 GNDA.n2103 GNDA.n2073 0.00166081
R21442 GNDA.n2127 GNDA.n2106 0.00166081
R21443 GNDA.n2105 GNDA.n2072 0.00166081
R21444 GNDA.n2128 GNDA.n2108 0.00166081
R21445 GNDA.n2107 GNDA.n2071 0.00166081
R21446 GNDA.n2129 GNDA.n2110 0.00166081
R21447 GNDA.n2109 GNDA.n2070 0.00166081
R21448 GNDA.n2130 GNDA.n2112 0.00166081
R21449 GNDA.n2111 GNDA.n2069 0.00166081
R21450 GNDA.n2131 GNDA.n2114 0.00166081
R21451 GNDA.n2113 GNDA.n2068 0.00166081
R21452 GNDA.n2132 GNDA.n2116 0.00166081
R21453 GNDA.n2115 GNDA.n2067 0.00166081
R21454 GNDA.n2376 GNDA.n2134 0.00166081
R21455 GNDA.n2469 GNDA.n2468 0.00166081
R21456 GNDA.n2435 GNDA.n1900 0.00166081
R21457 GNDA.n2437 GNDA.n1899 0.00166081
R21458 GNDA.n2439 GNDA.n1898 0.00166081
R21459 GNDA.n2441 GNDA.n1897 0.00166081
R21460 GNDA.n2443 GNDA.n1896 0.00166081
R21461 GNDA.n2445 GNDA.n1895 0.00166081
R21462 GNDA.n2447 GNDA.n1894 0.00166081
R21463 GNDA.n2449 GNDA.n1893 0.00166081
R21464 GNDA.n2451 GNDA.n1892 0.00166081
R21465 GNDA.n2453 GNDA.n1891 0.00166081
R21466 GNDA.n2455 GNDA.n1890 0.00166081
R21467 GNDA.n2457 GNDA.n1889 0.00166081
R21468 GNDA.n2459 GNDA.n1888 0.00166081
R21469 GNDA.n2461 GNDA.n1887 0.00166081
R21470 GNDA.n2463 GNDA.n1886 0.00166081
R21471 GNDA.n2465 GNDA.n1885 0.00166081
R21472 GNDA.n2435 GNDA.n2434 0.00166081
R21473 GNDA.n2437 GNDA.n2436 0.00166081
R21474 GNDA.n2439 GNDA.n2438 0.00166081
R21475 GNDA.n2441 GNDA.n2440 0.00166081
R21476 GNDA.n2443 GNDA.n2442 0.00166081
R21477 GNDA.n2445 GNDA.n2444 0.00166081
R21478 GNDA.n2447 GNDA.n2446 0.00166081
R21479 GNDA.n2449 GNDA.n2448 0.00166081
R21480 GNDA.n2451 GNDA.n2450 0.00166081
R21481 GNDA.n2453 GNDA.n2452 0.00166081
R21482 GNDA.n2455 GNDA.n2454 0.00166081
R21483 GNDA.n2457 GNDA.n2456 0.00166081
R21484 GNDA.n2459 GNDA.n2458 0.00166081
R21485 GNDA.n2461 GNDA.n2460 0.00166081
R21486 GNDA.n2463 GNDA.n2462 0.00166081
R21487 GNDA.n2465 GNDA.n2464 0.00166081
R21488 GNDA.n1919 GNDA.n1884 0.00166081
R21489 GNDA.n1920 GNDA.n1883 0.00166081
R21490 GNDA.n1921 GNDA.n1917 0.00166081
R21491 GNDA.n1922 GNDA.n1882 0.00166081
R21492 GNDA.n1923 GNDA.n1916 0.00166081
R21493 GNDA.n1924 GNDA.n1881 0.00166081
R21494 GNDA.n1925 GNDA.n1915 0.00166081
R21495 GNDA.n1926 GNDA.n1880 0.00166081
R21496 GNDA.n1927 GNDA.n1914 0.00166081
R21497 GNDA.n1928 GNDA.n1879 0.00166081
R21498 GNDA.n1929 GNDA.n1913 0.00166081
R21499 GNDA.n1930 GNDA.n1878 0.00166081
R21500 GNDA.n1931 GNDA.n1912 0.00166081
R21501 GNDA.n1932 GNDA.n1877 0.00166081
R21502 GNDA.n1933 GNDA.n1911 0.00166081
R21503 GNDA.n1934 GNDA.n1876 0.00166081
R21504 GNDA.n1935 GNDA.n1910 0.00166081
R21505 GNDA.n1936 GNDA.n1875 0.00166081
R21506 GNDA.n1937 GNDA.n1909 0.00166081
R21507 GNDA.n1938 GNDA.n1874 0.00166081
R21508 GNDA.n1939 GNDA.n1908 0.00166081
R21509 GNDA.n1940 GNDA.n1873 0.00166081
R21510 GNDA.n1941 GNDA.n1907 0.00166081
R21511 GNDA.n1942 GNDA.n1872 0.00166081
R21512 GNDA.n1943 GNDA.n1906 0.00166081
R21513 GNDA.n1944 GNDA.n1871 0.00166081
R21514 GNDA.n1945 GNDA.n1905 0.00166081
R21515 GNDA.n1946 GNDA.n1870 0.00166081
R21516 GNDA.n1947 GNDA.n1904 0.00166081
R21517 GNDA.n1948 GNDA.n1869 0.00166081
R21518 GNDA.n1949 GNDA.n1903 0.00166081
R21519 GNDA.n1950 GNDA.n1868 0.00166081
R21520 GNDA.n1951 GNDA.n1902 0.00166081
R21521 GNDA.n1901 GNDA.n1867 0.00166081
R21522 GNDA.n2344 GNDA.n2065 0.00166081
R21523 GNDA.n2346 GNDA.n2064 0.00166081
R21524 GNDA.n2348 GNDA.n2063 0.00166081
R21525 GNDA.n2350 GNDA.n2062 0.00166081
R21526 GNDA.n2352 GNDA.n2061 0.00166081
R21527 GNDA.n2354 GNDA.n2060 0.00166081
R21528 GNDA.n2356 GNDA.n2059 0.00166081
R21529 GNDA.n2358 GNDA.n2058 0.00166081
R21530 GNDA.n2360 GNDA.n2057 0.00166081
R21531 GNDA.n2362 GNDA.n2056 0.00166081
R21532 GNDA.n2364 GNDA.n2055 0.00166081
R21533 GNDA.n2366 GNDA.n2054 0.00166081
R21534 GNDA.n2368 GNDA.n2053 0.00166081
R21535 GNDA.n2370 GNDA.n2052 0.00166081
R21536 GNDA.n2372 GNDA.n2051 0.00166081
R21537 GNDA.n2374 GNDA.n2050 0.00166081
R21538 GNDA.n2378 GNDA.n2049 0.00166081
R21539 GNDA.n2346 GNDA.n2345 0.00166081
R21540 GNDA.n2348 GNDA.n2347 0.00166081
R21541 GNDA.n2350 GNDA.n2349 0.00166081
R21542 GNDA.n2352 GNDA.n2351 0.00166081
R21543 GNDA.n2354 GNDA.n2353 0.00166081
R21544 GNDA.n2356 GNDA.n2355 0.00166081
R21545 GNDA.n2358 GNDA.n2357 0.00166081
R21546 GNDA.n2360 GNDA.n2359 0.00166081
R21547 GNDA.n2362 GNDA.n2361 0.00166081
R21548 GNDA.n2364 GNDA.n2363 0.00166081
R21549 GNDA.n2366 GNDA.n2365 0.00166081
R21550 GNDA.n2368 GNDA.n2367 0.00166081
R21551 GNDA.n2370 GNDA.n2369 0.00166081
R21552 GNDA.n2372 GNDA.n2371 0.00166081
R21553 GNDA.n2374 GNDA.n2373 0.00166081
R21554 GNDA.n2117 GNDA.n2083 0.00166081
R21555 GNDA.n2086 GNDA.n2085 0.00166081
R21556 GNDA.n2118 GNDA.n2082 0.00166081
R21557 GNDA.n2088 GNDA.n2087 0.00166081
R21558 GNDA.n2119 GNDA.n2081 0.00166081
R21559 GNDA.n2090 GNDA.n2089 0.00166081
R21560 GNDA.n2120 GNDA.n2080 0.00166081
R21561 GNDA.n2092 GNDA.n2091 0.00166081
R21562 GNDA.n2121 GNDA.n2079 0.00166081
R21563 GNDA.n2094 GNDA.n2093 0.00166081
R21564 GNDA.n2122 GNDA.n2078 0.00166081
R21565 GNDA.n2096 GNDA.n2095 0.00166081
R21566 GNDA.n2123 GNDA.n2077 0.00166081
R21567 GNDA.n2098 GNDA.n2097 0.00166081
R21568 GNDA.n2124 GNDA.n2076 0.00166081
R21569 GNDA.n2100 GNDA.n2099 0.00166081
R21570 GNDA.n2125 GNDA.n2075 0.00166081
R21571 GNDA.n2102 GNDA.n2101 0.00166081
R21572 GNDA.n2126 GNDA.n2074 0.00166081
R21573 GNDA.n2104 GNDA.n2103 0.00166081
R21574 GNDA.n2127 GNDA.n2073 0.00166081
R21575 GNDA.n2106 GNDA.n2105 0.00166081
R21576 GNDA.n2128 GNDA.n2072 0.00166081
R21577 GNDA.n2108 GNDA.n2107 0.00166081
R21578 GNDA.n2129 GNDA.n2071 0.00166081
R21579 GNDA.n2110 GNDA.n2109 0.00166081
R21580 GNDA.n2130 GNDA.n2070 0.00166081
R21581 GNDA.n2112 GNDA.n2111 0.00166081
R21582 GNDA.n2131 GNDA.n2069 0.00166081
R21583 GNDA.n2114 GNDA.n2113 0.00166081
R21584 GNDA.n2132 GNDA.n2068 0.00166081
R21585 GNDA.n2116 GNDA.n2115 0.00166081
R21586 GNDA.n2134 GNDA.n2067 0.00166081
R21587 GNDA.n2375 GNDA.n2084 0.00166081
R21588 GNDA.n2429 GNDA.n1967 0.00166081
R21589 GNDA.n2409 GNDA.n1968 0.00166081
R21590 GNDA.n2407 GNDA.n2033 0.00166081
R21591 GNDA.n2408 GNDA.n1969 0.00166081
R21592 GNDA.n2405 GNDA.n2034 0.00166081
R21593 GNDA.n2406 GNDA.n1970 0.00166081
R21594 GNDA.n2403 GNDA.n2035 0.00166081
R21595 GNDA.n2404 GNDA.n1971 0.00166081
R21596 GNDA.n2401 GNDA.n2036 0.00166081
R21597 GNDA.n2402 GNDA.n1972 0.00166081
R21598 GNDA.n2399 GNDA.n2037 0.00166081
R21599 GNDA.n2400 GNDA.n1973 0.00166081
R21600 GNDA.n2397 GNDA.n2038 0.00166081
R21601 GNDA.n2398 GNDA.n1974 0.00166081
R21602 GNDA.n2395 GNDA.n2039 0.00166081
R21603 GNDA.n2396 GNDA.n1975 0.00166081
R21604 GNDA.n2393 GNDA.n2040 0.00166081
R21605 GNDA.n2394 GNDA.n1976 0.00166081
R21606 GNDA.n2391 GNDA.n2041 0.00166081
R21607 GNDA.n2392 GNDA.n1977 0.00166081
R21608 GNDA.n2389 GNDA.n2042 0.00166081
R21609 GNDA.n2390 GNDA.n1978 0.00166081
R21610 GNDA.n2387 GNDA.n2043 0.00166081
R21611 GNDA.n2388 GNDA.n1979 0.00166081
R21612 GNDA.n2385 GNDA.n2044 0.00166081
R21613 GNDA.n2386 GNDA.n1980 0.00166081
R21614 GNDA.n2383 GNDA.n2045 0.00166081
R21615 GNDA.n2384 GNDA.n1981 0.00166081
R21616 GNDA.n2381 GNDA.n2046 0.00166081
R21617 GNDA.n2382 GNDA.n1982 0.00166081
R21618 GNDA.n2379 GNDA.n2047 0.00166081
R21619 GNDA.n2380 GNDA.n1983 0.00166081
R21620 GNDA.n2048 GNDA.n2001 0.00166081
R21621 GNDA.n2048 GNDA.n1983 0.00166081
R21622 GNDA.n2047 GNDA.n1982 0.00166081
R21623 GNDA.n2046 GNDA.n1981 0.00166081
R21624 GNDA.n2045 GNDA.n1980 0.00166081
R21625 GNDA.n2044 GNDA.n1979 0.00166081
R21626 GNDA.n2043 GNDA.n1978 0.00166081
R21627 GNDA.n2042 GNDA.n1977 0.00166081
R21628 GNDA.n2041 GNDA.n1976 0.00166081
R21629 GNDA.n2040 GNDA.n1975 0.00166081
R21630 GNDA.n2039 GNDA.n1974 0.00166081
R21631 GNDA.n2038 GNDA.n1973 0.00166081
R21632 GNDA.n2037 GNDA.n1972 0.00166081
R21633 GNDA.n2036 GNDA.n1971 0.00166081
R21634 GNDA.n2035 GNDA.n1970 0.00166081
R21635 GNDA.n2034 GNDA.n1969 0.00166081
R21636 GNDA.n2033 GNDA.n1968 0.00166081
R21637 GNDA.n2425 GNDA.n1967 0.00166081
R21638 GNDA.n2432 GNDA.n1984 0.00166081
R21639 GNDA.n2380 GNDA.n2379 0.00166081
R21640 GNDA.n2382 GNDA.n2381 0.00166081
R21641 GNDA.n2384 GNDA.n2383 0.00166081
R21642 GNDA.n2386 GNDA.n2385 0.00166081
R21643 GNDA.n2388 GNDA.n2387 0.00166081
R21644 GNDA.n2390 GNDA.n2389 0.00166081
R21645 GNDA.n2392 GNDA.n2391 0.00166081
R21646 GNDA.n2394 GNDA.n2393 0.00166081
R21647 GNDA.n2396 GNDA.n2395 0.00166081
R21648 GNDA.n2398 GNDA.n2397 0.00166081
R21649 GNDA.n2400 GNDA.n2399 0.00166081
R21650 GNDA.n2402 GNDA.n2401 0.00166081
R21651 GNDA.n2404 GNDA.n2403 0.00166081
R21652 GNDA.n2406 GNDA.n2405 0.00166081
R21653 GNDA.n2408 GNDA.n2407 0.00166081
R21654 GNDA.n2426 GNDA.n1984 0.00166081
R21655 GNDA.n2431 GNDA.n2001 0.00166081
R21656 GNDA.n2428 GNDA.n2427 0.00166081
R21657 GNDA.n2410 GNDA.n2000 0.00166081
R21658 GNDA.n2032 GNDA.n2002 0.00166081
R21659 GNDA.n2411 GNDA.n1999 0.00166081
R21660 GNDA.n2031 GNDA.n2003 0.00166081
R21661 GNDA.n2412 GNDA.n1998 0.00166081
R21662 GNDA.n2030 GNDA.n2004 0.00166081
R21663 GNDA.n2413 GNDA.n1997 0.00166081
R21664 GNDA.n2029 GNDA.n2005 0.00166081
R21665 GNDA.n2414 GNDA.n1996 0.00166081
R21666 GNDA.n2028 GNDA.n2006 0.00166081
R21667 GNDA.n2415 GNDA.n1995 0.00166081
R21668 GNDA.n2027 GNDA.n2007 0.00166081
R21669 GNDA.n2416 GNDA.n1994 0.00166081
R21670 GNDA.n2026 GNDA.n2008 0.00166081
R21671 GNDA.n2417 GNDA.n1993 0.00166081
R21672 GNDA.n2025 GNDA.n2009 0.00166081
R21673 GNDA.n2418 GNDA.n1992 0.00166081
R21674 GNDA.n2024 GNDA.n2010 0.00166081
R21675 GNDA.n2419 GNDA.n1991 0.00166081
R21676 GNDA.n2023 GNDA.n2011 0.00166081
R21677 GNDA.n2420 GNDA.n1990 0.00166081
R21678 GNDA.n2022 GNDA.n2012 0.00166081
R21679 GNDA.n2421 GNDA.n1989 0.00166081
R21680 GNDA.n2021 GNDA.n2013 0.00166081
R21681 GNDA.n2422 GNDA.n1988 0.00166081
R21682 GNDA.n2020 GNDA.n2014 0.00166081
R21683 GNDA.n2423 GNDA.n1987 0.00166081
R21684 GNDA.n2019 GNDA.n2015 0.00166081
R21685 GNDA.n2424 GNDA.n1986 0.00166081
R21686 GNDA.n2018 GNDA.n2016 0.00166081
R21687 GNDA.n2017 GNDA.n1985 0.00166081
R21688 two_stage_opamp_dummy_magic_24_0.Vb2.n0 two_stage_opamp_dummy_magic_24_0.Vb2.t20 752.422
R21689 two_stage_opamp_dummy_magic_24_0.Vb2.n3 two_stage_opamp_dummy_magic_24_0.Vb2.t15 752.422
R21690 two_stage_opamp_dummy_magic_24_0.Vb2.n0 two_stage_opamp_dummy_magic_24_0.Vb2.t16 752.234
R21691 two_stage_opamp_dummy_magic_24_0.Vb2.n0 two_stage_opamp_dummy_magic_24_0.Vb2.t22 752.234
R21692 two_stage_opamp_dummy_magic_24_0.Vb2.n1 two_stage_opamp_dummy_magic_24_0.Vb2.t26 752.234
R21693 two_stage_opamp_dummy_magic_24_0.Vb2.n1 two_stage_opamp_dummy_magic_24_0.Vb2.t28 752.234
R21694 two_stage_opamp_dummy_magic_24_0.Vb2.n1 two_stage_opamp_dummy_magic_24_0.Vb2.t30 752.234
R21695 two_stage_opamp_dummy_magic_24_0.Vb2.n1 two_stage_opamp_dummy_magic_24_0.Vb2.t14 752.234
R21696 two_stage_opamp_dummy_magic_24_0.Vb2.n2 two_stage_opamp_dummy_magic_24_0.Vb2.t18 752.234
R21697 two_stage_opamp_dummy_magic_24_0.Vb2.n2 two_stage_opamp_dummy_magic_24_0.Vb2.t24 752.234
R21698 two_stage_opamp_dummy_magic_24_0.Vb2.n2 two_stage_opamp_dummy_magic_24_0.Vb2.t27 752.234
R21699 two_stage_opamp_dummy_magic_24_0.Vb2.n5 two_stage_opamp_dummy_magic_24_0.Vb2.t12 752.234
R21700 two_stage_opamp_dummy_magic_24_0.Vb2.n5 two_stage_opamp_dummy_magic_24_0.Vb2.t17 752.234
R21701 two_stage_opamp_dummy_magic_24_0.Vb2.n4 two_stage_opamp_dummy_magic_24_0.Vb2.t23 752.234
R21702 two_stage_opamp_dummy_magic_24_0.Vb2.n4 two_stage_opamp_dummy_magic_24_0.Vb2.t19 752.234
R21703 two_stage_opamp_dummy_magic_24_0.Vb2.n4 two_stage_opamp_dummy_magic_24_0.Vb2.t25 752.234
R21704 two_stage_opamp_dummy_magic_24_0.Vb2.n4 two_stage_opamp_dummy_magic_24_0.Vb2.t29 752.234
R21705 two_stage_opamp_dummy_magic_24_0.Vb2.n3 two_stage_opamp_dummy_magic_24_0.Vb2.t32 752.234
R21706 two_stage_opamp_dummy_magic_24_0.Vb2.n3 two_stage_opamp_dummy_magic_24_0.Vb2.t13 752.234
R21707 two_stage_opamp_dummy_magic_24_0.Vb2.n3 two_stage_opamp_dummy_magic_24_0.Vb2.t11 752.234
R21708 two_stage_opamp_dummy_magic_24_0.Vb2.n13 two_stage_opamp_dummy_magic_24_0.Vb2.t21 746.673
R21709 two_stage_opamp_dummy_magic_24_0.Vb2.n17 two_stage_opamp_dummy_magic_24_0.Vb2.t4 721.625
R21710 two_stage_opamp_dummy_magic_24_0.Vb2.n16 two_stage_opamp_dummy_magic_24_0.Vb2.t31 563.451
R21711 two_stage_opamp_dummy_magic_24_0.Vb2.n8 two_stage_opamp_dummy_magic_24_0.Vb2.n6 140.546
R21712 two_stage_opamp_dummy_magic_24_0.Vb2.n12 two_stage_opamp_dummy_magic_24_0.Vb2.n11 139.297
R21713 two_stage_opamp_dummy_magic_24_0.Vb2.n10 two_stage_opamp_dummy_magic_24_0.Vb2.n9 139.297
R21714 two_stage_opamp_dummy_magic_24_0.Vb2.n8 two_stage_opamp_dummy_magic_24_0.Vb2.n7 139.297
R21715 two_stage_opamp_dummy_magic_24_0.Vb2.n13 two_stage_opamp_dummy_magic_24_0.Vb2.n12 84.1349
R21716 two_stage_opamp_dummy_magic_24_0.Vb2.n18 two_stage_opamp_dummy_magic_24_0.Vb2.n17 67.013
R21717 two_stage_opamp_dummy_magic_24_0.Vb2.n11 two_stage_opamp_dummy_magic_24_0.Vb2.t3 24.0005
R21718 two_stage_opamp_dummy_magic_24_0.Vb2.n11 two_stage_opamp_dummy_magic_24_0.Vb2.t7 24.0005
R21719 two_stage_opamp_dummy_magic_24_0.Vb2.n9 two_stage_opamp_dummy_magic_24_0.Vb2.t8 24.0005
R21720 two_stage_opamp_dummy_magic_24_0.Vb2.n9 two_stage_opamp_dummy_magic_24_0.Vb2.t6 24.0005
R21721 two_stage_opamp_dummy_magic_24_0.Vb2.n7 two_stage_opamp_dummy_magic_24_0.Vb2.t9 24.0005
R21722 two_stage_opamp_dummy_magic_24_0.Vb2.n7 two_stage_opamp_dummy_magic_24_0.Vb2.t0 24.0005
R21723 two_stage_opamp_dummy_magic_24_0.Vb2.n6 two_stage_opamp_dummy_magic_24_0.Vb2.t10 24.0005
R21724 two_stage_opamp_dummy_magic_24_0.Vb2.n6 two_stage_opamp_dummy_magic_24_0.Vb2.t2 24.0005
R21725 two_stage_opamp_dummy_magic_24_0.Vb2.n15 two_stage_opamp_dummy_magic_24_0.Vb2.n14 15.188
R21726 two_stage_opamp_dummy_magic_24_0.Vb2.n18 two_stage_opamp_dummy_magic_24_0.Vb2.t5 11.2576
R21727 two_stage_opamp_dummy_magic_24_0.Vb2.t1 two_stage_opamp_dummy_magic_24_0.Vb2.n18 11.2576
R21728 two_stage_opamp_dummy_magic_24_0.Vb2.n17 two_stage_opamp_dummy_magic_24_0.Vb2.n16 7.35988
R21729 two_stage_opamp_dummy_magic_24_0.Vb2.n10 two_stage_opamp_dummy_magic_24_0.Vb2.n8 5.8755
R21730 two_stage_opamp_dummy_magic_24_0.Vb2.n15 two_stage_opamp_dummy_magic_24_0.Vb2.n13 4.55362
R21731 two_stage_opamp_dummy_magic_24_0.Vb2.n12 two_stage_opamp_dummy_magic_24_0.Vb2.n10 1.2505
R21732 two_stage_opamp_dummy_magic_24_0.Vb2.n16 two_stage_opamp_dummy_magic_24_0.Vb2.n15 1.14112
R21733 two_stage_opamp_dummy_magic_24_0.Vb2.n14 two_stage_opamp_dummy_magic_24_0.Vb2.n5 0.90675
R21734 two_stage_opamp_dummy_magic_24_0.Vb2.n4 two_stage_opamp_dummy_magic_24_0.Vb2.n3 0.7505
R21735 two_stage_opamp_dummy_magic_24_0.Vb2.n5 two_stage_opamp_dummy_magic_24_0.Vb2.n4 0.7505
R21736 two_stage_opamp_dummy_magic_24_0.Vb2.n2 two_stage_opamp_dummy_magic_24_0.Vb2.n1 0.7505
R21737 two_stage_opamp_dummy_magic_24_0.Vb2.n1 two_stage_opamp_dummy_magic_24_0.Vb2.n0 0.7505
R21738 two_stage_opamp_dummy_magic_24_0.Vb2.n14 two_stage_opamp_dummy_magic_24_0.Vb2.n2 0.6255
R21739 two_stage_opamp_dummy_magic_24_0.X.n43 two_stage_opamp_dummy_magic_24_0.X.t51 1172.87
R21740 two_stage_opamp_dummy_magic_24_0.X.n39 two_stage_opamp_dummy_magic_24_0.X.t46 1172.87
R21741 two_stage_opamp_dummy_magic_24_0.X.n43 two_stage_opamp_dummy_magic_24_0.X.t38 996.134
R21742 two_stage_opamp_dummy_magic_24_0.X.n44 two_stage_opamp_dummy_magic_24_0.X.t26 996.134
R21743 two_stage_opamp_dummy_magic_24_0.X.n45 two_stage_opamp_dummy_magic_24_0.X.t37 996.134
R21744 two_stage_opamp_dummy_magic_24_0.X.n46 two_stage_opamp_dummy_magic_24_0.X.t25 996.134
R21745 two_stage_opamp_dummy_magic_24_0.X.n42 two_stage_opamp_dummy_magic_24_0.X.t41 996.134
R21746 two_stage_opamp_dummy_magic_24_0.X.n41 two_stage_opamp_dummy_magic_24_0.X.t29 996.134
R21747 two_stage_opamp_dummy_magic_24_0.X.n40 two_stage_opamp_dummy_magic_24_0.X.t44 996.134
R21748 two_stage_opamp_dummy_magic_24_0.X.n39 two_stage_opamp_dummy_magic_24_0.X.t31 996.134
R21749 two_stage_opamp_dummy_magic_24_0.X.n10 two_stage_opamp_dummy_magic_24_0.X.t47 690.867
R21750 two_stage_opamp_dummy_magic_24_0.X.n9 two_stage_opamp_dummy_magic_24_0.X.t43 690.867
R21751 two_stage_opamp_dummy_magic_24_0.X.n19 two_stage_opamp_dummy_magic_24_0.X.t48 530.201
R21752 two_stage_opamp_dummy_magic_24_0.X.n18 two_stage_opamp_dummy_magic_24_0.X.t45 530.201
R21753 two_stage_opamp_dummy_magic_24_0.X.n16 two_stage_opamp_dummy_magic_24_0.X.t40 514.134
R21754 two_stage_opamp_dummy_magic_24_0.X.n15 two_stage_opamp_dummy_magic_24_0.X.t54 514.134
R21755 two_stage_opamp_dummy_magic_24_0.X.n14 two_stage_opamp_dummy_magic_24_0.X.t36 514.134
R21756 two_stage_opamp_dummy_magic_24_0.X.n13 two_stage_opamp_dummy_magic_24_0.X.t49 514.134
R21757 two_stage_opamp_dummy_magic_24_0.X.n12 two_stage_opamp_dummy_magic_24_0.X.t32 514.134
R21758 two_stage_opamp_dummy_magic_24_0.X.n11 two_stage_opamp_dummy_magic_24_0.X.t50 514.134
R21759 two_stage_opamp_dummy_magic_24_0.X.n10 two_stage_opamp_dummy_magic_24_0.X.t33 514.134
R21760 two_stage_opamp_dummy_magic_24_0.X.n9 two_stage_opamp_dummy_magic_24_0.X.t28 514.134
R21761 two_stage_opamp_dummy_magic_24_0.X.n19 two_stage_opamp_dummy_magic_24_0.X.t35 353.467
R21762 two_stage_opamp_dummy_magic_24_0.X.n20 two_stage_opamp_dummy_magic_24_0.X.t53 353.467
R21763 two_stage_opamp_dummy_magic_24_0.X.n21 two_stage_opamp_dummy_magic_24_0.X.t34 353.467
R21764 two_stage_opamp_dummy_magic_24_0.X.n22 two_stage_opamp_dummy_magic_24_0.X.t52 353.467
R21765 two_stage_opamp_dummy_magic_24_0.X.n23 two_stage_opamp_dummy_magic_24_0.X.t39 353.467
R21766 two_stage_opamp_dummy_magic_24_0.X.n24 two_stage_opamp_dummy_magic_24_0.X.t27 353.467
R21767 two_stage_opamp_dummy_magic_24_0.X.n25 two_stage_opamp_dummy_magic_24_0.X.t42 353.467
R21768 two_stage_opamp_dummy_magic_24_0.X.n18 two_stage_opamp_dummy_magic_24_0.X.t30 353.467
R21769 two_stage_opamp_dummy_magic_24_0.X.n42 two_stage_opamp_dummy_magic_24_0.X.n41 176.733
R21770 two_stage_opamp_dummy_magic_24_0.X.n41 two_stage_opamp_dummy_magic_24_0.X.n40 176.733
R21771 two_stage_opamp_dummy_magic_24_0.X.n40 two_stage_opamp_dummy_magic_24_0.X.n39 176.733
R21772 two_stage_opamp_dummy_magic_24_0.X.n44 two_stage_opamp_dummy_magic_24_0.X.n43 176.733
R21773 two_stage_opamp_dummy_magic_24_0.X.n45 two_stage_opamp_dummy_magic_24_0.X.n44 176.733
R21774 two_stage_opamp_dummy_magic_24_0.X.n46 two_stage_opamp_dummy_magic_24_0.X.n45 176.733
R21775 two_stage_opamp_dummy_magic_24_0.X.n20 two_stage_opamp_dummy_magic_24_0.X.n19 176.733
R21776 two_stage_opamp_dummy_magic_24_0.X.n21 two_stage_opamp_dummy_magic_24_0.X.n20 176.733
R21777 two_stage_opamp_dummy_magic_24_0.X.n22 two_stage_opamp_dummy_magic_24_0.X.n21 176.733
R21778 two_stage_opamp_dummy_magic_24_0.X.n23 two_stage_opamp_dummy_magic_24_0.X.n22 176.733
R21779 two_stage_opamp_dummy_magic_24_0.X.n24 two_stage_opamp_dummy_magic_24_0.X.n23 176.733
R21780 two_stage_opamp_dummy_magic_24_0.X.n25 two_stage_opamp_dummy_magic_24_0.X.n24 176.733
R21781 two_stage_opamp_dummy_magic_24_0.X.n11 two_stage_opamp_dummy_magic_24_0.X.n10 176.733
R21782 two_stage_opamp_dummy_magic_24_0.X.n12 two_stage_opamp_dummy_magic_24_0.X.n11 176.733
R21783 two_stage_opamp_dummy_magic_24_0.X.n13 two_stage_opamp_dummy_magic_24_0.X.n12 176.733
R21784 two_stage_opamp_dummy_magic_24_0.X.n14 two_stage_opamp_dummy_magic_24_0.X.n13 176.733
R21785 two_stage_opamp_dummy_magic_24_0.X.n15 two_stage_opamp_dummy_magic_24_0.X.n14 176.733
R21786 two_stage_opamp_dummy_magic_24_0.X.n16 two_stage_opamp_dummy_magic_24_0.X.n15 176.733
R21787 two_stage_opamp_dummy_magic_24_0.X.n27 two_stage_opamp_dummy_magic_24_0.X.n26 165.472
R21788 two_stage_opamp_dummy_magic_24_0.X.n27 two_stage_opamp_dummy_magic_24_0.X.n17 165.472
R21789 two_stage_opamp_dummy_magic_24_0.X.n49 two_stage_opamp_dummy_magic_24_0.X.n48 152
R21790 two_stage_opamp_dummy_magic_24_0.X.n50 two_stage_opamp_dummy_magic_24_0.X.n49 131.571
R21791 two_stage_opamp_dummy_magic_24_0.X.n49 two_stage_opamp_dummy_magic_24_0.X.n47 124.517
R21792 two_stage_opamp_dummy_magic_24_0.X.n78 two_stage_opamp_dummy_magic_24_0.X.n27 74.5362
R21793 two_stage_opamp_dummy_magic_24_0.X.n73 two_stage_opamp_dummy_magic_24_0.X.n72 66.0338
R21794 two_stage_opamp_dummy_magic_24_0.X.n70 two_stage_opamp_dummy_magic_24_0.X.n69 66.0338
R21795 two_stage_opamp_dummy_magic_24_0.X.n67 two_stage_opamp_dummy_magic_24_0.X.n66 66.0338
R21796 two_stage_opamp_dummy_magic_24_0.X.n63 two_stage_opamp_dummy_magic_24_0.X.n62 66.0338
R21797 two_stage_opamp_dummy_magic_24_0.X.n60 two_stage_opamp_dummy_magic_24_0.X.n59 66.0338
R21798 two_stage_opamp_dummy_magic_24_0.X.n57 two_stage_opamp_dummy_magic_24_0.X.n56 66.0338
R21799 two_stage_opamp_dummy_magic_24_0.X.n92 two_stage_opamp_dummy_magic_24_0.X.n90 54.7984
R21800 two_stage_opamp_dummy_magic_24_0.X.n100 two_stage_opamp_dummy_magic_24_0.X.n99 54.4547
R21801 two_stage_opamp_dummy_magic_24_0.X.n98 two_stage_opamp_dummy_magic_24_0.X.n97 54.4547
R21802 two_stage_opamp_dummy_magic_24_0.X.n96 two_stage_opamp_dummy_magic_24_0.X.n95 54.4547
R21803 two_stage_opamp_dummy_magic_24_0.X.n94 two_stage_opamp_dummy_magic_24_0.X.n93 54.4547
R21804 two_stage_opamp_dummy_magic_24_0.X.n92 two_stage_opamp_dummy_magic_24_0.X.n91 54.4547
R21805 two_stage_opamp_dummy_magic_24_0.X.n33 two_stage_opamp_dummy_magic_24_0.X.t19 41.0384
R21806 two_stage_opamp_dummy_magic_24_0.X.n47 two_stage_opamp_dummy_magic_24_0.X.n42 40.1672
R21807 two_stage_opamp_dummy_magic_24_0.X.n47 two_stage_opamp_dummy_magic_24_0.X.n46 40.1672
R21808 two_stage_opamp_dummy_magic_24_0.X.n26 two_stage_opamp_dummy_magic_24_0.X.n18 40.1672
R21809 two_stage_opamp_dummy_magic_24_0.X.n26 two_stage_opamp_dummy_magic_24_0.X.n25 40.1672
R21810 two_stage_opamp_dummy_magic_24_0.X.n17 two_stage_opamp_dummy_magic_24_0.X.n9 40.1672
R21811 two_stage_opamp_dummy_magic_24_0.X.n17 two_stage_opamp_dummy_magic_24_0.X.n16 40.1672
R21812 two_stage_opamp_dummy_magic_24_0.X.n51 two_stage_opamp_dummy_magic_24_0.X.n50 16.3217
R21813 two_stage_opamp_dummy_magic_24_0.X.n99 two_stage_opamp_dummy_magic_24_0.X.t18 16.0005
R21814 two_stage_opamp_dummy_magic_24_0.X.n99 two_stage_opamp_dummy_magic_24_0.X.t2 16.0005
R21815 two_stage_opamp_dummy_magic_24_0.X.n97 two_stage_opamp_dummy_magic_24_0.X.t1 16.0005
R21816 two_stage_opamp_dummy_magic_24_0.X.n97 two_stage_opamp_dummy_magic_24_0.X.t20 16.0005
R21817 two_stage_opamp_dummy_magic_24_0.X.n95 two_stage_opamp_dummy_magic_24_0.X.t15 16.0005
R21818 two_stage_opamp_dummy_magic_24_0.X.n95 two_stage_opamp_dummy_magic_24_0.X.t0 16.0005
R21819 two_stage_opamp_dummy_magic_24_0.X.n93 two_stage_opamp_dummy_magic_24_0.X.t4 16.0005
R21820 two_stage_opamp_dummy_magic_24_0.X.n93 two_stage_opamp_dummy_magic_24_0.X.t17 16.0005
R21821 two_stage_opamp_dummy_magic_24_0.X.n91 two_stage_opamp_dummy_magic_24_0.X.t16 16.0005
R21822 two_stage_opamp_dummy_magic_24_0.X.n91 two_stage_opamp_dummy_magic_24_0.X.t24 16.0005
R21823 two_stage_opamp_dummy_magic_24_0.X.n90 two_stage_opamp_dummy_magic_24_0.X.t3 16.0005
R21824 two_stage_opamp_dummy_magic_24_0.X.n90 two_stage_opamp_dummy_magic_24_0.X.t23 16.0005
R21825 two_stage_opamp_dummy_magic_24_0.X.n48 two_stage_opamp_dummy_magic_24_0.X.n38 12.8005
R21826 two_stage_opamp_dummy_magic_24_0.X.n72 two_stage_opamp_dummy_magic_24_0.X.t22 11.2576
R21827 two_stage_opamp_dummy_magic_24_0.X.n72 two_stage_opamp_dummy_magic_24_0.X.t11 11.2576
R21828 two_stage_opamp_dummy_magic_24_0.X.n69 two_stage_opamp_dummy_magic_24_0.X.t14 11.2576
R21829 two_stage_opamp_dummy_magic_24_0.X.n69 two_stage_opamp_dummy_magic_24_0.X.t12 11.2576
R21830 two_stage_opamp_dummy_magic_24_0.X.n66 two_stage_opamp_dummy_magic_24_0.X.t5 11.2576
R21831 two_stage_opamp_dummy_magic_24_0.X.n66 two_stage_opamp_dummy_magic_24_0.X.t6 11.2576
R21832 two_stage_opamp_dummy_magic_24_0.X.n62 two_stage_opamp_dummy_magic_24_0.X.t7 11.2576
R21833 two_stage_opamp_dummy_magic_24_0.X.n62 two_stage_opamp_dummy_magic_24_0.X.t9 11.2576
R21834 two_stage_opamp_dummy_magic_24_0.X.n59 two_stage_opamp_dummy_magic_24_0.X.t8 11.2576
R21835 two_stage_opamp_dummy_magic_24_0.X.n59 two_stage_opamp_dummy_magic_24_0.X.t10 11.2576
R21836 two_stage_opamp_dummy_magic_24_0.X.n56 two_stage_opamp_dummy_magic_24_0.X.t13 11.2576
R21837 two_stage_opamp_dummy_magic_24_0.X.n56 two_stage_opamp_dummy_magic_24_0.X.t21 11.2576
R21838 two_stage_opamp_dummy_magic_24_0.X.n101 two_stage_opamp_dummy_magic_24_0.X.n100 10.9224
R21839 two_stage_opamp_dummy_magic_24_0.X.n48 two_stage_opamp_dummy_magic_24_0.X.n36 9.36264
R21840 two_stage_opamp_dummy_magic_24_0.X.n38 two_stage_opamp_dummy_magic_24_0.X.n37 9.3005
R21841 two_stage_opamp_dummy_magic_24_0.X.n85 two_stage_opamp_dummy_magic_24_0.X.n3 5.96925
R21842 two_stage_opamp_dummy_magic_24_0.X.n58 two_stage_opamp_dummy_magic_24_0.X.n57 5.91717
R21843 two_stage_opamp_dummy_magic_24_0.X.n73 two_stage_opamp_dummy_magic_24_0.X.n71 5.91717
R21844 two_stage_opamp_dummy_magic_24_0.X.n102 two_stage_opamp_dummy_magic_24_0.X.n101 5.68397
R21845 two_stage_opamp_dummy_magic_24_0.X.n61 two_stage_opamp_dummy_magic_24_0.X.n57 5.66717
R21846 two_stage_opamp_dummy_magic_24_0.X.n85 two_stage_opamp_dummy_magic_24_0.X.n84 5.6255
R21847 two_stage_opamp_dummy_magic_24_0.X.n86 two_stage_opamp_dummy_magic_24_0.X.n2 5.6255
R21848 two_stage_opamp_dummy_magic_24_0.X.n105 two_stage_opamp_dummy_magic_24_0.X.n87 5.6255
R21849 two_stage_opamp_dummy_magic_24_0.X.n89 two_stage_opamp_dummy_magic_24_0.X.n88 5.6255
R21850 two_stage_opamp_dummy_magic_24_0.X.n50 two_stage_opamp_dummy_magic_24_0.X.n38 5.33141
R21851 two_stage_opamp_dummy_magic_24_0.X.n70 two_stage_opamp_dummy_magic_24_0.X.n54 5.29217
R21852 two_stage_opamp_dummy_magic_24_0.X.n71 two_stage_opamp_dummy_magic_24_0.X.n70 5.29217
R21853 two_stage_opamp_dummy_magic_24_0.X.n67 two_stage_opamp_dummy_magic_24_0.X.n65 5.29217
R21854 two_stage_opamp_dummy_magic_24_0.X.n68 two_stage_opamp_dummy_magic_24_0.X.n67 5.29217
R21855 two_stage_opamp_dummy_magic_24_0.X.n64 two_stage_opamp_dummy_magic_24_0.X.n63 5.29217
R21856 two_stage_opamp_dummy_magic_24_0.X.n63 two_stage_opamp_dummy_magic_24_0.X.n55 5.29217
R21857 two_stage_opamp_dummy_magic_24_0.X.n61 two_stage_opamp_dummy_magic_24_0.X.n60 5.29217
R21858 two_stage_opamp_dummy_magic_24_0.X.n60 two_stage_opamp_dummy_magic_24_0.X.n58 5.29217
R21859 two_stage_opamp_dummy_magic_24_0.X.n74 two_stage_opamp_dummy_magic_24_0.X.n73 5.29217
R21860 two_stage_opamp_dummy_magic_24_0.X.n77 two_stage_opamp_dummy_magic_24_0.X.n53 4.5005
R21861 two_stage_opamp_dummy_magic_24_0.X.n79 two_stage_opamp_dummy_magic_24_0.X.n78 4.5005
R21862 two_stage_opamp_dummy_magic_24_0.X.n78 two_stage_opamp_dummy_magic_24_0.X.n77 4.5005
R21863 two_stage_opamp_dummy_magic_24_0.X.n52 two_stage_opamp_dummy_magic_24_0.X.n51 4.5005
R21864 two_stage_opamp_dummy_magic_24_0.X.n30 two_stage_opamp_dummy_magic_24_0.X.n29 4.5005
R21865 two_stage_opamp_dummy_magic_24_0.X.n75 two_stage_opamp_dummy_magic_24_0.X.n74 4.49606
R21866 two_stage_opamp_dummy_magic_24_0.X.n32 two_stage_opamp_dummy_magic_24_0.X.n31 2.26187
R21867 two_stage_opamp_dummy_magic_24_0.X.n31 two_stage_opamp_dummy_magic_24_0.X.n28 2.26187
R21868 two_stage_opamp_dummy_magic_24_0.X.n79 two_stage_opamp_dummy_magic_24_0.X.n7 2.24063
R21869 two_stage_opamp_dummy_magic_24_0.X.n8 two_stage_opamp_dummy_magic_24_0.X.n6 2.24063
R21870 two_stage_opamp_dummy_magic_24_0.X.n76 two_stage_opamp_dummy_magic_24_0.X.n75 2.24063
R21871 two_stage_opamp_dummy_magic_24_0.X.n33 two_stage_opamp_dummy_magic_24_0.X.n32 2.24063
R21872 two_stage_opamp_dummy_magic_24_0.X.n35 two_stage_opamp_dummy_magic_24_0.X.n34 2.24063
R21873 two_stage_opamp_dummy_magic_24_0.X.n52 two_stage_opamp_dummy_magic_24_0.X.n36 2.22018
R21874 two_stage_opamp_dummy_magic_24_0.X.n104 two_stage_opamp_dummy_magic_24_0.X.n103 1.5005
R21875 two_stage_opamp_dummy_magic_24_0.X.n105 two_stage_opamp_dummy_magic_24_0.X.n1 1.5005
R21876 two_stage_opamp_dummy_magic_24_0.X.n107 two_stage_opamp_dummy_magic_24_0.X.n106 1.5005
R21877 two_stage_opamp_dummy_magic_24_0.X.n2 two_stage_opamp_dummy_magic_24_0.X.n0 1.5005
R21878 two_stage_opamp_dummy_magic_24_0.X.n82 two_stage_opamp_dummy_magic_24_0.X.n5 1.5005
R21879 two_stage_opamp_dummy_magic_24_0.X.n84 two_stage_opamp_dummy_magic_24_0.X.n83 1.5005
R21880 two_stage_opamp_dummy_magic_24_0.X.n81 two_stage_opamp_dummy_magic_24_0.X.n4 1.5005
R21881 two_stage_opamp_dummy_magic_24_0.X.n80 two_stage_opamp_dummy_magic_24_0.X.n3 1.5005
R21882 two_stage_opamp_dummy_magic_24_0.X.n52 two_stage_opamp_dummy_magic_24_0.X.n35 0.682792
R21883 two_stage_opamp_dummy_magic_24_0.X.n80 two_stage_opamp_dummy_magic_24_0.X.n79 0.630708
R21884 two_stage_opamp_dummy_magic_24_0.X.n58 two_stage_opamp_dummy_magic_24_0.X.n55 0.6255
R21885 two_stage_opamp_dummy_magic_24_0.X.n68 two_stage_opamp_dummy_magic_24_0.X.n55 0.6255
R21886 two_stage_opamp_dummy_magic_24_0.X.n71 two_stage_opamp_dummy_magic_24_0.X.n68 0.6255
R21887 two_stage_opamp_dummy_magic_24_0.X.n103 two_stage_opamp_dummy_magic_24_0.X.n102 0.564601
R21888 two_stage_opamp_dummy_magic_24_0.X.n77 two_stage_opamp_dummy_magic_24_0.X.n52 0.46925
R21889 two_stage_opamp_dummy_magic_24_0.X.n74 two_stage_opamp_dummy_magic_24_0.X.n54 0.3755
R21890 two_stage_opamp_dummy_magic_24_0.X.n65 two_stage_opamp_dummy_magic_24_0.X.n54 0.3755
R21891 two_stage_opamp_dummy_magic_24_0.X.n65 two_stage_opamp_dummy_magic_24_0.X.n64 0.3755
R21892 two_stage_opamp_dummy_magic_24_0.X.n64 two_stage_opamp_dummy_magic_24_0.X.n61 0.3755
R21893 two_stage_opamp_dummy_magic_24_0.X.n94 two_stage_opamp_dummy_magic_24_0.X.n92 0.34425
R21894 two_stage_opamp_dummy_magic_24_0.X.n96 two_stage_opamp_dummy_magic_24_0.X.n94 0.34425
R21895 two_stage_opamp_dummy_magic_24_0.X.n98 two_stage_opamp_dummy_magic_24_0.X.n96 0.34425
R21896 two_stage_opamp_dummy_magic_24_0.X.n100 two_stage_opamp_dummy_magic_24_0.X.n98 0.34425
R21897 two_stage_opamp_dummy_magic_24_0.X.n86 two_stage_opamp_dummy_magic_24_0.X.n85 0.34425
R21898 two_stage_opamp_dummy_magic_24_0.X.n87 two_stage_opamp_dummy_magic_24_0.X.n86 0.34425
R21899 two_stage_opamp_dummy_magic_24_0.X.n89 two_stage_opamp_dummy_magic_24_0.X.n87 0.34425
R21900 two_stage_opamp_dummy_magic_24_0.X.n101 two_stage_opamp_dummy_magic_24_0.X.n89 0.34425
R21901 two_stage_opamp_dummy_magic_24_0.X.n51 two_stage_opamp_dummy_magic_24_0.X.n37 0.1255
R21902 two_stage_opamp_dummy_magic_24_0.X.n37 two_stage_opamp_dummy_magic_24_0.X.n36 0.0626438
R21903 two_stage_opamp_dummy_magic_24_0.X.n4 two_stage_opamp_dummy_magic_24_0.X.n3 0.0577917
R21904 two_stage_opamp_dummy_magic_24_0.X.n84 two_stage_opamp_dummy_magic_24_0.X.n4 0.0577917
R21905 two_stage_opamp_dummy_magic_24_0.X.n84 two_stage_opamp_dummy_magic_24_0.X.n5 0.0577917
R21906 two_stage_opamp_dummy_magic_24_0.X.n5 two_stage_opamp_dummy_magic_24_0.X.n2 0.0577917
R21907 two_stage_opamp_dummy_magic_24_0.X.n106 two_stage_opamp_dummy_magic_24_0.X.n2 0.0577917
R21908 two_stage_opamp_dummy_magic_24_0.X.n106 two_stage_opamp_dummy_magic_24_0.X.n105 0.0577917
R21909 two_stage_opamp_dummy_magic_24_0.X.n105 two_stage_opamp_dummy_magic_24_0.X.n104 0.0577917
R21910 two_stage_opamp_dummy_magic_24_0.X.n104 two_stage_opamp_dummy_magic_24_0.X.n88 0.0577917
R21911 two_stage_opamp_dummy_magic_24_0.X.n81 two_stage_opamp_dummy_magic_24_0.X.n80 0.0577917
R21912 two_stage_opamp_dummy_magic_24_0.X.n83 two_stage_opamp_dummy_magic_24_0.X.n81 0.0577917
R21913 two_stage_opamp_dummy_magic_24_0.X.n83 two_stage_opamp_dummy_magic_24_0.X.n82 0.0577917
R21914 two_stage_opamp_dummy_magic_24_0.X.n82 two_stage_opamp_dummy_magic_24_0.X.n0 0.0577917
R21915 two_stage_opamp_dummy_magic_24_0.X.n107 two_stage_opamp_dummy_magic_24_0.X.n1 0.0577917
R21916 two_stage_opamp_dummy_magic_24_0.X.n103 two_stage_opamp_dummy_magic_24_0.X.n1 0.0577917
R21917 two_stage_opamp_dummy_magic_24_0.X.n102 two_stage_opamp_dummy_magic_24_0.X.n88 0.054517
R21918 two_stage_opamp_dummy_magic_24_0.X.n79 two_stage_opamp_dummy_magic_24_0.X.n6 0.0421667
R21919 two_stage_opamp_dummy_magic_24_0.X two_stage_opamp_dummy_magic_24_0.X.n107 0.0369583
R21920 two_stage_opamp_dummy_magic_24_0.X.n75 two_stage_opamp_dummy_magic_24_0.X.n7 0.0217373
R21921 two_stage_opamp_dummy_magic_24_0.X.n78 two_stage_opamp_dummy_magic_24_0.X.n8 0.0217373
R21922 two_stage_opamp_dummy_magic_24_0.X.n35 two_stage_opamp_dummy_magic_24_0.X.n28 0.0217373
R21923 two_stage_opamp_dummy_magic_24_0.X.n53 two_stage_opamp_dummy_magic_24_0.X.n7 0.0217373
R21924 two_stage_opamp_dummy_magic_24_0.X.n53 two_stage_opamp_dummy_magic_24_0.X.n8 0.0217373
R21925 two_stage_opamp_dummy_magic_24_0.X.n31 two_stage_opamp_dummy_magic_24_0.X.n29 0.0217373
R21926 two_stage_opamp_dummy_magic_24_0.X.n30 two_stage_opamp_dummy_magic_24_0.X.n28 0.0217373
R21927 two_stage_opamp_dummy_magic_24_0.X.n32 two_stage_opamp_dummy_magic_24_0.X.n30 0.0217373
R21928 two_stage_opamp_dummy_magic_24_0.X.n77 two_stage_opamp_dummy_magic_24_0.X.n76 0.0217373
R21929 two_stage_opamp_dummy_magic_24_0.X.n76 two_stage_opamp_dummy_magic_24_0.X.n6 0.0217373
R21930 two_stage_opamp_dummy_magic_24_0.X.n34 two_stage_opamp_dummy_magic_24_0.X.n29 0.0217373
R21931 two_stage_opamp_dummy_magic_24_0.X.n34 two_stage_opamp_dummy_magic_24_0.X.n33 0.0217373
R21932 two_stage_opamp_dummy_magic_24_0.X two_stage_opamp_dummy_magic_24_0.X.n0 0.0213333
R21933 two_stage_opamp_dummy_magic_24_0.Vb1.n9 two_stage_opamp_dummy_magic_24_0.Vb1.t22 484.385
R21934 two_stage_opamp_dummy_magic_24_0.Vb1.n7 two_stage_opamp_dummy_magic_24_0.Vb1.t16 484.212
R21935 two_stage_opamp_dummy_magic_24_0.Vb1.n7 two_stage_opamp_dummy_magic_24_0.Vb1.t27 484.212
R21936 two_stage_opamp_dummy_magic_24_0.Vb1.n7 two_stage_opamp_dummy_magic_24_0.Vb1.t14 484.212
R21937 two_stage_opamp_dummy_magic_24_0.Vb1.n7 two_stage_opamp_dummy_magic_24_0.Vb1.t26 484.212
R21938 two_stage_opamp_dummy_magic_24_0.Vb1.n6 two_stage_opamp_dummy_magic_24_0.Vb1.t13 484.212
R21939 two_stage_opamp_dummy_magic_24_0.Vb1.n6 two_stage_opamp_dummy_magic_24_0.Vb1.t24 484.212
R21940 two_stage_opamp_dummy_magic_24_0.Vb1.n6 two_stage_opamp_dummy_magic_24_0.Vb1.t19 484.212
R21941 two_stage_opamp_dummy_magic_24_0.Vb1.n6 two_stage_opamp_dummy_magic_24_0.Vb1.t25 484.212
R21942 two_stage_opamp_dummy_magic_24_0.Vb1.n8 two_stage_opamp_dummy_magic_24_0.Vb1.t32 484.212
R21943 two_stage_opamp_dummy_magic_24_0.Vb1.n8 two_stage_opamp_dummy_magic_24_0.Vb1.t23 484.212
R21944 two_stage_opamp_dummy_magic_24_0.Vb1.n11 two_stage_opamp_dummy_magic_24_0.Vb1.t21 484.212
R21945 two_stage_opamp_dummy_magic_24_0.Vb1.n11 two_stage_opamp_dummy_magic_24_0.Vb1.t31 484.212
R21946 two_stage_opamp_dummy_magic_24_0.Vb1.n10 two_stage_opamp_dummy_magic_24_0.Vb1.t20 484.212
R21947 two_stage_opamp_dummy_magic_24_0.Vb1.n10 two_stage_opamp_dummy_magic_24_0.Vb1.t29 484.212
R21948 two_stage_opamp_dummy_magic_24_0.Vb1.n10 two_stage_opamp_dummy_magic_24_0.Vb1.t17 484.212
R21949 two_stage_opamp_dummy_magic_24_0.Vb1.n10 two_stage_opamp_dummy_magic_24_0.Vb1.t30 484.212
R21950 two_stage_opamp_dummy_magic_24_0.Vb1.n9 two_stage_opamp_dummy_magic_24_0.Vb1.t18 484.212
R21951 two_stage_opamp_dummy_magic_24_0.Vb1.n9 two_stage_opamp_dummy_magic_24_0.Vb1.t28 484.212
R21952 two_stage_opamp_dummy_magic_24_0.Vb1.n9 two_stage_opamp_dummy_magic_24_0.Vb1.t15 484.212
R21953 two_stage_opamp_dummy_magic_24_0.Vb1.n14 two_stage_opamp_dummy_magic_24_0.Vb1.t8 449.868
R21954 two_stage_opamp_dummy_magic_24_0.Vb1.n13 two_stage_opamp_dummy_magic_24_0.Vb1.t4 449.868
R21955 two_stage_opamp_dummy_magic_24_0.Vb1.n14 two_stage_opamp_dummy_magic_24_0.Vb1.t6 273.134
R21956 two_stage_opamp_dummy_magic_24_0.Vb1.n13 two_stage_opamp_dummy_magic_24_0.Vb1.t2 273.134
R21957 two_stage_opamp_dummy_magic_24_0.Vb1.n3 two_stage_opamp_dummy_magic_24_0.Vb1.t12 166.847
R21958 two_stage_opamp_dummy_magic_24_0.Vb1.t12 two_stage_opamp_dummy_magic_24_0.Vb1.n5 166.847
R21959 two_stage_opamp_dummy_magic_24_0.Vb1.n0 two_stage_opamp_dummy_magic_24_0.Vb1.n15 161.3
R21960 two_stage_opamp_dummy_magic_24_0.Vb1 two_stage_opamp_dummy_magic_24_0.Vb1.n12 151.863
R21961 two_stage_opamp_dummy_magic_24_0.Vb1.n0 two_stage_opamp_dummy_magic_24_0.Vb1.n18 49.3505
R21962 two_stage_opamp_dummy_magic_24_0.Vb1.n17 two_stage_opamp_dummy_magic_24_0.Vb1.n16 49.3505
R21963 two_stage_opamp_dummy_magic_24_0.Vb1.n15 two_stage_opamp_dummy_magic_24_0.Vb1.n14 45.5227
R21964 two_stage_opamp_dummy_magic_24_0.Vb1.n15 two_stage_opamp_dummy_magic_24_0.Vb1.n13 45.5227
R21965 two_stage_opamp_dummy_magic_24_0.Vb1 two_stage_opamp_dummy_magic_24_0.Vb1.n20 37.089
R21966 two_stage_opamp_dummy_magic_24_0.Vb1.n12 two_stage_opamp_dummy_magic_24_0.Vb1.t11 19.7005
R21967 two_stage_opamp_dummy_magic_24_0.Vb1.n12 two_stage_opamp_dummy_magic_24_0.Vb1.t10 19.7005
R21968 two_stage_opamp_dummy_magic_24_0.Vb1.n18 two_stage_opamp_dummy_magic_24_0.Vb1.t3 16.0005
R21969 two_stage_opamp_dummy_magic_24_0.Vb1.n18 two_stage_opamp_dummy_magic_24_0.Vb1.t7 16.0005
R21970 two_stage_opamp_dummy_magic_24_0.Vb1.n16 two_stage_opamp_dummy_magic_24_0.Vb1.t0 16.0005
R21971 two_stage_opamp_dummy_magic_24_0.Vb1.n16 two_stage_opamp_dummy_magic_24_0.Vb1.t5 16.0005
R21972 two_stage_opamp_dummy_magic_24_0.Vb1.n19 two_stage_opamp_dummy_magic_24_0.Vb1.t9 16.0005
R21973 two_stage_opamp_dummy_magic_24_0.Vb1.n19 two_stage_opamp_dummy_magic_24_0.Vb1.t1 16.0005
R21974 two_stage_opamp_dummy_magic_24_0.Vb1.n1 two_stage_opamp_dummy_magic_24_0.Vb1.n0 4.938
R21975 two_stage_opamp_dummy_magic_24_0.Vb1.n19 two_stage_opamp_dummy_magic_24_0.Vb1.n2 51.6321
R21976 two_stage_opamp_dummy_magic_24_0.Vb1.n17 two_stage_opamp_dummy_magic_24_0.Vb1.n5 4.938
R21977 two_stage_opamp_dummy_magic_24_0.Vb1.n3 two_stage_opamp_dummy_magic_24_0.Vb1.n17 4.938
R21978 two_stage_opamp_dummy_magic_24_0.Vb1.n0 two_stage_opamp_dummy_magic_24_0.Vb1.n4 4.938
R21979 two_stage_opamp_dummy_magic_24_0.Vb1.n1 two_stage_opamp_dummy_magic_24_0.Vb1.n2 0.376365
R21980 two_stage_opamp_dummy_magic_24_0.Vb1.n20 two_stage_opamp_dummy_magic_24_0.Vb1.n1 4.88363
R21981 two_stage_opamp_dummy_magic_24_0.Vb1.n20 two_stage_opamp_dummy_magic_24_0.Vb1.n7 2.99226
R21982 two_stage_opamp_dummy_magic_24_0.Vb1.n7 two_stage_opamp_dummy_magic_24_0.Vb1.n6 1.03175
R21983 two_stage_opamp_dummy_magic_24_0.Vb1 two_stage_opamp_dummy_magic_24_0.Vb1.n11 0.852062
R21984 two_stage_opamp_dummy_magic_24_0.Vb1.n8 two_stage_opamp_dummy_magic_24_0.Vb1 0.852062
R21985 two_stage_opamp_dummy_magic_24_0.Vb1.n2 two_stage_opamp_dummy_magic_24_0.Vb1.n4 0.376365
R21986 two_stage_opamp_dummy_magic_24_0.Vb1.n10 two_stage_opamp_dummy_magic_24_0.Vb1.n9 0.688
R21987 two_stage_opamp_dummy_magic_24_0.Vb1.n11 two_stage_opamp_dummy_magic_24_0.Vb1.n10 0.688
R21988 two_stage_opamp_dummy_magic_24_0.Vb1.n1 two_stage_opamp_dummy_magic_24_0.Vb1.n5 0.688
R21989 two_stage_opamp_dummy_magic_24_0.Vb1.n4 two_stage_opamp_dummy_magic_24_0.Vb1.n3 0.688
R21990 two_stage_opamp_dummy_magic_24_0.Vb1.n6 two_stage_opamp_dummy_magic_24_0.Vb1.n8 0.516125
R21991 two_stage_opamp_dummy_magic_24_0.Vb1_2.n1 two_stage_opamp_dummy_magic_24_0.Vb1_2.t4 65.3505
R21992 two_stage_opamp_dummy_magic_24_0.Vb1_2.n3 two_stage_opamp_dummy_magic_24_0.Vb1_2.n2 49.3505
R21993 two_stage_opamp_dummy_magic_24_0.Vb1_2.n6 two_stage_opamp_dummy_magic_24_0.Vb1_2.n5 49.3505
R21994 two_stage_opamp_dummy_magic_24_0.Vb1_2.n2 two_stage_opamp_dummy_magic_24_0.Vb1_2.t2 16.0005
R21995 two_stage_opamp_dummy_magic_24_0.Vb1_2.n2 two_stage_opamp_dummy_magic_24_0.Vb1_2.t0 16.0005
R21996 two_stage_opamp_dummy_magic_24_0.Vb1_2.t3 two_stage_opamp_dummy_magic_24_0.Vb1_2.n6 16.0005
R21997 two_stage_opamp_dummy_magic_24_0.Vb1_2.n6 two_stage_opamp_dummy_magic_24_0.Vb1_2.t1 16.0005
R21998 two_stage_opamp_dummy_magic_24_0.Vb1_2.n1 two_stage_opamp_dummy_magic_24_0.Vb1_2.n0 6.41717
R21999 two_stage_opamp_dummy_magic_24_0.Vb1_2.n4 two_stage_opamp_dummy_magic_24_0.Vb1_2.n1 5.85467
R22000 two_stage_opamp_dummy_magic_24_0.Vb1_2.n3 two_stage_opamp_dummy_magic_24_0.Vb1_2.n0 5.72967
R22001 two_stage_opamp_dummy_magic_24_0.Vb1_2.n4 two_stage_opamp_dummy_magic_24_0.Vb1_2.n3 5.51092
R22002 two_stage_opamp_dummy_magic_24_0.Vb1_2.n5 two_stage_opamp_dummy_magic_24_0.Vb1_2.n0 5.16717
R22003 two_stage_opamp_dummy_magic_24_0.Vb1_2.n5 two_stage_opamp_dummy_magic_24_0.Vb1_2.n4 5.16717
R22004 two_stage_opamp_dummy_magic_24_0.Y.n64 two_stage_opamp_dummy_magic_24_0.Y.t48 1172.87
R22005 two_stage_opamp_dummy_magic_24_0.Y.n60 two_stage_opamp_dummy_magic_24_0.Y.t39 1172.87
R22006 two_stage_opamp_dummy_magic_24_0.Y.n64 two_stage_opamp_dummy_magic_24_0.Y.t40 996.134
R22007 two_stage_opamp_dummy_magic_24_0.Y.n65 two_stage_opamp_dummy_magic_24_0.Y.t28 996.134
R22008 two_stage_opamp_dummy_magic_24_0.Y.n66 two_stage_opamp_dummy_magic_24_0.Y.t44 996.134
R22009 two_stage_opamp_dummy_magic_24_0.Y.n67 two_stage_opamp_dummy_magic_24_0.Y.t30 996.134
R22010 two_stage_opamp_dummy_magic_24_0.Y.n63 two_stage_opamp_dummy_magic_24_0.Y.t47 996.134
R22011 two_stage_opamp_dummy_magic_24_0.Y.n62 two_stage_opamp_dummy_magic_24_0.Y.t52 996.134
R22012 two_stage_opamp_dummy_magic_24_0.Y.n61 two_stage_opamp_dummy_magic_24_0.Y.t35 996.134
R22013 two_stage_opamp_dummy_magic_24_0.Y.n60 two_stage_opamp_dummy_magic_24_0.Y.t25 996.134
R22014 two_stage_opamp_dummy_magic_24_0.Y.n36 two_stage_opamp_dummy_magic_24_0.Y.t43 690.867
R22015 two_stage_opamp_dummy_magic_24_0.Y.n29 two_stage_opamp_dummy_magic_24_0.Y.t33 690.867
R22016 two_stage_opamp_dummy_magic_24_0.Y.n45 two_stage_opamp_dummy_magic_24_0.Y.t46 530.201
R22017 two_stage_opamp_dummy_magic_24_0.Y.n38 two_stage_opamp_dummy_magic_24_0.Y.t36 530.201
R22018 two_stage_opamp_dummy_magic_24_0.Y.n36 two_stage_opamp_dummy_magic_24_0.Y.t34 514.134
R22019 two_stage_opamp_dummy_magic_24_0.Y.n29 two_stage_opamp_dummy_magic_24_0.Y.t51 514.134
R22020 two_stage_opamp_dummy_magic_24_0.Y.n30 two_stage_opamp_dummy_magic_24_0.Y.t31 514.134
R22021 two_stage_opamp_dummy_magic_24_0.Y.n31 two_stage_opamp_dummy_magic_24_0.Y.t49 514.134
R22022 two_stage_opamp_dummy_magic_24_0.Y.n32 two_stage_opamp_dummy_magic_24_0.Y.t42 514.134
R22023 two_stage_opamp_dummy_magic_24_0.Y.n33 two_stage_opamp_dummy_magic_24_0.Y.t27 514.134
R22024 two_stage_opamp_dummy_magic_24_0.Y.n34 two_stage_opamp_dummy_magic_24_0.Y.t38 514.134
R22025 two_stage_opamp_dummy_magic_24_0.Y.n35 two_stage_opamp_dummy_magic_24_0.Y.t54 514.134
R22026 two_stage_opamp_dummy_magic_24_0.Y.n45 two_stage_opamp_dummy_magic_24_0.Y.t37 353.467
R22027 two_stage_opamp_dummy_magic_24_0.Y.n44 two_stage_opamp_dummy_magic_24_0.Y.t26 353.467
R22028 two_stage_opamp_dummy_magic_24_0.Y.n43 two_stage_opamp_dummy_magic_24_0.Y.t41 353.467
R22029 two_stage_opamp_dummy_magic_24_0.Y.n42 two_stage_opamp_dummy_magic_24_0.Y.t29 353.467
R22030 two_stage_opamp_dummy_magic_24_0.Y.n41 two_stage_opamp_dummy_magic_24_0.Y.t45 353.467
R22031 two_stage_opamp_dummy_magic_24_0.Y.n40 two_stage_opamp_dummy_magic_24_0.Y.t50 353.467
R22032 two_stage_opamp_dummy_magic_24_0.Y.n39 two_stage_opamp_dummy_magic_24_0.Y.t32 353.467
R22033 two_stage_opamp_dummy_magic_24_0.Y.n38 two_stage_opamp_dummy_magic_24_0.Y.t53 353.467
R22034 two_stage_opamp_dummy_magic_24_0.Y.n63 two_stage_opamp_dummy_magic_24_0.Y.n62 176.733
R22035 two_stage_opamp_dummy_magic_24_0.Y.n62 two_stage_opamp_dummy_magic_24_0.Y.n61 176.733
R22036 two_stage_opamp_dummy_magic_24_0.Y.n61 two_stage_opamp_dummy_magic_24_0.Y.n60 176.733
R22037 two_stage_opamp_dummy_magic_24_0.Y.n65 two_stage_opamp_dummy_magic_24_0.Y.n64 176.733
R22038 two_stage_opamp_dummy_magic_24_0.Y.n66 two_stage_opamp_dummy_magic_24_0.Y.n65 176.733
R22039 two_stage_opamp_dummy_magic_24_0.Y.n67 two_stage_opamp_dummy_magic_24_0.Y.n66 176.733
R22040 two_stage_opamp_dummy_magic_24_0.Y.n44 two_stage_opamp_dummy_magic_24_0.Y.n43 176.733
R22041 two_stage_opamp_dummy_magic_24_0.Y.n43 two_stage_opamp_dummy_magic_24_0.Y.n42 176.733
R22042 two_stage_opamp_dummy_magic_24_0.Y.n42 two_stage_opamp_dummy_magic_24_0.Y.n41 176.733
R22043 two_stage_opamp_dummy_magic_24_0.Y.n41 two_stage_opamp_dummy_magic_24_0.Y.n40 176.733
R22044 two_stage_opamp_dummy_magic_24_0.Y.n40 two_stage_opamp_dummy_magic_24_0.Y.n39 176.733
R22045 two_stage_opamp_dummy_magic_24_0.Y.n39 two_stage_opamp_dummy_magic_24_0.Y.n38 176.733
R22046 two_stage_opamp_dummy_magic_24_0.Y.n35 two_stage_opamp_dummy_magic_24_0.Y.n34 176.733
R22047 two_stage_opamp_dummy_magic_24_0.Y.n34 two_stage_opamp_dummy_magic_24_0.Y.n33 176.733
R22048 two_stage_opamp_dummy_magic_24_0.Y.n33 two_stage_opamp_dummy_magic_24_0.Y.n32 176.733
R22049 two_stage_opamp_dummy_magic_24_0.Y.n32 two_stage_opamp_dummy_magic_24_0.Y.n31 176.733
R22050 two_stage_opamp_dummy_magic_24_0.Y.n31 two_stage_opamp_dummy_magic_24_0.Y.n30 176.733
R22051 two_stage_opamp_dummy_magic_24_0.Y.n30 two_stage_opamp_dummy_magic_24_0.Y.n29 176.733
R22052 two_stage_opamp_dummy_magic_24_0.Y.n47 two_stage_opamp_dummy_magic_24_0.Y.n46 165.472
R22053 two_stage_opamp_dummy_magic_24_0.Y.n47 two_stage_opamp_dummy_magic_24_0.Y.n37 165.472
R22054 two_stage_opamp_dummy_magic_24_0.Y.n70 two_stage_opamp_dummy_magic_24_0.Y.n69 152
R22055 two_stage_opamp_dummy_magic_24_0.Y.n71 two_stage_opamp_dummy_magic_24_0.Y.n70 131.571
R22056 two_stage_opamp_dummy_magic_24_0.Y.n70 two_stage_opamp_dummy_magic_24_0.Y.n68 124.517
R22057 two_stage_opamp_dummy_magic_24_0.Y.n98 two_stage_opamp_dummy_magic_24_0.Y.n47 74.5372
R22058 two_stage_opamp_dummy_magic_24_0.Y.n77 two_stage_opamp_dummy_magic_24_0.Y.n76 66.0338
R22059 two_stage_opamp_dummy_magic_24_0.Y.n80 two_stage_opamp_dummy_magic_24_0.Y.n79 66.0338
R22060 two_stage_opamp_dummy_magic_24_0.Y.n83 two_stage_opamp_dummy_magic_24_0.Y.n82 66.0338
R22061 two_stage_opamp_dummy_magic_24_0.Y.n87 two_stage_opamp_dummy_magic_24_0.Y.n86 66.0338
R22062 two_stage_opamp_dummy_magic_24_0.Y.n90 two_stage_opamp_dummy_magic_24_0.Y.n89 66.0338
R22063 two_stage_opamp_dummy_magic_24_0.Y.n93 two_stage_opamp_dummy_magic_24_0.Y.n92 66.0338
R22064 two_stage_opamp_dummy_magic_24_0.Y.n8 two_stage_opamp_dummy_magic_24_0.Y.n6 54.7984
R22065 two_stage_opamp_dummy_magic_24_0.Y.n8 two_stage_opamp_dummy_magic_24_0.Y.n7 54.4547
R22066 two_stage_opamp_dummy_magic_24_0.Y.n10 two_stage_opamp_dummy_magic_24_0.Y.n9 54.4547
R22067 two_stage_opamp_dummy_magic_24_0.Y.n12 two_stage_opamp_dummy_magic_24_0.Y.n11 54.4547
R22068 two_stage_opamp_dummy_magic_24_0.Y.n14 two_stage_opamp_dummy_magic_24_0.Y.n13 54.4547
R22069 two_stage_opamp_dummy_magic_24_0.Y.n16 two_stage_opamp_dummy_magic_24_0.Y.n15 54.4547
R22070 two_stage_opamp_dummy_magic_24_0.Y.n54 two_stage_opamp_dummy_magic_24_0.Y.t12 41.0384
R22071 two_stage_opamp_dummy_magic_24_0.Y.n68 two_stage_opamp_dummy_magic_24_0.Y.n63 40.1672
R22072 two_stage_opamp_dummy_magic_24_0.Y.n68 two_stage_opamp_dummy_magic_24_0.Y.n67 40.1672
R22073 two_stage_opamp_dummy_magic_24_0.Y.n46 two_stage_opamp_dummy_magic_24_0.Y.n44 40.1672
R22074 two_stage_opamp_dummy_magic_24_0.Y.n46 two_stage_opamp_dummy_magic_24_0.Y.n45 40.1672
R22075 two_stage_opamp_dummy_magic_24_0.Y.n37 two_stage_opamp_dummy_magic_24_0.Y.n35 40.1672
R22076 two_stage_opamp_dummy_magic_24_0.Y.n37 two_stage_opamp_dummy_magic_24_0.Y.n36 40.1672
R22077 two_stage_opamp_dummy_magic_24_0.Y.n72 two_stage_opamp_dummy_magic_24_0.Y.n71 16.3217
R22078 two_stage_opamp_dummy_magic_24_0.Y.n6 two_stage_opamp_dummy_magic_24_0.Y.t20 16.0005
R22079 two_stage_opamp_dummy_magic_24_0.Y.n6 two_stage_opamp_dummy_magic_24_0.Y.t1 16.0005
R22080 two_stage_opamp_dummy_magic_24_0.Y.n7 two_stage_opamp_dummy_magic_24_0.Y.t21 16.0005
R22081 two_stage_opamp_dummy_magic_24_0.Y.n7 two_stage_opamp_dummy_magic_24_0.Y.t14 16.0005
R22082 two_stage_opamp_dummy_magic_24_0.Y.n9 two_stage_opamp_dummy_magic_24_0.Y.t22 16.0005
R22083 two_stage_opamp_dummy_magic_24_0.Y.n9 two_stage_opamp_dummy_magic_24_0.Y.t15 16.0005
R22084 two_stage_opamp_dummy_magic_24_0.Y.n11 two_stage_opamp_dummy_magic_24_0.Y.t19 16.0005
R22085 two_stage_opamp_dummy_magic_24_0.Y.n11 two_stage_opamp_dummy_magic_24_0.Y.t17 16.0005
R22086 two_stage_opamp_dummy_magic_24_0.Y.n13 two_stage_opamp_dummy_magic_24_0.Y.t13 16.0005
R22087 two_stage_opamp_dummy_magic_24_0.Y.n13 two_stage_opamp_dummy_magic_24_0.Y.t16 16.0005
R22088 two_stage_opamp_dummy_magic_24_0.Y.n15 two_stage_opamp_dummy_magic_24_0.Y.t0 16.0005
R22089 two_stage_opamp_dummy_magic_24_0.Y.n15 two_stage_opamp_dummy_magic_24_0.Y.t18 16.0005
R22090 two_stage_opamp_dummy_magic_24_0.Y.n69 two_stage_opamp_dummy_magic_24_0.Y.n59 12.8005
R22091 two_stage_opamp_dummy_magic_24_0.Y.n76 two_stage_opamp_dummy_magic_24_0.Y.t23 11.2576
R22092 two_stage_opamp_dummy_magic_24_0.Y.n76 two_stage_opamp_dummy_magic_24_0.Y.t4 11.2576
R22093 two_stage_opamp_dummy_magic_24_0.Y.n79 two_stage_opamp_dummy_magic_24_0.Y.t6 11.2576
R22094 two_stage_opamp_dummy_magic_24_0.Y.n79 two_stage_opamp_dummy_magic_24_0.Y.t9 11.2576
R22095 two_stage_opamp_dummy_magic_24_0.Y.n82 two_stage_opamp_dummy_magic_24_0.Y.t11 11.2576
R22096 two_stage_opamp_dummy_magic_24_0.Y.n82 two_stage_opamp_dummy_magic_24_0.Y.t2 11.2576
R22097 two_stage_opamp_dummy_magic_24_0.Y.n86 two_stage_opamp_dummy_magic_24_0.Y.t3 11.2576
R22098 two_stage_opamp_dummy_magic_24_0.Y.n86 two_stage_opamp_dummy_magic_24_0.Y.t5 11.2576
R22099 two_stage_opamp_dummy_magic_24_0.Y.n89 two_stage_opamp_dummy_magic_24_0.Y.t7 11.2576
R22100 two_stage_opamp_dummy_magic_24_0.Y.n89 two_stage_opamp_dummy_magic_24_0.Y.t10 11.2576
R22101 two_stage_opamp_dummy_magic_24_0.Y.n92 two_stage_opamp_dummy_magic_24_0.Y.t8 11.2576
R22102 two_stage_opamp_dummy_magic_24_0.Y.n92 two_stage_opamp_dummy_magic_24_0.Y.t24 11.2576
R22103 two_stage_opamp_dummy_magic_24_0.Y.n17 two_stage_opamp_dummy_magic_24_0.Y.n16 10.9224
R22104 two_stage_opamp_dummy_magic_24_0.Y.n69 two_stage_opamp_dummy_magic_24_0.Y.n57 9.36264
R22105 two_stage_opamp_dummy_magic_24_0.Y.n59 two_stage_opamp_dummy_magic_24_0.Y.n58 9.3005
R22106 two_stage_opamp_dummy_magic_24_0.Y.n101 two_stage_opamp_dummy_magic_24_0.Y.n25 5.96925
R22107 two_stage_opamp_dummy_magic_24_0.Y.n93 two_stage_opamp_dummy_magic_24_0.Y.n91 5.91717
R22108 two_stage_opamp_dummy_magic_24_0.Y.n78 two_stage_opamp_dummy_magic_24_0.Y.n77 5.91717
R22109 two_stage_opamp_dummy_magic_24_0.Y.n18 two_stage_opamp_dummy_magic_24_0.Y.n17 5.68397
R22110 two_stage_opamp_dummy_magic_24_0.Y.n81 two_stage_opamp_dummy_magic_24_0.Y.n77 5.66717
R22111 two_stage_opamp_dummy_magic_24_0.Y.n19 two_stage_opamp_dummy_magic_24_0.Y.n5 5.6255
R22112 two_stage_opamp_dummy_magic_24_0.Y.n21 two_stage_opamp_dummy_magic_24_0.Y.n4 5.6255
R22113 two_stage_opamp_dummy_magic_24_0.Y.n107 two_stage_opamp_dummy_magic_24_0.Y.n1 5.6255
R22114 two_stage_opamp_dummy_magic_24_0.Y.n103 two_stage_opamp_dummy_magic_24_0.Y.n25 5.6255
R22115 two_stage_opamp_dummy_magic_24_0.Y.n71 two_stage_opamp_dummy_magic_24_0.Y.n59 5.33141
R22116 two_stage_opamp_dummy_magic_24_0.Y.n81 two_stage_opamp_dummy_magic_24_0.Y.n80 5.29217
R22117 two_stage_opamp_dummy_magic_24_0.Y.n80 two_stage_opamp_dummy_magic_24_0.Y.n78 5.29217
R22118 two_stage_opamp_dummy_magic_24_0.Y.n84 two_stage_opamp_dummy_magic_24_0.Y.n83 5.29217
R22119 two_stage_opamp_dummy_magic_24_0.Y.n83 two_stage_opamp_dummy_magic_24_0.Y.n75 5.29217
R22120 two_stage_opamp_dummy_magic_24_0.Y.n87 two_stage_opamp_dummy_magic_24_0.Y.n85 5.29217
R22121 two_stage_opamp_dummy_magic_24_0.Y.n88 two_stage_opamp_dummy_magic_24_0.Y.n87 5.29217
R22122 two_stage_opamp_dummy_magic_24_0.Y.n90 two_stage_opamp_dummy_magic_24_0.Y.n74 5.29217
R22123 two_stage_opamp_dummy_magic_24_0.Y.n91 two_stage_opamp_dummy_magic_24_0.Y.n90 5.29217
R22124 two_stage_opamp_dummy_magic_24_0.Y.n94 two_stage_opamp_dummy_magic_24_0.Y.n93 5.29217
R22125 two_stage_opamp_dummy_magic_24_0.Y.n99 two_stage_opamp_dummy_magic_24_0.Y.n26 4.5005
R22126 two_stage_opamp_dummy_magic_24_0.Y.n98 two_stage_opamp_dummy_magic_24_0.Y.n97 4.5005
R22127 two_stage_opamp_dummy_magic_24_0.Y.n99 two_stage_opamp_dummy_magic_24_0.Y.n98 4.5005
R22128 two_stage_opamp_dummy_magic_24_0.Y.n73 two_stage_opamp_dummy_magic_24_0.Y.n72 4.5005
R22129 two_stage_opamp_dummy_magic_24_0.Y.n51 two_stage_opamp_dummy_magic_24_0.Y.n50 4.5005
R22130 two_stage_opamp_dummy_magic_24_0.Y.n95 two_stage_opamp_dummy_magic_24_0.Y.n94 4.49527
R22131 two_stage_opamp_dummy_magic_24_0.Y.n52 two_stage_opamp_dummy_magic_24_0.Y.n49 2.26187
R22132 two_stage_opamp_dummy_magic_24_0.Y.n53 two_stage_opamp_dummy_magic_24_0.Y.n52 2.26187
R22133 two_stage_opamp_dummy_magic_24_0.Y.n97 two_stage_opamp_dummy_magic_24_0.Y.n96 2.24063
R22134 two_stage_opamp_dummy_magic_24_0.Y.n48 two_stage_opamp_dummy_magic_24_0.Y.n28 2.24063
R22135 two_stage_opamp_dummy_magic_24_0.Y.n56 two_stage_opamp_dummy_magic_24_0.Y.n49 2.24063
R22136 two_stage_opamp_dummy_magic_24_0.Y.n95 two_stage_opamp_dummy_magic_24_0.Y.n27 2.24063
R22137 two_stage_opamp_dummy_magic_24_0.Y.n55 two_stage_opamp_dummy_magic_24_0.Y.n54 2.24063
R22138 two_stage_opamp_dummy_magic_24_0.Y.n73 two_stage_opamp_dummy_magic_24_0.Y.n57 2.22018
R22139 two_stage_opamp_dummy_magic_24_0.Y.n101 two_stage_opamp_dummy_magic_24_0.Y.n100 1.5005
R22140 two_stage_opamp_dummy_magic_24_0.Y.n102 two_stage_opamp_dummy_magic_24_0.Y.n24 1.5005
R22141 two_stage_opamp_dummy_magic_24_0.Y.n104 two_stage_opamp_dummy_magic_24_0.Y.n103 1.5005
R22142 two_stage_opamp_dummy_magic_24_0.Y.n105 two_stage_opamp_dummy_magic_24_0.Y.n2 1.5005
R22143 two_stage_opamp_dummy_magic_24_0.Y.n107 two_stage_opamp_dummy_magic_24_0.Y.n106 1.5005
R22144 two_stage_opamp_dummy_magic_24_0.Y.n23 two_stage_opamp_dummy_magic_24_0.Y.n0 1.5005
R22145 two_stage_opamp_dummy_magic_24_0.Y.n22 two_stage_opamp_dummy_magic_24_0.Y.n21 1.5005
R22146 two_stage_opamp_dummy_magic_24_0.Y.n20 two_stage_opamp_dummy_magic_24_0.Y.n3 1.5005
R22147 two_stage_opamp_dummy_magic_24_0.Y.n73 two_stage_opamp_dummy_magic_24_0.Y.n56 0.682792
R22148 two_stage_opamp_dummy_magic_24_0.Y.n100 two_stage_opamp_dummy_magic_24_0.Y.n99 0.630708
R22149 two_stage_opamp_dummy_magic_24_0.Y.n91 two_stage_opamp_dummy_magic_24_0.Y.n88 0.6255
R22150 two_stage_opamp_dummy_magic_24_0.Y.n88 two_stage_opamp_dummy_magic_24_0.Y.n75 0.6255
R22151 two_stage_opamp_dummy_magic_24_0.Y.n78 two_stage_opamp_dummy_magic_24_0.Y.n75 0.6255
R22152 two_stage_opamp_dummy_magic_24_0.Y.n18 two_stage_opamp_dummy_magic_24_0.Y.n3 0.564601
R22153 two_stage_opamp_dummy_magic_24_0.Y.n97 two_stage_opamp_dummy_magic_24_0.Y.n73 0.46925
R22154 two_stage_opamp_dummy_magic_24_0.Y.n84 two_stage_opamp_dummy_magic_24_0.Y.n81 0.3755
R22155 two_stage_opamp_dummy_magic_24_0.Y.n85 two_stage_opamp_dummy_magic_24_0.Y.n84 0.3755
R22156 two_stage_opamp_dummy_magic_24_0.Y.n85 two_stage_opamp_dummy_magic_24_0.Y.n74 0.3755
R22157 two_stage_opamp_dummy_magic_24_0.Y.n94 two_stage_opamp_dummy_magic_24_0.Y.n74 0.3755
R22158 two_stage_opamp_dummy_magic_24_0.Y.n16 two_stage_opamp_dummy_magic_24_0.Y.n14 0.34425
R22159 two_stage_opamp_dummy_magic_24_0.Y.n14 two_stage_opamp_dummy_magic_24_0.Y.n12 0.34425
R22160 two_stage_opamp_dummy_magic_24_0.Y.n12 two_stage_opamp_dummy_magic_24_0.Y.n10 0.34425
R22161 two_stage_opamp_dummy_magic_24_0.Y.n10 two_stage_opamp_dummy_magic_24_0.Y.n8 0.34425
R22162 two_stage_opamp_dummy_magic_24_0.Y.n17 two_stage_opamp_dummy_magic_24_0.Y.n5 0.34425
R22163 two_stage_opamp_dummy_magic_24_0.Y.n5 two_stage_opamp_dummy_magic_24_0.Y.n4 0.34425
R22164 two_stage_opamp_dummy_magic_24_0.Y.n4 two_stage_opamp_dummy_magic_24_0.Y.n1 0.34425
R22165 two_stage_opamp_dummy_magic_24_0.Y.n25 two_stage_opamp_dummy_magic_24_0.Y.n1 0.34425
R22166 two_stage_opamp_dummy_magic_24_0.Y.n72 two_stage_opamp_dummy_magic_24_0.Y.n58 0.1255
R22167 two_stage_opamp_dummy_magic_24_0.Y.n58 two_stage_opamp_dummy_magic_24_0.Y.n57 0.0626438
R22168 two_stage_opamp_dummy_magic_24_0.Y.n20 two_stage_opamp_dummy_magic_24_0.Y.n19 0.0577917
R22169 two_stage_opamp_dummy_magic_24_0.Y.n21 two_stage_opamp_dummy_magic_24_0.Y.n20 0.0577917
R22170 two_stage_opamp_dummy_magic_24_0.Y.n21 two_stage_opamp_dummy_magic_24_0.Y.n0 0.0577917
R22171 two_stage_opamp_dummy_magic_24_0.Y.n107 two_stage_opamp_dummy_magic_24_0.Y.n2 0.0577917
R22172 two_stage_opamp_dummy_magic_24_0.Y.n103 two_stage_opamp_dummy_magic_24_0.Y.n2 0.0577917
R22173 two_stage_opamp_dummy_magic_24_0.Y.n103 two_stage_opamp_dummy_magic_24_0.Y.n102 0.0577917
R22174 two_stage_opamp_dummy_magic_24_0.Y.n102 two_stage_opamp_dummy_magic_24_0.Y.n101 0.0577917
R22175 two_stage_opamp_dummy_magic_24_0.Y.n22 two_stage_opamp_dummy_magic_24_0.Y.n3 0.0577917
R22176 two_stage_opamp_dummy_magic_24_0.Y.n23 two_stage_opamp_dummy_magic_24_0.Y.n22 0.0577917
R22177 two_stage_opamp_dummy_magic_24_0.Y.n106 two_stage_opamp_dummy_magic_24_0.Y.n23 0.0577917
R22178 two_stage_opamp_dummy_magic_24_0.Y.n106 two_stage_opamp_dummy_magic_24_0.Y.n105 0.0577917
R22179 two_stage_opamp_dummy_magic_24_0.Y.n105 two_stage_opamp_dummy_magic_24_0.Y.n104 0.0577917
R22180 two_stage_opamp_dummy_magic_24_0.Y.n104 two_stage_opamp_dummy_magic_24_0.Y.n24 0.0577917
R22181 two_stage_opamp_dummy_magic_24_0.Y.n100 two_stage_opamp_dummy_magic_24_0.Y.n24 0.0577917
R22182 two_stage_opamp_dummy_magic_24_0.Y.n19 two_stage_opamp_dummy_magic_24_0.Y.n18 0.054517
R22183 two_stage_opamp_dummy_magic_24_0.Y.n97 two_stage_opamp_dummy_magic_24_0.Y.n48 0.0421667
R22184 two_stage_opamp_dummy_magic_24_0.Y two_stage_opamp_dummy_magic_24_0.Y.n0 0.0369583
R22185 two_stage_opamp_dummy_magic_24_0.Y.n96 two_stage_opamp_dummy_magic_24_0.Y.n95 0.0217373
R22186 two_stage_opamp_dummy_magic_24_0.Y.n98 two_stage_opamp_dummy_magic_24_0.Y.n28 0.0217373
R22187 two_stage_opamp_dummy_magic_24_0.Y.n96 two_stage_opamp_dummy_magic_24_0.Y.n26 0.0217373
R22188 two_stage_opamp_dummy_magic_24_0.Y.n28 two_stage_opamp_dummy_magic_24_0.Y.n26 0.0217373
R22189 two_stage_opamp_dummy_magic_24_0.Y.n51 two_stage_opamp_dummy_magic_24_0.Y.n49 0.0217373
R22190 two_stage_opamp_dummy_magic_24_0.Y.n52 two_stage_opamp_dummy_magic_24_0.Y.n50 0.0217373
R22191 two_stage_opamp_dummy_magic_24_0.Y.n99 two_stage_opamp_dummy_magic_24_0.Y.n27 0.0217373
R22192 two_stage_opamp_dummy_magic_24_0.Y.n55 two_stage_opamp_dummy_magic_24_0.Y.n50 0.0217373
R22193 two_stage_opamp_dummy_magic_24_0.Y.n48 two_stage_opamp_dummy_magic_24_0.Y.n27 0.0217373
R22194 two_stage_opamp_dummy_magic_24_0.Y.n53 two_stage_opamp_dummy_magic_24_0.Y.n51 0.0217373
R22195 two_stage_opamp_dummy_magic_24_0.Y.n54 two_stage_opamp_dummy_magic_24_0.Y.n53 0.0217373
R22196 two_stage_opamp_dummy_magic_24_0.Y.n56 two_stage_opamp_dummy_magic_24_0.Y.n55 0.0217373
R22197 two_stage_opamp_dummy_magic_24_0.Y two_stage_opamp_dummy_magic_24_0.Y.n107 0.0213333
R22198 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n0 345.264
R22199 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n1 344.7
R22200 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n3 292.5
R22201 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n22 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t16 121.931
R22202 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n7 118.861
R22203 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n9 118.861
R22204 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n13 118.861
R22205 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n17 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n16 118.861
R22206 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n20 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n19 118.861
R22207 bgr_11_0.V_CMFB_S3 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n22 76.063
R22208 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n2 52.763
R22209 bgr_11_0.V_CMFB_S3 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n4 51.8547
R22210 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t2 39.4005
R22211 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t5 39.4005
R22212 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t1 39.4005
R22213 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t0 39.4005
R22214 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t4 39.4005
R22215 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t3 39.4005
R22216 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t8 19.7005
R22217 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t11 19.7005
R22218 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t15 19.7005
R22219 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t10 19.7005
R22220 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t14 19.7005
R22221 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t9 19.7005
R22222 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t7 19.7005
R22223 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t13 19.7005
R22224 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n19 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t6 19.7005
R22225 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n19 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t12 19.7005
R22226 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n22 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n21 5.90675
R22227 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n8 5.60467
R22228 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n20 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n18 5.54217
R22229 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n6 5.54217
R22230 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n10 5.04217
R22231 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n12 5.04217
R22232 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n17 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n5 5.04217
R22233 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n21 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n20 5.04217
R22234 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n6 4.97967
R22235 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n14 4.97967
R22236 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n18 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n17 4.97967
R22237 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n18 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n15 0.563
R22238 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n6 0.563
R22239 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n11 0.563
R22240 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n5 0.563
R22241 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n21 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n5 0.563
R22242 bgr_11_0.V_TOP.n23 bgr_11_0.V_TOP.n21 344.178
R22243 bgr_11_0.V_TOP.n23 bgr_11_0.V_TOP.n22 334.772
R22244 bgr_11_0.V_TOP.n1 bgr_11_0.V_TOP.t37 312.798
R22245 bgr_11_0.V_TOP bgr_11_0.V_TOP.t21 312.639
R22246 bgr_11_0.V_TOP.n36 bgr_11_0.V_TOP.t45 312.5
R22247 bgr_11_0.V_TOP.n42 bgr_11_0.V_TOP.t33 310.401
R22248 bgr_11_0.V_TOP.n41 bgr_11_0.V_TOP.t42 310.401
R22249 bgr_11_0.V_TOP.n40 bgr_11_0.V_TOP.t49 310.401
R22250 bgr_11_0.V_TOP.n39 bgr_11_0.V_TOP.t26 310.401
R22251 bgr_11_0.V_TOP.n38 bgr_11_0.V_TOP.t25 310.401
R22252 bgr_11_0.V_TOP.n37 bgr_11_0.V_TOP.t36 310.401
R22253 bgr_11_0.V_TOP.n5 bgr_11_0.V_TOP.t27 310.401
R22254 bgr_11_0.V_TOP.n4 bgr_11_0.V_TOP.t39 310.401
R22255 bgr_11_0.V_TOP.n3 bgr_11_0.V_TOP.t48 310.401
R22256 bgr_11_0.V_TOP.n2 bgr_11_0.V_TOP.t23 310.401
R22257 bgr_11_0.V_TOP.n1 bgr_11_0.V_TOP.t38 310.401
R22258 bgr_11_0.V_TOP.n34 bgr_11_0.V_TOP.t14 308
R22259 bgr_11_0.V_TOP.n7 bgr_11_0.V_TOP.t29 305.901
R22260 bgr_11_0.V_TOP.n31 bgr_11_0.V_TOP.n30 301.933
R22261 bgr_11_0.V_TOP.n29 bgr_11_0.V_TOP.n28 301.933
R22262 bgr_11_0.V_TOP.n27 bgr_11_0.V_TOP.n26 301.933
R22263 bgr_11_0.V_TOP.n24 bgr_11_0.V_TOP.n20 297.433
R22264 bgr_11_0.V_TOP.n19 bgr_11_0.V_TOP.t6 108.424
R22265 bgr_11_0.V_TOP.n32 bgr_11_0.V_TOP.t9 99.5675
R22266 bgr_11_0.V_TOP.n22 bgr_11_0.V_TOP.t11 39.4005
R22267 bgr_11_0.V_TOP.n22 bgr_11_0.V_TOP.t4 39.4005
R22268 bgr_11_0.V_TOP.n21 bgr_11_0.V_TOP.t0 39.4005
R22269 bgr_11_0.V_TOP.n21 bgr_11_0.V_TOP.t13 39.4005
R22270 bgr_11_0.V_TOP.n20 bgr_11_0.V_TOP.t12 39.4005
R22271 bgr_11_0.V_TOP.n20 bgr_11_0.V_TOP.t3 39.4005
R22272 bgr_11_0.V_TOP.n30 bgr_11_0.V_TOP.t5 39.4005
R22273 bgr_11_0.V_TOP.n30 bgr_11_0.V_TOP.t10 39.4005
R22274 bgr_11_0.V_TOP.n28 bgr_11_0.V_TOP.t8 39.4005
R22275 bgr_11_0.V_TOP.n28 bgr_11_0.V_TOP.t2 39.4005
R22276 bgr_11_0.V_TOP.n26 bgr_11_0.V_TOP.t7 39.4005
R22277 bgr_11_0.V_TOP.n26 bgr_11_0.V_TOP.t1 39.4005
R22278 bgr_11_0.V_TOP.n19 bgr_11_0.V_TOP.n18 29.1779
R22279 bgr_11_0.V_TOP.n25 bgr_11_0.V_TOP.n19 16.5063
R22280 bgr_11_0.V_TOP.n32 bgr_11_0.V_TOP.n31 4.90675
R22281 bgr_11_0.V_TOP.n8 bgr_11_0.V_TOP.t24 4.8295
R22282 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.t46 4.8295
R22283 bgr_11_0.V_TOP.n10 bgr_11_0.V_TOP.t34 4.8295
R22284 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.t18 4.8295
R22285 bgr_11_0.V_TOP.n12 bgr_11_0.V_TOP.t22 4.8295
R22286 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.t44 4.8295
R22287 bgr_11_0.V_TOP.n14 bgr_11_0.V_TOP.t47 4.8295
R22288 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.t35 4.8295
R22289 bgr_11_0.V_TOP.n16 bgr_11_0.V_TOP.t41 4.8295
R22290 bgr_11_0.V_TOP.n8 bgr_11_0.V_TOP.t32 4.5005
R22291 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.t19 4.5005
R22292 bgr_11_0.V_TOP.n10 bgr_11_0.V_TOP.t40 4.5005
R22293 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.t31 4.5005
R22294 bgr_11_0.V_TOP.n12 bgr_11_0.V_TOP.t30 4.5005
R22295 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.t17 4.5005
R22296 bgr_11_0.V_TOP.n14 bgr_11_0.V_TOP.t16 4.5005
R22297 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.t43 4.5005
R22298 bgr_11_0.V_TOP.n18 bgr_11_0.V_TOP.t20 4.5005
R22299 bgr_11_0.V_TOP.n17 bgr_11_0.V_TOP.t28 4.5005
R22300 bgr_11_0.V_TOP.n16 bgr_11_0.V_TOP.t15 4.5005
R22301 bgr_11_0.V_TOP.n7 bgr_11_0.V_TOP.n6 4.5005
R22302 bgr_11_0.V_TOP.n33 bgr_11_0.V_TOP.n0 4.5005
R22303 bgr_11_0.V_TOP.n35 bgr_11_0.V_TOP.n34 4.5005
R22304 bgr_11_0.V_TOP.n25 bgr_11_0.V_TOP.n24 4.5005
R22305 bgr_11_0.V_TOP.n24 bgr_11_0.V_TOP.n23 1.59425
R22306 bgr_11_0.V_TOP.n33 bgr_11_0.V_TOP.n32 1.21925
R22307 bgr_11_0.V_TOP.n27 bgr_11_0.V_TOP.n25 1.1255
R22308 bgr_11_0.V_TOP.n29 bgr_11_0.V_TOP.n27 1.1255
R22309 bgr_11_0.V_TOP.n31 bgr_11_0.V_TOP.n29 1.1255
R22310 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.n8 0.3295
R22311 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.n10 0.3295
R22312 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.n12 0.3295
R22313 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.n14 0.3295
R22314 bgr_11_0.V_TOP.n18 bgr_11_0.V_TOP.n17 0.3295
R22315 bgr_11_0.V_TOP.n17 bgr_11_0.V_TOP.n16 0.3295
R22316 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.n9 0.2825
R22317 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.n11 0.2825
R22318 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.n13 0.2825
R22319 bgr_11_0.V_TOP.n16 bgr_11_0.V_TOP.n15 0.2825
R22320 bgr_11_0.V_TOP.n2 bgr_11_0.V_TOP.n1 0.28175
R22321 bgr_11_0.V_TOP.n3 bgr_11_0.V_TOP.n2 0.28175
R22322 bgr_11_0.V_TOP.n4 bgr_11_0.V_TOP.n3 0.28175
R22323 bgr_11_0.V_TOP.n5 bgr_11_0.V_TOP.n4 0.28175
R22324 bgr_11_0.V_TOP.n6 bgr_11_0.V_TOP.n5 0.28175
R22325 bgr_11_0.V_TOP.n36 bgr_11_0.V_TOP.n35 0.28175
R22326 bgr_11_0.V_TOP.n37 bgr_11_0.V_TOP.n36 0.28175
R22327 bgr_11_0.V_TOP.n38 bgr_11_0.V_TOP.n37 0.28175
R22328 bgr_11_0.V_TOP.n39 bgr_11_0.V_TOP.n38 0.28175
R22329 bgr_11_0.V_TOP.n40 bgr_11_0.V_TOP.n39 0.28175
R22330 bgr_11_0.V_TOP.n41 bgr_11_0.V_TOP.n40 0.28175
R22331 bgr_11_0.V_TOP.n42 bgr_11_0.V_TOP.n41 0.28175
R22332 bgr_11_0.V_TOP.n6 bgr_11_0.V_TOP.n0 0.141125
R22333 bgr_11_0.V_TOP.n35 bgr_11_0.V_TOP.n0 0.141125
R22334 bgr_11_0.V_TOP bgr_11_0.V_TOP.n42 0.141125
R22335 bgr_11_0.V_TOP.n33 bgr_11_0.V_TOP.n7 0.141125
R22336 bgr_11_0.V_TOP.n34 bgr_11_0.V_TOP.n33 0.141125
R22337 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t7 651.405
R22338 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t8 648.03
R22339 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t9 537.922
R22340 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t4 117.243
R22341 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n1 107.266
R22342 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n4 105.016
R22343 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n2 105.016
R22344 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t2 13.1338
R22345 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t6 13.1338
R22346 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t3 13.1338
R22347 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t0 13.1338
R22348 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t5 13.1338
R22349 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t1 13.1338
R22350 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n5 7.32862
R22351 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n6 3.98488
R22352 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n3 2.2505
R22353 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n0 1.73488
R22354 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n7 1.53175
R22355 bgr_11_0.1st_Vout_1.n12 bgr_11_0.1st_Vout_1.t29 363.909
R22356 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.t13 351.88
R22357 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.n22 299.25
R22358 bgr_11_0.1st_Vout_1.n14 bgr_11_0.1st_Vout_1.n13 299.25
R22359 bgr_11_0.1st_Vout_1.n18 bgr_11_0.1st_Vout_1.n17 297.807
R22360 bgr_11_0.1st_Vout_1.n20 bgr_11_0.1st_Vout_1.t30 194.809
R22361 bgr_11_0.1st_Vout_1.n20 bgr_11_0.1st_Vout_1.t10 194.809
R22362 bgr_11_0.1st_Vout_1.n15 bgr_11_0.1st_Vout_1.t28 194.809
R22363 bgr_11_0.1st_Vout_1.n15 bgr_11_0.1st_Vout_1.t19 194.809
R22364 bgr_11_0.1st_Vout_1.n21 bgr_11_0.1st_Vout_1.n20 163.097
R22365 bgr_11_0.1st_Vout_1.n16 bgr_11_0.1st_Vout_1.n15 163.097
R22366 bgr_11_0.1st_Vout_1.n18 bgr_11_0.1st_Vout_1.t2 49.4474
R22367 bgr_11_0.1st_Vout_1.n22 bgr_11_0.1st_Vout_1.t1 39.4005
R22368 bgr_11_0.1st_Vout_1.n22 bgr_11_0.1st_Vout_1.t3 39.4005
R22369 bgr_11_0.1st_Vout_1.n13 bgr_11_0.1st_Vout_1.t5 39.4005
R22370 bgr_11_0.1st_Vout_1.n13 bgr_11_0.1st_Vout_1.t4 39.4005
R22371 bgr_11_0.1st_Vout_1.n17 bgr_11_0.1st_Vout_1.t6 39.4005
R22372 bgr_11_0.1st_Vout_1.n17 bgr_11_0.1st_Vout_1.t0 39.4005
R22373 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t27 4.8295
R22374 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t14 4.8295
R22375 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.t32 4.8295
R22376 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t22 4.8295
R22377 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.t25 4.8295
R22378 bgr_11_0.1st_Vout_1.n5 bgr_11_0.1st_Vout_1.t12 4.8295
R22379 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.t16 4.8295
R22380 bgr_11_0.1st_Vout_1.n7 bgr_11_0.1st_Vout_1.t7 4.8295
R22381 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.t24 4.8295
R22382 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t18 4.5005
R22383 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t23 4.5005
R22384 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.t26 4.5005
R22385 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t31 4.5005
R22386 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.t17 4.5005
R22387 bgr_11_0.1st_Vout_1.n5 bgr_11_0.1st_Vout_1.t21 4.5005
R22388 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.t8 4.5005
R22389 bgr_11_0.1st_Vout_1.n7 bgr_11_0.1st_Vout_1.t11 4.5005
R22390 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.t15 4.5005
R22391 bgr_11_0.1st_Vout_1.n10 bgr_11_0.1st_Vout_1.t20 4.5005
R22392 bgr_11_0.1st_Vout_1.n11 bgr_11_0.1st_Vout_1.t9 4.5005
R22393 bgr_11_0.1st_Vout_1.n19 bgr_11_0.1st_Vout_1.n18 1.44719
R22394 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.n1 0.3295
R22395 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.n3 0.3295
R22396 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.n5 0.3295
R22397 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.n7 0.3295
R22398 bgr_11_0.1st_Vout_1.n10 bgr_11_0.1st_Vout_1.n9 0.3295
R22399 bgr_11_0.1st_Vout_1.n11 bgr_11_0.1st_Vout_1.n10 0.3295
R22400 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.n2 0.2825
R22401 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.n4 0.2825
R22402 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.n6 0.2825
R22403 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.n8 0.2825
R22404 bgr_11_0.1st_Vout_1.n19 bgr_11_0.1st_Vout_1.n16 0.2505
R22405 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.n21 0.2505
R22406 bgr_11_0.1st_Vout_1.n14 bgr_11_0.1st_Vout_1.n12 0.21925
R22407 bgr_11_0.1st_Vout_1.n16 bgr_11_0.1st_Vout_1.n14 0.1255
R22408 bgr_11_0.1st_Vout_1.n21 bgr_11_0.1st_Vout_1.n19 0.1255
R22409 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.n0 0.09425
R22410 bgr_11_0.1st_Vout_1.n12 bgr_11_0.1st_Vout_1.n11 10.102
R22411 bgr_11_0.cap_res1.t20 bgr_11_0.cap_res1.t13 121.983
R22412 bgr_11_0.cap_res1.t9 bgr_11_0.cap_res1.t17 0.1603
R22413 bgr_11_0.cap_res1.t16 bgr_11_0.cap_res1.t19 0.1603
R22414 bgr_11_0.cap_res1.t8 bgr_11_0.cap_res1.t15 0.1603
R22415 bgr_11_0.cap_res1.t1 bgr_11_0.cap_res1.t7 0.1603
R22416 bgr_11_0.cap_res1.t6 bgr_11_0.cap_res1.t14 0.1603
R22417 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t10 0.159278
R22418 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t3 0.159278
R22419 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t11 0.159278
R22420 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t18 0.159278
R22421 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t9 0.1368
R22422 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t5 0.1368
R22423 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t16 0.1368
R22424 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t12 0.1368
R22425 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t8 0.1368
R22426 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t4 0.1368
R22427 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t1 0.1368
R22428 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t0 0.1368
R22429 bgr_11_0.cap_res1.n0 bgr_11_0.cap_res1.t6 0.1368
R22430 bgr_11_0.cap_res1.n0 bgr_11_0.cap_res1.t2 0.1368
R22431 bgr_11_0.cap_res1.t10 bgr_11_0.cap_res1.n0 0.00152174
R22432 bgr_11_0.cap_res1.t3 bgr_11_0.cap_res1.n1 0.00152174
R22433 bgr_11_0.cap_res1.t11 bgr_11_0.cap_res1.n2 0.00152174
R22434 bgr_11_0.cap_res1.t18 bgr_11_0.cap_res1.n3 0.00152174
R22435 bgr_11_0.cap_res1.t13 bgr_11_0.cap_res1.n4 0.00152174
R22436 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t3 119.785
R22437 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n0 107.121
R22438 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n1 97.4332
R22439 bgr_11_0.V_CMFB_S4 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n20 70.4693
R22440 bgr_11_0.V_CMFB_S4 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n2 39.7505
R22441 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n5 24.288
R22442 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n7 24.288
R22443 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n11 24.288
R22444 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n14 24.288
R22445 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n17 24.288
R22446 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t2 24.0005
R22447 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t0 24.0005
R22448 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t1 24.0005
R22449 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t4 24.0005
R22450 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t8 8.0005
R22451 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t11 8.0005
R22452 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t5 8.0005
R22453 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t10 8.0005
R22454 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t14 8.0005
R22455 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t9 8.0005
R22456 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t7 8.0005
R22457 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t13 8.0005
R22458 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t6 8.0005
R22459 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t12 8.0005
R22460 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n16 5.7505
R22461 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n4 5.7505
R22462 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n6 5.7505
R22463 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n19 5.6255
R22464 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n8 5.188
R22465 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n4 5.188
R22466 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n10 5.188
R22467 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n12 5.188
R22468 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n3 5.188
R22469 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n15 5.188
R22470 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n18 5.188
R22471 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n13 0.563
R22472 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n4 0.563
R22473 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n9 0.563
R22474 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n3 0.563
R22475 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n3 0.563
R22476 bgr_11_0.NFET_GATE_10uA.n3 bgr_11_0.NFET_GATE_10uA.t18 369.534
R22477 bgr_11_0.NFET_GATE_10uA.n2 bgr_11_0.NFET_GATE_10uA.t20 369.534
R22478 bgr_11_0.NFET_GATE_10uA.n8 bgr_11_0.NFET_GATE_10uA.t22 369.534
R22479 bgr_11_0.NFET_GATE_10uA.n7 bgr_11_0.NFET_GATE_10uA.t19 369.534
R22480 bgr_11_0.NFET_GATE_10uA.n14 bgr_11_0.NFET_GATE_10uA.t12 369.534
R22481 bgr_11_0.NFET_GATE_10uA.n11 bgr_11_0.NFET_GATE_10uA.t10 369.534
R22482 bgr_11_0.NFET_GATE_10uA.n17 bgr_11_0.NFET_GATE_10uA.t1 369.534
R22483 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n1 360.288
R22484 bgr_11_0.NFET_GATE_10uA.n18 bgr_11_0.NFET_GATE_10uA.t6 249.034
R22485 bgr_11_0.NFET_GATE_10uA.n5 bgr_11_0.NFET_GATE_10uA.t17 192.8
R22486 bgr_11_0.NFET_GATE_10uA.n4 bgr_11_0.NFET_GATE_10uA.t5 192.8
R22487 bgr_11_0.NFET_GATE_10uA.n3 bgr_11_0.NFET_GATE_10uA.t11 192.8
R22488 bgr_11_0.NFET_GATE_10uA.n2 bgr_11_0.NFET_GATE_10uA.t8 192.8
R22489 bgr_11_0.NFET_GATE_10uA.n8 bgr_11_0.NFET_GATE_10uA.t14 192.8
R22490 bgr_11_0.NFET_GATE_10uA.n7 bgr_11_0.NFET_GATE_10uA.t7 192.8
R22491 bgr_11_0.NFET_GATE_10uA.n14 bgr_11_0.NFET_GATE_10uA.t9 192.8
R22492 bgr_11_0.NFET_GATE_10uA.n11 bgr_11_0.NFET_GATE_10uA.t16 192.8
R22493 bgr_11_0.NFET_GATE_10uA.n12 bgr_11_0.NFET_GATE_10uA.t15 192.8
R22494 bgr_11_0.NFET_GATE_10uA.n13 bgr_11_0.NFET_GATE_10uA.t21 192.8
R22495 bgr_11_0.NFET_GATE_10uA.n17 bgr_11_0.NFET_GATE_10uA.t13 192.8
R22496 bgr_11_0.NFET_GATE_10uA.n5 bgr_11_0.NFET_GATE_10uA.n4 176.733
R22497 bgr_11_0.NFET_GATE_10uA.n4 bgr_11_0.NFET_GATE_10uA.n3 176.733
R22498 bgr_11_0.NFET_GATE_10uA.n12 bgr_11_0.NFET_GATE_10uA.n11 176.733
R22499 bgr_11_0.NFET_GATE_10uA.n13 bgr_11_0.NFET_GATE_10uA.n12 176.733
R22500 bgr_11_0.NFET_GATE_10uA.n10 bgr_11_0.NFET_GATE_10uA.n6 167.843
R22501 bgr_11_0.NFET_GATE_10uA.n10 bgr_11_0.NFET_GATE_10uA.n9 166.343
R22502 bgr_11_0.NFET_GATE_10uA.n16 bgr_11_0.NFET_GATE_10uA.n15 166.343
R22503 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n18 166.343
R22504 bgr_11_0.NFET_GATE_10uA.n19 bgr_11_0.NFET_GATE_10uA.n0 141.752
R22505 bgr_11_0.NFET_GATE_10uA.n6 bgr_11_0.NFET_GATE_10uA.n5 56.2338
R22506 bgr_11_0.NFET_GATE_10uA.n6 bgr_11_0.NFET_GATE_10uA.n2 56.2338
R22507 bgr_11_0.NFET_GATE_10uA.n9 bgr_11_0.NFET_GATE_10uA.n8 56.2338
R22508 bgr_11_0.NFET_GATE_10uA.n9 bgr_11_0.NFET_GATE_10uA.n7 56.2338
R22509 bgr_11_0.NFET_GATE_10uA.n15 bgr_11_0.NFET_GATE_10uA.n14 56.2338
R22510 bgr_11_0.NFET_GATE_10uA.n15 bgr_11_0.NFET_GATE_10uA.n13 56.2338
R22511 bgr_11_0.NFET_GATE_10uA.n18 bgr_11_0.NFET_GATE_10uA.n17 56.2338
R22512 bgr_11_0.NFET_GATE_10uA.n1 bgr_11_0.NFET_GATE_10uA.t4 39.4005
R22513 bgr_11_0.NFET_GATE_10uA.n1 bgr_11_0.NFET_GATE_10uA.t3 39.4005
R22514 bgr_11_0.NFET_GATE_10uA.t0 bgr_11_0.NFET_GATE_10uA.n19 24.0005
R22515 bgr_11_0.NFET_GATE_10uA.n19 bgr_11_0.NFET_GATE_10uA.t2 24.0005
R22516 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n16 2.01612
R22517 bgr_11_0.NFET_GATE_10uA.n16 bgr_11_0.NFET_GATE_10uA.n10 1.5005
R22518 two_stage_opamp_dummy_magic_24_0.V_err_gate.n2 two_stage_opamp_dummy_magic_24_0.V_err_gate.t8 479.322
R22519 two_stage_opamp_dummy_magic_24_0.V_err_gate.n2 two_stage_opamp_dummy_magic_24_0.V_err_gate.t6 479.322
R22520 two_stage_opamp_dummy_magic_24_0.V_err_gate.n6 two_stage_opamp_dummy_magic_24_0.V_err_gate.t7 479.322
R22521 two_stage_opamp_dummy_magic_24_0.V_err_gate.n6 two_stage_opamp_dummy_magic_24_0.V_err_gate.t9 479.322
R22522 two_stage_opamp_dummy_magic_24_0.V_err_gate.n3 two_stage_opamp_dummy_magic_24_0.V_err_gate.n1 178.625
R22523 two_stage_opamp_dummy_magic_24_0.V_err_gate.n5 two_stage_opamp_dummy_magic_24_0.V_err_gate.n4 177.987
R22524 two_stage_opamp_dummy_magic_24_0.V_err_gate two_stage_opamp_dummy_magic_24_0.V_err_gate.n0 170.357
R22525 two_stage_opamp_dummy_magic_24_0.V_err_gate.n3 two_stage_opamp_dummy_magic_24_0.V_err_gate.n2 165.8
R22526 two_stage_opamp_dummy_magic_24_0.V_err_gate two_stage_opamp_dummy_magic_24_0.V_err_gate.n6 165.8
R22527 two_stage_opamp_dummy_magic_24_0.V_err_gate.n0 two_stage_opamp_dummy_magic_24_0.V_err_gate.t2 24.0005
R22528 two_stage_opamp_dummy_magic_24_0.V_err_gate.n0 two_stage_opamp_dummy_magic_24_0.V_err_gate.t3 24.0005
R22529 two_stage_opamp_dummy_magic_24_0.V_err_gate.n4 two_stage_opamp_dummy_magic_24_0.V_err_gate.t4 15.7605
R22530 two_stage_opamp_dummy_magic_24_0.V_err_gate.n4 two_stage_opamp_dummy_magic_24_0.V_err_gate.t1 15.7605
R22531 two_stage_opamp_dummy_magic_24_0.V_err_gate.n1 two_stage_opamp_dummy_magic_24_0.V_err_gate.t0 15.7605
R22532 two_stage_opamp_dummy_magic_24_0.V_err_gate.n1 two_stage_opamp_dummy_magic_24_0.V_err_gate.t5 15.7605
R22533 two_stage_opamp_dummy_magic_24_0.V_err_gate two_stage_opamp_dummy_magic_24_0.V_err_gate.n5 1.76612
R22534 two_stage_opamp_dummy_magic_24_0.V_err_gate.n5 two_stage_opamp_dummy_magic_24_0.V_err_gate.n3 0.641125
R22535 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t28 610.534
R22536 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t18 610.534
R22537 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t16 433.8
R22538 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t21 433.8
R22539 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t30 433.8
R22540 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t19 433.8
R22541 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t26 433.8
R22542 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t14 433.8
R22543 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t24 433.8
R22544 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t12 433.8
R22545 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t29 433.8
R22546 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t31 433.8
R22547 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t20 433.8
R22548 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t27 433.8
R22549 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t15 433.8
R22550 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t25 433.8
R22551 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t13 433.8
R22552 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t23 433.8
R22553 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t17 433.8
R22554 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t22 433.8
R22555 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n31 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n23 287.264
R22556 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n25 287.264
R22557 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n28 287.264
R22558 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n24 287.264
R22559 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n10 176.733
R22560 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n9 176.733
R22561 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n8 176.733
R22562 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n7 176.733
R22563 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n6 176.733
R22564 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n5 176.733
R22565 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n4 176.733
R22566 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n3 176.733
R22567 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n13 176.733
R22568 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n14 176.733
R22569 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n15 176.733
R22570 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n16 176.733
R22571 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n17 176.733
R22572 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n18 176.733
R22573 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n20 176.733
R22574 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.V_tail_gate.n12 161.754
R22575 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.V_tail_gate.n22 161.754
R22576 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n2 63.1128
R22577 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n0 63.112
R22578 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n31 63.112
R22579 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n31 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n30 52.5725
R22580 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n2 52.5725
R22581 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n26 52.01
R22582 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n30 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n29 52.01
R22583 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.V_tail_gate.n32 50.4989
R22584 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.V_tail_gate.n33 50.4989
R22585 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_24_0.V_tail_gate 46.7517
R22586 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n11 45.5227
R22587 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n19 45.5227
R22588 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n21 45.5227
R22589 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n12 45.5227
R22590 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t8 39.4005
R22591 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t4 39.4005
R22592 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t10 39.4005
R22593 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t7 39.4005
R22594 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t9 39.4005
R22595 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t5 39.4005
R22596 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t6 39.4005
R22597 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t11 39.4005
R22598 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.V_tail_gate.n1 16.3608
R22599 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n32 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t0 16.0005
R22600 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n32 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t2 16.0005
R22601 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n33 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t3 16.0005
R22602 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n33 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t1 16.0005
R22603 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.V_tail_gate.n0 7.03346
R22604 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n30 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n27 0.563
R22605 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n1 0.340713
R22606 bgr_11_0.START_UP_NFET1 bgr_11_0.START_UP_NFET1.t0 141.653
R22607 bgr_11_0.V_mir1.n11 bgr_11_0.V_mir1.t18 310.488
R22608 bgr_11_0.V_mir1.n5 bgr_11_0.V_mir1.t13 310.488
R22609 bgr_11_0.V_mir1.n0 bgr_11_0.V_mir1.t17 310.488
R22610 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.n8 297.433
R22611 bgr_11_0.V_mir1.n4 bgr_11_0.V_mir1.n3 297.433
R22612 bgr_11_0.V_mir1.n15 bgr_11_0.V_mir1.n14 297.433
R22613 bgr_11_0.V_mir1.n13 bgr_11_0.V_mir1.t11 184.097
R22614 bgr_11_0.V_mir1.n7 bgr_11_0.V_mir1.t9 184.097
R22615 bgr_11_0.V_mir1.n2 bgr_11_0.V_mir1.t7 184.097
R22616 bgr_11_0.V_mir1.n12 bgr_11_0.V_mir1.n11 167.094
R22617 bgr_11_0.V_mir1.n6 bgr_11_0.V_mir1.n5 167.094
R22618 bgr_11_0.V_mir1.n1 bgr_11_0.V_mir1.n0 167.094
R22619 bgr_11_0.V_mir1.n14 bgr_11_0.V_mir1.n13 161.3
R22620 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.n7 161.3
R22621 bgr_11_0.V_mir1.n4 bgr_11_0.V_mir1.n2 161.3
R22622 bgr_11_0.V_mir1.n11 bgr_11_0.V_mir1.t14 120.501
R22623 bgr_11_0.V_mir1.n12 bgr_11_0.V_mir1.t5 120.501
R22624 bgr_11_0.V_mir1.n5 bgr_11_0.V_mir1.t15 120.501
R22625 bgr_11_0.V_mir1.n6 bgr_11_0.V_mir1.t3 120.501
R22626 bgr_11_0.V_mir1.n0 bgr_11_0.V_mir1.t16 120.501
R22627 bgr_11_0.V_mir1.n1 bgr_11_0.V_mir1.t1 120.501
R22628 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.t0 50.2004
R22629 bgr_11_0.V_mir1.n13 bgr_11_0.V_mir1.n12 40.7027
R22630 bgr_11_0.V_mir1.n7 bgr_11_0.V_mir1.n6 40.7027
R22631 bgr_11_0.V_mir1.n2 bgr_11_0.V_mir1.n1 40.7027
R22632 bgr_11_0.V_mir1.n8 bgr_11_0.V_mir1.t10 39.4005
R22633 bgr_11_0.V_mir1.n8 bgr_11_0.V_mir1.t4 39.4005
R22634 bgr_11_0.V_mir1.n3 bgr_11_0.V_mir1.t8 39.4005
R22635 bgr_11_0.V_mir1.n3 bgr_11_0.V_mir1.t2 39.4005
R22636 bgr_11_0.V_mir1.t12 bgr_11_0.V_mir1.n15 39.4005
R22637 bgr_11_0.V_mir1.n15 bgr_11_0.V_mir1.t6 39.4005
R22638 bgr_11_0.V_mir1.n10 bgr_11_0.V_mir1.n4 6.6255
R22639 bgr_11_0.V_mir1.n14 bgr_11_0.V_mir1.n10 6.6255
R22640 bgr_11_0.V_mir1.n10 bgr_11_0.V_mir1.n9 4.5005
R22641 two_stage_opamp_dummy_magic_24_0.V_tot.n2 two_stage_opamp_dummy_magic_24_0.V_tot.t4 648.343
R22642 two_stage_opamp_dummy_magic_24_0.V_tot.n1 two_stage_opamp_dummy_magic_24_0.V_tot.t5 648.343
R22643 two_stage_opamp_dummy_magic_24_0.V_tot.n3 two_stage_opamp_dummy_magic_24_0.V_tot.t3 117.591
R22644 two_stage_opamp_dummy_magic_24_0.V_tot.n0 two_stage_opamp_dummy_magic_24_0.V_tot.t2 117.591
R22645 two_stage_opamp_dummy_magic_24_0.V_tot.n0 two_stage_opamp_dummy_magic_24_0.V_tot.t1 108.424
R22646 two_stage_opamp_dummy_magic_24_0.V_tot.t0 two_stage_opamp_dummy_magic_24_0.V_tot.n3 108.424
R22647 two_stage_opamp_dummy_magic_24_0.V_tot.n1 two_stage_opamp_dummy_magic_24_0.V_tot.n0 43.0496
R22648 two_stage_opamp_dummy_magic_24_0.V_tot.n3 two_stage_opamp_dummy_magic_24_0.V_tot.n2 43.0496
R22649 two_stage_opamp_dummy_magic_24_0.V_tot.n2 two_stage_opamp_dummy_magic_24_0.V_tot.n1 1.563
R22650 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t5 573.044
R22651 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t1 433.8
R22652 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n0 184.643
R22653 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n1 163.978
R22654 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n2 33.0088
R22655 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t3 15.7605
R22656 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t4 15.7605
R22657 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t2 9.6005
R22658 two_stage_opamp_dummy_magic_24_0.err_amp_mir.t0 two_stage_opamp_dummy_magic_24_0.err_amp_mir.n3 9.6005
R22659 two_stage_opamp_dummy_magic_24_0.V_err_p.n1 two_stage_opamp_dummy_magic_24_0.V_err_p.n0 365.07
R22660 two_stage_opamp_dummy_magic_24_0.V_err_p.n0 two_stage_opamp_dummy_magic_24_0.V_err_p.t3 15.7605
R22661 two_stage_opamp_dummy_magic_24_0.V_err_p.n0 two_stage_opamp_dummy_magic_24_0.V_err_p.t1 15.7605
R22662 two_stage_opamp_dummy_magic_24_0.V_err_p.n1 two_stage_opamp_dummy_magic_24_0.V_err_p.t0 15.7605
R22663 two_stage_opamp_dummy_magic_24_0.V_err_p.t2 two_stage_opamp_dummy_magic_24_0.V_err_p.n1 15.7605
R22664 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n0 344.837
R22665 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n1 344.274
R22666 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n3 292.5
R22667 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n22 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t10 121.785
R22668 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n7 118.861
R22669 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n9 118.861
R22670 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n13 118.861
R22671 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n17 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n16 118.861
R22672 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n20 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n19 118.861
R22673 bgr_11_0.V_CMFB_S1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n22 78.0317
R22674 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n2 52.3363
R22675 bgr_11_0.V_CMFB_S1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n4 52.2813
R22676 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t15 39.4005
R22677 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t12 39.4005
R22678 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t14 39.4005
R22679 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t13 39.4005
R22680 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t11 39.4005
R22681 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t16 39.4005
R22682 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t8 19.7005
R22683 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t3 19.7005
R22684 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t9 19.7005
R22685 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t4 19.7005
R22686 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t1 19.7005
R22687 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t5 19.7005
R22688 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t0 19.7005
R22689 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t7 19.7005
R22690 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n19 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t2 19.7005
R22691 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n19 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t6 19.7005
R22692 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n22 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n21 5.90675
R22693 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n8 5.60467
R22694 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n20 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n18 5.54217
R22695 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n6 5.54217
R22696 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n10 5.04217
R22697 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n12 5.04217
R22698 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n17 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n5 5.04217
R22699 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n21 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n20 5.04217
R22700 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n6 4.97967
R22701 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n14 4.97967
R22702 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n18 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n17 4.97967
R22703 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n18 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n15 0.563
R22704 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n6 0.563
R22705 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n11 0.563
R22706 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n5 0.563
R22707 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n21 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n5 0.563
R22708 a_6350_30238.t0 a_6350_30238.t1 178.133
R22709 bgr_11_0.Vin+ bgr_11_0.Vin+.t6 529.879
R22710 bgr_11_0.Vin+.n0 bgr_11_0.Vin+.t4 148.653
R22711 bgr_11_0.Vin+.n0 bgr_11_0.Vin+.t5 125.418
R22712 bgr_11_0.Vin+.n3 bgr_11_0.Vin+.n1 106.609
R22713 bgr_11_0.Vin+.n3 bgr_11_0.Vin+.n2 104.484
R22714 bgr_11_0.Vin+.n4 bgr_11_0.Vin+.n0 25.0809
R22715 bgr_11_0.Vin+.n4 bgr_11_0.Vin+.n3 18.7817
R22716 bgr_11_0.Vin+.n2 bgr_11_0.Vin+.t2 13.1338
R22717 bgr_11_0.Vin+.n2 bgr_11_0.Vin+.t1 13.1338
R22718 bgr_11_0.Vin+.n1 bgr_11_0.Vin+.t0 13.1338
R22719 bgr_11_0.Vin+.n1 bgr_11_0.Vin+.t3 13.1338
R22720 bgr_11_0.Vin+ bgr_11_0.Vin+.n4 6.53175
R22721 a_6540_22450.n11 a_6540_22450.t18 310.488
R22722 a_6540_22450.n5 a_6540_22450.t13 310.488
R22723 a_6540_22450.n0 a_6540_22450.t14 310.488
R22724 a_6540_22450.n9 a_6540_22450.n8 297.433
R22725 a_6540_22450.n4 a_6540_22450.n3 297.433
R22726 a_6540_22450.n15 a_6540_22450.n14 297.433
R22727 a_6540_22450.n13 a_6540_22450.t7 184.097
R22728 a_6540_22450.n7 a_6540_22450.t5 184.097
R22729 a_6540_22450.n2 a_6540_22450.t3 184.097
R22730 a_6540_22450.n12 a_6540_22450.n11 167.094
R22731 a_6540_22450.n6 a_6540_22450.n5 167.094
R22732 a_6540_22450.n1 a_6540_22450.n0 167.094
R22733 a_6540_22450.n14 a_6540_22450.n13 161.3
R22734 a_6540_22450.n9 a_6540_22450.n7 161.3
R22735 a_6540_22450.n4 a_6540_22450.n2 161.3
R22736 a_6540_22450.n11 a_6540_22450.t15 120.501
R22737 a_6540_22450.n12 a_6540_22450.t11 120.501
R22738 a_6540_22450.n5 a_6540_22450.t17 120.501
R22739 a_6540_22450.n6 a_6540_22450.t1 120.501
R22740 a_6540_22450.n0 a_6540_22450.t16 120.501
R22741 a_6540_22450.n1 a_6540_22450.t9 120.501
R22742 a_6540_22450.n9 a_6540_22450.t0 50.2004
R22743 a_6540_22450.n13 a_6540_22450.n12 40.7027
R22744 a_6540_22450.n7 a_6540_22450.n6 40.7027
R22745 a_6540_22450.n2 a_6540_22450.n1 40.7027
R22746 a_6540_22450.n8 a_6540_22450.t2 39.4005
R22747 a_6540_22450.n8 a_6540_22450.t6 39.4005
R22748 a_6540_22450.n3 a_6540_22450.t10 39.4005
R22749 a_6540_22450.n3 a_6540_22450.t4 39.4005
R22750 a_6540_22450.t12 a_6540_22450.n15 39.4005
R22751 a_6540_22450.n15 a_6540_22450.t8 39.4005
R22752 a_6540_22450.n10 a_6540_22450.n4 6.6255
R22753 a_6540_22450.n14 a_6540_22450.n10 6.6255
R22754 a_6540_22450.n10 a_6540_22450.n9 4.5005
R22755 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t10 119.785
R22756 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n0 107.121
R22757 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n1 97.4332
R22758 bgr_11_0.V_CMFB_S2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n20 66.3443
R22759 bgr_11_0.V_CMFB_S2 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n2 30.9724
R22760 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n5 24.288
R22761 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n7 24.288
R22762 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n11 24.288
R22763 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n14 24.288
R22764 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n17 24.288
R22765 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t14 24.0005
R22766 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t11 24.0005
R22767 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t12 24.0005
R22768 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t13 24.0005
R22769 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t9 8.0005
R22770 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t4 8.0005
R22771 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t0 8.0005
R22772 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t5 8.0005
R22773 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t2 8.0005
R22774 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t6 8.0005
R22775 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t1 8.0005
R22776 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t8 8.0005
R22777 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t3 8.0005
R22778 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t7 8.0005
R22779 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n16 5.7505
R22780 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n4 5.7505
R22781 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n6 5.7505
R22782 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n19 5.6255
R22783 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n8 5.188
R22784 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n4 5.188
R22785 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n10 5.188
R22786 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n12 5.188
R22787 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n3 5.188
R22788 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n15 5.188
R22789 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n18 5.188
R22790 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n13 0.563
R22791 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n4 0.563
R22792 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n9 0.563
R22793 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n3 0.563
R22794 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n3 0.563
R22795 VIN-.n0 VIN-.t7 1097.62
R22796 VIN- VIN-.n9 433.019
R22797 VIN-.n9 VIN-.t10 273.134
R22798 VIN-.n0 VIN-.t9 273.134
R22799 VIN-.n1 VIN-.t3 273.134
R22800 VIN-.n2 VIN-.t8 273.134
R22801 VIN-.n3 VIN-.t1 273.134
R22802 VIN-.n4 VIN-.t5 273.134
R22803 VIN-.n5 VIN-.t2 273.134
R22804 VIN-.n6 VIN-.t6 273.134
R22805 VIN-.n7 VIN-.t0 273.134
R22806 VIN-.n8 VIN-.t4 273.134
R22807 VIN-.n9 VIN-.n8 176.733
R22808 VIN-.n8 VIN-.n7 176.733
R22809 VIN-.n7 VIN-.n6 176.733
R22810 VIN-.n6 VIN-.n5 176.733
R22811 VIN-.n5 VIN-.n4 176.733
R22812 VIN-.n4 VIN-.n3 176.733
R22813 VIN-.n3 VIN-.n2 176.733
R22814 VIN-.n2 VIN-.n1 176.733
R22815 VIN-.n1 VIN-.n0 176.733
R22816 two_stage_opamp_dummy_magic_24_0.VD1.n1 two_stage_opamp_dummy_magic_24_0.VD1.n0 49.7255
R22817 two_stage_opamp_dummy_magic_24_0.VD1.n25 two_stage_opamp_dummy_magic_24_0.VD1.n24 49.7255
R22818 two_stage_opamp_dummy_magic_24_0.VD1.n27 two_stage_opamp_dummy_magic_24_0.VD1.n9 49.7255
R22819 two_stage_opamp_dummy_magic_24_0.VD1.n21 two_stage_opamp_dummy_magic_24_0.VD1.n12 49.7255
R22820 two_stage_opamp_dummy_magic_24_0.VD1.n11 two_stage_opamp_dummy_magic_24_0.VD1.n10 49.7255
R22821 two_stage_opamp_dummy_magic_24_0.VD1.n15 two_stage_opamp_dummy_magic_24_0.VD1.n14 49.3505
R22822 two_stage_opamp_dummy_magic_24_0.VD1.n8 two_stage_opamp_dummy_magic_24_0.VD1.n7 49.3505
R22823 two_stage_opamp_dummy_magic_24_0.VD1.n31 two_stage_opamp_dummy_magic_24_0.VD1.n30 49.3505
R22824 two_stage_opamp_dummy_magic_24_0.VD1.n35 two_stage_opamp_dummy_magic_24_0.VD1.n34 49.3505
R22825 two_stage_opamp_dummy_magic_24_0.VD1.n5 two_stage_opamp_dummy_magic_24_0.VD1.n4 49.3505
R22826 two_stage_opamp_dummy_magic_24_0.VD1.n18 two_stage_opamp_dummy_magic_24_0.VD1.n17 49.3505
R22827 two_stage_opamp_dummy_magic_24_0.VD1.n14 two_stage_opamp_dummy_magic_24_0.VD1.t1 16.0005
R22828 two_stage_opamp_dummy_magic_24_0.VD1.n14 two_stage_opamp_dummy_magic_24_0.VD1.t12 16.0005
R22829 two_stage_opamp_dummy_magic_24_0.VD1.n7 two_stage_opamp_dummy_magic_24_0.VD1.t13 16.0005
R22830 two_stage_opamp_dummy_magic_24_0.VD1.n7 two_stage_opamp_dummy_magic_24_0.VD1.t0 16.0005
R22831 two_stage_opamp_dummy_magic_24_0.VD1.n30 two_stage_opamp_dummy_magic_24_0.VD1.t14 16.0005
R22832 two_stage_opamp_dummy_magic_24_0.VD1.n30 two_stage_opamp_dummy_magic_24_0.VD1.t18 16.0005
R22833 two_stage_opamp_dummy_magic_24_0.VD1.n34 two_stage_opamp_dummy_magic_24_0.VD1.t16 16.0005
R22834 two_stage_opamp_dummy_magic_24_0.VD1.n34 two_stage_opamp_dummy_magic_24_0.VD1.t20 16.0005
R22835 two_stage_opamp_dummy_magic_24_0.VD1.n4 two_stage_opamp_dummy_magic_24_0.VD1.t15 16.0005
R22836 two_stage_opamp_dummy_magic_24_0.VD1.n4 two_stage_opamp_dummy_magic_24_0.VD1.t19 16.0005
R22837 two_stage_opamp_dummy_magic_24_0.VD1.n0 two_stage_opamp_dummy_magic_24_0.VD1.t3 16.0005
R22838 two_stage_opamp_dummy_magic_24_0.VD1.n0 two_stage_opamp_dummy_magic_24_0.VD1.t10 16.0005
R22839 two_stage_opamp_dummy_magic_24_0.VD1.n24 two_stage_opamp_dummy_magic_24_0.VD1.t4 16.0005
R22840 two_stage_opamp_dummy_magic_24_0.VD1.n24 two_stage_opamp_dummy_magic_24_0.VD1.t8 16.0005
R22841 two_stage_opamp_dummy_magic_24_0.VD1.n9 two_stage_opamp_dummy_magic_24_0.VD1.t2 16.0005
R22842 two_stage_opamp_dummy_magic_24_0.VD1.n9 two_stage_opamp_dummy_magic_24_0.VD1.t7 16.0005
R22843 two_stage_opamp_dummy_magic_24_0.VD1.n12 two_stage_opamp_dummy_magic_24_0.VD1.t5 16.0005
R22844 two_stage_opamp_dummy_magic_24_0.VD1.n12 two_stage_opamp_dummy_magic_24_0.VD1.t9 16.0005
R22845 two_stage_opamp_dummy_magic_24_0.VD1.n17 two_stage_opamp_dummy_magic_24_0.VD1.t17 16.0005
R22846 two_stage_opamp_dummy_magic_24_0.VD1.n17 two_stage_opamp_dummy_magic_24_0.VD1.t21 16.0005
R22847 two_stage_opamp_dummy_magic_24_0.VD1.n10 two_stage_opamp_dummy_magic_24_0.VD1.t6 16.0005
R22848 two_stage_opamp_dummy_magic_24_0.VD1.n10 two_stage_opamp_dummy_magic_24_0.VD1.t11 16.0005
R22849 two_stage_opamp_dummy_magic_24_0.VD1.n25 two_stage_opamp_dummy_magic_24_0.VD1.n3 6.29217
R22850 two_stage_opamp_dummy_magic_24_0.VD1.n28 two_stage_opamp_dummy_magic_24_0.VD1.n27 6.29217
R22851 two_stage_opamp_dummy_magic_24_0.VD1.n21 two_stage_opamp_dummy_magic_24_0.VD1.n20 6.29217
R22852 two_stage_opamp_dummy_magic_24_0.VD1.n13 two_stage_opamp_dummy_magic_24_0.VD1.n11 6.29217
R22853 two_stage_opamp_dummy_magic_24_0.VD1.n32 two_stage_opamp_dummy_magic_24_0.VD1.n8 5.438
R22854 two_stage_opamp_dummy_magic_24_0.VD1.n16 two_stage_opamp_dummy_magic_24_0.VD1.n15 5.438
R22855 two_stage_opamp_dummy_magic_24_0.VD1.n28 two_stage_opamp_dummy_magic_24_0.VD1.n8 5.31821
R22856 two_stage_opamp_dummy_magic_24_0.VD1.n15 two_stage_opamp_dummy_magic_24_0.VD1.n13 5.31821
R22857 two_stage_opamp_dummy_magic_24_0.VD1.n31 two_stage_opamp_dummy_magic_24_0.VD1.n29 5.08383
R22858 two_stage_opamp_dummy_magic_24_0.VD1.n36 two_stage_opamp_dummy_magic_24_0.VD1.n35 5.08383
R22859 two_stage_opamp_dummy_magic_24_0.VD1.n5 two_stage_opamp_dummy_magic_24_0.VD1.n2 5.08383
R22860 two_stage_opamp_dummy_magic_24_0.VD1.n19 two_stage_opamp_dummy_magic_24_0.VD1.n18 5.08383
R22861 two_stage_opamp_dummy_magic_24_0.VD1.n27 two_stage_opamp_dummy_magic_24_0.VD1.n26 5.063
R22862 two_stage_opamp_dummy_magic_24_0.VD1.n22 two_stage_opamp_dummy_magic_24_0.VD1.n11 5.063
R22863 two_stage_opamp_dummy_magic_24_0.VD1.n32 two_stage_opamp_dummy_magic_24_0.VD1.n31 4.8755
R22864 two_stage_opamp_dummy_magic_24_0.VD1.n35 two_stage_opamp_dummy_magic_24_0.VD1.n33 4.8755
R22865 two_stage_opamp_dummy_magic_24_0.VD1.n6 two_stage_opamp_dummy_magic_24_0.VD1.n5 4.8755
R22866 two_stage_opamp_dummy_magic_24_0.VD1.n18 two_stage_opamp_dummy_magic_24_0.VD1.n16 4.8755
R22867 two_stage_opamp_dummy_magic_24_0.VD1 two_stage_opamp_dummy_magic_24_0.VD1.n37 4.60467
R22868 two_stage_opamp_dummy_magic_24_0.VD1.n26 two_stage_opamp_dummy_magic_24_0.VD1.n25 4.5005
R22869 two_stage_opamp_dummy_magic_24_0.VD1.n23 two_stage_opamp_dummy_magic_24_0.VD1.n1 4.5005
R22870 two_stage_opamp_dummy_magic_24_0.VD1.n22 two_stage_opamp_dummy_magic_24_0.VD1.n21 4.5005
R22871 two_stage_opamp_dummy_magic_24_0.VD1 two_stage_opamp_dummy_magic_24_0.VD1.n1 1.688
R22872 two_stage_opamp_dummy_magic_24_0.VD1.n26 two_stage_opamp_dummy_magic_24_0.VD1.n23 0.563
R22873 two_stage_opamp_dummy_magic_24_0.VD1.n23 two_stage_opamp_dummy_magic_24_0.VD1.n22 0.563
R22874 two_stage_opamp_dummy_magic_24_0.VD1.n33 two_stage_opamp_dummy_magic_24_0.VD1.n32 0.563
R22875 two_stage_opamp_dummy_magic_24_0.VD1.n33 two_stage_opamp_dummy_magic_24_0.VD1.n6 0.563
R22876 two_stage_opamp_dummy_magic_24_0.VD1.n16 two_stage_opamp_dummy_magic_24_0.VD1.n6 0.563
R22877 two_stage_opamp_dummy_magic_24_0.VD1.n19 two_stage_opamp_dummy_magic_24_0.VD1.n13 0.234875
R22878 two_stage_opamp_dummy_magic_24_0.VD1.n20 two_stage_opamp_dummy_magic_24_0.VD1.n19 0.234875
R22879 two_stage_opamp_dummy_magic_24_0.VD1.n20 two_stage_opamp_dummy_magic_24_0.VD1.n2 0.234875
R22880 two_stage_opamp_dummy_magic_24_0.VD1.n37 two_stage_opamp_dummy_magic_24_0.VD1.n2 0.234875
R22881 two_stage_opamp_dummy_magic_24_0.VD1.n37 two_stage_opamp_dummy_magic_24_0.VD1.n36 0.234875
R22882 two_stage_opamp_dummy_magic_24_0.VD1.n36 two_stage_opamp_dummy_magic_24_0.VD1.n3 0.234875
R22883 two_stage_opamp_dummy_magic_24_0.VD1.n29 two_stage_opamp_dummy_magic_24_0.VD1.n3 0.234875
R22884 two_stage_opamp_dummy_magic_24_0.VD1.n29 two_stage_opamp_dummy_magic_24_0.VD1.n28 0.234875
R22885 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t8 447.279
R22886 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t4 446.967
R22887 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t9 446.967
R22888 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t7 446.967
R22889 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t5 344.772
R22890 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n8 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t6 281.168
R22891 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t3 281.168
R22892 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t2 281.168
R22893 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n8 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n7 205.946
R22894 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n6 205.946
R22895 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n4 165.8
R22896 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n9 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n8 165.8
R22897 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n10 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t1 108.615
R22898 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t0 108.615
R22899 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n5 63.4857
R22900 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n4 51.5193
R22901 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n10 15.6567
R22902 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n3 10.5317
R22903 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n10 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n9 6.0005
R22904 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n2 6.0005
R22905 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n9 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n4 0.313
R22906 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n1 0.313
R22907 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n0 0.313
R22908 bgr_11_0.cap_res2.t0 bgr_11_0.cap_res2.t15 121.931
R22909 bgr_11_0.cap_res2.t10 bgr_11_0.cap_res2.t4 0.1603
R22910 bgr_11_0.cap_res2.t14 bgr_11_0.cap_res2.t9 0.1603
R22911 bgr_11_0.cap_res2.t8 bgr_11_0.cap_res2.t3 0.1603
R22912 bgr_11_0.cap_res2.t2 bgr_11_0.cap_res2.t16 0.1603
R22913 bgr_11_0.cap_res2.t6 bgr_11_0.cap_res2.t1 0.1603
R22914 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t11 0.159278
R22915 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t7 0.159278
R22916 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t13 0.159278
R22917 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t19 0.159278
R22918 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t20 0.1368
R22919 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t10 0.1368
R22920 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t5 0.1368
R22921 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t14 0.1368
R22922 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t18 0.1368
R22923 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t8 0.1368
R22924 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t12 0.1368
R22925 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t2 0.1368
R22926 bgr_11_0.cap_res2.n0 bgr_11_0.cap_res2.t17 0.1368
R22927 bgr_11_0.cap_res2.n0 bgr_11_0.cap_res2.t6 0.1368
R22928 bgr_11_0.cap_res2.t11 bgr_11_0.cap_res2.n0 0.00152174
R22929 bgr_11_0.cap_res2.t7 bgr_11_0.cap_res2.n1 0.00152174
R22930 bgr_11_0.cap_res2.t13 bgr_11_0.cap_res2.n2 0.00152174
R22931 bgr_11_0.cap_res2.t19 bgr_11_0.cap_res2.n3 0.00152174
R22932 bgr_11_0.cap_res2.t15 bgr_11_0.cap_res2.n4 0.00152174
R22933 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 807.99
R22934 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 172.969
R22935 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n142 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 84.0884
R22936 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 83.5719
R22937 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 83.5719
R22938 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 83.5719
R22939 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 83.5719
R22940 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 83.5719
R22941 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 83.5719
R22942 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 83.5719
R22943 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 83.5719
R22944 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 83.5719
R22945 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 83.5719
R22946 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 83.5719
R22947 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 83.5719
R22948 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 83.5719
R22949 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 83.5719
R22950 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 83.5719
R22951 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 83.5719
R22952 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 83.5719
R22953 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 83.5719
R22954 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 83.5719
R22955 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 83.5719
R22956 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 83.5719
R22957 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R22958 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 83.5719
R22959 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 73.8495
R22960 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 73.8495
R22961 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 73.3165
R22962 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 73.3165
R22963 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 73.3165
R22964 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 73.3165
R22965 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 73.3165
R22966 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 73.19
R22967 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 73.19
R22968 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 73.19
R22969 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 73.19
R22970 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 73.19
R22971 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 73.19
R22972 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 65.0299
R22973 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 65.0299
R22974 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 26.074
R22975 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 26.074
R22976 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 26.074
R22977 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 26.074
R22978 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 26.074
R22979 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 26.074
R22980 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 26.074
R22981 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 26.074
R22982 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 26.074
R22983 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 26.074
R22984 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 25.7843
R22985 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 25.7843
R22986 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 25.7843
R22987 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 25.7843
R22988 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 25.7843
R22989 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 25.7843
R22990 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 9.3005
R22991 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 9.3005
R22992 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R22993 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 9.3005
R22994 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 9.3005
R22995 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R22996 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 9.3005
R22997 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 9.3005
R22998 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 9.3005
R22999 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 9.3005
R23000 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R23001 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 9.3005
R23002 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 9.3005
R23003 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 9.3005
R23004 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 9.3005
R23005 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R23006 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 9.3005
R23007 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 9.3005
R23008 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 9.3005
R23009 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R23010 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 9.3005
R23011 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 9.3005
R23012 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 9.3005
R23013 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 9.3005
R23014 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R23015 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 9.3005
R23016 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 9.3005
R23017 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 9.3005
R23018 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 9.3005
R23019 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 9.3005
R23020 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 9.3005
R23021 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 9.3005
R23022 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 9.3005
R23023 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 9.3005
R23024 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 9.3005
R23025 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 9.3005
R23026 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 9.3005
R23027 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 9.3005
R23028 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 9.3005
R23029 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 9.3005
R23030 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 9.3005
R23031 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 9.3005
R23032 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 9.3005
R23033 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 9.3005
R23034 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 9.3005
R23035 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 9.3005
R23036 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 9.3005
R23037 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 9.3005
R23038 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 9.3005
R23039 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 9.3005
R23040 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 9.3005
R23041 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 9.3005
R23042 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 9.3005
R23043 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 9.3005
R23044 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 4.64654
R23045 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 4.64654
R23046 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 4.64654
R23047 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 4.64654
R23048 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 4.64654
R23049 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 4.64654
R23050 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 4.64654
R23051 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 4.64654
R23052 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 4.64654
R23053 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 2.36206
R23054 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 2.36206
R23055 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 2.36206
R23056 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 2.36206
R23057 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 2.19742
R23058 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 2.19742
R23059 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 2.19742
R23060 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 1.56363
R23061 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 1.56363
R23062 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 1.5505
R23063 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 1.5505
R23064 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 1.5505
R23065 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 1.5505
R23066 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 1.5505
R23067 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 1.5505
R23068 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 1.5505
R23069 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 1.5505
R23070 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 1.5505
R23071 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 1.5505
R23072 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 1.5505
R23073 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 1.5505
R23074 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 1.5505
R23075 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 1.5505
R23076 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 1.5505
R23077 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 1.5505
R23078 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n143 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n142 1.5505
R23079 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n145 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n144 1.5505
R23080 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R23081 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 1.25468
R23082 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.25468
R23083 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 1.25468
R23084 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 1.25468
R23085 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 1.25468
R23086 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.25468
R23087 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 1.19225
R23088 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 1.19225
R23089 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 1.19225
R23090 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 1.19225
R23091 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 1.19225
R23092 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n142 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.14402
R23093 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.07024
R23094 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 1.07024
R23095 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 1.07024
R23096 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 1.07024
R23097 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.07024
R23098 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 1.07024
R23099 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 1.0237
R23100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.0237
R23101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 1.0237
R23102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 1.0237
R23103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 1.0237
R23104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.0237
R23105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 0.885803
R23106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 0.885803
R23107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 0.885803
R23108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.885803
R23109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 0.885803
R23110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 0.885803
R23111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.885803
R23112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.885803
R23113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 0.812055
R23114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.812055
R23115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 0.77514
R23116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 0.77514
R23117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 0.77514
R23118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 0.77514
R23119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 0.77514
R23120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.77514
R23121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.77514
R23122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 0.77514
R23123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R23124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 0.756696
R23125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 0.756696
R23126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.756696
R23127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R23128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R23129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R23130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.756696
R23131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 0.711459
R23132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.711459
R23133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n145 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 0.701365
R23134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.647417
R23135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 0.647417
R23136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 0.590702
R23137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 0.590702
R23138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 0.590702
R23139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.590702
R23140 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 0.590702
R23141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 0.590702
R23142 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.576566
R23143 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.576566
R23144 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.530034
R23145 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 0.530034
R23146 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 0.290206
R23147 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 0.290206
R23148 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 0.290206
R23149 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.290206
R23150 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 0.290206
R23151 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 0.290206
R23152 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 0.290206
R23153 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 0.290206
R23154 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R23155 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R23156 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R23157 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R23158 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 0.203382
R23159 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n145 0.203382
R23160 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 0.154071
R23161 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.154071
R23162 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n143 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.154071
R23163 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 0.154071
R23164 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 0.137464
R23165 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 0.137464
R23166 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 0.134964
R23167 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 0.134964
R23168 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 0.0183571
R23169 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 0.0183571
R23170 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.0183571
R23171 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.0183571
R23172 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 0.0183571
R23173 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.0183571
R23174 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.0183571
R23175 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 0.0183571
R23176 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.0183571
R23177 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n144 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R23178 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n144 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n143 0.0183571
R23179 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R23180 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 0.0183571
R23181 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.0183571
R23182 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.0183571
R23183 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.0183571
R23184 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 0.0183571
R23185 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.0183571
R23186 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.0106786
R23187 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.0106786
R23188 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.0106786
R23189 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 0.00992001
R23190 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 0.00992001
R23191 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00992001
R23192 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 0.00992001
R23193 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 0.00992001
R23194 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00992001
R23195 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 0.00992001
R23196 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 0.00992001
R23197 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 0.00992001
R23198 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 0.00992001
R23199 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 0.00992001
R23200 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.00992001
R23201 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 0.00992001
R23202 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.00992001
R23203 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 0.00992001
R23204 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.00992001
R23205 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 0.00992001
R23206 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 0.00992001
R23207 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 0.00817857
R23208 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 0.00817857
R23209 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.00817857
R23210 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.00817857
R23211 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 0.00817857
R23212 two_stage_opamp_dummy_magic_24_0.Vb2_2.n2 two_stage_opamp_dummy_magic_24_0.Vb2_2.t6 661.375
R23213 two_stage_opamp_dummy_magic_24_0.Vb2_2.n4 two_stage_opamp_dummy_magic_24_0.Vb2_2.t3 661.375
R23214 two_stage_opamp_dummy_magic_24_0.Vb2_2.t7 two_stage_opamp_dummy_magic_24_0.Vb2_2.n0 213.131
R23215 two_stage_opamp_dummy_magic_24_0.Vb2_2.n3 two_stage_opamp_dummy_magic_24_0.Vb2_2.t4 213.131
R23216 two_stage_opamp_dummy_magic_24_0.Vb2_2.n6 two_stage_opamp_dummy_magic_24_0.Vb2_2.n1 155.123
R23217 two_stage_opamp_dummy_magic_24_0.Vb2_2.t0 two_stage_opamp_dummy_magic_24_0.Vb2_2.t7 146.155
R23218 two_stage_opamp_dummy_magic_24_0.Vb2_2.t4 two_stage_opamp_dummy_magic_24_0.Vb2_2.t0 146.155
R23219 two_stage_opamp_dummy_magic_24_0.Vb2_2.t8 two_stage_opamp_dummy_magic_24_0.Vb2_2.n0 76.2576
R23220 two_stage_opamp_dummy_magic_24_0.Vb2_2.n3 two_stage_opamp_dummy_magic_24_0.Vb2_2.t5 76.2576
R23221 two_stage_opamp_dummy_magic_24_0.Vb2_2.n7 two_stage_opamp_dummy_magic_24_0.Vb2_2.n6 66.4336
R23222 two_stage_opamp_dummy_magic_24_0.Vb2_2.n1 two_stage_opamp_dummy_magic_24_0.Vb2_2.t9 21.8894
R23223 two_stage_opamp_dummy_magic_24_0.Vb2_2.n1 two_stage_opamp_dummy_magic_24_0.Vb2_2.t2 21.8894
R23224 two_stage_opamp_dummy_magic_24_0.Vb2_2.t8 two_stage_opamp_dummy_magic_24_0.Vb2_2.n7 11.2576
R23225 two_stage_opamp_dummy_magic_24_0.Vb2_2.n7 two_stage_opamp_dummy_magic_24_0.Vb2_2.t1 11.2576
R23226 two_stage_opamp_dummy_magic_24_0.Vb2_2.n5 two_stage_opamp_dummy_magic_24_0.Vb2_2.n4 5.1255
R23227 two_stage_opamp_dummy_magic_24_0.Vb2_2.n6 two_stage_opamp_dummy_magic_24_0.Vb2_2.n5 4.92976
R23228 two_stage_opamp_dummy_magic_24_0.Vb2_2.n5 two_stage_opamp_dummy_magic_24_0.Vb2_2.n2 4.7505
R23229 two_stage_opamp_dummy_magic_24_0.Vb2_2.n4 two_stage_opamp_dummy_magic_24_0.Vb2_2.n3 1.888
R23230 two_stage_opamp_dummy_magic_24_0.Vb2_2.n2 two_stage_opamp_dummy_magic_24_0.Vb2_2.n0 1.888
R23231 two_stage_opamp_dummy_magic_24_0.V_err_mir_p two_stage_opamp_dummy_magic_24_0.V_err_mir_p.n0 187.315
R23232 two_stage_opamp_dummy_magic_24_0.V_err_mir_p two_stage_opamp_dummy_magic_24_0.V_err_mir_p.n1 177.755
R23233 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.t1 15.7605
R23234 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.t3 15.7605
R23235 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.t2 15.7605
R23236 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_24_0.V_err_mir_p.t0 15.7605
R23237 a_13940_n594.t0 a_13940_n594.t1 169.905
R23238 two_stage_opamp_dummy_magic_24_0.V_p_mir.n0 two_stage_opamp_dummy_magic_24_0.V_p_mir.t3 16.0005
R23239 two_stage_opamp_dummy_magic_24_0.V_p_mir.n0 two_stage_opamp_dummy_magic_24_0.V_p_mir.t2 16.0005
R23240 two_stage_opamp_dummy_magic_24_0.V_p_mir.t1 two_stage_opamp_dummy_magic_24_0.V_p_mir.n1 9.6005
R23241 two_stage_opamp_dummy_magic_24_0.V_p_mir.n1 two_stage_opamp_dummy_magic_24_0.V_p_mir.t0 9.6005
R23242 two_stage_opamp_dummy_magic_24_0.V_p_mir.n1 two_stage_opamp_dummy_magic_24_0.V_p_mir.n0 89.9887
R23243 a_13840_3288.t0 a_13840_3288.t1 294.339
R23244 bgr_11_0.START_UP.n4 bgr_11_0.START_UP.t7 238.322
R23245 bgr_11_0.START_UP.n4 bgr_11_0.START_UP.t6 238.322
R23246 bgr_11_0.START_UP.n5 bgr_11_0.START_UP.n4 167.332
R23247 bgr_11_0.START_UP.n0 bgr_11_0.START_UP.t5 130.001
R23248 bgr_11_0.START_UP.n3 bgr_11_0.START_UP.n1 111.796
R23249 bgr_11_0.START_UP.n3 bgr_11_0.START_UP.n2 105.171
R23250 bgr_11_0.START_UP.n0 bgr_11_0.START_UP.t4 81.7074
R23251 bgr_11_0.START_UP bgr_11_0.START_UP.n0 36.8552
R23252 bgr_11_0.START_UP bgr_11_0.START_UP.n5 15.3755
R23253 bgr_11_0.START_UP.n1 bgr_11_0.START_UP.t0 13.1338
R23254 bgr_11_0.START_UP.n1 bgr_11_0.START_UP.t2 13.1338
R23255 bgr_11_0.START_UP.n2 bgr_11_0.START_UP.t1 13.1338
R23256 bgr_11_0.START_UP.n2 bgr_11_0.START_UP.t3 13.1338
R23257 bgr_11_0.START_UP.n5 bgr_11_0.START_UP.n3 4.21925
R23258 a_11420_30238.t0 a_11420_30238.t1 178.133
R23259 bgr_11_0.Vin-.n8 bgr_11_0.Vin-.t8 539.797
R23260 bgr_11_0.Vin-.n7 bgr_11_0.Vin-.n6 351.865
R23261 bgr_11_0.Vin-.n18 bgr_11_0.Vin-.n17 141.667
R23262 bgr_11_0.Vin-.n9 bgr_11_0.Vin-.t7 117.817
R23263 bgr_11_0.Vin-.n5 bgr_11_0.Vin-.n3 109.204
R23264 bgr_11_0.Vin-.n5 bgr_11_0.Vin-.n4 104.829
R23265 bgr_11_0.Vin-.n19 bgr_11_0.Vin-.n18 84.0884
R23266 bgr_11_0.Vin-.n14 bgr_11_0.Vin-.n13 83.5719
R23267 bgr_11_0.Vin-.n15 bgr_11_0.Vin-.n0 83.5719
R23268 bgr_11_0.Vin-.n16 bgr_11_0.Vin-.n1 83.5719
R23269 bgr_11_0.Vin-.n11 bgr_11_0.Vin-.t4 65.0299
R23270 bgr_11_0.Vin-.n6 bgr_11_0.Vin-.t6 39.4005
R23271 bgr_11_0.Vin-.n6 bgr_11_0.Vin-.t5 39.4005
R23272 bgr_11_0.Vin-.n15 bgr_11_0.Vin-.n14 26.074
R23273 bgr_11_0.Vin-.n16 bgr_11_0.Vin-.n15 26.074
R23274 bgr_11_0.Vin-.n18 bgr_11_0.Vin-.n16 26.074
R23275 bgr_11_0.Vin-.n10 bgr_11_0.Vin-.n9 24.3755
R23276 bgr_11_0.Vin-.n9 bgr_11_0.Vin-.n8 17.6255
R23277 bgr_11_0.Vin-.n4 bgr_11_0.Vin-.t1 13.1338
R23278 bgr_11_0.Vin-.n4 bgr_11_0.Vin-.t2 13.1338
R23279 bgr_11_0.Vin-.n3 bgr_11_0.Vin-.t3 13.1338
R23280 bgr_11_0.Vin-.n3 bgr_11_0.Vin-.t0 13.1338
R23281 bgr_11_0.Vin-.n8 bgr_11_0.Vin-.n7 11.6567
R23282 bgr_11_0.Vin-.n7 bgr_11_0.Vin-.n5 3.8755
R23283 bgr_11_0.Vin-.n20 bgr_11_0.Vin-.n19 1.56836
R23284 bgr_11_0.Vin-.n13 bgr_11_0.Vin-.n11 1.56363
R23285 bgr_11_0.Vin-.n21 bgr_11_0.Vin-.n20 1.5505
R23286 bgr_11_0.Vin-.n12 bgr_11_0.Vin-.n2 1.5505
R23287 bgr_11_0.Vin-.n19 bgr_11_0.Vin-.n1 1.14402
R23288 bgr_11_0.Vin-.n12 bgr_11_0.Vin-.n0 0.885803
R23289 bgr_11_0.Vin-.n13 bgr_11_0.Vin-.n12 0.77514
R23290 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_11_0.Vin-.n0 0.756696
R23291 bgr_11_0.Vin-.n21 bgr_11_0.Vin-.n1 0.701365
R23292 bgr_11_0.Vin-.n11 bgr_11_0.Vin-.n10 0.530034
R23293 bgr_11_0.Vin-.n14 bgr_11_0.Vin-.t4 0.290206
R23294 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_11_0.Vin-.n21 0.203382
R23295 bgr_11_0.Vin-.n20 bgr_11_0.Vin-.n2 0.0183571
R23296 bgr_11_0.Vin-.n10 bgr_11_0.Vin-.n2 0.00817857
R23297 a_11300_30238.t0 a_11300_30238.t1 222.28
R23298 a_11950_28880.t0 a_11950_28880.t1 178.133
R23299 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t3 661.375
R23300 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t0 661.375
R23301 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n6 213.131
R23302 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t4 213.131
R23303 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t7 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t1 146.155
R23304 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t7 146.155
R23305 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t2 76.2576
R23306 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n7 76.2576
R23307 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n1 72.5885
R23308 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n2 66.4444
R23309 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t8 11.2576
R23310 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t5 11.2576
R23311 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t10 11.2576
R23312 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.t9 11.2576
R23313 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n4 5.1255
R23314 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n3 4.91892
R23315 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n0 4.7505
R23316 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n5 1.888
R23317 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_24_0.Vb2_Vb3.n0 1.888
R23318 a_3690_3288.t0 a_3690_3288.t1 294.339
R23319 a_13960_3288.t0 a_13960_3288.t1 169.905
R23320 a_3830_n594.t0 a_3830_n594.t1 169.905
R23321 two_stage_opamp_dummy_magic_24_0.err_amp_out.n1 two_stage_opamp_dummy_magic_24_0.err_amp_out.t4 1282.55
R23322 two_stage_opamp_dummy_magic_24_0.err_amp_out.n1 two_stage_opamp_dummy_magic_24_0.err_amp_out.n0 179.382
R23323 two_stage_opamp_dummy_magic_24_0.err_amp_out.n2 two_stage_opamp_dummy_magic_24_0.err_amp_out.n1 39.3422
R23324 two_stage_opamp_dummy_magic_24_0.err_amp_out.n0 two_stage_opamp_dummy_magic_24_0.err_amp_out.t3 15.7605
R23325 two_stage_opamp_dummy_magic_24_0.err_amp_out.n0 two_stage_opamp_dummy_magic_24_0.err_amp_out.t0 15.7605
R23326 two_stage_opamp_dummy_magic_24_0.err_amp_out.t1 two_stage_opamp_dummy_magic_24_0.err_amp_out.n2 9.6005
R23327 two_stage_opamp_dummy_magic_24_0.err_amp_out.n2 two_stage_opamp_dummy_magic_24_0.err_amp_out.t2 9.6005
R23328 a_11300_28630.t0 a_11300_28630.t1 178.133
R23329 bgr_11_0.V_p_1.n0 bgr_11_0.V_p_1.t2 99.8322
R23330 bgr_11_0.V_p_1.t0 bgr_11_0.V_p_1.n0 9.6005
R23331 bgr_11_0.V_p_1.n0 bgr_11_0.V_p_1.t1 9.6005
R23332 a_5700_30088.t0 a_5700_30088.t1 178.133
R23333 a_5820_28824.t0 a_5820_28824.t1 178.133
R23334 a_6470_28630.t0 a_6470_28630.t1 178.133
R23335 a_12070_30088.t0 a_12070_30088.t1 178.133
R23336 a_3810_3288.t0 a_3810_3288.t1 169.905
R23337 bgr_11_0.V_CUR_REF_REG bgr_11_0.V_CUR_REF_REG.t3 701.501
R23338 bgr_11_0.V_CUR_REF_REG.n1 bgr_11_0.V_CUR_REF_REG.n0 357.647
R23339 bgr_11_0.V_CUR_REF_REG.n1 bgr_11_0.V_CUR_REF_REG.t0 135.239
R23340 bgr_11_0.V_CUR_REF_REG.n0 bgr_11_0.V_CUR_REF_REG.t1 39.4005
R23341 bgr_11_0.V_CUR_REF_REG.n0 bgr_11_0.V_CUR_REF_REG.t2 39.4005
R23342 bgr_11_0.V_CUR_REF_REG bgr_11_0.V_CUR_REF_REG.n1 5.79738
R23343 bgr_11_0.V_p_2.n0 bgr_11_0.V_p_2.t2 142.558
R23344 bgr_11_0.V_p_2.t0 bgr_11_0.V_p_2.n0 9.6005
R23345 bgr_11_0.V_p_2.n0 bgr_11_0.V_p_2.t1 9.6005
C0 VOUT+ VOUT- 0.118487f
C1 a_4440_7230# VDDA 0.098742f
C2 two_stage_opamp_dummy_magic_24_0.cap_res_Y VDDA 7.86427f
C3 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.V_TOP 0.04106f
C4 bgr_11_0.PFET_GATE_10uA bgr_11_0.V_CUR_REF_REG 0.347737f
C5 bgr_11_0.V_CUR_REF_REG two_stage_opamp_dummy_magic_24_0.Vb3 1.51248f
C6 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_24_0.Vb1 0.091782f
C7 two_stage_opamp_dummy_magic_24_0.Vb3 a_5760_7230# 0.01595f
C8 two_stage_opamp_dummy_magic_24_0.X VDDA 6.95716f
C9 two_stage_opamp_dummy_magic_24_0.V_tail_gate VDDA 7.953129f
C10 two_stage_opamp_dummy_magic_24_0.Vb3 two_stage_opamp_dummy_magic_24_0.Vb1 0.292093f
C11 two_stage_opamp_dummy_magic_24_0.Vb1 m2_6870_1200# 0.051771f
C12 two_stage_opamp_dummy_magic_24_0.cap_res_Y two_stage_opamp_dummy_magic_24_0.cap_res_X 0.345243f
C13 two_stage_opamp_dummy_magic_24_0.V_err_gate two_stage_opamp_dummy_magic_24_0.X 0.091085f
C14 two_stage_opamp_dummy_magic_24_0.V_err_gate two_stage_opamp_dummy_magic_24_0.V_tail_gate 0.169255f
C15 two_stage_opamp_dummy_magic_24_0.Y VDDA 6.99024f
C16 two_stage_opamp_dummy_magic_24_0.cap_res_Y VOUT+ 50.921898f
C17 two_stage_opamp_dummy_magic_24_0.X two_stage_opamp_dummy_magic_24_0.cap_res_X 0.056362f
C18 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.cap_res_X 2.08159f
C19 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref two_stage_opamp_dummy_magic_24_0.cap_res_Y 0.157188f
C20 bgr_11_0.V_TOP VDDA 16.3436f
C21 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter two_stage_opamp_dummy_magic_24_0.Vb3 0.016733f
C22 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage m2_6870_1200# 0.04f
C23 bgr_11_0.V_TOP two_stage_opamp_dummy_magic_24_0.V_err_gate 0.104556f
C24 two_stage_opamp_dummy_magic_24_0.V_tail_gate VOUT+ 1.318f
C25 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref two_stage_opamp_dummy_magic_24_0.V_tail_gate 0.130497f
C26 two_stage_opamp_dummy_magic_24_0.Y VOUT+ 3.89657f
C27 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref two_stage_opamp_dummy_magic_24_0.Y 0.087335f
C28 two_stage_opamp_dummy_magic_24_0.cap_res_Y VOUT- 0.011897f
C29 bgr_11_0.V_TOP bgr_11_0.START_UP 1.37378f
C30 bgr_11_0.PFET_GATE_10uA VDDA 10.121f
C31 two_stage_opamp_dummy_magic_24_0.VD2 VIN+ 0.533278f
C32 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref bgr_11_0.V_TOP 0.939477f
C33 two_stage_opamp_dummy_magic_24_0.V_tail_gate VOUT- 1.318f
C34 two_stage_opamp_dummy_magic_24_0.X VOUT- 3.89657f
C35 two_stage_opamp_dummy_magic_24_0.Vb3 VDDA 9.376019f
C36 bgr_11_0.Vin+ bgr_11_0.1st_Vout_1 0.275724f
C37 two_stage_opamp_dummy_magic_24_0.Vb3 two_stage_opamp_dummy_magic_24_0.V_err_gate 0.150414f
C38 bgr_11_0.START_UP_NFET1 VDDA 0.18791f
C39 bgr_11_0.Vin+ bgr_11_0.V_CUR_REF_REG 1.57077f
C40 two_stage_opamp_dummy_magic_24_0.X two_stage_opamp_dummy_magic_24_0.VD1 4.16017f
C41 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.VD1 0.015748f
C42 two_stage_opamp_dummy_magic_24_0.VD1 VIN- 0.533278f
C43 two_stage_opamp_dummy_magic_24_0.Vb3 two_stage_opamp_dummy_magic_24_0.cap_res_X 0.142f
C44 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.VD2 0.016362f
C45 two_stage_opamp_dummy_magic_24_0.V_tail_gate VIN+ 0.061031f
C46 two_stage_opamp_dummy_magic_24_0.Y two_stage_opamp_dummy_magic_24_0.VD2 4.16017f
C47 two_stage_opamp_dummy_magic_24_0.Vb3 VOUT+ 0.041713f
C48 VIN+ VIN- 0.075694f
C49 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_24_0.V_err_amp_ref 0.808133f
C50 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref two_stage_opamp_dummy_magic_24_0.Vb3 2.49744f
C51 bgr_11_0.V_CUR_REF_REG two_stage_opamp_dummy_magic_24_0.Vb1 0.051702f
C52 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.cap_res_Y 2.08159f
C53 bgr_11_0.START_UP_NFET1 bgr_11_0.START_UP 0.145663f
C54 two_stage_opamp_dummy_magic_24_0.Y two_stage_opamp_dummy_magic_24_0.cap_res_Y 0.056362f
C55 bgr_11_0.Vin+ bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 1.06291f
C56 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.X 0.030556f
C57 two_stage_opamp_dummy_magic_24_0.V_tail_gate VIN- 0.05849f
C58 two_stage_opamp_dummy_magic_24_0.Vb3 VOUT- 0.052551f
C59 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.V_CUR_REF_REG 0.779503f
C60 two_stage_opamp_dummy_magic_24_0.Y two_stage_opamp_dummy_magic_24_0.X 0.148787f
C61 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.Y 0.030556f
C62 two_stage_opamp_dummy_magic_24_0.Vb1 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage 0.141498f
C63 bgr_11_0.V_TOP two_stage_opamp_dummy_magic_24_0.V_tail_gate 0.028061f
C64 bgr_11_0.Vin+ VDDA 1.72765f
C65 bgr_11_0.1st_Vout_1 VDDA 2.67125f
C66 bgr_11_0.Vin+ two_stage_opamp_dummy_magic_24_0.V_err_gate 0.066808f
C67 two_stage_opamp_dummy_magic_24_0.V_err_gate bgr_11_0.1st_Vout_1 0.134861f
C68 bgr_11_0.V_CUR_REF_REG VDDA 3.77153f
C69 two_stage_opamp_dummy_magic_24_0.Vb3 a_4440_7230# 0.012f
C70 two_stage_opamp_dummy_magic_24_0.Vb3 two_stage_opamp_dummy_magic_24_0.cap_res_Y 0.033021f
C71 two_stage_opamp_dummy_magic_24_0.V_err_mir_p VDDA 0.684276f
C72 bgr_11_0.V_CUR_REF_REG two_stage_opamp_dummy_magic_24_0.V_err_gate 0.375039f
C73 a_5760_7230# VDDA 0.09634f
C74 two_stage_opamp_dummy_magic_24_0.V_err_gate two_stage_opamp_dummy_magic_24_0.V_err_mir_p 0.429395f
C75 two_stage_opamp_dummy_magic_24_0.Vb1 VDDA 11.858f
C76 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_24_0.V_tail_gate 0.582654f
C77 bgr_11_0.Vin+ bgr_11_0.START_UP 0.170134f
C78 bgr_11_0.START_UP bgr_11_0.1st_Vout_1 0.13011f
C79 two_stage_opamp_dummy_magic_24_0.Vb3 two_stage_opamp_dummy_magic_24_0.X 0.561365f
C80 two_stage_opamp_dummy_magic_24_0.Vb3 two_stage_opamp_dummy_magic_24_0.V_tail_gate 1.24656f
C81 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref bgr_11_0.Vin+ 0.25235f
C82 two_stage_opamp_dummy_magic_24_0.Vb3 two_stage_opamp_dummy_magic_24_0.Y 0.547856f
C83 two_stage_opamp_dummy_magic_24_0.Vb1 two_stage_opamp_dummy_magic_24_0.cap_res_X 0.05001f
C84 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter VDDA 0.023423f
C85 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage VDDA 0.013713f
C86 bgr_11_0.PFET_GATE_10uA bgr_11_0.V_TOP 0.198568f
C87 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref bgr_11_0.V_CUR_REF_REG 2.48242f
C88 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref two_stage_opamp_dummy_magic_24_0.V_err_mir_p 0.047104f
C89 two_stage_opamp_dummy_magic_24_0.Vb1 VOUT+ 0.110554f
C90 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref two_stage_opamp_dummy_magic_24_0.Vb1 3.27173f
C91 two_stage_opamp_dummy_magic_24_0.cap_res_X two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage 0.04898f
C92 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage VOUT+ 4.76385f
C93 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_24_0.Vb3 2.32805f
C94 two_stage_opamp_dummy_magic_24_0.V_err_gate VDDA 3.06287f
C95 two_stage_opamp_dummy_magic_24_0.Vb1 two_stage_opamp_dummy_magic_24_0.VD1 0.556058f
C96 bgr_11_0.PFET_GATE_10uA bgr_11_0.START_UP_NFET1 0.010791f
C97 two_stage_opamp_dummy_magic_24_0.cap_res_X VDDA 7.8698f
C98 two_stage_opamp_dummy_magic_24_0.Vb1 two_stage_opamp_dummy_magic_24_0.VD2 0.558539f
C99 two_stage_opamp_dummy_magic_24_0.V_err_gate two_stage_opamp_dummy_magic_24_0.cap_res_X 0.183227f
C100 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage VOUT- 4.73805f
C101 bgr_11_0.START_UP VDDA 2.28936f
C102 two_stage_opamp_dummy_magic_24_0.Vb1 VIN+ 0.016303f
C103 bgr_11_0.Vin+ two_stage_opamp_dummy_magic_24_0.V_tail_gate 0.014649f
C104 VDDA VOUT+ 15.3097f
C105 two_stage_opamp_dummy_magic_24_0.V_err_gate bgr_11_0.START_UP 0.743841f
C106 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref VDDA 6.679029f
C107 two_stage_opamp_dummy_magic_24_0.Vb1 two_stage_opamp_dummy_magic_24_0.cap_res_Y 0.218019f
C108 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref two_stage_opamp_dummy_magic_24_0.V_err_gate 0.742005f
C109 bgr_11_0.V_CUR_REF_REG two_stage_opamp_dummy_magic_24_0.V_tail_gate 0.403953f
C110 two_stage_opamp_dummy_magic_24_0.cap_res_X VOUT+ 0.011897f
C111 bgr_11_0.Vin+ bgr_11_0.V_TOP 1.8967f
C112 bgr_11_0.V_TOP bgr_11_0.1st_Vout_1 2.6266f
C113 two_stage_opamp_dummy_magic_24_0.Vb1 two_stage_opamp_dummy_magic_24_0.V_tail_gate 0.630007f
C114 two_stage_opamp_dummy_magic_24_0.Vb1 two_stage_opamp_dummy_magic_24_0.X 1.58533f
C115 two_stage_opamp_dummy_magic_24_0.Vb1 VIN- 0.011528f
C116 VDDA VOUT- 15.3172f
C117 two_stage_opamp_dummy_magic_24_0.Vb1 two_stage_opamp_dummy_magic_24_0.Y 1.94718f
C118 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref bgr_11_0.START_UP 1.39993f
C119 two_stage_opamp_dummy_magic_24_0.V_err_gate VOUT- 0.020883f
C120 bgr_11_0.V_CUR_REF_REG bgr_11_0.V_TOP 0.308375f
C121 two_stage_opamp_dummy_magic_24_0.cap_res_Y two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage 0.04898f
C122 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref VOUT+ 0.020461f
C123 two_stage_opamp_dummy_magic_24_0.cap_res_X VOUT- 50.9233f
C124 two_stage_opamp_dummy_magic_24_0.V_tail_gate two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage 3.23133f
C125 VIN- GNDA 1.84317f
C126 VIN+ GNDA 1.84009f
C127 VOUT- GNDA 25.807001f
C128 VOUT+ GNDA 25.770336f
C129 VDDA GNDA 0.375312p
C130 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage GNDA 9.68961f
C131 two_stage_opamp_dummy_magic_24_0.VD1 GNDA 2.8949f
C132 two_stage_opamp_dummy_magic_24_0.VD2 GNDA 2.89089f
C133 two_stage_opamp_dummy_magic_24_0.cap_res_X GNDA 41.580433f
C134 two_stage_opamp_dummy_magic_24_0.V_err_mir_p GNDA 0.103495f
C135 two_stage_opamp_dummy_magic_24_0.cap_res_Y GNDA 41.53443f
C136 two_stage_opamp_dummy_magic_24_0.X GNDA 12.416237f
C137 two_stage_opamp_dummy_magic_24_0.Y GNDA 12.095636f
C138 a_5760_7230# GNDA 0.045515f
C139 a_4440_7230# GNDA 0.046297f
C140 two_stage_opamp_dummy_magic_24_0.V_tail_gate GNDA 40.157658f
C141 two_stage_opamp_dummy_magic_24_0.Vb1 GNDA 15.314911f
C142 bgr_11_0.1st_Vout_1 GNDA 11.637372f
C143 bgr_11_0.START_UP GNDA 6.621171f
C144 bgr_11_0.START_UP_NFET1 GNDA 5.23563f
C145 two_stage_opamp_dummy_magic_24_0.V_err_gate GNDA 12.054708f
C146 two_stage_opamp_dummy_magic_24_0.Vb3 GNDA 15.874961f
C147 bgr_11_0.V_TOP GNDA 10.653124f
C148 bgr_11_0.V_CUR_REF_REG GNDA 4.877919f
C149 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA 16.830502f
C150 bgr_11_0.Vin+ GNDA 4.647377f
C151 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref GNDA 11.94606f
C152 bgr_11_0.PFET_GATE_10uA GNDA 8.898536f
C153 bgr_11_0.V_CUR_REF_REG.t3 GNDA 0.066747f
C154 bgr_11_0.V_CUR_REF_REG.t0 GNDA 0.452298f
C155 bgr_11_0.V_CUR_REF_REG.t1 GNDA 0.013056f
C156 bgr_11_0.V_CUR_REF_REG.t2 GNDA 0.013056f
C157 bgr_11_0.V_CUR_REF_REG.n0 GNDA 0.100023f
C158 bgr_11_0.V_CUR_REF_REG.n1 GNDA 5.13907f
C159 two_stage_opamp_dummy_magic_24_0.err_amp_out.t2 GNDA 0.035995f
C160 two_stage_opamp_dummy_magic_24_0.err_amp_out.t4 GNDA 0.085538f
C161 two_stage_opamp_dummy_magic_24_0.err_amp_out.t3 GNDA 0.035995f
C162 two_stage_opamp_dummy_magic_24_0.err_amp_out.t0 GNDA 0.035995f
C163 two_stage_opamp_dummy_magic_24_0.err_amp_out.n0 GNDA 0.112847f
C164 two_stage_opamp_dummy_magic_24_0.err_amp_out.n1 GNDA 1.73725f
C165 two_stage_opamp_dummy_magic_24_0.err_amp_out.n2 GNDA 0.120386f
C166 two_stage_opamp_dummy_magic_24_0.err_amp_out.t1 GNDA 0.035995f
C167 bgr_11_0.Vin-.n0 GNDA 0.07858f
C168 bgr_11_0.Vin-.n1 GNDA 0.088293f
C169 bgr_11_0.Vin-.n2 GNDA 0.12735f
C170 bgr_11_0.Vin-.t4 GNDA 0.294736f
C171 bgr_11_0.Vin-.t3 GNDA 0.030534f
C172 bgr_11_0.Vin-.t0 GNDA 0.030534f
C173 bgr_11_0.Vin-.n3 GNDA 0.085799f
C174 bgr_11_0.Vin-.t1 GNDA 0.030534f
C175 bgr_11_0.Vin-.t2 GNDA 0.030534f
C176 bgr_11_0.Vin-.n4 GNDA 0.074088f
C177 bgr_11_0.Vin-.n5 GNDA 0.633984f
C178 bgr_11_0.Vin-.t6 GNDA 0.010178f
C179 bgr_11_0.Vin-.t5 GNDA 0.010178f
C180 bgr_11_0.Vin-.n6 GNDA 0.031534f
C181 bgr_11_0.Vin-.n7 GNDA 0.428495f
C182 bgr_11_0.Vin-.t8 GNDA 0.049457f
C183 bgr_11_0.Vin-.n8 GNDA 0.623119f
C184 bgr_11_0.Vin-.t7 GNDA 0.128901f
C185 bgr_11_0.Vin-.n9 GNDA 0.734405f
C186 bgr_11_0.Vin-.n10 GNDA 1.36082f
C187 bgr_11_0.Vin-.n11 GNDA 0.531118f
C188 bgr_11_0.Vin-.n12 GNDA 0.079463f
C189 bgr_11_0.Vin-.n13 GNDA 0.13464f
C190 bgr_11_0.Vin-.n14 GNDA 0.078726f
C191 bgr_11_0.Vin-.n15 GNDA 0.155721f
C192 bgr_11_0.Vin-.n16 GNDA 0.155721f
C193 bgr_11_0.Vin-.n17 GNDA -0.303656f
C194 bgr_11_0.Vin-.n18 GNDA 0.501878f
C195 bgr_11_0.Vin-.n19 GNDA 0.240599f
C196 bgr_11_0.Vin-.n20 GNDA 0.454563f
C197 bgr_11_0.Vin-.n21 GNDA 0.043263f
C198 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter GNDA 0.045912f
C199 bgr_11_0.START_UP.t4 GNDA 1.72724f
C200 bgr_11_0.START_UP.t5 GNDA 0.045404f
C201 bgr_11_0.START_UP.n0 GNDA 1.15615f
C202 bgr_11_0.START_UP.t0 GNDA 0.04333f
C203 bgr_11_0.START_UP.t2 GNDA 0.04333f
C204 bgr_11_0.START_UP.n1 GNDA 0.135247f
C205 bgr_11_0.START_UP.t1 GNDA 0.04333f
C206 bgr_11_0.START_UP.t3 GNDA 0.04333f
C207 bgr_11_0.START_UP.n2 GNDA 0.106737f
C208 bgr_11_0.START_UP.n3 GNDA 1.0283f
C209 bgr_11_0.START_UP.t6 GNDA 0.016282f
C210 bgr_11_0.START_UP.t7 GNDA 0.016282f
C211 bgr_11_0.START_UP.n4 GNDA 0.046713f
C212 bgr_11_0.START_UP.n5 GNDA 0.477587f
C213 bgr_11_0.cap_res2.t4 GNDA 0.334798f
C214 bgr_11_0.cap_res2.t10 GNDA 0.336011f
C215 bgr_11_0.cap_res2.t20 GNDA 0.318043f
C216 bgr_11_0.cap_res2.t9 GNDA 0.334798f
C217 bgr_11_0.cap_res2.t14 GNDA 0.336011f
C218 bgr_11_0.cap_res2.t5 GNDA 0.318043f
C219 bgr_11_0.cap_res2.t3 GNDA 0.334798f
C220 bgr_11_0.cap_res2.t8 GNDA 0.336011f
C221 bgr_11_0.cap_res2.t18 GNDA 0.318043f
C222 bgr_11_0.cap_res2.t16 GNDA 0.334798f
C223 bgr_11_0.cap_res2.t2 GNDA 0.336011f
C224 bgr_11_0.cap_res2.t12 GNDA 0.318043f
C225 bgr_11_0.cap_res2.t1 GNDA 0.334798f
C226 bgr_11_0.cap_res2.t6 GNDA 0.336011f
C227 bgr_11_0.cap_res2.t17 GNDA 0.318043f
C228 bgr_11_0.cap_res2.n0 GNDA 0.224415f
C229 bgr_11_0.cap_res2.t11 GNDA 0.178714f
C230 bgr_11_0.cap_res2.n1 GNDA 0.243496f
C231 bgr_11_0.cap_res2.t7 GNDA 0.178714f
C232 bgr_11_0.cap_res2.n2 GNDA 0.243496f
C233 bgr_11_0.cap_res2.t13 GNDA 0.178714f
C234 bgr_11_0.cap_res2.n3 GNDA 0.243496f
C235 bgr_11_0.cap_res2.t19 GNDA 0.178714f
C236 bgr_11_0.cap_res2.n4 GNDA 0.243496f
C237 bgr_11_0.cap_res2.t15 GNDA 0.360089f
C238 bgr_11_0.cap_res2.t0 GNDA 0.082395f
C239 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t0 GNDA 0.204065f
C240 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t8 GNDA 0.64181f
C241 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t4 GNDA 0.641633f
C242 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n0 GNDA 0.528383f
C243 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t9 GNDA 0.641633f
C244 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n1 GNDA 0.275151f
C245 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t7 GNDA 0.641633f
C246 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n2 GNDA 0.554173f
C247 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n3 GNDA 0.656492f
C248 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t1 GNDA 0.204065f
C249 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n4 GNDA 0.358405f
C250 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t6 GNDA 0.554419f
C251 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t3 GNDA 0.554419f
C252 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t2 GNDA 0.554419f
C253 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.t5 GNDA 0.599502f
C254 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n5 GNDA 0.200699f
C255 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n6 GNDA 0.249608f
C256 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n7 GNDA 0.249608f
C257 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n8 GNDA 0.244173f
C258 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n9 GNDA 0.406273f
C259 two_stage_opamp_dummy_magic_24_0.V_b_2nd_stage.n10 GNDA 1.16109f
C260 two_stage_opamp_dummy_magic_24_0.VD1.t3 GNDA 0.044096f
C261 two_stage_opamp_dummy_magic_24_0.VD1.t10 GNDA 0.044096f
C262 two_stage_opamp_dummy_magic_24_0.VD1.n0 GNDA 0.097626f
C263 two_stage_opamp_dummy_magic_24_0.VD1.n1 GNDA 0.458534f
C264 two_stage_opamp_dummy_magic_24_0.VD1.n2 GNDA 0.066168f
C265 two_stage_opamp_dummy_magic_24_0.VD1.n3 GNDA 0.109634f
C266 two_stage_opamp_dummy_magic_24_0.VD1.t15 GNDA 0.044096f
C267 two_stage_opamp_dummy_magic_24_0.VD1.t19 GNDA 0.044096f
C268 two_stage_opamp_dummy_magic_24_0.VD1.n4 GNDA 0.095949f
C269 two_stage_opamp_dummy_magic_24_0.VD1.n5 GNDA 0.369685f
C270 two_stage_opamp_dummy_magic_24_0.VD1.n6 GNDA 0.09378f
C271 two_stage_opamp_dummy_magic_24_0.VD1.t13 GNDA 0.044096f
C272 two_stage_opamp_dummy_magic_24_0.VD1.t0 GNDA 0.044096f
C273 two_stage_opamp_dummy_magic_24_0.VD1.n7 GNDA 0.095949f
C274 two_stage_opamp_dummy_magic_24_0.VD1.n8 GNDA 0.379992f
C275 two_stage_opamp_dummy_magic_24_0.VD1.t2 GNDA 0.044096f
C276 two_stage_opamp_dummy_magic_24_0.VD1.t7 GNDA 0.044096f
C277 two_stage_opamp_dummy_magic_24_0.VD1.n9 GNDA 0.097626f
C278 two_stage_opamp_dummy_magic_24_0.VD1.t6 GNDA 0.044096f
C279 two_stage_opamp_dummy_magic_24_0.VD1.t11 GNDA 0.044096f
C280 two_stage_opamp_dummy_magic_24_0.VD1.n10 GNDA 0.097626f
C281 two_stage_opamp_dummy_magic_24_0.VD1.n11 GNDA 0.625445f
C282 two_stage_opamp_dummy_magic_24_0.VD1.t5 GNDA 0.044096f
C283 two_stage_opamp_dummy_magic_24_0.VD1.t9 GNDA 0.044096f
C284 two_stage_opamp_dummy_magic_24_0.VD1.n12 GNDA 0.097626f
C285 two_stage_opamp_dummy_magic_24_0.VD1.n13 GNDA 0.168952f
C286 two_stage_opamp_dummy_magic_24_0.VD1.t1 GNDA 0.044096f
C287 two_stage_opamp_dummy_magic_24_0.VD1.t12 GNDA 0.044096f
C288 two_stage_opamp_dummy_magic_24_0.VD1.n14 GNDA 0.095949f
C289 two_stage_opamp_dummy_magic_24_0.VD1.n15 GNDA 0.379992f
C290 two_stage_opamp_dummy_magic_24_0.VD1.n16 GNDA 0.15941f
C291 two_stage_opamp_dummy_magic_24_0.VD1.t17 GNDA 0.044096f
C292 two_stage_opamp_dummy_magic_24_0.VD1.t21 GNDA 0.044096f
C293 two_stage_opamp_dummy_magic_24_0.VD1.n17 GNDA 0.095949f
C294 two_stage_opamp_dummy_magic_24_0.VD1.n18 GNDA 0.369685f
C295 two_stage_opamp_dummy_magic_24_0.VD1.n19 GNDA 0.066168f
C296 two_stage_opamp_dummy_magic_24_0.VD1.n20 GNDA 0.109634f
C297 two_stage_opamp_dummy_magic_24_0.VD1.n21 GNDA 0.617932f
C298 two_stage_opamp_dummy_magic_24_0.VD1.n22 GNDA 0.148295f
C299 two_stage_opamp_dummy_magic_24_0.VD1.n23 GNDA 0.088193f
C300 two_stage_opamp_dummy_magic_24_0.VD1.t4 GNDA 0.044096f
C301 two_stage_opamp_dummy_magic_24_0.VD1.t8 GNDA 0.044096f
C302 two_stage_opamp_dummy_magic_24_0.VD1.n24 GNDA 0.097626f
C303 two_stage_opamp_dummy_magic_24_0.VD1.n25 GNDA 0.617932f
C304 two_stage_opamp_dummy_magic_24_0.VD1.n26 GNDA 0.148295f
C305 two_stage_opamp_dummy_magic_24_0.VD1.n27 GNDA 0.625445f
C306 two_stage_opamp_dummy_magic_24_0.VD1.n28 GNDA 0.168952f
C307 two_stage_opamp_dummy_magic_24_0.VD1.n29 GNDA 0.066168f
C308 two_stage_opamp_dummy_magic_24_0.VD1.t14 GNDA 0.044096f
C309 two_stage_opamp_dummy_magic_24_0.VD1.t18 GNDA 0.044096f
C310 two_stage_opamp_dummy_magic_24_0.VD1.n30 GNDA 0.095949f
C311 two_stage_opamp_dummy_magic_24_0.VD1.n31 GNDA 0.369685f
C312 two_stage_opamp_dummy_magic_24_0.VD1.n32 GNDA 0.15941f
C313 two_stage_opamp_dummy_magic_24_0.VD1.n33 GNDA 0.09378f
C314 two_stage_opamp_dummy_magic_24_0.VD1.t16 GNDA 0.044096f
C315 two_stage_opamp_dummy_magic_24_0.VD1.t20 GNDA 0.044096f
C316 two_stage_opamp_dummy_magic_24_0.VD1.n34 GNDA 0.095949f
C317 two_stage_opamp_dummy_magic_24_0.VD1.n35 GNDA 0.369685f
C318 two_stage_opamp_dummy_magic_24_0.VD1.n36 GNDA 0.066168f
C319 two_stage_opamp_dummy_magic_24_0.VD1.n37 GNDA 0.051213f
C320 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t14 GNDA 0.029249f
C321 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t11 GNDA 0.029249f
C322 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n0 GNDA 0.091984f
C323 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t12 GNDA 0.029249f
C324 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t13 GNDA 0.029249f
C325 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n1 GNDA 0.062742f
C326 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n2 GNDA 2.77401f
C327 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t10 GNDA 0.358459f
C328 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n3 GNDA 0.101738f
C329 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n4 GNDA 0.175052f
C330 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t9 GNDA 0.087748f
C331 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t4 GNDA 0.087748f
C332 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n5 GNDA 0.187676f
C333 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n6 GNDA 0.587049f
C334 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t0 GNDA 0.087748f
C335 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t5 GNDA 0.087748f
C336 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n7 GNDA 0.187676f
C337 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n8 GNDA 0.571149f
C338 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n9 GNDA 0.175052f
C339 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n10 GNDA 0.101738f
C340 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t2 GNDA 0.087748f
C341 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t6 GNDA 0.087748f
C342 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n11 GNDA 0.187676f
C343 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n12 GNDA 0.571149f
C344 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n13 GNDA 0.101738f
C345 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t1 GNDA 0.087748f
C346 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t8 GNDA 0.087748f
C347 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n14 GNDA 0.187676f
C348 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n15 GNDA 0.571149f
C349 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n16 GNDA 0.175052f
C350 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t3 GNDA 0.087748f
C351 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.t7 GNDA 0.087748f
C352 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n17 GNDA 0.187676f
C353 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n18 GNDA 0.579099f
C354 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n19 GNDA 0.202941f
C355 two_stage_opamp_dummy_magic_24_0.V_CMFB_S2.n20 GNDA 3.08039f
C356 bgr_11_0.V_CMFB_S2 GNDA 5.78665f
C357 bgr_11_0.Vin+.t5 GNDA 0.221779f
C358 bgr_11_0.Vin+.t4 GNDA 0.096124f
C359 bgr_11_0.Vin+.n0 GNDA 1.46352f
C360 bgr_11_0.Vin+.t0 GNDA 0.033039f
C361 bgr_11_0.Vin+.t3 GNDA 0.033039f
C362 bgr_11_0.Vin+.n1 GNDA 0.084276f
C363 bgr_11_0.Vin+.t2 GNDA 0.033039f
C364 bgr_11_0.Vin+.t1 GNDA 0.033039f
C365 bgr_11_0.Vin+.n2 GNDA 0.078979f
C366 bgr_11_0.Vin+.n3 GNDA 0.79622f
C367 bgr_11_0.Vin+.n4 GNDA 0.652102f
C368 bgr_11_0.Vin+.t6 GNDA 0.052809f
C369 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t11 GNDA 0.020236f
C370 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t16 GNDA 0.020236f
C371 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n0 GNDA 0.050725f
C372 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t14 GNDA 0.020236f
C373 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t13 GNDA 0.020236f
C374 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n1 GNDA 0.050457f
C375 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n2 GNDA 0.448463f
C376 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t15 GNDA 0.020236f
C377 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t12 GNDA 0.020236f
C378 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n3 GNDA 0.040472f
C379 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n4 GNDA 0.075881f
C380 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t10 GNDA 0.255502f
C381 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n5 GNDA 0.063925f
C382 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n6 GNDA 0.113072f
C383 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t8 GNDA 0.040472f
C384 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t3 GNDA 0.040472f
C385 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n7 GNDA 0.082749f
C386 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n8 GNDA 0.277952f
C387 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t9 GNDA 0.040472f
C388 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t4 GNDA 0.040472f
C389 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n9 GNDA 0.082749f
C390 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n10 GNDA 0.26767f
C391 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n11 GNDA 0.108691f
C392 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n12 GNDA 0.063925f
C393 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t1 GNDA 0.040472f
C394 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t5 GNDA 0.040472f
C395 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n13 GNDA 0.082749f
C396 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n14 GNDA 0.26767f
C397 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n15 GNDA 0.066263f
C398 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t0 GNDA 0.040472f
C399 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t7 GNDA 0.040472f
C400 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n16 GNDA 0.082749f
C401 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n17 GNDA 0.26767f
C402 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n18 GNDA 0.113072f
C403 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t2 GNDA 0.040472f
C404 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.t6 GNDA 0.040472f
C405 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n19 GNDA 0.082749f
C406 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n20 GNDA 0.272958f
C407 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n21 GNDA 0.14752f
C408 two_stage_opamp_dummy_magic_24_0.V_CMFB_S1.n22 GNDA 2.42805f
C409 bgr_11_0.V_CMFB_S1 GNDA 2.38018f
C410 two_stage_opamp_dummy_magic_24_0.V_tot.t3 GNDA 0.204389f
C411 two_stage_opamp_dummy_magic_24_0.V_tot.t2 GNDA 0.204389f
C412 two_stage_opamp_dummy_magic_24_0.V_tot.t1 GNDA 0.191871f
C413 two_stage_opamp_dummy_magic_24_0.V_tot.n0 GNDA 1.15943f
C414 two_stage_opamp_dummy_magic_24_0.V_tot.t5 GNDA 0.058137f
C415 two_stage_opamp_dummy_magic_24_0.V_tot.n1 GNDA 1.08618f
C416 two_stage_opamp_dummy_magic_24_0.V_tot.t4 GNDA 0.058137f
C417 two_stage_opamp_dummy_magic_24_0.V_tot.n2 GNDA 1.08618f
C418 two_stage_opamp_dummy_magic_24_0.V_tot.n3 GNDA 1.15943f
C419 two_stage_opamp_dummy_magic_24_0.V_tot.t0 GNDA 0.191871f
C420 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n0 GNDA 6.31386f
C421 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n1 GNDA 5.3586f
C422 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n2 GNDA 0.134403f
C423 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t29 GNDA 0.016295f
C424 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t12 GNDA 0.016295f
C425 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t24 GNDA 0.016295f
C426 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t14 GNDA 0.016295f
C427 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t26 GNDA 0.016295f
C428 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t19 GNDA 0.016295f
C429 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t30 GNDA 0.016295f
C430 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t21 GNDA 0.016295f
C431 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t16 GNDA 0.016295f
C432 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t28 GNDA 0.019019f
C433 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n3 GNDA 0.017932f
C434 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n4 GNDA 0.011246f
C435 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n5 GNDA 0.011246f
C436 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n6 GNDA 0.011246f
C437 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n7 GNDA 0.011246f
C438 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n8 GNDA 0.011246f
C439 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n9 GNDA 0.011246f
C440 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n10 GNDA 0.011246f
C441 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n11 GNDA 0.010524f
C442 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t31 GNDA 0.016295f
C443 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t20 GNDA 0.016295f
C444 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t27 GNDA 0.016295f
C445 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t15 GNDA 0.016295f
C446 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t25 GNDA 0.016295f
C447 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t13 GNDA 0.016295f
C448 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t23 GNDA 0.016295f
C449 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t18 GNDA 0.019019f
C450 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n13 GNDA 0.017932f
C451 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n14 GNDA 0.011246f
C452 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n15 GNDA 0.011246f
C453 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n16 GNDA 0.011246f
C454 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n17 GNDA 0.011246f
C455 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n18 GNDA 0.011246f
C456 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n19 GNDA 0.010524f
C457 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t22 GNDA 0.016295f
C458 two_stage_opamp_dummy_magic_24_0.V_tail_gate.t17 GNDA 0.016295f
C459 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n20 GNDA 0.010524f
C460 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n21 GNDA 0.010524f
C461 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n23 GNDA 0.01224f
C462 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n24 GNDA 0.01224f
C463 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n25 GNDA 0.01224f
C464 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n26 GNDA 0.134041f
C465 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n27 GNDA 0.070082f
C466 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n28 GNDA 0.01224f
C467 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n29 GNDA 0.022226f
C468 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n30 GNDA 0.070082f
C469 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n31 GNDA 0.134395f
C470 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n32 GNDA 0.021933f
C471 two_stage_opamp_dummy_magic_24_0.V_tail_gate.n33 GNDA 0.021933f
C472 two_stage_opamp_dummy_magic_24_0.V_err_gate.t2 GNDA 0.02046f
C473 two_stage_opamp_dummy_magic_24_0.V_err_gate.t3 GNDA 0.02046f
C474 two_stage_opamp_dummy_magic_24_0.V_err_gate.n0 GNDA 0.25059f
C475 two_stage_opamp_dummy_magic_24_0.V_err_gate.t0 GNDA 0.051151f
C476 two_stage_opamp_dummy_magic_24_0.V_err_gate.t5 GNDA 0.051151f
C477 two_stage_opamp_dummy_magic_24_0.V_err_gate.n1 GNDA 0.156712f
C478 two_stage_opamp_dummy_magic_24_0.V_err_gate.t6 GNDA 0.057118f
C479 two_stage_opamp_dummy_magic_24_0.V_err_gate.t8 GNDA 0.057118f
C480 two_stage_opamp_dummy_magic_24_0.V_err_gate.n2 GNDA 0.085796f
C481 two_stage_opamp_dummy_magic_24_0.V_err_gate.n3 GNDA 0.316651f
C482 two_stage_opamp_dummy_magic_24_0.V_err_gate.t4 GNDA 0.051151f
C483 two_stage_opamp_dummy_magic_24_0.V_err_gate.t1 GNDA 0.051151f
C484 two_stage_opamp_dummy_magic_24_0.V_err_gate.n4 GNDA 0.156033f
C485 two_stage_opamp_dummy_magic_24_0.V_err_gate.n5 GNDA 0.242282f
C486 two_stage_opamp_dummy_magic_24_0.V_err_gate.t9 GNDA 0.057118f
C487 two_stage_opamp_dummy_magic_24_0.V_err_gate.t7 GNDA 0.057118f
C488 two_stage_opamp_dummy_magic_24_0.V_err_gate.n6 GNDA 0.085796f
C489 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t2 GNDA 0.027485f
C490 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t0 GNDA 0.027485f
C491 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n0 GNDA 0.086437f
C492 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t1 GNDA 0.027485f
C493 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t4 GNDA 0.027485f
C494 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n1 GNDA 0.058958f
C495 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n2 GNDA 1.83575f
C496 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t3 GNDA 0.33684f
C497 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n3 GNDA 0.095602f
C498 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n4 GNDA 0.164494f
C499 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t8 GNDA 0.082456f
C500 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t11 GNDA 0.082456f
C501 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n5 GNDA 0.176357f
C502 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n6 GNDA 0.551643f
C503 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t5 GNDA 0.082456f
C504 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t10 GNDA 0.082456f
C505 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n7 GNDA 0.176357f
C506 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n8 GNDA 0.536702f
C507 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n9 GNDA 0.164494f
C508 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n10 GNDA 0.095602f
C509 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t14 GNDA 0.082456f
C510 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t9 GNDA 0.082456f
C511 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n11 GNDA 0.176357f
C512 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n12 GNDA 0.536702f
C513 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n13 GNDA 0.095602f
C514 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t7 GNDA 0.082456f
C515 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t13 GNDA 0.082456f
C516 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n14 GNDA 0.176357f
C517 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n15 GNDA 0.536702f
C518 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n16 GNDA 0.164494f
C519 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t6 GNDA 0.082456f
C520 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.t12 GNDA 0.082456f
C521 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n17 GNDA 0.176357f
C522 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n18 GNDA 0.544172f
C523 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n19 GNDA 0.190701f
C524 two_stage_opamp_dummy_magic_24_0.V_CMFB_S4.n20 GNDA 2.95799f
C525 bgr_11_0.V_CMFB_S4 GNDA 4.43084f
C526 bgr_11_0.cap_res1.t5 GNDA 0.339883f
C527 bgr_11_0.cap_res1.t17 GNDA 0.357788f
C528 bgr_11_0.cap_res1.t9 GNDA 0.359085f
C529 bgr_11_0.cap_res1.t12 GNDA 0.339883f
C530 bgr_11_0.cap_res1.t19 GNDA 0.357788f
C531 bgr_11_0.cap_res1.t16 GNDA 0.359085f
C532 bgr_11_0.cap_res1.t4 GNDA 0.339883f
C533 bgr_11_0.cap_res1.t15 GNDA 0.357788f
C534 bgr_11_0.cap_res1.t8 GNDA 0.359085f
C535 bgr_11_0.cap_res1.t0 GNDA 0.339883f
C536 bgr_11_0.cap_res1.t7 GNDA 0.357788f
C537 bgr_11_0.cap_res1.t1 GNDA 0.359085f
C538 bgr_11_0.cap_res1.t2 GNDA 0.339883f
C539 bgr_11_0.cap_res1.t14 GNDA 0.357788f
C540 bgr_11_0.cap_res1.t6 GNDA 0.359085f
C541 bgr_11_0.cap_res1.n0 GNDA 0.239826f
C542 bgr_11_0.cap_res1.t10 GNDA 0.190986f
C543 bgr_11_0.cap_res1.n1 GNDA 0.260216f
C544 bgr_11_0.cap_res1.t3 GNDA 0.190986f
C545 bgr_11_0.cap_res1.n2 GNDA 0.260216f
C546 bgr_11_0.cap_res1.t11 GNDA 0.190986f
C547 bgr_11_0.cap_res1.n3 GNDA 0.260216f
C548 bgr_11_0.cap_res1.t18 GNDA 0.190986f
C549 bgr_11_0.cap_res1.n4 GNDA 0.260216f
C550 bgr_11_0.cap_res1.t13 GNDA 0.383393f
C551 bgr_11_0.cap_res1.t20 GNDA 0.088196f
C552 bgr_11_0.1st_Vout_1.n0 GNDA 0.191219f
C553 bgr_11_0.1st_Vout_1.t27 GNDA 0.240974f
C554 bgr_11_0.1st_Vout_1.t18 GNDA 0.236938f
C555 bgr_11_0.1st_Vout_1.t14 GNDA 0.240974f
C556 bgr_11_0.1st_Vout_1.t23 GNDA 0.236938f
C557 bgr_11_0.1st_Vout_1.n1 GNDA 0.158859f
C558 bgr_11_0.1st_Vout_1.n2 GNDA 0.203285f
C559 bgr_11_0.1st_Vout_1.t32 GNDA 0.240974f
C560 bgr_11_0.1st_Vout_1.t26 GNDA 0.236938f
C561 bgr_11_0.1st_Vout_1.t22 GNDA 0.240974f
C562 bgr_11_0.1st_Vout_1.t31 GNDA 0.236938f
C563 bgr_11_0.1st_Vout_1.n3 GNDA 0.158859f
C564 bgr_11_0.1st_Vout_1.n4 GNDA 0.247711f
C565 bgr_11_0.1st_Vout_1.t25 GNDA 0.240974f
C566 bgr_11_0.1st_Vout_1.t17 GNDA 0.236938f
C567 bgr_11_0.1st_Vout_1.t12 GNDA 0.240974f
C568 bgr_11_0.1st_Vout_1.t21 GNDA 0.236938f
C569 bgr_11_0.1st_Vout_1.n5 GNDA 0.158859f
C570 bgr_11_0.1st_Vout_1.n6 GNDA 0.247711f
C571 bgr_11_0.1st_Vout_1.t16 GNDA 0.240974f
C572 bgr_11_0.1st_Vout_1.t8 GNDA 0.236938f
C573 bgr_11_0.1st_Vout_1.t7 GNDA 0.240974f
C574 bgr_11_0.1st_Vout_1.t11 GNDA 0.236938f
C575 bgr_11_0.1st_Vout_1.n7 GNDA 0.158859f
C576 bgr_11_0.1st_Vout_1.n8 GNDA 0.247711f
C577 bgr_11_0.1st_Vout_1.t24 GNDA 0.240974f
C578 bgr_11_0.1st_Vout_1.t15 GNDA 0.236938f
C579 bgr_11_0.1st_Vout_1.n9 GNDA 0.203285f
C580 bgr_11_0.1st_Vout_1.t20 GNDA 0.236938f
C581 bgr_11_0.1st_Vout_1.n10 GNDA 0.10366f
C582 bgr_11_0.1st_Vout_1.t9 GNDA 0.236938f
C583 bgr_11_0.1st_Vout_1.n11 GNDA 2.00975f
C584 bgr_11_0.1st_Vout_1.t29 GNDA 0.01424f
C585 bgr_11_0.1st_Vout_1.n12 GNDA 3.07165f
C586 bgr_11_0.1st_Vout_1.n13 GNDA 0.012548f
C587 bgr_11_0.1st_Vout_1.n14 GNDA 0.191219f
C588 bgr_11_0.1st_Vout_1.n15 GNDA 0.017467f
C589 bgr_11_0.1st_Vout_1.n16 GNDA 0.173289f
C590 bgr_11_0.1st_Vout_1.n17 GNDA 0.012189f
C591 bgr_11_0.1st_Vout_1.t2 GNDA 0.054022f
C592 bgr_11_0.1st_Vout_1.n18 GNDA 0.173688f
C593 bgr_11_0.1st_Vout_1.n19 GNDA 0.127946f
C594 bgr_11_0.1st_Vout_1.n20 GNDA 0.017467f
C595 bgr_11_0.1st_Vout_1.n21 GNDA 0.173289f
C596 bgr_11_0.1st_Vout_1.n22 GNDA 0.012548f
C597 bgr_11_0.1st_Vout_1.t13 GNDA 0.013988f
C598 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t4 GNDA 0.36259f
C599 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t9 GNDA 0.11469f
C600 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n0 GNDA 3.72935f
C601 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t5 GNDA 0.068611f
C602 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t1 GNDA 0.068611f
C603 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n1 GNDA 0.191389f
C604 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t3 GNDA 0.068611f
C605 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t0 GNDA 0.068611f
C606 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n2 GNDA 0.172263f
C607 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n3 GNDA 2.11548f
C608 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t2 GNDA 0.068611f
C609 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t6 GNDA 0.068611f
C610 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n4 GNDA 0.172263f
C611 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n5 GNDA 1.57287f
C612 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n6 GNDA 1.00387f
C613 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t7 GNDA 0.078854f
C614 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.t8 GNDA 0.077505f
C615 two_stage_opamp_dummy_magic_24_0.V_err_amp_ref.n7 GNDA 0.570406f
C616 bgr_11_0.V_TOP.n0 GNDA 0.016831f
C617 bgr_11_0.V_TOP.t29 GNDA 0.128711f
C618 bgr_11_0.V_TOP.t37 GNDA 0.128973f
C619 bgr_11_0.V_TOP.t38 GNDA 0.129529f
C620 bgr_11_0.V_TOP.n1 GNDA 0.162971f
C621 bgr_11_0.V_TOP.t23 GNDA 0.129529f
C622 bgr_11_0.V_TOP.n2 GNDA 0.089272f
C623 bgr_11_0.V_TOP.t48 GNDA 0.129529f
C624 bgr_11_0.V_TOP.n3 GNDA 0.089272f
C625 bgr_11_0.V_TOP.t39 GNDA 0.129529f
C626 bgr_11_0.V_TOP.n4 GNDA 0.089272f
C627 bgr_11_0.V_TOP.t27 GNDA 0.129529f
C628 bgr_11_0.V_TOP.n5 GNDA 0.089272f
C629 bgr_11_0.V_TOP.n6 GNDA 0.025246f
C630 bgr_11_0.V_TOP.n7 GNDA 0.057364f
C631 bgr_11_0.V_TOP.t9 GNDA 0.129887f
C632 bgr_11_0.V_TOP.t20 GNDA 0.374019f
C633 bgr_11_0.V_TOP.t24 GNDA 0.38039f
C634 bgr_11_0.V_TOP.t32 GNDA 0.374019f
C635 bgr_11_0.V_TOP.n8 GNDA 0.250768f
C636 bgr_11_0.V_TOP.t19 GNDA 0.374019f
C637 bgr_11_0.V_TOP.t46 GNDA 0.38039f
C638 bgr_11_0.V_TOP.n9 GNDA 0.320897f
C639 bgr_11_0.V_TOP.t34 GNDA 0.38039f
C640 bgr_11_0.V_TOP.t40 GNDA 0.374019f
C641 bgr_11_0.V_TOP.n10 GNDA 0.250768f
C642 bgr_11_0.V_TOP.t31 GNDA 0.374019f
C643 bgr_11_0.V_TOP.t18 GNDA 0.38039f
C644 bgr_11_0.V_TOP.n11 GNDA 0.391025f
C645 bgr_11_0.V_TOP.t22 GNDA 0.38039f
C646 bgr_11_0.V_TOP.t30 GNDA 0.374019f
C647 bgr_11_0.V_TOP.n12 GNDA 0.250768f
C648 bgr_11_0.V_TOP.t17 GNDA 0.374019f
C649 bgr_11_0.V_TOP.t44 GNDA 0.38039f
C650 bgr_11_0.V_TOP.n13 GNDA 0.391025f
C651 bgr_11_0.V_TOP.t47 GNDA 0.38039f
C652 bgr_11_0.V_TOP.t16 GNDA 0.374019f
C653 bgr_11_0.V_TOP.n14 GNDA 0.250768f
C654 bgr_11_0.V_TOP.t43 GNDA 0.374019f
C655 bgr_11_0.V_TOP.t35 GNDA 0.38039f
C656 bgr_11_0.V_TOP.n15 GNDA 0.391025f
C657 bgr_11_0.V_TOP.t41 GNDA 0.38039f
C658 bgr_11_0.V_TOP.t15 GNDA 0.374019f
C659 bgr_11_0.V_TOP.n16 GNDA 0.320897f
C660 bgr_11_0.V_TOP.t28 GNDA 0.374019f
C661 bgr_11_0.V_TOP.n17 GNDA 0.163634f
C662 bgr_11_0.V_TOP.n18 GNDA 0.875119f
C663 bgr_11_0.V_TOP.t6 GNDA 0.105245f
C664 bgr_11_0.V_TOP.n19 GNDA 1.42428f
C665 bgr_11_0.V_TOP.n20 GNDA 0.019145f
C666 bgr_11_0.V_TOP.n21 GNDA 0.024925f
C667 bgr_11_0.V_TOP.n22 GNDA 0.022551f
C668 bgr_11_0.V_TOP.n23 GNDA 0.25922f
C669 bgr_11_0.V_TOP.n24 GNDA 0.158514f
C670 bgr_11_0.V_TOP.n25 GNDA 0.655866f
C671 bgr_11_0.V_TOP.n26 GNDA 0.020198f
C672 bgr_11_0.V_TOP.n27 GNDA 0.198604f
C673 bgr_11_0.V_TOP.n28 GNDA 0.020198f
C674 bgr_11_0.V_TOP.n29 GNDA 0.204214f
C675 bgr_11_0.V_TOP.n30 GNDA 0.020198f
C676 bgr_11_0.V_TOP.n31 GNDA 0.190361f
C677 bgr_11_0.V_TOP.n32 GNDA 0.391697f
C678 bgr_11_0.V_TOP.n33 GNDA 0.089765f
C679 bgr_11_0.V_TOP.t14 GNDA 0.127788f
C680 bgr_11_0.V_TOP.n34 GNDA 0.052677f
C681 bgr_11_0.V_TOP.n35 GNDA 0.025246f
C682 bgr_11_0.V_TOP.t45 GNDA 0.128533f
C683 bgr_11_0.V_TOP.n36 GNDA 0.084658f
C684 bgr_11_0.V_TOP.t36 GNDA 0.129529f
C685 bgr_11_0.V_TOP.n37 GNDA 0.089272f
C686 bgr_11_0.V_TOP.t25 GNDA 0.129529f
C687 bgr_11_0.V_TOP.n38 GNDA 0.089272f
C688 bgr_11_0.V_TOP.t26 GNDA 0.129529f
C689 bgr_11_0.V_TOP.n39 GNDA 0.089272f
C690 bgr_11_0.V_TOP.t49 GNDA 0.129529f
C691 bgr_11_0.V_TOP.n40 GNDA 0.089272f
C692 bgr_11_0.V_TOP.t42 GNDA 0.129529f
C693 bgr_11_0.V_TOP.n41 GNDA 0.089272f
C694 bgr_11_0.V_TOP.t33 GNDA 0.129529f
C695 bgr_11_0.V_TOP.n42 GNDA 0.080857f
C696 bgr_11_0.V_TOP.t21 GNDA 0.128562f
C697 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t4 GNDA 0.02058f
C698 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t3 GNDA 0.02058f
C699 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n0 GNDA 0.051609f
C700 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t1 GNDA 0.02058f
C701 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t0 GNDA 0.02058f
C702 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n1 GNDA 0.051337f
C703 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n2 GNDA 0.456371f
C704 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t2 GNDA 0.02058f
C705 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t5 GNDA 0.02058f
C706 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n3 GNDA 0.04116f
C707 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n4 GNDA 0.077143f
C708 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t16 GNDA 0.259571f
C709 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n5 GNDA 0.065012f
C710 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n6 GNDA 0.114994f
C711 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t8 GNDA 0.04116f
C712 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t11 GNDA 0.04116f
C713 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n7 GNDA 0.084156f
C714 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n8 GNDA 0.282677f
C715 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t15 GNDA 0.04116f
C716 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t10 GNDA 0.04116f
C717 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n9 GNDA 0.084156f
C718 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n10 GNDA 0.27222f
C719 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n11 GNDA 0.110539f
C720 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n12 GNDA 0.065012f
C721 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t14 GNDA 0.04116f
C722 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t9 GNDA 0.04116f
C723 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n13 GNDA 0.084156f
C724 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n14 GNDA 0.27222f
C725 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n15 GNDA 0.067389f
C726 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t7 GNDA 0.04116f
C727 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t13 GNDA 0.04116f
C728 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n16 GNDA 0.084156f
C729 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n17 GNDA 0.27222f
C730 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n18 GNDA 0.114994f
C731 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t6 GNDA 0.04116f
C732 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.t12 GNDA 0.04116f
C733 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n19 GNDA 0.084156f
C734 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n20 GNDA 0.277598f
C735 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n21 GNDA 0.150028f
C736 two_stage_opamp_dummy_magic_24_0.V_CMFB_S3.n22 GNDA 2.49812f
C737 bgr_11_0.V_CMFB_S3 GNDA 2.64392f
C738 two_stage_opamp_dummy_magic_24_0.Y.n0 GNDA 0.080895f
C739 two_stage_opamp_dummy_magic_24_0.Y.n1 GNDA 0.089884f
C740 two_stage_opamp_dummy_magic_24_0.Y.n2 GNDA 0.098872f
C741 two_stage_opamp_dummy_magic_24_0.Y.n3 GNDA 0.338887f
C742 two_stage_opamp_dummy_magic_24_0.Y.n4 GNDA 0.089884f
C743 two_stage_opamp_dummy_magic_24_0.Y.n5 GNDA 0.089884f
C744 two_stage_opamp_dummy_magic_24_0.Y.t20 GNDA 0.022471f
C745 two_stage_opamp_dummy_magic_24_0.Y.t1 GNDA 0.022471f
C746 two_stage_opamp_dummy_magic_24_0.Y.n6 GNDA 0.066035f
C747 two_stage_opamp_dummy_magic_24_0.Y.t21 GNDA 0.022471f
C748 two_stage_opamp_dummy_magic_24_0.Y.t14 GNDA 0.022471f
C749 two_stage_opamp_dummy_magic_24_0.Y.n7 GNDA 0.064754f
C750 two_stage_opamp_dummy_magic_24_0.Y.n8 GNDA 0.427989f
C751 two_stage_opamp_dummy_magic_24_0.Y.t22 GNDA 0.022471f
C752 two_stage_opamp_dummy_magic_24_0.Y.t15 GNDA 0.022471f
C753 two_stage_opamp_dummy_magic_24_0.Y.n9 GNDA 0.064754f
C754 two_stage_opamp_dummy_magic_24_0.Y.n10 GNDA 0.225121f
C755 two_stage_opamp_dummy_magic_24_0.Y.t19 GNDA 0.022471f
C756 two_stage_opamp_dummy_magic_24_0.Y.t17 GNDA 0.022471f
C757 two_stage_opamp_dummy_magic_24_0.Y.n11 GNDA 0.064754f
C758 two_stage_opamp_dummy_magic_24_0.Y.n12 GNDA 0.225121f
C759 two_stage_opamp_dummy_magic_24_0.Y.t13 GNDA 0.022471f
C760 two_stage_opamp_dummy_magic_24_0.Y.t16 GNDA 0.022471f
C761 two_stage_opamp_dummy_magic_24_0.Y.n13 GNDA 0.064754f
C762 two_stage_opamp_dummy_magic_24_0.Y.n14 GNDA 0.225121f
C763 two_stage_opamp_dummy_magic_24_0.Y.t0 GNDA 0.022471f
C764 two_stage_opamp_dummy_magic_24_0.Y.t18 GNDA 0.022471f
C765 two_stage_opamp_dummy_magic_24_0.Y.n15 GNDA 0.064754f
C766 two_stage_opamp_dummy_magic_24_0.Y.n16 GNDA 0.400394f
C767 two_stage_opamp_dummy_magic_24_0.Y.n17 GNDA 0.268572f
C768 two_stage_opamp_dummy_magic_24_0.Y.n18 GNDA 0.395173f
C769 two_stage_opamp_dummy_magic_24_0.Y.n19 GNDA 0.335138f
C770 two_stage_opamp_dummy_magic_24_0.Y.n20 GNDA 0.098872f
C771 two_stage_opamp_dummy_magic_24_0.Y.n21 GNDA 0.302609f
C772 two_stage_opamp_dummy_magic_24_0.Y.n22 GNDA 0.098872f
C773 two_stage_opamp_dummy_magic_24_0.Y.n23 GNDA 0.098872f
C774 two_stage_opamp_dummy_magic_24_0.Y.n24 GNDA 0.098872f
C775 two_stage_opamp_dummy_magic_24_0.Y.n25 GNDA 0.154826f
C776 two_stage_opamp_dummy_magic_24_0.Y.n26 GNDA 0.071907f
C777 two_stage_opamp_dummy_magic_24_0.Y.t54 GNDA 0.048313f
C778 two_stage_opamp_dummy_magic_24_0.Y.t38 GNDA 0.048313f
C779 two_stage_opamp_dummy_magic_24_0.Y.t27 GNDA 0.048313f
C780 two_stage_opamp_dummy_magic_24_0.Y.t42 GNDA 0.048313f
C781 two_stage_opamp_dummy_magic_24_0.Y.t49 GNDA 0.048313f
C782 two_stage_opamp_dummy_magic_24_0.Y.t31 GNDA 0.048313f
C783 two_stage_opamp_dummy_magic_24_0.Y.t51 GNDA 0.048313f
C784 two_stage_opamp_dummy_magic_24_0.Y.t33 GNDA 0.054923f
C785 two_stage_opamp_dummy_magic_24_0.Y.n29 GNDA 0.049567f
C786 two_stage_opamp_dummy_magic_24_0.Y.n30 GNDA 0.030336f
C787 two_stage_opamp_dummy_magic_24_0.Y.n31 GNDA 0.030336f
C788 two_stage_opamp_dummy_magic_24_0.Y.n32 GNDA 0.030336f
C789 two_stage_opamp_dummy_magic_24_0.Y.n33 GNDA 0.030336f
C790 two_stage_opamp_dummy_magic_24_0.Y.n34 GNDA 0.030336f
C791 two_stage_opamp_dummy_magic_24_0.Y.n35 GNDA 0.025561f
C792 two_stage_opamp_dummy_magic_24_0.Y.t34 GNDA 0.048313f
C793 two_stage_opamp_dummy_magic_24_0.Y.t43 GNDA 0.054923f
C794 two_stage_opamp_dummy_magic_24_0.Y.n36 GNDA 0.044792f
C795 two_stage_opamp_dummy_magic_24_0.Y.n37 GNDA 0.012412f
C796 two_stage_opamp_dummy_magic_24_0.Y.t26 GNDA 0.031459f
C797 two_stage_opamp_dummy_magic_24_0.Y.t41 GNDA 0.031459f
C798 two_stage_opamp_dummy_magic_24_0.Y.t29 GNDA 0.031459f
C799 two_stage_opamp_dummy_magic_24_0.Y.t45 GNDA 0.031459f
C800 two_stage_opamp_dummy_magic_24_0.Y.t50 GNDA 0.031459f
C801 two_stage_opamp_dummy_magic_24_0.Y.t32 GNDA 0.031459f
C802 two_stage_opamp_dummy_magic_24_0.Y.t53 GNDA 0.031459f
C803 two_stage_opamp_dummy_magic_24_0.Y.t36 GNDA 0.038201f
C804 two_stage_opamp_dummy_magic_24_0.Y.n38 GNDA 0.038201f
C805 two_stage_opamp_dummy_magic_24_0.Y.n39 GNDA 0.024718f
C806 two_stage_opamp_dummy_magic_24_0.Y.n40 GNDA 0.024718f
C807 two_stage_opamp_dummy_magic_24_0.Y.n41 GNDA 0.024718f
C808 two_stage_opamp_dummy_magic_24_0.Y.n42 GNDA 0.024718f
C809 two_stage_opamp_dummy_magic_24_0.Y.n43 GNDA 0.024718f
C810 two_stage_opamp_dummy_magic_24_0.Y.n44 GNDA 0.019943f
C811 two_stage_opamp_dummy_magic_24_0.Y.t37 GNDA 0.031459f
C812 two_stage_opamp_dummy_magic_24_0.Y.t46 GNDA 0.038201f
C813 two_stage_opamp_dummy_magic_24_0.Y.n45 GNDA 0.033425f
C814 two_stage_opamp_dummy_magic_24_0.Y.n46 GNDA 0.012412f
C815 two_stage_opamp_dummy_magic_24_0.Y.n47 GNDA 0.077428f
C816 two_stage_opamp_dummy_magic_24_0.Y.n48 GNDA 0.071907f
C817 two_stage_opamp_dummy_magic_24_0.Y.n49 GNDA 0.071232f
C818 two_stage_opamp_dummy_magic_24_0.Y.n50 GNDA 0.071907f
C819 two_stage_opamp_dummy_magic_24_0.Y.t12 GNDA 0.621783f
C820 two_stage_opamp_dummy_magic_24_0.Y.n51 GNDA 0.071907f
C821 two_stage_opamp_dummy_magic_24_0.Y.n52 GNDA 0.071907f
C822 two_stage_opamp_dummy_magic_24_0.Y.n54 GNDA 0.66715f
C823 two_stage_opamp_dummy_magic_24_0.Y.n56 GNDA 0.624692f
C824 two_stage_opamp_dummy_magic_24_0.Y.n57 GNDA 0.02381f
C825 two_stage_opamp_dummy_magic_24_0.Y.n58 GNDA 0.023969f
C826 two_stage_opamp_dummy_magic_24_0.Y.n59 GNDA 0.023969f
C827 two_stage_opamp_dummy_magic_24_0.Y.t47 GNDA 0.098872f
C828 two_stage_opamp_dummy_magic_24_0.Y.t52 GNDA 0.098872f
C829 two_stage_opamp_dummy_magic_24_0.Y.t35 GNDA 0.098872f
C830 two_stage_opamp_dummy_magic_24_0.Y.t25 GNDA 0.098872f
C831 two_stage_opamp_dummy_magic_24_0.Y.t39 GNDA 0.105306f
C832 two_stage_opamp_dummy_magic_24_0.Y.n60 GNDA 0.08345f
C833 two_stage_opamp_dummy_magic_24_0.Y.n61 GNDA 0.047189f
C834 two_stage_opamp_dummy_magic_24_0.Y.n62 GNDA 0.047189f
C835 two_stage_opamp_dummy_magic_24_0.Y.n63 GNDA 0.042414f
C836 two_stage_opamp_dummy_magic_24_0.Y.t30 GNDA 0.098872f
C837 two_stage_opamp_dummy_magic_24_0.Y.t44 GNDA 0.098872f
C838 two_stage_opamp_dummy_magic_24_0.Y.t28 GNDA 0.098872f
C839 two_stage_opamp_dummy_magic_24_0.Y.t40 GNDA 0.098872f
C840 two_stage_opamp_dummy_magic_24_0.Y.t48 GNDA 0.105306f
C841 two_stage_opamp_dummy_magic_24_0.Y.n64 GNDA 0.08345f
C842 two_stage_opamp_dummy_magic_24_0.Y.n65 GNDA 0.047189f
C843 two_stage_opamp_dummy_magic_24_0.Y.n66 GNDA 0.047189f
C844 two_stage_opamp_dummy_magic_24_0.Y.n67 GNDA 0.042414f
C845 two_stage_opamp_dummy_magic_24_0.Y.n68 GNDA 0.010184f
C846 two_stage_opamp_dummy_magic_24_0.Y.n69 GNDA 0.024128f
C847 two_stage_opamp_dummy_magic_24_0.Y.n70 GNDA 0.056796f
C848 two_stage_opamp_dummy_magic_24_0.Y.n71 GNDA 0.032394f
C849 two_stage_opamp_dummy_magic_24_0.Y.n72 GNDA 0.036763f
C850 two_stage_opamp_dummy_magic_24_0.Y.n73 GNDA 0.993216f
C851 two_stage_opamp_dummy_magic_24_0.Y.n74 GNDA 0.080841f
C852 two_stage_opamp_dummy_magic_24_0.Y.n75 GNDA 0.056872f
C853 two_stage_opamp_dummy_magic_24_0.Y.t23 GNDA 0.052432f
C854 two_stage_opamp_dummy_magic_24_0.Y.t4 GNDA 0.052432f
C855 two_stage_opamp_dummy_magic_24_0.Y.n76 GNDA 0.107256f
C856 two_stage_opamp_dummy_magic_24_0.Y.n77 GNDA 0.346283f
C857 two_stage_opamp_dummy_magic_24_0.Y.n78 GNDA 0.097017f
C858 two_stage_opamp_dummy_magic_24_0.Y.t6 GNDA 0.052432f
C859 two_stage_opamp_dummy_magic_24_0.Y.t9 GNDA 0.052432f
C860 two_stage_opamp_dummy_magic_24_0.Y.n79 GNDA 0.107256f
C861 two_stage_opamp_dummy_magic_24_0.Y.n80 GNDA 0.337778f
C862 two_stage_opamp_dummy_magic_24_0.Y.n81 GNDA 0.133949f
C863 two_stage_opamp_dummy_magic_24_0.Y.t11 GNDA 0.052432f
C864 two_stage_opamp_dummy_magic_24_0.Y.t2 GNDA 0.052432f
C865 two_stage_opamp_dummy_magic_24_0.Y.n82 GNDA 0.107256f
C866 two_stage_opamp_dummy_magic_24_0.Y.n83 GNDA 0.337778f
C867 two_stage_opamp_dummy_magic_24_0.Y.n84 GNDA 0.080841f
C868 two_stage_opamp_dummy_magic_24_0.Y.n85 GNDA 0.080841f
C869 two_stage_opamp_dummy_magic_24_0.Y.t3 GNDA 0.052432f
C870 two_stage_opamp_dummy_magic_24_0.Y.t5 GNDA 0.052432f
C871 two_stage_opamp_dummy_magic_24_0.Y.n86 GNDA 0.107256f
C872 two_stage_opamp_dummy_magic_24_0.Y.n87 GNDA 0.337778f
C873 two_stage_opamp_dummy_magic_24_0.Y.n88 GNDA 0.056872f
C874 two_stage_opamp_dummy_magic_24_0.Y.t7 GNDA 0.052432f
C875 two_stage_opamp_dummy_magic_24_0.Y.t10 GNDA 0.052432f
C876 two_stage_opamp_dummy_magic_24_0.Y.n89 GNDA 0.107256f
C877 two_stage_opamp_dummy_magic_24_0.Y.n90 GNDA 0.337778f
C878 two_stage_opamp_dummy_magic_24_0.Y.n91 GNDA 0.097017f
C879 two_stage_opamp_dummy_magic_24_0.Y.t8 GNDA 0.052432f
C880 two_stage_opamp_dummy_magic_24_0.Y.t24 GNDA 0.052432f
C881 two_stage_opamp_dummy_magic_24_0.Y.n92 GNDA 0.107256f
C882 two_stage_opamp_dummy_magic_24_0.Y.n93 GNDA 0.34252f
C883 two_stage_opamp_dummy_magic_24_0.Y.n94 GNDA 0.599255f
C884 two_stage_opamp_dummy_magic_24_0.Y.n95 GNDA 1.82456f
C885 two_stage_opamp_dummy_magic_24_0.Y.n97 GNDA 0.44043f
C886 two_stage_opamp_dummy_magic_24_0.Y.n98 GNDA 2.12499f
C887 two_stage_opamp_dummy_magic_24_0.Y.n99 GNDA 0.57975f
C888 two_stage_opamp_dummy_magic_24_0.Y.n100 GNDA 0.593233f
C889 two_stage_opamp_dummy_magic_24_0.Y.n101 GNDA 0.293095f
C890 two_stage_opamp_dummy_magic_24_0.Y.n102 GNDA 0.098872f
C891 two_stage_opamp_dummy_magic_24_0.Y.n103 GNDA 0.302609f
C892 two_stage_opamp_dummy_magic_24_0.Y.n104 GNDA 0.098872f
C893 two_stage_opamp_dummy_magic_24_0.Y.n105 GNDA 0.098872f
C894 two_stage_opamp_dummy_magic_24_0.Y.n106 GNDA 0.098872f
C895 two_stage_opamp_dummy_magic_24_0.Y.n107 GNDA 0.271149f
C896 two_stage_opamp_dummy_magic_24_0.Vb1_2.t1 GNDA 0.046205f
C897 two_stage_opamp_dummy_magic_24_0.Vb1_2.n0 GNDA 0.312531f
C898 two_stage_opamp_dummy_magic_24_0.Vb1_2.t4 GNDA 0.157018f
C899 two_stage_opamp_dummy_magic_24_0.Vb1_2.n1 GNDA 0.539239f
C900 two_stage_opamp_dummy_magic_24_0.Vb1_2.t2 GNDA 0.046205f
C901 two_stage_opamp_dummy_magic_24_0.Vb1_2.t0 GNDA 0.046205f
C902 two_stage_opamp_dummy_magic_24_0.Vb1_2.n2 GNDA 0.100536f
C903 two_stage_opamp_dummy_magic_24_0.Vb1_2.n3 GNDA 0.474689f
C904 two_stage_opamp_dummy_magic_24_0.Vb1_2.n4 GNDA 0.470919f
C905 two_stage_opamp_dummy_magic_24_0.Vb1_2.n5 GNDA 0.459714f
C906 two_stage_opamp_dummy_magic_24_0.Vb1_2.n6 GNDA 0.100536f
C907 two_stage_opamp_dummy_magic_24_0.Vb1_2.t3 GNDA 0.046205f
C908 two_stage_opamp_dummy_magic_24_0.Vb1.n0 GNDA 0.237532f
C909 two_stage_opamp_dummy_magic_24_0.Vb1.n1 GNDA 3.87535f
C910 two_stage_opamp_dummy_magic_24_0.Vb1.n2 GNDA 0.198304f
C911 two_stage_opamp_dummy_magic_24_0.Vb1.n3 GNDA 0.337191f
C912 two_stage_opamp_dummy_magic_24_0.Vb1.n4 GNDA 0.162417f
C913 two_stage_opamp_dummy_magic_24_0.Vb1.n5 GNDA 0.337191f
C914 two_stage_opamp_dummy_magic_24_0.Vb1.n6 GNDA 0.415806f
C915 two_stage_opamp_dummy_magic_24_0.Vb1.n7 GNDA 0.56577f
C916 two_stage_opamp_dummy_magic_24_0.Vb1.n8 GNDA 0.282752f
C917 two_stage_opamp_dummy_magic_24_0.Vb1.n9 GNDA 0.408201f
C918 two_stage_opamp_dummy_magic_24_0.Vb1.n10 GNDA 0.415806f
C919 two_stage_opamp_dummy_magic_24_0.Vb1.n11 GNDA 0.282752f
C920 two_stage_opamp_dummy_magic_24_0.Vb1.t11 GNDA 0.034413f
C921 two_stage_opamp_dummy_magic_24_0.Vb1.t10 GNDA 0.034413f
C922 two_stage_opamp_dummy_magic_24_0.Vb1.n12 GNDA 0.078293f
C923 two_stage_opamp_dummy_magic_24_0.Vb1.t2 GNDA 0.026455f
C924 two_stage_opamp_dummy_magic_24_0.Vb1.t4 GNDA 0.034313f
C925 two_stage_opamp_dummy_magic_24_0.Vb1.n13 GNDA 0.035278f
C926 two_stage_opamp_dummy_magic_24_0.Vb1.t6 GNDA 0.026455f
C927 two_stage_opamp_dummy_magic_24_0.Vb1.t8 GNDA 0.034313f
C928 two_stage_opamp_dummy_magic_24_0.Vb1.n14 GNDA 0.035278f
C929 two_stage_opamp_dummy_magic_24_0.Vb1.n15 GNDA 0.026296f
C930 two_stage_opamp_dummy_magic_24_0.Vb1.t12 GNDA 0.992567f
C931 two_stage_opamp_dummy_magic_24_0.Vb1.t0 GNDA 0.02581f
C932 two_stage_opamp_dummy_magic_24_0.Vb1.t5 GNDA 0.02581f
C933 two_stage_opamp_dummy_magic_24_0.Vb1.n16 GNDA 0.056159f
C934 two_stage_opamp_dummy_magic_24_0.Vb1.n17 GNDA 0.207472f
C935 two_stage_opamp_dummy_magic_24_0.Vb1.t3 GNDA 0.02581f
C936 two_stage_opamp_dummy_magic_24_0.Vb1.t7 GNDA 0.02581f
C937 two_stage_opamp_dummy_magic_24_0.Vb1.n18 GNDA 0.056159f
C938 two_stage_opamp_dummy_magic_24_0.Vb1.t9 GNDA 0.02581f
C939 two_stage_opamp_dummy_magic_24_0.Vb1.t1 GNDA 0.02581f
C940 two_stage_opamp_dummy_magic_24_0.Vb1.n19 GNDA 0.065328f
C941 two_stage_opamp_dummy_magic_24_0.Vb1.t22 GNDA 0.04079f
C942 two_stage_opamp_dummy_magic_24_0.Vb1.t15 GNDA 0.040756f
C943 two_stage_opamp_dummy_magic_24_0.Vb1.t28 GNDA 0.040756f
C944 two_stage_opamp_dummy_magic_24_0.Vb1.t18 GNDA 0.040756f
C945 two_stage_opamp_dummy_magic_24_0.Vb1.t30 GNDA 0.040756f
C946 two_stage_opamp_dummy_magic_24_0.Vb1.t17 GNDA 0.040756f
C947 two_stage_opamp_dummy_magic_24_0.Vb1.t29 GNDA 0.040756f
C948 two_stage_opamp_dummy_magic_24_0.Vb1.t20 GNDA 0.040756f
C949 two_stage_opamp_dummy_magic_24_0.Vb1.t31 GNDA 0.040756f
C950 two_stage_opamp_dummy_magic_24_0.Vb1.t21 GNDA 0.040756f
C951 two_stage_opamp_dummy_magic_24_0.Vb1.t23 GNDA 0.040756f
C952 two_stage_opamp_dummy_magic_24_0.Vb1.t32 GNDA 0.040756f
C953 two_stage_opamp_dummy_magic_24_0.Vb1.t25 GNDA 0.040756f
C954 two_stage_opamp_dummy_magic_24_0.Vb1.t19 GNDA 0.040756f
C955 two_stage_opamp_dummy_magic_24_0.Vb1.t24 GNDA 0.040756f
C956 two_stage_opamp_dummy_magic_24_0.Vb1.t13 GNDA 0.040756f
C957 two_stage_opamp_dummy_magic_24_0.Vb1.t26 GNDA 0.040756f
C958 two_stage_opamp_dummy_magic_24_0.Vb1.t14 GNDA 0.040756f
C959 two_stage_opamp_dummy_magic_24_0.Vb1.t27 GNDA 0.040756f
C960 two_stage_opamp_dummy_magic_24_0.Vb1.t16 GNDA 0.040756f
C961 two_stage_opamp_dummy_magic_24_0.Vb1.n20 GNDA 4.98332f
C962 two_stage_opamp_dummy_magic_24_0.X.n0 GNDA 0.067413f
C963 two_stage_opamp_dummy_magic_24_0.X.n1 GNDA 0.098872f
C964 two_stage_opamp_dummy_magic_24_0.X.n2 GNDA 0.302609f
C965 two_stage_opamp_dummy_magic_24_0.X.n3 GNDA 0.293095f
C966 two_stage_opamp_dummy_magic_24_0.X.n4 GNDA 0.098872f
C967 two_stage_opamp_dummy_magic_24_0.X.n5 GNDA 0.098872f
C968 two_stage_opamp_dummy_magic_24_0.X.n6 GNDA 0.071907f
C969 two_stage_opamp_dummy_magic_24_0.X.t28 GNDA 0.048313f
C970 two_stage_opamp_dummy_magic_24_0.X.t43 GNDA 0.054923f
C971 two_stage_opamp_dummy_magic_24_0.X.n9 GNDA 0.044792f
C972 two_stage_opamp_dummy_magic_24_0.X.t40 GNDA 0.048313f
C973 two_stage_opamp_dummy_magic_24_0.X.t54 GNDA 0.048313f
C974 two_stage_opamp_dummy_magic_24_0.X.t36 GNDA 0.048313f
C975 two_stage_opamp_dummy_magic_24_0.X.t49 GNDA 0.048313f
C976 two_stage_opamp_dummy_magic_24_0.X.t32 GNDA 0.048313f
C977 two_stage_opamp_dummy_magic_24_0.X.t50 GNDA 0.048313f
C978 two_stage_opamp_dummy_magic_24_0.X.t33 GNDA 0.048313f
C979 two_stage_opamp_dummy_magic_24_0.X.t47 GNDA 0.054923f
C980 two_stage_opamp_dummy_magic_24_0.X.n10 GNDA 0.049567f
C981 two_stage_opamp_dummy_magic_24_0.X.n11 GNDA 0.030336f
C982 two_stage_opamp_dummy_magic_24_0.X.n12 GNDA 0.030336f
C983 two_stage_opamp_dummy_magic_24_0.X.n13 GNDA 0.030336f
C984 two_stage_opamp_dummy_magic_24_0.X.n14 GNDA 0.030336f
C985 two_stage_opamp_dummy_magic_24_0.X.n15 GNDA 0.030336f
C986 two_stage_opamp_dummy_magic_24_0.X.n16 GNDA 0.025561f
C987 two_stage_opamp_dummy_magic_24_0.X.n17 GNDA 0.012412f
C988 two_stage_opamp_dummy_magic_24_0.X.t30 GNDA 0.031459f
C989 two_stage_opamp_dummy_magic_24_0.X.t45 GNDA 0.038201f
C990 two_stage_opamp_dummy_magic_24_0.X.n18 GNDA 0.033425f
C991 two_stage_opamp_dummy_magic_24_0.X.t42 GNDA 0.031459f
C992 two_stage_opamp_dummy_magic_24_0.X.t27 GNDA 0.031459f
C993 two_stage_opamp_dummy_magic_24_0.X.t39 GNDA 0.031459f
C994 two_stage_opamp_dummy_magic_24_0.X.t52 GNDA 0.031459f
C995 two_stage_opamp_dummy_magic_24_0.X.t34 GNDA 0.031459f
C996 two_stage_opamp_dummy_magic_24_0.X.t53 GNDA 0.031459f
C997 two_stage_opamp_dummy_magic_24_0.X.t35 GNDA 0.031459f
C998 two_stage_opamp_dummy_magic_24_0.X.t48 GNDA 0.038201f
C999 two_stage_opamp_dummy_magic_24_0.X.n19 GNDA 0.038201f
C1000 two_stage_opamp_dummy_magic_24_0.X.n20 GNDA 0.024718f
C1001 two_stage_opamp_dummy_magic_24_0.X.n21 GNDA 0.024718f
C1002 two_stage_opamp_dummy_magic_24_0.X.n22 GNDA 0.024718f
C1003 two_stage_opamp_dummy_magic_24_0.X.n23 GNDA 0.024718f
C1004 two_stage_opamp_dummy_magic_24_0.X.n24 GNDA 0.024718f
C1005 two_stage_opamp_dummy_magic_24_0.X.n25 GNDA 0.019943f
C1006 two_stage_opamp_dummy_magic_24_0.X.n26 GNDA 0.012412f
C1007 two_stage_opamp_dummy_magic_24_0.X.n27 GNDA 0.077423f
C1008 two_stage_opamp_dummy_magic_24_0.X.n29 GNDA 0.071907f
C1009 two_stage_opamp_dummy_magic_24_0.X.t19 GNDA 0.621783f
C1010 two_stage_opamp_dummy_magic_24_0.X.n30 GNDA 0.071907f
C1011 two_stage_opamp_dummy_magic_24_0.X.n31 GNDA 0.071907f
C1012 two_stage_opamp_dummy_magic_24_0.X.n32 GNDA 0.071232f
C1013 two_stage_opamp_dummy_magic_24_0.X.n33 GNDA 0.66715f
C1014 two_stage_opamp_dummy_magic_24_0.X.n35 GNDA 0.624692f
C1015 two_stage_opamp_dummy_magic_24_0.X.n36 GNDA 0.02381f
C1016 two_stage_opamp_dummy_magic_24_0.X.n37 GNDA 0.023969f
C1017 two_stage_opamp_dummy_magic_24_0.X.n38 GNDA 0.023969f
C1018 two_stage_opamp_dummy_magic_24_0.X.t41 GNDA 0.098872f
C1019 two_stage_opamp_dummy_magic_24_0.X.t29 GNDA 0.098872f
C1020 two_stage_opamp_dummy_magic_24_0.X.t44 GNDA 0.098872f
C1021 two_stage_opamp_dummy_magic_24_0.X.t31 GNDA 0.098872f
C1022 two_stage_opamp_dummy_magic_24_0.X.t46 GNDA 0.105306f
C1023 two_stage_opamp_dummy_magic_24_0.X.n39 GNDA 0.08345f
C1024 two_stage_opamp_dummy_magic_24_0.X.n40 GNDA 0.047189f
C1025 two_stage_opamp_dummy_magic_24_0.X.n41 GNDA 0.047189f
C1026 two_stage_opamp_dummy_magic_24_0.X.n42 GNDA 0.042414f
C1027 two_stage_opamp_dummy_magic_24_0.X.t25 GNDA 0.098872f
C1028 two_stage_opamp_dummy_magic_24_0.X.t37 GNDA 0.098872f
C1029 two_stage_opamp_dummy_magic_24_0.X.t26 GNDA 0.098872f
C1030 two_stage_opamp_dummy_magic_24_0.X.t38 GNDA 0.098872f
C1031 two_stage_opamp_dummy_magic_24_0.X.t51 GNDA 0.105306f
C1032 two_stage_opamp_dummy_magic_24_0.X.n43 GNDA 0.08345f
C1033 two_stage_opamp_dummy_magic_24_0.X.n44 GNDA 0.047189f
C1034 two_stage_opamp_dummy_magic_24_0.X.n45 GNDA 0.047189f
C1035 two_stage_opamp_dummy_magic_24_0.X.n46 GNDA 0.042414f
C1036 two_stage_opamp_dummy_magic_24_0.X.n47 GNDA 0.010184f
C1037 two_stage_opamp_dummy_magic_24_0.X.n48 GNDA 0.024128f
C1038 two_stage_opamp_dummy_magic_24_0.X.n49 GNDA 0.056796f
C1039 two_stage_opamp_dummy_magic_24_0.X.n50 GNDA 0.032394f
C1040 two_stage_opamp_dummy_magic_24_0.X.n51 GNDA 0.036763f
C1041 two_stage_opamp_dummy_magic_24_0.X.n52 GNDA 0.993216f
C1042 two_stage_opamp_dummy_magic_24_0.X.n53 GNDA 0.071907f
C1043 two_stage_opamp_dummy_magic_24_0.X.n54 GNDA 0.080841f
C1044 two_stage_opamp_dummy_magic_24_0.X.n55 GNDA 0.056872f
C1045 two_stage_opamp_dummy_magic_24_0.X.t13 GNDA 0.052432f
C1046 two_stage_opamp_dummy_magic_24_0.X.t21 GNDA 0.052432f
C1047 two_stage_opamp_dummy_magic_24_0.X.n56 GNDA 0.107256f
C1048 two_stage_opamp_dummy_magic_24_0.X.n57 GNDA 0.346283f
C1049 two_stage_opamp_dummy_magic_24_0.X.n58 GNDA 0.097017f
C1050 two_stage_opamp_dummy_magic_24_0.X.t8 GNDA 0.052432f
C1051 two_stage_opamp_dummy_magic_24_0.X.t10 GNDA 0.052432f
C1052 two_stage_opamp_dummy_magic_24_0.X.n59 GNDA 0.107256f
C1053 two_stage_opamp_dummy_magic_24_0.X.n60 GNDA 0.337778f
C1054 two_stage_opamp_dummy_magic_24_0.X.n61 GNDA 0.133949f
C1055 two_stage_opamp_dummy_magic_24_0.X.t7 GNDA 0.052432f
C1056 two_stage_opamp_dummy_magic_24_0.X.t9 GNDA 0.052432f
C1057 two_stage_opamp_dummy_magic_24_0.X.n62 GNDA 0.107256f
C1058 two_stage_opamp_dummy_magic_24_0.X.n63 GNDA 0.337778f
C1059 two_stage_opamp_dummy_magic_24_0.X.n64 GNDA 0.080841f
C1060 two_stage_opamp_dummy_magic_24_0.X.n65 GNDA 0.080841f
C1061 two_stage_opamp_dummy_magic_24_0.X.t5 GNDA 0.052432f
C1062 two_stage_opamp_dummy_magic_24_0.X.t6 GNDA 0.052432f
C1063 two_stage_opamp_dummy_magic_24_0.X.n66 GNDA 0.107256f
C1064 two_stage_opamp_dummy_magic_24_0.X.n67 GNDA 0.337778f
C1065 two_stage_opamp_dummy_magic_24_0.X.n68 GNDA 0.056872f
C1066 two_stage_opamp_dummy_magic_24_0.X.t14 GNDA 0.052432f
C1067 two_stage_opamp_dummy_magic_24_0.X.t12 GNDA 0.052432f
C1068 two_stage_opamp_dummy_magic_24_0.X.n69 GNDA 0.107256f
C1069 two_stage_opamp_dummy_magic_24_0.X.n70 GNDA 0.337778f
C1070 two_stage_opamp_dummy_magic_24_0.X.n71 GNDA 0.097017f
C1071 two_stage_opamp_dummy_magic_24_0.X.t22 GNDA 0.052432f
C1072 two_stage_opamp_dummy_magic_24_0.X.t11 GNDA 0.052432f
C1073 two_stage_opamp_dummy_magic_24_0.X.n72 GNDA 0.107256f
C1074 two_stage_opamp_dummy_magic_24_0.X.n73 GNDA 0.34252f
C1075 two_stage_opamp_dummy_magic_24_0.X.n74 GNDA 0.599223f
C1076 two_stage_opamp_dummy_magic_24_0.X.n75 GNDA 1.82459f
C1077 two_stage_opamp_dummy_magic_24_0.X.n77 GNDA 0.44043f
C1078 two_stage_opamp_dummy_magic_24_0.X.n78 GNDA 2.125f
C1079 two_stage_opamp_dummy_magic_24_0.X.n79 GNDA 0.57975f
C1080 two_stage_opamp_dummy_magic_24_0.X.n80 GNDA 0.593233f
C1081 two_stage_opamp_dummy_magic_24_0.X.n81 GNDA 0.098872f
C1082 two_stage_opamp_dummy_magic_24_0.X.n82 GNDA 0.098872f
C1083 two_stage_opamp_dummy_magic_24_0.X.n83 GNDA 0.098872f
C1084 two_stage_opamp_dummy_magic_24_0.X.n84 GNDA 0.302609f
C1085 two_stage_opamp_dummy_magic_24_0.X.n85 GNDA 0.154826f
C1086 two_stage_opamp_dummy_magic_24_0.X.n86 GNDA 0.089884f
C1087 two_stage_opamp_dummy_magic_24_0.X.n87 GNDA 0.089884f
C1088 two_stage_opamp_dummy_magic_24_0.X.n88 GNDA 0.335139f
C1089 two_stage_opamp_dummy_magic_24_0.X.n89 GNDA 0.089884f
C1090 two_stage_opamp_dummy_magic_24_0.X.t3 GNDA 0.022471f
C1091 two_stage_opamp_dummy_magic_24_0.X.t23 GNDA 0.022471f
C1092 two_stage_opamp_dummy_magic_24_0.X.n90 GNDA 0.066035f
C1093 two_stage_opamp_dummy_magic_24_0.X.t16 GNDA 0.022471f
C1094 two_stage_opamp_dummy_magic_24_0.X.t24 GNDA 0.022471f
C1095 two_stage_opamp_dummy_magic_24_0.X.n91 GNDA 0.064754f
C1096 two_stage_opamp_dummy_magic_24_0.X.n92 GNDA 0.427989f
C1097 two_stage_opamp_dummy_magic_24_0.X.t4 GNDA 0.022471f
C1098 two_stage_opamp_dummy_magic_24_0.X.t17 GNDA 0.022471f
C1099 two_stage_opamp_dummy_magic_24_0.X.n93 GNDA 0.064754f
C1100 two_stage_opamp_dummy_magic_24_0.X.n94 GNDA 0.225121f
C1101 two_stage_opamp_dummy_magic_24_0.X.t15 GNDA 0.022471f
C1102 two_stage_opamp_dummy_magic_24_0.X.t0 GNDA 0.022471f
C1103 two_stage_opamp_dummy_magic_24_0.X.n95 GNDA 0.064754f
C1104 two_stage_opamp_dummy_magic_24_0.X.n96 GNDA 0.225121f
C1105 two_stage_opamp_dummy_magic_24_0.X.t1 GNDA 0.022471f
C1106 two_stage_opamp_dummy_magic_24_0.X.t20 GNDA 0.022471f
C1107 two_stage_opamp_dummy_magic_24_0.X.n97 GNDA 0.064754f
C1108 two_stage_opamp_dummy_magic_24_0.X.n98 GNDA 0.225121f
C1109 two_stage_opamp_dummy_magic_24_0.X.t18 GNDA 0.022471f
C1110 two_stage_opamp_dummy_magic_24_0.X.t2 GNDA 0.022471f
C1111 two_stage_opamp_dummy_magic_24_0.X.n99 GNDA 0.064754f
C1112 two_stage_opamp_dummy_magic_24_0.X.n100 GNDA 0.400394f
C1113 two_stage_opamp_dummy_magic_24_0.X.n101 GNDA 0.268572f
C1114 two_stage_opamp_dummy_magic_24_0.X.n102 GNDA 0.395173f
C1115 two_stage_opamp_dummy_magic_24_0.X.n103 GNDA 0.338887f
C1116 two_stage_opamp_dummy_magic_24_0.X.n104 GNDA 0.098872f
C1117 two_stage_opamp_dummy_magic_24_0.X.n105 GNDA 0.302609f
C1118 two_stage_opamp_dummy_magic_24_0.X.n106 GNDA 0.098872f
C1119 two_stage_opamp_dummy_magic_24_0.X.n107 GNDA 0.080895f
C1120 two_stage_opamp_dummy_magic_24_0.Vb2.n0 GNDA 0.369264f
C1121 two_stage_opamp_dummy_magic_24_0.Vb2.n1 GNDA 0.506091f
C1122 two_stage_opamp_dummy_magic_24_0.Vb2.n2 GNDA 0.427517f
C1123 two_stage_opamp_dummy_magic_24_0.Vb2.n3 GNDA 0.495787f
C1124 two_stage_opamp_dummy_magic_24_0.Vb2.n4 GNDA 0.506091f
C1125 two_stage_opamp_dummy_magic_24_0.Vb2.n5 GNDA 0.331819f
C1126 two_stage_opamp_dummy_magic_24_0.Vb2.t5 GNDA 0.059937f
C1127 two_stage_opamp_dummy_magic_24_0.Vb2.t10 GNDA 0.017125f
C1128 two_stage_opamp_dummy_magic_24_0.Vb2.t2 GNDA 0.017125f
C1129 two_stage_opamp_dummy_magic_24_0.Vb2.n6 GNDA 0.057417f
C1130 two_stage_opamp_dummy_magic_24_0.Vb2.t9 GNDA 0.017125f
C1131 two_stage_opamp_dummy_magic_24_0.Vb2.t0 GNDA 0.017125f
C1132 two_stage_opamp_dummy_magic_24_0.Vb2.n7 GNDA 0.055842f
C1133 two_stage_opamp_dummy_magic_24_0.Vb2.n8 GNDA 0.510081f
C1134 two_stage_opamp_dummy_magic_24_0.Vb2.t8 GNDA 0.017125f
C1135 two_stage_opamp_dummy_magic_24_0.Vb2.t6 GNDA 0.017125f
C1136 two_stage_opamp_dummy_magic_24_0.Vb2.n9 GNDA 0.055842f
C1137 two_stage_opamp_dummy_magic_24_0.Vb2.n10 GNDA 0.334602f
C1138 two_stage_opamp_dummy_magic_24_0.Vb2.t3 GNDA 0.017125f
C1139 two_stage_opamp_dummy_magic_24_0.Vb2.t7 GNDA 0.017125f
C1140 two_stage_opamp_dummy_magic_24_0.Vb2.n11 GNDA 0.055842f
C1141 two_stage_opamp_dummy_magic_24_0.Vb2.n12 GNDA 2.20313f
C1142 two_stage_opamp_dummy_magic_24_0.Vb2.t21 GNDA 0.11016f
C1143 two_stage_opamp_dummy_magic_24_0.Vb2.n13 GNDA 2.01397f
C1144 two_stage_opamp_dummy_magic_24_0.Vb2.t15 GNDA 0.109827f
C1145 two_stage_opamp_dummy_magic_24_0.Vb2.t11 GNDA 0.109798f
C1146 two_stage_opamp_dummy_magic_24_0.Vb2.t13 GNDA 0.109798f
C1147 two_stage_opamp_dummy_magic_24_0.Vb2.t32 GNDA 0.109798f
C1148 two_stage_opamp_dummy_magic_24_0.Vb2.t29 GNDA 0.109798f
C1149 two_stage_opamp_dummy_magic_24_0.Vb2.t25 GNDA 0.109798f
C1150 two_stage_opamp_dummy_magic_24_0.Vb2.t19 GNDA 0.109798f
C1151 two_stage_opamp_dummy_magic_24_0.Vb2.t23 GNDA 0.109798f
C1152 two_stage_opamp_dummy_magic_24_0.Vb2.t17 GNDA 0.109798f
C1153 two_stage_opamp_dummy_magic_24_0.Vb2.t12 GNDA 0.109798f
C1154 two_stage_opamp_dummy_magic_24_0.Vb2.t20 GNDA 0.109827f
C1155 two_stage_opamp_dummy_magic_24_0.Vb2.t16 GNDA 0.109798f
C1156 two_stage_opamp_dummy_magic_24_0.Vb2.t22 GNDA 0.109798f
C1157 two_stage_opamp_dummy_magic_24_0.Vb2.t26 GNDA 0.109798f
C1158 two_stage_opamp_dummy_magic_24_0.Vb2.t28 GNDA 0.109798f
C1159 two_stage_opamp_dummy_magic_24_0.Vb2.t30 GNDA 0.109798f
C1160 two_stage_opamp_dummy_magic_24_0.Vb2.t14 GNDA 0.109798f
C1161 two_stage_opamp_dummy_magic_24_0.Vb2.t18 GNDA 0.109798f
C1162 two_stage_opamp_dummy_magic_24_0.Vb2.t24 GNDA 0.109798f
C1163 two_stage_opamp_dummy_magic_24_0.Vb2.t27 GNDA 0.109798f
C1164 two_stage_opamp_dummy_magic_24_0.Vb2.n14 GNDA 0.361332f
C1165 two_stage_opamp_dummy_magic_24_0.Vb2.n15 GNDA 0.369911f
C1166 two_stage_opamp_dummy_magic_24_0.Vb2.t31 GNDA 0.067192f
C1167 two_stage_opamp_dummy_magic_24_0.Vb2.n16 GNDA 0.257952f
C1168 two_stage_opamp_dummy_magic_24_0.Vb2.t4 GNDA 0.111885f
C1169 two_stage_opamp_dummy_magic_24_0.Vb2.n17 GNDA 0.518097f
C1170 two_stage_opamp_dummy_magic_24_0.Vb2.n18 GNDA 0.12728f
C1171 two_stage_opamp_dummy_magic_24_0.Vb2.t1 GNDA 0.059937f
C1172 two_stage_opamp_dummy_magic_24_0.VD2.t21 GNDA 0.044096f
C1173 two_stage_opamp_dummy_magic_24_0.VD2.t20 GNDA 0.044096f
C1174 two_stage_opamp_dummy_magic_24_0.VD2.n0 GNDA 0.097626f
C1175 two_stage_opamp_dummy_magic_24_0.VD2.n1 GNDA 0.458534f
C1176 two_stage_opamp_dummy_magic_24_0.VD2.n2 GNDA 0.066168f
C1177 two_stage_opamp_dummy_magic_24_0.VD2.n3 GNDA 0.109634f
C1178 two_stage_opamp_dummy_magic_24_0.VD2.t4 GNDA 0.044096f
C1179 two_stage_opamp_dummy_magic_24_0.VD2.t2 GNDA 0.044096f
C1180 two_stage_opamp_dummy_magic_24_0.VD2.n4 GNDA 0.095949f
C1181 two_stage_opamp_dummy_magic_24_0.VD2.n5 GNDA 0.369685f
C1182 two_stage_opamp_dummy_magic_24_0.VD2.n6 GNDA 0.09378f
C1183 two_stage_opamp_dummy_magic_24_0.VD2.t5 GNDA 0.044096f
C1184 two_stage_opamp_dummy_magic_24_0.VD2.t12 GNDA 0.044096f
C1185 two_stage_opamp_dummy_magic_24_0.VD2.n7 GNDA 0.095949f
C1186 two_stage_opamp_dummy_magic_24_0.VD2.n8 GNDA 0.379992f
C1187 two_stage_opamp_dummy_magic_24_0.VD2.t13 GNDA 0.044096f
C1188 two_stage_opamp_dummy_magic_24_0.VD2.t14 GNDA 0.044096f
C1189 two_stage_opamp_dummy_magic_24_0.VD2.n9 GNDA 0.097626f
C1190 two_stage_opamp_dummy_magic_24_0.VD2.t18 GNDA 0.044096f
C1191 two_stage_opamp_dummy_magic_24_0.VD2.t16 GNDA 0.044096f
C1192 two_stage_opamp_dummy_magic_24_0.VD2.n10 GNDA 0.097626f
C1193 two_stage_opamp_dummy_magic_24_0.VD2.n11 GNDA 0.625445f
C1194 two_stage_opamp_dummy_magic_24_0.VD2.t15 GNDA 0.044096f
C1195 two_stage_opamp_dummy_magic_24_0.VD2.t17 GNDA 0.044096f
C1196 two_stage_opamp_dummy_magic_24_0.VD2.n12 GNDA 0.097626f
C1197 two_stage_opamp_dummy_magic_24_0.VD2.n13 GNDA 0.168952f
C1198 two_stage_opamp_dummy_magic_24_0.VD2.t19 GNDA 0.044096f
C1199 two_stage_opamp_dummy_magic_24_0.VD2.t3 GNDA 0.044096f
C1200 two_stage_opamp_dummy_magic_24_0.VD2.n14 GNDA 0.095949f
C1201 two_stage_opamp_dummy_magic_24_0.VD2.n15 GNDA 0.379992f
C1202 two_stage_opamp_dummy_magic_24_0.VD2.n16 GNDA 0.15941f
C1203 two_stage_opamp_dummy_magic_24_0.VD2.t8 GNDA 0.044096f
C1204 two_stage_opamp_dummy_magic_24_0.VD2.t1 GNDA 0.044096f
C1205 two_stage_opamp_dummy_magic_24_0.VD2.n17 GNDA 0.095949f
C1206 two_stage_opamp_dummy_magic_24_0.VD2.n18 GNDA 0.369685f
C1207 two_stage_opamp_dummy_magic_24_0.VD2.n19 GNDA 0.066168f
C1208 two_stage_opamp_dummy_magic_24_0.VD2.n20 GNDA 0.109634f
C1209 two_stage_opamp_dummy_magic_24_0.VD2.n21 GNDA 0.617932f
C1210 two_stage_opamp_dummy_magic_24_0.VD2.n22 GNDA 0.148295f
C1211 two_stage_opamp_dummy_magic_24_0.VD2.n23 GNDA 0.088193f
C1212 two_stage_opamp_dummy_magic_24_0.VD2.t10 GNDA 0.044096f
C1213 two_stage_opamp_dummy_magic_24_0.VD2.t11 GNDA 0.044096f
C1214 two_stage_opamp_dummy_magic_24_0.VD2.n24 GNDA 0.097626f
C1215 two_stage_opamp_dummy_magic_24_0.VD2.n25 GNDA 0.617932f
C1216 two_stage_opamp_dummy_magic_24_0.VD2.n26 GNDA 0.148295f
C1217 two_stage_opamp_dummy_magic_24_0.VD2.n27 GNDA 0.625445f
C1218 two_stage_opamp_dummy_magic_24_0.VD2.n28 GNDA 0.168952f
C1219 two_stage_opamp_dummy_magic_24_0.VD2.n29 GNDA 0.066168f
C1220 two_stage_opamp_dummy_magic_24_0.VD2.t6 GNDA 0.044096f
C1221 two_stage_opamp_dummy_magic_24_0.VD2.t9 GNDA 0.044096f
C1222 two_stage_opamp_dummy_magic_24_0.VD2.n30 GNDA 0.095949f
C1223 two_stage_opamp_dummy_magic_24_0.VD2.n31 GNDA 0.369685f
C1224 two_stage_opamp_dummy_magic_24_0.VD2.n32 GNDA 0.15941f
C1225 two_stage_opamp_dummy_magic_24_0.VD2.n33 GNDA 0.09378f
C1226 two_stage_opamp_dummy_magic_24_0.VD2.t7 GNDA 0.044096f
C1227 two_stage_opamp_dummy_magic_24_0.VD2.t0 GNDA 0.044096f
C1228 two_stage_opamp_dummy_magic_24_0.VD2.n34 GNDA 0.095949f
C1229 two_stage_opamp_dummy_magic_24_0.VD2.n35 GNDA 0.369685f
C1230 two_stage_opamp_dummy_magic_24_0.VD2.n36 GNDA 0.066168f
C1231 two_stage_opamp_dummy_magic_24_0.VD2.n37 GNDA 0.051213f
C1232 two_stage_opamp_dummy_magic_24_0.V_source.n0 GNDA 2.47562f
C1233 two_stage_opamp_dummy_magic_24_0.V_source.n1 GNDA 1.13517f
C1234 two_stage_opamp_dummy_magic_24_0.V_source.n2 GNDA 0.181494f
C1235 two_stage_opamp_dummy_magic_24_0.V_source.n3 GNDA 0.152087f
C1236 two_stage_opamp_dummy_magic_24_0.V_source.n4 GNDA 0.152087f
C1237 two_stage_opamp_dummy_magic_24_0.V_source.n5 GNDA 0.196728f
C1238 two_stage_opamp_dummy_magic_24_0.V_source.n6 GNDA 1.54673f
C1239 two_stage_opamp_dummy_magic_24_0.V_source.n7 GNDA 1.57791f
C1240 two_stage_opamp_dummy_magic_24_0.V_source.n8 GNDA 0.222303f
C1241 two_stage_opamp_dummy_magic_24_0.V_source.t28 GNDA 0.087573f
C1242 two_stage_opamp_dummy_magic_24_0.V_source.n9 GNDA 0.184699f
C1243 two_stage_opamp_dummy_magic_24_0.V_source.t23 GNDA 0.026431f
C1244 two_stage_opamp_dummy_magic_24_0.V_source.t4 GNDA 0.026431f
C1245 two_stage_opamp_dummy_magic_24_0.V_source.n10 GNDA 0.056505f
C1246 two_stage_opamp_dummy_magic_24_0.V_source.t20 GNDA 0.026431f
C1247 two_stage_opamp_dummy_magic_24_0.V_source.t19 GNDA 0.026431f
C1248 two_stage_opamp_dummy_magic_24_0.V_source.n11 GNDA 0.056505f
C1249 two_stage_opamp_dummy_magic_24_0.V_source.n12 GNDA 0.179106f
C1250 two_stage_opamp_dummy_magic_24_0.V_source.t39 GNDA 0.026431f
C1251 two_stage_opamp_dummy_magic_24_0.V_source.t40 GNDA 0.026431f
C1252 two_stage_opamp_dummy_magic_24_0.V_source.n13 GNDA 0.056505f
C1253 two_stage_opamp_dummy_magic_24_0.V_source.n14 GNDA 0.179106f
C1254 two_stage_opamp_dummy_magic_24_0.V_source.t2 GNDA 0.026431f
C1255 two_stage_opamp_dummy_magic_24_0.V_source.t25 GNDA 0.026431f
C1256 two_stage_opamp_dummy_magic_24_0.V_source.n15 GNDA 0.056505f
C1257 two_stage_opamp_dummy_magic_24_0.V_source.n16 GNDA 0.179106f
C1258 two_stage_opamp_dummy_magic_24_0.V_source.n17 GNDA 0.057658f
C1259 two_stage_opamp_dummy_magic_24_0.V_source.t29 GNDA 0.015858f
C1260 two_stage_opamp_dummy_magic_24_0.V_source.t21 GNDA 0.015858f
C1261 two_stage_opamp_dummy_magic_24_0.V_source.n18 GNDA 0.034506f
C1262 two_stage_opamp_dummy_magic_24_0.V_source.n19 GNDA 0.144821f
C1263 two_stage_opamp_dummy_magic_24_0.V_source.t15 GNDA 0.015858f
C1264 two_stage_opamp_dummy_magic_24_0.V_source.t33 GNDA 0.015858f
C1265 two_stage_opamp_dummy_magic_24_0.V_source.n20 GNDA 0.034506f
C1266 two_stage_opamp_dummy_magic_24_0.V_source.n21 GNDA 0.139811f
C1267 two_stage_opamp_dummy_magic_24_0.V_source.t37 GNDA 0.015858f
C1268 two_stage_opamp_dummy_magic_24_0.V_source.t26 GNDA 0.015858f
C1269 two_stage_opamp_dummy_magic_24_0.V_source.n22 GNDA 0.034506f
C1270 two_stage_opamp_dummy_magic_24_0.V_source.n23 GNDA 0.139811f
C1271 two_stage_opamp_dummy_magic_24_0.V_source.n24 GNDA 0.033895f
C1272 two_stage_opamp_dummy_magic_24_0.V_source.n25 GNDA 0.033895f
C1273 two_stage_opamp_dummy_magic_24_0.V_source.t38 GNDA 0.015858f
C1274 two_stage_opamp_dummy_magic_24_0.V_source.t36 GNDA 0.015858f
C1275 two_stage_opamp_dummy_magic_24_0.V_source.n26 GNDA 0.034506f
C1276 two_stage_opamp_dummy_magic_24_0.V_source.n27 GNDA 0.104721f
C1277 two_stage_opamp_dummy_magic_24_0.V_source.t27 GNDA 0.015858f
C1278 two_stage_opamp_dummy_magic_24_0.V_source.t30 GNDA 0.015858f
C1279 two_stage_opamp_dummy_magic_24_0.V_source.n28 GNDA 0.034506f
C1280 two_stage_opamp_dummy_magic_24_0.V_source.n29 GNDA 0.104721f
C1281 two_stage_opamp_dummy_magic_24_0.V_source.n30 GNDA 0.085699f
C1282 two_stage_opamp_dummy_magic_24_0.V_source.t12 GNDA 0.015858f
C1283 two_stage_opamp_dummy_magic_24_0.V_source.t7 GNDA 0.015858f
C1284 two_stage_opamp_dummy_magic_24_0.V_source.n31 GNDA 0.034506f
C1285 two_stage_opamp_dummy_magic_24_0.V_source.n32 GNDA 0.104721f
C1286 two_stage_opamp_dummy_magic_24_0.V_source.n33 GNDA 0.085699f
C1287 two_stage_opamp_dummy_magic_24_0.V_source.t14 GNDA 0.015858f
C1288 two_stage_opamp_dummy_magic_24_0.V_source.t13 GNDA 0.015858f
C1289 two_stage_opamp_dummy_magic_24_0.V_source.n34 GNDA 0.034506f
C1290 two_stage_opamp_dummy_magic_24_0.V_source.n35 GNDA 0.104721f
C1291 two_stage_opamp_dummy_magic_24_0.V_source.n36 GNDA 0.033895f
C1292 two_stage_opamp_dummy_magic_24_0.V_source.t9 GNDA 0.015858f
C1293 two_stage_opamp_dummy_magic_24_0.V_source.t11 GNDA 0.015858f
C1294 two_stage_opamp_dummy_magic_24_0.V_source.n37 GNDA 0.034506f
C1295 two_stage_opamp_dummy_magic_24_0.V_source.n38 GNDA 0.144821f
C1296 two_stage_opamp_dummy_magic_24_0.V_source.t6 GNDA 0.015858f
C1297 two_stage_opamp_dummy_magic_24_0.V_source.t10 GNDA 0.015858f
C1298 two_stage_opamp_dummy_magic_24_0.V_source.n39 GNDA 0.034506f
C1299 two_stage_opamp_dummy_magic_24_0.V_source.n40 GNDA 0.139811f
C1300 two_stage_opamp_dummy_magic_24_0.V_source.n41 GNDA 0.057658f
C1301 two_stage_opamp_dummy_magic_24_0.V_source.n42 GNDA 0.033895f
C1302 two_stage_opamp_dummy_magic_24_0.V_source.t8 GNDA 0.015858f
C1303 two_stage_opamp_dummy_magic_24_0.V_source.t5 GNDA 0.015858f
C1304 two_stage_opamp_dummy_magic_24_0.V_source.n43 GNDA 0.034506f
C1305 two_stage_opamp_dummy_magic_24_0.V_source.n44 GNDA 0.139811f
C1306 two_stage_opamp_dummy_magic_24_0.V_source.n45 GNDA 0.181494f
C1307 two_stage_opamp_dummy_magic_24_0.V_source.t1 GNDA 0.026431f
C1308 two_stage_opamp_dummy_magic_24_0.V_source.t17 GNDA 0.026431f
C1309 two_stage_opamp_dummy_magic_24_0.V_source.n46 GNDA 0.056505f
C1310 two_stage_opamp_dummy_magic_24_0.V_source.n47 GNDA 0.179106f
C1311 two_stage_opamp_dummy_magic_24_0.V_source.t3 GNDA 0.026431f
C1312 two_stage_opamp_dummy_magic_24_0.V_source.t32 GNDA 0.026431f
C1313 two_stage_opamp_dummy_magic_24_0.V_source.n48 GNDA 0.056505f
C1314 two_stage_opamp_dummy_magic_24_0.V_source.t34 GNDA 0.026431f
C1315 two_stage_opamp_dummy_magic_24_0.V_source.t0 GNDA 0.026431f
C1316 two_stage_opamp_dummy_magic_24_0.V_source.n49 GNDA 0.056505f
C1317 two_stage_opamp_dummy_magic_24_0.V_source.n50 GNDA 0.179108f
C1318 two_stage_opamp_dummy_magic_24_0.V_source.t35 GNDA 0.026431f
C1319 two_stage_opamp_dummy_magic_24_0.V_source.t18 GNDA 0.026431f
C1320 two_stage_opamp_dummy_magic_24_0.V_source.n51 GNDA 0.056505f
C1321 two_stage_opamp_dummy_magic_24_0.V_source.n52 GNDA 0.214753f
C1322 two_stage_opamp_dummy_magic_24_0.V_source.t16 GNDA 0.026431f
C1323 two_stage_opamp_dummy_magic_24_0.V_source.t31 GNDA 0.026431f
C1324 two_stage_opamp_dummy_magic_24_0.V_source.n53 GNDA 0.056505f
C1325 two_stage_opamp_dummy_magic_24_0.V_source.n54 GNDA 0.214753f
C1326 two_stage_opamp_dummy_magic_24_0.V_source.t22 GNDA 0.026431f
C1327 two_stage_opamp_dummy_magic_24_0.V_source.t24 GNDA 0.026431f
C1328 two_stage_opamp_dummy_magic_24_0.V_source.n55 GNDA 0.056505f
C1329 two_stage_opamp_dummy_magic_24_0.V_source.n56 GNDA 0.214753f
C1330 two_stage_opamp_dummy_magic_24_0.V_source.n57 GNDA 0.081313f
C1331 two_stage_opamp_dummy_magic_24_0.V_source.n58 GNDA 0.139041f
C1332 two_stage_opamp_dummy_magic_24_0.VD3.t22 GNDA 0.047635f
C1333 two_stage_opamp_dummy_magic_24_0.VD3.n0 GNDA 0.4991f
C1334 two_stage_opamp_dummy_magic_24_0.VD3.t20 GNDA 0.047635f
C1335 two_stage_opamp_dummy_magic_24_0.VD3.t24 GNDA 0.047635f
C1336 two_stage_opamp_dummy_magic_24_0.VD3.n1 GNDA 0.097442f
C1337 two_stage_opamp_dummy_magic_24_0.VD3.n2 GNDA 0.360761f
C1338 two_stage_opamp_dummy_magic_24_0.VD3.n3 GNDA 0.856409f
C1339 two_stage_opamp_dummy_magic_24_0.VD3.t26 GNDA 0.047635f
C1340 two_stage_opamp_dummy_magic_24_0.VD3.t29 GNDA 0.047635f
C1341 two_stage_opamp_dummy_magic_24_0.VD3.n4 GNDA 0.097442f
C1342 two_stage_opamp_dummy_magic_24_0.VD3.n5 GNDA 0.345318f
C1343 two_stage_opamp_dummy_magic_24_0.VD3.n6 GNDA 0.088141f
C1344 two_stage_opamp_dummy_magic_24_0.VD3.n7 GNDA 0.088141f
C1345 two_stage_opamp_dummy_magic_24_0.VD3.t1 GNDA 0.047635f
C1346 two_stage_opamp_dummy_magic_24_0.VD3.t7 GNDA 0.047635f
C1347 two_stage_opamp_dummy_magic_24_0.VD3.n8 GNDA 0.107177f
C1348 two_stage_opamp_dummy_magic_24_0.VD3.n9 GNDA 0.818982f
C1349 two_stage_opamp_dummy_magic_24_0.VD3.t3 GNDA 0.047635f
C1350 two_stage_opamp_dummy_magic_24_0.VD3.t19 GNDA 0.047635f
C1351 two_stage_opamp_dummy_magic_24_0.VD3.n10 GNDA 0.107177f
C1352 two_stage_opamp_dummy_magic_24_0.VD3.n11 GNDA 0.818982f
C1353 two_stage_opamp_dummy_magic_24_0.VD3.t11 GNDA 0.047635f
C1354 two_stage_opamp_dummy_magic_24_0.VD3.t35 GNDA 0.047635f
C1355 two_stage_opamp_dummy_magic_24_0.VD3.n12 GNDA 0.107177f
C1356 two_stage_opamp_dummy_magic_24_0.VD3.n13 GNDA 0.818982f
C1357 two_stage_opamp_dummy_magic_24_0.VD3.t33 GNDA 0.047635f
C1358 two_stage_opamp_dummy_magic_24_0.VD3.t9 GNDA 0.047635f
C1359 two_stage_opamp_dummy_magic_24_0.VD3.n14 GNDA 0.107177f
C1360 two_stage_opamp_dummy_magic_24_0.VD3.n15 GNDA 0.818982f
C1361 two_stage_opamp_dummy_magic_24_0.VD3.t37 GNDA 0.047635f
C1362 two_stage_opamp_dummy_magic_24_0.VD3.t5 GNDA 0.047635f
C1363 two_stage_opamp_dummy_magic_24_0.VD3.n16 GNDA 0.107177f
C1364 two_stage_opamp_dummy_magic_24_0.VD3.n17 GNDA 1.10922f
C1365 two_stage_opamp_dummy_magic_24_0.VD3.t12 GNDA 0.083395f
C1366 two_stage_opamp_dummy_magic_24_0.VD3.n18 GNDA 0.269335f
C1367 two_stage_opamp_dummy_magic_24_0.VD3.t14 GNDA 0.169444f
C1368 two_stage_opamp_dummy_magic_24_0.VD3.n19 GNDA 0.543026f
C1369 two_stage_opamp_dummy_magic_24_0.VD3.t13 GNDA 0.406036f
C1370 two_stage_opamp_dummy_magic_24_0.VD3.t4 GNDA 0.318474f
C1371 two_stage_opamp_dummy_magic_24_0.VD3.t36 GNDA 0.318474f
C1372 two_stage_opamp_dummy_magic_24_0.VD3.t8 GNDA 0.318474f
C1373 two_stage_opamp_dummy_magic_24_0.VD3.t32 GNDA 0.318474f
C1374 two_stage_opamp_dummy_magic_24_0.VD3.t34 GNDA 0.318474f
C1375 two_stage_opamp_dummy_magic_24_0.VD3.t10 GNDA 0.318474f
C1376 two_stage_opamp_dummy_magic_24_0.VD3.t18 GNDA 0.318474f
C1377 two_stage_opamp_dummy_magic_24_0.VD3.t2 GNDA 0.318474f
C1378 two_stage_opamp_dummy_magic_24_0.VD3.t6 GNDA 0.318474f
C1379 two_stage_opamp_dummy_magic_24_0.VD3.t0 GNDA 0.318474f
C1380 two_stage_opamp_dummy_magic_24_0.VD3.t16 GNDA 0.406036f
C1381 two_stage_opamp_dummy_magic_24_0.VD3.t17 GNDA 0.169444f
C1382 two_stage_opamp_dummy_magic_24_0.VD3.n20 GNDA 0.543026f
C1383 two_stage_opamp_dummy_magic_24_0.VD3.t15 GNDA 0.083395f
C1384 two_stage_opamp_dummy_magic_24_0.VD3.n21 GNDA 0.253348f
C1385 two_stage_opamp_dummy_magic_24_0.VD3.n22 GNDA 1.47396f
C1386 two_stage_opamp_dummy_magic_24_0.VD3.t28 GNDA 0.047635f
C1387 two_stage_opamp_dummy_magic_24_0.VD3.t21 GNDA 0.047635f
C1388 two_stage_opamp_dummy_magic_24_0.VD3.n23 GNDA 0.097442f
C1389 two_stage_opamp_dummy_magic_24_0.VD3.n24 GNDA 0.349626f
C1390 two_stage_opamp_dummy_magic_24_0.VD3.n25 GNDA 1.53618f
C1391 two_stage_opamp_dummy_magic_24_0.VD3.t27 GNDA 0.047635f
C1392 two_stage_opamp_dummy_magic_24_0.VD3.t30 GNDA 0.047635f
C1393 two_stage_opamp_dummy_magic_24_0.VD3.n26 GNDA 0.097442f
C1394 two_stage_opamp_dummy_magic_24_0.VD3.n27 GNDA 0.345318f
C1395 two_stage_opamp_dummy_magic_24_0.VD3.n28 GNDA 0.4991f
C1396 two_stage_opamp_dummy_magic_24_0.VD3.n29 GNDA 0.4991f
C1397 two_stage_opamp_dummy_magic_24_0.VD3.t23 GNDA 0.047635f
C1398 two_stage_opamp_dummy_magic_24_0.VD3.t25 GNDA 0.047635f
C1399 two_stage_opamp_dummy_magic_24_0.VD3.n30 GNDA 0.097442f
C1400 two_stage_opamp_dummy_magic_24_0.VD3.n31 GNDA 0.345318f
C1401 two_stage_opamp_dummy_magic_24_0.VD3.n32 GNDA 0.051668f
C1402 two_stage_opamp_dummy_magic_24_0.VD3.n33 GNDA 0.051668f
C1403 two_stage_opamp_dummy_magic_24_0.VD3.n34 GNDA 0.345318f
C1404 two_stage_opamp_dummy_magic_24_0.VD3.n35 GNDA 0.097442f
C1405 two_stage_opamp_dummy_magic_24_0.VD3.t31 GNDA 0.047635f
C1406 two_stage_opamp_dummy_magic_24_0.VD4.t6 GNDA 0.047168f
C1407 two_stage_opamp_dummy_magic_24_0.VD4.n0 GNDA 0.848035f
C1408 two_stage_opamp_dummy_magic_24_0.VD4.n1 GNDA 0.051162f
C1409 two_stage_opamp_dummy_magic_24_0.VD4.t3 GNDA 0.047168f
C1410 two_stage_opamp_dummy_magic_24_0.VD4.t14 GNDA 0.047168f
C1411 two_stage_opamp_dummy_magic_24_0.VD4.n2 GNDA 0.106127f
C1412 two_stage_opamp_dummy_magic_24_0.VD4.n3 GNDA 0.810952f
C1413 two_stage_opamp_dummy_magic_24_0.VD4.t29 GNDA 0.167783f
C1414 two_stage_opamp_dummy_magic_24_0.VD4.t5 GNDA 0.047168f
C1415 two_stage_opamp_dummy_magic_24_0.VD4.t1 GNDA 0.047168f
C1416 two_stage_opamp_dummy_magic_24_0.VD4.n4 GNDA 0.106127f
C1417 two_stage_opamp_dummy_magic_24_0.VD4.n5 GNDA 0.810952f
C1418 two_stage_opamp_dummy_magic_24_0.VD4.t16 GNDA 0.047168f
C1419 two_stage_opamp_dummy_magic_24_0.VD4.t10 GNDA 0.047168f
C1420 two_stage_opamp_dummy_magic_24_0.VD4.n6 GNDA 0.106127f
C1421 two_stage_opamp_dummy_magic_24_0.VD4.n7 GNDA 0.810952f
C1422 two_stage_opamp_dummy_magic_24_0.VD4.t34 GNDA 0.047168f
C1423 two_stage_opamp_dummy_magic_24_0.VD4.t8 GNDA 0.047168f
C1424 two_stage_opamp_dummy_magic_24_0.VD4.n8 GNDA 0.106127f
C1425 two_stage_opamp_dummy_magic_24_0.VD4.n9 GNDA 0.810952f
C1426 two_stage_opamp_dummy_magic_24_0.VD4.t12 GNDA 0.047168f
C1427 two_stage_opamp_dummy_magic_24_0.VD4.t37 GNDA 0.047168f
C1428 two_stage_opamp_dummy_magic_24_0.VD4.n10 GNDA 0.106127f
C1429 two_stage_opamp_dummy_magic_24_0.VD4.n11 GNDA 1.09834f
C1430 two_stage_opamp_dummy_magic_24_0.VD4.t27 GNDA 0.082577f
C1431 two_stage_opamp_dummy_magic_24_0.VD4.n12 GNDA 0.266695f
C1432 two_stage_opamp_dummy_magic_24_0.VD4.n13 GNDA 0.537702f
C1433 two_stage_opamp_dummy_magic_24_0.VD4.t28 GNDA 0.402055f
C1434 two_stage_opamp_dummy_magic_24_0.VD4.t11 GNDA 0.315351f
C1435 two_stage_opamp_dummy_magic_24_0.VD4.t36 GNDA 0.315351f
C1436 two_stage_opamp_dummy_magic_24_0.VD4.t33 GNDA 0.315351f
C1437 two_stage_opamp_dummy_magic_24_0.VD4.t7 GNDA 0.315351f
C1438 two_stage_opamp_dummy_magic_24_0.VD4.t15 GNDA 0.315351f
C1439 two_stage_opamp_dummy_magic_24_0.VD4.t9 GNDA 0.315351f
C1440 two_stage_opamp_dummy_magic_24_0.VD4.t4 GNDA 0.315351f
C1441 two_stage_opamp_dummy_magic_24_0.VD4.t0 GNDA 0.315351f
C1442 two_stage_opamp_dummy_magic_24_0.VD4.t2 GNDA 0.315351f
C1443 two_stage_opamp_dummy_magic_24_0.VD4.t13 GNDA 0.315351f
C1444 two_stage_opamp_dummy_magic_24_0.VD4.t31 GNDA 0.402055f
C1445 two_stage_opamp_dummy_magic_24_0.VD4.t32 GNDA 0.167783f
C1446 two_stage_opamp_dummy_magic_24_0.VD4.n14 GNDA 0.537702f
C1447 two_stage_opamp_dummy_magic_24_0.VD4.t30 GNDA 0.082577f
C1448 two_stage_opamp_dummy_magic_24_0.VD4.n15 GNDA 0.250864f
C1449 two_stage_opamp_dummy_magic_24_0.VD4.n16 GNDA 1.45951f
C1450 two_stage_opamp_dummy_magic_24_0.VD4.n17 GNDA 1.52108f
C1451 two_stage_opamp_dummy_magic_24_0.VD4.t35 GNDA 0.047168f
C1452 two_stage_opamp_dummy_magic_24_0.VD4.t20 GNDA 0.047168f
C1453 two_stage_opamp_dummy_magic_24_0.VD4.n18 GNDA 0.096487f
C1454 two_stage_opamp_dummy_magic_24_0.VD4.n19 GNDA 0.346235f
C1455 two_stage_opamp_dummy_magic_24_0.VD4.n20 GNDA 0.087277f
C1456 two_stage_opamp_dummy_magic_24_0.VD4.t23 GNDA 0.047168f
C1457 two_stage_opamp_dummy_magic_24_0.VD4.t17 GNDA 0.047168f
C1458 two_stage_opamp_dummy_magic_24_0.VD4.n21 GNDA 0.096487f
C1459 two_stage_opamp_dummy_magic_24_0.VD4.n22 GNDA 0.341932f
C1460 two_stage_opamp_dummy_magic_24_0.VD4.n23 GNDA 0.494207f
C1461 two_stage_opamp_dummy_magic_24_0.VD4.t25 GNDA 0.047168f
C1462 two_stage_opamp_dummy_magic_24_0.VD4.t18 GNDA 0.047168f
C1463 two_stage_opamp_dummy_magic_24_0.VD4.n24 GNDA 0.096487f
C1464 two_stage_opamp_dummy_magic_24_0.VD4.n25 GNDA 0.341932f
C1465 two_stage_opamp_dummy_magic_24_0.VD4.n26 GNDA 0.494207f
C1466 two_stage_opamp_dummy_magic_24_0.VD4.n27 GNDA 0.494207f
C1467 two_stage_opamp_dummy_magic_24_0.VD4.t19 GNDA 0.047168f
C1468 two_stage_opamp_dummy_magic_24_0.VD4.t21 GNDA 0.047168f
C1469 two_stage_opamp_dummy_magic_24_0.VD4.n28 GNDA 0.096487f
C1470 two_stage_opamp_dummy_magic_24_0.VD4.n29 GNDA 0.341932f
C1471 two_stage_opamp_dummy_magic_24_0.VD4.n30 GNDA 0.051162f
C1472 two_stage_opamp_dummy_magic_24_0.VD4.t24 GNDA 0.047168f
C1473 two_stage_opamp_dummy_magic_24_0.VD4.t22 GNDA 0.047168f
C1474 two_stage_opamp_dummy_magic_24_0.VD4.n31 GNDA 0.096487f
C1475 two_stage_opamp_dummy_magic_24_0.VD4.n32 GNDA 0.341932f
C1476 two_stage_opamp_dummy_magic_24_0.VD4.n33 GNDA 0.087277f
C1477 two_stage_opamp_dummy_magic_24_0.VD4.n34 GNDA 0.357202f
C1478 two_stage_opamp_dummy_magic_24_0.VD4.n35 GNDA 0.096487f
C1479 two_stage_opamp_dummy_magic_24_0.VD4.t26 GNDA 0.047168f
C1480 two_stage_opamp_dummy_magic_24_0.Vb3.n0 GNDA 0.620039f
C1481 two_stage_opamp_dummy_magic_24_0.Vb3.n1 GNDA 0.687551f
C1482 two_stage_opamp_dummy_magic_24_0.Vb3.n2 GNDA 0.620039f
C1483 two_stage_opamp_dummy_magic_24_0.Vb3.n3 GNDA 0.687551f
C1484 two_stage_opamp_dummy_magic_24_0.Vb3.n4 GNDA 0.764393f
C1485 two_stage_opamp_dummy_magic_24_0.Vb3.n5 GNDA 0.71517f
C1486 two_stage_opamp_dummy_magic_24_0.Vb3.t26 GNDA 0.133081f
C1487 two_stage_opamp_dummy_magic_24_0.Vb3.t22 GNDA 0.133743f
C1488 two_stage_opamp_dummy_magic_24_0.Vb3.t20 GNDA 0.133708f
C1489 two_stage_opamp_dummy_magic_24_0.Vb3.t15 GNDA 0.133708f
C1490 two_stage_opamp_dummy_magic_24_0.Vb3.t9 GNDA 0.133708f
C1491 two_stage_opamp_dummy_magic_24_0.Vb3.t16 GNDA 0.133743f
C1492 two_stage_opamp_dummy_magic_24_0.Vb3.t13 GNDA 0.133708f
C1493 two_stage_opamp_dummy_magic_24_0.Vb3.t19 GNDA 0.133708f
C1494 two_stage_opamp_dummy_magic_24_0.Vb3.t21 GNDA 0.133708f
C1495 two_stage_opamp_dummy_magic_24_0.Vb3.t23 GNDA 0.133081f
C1496 two_stage_opamp_dummy_magic_24_0.Vb3.t27 GNDA 0.133081f
C1497 two_stage_opamp_dummy_magic_24_0.Vb3.t18 GNDA 0.133743f
C1498 two_stage_opamp_dummy_magic_24_0.Vb3.t12 GNDA 0.133708f
C1499 two_stage_opamp_dummy_magic_24_0.Vb3.t28 GNDA 0.133708f
C1500 two_stage_opamp_dummy_magic_24_0.Vb3.t10 GNDA 0.133708f
C1501 two_stage_opamp_dummy_magic_24_0.Vb3.t8 GNDA 0.133743f
C1502 two_stage_opamp_dummy_magic_24_0.Vb3.t14 GNDA 0.133708f
C1503 two_stage_opamp_dummy_magic_24_0.Vb3.t11 GNDA 0.133708f
C1504 two_stage_opamp_dummy_magic_24_0.Vb3.t17 GNDA 0.133708f
C1505 two_stage_opamp_dummy_magic_24_0.Vb3.t25 GNDA 0.133081f
C1506 two_stage_opamp_dummy_magic_24_0.Vb3.t1 GNDA 0.072988f
C1507 two_stage_opamp_dummy_magic_24_0.Vb3.t2 GNDA 0.072988f
C1508 two_stage_opamp_dummy_magic_24_0.Vb3.n6 GNDA 0.201297f
C1509 two_stage_opamp_dummy_magic_24_0.Vb3.t6 GNDA 0.020854f
C1510 two_stage_opamp_dummy_magic_24_0.Vb3.t0 GNDA 0.020854f
C1511 two_stage_opamp_dummy_magic_24_0.Vb3.n7 GNDA 0.067172f
C1512 two_stage_opamp_dummy_magic_24_0.Vb3.t7 GNDA 0.020854f
C1513 two_stage_opamp_dummy_magic_24_0.Vb3.t5 GNDA 0.020854f
C1514 two_stage_opamp_dummy_magic_24_0.Vb3.n8 GNDA 0.067172f
C1515 two_stage_opamp_dummy_magic_24_0.Vb3.n9 GNDA 0.370316f
C1516 two_stage_opamp_dummy_magic_24_0.Vb3.t3 GNDA 0.020854f
C1517 two_stage_opamp_dummy_magic_24_0.Vb3.t4 GNDA 0.020854f
C1518 two_stage_opamp_dummy_magic_24_0.Vb3.n10 GNDA 0.062987f
C1519 two_stage_opamp_dummy_magic_24_0.Vb3.n11 GNDA 1.18209f
C1520 two_stage_opamp_dummy_magic_24_0.Vb3.n12 GNDA 2.08726f
C1521 two_stage_opamp_dummy_magic_24_0.Vb3.t24 GNDA 0.134847f
C1522 two_stage_opamp_dummy_magic_24_0.Vb3.n13 GNDA 0.537965f
C1523 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t42 GNDA 0.412258f
C1524 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t84 GNDA 0.434383f
C1525 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t60 GNDA 0.413752f
C1526 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t65 GNDA 0.412258f
C1527 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t99 GNDA 0.221432f
C1528 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n0 GNDA 0.255706f
C1529 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t88 GNDA 0.412258f
C1530 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t101 GNDA 0.434383f
C1531 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t0 GNDA 0.221432f
C1532 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n1 GNDA 0.235076f
C1533 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t130 GNDA 0.412258f
C1534 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t5 GNDA 0.434383f
C1535 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t35 GNDA 0.221432f
C1536 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n2 GNDA 0.235076f
C1537 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t33 GNDA 0.412258f
C1538 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t127 GNDA 0.434383f
C1539 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t16 GNDA 0.221432f
C1540 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n3 GNDA 0.235076f
C1541 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t12 GNDA 0.412258f
C1542 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t79 GNDA 0.413752f
C1543 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t32 GNDA 0.412258f
C1544 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t73 GNDA 0.413752f
C1545 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t123 GNDA 0.412258f
C1546 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t39 GNDA 0.413752f
C1547 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t17 GNDA 0.412258f
C1548 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t46 GNDA 0.413752f
C1549 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t129 GNDA 0.412258f
C1550 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t75 GNDA 0.413752f
C1551 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t50 GNDA 0.412258f
C1552 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t90 GNDA 0.413752f
C1553 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t24 GNDA 0.412258f
C1554 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t119 GNDA 0.413752f
C1555 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t23 GNDA 0.412258f
C1556 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t52 GNDA 0.413752f
C1557 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t135 GNDA 0.412258f
C1558 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t80 GNDA 0.413752f
C1559 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t58 GNDA 0.412258f
C1560 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t95 GNDA 0.413752f
C1561 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t30 GNDA 0.412258f
C1562 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t125 GNDA 0.413752f
C1563 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t97 GNDA 0.412258f
C1564 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t137 GNDA 0.413752f
C1565 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t66 GNDA 0.412258f
C1566 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t21 GNDA 0.413752f
C1567 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t64 GNDA 0.412258f
C1568 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t98 GNDA 0.413752f
C1569 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t31 GNDA 0.412258f
C1570 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t131 GNDA 0.413752f
C1571 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t107 GNDA 0.412258f
C1572 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t4 GNDA 0.413752f
C1573 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t74 GNDA 0.412258f
C1574 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t28 GNDA 0.413752f
C1575 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t7 GNDA 0.412258f
C1576 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t38 GNDA 0.413752f
C1577 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t117 GNDA 0.412258f
C1578 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t61 GNDA 0.413752f
C1579 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t40 GNDA 0.412258f
C1580 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t82 GNDA 0.413752f
C1581 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t13 GNDA 0.412258f
C1582 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t102 GNDA 0.413752f
C1583 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t11 GNDA 0.412258f
C1584 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t41 GNDA 0.413752f
C1585 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t124 GNDA 0.412258f
C1586 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t69 GNDA 0.413752f
C1587 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t45 GNDA 0.412258f
C1588 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t85 GNDA 0.413752f
C1589 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t19 GNDA 0.412258f
C1590 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t112 GNDA 0.413752f
C1591 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t89 GNDA 0.412258f
C1592 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t133 GNDA 0.413752f
C1593 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t55 GNDA 0.412258f
C1594 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t9 GNDA 0.413752f
C1595 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t51 GNDA 0.412258f
C1596 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t91 GNDA 0.413752f
C1597 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t25 GNDA 0.412258f
C1598 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t120 GNDA 0.413752f
C1599 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t115 GNDA 0.412258f
C1600 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t59 GNDA 0.413752f
C1601 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t108 GNDA 0.412258f
C1602 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t43 GNDA 0.413752f
C1603 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t105 GNDA 0.412258f
C1604 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t2 GNDA 0.413752f
C1605 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t72 GNDA 0.412258f
C1606 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t26 GNDA 0.413752f
C1607 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t1 GNDA 0.412258f
C1608 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t34 GNDA 0.413752f
C1609 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t109 GNDA 0.412258f
C1610 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t56 GNDA 0.413752f
C1611 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t44 GNDA 0.412258f
C1612 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t87 GNDA 0.432471f
C1613 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t86 GNDA 0.412258f
C1614 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t134 GNDA 0.221432f
C1615 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n4 GNDA 0.236987f
C1616 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t62 GNDA 0.412258f
C1617 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t103 GNDA 0.221432f
C1618 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n5 GNDA 0.235076f
C1619 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t100 GNDA 0.412258f
C1620 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t6 GNDA 0.221432f
C1621 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n6 GNDA 0.235076f
C1622 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t3 GNDA 0.412258f
C1623 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t37 GNDA 0.221432f
C1624 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n7 GNDA 0.235076f
C1625 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t36 GNDA 0.412258f
C1626 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t78 GNDA 0.221432f
C1627 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n8 GNDA 0.235076f
C1628 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t18 GNDA 0.412258f
C1629 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t54 GNDA 0.221432f
C1630 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n9 GNDA 0.235076f
C1631 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t49 GNDA 0.412258f
C1632 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t94 GNDA 0.221432f
C1633 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n10 GNDA 0.235076f
C1634 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t93 GNDA 0.412258f
C1635 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t136 GNDA 0.221432f
C1636 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n11 GNDA 0.235076f
C1637 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t71 GNDA 0.412258f
C1638 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t114 GNDA 0.221432f
C1639 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n12 GNDA 0.235076f
C1640 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t111 GNDA 0.412258f
C1641 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t8 GNDA 0.221432f
C1642 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n13 GNDA 0.235076f
C1643 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t47 GNDA 0.412258f
C1644 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t128 GNDA 0.413752f
C1645 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t14 GNDA 0.412258f
C1646 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t83 GNDA 0.413752f
C1647 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t118 GNDA 0.199307f
C1648 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n14 GNDA 0.257077f
C1649 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t15 GNDA 0.220062f
C1650 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n15 GNDA 0.279201f
C1651 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t57 GNDA 0.220062f
C1652 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n16 GNDA 0.299832f
C1653 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t27 GNDA 0.220062f
C1654 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n17 GNDA 0.299832f
C1655 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t96 GNDA 0.220062f
C1656 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n18 GNDA 0.299832f
C1657 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t122 GNDA 0.220062f
C1658 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n19 GNDA 0.299832f
C1659 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t10 GNDA 0.220062f
C1660 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n20 GNDA 0.299832f
C1661 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t113 GNDA 0.220062f
C1662 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n21 GNDA 0.299832f
C1663 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t70 GNDA 0.220062f
C1664 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n22 GNDA 0.299832f
C1665 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t106 GNDA 0.220062f
C1666 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n23 GNDA 0.299832f
C1667 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t63 GNDA 0.220062f
C1668 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n24 GNDA 0.299832f
C1669 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t29 GNDA 0.220062f
C1670 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n25 GNDA 0.299832f
C1671 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t132 GNDA 0.220062f
C1672 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n26 GNDA 0.299832f
C1673 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t22 GNDA 0.220062f
C1674 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n27 GNDA 0.299832f
C1675 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t126 GNDA 0.220062f
C1676 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n28 GNDA 0.299832f
C1677 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t81 GNDA 0.220062f
C1678 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n29 GNDA 0.299832f
C1679 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t121 GNDA 0.220062f
C1680 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n30 GNDA 0.299832f
C1681 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t76 GNDA 0.220062f
C1682 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n31 GNDA 0.299832f
C1683 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t77 GNDA 0.220062f
C1684 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n32 GNDA 0.299832f
C1685 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t116 GNDA 0.220062f
C1686 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n33 GNDA 0.276337f
C1687 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t110 GNDA 0.413752f
C1688 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t67 GNDA 0.413752f
C1689 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t104 GNDA 0.412258f
C1690 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t53 GNDA 0.434383f
C1691 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t92 GNDA 0.221432f
C1692 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n34 GNDA 0.255706f
C1693 two_stage_opamp_dummy_magic_24_0.cap_res_Y.n35 GNDA 0.235076f
C1694 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t48 GNDA 0.221432f
C1695 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t20 GNDA 0.434383f
C1696 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t68 GNDA 0.590705f
C1697 two_stage_opamp_dummy_magic_24_0.cap_res_Y.t138 GNDA 0.355571f
C1698 VOUT+.n0 GNDA 0.037005f
C1699 VOUT+.t13 GNDA 0.053966f
C1700 VOUT+.t3 GNDA 0.053966f
C1701 VOUT+.n1 GNDA 0.115952f
C1702 VOUT+.n2 GNDA 0.284645f
C1703 VOUT+.n3 GNDA 0.037005f
C1704 VOUT+.n4 GNDA 0.245519f
C1705 VOUT+.t8 GNDA 0.053966f
C1706 VOUT+.t14 GNDA 0.053966f
C1707 VOUT+.n5 GNDA 0.115952f
C1708 VOUT+.n6 GNDA 0.29362f
C1709 VOUT+.n7 GNDA 0.164964f
C1710 VOUT+.t10 GNDA 0.053966f
C1711 VOUT+.t9 GNDA 0.053966f
C1712 VOUT+.n8 GNDA 0.115952f
C1713 VOUT+.n9 GNDA 0.279953f
C1714 VOUT+.n10 GNDA 0.131606f
C1715 VOUT+.n11 GNDA 0.037005f
C1716 VOUT+.n12 GNDA 0.190951f
C1717 VOUT+.n13 GNDA 0.037005f
C1718 VOUT+.n14 GNDA 0.037005f
C1719 VOUT+.n15 GNDA 0.037005f
C1720 VOUT+.n16 GNDA 0.037005f
C1721 VOUT+.n17 GNDA 0.084996f
C1722 VOUT+.n18 GNDA 0.099452f
C1723 VOUT+.n19 GNDA 0.077094f
C1724 VOUT+.n22 GNDA 0.039318f
C1725 VOUT+.n24 GNDA 0.039318f
C1726 VOUT+.n27 GNDA 0.057821f
C1727 VOUT+.n28 GNDA 0.096368f
C1728 VOUT+.n29 GNDA 0.061259f
C1729 VOUT+.n30 GNDA 0.057821f
C1730 VOUT+.n32 GNDA 0.039318f
C1731 VOUT+.n33 GNDA 0.036659f
C1732 VOUT+.n34 GNDA 0.039318f
C1733 VOUT+.n35 GNDA 0.050882f
C1734 VOUT+.n36 GNDA 0.073411f
C1735 VOUT+.n37 GNDA 0.071441f
C1736 VOUT+.n38 GNDA 0.050882f
C1737 VOUT+.n39 GNDA 0.050882f
C1738 VOUT+.n40 GNDA 0.071441f
C1739 VOUT+.n41 GNDA 0.071441f
C1740 VOUT+.n42 GNDA 0.050882f
C1741 VOUT+.n43 GNDA 0.081459f
C1742 VOUT+.t11 GNDA 0.046257f
C1743 VOUT+.t0 GNDA 0.046257f
C1744 VOUT+.n44 GNDA 0.09478f
C1745 VOUT+.n45 GNDA 0.244654f
C1746 VOUT+.t4 GNDA 0.046257f
C1747 VOUT+.t12 GNDA 0.046257f
C1748 VOUT+.n46 GNDA 0.09478f
C1749 VOUT+.n47 GNDA 0.244654f
C1750 VOUT+.t16 GNDA 0.046257f
C1751 VOUT+.t7 GNDA 0.046257f
C1752 VOUT+.n48 GNDA 0.09478f
C1753 VOUT+.n49 GNDA 0.242189f
C1754 VOUT+.n50 GNDA 0.05882f
C1755 VOUT+.t1 GNDA 0.046257f
C1756 VOUT+.t5 GNDA 0.046257f
C1757 VOUT+.n51 GNDA 0.09478f
C1758 VOUT+.n52 GNDA 0.242189f
C1759 VOUT+.n53 GNDA 0.033341f
C1760 VOUT+.t6 GNDA 0.046257f
C1761 VOUT+.t17 GNDA 0.046257f
C1762 VOUT+.n54 GNDA 0.09478f
C1763 VOUT+.n55 GNDA 0.242189f
C1764 VOUT+.n56 GNDA 0.033341f
C1765 VOUT+.n57 GNDA 0.05882f
C1766 VOUT+.t15 GNDA 0.046257f
C1767 VOUT+.t18 GNDA 0.046257f
C1768 VOUT+.n58 GNDA 0.09478f
C1769 VOUT+.n59 GNDA 0.242189f
C1770 VOUT+.n60 GNDA 0.03889f
C1771 VOUT+.n61 GNDA 0.023128f
C1772 VOUT+.n62 GNDA 0.023128f
C1773 VOUT+.n63 GNDA 0.03889f
C1774 VOUT+.n64 GNDA 0.071441f
C1775 VOUT+.n65 GNDA 0.100003f
C1776 VOUT+.n66 GNDA 0.124608f
C1777 VOUT+.n67 GNDA 0.1744f
C1778 VOUT+.n68 GNDA 0.050882f
C1779 VOUT+.n69 GNDA 0.083262f
C1780 VOUT+.n70 GNDA 0.050882f
C1781 VOUT+.n71 GNDA 0.083262f
C1782 VOUT+.n72 GNDA 0.050882f
C1783 VOUT+.n73 GNDA 0.050882f
C1784 VOUT+.n74 GNDA 0.050882f
C1785 VOUT+.n75 GNDA 0.083262f
C1786 VOUT+.n76 GNDA 0.050882f
C1787 VOUT+.n77 GNDA 0.076323f
C1788 VOUT+.n78 GNDA 0.24516f
C1789 VOUT+.n80 GNDA 0.077094f
C1790 VOUT+.n81 GNDA 0.039318f
C1791 VOUT+.n83 GNDA 0.039318f
C1792 VOUT+.n86 GNDA 0.077094f
C1793 VOUT+.n87 GNDA 0.238221f
C1794 VOUT+.n88 GNDA 0.549297f
C1795 VOUT+.n91 GNDA 0.057821f
C1796 VOUT+.n92 GNDA 0.057821f
C1797 VOUT+.n93 GNDA 0.057821f
C1798 VOUT+.n94 GNDA 0.057821f
C1799 VOUT+.n95 GNDA 0.169598f
C1800 VOUT+.n96 GNDA 0.057821f
C1801 VOUT+.t38 GNDA 0.308377f
C1802 VOUT+.t142 GNDA 0.31363f
C1803 VOUT+.t73 GNDA 0.308377f
C1804 VOUT+.n97 GNDA 0.206757f
C1805 VOUT+.n98 GNDA 0.134915f
C1806 VOUT+.t45 GNDA 0.312972f
C1807 VOUT+.t85 GNDA 0.312972f
C1808 VOUT+.t63 GNDA 0.312972f
C1809 VOUT+.t107 GNDA 0.312972f
C1810 VOUT+.t138 GNDA 0.312972f
C1811 VOUT+.t120 GNDA 0.312972f
C1812 VOUT+.t153 GNDA 0.312972f
C1813 VOUT+.t56 GNDA 0.312972f
C1814 VOUT+.t94 GNDA 0.312972f
C1815 VOUT+.t70 GNDA 0.312972f
C1816 VOUT+.t112 GNDA 0.312972f
C1817 VOUT+.t69 GNDA 0.308377f
C1818 VOUT+.n99 GNDA 0.207415f
C1819 VOUT+.t22 GNDA 0.308377f
C1820 VOUT+.n100 GNDA 0.265235f
C1821 VOUT+.t53 GNDA 0.308377f
C1822 VOUT+.n101 GNDA 0.265235f
C1823 VOUT+.t150 GNDA 0.308377f
C1824 VOUT+.n102 GNDA 0.265235f
C1825 VOUT+.t119 GNDA 0.308377f
C1826 VOUT+.n103 GNDA 0.265235f
C1827 VOUT+.t78 GNDA 0.308377f
C1828 VOUT+.n104 GNDA 0.265235f
C1829 VOUT+.t102 GNDA 0.308377f
C1830 VOUT+.n105 GNDA 0.265235f
C1831 VOUT+.t62 GNDA 0.308377f
C1832 VOUT+.n106 GNDA 0.265235f
C1833 VOUT+.t20 GNDA 0.308377f
C1834 VOUT+.n107 GNDA 0.265235f
C1835 VOUT+.t42 GNDA 0.308377f
C1836 VOUT+.n108 GNDA 0.265235f
C1837 VOUT+.t148 GNDA 0.308377f
C1838 VOUT+.n109 GNDA 0.265235f
C1839 VOUT+.t141 GNDA 0.308377f
C1840 VOUT+.t109 GNDA 0.31363f
C1841 VOUT+.t28 GNDA 0.308377f
C1842 VOUT+.n110 GNDA 0.206757f
C1843 VOUT+.n111 GNDA 0.250556f
C1844 VOUT+.t155 GNDA 0.31363f
C1845 VOUT+.t122 GNDA 0.308377f
C1846 VOUT+.n112 GNDA 0.206757f
C1847 VOUT+.t99 GNDA 0.308377f
C1848 VOUT+.t47 GNDA 0.31363f
C1849 VOUT+.t100 GNDA 0.308377f
C1850 VOUT+.n113 GNDA 0.206757f
C1851 VOUT+.n114 GNDA 0.250556f
C1852 VOUT+.t51 GNDA 0.31363f
C1853 VOUT+.t154 GNDA 0.308377f
C1854 VOUT+.n115 GNDA 0.206757f
C1855 VOUT+.t129 GNDA 0.308377f
C1856 VOUT+.t84 GNDA 0.31363f
C1857 VOUT+.t130 GNDA 0.308377f
C1858 VOUT+.n116 GNDA 0.206757f
C1859 VOUT+.n117 GNDA 0.250556f
C1860 VOUT+.t41 GNDA 0.31363f
C1861 VOUT+.t97 GNDA 0.308377f
C1862 VOUT+.n118 GNDA 0.206757f
C1863 VOUT+.t60 GNDA 0.308377f
C1864 VOUT+.t48 GNDA 0.31363f
C1865 VOUT+.t113 GNDA 0.308377f
C1866 VOUT+.n119 GNDA 0.206757f
C1867 VOUT+.n120 GNDA 0.250556f
C1868 VOUT+.t105 GNDA 0.31363f
C1869 VOUT+.t65 GNDA 0.308377f
C1870 VOUT+.n121 GNDA 0.206757f
C1871 VOUT+.t34 GNDA 0.308377f
C1872 VOUT+.t131 GNDA 0.31363f
C1873 VOUT+.t36 GNDA 0.308377f
C1874 VOUT+.n122 GNDA 0.206757f
C1875 VOUT+.n123 GNDA 0.250556f
C1876 VOUT+.t67 GNDA 0.31363f
C1877 VOUT+.t23 GNDA 0.308377f
C1878 VOUT+.n124 GNDA 0.206757f
C1879 VOUT+.t146 GNDA 0.308377f
C1880 VOUT+.t101 GNDA 0.31363f
C1881 VOUT+.t147 GNDA 0.308377f
C1882 VOUT+.n125 GNDA 0.206757f
C1883 VOUT+.n126 GNDA 0.250556f
C1884 VOUT+.t111 GNDA 0.31363f
C1885 VOUT+.t71 GNDA 0.308377f
C1886 VOUT+.n127 GNDA 0.206757f
C1887 VOUT+.t43 GNDA 0.308377f
C1888 VOUT+.t137 GNDA 0.31363f
C1889 VOUT+.t44 GNDA 0.308377f
C1890 VOUT+.n128 GNDA 0.206757f
C1891 VOUT+.n129 GNDA 0.250556f
C1892 VOUT+.t52 GNDA 0.31363f
C1893 VOUT+.t103 GNDA 0.308377f
C1894 VOUT+.n130 GNDA 0.201938f
C1895 VOUT+.t88 GNDA 0.31363f
C1896 VOUT+.t136 GNDA 0.308377f
C1897 VOUT+.n131 GNDA 0.201938f
C1898 VOUT+.t123 GNDA 0.31363f
C1899 VOUT+.t29 GNDA 0.308377f
C1900 VOUT+.n132 GNDA 0.201938f
C1901 VOUT+.t26 GNDA 0.31363f
C1902 VOUT+.t151 GNDA 0.308377f
C1903 VOUT+.n133 GNDA 0.201938f
C1904 VOUT+.t68 GNDA 0.31363f
C1905 VOUT+.t55 GNDA 0.308377f
C1906 VOUT+.n134 GNDA 0.203866f
C1907 VOUT+.t91 GNDA 0.31323f
C1908 VOUT+.t114 GNDA 0.31363f
C1909 VOUT+.t72 GNDA 0.308377f
C1910 VOUT+.n135 GNDA 0.206757f
C1911 VOUT+.t96 GNDA 0.308377f
C1912 VOUT+.n136 GNDA 0.134915f
C1913 VOUT+.t57 GNDA 0.308377f
C1914 VOUT+.n137 GNDA 0.268832f
C1915 VOUT+.t156 GNDA 0.308377f
C1916 VOUT+.n138 GNDA 0.199481f
C1917 VOUT+.t121 GNDA 0.308377f
C1918 VOUT+.n139 GNDA 0.197554f
C1919 VOUT+.t140 GNDA 0.308377f
C1920 VOUT+.n140 GNDA 0.197554f
C1921 VOUT+.t108 GNDA 0.308377f
C1922 VOUT+.n141 GNDA 0.197554f
C1923 VOUT+.t64 GNDA 0.308377f
C1924 VOUT+.n142 GNDA 0.197554f
C1925 VOUT+.t89 GNDA 0.308377f
C1926 VOUT+.n143 GNDA 0.134915f
C1927 VOUT+.t46 GNDA 0.308377f
C1928 VOUT+.n144 GNDA 0.134915f
C1929 VOUT+.t40 GNDA 0.308377f
C1930 VOUT+.t144 GNDA 0.31363f
C1931 VOUT+.t77 GNDA 0.308377f
C1932 VOUT+.n145 GNDA 0.206757f
C1933 VOUT+.n146 GNDA 0.192736f
C1934 VOUT+.t124 GNDA 0.31363f
C1935 VOUT+.t83 GNDA 0.308377f
C1936 VOUT+.n147 GNDA 0.206757f
C1937 VOUT+.t79 GNDA 0.308377f
C1938 VOUT+.t33 GNDA 0.31363f
C1939 VOUT+.t117 GNDA 0.308377f
C1940 VOUT+.n148 GNDA 0.206757f
C1941 VOUT+.n149 GNDA 0.250556f
C1942 VOUT+.t139 GNDA 0.31363f
C1943 VOUT+.t110 GNDA 0.308377f
C1944 VOUT+.n150 GNDA 0.206757f
C1945 VOUT+.t80 GNDA 0.308377f
C1946 VOUT+.t27 GNDA 0.31363f
C1947 VOUT+.t81 GNDA 0.308377f
C1948 VOUT+.n151 GNDA 0.206757f
C1949 VOUT+.n152 GNDA 0.250556f
C1950 VOUT+.t106 GNDA 0.31363f
C1951 VOUT+.t66 GNDA 0.308377f
C1952 VOUT+.n153 GNDA 0.206757f
C1953 VOUT+.t35 GNDA 0.308377f
C1954 VOUT+.t132 GNDA 0.31363f
C1955 VOUT+.t37 GNDA 0.308377f
C1956 VOUT+.n154 GNDA 0.206757f
C1957 VOUT+.n155 GNDA 0.250556f
C1958 VOUT+.t133 GNDA 0.31363f
C1959 VOUT+.t104 GNDA 0.308377f
C1960 VOUT+.n156 GNDA 0.206757f
C1961 VOUT+.t75 GNDA 0.308377f
C1962 VOUT+.t21 GNDA 0.31363f
C1963 VOUT+.t76 GNDA 0.308377f
C1964 VOUT+.n157 GNDA 0.206757f
C1965 VOUT+.n158 GNDA 0.250556f
C1966 VOUT+.t98 GNDA 0.31363f
C1967 VOUT+.t61 GNDA 0.308377f
C1968 VOUT+.n159 GNDA 0.206757f
C1969 VOUT+.t30 GNDA 0.308377f
C1970 VOUT+.t126 GNDA 0.31363f
C1971 VOUT+.t31 GNDA 0.308377f
C1972 VOUT+.n160 GNDA 0.206757f
C1973 VOUT+.n161 GNDA 0.250556f
C1974 VOUT+.t59 GNDA 0.31363f
C1975 VOUT+.t19 GNDA 0.308377f
C1976 VOUT+.n162 GNDA 0.206757f
C1977 VOUT+.t134 GNDA 0.308377f
C1978 VOUT+.t90 GNDA 0.31363f
C1979 VOUT+.t135 GNDA 0.308377f
C1980 VOUT+.n163 GNDA 0.206757f
C1981 VOUT+.n164 GNDA 0.250556f
C1982 VOUT+.t92 GNDA 0.31363f
C1983 VOUT+.t58 GNDA 0.308377f
C1984 VOUT+.n165 GNDA 0.206757f
C1985 VOUT+.t24 GNDA 0.308377f
C1986 VOUT+.t125 GNDA 0.31363f
C1987 VOUT+.t25 GNDA 0.308377f
C1988 VOUT+.n166 GNDA 0.206757f
C1989 VOUT+.n167 GNDA 0.250556f
C1990 VOUT+.t49 GNDA 0.31363f
C1991 VOUT+.t152 GNDA 0.308377f
C1992 VOUT+.n168 GNDA 0.206757f
C1993 VOUT+.t127 GNDA 0.308377f
C1994 VOUT+.t82 GNDA 0.31363f
C1995 VOUT+.t128 GNDA 0.308377f
C1996 VOUT+.n169 GNDA 0.206757f
C1997 VOUT+.n170 GNDA 0.250556f
C1998 VOUT+.t149 GNDA 0.31363f
C1999 VOUT+.t118 GNDA 0.308377f
C2000 VOUT+.n171 GNDA 0.206757f
C2001 VOUT+.t93 GNDA 0.308377f
C2002 VOUT+.t39 GNDA 0.31363f
C2003 VOUT+.t95 GNDA 0.308377f
C2004 VOUT+.n172 GNDA 0.206757f
C2005 VOUT+.n173 GNDA 0.250556f
C2006 VOUT+.t116 GNDA 0.31363f
C2007 VOUT+.t74 GNDA 0.308377f
C2008 VOUT+.n174 GNDA 0.206757f
C2009 VOUT+.t50 GNDA 0.308377f
C2010 VOUT+.t143 GNDA 0.31363f
C2011 VOUT+.t54 GNDA 0.308377f
C2012 VOUT+.n175 GNDA 0.206757f
C2013 VOUT+.n176 GNDA 0.250556f
C2014 VOUT+.t32 GNDA 0.31363f
C2015 VOUT+.t87 GNDA 0.308377f
C2016 VOUT+.n177 GNDA 0.206757f
C2017 VOUT+.t86 GNDA 0.308377f
C2018 VOUT+.n178 GNDA 0.250556f
C2019 VOUT+.t115 GNDA 0.308377f
C2020 VOUT+.n179 GNDA 0.132024f
C2021 VOUT+.t145 GNDA 0.308377f
C2022 VOUT+.n180 GNDA 0.344033f
C2023 VOUT+.n181 GNDA 0.283322f
C2024 VOUT+.n182 GNDA 0.057821f
C2025 VOUT+.n183 GNDA 0.057821f
C2026 VOUT+.n185 GNDA 0.558934f
C2027 VOUT+.n186 GNDA 0.058247f
C2028 VOUT+.n187 GNDA 1.09859f
C2029 VOUT+.n188 GNDA 0.039318f
C2030 VOUT+.n190 GNDA 0.037005f
C2031 VOUT+.n191 GNDA 1.08896f
C2032 VOUT+.n193 GNDA 0.039318f
C2033 VOUT+.n194 GNDA 0.077094f
C2034 VOUT+.n195 GNDA 0.104077f
C2035 VOUT+.t2 GNDA 0.088338f
C2036 VOUT+.n196 GNDA 0.271885f
C2037 two_stage_opamp_dummy_magic_24_0.cap_res_X.t57 GNDA 0.412258f
C2038 two_stage_opamp_dummy_magic_24_0.cap_res_X.t93 GNDA 0.413752f
C2039 two_stage_opamp_dummy_magic_24_0.cap_res_X.t25 GNDA 0.412258f
C2040 two_stage_opamp_dummy_magic_24_0.cap_res_X.t62 GNDA 0.413752f
C2041 two_stage_opamp_dummy_magic_24_0.cap_res_X.t115 GNDA 0.412258f
C2042 two_stage_opamp_dummy_magic_24_0.cap_res_X.t79 GNDA 0.413752f
C2043 two_stage_opamp_dummy_magic_24_0.cap_res_X.t54 GNDA 0.412258f
C2044 two_stage_opamp_dummy_magic_24_0.cap_res_X.t88 GNDA 0.413752f
C2045 two_stage_opamp_dummy_magic_24_0.cap_res_X.t71 GNDA 0.412258f
C2046 two_stage_opamp_dummy_magic_24_0.cap_res_X.t37 GNDA 0.413752f
C2047 two_stage_opamp_dummy_magic_24_0.cap_res_X.t90 GNDA 0.412258f
C2048 two_stage_opamp_dummy_magic_24_0.cap_res_X.t130 GNDA 0.413752f
C2049 two_stage_opamp_dummy_magic_24_0.cap_res_X.t109 GNDA 0.412258f
C2050 two_stage_opamp_dummy_magic_24_0.cap_res_X.t75 GNDA 0.413752f
C2051 two_stage_opamp_dummy_magic_24_0.cap_res_X.t59 GNDA 0.412258f
C2052 two_stage_opamp_dummy_magic_24_0.cap_res_X.t92 GNDA 0.413752f
C2053 two_stage_opamp_dummy_magic_24_0.cap_res_X.t77 GNDA 0.412258f
C2054 two_stage_opamp_dummy_magic_24_0.cap_res_X.t44 GNDA 0.413752f
C2055 two_stage_opamp_dummy_magic_24_0.cap_res_X.t96 GNDA 0.412258f
C2056 two_stage_opamp_dummy_magic_24_0.cap_res_X.t133 GNDA 0.413752f
C2057 two_stage_opamp_dummy_magic_24_0.cap_res_X.t114 GNDA 0.412258f
C2058 two_stage_opamp_dummy_magic_24_0.cap_res_X.t81 GNDA 0.413752f
C2059 two_stage_opamp_dummy_magic_24_0.cap_res_X.t138 GNDA 0.412258f
C2060 two_stage_opamp_dummy_magic_24_0.cap_res_X.t34 GNDA 0.413752f
C2061 two_stage_opamp_dummy_magic_24_0.cap_res_X.t15 GNDA 0.412258f
C2062 two_stage_opamp_dummy_magic_24_0.cap_res_X.t120 GNDA 0.413752f
C2063 two_stage_opamp_dummy_magic_24_0.cap_res_X.t102 GNDA 0.412258f
C2064 two_stage_opamp_dummy_magic_24_0.cap_res_X.t1 GNDA 0.413752f
C2065 two_stage_opamp_dummy_magic_24_0.cap_res_X.t121 GNDA 0.412258f
C2066 two_stage_opamp_dummy_magic_24_0.cap_res_X.t85 GNDA 0.413752f
C2067 two_stage_opamp_dummy_magic_24_0.cap_res_X.t6 GNDA 0.412258f
C2068 two_stage_opamp_dummy_magic_24_0.cap_res_X.t42 GNDA 0.413752f
C2069 two_stage_opamp_dummy_magic_24_0.cap_res_X.t23 GNDA 0.412258f
C2070 two_stage_opamp_dummy_magic_24_0.cap_res_X.t126 GNDA 0.413752f
C2071 two_stage_opamp_dummy_magic_24_0.cap_res_X.t46 GNDA 0.412258f
C2072 two_stage_opamp_dummy_magic_24_0.cap_res_X.t80 GNDA 0.413752f
C2073 two_stage_opamp_dummy_magic_24_0.cap_res_X.t60 GNDA 0.412258f
C2074 two_stage_opamp_dummy_magic_24_0.cap_res_X.t28 GNDA 0.413752f
C2075 two_stage_opamp_dummy_magic_24_0.cap_res_X.t83 GNDA 0.412258f
C2076 two_stage_opamp_dummy_magic_24_0.cap_res_X.t117 GNDA 0.413752f
C2077 two_stage_opamp_dummy_magic_24_0.cap_res_X.t98 GNDA 0.412258f
C2078 two_stage_opamp_dummy_magic_24_0.cap_res_X.t64 GNDA 0.413752f
C2079 two_stage_opamp_dummy_magic_24_0.cap_res_X.t49 GNDA 0.412258f
C2080 two_stage_opamp_dummy_magic_24_0.cap_res_X.t84 GNDA 0.413752f
C2081 two_stage_opamp_dummy_magic_24_0.cap_res_X.t65 GNDA 0.412258f
C2082 two_stage_opamp_dummy_magic_24_0.cap_res_X.t33 GNDA 0.413752f
C2083 two_stage_opamp_dummy_magic_24_0.cap_res_X.t87 GNDA 0.412258f
C2084 two_stage_opamp_dummy_magic_24_0.cap_res_X.t123 GNDA 0.413752f
C2085 two_stage_opamp_dummy_magic_24_0.cap_res_X.t104 GNDA 0.412258f
C2086 two_stage_opamp_dummy_magic_24_0.cap_res_X.t70 GNDA 0.413752f
C2087 two_stage_opamp_dummy_magic_24_0.cap_res_X.t128 GNDA 0.412258f
C2088 two_stage_opamp_dummy_magic_24_0.cap_res_X.t24 GNDA 0.413752f
C2089 two_stage_opamp_dummy_magic_24_0.cap_res_X.t7 GNDA 0.412258f
C2090 two_stage_opamp_dummy_magic_24_0.cap_res_X.t108 GNDA 0.413752f
C2091 two_stage_opamp_dummy_magic_24_0.cap_res_X.t91 GNDA 0.412258f
C2092 two_stage_opamp_dummy_magic_24_0.cap_res_X.t129 GNDA 0.413752f
C2093 two_stage_opamp_dummy_magic_24_0.cap_res_X.t110 GNDA 0.412258f
C2094 two_stage_opamp_dummy_magic_24_0.cap_res_X.t76 GNDA 0.413752f
C2095 two_stage_opamp_dummy_magic_24_0.cap_res_X.t95 GNDA 0.412258f
C2096 two_stage_opamp_dummy_magic_24_0.cap_res_X.t47 GNDA 0.413752f
C2097 two_stage_opamp_dummy_magic_24_0.cap_res_X.t127 GNDA 0.412258f
C2098 two_stage_opamp_dummy_magic_24_0.cap_res_X.t43 GNDA 0.413752f
C2099 two_stage_opamp_dummy_magic_24_0.cap_res_X.t4 GNDA 0.412258f
C2100 two_stage_opamp_dummy_magic_24_0.cap_res_X.t41 GNDA 0.413752f
C2101 two_stage_opamp_dummy_magic_24_0.cap_res_X.t21 GNDA 0.412258f
C2102 two_stage_opamp_dummy_magic_24_0.cap_res_X.t124 GNDA 0.413752f
C2103 two_stage_opamp_dummy_magic_24_0.cap_res_X.t40 GNDA 0.412258f
C2104 two_stage_opamp_dummy_magic_24_0.cap_res_X.t72 GNDA 0.413752f
C2105 two_stage_opamp_dummy_magic_24_0.cap_res_X.t55 GNDA 0.412258f
C2106 two_stage_opamp_dummy_magic_24_0.cap_res_X.t20 GNDA 0.413752f
C2107 two_stage_opamp_dummy_magic_24_0.cap_res_X.t99 GNDA 0.412258f
C2108 two_stage_opamp_dummy_magic_24_0.cap_res_X.t137 GNDA 0.413752f
C2109 two_stage_opamp_dummy_magic_24_0.cap_res_X.t11 GNDA 0.412258f
C2110 two_stage_opamp_dummy_magic_24_0.cap_res_X.t53 GNDA 0.432471f
C2111 two_stage_opamp_dummy_magic_24_0.cap_res_X.t38 GNDA 0.412258f
C2112 two_stage_opamp_dummy_magic_24_0.cap_res_X.t78 GNDA 0.221432f
C2113 two_stage_opamp_dummy_magic_24_0.cap_res_X.n0 GNDA 0.236987f
C2114 two_stage_opamp_dummy_magic_24_0.cap_res_X.t18 GNDA 0.412258f
C2115 two_stage_opamp_dummy_magic_24_0.cap_res_X.t56 GNDA 0.221432f
C2116 two_stage_opamp_dummy_magic_24_0.cap_res_X.n1 GNDA 0.235076f
C2117 two_stage_opamp_dummy_magic_24_0.cap_res_X.t119 GNDA 0.412258f
C2118 two_stage_opamp_dummy_magic_24_0.cap_res_X.t22 GNDA 0.221432f
C2119 two_stage_opamp_dummy_magic_24_0.cap_res_X.n2 GNDA 0.235076f
C2120 two_stage_opamp_dummy_magic_24_0.cap_res_X.t3 GNDA 0.412258f
C2121 two_stage_opamp_dummy_magic_24_0.cap_res_X.t45 GNDA 0.221432f
C2122 two_stage_opamp_dummy_magic_24_0.cap_res_X.n3 GNDA 0.235076f
C2123 two_stage_opamp_dummy_magic_24_0.cap_res_X.t101 GNDA 0.412258f
C2124 two_stage_opamp_dummy_magic_24_0.cap_res_X.t5 GNDA 0.221432f
C2125 two_stage_opamp_dummy_magic_24_0.cap_res_X.n4 GNDA 0.235076f
C2126 two_stage_opamp_dummy_magic_24_0.cap_res_X.t66 GNDA 0.412258f
C2127 two_stage_opamp_dummy_magic_24_0.cap_res_X.t106 GNDA 0.221432f
C2128 two_stage_opamp_dummy_magic_24_0.cap_res_X.n5 GNDA 0.235076f
C2129 two_stage_opamp_dummy_magic_24_0.cap_res_X.t30 GNDA 0.412258f
C2130 two_stage_opamp_dummy_magic_24_0.cap_res_X.t68 GNDA 0.221432f
C2131 two_stage_opamp_dummy_magic_24_0.cap_res_X.n6 GNDA 0.235076f
C2132 two_stage_opamp_dummy_magic_24_0.cap_res_X.t50 GNDA 0.412258f
C2133 two_stage_opamp_dummy_magic_24_0.cap_res_X.t89 GNDA 0.221432f
C2134 two_stage_opamp_dummy_magic_24_0.cap_res_X.n7 GNDA 0.235076f
C2135 two_stage_opamp_dummy_magic_24_0.cap_res_X.t9 GNDA 0.412258f
C2136 two_stage_opamp_dummy_magic_24_0.cap_res_X.t52 GNDA 0.221432f
C2137 two_stage_opamp_dummy_magic_24_0.cap_res_X.n8 GNDA 0.235076f
C2138 two_stage_opamp_dummy_magic_24_0.cap_res_X.t112 GNDA 0.412258f
C2139 two_stage_opamp_dummy_magic_24_0.cap_res_X.t13 GNDA 0.221432f
C2140 two_stage_opamp_dummy_magic_24_0.cap_res_X.n9 GNDA 0.235076f
C2141 two_stage_opamp_dummy_magic_24_0.cap_res_X.t61 GNDA 0.412258f
C2142 two_stage_opamp_dummy_magic_24_0.cap_res_X.t94 GNDA 0.413752f
C2143 two_stage_opamp_dummy_magic_24_0.cap_res_X.t135 GNDA 0.199307f
C2144 two_stage_opamp_dummy_magic_24_0.cap_res_X.n10 GNDA 0.257077f
C2145 two_stage_opamp_dummy_magic_24_0.cap_res_X.t39 GNDA 0.220062f
C2146 two_stage_opamp_dummy_magic_24_0.cap_res_X.n11 GNDA 0.279201f
C2147 two_stage_opamp_dummy_magic_24_0.cap_res_X.t107 GNDA 0.220062f
C2148 two_stage_opamp_dummy_magic_24_0.cap_res_X.n12 GNDA 0.299832f
C2149 two_stage_opamp_dummy_magic_24_0.cap_res_X.t73 GNDA 0.220062f
C2150 two_stage_opamp_dummy_magic_24_0.cap_res_X.n13 GNDA 0.299832f
C2151 two_stage_opamp_dummy_magic_24_0.cap_res_X.t136 GNDA 0.220062f
C2152 two_stage_opamp_dummy_magic_24_0.cap_res_X.n14 GNDA 0.299832f
C2153 two_stage_opamp_dummy_magic_24_0.cap_res_X.t27 GNDA 0.220062f
C2154 two_stage_opamp_dummy_magic_24_0.cap_res_X.n15 GNDA 0.299832f
C2155 two_stage_opamp_dummy_magic_24_0.cap_res_X.t58 GNDA 0.220062f
C2156 two_stage_opamp_dummy_magic_24_0.cap_res_X.n16 GNDA 0.299832f
C2157 two_stage_opamp_dummy_magic_24_0.cap_res_X.t19 GNDA 0.220062f
C2158 two_stage_opamp_dummy_magic_24_0.cap_res_X.n17 GNDA 0.299832f
C2159 two_stage_opamp_dummy_magic_24_0.cap_res_X.t118 GNDA 0.220062f
C2160 two_stage_opamp_dummy_magic_24_0.cap_res_X.n18 GNDA 0.299832f
C2161 two_stage_opamp_dummy_magic_24_0.cap_res_X.t14 GNDA 0.220062f
C2162 two_stage_opamp_dummy_magic_24_0.cap_res_X.n19 GNDA 0.299832f
C2163 two_stage_opamp_dummy_magic_24_0.cap_res_X.t113 GNDA 0.220062f
C2164 two_stage_opamp_dummy_magic_24_0.cap_res_X.n20 GNDA 0.299832f
C2165 two_stage_opamp_dummy_magic_24_0.cap_res_X.t74 GNDA 0.220062f
C2166 two_stage_opamp_dummy_magic_24_0.cap_res_X.n21 GNDA 0.299832f
C2167 two_stage_opamp_dummy_magic_24_0.cap_res_X.t36 GNDA 0.220062f
C2168 two_stage_opamp_dummy_magic_24_0.cap_res_X.n22 GNDA 0.299832f
C2169 two_stage_opamp_dummy_magic_24_0.cap_res_X.t69 GNDA 0.220062f
C2170 two_stage_opamp_dummy_magic_24_0.cap_res_X.n23 GNDA 0.299832f
C2171 two_stage_opamp_dummy_magic_24_0.cap_res_X.t31 GNDA 0.220062f
C2172 two_stage_opamp_dummy_magic_24_0.cap_res_X.n24 GNDA 0.299832f
C2173 two_stage_opamp_dummy_magic_24_0.cap_res_X.t131 GNDA 0.220062f
C2174 two_stage_opamp_dummy_magic_24_0.cap_res_X.n25 GNDA 0.299832f
C2175 two_stage_opamp_dummy_magic_24_0.cap_res_X.t26 GNDA 0.220062f
C2176 two_stage_opamp_dummy_magic_24_0.cap_res_X.n26 GNDA 0.299832f
C2177 two_stage_opamp_dummy_magic_24_0.cap_res_X.t125 GNDA 0.220062f
C2178 two_stage_opamp_dummy_magic_24_0.cap_res_X.n27 GNDA 0.299832f
C2179 two_stage_opamp_dummy_magic_24_0.cap_res_X.t97 GNDA 0.220062f
C2180 two_stage_opamp_dummy_magic_24_0.cap_res_X.n28 GNDA 0.299832f
C2181 two_stage_opamp_dummy_magic_24_0.cap_res_X.t134 GNDA 0.220062f
C2182 two_stage_opamp_dummy_magic_24_0.cap_res_X.n29 GNDA 0.276337f
C2183 two_stage_opamp_dummy_magic_24_0.cap_res_X.t111 GNDA 0.413752f
C2184 two_stage_opamp_dummy_magic_24_0.cap_res_X.t8 GNDA 0.413752f
C2185 two_stage_opamp_dummy_magic_24_0.cap_res_X.t103 GNDA 0.412258f
C2186 two_stage_opamp_dummy_magic_24_0.cap_res_X.t12 GNDA 0.434383f
C2187 two_stage_opamp_dummy_magic_24_0.cap_res_X.t48 GNDA 0.221432f
C2188 two_stage_opamp_dummy_magic_24_0.cap_res_X.n30 GNDA 0.255706f
C2189 two_stage_opamp_dummy_magic_24_0.cap_res_X.t10 GNDA 0.412258f
C2190 two_stage_opamp_dummy_magic_24_0.cap_res_X.t35 GNDA 0.434383f
C2191 two_stage_opamp_dummy_magic_24_0.cap_res_X.t17 GNDA 0.413752f
C2192 two_stage_opamp_dummy_magic_24_0.cap_res_X.t82 GNDA 0.412258f
C2193 two_stage_opamp_dummy_magic_24_0.cap_res_X.t116 GNDA 0.221432f
C2194 two_stage_opamp_dummy_magic_24_0.cap_res_X.n31 GNDA 0.255706f
C2195 two_stage_opamp_dummy_magic_24_0.cap_res_X.t122 GNDA 0.412258f
C2196 two_stage_opamp_dummy_magic_24_0.cap_res_X.t105 GNDA 0.434383f
C2197 two_stage_opamp_dummy_magic_24_0.cap_res_X.t2 GNDA 0.221432f
C2198 two_stage_opamp_dummy_magic_24_0.cap_res_X.n32 GNDA 0.235076f
C2199 two_stage_opamp_dummy_magic_24_0.cap_res_X.t86 GNDA 0.412258f
C2200 two_stage_opamp_dummy_magic_24_0.cap_res_X.t67 GNDA 0.434383f
C2201 two_stage_opamp_dummy_magic_24_0.cap_res_X.t100 GNDA 0.221432f
C2202 two_stage_opamp_dummy_magic_24_0.cap_res_X.n33 GNDA 0.235076f
C2203 two_stage_opamp_dummy_magic_24_0.cap_res_X.t51 GNDA 0.412258f
C2204 two_stage_opamp_dummy_magic_24_0.cap_res_X.t32 GNDA 0.434383f
C2205 two_stage_opamp_dummy_magic_24_0.cap_res_X.t63 GNDA 0.221432f
C2206 two_stage_opamp_dummy_magic_24_0.cap_res_X.n34 GNDA 0.235076f
C2207 two_stage_opamp_dummy_magic_24_0.cap_res_X.n35 GNDA 0.235076f
C2208 two_stage_opamp_dummy_magic_24_0.cap_res_X.t29 GNDA 0.221432f
C2209 two_stage_opamp_dummy_magic_24_0.cap_res_X.t132 GNDA 0.434383f
C2210 two_stage_opamp_dummy_magic_24_0.cap_res_X.t16 GNDA 0.590705f
C2211 two_stage_opamp_dummy_magic_24_0.cap_res_X.t0 GNDA 0.355569f
C2212 VOUT-.n1 GNDA 0.076987f
C2213 VOUT-.n4 GNDA 0.057741f
C2214 VOUT-.n5 GNDA 0.096234f
C2215 VOUT-.n6 GNDA 0.057741f
C2216 VOUT-.n7 GNDA 0.057741f
C2217 VOUT-.n9 GNDA 0.039264f
C2218 VOUT-.n11 GNDA 0.039264f
C2219 VOUT-.n13 GNDA 0.076987f
C2220 VOUT-.n14 GNDA 0.039264f
C2221 VOUT-.n16 GNDA 0.039264f
C2222 VOUT-.n18 GNDA 0.050812f
C2223 VOUT-.n19 GNDA 0.073309f
C2224 VOUT-.n20 GNDA 0.071342f
C2225 VOUT-.n21 GNDA 0.050812f
C2226 VOUT-.n22 GNDA 0.050812f
C2227 VOUT-.n23 GNDA 0.071342f
C2228 VOUT-.n24 GNDA 0.071342f
C2229 VOUT-.n25 GNDA 0.050812f
C2230 VOUT-.n26 GNDA 0.081345f
C2231 VOUT-.t10 GNDA 0.046192f
C2232 VOUT-.t1 GNDA 0.046192f
C2233 VOUT-.n27 GNDA 0.094648f
C2234 VOUT-.n28 GNDA 0.244315f
C2235 VOUT-.t0 GNDA 0.046192f
C2236 VOUT-.t14 GNDA 0.046192f
C2237 VOUT-.n29 GNDA 0.094648f
C2238 VOUT-.n30 GNDA 0.241853f
C2239 VOUT-.n31 GNDA 0.058739f
C2240 VOUT-.t13 GNDA 0.046192f
C2241 VOUT-.t2 GNDA 0.046192f
C2242 VOUT-.n32 GNDA 0.094648f
C2243 VOUT-.n33 GNDA 0.241853f
C2244 VOUT-.n34 GNDA 0.033295f
C2245 VOUT-.t16 GNDA 0.046192f
C2246 VOUT-.t3 GNDA 0.046192f
C2247 VOUT-.n35 GNDA 0.094648f
C2248 VOUT-.n36 GNDA 0.241853f
C2249 VOUT-.n37 GNDA 0.033295f
C2250 VOUT-.t18 GNDA 0.046192f
C2251 VOUT-.t11 GNDA 0.046192f
C2252 VOUT-.n38 GNDA 0.094648f
C2253 VOUT-.n39 GNDA 0.244315f
C2254 VOUT-.n40 GNDA 0.058739f
C2255 VOUT-.t4 GNDA 0.046192f
C2256 VOUT-.t8 GNDA 0.046192f
C2257 VOUT-.n41 GNDA 0.094648f
C2258 VOUT-.n42 GNDA 0.241853f
C2259 VOUT-.n43 GNDA 0.038836f
C2260 VOUT-.n44 GNDA 0.023096f
C2261 VOUT-.n45 GNDA 0.023096f
C2262 VOUT-.n46 GNDA 0.038836f
C2263 VOUT-.n47 GNDA 0.071342f
C2264 VOUT-.n48 GNDA 0.099864f
C2265 VOUT-.n49 GNDA 0.124435f
C2266 VOUT-.n50 GNDA 0.174158f
C2267 VOUT-.n51 GNDA 0.050812f
C2268 VOUT-.n52 GNDA 0.083146f
C2269 VOUT-.n53 GNDA 0.050812f
C2270 VOUT-.n54 GNDA 0.083146f
C2271 VOUT-.n55 GNDA 0.050812f
C2272 VOUT-.n56 GNDA 0.050812f
C2273 VOUT-.n57 GNDA 0.050812f
C2274 VOUT-.n58 GNDA 0.083146f
C2275 VOUT-.n59 GNDA 0.050812f
C2276 VOUT-.n60 GNDA 0.076218f
C2277 VOUT-.n61 GNDA 0.24482f
C2278 VOUT-.n62 GNDA 0.237891f
C2279 VOUT-.n64 GNDA 0.076987f
C2280 VOUT-.n65 GNDA 0.036954f
C2281 VOUT-.n66 GNDA 0.548535f
C2282 VOUT-.n69 GNDA 0.057741f
C2283 VOUT-.n70 GNDA 0.057741f
C2284 VOUT-.t96 GNDA 0.313195f
C2285 VOUT-.t63 GNDA 0.30795f
C2286 VOUT-.n71 GNDA 0.20647f
C2287 VOUT-.t22 GNDA 0.30795f
C2288 VOUT-.n72 GNDA 0.134728f
C2289 VOUT-.t58 GNDA 0.313195f
C2290 VOUT-.t20 GNDA 0.30795f
C2291 VOUT-.n73 GNDA 0.20647f
C2292 VOUT-.t118 GNDA 0.30795f
C2293 VOUT-.t45 GNDA 0.312538f
C2294 VOUT-.t148 GNDA 0.312538f
C2295 VOUT-.t107 GNDA 0.312538f
C2296 VOUT-.t127 GNDA 0.312538f
C2297 VOUT-.t91 GNDA 0.312538f
C2298 VOUT-.t56 GNDA 0.312538f
C2299 VOUT-.t154 GNDA 0.312538f
C2300 VOUT-.t38 GNDA 0.312538f
C2301 VOUT-.t139 GNDA 0.312538f
C2302 VOUT-.t119 GNDA 0.312538f
C2303 VOUT-.t146 GNDA 0.312538f
C2304 VOUT-.t104 GNDA 0.30795f
C2305 VOUT-.n74 GNDA 0.207127f
C2306 VOUT-.t79 GNDA 0.30795f
C2307 VOUT-.n75 GNDA 0.264867f
C2308 VOUT-.t101 GNDA 0.30795f
C2309 VOUT-.n76 GNDA 0.264867f
C2310 VOUT-.t135 GNDA 0.30795f
C2311 VOUT-.n77 GNDA 0.264867f
C2312 VOUT-.t112 GNDA 0.30795f
C2313 VOUT-.n78 GNDA 0.264867f
C2314 VOUT-.t152 GNDA 0.30795f
C2315 VOUT-.n79 GNDA 0.264867f
C2316 VOUT-.t51 GNDA 0.30795f
C2317 VOUT-.n80 GNDA 0.264867f
C2318 VOUT-.t89 GNDA 0.30795f
C2319 VOUT-.n81 GNDA 0.264867f
C2320 VOUT-.t68 GNDA 0.30795f
C2321 VOUT-.n82 GNDA 0.264867f
C2322 VOUT-.t105 GNDA 0.30795f
C2323 VOUT-.n83 GNDA 0.264867f
C2324 VOUT-.t144 GNDA 0.30795f
C2325 VOUT-.n84 GNDA 0.264867f
C2326 VOUT-.n85 GNDA 0.250209f
C2327 VOUT-.t117 GNDA 0.313195f
C2328 VOUT-.t85 GNDA 0.30795f
C2329 VOUT-.n86 GNDA 0.20647f
C2330 VOUT-.t50 GNDA 0.30795f
C2331 VOUT-.t102 GNDA 0.313195f
C2332 VOUT-.t137 GNDA 0.30795f
C2333 VOUT-.n87 GNDA 0.20647f
C2334 VOUT-.n88 GNDA 0.250209f
C2335 VOUT-.t153 GNDA 0.313195f
C2336 VOUT-.t116 GNDA 0.30795f
C2337 VOUT-.n89 GNDA 0.20647f
C2338 VOUT-.t84 GNDA 0.30795f
C2339 VOUT-.t136 GNDA 0.313195f
C2340 VOUT-.t33 GNDA 0.30795f
C2341 VOUT-.n90 GNDA 0.20647f
C2342 VOUT-.n91 GNDA 0.250209f
C2343 VOUT-.t62 GNDA 0.313195f
C2344 VOUT-.t110 GNDA 0.30795f
C2345 VOUT-.n92 GNDA 0.20647f
C2346 VOUT-.t21 GNDA 0.30795f
C2347 VOUT-.t30 GNDA 0.313195f
C2348 VOUT-.t114 GNDA 0.30795f
C2349 VOUT-.n93 GNDA 0.20647f
C2350 VOUT-.n94 GNDA 0.250209f
C2351 VOUT-.t66 GNDA 0.313195f
C2352 VOUT-.t28 GNDA 0.30795f
C2353 VOUT-.n95 GNDA 0.20647f
C2354 VOUT-.t130 GNDA 0.30795f
C2355 VOUT-.t47 GNDA 0.313195f
C2356 VOUT-.t81 GNDA 0.30795f
C2357 VOUT-.n96 GNDA 0.20647f
C2358 VOUT-.n97 GNDA 0.250209f
C2359 VOUT-.t29 GNDA 0.313195f
C2360 VOUT-.t133 GNDA 0.30795f
C2361 VOUT-.n98 GNDA 0.20647f
C2362 VOUT-.t99 GNDA 0.30795f
C2363 VOUT-.t150 GNDA 0.313195f
C2364 VOUT-.t49 GNDA 0.30795f
C2365 VOUT-.n99 GNDA 0.20647f
C2366 VOUT-.n100 GNDA 0.250209f
C2367 VOUT-.t70 GNDA 0.313195f
C2368 VOUT-.t34 GNDA 0.30795f
C2369 VOUT-.n101 GNDA 0.20647f
C2370 VOUT-.t138 GNDA 0.30795f
C2371 VOUT-.t53 GNDA 0.313195f
C2372 VOUT-.t87 GNDA 0.30795f
C2373 VOUT-.n102 GNDA 0.20647f
C2374 VOUT-.n103 GNDA 0.250209f
C2375 VOUT-.t100 GNDA 0.313195f
C2376 VOUT-.t64 GNDA 0.30795f
C2377 VOUT-.n104 GNDA 0.20647f
C2378 VOUT-.t23 GNDA 0.30795f
C2379 VOUT-.t54 GNDA 0.313195f
C2380 VOUT-.t145 GNDA 0.30795f
C2381 VOUT-.n105 GNDA 0.201658f
C2382 VOUT-.t141 GNDA 0.313195f
C2383 VOUT-.t25 GNDA 0.30795f
C2384 VOUT-.n106 GNDA 0.201658f
C2385 VOUT-.t106 GNDA 0.313195f
C2386 VOUT-.t125 GNDA 0.30795f
C2387 VOUT-.n107 GNDA 0.201658f
C2388 VOUT-.t71 GNDA 0.313195f
C2389 VOUT-.t90 GNDA 0.30795f
C2390 VOUT-.n108 GNDA 0.201658f
C2391 VOUT-.t35 GNDA 0.313195f
C2392 VOUT-.t52 GNDA 0.30795f
C2393 VOUT-.n109 GNDA 0.203583f
C2394 VOUT-.t75 GNDA 0.312796f
C2395 VOUT-.t147 GNDA 0.313195f
C2396 VOUT-.t122 GNDA 0.30795f
C2397 VOUT-.n110 GNDA 0.20647f
C2398 VOUT-.t140 GNDA 0.30795f
C2399 VOUT-.n111 GNDA 0.134728f
C2400 VOUT-.t41 GNDA 0.30795f
C2401 VOUT-.n112 GNDA 0.268459f
C2402 VOUT-.t155 GNDA 0.30795f
C2403 VOUT-.n113 GNDA 0.199205f
C2404 VOUT-.t57 GNDA 0.30795f
C2405 VOUT-.n114 GNDA 0.19728f
C2406 VOUT-.t94 GNDA 0.30795f
C2407 VOUT-.n115 GNDA 0.19728f
C2408 VOUT-.t128 GNDA 0.30795f
C2409 VOUT-.n116 GNDA 0.19728f
C2410 VOUT-.t109 GNDA 0.30795f
C2411 VOUT-.n117 GNDA 0.19728f
C2412 VOUT-.t149 GNDA 0.30795f
C2413 VOUT-.n118 GNDA 0.134728f
C2414 VOUT-.t46 GNDA 0.30795f
C2415 VOUT-.n119 GNDA 0.134728f
C2416 VOUT-.n120 GNDA 0.192468f
C2417 VOUT-.t132 GNDA 0.313195f
C2418 VOUT-.t95 GNDA 0.30795f
C2419 VOUT-.n121 GNDA 0.20647f
C2420 VOUT-.t60 GNDA 0.30795f
C2421 VOUT-.t42 GNDA 0.313195f
C2422 VOUT-.t78 GNDA 0.30795f
C2423 VOUT-.n122 GNDA 0.20647f
C2424 VOUT-.n123 GNDA 0.250209f
C2425 VOUT-.t103 GNDA 0.313195f
C2426 VOUT-.t69 GNDA 0.30795f
C2427 VOUT-.n124 GNDA 0.20647f
C2428 VOUT-.t32 GNDA 0.30795f
C2429 VOUT-.t86 GNDA 0.313195f
C2430 VOUT-.t120 GNDA 0.30795f
C2431 VOUT-.n125 GNDA 0.20647f
C2432 VOUT-.n126 GNDA 0.250209f
C2433 VOUT-.t67 GNDA 0.313195f
C2434 VOUT-.t27 GNDA 0.30795f
C2435 VOUT-.n127 GNDA 0.20647f
C2436 VOUT-.t131 GNDA 0.30795f
C2437 VOUT-.t48 GNDA 0.313195f
C2438 VOUT-.t82 GNDA 0.30795f
C2439 VOUT-.n128 GNDA 0.20647f
C2440 VOUT-.n129 GNDA 0.250209f
C2441 VOUT-.t98 GNDA 0.313195f
C2442 VOUT-.t65 GNDA 0.30795f
C2443 VOUT-.n130 GNDA 0.20647f
C2444 VOUT-.t26 GNDA 0.30795f
C2445 VOUT-.t80 GNDA 0.313195f
C2446 VOUT-.t113 GNDA 0.30795f
C2447 VOUT-.n131 GNDA 0.20647f
C2448 VOUT-.n132 GNDA 0.250209f
C2449 VOUT-.t61 GNDA 0.313195f
C2450 VOUT-.t24 GNDA 0.30795f
C2451 VOUT-.n133 GNDA 0.20647f
C2452 VOUT-.t126 GNDA 0.30795f
C2453 VOUT-.t43 GNDA 0.313195f
C2454 VOUT-.t76 GNDA 0.30795f
C2455 VOUT-.n134 GNDA 0.20647f
C2456 VOUT-.n135 GNDA 0.250209f
C2457 VOUT-.t19 GNDA 0.313195f
C2458 VOUT-.t123 GNDA 0.30795f
C2459 VOUT-.n136 GNDA 0.20647f
C2460 VOUT-.t88 GNDA 0.30795f
C2461 VOUT-.t142 GNDA 0.313195f
C2462 VOUT-.t37 GNDA 0.30795f
C2463 VOUT-.n137 GNDA 0.20647f
C2464 VOUT-.n138 GNDA 0.250209f
C2465 VOUT-.t55 GNDA 0.313195f
C2466 VOUT-.t156 GNDA 0.30795f
C2467 VOUT-.n139 GNDA 0.20647f
C2468 VOUT-.t121 GNDA 0.30795f
C2469 VOUT-.t36 GNDA 0.313195f
C2470 VOUT-.t72 GNDA 0.30795f
C2471 VOUT-.n140 GNDA 0.20647f
C2472 VOUT-.n141 GNDA 0.250209f
C2473 VOUT-.t151 GNDA 0.313195f
C2474 VOUT-.t115 GNDA 0.30795f
C2475 VOUT-.n142 GNDA 0.20647f
C2476 VOUT-.t83 GNDA 0.30795f
C2477 VOUT-.t134 GNDA 0.313195f
C2478 VOUT-.t31 GNDA 0.30795f
C2479 VOUT-.n143 GNDA 0.20647f
C2480 VOUT-.n144 GNDA 0.250209f
C2481 VOUT-.t111 GNDA 0.313195f
C2482 VOUT-.t77 GNDA 0.30795f
C2483 VOUT-.n145 GNDA 0.20647f
C2484 VOUT-.t44 GNDA 0.30795f
C2485 VOUT-.t97 GNDA 0.313195f
C2486 VOUT-.t129 GNDA 0.30795f
C2487 VOUT-.n146 GNDA 0.20647f
C2488 VOUT-.n147 GNDA 0.250209f
C2489 VOUT-.t74 GNDA 0.313195f
C2490 VOUT-.t40 GNDA 0.30795f
C2491 VOUT-.n148 GNDA 0.20647f
C2492 VOUT-.t143 GNDA 0.30795f
C2493 VOUT-.t59 GNDA 0.313195f
C2494 VOUT-.t93 GNDA 0.30795f
C2495 VOUT-.n149 GNDA 0.20647f
C2496 VOUT-.n150 GNDA 0.250209f
C2497 VOUT-.t108 GNDA 0.313195f
C2498 VOUT-.t73 GNDA 0.30795f
C2499 VOUT-.n151 GNDA 0.20647f
C2500 VOUT-.t39 GNDA 0.30795f
C2501 VOUT-.n152 GNDA 0.250209f
C2502 VOUT-.t124 GNDA 0.30795f
C2503 VOUT-.n153 GNDA 0.131345f
C2504 VOUT-.t92 GNDA 0.30795f
C2505 VOUT-.n154 GNDA 0.347901f
C2506 VOUT-.n155 GNDA 0.282929f
C2507 VOUT-.n156 GNDA 0.057741f
C2508 VOUT-.n157 GNDA 0.057741f
C2509 VOUT-.n158 GNDA 0.057741f
C2510 VOUT-.n159 GNDA 0.169362f
C2511 VOUT-.n160 GNDA 0.061174f
C2512 VOUT-.n161 GNDA 0.058167f
C2513 VOUT-.n163 GNDA 0.558159f
C2514 VOUT-.n164 GNDA 0.057741f
C2515 VOUT-.n165 GNDA 1.09707f
C2516 VOUT-.n169 GNDA 0.039264f
C2517 VOUT-.n170 GNDA 0.039264f
C2518 VOUT-.n171 GNDA 0.036954f
C2519 VOUT-.n172 GNDA 0.076987f
C2520 VOUT-.n173 GNDA 0.039264f
C2521 VOUT-.n174 GNDA 0.039264f
C2522 VOUT-.n176 GNDA 1.08745f
C2523 VOUT-.n177 GNDA 0.103933f
C2524 VOUT-.t7 GNDA 0.088216f
C2525 VOUT-.n178 GNDA 0.271508f
C2526 VOUT-.n179 GNDA 0.036954f
C2527 VOUT-.t17 GNDA 0.053891f
C2528 VOUT-.t9 GNDA 0.053891f
C2529 VOUT-.n180 GNDA 0.115791f
C2530 VOUT-.n181 GNDA 0.28425f
C2531 VOUT-.n182 GNDA 0.036954f
C2532 VOUT-.n183 GNDA 0.245179f
C2533 VOUT-.t5 GNDA 0.053891f
C2534 VOUT-.t15 GNDA 0.053891f
C2535 VOUT-.n184 GNDA 0.115791f
C2536 VOUT-.n185 GNDA 0.293212f
C2537 VOUT-.n186 GNDA 0.164735f
C2538 VOUT-.t6 GNDA 0.053891f
C2539 VOUT-.t12 GNDA 0.053891f
C2540 VOUT-.n187 GNDA 0.115791f
C2541 VOUT-.n188 GNDA 0.279565f
C2542 VOUT-.n189 GNDA 0.131424f
C2543 VOUT-.n190 GNDA 0.036954f
C2544 VOUT-.n191 GNDA 0.190686f
C2545 VOUT-.n192 GNDA 0.036954f
C2546 VOUT-.n193 GNDA 0.036954f
C2547 VOUT-.n194 GNDA 0.036954f
C2548 VOUT-.n195 GNDA 0.036954f
C2549 VOUT-.n196 GNDA 0.084879f
C2550 VOUT-.n197 GNDA 0.099314f
C2551 VDDA.n16 GNDA 0.142987f
C2552 VDDA.n17 GNDA 0.174762f
C2553 VDDA.n18 GNDA 0.142987f
C2554 VDDA.n19 GNDA 1.11212f
C2555 VDDA.n93 GNDA 0.023235f
C2556 VDDA.n192 GNDA 0.018469f
C2557 VDDA.n197 GNDA 2.02565f
C2558 VDDA.n271 GNDA 0.023235f
C2559 VDDA.n366 GNDA 0.046891f
C2560 VDDA.t73 GNDA 0.012362f
C2561 VDDA.n367 GNDA 0.039542f
C2562 VDDA.n372 GNDA 0.031874f
C2563 VDDA.n373 GNDA 0.013002f
C2564 VDDA.n374 GNDA 0.019424f
C2565 VDDA.t278 GNDA 0.017293f
C2566 VDDA.t27 GNDA 0.013107f
C2567 VDDA.t266 GNDA 0.017293f
C2568 VDDA.n375 GNDA 0.019424f
C2569 VDDA.n376 GNDA 0.012766f
C2570 VDDA.n377 GNDA 0.025975f
C2571 VDDA.n378 GNDA 0.041308f
C2572 VDDA.t273 GNDA 0.015838f
C2573 VDDA.n380 GNDA 0.016112f
C2574 VDDA.n381 GNDA 0.039542f
C2575 VDDA.t272 GNDA 0.029624f
C2576 VDDA.t78 GNDA 0.023235f
C2577 VDDA.t297 GNDA 0.029624f
C2578 VDDA.t298 GNDA 0.012362f
C2579 VDDA.n382 GNDA 0.039542f
C2580 VDDA.n383 GNDA 0.015876f
C2581 VDDA.n384 GNDA 0.02766f
C2582 VDDA.n385 GNDA 0.025856f
C2583 VDDA.n386 GNDA 0.157447f
C2584 VDDA.n391 GNDA 0.015331f
C2585 VDDA.n392 GNDA 0.05229f
C2586 VDDA.n393 GNDA 0.015331f
C2587 VDDA.n394 GNDA 0.05229f
C2588 VDDA.n395 GNDA 0.015331f
C2589 VDDA.n396 GNDA 0.05229f
C2590 VDDA.n397 GNDA 0.015331f
C2591 VDDA.n398 GNDA 0.05229f
C2592 VDDA.n399 GNDA 0.015331f
C2593 VDDA.n400 GNDA 0.061595f
C2594 VDDA.n401 GNDA 0.019317f
C2595 VDDA.t348 GNDA 0.020967f
C2596 VDDA.n402 GNDA 0.070136f
C2597 VDDA.t347 GNDA 0.045425f
C2598 VDDA.t115 GNDA 0.034952f
C2599 VDDA.t149 GNDA 0.034952f
C2600 VDDA.t402 GNDA 0.034952f
C2601 VDDA.t128 GNDA 0.034952f
C2602 VDDA.t16 GNDA 0.034952f
C2603 VDDA.t415 GNDA 0.034952f
C2604 VDDA.t130 GNDA 0.034952f
C2605 VDDA.t417 GNDA 0.034952f
C2606 VDDA.t380 GNDA 0.034952f
C2607 VDDA.t8 GNDA 0.034952f
C2608 VDDA.t332 GNDA 0.045425f
C2609 VDDA.t333 GNDA 0.020967f
C2610 VDDA.n403 GNDA 0.070136f
C2611 VDDA.n404 GNDA 0.018737f
C2612 VDDA.n405 GNDA 0.022694f
C2613 VDDA.n417 GNDA 0.065197f
C2614 VDDA.n419 GNDA 0.034749f
C2615 VDDA.n421 GNDA 0.034749f
C2616 VDDA.n423 GNDA 0.034749f
C2617 VDDA.n425 GNDA 0.046665f
C2618 VDDA.n426 GNDA 0.020852f
C2619 VDDA.n428 GNDA 0.063748f
C2620 VDDA.n430 GNDA 0.063748f
C2621 VDDA.n432 GNDA 0.025802f
C2622 VDDA.n433 GNDA 0.021766f
C2623 VDDA.t359 GNDA 0.017651f
C2624 VDDA.t410 GNDA 0.013107f
C2625 VDDA.t144 GNDA 0.013107f
C2626 VDDA.t147 GNDA 0.013107f
C2627 VDDA.t401 GNDA 0.013107f
C2628 VDDA.t173 GNDA 0.013107f
C2629 VDDA.t404 GNDA 0.013107f
C2630 VDDA.t18 GNDA 0.013107f
C2631 VDDA.t160 GNDA 0.013107f
C2632 VDDA.t101 GNDA 0.013107f
C2633 VDDA.t146 GNDA 0.013107f
C2634 VDDA.t344 GNDA 0.017651f
C2635 VDDA.n434 GNDA 0.021766f
C2636 VDDA.n435 GNDA 0.015601f
C2637 VDDA.n436 GNDA 0.090555f
C2638 VDDA.n437 GNDA 0.017576f
C2639 VDDA.n439 GNDA 0.067323f
C2640 VDDA.n441 GNDA 0.029388f
C2641 VDDA.t288 GNDA 0.017638f
C2642 VDDA.n452 GNDA 0.077749f
C2643 VDDA.n453 GNDA 0.046891f
C2644 VDDA.n455 GNDA 0.025931f
C2645 VDDA.t286 GNDA 0.012362f
C2646 VDDA.n459 GNDA 0.039321f
C2647 VDDA.n464 GNDA 1.11212f
C2648 VDDA.n538 GNDA 0.023235f
C2649 VDDA.n636 GNDA 0.018469f
C2650 VDDA.n692 GNDA 0.023235f
C2651 VDDA.n809 GNDA 0.126007f
C2652 VDDA.n810 GNDA 0.127497f
C2653 VDDA.n813 GNDA 0.746709f
C2654 VDDA.n879 GNDA 0.023235f
C2655 VDDA.n973 GNDA 1.11212f
C2656 VDDA.n976 GNDA 0.127497f
C2657 VDDA.n977 GNDA 0.126007f
C2658 VDDA.n979 GNDA 0.018469f
C2659 VDDA.n981 GNDA 0.018469f
C2660 VDDA.n1027 GNDA 0.023235f
C2661 VDDA.n1147 GNDA 0.127497f
C2662 VDDA.n1148 GNDA 0.126007f
C2663 VDDA.n1150 GNDA 0.018469f
C2664 VDDA.n1152 GNDA 0.018469f
C2665 VDDA.n1154 GNDA 0.018469f
C2666 VDDA.n1157 GNDA 0.126007f
C2667 VDDA.n1158 GNDA 0.127497f
C2668 VDDA.n1161 GNDA 1.66818f
C2669 VDDA.n1227 GNDA 0.023235f
C2670 VDDA.n1368 GNDA 0.270086f
C2671 VDDA.n1393 GNDA 0.02412f
C2672 VDDA.n1404 GNDA 0.027164f
C2673 VDDA.t181 GNDA 0.055507f
C2674 VDDA.t52 GNDA 0.055708f
C2675 VDDA.t69 GNDA 0.052729f
C2676 VDDA.t395 GNDA 0.055507f
C2677 VDDA.t392 GNDA 0.055708f
C2678 VDDA.t99 GNDA 0.052729f
C2679 VDDA.t55 GNDA 0.055507f
C2680 VDDA.t137 GNDA 0.055708f
C2681 VDDA.t387 GNDA 0.052729f
C2682 VDDA.t98 GNDA 0.055507f
C2683 VDDA.t68 GNDA 0.055708f
C2684 VDDA.t58 GNDA 0.052729f
C2685 VDDA.t139 GNDA 0.055507f
C2686 VDDA.t174 GNDA 0.055708f
C2687 VDDA.t394 GNDA 0.052729f
C2688 VDDA.n1458 GNDA 0.037206f
C2689 VDDA.t59 GNDA 0.029629f
C2690 VDDA.n1459 GNDA 0.04037f
C2691 VDDA.t138 GNDA 0.029629f
C2692 VDDA.n1460 GNDA 0.04037f
C2693 VDDA.t393 GNDA 0.029629f
C2694 VDDA.n1461 GNDA 0.04037f
C2695 VDDA.t163 GNDA 0.029629f
C2696 VDDA.n1462 GNDA 0.04037f
C2697 VDDA.t386 GNDA 0.158759f
C2698 VDDA.n1463 GNDA 0.672277f
C2699 VDDA.n1577 GNDA 0.023235f
C2700 VDDA.n1580 GNDA 2.39106f
C2701 VDDA.n1581 GNDA 1.57285f
C2702 VDDA.n1653 GNDA 0.021695f
C2703 VDDA.n1766 GNDA 0.030931f
C2704 VDDA.n1767 GNDA 0.015101f
C2705 VDDA.n1777 GNDA 0.017576f
C2706 VDDA.t325 GNDA 0.014597f
C2707 VDDA.t216 GNDA 0.013107f
C2708 VDDA.t291 GNDA 0.014597f
C2709 VDDA.n1785 GNDA 0.017576f
C2710 VDDA.n1790 GNDA 0.015955f
C2711 VDDA.n1791 GNDA 0.017577f
C2712 VDDA.n1905 GNDA 0.010353f
C2713 VDDA.n1908 GNDA 5.504991f
C2714 VDDA.t419 GNDA 0.117301f
C2715 VDDA.t421 GNDA 0.117301f
C2716 VDDA.t422 GNDA 0.111442f
C2717 VDDA.n1941 GNDA 0.215691f
C2718 VDDA.n1942 GNDA 0.113885f
C2719 VDDA.t420 GNDA 0.110083f
C2720 VDDA.n1943 GNDA 0.14778f
C2721 VDDA.n1944 GNDA 0.078147f
C2722 VDDA.n1949 GNDA 0.056301f
C2723 VDDA.n1950 GNDA 0.056301f
C2724 VDDA.n1952 GNDA 0.026545f
C2725 VDDA.n1956 GNDA 0.026545f
C2726 VDDA.n1958 GNDA 0.026545f
C2727 VDDA.n1960 GNDA 0.026545f
C2728 VDDA.n1962 GNDA 0.026545f
C2729 VDDA.n1964 GNDA 0.026545f
C2730 VDDA.n1966 GNDA 0.026545f
C2731 VDDA.n1968 GNDA 0.026545f
C2732 VDDA.n1970 GNDA 0.026545f
C2733 VDDA.n1972 GNDA 0.026545f
C2734 VDDA.n1976 GNDA 0.026545f
C2735 VDDA.n1978 GNDA 0.026545f
C2736 VDDA.n1980 GNDA 0.026545f
C2737 VDDA.n1982 GNDA 0.026545f
C2738 VDDA.n1984 GNDA 0.026545f
C2739 VDDA.n1986 GNDA 0.026545f
C2740 VDDA.n1988 GNDA 0.026545f
C2741 VDDA.n1990 GNDA 0.036171f
C2742 VDDA.n1991 GNDA 0.011609f
C2743 VDDA.n1994 GNDA 0.01224f
C2744 VDDA.t254 GNDA 0.010305f
C2745 VDDA.t275 GNDA 0.012674f
C2746 VDDA.n1995 GNDA 0.010566f
C2747 VDDA.n1999 GNDA 0.026985f
C2748 VDDA.n2000 GNDA 0.026985f
C2749 VDDA.n2001 GNDA 0.010932f
C2750 VDDA.n2004 GNDA 0.01285f
C2751 VDDA.t257 GNDA 0.010389f
C2752 VDDA.t318 GNDA 0.012481f
C2753 VDDA.n2005 GNDA 0.010064f
C2754 VDDA.n2009 GNDA 0.05737f
C2755 VDDA.n2010 GNDA 0.051833f
C2756 VDDA.n2015 GNDA 0.040811f
C2757 VDDA.n2016 GNDA 0.040811f
C2758 VDDA.t262 GNDA 0.014205f
C2759 VDDA.n2018 GNDA 0.011591f
C2760 VDDA.n2019 GNDA 0.011591f
C2761 VDDA.n2020 GNDA 0.011591f
C2762 VDDA.n2021 GNDA 0.011591f
C2763 VDDA.n2022 GNDA 0.011591f
C2764 VDDA.n2023 GNDA 0.011591f
C2765 VDDA.n2024 GNDA 0.011591f
C2766 VDDA.n2025 GNDA 0.011591f
C2767 VDDA.n2051 GNDA 0.027853f
C2768 VDDA.t263 GNDA 0.029541f
C2769 VDDA.t166 GNDA 0.030385f
C2770 VDDA.t94 GNDA 0.030385f
C2771 VDDA.t56 GNDA 0.030385f
C2772 VDDA.t39 GNDA 0.030385f
C2773 VDDA.t96 GNDA 0.030385f
C2774 VDDA.t179 GNDA 0.030385f
C2775 VDDA.t53 GNDA 0.030385f
C2776 VDDA.t384 GNDA 0.030385f
C2777 VDDA.t388 GNDA 0.030385f
C2778 VDDA.t164 GNDA 0.030385f
C2779 VDDA.t140 GNDA 0.030385f
C2780 VDDA.t177 GNDA 0.030385f
C2781 VDDA.t41 GNDA 0.030385f
C2782 VDDA.t161 GNDA 0.030385f
C2783 VDDA.t175 GNDA 0.030385f
C2784 VDDA.t182 GNDA 0.030385f
C2785 VDDA.t338 GNDA 0.029541f
C2786 VDDA.n2068 GNDA 0.027853f
C2787 VDDA.t337 GNDA 0.014205f
C2788 VDDA.n2072 GNDA 0.056768f
C2789 VDDA.n2073 GNDA 0.039845f
C2790 VDDA.n2074 GNDA 0.039845f
C2791 VDDA.n2075 GNDA 0.039845f
C2792 VDDA.n2076 GNDA 0.039845f
C2793 VDDA.n2077 GNDA 0.039845f
C2794 VDDA.n2078 GNDA 0.039845f
C2795 VDDA.n2079 GNDA 0.039845f
C2796 VDDA.n2080 GNDA 0.033599f
C2797 VDDA.n2081 GNDA 0.038312f
C2798 VDDA.n2083 GNDA 0.018223f
C2799 VDDA.t335 GNDA 0.012314f
C2800 VDDA.t294 GNDA 0.012049f
C2801 VDDA.n2084 GNDA 0.0174f
C2802 VDDA.n2086 GNDA 0.069888f
C2803 VDDA.n2087 GNDA 0.052726f
C2804 VDDA.n2092 GNDA 0.019065f
C2805 VDDA.n2093 GNDA 0.019065f
C2806 VDDA.n2096 GNDA 0.017304f
C2807 VDDA.t315 GNDA 0.012048f
C2808 VDDA.t251 GNDA 0.012048f
C2809 VDDA.n2097 GNDA 0.017304f
C2810 VDDA.n2102 GNDA 0.010336f
C2811 VDDA.t269 GNDA 0.010893f
C2812 VDDA.t341 GNDA 0.010893f
C2813 VDDA.n2103 GNDA 0.010336f
C2814 VDDA.n2111 GNDA 0.017304f
C2815 VDDA.t300 GNDA 0.012048f
C2816 VDDA.t321 GNDA 0.012048f
C2817 VDDA.n2112 GNDA 0.017304f
C2818 VDDA.n2117 GNDA 0.010338f
C2819 VDDA.t282 GNDA 0.010893f
C2820 VDDA.t306 GNDA 0.010893f
C2821 VDDA.n2118 GNDA 0.010338f
C2822 VDDA.n2120 GNDA 0.034994f
C2823 VDDA.n2121 GNDA 0.022085f
C2824 VDDA.n2122 GNDA 0.027343f
C2825 VDDA.n2123 GNDA 0.024662f
C2826 VDDA.n2124 GNDA 0.019409f
C2827 VDDA.n2125 GNDA 0.02209f
C2828 VDDA.n2126 GNDA 0.02209f
C2829 VDDA.n2127 GNDA 0.02209f
C2830 VDDA.n2128 GNDA 0.019409f
C2831 VDDA.n2129 GNDA 0.024662f
C2832 VDDA.n2130 GNDA 0.027343f
C2833 VDDA.n2131 GNDA 0.022084f
C2834 VDDA.n2132 GNDA 0.022084f
C2835 VDDA.n2133 GNDA 0.027343f
C2836 VDDA.n2134 GNDA 0.027939f
C2837 VDDA.n2135 GNDA 0.023282f
C2838 VDDA.n2136 GNDA 0.05743f
C2839 VDDA.n2137 GNDA 0.048556f
C2840 VDDA.n2142 GNDA 0.028002f
C2841 VDDA.n2144 GNDA 0.029789f
C2842 VDDA.n2254 GNDA 0.023235f
C2843 VDDA.n2257 GNDA 6.23584f
C2844 VDDA.n2258 GNDA 2.0177f
C2845 VDDA.n2261 GNDA 0.127497f
C2846 VDDA.n2262 GNDA 0.126007f
C2847 VDDA.n2264 GNDA 0.039321f
C2848 VDDA.n2266 GNDA 0.030385f
C2849 VDDA.n2267 GNDA 0.053444f
C2850 VDDA.n2269 GNDA 0.023839f
C2851 VDDA.n2271 GNDA 0.033546f
C2852 VDDA.n2274 GNDA 0.023839f
C2853 VDDA.n2276 GNDA 0.025931f
C2854 VDDA.n2277 GNDA 0.020241f
C2855 VDDA.n2279 GNDA 0.039843f
C2856 VDDA.t285 GNDA 0.029624f
C2857 VDDA.t113 GNDA 0.023235f
C2858 VDDA.t122 GNDA 0.023235f
C2859 VDDA.t76 GNDA 0.023235f
C2860 VDDA.t107 GNDA 0.023235f
C2861 VDDA.t92 GNDA 0.023235f
C2862 VDDA.t6 GNDA 0.023235f
C2863 VDDA.t88 GNDA 0.023235f
C2864 VDDA.t363 GNDA 0.023235f
C2865 VDDA.t368 GNDA 0.023235f
C2866 VDDA.t370 GNDA 0.023235f
C2867 VDDA.t353 GNDA 0.029624f
C2868 VDDA.t354 GNDA 0.012362f
C2869 VDDA.n2280 GNDA 0.039843f
C2870 VDDA.n2282 GNDA 0.020241f
C2871 VDDA.n2283 GNDA 0.038847f
C2872 VDDA.n2288 GNDA 0.015788f
C2873 VDDA.n2289 GNDA 0.05511f
C2874 VDDA.n2291 GNDA 0.015331f
C2875 VDDA.n2292 GNDA 0.05229f
C2876 VDDA.t304 GNDA 0.020967f
C2877 VDDA.n2293 GNDA 0.015331f
C2878 VDDA.n2294 GNDA 0.05229f
C2879 VDDA.n2295 GNDA 0.015331f
C2880 VDDA.n2296 GNDA 0.05229f
C2881 VDDA.n2297 GNDA 0.015331f
C2882 VDDA.n2298 GNDA 0.05229f
C2883 VDDA.n2299 GNDA 0.015331f
C2884 VDDA.n2300 GNDA 0.061595f
C2885 VDDA.n2301 GNDA 0.019317f
C2886 VDDA.n2302 GNDA 0.070136f
C2887 VDDA.t303 GNDA 0.045425f
C2888 VDDA.t109 GNDA 0.034952f
C2889 VDDA.t63 GNDA 0.034731f
C2890 VDDA.t374 GNDA 0.034478f
C2891 VDDA.t372 GNDA 0.034952f
C2892 VDDA.t111 GNDA 0.034952f
C2893 VDDA.t398 GNDA 0.034952f
C2894 VDDA.t134 GNDA 0.034952f
C2895 VDDA.t142 GNDA 0.034952f
C2896 VDDA.t171 GNDA 0.034952f
C2897 VDDA.t411 GNDA 0.034952f
C2898 VDDA.t312 GNDA 0.045425f
C2899 VDDA.t313 GNDA 0.020967f
C2900 VDDA.n2303 GNDA 0.070136f
C2901 VDDA.n2304 GNDA 0.018737f
C2902 VDDA.n2305 GNDA 0.022694f
C2903 VDDA.n2314 GNDA 0.064944f
C2904 VDDA.n2316 GNDA 0.034622f
C2905 VDDA.n2318 GNDA 0.034622f
C2906 VDDA.n2320 GNDA 0.034622f
C2907 VDDA.n2322 GNDA 0.046538f
C2908 VDDA.n2323 GNDA 0.020852f
C2909 VDDA.n2327 GNDA 0.06345f
C2910 VDDA.n2328 GNDA 0.025802f
C2911 VDDA.n2329 GNDA 0.021766f
C2912 VDDA.t309 GNDA 0.017651f
C2913 VDDA.t396 GNDA 0.013107f
C2914 VDDA.t5 GNDA 0.013107f
C2915 VDDA.t13 GNDA 0.013107f
C2916 VDDA.t152 GNDA 0.013107f
C2917 VDDA.t367 GNDA 0.013107f
C2918 VDDA.t133 GNDA 0.013107f
C2919 VDDA.t15 GNDA 0.013107f
C2920 VDDA.t413 GNDA 0.013107f
C2921 VDDA.t127 GNDA 0.013107f
C2922 VDDA.t397 GNDA 0.013107f
C2923 VDDA.t329 GNDA 0.017651f
C2924 VDDA.n2330 GNDA 0.021766f
C2925 VDDA.n2331 GNDA 0.015601f
C2926 VDDA.n2332 GNDA 0.090555f
C2927 VDDA.n2333 GNDA 0.017576f
C2928 VDDA.n2335 GNDA 0.06345f
C2929 VDDA.n2338 GNDA 0.067323f
C2930 VDDA.n2339 GNDA 0.067323f
C2931 VDDA.n2341 GNDA 0.017576f
C2932 VDDA.n2343 GNDA 0.05511f
C2933 VDDA.n2345 GNDA 0.055705f
C2934 VDDA.t35 GNDA 0.015838f
C2935 VDDA.t29 GNDA 0.015838f
C2936 VDDA.t192 GNDA 0.015838f
C2937 VDDA.t12 GNDA 0.015838f
C2938 VDDA.t260 GNDA 0.017638f
C2939 VDDA.n2355 GNDA 0.021237f
C2940 VDDA.n2361 GNDA 0.06726f
C2941 VDDA.n2363 GNDA 0.029388f
C2942 VDDA.n2364 GNDA 0.018705f
C2943 VDDA.n2365 GNDA 0.018705f
C2944 VDDA.n2381 GNDA 0.019437f
C2945 VDDA.t350 GNDA 0.017638f
C2946 VDDA.t103 GNDA 0.015838f
C2947 VDDA.t118 GNDA 0.015838f
C2948 VDDA.t25 GNDA 0.015838f
C2949 VDDA.t36 GNDA 0.015838f
C2950 VDDA.t356 GNDA 0.017638f
C2951 VDDA.n2389 GNDA 0.021237f
C2952 VDDA.n2393 GNDA 0.067261f
C2953 VDDA.n2394 GNDA 0.055705f
C2954 VDDA.n2395 GNDA 0.067323f
C2955 VDDA.n2396 GNDA 0.017576f
C2956 VDDA.n2398 GNDA 0.05511f
C2957 VDDA.n2399 GNDA 0.05511f
C2958 VDDA.n2401 GNDA 0.077749f
C2959 VDDA.n2403 GNDA 0.015788f
C2960 VDDA.n2404 GNDA 0.038848f
C2961 VDDA.t72 GNDA 0.029624f
C2962 VDDA.t361 GNDA 0.023235f
C2963 VDDA.t74 GNDA 0.023235f
C2964 VDDA.t80 GNDA 0.023235f
C2965 VDDA.t3 GNDA 0.023235f
C2966 VDDA.t90 GNDA 0.023235f
C2967 VDDA.t378 GNDA 0.023235f
C2968 VDDA.t86 GNDA 0.023235f
C2969 VDDA.t376 GNDA 0.023235f
C2970 VDDA.t120 GNDA 0.023235f
C2971 VDDA.t1 GNDA 0.023235f
C2972 VDDA.t408 GNDA 0.029624f
C2973 VDDA.t409 GNDA 0.012362f
C2974 VDDA.n2405 GNDA 0.039542f
C2975 VDDA.n2406 GNDA 0.020419f
C2976 VDDA.n2408 GNDA 0.025931f
C2977 VDDA.n2410 GNDA 0.023839f
C2978 VDDA.n2412 GNDA 0.033546f
C2979 VDDA.n2415 GNDA 0.023839f
C2980 VDDA.n2417 GNDA 0.025931f
C2981 VDDA.n2418 GNDA 0.020419f
C2982 VDDA.n2419 GNDA 0.053445f
C2983 VDDA.n2465 GNDA 0.023235f
C2984 VDDA.n2585 GNDA 0.127497f
C2985 VDDA.n2586 GNDA 0.126007f
C2986 VDDA.n2588 GNDA 0.030385f
C2987 VDDA.n2590 GNDA 0.039321f
C2988 VDDA.n2592 GNDA 0.039321f
C2989 VDDA.n2595 GNDA 0.126007f
C2990 VDDA.n2596 GNDA 0.127497f
C2991 VDDA.n2599 GNDA 1.66818f
C2992 VDDA.n2665 GNDA 0.023235f
C2993 VDDA.n2759 GNDA 1.11212f
C2994 VDDA.n2762 GNDA 0.127497f
C2995 VDDA.n2763 GNDA 0.126007f
C2996 VDDA.n2765 GNDA 0.018469f
C2997 VDDA.n2767 GNDA 0.018469f
C2998 VDDA.n2813 GNDA 0.023235f
C2999 VDDA.n2933 GNDA 0.127497f
C3000 VDDA.n2934 GNDA 0.126007f
C3001 VDDA.n2936 GNDA 0.018469f
C3002 VDDA.n2938 GNDA 0.018469f
C3003 VDDA.n2939 GNDA 0.018469f
C3004 VDDA.n2943 GNDA 0.126007f
C3005 VDDA.n2944 GNDA 0.127497f
C3006 VDDA.n2947 GNDA 59.573902f
C3007 VDDA.n2948 GNDA 0.071493f
C3008 VDDA.n2949 GNDA 0.071493f
C3009 VDDA.n2950 GNDA 0.071493f
C3010 VDDA.n2951 GNDA 0.071493f
C3011 VDDA.n2952 GNDA 0.071493f
C3012 VDDA.n2953 GNDA 0.071493f
C3013 VDDA.n2954 GNDA 0.071493f
C3014 VDDA.n2955 GNDA 0.071493f
C3015 VDDA.n2956 GNDA 0.071493f
C3016 VDDA.n2957 GNDA 0.071493f
C3017 VDDA.n2958 GNDA 0.071493f
C3018 VDDA.n2959 GNDA 0.071493f
C3019 VDDA.n2960 GNDA 0.071493f
C3020 VDDA.n2961 GNDA 0.071493f
C3021 VDDA.n2962 GNDA 0.071493f
C3022 VDDA.n2963 GNDA 0.071493f
C3023 VDDA.n2964 GNDA 0.071493f
C3024 VDDA.n2965 GNDA 0.091353f
C3025 VDDA.n2966 GNDA 0.071493f
C3026 VDDA.n2967 GNDA 0.071493f
C3027 VDDA.n2968 GNDA 0.071493f
C3028 VDDA.n2969 GNDA 0.071493f
C3029 VDDA.n2970 GNDA 0.071493f
C3030 VDDA.n2971 GNDA 0.071493f
C3031 VDDA.n2972 GNDA 0.071493f
C3032 VDDA.n2973 GNDA 0.071493f
C3033 VDDA.n2974 GNDA 0.071493f
C3034 VDDA.n2975 GNDA 0.071493f
C3035 VDDA.n2976 GNDA 0.071493f
C3036 VDDA.n2977 GNDA 0.071493f
C3037 VDDA.n2978 GNDA 0.071493f
C3038 VDDA.n2979 GNDA 0.071493f
C3039 VDDA.n2980 GNDA 0.071493f
C3040 VDDA.n2981 GNDA 0.071493f
C3041 VDDA.n2982 GNDA 0.142987f
C3042 VDDA.n2984 GNDA 0.071493f
C3043 VDDA.n2987 GNDA 0.071493f
C3044 VDDA.n2990 GNDA 0.071493f
C3045 VDDA.n2993 GNDA 0.071493f
C3046 VDDA.n2996 GNDA 0.071493f
C3047 VDDA.n2999 GNDA 0.071493f
C3048 VDDA.n3002 GNDA 0.071493f
C3049 VDDA.n3005 GNDA 0.071493f
C3050 VDDA.n3008 GNDA 0.071493f
C3051 VDDA.n3011 GNDA 0.071493f
C3052 VDDA.n3014 GNDA 0.071493f
C3053 VDDA.n3017 GNDA 0.071493f
C3054 VDDA.n3020 GNDA 0.071493f
C3055 VDDA.n3023 GNDA 0.071493f
C3056 VDDA.n3026 GNDA 0.071493f
C3057 VDDA.n3029 GNDA 0.071493f
C3058 VDDA.n3032 GNDA 0.071493f
C3059 VDDA.n3035 GNDA 0.091353f
C3060 VDDA.n3038 GNDA 0.071493f
C3061 VDDA.n3041 GNDA 0.071493f
C3062 VDDA.n3044 GNDA 0.071493f
C3063 VDDA.n3047 GNDA 0.071493f
C3064 VDDA.n3050 GNDA 0.071493f
C3065 VDDA.n3053 GNDA 0.071493f
C3066 VDDA.n3056 GNDA 0.071493f
C3067 VDDA.n3059 GNDA 0.071493f
C3068 VDDA.n3062 GNDA 0.071493f
C3069 VDDA.n3065 GNDA 0.071493f
C3070 VDDA.n3068 GNDA 0.071493f
C3071 VDDA.n3071 GNDA 0.071493f
C3072 VDDA.n3074 GNDA 0.071493f
C3073 VDDA.n3077 GNDA 0.071493f
C3074 VDDA.n3080 GNDA 0.071493f
C3075 VDDA.n3083 GNDA 0.071493f
C3076 VDDA.n3086 GNDA 0.142987f
C3077 VDDA.n3087 GNDA 0.142987f
C3078 VDDA.n3088 GNDA 0.142987f
C3079 VDDA.n3089 GNDA 0.142987f
C3080 VDDA.n3090 GNDA 0.142987f
C3081 VDDA.n3091 GNDA 0.142987f
C3082 VDDA.n3092 GNDA 0.142987f
C3083 VDDA.n3093 GNDA 0.142987f
C3084 VDDA.n3094 GNDA 0.142987f
C3085 VDDA.n3095 GNDA 0.142987f
C3086 VDDA.n3096 GNDA 0.142987f
C3087 VDDA.n3097 GNDA 0.142987f
C3088 VDDA.n3098 GNDA 0.142987f
C3089 VDDA.n3099 GNDA 0.142987f
C3090 VDDA.n3100 GNDA 0.142987f
C3091 VDDA.n3103 GNDA 0.142987f
C3092 VDDA.n3105 GNDA 0.142987f
C3093 VDDA.n3107 GNDA 0.142987f
C3094 VDDA.n3109 GNDA 0.142987f
C3095 VDDA.n3111 GNDA 0.142987f
C3096 VDDA.n3113 GNDA 0.142987f
C3097 VDDA.n3115 GNDA 0.142987f
C3098 VDDA.n3117 GNDA 0.142987f
C3099 VDDA.n3119 GNDA 0.142987f
C3100 VDDA.n3121 GNDA 0.142987f
C3101 VDDA.n3123 GNDA 0.142987f
C3102 VDDA.n3125 GNDA 0.142987f
C3103 VDDA.n3127 GNDA 0.142987f
C3104 VDDA.n3129 GNDA 0.142987f
C3105 VDDA.n3131 GNDA 0.142987f
C3106 VDDA.n3132 GNDA 0.087381f
C3107 VDDA.n3133 GNDA 59.089302f
C3108 VDDA.n3134 GNDA 0.466693f
C3109 bgr_11_0.PFET_GATE_10uA.t28 GNDA 0.023614f
C3110 bgr_11_0.PFET_GATE_10uA.t20 GNDA 0.023614f
C3111 bgr_11_0.PFET_GATE_10uA.n0 GNDA 0.082684f
C3112 bgr_11_0.PFET_GATE_10uA.t13 GNDA 0.020346f
C3113 bgr_11_0.PFET_GATE_10uA.t24 GNDA 0.030076f
C3114 bgr_11_0.PFET_GATE_10uA.n1 GNDA 0.03314f
C3115 bgr_11_0.PFET_GATE_10uA.t17 GNDA 0.020346f
C3116 bgr_11_0.PFET_GATE_10uA.t25 GNDA 0.030076f
C3117 bgr_11_0.PFET_GATE_10uA.n2 GNDA 0.03314f
C3118 bgr_11_0.PFET_GATE_10uA.n3 GNDA 0.032464f
C3119 bgr_11_0.PFET_GATE_10uA.n4 GNDA 1.03417f
C3120 bgr_11_0.PFET_GATE_10uA.t3 GNDA 0.363431f
C3121 bgr_11_0.PFET_GATE_10uA.t0 GNDA 0.324056f
C3122 bgr_11_0.PFET_GATE_10uA.t2 GNDA 0.020867f
C3123 bgr_11_0.PFET_GATE_10uA.t7 GNDA 0.020867f
C3124 bgr_11_0.PFET_GATE_10uA.n5 GNDA 0.045075f
C3125 bgr_11_0.PFET_GATE_10uA.n6 GNDA 1.1187f
C3126 bgr_11_0.PFET_GATE_10uA.t9 GNDA 0.020867f
C3127 bgr_11_0.PFET_GATE_10uA.t5 GNDA 0.020867f
C3128 bgr_11_0.PFET_GATE_10uA.n7 GNDA 0.045075f
C3129 bgr_11_0.PFET_GATE_10uA.n8 GNDA 0.455737f
C3130 bgr_11_0.PFET_GATE_10uA.t8 GNDA 0.020867f
C3131 bgr_11_0.PFET_GATE_10uA.t4 GNDA 0.020867f
C3132 bgr_11_0.PFET_GATE_10uA.n9 GNDA 0.045075f
C3133 bgr_11_0.PFET_GATE_10uA.n10 GNDA 0.446347f
C3134 bgr_11_0.PFET_GATE_10uA.t6 GNDA 0.020867f
C3135 bgr_11_0.PFET_GATE_10uA.t1 GNDA 0.020867f
C3136 bgr_11_0.PFET_GATE_10uA.n11 GNDA 0.045075f
C3137 bgr_11_0.PFET_GATE_10uA.n12 GNDA 0.700571f
C3138 bgr_11_0.PFET_GATE_10uA.n13 GNDA 2.98162f
C3139 bgr_11_0.PFET_GATE_10uA.t26 GNDA 0.074194f
C3140 bgr_11_0.PFET_GATE_10uA.n14 GNDA 1.61003f
C3141 bgr_11_0.PFET_GATE_10uA.t15 GNDA 0.020346f
C3142 bgr_11_0.PFET_GATE_10uA.t10 GNDA 0.030076f
C3143 bgr_11_0.PFET_GATE_10uA.n15 GNDA 0.03314f
C3144 bgr_11_0.PFET_GATE_10uA.t21 GNDA 0.020346f
C3145 bgr_11_0.PFET_GATE_10uA.t11 GNDA 0.030076f
C3146 bgr_11_0.PFET_GATE_10uA.n16 GNDA 0.03314f
C3147 bgr_11_0.PFET_GATE_10uA.n17 GNDA 0.031974f
C3148 bgr_11_0.PFET_GATE_10uA.n18 GNDA 1.29057f
C3149 bgr_11_0.PFET_GATE_10uA.t14 GNDA 0.020346f
C3150 bgr_11_0.PFET_GATE_10uA.t19 GNDA 0.020346f
C3151 bgr_11_0.PFET_GATE_10uA.t18 GNDA 0.020346f
C3152 bgr_11_0.PFET_GATE_10uA.t27 GNDA 0.030076f
C3153 bgr_11_0.PFET_GATE_10uA.n19 GNDA 0.037221f
C3154 bgr_11_0.PFET_GATE_10uA.n20 GNDA 0.026606f
C3155 bgr_11_0.PFET_GATE_10uA.n21 GNDA 0.020737f
C3156 bgr_11_0.PFET_GATE_10uA.t23 GNDA 0.020346f
C3157 bgr_11_0.PFET_GATE_10uA.t16 GNDA 0.020346f
C3158 bgr_11_0.PFET_GATE_10uA.t12 GNDA 0.020346f
C3159 bgr_11_0.PFET_GATE_10uA.t22 GNDA 0.030076f
C3160 bgr_11_0.PFET_GATE_10uA.n22 GNDA 0.037221f
C3161 bgr_11_0.PFET_GATE_10uA.n23 GNDA 0.026606f
C3162 bgr_11_0.PFET_GATE_10uA.n24 GNDA 0.020737f
C3163 bgr_11_0.PFET_GATE_10uA.n25 GNDA 0.059033f
C3164 bgr_11_0.1st_Vout_2.n0 GNDA 1.07305f
C3165 bgr_11_0.1st_Vout_2.n1 GNDA 0.297625f
C3166 bgr_11_0.1st_Vout_2.n2 GNDA 0.668271f
C3167 bgr_11_0.1st_Vout_2.n3 GNDA 0.091542f
C3168 bgr_11_0.1st_Vout_2.n4 GNDA 0.158156f
C3169 bgr_11_0.1st_Vout_2.t14 GNDA 0.011681f
C3170 bgr_11_0.1st_Vout_2.n6 GNDA 0.010675f
C3171 bgr_11_0.1st_Vout_2.n7 GNDA 0.115898f
C3172 bgr_11_0.1st_Vout_2.n8 GNDA 0.0146f
C3173 bgr_11_0.1st_Vout_2.t15 GNDA 0.011528f
C3174 bgr_11_0.1st_Vout_2.t29 GNDA 0.194725f
C3175 bgr_11_0.1st_Vout_2.t32 GNDA 0.198042f
C3176 bgr_11_0.1st_Vout_2.t27 GNDA 0.194725f
C3177 bgr_11_0.1st_Vout_2.t20 GNDA 0.194725f
C3178 bgr_11_0.1st_Vout_2.t12 GNDA 0.198042f
C3179 bgr_11_0.1st_Vout_2.t13 GNDA 0.198042f
C3180 bgr_11_0.1st_Vout_2.t31 GNDA 0.194725f
C3181 bgr_11_0.1st_Vout_2.t25 GNDA 0.194725f
C3182 bgr_11_0.1st_Vout_2.t19 GNDA 0.198042f
C3183 bgr_11_0.1st_Vout_2.t30 GNDA 0.198042f
C3184 bgr_11_0.1st_Vout_2.t24 GNDA 0.194725f
C3185 bgr_11_0.1st_Vout_2.t18 GNDA 0.194725f
C3186 bgr_11_0.1st_Vout_2.t11 GNDA 0.198042f
C3187 bgr_11_0.1st_Vout_2.t23 GNDA 0.198042f
C3188 bgr_11_0.1st_Vout_2.t17 GNDA 0.194725f
C3189 bgr_11_0.1st_Vout_2.t10 GNDA 0.194725f
C3190 bgr_11_0.1st_Vout_2.t28 GNDA 0.198042f
C3191 bgr_11_0.1st_Vout_2.t8 GNDA 0.198042f
C3192 bgr_11_0.1st_Vout_2.t16 GNDA 0.194725f
C3193 bgr_11_0.1st_Vout_2.t22 GNDA 0.194725f
C3194 bgr_11_0.1st_Vout_2.n9 GNDA 0.641071f
C3195 bgr_11_0.1st_Vout_2.n10 GNDA 0.010675f
C3196 bgr_11_0.1st_Vout_2.n11 GNDA 0.0146f
C3197 bgr_11_0.1st_Vout_2.n12 GNDA 0.14235f
C3198 bgr_11_0.1st_Vout_2.t4 GNDA 0.044569f
.ends

