magic
tech sky130A
magscale 1 2
timestamp 1737739666
<< nwell >>
rect -38 -838 314 -517
rect 592 -838 944 -517
rect 1222 -838 1574 -517
rect 1852 -838 2204 -517
rect 2482 -838 2834 -517
rect 3112 -838 3464 -517
rect 3742 -838 4094 -517
rect 4372 -838 4724 -517
<< pwell >>
rect 212 -277 246 -239
rect 842 -277 876 -239
rect 1472 -277 1506 -239
rect 2102 -277 2136 -239
rect 2732 -277 2766 -239
rect 3362 -277 3396 -239
rect 3992 -277 4026 -239
rect 4622 -277 4656 -239
rect 5 -459 275 -277
rect 635 -459 905 -277
rect 1265 -459 1535 -277
rect 1895 -459 2165 -277
rect 2525 -459 2795 -277
rect 3155 -459 3425 -277
rect 3785 -459 4055 -277
rect 4415 -459 4685 -277
<< locali >>
rect 107 -435 173 -307
rect 737 -435 803 -307
rect 1367 -435 1433 -307
rect 1997 -435 2063 -307
rect 2627 -435 2693 -307
rect 3257 -435 3323 -307
rect 3887 -435 3953 -307
rect 4517 -435 4583 -307
rect 17 -521 87 -471
rect 121 -555 155 -435
rect 189 -521 259 -471
rect 647 -521 717 -471
rect 751 -555 785 -435
rect 819 -521 889 -471
rect 1277 -521 1347 -471
rect 1381 -555 1415 -435
rect 1449 -521 1519 -471
rect 1907 -521 1977 -471
rect 2011 -555 2045 -435
rect 2079 -521 2149 -471
rect 2537 -521 2607 -471
rect 2641 -555 2675 -435
rect 2709 -521 2779 -471
rect 3167 -521 3237 -471
rect 3271 -555 3305 -435
rect 3339 -521 3409 -471
rect 3797 -521 3867 -471
rect 3901 -555 3935 -435
rect 3969 -521 4039 -471
rect 4427 -521 4497 -471
rect 4531 -555 4565 -435
rect 4599 -521 4669 -471
rect 121 -589 257 -555
rect 751 -589 887 -555
rect 1381 -589 1517 -555
rect 2011 -589 2147 -555
rect 2641 -589 2777 -555
rect 3271 -589 3407 -555
rect 3901 -589 4037 -555
rect 4531 -589 4667 -555
rect 191 -746 257 -589
rect 821 -746 887 -589
rect 1451 -746 1517 -589
rect 2081 -746 2147 -589
rect 2711 -746 2777 -589
rect 3341 -746 3407 -589
rect 3971 -746 4037 -589
rect 4601 -746 4667 -589
<< metal1 >>
rect 0 -304 276 -208
rect 630 -304 906 -208
rect 1260 -304 1536 -208
rect 1890 -304 2166 -208
rect 2520 -304 2796 -208
rect 3150 -304 3426 -208
rect 3780 -304 4056 -208
rect 4410 -304 4686 -208
rect 0 -848 276 -752
rect 630 -848 906 -752
rect 1260 -848 1536 -752
rect 1890 -848 2166 -752
rect 2520 -848 2796 -752
rect 3150 -848 3426 -752
rect 3780 -848 4056 -752
rect 4410 -848 4686 -752
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_0
timestamp 1737724875
transform 1 0 0 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_1
timestamp 1737724875
transform 1 0 630 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_2
timestamp 1737724875
transform 1 0 1260 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_3
timestamp 1737724875
transform 1 0 1890 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_4
timestamp 1737724875
transform 1 0 2520 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_5
timestamp 1737724875
transform 1 0 3150 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_6
timestamp 1737724875
transform 1 0 3780 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_7
timestamp 1737724875
transform 1 0 4410 0 1 0
box -38 -48 314 592
<< labels >>
rlabel locali s 4601 -746 4667 -589 2 Y
port 7 nsew signal output
rlabel locali s 4531 -589 4667 -555 2 Y
port 7 nsew signal output
rlabel locali s 4531 -555 4565 -435 2 Y
port 7 nsew signal output
rlabel locali s 4517 -435 4583 -307 2 Y
port 7 nsew signal output
rlabel metal1 s 4410 -848 4686 -752 2 VPWR
port 6 nsew power bidirectional abutment
rlabel nwell s 4372 -838 4724 -517 2 VPB
port 5 nsew power bidirectional
rlabel pwell s 4415 -459 4685 -277 2 VNB
port 4 nsew ground bidirectional
rlabel pwell s 4622 -277 4656 -239 2 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 4410 -304 4686 -208 4 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 4599 -521 4669 -471 2 B
port 2 nsew signal input
rlabel locali s 4427 -521 4497 -471 2 A
port 1 nsew signal input
rlabel locali s 3971 -746 4037 -589 2 Y
port 7 nsew signal output
rlabel locali s 3901 -589 4037 -555 2 Y
port 7 nsew signal output
rlabel locali s 3901 -555 3935 -435 2 Y
port 7 nsew signal output
rlabel locali s 3887 -435 3953 -307 2 Y
port 7 nsew signal output
rlabel metal1 s 3780 -848 4056 -752 2 VPWR
port 6 nsew power bidirectional abutment
rlabel nwell s 3742 -838 4094 -517 2 VPB
port 5 nsew power bidirectional
rlabel pwell s 3785 -459 4055 -277 2 VNB
port 4 nsew ground bidirectional
rlabel pwell s 3992 -277 4026 -239 2 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 3780 -304 4056 -208 4 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 3969 -521 4039 -471 2 B
port 2 nsew signal input
rlabel locali s 3797 -521 3867 -471 2 A
port 1 nsew signal input
rlabel locali s 3341 -746 3407 -589 2 Y
port 7 nsew signal output
rlabel locali s 3271 -589 3407 -555 2 Y
port 7 nsew signal output
rlabel locali s 3271 -555 3305 -435 2 Y
port 7 nsew signal output
rlabel locali s 3257 -435 3323 -307 2 Y
port 7 nsew signal output
rlabel metal1 s 3150 -848 3426 -752 2 VPWR
port 6 nsew power bidirectional abutment
rlabel nwell s 3112 -838 3464 -517 2 VPB
port 5 nsew power bidirectional
rlabel pwell s 3155 -459 3425 -277 2 VNB
port 4 nsew ground bidirectional
rlabel pwell s 3362 -277 3396 -239 2 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 3150 -304 3426 -208 4 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 3339 -521 3409 -471 2 B
port 2 nsew signal input
rlabel locali s 3167 -521 3237 -471 2 A
port 1 nsew signal input
rlabel locali s 2711 -746 2777 -589 2 Y
port 7 nsew signal output
rlabel locali s 2641 -589 2777 -555 2 Y
port 7 nsew signal output
rlabel locali s 2641 -555 2675 -435 2 Y
port 7 nsew signal output
rlabel locali s 2627 -435 2693 -307 2 Y
port 7 nsew signal output
rlabel metal1 s 2520 -848 2796 -752 2 VPWR
port 6 nsew power bidirectional abutment
rlabel nwell s 2482 -838 2834 -517 2 VPB
port 5 nsew power bidirectional
rlabel pwell s 2525 -459 2795 -277 2 VNB
port 4 nsew ground bidirectional
rlabel pwell s 2732 -277 2766 -239 2 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 2520 -304 2796 -208 4 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 2709 -521 2779 -471 2 B
port 2 nsew signal input
rlabel locali s 2537 -521 2607 -471 2 A
port 1 nsew signal input
rlabel locali s 2081 -746 2147 -589 2 Y
port 7 nsew signal output
rlabel locali s 2011 -589 2147 -555 2 Y
port 7 nsew signal output
rlabel locali s 2011 -555 2045 -435 2 Y
port 7 nsew signal output
rlabel locali s 1997 -435 2063 -307 2 Y
port 7 nsew signal output
rlabel metal1 s 1890 -848 2166 -752 2 VPWR
port 6 nsew power bidirectional abutment
rlabel nwell s 1852 -838 2204 -517 2 VPB
port 5 nsew power bidirectional
rlabel pwell s 1895 -459 2165 -277 2 VNB
port 4 nsew ground bidirectional
rlabel pwell s 2102 -277 2136 -239 2 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 1890 -304 2166 -208 4 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 2079 -521 2149 -471 2 B
port 2 nsew signal input
rlabel locali s 1907 -521 1977 -471 2 A
port 1 nsew signal input
rlabel locali s 1451 -746 1517 -589 2 Y
port 7 nsew signal output
rlabel locali s 1381 -589 1517 -555 2 Y
port 7 nsew signal output
rlabel locali s 1381 -555 1415 -435 2 Y
port 7 nsew signal output
rlabel locali s 1367 -435 1433 -307 2 Y
port 7 nsew signal output
rlabel metal1 s 1260 -848 1536 -752 2 VPWR
port 6 nsew power bidirectional abutment
rlabel nwell s 1222 -838 1574 -517 2 VPB
port 5 nsew power bidirectional
rlabel pwell s 1265 -459 1535 -277 2 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1472 -277 1506 -239 2 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 1260 -304 1536 -208 4 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1449 -521 1519 -471 2 B
port 2 nsew signal input
rlabel locali s 1277 -521 1347 -471 2 A
port 1 nsew signal input
rlabel locali s 821 -746 887 -589 2 Y
port 7 nsew signal output
rlabel locali s 751 -589 887 -555 2 Y
port 7 nsew signal output
rlabel locali s 751 -555 785 -435 2 Y
port 7 nsew signal output
rlabel locali s 737 -435 803 -307 2 Y
port 7 nsew signal output
rlabel metal1 s 630 -848 906 -752 2 VPWR
port 6 nsew power bidirectional abutment
rlabel nwell s 592 -838 944 -517 2 VPB
port 5 nsew power bidirectional
rlabel pwell s 635 -459 905 -277 2 VNB
port 4 nsew ground bidirectional
rlabel pwell s 842 -277 876 -239 2 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 630 -304 906 -208 4 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 819 -521 889 -471 2 B
port 2 nsew signal input
rlabel locali s 647 -521 717 -471 2 A
port 1 nsew signal input
rlabel locali s 191 -746 257 -589 2 Y
port 7 nsew signal output
rlabel locali s 121 -589 257 -555 2 Y
port 7 nsew signal output
rlabel locali s 121 -555 155 -435 2 Y
port 7 nsew signal output
rlabel locali s 107 -435 173 -307 2 Y
port 7 nsew signal output
rlabel metal1 s 0 -848 276 -752 2 VPWR
port 6 nsew power bidirectional abutment
rlabel nwell s -38 -838 314 -517 2 VPB
port 5 nsew power bidirectional
rlabel pwell s 5 -459 275 -277 2 VNB
port 4 nsew ground bidirectional
rlabel pwell s 212 -277 246 -239 2 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 -304 276 -208 4 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 189 -521 259 -471 2 B
port 2 nsew signal input
rlabel locali s 17 -521 87 -471 2 A
port 1 nsew signal input
<< end >>
