* PEX produced on Tue Jul  8 11:45:19 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 GNDA.t214 bgr_0.NFET_GATE_10uA.t5 two_stage_opamp_dummy_magic_0.Vb3.t4 GNDA.t213 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1 bgr_0.V_TOP.t13 VDDA.t430 VDDA.t432 VDDA.t431 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X2 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 GNDA.t57 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X3 two_stage_opamp_dummy_magic_0.VD2.t16 GNDA.t306 GNDA.t308 GNDA.t307 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X4 VOUT-.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5 VDDA.t468 bgr_0.V_TOP.t14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 VDDA.t467 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 two_stage_opamp_dummy_magic_0.Y.t25 GNDA.t60 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X7 VOUT-.t20 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8 VOUT-.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 bgr_0.Vin+.t5 bgr_0.V_TOP.t15 VDDA.t108 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X10 VDDA.t271 bgr_0.V_mir1.t17 bgr_0.1st_Vout_1.t5 VDDA.t270 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X11 two_stage_opamp_dummy_magic_0.V_err_gate.t4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X12 VOUT-.t22 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 bgr_0.1st_Vout_2.t11 bgr_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X14 VOUT-.t23 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 two_stage_opamp_dummy_magic_0.Y.t20 two_stage_opamp_dummy_magic_0.Vb2.t11 two_stage_opamp_dummy_magic_0.VD4.t25 two_stage_opamp_dummy_magic_0.VD4.t24 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X16 VDDA.t24 two_stage_opamp_dummy_magic_0.X.t25 VOUT+.t11 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X17 two_stage_opamp_dummy_magic_0.Y.t22 two_stage_opamp_dummy_magic_0.Vb1.t6 two_stage_opamp_dummy_magic_0.VD2.t19 GNDA.t331 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X18 bgr_0.1st_Vout_2.t10 bgr_0.V_CUR_REF_REG.t3 bgr_0.V_p_2.t9 GNDA.t355 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X19 VOUT-.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 VOUT-.t25 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 a_6810_23838.t1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 GNDA.t337 sky130_fd_pr__res_xhigh_po_0p35 l=4.2
X22 a_7460_23988.t0 bgr_0.Vin+.t0 GNDA.t110 sky130_fd_pr__res_xhigh_po_0p35 l=6
X23 VDDA.t229 two_stage_opamp_dummy_magic_0.X.t26 VOUT+.t10 VDDA.t228 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X24 VOUT-.t26 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 VOUT+.t16 GNDA.t303 GNDA.t305 GNDA.t304 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X26 bgr_0.1st_Vout_2.t12 bgr_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 VDDA.t429 VDDA.t427 bgr_0.NFET_GATE_10uA.t3 VDDA.t428 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X28 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 bgr_0.PFET_GATE_10uA.t10 VDDA.t214 VDDA.t213 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X29 VDDA.t182 two_stage_opamp_dummy_magic_0.V_err_gate.t14 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 VDDA.t181 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X30 VDDA.t196 bgr_0.PFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 VDDA.t195 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X31 VOUT+.t19 two_stage_opamp_dummy_magic_0.cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 VOUT+.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 VOUT+.t21 two_stage_opamp_dummy_magic_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 VOUT-.t27 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 bgr_0.1st_Vout_1.t11 bgr_0.cap_res1.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 VOUT-.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 VOUT-.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 bgr_0.1st_Vout_2.t6 bgr_0.V_mir2.t17 VDDA.t237 VDDA.t236 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X39 VDDA.t110 bgr_0.V_TOP.t16 bgr_0.Vin-.t7 VDDA.t109 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X40 VOUT+.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X41 two_stage_opamp_dummy_magic_0.V_p_mir.t1 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 GNDA.t147 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X42 VOUT-.t3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 GNDA.t32 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X43 bgr_0.1st_Vout_1.t10 bgr_0.Vin+.t6 bgr_0.V_p_1.t9 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X44 VDDA.t58 two_stage_opamp_dummy_magic_0.Y.t26 VOUT-.t5 VDDA.t57 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X45 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 two_stage_opamp_dummy_magic_0.X.t27 VDDA.t241 GNDA.t150 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X46 VOUT-.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 bgr_0.cap_res2.t20 bgr_0.PFET_GATE_10uA.t6 GNDA.t148 sky130_fd_pr__res_high_po_0p35 l=2.05
X48 VDDA.t426 VDDA.t424 two_stage_opamp_dummy_magic_0.V_err_gate.t11 VDDA.t425 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X49 bgr_0.1st_Vout_1.t12 bgr_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 two_stage_opamp_dummy_magic_0.V_err_p.t18 two_stage_opamp_dummy_magic_0.V_err_gate.t15 VDDA.t15 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X51 VOUT-.t31 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 VOUT+.t23 two_stage_opamp_dummy_magic_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X53 a_14560_5068.t1 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA.t67 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X54 two_stage_opamp_dummy_magic_0.Y.t0 two_stage_opamp_dummy_magic_0.Vb2.t12 two_stage_opamp_dummy_magic_0.VD4.t23 two_stage_opamp_dummy_magic_0.VD4.t22 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X55 two_stage_opamp_dummy_magic_0.V_err_p.t6 two_stage_opamp_dummy_magic_0.V_tot.t4 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X56 two_stage_opamp_dummy_magic_0.X.t23 two_stage_opamp_dummy_magic_0.Vb1.t7 two_stage_opamp_dummy_magic_0.VD1.t10 GNDA.t344 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X57 VOUT+.t24 two_stage_opamp_dummy_magic_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X58 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 two_stage_opamp_dummy_magic_0.X.t28 GNDA.t113 VDDA.t187 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X59 VDDA.t83 bgr_0.1st_Vout_1.t13 bgr_0.V_TOP.t0 VDDA.t82 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X60 bgr_0.V_TOP.t17 VDDA.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 VOUT+.t25 two_stage_opamp_dummy_magic_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X62 GNDA.t26 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 two_stage_opamp_dummy_magic_0.V_source.t20 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X63 GNDA.t38 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 two_stage_opamp_dummy_magic_0.V_source.t19 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X64 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 two_stage_opamp_dummy_magic_0.Y.t27 VDDA.t59 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X65 two_stage_opamp_dummy_magic_0.VD1.t20 VIN-.t0 two_stage_opamp_dummy_magic_0.V_source.t36 GNDA.t321 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X66 GNDA.t302 GNDA.t300 bgr_0.NFET_GATE_10uA.t0 GNDA.t301 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X67 bgr_0.START_UP.t5 bgr_0.V_TOP.t18 VDDA.t76 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X68 two_stage_opamp_dummy_magic_0.V_err_p.t17 two_stage_opamp_dummy_magic_0.V_err_gate.t16 VDDA.t17 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X69 VOUT+.t26 two_stage_opamp_dummy_magic_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X70 two_stage_opamp_dummy_magic_0.V_err_gate.t9 bgr_0.NFET_GATE_10uA.t6 GNDA.t212 GNDA.t211 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X71 bgr_0.1st_Vout_1.t8 bgr_0.Vin+.t7 bgr_0.V_p_1.t8 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X72 VOUT-.t32 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X73 VOUT+.t27 two_stage_opamp_dummy_magic_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 two_stage_opamp_dummy_magic_0.err_amp_out.t9 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 GNDA.t154 GNDA.t153 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X75 VOUT+.t28 two_stage_opamp_dummy_magic_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 VOUT+.t29 two_stage_opamp_dummy_magic_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X77 VOUT-.t33 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X78 bgr_0.1st_Vout_1.t14 bgr_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 two_stage_opamp_dummy_magic_0.VD1.t12 VIN-.t1 two_stage_opamp_dummy_magic_0.V_source.t26 GNDA.t140 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X80 bgr_0.V_TOP.t19 VDDA.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X81 bgr_0.V_mir2.t16 bgr_0.V_mir2.t15 VDDA.t85 VDDA.t84 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X82 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 VDDA.t421 VDDA.t423 VDDA.t422 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X83 VOUT+.t30 two_stage_opamp_dummy_magic_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 bgr_0.PFET_GATE_10uA.t12 VDDA.t247 VDDA.t246 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X85 two_stage_opamp_dummy_magic_0.err_amp_out.t8 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 GNDA.t127 GNDA.t126 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X86 VDDA.t224 bgr_0.PFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 VDDA.t223 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X87 GNDA.t299 GNDA.t297 two_stage_opamp_dummy_magic_0.X.t19 GNDA.t298 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X88 VOUT-.t34 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 bgr_0.V_TOP.t20 VDDA.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X90 bgr_0.1st_Vout_2.t3 bgr_0.V_CUR_REF_REG.t4 bgr_0.V_p_2.t8 GNDA.t96 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X91 two_stage_opamp_dummy_magic_0.Y.t19 GNDA.t294 GNDA.t296 GNDA.t295 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X92 VDDA.t203 two_stage_opamp_dummy_magic_0.X.t29 VOUT+.t9 VDDA.t202 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X93 GNDA.t293 GNDA.t291 two_stage_opamp_dummy_magic_0.VD1.t16 GNDA.t292 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X94 VOUT+.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 two_stage_opamp_dummy_magic_0.VD3.t31 VDDA.t418 VDDA.t420 VDDA.t419 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X96 VOUT+.t32 two_stage_opamp_dummy_magic_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 VOUT+.t0 a_14240_2076.t0 GNDA.t4 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X98 VOUT-.t35 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X99 VOUT+.t33 two_stage_opamp_dummy_magic_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 two_stage_opamp_dummy_magic_0.VD3.t37 two_stage_opamp_dummy_magic_0.VD3.t35 two_stage_opamp_dummy_magic_0.X.t24 two_stage_opamp_dummy_magic_0.VD3.t36 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X101 VDDA.t100 two_stage_opamp_dummy_magic_0.V_err_gate.t17 two_stage_opamp_dummy_magic_0.V_err_p.t16 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X102 VOUT-.t36 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X103 bgr_0.PFET_GATE_10uA.t5 bgr_0.1st_Vout_2.t13 VDDA.t460 VDDA.t459 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X104 GNDA.t290 GNDA.t288 two_stage_opamp_dummy_magic_0.VD1.t15 GNDA.t289 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X105 VOUT+.t34 two_stage_opamp_dummy_magic_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X106 bgr_0.V_TOP.t21 VDDA.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 two_stage_opamp_dummy_magic_0.X.t30 VDDA.t86 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X108 two_stage_opamp_dummy_magic_0.V_source.t18 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 GNDA.t112 GNDA.t111 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X109 bgr_0.START_UP_NFET1.t0 bgr_0.START_UP_NFET1 GNDA.t333 GNDA.t332 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X110 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 two_stage_opamp_dummy_magic_0.X.t31 VDDA.t25 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X111 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t18 VDDA.t102 VDDA.t101 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X112 a_5190_5068.t0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 GNDA.t86 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X113 VOUT-.t37 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 bgr_0.V_TOP.t22 VDDA.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 GNDA.t210 bgr_0.NFET_GATE_10uA.t7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 GNDA.t209 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X116 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 bgr_0.NFET_GATE_10uA.t8 GNDA.t208 GNDA.t207 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X117 VOUT+.t35 two_stage_opamp_dummy_magic_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X118 VOUT+.t36 two_stage_opamp_dummy_magic_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 GNDA.t103 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 two_stage_opamp_dummy_magic_0.V_source.t17 GNDA.t102 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X120 two_stage_opamp_dummy_magic_0.VD3.t29 two_stage_opamp_dummy_magic_0.Vb3.t8 VDDA.t313 VDDA.t312 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X121 VOUT+.t37 two_stage_opamp_dummy_magic_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 VOUT+.t38 two_stage_opamp_dummy_magic_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 VOUT+.t39 two_stage_opamp_dummy_magic_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 bgr_0.1st_Vout_2.t14 bgr_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 VOUT-.t38 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 VOUT-.t39 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X127 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 two_stage_opamp_dummy_magic_0.Y.t28 VDDA.t94 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X128 VOUT-.t40 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 VOUT-.t41 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 GNDA.t101 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X131 GNDA.t317 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 VOUT-.t17 GNDA.t316 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X132 VOUT-.t42 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 a_12530_23988.t0 bgr_0.Vin-.t0 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=6
X134 two_stage_opamp_dummy_magic_0.VD4.t35 two_stage_opamp_dummy_magic_0.Vb3.t9 VDDA.t311 VDDA.t310 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X135 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 two_stage_opamp_dummy_magic_0.Y.t29 GNDA.t59 VDDA.t95 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X136 bgr_0.1st_Vout_2.t2 bgr_0.V_mir2.t18 VDDA.t98 VDDA.t97 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X137 two_stage_opamp_dummy_magic_0.VD4.t21 two_stage_opamp_dummy_magic_0.Vb2.t13 two_stage_opamp_dummy_magic_0.Y.t11 two_stage_opamp_dummy_magic_0.VD4.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X138 VOUT+.t40 two_stage_opamp_dummy_magic_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 two_stage_opamp_dummy_magic_0.VD1.t9 two_stage_opamp_dummy_magic_0.Vb1.t8 two_stage_opamp_dummy_magic_0.X.t16 GNDA.t119 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X140 VOUT+.t41 two_stage_opamp_dummy_magic_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X141 bgr_0.1st_Vout_2.t15 bgr_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X142 two_stage_opamp_dummy_magic_0.Y.t6 two_stage_opamp_dummy_magic_0.Vb1.t9 two_stage_opamp_dummy_magic_0.VD2.t6 GNDA.t88 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X143 VOUT+.t42 two_stage_opamp_dummy_magic_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 VOUT-.t43 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 two_stage_opamp_dummy_magic_0.V_source.t25 VIN+.t0 two_stage_opamp_dummy_magic_0.VD2.t11 GNDA.t139 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X146 VOUT+.t43 two_stage_opamp_dummy_magic_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 VOUT-.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 VOUT-.t45 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 bgr_0.1st_Vout_1.t15 bgr_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 bgr_0.V_mir1.t15 bgr_0.Vin-.t8 bgr_0.V_p_1.t4 GNDA.t173 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X151 bgr_0.V_mir1.t13 bgr_0.V_mir1.t12 VDDA.t61 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X152 GNDA.t74 a_7580_22380.t0 GNDA.t73 sky130_fd_pr__res_xhigh_po_0p35 l=6
X153 GNDA.t99 two_stage_opamp_dummy_magic_0.Y.t30 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 VDDA.t149 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X154 two_stage_opamp_dummy_magic_0.V_source.t37 VIN+.t1 two_stage_opamp_dummy_magic_0.VD2.t18 GNDA.t322 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X155 VOUT+.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X156 VOUT+.t45 two_stage_opamp_dummy_magic_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 VDDA.t151 two_stage_opamp_dummy_magic_0.Y.t31 VOUT-.t8 VDDA.t150 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X158 VOUT-.t46 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 two_stage_opamp_dummy_magic_0.X.t32 VDDA.t438 GNDA.t319 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X160 VOUT+.t46 two_stage_opamp_dummy_magic_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X161 VOUT+.t47 two_stage_opamp_dummy_magic_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 two_stage_opamp_dummy_magic_0.V_source.t23 two_stage_opamp_dummy_magic_0.Vb1.t1 two_stage_opamp_dummy_magic_0.Vb1.t2 GNDA.t72 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=3.1
X163 two_stage_opamp_dummy_magic_0.V_source.t16 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 GNDA.t105 GNDA.t104 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X164 VDDA.t32 bgr_0.PFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_0.Vb1.t0 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X165 two_stage_opamp_dummy_magic_0.VD3.t28 two_stage_opamp_dummy_magic_0.Vb3.t10 VDDA.t309 VDDA.t308 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X166 VOUT+.t48 two_stage_opamp_dummy_magic_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X167 two_stage_opamp_dummy_magic_0.VD4.t19 two_stage_opamp_dummy_magic_0.Vb2.t14 two_stage_opamp_dummy_magic_0.Y.t2 two_stage_opamp_dummy_magic_0.VD4.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X168 bgr_0.V_TOP.t23 VDDA.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X169 VDDA.t417 VDDA.t415 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 VDDA.t416 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X170 VOUT+.t49 two_stage_opamp_dummy_magic_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 VOUT+.t50 two_stage_opamp_dummy_magic_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X172 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 bgr_0.PFET_GATE_10uA.t15 VDDA.t2 VDDA.t1 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X173 GNDA.t287 GNDA.t285 two_stage_opamp_dummy_magic_0.Y.t18 GNDA.t286 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X174 VOUT-.t47 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 VOUT-.t48 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 bgr_0.V_mir1.t1 bgr_0.Vin-.t9 bgr_0.V_p_1.t3 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X177 VOUT-.t49 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X178 GNDA.t109 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 two_stage_opamp_dummy_magic_0.V_source.t15 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X179 VOUT-.t50 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X180 bgr_0.START_UP.t4 bgr_0.V_TOP.t24 VDDA.t142 VDDA.t141 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X181 bgr_0.PFET_GATE_10uA.t4 bgr_0.1st_Vout_2.t16 VDDA.t226 VDDA.t225 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X182 VDDA.t267 bgr_0.V_mir1.t18 bgr_0.1st_Vout_1.t4 VDDA.t266 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X183 VOUT-.t51 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X184 VOUT+.t51 two_stage_opamp_dummy_magic_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 VOUT-.t4 two_stage_opamp_dummy_magic_0.Y.t32 VDDA.t55 VDDA.t54 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X186 VOUT+.t52 two_stage_opamp_dummy_magic_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X187 GNDA.t323 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 two_stage_opamp_dummy_magic_0.V_source.t14 GNDA.t283 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X188 two_stage_opamp_dummy_magic_0.Vb2.t7 bgr_0.NFET_GATE_10uA.t9 GNDA.t206 GNDA.t205 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X189 GNDA.t204 bgr_0.NFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_0.Vb2.t6 GNDA.t203 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X190 VOUT-.t52 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 bgr_0.V_TOP.t25 VDDA.t143 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 GNDA.t202 bgr_0.NFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_0.Vb2.t5 GNDA.t201 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X193 VDDA.t414 VDDA.t412 two_stage_opamp_dummy_magic_0.V_err_p.t21 VDDA.t413 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X194 two_stage_opamp_dummy_magic_0.VD1.t8 two_stage_opamp_dummy_magic_0.Vb1.t10 two_stage_opamp_dummy_magic_0.X.t3 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X195 VOUT-.t53 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 VOUT+.t53 two_stage_opamp_dummy_magic_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 two_stage_opamp_dummy_magic_0.err_amp_out.t4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 two_stage_opamp_dummy_magic_0.V_err_p.t1 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X198 VOUT-.t54 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 VOUT-.t55 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X200 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 a_14240_2076.t1 GNDA.t17 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X201 VDDA.t307 two_stage_opamp_dummy_magic_0.Vb3.t11 two_stage_opamp_dummy_magic_0.VD3.t27 VDDA.t306 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X202 GNDA.t107 two_stage_opamp_dummy_magic_0.X.t33 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 VDDA.t156 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X203 VOUT-.t56 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X204 two_stage_opamp_dummy_magic_0.V_source.t13 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 GNDA.t24 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X205 VDDA.t145 bgr_0.V_TOP.t26 bgr_0.Vin+.t4 VDDA.t144 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X206 bgr_0.1st_Vout_2.t5 bgr_0.V_mir2.t19 VDDA.t155 VDDA.t154 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X207 bgr_0.V_TOP.t1 bgr_0.1st_Vout_1.t16 VDDA.t158 VDDA.t157 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X208 bgr_0.V_CUR_REF_REG.t2 VDDA.t409 VDDA.t411 VDDA.t410 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X209 two_stage_opamp_dummy_magic_0.VD4.t5 two_stage_opamp_dummy_magic_0.VD4.t3 two_stage_opamp_dummy_magic_0.Y.t17 two_stage_opamp_dummy_magic_0.VD4.t4 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X210 VDDA.t305 two_stage_opamp_dummy_magic_0.Vb3.t12 two_stage_opamp_dummy_magic_0.VD4.t34 VDDA.t304 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X211 VOUT+.t54 two_stage_opamp_dummy_magic_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 VOUT+.t55 two_stage_opamp_dummy_magic_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 VOUT+.t56 two_stage_opamp_dummy_magic_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X214 VOUT-.t57 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X215 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 bgr_0.PFET_GATE_10uA.t16 VDDA.t222 VDDA.t221 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X216 VOUT+.t57 two_stage_opamp_dummy_magic_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 two_stage_opamp_dummy_magic_0.V_source.t2 VIN+.t2 two_stage_opamp_dummy_magic_0.VD2.t2 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X218 VOUT-.t58 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X219 GNDA.t39 two_stage_opamp_dummy_magic_0.Y.t33 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X220 two_stage_opamp_dummy_magic_0.V_source.t24 VIN-.t2 two_stage_opamp_dummy_magic_0.VD1.t11 GNDA.t138 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X221 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 GNDA.t282 GNDA.t284 GNDA.t283 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X222 VOUT-.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 VOUT-.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X224 bgr_0.1st_Vout_2.t17 bgr_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X225 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 two_stage_opamp_dummy_magic_0.V_err_gate.t3 VDDA.t148 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X226 two_stage_opamp_dummy_magic_0.V_source.t12 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 GNDA.t136 GNDA.t135 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X227 bgr_0.Vin+.t1 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 GNDA.t120 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X228 VOUT-.t61 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 VOUT-.t62 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 VOUT+.t58 two_stage_opamp_dummy_magic_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X231 VOUT+.t59 two_stage_opamp_dummy_magic_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 bgr_0.1st_Vout_2.t18 bgr_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X233 bgr_0.Vin+.t3 bgr_0.V_TOP.t27 VDDA.t164 VDDA.t163 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X234 VDDA.t303 two_stage_opamp_dummy_magic_0.Vb3.t13 two_stage_opamp_dummy_magic_0.VD3.t26 VDDA.t302 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X235 VDDA.t408 VDDA.t406 bgr_0.PFET_GATE_10uA.t9 VDDA.t407 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X236 VOUT+.t8 two_stage_opamp_dummy_magic_0.X.t34 VDDA.t452 VDDA.t451 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X237 two_stage_opamp_dummy_magic_0.VD2.t4 two_stage_opamp_dummy_magic_0.Vb1.t11 two_stage_opamp_dummy_magic_0.Y.t4 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X238 VOUT-.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 VDDA.t166 bgr_0.V_TOP.t28 bgr_0.Vin+.t2 VDDA.t165 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X240 VOUT-.t64 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 GNDA.t354 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 two_stage_opamp_dummy_magic_0.V_source.t11 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X242 bgr_0.1st_Vout_1.t17 bgr_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X243 GNDA.t347 a_12410_22380.t1 GNDA.t346 sky130_fd_pr__res_xhigh_po_0p35 l=6
X244 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 two_stage_opamp_dummy_magic_0.Y.t34 VDDA.t3 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X245 GNDA.t200 bgr_0.NFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_0.Vb3.t7 GNDA.t199 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X246 two_stage_opamp_dummy_magic_0.V_err_p.t20 VDDA.t403 VDDA.t405 VDDA.t404 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X247 VOUT+.t60 two_stage_opamp_dummy_magic_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X248 VOUT+.t61 two_stage_opamp_dummy_magic_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X249 VDDA.t301 two_stage_opamp_dummy_magic_0.Vb3.t14 two_stage_opamp_dummy_magic_0.VD4.t33 VDDA.t300 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X250 VOUT-.t65 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X251 VOUT-.t66 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X252 VOUT+.t62 two_stage_opamp_dummy_magic_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 bgr_0.cap_res1.t0 bgr_0.V_TOP.t2 GNDA.t125 sky130_fd_pr__res_high_po_0p35 l=2.05
X254 two_stage_opamp_dummy_magic_0.Vb3.t6 bgr_0.NFET_GATE_10uA.t13 GNDA.t198 GNDA.t197 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X255 bgr_0.V_mir2.t14 bgr_0.V_mir2.t13 VDDA.t250 VDDA.t249 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X256 VOUT+.t63 two_stage_opamp_dummy_magic_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X257 VDDA.t402 VDDA.t400 bgr_0.V_TOP.t12 VDDA.t401 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X258 VOUT-.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X259 VOUT-.t68 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X260 VDDA.t299 two_stage_opamp_dummy_magic_0.Vb3.t15 two_stage_opamp_dummy_magic_0.VD3.t25 VDDA.t298 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X261 VOUT-.t0 two_stage_opamp_dummy_magic_0.Y.t35 VDDA.t5 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X262 bgr_0.1st_Vout_1.t18 bgr_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 two_stage_opamp_dummy_magic_0.Y.t12 two_stage_opamp_dummy_magic_0.Vb2.t15 two_stage_opamp_dummy_magic_0.VD4.t17 two_stage_opamp_dummy_magic_0.VD4.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X264 VOUT+.t64 two_stage_opamp_dummy_magic_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 VOUT-.t69 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 bgr_0.V_TOP.t29 VDDA.t168 VDDA.t167 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X267 VDDA.t104 two_stage_opamp_dummy_magic_0.V_err_gate.t19 two_stage_opamp_dummy_magic_0.V_err_p.t15 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X268 bgr_0.1st_Vout_2.t19 bgr_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 sky130_fd_pr__pfet_01v8 ad=1.44 pd=8 as=0 ps=0 w=3.6 l=0.2
X270 VOUT+.t65 two_stage_opamp_dummy_magic_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 GNDA.t34 a_13060_22630.t0 GNDA.t33 sky130_fd_pr__res_xhigh_po_0p35 l=4
X272 VDDA.t106 two_stage_opamp_dummy_magic_0.V_err_gate.t20 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X273 two_stage_opamp_dummy_magic_0.VD1.t7 two_stage_opamp_dummy_magic_0.Vb1.t12 two_stage_opamp_dummy_magic_0.X.t22 GNDA.t330 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X274 VOUT-.t70 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X275 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 two_stage_opamp_dummy_magic_0.V_tot.t5 two_stage_opamp_dummy_magic_0.V_err_p.t0 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X276 bgr_0.1st_Vout_1.t3 bgr_0.V_mir1.t19 VDDA.t269 VDDA.t268 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X277 GNDA.t326 two_stage_opamp_dummy_magic_0.X.t35 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 VDDA.t444 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X278 bgr_0.1st_Vout_1.t19 bgr_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X279 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 VIN+.t3 two_stage_opamp_dummy_magic_0.V_p_mir.t3 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X280 two_stage_opamp_dummy_magic_0.V_source.t27 VIN-.t3 two_stage_opamp_dummy_magic_0.VD1.t13 GNDA.t142 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X281 VOUT+.t66 two_stage_opamp_dummy_magic_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X282 VDDA.t113 two_stage_opamp_dummy_magic_0.Y.t36 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 GNDA.t75 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X283 VOUT-.t71 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 VOUT+.t67 two_stage_opamp_dummy_magic_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X285 VOUT+.t68 two_stage_opamp_dummy_magic_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 bgr_0.NFET_GATE_10uA.t4 bgr_0.PFET_GATE_10uA.t17 VDDA.t441 VDDA.t440 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X287 VDDA.t93 bgr_0.PFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X288 VOUT-.t72 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X289 VOUT-.t73 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X290 bgr_0.1st_Vout_1.t20 bgr_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X291 bgr_0.V_p_2.t2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 bgr_0.V_mir2.t4 GNDA.t82 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X292 two_stage_opamp_dummy_magic_0.V_source.t40 VIN-.t4 two_stage_opamp_dummy_magic_0.VD1.t21 GNDA.t350 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X293 two_stage_opamp_dummy_magic_0.Y.t16 two_stage_opamp_dummy_magic_0.Vb2.t16 two_stage_opamp_dummy_magic_0.VD4.t15 two_stage_opamp_dummy_magic_0.VD4.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X294 VDDA.t297 two_stage_opamp_dummy_magic_0.Vb3.t16 two_stage_opamp_dummy_magic_0.VD3.t24 VDDA.t296 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X295 GNDA.t76 two_stage_opamp_dummy_magic_0.Y.t37 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 VDDA.t114 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X296 VDDA.t138 bgr_0.V_TOP.t30 bgr_0.START_UP.t3 VDDA.t137 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X297 two_stage_opamp_dummy_magic_0.VD4.t37 VDDA.t397 VDDA.t399 VDDA.t398 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X298 GNDA.t149 two_stage_opamp_dummy_magic_0.Y.t38 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 VDDA.t238 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X299 VOUT-.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 VOUT+.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 VOUT+.t70 two_stage_opamp_dummy_magic_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 two_stage_opamp_dummy_magic_0.V_tot.t6 two_stage_opamp_dummy_magic_0.V_err_gate.t13 VDDA.t450 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X303 VOUT-.t75 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 VOUT-.t76 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X305 bgr_0.V_TOP.t31 VDDA.t139 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X306 bgr_0.V_TOP.t7 bgr_0.1st_Vout_1.t21 VDDA.t257 VDDA.t256 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X307 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 two_stage_opamp_dummy_magic_0.V_tot.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t6 VDDA.t112 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X308 VOUT+.t1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 GNDA.t7 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X309 VOUT+.t7 two_stage_opamp_dummy_magic_0.X.t36 VDDA.t160 VDDA.t159 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X310 VOUT-.t77 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X311 VOUT+.t71 two_stage_opamp_dummy_magic_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X312 VOUT+.t72 two_stage_opamp_dummy_magic_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 VOUT+.t73 two_stage_opamp_dummy_magic_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 VOUT+.t74 two_stage_opamp_dummy_magic_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 bgr_0.V_TOP.t8 bgr_0.1st_Vout_1.t22 VDDA.t259 VDDA.t258 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X316 VOUT-.t78 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 VOUT-.t79 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 VOUT-.t80 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 bgr_0.NFET_GATE_10uA.t2 bgr_0.NFET_GATE_10uA.t1 GNDA.t196 GNDA.t195 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X320 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 two_stage_opamp_dummy_magic_0.V_err_gate.t21 VDDA.t178 VDDA.t177 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X321 GNDA.t194 bgr_0.NFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_0.Vb3.t5 GNDA.t193 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X322 VOUT-.t81 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 bgr_0.V_TOP.t32 VDDA.t140 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X324 two_stage_opamp_dummy_magic_0.VD3.t19 two_stage_opamp_dummy_magic_0.Vb2.t17 two_stage_opamp_dummy_magic_0.X.t10 two_stage_opamp_dummy_magic_0.VD3.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X325 VOUT-.t10 two_stage_opamp_dummy_magic_0.Y.t39 VDDA.t240 VDDA.t239 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X326 VOUT-.t6 two_stage_opamp_dummy_magic_0.Y.t40 VDDA.t80 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X327 bgr_0.1st_Vout_2.t20 bgr_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 VDDA.t87 two_stage_opamp_dummy_magic_0.X.t37 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X329 VOUT+.t75 two_stage_opamp_dummy_magic_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 VOUT+.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X331 VOUT+.t14 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 GNDA.t160 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X332 VOUT-.t82 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X333 VDDA.t180 two_stage_opamp_dummy_magic_0.V_err_gate.t22 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 VDDA.t179 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X334 two_stage_opamp_dummy_magic_0.VD3.t23 two_stage_opamp_dummy_magic_0.Vb3.t17 VDDA.t295 VDDA.t294 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X335 VDDA.t212 bgr_0.PFET_GATE_10uA.t19 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 VDDA.t211 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X336 VOUT+.t77 two_stage_opamp_dummy_magic_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X337 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 two_stage_opamp_dummy_magic_0.V_tot.t8 two_stage_opamp_dummy_magic_0.V_err_p.t19 VDDA.t197 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X338 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 GNDA.t353 GNDA.t352 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X339 two_stage_opamp_dummy_magic_0.VD1.t6 two_stage_opamp_dummy_magic_0.Vb1.t13 two_stage_opamp_dummy_magic_0.X.t0 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X340 bgr_0.1st_Vout_1.t23 bgr_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X341 bgr_0.V_mir1.t11 bgr_0.V_mir1.t10 VDDA.t22 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X342 VDDA.t134 bgr_0.V_TOP.t33 bgr_0.START_UP.t2 VDDA.t133 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X343 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_0.Y.t1 GNDA.t12 sky130_fd_pr__res_high_po_1p41 l=1.41
X344 two_stage_opamp_dummy_magic_0.err_amp_out.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 two_stage_opamp_dummy_magic_0.V_err_p.t3 VDDA.t121 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X345 VOUT+.t78 two_stage_opamp_dummy_magic_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X346 bgr_0.1st_Vout_2.t21 bgr_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X347 GNDA.t132 two_stage_opamp_dummy_magic_0.X.t38 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 VDDA.t230 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X348 VOUT+.t79 two_stage_opamp_dummy_magic_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X349 VOUT-.t83 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 VOUT-.t84 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 two_stage_opamp_dummy_magic_0.V_source.t28 VIN+.t4 two_stage_opamp_dummy_magic_0.VD2.t13 GNDA.t161 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X352 VOUT-.t85 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X353 a_6810_23838.t0 a_6930_22590.t1 GNDA.t137 sky130_fd_pr__res_xhigh_po_0p35 l=4.2
X354 a_7460_23988.t1 a_7580_22380.t1 GNDA.t141 sky130_fd_pr__res_xhigh_po_0p35 l=6
X355 bgr_0.V_p_2.t7 bgr_0.V_CUR_REF_REG.t5 bgr_0.1st_Vout_2.t4 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X356 two_stage_opamp_dummy_magic_0.VD4.t32 two_stage_opamp_dummy_magic_0.Vb3.t18 VDDA.t293 VDDA.t292 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X357 VDDA.t81 two_stage_opamp_dummy_magic_0.Y.t41 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X358 VOUT+.t80 two_stage_opamp_dummy_magic_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 GNDA.t281 GNDA.t279 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 GNDA.t280 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X360 two_stage_opamp_dummy_magic_0.V_source.t39 VIN+.t5 two_stage_opamp_dummy_magic_0.VD2.t20 GNDA.t339 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X361 bgr_0.1st_Vout_2.t22 bgr_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X362 GNDA.t131 two_stage_opamp_dummy_magic_0.Y.t42 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 VDDA.t216 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X363 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 VDDA.t394 VDDA.t396 VDDA.t395 sky130_fd_pr__pfet_01v8 ad=0.71 pd=3.95 as=1.42 ps=7.9 w=3.55 l=0.2
X364 bgr_0.1st_Vout_1.t9 bgr_0.Vin+.t8 bgr_0.V_p_1.t7 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X365 VDDA.t39 bgr_0.V_mir2.t20 bgr_0.1st_Vout_2.t0 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X366 VOUT+.t81 two_stage_opamp_dummy_magic_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X367 VOUT+.t82 two_stage_opamp_dummy_magic_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X368 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 two_stage_opamp_dummy_magic_0.V_err_gate.t2 VDDA.t119 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X369 bgr_0.1st_Vout_1.t24 bgr_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X370 GNDA.t219 GNDA.t278 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X371 VOUT+.t83 two_stage_opamp_dummy_magic_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 bgr_0.1st_Vout_2.t23 bgr_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 VOUT+.t84 two_stage_opamp_dummy_magic_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X374 GNDA.t192 bgr_0.NFET_GATE_10uA.t15 two_stage_opamp_dummy_magic_0.Vb2.t4 GNDA.t191 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X375 two_stage_opamp_dummy_magic_0.Vb2.t3 bgr_0.NFET_GATE_10uA.t16 GNDA.t190 GNDA.t189 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X376 two_stage_opamp_dummy_magic_0.VD2.t9 two_stage_opamp_dummy_magic_0.Vb1.t14 two_stage_opamp_dummy_magic_0.Y.t9 GNDA.t118 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X377 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 GNDA.t271 GNDA.t273 GNDA.t272 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X378 VOUT-.t86 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 GNDA.t219 GNDA.t277 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X380 GNDA.t276 GNDA.t274 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 GNDA.t275 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X381 GNDA.t270 GNDA.t268 two_stage_opamp_dummy_magic_0.Vb2.t9 GNDA.t269 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X382 VOUT+.t85 two_stage_opamp_dummy_magic_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 VOUT+.t6 two_stage_opamp_dummy_magic_0.X.t39 VDDA.t189 VDDA.t188 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X384 VOUT-.t87 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X385 bgr_0.PFET_GATE_10uA.t8 VDDA.t391 VDDA.t393 VDDA.t392 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X386 two_stage_opamp_dummy_magic_0.VD4.t31 two_stage_opamp_dummy_magic_0.Vb3.t19 VDDA.t291 VDDA.t290 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X387 bgr_0.1st_Vout_1.t2 bgr_0.V_mir1.t20 VDDA.t263 VDDA.t262 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X388 VOUT+.t86 two_stage_opamp_dummy_magic_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X389 two_stage_opamp_dummy_magic_0.V_err_p.t14 two_stage_opamp_dummy_magic_0.V_err_gate.t23 VDDA.t184 VDDA.t183 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X390 bgr_0.V_p_2.t6 bgr_0.V_CUR_REF_REG.t6 bgr_0.1st_Vout_2.t8 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X391 two_stage_opamp_dummy_magic_0.VD4.t13 two_stage_opamp_dummy_magic_0.Vb2.t18 two_stage_opamp_dummy_magic_0.Y.t10 two_stage_opamp_dummy_magic_0.VD4.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X392 VOUT+.t87 two_stage_opamp_dummy_magic_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X393 GNDA.t45 VDDA.t469 bgr_0.V_p_2.t10 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X394 VOUT-.t88 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X395 GNDA.t219 GNDA.t220 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X396 VOUT+.t88 two_stage_opamp_dummy_magic_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X397 two_stage_opamp_dummy_magic_0.Vb3.t1 two_stage_opamp_dummy_magic_0.Vb2.t19 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4 as=0.72 ps=4 w=3.6 l=0.2
X398 VOUT-.t9 two_stage_opamp_dummy_magic_0.Y.t43 VDDA.t218 VDDA.t217 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X399 VOUT-.t89 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 VDDA.t456 two_stage_opamp_dummy_magic_0.X.t40 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA.t342 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X401 GNDA.t219 GNDA.t267 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X402 VOUT+.t89 two_stage_opamp_dummy_magic_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 VDDA.t186 two_stage_opamp_dummy_magic_0.V_err_gate.t24 two_stage_opamp_dummy_magic_0.V_err_p.t13 VDDA.t185 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X404 VDDA.t199 bgr_0.V_mir2.t11 bgr_0.V_mir2.t12 VDDA.t198 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X405 two_stage_opamp_dummy_magic_0.err_amp_out.t2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 two_stage_opamp_dummy_magic_0.V_err_p.t4 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X406 two_stage_opamp_dummy_magic_0.err_amp_out.t10 GNDA.t264 GNDA.t266 GNDA.t265 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X407 two_stage_opamp_dummy_magic_0.VD1.t5 two_stage_opamp_dummy_magic_0.Vb1.t15 two_stage_opamp_dummy_magic_0.X.t17 GNDA.t145 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X408 GNDA.t327 two_stage_opamp_dummy_magic_0.X.t41 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 VDDA.t445 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X409 VOUT-.t90 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 VOUT-.t91 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 GNDA.t151 two_stage_opamp_dummy_magic_0.X.t42 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 VDDA.t242 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X412 bgr_0.V_p_2.t5 bgr_0.V_CUR_REF_REG.t7 bgr_0.1st_Vout_2.t9 GNDA.t345 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X413 VOUT-.t92 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 two_stage_opamp_dummy_magic_0.V_source.t38 two_stage_opamp_dummy_magic_0.err_amp_out.t12 GNDA.t325 GNDA.t324 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X415 VDDA.t71 two_stage_opamp_dummy_magic_0.Y.t44 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X416 two_stage_opamp_dummy_magic_0.V_source.t30 VIN-.t5 two_stage_opamp_dummy_magic_0.VD1.t14 GNDA.t164 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X417 a_13180_23838.t0 bgr_0.V_CUR_REF_REG.t0 GNDA.t30 sky130_fd_pr__res_xhigh_po_0p35 l=4
X418 VDDA.t174 two_stage_opamp_dummy_magic_0.V_err_gate.t25 two_stage_opamp_dummy_magic_0.V_err_p.t12 VDDA.t173 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X419 VDDA.t72 two_stage_opamp_dummy_magic_0.Y.t45 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X420 GNDA.t166 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 VOUT-.t11 GNDA.t165 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X421 two_stage_opamp_dummy_magic_0.VD3.t22 two_stage_opamp_dummy_magic_0.Vb3.t20 VDDA.t289 VDDA.t288 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X422 VOUT+.t90 two_stage_opamp_dummy_magic_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 bgr_0.V_TOP.t34 VDDA.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X424 two_stage_opamp_dummy_magic_0.X.t2 two_stage_opamp_dummy_magic_0.VD3.t32 two_stage_opamp_dummy_magic_0.VD3.t34 two_stage_opamp_dummy_magic_0.VD3.t33 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X425 GNDA.t129 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 two_stage_opamp_dummy_magic_0.err_amp_out.t7 GNDA.t128 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X426 VOUT+.t91 two_stage_opamp_dummy_magic_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 VOUT+.t92 two_stage_opamp_dummy_magic_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 VOUT+.t93 two_stage_opamp_dummy_magic_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X429 VOUT+.t94 two_stage_opamp_dummy_magic_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X430 VOUT+.t95 two_stage_opamp_dummy_magic_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 GNDA.t64 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 VOUT+.t12 GNDA.t63 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X432 VOUT-.t93 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 bgr_0.V_TOP.t35 VDDA.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 VDDA.t192 bgr_0.1st_Vout_2.t24 bgr_0.PFET_GATE_10uA.t3 VDDA.t191 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X435 VDDA.t390 VDDA.t388 two_stage_opamp_dummy_magic_0.Vb1.t4 VDDA.t389 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X436 VOUT-.t94 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 two_stage_opamp_dummy_magic_0.Vb1.t3 VDDA.t385 VDDA.t387 VDDA.t386 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X438 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 two_stage_opamp_dummy_magic_0.V_err_gate.t26 VDDA.t176 VDDA.t175 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X439 VOUT+.t96 two_stage_opamp_dummy_magic_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 two_stage_opamp_dummy_magic_0.V_tot.t9 two_stage_opamp_dummy_magic_0.V_err_gate.t7 VDDA.t251 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X441 VOUT-.t95 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X442 VOUT-.t96 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X443 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 bgr_0.PFET_GATE_10uA.t20 VDDA.t245 VDDA.t244 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X444 VOUT+.t97 two_stage_opamp_dummy_magic_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 VOUT+.t98 two_stage_opamp_dummy_magic_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X446 GNDA.t259 GNDA.t257 VOUT-.t13 GNDA.t258 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X447 VDDA.t449 bgr_0.PFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 VDDA.t448 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X448 two_stage_opamp_dummy_magic_0.VD2.t10 two_stage_opamp_dummy_magic_0.Vb1.t16 two_stage_opamp_dummy_magic_0.Y.t14 GNDA.t134 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X449 VOUT+.t5 two_stage_opamp_dummy_magic_0.X.t43 VDDA.t466 VDDA.t465 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X450 VOUT+.t4 two_stage_opamp_dummy_magic_0.X.t44 VDDA.t205 VDDA.t204 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X451 VOUT+.t99 two_stage_opamp_dummy_magic_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 bgr_0.V_TOP.t36 VDDA.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X453 VOUT+.t100 two_stage_opamp_dummy_magic_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X454 two_stage_opamp_dummy_magic_0.X.t4 two_stage_opamp_dummy_magic_0.Vb2.t20 two_stage_opamp_dummy_magic_0.VD3.t17 two_stage_opamp_dummy_magic_0.VD3.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X455 bgr_0.Vin-.t6 bgr_0.V_TOP.t37 VDDA.t130 VDDA.t129 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X456 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t27 VDDA.t48 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X457 VOUT+.t101 two_stage_opamp_dummy_magic_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X458 VOUT-.t97 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 VOUT-.t98 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 VOUT-.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 GNDA.t263 GNDA.t260 GNDA.t262 GNDA.t261 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X462 GNDA.t188 bgr_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 GNDA.t187 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X463 bgr_0.1st_Vout_1.t1 bgr_0.V_mir1.t21 VDDA.t265 VDDA.t264 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X464 GNDA.t315 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 two_stage_opamp_dummy_magic_0.V_source.t10 GNDA.t314 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X465 two_stage_opamp_dummy_magic_0.Vb2.t8 GNDA.t254 GNDA.t256 GNDA.t255 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X466 VDDA.t88 two_stage_opamp_dummy_magic_0.X.t45 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X467 VOUT-.t100 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X468 VOUT-.t101 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X469 bgr_0.1st_Vout_1.t25 bgr_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 two_stage_opamp_dummy_magic_0.V_err_gate.t1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 VDDA.t146 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X471 VOUT+.t102 two_stage_opamp_dummy_magic_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 bgr_0.1st_Vout_2.t25 bgr_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X473 VDDA.t50 two_stage_opamp_dummy_magic_0.V_err_gate.t28 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X474 VOUT-.t102 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X475 VDDA.t287 two_stage_opamp_dummy_magic_0.Vb3.t21 two_stage_opamp_dummy_magic_0.VD4.t30 VDDA.t286 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X476 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 VDDA.t382 VDDA.t384 VDDA.t383 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X477 GNDA.t168 VDDA.t379 VDDA.t381 VDDA.t380 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X478 bgr_0.1st_Vout_1.t26 bgr_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X479 two_stage_opamp_dummy_magic_0.V_source.t9 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 GNDA.t335 GNDA.t334 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X480 VOUT+.t103 two_stage_opamp_dummy_magic_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X481 VOUT+.t104 two_stage_opamp_dummy_magic_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 VOUT+.t105 two_stage_opamp_dummy_magic_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 two_stage_opamp_dummy_magic_0.V_source.t1 VIN+.t6 two_stage_opamp_dummy_magic_0.VD2.t1 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X484 VDDA.t126 two_stage_opamp_dummy_magic_0.Y.t46 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 GNDA.t84 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X485 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 bgr_0.PFET_GATE_10uA.t22 VDDA.t458 VDDA.t457 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X486 VOUT+.t106 two_stage_opamp_dummy_magic_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X487 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 bgr_0.V_TOP.t38 VDDA.t132 VDDA.t131 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X488 VOUT-.t103 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X489 VDDA.t70 bgr_0.V_mir2.t9 bgr_0.V_mir2.t10 VDDA.t69 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X490 GNDA.t156 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 GNDA.t155 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X491 VOUT-.t104 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X492 VDDA.t65 bgr_0.V_mir1.t8 bgr_0.V_mir1.t9 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X493 VDDA.t194 bgr_0.PFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 VDDA.t193 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X494 VDDA.t283 two_stage_opamp_dummy_magic_0.Vb3.t22 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 VDDA.t282 sky130_fd_pr__pfet_01v8 ad=0.71 pd=3.95 as=0.71 ps=3.95 w=3.55 l=0.2
X495 bgr_0.V_p_1.t2 bgr_0.Vin-.t10 bgr_0.V_mir1.t0 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X496 VOUT-.t105 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X497 bgr_0.1st_Vout_1.t27 bgr_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 bgr_0.1st_Vout_2.t26 bgr_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X499 VOUT-.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X500 bgr_0.V_TOP.t11 VDDA.t376 VDDA.t378 VDDA.t377 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X501 GNDA.t158 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 GNDA.t157 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X502 two_stage_opamp_dummy_magic_0.X.t21 two_stage_opamp_dummy_magic_0.Vb1.t17 two_stage_opamp_dummy_magic_0.VD1.t4 GNDA.t329 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X503 VDDA.t285 two_stage_opamp_dummy_magic_0.Vb3.t23 two_stage_opamp_dummy_magic_0.VD4.t29 VDDA.t284 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X504 two_stage_opamp_dummy_magic_0.X.t13 two_stage_opamp_dummy_magic_0.Vb2.t21 two_stage_opamp_dummy_magic_0.VD3.t15 two_stage_opamp_dummy_magic_0.VD3.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X505 VOUT-.t107 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X506 bgr_0.1st_Vout_1.t28 bgr_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X507 VOUT+.t107 two_stage_opamp_dummy_magic_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X508 VOUT+.t18 VDDA.t373 VDDA.t375 VDDA.t374 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X509 two_stage_opamp_dummy_magic_0.VD2.t21 two_stage_opamp_dummy_magic_0.Vb1.t18 two_stage_opamp_dummy_magic_0.Y.t24 GNDA.t343 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X510 VDDA.t372 VDDA.t370 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 VDDA.t371 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X511 VOUT+.t108 two_stage_opamp_dummy_magic_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X512 VOUT+.t109 two_stage_opamp_dummy_magic_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X513 VOUT-.t12 GNDA.t251 GNDA.t253 GNDA.t252 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X514 two_stage_opamp_dummy_magic_0.VD1.t0 VIN-.t6 two_stage_opamp_dummy_magic_0.V_source.t21 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X515 bgr_0.V_p_1.t1 bgr_0.Vin-.t11 bgr_0.V_mir1.t16 GNDA.t174 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X516 VOUT-.t108 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X517 VOUT-.t109 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X518 VOUT+.t110 two_stage_opamp_dummy_magic_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X519 VOUT-.t110 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X520 VOUT-.t111 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X521 VOUT-.t112 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X522 bgr_0.1st_Vout_1.t29 bgr_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 two_stage_opamp_dummy_magic_0.Vb3.t0 GNDA.t248 GNDA.t250 GNDA.t249 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X524 VOUT-.t113 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 bgr_0.Vin-.t1 bgr_0.START_UP.t6 bgr_0.V_TOP.t3 VDDA.t227 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X526 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 two_stage_opamp_dummy_magic_0.Vb3.t2 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 sky130_fd_pr__pfet_01v8 ad=1.44 pd=8 as=0.72 ps=4 w=3.6 l=0.2
X527 bgr_0.V_TOP.t4 bgr_0.START_UP.t7 bgr_0.Vin-.t2 VDDA.t248 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X528 two_stage_opamp_dummy_magic_0.VD1.t19 VIN-.t7 two_stage_opamp_dummy_magic_0.V_source.t35 GNDA.t318 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X529 VOUT+.t111 two_stage_opamp_dummy_magic_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X530 VOUT-.t114 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X531 VOUT-.t115 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 VDDA.t28 bgr_0.1st_Vout_2.t27 bgr_0.PFET_GATE_10uA.t2 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X533 bgr_0.V_mir1.t7 bgr_0.V_mir1.t6 VDDA.t437 VDDA.t436 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X534 VDDA.t439 two_stage_opamp_dummy_magic_0.X.t46 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 GNDA.t320 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X535 VOUT+.t112 two_stage_opamp_dummy_magic_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X536 VOUT+.t113 two_stage_opamp_dummy_magic_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X537 GNDA.t349 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 two_stage_opamp_dummy_magic_0.V_source.t8 GNDA.t348 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X538 VDDA.t231 two_stage_opamp_dummy_magic_0.X.t47 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 GNDA.t133 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X539 GNDA.t219 GNDA.t218 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X540 bgr_0.START_UP.t1 bgr_0.START_UP.t0 bgr_0.START_UP_NFET1.t0 GNDA.t162 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X541 VOUT-.t16 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 GNDA.t313 GNDA.t312 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X542 bgr_0.V_p_2.t0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 bgr_0.V_mir2.t3 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X543 two_stage_opamp_dummy_magic_0.cap_res_X.t0 two_stage_opamp_dummy_magic_0.X.t1 GNDA.t71 sky130_fd_pr__res_high_po_1p41 l=1.41
X544 VOUT-.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X545 VOUT+.t114 two_stage_opamp_dummy_magic_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X546 VOUT-.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 VOUT-.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X548 VDDA.t369 VDDA.t367 two_stage_opamp_dummy_magic_0.VD3.t30 VDDA.t368 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X549 VOUT+.t115 two_stage_opamp_dummy_magic_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X550 bgr_0.1st_Vout_2.t28 bgr_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X551 two_stage_opamp_dummy_magic_0.V_source.t7 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 GNDA.t122 GNDA.t121 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X552 two_stage_opamp_dummy_magic_0.VD3.t13 two_stage_opamp_dummy_magic_0.Vb2.t22 two_stage_opamp_dummy_magic_0.X.t7 two_stage_opamp_dummy_magic_0.VD3.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X553 VOUT-.t119 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X554 VDDA.t220 bgr_0.PFET_GATE_10uA.t24 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 VDDA.t219 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X555 VDDA.t435 bgr_0.V_mir2.t21 bgr_0.1st_Vout_2.t7 VDDA.t434 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X556 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 bgr_0.PFET_GATE_10uA.t25 VDDA.t30 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X557 VOUT+.t116 two_stage_opamp_dummy_magic_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X558 VOUT+.t117 two_stage_opamp_dummy_magic_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X559 bgr_0.V_p_1.t0 bgr_0.Vin-.t12 bgr_0.V_mir1.t14 GNDA.t167 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X560 GNDA.t219 GNDA.t231 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X561 GNDA.t14 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 two_stage_opamp_dummy_magic_0.err_amp_out.t6 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X562 bgr_0.1st_Vout_2.t29 bgr_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X563 VDDA.t366 VDDA.t364 two_stage_opamp_dummy_magic_0.VD4.t36 VDDA.t365 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X564 VOUT+.t118 two_stage_opamp_dummy_magic_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X565 VOUT+.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X566 VOUT-.t120 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X567 GNDA.t52 VDDA.t361 VDDA.t363 VDDA.t362 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X568 VOUT+.t120 two_stage_opamp_dummy_magic_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X569 VOUT-.t121 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 bgr_0.1st_Vout_1.t30 bgr_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X571 GNDA.t219 GNDA.t230 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X572 VOUT-.t122 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X573 VOUT+.t121 two_stage_opamp_dummy_magic_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X574 VDDA.t360 VDDA.t358 two_stage_opamp_dummy_magic_0.err_amp_out.t11 VDDA.t359 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X575 two_stage_opamp_dummy_magic_0.X.t15 two_stage_opamp_dummy_magic_0.Vb1.t19 two_stage_opamp_dummy_magic_0.VD1.t3 GNDA.t117 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X576 VOUT-.t123 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X577 GNDA.t219 GNDA.t247 bgr_0.Vin-.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X578 VDDA.t357 VDDA.t355 GNDA.t172 VDDA.t356 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X579 VOUT-.t124 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X580 bgr_0.1st_Vout_2.t30 bgr_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X581 two_stage_opamp_dummy_magic_0.VD2.t5 two_stage_opamp_dummy_magic_0.Vb1.t20 two_stage_opamp_dummy_magic_0.Y.t5 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X582 two_stage_opamp_dummy_magic_0.VD3.t11 two_stage_opamp_dummy_magic_0.Vb2.t23 two_stage_opamp_dummy_magic_0.X.t6 two_stage_opamp_dummy_magic_0.VD3.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X583 VOUT-.t125 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X584 GNDA.t186 bgr_0.NFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_0.V_err_gate.t8 GNDA.t185 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X585 bgr_0.Vin-.t5 bgr_0.V_TOP.t39 VDDA.t462 VDDA.t461 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X586 two_stage_opamp_dummy_magic_0.Y.t23 two_stage_opamp_dummy_magic_0.Vb2.t24 two_stage_opamp_dummy_magic_0.VD4.t11 two_stage_opamp_dummy_magic_0.VD4.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X587 a_12530_23988.t1 a_12410_22380.t0 GNDA.t78 sky130_fd_pr__res_xhigh_po_0p35 l=6
X588 two_stage_opamp_dummy_magic_0.Vb3.t3 bgr_0.NFET_GATE_10uA.t19 GNDA.t184 GNDA.t183 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X589 bgr_0.1st_Vout_2.t31 bgr_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X590 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 two_stage_opamp_dummy_magic_0.Y.t47 GNDA.t85 VDDA.t127 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X591 two_stage_opamp_dummy_magic_0.VD2.t0 VIN+.t7 two_stage_opamp_dummy_magic_0.V_source.t0 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X592 VOUT+.t122 two_stage_opamp_dummy_magic_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X593 VDDA.t10 bgr_0.V_mir2.t7 bgr_0.V_mir2.t8 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X594 GNDA.t70 a_6930_22590.t0 GNDA.t69 sky130_fd_pr__res_xhigh_po_0p35 l=4.2
X595 VOUT-.t15 VDDA.t352 VDDA.t354 VDDA.t353 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X596 VDDA.t317 GNDA.t244 GNDA.t246 GNDA.t245 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X597 VOUT-.t126 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X598 bgr_0.1st_Vout_1.t31 bgr_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X599 bgr_0.1st_Vout_2.t32 bgr_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X600 GNDA.t95 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 two_stage_opamp_dummy_magic_0.V_source.t6 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X601 two_stage_opamp_dummy_magic_0.V_err_gate.t5 two_stage_opamp_dummy_magic_0.V_tot.t10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X602 VOUT+.t123 two_stage_opamp_dummy_magic_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X603 two_stage_opamp_dummy_magic_0.VD4.t28 two_stage_opamp_dummy_magic_0.Vb3.t24 VDDA.t281 VDDA.t280 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X604 two_stage_opamp_dummy_magic_0.VD3.t9 two_stage_opamp_dummy_magic_0.Vb2.t25 two_stage_opamp_dummy_magic_0.X.t5 two_stage_opamp_dummy_magic_0.VD3.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X605 VDDA.t351 VDDA.t349 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 VDDA.t350 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X606 VOUT-.t127 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X607 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 bgr_0.PFET_GATE_10uA.t26 VDDA.t162 VDDA.t161 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X608 VOUT+.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X609 VOUT+.t125 two_stage_opamp_dummy_magic_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X610 a_13180_23838.t1 a_13060_22630.t1 GNDA.t115 sky130_fd_pr__res_xhigh_po_0p35 l=4
X611 two_stage_opamp_dummy_magic_0.Y.t7 two_stage_opamp_dummy_magic_0.Vb1.t21 two_stage_opamp_dummy_magic_0.VD2.t7 GNDA.t92 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X612 VDDA.t348 VDDA.t346 VOUT+.t17 VDDA.t347 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X613 VOUT-.t128 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X614 bgr_0.V_p_1.t6 bgr_0.Vin+.t9 bgr_0.1st_Vout_1.t6 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X615 VDDA.t261 bgr_0.V_mir1.t22 bgr_0.1st_Vout_1.t0 VDDA.t260 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X616 two_stage_opamp_dummy_magic_0.V_source.t5 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 GNDA.t50 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X617 VDDA.t345 VDDA.t342 VDDA.t344 VDDA.t343 sky130_fd_pr__pfet_01v8 ad=0.24 pd=2 as=0 ps=0 w=0.6 l=0.2
X618 bgr_0.V_TOP.t40 VDDA.t463 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X619 VDDA.t341 VDDA.t339 VDDA.t341 VDDA.t340 sky130_fd_pr__pfet_01v8 ad=0.71 pd=3.95 as=0 ps=0 w=3.55 l=0.2
X620 VOUT+.t126 two_stage_opamp_dummy_magic_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X621 VOUT+.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X622 VOUT+.t128 two_stage_opamp_dummy_magic_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X623 VDDA.t124 two_stage_opamp_dummy_magic_0.Y.t48 VOUT-.t7 VDDA.t123 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X624 VOUT-.t129 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X625 VOUT+.t129 two_stage_opamp_dummy_magic_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X626 two_stage_opamp_dummy_magic_0.V_source.t4 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 GNDA.t36 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X627 two_stage_opamp_dummy_magic_0.VD3.t7 two_stage_opamp_dummy_magic_0.Vb2.t26 two_stage_opamp_dummy_magic_0.X.t9 two_stage_opamp_dummy_magic_0.VD3.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X628 two_stage_opamp_dummy_magic_0.VD4.t27 two_stage_opamp_dummy_magic_0.Vb3.t25 VDDA.t279 VDDA.t278 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X629 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 a_5710_2076.t0 GNDA.t336 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X630 two_stage_opamp_dummy_magic_0.V_err_p.t11 two_stage_opamp_dummy_magic_0.V_err_gate.t29 VDDA.t41 VDDA.t40 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X631 VOUT-.t130 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X632 VOUT-.t131 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X633 two_stage_opamp_dummy_magic_0.X.t20 two_stage_opamp_dummy_magic_0.Vb1.t22 two_stage_opamp_dummy_magic_0.VD1.t2 GNDA.t328 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X634 bgr_0.V_TOP.t41 VDDA.t464 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X635 bgr_0.V_p_1.t5 bgr_0.Vin+.t10 bgr_0.1st_Vout_1.t7 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X636 VDDA.t338 VDDA.t336 bgr_0.V_TOP.t10 VDDA.t337 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X637 VOUT+.t130 two_stage_opamp_dummy_magic_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X638 two_stage_opamp_dummy_magic_0.Vb2.t2 bgr_0.NFET_GATE_10uA.t20 GNDA.t182 GNDA.t181 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X639 GNDA.t180 bgr_0.NFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 GNDA.t179 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X640 two_stage_opamp_dummy_magic_0.V_err_p.t8 two_stage_opamp_dummy_magic_0.V_tot.t11 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X641 VOUT+.t131 two_stage_opamp_dummy_magic_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X642 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 two_stage_opamp_dummy_magic_0.X.t48 GNDA.t2 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X643 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 bgr_0.NFET_GATE_10uA.t22 GNDA.t178 GNDA.t177 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X644 bgr_0.V_TOP.t42 VDDA.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X645 two_stage_opamp_dummy_magic_0.VD2.t17 VIN+.t8 two_stage_opamp_dummy_magic_0.V_source.t32 GNDA.t309 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X646 GNDA.t243 GNDA.t242 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X647 a_5310_5068.t0 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA.t123 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X648 bgr_0.V_TOP.t43 VDDA.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X649 VOUT+.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X650 VOUT+.t133 two_stage_opamp_dummy_magic_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X651 VDDA.t74 bgr_0.V_mir2.t22 bgr_0.1st_Vout_2.t1 VDDA.t73 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X652 VOUT+.t134 two_stage_opamp_dummy_magic_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X653 VDDA.t255 bgr_0.1st_Vout_1.t32 bgr_0.V_TOP.t6 VDDA.t254 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X654 VOUT-.t132 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X655 VOUT+.t135 two_stage_opamp_dummy_magic_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X656 VOUT+.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X657 two_stage_opamp_dummy_magic_0.VD2.t14 VIN+.t9 two_stage_opamp_dummy_magic_0.V_source.t29 GNDA.t163 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X658 a_14560_5068.t0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 GNDA.t1 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X659 two_stage_opamp_dummy_magic_0.VD3.t21 two_stage_opamp_dummy_magic_0.Vb3.t26 VDDA.t277 VDDA.t276 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X660 VOUT-.t133 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X661 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 two_stage_opamp_dummy_magic_0.Y.t49 GNDA.t83 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X662 VDDA.t335 VDDA.t333 GNDA.t43 VDDA.t334 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X663 GNDA.t90 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 two_stage_opamp_dummy_magic_0.V_p_mir.t0 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X664 two_stage_opamp_dummy_magic_0.V_err_gate.t0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 VDDA.t118 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X665 bgr_0.V_TOP.t44 VDDA.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X666 VDDA.t332 VDDA.t330 two_stage_opamp_dummy_magic_0.Vb2.t10 VDDA.t331 sky130_fd_pr__pfet_01v8 ad=0.24 pd=2 as=0.12 ps=1 w=0.6 l=0.2
X667 two_stage_opamp_dummy_magic_0.X.t8 two_stage_opamp_dummy_magic_0.Vb2.t27 two_stage_opamp_dummy_magic_0.VD3.t5 two_stage_opamp_dummy_magic_0.VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X668 two_stage_opamp_dummy_magic_0.Y.t3 two_stage_opamp_dummy_magic_0.Vb1.t23 two_stage_opamp_dummy_magic_0.VD2.t3 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X669 VDDA.t233 two_stage_opamp_dummy_magic_0.X.t49 VOUT+.t3 VDDA.t232 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X670 bgr_0.V_TOP.t45 VDDA.t207 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X671 bgr_0.V_mir2.t6 bgr_0.V_mir2.t5 VDDA.t12 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X672 VDDA.t37 bgr_0.V_mir1.t4 bgr_0.V_mir1.t5 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X673 VOUT+.t137 two_stage_opamp_dummy_magic_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X674 two_stage_opamp_dummy_magic_0.VD4.t9 two_stage_opamp_dummy_magic_0.Vb2.t28 two_stage_opamp_dummy_magic_0.Y.t21 two_stage_opamp_dummy_magic_0.VD4.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X675 VOUT+.t138 two_stage_opamp_dummy_magic_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X676 two_stage_opamp_dummy_magic_0.V_source.t3 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 GNDA.t79 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X677 VDDA.t316 GNDA.t239 GNDA.t241 GNDA.t240 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X678 VOUT+.t139 two_stage_opamp_dummy_magic_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X679 bgr_0.V_mir2.t2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 bgr_0.V_p_2.t1 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X680 VDDA.t43 two_stage_opamp_dummy_magic_0.V_err_gate.t30 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 VDDA.t42 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X681 VOUT-.t134 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X682 VOUT-.t135 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X683 bgr_0.PFET_GATE_10uA.t7 VDDA.t470 GNDA.t169 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X684 VOUT-.t136 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X685 VDDA.t7 two_stage_opamp_dummy_magic_0.Y.t50 VOUT-.t1 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X686 bgr_0.1st_Vout_1.t33 bgr_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X687 VDDA.t329 VDDA.t327 VOUT-.t14 VDDA.t328 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X688 VOUT+.t140 two_stage_opamp_dummy_magic_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X689 GNDA.t238 GNDA.t236 VDDA.t315 GNDA.t237 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X690 two_stage_opamp_dummy_magic_0.Vb1.t5 bgr_0.PFET_GATE_10uA.t27 VDDA.t447 VDDA.t446 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X691 VDDA.t209 bgr_0.V_TOP.t46 bgr_0.Vin-.t4 VDDA.t208 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X692 VOUT-.t137 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X693 two_stage_opamp_dummy_magic_0.V_err_p.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t31 VDDA.t170 VDDA.t169 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X694 bgr_0.PFET_GATE_10uA.t1 bgr_0.1st_Vout_2.t33 VDDA.t201 VDDA.t200 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X695 two_stage_opamp_dummy_magic_0.X.t14 two_stage_opamp_dummy_magic_0.Vb1.t24 two_stage_opamp_dummy_magic_0.VD1.t1 GNDA.t116 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X696 VOUT-.t138 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X697 VDDA.t454 bgr_0.PFET_GATE_10uA.t28 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 VDDA.t453 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X698 two_stage_opamp_dummy_magic_0.V_err_p.t7 two_stage_opamp_dummy_magic_0.V_tot.t12 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X699 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 VDDA.t324 VDDA.t326 VDDA.t325 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X700 two_stage_opamp_dummy_magic_0.V_err_p.t2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 two_stage_opamp_dummy_magic_0.err_amp_out.t1 VDDA.t117 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X701 VOUT+.t141 two_stage_opamp_dummy_magic_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X702 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 two_stage_opamp_dummy_magic_0.X.t50 GNDA.t20 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X703 a_14680_5068.t0 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA.t106 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X704 two_stage_opamp_dummy_magic_0.VD4.t7 two_stage_opamp_dummy_magic_0.Vb2.t29 two_stage_opamp_dummy_magic_0.Y.t13 two_stage_opamp_dummy_magic_0.VD4.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X705 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 two_stage_opamp_dummy_magic_0.Y.t51 VDDA.t8 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X706 two_stage_opamp_dummy_magic_0.V_p_mir.t2 VIN-.t8 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X707 two_stage_opamp_dummy_magic_0.VD1.t18 VIN-.t9 two_stage_opamp_dummy_magic_0.V_source.t34 GNDA.t311 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X708 VOUT+.t142 two_stage_opamp_dummy_magic_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X709 VOUT-.t139 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X710 VDDA.t67 bgr_0.1st_Vout_2.t34 bgr_0.PFET_GATE_10uA.t0 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X711 VOUT-.t140 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X712 VOUT-.t141 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X713 GNDA.t66 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 VOUT+.t13 GNDA.t65 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X714 VOUT-.t142 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X715 VOUT-.t143 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X716 bgr_0.1st_Vout_1.t34 bgr_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X717 a_5190_5068.t1 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA.t341 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X718 bgr_0.1st_Vout_2.t35 bgr_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X719 VOUT+.t143 two_stage_opamp_dummy_magic_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X720 bgr_0.V_mir2.t1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 bgr_0.V_p_2.t4 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X721 two_stage_opamp_dummy_magic_0.VD1.t17 VIN-.t10 two_stage_opamp_dummy_magic_0.V_source.t33 GNDA.t310 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X722 two_stage_opamp_dummy_magic_0.X.t11 two_stage_opamp_dummy_magic_0.Vb2.t30 two_stage_opamp_dummy_magic_0.VD3.t3 two_stage_opamp_dummy_magic_0.VD3.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X723 VDDA.t275 two_stage_opamp_dummy_magic_0.Vb3.t27 two_stage_opamp_dummy_magic_0.VD4.t26 VDDA.t274 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X724 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 two_stage_opamp_dummy_magic_0.Y.t52 GNDA.t11 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X725 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 bgr_0.NFET_GATE_10uA.t23 GNDA.t176 GNDA.t175 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X726 VOUT+.t144 two_stage_opamp_dummy_magic_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X727 GNDA.t219 GNDA.t235 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X728 VOUT+.t145 two_stage_opamp_dummy_magic_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X729 two_stage_opamp_dummy_magic_0.V_err_gate.t10 VDDA.t321 VDDA.t323 VDDA.t322 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X730 VOUT-.t144 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X731 bgr_0.1st_Vout_1.t35 bgr_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X732 two_stage_opamp_dummy_magic_0.V_err_gate.t12 two_stage_opamp_dummy_magic_0.V_tot.t13 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 VDDA.t433 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X733 VOUT+.t146 two_stage_opamp_dummy_magic_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X734 VDDA.t253 bgr_0.1st_Vout_1.t36 bgr_0.V_TOP.t5 VDDA.t252 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X735 GNDA.t170 VDDA.t471 bgr_0.V_TOP.t9 GNDA.t167 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X736 two_stage_opamp_dummy_magic_0.Y.t15 two_stage_opamp_dummy_magic_0.Vb1.t25 two_stage_opamp_dummy_magic_0.VD2.t12 GNDA.t144 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X737 bgr_0.V_TOP.t47 VDDA.t210 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X738 two_stage_opamp_dummy_magic_0.Vb2.t1 two_stage_opamp_dummy_magic_0.Vb2.t0 VDDA.t116 VDDA.t115 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1 as=0.12 ps=1 w=0.6 l=0.2
X739 GNDA.t234 GNDA.t232 VOUT+.t15 GNDA.t233 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X740 VDDA.t235 two_stage_opamp_dummy_magic_0.X.t51 VOUT+.t2 VDDA.t234 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X741 VOUT+.t147 two_stage_opamp_dummy_magic_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X742 VDDA.t90 bgr_0.V_TOP.t48 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 VDDA.t89 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X743 VOUT-.t145 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X744 VOUT-.t146 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X745 VOUT-.t147 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X746 VOUT+.t148 two_stage_opamp_dummy_magic_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X747 VOUT+.t149 two_stage_opamp_dummy_magic_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X748 bgr_0.V_mir2.t0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 bgr_0.V_p_2.t3 GNDA.t338 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X749 VOUT-.t148 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X750 VDDA.t153 bgr_0.PFET_GATE_10uA.t29 bgr_0.V_CUR_REF_REG.t1 VDDA.t152 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X751 VDDA.t172 two_stage_opamp_dummy_magic_0.V_err_gate.t32 two_stage_opamp_dummy_magic_0.V_err_p.t9 VDDA.t171 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X752 two_stage_opamp_dummy_magic_0.Y.t8 two_stage_opamp_dummy_magic_0.VD4.t0 two_stage_opamp_dummy_magic_0.VD4.t2 two_stage_opamp_dummy_magic_0.VD4.t1 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X753 VOUT-.t149 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X754 VOUT+.t150 two_stage_opamp_dummy_magic_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X755 VOUT-.t150 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X756 two_stage_opamp_dummy_magic_0.X.t12 two_stage_opamp_dummy_magic_0.Vb2.t31 two_stage_opamp_dummy_magic_0.VD3.t1 two_stage_opamp_dummy_magic_0.VD3.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X757 VOUT+.t151 two_stage_opamp_dummy_magic_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X758 VOUT-.t18 a_5710_2076.t1 GNDA.t340 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X759 VDDA.t20 two_stage_opamp_dummy_magic_0.Y.t53 VOUT-.t2 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X760 VOUT-.t151 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X761 VOUT+.t152 two_stage_opamp_dummy_magic_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X762 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 two_stage_opamp_dummy_magic_0.X.t52 VDDA.t243 GNDA.t152 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X763 VOUT+.t153 two_stage_opamp_dummy_magic_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X764 bgr_0.V_p_1.t10 VDDA.t472 GNDA.t171 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X765 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 two_stage_opamp_dummy_magic_0.V_err_gate.t33 VDDA.t63 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X766 VOUT-.t152 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X767 bgr_0.V_TOP.t49 VDDA.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X768 two_stage_opamp_dummy_magic_0.X.t18 GNDA.t227 GNDA.t229 GNDA.t228 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X769 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 VDDA.t318 VDDA.t320 VDDA.t319 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X770 two_stage_opamp_dummy_magic_0.V_err_p.t5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 two_stage_opamp_dummy_magic_0.err_amp_out.t0 VDDA.t455 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X771 GNDA.t16 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 two_stage_opamp_dummy_magic_0.err_amp_out.t5 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X772 VOUT-.t153 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X773 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 two_stage_opamp_dummy_magic_0.X.t53 GNDA.t114 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X774 VOUT-.t154 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X775 VOUT+.t154 two_stage_opamp_dummy_magic_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X776 VOUT+.t155 two_stage_opamp_dummy_magic_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X777 bgr_0.1st_Vout_2.t36 bgr_0.cap_res2.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X778 a_5310_5068.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 GNDA.t351 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X779 VDDA.t443 bgr_0.V_mir1.t2 bgr_0.V_mir1.t3 VDDA.t442 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X780 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 two_stage_opamp_dummy_magic_0.X.t54 GNDA.t124 VDDA.t206 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X781 VOUT-.t155 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X782 GNDA.t226 GNDA.t224 two_stage_opamp_dummy_magic_0.V_source.t31 GNDA.t225 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X783 two_stage_opamp_dummy_magic_0.VD2.t15 GNDA.t221 GNDA.t223 GNDA.t222 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X784 VOUT-.t156 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X785 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 two_stage_opamp_dummy_magic_0.Y.t54 VDDA.t215 GNDA.t130 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X786 GNDA.t217 GNDA.t215 VDDA.t314 GNDA.t216 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X787 two_stage_opamp_dummy_magic_0.VD2.t8 VIN+.t10 two_stage_opamp_dummy_magic_0.V_source.t22 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X788 a_14680_5068.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 GNDA.t143 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X789 VDDA.t273 two_stage_opamp_dummy_magic_0.Vb3.t28 two_stage_opamp_dummy_magic_0.VD3.t20 VDDA.t272 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X790 VOUT+.t156 two_stage_opamp_dummy_magic_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.t1 384.967
R1 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t10 369.534
R2 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t22 369.534
R3 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t7 369.534
R4 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t16 369.534
R5 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t12 369.534
R6 bgr_0.NFET_GATE_10uA.t1 bgr_0.NFET_GATE_10uA.n18 369.534
R7 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n20 366.553
R8 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.t9 192.8
R9 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.t17 192.8
R10 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t23 192.8
R11 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t11 192.8
R12 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t20 192.8
R13 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t21 192.8
R14 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.t8 192.8
R15 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.t15 192.8
R16 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.t19 192.8
R17 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.t5 192.8
R18 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t13 192.8
R19 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.t18 192.8
R20 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.t6 192.8
R21 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.t14 192.8
R22 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.n11 176.733
R23 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.n10 176.733
R24 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.n4 176.733
R25 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.n5 176.733
R26 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.n2 176.733
R27 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.n1 176.733
R28 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.n17 176.733
R29 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.n16 176.733
R30 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n13 169.852
R31 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n8 169.852
R32 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n14 166.133
R33 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.n0 126.877
R34 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n12 56.2338
R35 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n9 56.2338
R36 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n7 56.2338
R37 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n6 56.2338
R38 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n3 56.2338
R39 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.n15 56.2338
R40 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t3 39.4005
R41 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t4 39.4005
R42 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n19 30.6442
R43 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t0 24.0005
R44 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t2 24.0005
R45 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.t22 661.375
R46 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.t12 611.739
R47 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.t25 611.739
R48 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.t11 611.739
R49 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.t20 611.739
R50 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.t18 421.75
R51 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.t21 421.75
R52 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.t24 421.75
R53 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.t27 421.75
R54 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.t23 421.75
R55 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.t19 421.75
R56 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.t14 421.75
R57 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.t9 421.75
R58 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.t17 421.75
R59 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.t15 421.75
R60 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.t26 421.75
R61 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.t28 421.75
R62 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.t16 421.75
R63 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.t10 421.75
R64 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.t13 421.75
R65 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.t8 421.75
R66 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.n23 176.25
R67 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.n14 175.696
R68 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.n5 174.964
R69 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.n19 167.094
R70 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.n20 167.094
R71 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.n21 167.094
R72 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.n15 167.094
R73 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.n16 167.094
R74 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.n17 167.094
R75 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.n10 167.094
R76 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.n11 167.094
R77 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.n12 167.094
R78 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.n6 167.094
R79 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.n7 167.094
R80 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.n8 167.094
R81 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.n0 139.639
R82 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.n1 139.638
R83 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.n3 134.577
R84 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.n22 47.1294
R85 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.n18 47.1294
R86 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.n13 47.1294
R87 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.n9 47.1294
R88 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb3.n4 41.063
R89 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb3.n26 37.1567
R90 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.t4 24.0005
R91 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.t6 24.0005
R92 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.t7 24.0005
R93 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.t0 24.0005
R94 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t5 24.0005
R95 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t3 24.0005
R96 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t2 10.9449
R97 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t1 10.9449
R98 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.n24 9.5005
R99 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.n25 6.28175
R100 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.n2 4.5005
R101 GNDA.n2066 GNDA.n29 227083
R102 GNDA.n2408 GNDA.n159 176550
R103 GNDA.n2408 GNDA.n160 127050
R104 GNDA.n2154 GNDA.n2153 39792.7
R105 GNDA.n2156 GNDA.n2155 32716.6
R106 GNDA.n2426 GNDA.n2425 30529.2
R107 GNDA.n2148 GNDA.n2068 29344.6
R108 GNDA.n2149 GNDA.n2148 28430.8
R109 GNDA.n2425 GNDA.n79 28430.8
R110 GNDA.n2067 GNDA.n2066 26656.2
R111 GNDA.n2153 GNDA.n2058 26648.4
R112 GNDA.n2149 GNDA.n2065 23523.1
R113 GNDA.n2065 GNDA.n79 23523.1
R114 GNDA.n2065 GNDA.n2064 19630.8
R115 GNDA.n2150 GNDA.n2149 18164.1
R116 GNDA.n2062 GNDA.n79 18118.3
R117 GNDA.n2155 GNDA.n2152 15840.2
R118 GNDA.n2156 GNDA.n2059 15312.1
R119 GNDA.n2155 GNDA.n2154 15051.6
R120 GNDA.n2152 GNDA.n2151 14764.7
R121 GNDA.n2059 GNDA.n2058 14331.7
R122 GNDA.n2157 GNDA.n2156 14285.8
R123 GNDA.n2183 GNDA.n176 12361.8
R124 GNDA.n2387 GNDA.n176 12312.5
R125 GNDA.n2066 GNDA.n79 11934.7
R126 GNDA.n2183 GNDA.n175 11918.5
R127 GNDA.n2387 GNDA.n175 11869.2
R128 GNDA.n2063 GNDA.n2062 11314.3
R129 GNDA.n2151 GNDA.n2150 11314.3
R130 GNDA.n2063 GNDA.n2061 10529
R131 GNDA.n40 GNDA.n39 10441
R132 GNDA.n41 GNDA.n39 10441
R133 GNDA.n2438 GNDA.n40 10441
R134 GNDA.n2438 GNDA.n41 10441
R135 GNDA.n2153 GNDA.t219 10371.4
R136 GNDA.n2061 GNDA.n159 9741.28
R137 GNDA.n2452 GNDA.n30 9259
R138 GNDA.n2369 GNDA.n2368 9062
R139 GNDA.n2452 GNDA.n31 8914.25
R140 GNDA.n2150 GNDA.n2060 8145.95
R141 GNDA.n2160 GNDA.n2058 7953.85
R142 GNDA.n186 GNDA.n184 7880
R143 GNDA.n2377 GNDA.n184 7880
R144 GNDA.n2186 GNDA.n307 7880
R145 GNDA.n2190 GNDA.n307 7880
R146 GNDA.n2374 GNDA.n186 7830.75
R147 GNDA.n2377 GNDA.n2374 7830.75
R148 GNDA.n2190 GNDA.n308 7830.75
R149 GNDA.n2186 GNDA.n308 7830.75
R150 GNDA.n144 GNDA.n132 7732.25
R151 GNDA.n144 GNDA.n100 7732.25
R152 GNDA.n146 GNDA.n132 7732.25
R153 GNDA.n146 GNDA.n100 7732.25
R154 GNDA.n2132 GNDA.n2105 7732.25
R155 GNDA.n2132 GNDA.n2106 7732.25
R156 GNDA.n2118 GNDA.n2105 7732.25
R157 GNDA.n2118 GNDA.n2106 7732.25
R158 GNDA.n2062 GNDA.n160 7472.73
R159 GNDA.n2390 GNDA.n170 7289
R160 GNDA.n2181 GNDA.n312 7289
R161 GNDA.n2394 GNDA.n170 7239.75
R162 GNDA.n2177 GNDA.n312 7239.75
R163 GNDA.n2151 GNDA.n2064 7071.43
R164 GNDA.n2390 GNDA.n169 6845.75
R165 GNDA.n2181 GNDA.n311 6845.75
R166 GNDA.n2394 GNDA.n169 6796.5
R167 GNDA.n2177 GNDA.n311 6796.5
R168 GNDA.n2398 GNDA.n167 6254.75
R169 GNDA.n2399 GNDA.n2398 6205.5
R170 GNDA.n167 GNDA.n166 6107
R171 GNDA.n2173 GNDA.n2051 6107
R172 GNDA.n2399 GNDA.n166 6057.75
R173 GNDA.n2052 GNDA.n2051 6057.75
R174 GNDA.n2173 GNDA.n2172 6057.75
R175 GNDA.n2172 GNDA.n2052 6008.5
R176 GNDA.n2140 GNDA.n2074 6008.5
R177 GNDA.n2416 GNDA.n88 5860.75
R178 GNDA.n2416 GNDA.n89 5811.5
R179 GNDA.n2092 GNDA.n2074 5762.25
R180 GNDA.n2068 GNDA.n2067 5446.53
R181 GNDA.n2427 GNDA.n76 5319
R182 GNDA.n2126 GNDA.n2120 5319
R183 GNDA.n2140 GNDA.n2075 5319
R184 GNDA.n2418 GNDA.n88 5319
R185 GNDA.n2092 GNDA.n2075 5269.75
R186 GNDA.n2418 GNDA.n89 5269.75
R187 GNDA.n2445 GNDA.n30 5171.25
R188 GNDA.n2447 GNDA.n31 5171.25
R189 GNDA.n2147 GNDA.n2070 5171.25
R190 GNDA.n150 GNDA.n94 5171.25
R191 GNDA.n2143 GNDA.n2070 5122
R192 GNDA.n154 GNDA.n94 5122
R193 GNDA.n2372 GNDA.n2368 4974.25
R194 GNDA.n1910 GNDA.n444 4974.25
R195 GNDA.n1909 GNDA.n444 4974.25
R196 GNDA.n2147 GNDA.n2071 4944.7
R197 GNDA.n150 GNDA.n96 4944.7
R198 GNDA.n61 GNDA.n37 4925
R199 GNDA.n68 GNDA.n37 4925
R200 GNDA.n2143 GNDA.n2071 4895.45
R201 GNDA.n154 GNDA.n96 4895.45
R202 GNDA.n61 GNDA.n38 4728
R203 GNDA.n68 GNDA.n38 4728
R204 GNDA.n1801 GNDA.n513 4678.75
R205 GNDA.n1790 GNDA.n513 4629.5
R206 GNDA.n1801 GNDA.n514 4629.5
R207 GNDA.n1790 GNDA.n514 4580.25
R208 GNDA.n2402 GNDA.n163 4580.25
R209 GNDA.n2406 GNDA.n163 4580.25
R210 GNDA.n2162 GNDA.n2056 4580.25
R211 GNDA.n2168 GNDA.n2056 4580.25
R212 GNDA.n1797 GNDA.n522 4531
R213 GNDA.n1797 GNDA.n1796 4531
R214 GNDA.n523 GNDA.n522 4531
R215 GNDA.n1796 GNDA.n523 4531
R216 GNDA.n1915 GNDA.n1909 4531
R217 GNDA.n1915 GNDA.n1910 4531
R218 GNDA.n2402 GNDA.n162 4481.75
R219 GNDA.n2406 GNDA.n162 4481.75
R220 GNDA.n2162 GNDA.n2055 4481.75
R221 GNDA.n2168 GNDA.n2055 4481.75
R222 GNDA.n2064 GNDA.n2063 4242.86
R223 GNDA.n2149 GNDA.n2067 3964.58
R224 GNDA.n139 GNDA.n82 3619.88
R225 GNDA.n2110 GNDA.n2108 3619.88
R226 GNDA.n2445 GNDA.n35 3595.25
R227 GNDA.n2455 GNDA.n26 3447.5
R228 GNDA.n2408 GNDA.n2407 3410.1
R229 GNDA.n2441 GNDA.n26 3398.25
R230 GNDA.n2455 GNDA.n27 3349
R231 GNDA.n2441 GNDA.n27 3299.75
R232 GNDA.n2447 GNDA.n35 3250.5
R233 GNDA.n2409 GNDA.n2408 3002.94
R234 GNDA.n135 GNDA.n82 2437.88
R235 GNDA.n2108 GNDA.n2098 2437.88
R236 GNDA.n2089 GNDA.n2078 2326.02
R237 GNDA.n2081 GNDA.n2078 2326.02
R238 GNDA.n158 GNDA.n92 2326.02
R239 GNDA.n2411 GNDA.n158 2326.02
R240 GNDA.n2091 GNDA.n2060 2270.39
R241 GNDA.n646 GNDA.n530 2142.38
R242 GNDA.n1921 GNDA.n438 2142.38
R243 GNDA.n2159 GNDA.n2059 1965.33
R244 GNDA.n2158 GNDA.n2157 1906.86
R245 GNDA.n1793 GNDA.n530 1846.88
R246 GNDA.n511 GNDA.n438 1846.88
R247 GNDA.n2154 GNDA.n159 1791
R248 GNDA.n2061 GNDA.n160 1600
R249 GNDA.n2423 GNDA.n82 1456.78
R250 GNDA.n2108 GNDA.n2097 1456.78
R251 GNDA.n2161 GNDA.n2160 1445.81
R252 GNDA.n2159 GNDA.n2158 1238.02
R253 GNDA.n2309 GNDA.n2308 1214.72
R254 GNDA.n2308 GNDA.n2307 1214.72
R255 GNDA.n2307 GNDA.n248 1214.72
R256 GNDA.n2301 GNDA.n248 1214.72
R257 GNDA.n2301 GNDA.n2300 1214.72
R258 GNDA.n2297 GNDA.n256 1214.72
R259 GNDA.n262 GNDA.n256 1214.72
R260 GNDA.n2290 GNDA.n262 1214.72
R261 GNDA.n2290 GNDA.n2289 1214.72
R262 GNDA.n2289 GNDA.n2288 1214.72
R263 GNDA.n1968 GNDA.n398 1214.72
R264 GNDA.n1974 GNDA.n398 1214.72
R265 GNDA.n1975 GNDA.n1974 1214.72
R266 GNDA.n1975 GNDA.n394 1214.72
R267 GNDA.n1981 GNDA.n394 1214.72
R268 GNDA.n1983 GNDA.n389 1214.72
R269 GNDA.n1989 GNDA.n389 1214.72
R270 GNDA.n1990 GNDA.n1989 1214.72
R271 GNDA.n1990 GNDA.n385 1214.72
R272 GNDA.n1996 GNDA.n385 1214.72
R273 GNDA.n2127 GNDA.n2068 1184.62
R274 GNDA.n2085 GNDA.n2078 1114.8
R275 GNDA.n158 GNDA.n157 1114.8
R276 GNDA.n2160 GNDA.n2159 1017.76
R277 GNDA.n530 GNDA.n529 991.841
R278 GNDA.n1918 GNDA.n438 991.841
R279 GNDA.n2152 GNDA.n2061 924.639
R280 GNDA.n2300 GNDA.t219 823.313
R281 GNDA.n1981 GNDA.t219 823.313
R282 GNDA.n2385 GNDA.n178 803.201
R283 GNDA.n2386 GNDA.n2385 800
R284 GNDA.n178 GNDA.n177 774.4
R285 GNDA.n2386 GNDA.n177 771.201
R286 GNDA.n2099 GNDA.t244 734.418
R287 GNDA.n2095 GNDA.t236 734.418
R288 GNDA.n84 GNDA.t239 734.418
R289 GNDA.n136 GNDA.t215 734.418
R290 GNDA.n2429 GNDA.n2428 691.201
R291 GNDA.n2125 GNDA.n72 691.201
R292 GNDA.n33 GNDA.t260 682.201
R293 GNDA.n2437 GNDA.n2436 678.4
R294 GNDA.n2437 GNDA.n42 672
R295 GNDA.n2041 GNDA.n335 669.307
R296 GNDA.n102 GNDA.t224 666.134
R297 GNDA.n2088 GNDA.n2082 617.601
R298 GNDA.n2412 GNDA.n91 617.601
R299 GNDA.n2451 GNDA.n32 601.601
R300 GNDA.n541 GNDA.n539 598.37
R301 GNDA.n506 GNDA.n505 596.981
R302 GNDA.t298 GNDA.n2127 592.308
R303 GNDA.n2426 GNDA.t295 592.308
R304 GNDA.n1646 GNDA.n1645 585
R305 GNDA.n1648 GNDA.n1647 585
R306 GNDA.n1650 GNDA.n1649 585
R307 GNDA.n1652 GNDA.n1651 585
R308 GNDA.n1654 GNDA.n1653 585
R309 GNDA.n1656 GNDA.n1655 585
R310 GNDA.n1658 GNDA.n1657 585
R311 GNDA.n1660 GNDA.n1659 585
R312 GNDA.n1662 GNDA.n1661 585
R313 GNDA.n1664 GNDA.n1663 585
R314 GNDA.n1665 GNDA.n429 585
R315 GNDA.n1923 GNDA.n429 585
R316 GNDA.n1667 GNDA.n1666 585
R317 GNDA.n1668 GNDA.n1667 585
R318 GNDA.n1927 GNDA.n415 585
R319 GNDA.n1926 GNDA.n1925 585
R320 GNDA.n417 GNDA.n416 585
R321 GNDA.n784 GNDA.n783 585
R322 GNDA.n786 GNDA.n785 585
R323 GNDA.n788 GNDA.n787 585
R324 GNDA.n790 GNDA.n789 585
R325 GNDA.n792 GNDA.n791 585
R326 GNDA.n794 GNDA.n793 585
R327 GNDA.n796 GNDA.n795 585
R328 GNDA.n797 GNDA.n422 585
R329 GNDA.n1923 GNDA.n422 585
R330 GNDA.n799 GNDA.n798 585
R331 GNDA.n799 GNDA.n782 585
R332 GNDA.n1923 GNDA.n437 585
R333 GNDA.n481 GNDA.n480 585
R334 GNDA.n483 GNDA.n482 585
R335 GNDA.n485 GNDA.n484 585
R336 GNDA.n487 GNDA.n486 585
R337 GNDA.n489 GNDA.n488 585
R338 GNDA.n491 GNDA.n490 585
R339 GNDA.n493 GNDA.n492 585
R340 GNDA.n495 GNDA.n494 585
R341 GNDA.n497 GNDA.n496 585
R342 GNDA.n499 GNDA.n498 585
R343 GNDA.n501 GNDA.n500 585
R344 GNDA.n2287 GNDA.n2286 585
R345 GNDA.n2288 GNDA.n2287 585
R346 GNDA.n263 GNDA.n260 585
R347 GNDA.n2289 GNDA.n263 585
R348 GNDA.n2292 GNDA.n259 585
R349 GNDA.n2290 GNDA.n259 585
R350 GNDA.n2293 GNDA.n258 585
R351 GNDA.n262 GNDA.n258 585
R352 GNDA.n2294 GNDA.n254 585
R353 GNDA.n256 GNDA.n254 585
R354 GNDA.n2298 GNDA.n255 585
R355 GNDA.n2298 GNDA.n2297 585
R356 GNDA.n2299 GNDA.n252 585
R357 GNDA.n2300 GNDA.n2299 585
R358 GNDA.n2303 GNDA.n251 585
R359 GNDA.n2301 GNDA.n251 585
R360 GNDA.n2304 GNDA.n250 585
R361 GNDA.n250 GNDA.n248 585
R362 GNDA.n2305 GNDA.n247 585
R363 GNDA.n2307 GNDA.n247 585
R364 GNDA.n246 GNDA.n243 585
R365 GNDA.n2308 GNDA.n246 585
R366 GNDA.n2311 GNDA.n224 585
R367 GNDA.n2309 GNDA.n224 585
R368 GNDA.n2311 GNDA.n2310 585
R369 GNDA.n2310 GNDA.n2309 585
R370 GNDA.n245 GNDA.n243 585
R371 GNDA.n2308 GNDA.n245 585
R372 GNDA.n2306 GNDA.n2305 585
R373 GNDA.n2307 GNDA.n2306 585
R374 GNDA.n2304 GNDA.n249 585
R375 GNDA.n249 GNDA.n248 585
R376 GNDA.n2303 GNDA.n2302 585
R377 GNDA.n2302 GNDA.n2301 585
R378 GNDA.n253 GNDA.n252 585
R379 GNDA.n2300 GNDA.n253 585
R380 GNDA.n2296 GNDA.n255 585
R381 GNDA.n2297 GNDA.n2296 585
R382 GNDA.n2295 GNDA.n2294 585
R383 GNDA.n2295 GNDA.n256 585
R384 GNDA.n2293 GNDA.n257 585
R385 GNDA.n262 GNDA.n257 585
R386 GNDA.n2292 GNDA.n2291 585
R387 GNDA.n2291 GNDA.n2290 585
R388 GNDA.n261 GNDA.n260 585
R389 GNDA.n2289 GNDA.n261 585
R390 GNDA.n2286 GNDA.n264 585
R391 GNDA.n2288 GNDA.n264 585
R392 GNDA.n1714 GNDA.n1200 585
R393 GNDA.n1716 GNDA.n1191 585
R394 GNDA.n1717 GNDA.n1190 585
R395 GNDA.n1720 GNDA.n1189 585
R396 GNDA.n1721 GNDA.n1188 585
R397 GNDA.n1724 GNDA.n1187 585
R398 GNDA.n1725 GNDA.n1186 585
R399 GNDA.n1728 GNDA.n1185 585
R400 GNDA.n1729 GNDA.n1184 585
R401 GNDA.n1730 GNDA.n1183 585
R402 GNDA.n1192 GNDA.n1174 585
R403 GNDA.n1735 GNDA.n1171 585
R404 GNDA.n1735 GNDA.n1734 585
R405 GNDA.n1176 GNDA.n1174 585
R406 GNDA.n1731 GNDA.n1730 585
R407 GNDA.n1732 GNDA.n1731 585
R408 GNDA.n1729 GNDA.n1182 585
R409 GNDA.n1728 GNDA.n1727 585
R410 GNDA.n1726 GNDA.n1725 585
R411 GNDA.n1724 GNDA.n1723 585
R412 GNDA.n1722 GNDA.n1721 585
R413 GNDA.n1720 GNDA.n1719 585
R414 GNDA.n1718 GNDA.n1717 585
R415 GNDA.n1716 GNDA.n1715 585
R416 GNDA.n1714 GNDA.n1181 585
R417 GNDA.n1732 GNDA.n1181 585
R418 GNDA.n1995 GNDA.n384 585
R419 GNDA.n1996 GNDA.n1995 585
R420 GNDA.n1994 GNDA.n1993 585
R421 GNDA.n1994 GNDA.n385 585
R422 GNDA.n1992 GNDA.n386 585
R423 GNDA.n1990 GNDA.n386 585
R424 GNDA.n1988 GNDA.n387 585
R425 GNDA.n1989 GNDA.n1988 585
R426 GNDA.n1987 GNDA.n1986 585
R427 GNDA.n1987 GNDA.n389 585
R428 GNDA.n391 GNDA.n390 585
R429 GNDA.n1983 GNDA.n390 585
R430 GNDA.n1980 GNDA.n393 585
R431 GNDA.n1981 GNDA.n1980 585
R432 GNDA.n1979 GNDA.n1978 585
R433 GNDA.n1979 GNDA.n394 585
R434 GNDA.n1977 GNDA.n395 585
R435 GNDA.n1975 GNDA.n395 585
R436 GNDA.n1973 GNDA.n396 585
R437 GNDA.n1974 GNDA.n1973 585
R438 GNDA.n1972 GNDA.n1971 585
R439 GNDA.n1972 GNDA.n398 585
R440 GNDA.n400 GNDA.n399 585
R441 GNDA.n1968 GNDA.n399 585
R442 GNDA.n1969 GNDA.n400 585
R443 GNDA.n1969 GNDA.n1968 585
R444 GNDA.n1971 GNDA.n1970 585
R445 GNDA.n1970 GNDA.n398 585
R446 GNDA.n397 GNDA.n396 585
R447 GNDA.n1974 GNDA.n397 585
R448 GNDA.n1977 GNDA.n1976 585
R449 GNDA.n1976 GNDA.n1975 585
R450 GNDA.n1978 GNDA.n392 585
R451 GNDA.n394 GNDA.n392 585
R452 GNDA.n1982 GNDA.n393 585
R453 GNDA.n1982 GNDA.n1981 585
R454 GNDA.n1984 GNDA.n391 585
R455 GNDA.n1984 GNDA.n1983 585
R456 GNDA.n1986 GNDA.n1985 585
R457 GNDA.n1985 GNDA.n389 585
R458 GNDA.n388 GNDA.n387 585
R459 GNDA.n1989 GNDA.n388 585
R460 GNDA.n1992 GNDA.n1991 585
R461 GNDA.n1991 GNDA.n1990 585
R462 GNDA.n1993 GNDA.n383 585
R463 GNDA.n385 GNDA.n383 585
R464 GNDA.n1997 GNDA.n384 585
R465 GNDA.n1997 GNDA.n1996 585
R466 GNDA.n1952 GNDA.n1951 585
R467 GNDA.n1951 GNDA.n402 585
R468 GNDA.n1950 GNDA.n405 585
R469 GNDA.n1950 GNDA.n1949 585
R470 GNDA.n1944 GNDA.n406 585
R471 GNDA.n1948 GNDA.n406 585
R472 GNDA.n1946 GNDA.n1945 585
R473 GNDA.n1947 GNDA.n1946 585
R474 GNDA.n1943 GNDA.n408 585
R475 GNDA.n408 GNDA.n407 585
R476 GNDA.n1942 GNDA.n1941 585
R477 GNDA.n1941 GNDA.n1940 585
R478 GNDA.n410 GNDA.n409 585
R479 GNDA.n1939 GNDA.n410 585
R480 GNDA.n1937 GNDA.n1936 585
R481 GNDA.n1938 GNDA.n1937 585
R482 GNDA.n1935 GNDA.n412 585
R483 GNDA.n412 GNDA.n411 585
R484 GNDA.n1934 GNDA.n1933 585
R485 GNDA.n1933 GNDA.n1932 585
R486 GNDA.n414 GNDA.n413 585
R487 GNDA.n1931 GNDA.n414 585
R488 GNDA.n1929 GNDA.n1928 585
R489 GNDA.n1930 GNDA.n1929 585
R490 GNDA.n2040 GNDA.n2039 585
R491 GNDA.n2038 GNDA.n336 585
R492 GNDA.n2038 GNDA.t219 585
R493 GNDA.n1738 GNDA.n1737 585
R494 GNDA.n1172 GNDA.n1170 585
R495 GNDA.n1626 GNDA.n1625 585
R496 GNDA.n1628 GNDA.n1627 585
R497 GNDA.n1630 GNDA.n1629 585
R498 GNDA.n1632 GNDA.n1631 585
R499 GNDA.n1634 GNDA.n1633 585
R500 GNDA.n1636 GNDA.n1635 585
R501 GNDA.n1638 GNDA.n1637 585
R502 GNDA.n1640 GNDA.n1639 585
R503 GNDA.n1642 GNDA.n1641 585
R504 GNDA.n1644 GNDA.n1643 585
R505 GNDA.n1485 GNDA.n1484 585
R506 GNDA.n1483 GNDA.n1482 585
R507 GNDA.n1481 GNDA.n1480 585
R508 GNDA.n1479 GNDA.n1478 585
R509 GNDA.n1477 GNDA.n1476 585
R510 GNDA.n1475 GNDA.n1474 585
R511 GNDA.n1473 GNDA.n1472 585
R512 GNDA.n1471 GNDA.n1470 585
R513 GNDA.n1469 GNDA.n1468 585
R514 GNDA.n1467 GNDA.n1466 585
R515 GNDA.n1465 GNDA.n1464 585
R516 GNDA.n1175 GNDA.n1173 585
R517 GNDA.n1742 GNDA.n1152 585
R518 GNDA.n1487 GNDA.n1153 585
R519 GNDA.n1489 GNDA.n1488 585
R520 GNDA.n1491 GNDA.n1490 585
R521 GNDA.n1493 GNDA.n1492 585
R522 GNDA.n1495 GNDA.n1494 585
R523 GNDA.n1497 GNDA.n1496 585
R524 GNDA.n1499 GNDA.n1498 585
R525 GNDA.n1501 GNDA.n1500 585
R526 GNDA.n1503 GNDA.n1502 585
R527 GNDA.n1505 GNDA.n1504 585
R528 GNDA.n1507 GNDA.n1506 585
R529 GNDA.n381 GNDA.n380 585
R530 GNDA.n1999 GNDA.n380 585
R531 GNDA.n1030 GNDA.n1029 585
R532 GNDA.n1027 GNDA.n781 585
R533 GNDA.n802 GNDA.n801 585
R534 GNDA.n1022 GNDA.n1021 585
R535 GNDA.n1020 GNDA.n1019 585
R536 GNDA.n946 GNDA.n806 585
R537 GNDA.n948 GNDA.n947 585
R538 GNDA.n953 GNDA.n952 585
R539 GNDA.n951 GNDA.n944 585
R540 GNDA.n959 GNDA.n958 585
R541 GNDA.n961 GNDA.n960 585
R542 GNDA.n942 GNDA.n941 585
R543 GNDA.n1998 GNDA.n381 585
R544 GNDA.n1999 GNDA.n1998 585
R545 GNDA.n939 GNDA.n382 585
R546 GNDA.n937 GNDA.n936 585
R547 GNDA.n935 GNDA.n934 585
R548 GNDA.n851 GNDA.n827 585
R549 GNDA.n853 GNDA.n852 585
R550 GNDA.n857 GNDA.n856 585
R551 GNDA.n859 GNDA.n858 585
R552 GNDA.n866 GNDA.n865 585
R553 GNDA.n864 GNDA.n849 585
R554 GNDA.n872 GNDA.n871 585
R555 GNDA.n874 GNDA.n873 585
R556 GNDA.n847 GNDA.n846 585
R557 GNDA.n2314 GNDA.n2313 585
R558 GNDA.n225 GNDA.n223 585
R559 GNDA.n461 GNDA.n460 585
R560 GNDA.n463 GNDA.n462 585
R561 GNDA.n465 GNDA.n464 585
R562 GNDA.n467 GNDA.n466 585
R563 GNDA.n469 GNDA.n468 585
R564 GNDA.n471 GNDA.n470 585
R565 GNDA.n473 GNDA.n472 585
R566 GNDA.n475 GNDA.n474 585
R567 GNDA.n477 GNDA.n476 585
R568 GNDA.n479 GNDA.n478 585
R569 GNDA.n2322 GNDA.n2321 585
R570 GNDA.n2320 GNDA.n2319 585
R571 GNDA.n2318 GNDA.n206 585
R572 GNDA.n226 GNDA.n207 585
R573 GNDA.n228 GNDA.n227 585
R574 GNDA.n230 GNDA.n229 585
R575 GNDA.n232 GNDA.n231 585
R576 GNDA.n234 GNDA.n233 585
R577 GNDA.n236 GNDA.n235 585
R578 GNDA.n238 GNDA.n237 585
R579 GNDA.n240 GNDA.n239 585
R580 GNDA.n244 GNDA.n241 585
R581 GNDA.n1132 GNDA.n1131 585
R582 GNDA.n1130 GNDA.n1129 585
R583 GNDA.n1128 GNDA.n1127 585
R584 GNDA.n1126 GNDA.n1125 585
R585 GNDA.n1124 GNDA.n1123 585
R586 GNDA.n1122 GNDA.n1121 585
R587 GNDA.n1120 GNDA.n1119 585
R588 GNDA.n1118 GNDA.n1117 585
R589 GNDA.n1116 GNDA.n1115 585
R590 GNDA.n1114 GNDA.n1113 585
R591 GNDA.n1112 GNDA.n1111 585
R592 GNDA.n1110 GNDA.n203 585
R593 GNDA.n1203 GNDA.n242 585
R594 GNDA.n1543 GNDA.n1203 585
R595 GNDA.n1671 GNDA.n1670 585
R596 GNDA.n1672 GNDA.n1559 585
R597 GNDA.n1682 GNDA.n1681 585
R598 GNDA.n1684 GNDA.n1558 585
R599 GNDA.n1687 GNDA.n1686 585
R600 GNDA.n1688 GNDA.n1554 585
R601 GNDA.n1697 GNDA.n1696 585
R602 GNDA.n1699 GNDA.n1553 585
R603 GNDA.n1702 GNDA.n1701 585
R604 GNDA.n1549 GNDA.n1548 585
R605 GNDA.n1709 GNDA.n1708 585
R606 GNDA.n1712 GNDA.n1711 585
R607 GNDA.n1544 GNDA.n242 585
R608 GNDA.n1544 GNDA.n1543 585
R609 GNDA.n1545 GNDA.n1201 585
R610 GNDA.n1409 GNDA.n1216 585
R611 GNDA.n1432 GNDA.n1431 585
R612 GNDA.n1429 GNDA.n1428 585
R613 GNDA.n1427 GNDA.n1426 585
R614 GNDA.n1422 GNDA.n1421 585
R615 GNDA.n1420 GNDA.n1419 585
R616 GNDA.n1415 GNDA.n1414 585
R617 GNDA.n1413 GNDA.n1335 585
R618 GNDA.n1440 GNDA.n1439 585
R619 GNDA.n1442 GNDA.n1441 585
R620 GNDA.n1445 GNDA.n1444 585
R621 GNDA.n1332 GNDA.n1219 585
R622 GNDA.n1330 GNDA.n1329 585
R623 GNDA.n1328 GNDA.n1327 585
R624 GNDA.n1244 GNDA.n1222 585
R625 GNDA.n1246 GNDA.n1245 585
R626 GNDA.n1250 GNDA.n1249 585
R627 GNDA.n1252 GNDA.n1251 585
R628 GNDA.n1259 GNDA.n1258 585
R629 GNDA.n1257 GNDA.n1242 585
R630 GNDA.n1265 GNDA.n1264 585
R631 GNDA.n1267 GNDA.n1266 585
R632 GNDA.n1151 GNDA.n1150 585
R633 GNDA.n1771 GNDA.n1770 585
R634 GNDA.n642 GNDA.n641 585
R635 GNDA.n1135 GNDA.n1134 585
R636 GNDA.n1137 GNDA.n1136 585
R637 GNDA.n1139 GNDA.n1138 585
R638 GNDA.n1141 GNDA.n1140 585
R639 GNDA.n1143 GNDA.n1142 585
R640 GNDA.n1145 GNDA.n1144 585
R641 GNDA.n1146 GNDA.n1109 585
R642 GNDA.n1148 GNDA.n1147 585
R643 GNDA.n1133 GNDA.n1108 585
R644 GNDA.n1768 GNDA.n1103 585
R645 GNDA.n1764 GNDA.n1763 585
R646 GNDA.n1762 GNDA.n1761 585
R647 GNDA.n1760 GNDA.n1759 585
R648 GNDA.n1758 GNDA.n1757 585
R649 GNDA.n1756 GNDA.n1755 585
R650 GNDA.n1754 GNDA.n1753 585
R651 GNDA.n1752 GNDA.n1751 585
R652 GNDA.n1750 GNDA.n1749 585
R653 GNDA.n1748 GNDA.n1747 585
R654 GNDA.n1746 GNDA.n1745 585
R655 GNDA.n1744 GNDA.n1743 585
R656 GNDA.n1768 GNDA.n1767 585
R657 GNDA.n1768 GNDA.n1096 585
R658 GNDA.n663 GNDA.n376 585
R659 GNDA.n768 GNDA.n767 585
R660 GNDA.n665 GNDA.n662 585
R661 GNDA.n762 GNDA.n761 585
R662 GNDA.n760 GNDA.n759 585
R663 GNDA.n678 GNDA.n669 585
R664 GNDA.n680 GNDA.n679 585
R665 GNDA.n684 GNDA.n683 585
R666 GNDA.n686 GNDA.n685 585
R667 GNDA.n687 GNDA.n657 585
R668 GNDA.n1035 GNDA.n1034 585
R669 GNDA.n1037 GNDA.n654 585
R670 GNDA.n1093 GNDA.n1092 585
R671 GNDA.n1091 GNDA.n1090 585
R672 GNDA.n1089 GNDA.n1088 585
R673 GNDA.n1087 GNDA.n1086 585
R674 GNDA.n1085 GNDA.n1084 585
R675 GNDA.n1083 GNDA.n1082 585
R676 GNDA.n1081 GNDA.n1080 585
R677 GNDA.n1079 GNDA.n1078 585
R678 GNDA.n1077 GNDA.n1076 585
R679 GNDA.n1075 GNDA.n1074 585
R680 GNDA.n1073 GNDA.n1072 585
R681 GNDA.n1071 GNDA.n1038 585
R682 GNDA.n1071 GNDA.n1070 585
R683 GNDA.n1065 GNDA.n1039 585
R684 GNDA.n1069 GNDA.n1039 585
R685 GNDA.n1067 GNDA.n1066 585
R686 GNDA.n1068 GNDA.n1067 585
R687 GNDA.n1064 GNDA.n1041 585
R688 GNDA.n1041 GNDA.n1040 585
R689 GNDA.n1063 GNDA.n1062 585
R690 GNDA.n1062 GNDA.n1061 585
R691 GNDA.n1043 GNDA.n1042 585
R692 GNDA.n1060 GNDA.n1043 585
R693 GNDA.n1058 GNDA.n1057 585
R694 GNDA.n1059 GNDA.n1058 585
R695 GNDA.n1056 GNDA.n1045 585
R696 GNDA.n1045 GNDA.n1044 585
R697 GNDA.n1055 GNDA.n1054 585
R698 GNDA.n1054 GNDA.n1053 585
R699 GNDA.n1047 GNDA.n1046 585
R700 GNDA.n1052 GNDA.n1047 585
R701 GNDA.n1050 GNDA.n1049 585
R702 GNDA.n1051 GNDA.n1050 585
R703 GNDA.n349 GNDA.n346 585
R704 GNDA.n1048 GNDA.n349 585
R705 GNDA.n2026 GNDA.n345 585
R706 GNDA.n345 GNDA.n344 585
R707 GNDA.n2028 GNDA.n2027 585
R708 GNDA.n2029 GNDA.n2028 585
R709 GNDA.n343 GNDA.n342 585
R710 GNDA.n2030 GNDA.n343 585
R711 GNDA.n2033 GNDA.n2032 585
R712 GNDA.n2032 GNDA.n2031 585
R713 GNDA.n2034 GNDA.n340 585
R714 GNDA.n340 GNDA.n338 585
R715 GNDA.n2036 GNDA.n2035 585
R716 GNDA.n2037 GNDA.n2036 585
R717 GNDA.n1955 GNDA.n339 585
R718 GNDA.n339 GNDA.n337 585
R719 GNDA.n1957 GNDA.n1956 585
R720 GNDA.n1958 GNDA.n1957 585
R721 GNDA.n1961 GNDA.n1960 585
R722 GNDA.n1960 GNDA.n1959 585
R723 GNDA.n1962 GNDA.n404 585
R724 GNDA.n404 GNDA.n403 585
R725 GNDA.n1964 GNDA.n1963 585
R726 GNDA.n1965 GNDA.n1964 585
R727 GNDA.n1954 GNDA.n401 585
R728 GNDA.n1966 GNDA.n401 585
R729 GNDA.n2002 GNDA.n374 585
R730 GNDA.n2003 GNDA.n365 585
R731 GNDA.n2006 GNDA.n364 585
R732 GNDA.n2007 GNDA.n363 585
R733 GNDA.n2010 GNDA.n362 585
R734 GNDA.n2011 GNDA.n361 585
R735 GNDA.n2014 GNDA.n360 585
R736 GNDA.n2016 GNDA.n359 585
R737 GNDA.n2017 GNDA.n358 585
R738 GNDA.n2018 GNDA.n357 585
R739 GNDA.n366 GNDA.n348 585
R740 GNDA.n2024 GNDA.n347 585
R741 GNDA.n379 GNDA.n377 585
R742 GNDA.n1999 GNDA.n379 585
R743 GNDA.n2024 GNDA.n2023 585
R744 GNDA.n350 GNDA.n348 585
R745 GNDA.n2019 GNDA.n2018 585
R746 GNDA.n2017 GNDA.n356 585
R747 GNDA.n2016 GNDA.n2015 585
R748 GNDA.n2014 GNDA.n2013 585
R749 GNDA.n2012 GNDA.n2011 585
R750 GNDA.n2010 GNDA.n2009 585
R751 GNDA.n2008 GNDA.n2007 585
R752 GNDA.n2006 GNDA.n2005 585
R753 GNDA.n2004 GNDA.n2003 585
R754 GNDA.n2002 GNDA.n2001 585
R755 GNDA.n2000 GNDA.n377 585
R756 GNDA.n2000 GNDA.n1999 585
R757 GNDA.n1535 GNDA.n1447 585
R758 GNDA.n1538 GNDA.n1537 585
R759 GNDA.n1451 GNDA.n1450 585
R760 GNDA.n1531 GNDA.n1530 585
R761 GNDA.n1457 GNDA.n1456 585
R762 GNDA.n1524 GNDA.n1523 585
R763 GNDA.n1522 GNDA.n1521 585
R764 GNDA.n1520 GNDA.n1461 585
R765 GNDA.n1460 GNDA.n1459 585
R766 GNDA.n1514 GNDA.n1513 585
R767 GNDA.n1512 GNDA.n1511 585
R768 GNDA.n1510 GNDA.n1486 585
R769 GNDA.n1218 GNDA.n1217 585
R770 GNDA.n1543 GNDA.n1217 585
R771 GNDA.n1510 GNDA.n1509 585
R772 GNDA.n1511 GNDA.n1462 585
R773 GNDA.n1515 GNDA.n1514 585
R774 GNDA.n1517 GNDA.n1459 585
R775 GNDA.n1520 GNDA.n1519 585
R776 GNDA.n1521 GNDA.n1458 585
R777 GNDA.n1525 GNDA.n1524 585
R778 GNDA.n1527 GNDA.n1457 585
R779 GNDA.n1530 GNDA.n1529 585
R780 GNDA.n1450 GNDA.n1449 585
R781 GNDA.n1539 GNDA.n1538 585
R782 GNDA.n1541 GNDA.n1447 585
R783 GNDA.n1542 GNDA.n1218 585
R784 GNDA.n1543 GNDA.n1542 585
R785 GNDA.n196 GNDA.n190 585
R786 GNDA.n2341 GNDA.n2340 585
R787 GNDA.n2342 GNDA.n2332 585
R788 GNDA.n2345 GNDA.n2331 585
R789 GNDA.n2346 GNDA.n2330 585
R790 GNDA.n2349 GNDA.n2329 585
R791 GNDA.n2350 GNDA.n2328 585
R792 GNDA.n2353 GNDA.n2327 585
R793 GNDA.n2355 GNDA.n2326 585
R794 GNDA.n2356 GNDA.n2325 585
R795 GNDA.n2357 GNDA.n2324 585
R796 GNDA.n2358 GNDA.n2323 585
R797 GNDA.n2359 GNDA.n2358 585
R798 GNDA.n2357 GNDA.n202 585
R799 GNDA.n2356 GNDA.n201 585
R800 GNDA.n2361 GNDA.n201 585
R801 GNDA.n2355 GNDA.n2354 585
R802 GNDA.n2353 GNDA.n2352 585
R803 GNDA.n2351 GNDA.n2350 585
R804 GNDA.n2349 GNDA.n2348 585
R805 GNDA.n2347 GNDA.n2346 585
R806 GNDA.n2345 GNDA.n2344 585
R807 GNDA.n2343 GNDA.n2342 585
R808 GNDA.n2341 GNDA.n195 585
R809 GNDA.n2362 GNDA.n196 585
R810 GNDA.n2362 GNDA.n2361 585
R811 GNDA.n2284 GNDA.n266 585
R812 GNDA.n510 GNDA.n266 585
R813 GNDA.n505 GNDA.n504 585
R814 GNDA.n1884 GNDA.n1883 585
R815 GNDA.n1883 GNDA.n1882 585
R816 GNDA.n457 GNDA.n456 585
R817 GNDA.n1881 GNDA.n456 585
R818 GNDA.n1892 GNDA.n1891 585
R819 GNDA.n1893 GNDA.n1892 585
R820 GNDA.n455 GNDA.n454 585
R821 GNDA.n1894 GNDA.n455 585
R822 GNDA.n1897 GNDA.n1896 585
R823 GNDA.n1896 GNDA.n1895 585
R824 GNDA.n451 GNDA.n446 585
R825 GNDA.n446 GNDA.n445 585
R826 GNDA.n1907 GNDA.n1906 585
R827 GNDA.n1908 GNDA.n1907 585
R828 GNDA.n449 GNDA.n447 585
R829 GNDA.n507 GNDA.n447 585
R830 GNDA.n1806 GNDA.n509 585
R831 GNDA.n509 GNDA.n508 585
R832 GNDA.n1879 GNDA.n1878 585
R833 GNDA.n1880 GNDA.n1879 585
R834 GNDA.n1804 GNDA.n268 585
R835 GNDA.n1804 GNDA.n1803 585
R836 GNDA.n2365 GNDA.n2364 585
R837 GNDA.n2366 GNDA.n2365 585
R838 GNDA.n2284 GNDA.n2283 585
R839 GNDA.n2283 GNDA.n269 585
R840 GNDA.n2282 GNDA.n267 585
R841 GNDA.n2282 GNDA.n2281 585
R842 GNDA.n2269 GNDA.n270 585
R843 GNDA.n2280 GNDA.n270 585
R844 GNDA.n2278 GNDA.n2277 585
R845 GNDA.n2279 GNDA.n2278 585
R846 GNDA.n274 GNDA.n272 585
R847 GNDA.n305 GNDA.n272 585
R848 GNDA.n304 GNDA.n303 585
R849 GNDA.n306 GNDA.n304 585
R850 GNDA.n2193 GNDA.n299 585
R851 GNDA.n2193 GNDA.n2192 585
R852 GNDA.n2198 GNDA.n2197 585
R853 GNDA.n2197 GNDA.n2196 585
R854 GNDA.n2203 GNDA.n298 585
R855 GNDA.n2194 GNDA.n298 585
R856 GNDA.n2209 GNDA.n2208 585
R857 GNDA.n2210 GNDA.n2209 585
R858 GNDA.n297 GNDA.n296 585
R859 GNDA.n2211 GNDA.n297 585
R860 GNDA.n2215 GNDA.n2214 585
R861 GNDA.n2214 GNDA.n2213 585
R862 GNDA.n294 GNDA.n191 585
R863 GNDA.n2212 GNDA.n191 585
R864 GNDA.n2364 GNDA.n2363 585
R865 GNDA.n2363 GNDA.n193 585
R866 GNDA.n532 GNDA.n194 585
R867 GNDA.n1789 GNDA.n194 585
R868 GNDA.n1787 GNDA.n1786 585
R869 GNDA.n1788 GNDA.n1787 585
R870 GNDA.n534 GNDA.n531 585
R871 GNDA.n1778 GNDA.n531 585
R872 GNDA.n1781 GNDA.n1780 585
R873 GNDA.n1780 GNDA.n1779 585
R874 GNDA.n616 GNDA.n538 585
R875 GNDA.n538 GNDA.n187 585
R876 GNDA.n617 GNDA.n612 585
R877 GNDA.n612 GNDA.n611 585
R878 GNDA.n626 GNDA.n625 585
R879 GNDA.n627 GNDA.n626 585
R880 GNDA.n613 GNDA.n610 585
R881 GNDA.n628 GNDA.n610 585
R882 GNDA.n632 GNDA.n631 585
R883 GNDA.n631 GNDA.n630 585
R884 GNDA.n633 GNDA.n540 585
R885 GNDA.n629 GNDA.n540 585
R886 GNDA.n1776 GNDA.n1775 585
R887 GNDA.n1777 GNDA.n1776 585
R888 GNDA.n1773 GNDA.n541 585
R889 GNDA.n2136 GNDA.n2097 585
R890 GNDA.n2097 GNDA.n2069 585
R891 GNDA.n2423 GNDA.n2422 585
R892 GNDA.n2424 GNDA.n2423 585
R893 GNDA.n2135 GNDA.n2100 569.601
R894 GNDA.n137 GNDA.n83 569.601
R895 GNDA.n2101 GNDA.t232 535.191
R896 GNDA.n2103 GNDA.t303 535.191
R897 GNDA.n98 GNDA.t251 535.191
R898 GNDA.n140 GNDA.t257 535.191
R899 GNDA.n2288 GNDA.n265 512.884
R900 GNDA.n1996 GNDA.t219 512.884
R901 GNDA.n2379 GNDA.n2378 512
R902 GNDA.n2379 GNDA.n183 512
R903 GNDA.n2189 GNDA.n309 512
R904 GNDA.n2187 GNDA.n309 512
R905 GNDA.n2378 GNDA.n185 508.8
R906 GNDA.n185 GNDA.n183 508.8
R907 GNDA.n2189 GNDA.n2188 508.8
R908 GNDA.n2188 GNDA.n2187 508.8
R909 GNDA.n2117 GNDA.n2116 496
R910 GNDA.n147 GNDA.n101 496
R911 GNDA.n46 GNDA.t242 493.418
R912 GNDA.n47 GNDA.t221 493.418
R913 GNDA.n48 GNDA.t291 493.418
R914 GNDA.n43 GNDA.t306 493.418
R915 GNDA.n44 GNDA.t288 493.418
R916 GNDA.n45 GNDA.t282 493.418
R917 GNDA.n77 GNDA.t294 493.418
R918 GNDA.n73 GNDA.t285 493.418
R919 GNDA.n2122 GNDA.t227 493.418
R920 GNDA.n2121 GNDA.t297 493.418
R921 GNDA.n2117 GNDA.n2111 489.601
R922 GNDA.n148 GNDA.n147 489.601
R923 GNDA.n2392 GNDA.n2391 473.601
R924 GNDA.n2180 GNDA.n2179 473.601
R925 GNDA.n2393 GNDA.n2392 464
R926 GNDA.n2179 GNDA.n2178 464
R927 GNDA.n2130 GNDA.n2129 463.603
R928 GNDA.n134 GNDA.n133 463.603
R929 GNDA.n2391 GNDA.n171 438.401
R930 GNDA.n2180 GNDA.n2049 438.401
R931 GNDA.n2450 GNDA.n2449 428.8
R932 GNDA.n2393 GNDA.n171 428.8
R933 GNDA.n2178 GNDA.n2049 428.8
R934 GNDA.n2435 GNDA.n2434 422.401
R935 GNDA.n50 GNDA.n49 422.401
R936 GNDA.n78 GNDA.n74 422.401
R937 GNDA.n2124 GNDA.n2123 422.401
R938 GNDA.n441 GNDA.t271 413.084
R939 GNDA.n439 GNDA.t268 413.084
R940 GNDA.n519 GNDA.t248 413.084
R941 GNDA.n517 GNDA.t300 413.084
R942 GNDA.n643 GNDA.t254 413.084
R943 GNDA.n526 GNDA.t274 413.084
R944 GNDA.n173 GNDA.n168 400
R945 GNDA.n168 GNDA.n165 396.8
R946 GNDA.n2158 GNDA.n2060 396.284
R947 GNDA.n2297 GNDA.t219 391.411
R948 GNDA.n1983 GNDA.t219 391.411
R949 GNDA.n173 GNDA.n172 390.401
R950 GNDA.n2165 GNDA.n2050 390.401
R951 GNDA.n2139 GNDA.n2076 390.401
R952 GNDA.n172 GNDA.n165 387.2
R953 GNDA.n2166 GNDA.n2165 387.2
R954 GNDA.n2053 GNDA.n2050 387.2
R955 GNDA.n2166 GNDA.n2053 384
R956 GNDA.n2371 GNDA.n2369 381.642
R957 GNDA.n2415 GNDA.n86 380.8
R958 GNDA.t298 GNDA.t329 372.308
R959 GNDA.t329 GNDA.t119 372.308
R960 GNDA.t119 GNDA.t117 372.308
R961 GNDA.t117 GNDA.t145 372.308
R962 GNDA.t344 GNDA.t145 372.308
R963 GNDA.t344 GNDA.t93 372.308
R964 GNDA.t93 GNDA.t328 372.308
R965 GNDA.t155 GNDA.t100 372.308
R966 GNDA.t126 GNDA.t13 372.308
R967 GNDA.t343 GNDA.t88 372.308
R968 GNDA.t88 GNDA.t87 372.308
R969 GNDA.t144 GNDA.t118 372.308
R970 GNDA.t118 GNDA.t331 372.308
R971 GNDA.t331 GNDA.t134 372.308
R972 GNDA.t295 GNDA.t134 372.308
R973 GNDA.n2021 GNDA.n351 370.214
R974 GNDA.n372 GNDA.n351 365.957
R975 GNDA.n2093 GNDA.n2077 361.601
R976 GNDA.t330 GNDA.n36 355.385
R977 GNDA.n2119 GNDA.t153 355.385
R978 GNDA.n75 GNDA.t157 355.385
R979 GNDA.t21 GNDA.n28 355.385
R980 GNDA.t87 GNDA.n29 355.385
R981 GNDA.n2414 GNDA.n87 352
R982 GNDA.n2094 GNDA.n2093 342.401
R983 GNDA.n2419 GNDA.n87 342.401
R984 GNDA.n2444 GNDA.n32 336
R985 GNDA.n2449 GNDA.n2448 336
R986 GNDA.n2144 GNDA.n2073 332.8
R987 GNDA.n153 GNDA.n97 332.8
R988 GNDA.n63 GNDA.t264 332.75
R989 GNDA.n64 GNDA.t279 332.75
R990 GNDA.n372 GNDA.t219 327.661
R991 GNDA.n2338 GNDA.t219 172.876
R992 GNDA.n2372 GNDA.n2371 323.673
R993 GNDA.n2021 GNDA.t219 323.404
R994 GNDA.n2361 GNDA.t219 172.615
R995 GNDA.n1912 GNDA.n1911 323.2
R996 GNDA.n2146 GNDA.n2145 321.281
R997 GNDA.n152 GNDA.n151 321.281
R998 GNDA.n2145 GNDA.n2144 318.08
R999 GNDA.n153 GNDA.n152 318.08
R1000 GNDA.n1913 GNDA.n1912 316.8
R1001 GNDA.n2136 GNDA.n2135 310.401
R1002 GNDA.n2116 GNDA.n2104 310.401
R1003 GNDA.n2422 GNDA.n83 310.401
R1004 GNDA.n141 GNDA.n101 310.401
R1005 GNDA.n1800 GNDA.n515 304
R1006 GNDA.n2111 GNDA.n2102 304
R1007 GNDA.n148 GNDA.n99 304
R1008 GNDA.n70 GNDA.n69 300.8
R1009 GNDA.n70 GNDA.n62 300.8
R1010 GNDA.n516 GNDA.n515 300.8
R1011 GNDA.n2073 GNDA.n2072 300.8
R1012 GNDA.n149 GNDA.n97 300.8
R1013 GNDA.n2405 GNDA.n2404 297.601
R1014 GNDA.n2163 GNDA.n2057 297.601
R1015 GNDA.n2086 GNDA.n2082 296
R1016 GNDA.n91 GNDA.n90 296
R1017 GNDA.n1800 GNDA.n1799 294.401
R1018 GNDA.n525 GNDA.n524 294.401
R1019 GNDA.n1795 GNDA.n525 294.401
R1020 GNDA.n1914 GNDA.n1911 294.401
R1021 GNDA.n2147 GNDA.n2146 292.5
R1022 GNDA.n2148 GNDA.n2147 292.5
R1023 GNDA.n2145 GNDA.n2071 292.5
R1024 GNDA.n2079 GNDA.n2071 292.5
R1025 GNDA.n2144 GNDA.n2143 292.5
R1026 GNDA.n2143 GNDA.n2142 292.5
R1027 GNDA.n2073 GNDA.n2070 292.5
R1028 GNDA.n2079 GNDA.n2070 292.5
R1029 GNDA.n2076 GNDA.n2074 292.5
R1030 GNDA.n2083 GNDA.n2074 292.5
R1031 GNDA.n2140 GNDA.n2139 292.5
R1032 GNDA.n2141 GNDA.n2140 292.5
R1033 GNDA.n2094 GNDA.n2075 292.5
R1034 GNDA.n2083 GNDA.n2075 292.5
R1035 GNDA.n2093 GNDA.n2092 292.5
R1036 GNDA.n2092 GNDA.n2091 292.5
R1037 GNDA.n2086 GNDA.n2085 292.5
R1038 GNDA.n2085 GNDA.n2084 292.5
R1039 GNDA.n1911 GNDA.n1909 292.5
R1040 GNDA.n1909 GNDA.n310 292.5
R1041 GNDA.n2187 GNDA.n2186 292.5
R1042 GNDA.n2186 GNDA.n2185 292.5
R1043 GNDA.n2183 GNDA.n178 292.5
R1044 GNDA.n2184 GNDA.n2183 292.5
R1045 GNDA.n1921 GNDA.n1920 292.5
R1046 GNDA.n1922 GNDA.n1921 292.5
R1047 GNDA.n2168 GNDA.n2167 292.5
R1048 GNDA.n2169 GNDA.n2168 292.5
R1049 GNDA.n2057 GNDA.n2056 292.5
R1050 GNDA.n2056 GNDA.n2054 292.5
R1051 GNDA.n2163 GNDA.n2162 292.5
R1052 GNDA.n2162 GNDA.n2161 292.5
R1053 GNDA.n2164 GNDA.n2055 292.5
R1054 GNDA.n2055 GNDA.n2054 292.5
R1055 GNDA.n2173 GNDA.n2050 292.5
R1056 GNDA.n2174 GNDA.n2173 292.5
R1057 GNDA.n2172 GNDA.n2053 292.5
R1058 GNDA.n2172 GNDA.n2171 292.5
R1059 GNDA.n2166 GNDA.n2052 292.5
R1060 GNDA.n2170 GNDA.n2052 292.5
R1061 GNDA.n2165 GNDA.n2051 292.5
R1062 GNDA.n2171 GNDA.n2051 292.5
R1063 GNDA.n2181 GNDA.n2180 292.5
R1064 GNDA.n2182 GNDA.n2181 292.5
R1065 GNDA.n2179 GNDA.n312 292.5
R1066 GNDA.n2175 GNDA.n312 292.5
R1067 GNDA.n2178 GNDA.n2177 292.5
R1068 GNDA.n2177 GNDA.n2176 292.5
R1069 GNDA.n2049 GNDA.n311 292.5
R1070 GNDA.n2175 GNDA.n311 292.5
R1071 GNDA.n154 GNDA.n153 292.5
R1072 GNDA.n155 GNDA.n154 292.5
R1073 GNDA.n152 GNDA.n96 292.5
R1074 GNDA.n96 GNDA.n95 292.5
R1075 GNDA.n151 GNDA.n150 292.5
R1076 GNDA.n150 GNDA.n80 292.5
R1077 GNDA.n97 GNDA.n94 292.5
R1078 GNDA.n95 GNDA.n94 292.5
R1079 GNDA.n89 GNDA.n87 292.5
R1080 GNDA.n2409 GNDA.n89 292.5
R1081 GNDA.n2419 GNDA.n2418 292.5
R1082 GNDA.n2418 GNDA.n2417 292.5
R1083 GNDA.n88 GNDA.n86 292.5
R1084 GNDA.n93 GNDA.n88 292.5
R1085 GNDA.n2416 GNDA.n2415 292.5
R1086 GNDA.n2417 GNDA.n2416 292.5
R1087 GNDA.n157 GNDA.n90 292.5
R1088 GNDA.n157 GNDA.n156 292.5
R1089 GNDA.n2369 GNDA.n174 292.5
R1090 GNDA.n2378 GNDA.n2377 292.5
R1091 GNDA.n2377 GNDA.n2376 292.5
R1092 GNDA.n2387 GNDA.n2386 292.5
R1093 GNDA.n2388 GNDA.n2387 292.5
R1094 GNDA.n646 GNDA.n645 292.5
R1095 GNDA.n647 GNDA.n646 292.5
R1096 GNDA.n2406 GNDA.n2405 292.5
R1097 GNDA.n2407 GNDA.n2406 292.5
R1098 GNDA.n2404 GNDA.n163 292.5
R1099 GNDA.n163 GNDA.n161 292.5
R1100 GNDA.n2403 GNDA.n2402 292.5
R1101 GNDA.n2402 GNDA.n2401 292.5
R1102 GNDA.n164 GNDA.n162 292.5
R1103 GNDA.n162 GNDA.n161 292.5
R1104 GNDA.n2399 GNDA.n165 292.5
R1105 GNDA.n2400 GNDA.n2399 292.5
R1106 GNDA.n2398 GNDA.n168 292.5
R1107 GNDA.n2398 GNDA.n2397 292.5
R1108 GNDA.n173 GNDA.n167 292.5
R1109 GNDA.n2396 GNDA.n167 292.5
R1110 GNDA.n172 GNDA.n166 292.5
R1111 GNDA.n2397 GNDA.n166 292.5
R1112 GNDA.n2394 GNDA.n2393 292.5
R1113 GNDA.n2395 GNDA.n2394 292.5
R1114 GNDA.n2392 GNDA.n170 292.5
R1115 GNDA.n2375 GNDA.n170 292.5
R1116 GNDA.n2391 GNDA.n2390 292.5
R1117 GNDA.n2390 GNDA.n2389 292.5
R1118 GNDA.n171 GNDA.n169 292.5
R1119 GNDA.n2375 GNDA.n169 292.5
R1120 GNDA.n1913 GNDA.n1910 292.5
R1121 GNDA.n1910 GNDA.n271 292.5
R1122 GNDA.n1912 GNDA.n444 292.5
R1123 GNDA.n1916 GNDA.n444 292.5
R1124 GNDA.n1915 GNDA.n1914 292.5
R1125 GNDA.n1916 GNDA.n1915 292.5
R1126 GNDA.n2373 GNDA.n2372 292.5
R1127 GNDA.n2370 GNDA.n2368 292.5
R1128 GNDA.n2368 GNDA.n2367 292.5
R1129 GNDA.n2190 GNDA.n2189 292.5
R1130 GNDA.n2191 GNDA.n2190 292.5
R1131 GNDA.n2188 GNDA.n308 292.5
R1132 GNDA.n1916 GNDA.n308 292.5
R1133 GNDA.n309 GNDA.n307 292.5
R1134 GNDA.n1916 GNDA.n307 292.5
R1135 GNDA.n2374 GNDA.n185 292.5
R1136 GNDA.n2374 GNDA.n2373 292.5
R1137 GNDA.n186 GNDA.n183 292.5
R1138 GNDA.n2195 GNDA.n186 292.5
R1139 GNDA.n2379 GNDA.n184 292.5
R1140 GNDA.n2373 GNDA.n184 292.5
R1141 GNDA.n2385 GNDA.n176 292.5
R1142 GNDA.t219 GNDA.n176 292.5
R1143 GNDA.n177 GNDA.n175 292.5
R1144 GNDA.t219 GNDA.n175 292.5
R1145 GNDA.n511 GNDA.n443 292.5
R1146 GNDA.n512 GNDA.n511 292.5
R1147 GNDA.n1919 GNDA.n1918 292.5
R1148 GNDA.n1918 GNDA.n1917 292.5
R1149 GNDA.n1796 GNDA.n1795 292.5
R1150 GNDA.n1796 GNDA.n189 292.5
R1151 GNDA.n525 GNDA.n523 292.5
R1152 GNDA.n523 GNDA.t219 292.5
R1153 GNDA.n524 GNDA.n522 292.5
R1154 GNDA.n522 GNDA.n521 292.5
R1155 GNDA.n1798 GNDA.n1797 292.5
R1156 GNDA.n1797 GNDA.t219 292.5
R1157 GNDA.n529 GNDA.n528 292.5
R1158 GNDA.n529 GNDA.n188 292.5
R1159 GNDA.n1794 GNDA.n1793 292.5
R1160 GNDA.n1793 GNDA.n1792 292.5
R1161 GNDA.n1790 GNDA.n516 292.5
R1162 GNDA.n1791 GNDA.n1790 292.5
R1163 GNDA.n1799 GNDA.n514 292.5
R1164 GNDA.n514 GNDA.t219 292.5
R1165 GNDA.n1801 GNDA.n1800 292.5
R1166 GNDA.n1802 GNDA.n1801 292.5
R1167 GNDA.n515 GNDA.n513 292.5
R1168 GNDA.n513 GNDA.t219 292.5
R1169 GNDA.n2120 GNDA.n72 292.5
R1170 GNDA.n2120 GNDA.n2119 292.5
R1171 GNDA.n2126 GNDA.n2125 292.5
R1172 GNDA.n2127 GNDA.n2126 292.5
R1173 GNDA.n2428 GNDA.n2427 292.5
R1174 GNDA.n2427 GNDA.n2426 292.5
R1175 GNDA.n2429 GNDA.n76 292.5
R1176 GNDA.n76 GNDA.n75 292.5
R1177 GNDA.n69 GNDA.n68 292.5
R1178 GNDA.n68 GNDA.n28 292.5
R1179 GNDA.n70 GNDA.n38 292.5
R1180 GNDA.n2439 GNDA.n38 292.5
R1181 GNDA.n62 GNDA.n61 292.5
R1182 GNDA.n61 GNDA.n36 292.5
R1183 GNDA.n66 GNDA.n37 292.5
R1184 GNDA.n2439 GNDA.n37 292.5
R1185 GNDA.n2116 GNDA.n2106 292.5
R1186 GNDA.n2130 GNDA.n2106 292.5
R1187 GNDA.n2118 GNDA.n2117 292.5
R1188 GNDA.n2131 GNDA.n2118 292.5
R1189 GNDA.n2111 GNDA.n2105 292.5
R1190 GNDA.n2107 GNDA.n2105 292.5
R1191 GNDA.n2133 GNDA.n2132 292.5
R1192 GNDA.n2132 GNDA.n2131 292.5
R1193 GNDA.n2452 GNDA.n2451 292.5
R1194 GNDA.n2453 GNDA.n2452 292.5
R1195 GNDA.n2449 GNDA.n31 292.5
R1196 GNDA.n2439 GNDA.n31 292.5
R1197 GNDA.n2448 GNDA.n2447 292.5
R1198 GNDA.n2447 GNDA.n2446 292.5
R1199 GNDA.n2443 GNDA.n35 292.5
R1200 GNDA.n2128 GNDA.n35 292.5
R1201 GNDA.n2445 GNDA.n2444 292.5
R1202 GNDA.n2446 GNDA.n2445 292.5
R1203 GNDA.n32 GNDA.n30 292.5
R1204 GNDA.n2439 GNDA.n30 292.5
R1205 GNDA.n148 GNDA.n100 292.5
R1206 GNDA.n100 GNDA.n81 292.5
R1207 GNDA.n147 GNDA.n146 292.5
R1208 GNDA.n146 GNDA.n145 292.5
R1209 GNDA.n132 GNDA.n101 292.5
R1210 GNDA.n134 GNDA.n132 292.5
R1211 GNDA.n144 GNDA.n143 292.5
R1212 GNDA.n145 GNDA.n144 292.5
R1213 GNDA.n2436 GNDA.n41 292.5
R1214 GNDA.n133 GNDA.n41 292.5
R1215 GNDA.n2438 GNDA.n2437 292.5
R1216 GNDA.n2439 GNDA.n2438 292.5
R1217 GNDA.n42 GNDA.n40 292.5
R1218 GNDA.n2129 GNDA.n40 292.5
R1219 GNDA.n2432 GNDA.n39 292.5
R1220 GNDA.n2439 GNDA.n39 292.5
R1221 GNDA.n2135 GNDA.n2098 292.5
R1222 GNDA.t65 GNDA.n2098 292.5
R1223 GNDA.n2110 GNDA.n2109 292.5
R1224 GNDA.t65 GNDA.n2110 292.5
R1225 GNDA.n135 GNDA.n83 292.5
R1226 GNDA.t312 GNDA.n135 292.5
R1227 GNDA.n139 GNDA.n138 292.5
R1228 GNDA.t312 GNDA.n139 292.5
R1229 GNDA.n2456 GNDA.n2455 292.5
R1230 GNDA.n2455 GNDA.n2454 292.5
R1231 GNDA.n26 GNDA.n25 292.5
R1232 GNDA.n2439 GNDA.n26 292.5
R1233 GNDA.n2441 GNDA.n2440 292.5
R1234 GNDA.n2442 GNDA.n2441 292.5
R1235 GNDA.n27 GNDA.n24 292.5
R1236 GNDA.n2439 GNDA.n27 292.5
R1237 GNDA.n2405 GNDA.n164 291.2
R1238 GNDA.n2404 GNDA.n2403 291.2
R1239 GNDA.n2164 GNDA.n2163 291.2
R1240 GNDA.n2167 GNDA.n2057 291.2
R1241 GNDA.n1799 GNDA.n516 291.2
R1242 GNDA.n1914 GNDA.n1913 288
R1243 GNDA.n2403 GNDA.n164 284.8
R1244 GNDA.n2167 GNDA.n2164 284.8
R1245 GNDA.n442 GNDA.n440 281.601
R1246 GNDA.n644 GNDA.n527 281.601
R1247 GNDA.n1920 GNDA.n1919 278.401
R1248 GNDA.n645 GNDA.n528 278.401
R1249 GNDA.t28 GNDA.t162 271.649
R1250 GNDA.t332 GNDA.t44 271.649
R1251 GNDA.n1923 GNDA.n430 264.301
R1252 GNDA.n1923 GNDA.n423 264.301
R1253 GNDA.n503 GNDA.n502 264.301
R1254 GNDA.n1772 GNDA.n640 264.301
R1255 GNDA.n1766 GNDA.n1765 264.301
R1256 GNDA.n1095 GNDA.n1094 264.301
R1257 GNDA.n1131 GNDA.n1108 259.416
R1258 GNDA.n1743 GNDA.n1742 259.416
R1259 GNDA.n347 GNDA.n345 259.416
R1260 GNDA.n1486 GNDA.n1485 259.416
R1261 GNDA.n2323 GNDA.n2322 259.416
R1262 GNDA.n1951 GNDA.n399 259.416
R1263 GNDA.n1738 GNDA.n1171 259.416
R1264 GNDA.n2314 GNDA.n224 259.416
R1265 GNDA.n1072 GNDA.n1071 259.416
R1266 GNDA.n63 GNDA.t266 258.601
R1267 GNDA.n64 GNDA.t281 258.601
R1268 GNDA.n589 GNDA.n556 258.334
R1269 GNDA.n1306 GNDA.n1305 258.334
R1270 GNDA.n913 GNDA.n912 258.334
R1271 GNDA.n1391 GNDA.n1390 258.334
R1272 GNDA.n2254 GNDA.n2253 258.334
R1273 GNDA.n998 GNDA.n823 258.334
R1274 GNDA.n1610 GNDA.n1565 258.334
R1275 GNDA.n1840 GNDA.n1817 258.334
R1276 GNDA.n737 GNDA.n703 258.334
R1277 GNDA.n1923 GNDA.n424 254.34
R1278 GNDA.n1923 GNDA.n425 254.34
R1279 GNDA.n1923 GNDA.n426 254.34
R1280 GNDA.n1923 GNDA.n427 254.34
R1281 GNDA.n1923 GNDA.n428 254.34
R1282 GNDA.n1924 GNDA.n1923 254.34
R1283 GNDA.n1923 GNDA.n418 254.34
R1284 GNDA.n1923 GNDA.n419 254.34
R1285 GNDA.n1923 GNDA.n420 254.34
R1286 GNDA.n1923 GNDA.n421 254.34
R1287 GNDA.n1923 GNDA.n431 254.34
R1288 GNDA.n1923 GNDA.n432 254.34
R1289 GNDA.n1923 GNDA.n433 254.34
R1290 GNDA.n1923 GNDA.n434 254.34
R1291 GNDA.n1923 GNDA.n435 254.34
R1292 GNDA.n1923 GNDA.n436 254.34
R1293 GNDA.n1199 GNDA.n1198 254.34
R1294 GNDA.n1198 GNDA.n1197 254.34
R1295 GNDA.n1198 GNDA.n1196 254.34
R1296 GNDA.n1198 GNDA.n1195 254.34
R1297 GNDA.n1198 GNDA.n1194 254.34
R1298 GNDA.n1198 GNDA.n1193 254.34
R1299 GNDA.n1733 GNDA.n1732 254.34
R1300 GNDA.n1732 GNDA.n1177 254.34
R1301 GNDA.n1732 GNDA.n1178 254.34
R1302 GNDA.n1732 GNDA.n1179 254.34
R1303 GNDA.n1732 GNDA.n1180 254.34
R1304 GNDA.n1740 GNDA.n1739 254.34
R1305 GNDA.n1740 GNDA.n1169 254.34
R1306 GNDA.n1740 GNDA.n1168 254.34
R1307 GNDA.n1740 GNDA.n1167 254.34
R1308 GNDA.n1740 GNDA.n1166 254.34
R1309 GNDA.n1740 GNDA.n1165 254.34
R1310 GNDA.n1740 GNDA.n1164 254.34
R1311 GNDA.n1740 GNDA.n1163 254.34
R1312 GNDA.n1740 GNDA.n1162 254.34
R1313 GNDA.n1740 GNDA.n1161 254.34
R1314 GNDA.n1740 GNDA.n1160 254.34
R1315 GNDA.n1740 GNDA.n1159 254.34
R1316 GNDA.n1741 GNDA.n1740 254.34
R1317 GNDA.n1740 GNDA.n1158 254.34
R1318 GNDA.n1740 GNDA.n1157 254.34
R1319 GNDA.n1740 GNDA.n1156 254.34
R1320 GNDA.n1740 GNDA.n1155 254.34
R1321 GNDA.n1740 GNDA.n1154 254.34
R1322 GNDA.n1032 GNDA.n1031 254.34
R1323 GNDA.n1032 GNDA.n780 254.34
R1324 GNDA.n1032 GNDA.n779 254.34
R1325 GNDA.n1032 GNDA.n778 254.34
R1326 GNDA.n1032 GNDA.n777 254.34
R1327 GNDA.n1032 GNDA.n776 254.34
R1328 GNDA.n1032 GNDA.n775 254.34
R1329 GNDA.n1032 GNDA.n774 254.34
R1330 GNDA.n1032 GNDA.n773 254.34
R1331 GNDA.n1032 GNDA.n772 254.34
R1332 GNDA.n1032 GNDA.n771 254.34
R1333 GNDA.n1032 GNDA.n770 254.34
R1334 GNDA.n2316 GNDA.n2315 254.34
R1335 GNDA.n2316 GNDA.n222 254.34
R1336 GNDA.n2316 GNDA.n221 254.34
R1337 GNDA.n2316 GNDA.n220 254.34
R1338 GNDA.n2316 GNDA.n219 254.34
R1339 GNDA.n2316 GNDA.n218 254.34
R1340 GNDA.n2316 GNDA.n205 254.34
R1341 GNDA.n2317 GNDA.n2316 254.34
R1342 GNDA.n2316 GNDA.n217 254.34
R1343 GNDA.n2316 GNDA.n216 254.34
R1344 GNDA.n2316 GNDA.n215 254.34
R1345 GNDA.n2316 GNDA.n214 254.34
R1346 GNDA.n2316 GNDA.n213 254.34
R1347 GNDA.n2316 GNDA.n212 254.34
R1348 GNDA.n2316 GNDA.n211 254.34
R1349 GNDA.n2316 GNDA.n210 254.34
R1350 GNDA.n2316 GNDA.n209 254.34
R1351 GNDA.n2316 GNDA.n208 254.34
R1352 GNDA.n1669 GNDA.n1547 254.34
R1353 GNDA.n1683 GNDA.n1547 254.34
R1354 GNDA.n1685 GNDA.n1547 254.34
R1355 GNDA.n1698 GNDA.n1547 254.34
R1356 GNDA.n1700 GNDA.n1547 254.34
R1357 GNDA.n1710 GNDA.n1547 254.34
R1358 GNDA.n1547 GNDA.n1546 254.34
R1359 GNDA.n1547 GNDA.n1215 254.34
R1360 GNDA.n1547 GNDA.n1214 254.34
R1361 GNDA.n1547 GNDA.n1213 254.34
R1362 GNDA.n1547 GNDA.n1212 254.34
R1363 GNDA.n1547 GNDA.n1211 254.34
R1364 GNDA.n1547 GNDA.n1210 254.34
R1365 GNDA.n1547 GNDA.n1209 254.34
R1366 GNDA.n1547 GNDA.n1208 254.34
R1367 GNDA.n1547 GNDA.n1207 254.34
R1368 GNDA.n1547 GNDA.n1206 254.34
R1369 GNDA.n1547 GNDA.n1205 254.34
R1370 GNDA.n1769 GNDA.n1768 254.34
R1371 GNDA.n1768 GNDA.n1104 254.34
R1372 GNDA.n1768 GNDA.n1105 254.34
R1373 GNDA.n1768 GNDA.n1106 254.34
R1374 GNDA.n1768 GNDA.n1107 254.34
R1375 GNDA.n1768 GNDA.n1149 254.34
R1376 GNDA.n1768 GNDA.n1102 254.34
R1377 GNDA.n1768 GNDA.n1101 254.34
R1378 GNDA.n1768 GNDA.n1100 254.34
R1379 GNDA.n1768 GNDA.n1099 254.34
R1380 GNDA.n1768 GNDA.n1098 254.34
R1381 GNDA.n1768 GNDA.n1097 254.34
R1382 GNDA.n1032 GNDA.n769 254.34
R1383 GNDA.n1032 GNDA.n661 254.34
R1384 GNDA.n1032 GNDA.n660 254.34
R1385 GNDA.n1032 GNDA.n659 254.34
R1386 GNDA.n1032 GNDA.n658 254.34
R1387 GNDA.n1033 GNDA.n1032 254.34
R1388 GNDA.n1768 GNDA.n653 254.34
R1389 GNDA.n1768 GNDA.n652 254.34
R1390 GNDA.n1768 GNDA.n651 254.34
R1391 GNDA.n1768 GNDA.n650 254.34
R1392 GNDA.n1768 GNDA.n649 254.34
R1393 GNDA.n1768 GNDA.n648 254.34
R1394 GNDA.n373 GNDA.n372 254.34
R1395 GNDA.n372 GNDA.n371 254.34
R1396 GNDA.n372 GNDA.n370 254.34
R1397 GNDA.n372 GNDA.n369 254.34
R1398 GNDA.n372 GNDA.n368 254.34
R1399 GNDA.n372 GNDA.n367 254.34
R1400 GNDA.n2022 GNDA.n2021 254.34
R1401 GNDA.n2021 GNDA.n2020 254.34
R1402 GNDA.n2021 GNDA.n355 254.34
R1403 GNDA.n2021 GNDA.n354 254.34
R1404 GNDA.n2021 GNDA.n353 254.34
R1405 GNDA.n2021 GNDA.n352 254.34
R1406 GNDA.n1536 GNDA.n1534 254.34
R1407 GNDA.n1534 GNDA.n1532 254.34
R1408 GNDA.n1534 GNDA.n1455 254.34
R1409 GNDA.n1534 GNDA.n1454 254.34
R1410 GNDA.n1534 GNDA.n1453 254.34
R1411 GNDA.n1534 GNDA.n1452 254.34
R1412 GNDA.n1508 GNDA.n1448 254.34
R1413 GNDA.n1516 GNDA.n1448 254.34
R1414 GNDA.n1518 GNDA.n1448 254.34
R1415 GNDA.n1526 GNDA.n1448 254.34
R1416 GNDA.n1528 GNDA.n1448 254.34
R1417 GNDA.n1540 GNDA.n1448 254.34
R1418 GNDA.n2339 GNDA.n2338 254.34
R1419 GNDA.n2338 GNDA.n2337 254.34
R1420 GNDA.n2338 GNDA.n2336 254.34
R1421 GNDA.n2338 GNDA.n2335 254.34
R1422 GNDA.n2338 GNDA.n2334 254.34
R1423 GNDA.n2338 GNDA.n2333 254.34
R1424 GNDA.n2361 GNDA.n2360 254.34
R1425 GNDA.n2361 GNDA.n197 254.34
R1426 GNDA.n2361 GNDA.n198 254.34
R1427 GNDA.n2361 GNDA.n199 254.34
R1428 GNDA.n2361 GNDA.n200 254.34
R1429 GNDA.t219 GNDA.n335 250.349
R1430 GNDA.n2359 GNDA.n203 249.663
R1431 GNDA.n1509 GNDA.n1507 249.663
R1432 GNDA.n1969 GNDA.n401 249.663
R1433 GNDA.n1734 GNDA.n1175 249.663
R1434 GNDA.n2310 GNDA.n244 249.663
R1435 GNDA.n1929 GNDA.n415 249.663
R1436 GNDA.n1645 GNDA.n1644 249.663
R1437 GNDA.n480 GNDA.n479 249.663
R1438 GNDA.n2023 GNDA.n349 249.663
R1439 GNDA.n1919 GNDA.n443 240
R1440 GNDA.n1794 GNDA.n528 240
R1441 GNDA.n2137 GNDA.n2096 240
R1442 GNDA.n2421 GNDA.n85 240
R1443 GNDA.t330 GNDA.t280 236.923
R1444 GNDA.t116 GNDA.t56 236.923
R1445 GNDA.t22 GNDA.t128 236.923
R1446 GNDA.t228 GNDA.t153 236.923
R1447 GNDA.t157 GNDA.t286 236.923
R1448 GNDA.t352 GNDA.t92 236.923
R1449 GNDA.t41 GNDA.t15 236.923
R1450 GNDA.t21 GNDA.t265 236.923
R1451 GNDA.n2444 GNDA.n2443 233.601
R1452 GNDA.n57 GNDA.n55 227.096
R1453 GNDA.n54 GNDA.n52 227.096
R1454 GNDA.n57 GNDA.n56 226.534
R1455 GNDA.n54 GNDA.n53 226.534
R1456 GNDA.n2088 GNDA.n2087 225.601
R1457 GNDA.n2413 GNDA.n2412 225.601
R1458 GNDA.n2101 GNDA.t234 224.525
R1459 GNDA.n2103 GNDA.t305 224.525
R1460 GNDA.n98 GNDA.t253 224.525
R1461 GNDA.n140 GNDA.t259 224.525
R1462 GNDA.n2456 GNDA.n25 224
R1463 GNDA.n60 GNDA.n59 222.034
R1464 GNDA.n2440 GNDA.n25 220.8
R1465 GNDA.n66 GNDA.n65 211.201
R1466 GNDA.n67 GNDA.n66 211.201
R1467 GNDA.n2109 GNDA.n2096 211.201
R1468 GNDA.n2109 GNDA.n2100 211.201
R1469 GNDA.n138 GNDA.n137 211.201
R1470 GNDA.n138 GNDA.n85 211.201
R1471 GNDA.n2440 GNDA.n24 209.601
R1472 GNDA.n2457 GNDA.n2456 208
R1473 GNDA.n14 GNDA.n12 206.052
R1474 GNDA.n3 GNDA.n1 206.052
R1475 GNDA.n22 GNDA.n21 205.488
R1476 GNDA.n20 GNDA.n19 205.488
R1477 GNDA.n18 GNDA.n17 205.488
R1478 GNDA.n16 GNDA.n15 205.488
R1479 GNDA.n14 GNDA.n13 205.488
R1480 GNDA.n11 GNDA.n10 205.488
R1481 GNDA.n9 GNDA.n8 205.488
R1482 GNDA.n7 GNDA.n6 205.488
R1483 GNDA.n5 GNDA.n4 205.488
R1484 GNDA.n3 GNDA.n2 205.488
R1485 GNDA.n1103 GNDA.n541 197
R1486 GNDA.n1767 GNDA.n1150 197
R1487 GNDA.n2039 GNDA.n2038 197
R1488 GNDA.n846 GNDA.n379 197
R1489 GNDA.n1444 GNDA.n1217 197
R1490 GNDA.n2365 GNDA.n191 197
R1491 GNDA.n941 GNDA.n380 197
R1492 GNDA.n1711 GNDA.n1203 197
R1493 GNDA.n1804 GNDA.n266 197
R1494 GNDA.n1096 GNDA.n654 197
R1495 GNDA.n2082 GNDA.n2081 195
R1496 GNDA.n2081 GNDA.n2080 195
R1497 GNDA.n2089 GNDA.n2088 195
R1498 GNDA.n2090 GNDA.n2089 195
R1499 GNDA.n2412 GNDA.n2411 195
R1500 GNDA.n2411 GNDA.n2410 195
R1501 GNDA.n92 GNDA.n91 195
R1502 GNDA.n95 GNDA.n92 195
R1503 GNDA.n2133 GNDA.n2104 192
R1504 GNDA.n143 GNDA.n141 192
R1505 GNDA.n2363 GNDA.n194 187.249
R1506 GNDA.n1542 GNDA.n1219 187.249
R1507 GNDA.n1998 GNDA.n382 187.249
R1508 GNDA.n1545 GNDA.n1544 187.249
R1509 GNDA.n2283 GNDA.n2282 187.249
R1510 GNDA.n1030 GNDA.n782 187.249
R1511 GNDA.n1670 GNDA.n1668 187.249
R1512 GNDA.n505 GNDA.n437 187.249
R1513 GNDA.n2000 GNDA.n376 187.249
R1514 GNDA.n2439 GNDA.t100 186.155
R1515 GNDA.n2439 GNDA.t13 186.155
R1516 GNDA.n591 GNDA.n556 185
R1517 GNDA.n606 GNDA.n605 185
R1518 GNDA.n604 GNDA.n557 185
R1519 GNDA.n603 GNDA.n602 185
R1520 GNDA.n601 GNDA.n600 185
R1521 GNDA.n599 GNDA.n598 185
R1522 GNDA.n597 GNDA.n596 185
R1523 GNDA.n595 GNDA.n594 185
R1524 GNDA.n593 GNDA.n592 185
R1525 GNDA.n574 GNDA.n573 185
R1526 GNDA.n576 GNDA.n575 185
R1527 GNDA.n578 GNDA.n577 185
R1528 GNDA.n580 GNDA.n579 185
R1529 GNDA.n582 GNDA.n581 185
R1530 GNDA.n584 GNDA.n583 185
R1531 GNDA.n586 GNDA.n585 185
R1532 GNDA.n588 GNDA.n587 185
R1533 GNDA.n590 GNDA.n589 185
R1534 GNDA.n639 GNDA.n638 185
R1535 GNDA.n558 GNDA.n543 185
R1536 GNDA.n560 GNDA.n559 185
R1537 GNDA.n562 GNDA.n561 185
R1538 GNDA.n564 GNDA.n563 185
R1539 GNDA.n566 GNDA.n565 185
R1540 GNDA.n568 GNDA.n567 185
R1541 GNDA.n570 GNDA.n569 185
R1542 GNDA.n572 GNDA.n571 185
R1543 GNDA.n637 GNDA.n542 185
R1544 GNDA.n635 GNDA.n634 185
R1545 GNDA.n609 GNDA.n608 185
R1546 GNDA.n624 GNDA.n623 185
R1547 GNDA.n621 GNDA.n614 185
R1548 GNDA.n619 GNDA.n618 185
R1549 GNDA.n615 GNDA.n537 185
R1550 GNDA.n1783 GNDA.n1782 185
R1551 GNDA.n1785 GNDA.n1784 185
R1552 GNDA.n1307 GNDA.n1306 185
R1553 GNDA.n1309 GNDA.n1308 185
R1554 GNDA.n1311 GNDA.n1310 185
R1555 GNDA.n1313 GNDA.n1312 185
R1556 GNDA.n1315 GNDA.n1314 185
R1557 GNDA.n1317 GNDA.n1316 185
R1558 GNDA.n1319 GNDA.n1318 185
R1559 GNDA.n1321 GNDA.n1320 185
R1560 GNDA.n1322 GNDA.n1220 185
R1561 GNDA.n1289 GNDA.n1288 185
R1562 GNDA.n1291 GNDA.n1290 185
R1563 GNDA.n1293 GNDA.n1292 185
R1564 GNDA.n1295 GNDA.n1294 185
R1565 GNDA.n1297 GNDA.n1296 185
R1566 GNDA.n1299 GNDA.n1298 185
R1567 GNDA.n1301 GNDA.n1300 185
R1568 GNDA.n1303 GNDA.n1302 185
R1569 GNDA.n1305 GNDA.n1304 185
R1570 GNDA.n1271 GNDA.n1270 185
R1571 GNDA.n1273 GNDA.n1272 185
R1572 GNDA.n1275 GNDA.n1274 185
R1573 GNDA.n1277 GNDA.n1276 185
R1574 GNDA.n1279 GNDA.n1278 185
R1575 GNDA.n1281 GNDA.n1280 185
R1576 GNDA.n1283 GNDA.n1282 185
R1577 GNDA.n1285 GNDA.n1284 185
R1578 GNDA.n1287 GNDA.n1286 185
R1579 GNDA.n1269 GNDA.n1268 185
R1580 GNDA.n1263 GNDA.n1262 185
R1581 GNDA.n1261 GNDA.n1260 185
R1582 GNDA.n1256 GNDA.n1255 185
R1583 GNDA.n1254 GNDA.n1253 185
R1584 GNDA.n1248 GNDA.n1247 185
R1585 GNDA.n1243 GNDA.n1224 185
R1586 GNDA.n1326 GNDA.n1325 185
R1587 GNDA.n1223 GNDA.n1221 185
R1588 GNDA.n914 GNDA.n913 185
R1589 GNDA.n916 GNDA.n915 185
R1590 GNDA.n918 GNDA.n917 185
R1591 GNDA.n920 GNDA.n919 185
R1592 GNDA.n922 GNDA.n921 185
R1593 GNDA.n924 GNDA.n923 185
R1594 GNDA.n926 GNDA.n925 185
R1595 GNDA.n928 GNDA.n927 185
R1596 GNDA.n929 GNDA.n825 185
R1597 GNDA.n896 GNDA.n895 185
R1598 GNDA.n898 GNDA.n897 185
R1599 GNDA.n900 GNDA.n899 185
R1600 GNDA.n902 GNDA.n901 185
R1601 GNDA.n904 GNDA.n903 185
R1602 GNDA.n906 GNDA.n905 185
R1603 GNDA.n908 GNDA.n907 185
R1604 GNDA.n910 GNDA.n909 185
R1605 GNDA.n912 GNDA.n911 185
R1606 GNDA.n878 GNDA.n877 185
R1607 GNDA.n880 GNDA.n879 185
R1608 GNDA.n882 GNDA.n881 185
R1609 GNDA.n884 GNDA.n883 185
R1610 GNDA.n886 GNDA.n885 185
R1611 GNDA.n888 GNDA.n887 185
R1612 GNDA.n890 GNDA.n889 185
R1613 GNDA.n892 GNDA.n891 185
R1614 GNDA.n894 GNDA.n893 185
R1615 GNDA.n876 GNDA.n875 185
R1616 GNDA.n870 GNDA.n869 185
R1617 GNDA.n868 GNDA.n867 185
R1618 GNDA.n863 GNDA.n862 185
R1619 GNDA.n861 GNDA.n860 185
R1620 GNDA.n855 GNDA.n854 185
R1621 GNDA.n850 GNDA.n829 185
R1622 GNDA.n933 GNDA.n932 185
R1623 GNDA.n828 GNDA.n826 185
R1624 GNDA.n1392 GNDA.n1391 185
R1625 GNDA.n1394 GNDA.n1393 185
R1626 GNDA.n1396 GNDA.n1395 185
R1627 GNDA.n1398 GNDA.n1397 185
R1628 GNDA.n1400 GNDA.n1399 185
R1629 GNDA.n1402 GNDA.n1401 185
R1630 GNDA.n1404 GNDA.n1403 185
R1631 GNDA.n1406 GNDA.n1405 185
R1632 GNDA.n1407 GNDA.n1355 185
R1633 GNDA.n1374 GNDA.n1373 185
R1634 GNDA.n1376 GNDA.n1375 185
R1635 GNDA.n1378 GNDA.n1377 185
R1636 GNDA.n1380 GNDA.n1379 185
R1637 GNDA.n1382 GNDA.n1381 185
R1638 GNDA.n1384 GNDA.n1383 185
R1639 GNDA.n1386 GNDA.n1385 185
R1640 GNDA.n1388 GNDA.n1387 185
R1641 GNDA.n1390 GNDA.n1389 185
R1642 GNDA.n1347 GNDA.n1333 185
R1643 GNDA.n1358 GNDA.n1357 185
R1644 GNDA.n1360 GNDA.n1359 185
R1645 GNDA.n1362 GNDA.n1361 185
R1646 GNDA.n1364 GNDA.n1363 185
R1647 GNDA.n1366 GNDA.n1365 185
R1648 GNDA.n1368 GNDA.n1367 185
R1649 GNDA.n1370 GNDA.n1369 185
R1650 GNDA.n1372 GNDA.n1371 185
R1651 GNDA.n1337 GNDA.n1334 185
R1652 GNDA.n1438 GNDA.n1437 185
R1653 GNDA.n1412 GNDA.n1336 185
R1654 GNDA.n1418 GNDA.n1417 185
R1655 GNDA.n1416 GNDA.n1411 185
R1656 GNDA.n1425 GNDA.n1424 185
R1657 GNDA.n1423 GNDA.n1410 185
R1658 GNDA.n1430 GNDA.n1356 185
R1659 GNDA.n1434 GNDA.n1433 185
R1660 GNDA.n2255 GNDA.n2254 185
R1661 GNDA.n2257 GNDA.n2256 185
R1662 GNDA.n2259 GNDA.n2258 185
R1663 GNDA.n2261 GNDA.n2260 185
R1664 GNDA.n2263 GNDA.n2262 185
R1665 GNDA.n2265 GNDA.n2264 185
R1666 GNDA.n2267 GNDA.n2266 185
R1667 GNDA.n2268 GNDA.n293 185
R1668 GNDA.n2272 GNDA.n2271 185
R1669 GNDA.n2237 GNDA.n2236 185
R1670 GNDA.n2239 GNDA.n2238 185
R1671 GNDA.n2241 GNDA.n2240 185
R1672 GNDA.n2243 GNDA.n2242 185
R1673 GNDA.n2245 GNDA.n2244 185
R1674 GNDA.n2247 GNDA.n2246 185
R1675 GNDA.n2249 GNDA.n2248 185
R1676 GNDA.n2251 GNDA.n2250 185
R1677 GNDA.n2253 GNDA.n2252 185
R1678 GNDA.n2219 GNDA.n2218 185
R1679 GNDA.n2221 GNDA.n2220 185
R1680 GNDA.n2223 GNDA.n2222 185
R1681 GNDA.n2225 GNDA.n2224 185
R1682 GNDA.n2227 GNDA.n2226 185
R1683 GNDA.n2229 GNDA.n2228 185
R1684 GNDA.n2231 GNDA.n2230 185
R1685 GNDA.n2233 GNDA.n2232 185
R1686 GNDA.n2235 GNDA.n2234 185
R1687 GNDA.n2217 GNDA.n2216 185
R1688 GNDA.n2207 GNDA.n2206 185
R1689 GNDA.n2205 GNDA.n2204 185
R1690 GNDA.n2202 GNDA.n2201 185
R1691 GNDA.n2200 GNDA.n2199 185
R1692 GNDA.n302 GNDA.n301 185
R1693 GNDA.n300 GNDA.n276 185
R1694 GNDA.n2276 GNDA.n2275 185
R1695 GNDA.n275 GNDA.n273 185
R1696 GNDA.n1000 GNDA.n823 185
R1697 GNDA.n1014 GNDA.n1013 185
R1698 GNDA.n1012 GNDA.n824 185
R1699 GNDA.n1011 GNDA.n1010 185
R1700 GNDA.n1009 GNDA.n1008 185
R1701 GNDA.n1007 GNDA.n1006 185
R1702 GNDA.n1005 GNDA.n1004 185
R1703 GNDA.n1003 GNDA.n1002 185
R1704 GNDA.n1001 GNDA.n800 185
R1705 GNDA.n983 GNDA.n982 185
R1706 GNDA.n985 GNDA.n984 185
R1707 GNDA.n987 GNDA.n986 185
R1708 GNDA.n989 GNDA.n988 185
R1709 GNDA.n991 GNDA.n990 185
R1710 GNDA.n993 GNDA.n992 185
R1711 GNDA.n995 GNDA.n994 185
R1712 GNDA.n997 GNDA.n996 185
R1713 GNDA.n999 GNDA.n998 185
R1714 GNDA.n965 GNDA.n964 185
R1715 GNDA.n967 GNDA.n966 185
R1716 GNDA.n969 GNDA.n968 185
R1717 GNDA.n971 GNDA.n970 185
R1718 GNDA.n973 GNDA.n972 185
R1719 GNDA.n975 GNDA.n974 185
R1720 GNDA.n977 GNDA.n976 185
R1721 GNDA.n979 GNDA.n978 185
R1722 GNDA.n981 GNDA.n980 185
R1723 GNDA.n963 GNDA.n962 185
R1724 GNDA.n957 GNDA.n956 185
R1725 GNDA.n955 GNDA.n954 185
R1726 GNDA.n950 GNDA.n949 185
R1727 GNDA.n945 GNDA.n808 185
R1728 GNDA.n1018 GNDA.n1017 185
R1729 GNDA.n807 GNDA.n805 185
R1730 GNDA.n1024 GNDA.n1023 185
R1731 GNDA.n1026 GNDA.n1025 185
R1732 GNDA.n1610 GNDA.n1609 185
R1733 GNDA.n1612 GNDA.n1564 185
R1734 GNDA.n1615 GNDA.n1614 185
R1735 GNDA.n1616 GNDA.n1563 185
R1736 GNDA.n1618 GNDA.n1617 185
R1737 GNDA.n1620 GNDA.n1562 185
R1738 GNDA.n1623 GNDA.n1622 185
R1739 GNDA.n1624 GNDA.n1561 185
R1740 GNDA.n1675 GNDA.n1674 185
R1741 GNDA.n1592 GNDA.n1569 185
R1742 GNDA.n1594 GNDA.n1593 185
R1743 GNDA.n1596 GNDA.n1568 185
R1744 GNDA.n1599 GNDA.n1598 185
R1745 GNDA.n1600 GNDA.n1567 185
R1746 GNDA.n1602 GNDA.n1601 185
R1747 GNDA.n1604 GNDA.n1566 185
R1748 GNDA.n1607 GNDA.n1606 185
R1749 GNDA.n1608 GNDA.n1565 185
R1750 GNDA.n1576 GNDA.n1550 185
R1751 GNDA.n1577 GNDA.n1575 185
R1752 GNDA.n1579 GNDA.n1578 185
R1753 GNDA.n1581 GNDA.n1572 185
R1754 GNDA.n1583 GNDA.n1582 185
R1755 GNDA.n1584 GNDA.n1571 185
R1756 GNDA.n1586 GNDA.n1585 185
R1757 GNDA.n1588 GNDA.n1570 185
R1758 GNDA.n1591 GNDA.n1590 185
R1759 GNDA.n1707 GNDA.n1706 185
R1760 GNDA.n1704 GNDA.n1703 185
R1761 GNDA.n1552 GNDA.n1551 185
R1762 GNDA.n1695 GNDA.n1694 185
R1763 GNDA.n1692 GNDA.n1555 185
R1764 GNDA.n1690 GNDA.n1689 185
R1765 GNDA.n1557 GNDA.n1556 185
R1766 GNDA.n1680 GNDA.n1679 185
R1767 GNDA.n1677 GNDA.n1560 185
R1768 GNDA.n1838 GNDA.n1817 185
R1769 GNDA.n1837 GNDA.n1836 185
R1770 GNDA.n1835 GNDA.n1818 185
R1771 GNDA.n1833 GNDA.n1832 185
R1772 GNDA.n1831 GNDA.n1820 185
R1773 GNDA.n1830 GNDA.n1829 185
R1774 GNDA.n1827 GNDA.n1821 185
R1775 GNDA.n1825 GNDA.n1824 185
R1776 GNDA.n1823 GNDA.n1822 185
R1777 GNDA.n1856 GNDA.n1855 185
R1778 GNDA.n1854 GNDA.n1813 185
R1779 GNDA.n1853 GNDA.n1852 185
R1780 GNDA.n1850 GNDA.n1814 185
R1781 GNDA.n1848 GNDA.n1847 185
R1782 GNDA.n1846 GNDA.n1815 185
R1783 GNDA.n1845 GNDA.n1844 185
R1784 GNDA.n1842 GNDA.n1816 185
R1785 GNDA.n1840 GNDA.n1839 185
R1786 GNDA.n1876 GNDA.n1875 185
R1787 GNDA.n1871 GNDA.n1808 185
R1788 GNDA.n1870 GNDA.n1869 185
R1789 GNDA.n1868 GNDA.n1867 185
R1790 GNDA.n1866 GNDA.n1810 185
R1791 GNDA.n1864 GNDA.n1863 185
R1792 GNDA.n1862 GNDA.n1811 185
R1793 GNDA.n1861 GNDA.n1860 185
R1794 GNDA.n1858 GNDA.n1812 185
R1795 GNDA.n1874 GNDA.n1807 185
R1796 GNDA.n1805 GNDA.n450 185
R1797 GNDA.n1905 GNDA.n1904 185
R1798 GNDA.n1902 GNDA.n448 185
R1799 GNDA.n1901 GNDA.n452 185
R1800 GNDA.n1899 GNDA.n1898 185
R1801 GNDA.n1890 GNDA.n453 185
R1802 GNDA.n1889 GNDA.n1888 185
R1803 GNDA.n1886 GNDA.n1885 185
R1804 GNDA.n739 GNDA.n703 185
R1805 GNDA.n754 GNDA.n753 185
R1806 GNDA.n752 GNDA.n704 185
R1807 GNDA.n751 GNDA.n750 185
R1808 GNDA.n749 GNDA.n748 185
R1809 GNDA.n747 GNDA.n746 185
R1810 GNDA.n745 GNDA.n744 185
R1811 GNDA.n743 GNDA.n742 185
R1812 GNDA.n741 GNDA.n740 185
R1813 GNDA.n722 GNDA.n721 185
R1814 GNDA.n724 GNDA.n723 185
R1815 GNDA.n726 GNDA.n725 185
R1816 GNDA.n728 GNDA.n727 185
R1817 GNDA.n730 GNDA.n729 185
R1818 GNDA.n732 GNDA.n731 185
R1819 GNDA.n734 GNDA.n733 185
R1820 GNDA.n736 GNDA.n735 185
R1821 GNDA.n738 GNDA.n737 185
R1822 GNDA.n696 GNDA.n655 185
R1823 GNDA.n706 GNDA.n705 185
R1824 GNDA.n708 GNDA.n707 185
R1825 GNDA.n710 GNDA.n709 185
R1826 GNDA.n712 GNDA.n711 185
R1827 GNDA.n714 GNDA.n713 185
R1828 GNDA.n716 GNDA.n715 185
R1829 GNDA.n718 GNDA.n717 185
R1830 GNDA.n720 GNDA.n719 185
R1831 GNDA.n695 GNDA.n656 185
R1832 GNDA.n689 GNDA.n688 185
R1833 GNDA.n676 GNDA.n675 185
R1834 GNDA.n682 GNDA.n681 185
R1835 GNDA.n677 GNDA.n671 185
R1836 GNDA.n758 GNDA.n757 185
R1837 GNDA.n670 GNDA.n668 185
R1838 GNDA.n764 GNDA.n763 185
R1839 GNDA.n766 GNDA.n765 185
R1840 GNDA.n1967 GNDA.n402 183.948
R1841 GNDA.n351 GNDA.n344 183.948
R1842 GNDA.n2138 GNDA.n2094 182.4
R1843 GNDA.n2420 GNDA.n2419 182.4
R1844 GNDA.t245 GNDA.n2130 181.226
R1845 GNDA.t216 GNDA.n134 181.226
R1846 GNDA.n1967 GNDA.n1966 180.013
R1847 GNDA.n1048 GNDA.n351 180.013
R1848 GNDA.n2371 GNDA.n2370 178.119
R1849 GNDA.n1148 GNDA.n1109 175.546
R1850 GNDA.n1144 GNDA.n1143 175.546
R1851 GNDA.n1140 GNDA.n1139 175.546
R1852 GNDA.n1136 GNDA.n1135 175.546
R1853 GNDA.n1770 GNDA.n642 175.546
R1854 GNDA.n1787 GNDA.n194 175.546
R1855 GNDA.n1787 GNDA.n531 175.546
R1856 GNDA.n1780 GNDA.n531 175.546
R1857 GNDA.n1780 GNDA.n538 175.546
R1858 GNDA.n612 GNDA.n538 175.546
R1859 GNDA.n626 GNDA.n612 175.546
R1860 GNDA.n626 GNDA.n610 175.546
R1861 GNDA.n631 GNDA.n610 175.546
R1862 GNDA.n631 GNDA.n540 175.546
R1863 GNDA.n1776 GNDA.n540 175.546
R1864 GNDA.n1776 GNDA.n541 175.546
R1865 GNDA.n202 GNDA.n201 175.546
R1866 GNDA.n2354 GNDA.n201 175.546
R1867 GNDA.n2352 GNDA.n2351 175.546
R1868 GNDA.n2348 GNDA.n2347 175.546
R1869 GNDA.n2344 GNDA.n2343 175.546
R1870 GNDA.n2362 GNDA.n195 175.546
R1871 GNDA.n1113 GNDA.n1112 175.546
R1872 GNDA.n1117 GNDA.n1116 175.546
R1873 GNDA.n1121 GNDA.n1120 175.546
R1874 GNDA.n1125 GNDA.n1124 175.546
R1875 GNDA.n1129 GNDA.n1128 175.546
R1876 GNDA.n1747 GNDA.n1746 175.546
R1877 GNDA.n1751 GNDA.n1750 175.546
R1878 GNDA.n1755 GNDA.n1754 175.546
R1879 GNDA.n1759 GNDA.n1758 175.546
R1880 GNDA.n1763 GNDA.n1762 175.546
R1881 GNDA.n1329 GNDA.n1328 175.546
R1882 GNDA.n1245 GNDA.n1244 175.546
R1883 GNDA.n1251 GNDA.n1250 175.546
R1884 GNDA.n1258 GNDA.n1257 175.546
R1885 GNDA.n1266 GNDA.n1265 175.546
R1886 GNDA.n1515 GNDA.n1462 175.546
R1887 GNDA.n1519 GNDA.n1517 175.546
R1888 GNDA.n1525 GNDA.n1458 175.546
R1889 GNDA.n1529 GNDA.n1527 175.546
R1890 GNDA.n1539 GNDA.n1449 175.546
R1891 GNDA.n1504 GNDA.n1503 175.546
R1892 GNDA.n1500 GNDA.n1499 175.546
R1893 GNDA.n1496 GNDA.n1495 175.546
R1894 GNDA.n1492 GNDA.n1491 175.546
R1895 GNDA.n1488 GNDA.n1153 175.546
R1896 GNDA.n366 GNDA.n357 175.546
R1897 GNDA.n359 GNDA.n358 175.546
R1898 GNDA.n361 GNDA.n360 175.546
R1899 GNDA.n363 GNDA.n362 175.546
R1900 GNDA.n365 GNDA.n364 175.546
R1901 GNDA.n1964 GNDA.n401 175.546
R1902 GNDA.n1964 GNDA.n404 175.546
R1903 GNDA.n1960 GNDA.n404 175.546
R1904 GNDA.n1960 GNDA.n1957 175.546
R1905 GNDA.n1957 GNDA.n339 175.546
R1906 GNDA.n2036 GNDA.n339 175.546
R1907 GNDA.n2036 GNDA.n340 175.546
R1908 GNDA.n2032 GNDA.n340 175.546
R1909 GNDA.n2032 GNDA.n343 175.546
R1910 GNDA.n2028 GNDA.n343 175.546
R1911 GNDA.n2028 GNDA.n345 175.546
R1912 GNDA.n936 GNDA.n935 175.546
R1913 GNDA.n852 GNDA.n851 175.546
R1914 GNDA.n858 GNDA.n857 175.546
R1915 GNDA.n865 GNDA.n864 175.546
R1916 GNDA.n873 GNDA.n872 175.546
R1917 GNDA.n1970 GNDA.n1969 175.546
R1918 GNDA.n1970 GNDA.n397 175.546
R1919 GNDA.n1976 GNDA.n397 175.546
R1920 GNDA.n1976 GNDA.n392 175.546
R1921 GNDA.n1982 GNDA.n392 175.546
R1922 GNDA.n1984 GNDA.n1982 175.546
R1923 GNDA.n1985 GNDA.n1984 175.546
R1924 GNDA.n1985 GNDA.n388 175.546
R1925 GNDA.n1991 GNDA.n388 175.546
R1926 GNDA.n1991 GNDA.n383 175.546
R1927 GNDA.n1997 GNDA.n383 175.546
R1928 GNDA.n1513 GNDA.n1512 175.546
R1929 GNDA.n1461 GNDA.n1460 175.546
R1930 GNDA.n1523 GNDA.n1522 175.546
R1931 GNDA.n1531 GNDA.n1456 175.546
R1932 GNDA.n1537 GNDA.n1451 175.546
R1933 GNDA.n1466 GNDA.n1465 175.546
R1934 GNDA.n1470 GNDA.n1469 175.546
R1935 GNDA.n1474 GNDA.n1473 175.546
R1936 GNDA.n1478 GNDA.n1477 175.546
R1937 GNDA.n1482 GNDA.n1481 175.546
R1938 GNDA.n1431 GNDA.n1216 175.546
R1939 GNDA.n1428 GNDA.n1427 175.546
R1940 GNDA.n1421 GNDA.n1420 175.546
R1941 GNDA.n1414 GNDA.n1413 175.546
R1942 GNDA.n1441 GNDA.n1440 175.546
R1943 GNDA.n1731 GNDA.n1176 175.546
R1944 GNDA.n1731 GNDA.n1182 175.546
R1945 GNDA.n1727 GNDA.n1726 175.546
R1946 GNDA.n1723 GNDA.n1722 175.546
R1947 GNDA.n1719 GNDA.n1718 175.546
R1948 GNDA.n1715 GNDA.n1181 175.546
R1949 GNDA.n2325 GNDA.n2324 175.546
R1950 GNDA.n2327 GNDA.n2326 175.546
R1951 GNDA.n2329 GNDA.n2328 175.546
R1952 GNDA.n2331 GNDA.n2330 175.546
R1953 GNDA.n2340 GNDA.n2332 175.546
R1954 GNDA.n239 GNDA.n238 175.546
R1955 GNDA.n235 GNDA.n234 175.546
R1956 GNDA.n231 GNDA.n230 175.546
R1957 GNDA.n227 GNDA.n207 175.546
R1958 GNDA.n2319 GNDA.n2318 175.546
R1959 GNDA.n2282 GNDA.n270 175.546
R1960 GNDA.n2278 GNDA.n270 175.546
R1961 GNDA.n2278 GNDA.n272 175.546
R1962 GNDA.n304 GNDA.n272 175.546
R1963 GNDA.n2193 GNDA.n304 175.546
R1964 GNDA.n2197 GNDA.n2193 175.546
R1965 GNDA.n2197 GNDA.n298 175.546
R1966 GNDA.n2209 GNDA.n298 175.546
R1967 GNDA.n2209 GNDA.n297 175.546
R1968 GNDA.n2214 GNDA.n297 175.546
R1969 GNDA.n2214 GNDA.n191 175.546
R1970 GNDA.n2310 GNDA.n245 175.546
R1971 GNDA.n2306 GNDA.n245 175.546
R1972 GNDA.n2306 GNDA.n249 175.546
R1973 GNDA.n2302 GNDA.n249 175.546
R1974 GNDA.n2302 GNDA.n253 175.546
R1975 GNDA.n2296 GNDA.n253 175.546
R1976 GNDA.n2296 GNDA.n2295 175.546
R1977 GNDA.n2295 GNDA.n257 175.546
R1978 GNDA.n2291 GNDA.n257 175.546
R1979 GNDA.n2291 GNDA.n261 175.546
R1980 GNDA.n264 GNDA.n261 175.546
R1981 GNDA.n1972 GNDA.n399 175.546
R1982 GNDA.n1973 GNDA.n1972 175.546
R1983 GNDA.n1973 GNDA.n395 175.546
R1984 GNDA.n1979 GNDA.n395 175.546
R1985 GNDA.n1980 GNDA.n1979 175.546
R1986 GNDA.n1980 GNDA.n390 175.546
R1987 GNDA.n1987 GNDA.n390 175.546
R1988 GNDA.n1988 GNDA.n1987 175.546
R1989 GNDA.n1988 GNDA.n386 175.546
R1990 GNDA.n1994 GNDA.n386 175.546
R1991 GNDA.n1995 GNDA.n1994 175.546
R1992 GNDA.n1929 GNDA.n414 175.546
R1993 GNDA.n1933 GNDA.n414 175.546
R1994 GNDA.n1933 GNDA.n412 175.546
R1995 GNDA.n1937 GNDA.n412 175.546
R1996 GNDA.n1937 GNDA.n410 175.546
R1997 GNDA.n1941 GNDA.n410 175.546
R1998 GNDA.n1941 GNDA.n408 175.546
R1999 GNDA.n1946 GNDA.n408 175.546
R2000 GNDA.n1946 GNDA.n406 175.546
R2001 GNDA.n1950 GNDA.n406 175.546
R2002 GNDA.n1951 GNDA.n1950 175.546
R2003 GNDA.n801 GNDA.n781 175.546
R2004 GNDA.n1021 GNDA.n1020 175.546
R2005 GNDA.n947 GNDA.n946 175.546
R2006 GNDA.n952 GNDA.n951 175.546
R2007 GNDA.n960 GNDA.n959 175.546
R2008 GNDA.n1925 GNDA.n417 175.546
R2009 GNDA.n785 GNDA.n784 175.546
R2010 GNDA.n789 GNDA.n788 175.546
R2011 GNDA.n793 GNDA.n792 175.546
R2012 GNDA.n795 GNDA.n422 175.546
R2013 GNDA.n798 GNDA.n422 175.546
R2014 GNDA.n1192 GNDA.n1183 175.546
R2015 GNDA.n1185 GNDA.n1184 175.546
R2016 GNDA.n1187 GNDA.n1186 175.546
R2017 GNDA.n1189 GNDA.n1188 175.546
R2018 GNDA.n1191 GNDA.n1190 175.546
R2019 GNDA.n1641 GNDA.n1640 175.546
R2020 GNDA.n1637 GNDA.n1636 175.546
R2021 GNDA.n1633 GNDA.n1632 175.546
R2022 GNDA.n1629 GNDA.n1628 175.546
R2023 GNDA.n1625 GNDA.n1170 175.546
R2024 GNDA.n1682 GNDA.n1559 175.546
R2025 GNDA.n1686 GNDA.n1684 175.546
R2026 GNDA.n1697 GNDA.n1554 175.546
R2027 GNDA.n1701 GNDA.n1699 175.546
R2028 GNDA.n1709 GNDA.n1548 175.546
R2029 GNDA.n1649 GNDA.n1648 175.546
R2030 GNDA.n1653 GNDA.n1652 175.546
R2031 GNDA.n1657 GNDA.n1656 175.546
R2032 GNDA.n1661 GNDA.n1660 175.546
R2033 GNDA.n1663 GNDA.n429 175.546
R2034 GNDA.n1666 GNDA.n429 175.546
R2035 GNDA.n246 GNDA.n224 175.546
R2036 GNDA.n247 GNDA.n246 175.546
R2037 GNDA.n250 GNDA.n247 175.546
R2038 GNDA.n251 GNDA.n250 175.546
R2039 GNDA.n2299 GNDA.n251 175.546
R2040 GNDA.n2299 GNDA.n2298 175.546
R2041 GNDA.n2298 GNDA.n254 175.546
R2042 GNDA.n258 GNDA.n254 175.546
R2043 GNDA.n259 GNDA.n258 175.546
R2044 GNDA.n263 GNDA.n259 175.546
R2045 GNDA.n2287 GNDA.n263 175.546
R2046 GNDA.n476 GNDA.n475 175.546
R2047 GNDA.n472 GNDA.n471 175.546
R2048 GNDA.n468 GNDA.n467 175.546
R2049 GNDA.n464 GNDA.n463 175.546
R2050 GNDA.n460 GNDA.n223 175.546
R2051 GNDA.n1883 GNDA.n505 175.546
R2052 GNDA.n1883 GNDA.n456 175.546
R2053 GNDA.n1892 GNDA.n456 175.546
R2054 GNDA.n1892 GNDA.n455 175.546
R2055 GNDA.n1896 GNDA.n455 175.546
R2056 GNDA.n1896 GNDA.n446 175.546
R2057 GNDA.n1907 GNDA.n446 175.546
R2058 GNDA.n1907 GNDA.n447 175.546
R2059 GNDA.n509 GNDA.n447 175.546
R2060 GNDA.n1879 GNDA.n509 175.546
R2061 GNDA.n1879 GNDA.n1804 175.546
R2062 GNDA.n484 GNDA.n483 175.546
R2063 GNDA.n488 GNDA.n487 175.546
R2064 GNDA.n492 GNDA.n491 175.546
R2065 GNDA.n496 GNDA.n495 175.546
R2066 GNDA.n500 GNDA.n499 175.546
R2067 GNDA.n2019 GNDA.n350 175.546
R2068 GNDA.n2015 GNDA.n356 175.546
R2069 GNDA.n2013 GNDA.n2012 175.546
R2070 GNDA.n2009 GNDA.n2008 175.546
R2071 GNDA.n2005 GNDA.n2004 175.546
R2072 GNDA.n1050 GNDA.n349 175.546
R2073 GNDA.n1050 GNDA.n1047 175.546
R2074 GNDA.n1054 GNDA.n1047 175.546
R2075 GNDA.n1054 GNDA.n1045 175.546
R2076 GNDA.n1058 GNDA.n1045 175.546
R2077 GNDA.n1058 GNDA.n1043 175.546
R2078 GNDA.n1062 GNDA.n1043 175.546
R2079 GNDA.n1062 GNDA.n1041 175.546
R2080 GNDA.n1067 GNDA.n1041 175.546
R2081 GNDA.n1067 GNDA.n1039 175.546
R2082 GNDA.n1071 GNDA.n1039 175.546
R2083 GNDA.n768 GNDA.n662 175.546
R2084 GNDA.n761 GNDA.n760 175.546
R2085 GNDA.n679 GNDA.n678 175.546
R2086 GNDA.n685 GNDA.n684 175.546
R2087 GNDA.n1034 GNDA.n657 175.546
R2088 GNDA.n1076 GNDA.n1075 175.546
R2089 GNDA.n1080 GNDA.n1079 175.546
R2090 GNDA.n1084 GNDA.n1083 175.546
R2091 GNDA.n1088 GNDA.n1087 175.546
R2092 GNDA.n1092 GNDA.n1091 175.546
R2093 GNDA.n1534 GNDA.n1533 173.881
R2094 GNDA.n1198 GNDA.t219 172.876
R2095 GNDA.n1732 GNDA.t219 172.615
R2096 GNDA.n1533 GNDA.n1448 171.624
R2097 GNDA.n1798 GNDA.n520 169.601
R2098 GNDA.n1798 GNDA.n518 169.601
R2099 GNDA.n638 GNDA.n637 163.333
R2100 GNDA.n1270 GNDA.n1269 163.333
R2101 GNDA.n877 GNDA.n876 163.333
R2102 GNDA.n1347 GNDA.n1337 163.333
R2103 GNDA.n2218 GNDA.n2217 163.333
R2104 GNDA.n964 GNDA.n963 163.333
R2105 GNDA.n1706 GNDA.n1550 163.333
R2106 GNDA.n1875 GNDA.n1874 163.333
R2107 GNDA.n696 GNDA.n695 163.333
R2108 GNDA.n441 GNDA.t273 160.725
R2109 GNDA.n439 GNDA.t270 160.725
R2110 GNDA.n519 GNDA.t250 160.725
R2111 GNDA.n517 GNDA.t302 160.725
R2112 GNDA.n643 GNDA.t256 160.725
R2113 GNDA.n526 GNDA.t276 160.725
R2114 GNDA.n313 GNDA.t333 156.919
R2115 GNDA.n2443 GNDA.n34 156.8
R2116 GNDA.n2134 GNDA.n2102 153.601
R2117 GNDA.n142 GNDA.n99 153.601
R2118 GNDA.n2099 GNDA.t246 152.994
R2119 GNDA.n2095 GNDA.t238 152.994
R2120 GNDA.n84 GNDA.t241 152.994
R2121 GNDA.n136 GNDA.t217 152.994
R2122 GNDA.n2451 GNDA.n2450 150.4
R2123 GNDA.n2139 GNDA.n2138 150.4
R2124 GNDA.n2420 GNDA.n86 150.4
R2125 GNDA.n587 GNDA.n586 150
R2126 GNDA.n583 GNDA.n582 150
R2127 GNDA.n579 GNDA.n578 150
R2128 GNDA.n575 GNDA.n574 150
R2129 GNDA.n571 GNDA.n570 150
R2130 GNDA.n567 GNDA.n566 150
R2131 GNDA.n563 GNDA.n562 150
R2132 GNDA.n559 GNDA.n558 150
R2133 GNDA.n1784 GNDA.n1783 150
R2134 GNDA.n619 GNDA.n615 150
R2135 GNDA.n623 GNDA.n621 150
R2136 GNDA.n635 GNDA.n608 150
R2137 GNDA.n606 GNDA.n557 150
R2138 GNDA.n602 GNDA.n601 150
R2139 GNDA.n598 GNDA.n597 150
R2140 GNDA.n594 GNDA.n593 150
R2141 GNDA.n1302 GNDA.n1301 150
R2142 GNDA.n1298 GNDA.n1297 150
R2143 GNDA.n1294 GNDA.n1293 150
R2144 GNDA.n1290 GNDA.n1289 150
R2145 GNDA.n1286 GNDA.n1285 150
R2146 GNDA.n1282 GNDA.n1281 150
R2147 GNDA.n1278 GNDA.n1277 150
R2148 GNDA.n1274 GNDA.n1273 150
R2149 GNDA.n1325 GNDA.n1223 150
R2150 GNDA.n1247 GNDA.n1224 150
R2151 GNDA.n1255 GNDA.n1254 150
R2152 GNDA.n1262 GNDA.n1261 150
R2153 GNDA.n1310 GNDA.n1309 150
R2154 GNDA.n1314 GNDA.n1313 150
R2155 GNDA.n1318 GNDA.n1317 150
R2156 GNDA.n1322 GNDA.n1321 150
R2157 GNDA.n909 GNDA.n908 150
R2158 GNDA.n905 GNDA.n904 150
R2159 GNDA.n901 GNDA.n900 150
R2160 GNDA.n897 GNDA.n896 150
R2161 GNDA.n893 GNDA.n892 150
R2162 GNDA.n889 GNDA.n888 150
R2163 GNDA.n885 GNDA.n884 150
R2164 GNDA.n881 GNDA.n880 150
R2165 GNDA.n932 GNDA.n828 150
R2166 GNDA.n854 GNDA.n829 150
R2167 GNDA.n862 GNDA.n861 150
R2168 GNDA.n869 GNDA.n868 150
R2169 GNDA.n917 GNDA.n916 150
R2170 GNDA.n921 GNDA.n920 150
R2171 GNDA.n925 GNDA.n924 150
R2172 GNDA.n929 GNDA.n928 150
R2173 GNDA.n1387 GNDA.n1386 150
R2174 GNDA.n1383 GNDA.n1382 150
R2175 GNDA.n1379 GNDA.n1378 150
R2176 GNDA.n1375 GNDA.n1374 150
R2177 GNDA.n1371 GNDA.n1370 150
R2178 GNDA.n1367 GNDA.n1366 150
R2179 GNDA.n1363 GNDA.n1362 150
R2180 GNDA.n1359 GNDA.n1358 150
R2181 GNDA.n1434 GNDA.n1356 150
R2182 GNDA.n1424 GNDA.n1423 150
R2183 GNDA.n1417 GNDA.n1416 150
R2184 GNDA.n1437 GNDA.n1336 150
R2185 GNDA.n1395 GNDA.n1394 150
R2186 GNDA.n1399 GNDA.n1398 150
R2187 GNDA.n1403 GNDA.n1402 150
R2188 GNDA.n1405 GNDA.n1355 150
R2189 GNDA.n2250 GNDA.n2249 150
R2190 GNDA.n2246 GNDA.n2245 150
R2191 GNDA.n2242 GNDA.n2241 150
R2192 GNDA.n2238 GNDA.n2237 150
R2193 GNDA.n2234 GNDA.n2233 150
R2194 GNDA.n2230 GNDA.n2229 150
R2195 GNDA.n2226 GNDA.n2225 150
R2196 GNDA.n2222 GNDA.n2221 150
R2197 GNDA.n2275 GNDA.n275 150
R2198 GNDA.n301 GNDA.n276 150
R2199 GNDA.n2201 GNDA.n2200 150
R2200 GNDA.n2206 GNDA.n2205 150
R2201 GNDA.n2258 GNDA.n2257 150
R2202 GNDA.n2262 GNDA.n2261 150
R2203 GNDA.n2266 GNDA.n2265 150
R2204 GNDA.n2272 GNDA.n293 150
R2205 GNDA.n996 GNDA.n995 150
R2206 GNDA.n992 GNDA.n991 150
R2207 GNDA.n988 GNDA.n987 150
R2208 GNDA.n984 GNDA.n983 150
R2209 GNDA.n980 GNDA.n979 150
R2210 GNDA.n976 GNDA.n975 150
R2211 GNDA.n972 GNDA.n971 150
R2212 GNDA.n968 GNDA.n967 150
R2213 GNDA.n1025 GNDA.n1024 150
R2214 GNDA.n1017 GNDA.n807 150
R2215 GNDA.n949 GNDA.n808 150
R2216 GNDA.n956 GNDA.n955 150
R2217 GNDA.n1014 GNDA.n824 150
R2218 GNDA.n1010 GNDA.n1009 150
R2219 GNDA.n1006 GNDA.n1005 150
R2220 GNDA.n1002 GNDA.n1001 150
R2221 GNDA.n1606 GNDA.n1604 150
R2222 GNDA.n1602 GNDA.n1567 150
R2223 GNDA.n1598 GNDA.n1596 150
R2224 GNDA.n1594 GNDA.n1569 150
R2225 GNDA.n1590 GNDA.n1588 150
R2226 GNDA.n1586 GNDA.n1571 150
R2227 GNDA.n1582 GNDA.n1581 150
R2228 GNDA.n1579 GNDA.n1575 150
R2229 GNDA.n1679 GNDA.n1677 150
R2230 GNDA.n1690 GNDA.n1556 150
R2231 GNDA.n1694 GNDA.n1692 150
R2232 GNDA.n1704 GNDA.n1551 150
R2233 GNDA.n1614 GNDA.n1612 150
R2234 GNDA.n1618 GNDA.n1563 150
R2235 GNDA.n1622 GNDA.n1620 150
R2236 GNDA.n1675 GNDA.n1561 150
R2237 GNDA.n1844 GNDA.n1842 150
R2238 GNDA.n1848 GNDA.n1815 150
R2239 GNDA.n1852 GNDA.n1850 150
R2240 GNDA.n1856 GNDA.n1813 150
R2241 GNDA.n1860 GNDA.n1858 150
R2242 GNDA.n1864 GNDA.n1811 150
R2243 GNDA.n1867 GNDA.n1866 150
R2244 GNDA.n1871 GNDA.n1870 150
R2245 GNDA.n1888 GNDA.n1886 150
R2246 GNDA.n1899 GNDA.n453 150
R2247 GNDA.n1902 GNDA.n1901 150
R2248 GNDA.n1904 GNDA.n450 150
R2249 GNDA.n1836 GNDA.n1835 150
R2250 GNDA.n1833 GNDA.n1820 150
R2251 GNDA.n1829 GNDA.n1827 150
R2252 GNDA.n1825 GNDA.n1822 150
R2253 GNDA.n735 GNDA.n734 150
R2254 GNDA.n731 GNDA.n730 150
R2255 GNDA.n727 GNDA.n726 150
R2256 GNDA.n723 GNDA.n722 150
R2257 GNDA.n719 GNDA.n718 150
R2258 GNDA.n715 GNDA.n714 150
R2259 GNDA.n711 GNDA.n710 150
R2260 GNDA.n707 GNDA.n706 150
R2261 GNDA.n765 GNDA.n764 150
R2262 GNDA.n757 GNDA.n670 150
R2263 GNDA.n681 GNDA.n671 150
R2264 GNDA.n689 GNDA.n675 150
R2265 GNDA.n754 GNDA.n704 150
R2266 GNDA.n750 GNDA.n749 150
R2267 GNDA.n746 GNDA.n745 150
R2268 GNDA.n742 GNDA.n741 150
R2269 GNDA.n2129 GNDA.t292 147.511
R2270 GNDA.n133 GNDA.t307 147.511
R2271 GNDA.n316 GNDA.n314 139.638
R2272 GNDA.n332 GNDA.n331 139.077
R2273 GNDA.n330 GNDA.n329 139.077
R2274 GNDA.n328 GNDA.n327 139.077
R2275 GNDA.n326 GNDA.n325 139.077
R2276 GNDA.n324 GNDA.n323 139.077
R2277 GNDA.n322 GNDA.n321 139.077
R2278 GNDA.n320 GNDA.n319 139.077
R2279 GNDA.n318 GNDA.n317 139.077
R2280 GNDA.n316 GNDA.n315 139.077
R2281 GNDA.t116 GNDA.t280 135.386
R2282 GNDA.t22 GNDA.t56 135.386
R2283 GNDA.t228 GNDA.t128 135.386
R2284 GNDA.t286 GNDA.t352 135.386
R2285 GNDA.t15 GNDA.t92 135.386
R2286 GNDA.t41 GNDA.t265 135.386
R2287 GNDA.n2107 GNDA.n2069 134.867
R2288 GNDA.n2424 GNDA.n81 134.867
R2289 GNDA.n2436 GNDA.n2435 134.4
R2290 GNDA.n2429 GNDA.n74 134.4
R2291 GNDA.n2428 GNDA.n78 134.4
R2292 GNDA.n2125 GNDA.n2124 134.4
R2293 GNDA.n2123 GNDA.n72 134.4
R2294 GNDA.n1769 GNDA.n640 132.721
R2295 GNDA.n1766 GNDA.n1102 132.721
R2296 GNDA.n502 GNDA.n436 132.721
R2297 GNDA.n1095 GNDA.n653 132.721
R2298 GNDA.n49 GNDA.n42 128
R2299 GNDA.n2363 GNDA.n2362 124.832
R2300 GNDA.n1542 GNDA.n1541 124.832
R2301 GNDA.n379 GNDA.n374 124.832
R2302 GNDA.n1998 GNDA.n1997 124.832
R2303 GNDA.n1535 GNDA.n1217 124.832
R2304 GNDA.n1544 GNDA.n1181 124.832
R2305 GNDA.n2365 GNDA.n190 124.832
R2306 GNDA.n2283 GNDA.n264 124.832
R2307 GNDA.n1995 GNDA.n380 124.832
R2308 GNDA.n1203 GNDA.n1200 124.832
R2309 GNDA.n2287 GNDA.n266 124.832
R2310 GNDA.n2001 GNDA.n2000 124.832
R2311 GNDA.n1920 GNDA.n440 118.4
R2312 GNDA.n443 GNDA.n442 118.4
R2313 GNDA.n1795 GNDA.n520 118.4
R2314 GNDA.n524 GNDA.n518 118.4
R2315 GNDA.n1794 GNDA.n527 118.4
R2316 GNDA.n645 GNDA.n644 118.4
R2317 GNDA.n2044 GNDA.t70 115.105
R2318 GNDA.n2042 GNDA.t74 114.635
R2319 GNDA.n2047 GNDA.t34 114.635
R2320 GNDA.n2048 GNDA.t347 114.448
R2321 GNDA.n46 GNDA.t243 113.974
R2322 GNDA.n47 GNDA.t223 113.974
R2323 GNDA.n48 GNDA.t293 113.974
R2324 GNDA.n43 GNDA.t308 113.974
R2325 GNDA.n44 GNDA.t290 113.974
R2326 GNDA.n45 GNDA.t284 113.974
R2327 GNDA.n77 GNDA.t296 113.974
R2328 GNDA.n73 GNDA.t287 113.974
R2329 GNDA.n2122 GNDA.t229 113.974
R2330 GNDA.n2121 GNDA.t299 113.974
R2331 GNDA.n69 GNDA.n67 108.8
R2332 GNDA.n65 GNDA.n62 108.8
R2333 GNDA.n2316 GNDA.t219 47.6748
R2334 GNDA.n105 GNDA.n104 99.0842
R2335 GNDA.n107 GNDA.n106 99.0842
R2336 GNDA.n109 GNDA.n108 99.0842
R2337 GNDA.n111 GNDA.n110 99.0842
R2338 GNDA.n113 GNDA.n112 99.0842
R2339 GNDA.n115 GNDA.n114 99.0842
R2340 GNDA.n117 GNDA.n116 99.0842
R2341 GNDA.n119 GNDA.n118 99.0842
R2342 GNDA.n121 GNDA.n120 99.0842
R2343 GNDA.n123 GNDA.n122 99.0842
R2344 GNDA.n125 GNDA.n124 99.0842
R2345 GNDA.n2213 GNDA.n2212 96.988
R2346 GNDA.n1789 GNDA.n1788 96.988
R2347 GNDA.n2115 GNDA.n2112 95.101
R2348 GNDA.n131 GNDA.n130 95.101
R2349 GNDA.n102 GNDA.t226 94.8842
R2350 GNDA.n33 GNDA.t263 94.8842
R2351 GNDA.n1803 GNDA.t272 94.8327
R2352 GNDA.t301 GNDA.n2280 94.8327
R2353 GNDA.n2114 GNDA.n2113 94.601
R2354 GNDA.n129 GNDA.n128 94.601
R2355 GNDA.t54 GNDA.t237 92.7208
R2356 GNDA.t342 GNDA.t152 92.7208
R2357 GNDA.t55 GNDA.t150 92.7208
R2358 GNDA.t53 GNDA.t320 92.7208
R2359 GNDA.t108 GNDA.t49 92.7208
R2360 GNDA.t49 GNDA.t68 92.7208
R2361 GNDA.t283 GNDA.t48 92.7208
R2362 GNDA.t35 GNDA.t283 92.7208
R2363 GNDA.t84 GNDA.t40 92.7208
R2364 GNDA.t9 GNDA.t51 92.7208
R2365 GNDA.t130 GNDA.t46 92.7208
R2366 GNDA.t5 GNDA.t240 92.7208
R2367 GNDA.n1931 GNDA.n1930 88.5317
R2368 GNDA.n1932 GNDA.n1931 88.5317
R2369 GNDA.n1932 GNDA.n411 88.5317
R2370 GNDA.n1938 GNDA.n411 88.5317
R2371 GNDA.n1939 GNDA.n1938 88.5317
R2372 GNDA.n1940 GNDA.n407 88.5317
R2373 GNDA.n1947 GNDA.n407 88.5317
R2374 GNDA.n1948 GNDA.n1947 88.5317
R2375 GNDA.n1949 GNDA.n1948 88.5317
R2376 GNDA.n1949 GNDA.n402 88.5317
R2377 GNDA.n1966 GNDA.n1965 88.5317
R2378 GNDA.n1965 GNDA.n403 88.5317
R2379 GNDA.n1959 GNDA.n403 88.5317
R2380 GNDA.n1959 GNDA.n1958 88.5317
R2381 GNDA.n1958 GNDA.n337 88.5317
R2382 GNDA.n2037 GNDA.n338 88.5317
R2383 GNDA.n2031 GNDA.n338 88.5317
R2384 GNDA.n2031 GNDA.n2030 88.5317
R2385 GNDA.n2030 GNDA.n2029 88.5317
R2386 GNDA.n2029 GNDA.n344 88.5317
R2387 GNDA.n1051 GNDA.n1048 88.5317
R2388 GNDA.n1052 GNDA.n1051 88.5317
R2389 GNDA.n1053 GNDA.n1052 88.5317
R2390 GNDA.n1053 GNDA.n1044 88.5317
R2391 GNDA.n1059 GNDA.n1044 88.5317
R2392 GNDA.n1061 GNDA.n1060 88.5317
R2393 GNDA.n1061 GNDA.n1040 88.5317
R2394 GNDA.n1068 GNDA.n1040 88.5317
R2395 GNDA.n1069 GNDA.n1068 88.5317
R2396 GNDA.n1070 GNDA.n1069 88.5317
R2397 GNDA.t319 GNDA.t304 88.5063
R2398 GNDA.t47 GNDA.t258 88.5063
R2399 GNDA.t162 GNDA.t61 86.2116
R2400 GNDA.t332 GNDA.t355 86.2116
R2401 GNDA.n2381 GNDA.n2380 85.2845
R2402 GNDA.n181 GNDA.n180 85.2845
R2403 GNDA.n2039 GNDA.n335 84.306
R2404 GNDA.n521 GNDA.n269 82.9787
R2405 GNDA.n2191 GNDA.n306 82.9787
R2406 GNDA.n2366 GNDA.n189 81.9011
R2407 GNDA.n2309 GNDA.t219 80.9821
R2408 GNDA.n1968 GNDA.n1967 80.9821
R2409 GNDA.t233 GNDA.t54 80.0771
R2410 GNDA.t63 GNDA.t319 80.0771
R2411 GNDA.t31 GNDA.t47 80.0771
R2412 GNDA.t252 GNDA.t5 80.0771
R2413 GNDA.n2195 GNDA.n2194 78.6681
R2414 GNDA.n2182 GNDA.n310 78.6358
R2415 GNDA.n2389 GNDA.n174 78.6358
R2416 GNDA.t199 GNDA.n2211 77.5905
R2417 GNDA.n1533 GNDA.t219 76.3879
R2418 GNDA.n1149 GNDA.n1148 76.3222
R2419 GNDA.n1144 GNDA.n1107 76.3222
R2420 GNDA.n1140 GNDA.n1106 76.3222
R2421 GNDA.n1136 GNDA.n1105 76.3222
R2422 GNDA.n1104 GNDA.n642 76.3222
R2423 GNDA.n2360 GNDA.n2359 76.3222
R2424 GNDA.n2354 GNDA.n197 76.3222
R2425 GNDA.n2351 GNDA.n198 76.3222
R2426 GNDA.n2347 GNDA.n199 76.3222
R2427 GNDA.n2343 GNDA.n200 76.3222
R2428 GNDA.n1112 GNDA.n208 76.3222
R2429 GNDA.n1116 GNDA.n209 76.3222
R2430 GNDA.n1120 GNDA.n210 76.3222
R2431 GNDA.n1124 GNDA.n211 76.3222
R2432 GNDA.n1128 GNDA.n212 76.3222
R2433 GNDA.n1131 GNDA.n213 76.3222
R2434 GNDA.n1746 GNDA.n1097 76.3222
R2435 GNDA.n1750 GNDA.n1098 76.3222
R2436 GNDA.n1754 GNDA.n1099 76.3222
R2437 GNDA.n1758 GNDA.n1100 76.3222
R2438 GNDA.n1762 GNDA.n1101 76.3222
R2439 GNDA.n1219 GNDA.n1210 76.3222
R2440 GNDA.n1328 GNDA.n1209 76.3222
R2441 GNDA.n1245 GNDA.n1208 76.3222
R2442 GNDA.n1251 GNDA.n1207 76.3222
R2443 GNDA.n1257 GNDA.n1206 76.3222
R2444 GNDA.n1266 GNDA.n1205 76.3222
R2445 GNDA.n1509 GNDA.n1508 76.3222
R2446 GNDA.n1516 GNDA.n1515 76.3222
R2447 GNDA.n1519 GNDA.n1518 76.3222
R2448 GNDA.n1526 GNDA.n1525 76.3222
R2449 GNDA.n1529 GNDA.n1528 76.3222
R2450 GNDA.n1540 GNDA.n1539 76.3222
R2451 GNDA.n1504 GNDA.n1154 76.3222
R2452 GNDA.n1500 GNDA.n1155 76.3222
R2453 GNDA.n1496 GNDA.n1156 76.3222
R2454 GNDA.n1492 GNDA.n1157 76.3222
R2455 GNDA.n1488 GNDA.n1158 76.3222
R2456 GNDA.n1742 GNDA.n1741 76.3222
R2457 GNDA.n367 GNDA.n366 76.3222
R2458 GNDA.n368 GNDA.n358 76.3222
R2459 GNDA.n369 GNDA.n360 76.3222
R2460 GNDA.n370 GNDA.n362 76.3222
R2461 GNDA.n371 GNDA.n364 76.3222
R2462 GNDA.n374 GNDA.n373 76.3222
R2463 GNDA.n775 GNDA.n382 76.3222
R2464 GNDA.n935 GNDA.n774 76.3222
R2465 GNDA.n852 GNDA.n773 76.3222
R2466 GNDA.n858 GNDA.n772 76.3222
R2467 GNDA.n864 GNDA.n771 76.3222
R2468 GNDA.n873 GNDA.n770 76.3222
R2469 GNDA.n1512 GNDA.n1452 76.3222
R2470 GNDA.n1460 GNDA.n1453 76.3222
R2471 GNDA.n1522 GNDA.n1454 76.3222
R2472 GNDA.n1456 GNDA.n1455 76.3222
R2473 GNDA.n1532 GNDA.n1451 76.3222
R2474 GNDA.n1536 GNDA.n1535 76.3222
R2475 GNDA.n1465 GNDA.n1159 76.3222
R2476 GNDA.n1469 GNDA.n1160 76.3222
R2477 GNDA.n1473 GNDA.n1161 76.3222
R2478 GNDA.n1477 GNDA.n1162 76.3222
R2479 GNDA.n1481 GNDA.n1163 76.3222
R2480 GNDA.n1485 GNDA.n1164 76.3222
R2481 GNDA.n1546 GNDA.n1545 76.3222
R2482 GNDA.n1431 GNDA.n1215 76.3222
R2483 GNDA.n1427 GNDA.n1214 76.3222
R2484 GNDA.n1420 GNDA.n1213 76.3222
R2485 GNDA.n1413 GNDA.n1212 76.3222
R2486 GNDA.n1441 GNDA.n1211 76.3222
R2487 GNDA.n1734 GNDA.n1733 76.3222
R2488 GNDA.n1182 GNDA.n1177 76.3222
R2489 GNDA.n1726 GNDA.n1178 76.3222
R2490 GNDA.n1722 GNDA.n1179 76.3222
R2491 GNDA.n1718 GNDA.n1180 76.3222
R2492 GNDA.n2333 GNDA.n2324 76.3222
R2493 GNDA.n2334 GNDA.n2326 76.3222
R2494 GNDA.n2335 GNDA.n2328 76.3222
R2495 GNDA.n2336 GNDA.n2330 76.3222
R2496 GNDA.n2337 GNDA.n2332 76.3222
R2497 GNDA.n2339 GNDA.n190 76.3222
R2498 GNDA.n239 GNDA.n214 76.3222
R2499 GNDA.n235 GNDA.n215 76.3222
R2500 GNDA.n231 GNDA.n216 76.3222
R2501 GNDA.n227 GNDA.n217 76.3222
R2502 GNDA.n2318 GNDA.n2317 76.3222
R2503 GNDA.n2322 GNDA.n205 76.3222
R2504 GNDA.n1031 GNDA.n1030 76.3222
R2505 GNDA.n801 GNDA.n780 76.3222
R2506 GNDA.n1020 GNDA.n779 76.3222
R2507 GNDA.n947 GNDA.n778 76.3222
R2508 GNDA.n951 GNDA.n777 76.3222
R2509 GNDA.n960 GNDA.n776 76.3222
R2510 GNDA.n1924 GNDA.n415 76.3222
R2511 GNDA.n418 GNDA.n417 76.3222
R2512 GNDA.n785 GNDA.n419 76.3222
R2513 GNDA.n789 GNDA.n420 76.3222
R2514 GNDA.n793 GNDA.n421 76.3222
R2515 GNDA.n1193 GNDA.n1171 76.3222
R2516 GNDA.n1194 GNDA.n1183 76.3222
R2517 GNDA.n1195 GNDA.n1185 76.3222
R2518 GNDA.n1196 GNDA.n1187 76.3222
R2519 GNDA.n1197 GNDA.n1189 76.3222
R2520 GNDA.n1199 GNDA.n1191 76.3222
R2521 GNDA.n1641 GNDA.n1165 76.3222
R2522 GNDA.n1637 GNDA.n1166 76.3222
R2523 GNDA.n1633 GNDA.n1167 76.3222
R2524 GNDA.n1629 GNDA.n1168 76.3222
R2525 GNDA.n1625 GNDA.n1169 76.3222
R2526 GNDA.n1739 GNDA.n1738 76.3222
R2527 GNDA.n1670 GNDA.n1669 76.3222
R2528 GNDA.n1683 GNDA.n1682 76.3222
R2529 GNDA.n1686 GNDA.n1685 76.3222
R2530 GNDA.n1698 GNDA.n1697 76.3222
R2531 GNDA.n1701 GNDA.n1700 76.3222
R2532 GNDA.n1710 GNDA.n1709 76.3222
R2533 GNDA.n1645 GNDA.n424 76.3222
R2534 GNDA.n1649 GNDA.n425 76.3222
R2535 GNDA.n1653 GNDA.n426 76.3222
R2536 GNDA.n1657 GNDA.n427 76.3222
R2537 GNDA.n1661 GNDA.n428 76.3222
R2538 GNDA.n1648 GNDA.n424 76.3222
R2539 GNDA.n1652 GNDA.n425 76.3222
R2540 GNDA.n1656 GNDA.n426 76.3222
R2541 GNDA.n1660 GNDA.n427 76.3222
R2542 GNDA.n1663 GNDA.n428 76.3222
R2543 GNDA.n1925 GNDA.n1924 76.3222
R2544 GNDA.n784 GNDA.n418 76.3222
R2545 GNDA.n788 GNDA.n419 76.3222
R2546 GNDA.n792 GNDA.n420 76.3222
R2547 GNDA.n795 GNDA.n421 76.3222
R2548 GNDA.n476 GNDA.n218 76.3222
R2549 GNDA.n472 GNDA.n219 76.3222
R2550 GNDA.n468 GNDA.n220 76.3222
R2551 GNDA.n464 GNDA.n221 76.3222
R2552 GNDA.n460 GNDA.n222 76.3222
R2553 GNDA.n2315 GNDA.n2314 76.3222
R2554 GNDA.n480 GNDA.n431 76.3222
R2555 GNDA.n484 GNDA.n432 76.3222
R2556 GNDA.n488 GNDA.n433 76.3222
R2557 GNDA.n492 GNDA.n434 76.3222
R2558 GNDA.n496 GNDA.n435 76.3222
R2559 GNDA.n500 GNDA.n436 76.3222
R2560 GNDA.n483 GNDA.n431 76.3222
R2561 GNDA.n487 GNDA.n432 76.3222
R2562 GNDA.n491 GNDA.n433 76.3222
R2563 GNDA.n495 GNDA.n434 76.3222
R2564 GNDA.n499 GNDA.n435 76.3222
R2565 GNDA.n1200 GNDA.n1199 76.3222
R2566 GNDA.n1197 GNDA.n1190 76.3222
R2567 GNDA.n1196 GNDA.n1188 76.3222
R2568 GNDA.n1195 GNDA.n1186 76.3222
R2569 GNDA.n1194 GNDA.n1184 76.3222
R2570 GNDA.n1193 GNDA.n1192 76.3222
R2571 GNDA.n1733 GNDA.n1176 76.3222
R2572 GNDA.n1727 GNDA.n1177 76.3222
R2573 GNDA.n1723 GNDA.n1178 76.3222
R2574 GNDA.n1719 GNDA.n1179 76.3222
R2575 GNDA.n1715 GNDA.n1180 76.3222
R2576 GNDA.n1739 GNDA.n1170 76.3222
R2577 GNDA.n1628 GNDA.n1169 76.3222
R2578 GNDA.n1632 GNDA.n1168 76.3222
R2579 GNDA.n1636 GNDA.n1167 76.3222
R2580 GNDA.n1640 GNDA.n1166 76.3222
R2581 GNDA.n1644 GNDA.n1165 76.3222
R2582 GNDA.n1482 GNDA.n1164 76.3222
R2583 GNDA.n1478 GNDA.n1163 76.3222
R2584 GNDA.n1474 GNDA.n1162 76.3222
R2585 GNDA.n1470 GNDA.n1161 76.3222
R2586 GNDA.n1466 GNDA.n1160 76.3222
R2587 GNDA.n1175 GNDA.n1159 76.3222
R2588 GNDA.n1741 GNDA.n1153 76.3222
R2589 GNDA.n1491 GNDA.n1158 76.3222
R2590 GNDA.n1495 GNDA.n1157 76.3222
R2591 GNDA.n1499 GNDA.n1156 76.3222
R2592 GNDA.n1503 GNDA.n1155 76.3222
R2593 GNDA.n1507 GNDA.n1154 76.3222
R2594 GNDA.n1031 GNDA.n781 76.3222
R2595 GNDA.n1021 GNDA.n780 76.3222
R2596 GNDA.n946 GNDA.n779 76.3222
R2597 GNDA.n952 GNDA.n778 76.3222
R2598 GNDA.n959 GNDA.n777 76.3222
R2599 GNDA.n941 GNDA.n776 76.3222
R2600 GNDA.n936 GNDA.n775 76.3222
R2601 GNDA.n851 GNDA.n774 76.3222
R2602 GNDA.n857 GNDA.n773 76.3222
R2603 GNDA.n865 GNDA.n772 76.3222
R2604 GNDA.n872 GNDA.n771 76.3222
R2605 GNDA.n846 GNDA.n770 76.3222
R2606 GNDA.n2315 GNDA.n223 76.3222
R2607 GNDA.n463 GNDA.n222 76.3222
R2608 GNDA.n467 GNDA.n221 76.3222
R2609 GNDA.n471 GNDA.n220 76.3222
R2610 GNDA.n475 GNDA.n219 76.3222
R2611 GNDA.n479 GNDA.n218 76.3222
R2612 GNDA.n2319 GNDA.n205 76.3222
R2613 GNDA.n2317 GNDA.n207 76.3222
R2614 GNDA.n230 GNDA.n217 76.3222
R2615 GNDA.n234 GNDA.n216 76.3222
R2616 GNDA.n238 GNDA.n215 76.3222
R2617 GNDA.n244 GNDA.n214 76.3222
R2618 GNDA.n1129 GNDA.n213 76.3222
R2619 GNDA.n1125 GNDA.n212 76.3222
R2620 GNDA.n1121 GNDA.n211 76.3222
R2621 GNDA.n1117 GNDA.n210 76.3222
R2622 GNDA.n1113 GNDA.n209 76.3222
R2623 GNDA.n208 GNDA.n203 76.3222
R2624 GNDA.n1669 GNDA.n1559 76.3222
R2625 GNDA.n1684 GNDA.n1683 76.3222
R2626 GNDA.n1685 GNDA.n1554 76.3222
R2627 GNDA.n1699 GNDA.n1698 76.3222
R2628 GNDA.n1700 GNDA.n1548 76.3222
R2629 GNDA.n1711 GNDA.n1710 76.3222
R2630 GNDA.n1546 GNDA.n1216 76.3222
R2631 GNDA.n1428 GNDA.n1215 76.3222
R2632 GNDA.n1421 GNDA.n1214 76.3222
R2633 GNDA.n1414 GNDA.n1213 76.3222
R2634 GNDA.n1440 GNDA.n1212 76.3222
R2635 GNDA.n1444 GNDA.n1211 76.3222
R2636 GNDA.n1329 GNDA.n1210 76.3222
R2637 GNDA.n1244 GNDA.n1209 76.3222
R2638 GNDA.n1250 GNDA.n1208 76.3222
R2639 GNDA.n1258 GNDA.n1207 76.3222
R2640 GNDA.n1265 GNDA.n1206 76.3222
R2641 GNDA.n1205 GNDA.n1150 76.3222
R2642 GNDA.n1770 GNDA.n1769 76.3222
R2643 GNDA.n1135 GNDA.n1104 76.3222
R2644 GNDA.n1139 GNDA.n1105 76.3222
R2645 GNDA.n1143 GNDA.n1106 76.3222
R2646 GNDA.n1109 GNDA.n1107 76.3222
R2647 GNDA.n1149 GNDA.n1108 76.3222
R2648 GNDA.n1763 GNDA.n1102 76.3222
R2649 GNDA.n1759 GNDA.n1101 76.3222
R2650 GNDA.n1755 GNDA.n1100 76.3222
R2651 GNDA.n1751 GNDA.n1099 76.3222
R2652 GNDA.n1747 GNDA.n1098 76.3222
R2653 GNDA.n1743 GNDA.n1097 76.3222
R2654 GNDA.n2023 GNDA.n2022 76.3222
R2655 GNDA.n2020 GNDA.n2019 76.3222
R2656 GNDA.n2015 GNDA.n355 76.3222
R2657 GNDA.n2012 GNDA.n354 76.3222
R2658 GNDA.n2008 GNDA.n353 76.3222
R2659 GNDA.n2004 GNDA.n352 76.3222
R2660 GNDA.n769 GNDA.n376 76.3222
R2661 GNDA.n662 GNDA.n661 76.3222
R2662 GNDA.n760 GNDA.n660 76.3222
R2663 GNDA.n679 GNDA.n659 76.3222
R2664 GNDA.n685 GNDA.n658 76.3222
R2665 GNDA.n1034 GNDA.n1033 76.3222
R2666 GNDA.n1072 GNDA.n648 76.3222
R2667 GNDA.n1076 GNDA.n649 76.3222
R2668 GNDA.n1080 GNDA.n650 76.3222
R2669 GNDA.n1084 GNDA.n651 76.3222
R2670 GNDA.n1088 GNDA.n652 76.3222
R2671 GNDA.n1092 GNDA.n653 76.3222
R2672 GNDA.n769 GNDA.n768 76.3222
R2673 GNDA.n761 GNDA.n661 76.3222
R2674 GNDA.n678 GNDA.n660 76.3222
R2675 GNDA.n684 GNDA.n659 76.3222
R2676 GNDA.n658 GNDA.n657 76.3222
R2677 GNDA.n1033 GNDA.n654 76.3222
R2678 GNDA.n1091 GNDA.n652 76.3222
R2679 GNDA.n1087 GNDA.n651 76.3222
R2680 GNDA.n1083 GNDA.n650 76.3222
R2681 GNDA.n1079 GNDA.n649 76.3222
R2682 GNDA.n1075 GNDA.n648 76.3222
R2683 GNDA.n373 GNDA.n365 76.3222
R2684 GNDA.n371 GNDA.n363 76.3222
R2685 GNDA.n370 GNDA.n361 76.3222
R2686 GNDA.n369 GNDA.n359 76.3222
R2687 GNDA.n368 GNDA.n357 76.3222
R2688 GNDA.n367 GNDA.n347 76.3222
R2689 GNDA.n2022 GNDA.n350 76.3222
R2690 GNDA.n2020 GNDA.n356 76.3222
R2691 GNDA.n2013 GNDA.n355 76.3222
R2692 GNDA.n2009 GNDA.n354 76.3222
R2693 GNDA.n2005 GNDA.n353 76.3222
R2694 GNDA.n2001 GNDA.n352 76.3222
R2695 GNDA.n1537 GNDA.n1536 76.3222
R2696 GNDA.n1532 GNDA.n1531 76.3222
R2697 GNDA.n1523 GNDA.n1455 76.3222
R2698 GNDA.n1461 GNDA.n1454 76.3222
R2699 GNDA.n1513 GNDA.n1453 76.3222
R2700 GNDA.n1486 GNDA.n1452 76.3222
R2701 GNDA.n1508 GNDA.n1462 76.3222
R2702 GNDA.n1517 GNDA.n1516 76.3222
R2703 GNDA.n1518 GNDA.n1458 76.3222
R2704 GNDA.n1527 GNDA.n1526 76.3222
R2705 GNDA.n1528 GNDA.n1449 76.3222
R2706 GNDA.n1541 GNDA.n1540 76.3222
R2707 GNDA.n2340 GNDA.n2339 76.3222
R2708 GNDA.n2337 GNDA.n2331 76.3222
R2709 GNDA.n2336 GNDA.n2329 76.3222
R2710 GNDA.n2335 GNDA.n2327 76.3222
R2711 GNDA.n2334 GNDA.n2325 76.3222
R2712 GNDA.n2333 GNDA.n2323 76.3222
R2713 GNDA.n2360 GNDA.n202 76.3222
R2714 GNDA.n2352 GNDA.n197 76.3222
R2715 GNDA.n2348 GNDA.n198 76.3222
R2716 GNDA.n2344 GNDA.n199 76.3222
R2717 GNDA.n200 GNDA.n195 76.3222
R2718 GNDA.t292 GNDA.t298 75.8626
R2719 GNDA.t18 GNDA.t329 75.8626
R2720 GNDA.t98 GNDA.t117 75.8626
R2721 GNDA.t331 GNDA.t310 75.8626
R2722 GNDA.t339 GNDA.t134 75.8626
R2723 GNDA.t307 GNDA.t295 75.8626
R2724 GNDA.n574 GNDA.n547 74.5978
R2725 GNDA.n571 GNDA.n547 74.5978
R2726 GNDA.n1289 GNDA.n1230 74.5978
R2727 GNDA.n1286 GNDA.n1230 74.5978
R2728 GNDA.n896 GNDA.n835 74.5978
R2729 GNDA.n893 GNDA.n835 74.5978
R2730 GNDA.n1374 GNDA.n1343 74.5978
R2731 GNDA.n1371 GNDA.n1343 74.5978
R2732 GNDA.n2237 GNDA.n282 74.5978
R2733 GNDA.n2234 GNDA.n282 74.5978
R2734 GNDA.n983 GNDA.n813 74.5978
R2735 GNDA.n980 GNDA.n813 74.5978
R2736 GNDA.n1589 GNDA.n1569 74.5978
R2737 GNDA.n1590 GNDA.n1589 74.5978
R2738 GNDA.n1857 GNDA.n1856 74.5978
R2739 GNDA.n1858 GNDA.n1857 74.5978
R2740 GNDA.n722 GNDA.n691 74.5978
R2741 GNDA.n719 GNDA.n691 74.5978
R2742 GNDA.t195 GNDA.n2279 73.2799
R2743 GNDA.n2091 GNDA.t67 72.3996
R2744 GNDA.n2148 GNDA.t4 72.3996
R2745 GNDA.t340 GNDA.n80 72.3996
R2746 GNDA.t341 GNDA.n2409 72.3996
R2747 GNDA.t139 GNDA.n2128 71.648
R2748 GNDA.n155 GNDA.n93 70.0642
R2749 GNDA.n1784 GNDA.n535 69.3109
R2750 GNDA.n593 GNDA.n535 69.3109
R2751 GNDA.n1323 GNDA.n1223 69.3109
R2752 GNDA.n1323 GNDA.n1322 69.3109
R2753 GNDA.n930 GNDA.n828 69.3109
R2754 GNDA.n930 GNDA.n929 69.3109
R2755 GNDA.n1435 GNDA.n1434 69.3109
R2756 GNDA.n1435 GNDA.n1355 69.3109
R2757 GNDA.n2273 GNDA.n275 69.3109
R2758 GNDA.n2273 GNDA.n2272 69.3109
R2759 GNDA.n1025 GNDA.n803 69.3109
R2760 GNDA.n1001 GNDA.n803 69.3109
R2761 GNDA.n1677 GNDA.n1676 69.3109
R2762 GNDA.n1676 GNDA.n1675 69.3109
R2763 GNDA.n1886 GNDA.n458 69.3109
R2764 GNDA.n1822 GNDA.n458 69.3109
R2765 GNDA.n765 GNDA.n666 69.3109
R2766 GNDA.n741 GNDA.n666 69.3109
R2767 GNDA.n1881 GNDA.t189 66.8141
R2768 GNDA.t211 GNDA.n305 66.8141
R2769 GNDA.t278 GNDA.n607 65.8183
R2770 GNDA.t278 GNDA.n555 65.8183
R2771 GNDA.t278 GNDA.n554 65.8183
R2772 GNDA.t278 GNDA.n553 65.8183
R2773 GNDA.t278 GNDA.n546 65.8183
R2774 GNDA.t278 GNDA.n551 65.8183
R2775 GNDA.t278 GNDA.n545 65.8183
R2776 GNDA.t278 GNDA.n552 65.8183
R2777 GNDA.t278 GNDA.n544 65.8183
R2778 GNDA.t278 GNDA.n550 65.8183
R2779 GNDA.t278 GNDA.n549 65.8183
R2780 GNDA.t278 GNDA.n548 65.8183
R2781 GNDA.n636 GNDA.t278 65.8183
R2782 GNDA.n622 GNDA.t278 65.8183
R2783 GNDA.n620 GNDA.t278 65.8183
R2784 GNDA.t278 GNDA.n536 65.8183
R2785 GNDA.t277 GNDA.n1240 65.8183
R2786 GNDA.t277 GNDA.n1239 65.8183
R2787 GNDA.t277 GNDA.n1238 65.8183
R2788 GNDA.t277 GNDA.n1237 65.8183
R2789 GNDA.t277 GNDA.n1228 65.8183
R2790 GNDA.t277 GNDA.n1235 65.8183
R2791 GNDA.t277 GNDA.n1225 65.8183
R2792 GNDA.t277 GNDA.n1236 65.8183
R2793 GNDA.t277 GNDA.n1234 65.8183
R2794 GNDA.t277 GNDA.n1233 65.8183
R2795 GNDA.t277 GNDA.n1232 65.8183
R2796 GNDA.t277 GNDA.n1231 65.8183
R2797 GNDA.t277 GNDA.n1229 65.8183
R2798 GNDA.t277 GNDA.n1227 65.8183
R2799 GNDA.t277 GNDA.n1226 65.8183
R2800 GNDA.n1324 GNDA.t277 65.8183
R2801 GNDA.t235 GNDA.n845 65.8183
R2802 GNDA.t235 GNDA.n844 65.8183
R2803 GNDA.t235 GNDA.n843 65.8183
R2804 GNDA.t235 GNDA.n842 65.8183
R2805 GNDA.t235 GNDA.n833 65.8183
R2806 GNDA.t235 GNDA.n840 65.8183
R2807 GNDA.t235 GNDA.n830 65.8183
R2808 GNDA.t235 GNDA.n841 65.8183
R2809 GNDA.t235 GNDA.n839 65.8183
R2810 GNDA.t235 GNDA.n838 65.8183
R2811 GNDA.t235 GNDA.n837 65.8183
R2812 GNDA.t235 GNDA.n836 65.8183
R2813 GNDA.t235 GNDA.n834 65.8183
R2814 GNDA.t235 GNDA.n832 65.8183
R2815 GNDA.t235 GNDA.n831 65.8183
R2816 GNDA.n931 GNDA.t235 65.8183
R2817 GNDA.t247 GNDA.n1354 65.8183
R2818 GNDA.t247 GNDA.n1353 65.8183
R2819 GNDA.t247 GNDA.n1352 65.8183
R2820 GNDA.t247 GNDA.n1351 65.8183
R2821 GNDA.t247 GNDA.n1342 65.8183
R2822 GNDA.t247 GNDA.n1349 65.8183
R2823 GNDA.t247 GNDA.n1339 65.8183
R2824 GNDA.t247 GNDA.n1350 65.8183
R2825 GNDA.t247 GNDA.n1348 65.8183
R2826 GNDA.t247 GNDA.n1346 65.8183
R2827 GNDA.t247 GNDA.n1345 65.8183
R2828 GNDA.t247 GNDA.n1344 65.8183
R2829 GNDA.n1436 GNDA.t247 65.8183
R2830 GNDA.t247 GNDA.n1341 65.8183
R2831 GNDA.t247 GNDA.n1340 65.8183
R2832 GNDA.t247 GNDA.n1338 65.8183
R2833 GNDA.t230 GNDA.n292 65.8183
R2834 GNDA.t230 GNDA.n291 65.8183
R2835 GNDA.t230 GNDA.n290 65.8183
R2836 GNDA.t230 GNDA.n289 65.8183
R2837 GNDA.t230 GNDA.n280 65.8183
R2838 GNDA.t230 GNDA.n287 65.8183
R2839 GNDA.t230 GNDA.n277 65.8183
R2840 GNDA.t230 GNDA.n288 65.8183
R2841 GNDA.t230 GNDA.n286 65.8183
R2842 GNDA.t230 GNDA.n285 65.8183
R2843 GNDA.t230 GNDA.n284 65.8183
R2844 GNDA.t230 GNDA.n283 65.8183
R2845 GNDA.t230 GNDA.n281 65.8183
R2846 GNDA.t230 GNDA.n279 65.8183
R2847 GNDA.t230 GNDA.n278 65.8183
R2848 GNDA.n2274 GNDA.t230 65.8183
R2849 GNDA.t231 GNDA.n1015 65.8183
R2850 GNDA.t231 GNDA.n822 65.8183
R2851 GNDA.t231 GNDA.n821 65.8183
R2852 GNDA.t231 GNDA.n820 65.8183
R2853 GNDA.t231 GNDA.n811 65.8183
R2854 GNDA.t231 GNDA.n818 65.8183
R2855 GNDA.t231 GNDA.n809 65.8183
R2856 GNDA.t231 GNDA.n819 65.8183
R2857 GNDA.t231 GNDA.n817 65.8183
R2858 GNDA.t231 GNDA.n816 65.8183
R2859 GNDA.t231 GNDA.n815 65.8183
R2860 GNDA.t231 GNDA.n814 65.8183
R2861 GNDA.t231 GNDA.n812 65.8183
R2862 GNDA.t231 GNDA.n810 65.8183
R2863 GNDA.n1016 GNDA.t231 65.8183
R2864 GNDA.t231 GNDA.n804 65.8183
R2865 GNDA.n1611 GNDA.t267 65.8183
R2866 GNDA.n1613 GNDA.t267 65.8183
R2867 GNDA.n1619 GNDA.t267 65.8183
R2868 GNDA.n1621 GNDA.t267 65.8183
R2869 GNDA.n1595 GNDA.t267 65.8183
R2870 GNDA.n1597 GNDA.t267 65.8183
R2871 GNDA.n1603 GNDA.t267 65.8183
R2872 GNDA.n1605 GNDA.t267 65.8183
R2873 GNDA.n1574 GNDA.t267 65.8183
R2874 GNDA.n1580 GNDA.t267 65.8183
R2875 GNDA.n1573 GNDA.t267 65.8183
R2876 GNDA.n1587 GNDA.t267 65.8183
R2877 GNDA.n1705 GNDA.t267 65.8183
R2878 GNDA.n1693 GNDA.t267 65.8183
R2879 GNDA.n1691 GNDA.t267 65.8183
R2880 GNDA.n1678 GNDA.t267 65.8183
R2881 GNDA.n1819 GNDA.t220 65.8183
R2882 GNDA.n1834 GNDA.t220 65.8183
R2883 GNDA.n1828 GNDA.t220 65.8183
R2884 GNDA.n1826 GNDA.t220 65.8183
R2885 GNDA.n1851 GNDA.t220 65.8183
R2886 GNDA.n1849 GNDA.t220 65.8183
R2887 GNDA.n1843 GNDA.t220 65.8183
R2888 GNDA.n1841 GNDA.t220 65.8183
R2889 GNDA.n1872 GNDA.t220 65.8183
R2890 GNDA.n1809 GNDA.t220 65.8183
R2891 GNDA.n1865 GNDA.t220 65.8183
R2892 GNDA.n1859 GNDA.t220 65.8183
R2893 GNDA.n1873 GNDA.t220 65.8183
R2894 GNDA.n1903 GNDA.t220 65.8183
R2895 GNDA.n1900 GNDA.t220 65.8183
R2896 GNDA.n1887 GNDA.t220 65.8183
R2897 GNDA.t218 GNDA.n755 65.8183
R2898 GNDA.t218 GNDA.n702 65.8183
R2899 GNDA.t218 GNDA.n701 65.8183
R2900 GNDA.t218 GNDA.n700 65.8183
R2901 GNDA.t218 GNDA.n674 65.8183
R2902 GNDA.t218 GNDA.n698 65.8183
R2903 GNDA.t218 GNDA.n672 65.8183
R2904 GNDA.t218 GNDA.n699 65.8183
R2905 GNDA.t218 GNDA.n697 65.8183
R2906 GNDA.t218 GNDA.n694 65.8183
R2907 GNDA.t218 GNDA.n693 65.8183
R2908 GNDA.t218 GNDA.n692 65.8183
R2909 GNDA.t218 GNDA.n690 65.8183
R2910 GNDA.t218 GNDA.n673 65.8183
R2911 GNDA.n756 GNDA.t218 65.8183
R2912 GNDA.t218 GNDA.n667 65.8183
R2913 GNDA.n2433 GNDA.n2432 64.0005
R2914 GNDA.n2432 GNDA.n51 64.0005
R2915 GNDA.t159 GNDA.t342 63.2189
R2916 GNDA.t6 GNDA.t53 63.2189
R2917 GNDA.t165 GNDA.t84 63.2189
R2918 GNDA.t316 GNDA.t130 63.2189
R2919 GNDA.n2210 GNDA.t213 62.5036
R2920 GNDA.t203 GNDA.n629 62.5036
R2921 GNDA.t62 GNDA.n1894 61.4259
R2922 GNDA.t173 GNDA.n507 61.4259
R2923 GNDA.t179 GNDA.t77 59.2706
R2924 GNDA.t91 GNDA.t175 59.2706
R2925 GNDA.t228 GNDA.t108 59.0043
R2926 GNDA.t286 GNDA.t35 59.0043
R2927 GNDA.n2367 GNDA.n2366 58.193
R2928 GNDA.t278 GNDA.n535 57.8461
R2929 GNDA.t277 GNDA.n1323 57.8461
R2930 GNDA.t235 GNDA.n930 57.8461
R2931 GNDA.t247 GNDA.n1435 57.8461
R2932 GNDA.t230 GNDA.n2273 57.8461
R2933 GNDA.t231 GNDA.n803 57.8461
R2934 GNDA.n1676 GNDA.t267 57.8461
R2935 GNDA.n458 GNDA.t220 57.8461
R2936 GNDA.t218 GNDA.n666 57.8461
R2937 GNDA.n2087 GNDA.n2086 57.6005
R2938 GNDA.n2413 GNDA.n90 57.6005
R2939 GNDA.n2169 GNDA.n2054 57.1898
R2940 GNDA.n2407 GNDA.n161 57.1898
R2941 GNDA.n271 GNDA.n269 57.1154
R2942 GNDA.n1779 GNDA.t82 57.1154
R2943 GNDA.n628 GNDA.t96 57.1154
R2944 GNDA.n798 GNDA.n423 56.3995
R2945 GNDA.n1666 GNDA.n430 56.3995
R2946 GNDA.n1668 GNDA.n430 56.3995
R2947 GNDA.n782 GNDA.n423 56.3995
R2948 GNDA.n502 GNDA.n437 56.3995
R2949 GNDA.n1103 GNDA.n640 56.3995
R2950 GNDA.n1767 GNDA.n1766 56.3995
R2951 GNDA.n1096 GNDA.n1095 56.3995
R2952 GNDA.t197 GNDA.n2210 56.0377
R2953 GNDA.n2161 GNDA.t125 55.4026
R2954 GNDA.t30 GNDA.n2170 55.4026
R2955 GNDA.n2174 GNDA.t33 55.4026
R2956 GNDA.n2176 GNDA.t3 55.4026
R2957 GNDA.n2395 GNDA.t110 55.4026
R2958 GNDA.t69 GNDA.n2396 55.4026
R2959 GNDA.n2400 GNDA.t337 55.4026
R2960 GNDA.n2401 GNDA.t148 55.4026
R2961 GNDA.t278 GNDA.n547 55.2026
R2962 GNDA.t277 GNDA.n1230 55.2026
R2963 GNDA.t235 GNDA.n835 55.2026
R2964 GNDA.t247 GNDA.n1343 55.2026
R2965 GNDA.t230 GNDA.n282 55.2026
R2966 GNDA.t231 GNDA.n813 55.2026
R2967 GNDA.n1589 GNDA.t267 55.2026
R2968 GNDA.n1857 GNDA.t220 55.2026
R2969 GNDA.t218 GNDA.n691 55.2026
R2970 GNDA.n2131 GNDA.t133 54.7898
R2971 GNDA.n145 GNDA.t58 54.7898
R2972 GNDA.n2448 GNDA.n34 54.4005
R2973 GNDA.n589 GNDA.n552 53.3664
R2974 GNDA.n586 GNDA.n545 53.3664
R2975 GNDA.n582 GNDA.n551 53.3664
R2976 GNDA.n578 GNDA.n546 53.3664
R2977 GNDA.n567 GNDA.n548 53.3664
R2978 GNDA.n563 GNDA.n549 53.3664
R2979 GNDA.n559 GNDA.n550 53.3664
R2980 GNDA.n638 GNDA.n544 53.3664
R2981 GNDA.n1783 GNDA.n536 53.3664
R2982 GNDA.n620 GNDA.n619 53.3664
R2983 GNDA.n623 GNDA.n622 53.3664
R2984 GNDA.n636 GNDA.n635 53.3664
R2985 GNDA.n607 GNDA.n606 53.3664
R2986 GNDA.n557 GNDA.n555 53.3664
R2987 GNDA.n601 GNDA.n554 53.3664
R2988 GNDA.n597 GNDA.n553 53.3664
R2989 GNDA.n607 GNDA.n556 53.3664
R2990 GNDA.n602 GNDA.n555 53.3664
R2991 GNDA.n598 GNDA.n554 53.3664
R2992 GNDA.n594 GNDA.n553 53.3664
R2993 GNDA.n575 GNDA.n546 53.3664
R2994 GNDA.n579 GNDA.n551 53.3664
R2995 GNDA.n583 GNDA.n545 53.3664
R2996 GNDA.n587 GNDA.n552 53.3664
R2997 GNDA.n558 GNDA.n544 53.3664
R2998 GNDA.n562 GNDA.n550 53.3664
R2999 GNDA.n566 GNDA.n549 53.3664
R3000 GNDA.n570 GNDA.n548 53.3664
R3001 GNDA.n637 GNDA.n636 53.3664
R3002 GNDA.n622 GNDA.n608 53.3664
R3003 GNDA.n621 GNDA.n620 53.3664
R3004 GNDA.n615 GNDA.n536 53.3664
R3005 GNDA.n1305 GNDA.n1236 53.3664
R3006 GNDA.n1301 GNDA.n1225 53.3664
R3007 GNDA.n1297 GNDA.n1235 53.3664
R3008 GNDA.n1293 GNDA.n1228 53.3664
R3009 GNDA.n1282 GNDA.n1231 53.3664
R3010 GNDA.n1278 GNDA.n1232 53.3664
R3011 GNDA.n1274 GNDA.n1233 53.3664
R3012 GNDA.n1270 GNDA.n1234 53.3664
R3013 GNDA.n1325 GNDA.n1324 53.3664
R3014 GNDA.n1247 GNDA.n1226 53.3664
R3015 GNDA.n1255 GNDA.n1227 53.3664
R3016 GNDA.n1262 GNDA.n1229 53.3664
R3017 GNDA.n1309 GNDA.n1240 53.3664
R3018 GNDA.n1310 GNDA.n1239 53.3664
R3019 GNDA.n1314 GNDA.n1238 53.3664
R3020 GNDA.n1318 GNDA.n1237 53.3664
R3021 GNDA.n1306 GNDA.n1240 53.3664
R3022 GNDA.n1313 GNDA.n1239 53.3664
R3023 GNDA.n1317 GNDA.n1238 53.3664
R3024 GNDA.n1321 GNDA.n1237 53.3664
R3025 GNDA.n1290 GNDA.n1228 53.3664
R3026 GNDA.n1294 GNDA.n1235 53.3664
R3027 GNDA.n1298 GNDA.n1225 53.3664
R3028 GNDA.n1302 GNDA.n1236 53.3664
R3029 GNDA.n1273 GNDA.n1234 53.3664
R3030 GNDA.n1277 GNDA.n1233 53.3664
R3031 GNDA.n1281 GNDA.n1232 53.3664
R3032 GNDA.n1285 GNDA.n1231 53.3664
R3033 GNDA.n1269 GNDA.n1229 53.3664
R3034 GNDA.n1261 GNDA.n1227 53.3664
R3035 GNDA.n1254 GNDA.n1226 53.3664
R3036 GNDA.n1324 GNDA.n1224 53.3664
R3037 GNDA.n912 GNDA.n841 53.3664
R3038 GNDA.n908 GNDA.n830 53.3664
R3039 GNDA.n904 GNDA.n840 53.3664
R3040 GNDA.n900 GNDA.n833 53.3664
R3041 GNDA.n889 GNDA.n836 53.3664
R3042 GNDA.n885 GNDA.n837 53.3664
R3043 GNDA.n881 GNDA.n838 53.3664
R3044 GNDA.n877 GNDA.n839 53.3664
R3045 GNDA.n932 GNDA.n931 53.3664
R3046 GNDA.n854 GNDA.n831 53.3664
R3047 GNDA.n862 GNDA.n832 53.3664
R3048 GNDA.n869 GNDA.n834 53.3664
R3049 GNDA.n916 GNDA.n845 53.3664
R3050 GNDA.n917 GNDA.n844 53.3664
R3051 GNDA.n921 GNDA.n843 53.3664
R3052 GNDA.n925 GNDA.n842 53.3664
R3053 GNDA.n913 GNDA.n845 53.3664
R3054 GNDA.n920 GNDA.n844 53.3664
R3055 GNDA.n924 GNDA.n843 53.3664
R3056 GNDA.n928 GNDA.n842 53.3664
R3057 GNDA.n897 GNDA.n833 53.3664
R3058 GNDA.n901 GNDA.n840 53.3664
R3059 GNDA.n905 GNDA.n830 53.3664
R3060 GNDA.n909 GNDA.n841 53.3664
R3061 GNDA.n880 GNDA.n839 53.3664
R3062 GNDA.n884 GNDA.n838 53.3664
R3063 GNDA.n888 GNDA.n837 53.3664
R3064 GNDA.n892 GNDA.n836 53.3664
R3065 GNDA.n876 GNDA.n834 53.3664
R3066 GNDA.n868 GNDA.n832 53.3664
R3067 GNDA.n861 GNDA.n831 53.3664
R3068 GNDA.n931 GNDA.n829 53.3664
R3069 GNDA.n1390 GNDA.n1350 53.3664
R3070 GNDA.n1386 GNDA.n1339 53.3664
R3071 GNDA.n1382 GNDA.n1349 53.3664
R3072 GNDA.n1378 GNDA.n1342 53.3664
R3073 GNDA.n1367 GNDA.n1344 53.3664
R3074 GNDA.n1363 GNDA.n1345 53.3664
R3075 GNDA.n1359 GNDA.n1346 53.3664
R3076 GNDA.n1348 GNDA.n1347 53.3664
R3077 GNDA.n1356 GNDA.n1338 53.3664
R3078 GNDA.n1424 GNDA.n1340 53.3664
R3079 GNDA.n1417 GNDA.n1341 53.3664
R3080 GNDA.n1437 GNDA.n1436 53.3664
R3081 GNDA.n1394 GNDA.n1354 53.3664
R3082 GNDA.n1395 GNDA.n1353 53.3664
R3083 GNDA.n1399 GNDA.n1352 53.3664
R3084 GNDA.n1403 GNDA.n1351 53.3664
R3085 GNDA.n1391 GNDA.n1354 53.3664
R3086 GNDA.n1398 GNDA.n1353 53.3664
R3087 GNDA.n1402 GNDA.n1352 53.3664
R3088 GNDA.n1405 GNDA.n1351 53.3664
R3089 GNDA.n1375 GNDA.n1342 53.3664
R3090 GNDA.n1379 GNDA.n1349 53.3664
R3091 GNDA.n1383 GNDA.n1339 53.3664
R3092 GNDA.n1387 GNDA.n1350 53.3664
R3093 GNDA.n1358 GNDA.n1348 53.3664
R3094 GNDA.n1362 GNDA.n1346 53.3664
R3095 GNDA.n1366 GNDA.n1345 53.3664
R3096 GNDA.n1370 GNDA.n1344 53.3664
R3097 GNDA.n1436 GNDA.n1337 53.3664
R3098 GNDA.n1341 GNDA.n1336 53.3664
R3099 GNDA.n1416 GNDA.n1340 53.3664
R3100 GNDA.n1423 GNDA.n1338 53.3664
R3101 GNDA.n2253 GNDA.n288 53.3664
R3102 GNDA.n2249 GNDA.n277 53.3664
R3103 GNDA.n2245 GNDA.n287 53.3664
R3104 GNDA.n2241 GNDA.n280 53.3664
R3105 GNDA.n2230 GNDA.n283 53.3664
R3106 GNDA.n2226 GNDA.n284 53.3664
R3107 GNDA.n2222 GNDA.n285 53.3664
R3108 GNDA.n2218 GNDA.n286 53.3664
R3109 GNDA.n2275 GNDA.n2274 53.3664
R3110 GNDA.n301 GNDA.n278 53.3664
R3111 GNDA.n2201 GNDA.n279 53.3664
R3112 GNDA.n2206 GNDA.n281 53.3664
R3113 GNDA.n2257 GNDA.n292 53.3664
R3114 GNDA.n2258 GNDA.n291 53.3664
R3115 GNDA.n2262 GNDA.n290 53.3664
R3116 GNDA.n2266 GNDA.n289 53.3664
R3117 GNDA.n2254 GNDA.n292 53.3664
R3118 GNDA.n2261 GNDA.n291 53.3664
R3119 GNDA.n2265 GNDA.n290 53.3664
R3120 GNDA.n293 GNDA.n289 53.3664
R3121 GNDA.n2238 GNDA.n280 53.3664
R3122 GNDA.n2242 GNDA.n287 53.3664
R3123 GNDA.n2246 GNDA.n277 53.3664
R3124 GNDA.n2250 GNDA.n288 53.3664
R3125 GNDA.n2221 GNDA.n286 53.3664
R3126 GNDA.n2225 GNDA.n285 53.3664
R3127 GNDA.n2229 GNDA.n284 53.3664
R3128 GNDA.n2233 GNDA.n283 53.3664
R3129 GNDA.n2217 GNDA.n281 53.3664
R3130 GNDA.n2205 GNDA.n279 53.3664
R3131 GNDA.n2200 GNDA.n278 53.3664
R3132 GNDA.n2274 GNDA.n276 53.3664
R3133 GNDA.n998 GNDA.n819 53.3664
R3134 GNDA.n995 GNDA.n809 53.3664
R3135 GNDA.n991 GNDA.n818 53.3664
R3136 GNDA.n987 GNDA.n811 53.3664
R3137 GNDA.n976 GNDA.n814 53.3664
R3138 GNDA.n972 GNDA.n815 53.3664
R3139 GNDA.n968 GNDA.n816 53.3664
R3140 GNDA.n964 GNDA.n817 53.3664
R3141 GNDA.n1024 GNDA.n804 53.3664
R3142 GNDA.n1017 GNDA.n1016 53.3664
R3143 GNDA.n949 GNDA.n810 53.3664
R3144 GNDA.n956 GNDA.n812 53.3664
R3145 GNDA.n1015 GNDA.n1014 53.3664
R3146 GNDA.n824 GNDA.n822 53.3664
R3147 GNDA.n1009 GNDA.n821 53.3664
R3148 GNDA.n1005 GNDA.n820 53.3664
R3149 GNDA.n1015 GNDA.n823 53.3664
R3150 GNDA.n1010 GNDA.n822 53.3664
R3151 GNDA.n1006 GNDA.n821 53.3664
R3152 GNDA.n1002 GNDA.n820 53.3664
R3153 GNDA.n984 GNDA.n811 53.3664
R3154 GNDA.n988 GNDA.n818 53.3664
R3155 GNDA.n992 GNDA.n809 53.3664
R3156 GNDA.n996 GNDA.n819 53.3664
R3157 GNDA.n967 GNDA.n817 53.3664
R3158 GNDA.n971 GNDA.n816 53.3664
R3159 GNDA.n975 GNDA.n815 53.3664
R3160 GNDA.n979 GNDA.n814 53.3664
R3161 GNDA.n963 GNDA.n812 53.3664
R3162 GNDA.n955 GNDA.n810 53.3664
R3163 GNDA.n1016 GNDA.n808 53.3664
R3164 GNDA.n807 GNDA.n804 53.3664
R3165 GNDA.n1605 GNDA.n1565 53.3664
R3166 GNDA.n1604 GNDA.n1603 53.3664
R3167 GNDA.n1597 GNDA.n1567 53.3664
R3168 GNDA.n1596 GNDA.n1595 53.3664
R3169 GNDA.n1587 GNDA.n1586 53.3664
R3170 GNDA.n1582 GNDA.n1573 53.3664
R3171 GNDA.n1580 GNDA.n1579 53.3664
R3172 GNDA.n1574 GNDA.n1550 53.3664
R3173 GNDA.n1679 GNDA.n1678 53.3664
R3174 GNDA.n1691 GNDA.n1690 53.3664
R3175 GNDA.n1694 GNDA.n1693 53.3664
R3176 GNDA.n1705 GNDA.n1704 53.3664
R3177 GNDA.n1612 GNDA.n1611 53.3664
R3178 GNDA.n1614 GNDA.n1613 53.3664
R3179 GNDA.n1619 GNDA.n1618 53.3664
R3180 GNDA.n1622 GNDA.n1621 53.3664
R3181 GNDA.n1611 GNDA.n1610 53.3664
R3182 GNDA.n1613 GNDA.n1563 53.3664
R3183 GNDA.n1620 GNDA.n1619 53.3664
R3184 GNDA.n1621 GNDA.n1561 53.3664
R3185 GNDA.n1595 GNDA.n1594 53.3664
R3186 GNDA.n1598 GNDA.n1597 53.3664
R3187 GNDA.n1603 GNDA.n1602 53.3664
R3188 GNDA.n1606 GNDA.n1605 53.3664
R3189 GNDA.n1575 GNDA.n1574 53.3664
R3190 GNDA.n1581 GNDA.n1580 53.3664
R3191 GNDA.n1573 GNDA.n1571 53.3664
R3192 GNDA.n1588 GNDA.n1587 53.3664
R3193 GNDA.n1706 GNDA.n1705 53.3664
R3194 GNDA.n1693 GNDA.n1551 53.3664
R3195 GNDA.n1692 GNDA.n1691 53.3664
R3196 GNDA.n1678 GNDA.n1556 53.3664
R3197 GNDA.n1841 GNDA.n1840 53.3664
R3198 GNDA.n1844 GNDA.n1843 53.3664
R3199 GNDA.n1849 GNDA.n1848 53.3664
R3200 GNDA.n1852 GNDA.n1851 53.3664
R3201 GNDA.n1859 GNDA.n1811 53.3664
R3202 GNDA.n1866 GNDA.n1865 53.3664
R3203 GNDA.n1870 GNDA.n1809 53.3664
R3204 GNDA.n1875 GNDA.n1872 53.3664
R3205 GNDA.n1888 GNDA.n1887 53.3664
R3206 GNDA.n1900 GNDA.n1899 53.3664
R3207 GNDA.n1903 GNDA.n1902 53.3664
R3208 GNDA.n1873 GNDA.n450 53.3664
R3209 GNDA.n1836 GNDA.n1819 53.3664
R3210 GNDA.n1835 GNDA.n1834 53.3664
R3211 GNDA.n1828 GNDA.n1820 53.3664
R3212 GNDA.n1827 GNDA.n1826 53.3664
R3213 GNDA.n1819 GNDA.n1817 53.3664
R3214 GNDA.n1834 GNDA.n1833 53.3664
R3215 GNDA.n1829 GNDA.n1828 53.3664
R3216 GNDA.n1826 GNDA.n1825 53.3664
R3217 GNDA.n1851 GNDA.n1813 53.3664
R3218 GNDA.n1850 GNDA.n1849 53.3664
R3219 GNDA.n1843 GNDA.n1815 53.3664
R3220 GNDA.n1842 GNDA.n1841 53.3664
R3221 GNDA.n1872 GNDA.n1871 53.3664
R3222 GNDA.n1867 GNDA.n1809 53.3664
R3223 GNDA.n1865 GNDA.n1864 53.3664
R3224 GNDA.n1860 GNDA.n1859 53.3664
R3225 GNDA.n1874 GNDA.n1873 53.3664
R3226 GNDA.n1904 GNDA.n1903 53.3664
R3227 GNDA.n1901 GNDA.n1900 53.3664
R3228 GNDA.n1887 GNDA.n453 53.3664
R3229 GNDA.n737 GNDA.n699 53.3664
R3230 GNDA.n734 GNDA.n672 53.3664
R3231 GNDA.n730 GNDA.n698 53.3664
R3232 GNDA.n726 GNDA.n674 53.3664
R3233 GNDA.n715 GNDA.n692 53.3664
R3234 GNDA.n711 GNDA.n693 53.3664
R3235 GNDA.n707 GNDA.n694 53.3664
R3236 GNDA.n697 GNDA.n696 53.3664
R3237 GNDA.n764 GNDA.n667 53.3664
R3238 GNDA.n757 GNDA.n756 53.3664
R3239 GNDA.n681 GNDA.n673 53.3664
R3240 GNDA.n690 GNDA.n689 53.3664
R3241 GNDA.n755 GNDA.n754 53.3664
R3242 GNDA.n704 GNDA.n702 53.3664
R3243 GNDA.n749 GNDA.n701 53.3664
R3244 GNDA.n745 GNDA.n700 53.3664
R3245 GNDA.n755 GNDA.n703 53.3664
R3246 GNDA.n750 GNDA.n702 53.3664
R3247 GNDA.n746 GNDA.n701 53.3664
R3248 GNDA.n742 GNDA.n700 53.3664
R3249 GNDA.n723 GNDA.n674 53.3664
R3250 GNDA.n727 GNDA.n698 53.3664
R3251 GNDA.n731 GNDA.n672 53.3664
R3252 GNDA.n735 GNDA.n699 53.3664
R3253 GNDA.n706 GNDA.n697 53.3664
R3254 GNDA.n710 GNDA.n694 53.3664
R3255 GNDA.n714 GNDA.n693 53.3664
R3256 GNDA.n718 GNDA.n692 53.3664
R3257 GNDA.n695 GNDA.n690 53.3664
R3258 GNDA.n675 GNDA.n673 53.3664
R3259 GNDA.n756 GNDA.n671 53.3664
R3260 GNDA.n670 GNDA.n667 53.3664
R3261 GNDA.n305 GNDA.t185 51.7272
R3262 GNDA.n2142 GNDA.n2141 51.3805
R3263 GNDA.n2434 GNDA.n2433 51.2005
R3264 GNDA.n51 GNDA.n50 51.2005
R3265 GNDA.t81 GNDA.n193 50.6495
R3266 GNDA.n2148 GNDA.n2069 50.5752
R3267 GNDA.n2425 GNDA.n2424 50.5752
R3268 GNDA.n510 GNDA.t167 49.5719
R3269 GNDA.t269 GNDA.t174 48.4943
R3270 GNDA.n2367 GNDA.t249 48.4943
R3271 GNDA.t80 GNDA.t255 48.4943
R3272 GNDA.n59 GNDA.t101 48.0005
R3273 GNDA.n59 GNDA.t14 48.0005
R3274 GNDA.n56 GNDA.t127 48.0005
R3275 GNDA.n56 GNDA.t158 48.0005
R3276 GNDA.n55 GNDA.t353 48.0005
R3277 GNDA.n55 GNDA.t16 48.0005
R3278 GNDA.n53 GNDA.t154 48.0005
R3279 GNDA.n53 GNDA.t156 48.0005
R3280 GNDA.n52 GNDA.t57 48.0005
R3281 GNDA.n52 GNDA.t129 48.0005
R3282 GNDA.n1740 GNDA.t219 47.6748
R3283 GNDA.t65 GNDA.t55 46.3607
R3284 GNDA.t19 GNDA.t65 46.3607
R3285 GNDA.t68 GNDA.n2439 46.3607
R3286 GNDA.t75 GNDA.t312 46.3607
R3287 GNDA.t312 GNDA.t9 46.3607
R3288 GNDA.n2281 GNDA.n271 46.339
R3289 GNDA.n2196 GNDA.t219 46.339
R3290 GNDA.t219 GNDA.n1939 46.2335
R3291 GNDA.t219 GNDA.n337 46.2335
R3292 GNDA.t219 GNDA.n1059 46.2335
R3293 GNDA.n1882 GNDA.t269 45.2613
R3294 GNDA.n2279 GNDA.t185 45.2613
R3295 GNDA.n1779 GNDA.t201 45.2613
R3296 GNDA.n2192 GNDA.t120 44.1837
R3297 GNDA.t27 GNDA.t219 43.1061
R3298 GNDA.t167 GNDA.n265 43.1061
R3299 GNDA.t219 GNDA.t81 43.1061
R3300 GNDA.n1791 GNDA.t97 43.1061
R3301 GNDA.t345 GNDA.t219 43.1061
R3302 GNDA.t115 GNDA.t33 42.8925
R3303 GNDA.t137 GNDA.t69 42.8925
R3304 GNDA.n1940 GNDA.t219 42.2987
R3305 GNDA.t219 GNDA.n2037 42.2987
R3306 GNDA.n1060 GNDA.t219 42.2987
R3307 GNDA.t164 GNDA.t225 42.1461
R3308 GNDA.t8 GNDA.t37 42.1461
R3309 GNDA.t309 GNDA.t23 42.1461
R3310 GNDA.t142 GNDA.t25 42.1461
R3311 GNDA.t311 GNDA.t334 42.1461
R3312 GNDA.t161 GNDA.t102 42.1461
R3313 GNDA.t222 GNDA.t121 42.1461
R3314 GNDA.t314 GNDA.t289 42.1461
R3315 GNDA.t111 GNDA.t318 42.1461
R3316 GNDA.t348 GNDA.t322 42.1461
R3317 GNDA.t104 GNDA.t0 42.1461
R3318 GNDA.t94 GNDA.t138 42.1461
R3319 GNDA.t135 GNDA.t140 42.1461
R3320 GNDA.t89 GNDA.t10 42.1461
R3321 GNDA.t146 GNDA.t163 42.1461
R3322 GNDA.t261 GNDA.t350 42.1461
R3323 GNDA.n2171 GNDA.t30 41.1053
R3324 GNDA.t3 GNDA.n2175 41.1053
R3325 GNDA.n2375 GNDA.t110 41.1053
R3326 GNDA.n2397 GNDA.t337 41.1053
R3327 GNDA.n507 GNDA.t181 40.9508
R3328 GNDA.n2211 GNDA.t197 40.9508
R3329 GNDA.n1777 GNDA.t255 40.9508
R3330 GNDA.n2373 GNDA.n187 39.8731
R3331 GNDA.t96 GNDA.n627 39.8731
R3332 GNDA.t44 GNDA.n1777 39.8731
R3333 GNDA.n2131 GNDA.t19 37.9315
R3334 GNDA.n2446 GNDA.t321 37.9315
R3335 GNDA.t48 GNDA.t72 37.9315
R3336 GNDA.n145 GNDA.t75 37.9315
R3337 GNDA.t207 GNDA.t219 37.7179
R3338 GNDA.t187 GNDA.t219 37.7179
R3339 GNDA.n2185 GNDA.t346 37.531
R3340 GNDA.n2388 GNDA.t73 37.531
R3341 GNDA.n2376 GNDA.t73 37.531
R3342 GNDA.n2170 GNDA.n2169 35.7438
R3343 GNDA.n2176 GNDA.n2174 35.7438
R3344 GNDA.n2396 GNDA.n2395 35.7438
R3345 GNDA.n2401 GNDA.n2400 35.7438
R3346 GNDA.n23 GNDA.n22 35.688
R3347 GNDA.n2459 GNDA.n11 35.688
R3348 GNDA.n1882 GNDA.t28 35.5626
R3349 GNDA.n1895 GNDA.t62 35.5626
R3350 GNDA.n1916 GNDA.n1908 35.5626
R3351 GNDA.t71 GNDA.t143 34.5653
R3352 GNDA.t12 GNDA.t351 34.5653
R3353 GNDA.n445 GNDA.t191 34.4849
R3354 GNDA.n2194 GNDA.t213 34.4849
R3355 GNDA.n630 GNDA.t203 34.4849
R3356 GNDA.t346 GNDA.n2184 33.9566
R3357 GNDA.t225 GNDA.t145 33.717
R3358 GNDA.t324 GNDA.t344 33.717
R3359 GNDA.t37 GNDA.t93 33.717
R3360 GNDA.t23 GNDA.t328 33.717
R3361 GNDA.t25 GNDA.t330 33.717
R3362 GNDA.t334 GNDA.t116 33.717
R3363 GNDA.t121 GNDA.t228 33.717
R3364 GNDA.t286 GNDA.t314 33.717
R3365 GNDA.t41 GNDA.t348 33.717
R3366 GNDA.t21 GNDA.t104 33.717
R3367 GNDA.t343 GNDA.t94 33.717
R3368 GNDA.t88 GNDA.t135 33.717
R3369 GNDA.t87 GNDA.t89 33.717
R3370 GNDA.t144 GNDA.t146 33.717
R3371 GNDA.t118 GNDA.t261 33.717
R3372 GNDA.n378 GNDA.t219 32.9056
R3373 GNDA.n1204 GNDA.t219 32.9056
R3374 GNDA.t29 GNDA.n1802 32.3297
R3375 GNDA.n1802 GNDA.n512 32.3297
R3376 GNDA.n2403 GNDA.n165 32.0005
R3377 GNDA.n2167 GNDA.n2166 32.0005
R3378 GNDA.n2393 GNDA.n173 32.0005
R3379 GNDA.n2178 GNDA.n2050 32.0005
R3380 GNDA.n2090 GNDA.t106 30.3614
R3381 GNDA.t143 GNDA.n2083 30.3614
R3382 GNDA.n2079 GNDA.t4 30.3614
R3383 GNDA.n95 GNDA.t340 30.3614
R3384 GNDA.n2417 GNDA.t351 30.3614
R3385 GNDA.n2410 GNDA.t123 30.3614
R3386 GNDA.n1893 GNDA.t189 30.1744
R3387 GNDA.n306 GNDA.t211 30.1744
R3388 GNDA.n611 GNDA.t205 30.1744
R3389 GNDA.t150 GNDA.t159 29.5024
R3390 GNDA.t133 GNDA.t6 29.5024
R3391 GNDA.t58 GNDA.t165 29.5024
R3392 GNDA.t51 GNDA.t316 29.5024
R3393 GNDA.t77 GNDA.n1893 29.0968
R3394 GNDA.n1908 GNDA.t42 29.0968
R3395 GNDA.n1803 GNDA.t29 29.0968
R3396 GNDA.n2138 GNDA.n2137 28.538
R3397 GNDA.n2421 GNDA.n2420 28.538
R3398 GNDA.n149 GNDA.n148 28.163
R3399 GNDA.n2111 GNDA.n2072 28.038
R3400 GNDA.n524 GNDA.n443 27.8193
R3401 GNDA.n1795 GNDA.n1794 27.8193
R3402 GNDA.n591 GNDA.n590 27.5561
R3403 GNDA.n1307 GNDA.n1304 27.5561
R3404 GNDA.n914 GNDA.n911 27.5561
R3405 GNDA.n1392 GNDA.n1389 27.5561
R3406 GNDA.n2255 GNDA.n2252 27.5561
R3407 GNDA.n1000 GNDA.n999 27.5561
R3408 GNDA.n1609 GNDA.n1608 27.5561
R3409 GNDA.n1839 GNDA.n1838 27.5561
R3410 GNDA.n739 GNDA.n738 27.5561
R3411 GNDA.t181 GNDA.t42 26.9415
R3412 GNDA.t201 GNDA.t338 26.9415
R3413 GNDA.n573 GNDA.n572 26.6672
R3414 GNDA.n1288 GNDA.n1287 26.6672
R3415 GNDA.n895 GNDA.n894 26.6672
R3416 GNDA.n1373 GNDA.n1372 26.6672
R3417 GNDA.n2236 GNDA.n2235 26.6672
R3418 GNDA.n982 GNDA.n981 26.6672
R3419 GNDA.n1592 GNDA.n1591 26.6672
R3420 GNDA.n1855 GNDA.n1812 26.6672
R3421 GNDA.n721 GNDA.n720 26.6672
R3422 GNDA.t67 GNDA.n2090 25.6905
R3423 GNDA.n2083 GNDA.t106 25.6905
R3424 GNDA.n95 GNDA.t336 25.6905
R3425 GNDA.n2417 GNDA.t123 25.6905
R3426 GNDA.n2410 GNDA.t341 25.6905
R3427 GNDA.n2134 GNDA.n2133 25.6005
R3428 GNDA.n143 GNDA.n142 25.6005
R3429 GNDA.n645 GNDA.n334 24.8042
R3430 GNDA.t97 GNDA.n1789 24.7862
R3431 GNDA.t338 GNDA.n187 24.7862
R3432 GNDA.n630 GNDA.t91 24.7862
R3433 GNDA.n331 GNDA.t176 24.0005
R3434 GNDA.n331 GNDA.t204 24.0005
R3435 GNDA.n329 GNDA.t206 24.0005
R3436 GNDA.n329 GNDA.t188 24.0005
R3437 GNDA.n327 GNDA.t178 24.0005
R3438 GNDA.n327 GNDA.t202 24.0005
R3439 GNDA.n325 GNDA.t198 24.0005
R3440 GNDA.n325 GNDA.t200 24.0005
R3441 GNDA.n323 GNDA.t184 24.0005
R3442 GNDA.n323 GNDA.t214 24.0005
R3443 GNDA.n321 GNDA.t212 24.0005
R3444 GNDA.n321 GNDA.t194 24.0005
R3445 GNDA.n319 GNDA.t196 24.0005
R3446 GNDA.n319 GNDA.t186 24.0005
R3447 GNDA.n317 GNDA.t182 24.0005
R3448 GNDA.n317 GNDA.t210 24.0005
R3449 GNDA.n315 GNDA.t208 24.0005
R3450 GNDA.n315 GNDA.t192 24.0005
R3451 GNDA.n314 GNDA.t190 24.0005
R3452 GNDA.n314 GNDA.t180 24.0005
R3453 GNDA.n2280 GNDA.t195 23.7086
R3454 GNDA.t177 GNDA.n1778 23.7086
R3455 GNDA.n1070 GNDA.t219 23.6088
R3456 GNDA.n102 GNDA.n34 22.4005
R3457 GNDA.n2450 GNDA.n33 22.4005
R3458 GNDA.n2146 GNDA.n2072 22.4005
R3459 GNDA.n151 GNDA.n149 22.4005
R3460 GNDA.n2461 GNDA.n2460 21.7146
R3461 GNDA.n1917 GNDA.n1916 21.5533
R3462 GNDA.n1792 GNDA.n1791 21.5533
R3463 GNDA.n2373 GNDA.n188 21.5533
R3464 GNDA.n2184 GNDA.n2182 21.4465
R3465 GNDA.n67 GNDA.n63 21.3338
R3466 GNDA.n65 GNDA.n64 21.3338
R3467 GNDA.n51 GNDA.n46 21.3338
R3468 GNDA.n50 GNDA.n47 21.3338
R3469 GNDA.n49 GNDA.n48 21.3338
R3470 GNDA.n2435 GNDA.n43 21.3338
R3471 GNDA.n2434 GNDA.n44 21.3338
R3472 GNDA.n2433 GNDA.n45 21.3338
R3473 GNDA.n78 GNDA.n77 21.3338
R3474 GNDA.n74 GNDA.n73 21.3338
R3475 GNDA.n2123 GNDA.n2122 21.3338
R3476 GNDA.n2124 GNDA.n2121 21.3338
R3477 GNDA.n442 GNDA.n441 21.3338
R3478 GNDA.n440 GNDA.n439 21.3338
R3479 GNDA.n520 GNDA.n519 21.3338
R3480 GNDA.n518 GNDA.n517 21.3338
R3481 GNDA.n644 GNDA.n643 21.3338
R3482 GNDA.n527 GNDA.n526 21.3338
R3483 GNDA.n2100 GNDA.n2099 21.3338
R3484 GNDA.n2096 GNDA.n2095 21.3338
R3485 GNDA.n2102 GNDA.n2101 21.3338
R3486 GNDA.n2104 GNDA.n2103 21.3338
R3487 GNDA.n85 GNDA.n84 21.3338
R3488 GNDA.n137 GNDA.n136 21.3338
R3489 GNDA.n99 GNDA.n98 21.3338
R3490 GNDA.n141 GNDA.n140 21.3338
R3491 GNDA.t102 GNDA.n2442 21.0733
R3492 GNDA.n2454 GNDA.t92 21.0733
R3493 GNDA.n2084 GNDA.t1 21.0196
R3494 GNDA.n2142 GNDA.t1 21.0196
R3495 GNDA.n2141 GNDA.t17 21.0196
R3496 GNDA.n156 GNDA.t86 21.0196
R3497 GNDA.n2042 GNDA.n2041 21.0192
R3498 GNDA.n1799 GNDA.n1798 20.413
R3499 GNDA.n2414 GNDA.n2413 20.288
R3500 GNDA.n2087 GNDA.n2077 20.1943
R3501 GNDA.n2135 GNDA.n2134 19.7255
R3502 GNDA.n142 GNDA.n83 19.7255
R3503 GNDA.n21 GNDA.t59 19.7005
R3504 GNDA.n21 GNDA.t52 19.7005
R3505 GNDA.n19 GNDA.t83 19.7005
R3506 GNDA.n19 GNDA.t76 19.7005
R3507 GNDA.n17 GNDA.t85 19.7005
R3508 GNDA.n17 GNDA.t39 19.7005
R3509 GNDA.n15 GNDA.t60 19.7005
R3510 GNDA.n15 GNDA.t99 19.7005
R3511 GNDA.n13 GNDA.t11 19.7005
R3512 GNDA.n13 GNDA.t131 19.7005
R3513 GNDA.n12 GNDA.t43 19.7005
R3514 GNDA.n12 GNDA.t149 19.7005
R3515 GNDA.n10 GNDA.t172 19.7005
R3516 GNDA.n10 GNDA.t107 19.7005
R3517 GNDA.n8 GNDA.t2 19.7005
R3518 GNDA.n8 GNDA.t326 19.7005
R3519 GNDA.n6 GNDA.t20 19.7005
R3520 GNDA.n6 GNDA.t132 19.7005
R3521 GNDA.n4 GNDA.t124 19.7005
R3522 GNDA.n4 GNDA.t151 19.7005
R3523 GNDA.n2 GNDA.t114 19.7005
R3524 GNDA.n2 GNDA.t327 19.7005
R3525 GNDA.n1 GNDA.t113 19.7005
R3526 GNDA.n1 GNDA.t168 19.7005
R3527 GNDA.n1930 GNDA.t219 19.6741
R3528 GNDA.n508 GNDA.t209 19.398
R3529 GNDA.n2213 GNDA.t199 19.398
R3530 GNDA.n1768 GNDA.n647 19.3019
R3531 GNDA.n2381 GNDA.n2379 19.2005
R3532 GNDA.n309 GNDA.n181 19.2005
R3533 GNDA.n1923 GNDA.n1922 18.9444
R3534 GNDA.n2080 GNDA.n2079 18.6842
R3535 GNDA.n2425 GNDA.n80 18.6842
R3536 GNDA.n341 GNDA.n336 18.5605
R3537 GNDA.n2046 GNDA 18.1546
R3538 GNDA.n2389 GNDA.n2388 17.8721
R3539 GNDA.n2383 GNDA.n181 17.613
R3540 GNDA.n1133 GNDA.n1132 17.5843
R3541 GNDA.n1744 GNDA.n1152 17.5843
R3542 GNDA.n1073 GNDA.n1038 17.5843
R3543 GNDA.n1928 GNDA.n1927 16.9379
R3544 GNDA.n1646 GNDA.n1643 16.9379
R3545 GNDA.n481 GNDA.n478 16.9379
R3546 GNDA.t328 GNDA.n36 16.9236
R3547 GNDA.n2119 GNDA.t155 16.9236
R3548 GNDA.n75 GNDA.t126 16.9236
R3549 GNDA.t343 GNDA.n28 16.9236
R3550 GNDA.t144 GNDA.n29 16.9236
R3551 GNDA.t298 GNDA.t18 16.8587
R3552 GNDA.t329 GNDA.t139 16.8587
R3553 GNDA.t119 GNDA.t98 16.8587
R3554 GNDA.t117 GNDA.t164 16.8587
R3555 GNDA.t145 GNDA.t321 16.8587
R3556 GNDA.t344 GNDA.t8 16.8587
R3557 GNDA.t93 GNDA.t309 16.8587
R3558 GNDA.t328 GNDA.t142 16.8587
R3559 GNDA.t330 GNDA.t311 16.8587
R3560 GNDA.t116 GNDA.t161 16.8587
R3561 GNDA.t22 GNDA.t222 16.8587
R3562 GNDA.t289 GNDA.t92 16.8587
R3563 GNDA.t318 GNDA.t41 16.8587
R3564 GNDA.t322 GNDA.t21 16.8587
R3565 GNDA.t0 GNDA.t343 16.8587
R3566 GNDA.t138 GNDA.t88 16.8587
R3567 GNDA.t140 GNDA.t87 16.8587
R3568 GNDA.t10 GNDA.t144 16.8587
R3569 GNDA.t163 GNDA.t118 16.8587
R3570 GNDA.t350 GNDA.t331 16.8587
R3571 GNDA.t295 GNDA.t339 16.8587
R3572 GNDA.n2157 GNDA.n2152 16.7944
R3573 GNDA.n2312 GNDA.n242 16.7709
R3574 GNDA.n1736 GNDA.n381 16.7709
R3575 GNDA.n1463 GNDA.n377 16.7709
R3576 GNDA.n1218 GNDA.n204 16.7709
R3577 GNDA.t209 GNDA.t173 16.1651
R3578 GNDA.t82 GNDA.t177 16.1651
R3579 GNDA.n605 GNDA.n591 16.0005
R3580 GNDA.n605 GNDA.n604 16.0005
R3581 GNDA.n604 GNDA.n603 16.0005
R3582 GNDA.n603 GNDA.n600 16.0005
R3583 GNDA.n600 GNDA.n599 16.0005
R3584 GNDA.n599 GNDA.n596 16.0005
R3585 GNDA.n596 GNDA.n595 16.0005
R3586 GNDA.n595 GNDA.n592 16.0005
R3587 GNDA.n590 GNDA.n588 16.0005
R3588 GNDA.n588 GNDA.n585 16.0005
R3589 GNDA.n585 GNDA.n584 16.0005
R3590 GNDA.n584 GNDA.n581 16.0005
R3591 GNDA.n581 GNDA.n580 16.0005
R3592 GNDA.n580 GNDA.n577 16.0005
R3593 GNDA.n577 GNDA.n576 16.0005
R3594 GNDA.n576 GNDA.n573 16.0005
R3595 GNDA.n572 GNDA.n569 16.0005
R3596 GNDA.n569 GNDA.n568 16.0005
R3597 GNDA.n568 GNDA.n565 16.0005
R3598 GNDA.n565 GNDA.n564 16.0005
R3599 GNDA.n564 GNDA.n561 16.0005
R3600 GNDA.n561 GNDA.n560 16.0005
R3601 GNDA.n560 GNDA.n543 16.0005
R3602 GNDA.n639 GNDA.n543 16.0005
R3603 GNDA.n1308 GNDA.n1307 16.0005
R3604 GNDA.n1311 GNDA.n1308 16.0005
R3605 GNDA.n1312 GNDA.n1311 16.0005
R3606 GNDA.n1315 GNDA.n1312 16.0005
R3607 GNDA.n1316 GNDA.n1315 16.0005
R3608 GNDA.n1319 GNDA.n1316 16.0005
R3609 GNDA.n1320 GNDA.n1319 16.0005
R3610 GNDA.n1320 GNDA.n1220 16.0005
R3611 GNDA.n1304 GNDA.n1303 16.0005
R3612 GNDA.n1303 GNDA.n1300 16.0005
R3613 GNDA.n1300 GNDA.n1299 16.0005
R3614 GNDA.n1299 GNDA.n1296 16.0005
R3615 GNDA.n1296 GNDA.n1295 16.0005
R3616 GNDA.n1295 GNDA.n1292 16.0005
R3617 GNDA.n1292 GNDA.n1291 16.0005
R3618 GNDA.n1291 GNDA.n1288 16.0005
R3619 GNDA.n1287 GNDA.n1284 16.0005
R3620 GNDA.n1284 GNDA.n1283 16.0005
R3621 GNDA.n1283 GNDA.n1280 16.0005
R3622 GNDA.n1280 GNDA.n1279 16.0005
R3623 GNDA.n1279 GNDA.n1276 16.0005
R3624 GNDA.n1276 GNDA.n1275 16.0005
R3625 GNDA.n1275 GNDA.n1272 16.0005
R3626 GNDA.n1272 GNDA.n1271 16.0005
R3627 GNDA.n915 GNDA.n914 16.0005
R3628 GNDA.n918 GNDA.n915 16.0005
R3629 GNDA.n919 GNDA.n918 16.0005
R3630 GNDA.n922 GNDA.n919 16.0005
R3631 GNDA.n923 GNDA.n922 16.0005
R3632 GNDA.n926 GNDA.n923 16.0005
R3633 GNDA.n927 GNDA.n926 16.0005
R3634 GNDA.n927 GNDA.n825 16.0005
R3635 GNDA.n911 GNDA.n910 16.0005
R3636 GNDA.n910 GNDA.n907 16.0005
R3637 GNDA.n907 GNDA.n906 16.0005
R3638 GNDA.n906 GNDA.n903 16.0005
R3639 GNDA.n903 GNDA.n902 16.0005
R3640 GNDA.n902 GNDA.n899 16.0005
R3641 GNDA.n899 GNDA.n898 16.0005
R3642 GNDA.n898 GNDA.n895 16.0005
R3643 GNDA.n894 GNDA.n891 16.0005
R3644 GNDA.n891 GNDA.n890 16.0005
R3645 GNDA.n890 GNDA.n887 16.0005
R3646 GNDA.n887 GNDA.n886 16.0005
R3647 GNDA.n886 GNDA.n883 16.0005
R3648 GNDA.n883 GNDA.n882 16.0005
R3649 GNDA.n882 GNDA.n879 16.0005
R3650 GNDA.n879 GNDA.n878 16.0005
R3651 GNDA.n1393 GNDA.n1392 16.0005
R3652 GNDA.n1396 GNDA.n1393 16.0005
R3653 GNDA.n1397 GNDA.n1396 16.0005
R3654 GNDA.n1400 GNDA.n1397 16.0005
R3655 GNDA.n1401 GNDA.n1400 16.0005
R3656 GNDA.n1404 GNDA.n1401 16.0005
R3657 GNDA.n1406 GNDA.n1404 16.0005
R3658 GNDA.n1407 GNDA.n1406 16.0005
R3659 GNDA.n1389 GNDA.n1388 16.0005
R3660 GNDA.n1388 GNDA.n1385 16.0005
R3661 GNDA.n1385 GNDA.n1384 16.0005
R3662 GNDA.n1384 GNDA.n1381 16.0005
R3663 GNDA.n1381 GNDA.n1380 16.0005
R3664 GNDA.n1380 GNDA.n1377 16.0005
R3665 GNDA.n1377 GNDA.n1376 16.0005
R3666 GNDA.n1376 GNDA.n1373 16.0005
R3667 GNDA.n1372 GNDA.n1369 16.0005
R3668 GNDA.n1369 GNDA.n1368 16.0005
R3669 GNDA.n1368 GNDA.n1365 16.0005
R3670 GNDA.n1365 GNDA.n1364 16.0005
R3671 GNDA.n1364 GNDA.n1361 16.0005
R3672 GNDA.n1361 GNDA.n1360 16.0005
R3673 GNDA.n1360 GNDA.n1357 16.0005
R3674 GNDA.n1357 GNDA.n1333 16.0005
R3675 GNDA.n2256 GNDA.n2255 16.0005
R3676 GNDA.n2259 GNDA.n2256 16.0005
R3677 GNDA.n2260 GNDA.n2259 16.0005
R3678 GNDA.n2263 GNDA.n2260 16.0005
R3679 GNDA.n2264 GNDA.n2263 16.0005
R3680 GNDA.n2267 GNDA.n2264 16.0005
R3681 GNDA.n2268 GNDA.n2267 16.0005
R3682 GNDA.n2271 GNDA.n2268 16.0005
R3683 GNDA.n2252 GNDA.n2251 16.0005
R3684 GNDA.n2251 GNDA.n2248 16.0005
R3685 GNDA.n2248 GNDA.n2247 16.0005
R3686 GNDA.n2247 GNDA.n2244 16.0005
R3687 GNDA.n2244 GNDA.n2243 16.0005
R3688 GNDA.n2243 GNDA.n2240 16.0005
R3689 GNDA.n2240 GNDA.n2239 16.0005
R3690 GNDA.n2239 GNDA.n2236 16.0005
R3691 GNDA.n2235 GNDA.n2232 16.0005
R3692 GNDA.n2232 GNDA.n2231 16.0005
R3693 GNDA.n2231 GNDA.n2228 16.0005
R3694 GNDA.n2228 GNDA.n2227 16.0005
R3695 GNDA.n2227 GNDA.n2224 16.0005
R3696 GNDA.n2224 GNDA.n2223 16.0005
R3697 GNDA.n2223 GNDA.n2220 16.0005
R3698 GNDA.n2220 GNDA.n2219 16.0005
R3699 GNDA.n1013 GNDA.n1000 16.0005
R3700 GNDA.n1013 GNDA.n1012 16.0005
R3701 GNDA.n1012 GNDA.n1011 16.0005
R3702 GNDA.n1011 GNDA.n1008 16.0005
R3703 GNDA.n1008 GNDA.n1007 16.0005
R3704 GNDA.n1007 GNDA.n1004 16.0005
R3705 GNDA.n1004 GNDA.n1003 16.0005
R3706 GNDA.n1003 GNDA.n800 16.0005
R3707 GNDA.n999 GNDA.n997 16.0005
R3708 GNDA.n997 GNDA.n994 16.0005
R3709 GNDA.n994 GNDA.n993 16.0005
R3710 GNDA.n993 GNDA.n990 16.0005
R3711 GNDA.n990 GNDA.n989 16.0005
R3712 GNDA.n989 GNDA.n986 16.0005
R3713 GNDA.n986 GNDA.n985 16.0005
R3714 GNDA.n985 GNDA.n982 16.0005
R3715 GNDA.n981 GNDA.n978 16.0005
R3716 GNDA.n978 GNDA.n977 16.0005
R3717 GNDA.n977 GNDA.n974 16.0005
R3718 GNDA.n974 GNDA.n973 16.0005
R3719 GNDA.n973 GNDA.n970 16.0005
R3720 GNDA.n970 GNDA.n969 16.0005
R3721 GNDA.n969 GNDA.n966 16.0005
R3722 GNDA.n966 GNDA.n965 16.0005
R3723 GNDA.n1609 GNDA.n1564 16.0005
R3724 GNDA.n1615 GNDA.n1564 16.0005
R3725 GNDA.n1616 GNDA.n1615 16.0005
R3726 GNDA.n1617 GNDA.n1616 16.0005
R3727 GNDA.n1617 GNDA.n1562 16.0005
R3728 GNDA.n1623 GNDA.n1562 16.0005
R3729 GNDA.n1624 GNDA.n1623 16.0005
R3730 GNDA.n1674 GNDA.n1624 16.0005
R3731 GNDA.n1608 GNDA.n1607 16.0005
R3732 GNDA.n1607 GNDA.n1566 16.0005
R3733 GNDA.n1601 GNDA.n1566 16.0005
R3734 GNDA.n1601 GNDA.n1600 16.0005
R3735 GNDA.n1600 GNDA.n1599 16.0005
R3736 GNDA.n1599 GNDA.n1568 16.0005
R3737 GNDA.n1593 GNDA.n1568 16.0005
R3738 GNDA.n1593 GNDA.n1592 16.0005
R3739 GNDA.n1591 GNDA.n1570 16.0005
R3740 GNDA.n1585 GNDA.n1570 16.0005
R3741 GNDA.n1585 GNDA.n1584 16.0005
R3742 GNDA.n1584 GNDA.n1583 16.0005
R3743 GNDA.n1583 GNDA.n1572 16.0005
R3744 GNDA.n1578 GNDA.n1572 16.0005
R3745 GNDA.n1578 GNDA.n1577 16.0005
R3746 GNDA.n1577 GNDA.n1576 16.0005
R3747 GNDA.n2041 GNDA.n2040 16.0005
R3748 GNDA.n2040 GNDA.n336 16.0005
R3749 GNDA.n1838 GNDA.n1837 16.0005
R3750 GNDA.n1837 GNDA.n1818 16.0005
R3751 GNDA.n1832 GNDA.n1818 16.0005
R3752 GNDA.n1832 GNDA.n1831 16.0005
R3753 GNDA.n1831 GNDA.n1830 16.0005
R3754 GNDA.n1830 GNDA.n1821 16.0005
R3755 GNDA.n1824 GNDA.n1821 16.0005
R3756 GNDA.n1824 GNDA.n1823 16.0005
R3757 GNDA.n1839 GNDA.n1816 16.0005
R3758 GNDA.n1845 GNDA.n1816 16.0005
R3759 GNDA.n1846 GNDA.n1845 16.0005
R3760 GNDA.n1847 GNDA.n1846 16.0005
R3761 GNDA.n1847 GNDA.n1814 16.0005
R3762 GNDA.n1853 GNDA.n1814 16.0005
R3763 GNDA.n1854 GNDA.n1853 16.0005
R3764 GNDA.n1855 GNDA.n1854 16.0005
R3765 GNDA.n1861 GNDA.n1812 16.0005
R3766 GNDA.n1862 GNDA.n1861 16.0005
R3767 GNDA.n1863 GNDA.n1862 16.0005
R3768 GNDA.n1863 GNDA.n1810 16.0005
R3769 GNDA.n1868 GNDA.n1810 16.0005
R3770 GNDA.n1869 GNDA.n1868 16.0005
R3771 GNDA.n1869 GNDA.n1808 16.0005
R3772 GNDA.n1876 GNDA.n1808 16.0005
R3773 GNDA.n753 GNDA.n739 16.0005
R3774 GNDA.n753 GNDA.n752 16.0005
R3775 GNDA.n752 GNDA.n751 16.0005
R3776 GNDA.n751 GNDA.n748 16.0005
R3777 GNDA.n748 GNDA.n747 16.0005
R3778 GNDA.n747 GNDA.n744 16.0005
R3779 GNDA.n744 GNDA.n743 16.0005
R3780 GNDA.n743 GNDA.n740 16.0005
R3781 GNDA.n738 GNDA.n736 16.0005
R3782 GNDA.n736 GNDA.n733 16.0005
R3783 GNDA.n733 GNDA.n732 16.0005
R3784 GNDA.n732 GNDA.n729 16.0005
R3785 GNDA.n729 GNDA.n728 16.0005
R3786 GNDA.n728 GNDA.n725 16.0005
R3787 GNDA.n725 GNDA.n724 16.0005
R3788 GNDA.n724 GNDA.n721 16.0005
R3789 GNDA.n720 GNDA.n717 16.0005
R3790 GNDA.n717 GNDA.n716 16.0005
R3791 GNDA.n716 GNDA.n713 16.0005
R3792 GNDA.n713 GNDA.n712 16.0005
R3793 GNDA.n712 GNDA.n709 16.0005
R3794 GNDA.n709 GNDA.n708 16.0005
R3795 GNDA.n708 GNDA.n705 16.0005
R3796 GNDA.n705 GNDA.n655 16.0005
R3797 GNDA.n2370 GNDA.n179 15.363
R3798 GNDA.n1913 GNDA.n179 15.363
R3799 GNDA.t28 GNDA.n506 15.3002
R3800 GNDA.n2043 GNDA.n171 15.113
R3801 GNDA.n512 GNDA.n510 15.0874
R3802 GNDA.n2049 GNDA.n2048 14.6443
R3803 GNDA.n2458 GNDA.n2457 14.6443
R3804 GNDA.n1032 GNDA.n378 14.555
R3805 GNDA.n1547 GNDA.n1204 14.555
R3806 GNDA.t44 GNDA.n539 14.2266
R3807 GNDA.n2430 GNDA.n2429 14.2068
R3808 GNDA.n2430 GNDA.n72 14.2068
R3809 GNDA.n2117 GNDA.n2115 14.0505
R3810 GNDA.n147 GNDA.n131 14.0505
R3811 GNDA.n1792 GNDA.n193 14.0098
R3812 GNDA.n2382 GNDA.n2381 13.8005
R3813 GNDA.n126 GNDA.n33 13.8005
R3814 GNDA.n103 GNDA.n102 13.8005
R3815 GNDA.n2382 GNDA.n182 13.0042
R3816 GNDA.n1895 GNDA.t207 12.9322
R3817 GNDA.n2196 GNDA.t183 12.9322
R3818 GNDA.t175 GNDA.n628 12.9322
R3819 GNDA.n2077 GNDA.n2076 12.8005
R3820 GNDA.n2415 GNDA.n2414 12.8005
R3821 GNDA.t237 GNDA.n2107 12.6442
R3822 GNDA.t152 GNDA.t233 12.6442
R3823 GNDA.t320 GNDA.t63 12.6442
R3824 GNDA.n2442 GNDA.t22 12.6442
R3825 GNDA.n2454 GNDA.t111 12.6442
R3826 GNDA.t310 GNDA.n2453 12.6442
R3827 GNDA.t40 GNDA.t31 12.6442
R3828 GNDA.t46 GNDA.t252 12.6442
R3829 GNDA.t240 GNDA.n81 12.6442
R3830 GNDA.n333 GNDA.n332 12.0667
R3831 GNDA.n1147 GNDA.n1133 11.6369
R3832 GNDA.n1147 GNDA.n1146 11.6369
R3833 GNDA.n1146 GNDA.n1145 11.6369
R3834 GNDA.n1145 GNDA.n1142 11.6369
R3835 GNDA.n1142 GNDA.n1141 11.6369
R3836 GNDA.n1141 GNDA.n1138 11.6369
R3837 GNDA.n1138 GNDA.n1137 11.6369
R3838 GNDA.n1137 GNDA.n1134 11.6369
R3839 GNDA.n1134 GNDA.n641 11.6369
R3840 GNDA.n1771 GNDA.n641 11.6369
R3841 GNDA.n1111 GNDA.n1110 11.6369
R3842 GNDA.n1114 GNDA.n1111 11.6369
R3843 GNDA.n1115 GNDA.n1114 11.6369
R3844 GNDA.n1118 GNDA.n1115 11.6369
R3845 GNDA.n1119 GNDA.n1118 11.6369
R3846 GNDA.n1122 GNDA.n1119 11.6369
R3847 GNDA.n1123 GNDA.n1122 11.6369
R3848 GNDA.n1126 GNDA.n1123 11.6369
R3849 GNDA.n1127 GNDA.n1126 11.6369
R3850 GNDA.n1130 GNDA.n1127 11.6369
R3851 GNDA.n1132 GNDA.n1130 11.6369
R3852 GNDA.n1745 GNDA.n1744 11.6369
R3853 GNDA.n1748 GNDA.n1745 11.6369
R3854 GNDA.n1749 GNDA.n1748 11.6369
R3855 GNDA.n1752 GNDA.n1749 11.6369
R3856 GNDA.n1753 GNDA.n1752 11.6369
R3857 GNDA.n1756 GNDA.n1753 11.6369
R3858 GNDA.n1757 GNDA.n1756 11.6369
R3859 GNDA.n1760 GNDA.n1757 11.6369
R3860 GNDA.n1761 GNDA.n1760 11.6369
R3861 GNDA.n1764 GNDA.n1761 11.6369
R3862 GNDA.n1506 GNDA.n1505 11.6369
R3863 GNDA.n1505 GNDA.n1502 11.6369
R3864 GNDA.n1502 GNDA.n1501 11.6369
R3865 GNDA.n1501 GNDA.n1498 11.6369
R3866 GNDA.n1498 GNDA.n1497 11.6369
R3867 GNDA.n1497 GNDA.n1494 11.6369
R3868 GNDA.n1494 GNDA.n1493 11.6369
R3869 GNDA.n1493 GNDA.n1490 11.6369
R3870 GNDA.n1490 GNDA.n1489 11.6369
R3871 GNDA.n1489 GNDA.n1487 11.6369
R3872 GNDA.n1487 GNDA.n1152 11.6369
R3873 GNDA.n1464 GNDA.n1173 11.6369
R3874 GNDA.n1467 GNDA.n1464 11.6369
R3875 GNDA.n1468 GNDA.n1467 11.6369
R3876 GNDA.n1471 GNDA.n1468 11.6369
R3877 GNDA.n1472 GNDA.n1471 11.6369
R3878 GNDA.n1475 GNDA.n1472 11.6369
R3879 GNDA.n1476 GNDA.n1475 11.6369
R3880 GNDA.n1479 GNDA.n1476 11.6369
R3881 GNDA.n1480 GNDA.n1479 11.6369
R3882 GNDA.n1483 GNDA.n1480 11.6369
R3883 GNDA.n1484 GNDA.n1483 11.6369
R3884 GNDA.n1928 GNDA.n413 11.6369
R3885 GNDA.n1934 GNDA.n413 11.6369
R3886 GNDA.n1935 GNDA.n1934 11.6369
R3887 GNDA.n1936 GNDA.n1935 11.6369
R3888 GNDA.n1936 GNDA.n409 11.6369
R3889 GNDA.n1942 GNDA.n409 11.6369
R3890 GNDA.n1943 GNDA.n1942 11.6369
R3891 GNDA.n1945 GNDA.n1943 11.6369
R3892 GNDA.n1945 GNDA.n1944 11.6369
R3893 GNDA.n1944 GNDA.n405 11.6369
R3894 GNDA.n1952 GNDA.n405 11.6369
R3895 GNDA.n1927 GNDA.n1926 11.6369
R3896 GNDA.n1926 GNDA.n416 11.6369
R3897 GNDA.n783 GNDA.n416 11.6369
R3898 GNDA.n786 GNDA.n783 11.6369
R3899 GNDA.n787 GNDA.n786 11.6369
R3900 GNDA.n790 GNDA.n787 11.6369
R3901 GNDA.n791 GNDA.n790 11.6369
R3902 GNDA.n794 GNDA.n791 11.6369
R3903 GNDA.n796 GNDA.n794 11.6369
R3904 GNDA.n797 GNDA.n796 11.6369
R3905 GNDA.n1643 GNDA.n1642 11.6369
R3906 GNDA.n1642 GNDA.n1639 11.6369
R3907 GNDA.n1639 GNDA.n1638 11.6369
R3908 GNDA.n1638 GNDA.n1635 11.6369
R3909 GNDA.n1635 GNDA.n1634 11.6369
R3910 GNDA.n1634 GNDA.n1631 11.6369
R3911 GNDA.n1631 GNDA.n1630 11.6369
R3912 GNDA.n1630 GNDA.n1627 11.6369
R3913 GNDA.n1627 GNDA.n1626 11.6369
R3914 GNDA.n1626 GNDA.n1172 11.6369
R3915 GNDA.n1737 GNDA.n1172 11.6369
R3916 GNDA.n1647 GNDA.n1646 11.6369
R3917 GNDA.n1650 GNDA.n1647 11.6369
R3918 GNDA.n1651 GNDA.n1650 11.6369
R3919 GNDA.n1654 GNDA.n1651 11.6369
R3920 GNDA.n1655 GNDA.n1654 11.6369
R3921 GNDA.n1658 GNDA.n1655 11.6369
R3922 GNDA.n1659 GNDA.n1658 11.6369
R3923 GNDA.n1662 GNDA.n1659 11.6369
R3924 GNDA.n1664 GNDA.n1662 11.6369
R3925 GNDA.n1665 GNDA.n1664 11.6369
R3926 GNDA.n482 GNDA.n481 11.6369
R3927 GNDA.n485 GNDA.n482 11.6369
R3928 GNDA.n486 GNDA.n485 11.6369
R3929 GNDA.n489 GNDA.n486 11.6369
R3930 GNDA.n490 GNDA.n489 11.6369
R3931 GNDA.n493 GNDA.n490 11.6369
R3932 GNDA.n494 GNDA.n493 11.6369
R3933 GNDA.n497 GNDA.n494 11.6369
R3934 GNDA.n498 GNDA.n497 11.6369
R3935 GNDA.n501 GNDA.n498 11.6369
R3936 GNDA.n241 GNDA.n240 11.6369
R3937 GNDA.n240 GNDA.n237 11.6369
R3938 GNDA.n237 GNDA.n236 11.6369
R3939 GNDA.n236 GNDA.n233 11.6369
R3940 GNDA.n233 GNDA.n232 11.6369
R3941 GNDA.n232 GNDA.n229 11.6369
R3942 GNDA.n229 GNDA.n228 11.6369
R3943 GNDA.n228 GNDA.n226 11.6369
R3944 GNDA.n226 GNDA.n206 11.6369
R3945 GNDA.n2320 GNDA.n206 11.6369
R3946 GNDA.n2321 GNDA.n2320 11.6369
R3947 GNDA.n478 GNDA.n477 11.6369
R3948 GNDA.n477 GNDA.n474 11.6369
R3949 GNDA.n474 GNDA.n473 11.6369
R3950 GNDA.n473 GNDA.n470 11.6369
R3951 GNDA.n470 GNDA.n469 11.6369
R3952 GNDA.n469 GNDA.n466 11.6369
R3953 GNDA.n466 GNDA.n465 11.6369
R3954 GNDA.n465 GNDA.n462 11.6369
R3955 GNDA.n462 GNDA.n461 11.6369
R3956 GNDA.n461 GNDA.n225 11.6369
R3957 GNDA.n2313 GNDA.n225 11.6369
R3958 GNDA.n1074 GNDA.n1073 11.6369
R3959 GNDA.n1077 GNDA.n1074 11.6369
R3960 GNDA.n1078 GNDA.n1077 11.6369
R3961 GNDA.n1081 GNDA.n1078 11.6369
R3962 GNDA.n1082 GNDA.n1081 11.6369
R3963 GNDA.n1085 GNDA.n1082 11.6369
R3964 GNDA.n1086 GNDA.n1085 11.6369
R3965 GNDA.n1089 GNDA.n1086 11.6369
R3966 GNDA.n1090 GNDA.n1089 11.6369
R3967 GNDA.n1093 GNDA.n1090 11.6369
R3968 GNDA.n1049 GNDA.n346 11.6369
R3969 GNDA.n1049 GNDA.n1046 11.6369
R3970 GNDA.n1055 GNDA.n1046 11.6369
R3971 GNDA.n1056 GNDA.n1055 11.6369
R3972 GNDA.n1057 GNDA.n1056 11.6369
R3973 GNDA.n1057 GNDA.n1042 11.6369
R3974 GNDA.n1063 GNDA.n1042 11.6369
R3975 GNDA.n1064 GNDA.n1063 11.6369
R3976 GNDA.n1066 GNDA.n1064 11.6369
R3977 GNDA.n1066 GNDA.n1065 11.6369
R3978 GNDA.n1065 GNDA.n1038 11.6369
R3979 GNDA.n1963 GNDA.n1954 11.6369
R3980 GNDA.n1963 GNDA.n1962 11.6369
R3981 GNDA.n1962 GNDA.n1961 11.6369
R3982 GNDA.n1961 GNDA.n1956 11.6369
R3983 GNDA.n1956 GNDA.n1955 11.6369
R3984 GNDA.n2035 GNDA.n2034 11.6369
R3985 GNDA.n2034 GNDA.n2033 11.6369
R3986 GNDA.n2033 GNDA.n342 11.6369
R3987 GNDA.n2027 GNDA.n342 11.6369
R3988 GNDA.n2027 GNDA.n2026 11.6369
R3989 GNDA.n2432 GNDA.n2431 11.0505
R3990 GNDA.n521 GNDA.n265 10.7769
R3991 GNDA.t219 GNDA.n189 10.7769
R3992 GNDA.n103 GNDA.n0 9.938
R3993 GNDA.n2385 GNDA.n2384 9.78488
R3994 GNDA.n1923 GNDA.n310 9.65119
R3995 GNDA.n127 GNDA.n126 9.6255
R3996 GNDA.n104 GNDA.t325 9.6005
R3997 GNDA.n104 GNDA.t38 9.6005
R3998 GNDA.n106 GNDA.t24 9.6005
R3999 GNDA.n106 GNDA.t26 9.6005
R4000 GNDA.n108 GNDA.t335 9.6005
R4001 GNDA.n108 GNDA.t103 9.6005
R4002 GNDA.n110 GNDA.t122 9.6005
R4003 GNDA.n110 GNDA.t109 9.6005
R4004 GNDA.n112 GNDA.t50 9.6005
R4005 GNDA.n112 GNDA.t354 9.6005
R4006 GNDA.n114 GNDA.t79 9.6005
R4007 GNDA.n114 GNDA.t323 9.6005
R4008 GNDA.n116 GNDA.t36 9.6005
R4009 GNDA.n116 GNDA.t315 9.6005
R4010 GNDA.n118 GNDA.t112 9.6005
R4011 GNDA.n118 GNDA.t349 9.6005
R4012 GNDA.n120 GNDA.t105 9.6005
R4013 GNDA.n120 GNDA.t95 9.6005
R4014 GNDA.n122 GNDA.t136 9.6005
R4015 GNDA.n122 GNDA.t90 9.6005
R4016 GNDA.n124 GNDA.t147 9.6005
R4017 GNDA.n124 GNDA.t262 9.6005
R4018 GNDA.n2380 GNDA.t169 9.6005
R4019 GNDA.n2380 GNDA.t45 9.6005
R4020 GNDA.n180 GNDA.t171 9.6005
R4021 GNDA.n180 GNDA.t170 9.6005
R4022 GNDA.n71 GNDA.n70 9.3005
R4023 GNDA.n1768 GNDA.n174 9.29376
R4024 GNDA.n2046 GNDA 9.2432
R4025 GNDA.n1894 GNDA.t179 8.62161
R4026 GNDA.n2192 GNDA.t193 8.62161
R4027 GNDA.n627 GNDA.t187 8.62161
R4028 GNDA.n1999 GNDA.n378 8.60107
R4029 GNDA.n1543 GNDA.n1204 8.60107
R4030 GNDA.n2439 GNDA.t72 8.42962
R4031 GNDA.n1922 GNDA.t219 8.22146
R4032 GNDA.n647 GNDA.t219 8.22146
R4033 GNDA.n2384 GNDA.n179 7.71925
R4034 GNDA.n2045 GNDA.n2044 7.56675
R4035 GNDA.n2047 GNDA.n2046 7.56675
R4036 GNDA.t162 GNDA.n508 7.54397
R4037 GNDA.n611 GNDA.t345 7.54397
R4038 GNDA.n629 GNDA.t80 7.54397
R4039 GNDA.n2080 GNDA.t17 7.00687
R4040 GNDA.n2459 GNDA.n2458 6.7505
R4041 GNDA.n1484 GNDA.n1463 6.72373
R4042 GNDA.n1953 GNDA.n1952 6.72373
R4043 GNDA.n1737 GNDA.n1736 6.72373
R4044 GNDA.n2321 GNDA.n204 6.72373
R4045 GNDA.n2313 GNDA.n2312 6.72373
R4046 GNDA.n2026 GNDA.n2025 6.72373
R4047 GNDA.n2458 GNDA.n23 6.688
R4048 GNDA.n2114 GNDA.n0 6.563
R4049 GNDA.n129 GNDA.n127 6.563
R4050 GNDA.t120 GNDA.t219 6.46633
R4051 GNDA.n539 GNDA.t219 6.44277
R4052 GNDA.n2137 GNDA.n2136 6.4005
R4053 GNDA.n2422 GNDA.n2421 6.4005
R4054 GNDA GNDA.n2045 6.25048
R4055 GNDA.n1110 GNDA.n204 6.20656
R4056 GNDA.n1506 GNDA.n1463 6.20656
R4057 GNDA.n1736 GNDA.n1173 6.20656
R4058 GNDA.n2312 GNDA.n241 6.20656
R4059 GNDA.n2025 GNDA.n346 6.20656
R4060 GNDA.n1954 GNDA.n1953 6.20656
R4061 GNDA.n1955 GNDA.n341 6.07727
R4062 GNDA.n2035 GNDA.n341 5.5601
R4063 GNDA.n1774 GNDA.n639 5.51161
R4064 GNDA.n1271 GNDA.n1241 5.51161
R4065 GNDA.n878 GNDA.n848 5.51161
R4066 GNDA.n1443 GNDA.n1333 5.51161
R4067 GNDA.n2219 GNDA.n295 5.51161
R4068 GNDA.n965 GNDA.n943 5.51161
R4069 GNDA.n1576 GNDA.n1202 5.51161
R4070 GNDA.n1877 GNDA.n1876 5.51161
R4071 GNDA.n1036 GNDA.n655 5.51161
R4072 GNDA.n1917 GNDA.t191 5.3887
R4073 GNDA.t193 GNDA.n2191 5.3887
R4074 GNDA.t183 GNDA.n2195 5.3887
R4075 GNDA.t355 GNDA.t275 5.3887
R4076 GNDA.t205 GNDA.n188 5.3887
R4077 GNDA.n506 GNDA.t219 5.36915
R4078 GNDA.n2185 GNDA.t78 5.36199
R4079 GNDA.n2376 GNDA.t141 5.36199
R4080 GNDA.n1773 GNDA.n1772 5.1717
R4081 GNDA.n1765 GNDA.n1151 5.1717
R4082 GNDA.n1094 GNDA.n1037 5.1717
R4083 GNDA.n127 GNDA.n23 5.03175
R4084 GNDA.n1029 GNDA.n799 4.9157
R4085 GNDA.n1671 GNDA.n1667 4.9157
R4086 GNDA.n504 GNDA.n503 4.9157
R4087 GNDA.n60 GNDA.n58 4.5005
R4088 GNDA.n2431 GNDA.n2430 4.5005
R4089 GNDA.n2384 GNDA.n2383 4.5005
R4090 GNDA.n2460 GNDA.n2459 4.5005
R4091 GNDA.n2311 GNDA.n243 4.26717
R4092 GNDA.n2305 GNDA.n243 4.26717
R4093 GNDA.n2305 GNDA.n2304 4.26717
R4094 GNDA.n2304 GNDA.n2303 4.26717
R4095 GNDA.n2303 GNDA.n252 4.26717
R4096 GNDA.n255 GNDA.n252 4.26717
R4097 GNDA.n2294 GNDA.n255 4.26717
R4098 GNDA.n2294 GNDA.n2293 4.26717
R4099 GNDA.n2293 GNDA.n2292 4.26717
R4100 GNDA.n2292 GNDA.n260 4.26717
R4101 GNDA.n2286 GNDA.n260 4.26717
R4102 GNDA.n1735 GNDA.n1174 4.26717
R4103 GNDA.n1730 GNDA.n1174 4.26717
R4104 GNDA.n1730 GNDA.n1729 4.26717
R4105 GNDA.n1729 GNDA.n1728 4.26717
R4106 GNDA.n1728 GNDA.n1725 4.26717
R4107 GNDA.n1725 GNDA.n1724 4.26717
R4108 GNDA.n1724 GNDA.n1721 4.26717
R4109 GNDA.n1721 GNDA.n1720 4.26717
R4110 GNDA.n1720 GNDA.n1717 4.26717
R4111 GNDA.n1717 GNDA.n1716 4.26717
R4112 GNDA.n1716 GNDA.n1714 4.26717
R4113 GNDA.n1971 GNDA.n400 4.26717
R4114 GNDA.n1971 GNDA.n396 4.26717
R4115 GNDA.n1977 GNDA.n396 4.26717
R4116 GNDA.n1978 GNDA.n1977 4.26717
R4117 GNDA.n1978 GNDA.n393 4.26717
R4118 GNDA.n393 GNDA.n391 4.26717
R4119 GNDA.n1986 GNDA.n391 4.26717
R4120 GNDA.n1986 GNDA.n387 4.26717
R4121 GNDA.n1992 GNDA.n387 4.26717
R4122 GNDA.n1993 GNDA.n1992 4.26717
R4123 GNDA.n1993 GNDA.n384 4.26717
R4124 GNDA.n2024 GNDA.n348 4.26717
R4125 GNDA.n2018 GNDA.n348 4.26717
R4126 GNDA.n2018 GNDA.n2017 4.26717
R4127 GNDA.n2017 GNDA.n2016 4.26717
R4128 GNDA.n2016 GNDA.n2014 4.26717
R4129 GNDA.n2014 GNDA.n2011 4.26717
R4130 GNDA.n2011 GNDA.n2010 4.26717
R4131 GNDA.n2010 GNDA.n2007 4.26717
R4132 GNDA.n2007 GNDA.n2006 4.26717
R4133 GNDA.n2006 GNDA.n2003 4.26717
R4134 GNDA.n2003 GNDA.n2002 4.26717
R4135 GNDA.n1511 GNDA.n1510 4.26717
R4136 GNDA.n1514 GNDA.n1511 4.26717
R4137 GNDA.n1514 GNDA.n1459 4.26717
R4138 GNDA.n1520 GNDA.n1459 4.26717
R4139 GNDA.n1521 GNDA.n1520 4.26717
R4140 GNDA.n1524 GNDA.n1521 4.26717
R4141 GNDA.n1524 GNDA.n1457 4.26717
R4142 GNDA.n1530 GNDA.n1457 4.26717
R4143 GNDA.n1530 GNDA.n1450 4.26717
R4144 GNDA.n1538 GNDA.n1450 4.26717
R4145 GNDA.n1538 GNDA.n1447 4.26717
R4146 GNDA.n2358 GNDA.n2357 4.26717
R4147 GNDA.n2357 GNDA.n2356 4.26717
R4148 GNDA.n2356 GNDA.n2355 4.26717
R4149 GNDA.n2355 GNDA.n2353 4.26717
R4150 GNDA.n2353 GNDA.n2350 4.26717
R4151 GNDA.n2350 GNDA.n2349 4.26717
R4152 GNDA.n2349 GNDA.n2346 4.26717
R4153 GNDA.n2346 GNDA.n2345 4.26717
R4154 GNDA.n2345 GNDA.n2342 4.26717
R4155 GNDA.n2342 GNDA.n2341 4.26717
R4156 GNDA.n2341 GNDA.n196 4.26717
R4157 GNDA.t304 GNDA.t245 4.21506
R4158 GNDA.n2128 GNDA.t119 4.21506
R4159 GNDA.n2446 GNDA.t324 4.21506
R4160 GNDA.n2453 GNDA.t134 4.21506
R4161 GNDA.t258 GNDA.t216 4.21506
R4162 GNDA.n2312 GNDA.n2311 3.93531
R4163 GNDA.n1736 GNDA.n1735 3.93531
R4164 GNDA.n1953 GNDA.n400 3.93531
R4165 GNDA.n2025 GNDA.n2024 3.93531
R4166 GNDA.n1510 GNDA.n1463 3.93531
R4167 GNDA.n2358 GNDA.n204 3.93531
R4168 GNDA.n2383 GNDA.n2382 3.813
R4169 GNDA.n1786 GNDA.n1785 3.7893
R4170 GNDA.n1782 GNDA.n534 3.7893
R4171 GNDA.n1781 GNDA.n537 3.7893
R4172 GNDA.n618 GNDA.n616 3.7893
R4173 GNDA.n617 GNDA.n614 3.7893
R4174 GNDA.n613 GNDA.n609 3.7893
R4175 GNDA.n634 GNDA.n632 3.7893
R4176 GNDA.n633 GNDA.n542 3.7893
R4177 GNDA.n1330 GNDA.n1221 3.7893
R4178 GNDA.n1327 GNDA.n1326 3.7893
R4179 GNDA.n1243 GNDA.n1222 3.7893
R4180 GNDA.n1248 GNDA.n1246 3.7893
R4181 GNDA.n1253 GNDA.n1249 3.7893
R4182 GNDA.n1260 GNDA.n1259 3.7893
R4183 GNDA.n1263 GNDA.n1242 3.7893
R4184 GNDA.n1268 GNDA.n1264 3.7893
R4185 GNDA.n937 GNDA.n826 3.7893
R4186 GNDA.n934 GNDA.n933 3.7893
R4187 GNDA.n850 GNDA.n827 3.7893
R4188 GNDA.n855 GNDA.n853 3.7893
R4189 GNDA.n860 GNDA.n856 3.7893
R4190 GNDA.n867 GNDA.n866 3.7893
R4191 GNDA.n870 GNDA.n849 3.7893
R4192 GNDA.n875 GNDA.n871 3.7893
R4193 GNDA.n1433 GNDA.n1409 3.7893
R4194 GNDA.n1432 GNDA.n1430 3.7893
R4195 GNDA.n1429 GNDA.n1410 3.7893
R4196 GNDA.n1426 GNDA.n1425 3.7893
R4197 GNDA.n1422 GNDA.n1411 3.7893
R4198 GNDA.n1415 GNDA.n1412 3.7893
R4199 GNDA.n1438 GNDA.n1335 3.7893
R4200 GNDA.n1439 GNDA.n1334 3.7893
R4201 GNDA.n2269 GNDA.n273 3.7893
R4202 GNDA.n2277 GNDA.n2276 3.7893
R4203 GNDA.n300 GNDA.n274 3.7893
R4204 GNDA.n303 GNDA.n302 3.7893
R4205 GNDA.n2199 GNDA.n299 3.7893
R4206 GNDA.n2204 GNDA.n2203 3.7893
R4207 GNDA.n2208 GNDA.n2207 3.7893
R4208 GNDA.n2216 GNDA.n296 3.7893
R4209 GNDA.n1027 GNDA.n1026 3.7893
R4210 GNDA.n1023 GNDA.n802 3.7893
R4211 GNDA.n1022 GNDA.n805 3.7893
R4212 GNDA.n1019 GNDA.n1018 3.7893
R4213 GNDA.n945 GNDA.n806 3.7893
R4214 GNDA.n954 GNDA.n953 3.7893
R4215 GNDA.n957 GNDA.n944 3.7893
R4216 GNDA.n962 GNDA.n958 3.7893
R4217 GNDA.n1672 GNDA.n1560 3.7893
R4218 GNDA.n1681 GNDA.n1680 3.7893
R4219 GNDA.n1558 GNDA.n1557 3.7893
R4220 GNDA.n1689 GNDA.n1687 3.7893
R4221 GNDA.n1688 GNDA.n1555 3.7893
R4222 GNDA.n1553 GNDA.n1552 3.7893
R4223 GNDA.n1703 GNDA.n1702 3.7893
R4224 GNDA.n1707 GNDA.n1549 3.7893
R4225 GNDA.n1885 GNDA.n1884 3.7893
R4226 GNDA.n1889 GNDA.n457 3.7893
R4227 GNDA.n1891 GNDA.n1890 3.7893
R4228 GNDA.n1898 GNDA.n454 3.7893
R4229 GNDA.n1897 GNDA.n452 3.7893
R4230 GNDA.n1906 GNDA.n1905 3.7893
R4231 GNDA.n1805 GNDA.n449 3.7893
R4232 GNDA.n1807 GNDA.n1806 3.7893
R4233 GNDA.n767 GNDA.n766 3.7893
R4234 GNDA.n763 GNDA.n665 3.7893
R4235 GNDA.n762 GNDA.n668 3.7893
R4236 GNDA.n759 GNDA.n758 3.7893
R4237 GNDA.n677 GNDA.n669 3.7893
R4238 GNDA.n683 GNDA.n676 3.7893
R4239 GNDA.n688 GNDA.n686 3.7893
R4240 GNDA.n687 GNDA.n656 3.7893
R4241 GNDA GNDA.n624 3.7381
R4242 GNDA.n1256 GNDA 3.7381
R4243 GNDA.n863 GNDA 3.7381
R4244 GNDA GNDA.n1418 3.7381
R4245 GNDA.n2202 GNDA 3.7381
R4246 GNDA.n950 GNDA 3.7381
R4247 GNDA GNDA.n1695 3.7381
R4248 GNDA GNDA.n448 3.7381
R4249 GNDA.n682 GNDA 3.7381
R4250 GNDA.n2113 GNDA.t7 3.42907
R4251 GNDA.n2113 GNDA.t64 3.42907
R4252 GNDA.n2112 GNDA.t160 3.42907
R4253 GNDA.n2112 GNDA.t66 3.42907
R4254 GNDA.n130 GNDA.t313 3.42907
R4255 GNDA.n130 GNDA.t317 3.42907
R4256 GNDA.n128 GNDA.t32 3.42907
R4257 GNDA.n128 GNDA.t166 3.42907
R4258 GNDA.n2045 GNDA.n334 3.41975
R4259 GNDA.t174 GNDA.n1881 3.23342
R4260 GNDA.n445 GNDA.t27 3.23342
R4261 GNDA.t61 GNDA.n1880 3.23342
R4262 GNDA.n1778 GNDA.t332 3.23342
R4263 GNDA.n533 GNDA.n532 2.6629
R4264 GNDA.n1332 GNDA.n1331 2.6629
R4265 GNDA.n939 GNDA.n938 2.6629
R4266 GNDA.n847 GNDA.n375 2.6629
R4267 GNDA.n1408 GNDA.n1201 2.6629
R4268 GNDA.n1446 GNDA.n1445 2.6629
R4269 GNDA.n2270 GNDA.n267 2.6629
R4270 GNDA.n294 GNDA.n192 2.6629
R4271 GNDA.n1029 GNDA.n1028 2.6629
R4272 GNDA.n942 GNDA.n940 2.6629
R4273 GNDA.n1673 GNDA.n1671 2.6629
R4274 GNDA.n1713 GNDA.n1712 2.6629
R4275 GNDA.n504 GNDA.n459 2.6629
R4276 GNDA.n2285 GNDA.n268 2.6629
R4277 GNDA.n664 GNDA.n663 2.6629
R4278 GNDA.n532 GNDA.n192 2.4581
R4279 GNDA.n1774 GNDA.n1773 2.4581
R4280 GNDA.n1446 GNDA.n1332 2.4581
R4281 GNDA.n1241 GNDA.n1151 2.4581
R4282 GNDA.n940 GNDA.n939 2.4581
R4283 GNDA.n848 GNDA.n847 2.4581
R4284 GNDA.n1713 GNDA.n1201 2.4581
R4285 GNDA.n1445 GNDA.n1443 2.4581
R4286 GNDA.n2285 GNDA.n267 2.4581
R4287 GNDA.n295 GNDA.n294 2.4581
R4288 GNDA.n943 GNDA.n942 2.4581
R4289 GNDA.n1712 GNDA.n1202 2.4581
R4290 GNDA.n1877 GNDA.n268 2.4581
R4291 GNDA.n663 GNDA.n375 2.4581
R4292 GNDA.n1037 GNDA.n1036 2.4581
R4293 GNDA.n320 GNDA.n318 2.34425
R4294 GNDA.n328 GNDA.n326 2.34425
R4295 GNDA.t336 GNDA.n93 2.33596
R4296 GNDA.t86 GNDA.n155 2.33596
R4297 GNDA.n2286 GNDA.n2285 2.18124
R4298 GNDA.n1714 GNDA.n1713 2.18124
R4299 GNDA.n940 GNDA.n384 2.18124
R4300 GNDA.n2002 GNDA.n375 2.18124
R4301 GNDA.n1447 GNDA.n1446 2.18124
R4302 GNDA.n196 GNDA.n192 2.18124
R4303 GNDA.n1880 GNDA.t272 2.15578
R4304 GNDA.n2281 GNDA.t301 2.15578
R4305 GNDA.n2212 GNDA.t249 2.15578
R4306 GNDA.n1788 GNDA.t275 2.15578
R4307 GNDA.n1775 GNDA.n1774 2.1509
R4308 GNDA.n1267 GNDA.n1241 2.1509
R4309 GNDA.n874 GNDA.n848 2.1509
R4310 GNDA.n1443 GNDA.n1442 2.1509
R4311 GNDA.n2215 GNDA.n295 2.1509
R4312 GNDA.n961 GNDA.n943 2.1509
R4313 GNDA.n1708 GNDA.n1202 2.1509
R4314 GNDA.n1878 GNDA.n1877 2.1509
R4315 GNDA.n1036 GNDA.n1035 2.1509
R4316 GNDA.n592 GNDA.n533 2.13383
R4317 GNDA.n1331 GNDA.n1220 2.13383
R4318 GNDA.n938 GNDA.n825 2.13383
R4319 GNDA.n1408 GNDA.n1407 2.13383
R4320 GNDA.n2271 GNDA.n2270 2.13383
R4321 GNDA.n1028 GNDA.n800 2.13383
R4322 GNDA.n1674 GNDA.n1673 2.13383
R4323 GNDA.n1823 GNDA.n459 2.13383
R4324 GNDA.n740 GNDA.n664 2.13383
R4325 GNDA GNDA.n182 2.09787
R4326 GNDA.n2285 GNDA.n2284 2.08643
R4327 GNDA.n1713 GNDA.n242 2.08643
R4328 GNDA.n940 GNDA.n381 2.08643
R4329 GNDA.n377 GNDA.n375 2.08643
R4330 GNDA.n1446 GNDA.n1218 2.08643
R4331 GNDA.n2364 GNDA.n192 2.08643
R4332 GNDA.n1786 GNDA.n533 1.9461
R4333 GNDA.n1331 GNDA.n1330 1.9461
R4334 GNDA.n938 GNDA.n937 1.9461
R4335 GNDA.n1409 GNDA.n1408 1.9461
R4336 GNDA.n2270 GNDA.n2269 1.9461
R4337 GNDA.n1028 GNDA.n1027 1.9461
R4338 GNDA.n1673 GNDA.n1672 1.9461
R4339 GNDA.n1884 GNDA.n459 1.9461
R4340 GNDA.n767 GNDA.n664 1.9461
R4341 GNDA.t125 GNDA.n2054 1.78766
R4342 GNDA.n2171 GNDA.t115 1.78766
R4343 GNDA.n2175 GNDA.t78 1.78766
R4344 GNDA.t141 GNDA.n2375 1.78766
R4345 GNDA.n2397 GNDA.t137 1.78766
R4346 GNDA.t148 GNDA.n161 1.78766
R4347 GNDA.n2457 GNDA.n24 1.6005
R4348 GNDA.n2044 GNDA.n2043 1.5005
R4349 GNDA.n2048 GNDA.n2047 1.5005
R4350 GNDA.n1772 GNDA.n1771 1.47392
R4351 GNDA.n1765 GNDA.n1764 1.47392
R4352 GNDA.n799 GNDA.n797 1.47392
R4353 GNDA.n1667 GNDA.n1665 1.47392
R4354 GNDA.n503 GNDA.n501 1.47392
R4355 GNDA.n1094 GNDA.n1093 1.47392
R4356 GNDA.n2431 GNDA.n71 1.188
R4357 GNDA GNDA.n2461 0.9405
R4358 GNDA.n1785 GNDA.n534 0.8197
R4359 GNDA.n1782 GNDA.n1781 0.8197
R4360 GNDA.n616 GNDA.n537 0.8197
R4361 GNDA.n618 GNDA.n617 0.8197
R4362 GNDA.n624 GNDA.n613 0.8197
R4363 GNDA.n632 GNDA.n609 0.8197
R4364 GNDA.n634 GNDA.n633 0.8197
R4365 GNDA.n1775 GNDA.n542 0.8197
R4366 GNDA.n1327 GNDA.n1221 0.8197
R4367 GNDA.n1326 GNDA.n1222 0.8197
R4368 GNDA.n1246 GNDA.n1243 0.8197
R4369 GNDA.n1249 GNDA.n1248 0.8197
R4370 GNDA.n1259 GNDA.n1256 0.8197
R4371 GNDA.n1260 GNDA.n1242 0.8197
R4372 GNDA.n1264 GNDA.n1263 0.8197
R4373 GNDA.n1268 GNDA.n1267 0.8197
R4374 GNDA.n934 GNDA.n826 0.8197
R4375 GNDA.n933 GNDA.n827 0.8197
R4376 GNDA.n853 GNDA.n850 0.8197
R4377 GNDA.n856 GNDA.n855 0.8197
R4378 GNDA.n866 GNDA.n863 0.8197
R4379 GNDA.n867 GNDA.n849 0.8197
R4380 GNDA.n871 GNDA.n870 0.8197
R4381 GNDA.n875 GNDA.n874 0.8197
R4382 GNDA.n1433 GNDA.n1432 0.8197
R4383 GNDA.n1430 GNDA.n1429 0.8197
R4384 GNDA.n1426 GNDA.n1410 0.8197
R4385 GNDA.n1425 GNDA.n1422 0.8197
R4386 GNDA.n1418 GNDA.n1415 0.8197
R4387 GNDA.n1412 GNDA.n1335 0.8197
R4388 GNDA.n1439 GNDA.n1438 0.8197
R4389 GNDA.n1442 GNDA.n1334 0.8197
R4390 GNDA.n2277 GNDA.n273 0.8197
R4391 GNDA.n2276 GNDA.n274 0.8197
R4392 GNDA.n303 GNDA.n300 0.8197
R4393 GNDA.n302 GNDA.n299 0.8197
R4394 GNDA.n2203 GNDA.n2202 0.8197
R4395 GNDA.n2208 GNDA.n2204 0.8197
R4396 GNDA.n2207 GNDA.n296 0.8197
R4397 GNDA.n2216 GNDA.n2215 0.8197
R4398 GNDA.n1026 GNDA.n802 0.8197
R4399 GNDA.n1023 GNDA.n1022 0.8197
R4400 GNDA.n1019 GNDA.n805 0.8197
R4401 GNDA.n1018 GNDA.n806 0.8197
R4402 GNDA.n953 GNDA.n950 0.8197
R4403 GNDA.n954 GNDA.n944 0.8197
R4404 GNDA.n958 GNDA.n957 0.8197
R4405 GNDA.n962 GNDA.n961 0.8197
R4406 GNDA.n1681 GNDA.n1560 0.8197
R4407 GNDA.n1680 GNDA.n1558 0.8197
R4408 GNDA.n1687 GNDA.n1557 0.8197
R4409 GNDA.n1689 GNDA.n1688 0.8197
R4410 GNDA.n1695 GNDA.n1553 0.8197
R4411 GNDA.n1702 GNDA.n1552 0.8197
R4412 GNDA.n1703 GNDA.n1549 0.8197
R4413 GNDA.n1708 GNDA.n1707 0.8197
R4414 GNDA.n1885 GNDA.n457 0.8197
R4415 GNDA.n1891 GNDA.n1889 0.8197
R4416 GNDA.n1890 GNDA.n454 0.8197
R4417 GNDA.n1898 GNDA.n1897 0.8197
R4418 GNDA.n1906 GNDA.n448 0.8197
R4419 GNDA.n1905 GNDA.n449 0.8197
R4420 GNDA.n1806 GNDA.n1805 0.8197
R4421 GNDA.n1878 GNDA.n1807 0.8197
R4422 GNDA.n766 GNDA.n665 0.8197
R4423 GNDA.n763 GNDA.n762 0.8197
R4424 GNDA.n759 GNDA.n668 0.8197
R4425 GNDA.n758 GNDA.n669 0.8197
R4426 GNDA.n683 GNDA.n682 0.8197
R4427 GNDA.n686 GNDA.n676 0.8197
R4428 GNDA.n688 GNDA.n687 0.8197
R4429 GNDA.n1035 GNDA.n656 0.8197
R4430 GNDA.n105 GNDA.n103 0.59425
R4431 GNDA.n614 GNDA 0.5637
R4432 GNDA.n1253 GNDA 0.5637
R4433 GNDA.n860 GNDA 0.5637
R4434 GNDA GNDA.n1411 0.5637
R4435 GNDA.n2199 GNDA 0.5637
R4436 GNDA GNDA.n945 0.5637
R4437 GNDA.n1555 GNDA 0.5637
R4438 GNDA.n452 GNDA 0.5637
R4439 GNDA GNDA.n677 0.5637
R4440 GNDA.n16 GNDA.n14 0.563
R4441 GNDA.n18 GNDA.n16 0.563
R4442 GNDA.n20 GNDA.n18 0.563
R4443 GNDA.n22 GNDA.n20 0.563
R4444 GNDA.n58 GNDA.n57 0.563
R4445 GNDA.n58 GNDA.n54 0.563
R4446 GNDA.n318 GNDA.n316 0.563
R4447 GNDA.n322 GNDA.n320 0.563
R4448 GNDA.n324 GNDA.n322 0.563
R4449 GNDA.n326 GNDA.n324 0.563
R4450 GNDA.n330 GNDA.n328 0.563
R4451 GNDA.n332 GNDA.n330 0.563
R4452 GNDA.n5 GNDA.n3 0.563
R4453 GNDA.n7 GNDA.n5 0.563
R4454 GNDA.n9 GNDA.n7 0.563
R4455 GNDA.n11 GNDA.n9 0.563
R4456 GNDA.n125 GNDA.n123 0.563
R4457 GNDA.n123 GNDA.n121 0.563
R4458 GNDA.n121 GNDA.n119 0.563
R4459 GNDA.n119 GNDA.n117 0.563
R4460 GNDA.n117 GNDA.n115 0.563
R4461 GNDA.n115 GNDA.n113 0.563
R4462 GNDA.n113 GNDA.n111 0.563
R4463 GNDA.n111 GNDA.n109 0.563
R4464 GNDA.n109 GNDA.n107 0.563
R4465 GNDA.n107 GNDA.n105 0.563
R4466 GNDA.n2460 GNDA.n0 0.53175
R4467 GNDA.n2115 GNDA.n2114 0.5005
R4468 GNDA.n131 GNDA.n129 0.5005
R4469 GNDA.n2084 GNDA.t71 0.467591
R4470 GNDA.n156 GNDA.t12 0.467591
R4471 GNDA.n2043 GNDA.n2042 0.28175
R4472 GNDA.n126 GNDA.n125 0.28175
R4473 GNDA.n313 GNDA.n182 0.276625
R4474 GNDA.n625 GNDA 0.2565
R4475 GNDA GNDA.n1252 0.2565
R4476 GNDA GNDA.n859 0.2565
R4477 GNDA.n1419 GNDA 0.2565
R4478 GNDA GNDA.n2198 0.2565
R4479 GNDA.n948 GNDA 0.2565
R4480 GNDA.n1696 GNDA 0.2565
R4481 GNDA GNDA.n451 0.2565
R4482 GNDA.n680 GNDA 0.2565
R4483 GNDA.n71 GNDA.n60 0.2505
R4484 GNDA.n333 GNDA.n313 0.22375
R4485 GNDA.n334 GNDA.n333 0.100375
R4486 GNDA.n625 GNDA 0.0517
R4487 GNDA.n1252 GNDA 0.0517
R4488 GNDA.n859 GNDA 0.0517
R4489 GNDA.n1419 GNDA 0.0517
R4490 GNDA.n2198 GNDA 0.0517
R4491 GNDA GNDA.n948 0.0517
R4492 GNDA.n1696 GNDA 0.0517
R4493 GNDA.n451 GNDA 0.0517
R4494 GNDA GNDA.n680 0.0517
R4495 VDDA.n382 VDDA.n349 6600
R4496 VDDA.n384 VDDA.n349 6600
R4497 VDDA.n384 VDDA.n350 6570
R4498 VDDA.n382 VDDA.n350 6570
R4499 VDDA.n337 VDDA.n272 4710
R4500 VDDA.n337 VDDA.n273 4710
R4501 VDDA.n339 VDDA.n272 4710
R4502 VDDA.n339 VDDA.n273 4710
R4503 VDDA.n295 VDDA.n294 4710
R4504 VDDA.n297 VDDA.n294 4710
R4505 VDDA.n295 VDDA.n288 4710
R4506 VDDA.n297 VDDA.n288 4710
R4507 VDDA.n143 VDDA.n129 4605
R4508 VDDA.n145 VDDA.n129 4605
R4509 VDDA.n69 VDDA.n65 4605
R4510 VDDA.n69 VDDA.n66 4605
R4511 VDDA.n179 VDDA.n175 4590
R4512 VDDA.n179 VDDA.n176 4590
R4513 VDDA.n181 VDDA.n176 4590
R4514 VDDA.n181 VDDA.n175 4590
R4515 VDDA.n143 VDDA.n130 4575
R4516 VDDA.n145 VDDA.n130 4575
R4517 VDDA.n71 VDDA.n65 4575
R4518 VDDA.n71 VDDA.n66 4575
R4519 VDDA.n205 VDDA.n198 4020
R4520 VDDA.n207 VDDA.n198 4020
R4521 VDDA.n205 VDDA.n204 4020
R4522 VDDA.n207 VDDA.n204 4020
R4523 VDDA.n93 VDDA.n86 4020
R4524 VDDA.n95 VDDA.n86 4020
R4525 VDDA.n93 VDDA.n92 4020
R4526 VDDA.n95 VDDA.n92 4020
R4527 VDDA.n448 VDDA.n416 3420
R4528 VDDA.n448 VDDA.n417 3420
R4529 VDDA.n122 VDDA.n115 3390
R4530 VDDA.n124 VDDA.n115 3390
R4531 VDDA.n122 VDDA.n121 3390
R4532 VDDA.n124 VDDA.n121 3390
R4533 VDDA.n49 VDDA.n42 3390
R4534 VDDA.n51 VDDA.n42 3390
R4535 VDDA.n49 VDDA.n48 3390
R4536 VDDA.n51 VDDA.n48 3390
R4537 VDDA.n23 VDDA.n17 2940
R4538 VDDA.n25 VDDA.n17 2940
R4539 VDDA.n25 VDDA.n22 2940
R4540 VDDA.n23 VDDA.n22 2940
R4541 VDDA.n31 VDDA.n12 2940
R4542 VDDA.n33 VDDA.n12 2940
R4543 VDDA.n33 VDDA.n30 2940
R4544 VDDA.n31 VDDA.n30 2940
R4545 VDDA.n450 VDDA.n416 2760
R4546 VDDA.n450 VDDA.n417 2760
R4547 VDDA.n235 VDDA.n224 2520
R4548 VDDA.n232 VDDA.n225 2505
R4549 VDDA.n235 VDDA.n225 2475
R4550 VDDA.n232 VDDA.n224 2220
R4551 VDDA.n464 VDDA.n410 2145
R4552 VDDA.n464 VDDA.n411 2100
R4553 VDDA.n461 VDDA.n411 2100
R4554 VDDA.n429 VDDA.n422 2100
R4555 VDDA.n431 VDDA.n422 2100
R4556 VDDA.n431 VDDA.n423 2100
R4557 VDDA.n429 VDDA.n423 2100
R4558 VDDA.n461 VDDA.n410 2055
R4559 VDDA.n397 VDDA.n395 1770
R4560 VDDA.n399 VDDA.n395 1770
R4561 VDDA.n397 VDDA.n392 1770
R4562 VDDA.n399 VDDA.n392 1770
R4563 VDDA.n358 VDDA.n356 1770
R4564 VDDA.n360 VDDA.n356 1770
R4565 VDDA.n358 VDDA.n353 1770
R4566 VDDA.n360 VDDA.n353 1770
R4567 VDDA.n247 VDDA.n220 1575
R4568 VDDA.n246 VDDA.n220 1575
R4569 VDDA.n246 VDDA.n219 1545
R4570 VDDA.n247 VDDA.n219 1545
R4571 VDDA.n140 VDDA.t346 1216.42
R4572 VDDA.n148 VDDA.t373 1216.42
R4573 VDDA.n63 VDDA.t352 1216.42
R4574 VDDA.n74 VDDA.t327 1216.42
R4575 VDDA.n381 VDDA.n348 704
R4576 VDDA.n385 VDDA.n348 704
R4577 VDDA.n19 VDDA.t360 689.4
R4578 VDDA.n18 VDDA.t384 689.4
R4579 VDDA.n14 VDDA.t426 689.4
R4580 VDDA.n13 VDDA.t323 689.4
R4581 VDDA.n229 VDDA.t339 666.134
R4582 VDDA.n238 VDDA.t394 666.134
R4583 VDDA.n172 VDDA.t405 663.801
R4584 VDDA.n185 VDDA.t414 663.801
R4585 VDDA.n201 VDDA.t364 660.109
R4586 VDDA.n199 VDDA.t397 660.109
R4587 VDDA.n89 VDDA.t367 660.109
R4588 VDDA.n87 VDDA.t418 660.109
R4589 VDDA.t339 VDDA.n228 658.101
R4590 VDDA.n242 VDDA.t332 650.668
R4591 VDDA.n251 VDDA.t345 650.668
R4592 VDDA.n216 VDDA.n215 632.293
R4593 VDDA.n152 VDDA.n151 626.534
R4594 VDDA.n155 VDDA.n154 626.534
R4595 VDDA.n157 VDDA.n156 626.534
R4596 VDDA.n159 VDDA.n158 626.534
R4597 VDDA.n161 VDDA.n160 626.534
R4598 VDDA.n163 VDDA.n162 626.534
R4599 VDDA.n165 VDDA.n164 626.534
R4600 VDDA.n167 VDDA.n166 626.534
R4601 VDDA.n169 VDDA.n168 626.534
R4602 VDDA.n171 VDDA.n170 626.534
R4603 VDDA.n118 VDDA.t355 573.75
R4604 VDDA.n116 VDDA.t379 573.75
R4605 VDDA.n45 VDDA.t333 573.75
R4606 VDDA.n43 VDDA.t361 573.75
R4607 VDDA.n380 VDDA.n347 518.4
R4608 VDDA.n386 VDDA.n347 518.4
R4609 VDDA.n299 VDDA.n298 496
R4610 VDDA.n299 VDDA.n287 496
R4611 VDDA.n146 VDDA.n128 491.2
R4612 VDDA.n142 VDDA.n128 491.2
R4613 VDDA.n68 VDDA.n40 491.2
R4614 VDDA.n68 VDDA.n67 491.2
R4615 VDDA.n178 VDDA.n153 489.601
R4616 VDDA.n178 VDDA.n177 489.601
R4617 VDDA.n209 VDDA.n208 428.8
R4618 VDDA.n209 VDDA.n197 428.8
R4619 VDDA.n97 VDDA.n96 428.8
R4620 VDDA.n97 VDDA.n85 428.8
R4621 VDDA.n393 VDDA.t385 419.108
R4622 VDDA.n390 VDDA.t388 419.108
R4623 VDDA.n354 VDDA.t430 413.084
R4624 VDDA.n351 VDDA.t400 413.084
R4625 VDDA.n458 VDDA.t349 409.067
R4626 VDDA.n467 VDDA.t421 409.067
R4627 VDDA.n445 VDDA.t427 409.067
R4628 VDDA.n453 VDDA.t409 409.067
R4629 VDDA.n426 VDDA.t415 409.067
R4630 VDDA.n434 VDDA.t324 390.322
R4631 VDDA.t413 VDDA.n175 389.375
R4632 VDDA.t404 VDDA.n176 389.375
R4633 VDDA.t425 VDDA.n30 389.375
R4634 VDDA.t322 VDDA.n12 389.375
R4635 VDDA.n393 VDDA.t387 389.185
R4636 VDDA.n390 VDDA.t390 389.185
R4637 VDDA.n183 VDDA.n182 387.2
R4638 VDDA.n182 VDDA.n174 387.2
R4639 VDDA.n445 VDDA.t429 387.051
R4640 VDDA.n453 VDDA.t411 387.051
R4641 VDDA.n270 VDDA.t393 384.918
R4642 VDDA.n274 VDDA.t408 384.918
R4643 VDDA.n289 VDDA.t378 384.918
R4644 VDDA.n291 VDDA.t338 384.918
R4645 VDDA.n354 VDDA.t432 384.918
R4646 VDDA.n351 VDDA.t402 384.918
R4647 VDDA.t359 VDDA.n22 384.168
R4648 VDDA.t383 VDDA.n17 384.168
R4649 VDDA.n276 VDDA.n275 384
R4650 VDDA.n275 VDDA.n271 384
R4651 VDDA.n293 VDDA.n292 384
R4652 VDDA.n293 VDDA.n290 384
R4653 VDDA.n426 VDDA.t417 370.728
R4654 VDDA.n434 VDDA.t326 370.728
R4655 VDDA.n458 VDDA.t351 370.3
R4656 VDDA.n467 VDDA.t423 370.3
R4657 VDDA.n447 VDDA.n415 364.8
R4658 VDDA.n379 VDDA.t370 360.868
R4659 VDDA.n387 VDDA.t318 360.868
R4660 VDDA.n270 VDDA.t391 358.858
R4661 VDDA.n274 VDDA.t406 358.858
R4662 VDDA.n289 VDDA.t376 358.858
R4663 VDDA.n291 VDDA.t336 358.858
R4664 VDDA.n126 VDDA.n125 355.2
R4665 VDDA.n126 VDDA.n114 355.2
R4666 VDDA.n53 VDDA.n52 355.2
R4667 VDDA.n53 VDDA.n41 355.2
R4668 VDDA.t407 VDDA.n337 351.591
R4669 VDDA.n339 VDDA.t392 351.591
R4670 VDDA.t337 VDDA.n295 351.591
R4671 VDDA.n297 VDDA.t377 351.591
R4672 VDDA.t331 VDDA.n246 346.668
R4673 VDDA.n247 VDDA.t343 346.668
R4674 VDDA.n419 VDDA.n418 345.127
R4675 VDDA.n425 VDDA.n424 345.127
R4676 VDDA.n407 VDDA.n406 344.7
R4677 VDDA.n456 VDDA.n455 344.7
R4678 VDDA.t389 VDDA.n397 344.394
R4679 VDDA.n399 VDDA.t386 344.394
R4680 VDDA.t401 VDDA.n358 344.394
R4681 VDDA.n360 VDDA.t431 344.394
R4682 VDDA.t350 VDDA.n461 344.394
R4683 VDDA.n464 VDDA.t422 344.394
R4684 VDDA.n281 VDDA.n279 342.3
R4685 VDDA.n309 VDDA.n308 341.675
R4686 VDDA.n307 VDDA.n306 341.675
R4687 VDDA.n305 VDDA.n304 341.675
R4688 VDDA.n303 VDDA.n302 341.675
R4689 VDDA.n285 VDDA.n284 341.675
R4690 VDDA.n283 VDDA.n282 341.675
R4691 VDDA.n281 VDDA.n280 341.675
R4692 VDDA.t428 VDDA.n448 340.635
R4693 VDDA.n450 VDDA.t410 340.635
R4694 VDDA.t416 VDDA.n429 340.635
R4695 VDDA.n431 VDDA.t325 340.635
R4696 VDDA.n413 VDDA.n412 339.272
R4697 VDDA.n437 VDDA.n436 339.272
R4698 VDDA.n439 VDDA.n438 339.272
R4699 VDDA.n441 VDDA.n440 339.272
R4700 VDDA.n443 VDDA.n442 339.272
R4701 VDDA.n342 VDDA.n266 337.175
R4702 VDDA.n268 VDDA.n267 337.175
R4703 VDDA.n318 VDDA.n317 337.175
R4704 VDDA.n321 VDDA.n315 337.175
R4705 VDDA.n313 VDDA.n312 337.175
R4706 VDDA.n325 VDDA.n324 337.175
R4707 VDDA.n328 VDDA.n311 337.175
R4708 VDDA.n331 VDDA.n330 337.175
R4709 VDDA.n334 VDDA.n278 337.175
R4710 VDDA.n300 VDDA.n286 337.175
R4711 VDDA.n403 VDDA.n389 335.022
R4712 VDDA.n173 VDDA.t403 332.75
R4713 VDDA.n184 VDDA.t412 332.75
R4714 VDDA.n19 VDDA.t358 332.75
R4715 VDDA.n18 VDDA.t382 332.75
R4716 VDDA.n14 VDDA.t424 332.75
R4717 VDDA.n13 VDDA.t321 332.75
R4718 VDDA.n21 VDDA.n16 313.601
R4719 VDDA.n243 VDDA.t330 310.659
R4720 VDDA.n250 VDDA.t342 310.659
R4721 VDDA.n28 VDDA.n16 307.2
R4722 VDDA.n36 VDDA.n11 307.2
R4723 VDDA.n29 VDDA.n11 307.2
R4724 VDDA.n451 VDDA.n415 294.401
R4725 VDDA.t356 VDDA.n122 285.815
R4726 VDDA.n124 VDDA.t380 285.815
R4727 VDDA.t334 VDDA.n49 285.815
R4728 VDDA.n51 VDDA.t362 285.815
R4729 VDDA.t371 VDDA.n382 278.95
R4730 VDDA.n384 VDDA.t319 278.95
R4731 VDDA.n118 VDDA.t357 277.916
R4732 VDDA.n116 VDDA.t381 277.916
R4733 VDDA.n45 VDDA.t335 277.916
R4734 VDDA.n43 VDDA.t363 277.916
R4735 VDDA.n147 VDDA.n146 276.8
R4736 VDDA.n142 VDDA.n141 276.8
R4737 VDDA.n73 VDDA.n40 276.8
R4738 VDDA.n67 VDDA.n64 276.8
R4739 VDDA.n379 VDDA.t372 270.705
R4740 VDDA.n387 VDDA.t320 270.705
R4741 VDDA.n236 VDDA.n223 268.8
R4742 VDDA.n446 VDDA.n414 246.4
R4743 VDDA.t365 VDDA.n205 239.915
R4744 VDDA.n207 VDDA.t398 239.915
R4745 VDDA.t368 VDDA.n93 239.915
R4746 VDDA.n95 VDDA.t419 239.915
R4747 VDDA.n231 VDDA.n223 236.8
R4748 VDDA.n203 VDDA.n202 230.4
R4749 VDDA.n203 VDDA.n200 230.4
R4750 VDDA.n91 VDDA.n90 230.4
R4751 VDDA.n91 VDDA.n88 230.4
R4752 VDDA.n465 VDDA.n409 228.8
R4753 VDDA.n428 VDDA.n421 224
R4754 VDDA.n432 VDDA.n421 224
R4755 VDDA.n460 VDDA.n409 219.201
R4756 VDDA.n231 VDDA.n230 216
R4757 VDDA.n120 VDDA.n119 211.201
R4758 VDDA.n120 VDDA.n117 211.201
R4759 VDDA.n47 VDDA.n46 211.201
R4760 VDDA.n47 VDDA.n44 211.201
R4761 VDDA.n26 VDDA.n20 211.201
R4762 VDDA.n27 VDDA.n26 211.201
R4763 VDDA.n35 VDDA.n34 211.201
R4764 VDDA.n141 VDDA.n127 204.8
R4765 VDDA.n147 VDDA.n127 204.8
R4766 VDDA.n73 VDDA.n72 204.8
R4767 VDDA.n72 VDDA.n64 204.8
R4768 VDDA.n34 VDDA.n15 202.971
R4769 VDDA.n237 VDDA.n236 200
R4770 VDDA.n208 VDDA.n200 198.4
R4771 VDDA.n202 VDDA.n197 198.4
R4772 VDDA.n96 VDDA.n88 198.4
R4773 VDDA.n90 VDDA.n85 198.4
R4774 VDDA.t115 VDDA.t331 190
R4775 VDDA.t343 VDDA.t115 190
R4776 VDDA.n341 VDDA.n340 188.8
R4777 VDDA.n336 VDDA.n335 188.8
R4778 VDDA.n400 VDDA.n394 188.8
R4779 VDDA.n396 VDDA.n394 188.8
R4780 VDDA.n361 VDDA.n355 188.8
R4781 VDDA.n357 VDDA.n355 188.8
R4782 VDDA.t40 VDDA.t413 186.607
R4783 VDDA.t105 VDDA.t40 186.607
R4784 VDDA.t175 VDDA.t105 186.607
R4785 VDDA.t103 VDDA.t175 186.607
R4786 VDDA.t169 VDDA.t103 186.607
R4787 VDDA.t179 VDDA.t169 186.607
R4788 VDDA.t62 VDDA.t179 186.607
R4789 VDDA.t185 VDDA.t62 186.607
R4790 VDDA.t14 VDDA.t185 186.607
R4791 VDDA.t49 VDDA.t14 186.607
R4792 VDDA.t101 VDDA.t173 186.607
R4793 VDDA.t173 VDDA.t16 186.607
R4794 VDDA.t16 VDDA.t42 186.607
R4795 VDDA.t42 VDDA.t177 186.607
R4796 VDDA.t177 VDDA.t171 186.607
R4797 VDDA.t171 VDDA.t183 186.607
R4798 VDDA.t183 VDDA.t181 186.607
R4799 VDDA.t181 VDDA.t47 186.607
R4800 VDDA.t47 VDDA.t99 186.607
R4801 VDDA.t99 VDDA.t404 186.607
R4802 VDDA.t146 VDDA.t425 186.607
R4803 VDDA.t112 VDDA.t146 186.607
R4804 VDDA.t433 VDDA.t112 186.607
R4805 VDDA.t119 VDDA.t433 186.607
R4806 VDDA.t122 VDDA.t119 186.607
R4807 VDDA.t251 VDDA.t34 186.607
R4808 VDDA.t34 VDDA.t148 186.607
R4809 VDDA.t148 VDDA.t118 186.607
R4810 VDDA.t118 VDDA.t450 186.607
R4811 VDDA.t450 VDDA.t322 186.607
R4812 VDDA.t147 VDDA.t359 183.333
R4813 VDDA.t68 VDDA.t147 183.333
R4814 VDDA.t13 VDDA.t68 183.333
R4815 VDDA.t117 VDDA.t13 183.333
R4816 VDDA.t121 VDDA.t117 183.333
R4817 VDDA.t35 VDDA.t197 183.333
R4818 VDDA.t197 VDDA.t455 183.333
R4819 VDDA.t455 VDDA.t120 183.333
R4820 VDDA.t120 VDDA.t33 183.333
R4821 VDDA.t33 VDDA.t383 183.333
R4822 VDDA.n381 VDDA.n380 182.4
R4823 VDDA.n386 VDDA.n385 182.4
R4824 VDDA.n139 VDDA.t348 178.124
R4825 VDDA.n149 VDDA.t375 178.124
R4826 VDDA.n62 VDDA.t354 178.124
R4827 VDDA.n75 VDDA.t329 178.124
R4828 VDDA.n452 VDDA.n414 176
R4829 VDDA.n226 VDDA.n221 173.733
R4830 VDDA.t200 VDDA.t407 172.727
R4831 VDDA.t38 VDDA.t200 172.727
R4832 VDDA.t236 VDDA.t38 172.727
R4833 VDDA.t69 VDDA.t236 172.727
R4834 VDDA.t11 VDDA.t69 172.727
R4835 VDDA.t191 VDDA.t11 172.727
R4836 VDDA.t459 VDDA.t191 172.727
R4837 VDDA.t434 VDDA.t459 172.727
R4838 VDDA.t154 VDDA.t434 172.727
R4839 VDDA.t84 VDDA.t198 172.727
R4840 VDDA.t27 VDDA.t84 172.727
R4841 VDDA.t225 VDDA.t27 172.727
R4842 VDDA.t73 VDDA.t225 172.727
R4843 VDDA.t97 VDDA.t73 172.727
R4844 VDDA.t9 VDDA.t97 172.727
R4845 VDDA.t249 VDDA.t9 172.727
R4846 VDDA.t66 VDDA.t249 172.727
R4847 VDDA.t392 VDDA.t66 172.727
R4848 VDDA.t256 VDDA.t337 172.727
R4849 VDDA.t64 VDDA.t256 172.727
R4850 VDDA.t60 VDDA.t64 172.727
R4851 VDDA.t260 VDDA.t60 172.727
R4852 VDDA.t268 VDDA.t260 172.727
R4853 VDDA.t252 VDDA.t268 172.727
R4854 VDDA.t157 VDDA.t252 172.727
R4855 VDDA.t36 VDDA.t157 172.727
R4856 VDDA.t21 VDDA.t36 172.727
R4857 VDDA.t264 VDDA.t270 172.727
R4858 VDDA.t254 VDDA.t264 172.727
R4859 VDDA.t258 VDDA.t254 172.727
R4860 VDDA.t442 VDDA.t258 172.727
R4861 VDDA.t436 VDDA.t442 172.727
R4862 VDDA.t266 VDDA.t436 172.727
R4863 VDDA.t262 VDDA.t266 172.727
R4864 VDDA.t82 VDDA.t262 172.727
R4865 VDDA.t377 VDDA.t82 172.727
R4866 VDDA.n346 VDDA.n345 168.435
R4867 VDDA.n365 VDDA.n364 168.435
R4868 VDDA.n367 VDDA.n366 168.435
R4869 VDDA.n369 VDDA.n368 168.435
R4870 VDDA.n371 VDDA.n370 168.435
R4871 VDDA.n373 VDDA.n372 168.435
R4872 VDDA.n375 VDDA.n374 168.435
R4873 VDDA.n377 VDDA.n376 168.435
R4874 VDDA.n245 VDDA.n218 164.8
R4875 VDDA.n248 VDDA.n218 164.8
R4876 VDDA.t347 VDDA.n143 161.817
R4877 VDDA.n145 VDDA.t374 161.817
R4878 VDDA.t328 VDDA.n65 161.817
R4879 VDDA.t353 VDDA.n66 161.817
R4880 VDDA.n235 VDDA.t395 161.733
R4881 VDDA.n195 VDDA.n193 160.428
R4882 VDDA.n192 VDDA.n190 160.428
R4883 VDDA.n83 VDDA.n81 160.428
R4884 VDDA.n80 VDDA.n78 160.428
R4885 VDDA.t167 VDDA.t371 159.814
R4886 VDDA.t137 VDDA.t167 159.814
R4887 VDDA.t75 VDDA.t137 159.814
R4888 VDDA.t208 VDDA.t75 159.814
R4889 VDDA.t129 VDDA.t208 159.814
R4890 VDDA.t144 VDDA.t129 159.814
R4891 VDDA.t163 VDDA.t144 159.814
R4892 VDDA.t467 VDDA.t163 159.814
R4893 VDDA.t165 VDDA.t131 159.814
R4894 VDDA.t107 VDDA.t165 159.814
R4895 VDDA.t109 VDDA.t107 159.814
R4896 VDDA.t461 VDDA.t109 159.814
R4897 VDDA.t133 VDDA.t461 159.814
R4898 VDDA.t141 VDDA.t133 159.814
R4899 VDDA.t89 VDDA.t141 159.814
R4900 VDDA.t319 VDDA.t89 159.814
R4901 VDDA.n195 VDDA.n194 159.803
R4902 VDDA.n192 VDDA.n191 159.803
R4903 VDDA.n83 VDDA.n82 159.803
R4904 VDDA.n80 VDDA.n79 159.803
R4905 VDDA.t340 VDDA.n232 159.147
R4906 VDDA.t446 VDDA.t389 158.333
R4907 VDDA.t386 VDDA.t31 158.333
R4908 VDDA.t248 VDDA.t401 158.333
R4909 VDDA.t431 VDDA.t227 158.333
R4910 VDDA.t246 VDDA.t350 158.333
R4911 VDDA.t211 VDDA.t246 158.333
R4912 VDDA.t223 VDDA.t161 158.333
R4913 VDDA.t422 VDDA.t223 158.333
R4914 VDDA.t440 VDDA.t428 155.97
R4915 VDDA.t219 VDDA.t440 155.97
R4916 VDDA.t213 VDDA.t219 155.97
R4917 VDDA.t92 VDDA.t213 155.97
R4918 VDDA.t29 VDDA.t92 155.97
R4919 VDDA.t195 VDDA.t29 155.97
R4920 VDDA.t193 VDDA.t221 155.97
R4921 VDDA.t457 VDDA.t193 155.97
R4922 VDDA.t152 VDDA.t457 155.97
R4923 VDDA.t410 VDDA.t152 155.97
R4924 VDDA.t244 VDDA.t416 155.97
R4925 VDDA.t453 VDDA.t244 155.97
R4926 VDDA.t448 VDDA.t1 155.97
R4927 VDDA.t325 VDDA.t448 155.97
R4928 VDDA.n201 VDDA.t366 155.125
R4929 VDDA.n199 VDDA.t399 155.125
R4930 VDDA.n89 VDDA.t369 155.125
R4931 VDDA.n87 VDDA.t420 155.125
R4932 VDDA.n139 VDDA.n138 151.882
R4933 VDDA.n62 VDDA.n61 151.882
R4934 VDDA.n150 VDDA.n149 151.321
R4935 VDDA.n76 VDDA.n75 151.321
R4936 VDDA.n125 VDDA.n117 150.4
R4937 VDDA.n119 VDDA.n114 150.4
R4938 VDDA.n52 VDDA.n44 150.4
R4939 VDDA.n46 VDDA.n41 150.4
R4940 VDDA.n211 VDDA.n210 146.002
R4941 VDDA.n99 VDDA.n98 146.002
R4942 VDDA.n113 VDDA.n112 145.429
R4943 VDDA.n132 VDDA.n131 145.429
R4944 VDDA.n134 VDDA.n133 145.429
R4945 VDDA.n136 VDDA.n135 145.429
R4946 VDDA.n138 VDDA.n137 145.429
R4947 VDDA.n39 VDDA.n38 145.429
R4948 VDDA.n55 VDDA.n54 145.429
R4949 VDDA.n57 VDDA.n56 145.429
R4950 VDDA.n59 VDDA.n58 145.429
R4951 VDDA.n61 VDDA.n60 145.429
R4952 VDDA.n149 VDDA.n148 135.387
R4953 VDDA.n140 VDDA.n139 135.387
R4954 VDDA.n75 VDDA.n74 135.387
R4955 VDDA.n63 VDDA.n62 135.387
R4956 VDDA.t156 VDDA.t356 121.513
R4957 VDDA.t0 VDDA.t156 121.513
R4958 VDDA.t444 VDDA.t0 121.513
R4959 VDDA.t26 VDDA.t444 121.513
R4960 VDDA.t230 VDDA.t26 121.513
R4961 VDDA.t242 VDDA.t206 121.513
R4962 VDDA.t190 VDDA.t242 121.513
R4963 VDDA.t445 VDDA.t190 121.513
R4964 VDDA.t187 VDDA.t445 121.513
R4965 VDDA.t380 VDDA.t187 121.513
R4966 VDDA.t238 VDDA.t334 121.513
R4967 VDDA.t18 VDDA.t238 121.513
R4968 VDDA.t216 VDDA.t18 121.513
R4969 VDDA.t96 VDDA.t216 121.513
R4970 VDDA.t149 VDDA.t96 121.513
R4971 VDDA.t56 VDDA.t127 121.513
R4972 VDDA.t125 VDDA.t56 121.513
R4973 VDDA.t114 VDDA.t125 121.513
R4974 VDDA.t95 VDDA.t114 121.513
R4975 VDDA.t362 VDDA.t95 121.513
R4976 VDDA.n340 VDDA.n271 118.4
R4977 VDDA.n336 VDDA.n276 118.4
R4978 VDDA.n298 VDDA.n290 118.4
R4979 VDDA.n292 VDDA.n287 118.4
R4980 VDDA.n401 VDDA.n400 118.4
R4981 VDDA.n396 VDDA.n391 118.4
R4982 VDDA.n362 VDDA.n361 118.4
R4983 VDDA.n357 VDDA.n352 118.4
R4984 VDDA.n460 VDDA.n459 118.4
R4985 VDDA.n466 VDDA.n465 118.4
R4986 VDDA.n447 VDDA.n446 118.4
R4987 VDDA.n452 VDDA.n451 118.4
R4988 VDDA.n428 VDDA.n427 118.4
R4989 VDDA.n433 VDDA.n432 118.4
R4990 VDDA.n245 VDDA.n244 110.4
R4991 VDDA.n249 VDDA.n248 110.4
R4992 VDDA.n240 VDDA.n239 108.734
R4993 VDDA.n459 VDDA.n408 105.6
R4994 VDDA.n466 VDDA.n408 105.6
R4995 VDDA.n427 VDDA.n420 105.6
R4996 VDDA.n433 VDDA.n420 105.6
R4997 VDDA.n183 VDDA.n153 102.4
R4998 VDDA.n177 VDDA.n174 102.4
R4999 VDDA.n21 VDDA.n20 102.4
R5000 VDDA.t278 VDDA.t365 98.2764
R5001 VDDA.t284 VDDA.t278 98.2764
R5002 VDDA.t290 VDDA.t284 98.2764
R5003 VDDA.t300 VDDA.t290 98.2764
R5004 VDDA.t310 VDDA.t300 98.2764
R5005 VDDA.t280 VDDA.t274 98.2764
R5006 VDDA.t286 VDDA.t280 98.2764
R5007 VDDA.t292 VDDA.t286 98.2764
R5008 VDDA.t304 VDDA.t292 98.2764
R5009 VDDA.t398 VDDA.t304 98.2764
R5010 VDDA.t288 VDDA.t368 98.2764
R5011 VDDA.t296 VDDA.t288 98.2764
R5012 VDDA.t308 VDDA.t296 98.2764
R5013 VDDA.t302 VDDA.t308 98.2764
R5014 VDDA.t312 VDDA.t302 98.2764
R5015 VDDA.t276 VDDA.t272 98.2764
R5016 VDDA.t298 VDDA.t276 98.2764
R5017 VDDA.t294 VDDA.t298 98.2764
R5018 VDDA.t306 VDDA.t294 98.2764
R5019 VDDA.t419 VDDA.t306 98.2764
R5020 VDDA.n103 VDDA.n101 97.4034
R5021 VDDA.n2 VDDA.n0 97.4034
R5022 VDDA.n111 VDDA.n110 96.8409
R5023 VDDA.n109 VDDA.n108 96.8409
R5024 VDDA.n107 VDDA.n106 96.8409
R5025 VDDA.n105 VDDA.n104 96.8409
R5026 VDDA.n103 VDDA.n102 96.8409
R5027 VDDA.n10 VDDA.n9 96.8409
R5028 VDDA.n8 VDDA.n7 96.8409
R5029 VDDA.n6 VDDA.n5 96.8409
R5030 VDDA.n4 VDDA.n3 96.8409
R5031 VDDA.n2 VDDA.n1 96.8409
R5032 VDDA.t395 VDDA.t282 96.6107
R5033 VDDA.n28 VDDA.n27 96.0005
R5034 VDDA.n29 VDDA.n15 96.0005
R5035 VDDA.n36 VDDA.n35 96.0005
R5036 VDDA.n228 VDDA.n227 94.9338
R5037 VDDA.n180 VDDA.t49 93.3041
R5038 VDDA.n180 VDDA.t101 93.3041
R5039 VDDA.n32 VDDA.t122 93.3041
R5040 VDDA.n32 VDDA.t251 93.3041
R5041 VDDA.n219 VDDA.n218 92.5005
R5042 VDDA.t115 VDDA.n219 92.5005
R5043 VDDA.n220 VDDA.n217 92.5005
R5044 VDDA.t115 VDDA.n220 92.5005
R5045 VDDA.n224 VDDA.n223 92.5005
R5046 VDDA.n233 VDDA.n224 92.5005
R5047 VDDA.n225 VDDA.n222 92.5005
R5048 VDDA.n234 VDDA.n225 92.5005
R5049 VDDA.n208 VDDA.n207 92.5005
R5050 VDDA.n204 VDDA.n203 92.5005
R5051 VDDA.n206 VDDA.n204 92.5005
R5052 VDDA.n205 VDDA.n197 92.5005
R5053 VDDA.n209 VDDA.n198 92.5005
R5054 VDDA.n206 VDDA.n198 92.5005
R5055 VDDA.n175 VDDA.n153 92.5005
R5056 VDDA.n179 VDDA.n178 92.5005
R5057 VDDA.n180 VDDA.n179 92.5005
R5058 VDDA.n177 VDDA.n176 92.5005
R5059 VDDA.n182 VDDA.n181 92.5005
R5060 VDDA.n181 VDDA.n180 92.5005
R5061 VDDA.n125 VDDA.n124 92.5005
R5062 VDDA.n121 VDDA.n120 92.5005
R5063 VDDA.n123 VDDA.n121 92.5005
R5064 VDDA.n122 VDDA.n114 92.5005
R5065 VDDA.n126 VDDA.n115 92.5005
R5066 VDDA.n123 VDDA.n115 92.5005
R5067 VDDA.n130 VDDA.n127 92.5005
R5068 VDDA.n144 VDDA.n130 92.5005
R5069 VDDA.n129 VDDA.n128 92.5005
R5070 VDDA.n144 VDDA.n129 92.5005
R5071 VDDA.n96 VDDA.n95 92.5005
R5072 VDDA.n92 VDDA.n91 92.5005
R5073 VDDA.n94 VDDA.n92 92.5005
R5074 VDDA.n93 VDDA.n85 92.5005
R5075 VDDA.n97 VDDA.n86 92.5005
R5076 VDDA.n94 VDDA.n86 92.5005
R5077 VDDA.n52 VDDA.n51 92.5005
R5078 VDDA.n48 VDDA.n47 92.5005
R5079 VDDA.n50 VDDA.n48 92.5005
R5080 VDDA.n49 VDDA.n41 92.5005
R5081 VDDA.n53 VDDA.n42 92.5005
R5082 VDDA.n50 VDDA.n42 92.5005
R5083 VDDA.n72 VDDA.n71 92.5005
R5084 VDDA.n71 VDDA.n70 92.5005
R5085 VDDA.n69 VDDA.n68 92.5005
R5086 VDDA.n70 VDDA.n69 92.5005
R5087 VDDA.n23 VDDA.n16 92.5005
R5088 VDDA.n24 VDDA.n23 92.5005
R5089 VDDA.n22 VDDA.n21 92.5005
R5090 VDDA.n26 VDDA.n25 92.5005
R5091 VDDA.n25 VDDA.n24 92.5005
R5092 VDDA.n28 VDDA.n17 92.5005
R5093 VDDA.n31 VDDA.n11 92.5005
R5094 VDDA.n32 VDDA.n31 92.5005
R5095 VDDA.n30 VDDA.n29 92.5005
R5096 VDDA.n34 VDDA.n33 92.5005
R5097 VDDA.n33 VDDA.n32 92.5005
R5098 VDDA.n36 VDDA.n12 92.5005
R5099 VDDA.n323 VDDA.n273 92.5005
R5100 VDDA.n338 VDDA.n273 92.5005
R5101 VDDA.n340 VDDA.n339 92.5005
R5102 VDDA.n275 VDDA.n272 92.5005
R5103 VDDA.n338 VDDA.n272 92.5005
R5104 VDDA.n337 VDDA.n336 92.5005
R5105 VDDA.n298 VDDA.n297 92.5005
R5106 VDDA.n294 VDDA.n293 92.5005
R5107 VDDA.n296 VDDA.n294 92.5005
R5108 VDDA.n295 VDDA.n287 92.5005
R5109 VDDA.n299 VDDA.n288 92.5005
R5110 VDDA.n296 VDDA.n288 92.5005
R5111 VDDA.n400 VDDA.n399 92.5005
R5112 VDDA.n395 VDDA.n394 92.5005
R5113 VDDA.n398 VDDA.n395 92.5005
R5114 VDDA.n397 VDDA.n396 92.5005
R5115 VDDA.n402 VDDA.n392 92.5005
R5116 VDDA.n398 VDDA.n392 92.5005
R5117 VDDA.n382 VDDA.n381 92.5005
R5118 VDDA.n349 VDDA.n348 92.5005
R5119 VDDA.n383 VDDA.n349 92.5005
R5120 VDDA.n385 VDDA.n384 92.5005
R5121 VDDA.n350 VDDA.n347 92.5005
R5122 VDDA.n383 VDDA.n350 92.5005
R5123 VDDA.n361 VDDA.n360 92.5005
R5124 VDDA.n356 VDDA.n355 92.5005
R5125 VDDA.n359 VDDA.n356 92.5005
R5126 VDDA.n358 VDDA.n357 92.5005
R5127 VDDA.n363 VDDA.n353 92.5005
R5128 VDDA.n359 VDDA.n353 92.5005
R5129 VDDA.n461 VDDA.n460 92.5005
R5130 VDDA.n410 VDDA.n409 92.5005
R5131 VDDA.n462 VDDA.n410 92.5005
R5132 VDDA.n465 VDDA.n464 92.5005
R5133 VDDA.n411 VDDA.n408 92.5005
R5134 VDDA.n463 VDDA.n411 92.5005
R5135 VDDA.n448 VDDA.n447 92.5005
R5136 VDDA.n416 VDDA.n415 92.5005
R5137 VDDA.n449 VDDA.n416 92.5005
R5138 VDDA.n451 VDDA.n450 92.5005
R5139 VDDA.n417 VDDA.n414 92.5005
R5140 VDDA.n449 VDDA.n417 92.5005
R5141 VDDA.n429 VDDA.n428 92.5005
R5142 VDDA.n422 VDDA.n421 92.5005
R5143 VDDA.n430 VDDA.n422 92.5005
R5144 VDDA.n432 VDDA.n431 92.5005
R5145 VDDA.n423 VDDA.n420 92.5005
R5146 VDDA.n430 VDDA.n423 92.5005
R5147 VDDA.n24 VDDA.t121 91.6672
R5148 VDDA.n24 VDDA.t35 91.6672
R5149 VDDA.n239 VDDA.n238 88.5338
R5150 VDDA.n229 VDDA.n227 88.5338
R5151 VDDA.n338 VDDA.t154 86.3641
R5152 VDDA.t198 VDDA.n338 86.3641
R5153 VDDA.n296 VDDA.t21 86.3641
R5154 VDDA.t270 VDDA.n296 86.3641
R5155 VDDA.n383 VDDA.t467 79.907
R5156 VDDA.t131 VDDA.n383 79.907
R5157 VDDA.n398 VDDA.t446 79.1672
R5158 VDDA.t31 VDDA.n398 79.1672
R5159 VDDA.n359 VDDA.t248 79.1672
R5160 VDDA.t227 VDDA.n359 79.1672
R5161 VDDA.t161 VDDA.n463 79.1672
R5162 VDDA.n151 VDDA.t41 78.8005
R5163 VDDA.n151 VDDA.t106 78.8005
R5164 VDDA.n154 VDDA.t176 78.8005
R5165 VDDA.n154 VDDA.t104 78.8005
R5166 VDDA.n156 VDDA.t170 78.8005
R5167 VDDA.n156 VDDA.t180 78.8005
R5168 VDDA.n158 VDDA.t63 78.8005
R5169 VDDA.n158 VDDA.t186 78.8005
R5170 VDDA.n160 VDDA.t15 78.8005
R5171 VDDA.n160 VDDA.t50 78.8005
R5172 VDDA.n162 VDDA.t102 78.8005
R5173 VDDA.n162 VDDA.t174 78.8005
R5174 VDDA.n164 VDDA.t17 78.8005
R5175 VDDA.n164 VDDA.t43 78.8005
R5176 VDDA.n166 VDDA.t178 78.8005
R5177 VDDA.n166 VDDA.t172 78.8005
R5178 VDDA.n168 VDDA.t184 78.8005
R5179 VDDA.n168 VDDA.t182 78.8005
R5180 VDDA.n170 VDDA.t48 78.8005
R5181 VDDA.n170 VDDA.t100 78.8005
R5182 VDDA.n449 VDDA.t195 77.9856
R5183 VDDA.t221 VDDA.n449 77.9856
R5184 VDDA.n430 VDDA.t453 77.9856
R5185 VDDA.t1 VDDA.n430 77.9856
R5186 VDDA.n233 VDDA.t340 76.4836
R5187 VDDA.n227 VDDA.t341 76.0991
R5188 VDDA.n239 VDDA.t396 76.0991
R5189 VDDA.n215 VDDA.t116 65.6672
R5190 VDDA.n215 VDDA.t344 65.6672
R5191 VDDA.n237 VDDA.n222 64.0005
R5192 VDDA.n335 VDDA.n277 64.0005
R5193 VDDA.n327 VDDA.n277 64.0005
R5194 VDDA.n327 VDDA.n326 64.0005
R5195 VDDA.n326 VDDA.n323 64.0005
R5196 VDDA.n323 VDDA.n322 64.0005
R5197 VDDA.n322 VDDA.n314 64.0005
R5198 VDDA.n314 VDDA.n269 64.0005
R5199 VDDA.n341 VDDA.n269 64.0005
R5200 VDDA.n363 VDDA.n362 64.0005
R5201 VDDA.n363 VDDA.n352 64.0005
R5202 VDDA.t451 VDDA.t347 62.9523
R5203 VDDA.t232 VDDA.t451 62.9523
R5204 VDDA.t159 VDDA.t232 62.9523
R5205 VDDA.t234 VDDA.t159 62.9523
R5206 VDDA.t188 VDDA.t234 62.9523
R5207 VDDA.t204 VDDA.t228 62.9523
R5208 VDDA.t23 VDDA.t204 62.9523
R5209 VDDA.t465 VDDA.t23 62.9523
R5210 VDDA.t202 VDDA.t465 62.9523
R5211 VDDA.t374 VDDA.t202 62.9523
R5212 VDDA.t79 VDDA.t328 62.9523
R5213 VDDA.t19 VDDA.t79 62.9523
R5214 VDDA.t217 VDDA.t19 62.9523
R5215 VDDA.t57 VDDA.t217 62.9523
R5216 VDDA.t54 VDDA.t57 62.9523
R5217 VDDA.t123 VDDA.t4 62.9523
R5218 VDDA.t4 VDDA.t6 62.9523
R5219 VDDA.t6 VDDA.t239 62.9523
R5220 VDDA.t239 VDDA.t150 62.9523
R5221 VDDA.t150 VDDA.t353 62.9523
R5222 VDDA.n402 VDDA.n401 62.7205
R5223 VDDA.n402 VDDA.n391 62.7205
R5224 VDDA.n246 VDDA.n245 61.6672
R5225 VDDA.n248 VDDA.n247 61.6672
R5226 VDDA.n146 VDDA.n145 61.6672
R5227 VDDA.n143 VDDA.n142 61.6672
R5228 VDDA.n65 VDDA.n40 61.6672
R5229 VDDA.n67 VDDA.n66 61.6672
R5230 VDDA.n123 VDDA.t230 60.7563
R5231 VDDA.t206 VDDA.n123 60.7563
R5232 VDDA.n50 VDDA.t149 60.7563
R5233 VDDA.t127 VDDA.n50 60.7563
R5234 VDDA.n262 VDDA.t470 59.5681
R5235 VDDA.n261 VDDA.t471 59.5681
R5236 VDDA.n244 VDDA.n217 57.6005
R5237 VDDA.n249 VDDA.n217 57.6005
R5238 VDDA.n462 VDDA.t211 57.5763
R5239 VDDA.n261 VDDA.t472 51.8888
R5240 VDDA.n230 VDDA.n222 51.2005
R5241 VDDA.n206 VDDA.t310 49.1384
R5242 VDDA.t274 VDDA.n206 49.1384
R5243 VDDA.n94 VDDA.t312 49.1384
R5244 VDDA.t272 VDDA.n94 49.1384
R5245 VDDA.n263 VDDA.t469 48.9557
R5246 VDDA.n252 VDDA.n251 47.2938
R5247 VDDA.n242 VDDA.n241 42.7938
R5248 VDDA.n172 VDDA.n171 42.0963
R5249 VDDA.n186 VDDA.n185 41.5338
R5250 VDDA.n266 VDDA.t250 39.4005
R5251 VDDA.n266 VDDA.t67 39.4005
R5252 VDDA.n267 VDDA.t98 39.4005
R5253 VDDA.n267 VDDA.t10 39.4005
R5254 VDDA.n317 VDDA.t226 39.4005
R5255 VDDA.n317 VDDA.t74 39.4005
R5256 VDDA.n315 VDDA.t85 39.4005
R5257 VDDA.n315 VDDA.t28 39.4005
R5258 VDDA.n312 VDDA.t155 39.4005
R5259 VDDA.n312 VDDA.t199 39.4005
R5260 VDDA.n324 VDDA.t460 39.4005
R5261 VDDA.n324 VDDA.t435 39.4005
R5262 VDDA.n311 VDDA.t12 39.4005
R5263 VDDA.n311 VDDA.t192 39.4005
R5264 VDDA.n330 VDDA.t237 39.4005
R5265 VDDA.n330 VDDA.t70 39.4005
R5266 VDDA.n278 VDDA.t201 39.4005
R5267 VDDA.n278 VDDA.t39 39.4005
R5268 VDDA.n308 VDDA.t263 39.4005
R5269 VDDA.n308 VDDA.t83 39.4005
R5270 VDDA.n306 VDDA.t437 39.4005
R5271 VDDA.n306 VDDA.t267 39.4005
R5272 VDDA.n304 VDDA.t259 39.4005
R5273 VDDA.n304 VDDA.t443 39.4005
R5274 VDDA.n302 VDDA.t265 39.4005
R5275 VDDA.n302 VDDA.t255 39.4005
R5276 VDDA.n286 VDDA.t22 39.4005
R5277 VDDA.n286 VDDA.t271 39.4005
R5278 VDDA.n284 VDDA.t158 39.4005
R5279 VDDA.n284 VDDA.t37 39.4005
R5280 VDDA.n282 VDDA.t269 39.4005
R5281 VDDA.n282 VDDA.t253 39.4005
R5282 VDDA.n280 VDDA.t61 39.4005
R5283 VDDA.n280 VDDA.t261 39.4005
R5284 VDDA.n279 VDDA.t257 39.4005
R5285 VDDA.n279 VDDA.t65 39.4005
R5286 VDDA.n389 VDDA.t447 39.4005
R5287 VDDA.n389 VDDA.t32 39.4005
R5288 VDDA.n406 VDDA.t162 39.4005
R5289 VDDA.n406 VDDA.t224 39.4005
R5290 VDDA.n455 VDDA.t247 39.4005
R5291 VDDA.n455 VDDA.t212 39.4005
R5292 VDDA.n412 VDDA.t458 39.4005
R5293 VDDA.n412 VDDA.t153 39.4005
R5294 VDDA.n436 VDDA.t222 39.4005
R5295 VDDA.n436 VDDA.t194 39.4005
R5296 VDDA.n438 VDDA.t30 39.4005
R5297 VDDA.n438 VDDA.t196 39.4005
R5298 VDDA.n440 VDDA.t214 39.4005
R5299 VDDA.n440 VDDA.t93 39.4005
R5300 VDDA.n442 VDDA.t441 39.4005
R5301 VDDA.n442 VDDA.t220 39.4005
R5302 VDDA.n418 VDDA.t2 39.4005
R5303 VDDA.n418 VDDA.t449 39.4005
R5304 VDDA.n424 VDDA.t245 39.4005
R5305 VDDA.n424 VDDA.t454 39.4005
R5306 VDDA.n144 VDDA.t188 31.4764
R5307 VDDA.t228 VDDA.n144 31.4764
R5308 VDDA.n70 VDDA.t54 31.4764
R5309 VDDA.n70 VDDA.t123 31.4764
R5310 VDDA.n260 VDDA.n254 28.9706
R5311 VDDA.n29 VDDA.n28 28.663
R5312 VDDA.n251 VDDA.n250 27.3072
R5313 VDDA.n243 VDDA.n242 27.3072
R5314 VDDA.n185 VDDA.n184 25.6005
R5315 VDDA.n173 VDDA.n172 25.6005
R5316 VDDA.n250 VDDA.n249 24.5338
R5317 VDDA.n244 VDDA.n243 24.5338
R5318 VDDA.n238 VDDA.n237 24.5338
R5319 VDDA.n230 VDDA.n229 24.5338
R5320 VDDA.n463 VDDA.n462 21.5914
R5321 VDDA.n254 VDDA.n253 21.5392
R5322 VDDA.n202 VDDA.n201 21.3338
R5323 VDDA.n200 VDDA.n199 21.3338
R5324 VDDA.n184 VDDA.n183 21.3338
R5325 VDDA.n174 VDDA.n173 21.3338
R5326 VDDA.n119 VDDA.n118 21.3338
R5327 VDDA.n117 VDDA.n116 21.3338
R5328 VDDA.n148 VDDA.n147 21.3338
R5329 VDDA.n141 VDDA.n140 21.3338
R5330 VDDA.n90 VDDA.n89 21.3338
R5331 VDDA.n88 VDDA.n87 21.3338
R5332 VDDA.n46 VDDA.n45 21.3338
R5333 VDDA.n44 VDDA.n43 21.3338
R5334 VDDA.n74 VDDA.n73 21.3338
R5335 VDDA.n64 VDDA.n63 21.3338
R5336 VDDA.n20 VDDA.n19 21.3338
R5337 VDDA.n27 VDDA.n18 21.3338
R5338 VDDA.n15 VDDA.n14 21.3338
R5339 VDDA.n35 VDDA.n13 21.3338
R5340 VDDA.n271 VDDA.n270 21.3338
R5341 VDDA.n276 VDDA.n274 21.3338
R5342 VDDA.n290 VDDA.n289 21.3338
R5343 VDDA.n292 VDDA.n291 21.3338
R5344 VDDA.n401 VDDA.n393 21.3338
R5345 VDDA.n391 VDDA.n390 21.3338
R5346 VDDA.n362 VDDA.n354 21.3338
R5347 VDDA.n352 VDDA.n351 21.3338
R5348 VDDA.n260 VDDA.t464 19.9244
R5349 VDDA.n37 VDDA.n36 19.5505
R5350 VDDA.n127 VDDA.n126 19.538
R5351 VDDA.n72 VDDA.n53 19.538
R5352 VDDA.n211 VDDA.n209 19.2005
R5353 VDDA.n99 VDDA.n97 19.2005
R5354 VDDA.n387 VDDA.n386 19.2005
R5355 VDDA.n380 VDDA.n379 19.2005
R5356 VDDA.n467 VDDA.n466 19.2005
R5357 VDDA.n459 VDDA.n458 19.2005
R5358 VDDA.n453 VDDA.n452 19.2005
R5359 VDDA.n446 VDDA.n445 19.2005
R5360 VDDA.n434 VDDA.n433 19.2005
R5361 VDDA.n427 VDDA.n426 19.2005
R5362 VDDA.n236 VDDA.n235 16.8187
R5363 VDDA.n188 VDDA.n111 16.813
R5364 VDDA.n378 VDDA.n363 16.363
R5365 VDDA.t282 VDDA.n234 16.1022
R5366 VDDA.n426 VDDA.n425 14.363
R5367 VDDA.n232 VDDA.n231 14.2313
R5368 VDDA.n228 VDDA.n221 14.0505
R5369 VDDA.n379 VDDA.n378 13.8005
R5370 VDDA.n388 VDDA.n387 13.8005
R5371 VDDA.n458 VDDA.n457 13.8005
R5372 VDDA.n445 VDDA.n444 13.8005
R5373 VDDA.n435 VDDA.n434 13.8005
R5374 VDDA.n454 VDDA.n453 13.8005
R5375 VDDA.n468 VDDA.n467 13.8005
R5376 VDDA.n37 VDDA.n10 13.6255
R5377 VDDA.n213 VDDA.n189 13.5943
R5378 VDDA.n345 VDDA.t142 13.1338
R5379 VDDA.n345 VDDA.t90 13.1338
R5380 VDDA.n364 VDDA.t462 13.1338
R5381 VDDA.n364 VDDA.t134 13.1338
R5382 VDDA.n366 VDDA.t108 13.1338
R5383 VDDA.n366 VDDA.t110 13.1338
R5384 VDDA.n368 VDDA.t132 13.1338
R5385 VDDA.n368 VDDA.t166 13.1338
R5386 VDDA.n370 VDDA.t164 13.1338
R5387 VDDA.n370 VDDA.t468 13.1338
R5388 VDDA.n372 VDDA.t130 13.1338
R5389 VDDA.n372 VDDA.t145 13.1338
R5390 VDDA.n374 VDDA.t76 13.1338
R5391 VDDA.n374 VDDA.t209 13.1338
R5392 VDDA.n376 VDDA.t168 13.1338
R5393 VDDA.n376 VDDA.t138 13.1338
R5394 VDDA.n264 VDDA.n263 11.6572
R5395 VDDA.n469 VDDA.n468 11.4105
R5396 VDDA.n210 VDDA.t311 11.2576
R5397 VDDA.n210 VDDA.t275 11.2576
R5398 VDDA.n194 VDDA.t281 11.2576
R5399 VDDA.n194 VDDA.t287 11.2576
R5400 VDDA.n193 VDDA.t293 11.2576
R5401 VDDA.n193 VDDA.t305 11.2576
R5402 VDDA.n191 VDDA.t291 11.2576
R5403 VDDA.n191 VDDA.t301 11.2576
R5404 VDDA.n190 VDDA.t279 11.2576
R5405 VDDA.n190 VDDA.t285 11.2576
R5406 VDDA.n98 VDDA.t313 11.2576
R5407 VDDA.n98 VDDA.t273 11.2576
R5408 VDDA.n82 VDDA.t277 11.2576
R5409 VDDA.n82 VDDA.t299 11.2576
R5410 VDDA.n81 VDDA.t295 11.2576
R5411 VDDA.n81 VDDA.t307 11.2576
R5412 VDDA.n79 VDDA.t309 11.2576
R5413 VDDA.n79 VDDA.t303 11.2576
R5414 VDDA.n78 VDDA.t289 11.2576
R5415 VDDA.n78 VDDA.t297 11.2576
R5416 VDDA.t341 VDDA.n226 11.0991
R5417 VDDA.n226 VDDA.t283 11.0991
R5418 VDDA.n405 VDDA.n404 9.75871
R5419 VDDA.n344 VDDA.n343 9.723
R5420 VDDA.n189 VDDA.n188 9.5005
R5421 VDDA.n212 VDDA.n211 9.3005
R5422 VDDA.n100 VDDA.n99 9.3005
R5423 VDDA.n331 VDDA.n277 9.3005
R5424 VDDA.n328 VDDA.n327 9.3005
R5425 VDDA.n326 VDDA.n325 9.3005
R5426 VDDA.n323 VDDA.n313 9.3005
R5427 VDDA.n322 VDDA.n321 9.3005
R5428 VDDA.n318 VDDA.n314 9.3005
R5429 VDDA.n269 VDDA.n268 9.3005
R5430 VDDA.n342 VDDA.n341 9.3005
R5431 VDDA.n335 VDDA.n334 9.3005
R5432 VDDA.n300 VDDA.n299 9.3005
R5433 VDDA.n403 VDDA.n402 9.3005
R5434 VDDA.n241 VDDA.n240 9.2505
R5435 VDDA.n110 VDDA.t438 8.0005
R5436 VDDA.n110 VDDA.t317 8.0005
R5437 VDDA.n108 VDDA.t86 8.0005
R5438 VDDA.n108 VDDA.t439 8.0005
R5439 VDDA.n106 VDDA.t25 8.0005
R5440 VDDA.n106 VDDA.t231 8.0005
R5441 VDDA.n104 VDDA.t241 8.0005
R5442 VDDA.n104 VDDA.t88 8.0005
R5443 VDDA.n102 VDDA.t243 8.0005
R5444 VDDA.n102 VDDA.t456 8.0005
R5445 VDDA.n101 VDDA.t315 8.0005
R5446 VDDA.n101 VDDA.t87 8.0005
R5447 VDDA.n9 VDDA.t314 8.0005
R5448 VDDA.n9 VDDA.t72 8.0005
R5449 VDDA.n7 VDDA.t59 8.0005
R5450 VDDA.n7 VDDA.t126 8.0005
R5451 VDDA.n5 VDDA.t94 8.0005
R5452 VDDA.n5 VDDA.t113 8.0005
R5453 VDDA.n3 VDDA.t8 8.0005
R5454 VDDA.n3 VDDA.t81 8.0005
R5455 VDDA.n1 VDDA.t215 8.0005
R5456 VDDA.n1 VDDA.t71 8.0005
R5457 VDDA.n0 VDDA.t3 8.0005
R5458 VDDA.n0 VDDA.t316 8.0005
R5459 VDDA.n213 VDDA.n212 7.8755
R5460 VDDA.n189 VDDA.n100 7.84425
R5461 VDDA.n253 VDDA.n252 6.6255
R5462 VDDA.n112 VDDA.t466 6.56717
R5463 VDDA.n112 VDDA.t203 6.56717
R5464 VDDA.n131 VDDA.t205 6.56717
R5465 VDDA.n131 VDDA.t24 6.56717
R5466 VDDA.n133 VDDA.t189 6.56717
R5467 VDDA.n133 VDDA.t229 6.56717
R5468 VDDA.n135 VDDA.t160 6.56717
R5469 VDDA.n135 VDDA.t235 6.56717
R5470 VDDA.n137 VDDA.t452 6.56717
R5471 VDDA.n137 VDDA.t233 6.56717
R5472 VDDA.n38 VDDA.t80 6.56717
R5473 VDDA.n38 VDDA.t20 6.56717
R5474 VDDA.n54 VDDA.t218 6.56717
R5475 VDDA.n54 VDDA.t58 6.56717
R5476 VDDA.n56 VDDA.t55 6.56717
R5477 VDDA.n56 VDDA.t124 6.56717
R5478 VDDA.n58 VDDA.t5 6.56717
R5479 VDDA.n58 VDDA.t7 6.56717
R5480 VDDA.n60 VDDA.t240 6.56717
R5481 VDDA.n60 VDDA.t151 6.56717
R5482 VDDA.n77 VDDA.n76 5.438
R5483 VDDA.n241 VDDA.n216 5.1255
R5484 VDDA.n214 VDDA.n77 5.0005
R5485 VDDA.n264 VDDA.n260 4.5595
R5486 VDDA.n212 VDDA.n196 4.5005
R5487 VDDA.n188 VDDA.n187 4.5005
R5488 VDDA.n100 VDDA.n84 4.5005
R5489 VDDA.n214 VDDA.n213 4.5005
R5490 VDDA.n301 VDDA.n300 4.5005
R5491 VDDA.n334 VDDA.n333 4.5005
R5492 VDDA.n332 VDDA.n331 4.5005
R5493 VDDA.n329 VDDA.n328 4.5005
R5494 VDDA.n325 VDDA.n310 4.5005
R5495 VDDA.n316 VDDA.n313 4.5005
R5496 VDDA.n321 VDDA.n320 4.5005
R5497 VDDA.n319 VDDA.n318 4.5005
R5498 VDDA.n268 VDDA.n265 4.5005
R5499 VDDA.n343 VDDA.n342 4.5005
R5500 VDDA.n404 VDDA.n403 4.5005
R5501 VDDA.n262 VDDA.n261 4.12334
R5502 VDDA.n234 VDDA.n233 4.02592
R5503 VDDA.n470 VDDA.n469 3.71013
R5504 VDDA.n333 VDDA.n309 3.3755
R5505 VDDA.n77 VDDA.n37 3.09425
R5506 VDDA.n187 VDDA.n186 2.96925
R5507 VDDA.n263 VDDA.n262 2.93377
R5508 VDDA.n404 VDDA.n388 2.47371
R5509 VDDA.n253 VDDA.n214 1.938
R5510 VDDA.n444 VDDA.n435 1.813
R5511 VDDA.n457 VDDA.n454 1.813
R5512 VDDA VDDA.n470 1.7019
R5513 VDDA.n470 VDDA.n254 1.105
R5514 VDDA.n378 VDDA.n377 1.0005
R5515 VDDA.n377 VDDA.n375 1.0005
R5516 VDDA.n375 VDDA.n373 1.0005
R5517 VDDA.n373 VDDA.n371 1.0005
R5518 VDDA.n371 VDDA.n369 1.0005
R5519 VDDA.n369 VDDA.n367 1.0005
R5520 VDDA.n367 VDDA.n365 1.0005
R5521 VDDA.n365 VDDA.n346 1.0005
R5522 VDDA.n388 VDDA.n346 1.0005
R5523 VDDA.n187 VDDA.n150 0.90675
R5524 VDDA.n344 VDDA.n264 0.840625
R5525 VDDA.n405 VDDA.n344 0.74075
R5526 VDDA.n240 VDDA.n221 0.6255
R5527 VDDA.n196 VDDA.n195 0.6255
R5528 VDDA.n196 VDDA.n192 0.6255
R5529 VDDA.n84 VDDA.n83 0.6255
R5530 VDDA.n84 VDDA.n80 0.6255
R5531 VDDA.n283 VDDA.n281 0.6255
R5532 VDDA.n285 VDDA.n283 0.6255
R5533 VDDA.n301 VDDA.n285 0.6255
R5534 VDDA.n303 VDDA.n301 0.6255
R5535 VDDA.n305 VDDA.n303 0.6255
R5536 VDDA.n307 VDDA.n305 0.6255
R5537 VDDA.n309 VDDA.n307 0.6255
R5538 VDDA.n333 VDDA.n332 0.6255
R5539 VDDA.n332 VDDA.n329 0.6255
R5540 VDDA.n329 VDDA.n310 0.6255
R5541 VDDA.n316 VDDA.n310 0.6255
R5542 VDDA.n320 VDDA.n316 0.6255
R5543 VDDA.n320 VDDA.n319 0.6255
R5544 VDDA.n319 VDDA.n265 0.6255
R5545 VDDA.n343 VDDA.n265 0.6255
R5546 VDDA.n171 VDDA.n169 0.563
R5547 VDDA.n169 VDDA.n167 0.563
R5548 VDDA.n167 VDDA.n165 0.563
R5549 VDDA.n165 VDDA.n163 0.563
R5550 VDDA.n163 VDDA.n161 0.563
R5551 VDDA.n161 VDDA.n159 0.563
R5552 VDDA.n159 VDDA.n157 0.563
R5553 VDDA.n157 VDDA.n155 0.563
R5554 VDDA.n155 VDDA.n152 0.563
R5555 VDDA.n186 VDDA.n152 0.563
R5556 VDDA.n138 VDDA.n136 0.563
R5557 VDDA.n136 VDDA.n134 0.563
R5558 VDDA.n134 VDDA.n132 0.563
R5559 VDDA.n132 VDDA.n113 0.563
R5560 VDDA.n150 VDDA.n113 0.563
R5561 VDDA.n105 VDDA.n103 0.563
R5562 VDDA.n107 VDDA.n105 0.563
R5563 VDDA.n109 VDDA.n107 0.563
R5564 VDDA.n111 VDDA.n109 0.563
R5565 VDDA.n61 VDDA.n59 0.563
R5566 VDDA.n59 VDDA.n57 0.563
R5567 VDDA.n57 VDDA.n55 0.563
R5568 VDDA.n55 VDDA.n39 0.563
R5569 VDDA.n76 VDDA.n39 0.563
R5570 VDDA.n4 VDDA.n2 0.563
R5571 VDDA.n6 VDDA.n4 0.563
R5572 VDDA.n8 VDDA.n6 0.563
R5573 VDDA.n10 VDDA.n8 0.563
R5574 VDDA.n425 VDDA.n419 0.563
R5575 VDDA.n435 VDDA.n419 0.563
R5576 VDDA.n444 VDDA.n443 0.563
R5577 VDDA.n443 VDDA.n441 0.563
R5578 VDDA.n441 VDDA.n439 0.563
R5579 VDDA.n439 VDDA.n437 0.563
R5580 VDDA.n437 VDDA.n413 0.563
R5581 VDDA.n454 VDDA.n413 0.563
R5582 VDDA.n457 VDDA.n456 0.563
R5583 VDDA.n456 VDDA.n407 0.563
R5584 VDDA.n468 VDDA.n407 0.563
R5585 VDDA VDDA.n405 0.41175
R5586 VDDA.n252 VDDA.n216 0.2505
R5587 VDDA.t210 VDDA.t463 0.1603
R5588 VDDA.t46 VDDA.t111 0.1603
R5589 VDDA.t91 VDDA.t51 0.1603
R5590 VDDA.t143 VDDA.t78 0.1603
R5591 VDDA.t136 VDDA.t139 0.1603
R5592 VDDA.n256 VDDA.t140 0.159278
R5593 VDDA.n257 VDDA.t44 0.159278
R5594 VDDA.n258 VDDA.t53 0.159278
R5595 VDDA.n259 VDDA.t77 0.159278
R5596 VDDA.n259 VDDA.t135 0.1368
R5597 VDDA.n259 VDDA.t210 0.1368
R5598 VDDA.n258 VDDA.t52 0.1368
R5599 VDDA.n258 VDDA.t46 0.1368
R5600 VDDA.n257 VDDA.t128 0.1368
R5601 VDDA.n257 VDDA.t91 0.1368
R5602 VDDA.n256 VDDA.t207 0.1368
R5603 VDDA.n256 VDDA.t143 0.1368
R5604 VDDA.n255 VDDA.t45 0.1368
R5605 VDDA.n255 VDDA.t136 0.1368
R5606 VDDA.n469 VDDA 0.135625
R5607 VDDA.t140 VDDA.n255 0.00152174
R5608 VDDA.t44 VDDA.n256 0.00152174
R5609 VDDA.t53 VDDA.n257 0.00152174
R5610 VDDA.t77 VDDA.n258 0.00152174
R5611 VDDA.t464 VDDA.n259 0.00152174
R5612 bgr_0.V_TOP.n0 bgr_0.V_TOP.t29 369.534
R5613 bgr_0.V_TOP.n23 bgr_0.V_TOP.n21 339.961
R5614 bgr_0.V_TOP.n23 bgr_0.V_TOP.n22 339.272
R5615 bgr_0.V_TOP.n19 bgr_0.V_TOP.n18 339.272
R5616 bgr_0.V_TOP.n27 bgr_0.V_TOP.n26 339.272
R5617 bgr_0.V_TOP.n29 bgr_0.V_TOP.n28 339.272
R5618 bgr_0.V_TOP.n24 bgr_0.V_TOP.n20 334.772
R5619 bgr_0.V_TOP.n39 bgr_0.V_TOP.n38 224.934
R5620 bgr_0.V_TOP.n38 bgr_0.V_TOP.n37 224.934
R5621 bgr_0.V_TOP.n37 bgr_0.V_TOP.n36 224.934
R5622 bgr_0.V_TOP.n36 bgr_0.V_TOP.n35 224.934
R5623 bgr_0.V_TOP.n35 bgr_0.V_TOP.n34 224.934
R5624 bgr_0.V_TOP.n34 bgr_0.V_TOP.n33 224.934
R5625 bgr_0.V_TOP.n33 bgr_0.V_TOP.n32 224.934
R5626 bgr_0.V_TOP.n1 bgr_0.V_TOP.n0 224.934
R5627 bgr_0.V_TOP.n2 bgr_0.V_TOP.n1 224.934
R5628 bgr_0.V_TOP.n3 bgr_0.V_TOP.n2 224.934
R5629 bgr_0.V_TOP.n4 bgr_0.V_TOP.n3 224.934
R5630 bgr_0.V_TOP.n5 bgr_0.V_TOP.n4 224.934
R5631 bgr_0.V_TOP bgr_0.V_TOP.t48 214.222
R5632 bgr_0.V_TOP.n31 bgr_0.V_TOP.n30 163.175
R5633 bgr_0.V_TOP.n39 bgr_0.V_TOP.t24 144.601
R5634 bgr_0.V_TOP.n38 bgr_0.V_TOP.t33 144.601
R5635 bgr_0.V_TOP.n37 bgr_0.V_TOP.t39 144.601
R5636 bgr_0.V_TOP.n36 bgr_0.V_TOP.t16 144.601
R5637 bgr_0.V_TOP.n35 bgr_0.V_TOP.t15 144.601
R5638 bgr_0.V_TOP.n34 bgr_0.V_TOP.t28 144.601
R5639 bgr_0.V_TOP.n33 bgr_0.V_TOP.t38 144.601
R5640 bgr_0.V_TOP.n32 bgr_0.V_TOP.t14 144.601
R5641 bgr_0.V_TOP.n0 bgr_0.V_TOP.t30 144.601
R5642 bgr_0.V_TOP.n1 bgr_0.V_TOP.t18 144.601
R5643 bgr_0.V_TOP.n2 bgr_0.V_TOP.t46 144.601
R5644 bgr_0.V_TOP.n3 bgr_0.V_TOP.t37 144.601
R5645 bgr_0.V_TOP.n4 bgr_0.V_TOP.t26 144.601
R5646 bgr_0.V_TOP.n5 bgr_0.V_TOP.t27 144.601
R5647 bgr_0.V_TOP.n17 bgr_0.V_TOP.t2 108.424
R5648 bgr_0.V_TOP.n30 bgr_0.V_TOP.t9 95.4467
R5649 bgr_0.V_TOP bgr_0.V_TOP.n39 69.6227
R5650 bgr_0.V_TOP.n32 bgr_0.V_TOP.n31 69.6227
R5651 bgr_0.V_TOP.n31 bgr_0.V_TOP.n5 69.6227
R5652 bgr_0.V_TOP.n18 bgr_0.V_TOP.t10 39.4005
R5653 bgr_0.V_TOP.n18 bgr_0.V_TOP.t7 39.4005
R5654 bgr_0.V_TOP.n20 bgr_0.V_TOP.t5 39.4005
R5655 bgr_0.V_TOP.n20 bgr_0.V_TOP.t1 39.4005
R5656 bgr_0.V_TOP.n22 bgr_0.V_TOP.t3 39.4005
R5657 bgr_0.V_TOP.n22 bgr_0.V_TOP.t13 39.4005
R5658 bgr_0.V_TOP.n21 bgr_0.V_TOP.t12 39.4005
R5659 bgr_0.V_TOP.n21 bgr_0.V_TOP.t4 39.4005
R5660 bgr_0.V_TOP.n26 bgr_0.V_TOP.t6 39.4005
R5661 bgr_0.V_TOP.n26 bgr_0.V_TOP.t8 39.4005
R5662 bgr_0.V_TOP.n28 bgr_0.V_TOP.t0 39.4005
R5663 bgr_0.V_TOP.n28 bgr_0.V_TOP.t11 39.4005
R5664 bgr_0.V_TOP.n17 bgr_0.V_TOP.n16 37.1479
R5665 bgr_0.V_TOP.n19 bgr_0.V_TOP.n17 27.8371
R5666 bgr_0.V_TOP.n24 bgr_0.V_TOP.n23 8.313
R5667 bgr_0.V_TOP.n30 bgr_0.V_TOP.n29 5.188
R5668 bgr_0.V_TOP.n6 bgr_0.V_TOP.t31 4.8295
R5669 bgr_0.V_TOP.n7 bgr_0.V_TOP.t22 4.8295
R5670 bgr_0.V_TOP.n8 bgr_0.V_TOP.t20 4.8295
R5671 bgr_0.V_TOP.n9 bgr_0.V_TOP.t45 4.8295
R5672 bgr_0.V_TOP.n10 bgr_0.V_TOP.t42 4.8295
R5673 bgr_0.V_TOP.n11 bgr_0.V_TOP.t36 4.8295
R5674 bgr_0.V_TOP.n12 bgr_0.V_TOP.t17 4.8295
R5675 bgr_0.V_TOP.n13 bgr_0.V_TOP.t43 4.8295
R5676 bgr_0.V_TOP.n14 bgr_0.V_TOP.t34 4.8295
R5677 bgr_0.V_TOP.n6 bgr_0.V_TOP.t35 4.5005
R5678 bgr_0.V_TOP.n7 bgr_0.V_TOP.t32 4.5005
R5679 bgr_0.V_TOP.n8 bgr_0.V_TOP.t25 4.5005
R5680 bgr_0.V_TOP.n9 bgr_0.V_TOP.t21 4.5005
R5681 bgr_0.V_TOP.n10 bgr_0.V_TOP.t49 4.5005
R5682 bgr_0.V_TOP.n11 bgr_0.V_TOP.t44 4.5005
R5683 bgr_0.V_TOP.n12 bgr_0.V_TOP.t23 4.5005
R5684 bgr_0.V_TOP.n13 bgr_0.V_TOP.t19 4.5005
R5685 bgr_0.V_TOP.n16 bgr_0.V_TOP.t40 4.5005
R5686 bgr_0.V_TOP.n15 bgr_0.V_TOP.t47 4.5005
R5687 bgr_0.V_TOP.n14 bgr_0.V_TOP.t41 4.5005
R5688 bgr_0.V_TOP.n25 bgr_0.V_TOP.n24 4.5005
R5689 bgr_0.V_TOP.n29 bgr_0.V_TOP.n27 2.1255
R5690 bgr_0.V_TOP.n27 bgr_0.V_TOP.n25 2.1255
R5691 bgr_0.V_TOP.n25 bgr_0.V_TOP.n19 2.1255
R5692 bgr_0.V_TOP.n7 bgr_0.V_TOP.n6 0.3295
R5693 bgr_0.V_TOP.n9 bgr_0.V_TOP.n8 0.3295
R5694 bgr_0.V_TOP.n11 bgr_0.V_TOP.n10 0.3295
R5695 bgr_0.V_TOP.n13 bgr_0.V_TOP.n12 0.3295
R5696 bgr_0.V_TOP.n16 bgr_0.V_TOP.n15 0.3295
R5697 bgr_0.V_TOP.n15 bgr_0.V_TOP.n14 0.3295
R5698 bgr_0.V_TOP.n9 bgr_0.V_TOP.n7 0.2825
R5699 bgr_0.V_TOP.n11 bgr_0.V_TOP.n9 0.2825
R5700 bgr_0.V_TOP.n13 bgr_0.V_TOP.n11 0.2825
R5701 bgr_0.V_TOP.n14 bgr_0.V_TOP.n13 0.2825
R5702 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 628.034
R5703 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 626.784
R5704 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 622.284
R5705 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 289.2
R5706 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 289.2
R5707 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 227.252
R5708 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 212.733
R5709 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 212.733
R5710 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 176.733
R5711 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 176.733
R5712 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 176.733
R5713 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 176.733
R5714 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 176.733
R5715 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 152
R5716 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 152
R5717 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 112.468
R5718 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 112.468
R5719 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 112.468
R5720 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 112.468
R5721 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 112.468
R5722 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 112.468
R5723 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 112.468
R5724 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 112.468
R5725 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 78.8005
R5726 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 78.8005
R5727 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 78.8005
R5728 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 78.8005
R5729 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 78.8005
R5730 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 78.8005
R5731 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 48.0005
R5732 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 48.0005
R5733 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 48.0005
R5734 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 48.0005
R5735 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 48.0005
R5736 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 48.0005
R5737 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 45.5227
R5738 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 45.5227
R5739 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 45.5227
R5740 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 45.5227
R5741 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 15.488
R5742 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 14.1755
R5743 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 5.7505
R5744 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 5.28175
R5745 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 0.84425
R5746 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.n7 114.719
R5747 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.n6 114.719
R5748 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n10 114.156
R5749 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.n8 114.156
R5750 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.n0 112.456
R5751 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.n18 112.454
R5752 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n17 111.206
R5753 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.n3 111.206
R5754 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.n1 111.206
R5755 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n5 109.656
R5756 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.n14 106.706
R5757 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.t2 16.0005
R5758 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.t14 16.0005
R5759 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t6 16.0005
R5760 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t5 16.0005
R5761 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.t12 16.0005
R5762 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.t9 16.0005
R5763 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.t19 16.0005
R5764 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.t10 16.0005
R5765 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.t7 16.0005
R5766 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.t4 16.0005
R5767 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t3 16.0005
R5768 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t21 16.0005
R5769 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t18 16.0005
R5770 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t0 16.0005
R5771 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t13 16.0005
R5772 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t15 16.0005
R5773 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t1 16.0005
R5774 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t17 16.0005
R5775 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.t11 16.0005
R5776 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.t8 16.0005
R5777 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.t20 16.0005
R5778 two_stage_opamp_dummy_magic_0.VD2.t16 two_stage_opamp_dummy_magic_0.VD2.n19 16.0005
R5779 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n12 4.5005
R5780 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n15 4.5005
R5781 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n4 3.6255
R5782 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.n2 1.2505
R5783 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n16 1.2505
R5784 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.n13 0.78175
R5785 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n9 0.563
R5786 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.n11 0.563
R5787 VOUT-.n14 VOUT-.n6 145.989
R5788 VOUT-.n9 VOUT-.n7 145.989
R5789 VOUT-.n13 VOUT-.n12 145.427
R5790 VOUT-.n11 VOUT-.n10 145.427
R5791 VOUT-.n9 VOUT-.n8 145.427
R5792 VOUT-.n16 VOUT-.n15 140.927
R5793 VOUT-.n5 VOUT-.t18 113.192
R5794 VOUT-.n2 VOUT-.n0 95.7303
R5795 VOUT-.n4 VOUT-.n3 94.6053
R5796 VOUT-.n2 VOUT-.n1 94.6053
R5797 VOUT-.n96 VOUT-.n16 20.813
R5798 VOUT-.n96 VOUT-.n95 11.6871
R5799 VOUT- VOUT-.n96 8.34425
R5800 VOUT-.n15 VOUT-.t2 6.56717
R5801 VOUT-.n15 VOUT-.t9 6.56717
R5802 VOUT-.n12 VOUT-.t5 6.56717
R5803 VOUT-.n12 VOUT-.t4 6.56717
R5804 VOUT-.n10 VOUT-.t7 6.56717
R5805 VOUT-.n10 VOUT-.t0 6.56717
R5806 VOUT-.n8 VOUT-.t1 6.56717
R5807 VOUT-.n8 VOUT-.t10 6.56717
R5808 VOUT-.n7 VOUT-.t8 6.56717
R5809 VOUT-.n7 VOUT-.t15 6.56717
R5810 VOUT-.n6 VOUT-.t14 6.56717
R5811 VOUT-.n6 VOUT-.t6 6.56717
R5812 VOUT-.n43 VOUT-.t85 4.8295
R5813 VOUT-.n45 VOUT-.t131 4.8295
R5814 VOUT-.n47 VOUT-.t31 4.8295
R5815 VOUT-.n49 VOUT-.t62 4.8295
R5816 VOUT-.n51 VOUT-.t114 4.8295
R5817 VOUT-.n63 VOUT-.t40 4.8295
R5818 VOUT-.n65 VOUT-.t34 4.8295
R5819 VOUT-.n66 VOUT-.t136 4.8295
R5820 VOUT-.n68 VOUT-.t70 4.8295
R5821 VOUT-.n69 VOUT-.t36 4.8295
R5822 VOUT-.n71 VOUT-.t95 4.8295
R5823 VOUT-.n72 VOUT-.t66 4.8295
R5824 VOUT-.n74 VOUT-.t55 4.8295
R5825 VOUT-.n75 VOUT-.t29 4.8295
R5826 VOUT-.n77 VOUT-.t91 4.8295
R5827 VOUT-.n78 VOUT-.t58 4.8295
R5828 VOUT-.n80 VOUT-.t49 4.8295
R5829 VOUT-.n81 VOUT-.t20 4.8295
R5830 VOUT-.n83 VOUT-.t148 4.8295
R5831 VOUT-.n84 VOUT-.t122 4.8295
R5832 VOUT-.n86 VOUT-.t44 4.8295
R5833 VOUT-.n87 VOUT-.t152 4.8295
R5834 VOUT-.n89 VOUT-.t142 4.8295
R5835 VOUT-.n90 VOUT-.t116 4.8295
R5836 VOUT-.n17 VOUT-.t108 4.8295
R5837 VOUT-.n29 VOUT-.t28 4.8295
R5838 VOUT-.n31 VOUT-.t24 4.8295
R5839 VOUT-.n32 VOUT-.t129 4.8295
R5840 VOUT-.n34 VOUT-.t61 4.8295
R5841 VOUT-.n35 VOUT-.t32 4.8295
R5842 VOUT-.n37 VOUT-.t100 4.8295
R5843 VOUT-.n38 VOUT-.t71 4.8295
R5844 VOUT-.n40 VOUT-.t69 4.8295
R5845 VOUT-.n41 VOUT-.t35 4.8295
R5846 VOUT-.n92 VOUT-.t77 4.8295
R5847 VOUT-.n56 VOUT-.t26 4.8154
R5848 VOUT-.n55 VOUT-.t59 4.8154
R5849 VOUT-.n54 VOUT-.t37 4.8154
R5850 VOUT-.n53 VOUT-.t81 4.8154
R5851 VOUT-.n62 VOUT-.t132 4.806
R5852 VOUT-.n61 VOUT-.t115 4.806
R5853 VOUT-.n60 VOUT-.t146 4.806
R5854 VOUT-.n59 VOUT-.t46 4.806
R5855 VOUT-.n58 VOUT-.t87 4.806
R5856 VOUT-.n57 VOUT-.t65 4.806
R5857 VOUT-.n56 VOUT-.t102 4.806
R5858 VOUT-.n55 VOUT-.t134 4.806
R5859 VOUT-.n54 VOUT-.t120 4.806
R5860 VOUT-.n53 VOUT-.t155 4.806
R5861 VOUT-.n28 VOUT-.t48 4.806
R5862 VOUT-.n27 VOUT-.t92 4.806
R5863 VOUT-.n26 VOUT-.t42 4.806
R5864 VOUT-.n25 VOUT-.t130 4.806
R5865 VOUT-.n24 VOUT-.t84 4.806
R5866 VOUT-.n23 VOUT-.t125 4.806
R5867 VOUT-.n22 VOUT-.t74 4.806
R5868 VOUT-.n21 VOUT-.t23 4.806
R5869 VOUT-.n20 VOUT-.t64 4.806
R5870 VOUT-.n19 VOUT-.t150 4.806
R5871 VOUT-.n44 VOUT-.t96 4.5005
R5872 VOUT-.n43 VOUT-.t57 4.5005
R5873 VOUT-.n45 VOUT-.t104 4.5005
R5874 VOUT-.n46 VOUT-.t73 4.5005
R5875 VOUT-.n47 VOUT-.t138 4.5005
R5876 VOUT-.n48 VOUT-.t107 4.5005
R5877 VOUT-.n49 VOUT-.t41 4.5005
R5878 VOUT-.n50 VOUT-.t143 4.5005
R5879 VOUT-.n51 VOUT-.t21 4.5005
R5880 VOUT-.n52 VOUT-.t126 4.5005
R5881 VOUT-.n53 VOUT-.t119 4.5005
R5882 VOUT-.n54 VOUT-.t82 4.5005
R5883 VOUT-.n55 VOUT-.t97 4.5005
R5884 VOUT-.n56 VOUT-.t63 4.5005
R5885 VOUT-.n57 VOUT-.t27 4.5005
R5886 VOUT-.n58 VOUT-.t45 4.5005
R5887 VOUT-.n59 VOUT-.t144 4.5005
R5888 VOUT-.n60 VOUT-.t112 4.5005
R5889 VOUT-.n61 VOUT-.t76 4.5005
R5890 VOUT-.n62 VOUT-.t93 4.5005
R5891 VOUT-.n64 VOUT-.t56 4.5005
R5892 VOUT-.n63 VOUT-.t19 4.5005
R5893 VOUT-.n65 VOUT-.t52 4.5005
R5894 VOUT-.n67 VOUT-.t156 4.5005
R5895 VOUT-.n66 VOUT-.t121 4.5005
R5896 VOUT-.n68 VOUT-.t89 4.5005
R5897 VOUT-.n70 VOUT-.t50 4.5005
R5898 VOUT-.n69 VOUT-.t151 4.5005
R5899 VOUT-.n71 VOUT-.t43 4.5005
R5900 VOUT-.n73 VOUT-.t145 4.5005
R5901 VOUT-.n72 VOUT-.t118 4.5005
R5902 VOUT-.n74 VOUT-.t141 4.5005
R5903 VOUT-.n76 VOUT-.t111 4.5005
R5904 VOUT-.n75 VOUT-.t80 4.5005
R5905 VOUT-.n77 VOUT-.t39 4.5005
R5906 VOUT-.n79 VOUT-.t139 4.5005
R5907 VOUT-.n78 VOUT-.t109 4.5005
R5908 VOUT-.n80 VOUT-.t135 4.5005
R5909 VOUT-.n82 VOUT-.t103 4.5005
R5910 VOUT-.n81 VOUT-.t72 4.5005
R5911 VOUT-.n83 VOUT-.t99 4.5005
R5912 VOUT-.n85 VOUT-.t68 4.5005
R5913 VOUT-.n84 VOUT-.t33 4.5005
R5914 VOUT-.n86 VOUT-.t133 4.5005
R5915 VOUT-.n88 VOUT-.t98 4.5005
R5916 VOUT-.n87 VOUT-.t67 4.5005
R5917 VOUT-.n89 VOUT-.t94 4.5005
R5918 VOUT-.n91 VOUT-.t60 4.5005
R5919 VOUT-.n90 VOUT-.t30 4.5005
R5920 VOUT-.n18 VOUT-.t101 4.5005
R5921 VOUT-.n17 VOUT-.t149 4.5005
R5922 VOUT-.n19 VOUT-.t88 4.5005
R5923 VOUT-.n20 VOUT-.t51 4.5005
R5924 VOUT-.n21 VOUT-.t137 4.5005
R5925 VOUT-.n22 VOUT-.t106 4.5005
R5926 VOUT-.n23 VOUT-.t75 4.5005
R5927 VOUT-.n24 VOUT-.t25 4.5005
R5928 VOUT-.n25 VOUT-.t128 4.5005
R5929 VOUT-.n26 VOUT-.t90 4.5005
R5930 VOUT-.n27 VOUT-.t54 4.5005
R5931 VOUT-.n28 VOUT-.t140 4.5005
R5932 VOUT-.n30 VOUT-.t110 4.5005
R5933 VOUT-.n29 VOUT-.t79 4.5005
R5934 VOUT-.n31 VOUT-.t113 4.5005
R5935 VOUT-.n33 VOUT-.t78 4.5005
R5936 VOUT-.n32 VOUT-.t38 4.5005
R5937 VOUT-.n34 VOUT-.t147 4.5005
R5938 VOUT-.n36 VOUT-.t117 4.5005
R5939 VOUT-.n35 VOUT-.t83 4.5005
R5940 VOUT-.n37 VOUT-.t47 4.5005
R5941 VOUT-.n39 VOUT-.t153 4.5005
R5942 VOUT-.n38 VOUT-.t123 4.5005
R5943 VOUT-.n40 VOUT-.t154 4.5005
R5944 VOUT-.n42 VOUT-.t124 4.5005
R5945 VOUT-.n41 VOUT-.t86 4.5005
R5946 VOUT-.n95 VOUT-.t105 4.5005
R5947 VOUT-.n94 VOUT-.t53 4.5005
R5948 VOUT-.n93 VOUT-.t22 4.5005
R5949 VOUT-.n92 VOUT-.t127 4.5005
R5950 VOUT-.n16 VOUT-.n14 4.5005
R5951 VOUT-.n3 VOUT-.t17 3.42907
R5952 VOUT-.n3 VOUT-.t12 3.42907
R5953 VOUT-.n1 VOUT-.t11 3.42907
R5954 VOUT-.n1 VOUT-.t16 3.42907
R5955 VOUT-.n0 VOUT-.t13 3.42907
R5956 VOUT-.n0 VOUT-.t3 3.42907
R5957 VOUT- VOUT-.n5 2.84425
R5958 VOUT-.n5 VOUT-.n4 2.15675
R5959 VOUT-.n4 VOUT-.n2 1.1255
R5960 VOUT-.n11 VOUT-.n9 0.563
R5961 VOUT-.n13 VOUT-.n11 0.563
R5962 VOUT-.n14 VOUT-.n13 0.563
R5963 VOUT-.n44 VOUT-.n43 0.3295
R5964 VOUT-.n46 VOUT-.n45 0.3295
R5965 VOUT-.n48 VOUT-.n47 0.3295
R5966 VOUT-.n50 VOUT-.n49 0.3295
R5967 VOUT-.n52 VOUT-.n51 0.3295
R5968 VOUT-.n54 VOUT-.n53 0.3295
R5969 VOUT-.n55 VOUT-.n54 0.3295
R5970 VOUT-.n56 VOUT-.n55 0.3295
R5971 VOUT-.n57 VOUT-.n56 0.3295
R5972 VOUT-.n58 VOUT-.n57 0.3295
R5973 VOUT-.n59 VOUT-.n58 0.3295
R5974 VOUT-.n60 VOUT-.n59 0.3295
R5975 VOUT-.n61 VOUT-.n60 0.3295
R5976 VOUT-.n62 VOUT-.n61 0.3295
R5977 VOUT-.n64 VOUT-.n62 0.3295
R5978 VOUT-.n64 VOUT-.n63 0.3295
R5979 VOUT-.n67 VOUT-.n65 0.3295
R5980 VOUT-.n67 VOUT-.n66 0.3295
R5981 VOUT-.n70 VOUT-.n68 0.3295
R5982 VOUT-.n70 VOUT-.n69 0.3295
R5983 VOUT-.n73 VOUT-.n71 0.3295
R5984 VOUT-.n73 VOUT-.n72 0.3295
R5985 VOUT-.n76 VOUT-.n74 0.3295
R5986 VOUT-.n76 VOUT-.n75 0.3295
R5987 VOUT-.n79 VOUT-.n77 0.3295
R5988 VOUT-.n79 VOUT-.n78 0.3295
R5989 VOUT-.n82 VOUT-.n80 0.3295
R5990 VOUT-.n82 VOUT-.n81 0.3295
R5991 VOUT-.n85 VOUT-.n83 0.3295
R5992 VOUT-.n85 VOUT-.n84 0.3295
R5993 VOUT-.n88 VOUT-.n86 0.3295
R5994 VOUT-.n88 VOUT-.n87 0.3295
R5995 VOUT-.n91 VOUT-.n89 0.3295
R5996 VOUT-.n91 VOUT-.n90 0.3295
R5997 VOUT-.n18 VOUT-.n17 0.3295
R5998 VOUT-.n20 VOUT-.n19 0.3295
R5999 VOUT-.n21 VOUT-.n20 0.3295
R6000 VOUT-.n22 VOUT-.n21 0.3295
R6001 VOUT-.n23 VOUT-.n22 0.3295
R6002 VOUT-.n24 VOUT-.n23 0.3295
R6003 VOUT-.n25 VOUT-.n24 0.3295
R6004 VOUT-.n26 VOUT-.n25 0.3295
R6005 VOUT-.n27 VOUT-.n26 0.3295
R6006 VOUT-.n28 VOUT-.n27 0.3295
R6007 VOUT-.n30 VOUT-.n28 0.3295
R6008 VOUT-.n30 VOUT-.n29 0.3295
R6009 VOUT-.n33 VOUT-.n31 0.3295
R6010 VOUT-.n33 VOUT-.n32 0.3295
R6011 VOUT-.n36 VOUT-.n34 0.3295
R6012 VOUT-.n36 VOUT-.n35 0.3295
R6013 VOUT-.n39 VOUT-.n37 0.3295
R6014 VOUT-.n39 VOUT-.n38 0.3295
R6015 VOUT-.n42 VOUT-.n40 0.3295
R6016 VOUT-.n42 VOUT-.n41 0.3295
R6017 VOUT-.n95 VOUT-.n94 0.3295
R6018 VOUT-.n94 VOUT-.n93 0.3295
R6019 VOUT-.n93 VOUT-.n92 0.3295
R6020 VOUT-.n60 VOUT-.n46 0.306
R6021 VOUT-.n59 VOUT-.n48 0.306
R6022 VOUT-.n58 VOUT-.n50 0.306
R6023 VOUT-.n57 VOUT-.n52 0.306
R6024 VOUT-.n64 VOUT-.n44 0.2825
R6025 VOUT-.n67 VOUT-.n64 0.2825
R6026 VOUT-.n70 VOUT-.n67 0.2825
R6027 VOUT-.n73 VOUT-.n70 0.2825
R6028 VOUT-.n76 VOUT-.n73 0.2825
R6029 VOUT-.n79 VOUT-.n76 0.2825
R6030 VOUT-.n82 VOUT-.n79 0.2825
R6031 VOUT-.n85 VOUT-.n82 0.2825
R6032 VOUT-.n88 VOUT-.n85 0.2825
R6033 VOUT-.n91 VOUT-.n88 0.2825
R6034 VOUT-.n30 VOUT-.n18 0.2825
R6035 VOUT-.n33 VOUT-.n30 0.2825
R6036 VOUT-.n36 VOUT-.n33 0.2825
R6037 VOUT-.n39 VOUT-.n36 0.2825
R6038 VOUT-.n42 VOUT-.n39 0.2825
R6039 VOUT-.n93 VOUT-.n42 0.2825
R6040 VOUT-.n93 VOUT-.n91 0.2825
R6041 two_stage_opamp_dummy_magic_0.cap_res_Y two_stage_opamp_dummy_magic_0.cap_res_Y.t0 49.083
R6042 two_stage_opamp_dummy_magic_0.cap_res_Y two_stage_opamp_dummy_magic_0.cap_res_Y.t126 0.922875
R6043 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 0.1603
R6044 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 0.1603
R6045 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 0.1603
R6046 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 0.1603
R6047 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 0.1603
R6048 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 0.1603
R6049 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 0.1603
R6050 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 0.1603
R6051 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 0.1603
R6052 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 0.1603
R6053 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 0.1603
R6054 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 0.1603
R6055 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 0.1603
R6056 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 0.1603
R6057 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 0.1603
R6058 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 0.1603
R6059 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 0.1603
R6060 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 0.1603
R6061 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 0.1603
R6062 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 0.1603
R6063 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 0.1603
R6064 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 0.1603
R6065 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 0.1603
R6066 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 0.1603
R6067 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 0.1603
R6068 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 0.1603
R6069 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 0.1603
R6070 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 0.1603
R6071 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 0.1603
R6072 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 0.1603
R6073 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 0.1603
R6074 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 0.1603
R6075 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 0.1603
R6076 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 0.1603
R6077 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 0.1603
R6078 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 0.1603
R6079 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 0.1603
R6080 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 0.1603
R6081 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 0.1603
R6082 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 0.1603
R6083 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 0.1603
R6084 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 0.1603
R6085 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 0.1603
R6086 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 0.1603
R6087 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 0.1603
R6088 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 0.1603
R6089 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 0.1603
R6090 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 0.1603
R6091 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 0.1603
R6092 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 0.1603
R6093 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 0.1603
R6094 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 0.1603
R6095 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 0.1603
R6096 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 0.1603
R6097 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 0.1603
R6098 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 0.1603
R6099 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 0.1603
R6100 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 0.1603
R6101 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 0.159278
R6102 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 0.159278
R6103 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 0.159278
R6104 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 0.159278
R6105 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 0.159278
R6106 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 0.159278
R6107 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 0.159278
R6108 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 0.159278
R6109 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 0.159278
R6110 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 0.159278
R6111 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 0.159278
R6112 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 0.159278
R6113 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 0.159278
R6114 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 0.159278
R6115 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 0.159278
R6116 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 0.159278
R6117 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 0.159278
R6118 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 0.159278
R6119 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 0.159278
R6120 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 0.159278
R6121 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 0.159278
R6122 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 0.159278
R6123 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 0.159278
R6124 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 0.159278
R6125 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 0.159278
R6126 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 0.159278
R6127 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 0.159278
R6128 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 0.137822
R6129 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 0.1368
R6130 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 0.1368
R6131 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 0.1368
R6132 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 0.1368
R6133 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 0.1368
R6134 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 0.1368
R6135 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 0.1368
R6136 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 0.1368
R6137 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 0.1368
R6138 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 0.1368
R6139 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 0.1368
R6140 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 0.1368
R6141 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 0.1368
R6142 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 0.1368
R6143 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 0.1368
R6144 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 0.1368
R6145 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 0.1368
R6146 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 0.1368
R6147 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 0.1368
R6148 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 0.1368
R6149 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 0.1368
R6150 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 0.1368
R6151 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 0.1368
R6152 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 0.1368
R6153 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 0.1368
R6154 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 0.1368
R6155 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 0.1368
R6156 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 0.1368
R6157 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 0.1368
R6158 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 0.1368
R6159 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 0.1368
R6160 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 0.114322
R6161 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 0.1133
R6162 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 0.1133
R6163 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 0.1133
R6164 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 0.1133
R6165 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 0.1133
R6166 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 0.1133
R6167 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 0.1133
R6168 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 0.1133
R6169 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 0.1133
R6170 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 0.1133
R6171 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 0.1133
R6172 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 0.1133
R6173 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 0.1133
R6174 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 0.1133
R6175 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 0.1133
R6176 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 0.1133
R6177 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 0.1133
R6178 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 0.1133
R6179 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 0.1133
R6180 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 0.00152174
R6181 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 0.00152174
R6182 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 0.00152174
R6183 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 0.00152174
R6184 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 0.00152174
R6185 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 0.00152174
R6186 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 0.00152174
R6187 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 0.00152174
R6188 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 0.00152174
R6189 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 0.00152174
R6190 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 0.00152174
R6191 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 0.00152174
R6192 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 0.00152174
R6193 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 0.00152174
R6194 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 0.00152174
R6195 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 0.00152174
R6196 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 0.00152174
R6197 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 0.00152174
R6198 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 0.00152174
R6199 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 0.00152174
R6200 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 0.00152174
R6201 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 0.00152174
R6202 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 0.00152174
R6203 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 0.00152174
R6204 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 0.00152174
R6205 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 0.00152174
R6206 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 0.00152174
R6207 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 0.00152174
R6208 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 0.00152174
R6209 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 0.00152174
R6210 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 0.00152174
R6211 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 0.00152174
R6212 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 0.00152174
R6213 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 0.00152174
R6214 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 0.00152174
R6215 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 0.00152174
R6216 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 688.859
R6217 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 514.134
R6218 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 323.491
R6219 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 322.692
R6220 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 270.591
R6221 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 270.591
R6222 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 270.591
R6223 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 270.591
R6224 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 233.374
R6225 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 233.374
R6226 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 233.374
R6227 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 233.374
R6228 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 214.056
R6229 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 174.726
R6230 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 174.726
R6231 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 174.726
R6232 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 174.726
R6233 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 173.591
R6234 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 169.216
R6235 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 169.216
R6236 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 129.24
R6237 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 129.24
R6238 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 129.24
R6239 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 129.24
R6240 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 128.534
R6241 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 128.534
R6242 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 125.817
R6243 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 46.1567
R6244 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 13.1338
R6245 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 13.1338
R6246 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 13.1338
R6247 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 13.1338
R6248 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 13.1338
R6249 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 13.1338
R6250 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 10.0317
R6251 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 4.3755
R6252 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 3.688
R6253 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 3.03175
R6254 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 2.0005
R6255 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 1.2755
R6256 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 1.2755
R6257 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 0.8005
R6258 two_stage_opamp_dummy_magic_0.Y.n49 two_stage_opamp_dummy_magic_0.Y.t31 1172.87
R6259 two_stage_opamp_dummy_magic_0.Y.n43 two_stage_opamp_dummy_magic_0.Y.t40 1172.87
R6260 two_stage_opamp_dummy_magic_0.Y.n50 two_stage_opamp_dummy_magic_0.Y.t50 996.134
R6261 two_stage_opamp_dummy_magic_0.Y.n49 two_stage_opamp_dummy_magic_0.Y.t39 996.134
R6262 two_stage_opamp_dummy_magic_0.Y.n43 two_stage_opamp_dummy_magic_0.Y.t53 996.134
R6263 two_stage_opamp_dummy_magic_0.Y.n44 two_stage_opamp_dummy_magic_0.Y.t43 996.134
R6264 two_stage_opamp_dummy_magic_0.Y.n45 two_stage_opamp_dummy_magic_0.Y.t26 996.134
R6265 two_stage_opamp_dummy_magic_0.Y.n46 two_stage_opamp_dummy_magic_0.Y.t32 996.134
R6266 two_stage_opamp_dummy_magic_0.Y.n47 two_stage_opamp_dummy_magic_0.Y.t48 996.134
R6267 two_stage_opamp_dummy_magic_0.Y.n48 two_stage_opamp_dummy_magic_0.Y.t35 996.134
R6268 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.t34 690.867
R6269 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.t45 690.867
R6270 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.t29 530.201
R6271 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.t38 530.201
R6272 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.t44 514.134
R6273 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.t54 514.134
R6274 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.t41 514.134
R6275 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.t51 514.134
R6276 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.t36 514.134
R6277 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.t28 514.134
R6278 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.t46 514.134
R6279 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.t27 514.134
R6280 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.t42 353.467
R6281 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.t25 353.467
R6282 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.t30 353.467
R6283 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.t47 353.467
R6284 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.t33 353.467
R6285 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.t49 353.467
R6286 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.t37 353.467
R6287 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.t52 353.467
R6288 two_stage_opamp_dummy_magic_0.Y.n50 two_stage_opamp_dummy_magic_0.Y.n49 176.733
R6289 two_stage_opamp_dummy_magic_0.Y.n44 two_stage_opamp_dummy_magic_0.Y.n43 176.733
R6290 two_stage_opamp_dummy_magic_0.Y.n45 two_stage_opamp_dummy_magic_0.Y.n44 176.733
R6291 two_stage_opamp_dummy_magic_0.Y.n46 two_stage_opamp_dummy_magic_0.Y.n45 176.733
R6292 two_stage_opamp_dummy_magic_0.Y.n47 two_stage_opamp_dummy_magic_0.Y.n46 176.733
R6293 two_stage_opamp_dummy_magic_0.Y.n48 two_stage_opamp_dummy_magic_0.Y.n47 176.733
R6294 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.n28 176.733
R6295 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.n27 176.733
R6296 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.n26 176.733
R6297 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.n25 176.733
R6298 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.n24 176.733
R6299 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.n23 176.733
R6300 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.n37 176.733
R6301 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.n36 176.733
R6302 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.n35 176.733
R6303 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.n34 176.733
R6304 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.n33 176.733
R6305 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.n32 176.733
R6306 two_stage_opamp_dummy_magic_0.Y.n52 two_stage_opamp_dummy_magic_0.Y.n51 166.436
R6307 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n30 161.843
R6308 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n39 161.718
R6309 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.n11 160.427
R6310 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.n18 159.802
R6311 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.n16 159.802
R6312 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.n14 159.802
R6313 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.n12 159.802
R6314 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.n20 155.302
R6315 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.n8 114.689
R6316 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.n1 114.689
R6317 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.n6 114.126
R6318 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.n4 114.126
R6319 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.n2 114.126
R6320 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n0 109.626
R6321 two_stage_opamp_dummy_magic_0.Y.n51 two_stage_opamp_dummy_magic_0.Y.n50 51.9494
R6322 two_stage_opamp_dummy_magic_0.Y.n51 two_stage_opamp_dummy_magic_0.Y.n48 51.9494
R6323 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.n29 51.9494
R6324 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.n22 51.9494
R6325 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n38 51.9494
R6326 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n31 51.9494
R6327 two_stage_opamp_dummy_magic_0.Y.t1 two_stage_opamp_dummy_magic_0.Y.n52 49.3036
R6328 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.n21 17.4067
R6329 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.t14 16.0005
R6330 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.t19 16.0005
R6331 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.t5 16.0005
R6332 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.t15 16.0005
R6333 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.t24 16.0005
R6334 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.t6 16.0005
R6335 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.t4 16.0005
R6336 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.t3 16.0005
R6337 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t18 16.0005
R6338 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t7 16.0005
R6339 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t9 16.0005
R6340 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t22 16.0005
R6341 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.n40 13.9693
R6342 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.t21 11.2576
R6343 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.t8 11.2576
R6344 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.t11 11.2576
R6345 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.t20 11.2576
R6346 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.t10 11.2576
R6347 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.t12 11.2576
R6348 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.t13 11.2576
R6349 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.t23 11.2576
R6350 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.t2 11.2576
R6351 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.t0 11.2576
R6352 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t17 11.2576
R6353 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t16 11.2576
R6354 two_stage_opamp_dummy_magic_0.Y.n42 two_stage_opamp_dummy_magic_0.Y.n10 9.28175
R6355 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.n19 5.1255
R6356 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n9 4.5005
R6357 two_stage_opamp_dummy_magic_0.Y.n42 two_stage_opamp_dummy_magic_0.Y.n41 4.5005
R6358 two_stage_opamp_dummy_magic_0.Y.n52 two_stage_opamp_dummy_magic_0.Y.n42 3.40675
R6359 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.n13 0.6255
R6360 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.n15 0.6255
R6361 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.n17 0.6255
R6362 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.n3 0.563
R6363 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.n5 0.563
R6364 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.n7 0.563
R6365 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 345.264
R6366 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 344.7
R6367 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 292.5
R6368 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 206.052
R6369 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 205.488
R6370 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 205.488
R6371 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 205.488
R6372 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 205.488
R6373 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 122.504
R6374 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 52.763
R6375 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 51.7297
R6376 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 42.313
R6377 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 39.4005
R6378 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 39.4005
R6379 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 39.4005
R6380 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 39.4005
R6381 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 39.4005
R6382 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 39.4005
R6383 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 19.7005
R6384 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 19.7005
R6385 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 19.7005
R6386 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 19.7005
R6387 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 19.7005
R6388 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 19.7005
R6389 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 19.7005
R6390 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 19.7005
R6391 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 19.7005
R6392 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 19.7005
R6393 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 6.21925
R6394 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 0.563
R6395 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 0.563
R6396 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 0.563
R6397 bgr_0.Vin+.n3 bgr_0.Vin+.n2 526.183
R6398 bgr_0.Vin+.n1 bgr_0.Vin+.n0 514.134
R6399 bgr_0.Vin+.n0 bgr_0.Vin+.t8 303.259
R6400 bgr_0.Vin+.n5 bgr_0.Vin+.n3 227.169
R6401 bgr_0.Vin+.n0 bgr_0.Vin+.t9 174.726
R6402 bgr_0.Vin+.n1 bgr_0.Vin+.t6 174.726
R6403 bgr_0.Vin+.n2 bgr_0.Vin+.t10 174.726
R6404 bgr_0.Vin+.n7 bgr_0.Vin+.n6 168.435
R6405 bgr_0.Vin+.n5 bgr_0.Vin+.n4 168.435
R6406 bgr_0.Vin+.n8 bgr_0.Vin+.t1 158.989
R6407 bgr_0.Vin+.n2 bgr_0.Vin+.n1 128.534
R6408 bgr_0.Vin+.t0 bgr_0.Vin+.n8 119.067
R6409 bgr_0.Vin+.n3 bgr_0.Vin+.t7 96.4005
R6410 bgr_0.Vin+.n8 bgr_0.Vin+.n7 35.0317
R6411 bgr_0.Vin+.n6 bgr_0.Vin+.t2 13.1338
R6412 bgr_0.Vin+.n6 bgr_0.Vin+.t5 13.1338
R6413 bgr_0.Vin+.n4 bgr_0.Vin+.t4 13.1338
R6414 bgr_0.Vin+.n4 bgr_0.Vin+.t3 13.1338
R6415 bgr_0.Vin+.n7 bgr_0.Vin+.n5 2.1255
R6416 bgr_0.V_mir1.n20 bgr_0.V_mir1.n19 325.473
R6417 bgr_0.V_mir1.n13 bgr_0.V_mir1.n12 325.473
R6418 bgr_0.V_mir1.n4 bgr_0.V_mir1.n3 325.473
R6419 bgr_0.V_mir1.n16 bgr_0.V_mir1.t19 310.488
R6420 bgr_0.V_mir1.n9 bgr_0.V_mir1.t21 310.488
R6421 bgr_0.V_mir1.n0 bgr_0.V_mir1.t20 310.488
R6422 bgr_0.V_mir1.n7 bgr_0.V_mir1.t14 278.312
R6423 bgr_0.V_mir1.n7 bgr_0.V_mir1.n6 228.939
R6424 bgr_0.V_mir1.n8 bgr_0.V_mir1.n5 224.439
R6425 bgr_0.V_mir1.n18 bgr_0.V_mir1.t8 184.097
R6426 bgr_0.V_mir1.n11 bgr_0.V_mir1.t4 184.097
R6427 bgr_0.V_mir1.n2 bgr_0.V_mir1.t2 184.097
R6428 bgr_0.V_mir1.n17 bgr_0.V_mir1.n16 167.094
R6429 bgr_0.V_mir1.n10 bgr_0.V_mir1.n9 167.094
R6430 bgr_0.V_mir1.n1 bgr_0.V_mir1.n0 167.094
R6431 bgr_0.V_mir1.n13 bgr_0.V_mir1.n11 152
R6432 bgr_0.V_mir1.n4 bgr_0.V_mir1.n2 152
R6433 bgr_0.V_mir1.n19 bgr_0.V_mir1.n18 152
R6434 bgr_0.V_mir1.n16 bgr_0.V_mir1.t22 120.501
R6435 bgr_0.V_mir1.n17 bgr_0.V_mir1.t12 120.501
R6436 bgr_0.V_mir1.n9 bgr_0.V_mir1.t17 120.501
R6437 bgr_0.V_mir1.n10 bgr_0.V_mir1.t10 120.501
R6438 bgr_0.V_mir1.n0 bgr_0.V_mir1.t18 120.501
R6439 bgr_0.V_mir1.n1 bgr_0.V_mir1.t6 120.501
R6440 bgr_0.V_mir1.n6 bgr_0.V_mir1.t0 48.0005
R6441 bgr_0.V_mir1.n6 bgr_0.V_mir1.t15 48.0005
R6442 bgr_0.V_mir1.n5 bgr_0.V_mir1.t16 48.0005
R6443 bgr_0.V_mir1.n5 bgr_0.V_mir1.t1 48.0005
R6444 bgr_0.V_mir1.n18 bgr_0.V_mir1.n17 40.7027
R6445 bgr_0.V_mir1.n11 bgr_0.V_mir1.n10 40.7027
R6446 bgr_0.V_mir1.n2 bgr_0.V_mir1.n1 40.7027
R6447 bgr_0.V_mir1.n12 bgr_0.V_mir1.t5 39.4005
R6448 bgr_0.V_mir1.n12 bgr_0.V_mir1.t11 39.4005
R6449 bgr_0.V_mir1.n3 bgr_0.V_mir1.t3 39.4005
R6450 bgr_0.V_mir1.n3 bgr_0.V_mir1.t7 39.4005
R6451 bgr_0.V_mir1.n20 bgr_0.V_mir1.t9 39.4005
R6452 bgr_0.V_mir1.t13 bgr_0.V_mir1.n20 39.4005
R6453 bgr_0.V_mir1.n15 bgr_0.V_mir1.n4 15.8005
R6454 bgr_0.V_mir1.n19 bgr_0.V_mir1.n15 15.8005
R6455 bgr_0.V_mir1.n14 bgr_0.V_mir1.n13 9.3005
R6456 bgr_0.V_mir1.n8 bgr_0.V_mir1.n7 5.8755
R6457 bgr_0.V_mir1.n15 bgr_0.V_mir1.n14 4.5005
R6458 bgr_0.V_mir1.n14 bgr_0.V_mir1.n8 0.78175
R6459 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.t13 354.854
R6460 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t21 346.8
R6461 bgr_0.1st_Vout_1.n20 bgr_0.1st_Vout_1.n19 339.522
R6462 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.n6 339.522
R6463 bgr_0.1st_Vout_1.n15 bgr_0.1st_Vout_1.n14 335.022
R6464 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t8 275.909
R6465 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.n10 227.909
R6466 bgr_0.1st_Vout_1.n13 bgr_0.1st_Vout_1.n12 222.034
R6467 bgr_0.1st_Vout_1.n17 bgr_0.1st_Vout_1.t22 184.097
R6468 bgr_0.1st_Vout_1.n17 bgr_0.1st_Vout_1.t32 184.097
R6469 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t16 184.097
R6470 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t36 184.097
R6471 bgr_0.1st_Vout_1.n18 bgr_0.1st_Vout_1.n17 166.05
R6472 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.n8 166.05
R6473 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.n4 54.2759
R6474 bgr_0.1st_Vout_1.n12 bgr_0.1st_Vout_1.t7 48.0005
R6475 bgr_0.1st_Vout_1.n12 bgr_0.1st_Vout_1.t10 48.0005
R6476 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t6 48.0005
R6477 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t9 48.0005
R6478 bgr_0.1st_Vout_1.n19 bgr_0.1st_Vout_1.t4 39.4005
R6479 bgr_0.1st_Vout_1.n19 bgr_0.1st_Vout_1.t2 39.4005
R6480 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t0 39.4005
R6481 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t3 39.4005
R6482 bgr_0.1st_Vout_1.n14 bgr_0.1st_Vout_1.t5 39.4005
R6483 bgr_0.1st_Vout_1.n14 bgr_0.1st_Vout_1.t1 39.4005
R6484 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t11 4.8295
R6485 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t29 4.8295
R6486 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t31 4.8295
R6487 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t20 4.8295
R6488 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t24 4.8295
R6489 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t14 4.8295
R6490 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t30 4.8295
R6491 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t18 4.8295
R6492 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t23 4.8295
R6493 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t15 4.5005
R6494 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t35 4.5005
R6495 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t34 4.5005
R6496 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t28 4.5005
R6497 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t27 4.5005
R6498 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t19 4.5005
R6499 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t33 4.5005
R6500 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t26 4.5005
R6501 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t25 4.5005
R6502 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t17 4.5005
R6503 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t12 4.5005
R6504 bgr_0.1st_Vout_1.n13 bgr_0.1st_Vout_1.n11 4.5005
R6505 bgr_0.1st_Vout_1.n16 bgr_0.1st_Vout_1.n15 4.5005
R6506 bgr_0.1st_Vout_1.n20 bgr_0.1st_Vout_1.n18 1.3755
R6507 bgr_0.1st_Vout_1.n16 bgr_0.1st_Vout_1.n9 1.3755
R6508 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.n5 1.188
R6509 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n2 0.8935
R6510 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.n0 0.8935
R6511 bgr_0.1st_Vout_1.n15 bgr_0.1st_Vout_1.n13 0.78175
R6512 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.n3 0.6585
R6513 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.n1 0.6585
R6514 bgr_0.1st_Vout_1.n18 bgr_0.1st_Vout_1.n16 0.6255
R6515 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.n7 0.6255
R6516 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n20 0.438
R6517 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 632.186
R6518 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 630.264
R6519 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 630.264
R6520 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 630.264
R6521 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 628.003
R6522 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 628.003
R6523 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 626.753
R6524 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 626.753
R6525 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 625.756
R6526 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 622.231
R6527 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 78.8005
R6528 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 78.8005
R6529 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 78.8005
R6530 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 78.8005
R6531 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 78.8005
R6532 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 78.8005
R6533 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 78.8005
R6534 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 78.8005
R6535 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 78.8005
R6536 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 78.8005
R6537 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 78.8005
R6538 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 78.8005
R6539 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 78.8005
R6540 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 78.8005
R6541 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 78.8005
R6542 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 78.8005
R6543 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 78.8005
R6544 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 78.8005
R6545 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 78.8005
R6546 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 78.8005
R6547 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 8.22272
R6548 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 6.188
R6549 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n28 630.264
R6550 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n3 627.316
R6551 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n5 626.784
R6552 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n4 626.784
R6553 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n27 626.784
R6554 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate.n25 585
R6555 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.t17 289.2
R6556 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.t29 289.2
R6557 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.n22 176.733
R6558 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.n6 176.733
R6559 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.n7 176.733
R6560 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.n8 176.733
R6561 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.n9 176.733
R6562 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.n10 176.733
R6563 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.n11 176.733
R6564 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.n12 176.733
R6565 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.n13 176.733
R6566 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.n14 176.733
R6567 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.n15 176.733
R6568 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.n16 176.733
R6569 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.n17 176.733
R6570 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.n18 176.733
R6571 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.n19 176.733
R6572 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.n20 176.733
R6573 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n2 175.013
R6574 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n24 162.494
R6575 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.t14 112.468
R6576 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.t27 112.468
R6577 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.t20 112.468
R6578 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.t26 112.468
R6579 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.t19 112.468
R6580 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.t31 112.468
R6581 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.t22 112.468
R6582 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.t33 112.468
R6583 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.t24 112.468
R6584 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.t15 112.468
R6585 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.t28 112.468
R6586 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.t18 112.468
R6587 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.t25 112.468
R6588 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.t16 112.468
R6589 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.t30 112.468
R6590 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.t21 112.468
R6591 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.t32 112.468
R6592 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.t23 112.468
R6593 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.t7 78.8005
R6594 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.t5 78.8005
R6595 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.t3 78.8005
R6596 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.t0 78.8005
R6597 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.t13 78.8005
R6598 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.t10 78.8005
R6599 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t6 78.8005
R6600 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t12 78.8005
R6601 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.t11 78.8005
R6602 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.t1 78.8005
R6603 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate.t2 78.8005
R6604 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate.t4 78.8005
R6605 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n1 54.7817
R6606 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.n23 49.8072
R6607 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.n21 49.8072
R6608 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n26 41.7838
R6609 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate 39.8442
R6610 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.t8 24.0005
R6611 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.t9 24.0005
R6612 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n0 2.313
R6613 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.t33 355.293
R6614 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t34 346.8
R6615 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.n12 339.522
R6616 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n5 339.522
R6617 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n10 335.022
R6618 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t8 275.909
R6619 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.n7 227.909
R6620 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n9 222.034
R6621 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.t13 184.097
R6622 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.t24 184.097
R6623 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t16 184.097
R6624 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t27 184.097
R6625 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n11 166.05
R6626 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n6 166.05
R6627 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n4 52.9634
R6628 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.t9 48.0005
R6629 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.t3 48.0005
R6630 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t4 48.0005
R6631 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t10 48.0005
R6632 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t7 39.4005
R6633 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t5 39.4005
R6634 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t1 39.4005
R6635 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t2 39.4005
R6636 bgr_0.1st_Vout_2.t0 bgr_0.1st_Vout_2.n13 39.4005
R6637 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.t6 39.4005
R6638 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n3 5.28175
R6639 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t17 4.8295
R6640 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t35 4.8295
R6641 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t11 4.8295
R6642 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t26 4.8295
R6643 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t30 4.8295
R6644 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t19 4.8295
R6645 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t36 4.8295
R6646 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t25 4.8295
R6647 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t18 4.8295
R6648 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n8 4.5005
R6649 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t12 4.5005
R6650 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t32 4.5005
R6651 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t31 4.5005
R6652 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t23 4.5005
R6653 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t22 4.5005
R6654 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t15 4.5005
R6655 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t29 4.5005
R6656 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t21 4.5005
R6657 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t28 4.5005
R6658 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t20 4.5005
R6659 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t14 4.5005
R6660 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n0 3.188
R6661 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.n2 3.1025
R6662 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.n1 2.0005
R6663 bgr_0.cap_res2.t20 bgr_0.cap_res2.t17 121.245
R6664 bgr_0.cap_res2.t12 bgr_0.cap_res2.t6 0.1603
R6665 bgr_0.cap_res2.t5 bgr_0.cap_res2.t0 0.1603
R6666 bgr_0.cap_res2.t10 bgr_0.cap_res2.t4 0.1603
R6667 bgr_0.cap_res2.t3 bgr_0.cap_res2.t19 0.1603
R6668 bgr_0.cap_res2.t18 bgr_0.cap_res2.t15 0.1603
R6669 bgr_0.cap_res2.n1 bgr_0.cap_res2.t2 0.159278
R6670 bgr_0.cap_res2.n2 bgr_0.cap_res2.t9 0.159278
R6671 bgr_0.cap_res2.n3 bgr_0.cap_res2.t16 0.159278
R6672 bgr_0.cap_res2.n4 bgr_0.cap_res2.t11 0.159278
R6673 bgr_0.cap_res2.n4 bgr_0.cap_res2.t14 0.1368
R6674 bgr_0.cap_res2.n4 bgr_0.cap_res2.t12 0.1368
R6675 bgr_0.cap_res2.n3 bgr_0.cap_res2.t8 0.1368
R6676 bgr_0.cap_res2.n3 bgr_0.cap_res2.t5 0.1368
R6677 bgr_0.cap_res2.n2 bgr_0.cap_res2.t13 0.1368
R6678 bgr_0.cap_res2.n2 bgr_0.cap_res2.t10 0.1368
R6679 bgr_0.cap_res2.n1 bgr_0.cap_res2.t7 0.1368
R6680 bgr_0.cap_res2.n1 bgr_0.cap_res2.t3 0.1368
R6681 bgr_0.cap_res2.n0 bgr_0.cap_res2.t1 0.1368
R6682 bgr_0.cap_res2.n0 bgr_0.cap_res2.t18 0.1368
R6683 bgr_0.cap_res2.t2 bgr_0.cap_res2.n0 0.00152174
R6684 bgr_0.cap_res2.t9 bgr_0.cap_res2.n1 0.00152174
R6685 bgr_0.cap_res2.t16 bgr_0.cap_res2.n2 0.00152174
R6686 bgr_0.cap_res2.t11 bgr_0.cap_res2.n3 0.00152174
R6687 bgr_0.cap_res2.t17 bgr_0.cap_res2.n4 0.00152174
R6688 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.t19 673.034
R6689 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.n0 620.841
R6690 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.t28 611.739
R6691 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.t16 611.739
R6692 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.t22 611.739
R6693 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.t31 611.739
R6694 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.t11 421.75
R6695 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.t13 421.75
R6696 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.t15 421.75
R6697 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.t18 421.75
R6698 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.t14 421.75
R6699 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.t12 421.75
R6700 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.t29 421.75
R6701 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.t24 421.75
R6702 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.t27 421.75
R6703 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.t25 421.75
R6704 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.t30 421.75
R6705 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.t17 421.75
R6706 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.t26 421.75
R6707 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.t21 421.75
R6708 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.t23 421.75
R6709 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.t20 421.75
R6710 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.t0 284.55
R6711 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.n10 169.405
R6712 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.n19 168.843
R6713 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.n15 167.094
R6714 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.n16 167.094
R6715 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.n17 167.094
R6716 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.n11 167.094
R6717 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.n12 167.094
R6718 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.n13 167.094
R6719 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.n6 167.094
R6720 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.n7 167.094
R6721 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.n8 167.094
R6722 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.n2 167.094
R6723 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.n3 167.094
R6724 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.n4 167.094
R6725 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n27 140.857
R6726 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.n25 139.608
R6727 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.n23 139.608
R6728 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n28 139.608
R6729 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t10 65.6672
R6730 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t1 65.6672
R6731 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.n22 60.8755
R6732 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.n18 47.1294
R6733 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.n14 47.1294
R6734 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.n9 47.1294
R6735 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.n5 47.1294
R6736 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.t6 24.0005
R6737 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.t8 24.0005
R6738 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.t4 24.0005
R6739 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.t2 24.0005
R6740 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.t9 24.0005
R6741 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.t3 24.0005
R6742 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.t5 24.0005
R6743 two_stage_opamp_dummy_magic_0.Vb2.t7 two_stage_opamp_dummy_magic_0.Vb2.n29 24.0005
R6744 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.n1 17.8942
R6745 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.n20 13.0943
R6746 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n26 7.563
R6747 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.n21 4.5005
R6748 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.n24 1.2505
R6749 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n4 4020
R6750 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.n4 4020
R6751 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n10 4020
R6752 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.n10 4020
R6753 two_stage_opamp_dummy_magic_0.VD4.n7 two_stage_opamp_dummy_magic_0.VD4.t3 660.109
R6754 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.t0 660.109
R6755 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.n14 422.401
R6756 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.n3 422.401
R6757 two_stage_opamp_dummy_magic_0.VD4.t4 two_stage_opamp_dummy_magic_0.VD4.n11 239.915
R6758 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.t1 239.915
R6759 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.n8 230.4
R6760 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.n6 230.4
R6761 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.n6 198.4
R6762 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n3 198.4
R6763 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.n0 160.428
R6764 two_stage_opamp_dummy_magic_0.VD4.n25 two_stage_opamp_dummy_magic_0.VD4.n23 160.427
R6765 two_stage_opamp_dummy_magic_0.VD4.n22 two_stage_opamp_dummy_magic_0.VD4.n21 159.804
R6766 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.n19 159.803
R6767 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.n1 159.803
R6768 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.n32 159.802
R6769 two_stage_opamp_dummy_magic_0.VD4.n31 two_stage_opamp_dummy_magic_0.VD4.n30 159.802
R6770 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.n28 159.802
R6771 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n26 159.802
R6772 two_stage_opamp_dummy_magic_0.VD4.n25 two_stage_opamp_dummy_magic_0.VD4.n24 159.802
R6773 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.n16 155.303
R6774 two_stage_opamp_dummy_magic_0.VD4.n7 two_stage_opamp_dummy_magic_0.VD4.t5 155.125
R6775 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.t2 155.125
R6776 two_stage_opamp_dummy_magic_0.VD4.t14 two_stage_opamp_dummy_magic_0.VD4.t4 98.2764
R6777 two_stage_opamp_dummy_magic_0.VD4.t18 two_stage_opamp_dummy_magic_0.VD4.t14 98.2764
R6778 two_stage_opamp_dummy_magic_0.VD4.t22 two_stage_opamp_dummy_magic_0.VD4.t18 98.2764
R6779 two_stage_opamp_dummy_magic_0.VD4.t6 two_stage_opamp_dummy_magic_0.VD4.t22 98.2764
R6780 two_stage_opamp_dummy_magic_0.VD4.t10 two_stage_opamp_dummy_magic_0.VD4.t6 98.2764
R6781 two_stage_opamp_dummy_magic_0.VD4.t16 two_stage_opamp_dummy_magic_0.VD4.t12 98.2764
R6782 two_stage_opamp_dummy_magic_0.VD4.t20 two_stage_opamp_dummy_magic_0.VD4.t16 98.2764
R6783 two_stage_opamp_dummy_magic_0.VD4.t24 two_stage_opamp_dummy_magic_0.VD4.t20 98.2764
R6784 two_stage_opamp_dummy_magic_0.VD4.t8 two_stage_opamp_dummy_magic_0.VD4.t24 98.2764
R6785 two_stage_opamp_dummy_magic_0.VD4.t1 two_stage_opamp_dummy_magic_0.VD4.t8 98.2764
R6786 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.n13 92.5005
R6787 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.n9 92.5005
R6788 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n10 92.5005
R6789 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n3 92.5005
R6790 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.n4 92.5005
R6791 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n4 92.5005
R6792 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.t10 49.1384
R6793 two_stage_opamp_dummy_magic_0.VD4.t12 two_stage_opamp_dummy_magic_0.VD4.n12 49.1384
R6794 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n7 21.3338
R6795 two_stage_opamp_dummy_magic_0.VD4.n6 two_stage_opamp_dummy_magic_0.VD4.n5 21.3338
R6796 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.t36 11.2576
R6797 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.t27 11.2576
R6798 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.t29 11.2576
R6799 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.t31 11.2576
R6800 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.t33 11.2576
R6801 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.t35 11.2576
R6802 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.t26 11.2576
R6803 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.t28 11.2576
R6804 two_stage_opamp_dummy_magic_0.VD4.n24 two_stage_opamp_dummy_magic_0.VD4.t30 11.2576
R6805 two_stage_opamp_dummy_magic_0.VD4.n24 two_stage_opamp_dummy_magic_0.VD4.t32 11.2576
R6806 two_stage_opamp_dummy_magic_0.VD4.n23 two_stage_opamp_dummy_magic_0.VD4.t34 11.2576
R6807 two_stage_opamp_dummy_magic_0.VD4.n23 two_stage_opamp_dummy_magic_0.VD4.t37 11.2576
R6808 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.t17 11.2576
R6809 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.t21 11.2576
R6810 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.t11 11.2576
R6811 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.t13 11.2576
R6812 two_stage_opamp_dummy_magic_0.VD4.n1 two_stage_opamp_dummy_magic_0.VD4.t23 11.2576
R6813 two_stage_opamp_dummy_magic_0.VD4.n1 two_stage_opamp_dummy_magic_0.VD4.t7 11.2576
R6814 two_stage_opamp_dummy_magic_0.VD4.n0 two_stage_opamp_dummy_magic_0.VD4.t15 11.2576
R6815 two_stage_opamp_dummy_magic_0.VD4.n0 two_stage_opamp_dummy_magic_0.VD4.t19 11.2576
R6816 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.t25 11.2576
R6817 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.t9 11.2576
R6818 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.n15 9.5505
R6819 two_stage_opamp_dummy_magic_0.VD4 two_stage_opamp_dummy_magic_0.VD4.n33 8.5005
R6820 two_stage_opamp_dummy_magic_0.VD4 two_stage_opamp_dummy_magic_0.VD4.n22 5.938
R6821 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.n17 4.5005
R6822 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n25 0.6255
R6823 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.n27 0.6255
R6824 two_stage_opamp_dummy_magic_0.VD4.n31 two_stage_opamp_dummy_magic_0.VD4.n29 0.6255
R6825 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.n31 0.6255
R6826 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.n2 0.6255
R6827 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.n18 0.6255
R6828 two_stage_opamp_dummy_magic_0.VD4.n22 two_stage_opamp_dummy_magic_0.VD4.n20 0.6255
R6829 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.t29 1172.87
R6830 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t34 1172.87
R6831 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.t51 996.134
R6832 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.t39 996.134
R6833 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.t26 996.134
R6834 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.t44 996.134
R6835 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.t25 996.134
R6836 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.t43 996.134
R6837 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t49 996.134
R6838 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.t36 996.134
R6839 two_stage_opamp_dummy_magic_0.X.n48 two_stage_opamp_dummy_magic_0.X.t32 690.867
R6840 two_stage_opamp_dummy_magic_0.X.n41 two_stage_opamp_dummy_magic_0.X.t37 690.867
R6841 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.t28 530.201
R6842 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.t33 530.201
R6843 two_stage_opamp_dummy_magic_0.X.n48 two_stage_opamp_dummy_magic_0.X.t46 514.134
R6844 two_stage_opamp_dummy_magic_0.X.n47 two_stage_opamp_dummy_magic_0.X.t30 514.134
R6845 two_stage_opamp_dummy_magic_0.X.n46 two_stage_opamp_dummy_magic_0.X.t47 514.134
R6846 two_stage_opamp_dummy_magic_0.X.n45 two_stage_opamp_dummy_magic_0.X.t31 514.134
R6847 two_stage_opamp_dummy_magic_0.X.n44 two_stage_opamp_dummy_magic_0.X.t45 514.134
R6848 two_stage_opamp_dummy_magic_0.X.n43 two_stage_opamp_dummy_magic_0.X.t27 514.134
R6849 two_stage_opamp_dummy_magic_0.X.n42 two_stage_opamp_dummy_magic_0.X.t40 514.134
R6850 two_stage_opamp_dummy_magic_0.X.n41 two_stage_opamp_dummy_magic_0.X.t52 514.134
R6851 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.t41 353.467
R6852 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.t48 353.467
R6853 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.t35 353.467
R6854 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.t50 353.467
R6855 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.t38 353.467
R6856 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.t54 353.467
R6857 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.t42 353.467
R6858 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.t53 353.467
R6859 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.n17 176.733
R6860 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.n16 176.733
R6861 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.n15 176.733
R6862 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.n14 176.733
R6863 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.n13 176.733
R6864 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.n11 176.733
R6865 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.n32 176.733
R6866 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.n33 176.733
R6867 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.n34 176.733
R6868 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.n35 176.733
R6869 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.n36 176.733
R6870 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.n37 176.733
R6871 two_stage_opamp_dummy_magic_0.X.n42 two_stage_opamp_dummy_magic_0.X.n41 176.733
R6872 two_stage_opamp_dummy_magic_0.X.n43 two_stage_opamp_dummy_magic_0.X.n42 176.733
R6873 two_stage_opamp_dummy_magic_0.X.n44 two_stage_opamp_dummy_magic_0.X.n43 176.733
R6874 two_stage_opamp_dummy_magic_0.X.n45 two_stage_opamp_dummy_magic_0.X.n44 176.733
R6875 two_stage_opamp_dummy_magic_0.X.n46 two_stage_opamp_dummy_magic_0.X.n45 176.733
R6876 two_stage_opamp_dummy_magic_0.X.n47 two_stage_opamp_dummy_magic_0.X.n46 176.733
R6877 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.n19 166.436
R6878 two_stage_opamp_dummy_magic_0.X.n50 two_stage_opamp_dummy_magic_0.X.n40 161.843
R6879 two_stage_opamp_dummy_magic_0.X.n50 two_stage_opamp_dummy_magic_0.X.n49 161.718
R6880 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.n21 160.427
R6881 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.n28 159.802
R6882 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.n26 159.802
R6883 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.n24 159.802
R6884 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.n22 159.802
R6885 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.n30 155.302
R6886 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.n2 114.689
R6887 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.n1 114.689
R6888 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.n7 114.126
R6889 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.n5 114.126
R6890 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.n3 114.126
R6891 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n0 109.626
R6892 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n18 51.9494
R6893 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n12 51.9494
R6894 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n39 51.9494
R6895 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n38 51.9494
R6896 two_stage_opamp_dummy_magic_0.X.n49 two_stage_opamp_dummy_magic_0.X.n48 51.9494
R6897 two_stage_opamp_dummy_magic_0.X.n49 two_stage_opamp_dummy_magic_0.X.n47 51.9494
R6898 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.t1 49.3037
R6899 two_stage_opamp_dummy_magic_0.X.n51 two_stage_opamp_dummy_magic_0.X.n31 17.438
R6900 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.t17 16.0005
R6901 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.t23 16.0005
R6902 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.t3 16.0005
R6903 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.t20 16.0005
R6904 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.t22 16.0005
R6905 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.t14 16.0005
R6906 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.t0 16.0005
R6907 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.t18 16.0005
R6908 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t19 16.0005
R6909 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t21 16.0005
R6910 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t16 16.0005
R6911 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t15 16.0005
R6912 two_stage_opamp_dummy_magic_0.X.n51 two_stage_opamp_dummy_magic_0.X.n50 13.938
R6913 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.t24 11.2576
R6914 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.t12 11.2576
R6915 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.t9 11.2576
R6916 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.t13 11.2576
R6917 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.t6 11.2576
R6918 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.t4 11.2576
R6919 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.t10 11.2576
R6920 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.t11 11.2576
R6921 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.t5 11.2576
R6922 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.t8 11.2576
R6923 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.t7 11.2576
R6924 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.t2 11.2576
R6925 two_stage_opamp_dummy_magic_0.X.n53 two_stage_opamp_dummy_magic_0.X.n52 7.53175
R6926 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.n29 5.1255
R6927 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n9 4.5005
R6928 two_stage_opamp_dummy_magic_0.X.n52 two_stage_opamp_dummy_magic_0.X.n51 4.5005
R6929 two_stage_opamp_dummy_magic_0.X.n52 two_stage_opamp_dummy_magic_0.X.n20 3.3755
R6930 two_stage_opamp_dummy_magic_0.X.n53 two_stage_opamp_dummy_magic_0.X.n10 1.71925
R6931 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.n23 0.6255
R6932 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.n25 0.6255
R6933 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.n27 0.6255
R6934 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.n4 0.563
R6935 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.n6 0.563
R6936 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.n8 0.563
R6937 two_stage_opamp_dummy_magic_0.X two_stage_opamp_dummy_magic_0.X.n53 0.063
R6938 VOUT+.n2 VOUT+.n0 145.989
R6939 VOUT+.n8 VOUT+.n7 145.989
R6940 VOUT+.n6 VOUT+.n5 145.427
R6941 VOUT+.n4 VOUT+.n3 145.427
R6942 VOUT+.n2 VOUT+.n1 145.427
R6943 VOUT+.n10 VOUT+.n9 140.927
R6944 VOUT+.n96 VOUT+.t0 113.192
R6945 VOUT+.n93 VOUT+.n91 95.7303
R6946 VOUT+.n95 VOUT+.n94 94.6053
R6947 VOUT+.n93 VOUT+.n92 94.6053
R6948 VOUT+.n90 VOUT+.n10 20.813
R6949 VOUT+.n90 VOUT+.n89 11.6871
R6950 VOUT+ VOUT+.n90 8.34425
R6951 VOUT+.n9 VOUT+.t11 6.56717
R6952 VOUT+.n9 VOUT+.t5 6.56717
R6953 VOUT+.n7 VOUT+.t9 6.56717
R6954 VOUT+.n7 VOUT+.t18 6.56717
R6955 VOUT+.n5 VOUT+.t10 6.56717
R6956 VOUT+.n5 VOUT+.t4 6.56717
R6957 VOUT+.n3 VOUT+.t2 6.56717
R6958 VOUT+.n3 VOUT+.t6 6.56717
R6959 VOUT+.n1 VOUT+.t3 6.56717
R6960 VOUT+.n1 VOUT+.t7 6.56717
R6961 VOUT+.n0 VOUT+.t17 6.56717
R6962 VOUT+.n0 VOUT+.t8 6.56717
R6963 VOUT+.n37 VOUT+.t108 4.8295
R6964 VOUT+.n46 VOUT+.t65 4.8295
R6965 VOUT+.n44 VOUT+.t118 4.8295
R6966 VOUT+.n42 VOUT+.t151 4.8295
R6967 VOUT+.n40 VOUT+.t44 4.8295
R6968 VOUT+.n39 VOUT+.t67 4.8295
R6969 VOUT+.n59 VOUT+.t27 4.8295
R6970 VOUT+.n60 VOUT+.t76 4.8295
R6971 VOUT+.n62 VOUT+.t62 4.8295
R6972 VOUT+.n63 VOUT+.t112 4.8295
R6973 VOUT+.n65 VOUT+.t114 4.8295
R6974 VOUT+.n66 VOUT+.t99 4.8295
R6975 VOUT+.n68 VOUT+.t74 4.8295
R6976 VOUT+.n69 VOUT+.t55 4.8295
R6977 VOUT+.n71 VOUT+.t109 4.8295
R6978 VOUT+.n72 VOUT+.t91 4.8295
R6979 VOUT+.n74 VOUT+.t68 4.8295
R6980 VOUT+.n75 VOUT+.t52 4.8295
R6981 VOUT+.n77 VOUT+.t29 4.8295
R6982 VOUT+.n78 VOUT+.t153 4.8295
R6983 VOUT+.n80 VOUT+.t63 4.8295
R6984 VOUT+.n81 VOUT+.t46 4.8295
R6985 VOUT+.n83 VOUT+.t22 4.8295
R6986 VOUT+.n84 VOUT+.t146 4.8295
R6987 VOUT+.n11 VOUT+.t117 4.8295
R6988 VOUT+.n13 VOUT+.t72 4.8295
R6989 VOUT+.n25 VOUT+.t37 4.8295
R6990 VOUT+.n26 VOUT+.t20 4.8295
R6991 VOUT+.n28 VOUT+.t79 4.8295
R6992 VOUT+.n29 VOUT+.t60 4.8295
R6993 VOUT+.n31 VOUT+.t121 4.8295
R6994 VOUT+.n32 VOUT+.t104 4.8295
R6995 VOUT+.n34 VOUT+.t84 4.8295
R6996 VOUT+.n35 VOUT+.t66 4.8295
R6997 VOUT+.n86 VOUT+.t123 4.8295
R6998 VOUT+.n48 VOUT+.t95 4.8154
R6999 VOUT+.n49 VOUT+.t70 4.8154
R7000 VOUT+.n50 VOUT+.t110 4.8154
R7001 VOUT+.n51 VOUT+.t145 4.8154
R7002 VOUT+.n48 VOUT+.t32 4.806
R7003 VOUT+.n49 VOUT+.t150 4.806
R7004 VOUT+.n50 VOUT+.t50 4.806
R7005 VOUT+.n51 VOUT+.t87 4.806
R7006 VOUT+.n52 VOUT+.t125 4.806
R7007 VOUT+.n53 VOUT+.t105 4.806
R7008 VOUT+.n54 VOUT+.t140 4.806
R7009 VOUT+.n55 VOUT+.t36 4.806
R7010 VOUT+.n56 VOUT+.t156 4.806
R7011 VOUT+.n57 VOUT+.t53 4.806
R7012 VOUT+.n14 VOUT+.t73 4.806
R7013 VOUT+.n15 VOUT+.t116 4.806
R7014 VOUT+.n16 VOUT+.t64 4.806
R7015 VOUT+.n17 VOUT+.t154 4.806
R7016 VOUT+.n18 VOUT+.t106 4.806
R7017 VOUT+.n19 VOUT+.t143 4.806
R7018 VOUT+.n20 VOUT+.t96 4.806
R7019 VOUT+.n21 VOUT+.t42 4.806
R7020 VOUT+.n22 VOUT+.t86 4.806
R7021 VOUT+.n23 VOUT+.t34 4.806
R7022 VOUT+.n37 VOUT+.t69 4.5005
R7023 VOUT+.n38 VOUT+.t90 4.5005
R7024 VOUT+.n46 VOUT+.t80 4.5005
R7025 VOUT+.n47 VOUT+.t43 4.5005
R7026 VOUT+.n44 VOUT+.t56 4.5005
R7027 VOUT+.n45 VOUT+.t21 4.5005
R7028 VOUT+.n42 VOUT+.t98 4.5005
R7029 VOUT+.n43 VOUT+.t59 4.5005
R7030 VOUT+.n40 VOUT+.t136 4.5005
R7031 VOUT+.n41 VOUT+.t101 4.5005
R7032 VOUT+.n39 VOUT+.t30 4.5005
R7033 VOUT+.n58 VOUT+.t51 4.5005
R7034 VOUT+.n57 VOUT+.t155 4.5005
R7035 VOUT+.n56 VOUT+.t119 4.5005
R7036 VOUT+.n55 VOUT+.t139 4.5005
R7037 VOUT+.n54 VOUT+.t102 4.5005
R7038 VOUT+.n53 VOUT+.t61 4.5005
R7039 VOUT+.n52 VOUT+.t85 4.5005
R7040 VOUT+.n51 VOUT+.t45 4.5005
R7041 VOUT+.n50 VOUT+.t147 4.5005
R7042 VOUT+.n49 VOUT+.t111 4.5005
R7043 VOUT+.n48 VOUT+.t134 4.5005
R7044 VOUT+.n59 VOUT+.t130 4.5005
R7045 VOUT+.n61 VOUT+.t152 4.5005
R7046 VOUT+.n60 VOUT+.t115 4.5005
R7047 VOUT+.n62 VOUT+.t23 4.5005
R7048 VOUT+.n64 VOUT+.t47 4.5005
R7049 VOUT+.n63 VOUT+.t148 4.5005
R7050 VOUT+.n65 VOUT+.t78 4.5005
R7051 VOUT+.n67 VOUT+.t26 4.5005
R7052 VOUT+.n66 VOUT+.t132 4.5005
R7053 VOUT+.n68 VOUT+.t39 4.5005
R7054 VOUT+.n70 VOUT+.t128 4.5005
R7055 VOUT+.n69 VOUT+.t92 4.5005
R7056 VOUT+.n71 VOUT+.t71 4.5005
R7057 VOUT+.n73 VOUT+.t19 4.5005
R7058 VOUT+.n72 VOUT+.t126 4.5005
R7059 VOUT+.n74 VOUT+.t33 4.5005
R7060 VOUT+.n76 VOUT+.t122 4.5005
R7061 VOUT+.n75 VOUT+.t88 4.5005
R7062 VOUT+.n77 VOUT+.t135 4.5005
R7063 VOUT+.n79 VOUT+.t82 4.5005
R7064 VOUT+.n78 VOUT+.t48 4.5005
R7065 VOUT+.n80 VOUT+.t28 4.5005
R7066 VOUT+.n82 VOUT+.t120 4.5005
R7067 VOUT+.n81 VOUT+.t81 4.5005
R7068 VOUT+.n83 VOUT+.t129 4.5005
R7069 VOUT+.n85 VOUT+.t77 4.5005
R7070 VOUT+.n84 VOUT+.t40 4.5005
R7071 VOUT+.n11 VOUT+.t25 4.5005
R7072 VOUT+.n12 VOUT+.t124 4.5005
R7073 VOUT+.n13 VOUT+.t38 4.5005
R7074 VOUT+.n24 VOUT+.t127 4.5005
R7075 VOUT+.n23 VOUT+.t94 4.5005
R7076 VOUT+.n22 VOUT+.t54 4.5005
R7077 VOUT+.n21 VOUT+.t144 4.5005
R7078 VOUT+.n20 VOUT+.t113 4.5005
R7079 VOUT+.n19 VOUT+.t75 4.5005
R7080 VOUT+.n18 VOUT+.t24 4.5005
R7081 VOUT+.n17 VOUT+.t131 4.5005
R7082 VOUT+.n16 VOUT+.t97 4.5005
R7083 VOUT+.n15 VOUT+.t58 4.5005
R7084 VOUT+.n14 VOUT+.t149 4.5005
R7085 VOUT+.n25 VOUT+.t142 4.5005
R7086 VOUT+.n27 VOUT+.t93 4.5005
R7087 VOUT+.n26 VOUT+.t57 4.5005
R7088 VOUT+.n28 VOUT+.t41 4.5005
R7089 VOUT+.n30 VOUT+.t133 4.5005
R7090 VOUT+.n29 VOUT+.t100 4.5005
R7091 VOUT+.n31 VOUT+.t83 4.5005
R7092 VOUT+.n33 VOUT+.t31 4.5005
R7093 VOUT+.n32 VOUT+.t137 4.5005
R7094 VOUT+.n34 VOUT+.t49 4.5005
R7095 VOUT+.n36 VOUT+.t138 4.5005
R7096 VOUT+.n35 VOUT+.t103 4.5005
R7097 VOUT+.n86 VOUT+.t89 4.5005
R7098 VOUT+.n87 VOUT+.t35 4.5005
R7099 VOUT+.n88 VOUT+.t141 4.5005
R7100 VOUT+.n89 VOUT+.t107 4.5005
R7101 VOUT+.n10 VOUT+.n8 4.5005
R7102 VOUT+.n94 VOUT+.t15 3.42907
R7103 VOUT+.n94 VOUT+.t14 3.42907
R7104 VOUT+.n92 VOUT+.t13 3.42907
R7105 VOUT+.n92 VOUT+.t1 3.42907
R7106 VOUT+.n91 VOUT+.t12 3.42907
R7107 VOUT+.n91 VOUT+.t16 3.42907
R7108 VOUT+ VOUT+.n96 2.96925
R7109 VOUT+.n96 VOUT+.n95 2.03175
R7110 VOUT+.n95 VOUT+.n93 1.1255
R7111 VOUT+.n4 VOUT+.n2 0.563
R7112 VOUT+.n6 VOUT+.n4 0.563
R7113 VOUT+.n8 VOUT+.n6 0.563
R7114 VOUT+.n38 VOUT+.n37 0.3295
R7115 VOUT+.n47 VOUT+.n46 0.3295
R7116 VOUT+.n45 VOUT+.n44 0.3295
R7117 VOUT+.n43 VOUT+.n42 0.3295
R7118 VOUT+.n41 VOUT+.n40 0.3295
R7119 VOUT+.n58 VOUT+.n39 0.3295
R7120 VOUT+.n58 VOUT+.n57 0.3295
R7121 VOUT+.n57 VOUT+.n56 0.3295
R7122 VOUT+.n56 VOUT+.n55 0.3295
R7123 VOUT+.n55 VOUT+.n54 0.3295
R7124 VOUT+.n54 VOUT+.n53 0.3295
R7125 VOUT+.n53 VOUT+.n52 0.3295
R7126 VOUT+.n52 VOUT+.n51 0.3295
R7127 VOUT+.n51 VOUT+.n50 0.3295
R7128 VOUT+.n50 VOUT+.n49 0.3295
R7129 VOUT+.n49 VOUT+.n48 0.3295
R7130 VOUT+.n61 VOUT+.n59 0.3295
R7131 VOUT+.n61 VOUT+.n60 0.3295
R7132 VOUT+.n64 VOUT+.n62 0.3295
R7133 VOUT+.n64 VOUT+.n63 0.3295
R7134 VOUT+.n67 VOUT+.n65 0.3295
R7135 VOUT+.n67 VOUT+.n66 0.3295
R7136 VOUT+.n70 VOUT+.n68 0.3295
R7137 VOUT+.n70 VOUT+.n69 0.3295
R7138 VOUT+.n73 VOUT+.n71 0.3295
R7139 VOUT+.n73 VOUT+.n72 0.3295
R7140 VOUT+.n76 VOUT+.n74 0.3295
R7141 VOUT+.n76 VOUT+.n75 0.3295
R7142 VOUT+.n79 VOUT+.n77 0.3295
R7143 VOUT+.n79 VOUT+.n78 0.3295
R7144 VOUT+.n82 VOUT+.n80 0.3295
R7145 VOUT+.n82 VOUT+.n81 0.3295
R7146 VOUT+.n85 VOUT+.n83 0.3295
R7147 VOUT+.n85 VOUT+.n84 0.3295
R7148 VOUT+.n12 VOUT+.n11 0.3295
R7149 VOUT+.n24 VOUT+.n13 0.3295
R7150 VOUT+.n24 VOUT+.n23 0.3295
R7151 VOUT+.n23 VOUT+.n22 0.3295
R7152 VOUT+.n22 VOUT+.n21 0.3295
R7153 VOUT+.n21 VOUT+.n20 0.3295
R7154 VOUT+.n20 VOUT+.n19 0.3295
R7155 VOUT+.n19 VOUT+.n18 0.3295
R7156 VOUT+.n18 VOUT+.n17 0.3295
R7157 VOUT+.n17 VOUT+.n16 0.3295
R7158 VOUT+.n16 VOUT+.n15 0.3295
R7159 VOUT+.n15 VOUT+.n14 0.3295
R7160 VOUT+.n27 VOUT+.n25 0.3295
R7161 VOUT+.n27 VOUT+.n26 0.3295
R7162 VOUT+.n30 VOUT+.n28 0.3295
R7163 VOUT+.n30 VOUT+.n29 0.3295
R7164 VOUT+.n33 VOUT+.n31 0.3295
R7165 VOUT+.n33 VOUT+.n32 0.3295
R7166 VOUT+.n36 VOUT+.n34 0.3295
R7167 VOUT+.n36 VOUT+.n35 0.3295
R7168 VOUT+.n87 VOUT+.n86 0.3295
R7169 VOUT+.n88 VOUT+.n87 0.3295
R7170 VOUT+.n89 VOUT+.n88 0.3295
R7171 VOUT+.n52 VOUT+.n47 0.306
R7172 VOUT+.n53 VOUT+.n45 0.306
R7173 VOUT+.n54 VOUT+.n43 0.306
R7174 VOUT+.n55 VOUT+.n41 0.306
R7175 VOUT+.n58 VOUT+.n38 0.2825
R7176 VOUT+.n61 VOUT+.n58 0.2825
R7177 VOUT+.n64 VOUT+.n61 0.2825
R7178 VOUT+.n67 VOUT+.n64 0.2825
R7179 VOUT+.n70 VOUT+.n67 0.2825
R7180 VOUT+.n73 VOUT+.n70 0.2825
R7181 VOUT+.n76 VOUT+.n73 0.2825
R7182 VOUT+.n79 VOUT+.n76 0.2825
R7183 VOUT+.n82 VOUT+.n79 0.2825
R7184 VOUT+.n85 VOUT+.n82 0.2825
R7185 VOUT+.n24 VOUT+.n12 0.2825
R7186 VOUT+.n27 VOUT+.n24 0.2825
R7187 VOUT+.n30 VOUT+.n27 0.2825
R7188 VOUT+.n33 VOUT+.n30 0.2825
R7189 VOUT+.n36 VOUT+.n33 0.2825
R7190 VOUT+.n87 VOUT+.n36 0.2825
R7191 VOUT+.n87 VOUT+.n85 0.2825
R7192 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.t16 449.868
R7193 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.t21 449.868
R7194 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.t13 449.868
R7195 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.t17 449.868
R7196 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.n0 339.961
R7197 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.n1 339.272
R7198 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.t6 273.134
R7199 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.t14 273.134
R7200 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.t25 273.134
R7201 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.t20 273.134
R7202 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.t9 273.134
R7203 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.t18 273.134
R7204 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.t23 273.134
R7205 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.t11 273.134
R7206 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.t24 273.134
R7207 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.t12 273.134
R7208 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.t22 273.134
R7209 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.t10 273.134
R7210 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.t7 273.134
R7211 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.t15 273.134
R7212 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.t19 273.134
R7213 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.t8 273.134
R7214 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t2 184.665
R7215 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.n19 176.733
R7216 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.n18 176.733
R7217 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.n17 176.733
R7218 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.n13 176.733
R7219 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.n14 176.733
R7220 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.n15 176.733
R7221 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.n10 176.733
R7222 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.n9 176.733
R7223 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.n8 176.733
R7224 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.n4 176.733
R7225 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.n5 176.733
R7226 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.n6 176.733
R7227 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.n12 171.644
R7228 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.n21 165.8
R7229 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t1 62.0342
R7230 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.n20 56.2338
R7231 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.n16 56.2338
R7232 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.n11 56.2338
R7233 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.n7 56.2338
R7234 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t0 39.4005
R7235 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t3 39.4005
R7236 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t4 39.4005
R7237 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t5 39.4005
R7238 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb1.n23 35.662
R7239 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.n3 23.4681
R7240 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb1.n2 12.1255
R7241 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.n22 7.98488
R7242 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.n3 526.183
R7243 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.n1 514.134
R7244 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n0 360.586
R7245 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t5 303.259
R7246 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n4 210.169
R7247 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t3 174.726
R7248 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.t7 174.726
R7249 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.t4 174.726
R7250 bgr_0.V_CUR_REF_REG.t0 bgr_0.V_CUR_REF_REG.n5 153.474
R7251 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.n2 128.534
R7252 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t6 96.4005
R7253 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t1 39.4005
R7254 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t2 39.4005
R7255 bgr_0.V_p_2.n1 bgr_0.V_p_2.n2 229.562
R7256 bgr_0.V_p_2.n1 bgr_0.V_p_2.n5 228.939
R7257 bgr_0.V_p_2.n0 bgr_0.V_p_2.n4 228.939
R7258 bgr_0.V_p_2.n0 bgr_0.V_p_2.n3 228.939
R7259 bgr_0.V_p_2.n6 bgr_0.V_p_2.n1 228.938
R7260 bgr_0.V_p_2.n0 bgr_0.V_p_2.t10 98.2279
R7261 bgr_0.V_p_2.n5 bgr_0.V_p_2.t3 48.0005
R7262 bgr_0.V_p_2.n5 bgr_0.V_p_2.t5 48.0005
R7263 bgr_0.V_p_2.n4 bgr_0.V_p_2.t8 48.0005
R7264 bgr_0.V_p_2.n4 bgr_0.V_p_2.t0 48.0005
R7265 bgr_0.V_p_2.n3 bgr_0.V_p_2.t4 48.0005
R7266 bgr_0.V_p_2.n3 bgr_0.V_p_2.t6 48.0005
R7267 bgr_0.V_p_2.n2 bgr_0.V_p_2.t1 48.0005
R7268 bgr_0.V_p_2.n2 bgr_0.V_p_2.t7 48.0005
R7269 bgr_0.V_p_2.t9 bgr_0.V_p_2.n6 48.0005
R7270 bgr_0.V_p_2.n6 bgr_0.V_p_2.t2 48.0005
R7271 bgr_0.V_p_2.n1 bgr_0.V_p_2.n0 1.8755
R7272 a_6810_23838.t0 a_6810_23838.t1 178.133
R7273 a_7460_23988.t0 a_7460_23988.t1 178.133
R7274 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t13 369.534
R7275 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t12 369.534
R7276 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t29 369.534
R7277 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t17 369.534
R7278 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t21 369.534
R7279 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t20 369.534
R7280 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n6 341.397
R7281 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n9 339.272
R7282 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n7 339.272
R7283 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n12 334.772
R7284 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.t14 238.322
R7285 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.t27 238.322
R7286 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t26 192.8
R7287 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t19 192.8
R7288 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.t16 192.8
R7289 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.t23 192.8
R7290 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t22 192.8
R7291 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t24 192.8
R7292 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.t10 192.8
R7293 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.t18 192.8
R7294 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.t25 192.8
R7295 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.t11 192.8
R7296 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t15 192.8
R7297 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t28 192.8
R7298 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.n24 176.733
R7299 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.n23 176.733
R7300 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.n18 176.733
R7301 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.n19 176.733
R7302 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.n20 176.733
R7303 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.n21 176.733
R7304 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n2 171.321
R7305 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n5 168.166
R7306 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.n14 167.519
R7307 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n26 166.071
R7308 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.t6 137.48
R7309 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.t7 100.635
R7310 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n4 56.2338
R7311 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n3 56.2338
R7312 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n25 56.2338
R7313 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n22 56.2338
R7314 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n1 56.2338
R7315 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n0 56.2338
R7316 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t9 39.4005
R7317 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t1 39.4005
R7318 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t3 39.4005
R7319 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t5 39.4005
R7320 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t2 39.4005
R7321 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t4 39.4005
R7322 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t0 39.4005
R7323 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t8 39.4005
R7324 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n16 27.5005
R7325 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n13 9.53175
R7326 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n11 4.5005
R7327 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n17 2.34425
R7328 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n8 2.1255
R7329 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.n10 2.1255
R7330 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n15 1.688
R7331 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 610.534
R7332 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 610.534
R7333 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 433.8
R7334 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 433.8
R7335 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 433.8
R7336 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 433.8
R7337 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 433.8
R7338 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 433.8
R7339 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 433.8
R7340 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 433.8
R7341 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 433.8
R7342 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 433.8
R7343 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 433.8
R7344 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 433.8
R7345 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 433.8
R7346 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 433.8
R7347 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 433.8
R7348 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 433.8
R7349 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 433.8
R7350 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 433.8
R7351 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 339.836
R7352 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 339.834
R7353 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 339.272
R7354 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 287.264
R7355 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 221.293
R7356 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 176.733
R7357 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 176.733
R7358 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 176.733
R7359 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 176.733
R7360 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 176.733
R7361 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 176.733
R7362 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 176.733
R7363 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 176.733
R7364 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 176.733
R7365 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 176.733
R7366 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 176.733
R7367 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 176.733
R7368 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 176.733
R7369 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 176.733
R7370 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 176.733
R7371 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 176.733
R7372 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 117.825
R7373 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.V_tail_gate.n29 71.9693
R7374 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 65.2045
R7375 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 56.2338
R7376 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 56.2338
R7377 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 53.2453
R7378 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 52.01
R7379 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.V_tail_gate.n6 51.6642
R7380 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 39.4005
R7381 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 39.4005
R7382 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 39.4005
R7383 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 39.4005
R7384 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 39.4005
R7385 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 39.4005
R7386 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 39.4005
R7387 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 39.4005
R7388 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 16.0005
R7389 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 16.0005
R7390 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 16.0005
R7391 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 16.0005
R7392 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 0.563
R7393 two_stage_opamp_dummy_magic_0.cap_res_X.t0 two_stage_opamp_dummy_magic_0.cap_res_X.t6 50.0055
R7394 two_stage_opamp_dummy_magic_0.cap_res_X.t23 two_stage_opamp_dummy_magic_0.cap_res_X.t62 0.1603
R7395 two_stage_opamp_dummy_magic_0.cap_res_X.t46 two_stage_opamp_dummy_magic_0.cap_res_X.t87 0.1603
R7396 two_stage_opamp_dummy_magic_0.cap_res_X.t10 two_stage_opamp_dummy_magic_0.cap_res_X.t47 0.1603
R7397 two_stage_opamp_dummy_magic_0.cap_res_X.t112 two_stage_opamp_dummy_magic_0.cap_res_X.t12 0.1603
R7398 two_stage_opamp_dummy_magic_0.cap_res_X.t77 two_stage_opamp_dummy_magic_0.cap_res_X.t92 0.1603
R7399 two_stage_opamp_dummy_magic_0.cap_res_X.t114 two_stage_opamp_dummy_magic_0.cap_res_X.t77 0.1603
R7400 two_stage_opamp_dummy_magic_0.cap_res_X.t72 two_stage_opamp_dummy_magic_0.cap_res_X.t114 0.1603
R7401 two_stage_opamp_dummy_magic_0.cap_res_X.t101 two_stage_opamp_dummy_magic_0.cap_res_X.t39 0.1603
R7402 two_stage_opamp_dummy_magic_0.cap_res_X.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t101 0.1603
R7403 two_stage_opamp_dummy_magic_0.cap_res_X.t96 two_stage_opamp_dummy_magic_0.cap_res_X.t136 0.1603
R7404 two_stage_opamp_dummy_magic_0.cap_res_X.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t90 0.1603
R7405 two_stage_opamp_dummy_magic_0.cap_res_X.t88 two_stage_opamp_dummy_magic_0.cap_res_X.t49 0.1603
R7406 two_stage_opamp_dummy_magic_0.cap_res_X.t42 two_stage_opamp_dummy_magic_0.cap_res_X.t81 0.1603
R7407 two_stage_opamp_dummy_magic_0.cap_res_X.t27 two_stage_opamp_dummy_magic_0.cap_res_X.t130 0.1603
R7408 two_stage_opamp_dummy_magic_0.cap_res_X.t9 two_stage_opamp_dummy_magic_0.cap_res_X.t45 0.1603
R7409 two_stage_opamp_dummy_magic_0.cap_res_X.t134 two_stage_opamp_dummy_magic_0.cap_res_X.t95 0.1603
R7410 two_stage_opamp_dummy_magic_0.cap_res_X.t25 two_stage_opamp_dummy_magic_0.cap_res_X.t58 0.1603
R7411 two_stage_opamp_dummy_magic_0.cap_res_X.t79 two_stage_opamp_dummy_magic_0.cap_res_X.t43 0.1603
R7412 two_stage_opamp_dummy_magic_0.cap_res_X.t65 two_stage_opamp_dummy_magic_0.cap_res_X.t102 0.1603
R7413 two_stage_opamp_dummy_magic_0.cap_res_X.t118 two_stage_opamp_dummy_magic_0.cap_res_X.t83 0.1603
R7414 two_stage_opamp_dummy_magic_0.cap_res_X.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t66 0.1603
R7415 two_stage_opamp_dummy_magic_0.cap_res_X.t86 two_stage_opamp_dummy_magic_0.cap_res_X.t48 0.1603
R7416 two_stage_opamp_dummy_magic_0.cap_res_X.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t105 0.1603
R7417 two_stage_opamp_dummy_magic_0.cap_res_X.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t89 0.1603
R7418 two_stage_opamp_dummy_magic_0.cap_res_X.t109 two_stage_opamp_dummy_magic_0.cap_res_X.t4 0.1603
R7419 two_stage_opamp_dummy_magic_0.cap_res_X.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t128 0.1603
R7420 two_stage_opamp_dummy_magic_0.cap_res_X.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t111 0.1603
R7421 two_stage_opamp_dummy_magic_0.cap_res_X.t129 two_stage_opamp_dummy_magic_0.cap_res_X.t94 0.1603
R7422 two_stage_opamp_dummy_magic_0.cap_res_X.t117 two_stage_opamp_dummy_magic_0.cap_res_X.t11 0.1603
R7423 two_stage_opamp_dummy_magic_0.cap_res_X.t28 two_stage_opamp_dummy_magic_0.cap_res_X.t135 0.1603
R7424 two_stage_opamp_dummy_magic_0.cap_res_X.t16 two_stage_opamp_dummy_magic_0.cap_res_X.t50 0.1603
R7425 two_stage_opamp_dummy_magic_0.cap_res_X.t68 two_stage_opamp_dummy_magic_0.cap_res_X.t34 0.1603
R7426 two_stage_opamp_dummy_magic_0.cap_res_X.t54 two_stage_opamp_dummy_magic_0.cap_res_X.t91 0.1603
R7427 two_stage_opamp_dummy_magic_0.cap_res_X.t108 two_stage_opamp_dummy_magic_0.cap_res_X.t73 0.1603
R7428 two_stage_opamp_dummy_magic_0.cap_res_X.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t53 0.1603
R7429 two_stage_opamp_dummy_magic_0.cap_res_X.t74 two_stage_opamp_dummy_magic_0.cap_res_X.t36 0.1603
R7430 two_stage_opamp_dummy_magic_0.cap_res_X.t57 two_stage_opamp_dummy_magic_0.cap_res_X.t97 0.1603
R7431 two_stage_opamp_dummy_magic_0.cap_res_X.t116 two_stage_opamp_dummy_magic_0.cap_res_X.t78 0.1603
R7432 two_stage_opamp_dummy_magic_0.cap_res_X.t100 two_stage_opamp_dummy_magic_0.cap_res_X.t137 0.1603
R7433 two_stage_opamp_dummy_magic_0.cap_res_X.t15 two_stage_opamp_dummy_magic_0.cap_res_X.t120 0.1603
R7434 two_stage_opamp_dummy_magic_0.cap_res_X.t8 two_stage_opamp_dummy_magic_0.cap_res_X.t84 0.1603
R7435 two_stage_opamp_dummy_magic_0.cap_res_X.t99 two_stage_opamp_dummy_magic_0.cap_res_X.t41 0.1603
R7436 two_stage_opamp_dummy_magic_0.cap_res_X.t60 two_stage_opamp_dummy_magic_0.cap_res_X.t93 0.1603
R7437 two_stage_opamp_dummy_magic_0.cap_res_X.t26 two_stage_opamp_dummy_magic_0.cap_res_X.t3 0.1603
R7438 two_stage_opamp_dummy_magic_0.cap_res_X.t133 two_stage_opamp_dummy_magic_0.cap_res_X.t51 0.1603
R7439 two_stage_opamp_dummy_magic_0.cap_res_X.t82 two_stage_opamp_dummy_magic_0.cap_res_X.t14 0.1603
R7440 two_stage_opamp_dummy_magic_0.cap_res_X.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t61 0.1603
R7441 two_stage_opamp_dummy_magic_0.cap_res_X.t13 two_stage_opamp_dummy_magic_0.cap_res_X.t115 0.1603
R7442 two_stage_opamp_dummy_magic_0.cap_res_X.t103 two_stage_opamp_dummy_magic_0.cap_res_X.t71 0.1603
R7443 two_stage_opamp_dummy_magic_0.cap_res_X.t63 two_stage_opamp_dummy_magic_0.cap_res_X.t123 0.1603
R7444 two_stage_opamp_dummy_magic_0.cap_res_X.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t85 0.1603
R7445 two_stage_opamp_dummy_magic_0.cap_res_X.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t40 0.1603
R7446 two_stage_opamp_dummy_magic_0.cap_res_X.t21 two_stage_opamp_dummy_magic_0.cap_res_X.t113 0.1603
R7447 two_stage_opamp_dummy_magic_0.cap_res_X.t56 two_stage_opamp_dummy_magic_0.cap_res_X.t21 0.1603
R7448 two_stage_opamp_dummy_magic_0.cap_res_X.t18 two_stage_opamp_dummy_magic_0.cap_res_X.t56 0.1603
R7449 two_stage_opamp_dummy_magic_0.cap_res_X.t98 two_stage_opamp_dummy_magic_0.cap_res_X.t55 0.1603
R7450 two_stage_opamp_dummy_magic_0.cap_res_X.t59 two_stage_opamp_dummy_magic_0.cap_res_X.t98 0.1603
R7451 two_stage_opamp_dummy_magic_0.cap_res_X.t6 two_stage_opamp_dummy_magic_0.cap_res_X.t59 0.1603
R7452 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t125 0.159278
R7453 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t7 0.159278
R7454 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t107 0.159278
R7455 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t70 0.159278
R7456 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t32 0.159278
R7457 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t52 0.159278
R7458 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t67 0.159278
R7459 two_stage_opamp_dummy_magic_0.cap_res_X.t30 two_stage_opamp_dummy_magic_0.cap_res_X.n9 0.159278
R7460 two_stage_opamp_dummy_magic_0.cap_res_X.t64 two_stage_opamp_dummy_magic_0.cap_res_X.n10 0.159278
R7461 two_stage_opamp_dummy_magic_0.cap_res_X.t24 two_stage_opamp_dummy_magic_0.cap_res_X.n11 0.159278
R7462 two_stage_opamp_dummy_magic_0.cap_res_X.t126 two_stage_opamp_dummy_magic_0.cap_res_X.n12 0.159278
R7463 two_stage_opamp_dummy_magic_0.cap_res_X.t19 two_stage_opamp_dummy_magic_0.cap_res_X.n13 0.159278
R7464 two_stage_opamp_dummy_magic_0.cap_res_X.t122 two_stage_opamp_dummy_magic_0.cap_res_X.n14 0.159278
R7465 two_stage_opamp_dummy_magic_0.cap_res_X.t80 two_stage_opamp_dummy_magic_0.cap_res_X.n15 0.159278
R7466 two_stage_opamp_dummy_magic_0.cap_res_X.t37 two_stage_opamp_dummy_magic_0.cap_res_X.n16 0.159278
R7467 two_stage_opamp_dummy_magic_0.cap_res_X.t75 two_stage_opamp_dummy_magic_0.cap_res_X.n17 0.159278
R7468 two_stage_opamp_dummy_magic_0.cap_res_X.t35 two_stage_opamp_dummy_magic_0.cap_res_X.n18 0.159278
R7469 two_stage_opamp_dummy_magic_0.cap_res_X.t138 two_stage_opamp_dummy_magic_0.cap_res_X.n19 0.159278
R7470 two_stage_opamp_dummy_magic_0.cap_res_X.t29 two_stage_opamp_dummy_magic_0.cap_res_X.n20 0.159278
R7471 two_stage_opamp_dummy_magic_0.cap_res_X.t131 two_stage_opamp_dummy_magic_0.cap_res_X.n21 0.159278
R7472 two_stage_opamp_dummy_magic_0.cap_res_X.t110 two_stage_opamp_dummy_magic_0.cap_res_X.n22 0.159278
R7473 two_stage_opamp_dummy_magic_0.cap_res_X.t5 two_stage_opamp_dummy_magic_0.cap_res_X.n23 0.159278
R7474 two_stage_opamp_dummy_magic_0.cap_res_X.t106 two_stage_opamp_dummy_magic_0.cap_res_X.n24 0.159278
R7475 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t104 0.159278
R7476 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t1 0.159278
R7477 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t121 0.159278
R7478 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.t17 0.159278
R7479 two_stage_opamp_dummy_magic_0.cap_res_X.t67 two_stage_opamp_dummy_magic_0.cap_res_X.t88 0.137822
R7480 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t127 0.1368
R7481 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t42 0.1368
R7482 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t27 0.1368
R7483 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t9 0.1368
R7484 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t134 0.1368
R7485 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t25 0.1368
R7486 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t79 0.1368
R7487 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t65 0.1368
R7488 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t118 0.1368
R7489 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t31 0.1368
R7490 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t86 0.1368
R7491 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t69 0.1368
R7492 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t124 0.1368
R7493 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t109 0.1368
R7494 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t22 0.1368
R7495 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t76 0.1368
R7496 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t129 0.1368
R7497 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t117 0.1368
R7498 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t28 0.1368
R7499 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t16 0.1368
R7500 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t68 0.1368
R7501 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t54 0.1368
R7502 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t108 0.1368
R7503 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t20 0.1368
R7504 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t74 0.1368
R7505 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t57 0.1368
R7506 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t116 0.1368
R7507 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t100 0.1368
R7508 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t15 0.1368
R7509 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.t119 0.1368
R7510 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.t132 0.1368
R7511 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t8 0.114322
R7512 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.n29 0.1133
R7513 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.n30 0.1133
R7514 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.n31 0.1133
R7515 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.n32 0.1133
R7516 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.n33 0.1133
R7517 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.n0 0.1133
R7518 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.n1 0.1133
R7519 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.n2 0.1133
R7520 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.n3 0.1133
R7521 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.n4 0.1133
R7522 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.n5 0.1133
R7523 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.n6 0.1133
R7524 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.n7 0.1133
R7525 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.n8 0.1133
R7526 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.n25 0.1133
R7527 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.n26 0.1133
R7528 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.n27 0.1133
R7529 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n28 0.1133
R7530 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n34 0.1133
R7531 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t23 0.00152174
R7532 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t46 0.00152174
R7533 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t10 0.00152174
R7534 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t112 0.00152174
R7535 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t72 0.00152174
R7536 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t96 0.00152174
R7537 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t99 0.00152174
R7538 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.t60 0.00152174
R7539 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.t26 0.00152174
R7540 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.t133 0.00152174
R7541 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.t82 0.00152174
R7542 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.t44 0.00152174
R7543 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.t13 0.00152174
R7544 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.t103 0.00152174
R7545 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.t63 0.00152174
R7546 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.t33 0.00152174
R7547 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.t30 0.00152174
R7548 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t64 0.00152174
R7549 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t24 0.00152174
R7550 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t126 0.00152174
R7551 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t19 0.00152174
R7552 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t122 0.00152174
R7553 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t80 0.00152174
R7554 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t37 0.00152174
R7555 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t75 0.00152174
R7556 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t35 0.00152174
R7557 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t138 0.00152174
R7558 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t29 0.00152174
R7559 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t131 0.00152174
R7560 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t110 0.00152174
R7561 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t5 0.00152174
R7562 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t106 0.00152174
R7563 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t2 0.00152174
R7564 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t38 0.00152174
R7565 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t18 0.00152174
R7566 two_stage_opamp_dummy_magic_0.cap_res_X.t55 two_stage_opamp_dummy_magic_0.cap_res_X.n35 0.00152174
R7567 bgr_0.cap_res1.t0 bgr_0.cap_res1.t10 121.245
R7568 bgr_0.cap_res1.t16 bgr_0.cap_res1.t19 0.1603
R7569 bgr_0.cap_res1.t9 bgr_0.cap_res1.t15 0.1603
R7570 bgr_0.cap_res1.t14 bgr_0.cap_res1.t18 0.1603
R7571 bgr_0.cap_res1.t7 bgr_0.cap_res1.t13 0.1603
R7572 bgr_0.cap_res1.t1 bgr_0.cap_res1.t6 0.1603
R7573 bgr_0.cap_res1.n1 bgr_0.cap_res1.t17 0.159278
R7574 bgr_0.cap_res1.n2 bgr_0.cap_res1.t2 0.159278
R7575 bgr_0.cap_res1.n3 bgr_0.cap_res1.t8 0.159278
R7576 bgr_0.cap_res1.n4 bgr_0.cap_res1.t3 0.159278
R7577 bgr_0.cap_res1.n4 bgr_0.cap_res1.t16 0.1368
R7578 bgr_0.cap_res1.n4 bgr_0.cap_res1.t12 0.1368
R7579 bgr_0.cap_res1.n3 bgr_0.cap_res1.t9 0.1368
R7580 bgr_0.cap_res1.n3 bgr_0.cap_res1.t5 0.1368
R7581 bgr_0.cap_res1.n2 bgr_0.cap_res1.t14 0.1368
R7582 bgr_0.cap_res1.n2 bgr_0.cap_res1.t11 0.1368
R7583 bgr_0.cap_res1.n1 bgr_0.cap_res1.t7 0.1368
R7584 bgr_0.cap_res1.n1 bgr_0.cap_res1.t4 0.1368
R7585 bgr_0.cap_res1.n0 bgr_0.cap_res1.t1 0.1368
R7586 bgr_0.cap_res1.n0 bgr_0.cap_res1.t20 0.1368
R7587 bgr_0.cap_res1.t17 bgr_0.cap_res1.n0 0.00152174
R7588 bgr_0.cap_res1.t2 bgr_0.cap_res1.n1 0.00152174
R7589 bgr_0.cap_res1.t8 bgr_0.cap_res1.n2 0.00152174
R7590 bgr_0.cap_res1.t3 bgr_0.cap_res1.n3 0.00152174
R7591 bgr_0.cap_res1.t10 bgr_0.cap_res1.n4 0.00152174
R7592 bgr_0.V_mir2.n20 bgr_0.V_mir2.n19 325.473
R7593 bgr_0.V_mir2.n13 bgr_0.V_mir2.n12 325.473
R7594 bgr_0.V_mir2.n8 bgr_0.V_mir2.n7 325.473
R7595 bgr_0.V_mir2.n16 bgr_0.V_mir2.t21 310.488
R7596 bgr_0.V_mir2.n9 bgr_0.V_mir2.t22 310.488
R7597 bgr_0.V_mir2.n4 bgr_0.V_mir2.t20 310.488
R7598 bgr_0.V_mir2.n2 bgr_0.V_mir2.t2 278.312
R7599 bgr_0.V_mir2.n2 bgr_0.V_mir2.n1 228.939
R7600 bgr_0.V_mir2.n3 bgr_0.V_mir2.n0 224.439
R7601 bgr_0.V_mir2.n18 bgr_0.V_mir2.t15 184.097
R7602 bgr_0.V_mir2.n11 bgr_0.V_mir2.t13 184.097
R7603 bgr_0.V_mir2.n6 bgr_0.V_mir2.t5 184.097
R7604 bgr_0.V_mir2.n17 bgr_0.V_mir2.n16 167.094
R7605 bgr_0.V_mir2.n10 bgr_0.V_mir2.n9 167.094
R7606 bgr_0.V_mir2.n5 bgr_0.V_mir2.n4 167.094
R7607 bgr_0.V_mir2.n13 bgr_0.V_mir2.n11 152
R7608 bgr_0.V_mir2.n8 bgr_0.V_mir2.n6 152
R7609 bgr_0.V_mir2.n19 bgr_0.V_mir2.n18 152
R7610 bgr_0.V_mir2.n16 bgr_0.V_mir2.t19 120.501
R7611 bgr_0.V_mir2.n17 bgr_0.V_mir2.t11 120.501
R7612 bgr_0.V_mir2.n9 bgr_0.V_mir2.t18 120.501
R7613 bgr_0.V_mir2.n10 bgr_0.V_mir2.t7 120.501
R7614 bgr_0.V_mir2.n4 bgr_0.V_mir2.t17 120.501
R7615 bgr_0.V_mir2.n5 bgr_0.V_mir2.t9 120.501
R7616 bgr_0.V_mir2.n1 bgr_0.V_mir2.t4 48.0005
R7617 bgr_0.V_mir2.n1 bgr_0.V_mir2.t0 48.0005
R7618 bgr_0.V_mir2.n0 bgr_0.V_mir2.t3 48.0005
R7619 bgr_0.V_mir2.n0 bgr_0.V_mir2.t1 48.0005
R7620 bgr_0.V_mir2.n18 bgr_0.V_mir2.n17 40.7027
R7621 bgr_0.V_mir2.n11 bgr_0.V_mir2.n10 40.7027
R7622 bgr_0.V_mir2.n6 bgr_0.V_mir2.n5 40.7027
R7623 bgr_0.V_mir2.n12 bgr_0.V_mir2.t8 39.4005
R7624 bgr_0.V_mir2.n12 bgr_0.V_mir2.t14 39.4005
R7625 bgr_0.V_mir2.n7 bgr_0.V_mir2.t10 39.4005
R7626 bgr_0.V_mir2.n7 bgr_0.V_mir2.t6 39.4005
R7627 bgr_0.V_mir2.n20 bgr_0.V_mir2.t12 39.4005
R7628 bgr_0.V_mir2.t16 bgr_0.V_mir2.n20 39.4005
R7629 bgr_0.V_mir2.n14 bgr_0.V_mir2.n13 15.8005
R7630 bgr_0.V_mir2.n14 bgr_0.V_mir2.n8 15.8005
R7631 bgr_0.V_mir2.n19 bgr_0.V_mir2.n15 9.3005
R7632 bgr_0.V_mir2.n3 bgr_0.V_mir2.n2 5.8755
R7633 bgr_0.V_mir2.n15 bgr_0.V_mir2.n14 4.5005
R7634 bgr_0.V_mir2.n15 bgr_0.V_mir2.n3 0.78175
R7635 bgr_0.Vin-.n7 bgr_0.Vin-.t12 688.859
R7636 bgr_0.Vin-.n9 bgr_0.Vin-.n8 514.134
R7637 bgr_0.Vin-.n6 bgr_0.Vin-.n5 351.522
R7638 bgr_0.Vin-.n11 bgr_0.Vin-.n10 213.4
R7639 bgr_0.Vin-.n7 bgr_0.Vin-.t8 174.726
R7640 bgr_0.Vin-.n8 bgr_0.Vin-.t10 174.726
R7641 bgr_0.Vin-.n9 bgr_0.Vin-.t9 174.726
R7642 bgr_0.Vin-.n10 bgr_0.Vin-.t11 174.726
R7643 bgr_0.Vin-.n4 bgr_0.Vin-.n2 173.029
R7644 bgr_0.Vin-.n4 bgr_0.Vin-.n3 168.654
R7645 bgr_0.Vin-.n8 bgr_0.Vin-.n7 128.534
R7646 bgr_0.Vin-.n10 bgr_0.Vin-.n9 128.534
R7647 bgr_0.Vin-.n12 bgr_0.Vin-.t0 119.099
R7648 bgr_0.Vin-.n16 bgr_0.Vin-.n15 83.5719
R7649 bgr_0.Vin-.n1 bgr_0.Vin-.n0 83.5719
R7650 bgr_0.Vin-.n19 bgr_0.Vin-.n1 73.8495
R7651 bgr_0.Vin-.t3 bgr_0.Vin-.n14 65.0341
R7652 bgr_0.Vin-.n5 bgr_0.Vin-.t2 39.4005
R7653 bgr_0.Vin-.n5 bgr_0.Vin-.t1 39.4005
R7654 bgr_0.Vin-.n13 bgr_0.Vin-.n12 28.813
R7655 bgr_0.Vin-.n15 bgr_0.Vin-.n1 26.074
R7656 bgr_0.Vin-.n12 bgr_0.Vin-.n11 16.188
R7657 bgr_0.Vin-.n3 bgr_0.Vin-.t4 13.1338
R7658 bgr_0.Vin-.n3 bgr_0.Vin-.t6 13.1338
R7659 bgr_0.Vin-.n2 bgr_0.Vin-.t7 13.1338
R7660 bgr_0.Vin-.n2 bgr_0.Vin-.t5 13.1338
R7661 bgr_0.Vin-.n11 bgr_0.Vin-.n6 11.2193
R7662 bgr_0.Vin-.n6 bgr_0.Vin-.n4 3.8755
R7663 bgr_0.Vin-.n16 bgr_0.Vin-.n14 1.56483
R7664 bgr_0.Vin-.n18 bgr_0.Vin-.n17 1.5505
R7665 bgr_0.Vin-.n17 bgr_0.Vin-.n0 0.885803
R7666 bgr_0.Vin-.n17 bgr_0.Vin-.n16 0.77514
R7667 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_0.Vin-.n0 0.756696
R7668 bgr_0.Vin-.n19 bgr_0.Vin-.n18 0.711459
R7669 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_0.Vin-.n19 0.576566
R7670 bgr_0.Vin-.n14 bgr_0.Vin-.n13 0.531499
R7671 bgr_0.Vin-.n15 bgr_0.Vin-.t3 0.290206
R7672 bgr_0.Vin-.n18 bgr_0.Vin-.n13 0.00817857
R7673 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.n0 219.928
R7674 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t3 16.0005
R7675 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t2 16.0005
R7676 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.t0 9.6005
R7677 two_stage_opamp_dummy_magic_0.V_p_mir.t1 two_stage_opamp_dummy_magic_0.V_p_mir.n1 9.6005
R7678 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 525.38
R7679 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 525.38
R7680 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 366.856
R7681 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 366.856
R7682 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 281.168
R7683 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 281.168
R7684 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 281.168
R7685 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 281.168
R7686 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 244.214
R7687 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 244.214
R7688 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 166.03
R7689 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 166.03
R7690 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 117.974
R7691 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 117.849
R7692 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 85.6894
R7693 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 85.6894
R7694 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 36.813
R7695 bgr_0.V_p_1.n1 bgr_0.V_p_1.n5 229.562
R7696 bgr_0.V_p_1.n1 bgr_0.V_p_1.n4 228.939
R7697 bgr_0.V_p_1.n0 bgr_0.V_p_1.n3 228.939
R7698 bgr_0.V_p_1.n0 bgr_0.V_p_1.n2 228.939
R7699 bgr_0.V_p_1.n6 bgr_0.V_p_1.n1 228.938
R7700 bgr_0.V_p_1.n0 bgr_0.V_p_1.t10 98.2279
R7701 bgr_0.V_p_1.n5 bgr_0.V_p_1.t7 48.0005
R7702 bgr_0.V_p_1.n5 bgr_0.V_p_1.t0 48.0005
R7703 bgr_0.V_p_1.n4 bgr_0.V_p_1.t9 48.0005
R7704 bgr_0.V_p_1.n4 bgr_0.V_p_1.t2 48.0005
R7705 bgr_0.V_p_1.n3 bgr_0.V_p_1.t3 48.0005
R7706 bgr_0.V_p_1.n3 bgr_0.V_p_1.t5 48.0005
R7707 bgr_0.V_p_1.n2 bgr_0.V_p_1.t8 48.0005
R7708 bgr_0.V_p_1.n2 bgr_0.V_p_1.t1 48.0005
R7709 bgr_0.V_p_1.t4 bgr_0.V_p_1.n6 48.0005
R7710 bgr_0.V_p_1.n6 bgr_0.V_p_1.t6 48.0005
R7711 bgr_0.V_p_1.n1 bgr_0.V_p_1.n0 1.8755
R7712 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 144.827
R7713 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 134.577
R7714 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 120.66
R7715 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 97.4009
R7716 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 96.8384
R7717 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 96.8384
R7718 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 96.8384
R7719 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 96.8384
R7720 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 37.4067
R7721 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 35.2505
R7722 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 24.0005
R7723 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 24.0005
R7724 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 24.0005
R7725 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 24.0005
R7726 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 8.0005
R7727 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 8.0005
R7728 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 8.0005
R7729 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 8.0005
R7730 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 8.0005
R7731 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 8.0005
R7732 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 8.0005
R7733 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 8.0005
R7734 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 8.0005
R7735 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 8.0005
R7736 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 5.938
R7737 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 0.563
R7738 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 0.563
R7739 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 0.563
R7740 bgr_0.V_CMFB_S2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n13 0.047375
R7741 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n3 630.827
R7742 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n8 630.264
R7743 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n6 630.264
R7744 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n4 630.264
R7745 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n13 627.784
R7746 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n0 627.784
R7747 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.n2 627.168
R7748 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n16 626.534
R7749 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n14 626.534
R7750 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.n18 626.534
R7751 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n1 622.034
R7752 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.t12 78.8005
R7753 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.t17 78.8005
R7754 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t9 78.8005
R7755 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t14 78.8005
R7756 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t16 78.8005
R7757 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t20 78.8005
R7758 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t15 78.8005
R7759 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t10 78.8005
R7760 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.t19 78.8005
R7761 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.t5 78.8005
R7762 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t3 78.8005
R7763 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t7 78.8005
R7764 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t0 78.8005
R7765 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t2 78.8005
R7766 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.t1 78.8005
R7767 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.t8 78.8005
R7768 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t4 78.8005
R7769 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t6 78.8005
R7770 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t21 78.8005
R7771 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t11 78.8005
R7772 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.t13 78.8005
R7773 two_stage_opamp_dummy_magic_0.V_err_p.t18 two_stage_opamp_dummy_magic_0.V_err_p.n19 78.8005
R7774 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.n9 5.0005
R7775 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n11 4.5005
R7776 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n10 1.60845
R7777 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n15 1.2505
R7778 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n17 1.2505
R7779 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n12 1.2505
R7780 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n5 0.563
R7781 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n7 0.563
R7782 a_14560_5068.t0 a_14560_5068.t1 294.339
R7783 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.t6 327.623
R7784 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.t4 326.365
R7785 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t10 168.701
R7786 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t9 168.701
R7787 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.n1 167.05
R7788 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.n7 165.8
R7789 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.n5 165.8
R7790 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.n2 165.8
R7791 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.t13 157.989
R7792 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.t7 157.989
R7793 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.t8 157.989
R7794 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.t12 157.989
R7795 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.t5 157.989
R7796 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.t11 157.989
R7797 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.t1 117.591
R7798 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t2 117.591
R7799 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t3 108.424
R7800 two_stage_opamp_dummy_magic_0.V_tot.t0 two_stage_opamp_dummy_magic_0.V_tot.n11 108.424
R7801 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n0 37.5496
R7802 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.n10 37.1121
R7803 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n9 10.6255
R7804 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.n8 2.063
R7805 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.n6 1.26612
R7806 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.n3 1.15363
R7807 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.n4 1.12862
R7808 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.n9 114.719
R7809 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n4 114.719
R7810 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n5 114.156
R7811 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.n7 114.156
R7812 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n0 113.081
R7813 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n15 111.769
R7814 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n17 111.769
R7815 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VD1.n19 111.769
R7816 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n1 111.769
R7817 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n3 109.656
R7818 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n12 107.269
R7819 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t2 16.0005
R7820 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t7 16.0005
R7821 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.t15 16.0005
R7822 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.t19 16.0005
R7823 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t11 16.0005
R7824 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t12 16.0005
R7825 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.t21 16.0005
R7826 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.t17 16.0005
R7827 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t14 16.0005
R7828 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t20 16.0005
R7829 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t16 16.0005
R7830 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t0 16.0005
R7831 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t13 16.0005
R7832 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t18 16.0005
R7833 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.t1 16.0005
R7834 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.t6 16.0005
R7835 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t3 16.0005
R7836 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t5 16.0005
R7837 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t4 16.0005
R7838 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t9 16.0005
R7839 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t10 16.0005
R7840 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t8 16.0005
R7841 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n13 4.5005
R7842 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n10 4.5005
R7843 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n14 3.563
R7844 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n16 1.313
R7845 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n2 1.2505
R7846 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VD1.n18 1.2505
R7847 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.n8 0.563
R7848 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.n6 0.563
R7849 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n11 0.21925
R7850 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 344.837
R7851 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 344.274
R7852 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 292.5
R7853 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 206.052
R7854 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 205.488
R7855 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 205.488
R7856 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 205.488
R7857 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 205.488
R7858 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 122.504
R7859 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 52.3363
R7860 bgr_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 52.1563
R7861 bgr_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 42.313
R7862 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 39.4005
R7863 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 39.4005
R7864 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 39.4005
R7865 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 39.4005
R7866 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 39.4005
R7867 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 39.4005
R7868 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 19.7005
R7869 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 19.7005
R7870 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 19.7005
R7871 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 19.7005
R7872 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 19.7005
R7873 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 19.7005
R7874 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 19.7005
R7875 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 19.7005
R7876 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 19.7005
R7877 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 19.7005
R7878 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 6.21925
R7879 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 0.563
R7880 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 0.563
R7881 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 0.563
R7882 two_stage_opamp_dummy_magic_0.V_source.n9 two_stage_opamp_dummy_magic_0.V_source.t23 206.47
R7883 two_stage_opamp_dummy_magic_0.V_source.n28 two_stage_opamp_dummy_magic_0.V_source.n26 118.168
R7884 two_stage_opamp_dummy_magic_0.V_source.n21 two_stage_opamp_dummy_magic_0.V_source.n19 117.831
R7885 two_stage_opamp_dummy_magic_0.V_source.n34 two_stage_opamp_dummy_magic_0.V_source.n33 117.269
R7886 two_stage_opamp_dummy_magic_0.V_source.n32 two_stage_opamp_dummy_magic_0.V_source.n31 117.269
R7887 two_stage_opamp_dummy_magic_0.V_source.n30 two_stage_opamp_dummy_magic_0.V_source.n29 117.269
R7888 two_stage_opamp_dummy_magic_0.V_source.n28 two_stage_opamp_dummy_magic_0.V_source.n27 117.269
R7889 two_stage_opamp_dummy_magic_0.V_source.n25 two_stage_opamp_dummy_magic_0.V_source.n24 117.269
R7890 two_stage_opamp_dummy_magic_0.V_source.n23 two_stage_opamp_dummy_magic_0.V_source.n22 117.269
R7891 two_stage_opamp_dummy_magic_0.V_source.n21 two_stage_opamp_dummy_magic_0.V_source.n20 117.269
R7892 two_stage_opamp_dummy_magic_0.V_source.n36 two_stage_opamp_dummy_magic_0.V_source.n18 113.136
R7893 two_stage_opamp_dummy_magic_0.V_source.n2 two_stage_opamp_dummy_magic_0.V_source.n0 99.7407
R7894 two_stage_opamp_dummy_magic_0.V_source.n5 two_stage_opamp_dummy_magic_0.V_source.n3 99.647
R7895 two_stage_opamp_dummy_magic_0.V_source.n16 two_stage_opamp_dummy_magic_0.V_source.n15 99.0845
R7896 two_stage_opamp_dummy_magic_0.V_source.n14 two_stage_opamp_dummy_magic_0.V_source.n13 99.0845
R7897 two_stage_opamp_dummy_magic_0.V_source.n12 two_stage_opamp_dummy_magic_0.V_source.n11 99.0845
R7898 two_stage_opamp_dummy_magic_0.V_source.n7 two_stage_opamp_dummy_magic_0.V_source.n6 99.0845
R7899 two_stage_opamp_dummy_magic_0.V_source.n5 two_stage_opamp_dummy_magic_0.V_source.n4 99.0845
R7900 two_stage_opamp_dummy_magic_0.V_source.n2 two_stage_opamp_dummy_magic_0.V_source.n1 99.0845
R7901 two_stage_opamp_dummy_magic_0.V_source.n38 two_stage_opamp_dummy_magic_0.V_source.n37 94.5857
R7902 two_stage_opamp_dummy_magic_0.V_source.n9 two_stage_opamp_dummy_magic_0.V_source.n8 94.5845
R7903 two_stage_opamp_dummy_magic_0.V_source.n33 two_stage_opamp_dummy_magic_0.V_source.t35 16.0005
R7904 two_stage_opamp_dummy_magic_0.V_source.n33 two_stage_opamp_dummy_magic_0.V_source.t37 16.0005
R7905 two_stage_opamp_dummy_magic_0.V_source.n31 two_stage_opamp_dummy_magic_0.V_source.t0 16.0005
R7906 two_stage_opamp_dummy_magic_0.V_source.n31 two_stage_opamp_dummy_magic_0.V_source.t24 16.0005
R7907 two_stage_opamp_dummy_magic_0.V_source.n29 two_stage_opamp_dummy_magic_0.V_source.t26 16.0005
R7908 two_stage_opamp_dummy_magic_0.V_source.n29 two_stage_opamp_dummy_magic_0.V_source.t2 16.0005
R7909 two_stage_opamp_dummy_magic_0.V_source.n27 two_stage_opamp_dummy_magic_0.V_source.t29 16.0005
R7910 two_stage_opamp_dummy_magic_0.V_source.n27 two_stage_opamp_dummy_magic_0.V_source.t40 16.0005
R7911 two_stage_opamp_dummy_magic_0.V_source.n26 two_stage_opamp_dummy_magic_0.V_source.t33 16.0005
R7912 two_stage_opamp_dummy_magic_0.V_source.n26 two_stage_opamp_dummy_magic_0.V_source.t39 16.0005
R7913 two_stage_opamp_dummy_magic_0.V_source.n24 two_stage_opamp_dummy_magic_0.V_source.t32 16.0005
R7914 two_stage_opamp_dummy_magic_0.V_source.n24 two_stage_opamp_dummy_magic_0.V_source.t27 16.0005
R7915 two_stage_opamp_dummy_magic_0.V_source.n22 two_stage_opamp_dummy_magic_0.V_source.t36 16.0005
R7916 two_stage_opamp_dummy_magic_0.V_source.n22 two_stage_opamp_dummy_magic_0.V_source.t1 16.0005
R7917 two_stage_opamp_dummy_magic_0.V_source.n20 two_stage_opamp_dummy_magic_0.V_source.t22 16.0005
R7918 two_stage_opamp_dummy_magic_0.V_source.n20 two_stage_opamp_dummy_magic_0.V_source.t30 16.0005
R7919 two_stage_opamp_dummy_magic_0.V_source.n19 two_stage_opamp_dummy_magic_0.V_source.t21 16.0005
R7920 two_stage_opamp_dummy_magic_0.V_source.n19 two_stage_opamp_dummy_magic_0.V_source.t25 16.0005
R7921 two_stage_opamp_dummy_magic_0.V_source.n18 two_stage_opamp_dummy_magic_0.V_source.t34 16.0005
R7922 two_stage_opamp_dummy_magic_0.V_source.n18 two_stage_opamp_dummy_magic_0.V_source.t28 16.0005
R7923 two_stage_opamp_dummy_magic_0.V_source.n15 two_stage_opamp_dummy_magic_0.V_source.t17 9.6005
R7924 two_stage_opamp_dummy_magic_0.V_source.n15 two_stage_opamp_dummy_magic_0.V_source.t7 9.6005
R7925 two_stage_opamp_dummy_magic_0.V_source.n13 two_stage_opamp_dummy_magic_0.V_source.t15 9.6005
R7926 two_stage_opamp_dummy_magic_0.V_source.n13 two_stage_opamp_dummy_magic_0.V_source.t5 9.6005
R7927 two_stage_opamp_dummy_magic_0.V_source.n11 two_stage_opamp_dummy_magic_0.V_source.t11 9.6005
R7928 two_stage_opamp_dummy_magic_0.V_source.n11 two_stage_opamp_dummy_magic_0.V_source.t3 9.6005
R7929 two_stage_opamp_dummy_magic_0.V_source.n8 two_stage_opamp_dummy_magic_0.V_source.t14 9.6005
R7930 two_stage_opamp_dummy_magic_0.V_source.n8 two_stage_opamp_dummy_magic_0.V_source.t4 9.6005
R7931 two_stage_opamp_dummy_magic_0.V_source.n6 two_stage_opamp_dummy_magic_0.V_source.t10 9.6005
R7932 two_stage_opamp_dummy_magic_0.V_source.n6 two_stage_opamp_dummy_magic_0.V_source.t18 9.6005
R7933 two_stage_opamp_dummy_magic_0.V_source.n4 two_stage_opamp_dummy_magic_0.V_source.t8 9.6005
R7934 two_stage_opamp_dummy_magic_0.V_source.n4 two_stage_opamp_dummy_magic_0.V_source.t16 9.6005
R7935 two_stage_opamp_dummy_magic_0.V_source.n3 two_stage_opamp_dummy_magic_0.V_source.t6 9.6005
R7936 two_stage_opamp_dummy_magic_0.V_source.n3 two_stage_opamp_dummy_magic_0.V_source.t12 9.6005
R7937 two_stage_opamp_dummy_magic_0.V_source.n1 two_stage_opamp_dummy_magic_0.V_source.t19 9.6005
R7938 two_stage_opamp_dummy_magic_0.V_source.n1 two_stage_opamp_dummy_magic_0.V_source.t13 9.6005
R7939 two_stage_opamp_dummy_magic_0.V_source.n0 two_stage_opamp_dummy_magic_0.V_source.t31 9.6005
R7940 two_stage_opamp_dummy_magic_0.V_source.n0 two_stage_opamp_dummy_magic_0.V_source.t38 9.6005
R7941 two_stage_opamp_dummy_magic_0.V_source.t20 two_stage_opamp_dummy_magic_0.V_source.n38 9.6005
R7942 two_stage_opamp_dummy_magic_0.V_source.n38 two_stage_opamp_dummy_magic_0.V_source.t9 9.6005
R7943 two_stage_opamp_dummy_magic_0.V_source.n10 two_stage_opamp_dummy_magic_0.V_source.n9 4.5005
R7944 two_stage_opamp_dummy_magic_0.V_source.n36 two_stage_opamp_dummy_magic_0.V_source.n35 4.5005
R7945 two_stage_opamp_dummy_magic_0.V_source.n37 two_stage_opamp_dummy_magic_0.V_source.n17 4.5005
R7946 two_stage_opamp_dummy_magic_0.V_source.n35 two_stage_opamp_dummy_magic_0.V_source.n34 3.65675
R7947 two_stage_opamp_dummy_magic_0.V_source.n37 two_stage_opamp_dummy_magic_0.V_source.n36 1.28175
R7948 two_stage_opamp_dummy_magic_0.V_source.n7 two_stage_opamp_dummy_magic_0.V_source.n5 0.563
R7949 two_stage_opamp_dummy_magic_0.V_source.n10 two_stage_opamp_dummy_magic_0.V_source.n7 0.563
R7950 two_stage_opamp_dummy_magic_0.V_source.n12 two_stage_opamp_dummy_magic_0.V_source.n10 0.563
R7951 two_stage_opamp_dummy_magic_0.V_source.n14 two_stage_opamp_dummy_magic_0.V_source.n12 0.563
R7952 two_stage_opamp_dummy_magic_0.V_source.n16 two_stage_opamp_dummy_magic_0.V_source.n14 0.563
R7953 two_stage_opamp_dummy_magic_0.V_source.n17 two_stage_opamp_dummy_magic_0.V_source.n16 0.563
R7954 two_stage_opamp_dummy_magic_0.V_source.n17 two_stage_opamp_dummy_magic_0.V_source.n2 0.563
R7955 two_stage_opamp_dummy_magic_0.V_source.n30 two_stage_opamp_dummy_magic_0.V_source.n28 0.563
R7956 two_stage_opamp_dummy_magic_0.V_source.n32 two_stage_opamp_dummy_magic_0.V_source.n30 0.563
R7957 two_stage_opamp_dummy_magic_0.V_source.n34 two_stage_opamp_dummy_magic_0.V_source.n32 0.563
R7958 two_stage_opamp_dummy_magic_0.V_source.n23 two_stage_opamp_dummy_magic_0.V_source.n21 0.563
R7959 two_stage_opamp_dummy_magic_0.V_source.n25 two_stage_opamp_dummy_magic_0.V_source.n23 0.563
R7960 two_stage_opamp_dummy_magic_0.V_source.n35 two_stage_opamp_dummy_magic_0.V_source.n25 0.53175
R7961 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 144.827
R7962 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 134.577
R7963 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 120.66
R7964 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 97.4009
R7965 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 96.8384
R7966 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 96.8384
R7967 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 96.8384
R7968 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 96.8384
R7969 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 37.4067
R7970 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 35.2505
R7971 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 24.0005
R7972 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 24.0005
R7973 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 24.0005
R7974 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 24.0005
R7975 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 8.0005
R7976 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 8.0005
R7977 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 8.0005
R7978 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 8.0005
R7979 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 8.0005
R7980 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 8.0005
R7981 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 8.0005
R7982 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 8.0005
R7983 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 8.0005
R7984 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 8.0005
R7985 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 5.938
R7986 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 0.563
R7987 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 0.563
R7988 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 0.563
R7989 bgr_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n13 0.047375
R7990 VIN-.n4 VIN-.t8 485.021
R7991 VIN-.n1 VIN-.t6 484.159
R7992 VIN-.n5 VIN-.t7 483.358
R7993 VIN-.n8 VIN-.t10 431.536
R7994 VIN-.n2 VIN-.t9 431.536
R7995 VIN-.n6 VIN-.t1 431.257
R7996 VIN-.n0 VIN-.t0 431.257
R7997 VIN-.n6 VIN-.t2 289.908
R7998 VIN-.n0 VIN-.t5 289.908
R7999 VIN-.n8 VIN-.t4 279.183
R8000 VIN-.n2 VIN-.t3 279.183
R8001 VIN-.n7 VIN-.n6 233.374
R8002 VIN-.n1 VIN-.n0 233.374
R8003 VIN-.n9 VIN-.n8 188.989
R8004 VIN-.n3 VIN-.n2 188.989
R8005 VIN-.n4 VIN-.n3 2.463
R8006 VIN- VIN-.n9 1.78175
R8007 VIN-.n5 VIN-.n4 1.563
R8008 VIN-.n3 VIN-.n1 1.2755
R8009 VIN-.n9 VIN-.n7 1.2755
R8010 VIN-.n7 VIN-.n5 0.8005
R8011 bgr_0.START_UP.n4 bgr_0.START_UP.t6 238.322
R8012 bgr_0.START_UP.n4 bgr_0.START_UP.t7 238.322
R8013 bgr_0.START_UP.n3 bgr_0.START_UP.n1 175.56
R8014 bgr_0.START_UP.n3 bgr_0.START_UP.n2 168.936
R8015 bgr_0.START_UP.n5 bgr_0.START_UP.n4 166.925
R8016 bgr_0.START_UP.n0 bgr_0.START_UP.t1 130.001
R8017 bgr_0.START_UP.n0 bgr_0.START_UP.t0 81.7074
R8018 bgr_0.START_UP bgr_0.START_UP.n0 36.9489
R8019 bgr_0.START_UP bgr_0.START_UP.n5 13.4693
R8020 bgr_0.START_UP.n1 bgr_0.START_UP.t2 13.1338
R8021 bgr_0.START_UP.n1 bgr_0.START_UP.t4 13.1338
R8022 bgr_0.START_UP.n2 bgr_0.START_UP.t3 13.1338
R8023 bgr_0.START_UP.n2 bgr_0.START_UP.t5 13.1338
R8024 bgr_0.START_UP.n5 bgr_0.START_UP.n3 4.21925
R8025 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.t12 670.048
R8026 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.n0 631.982
R8027 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n3 627.128
R8028 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.n1 627.128
R8029 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.n7 226.534
R8030 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.n5 226.534
R8031 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n4 222.034
R8032 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t0 78.8005
R8033 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t2 78.8005
R8034 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t1 78.8005
R8035 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t3 78.8005
R8036 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t11 78.8005
R8037 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t4 78.8005
R8038 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.t6 48.0005
R8039 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.t8 48.0005
R8040 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.t5 48.0005
R8041 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.t10 48.0005
R8042 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.t7 48.0005
R8043 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.t9 48.0005
R8044 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n9 8.938
R8045 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n8 5.7505
R8046 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n2 1.313
R8047 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.n6 1.2505
R8048 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n1 4020
R8049 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.n1 4020
R8050 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n7 4020
R8051 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.n7 4020
R8052 two_stage_opamp_dummy_magic_0.VD3.n4 two_stage_opamp_dummy_magic_0.VD3.t35 660.109
R8053 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.t32 660.109
R8054 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.n11 422.401
R8055 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.n0 422.401
R8056 two_stage_opamp_dummy_magic_0.VD3.t36 two_stage_opamp_dummy_magic_0.VD3.n8 239.915
R8057 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.t33 239.915
R8058 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.n5 230.4
R8059 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.n3 230.4
R8060 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.n3 198.4
R8061 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.n0 198.4
R8062 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.n28 160.428
R8063 two_stage_opamp_dummy_magic_0.VD3.n15 two_stage_opamp_dummy_magic_0.VD3.n13 160.427
R8064 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.n29 159.803
R8065 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.n26 159.803
R8066 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n24 159.803
R8067 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n22 159.802
R8068 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.n20 159.802
R8069 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.n18 159.802
R8070 two_stage_opamp_dummy_magic_0.VD3.n17 two_stage_opamp_dummy_magic_0.VD3.n16 159.802
R8071 two_stage_opamp_dummy_magic_0.VD3.n15 two_stage_opamp_dummy_magic_0.VD3.n14 159.802
R8072 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.n32 155.304
R8073 two_stage_opamp_dummy_magic_0.VD3.n4 two_stage_opamp_dummy_magic_0.VD3.t37 155.125
R8074 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.t34 155.125
R8075 two_stage_opamp_dummy_magic_0.VD3.t0 two_stage_opamp_dummy_magic_0.VD3.t36 98.2764
R8076 two_stage_opamp_dummy_magic_0.VD3.t6 two_stage_opamp_dummy_magic_0.VD3.t0 98.2764
R8077 two_stage_opamp_dummy_magic_0.VD3.t14 two_stage_opamp_dummy_magic_0.VD3.t6 98.2764
R8078 two_stage_opamp_dummy_magic_0.VD3.t10 two_stage_opamp_dummy_magic_0.VD3.t14 98.2764
R8079 two_stage_opamp_dummy_magic_0.VD3.t16 two_stage_opamp_dummy_magic_0.VD3.t10 98.2764
R8080 two_stage_opamp_dummy_magic_0.VD3.t2 two_stage_opamp_dummy_magic_0.VD3.t18 98.2764
R8081 two_stage_opamp_dummy_magic_0.VD3.t8 two_stage_opamp_dummy_magic_0.VD3.t2 98.2764
R8082 two_stage_opamp_dummy_magic_0.VD3.t4 two_stage_opamp_dummy_magic_0.VD3.t8 98.2764
R8083 two_stage_opamp_dummy_magic_0.VD3.t12 two_stage_opamp_dummy_magic_0.VD3.t4 98.2764
R8084 two_stage_opamp_dummy_magic_0.VD3.t33 two_stage_opamp_dummy_magic_0.VD3.t12 98.2764
R8085 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.n10 92.5005
R8086 two_stage_opamp_dummy_magic_0.VD3.n7 two_stage_opamp_dummy_magic_0.VD3.n6 92.5005
R8087 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.n7 92.5005
R8088 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n0 92.5005
R8089 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.n1 92.5005
R8090 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.n1 92.5005
R8091 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.t16 49.1384
R8092 two_stage_opamp_dummy_magic_0.VD3.t18 two_stage_opamp_dummy_magic_0.VD3.n9 49.1384
R8093 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.n4 21.3338
R8094 two_stage_opamp_dummy_magic_0.VD3.n3 two_stage_opamp_dummy_magic_0.VD3.n2 21.3338
R8095 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n23 14.438
R8096 two_stage_opamp_dummy_magic_0.VD3.n29 two_stage_opamp_dummy_magic_0.VD3.t3 11.2576
R8097 two_stage_opamp_dummy_magic_0.VD3.n29 two_stage_opamp_dummy_magic_0.VD3.t9 11.2576
R8098 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.t5 11.2576
R8099 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.t13 11.2576
R8100 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.t15 11.2576
R8101 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.t11 11.2576
R8102 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.t1 11.2576
R8103 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.t7 11.2576
R8104 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.t27 11.2576
R8105 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.t31 11.2576
R8106 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.t25 11.2576
R8107 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.t23 11.2576
R8108 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.t20 11.2576
R8109 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.t21 11.2576
R8110 two_stage_opamp_dummy_magic_0.VD3.n16 two_stage_opamp_dummy_magic_0.VD3.t26 11.2576
R8111 two_stage_opamp_dummy_magic_0.VD3.n16 two_stage_opamp_dummy_magic_0.VD3.t29 11.2576
R8112 two_stage_opamp_dummy_magic_0.VD3.n14 two_stage_opamp_dummy_magic_0.VD3.t24 11.2576
R8113 two_stage_opamp_dummy_magic_0.VD3.n14 two_stage_opamp_dummy_magic_0.VD3.t28 11.2576
R8114 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.t30 11.2576
R8115 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.t22 11.2576
R8116 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.t17 11.2576
R8117 two_stage_opamp_dummy_magic_0.VD3.t19 two_stage_opamp_dummy_magic_0.VD3.n33 11.2576
R8118 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.n12 9.5505
R8119 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.n31 4.5005
R8120 two_stage_opamp_dummy_magic_0.VD3.n31 two_stage_opamp_dummy_magic_0.VD3.n30 0.6255
R8121 two_stage_opamp_dummy_magic_0.VD3.n17 two_stage_opamp_dummy_magic_0.VD3.n15 0.6255
R8122 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.n17 0.6255
R8123 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.n19 0.6255
R8124 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n21 0.6255
R8125 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.n25 0.6255
R8126 two_stage_opamp_dummy_magic_0.VD3.n31 two_stage_opamp_dummy_magic_0.VD3.n27 0.6255
R8127 a_14240_2076.t0 a_14240_2076.t1 169.905
R8128 bgr_0.START_UP_NFET1 bgr_0.START_UP_NFET1.t0 141.653
R8129 a_5190_5068.t0 a_5190_5068.t1 294.339
R8130 a_12530_23988.t0 a_12530_23988.t1 178.133
R8131 VIN+.n9 VIN+.t5 485.127
R8132 VIN+.n4 VIN+.t3 485.127
R8133 VIN+.n3 VIN+.t4 485.127
R8134 VIN+.n7 VIN+.t9 318.656
R8135 VIN+.n7 VIN+.t2 318.656
R8136 VIN+.n5 VIN+.t7 318.656
R8137 VIN+.n5 VIN+.t1 318.656
R8138 VIN+.n1 VIN+.t8 318.656
R8139 VIN+.n1 VIN+.t6 318.656
R8140 VIN+.n0 VIN+.t10 318.656
R8141 VIN+.n0 VIN+.t0 318.656
R8142 VIN+.n2 VIN+.n0 167.05
R8143 VIN+.n8 VIN+.n7 165.8
R8144 VIN+.n6 VIN+.n5 165.8
R8145 VIN+.n2 VIN+.n1 165.8
R8146 VIN+.n6 VIN+.n4 2.34425
R8147 VIN+.n4 VIN+.n3 1.3005
R8148 VIN+.n8 VIN+.n6 1.2505
R8149 VIN+.n3 VIN+.n2 1.15675
R8150 VIN+.n9 VIN+.n8 1.15675
R8151 VIN+ VIN+.n9 0.963
R8152 a_7580_22380.t0 a_7580_22380.t1 178.133
R8153 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 195.608
R8154 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 83.5719
R8155 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 83.5719
R8156 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 83.5719
R8157 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 83.5719
R8158 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 83.5719
R8159 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 83.5719
R8160 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 83.5719
R8161 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 83.5719
R8162 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 83.5719
R8163 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 83.5719
R8164 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 83.5719
R8165 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 83.5719
R8166 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 83.5719
R8167 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 83.5719
R8168 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 83.5719
R8169 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 83.5719
R8170 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 83.5719
R8171 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 83.5719
R8172 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 83.5719
R8173 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 83.5719
R8174 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R8175 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 83.5719
R8176 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 73.8495
R8177 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 73.8495
R8178 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 73.3165
R8179 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 73.3165
R8180 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 73.3165
R8181 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 73.3165
R8182 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 73.3165
R8183 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 73.3165
R8184 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 73.19
R8185 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 73.19
R8186 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 73.19
R8187 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 73.19
R8188 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 73.19
R8189 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 73.19
R8190 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 65.0299
R8191 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 65.0299
R8192 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 26.074
R8193 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 26.074
R8194 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 26.074
R8195 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 26.074
R8196 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 26.074
R8197 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 26.074
R8198 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 26.074
R8199 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 26.074
R8200 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 25.7843
R8201 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 25.7843
R8202 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 25.7843
R8203 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 25.7843
R8204 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 25.7843
R8205 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 25.7843
R8206 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R8207 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R8208 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8209 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R8210 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R8211 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8212 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R8213 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 9.3005
R8214 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R8215 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R8216 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8217 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R8218 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 9.3005
R8219 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 9.3005
R8220 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R8221 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8222 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R8223 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R8224 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R8225 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8226 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R8227 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R8228 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R8229 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R8230 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R8231 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 9.3005
R8232 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 9.3005
R8233 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 9.3005
R8234 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8235 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8236 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8237 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 9.3005
R8238 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8239 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8240 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8241 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 9.3005
R8242 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8243 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8244 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R8245 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8246 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8247 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R8248 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8249 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8250 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8251 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R8252 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8253 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8254 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 9.3005
R8255 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 9.3005
R8256 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R8257 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R8258 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R8259 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R8260 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 4.64654
R8261 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 4.64654
R8262 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 4.64654
R8263 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 4.64654
R8264 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 4.64654
R8265 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 4.64654
R8266 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 4.64654
R8267 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 4.64654
R8268 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 4.64654
R8269 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 2.36206
R8270 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 2.36206
R8271 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 2.36206
R8272 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 2.36206
R8273 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 2.19742
R8274 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 2.19742
R8275 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 2.19742
R8276 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 2.19742
R8277 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 1.56363
R8278 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.56363
R8279 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 1.5505
R8280 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R8281 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 1.5505
R8282 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 1.5505
R8283 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 1.5505
R8284 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 1.5505
R8285 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 1.5505
R8286 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 1.5505
R8287 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 1.5505
R8288 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 1.5505
R8289 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 1.5505
R8290 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 1.5505
R8291 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 1.5505
R8292 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 1.5505
R8293 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 1.5505
R8294 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 1.5505
R8295 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 1.5505
R8296 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 1.5505
R8297 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.25468
R8298 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 1.25468
R8299 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.25468
R8300 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.25468
R8301 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 1.25468
R8302 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 1.25468
R8303 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 1.19225
R8304 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 1.19225
R8305 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 1.19225
R8306 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 1.19225
R8307 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 1.19225
R8308 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.19225
R8309 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 1.07024
R8310 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 1.07024
R8311 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 1.07024
R8312 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 1.07024
R8313 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 1.07024
R8314 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.07024
R8315 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.0237
R8316 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 1.0237
R8317 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.0237
R8318 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.0237
R8319 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 1.0237
R8320 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 1.0237
R8321 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.885803
R8322 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 0.885803
R8323 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 0.885803
R8324 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 0.885803
R8325 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.885803
R8326 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.885803
R8327 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 0.885803
R8328 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.885803
R8329 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 0.812055
R8330 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 0.812055
R8331 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.77514
R8332 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.77514
R8333 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 0.77514
R8334 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.77514
R8335 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.77514
R8336 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 0.77514
R8337 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 0.77514
R8338 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 0.77514
R8339 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.756696
R8340 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R8341 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.756696
R8342 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 0.756696
R8343 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R8344 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.756696
R8345 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R8346 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.756696
R8347 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 0.711459
R8348 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.711459
R8349 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.647417
R8350 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 0.647417
R8351 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.590702
R8352 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 0.590702
R8353 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.590702
R8354 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 0.590702
R8355 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.590702
R8356 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 0.590702
R8357 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.576566
R8358 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.576566
R8359 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 0.530034
R8360 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 0.530034
R8361 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 0.290206
R8362 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 0.290206
R8363 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 0.290206
R8364 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 0.290206
R8365 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 0.290206
R8366 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 0.290206
R8367 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 0.290206
R8368 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 0.290206
R8369 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8370 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8371 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8372 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.203382
R8373 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8374 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 0.203382
R8375 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 0.154071
R8376 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 0.154071
R8377 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 0.154071
R8378 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 0.154071
R8379 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 0.137464
R8380 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 0.137464
R8381 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 0.134964
R8382 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 0.134964
R8383 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R8384 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 0.0183571
R8385 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R8386 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R8387 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 0.0183571
R8388 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R8389 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R8390 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 0.0183571
R8391 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0183571
R8392 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R8393 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R8394 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R8395 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R8396 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 0.0183571
R8397 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R8398 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R8399 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 0.0183571
R8400 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0183571
R8401 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0106786
R8402 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0106786
R8403 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.0106786
R8404 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 0.00992001
R8405 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 0.00992001
R8406 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R8407 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 0.00992001
R8408 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R8409 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R8410 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R8411 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 0.00992001
R8412 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 0.00992001
R8413 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 0.00992001
R8414 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R8415 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 0.00992001
R8416 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R8417 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R8418 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R8419 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R8420 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 0.00992001
R8421 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R8422 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.00817857
R8423 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00817857
R8424 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 0.00817857
R8425 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 0.00817857
R8426 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.00817857
R8427 a_12410_22380.t0 a_12410_22380.t1 178.133
R8428 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 2655
R8429 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 2595
R8430 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 2280
R8431 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 2250
R8432 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 672.159
R8433 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 672.159
R8434 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 276.8
R8435 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 240
R8436 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 206.4
R8437 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 204.8
R8438 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 179.933
R8439 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 170.3
R8440 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 160.517
R8441 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 160.517
R8442 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 110.425
R8443 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 110.05
R8444 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 95.7988
R8445 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 92.5005
R8446 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 92.5005
R8447 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 92.5005
R8448 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 92.5005
R8449 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 89.6005
R8450 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 89.6005
R8451 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 76.8005
R8452 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 75.9449
R8453 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 75.9449
R8454 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 47.8997
R8455 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 47.8997
R8456 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 38.4005
R8457 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 24.5338
R8458 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 24.5338
R8459 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 16.8187
R8460 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 16.8187
R8461 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 11.0991
R8462 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 11.0991
R8463 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 10.9449
R8464 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 10.9449
R8465 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 6.21925
R8466 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 4.5005
R8467 a_13060_22630.t0 a_13060_22630.t1 178.133
R8468 a_6930_22590.t0 a_6930_22590.t1 178.133
R8469 a_13180_23838.t0 a_13180_23838.t1 178.133
R8470 a_5710_2076.t0 a_5710_2076.t1 169.905
R8471 a_5310_5068.t0 a_5310_5068.t1 169.905
R8472 a_14680_5068.t0 a_14680_5068.t1 169.905
C0 VOUT- two_stage_opamp_dummy_magic_0.cap_res_Y 50.8385f
C1 VIN- two_stage_opamp_dummy_magic_0.VD1 0.85667f
C2 VOUT- VOUT+ 0.305434f
C3 VDDA bgr_0.V_TOP 15.1696f
C4 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_amp_ref 1.40619f
C5 VIN+ two_stage_opamp_dummy_magic_0.VD1 0.058217f
C6 VDDA two_stage_opamp_dummy_magic_0.err_amp_out 1.13079f
C7 bgr_0.START_UP two_stage_opamp_dummy_magic_0.V_err_amp_ref 1.36422f
C8 VDDA two_stage_opamp_dummy_magic_0.cap_res_Y 0.798008f
C9 two_stage_opamp_dummy_magic_0.VD4 two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.508546f
C10 m2_10730_16580# bgr_0.1st_Vout_1 0.075543f
C11 VDDA VOUT+ 6.65903f
C12 VDDA two_stage_opamp_dummy_magic_0.X 5.39586f
C13 VDDA bgr_0.START_UP_NFET1 0.148407f
C14 bgr_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_amp_ref 1.64432f
C15 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.X 0.425972f
C16 VOUT- two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.038796f
C17 VOUT+ two_stage_opamp_dummy_magic_0.cap_res_Y 0.028842f
C18 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_gate 3.51065f
C19 VOUT+ two_stage_opamp_dummy_magic_0.X 2.14019f
C20 bgr_0.NFET_GATE_10uA bgr_0.START_UP 1.60479f
C21 bgr_0.1st_Vout_1 bgr_0.NFET_GATE_10uA 0.038707f
C22 VDDA two_stage_opamp_dummy_magic_0.V_err_amp_ref 4.2739f
C23 bgr_0.1st_Vout_1 two_stage_opamp_dummy_magic_0.V_err_gate 0.041082f
C24 bgr_0.V_TOP two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.581165f
C25 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.VD4 0.013177f
C26 m2_10730_16580# VDDA 0.010446f
C27 bgr_0.NFET_GATE_10uA bgr_0.PFET_GATE_10uA 0.011883f
C28 m2_10730_16580# bgr_0.V_TOP 0.012f
C29 bgr_0.1st_Vout_1 bgr_0.START_UP 0.041693f
C30 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.Vb2_Vb3 0.069137f
C31 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.52226f
C32 two_stage_opamp_dummy_magic_0.cap_res_Y two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.238802f
C33 VIN- VIN+ 0.562828f
C34 VDDA bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.046803f
C35 bgr_0.V_TOP bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.055802f
C36 VDDA bgr_0.NFET_GATE_10uA 1.06707f
C37 bgr_0.V_TOP bgr_0.NFET_GATE_10uA 0.062551f
C38 VDDA two_stage_opamp_dummy_magic_0.V_err_gate 4.16561f
C39 m2_9370_16580# bgr_0.PFET_GATE_10uA 0.012f
C40 bgr_0.V_TOP two_stage_opamp_dummy_magic_0.V_err_gate 0.081361f
C41 VDDA bgr_0.START_UP 1.52151f
C42 bgr_0.V_TOP bgr_0.START_UP 0.812081f
C43 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.V_err_gate 0.261364f
C44 VDDA bgr_0.1st_Vout_1 2.13761f
C45 bgr_0.1st_Vout_1 bgr_0.V_TOP 2.47115f
C46 VDDA two_stage_opamp_dummy_magic_0.VD4 4.42804f
C47 VDDA two_stage_opamp_dummy_magic_0.Vb2_Vb3 0.987228f
C48 VDDA bgr_0.PFET_GATE_10uA 9.750259f
C49 bgr_0.V_TOP bgr_0.PFET_GATE_10uA 0.18077f
C50 bgr_0.NFET_GATE_10uA bgr_0.START_UP_NFET1 0.318695f
C51 VOUT+ two_stage_opamp_dummy_magic_0.V_err_gate 0.039202f
C52 two_stage_opamp_dummy_magic_0.X two_stage_opamp_dummy_magic_0.V_err_gate 0.128771f
C53 VDDA VOUT- 6.69956f
C54 bgr_0.START_UP_NFET1 bgr_0.START_UP 0.145663f
C55 m2_9370_16580# VDDA 0.010446f
C56 two_stage_opamp_dummy_magic_0.cap_res_Y two_stage_opamp_dummy_magic_0.VD4 0.036097f
C57 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.X 1.05328f
C58 two_stage_opamp_dummy_magic_0.cap_res_Y bgr_0.PFET_GATE_10uA 0.01025f
C59 VOUT+ two_stage_opamp_dummy_magic_0.Vb2_Vb3 0.039712f
C60 VIN+ GNDA 2.062214f
C61 VIN- GNDA 2.154258f
C62 VOUT+ GNDA 17.61802f
C63 VOUT- GNDA 17.631264f
C64 VDDA GNDA 0.158145p
C65 two_stage_opamp_dummy_magic_0.VD1 GNDA 2.42208f
C66 two_stage_opamp_dummy_magic_0.err_amp_out GNDA 2.678583f
C67 two_stage_opamp_dummy_magic_0.cap_res_Y GNDA 33.765926f
C68 two_stage_opamp_dummy_magic_0.X GNDA 5.494094f
C69 bgr_0.1st_Vout_1 GNDA 7.153163f
C70 bgr_0.START_UP GNDA 6.451247f
C71 bgr_0.START_UP_NFET1 GNDA 5.22875f
C72 two_stage_opamp_dummy_magic_0.V_err_gate GNDA 9.435944f
C73 bgr_0.NFET_GATE_10uA GNDA 8.19126f
C74 bgr_0.V_TOP GNDA 8.727081f
C75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA 18.0473f
C76 two_stage_opamp_dummy_magic_0.V_err_amp_ref GNDA 6.953361f
C77 bgr_0.PFET_GATE_10uA GNDA 5.555353f
C78 two_stage_opamp_dummy_magic_0.VD4 GNDA 6.43896f
C79 two_stage_opamp_dummy_magic_0.Vb2_Vb3 GNDA 3.47841f
C80 VIN+.t0 GNDA 0.042021f
C81 VIN+.t10 GNDA 0.042021f
C82 VIN+.n0 GNDA 0.086842f
C83 VIN+.t6 GNDA 0.042021f
C84 VIN+.t8 GNDA 0.042021f
C85 VIN+.n1 GNDA 0.085639f
C86 VIN+.n2 GNDA 0.361638f
C87 VIN+.t4 GNDA 0.059118f
C88 VIN+.n3 GNDA 0.216459f
C89 VIN+.t3 GNDA 0.059118f
C90 VIN+.n4 GNDA 0.263959f
C91 VIN+.t1 GNDA 0.042021f
C92 VIN+.t7 GNDA 0.042021f
C93 VIN+.n5 GNDA 0.085639f
C94 VIN+.n6 GNDA 0.249653f
C95 VIN+.t2 GNDA 0.042021f
C96 VIN+.t9 GNDA 0.042021f
C97 VIN+.n7 GNDA 0.085639f
C98 VIN+.n8 GNDA 0.202005f
C99 VIN+.t5 GNDA 0.059118f
C100 VIN+.n9 GNDA 0.202625f
C101 two_stage_opamp_dummy_magic_0.VD3.t17 GNDA 0.026025f
C102 two_stage_opamp_dummy_magic_0.VD3.n0 GNDA 0.073371f
C103 two_stage_opamp_dummy_magic_0.VD3.n1 GNDA 0.100747f
C104 two_stage_opamp_dummy_magic_0.VD3.t34 GNDA 0.128386f
C105 two_stage_opamp_dummy_magic_0.VD3.t32 GNDA 0.045318f
C106 two_stage_opamp_dummy_magic_0.VD3.n2 GNDA 0.083755f
C107 two_stage_opamp_dummy_magic_0.VD3.n3 GNDA 0.053992f
C108 two_stage_opamp_dummy_magic_0.VD3.t37 GNDA 0.128386f
C109 two_stage_opamp_dummy_magic_0.VD3.t35 GNDA 0.045318f
C110 two_stage_opamp_dummy_magic_0.VD3.n4 GNDA 0.083755f
C111 two_stage_opamp_dummy_magic_0.VD3.n5 GNDA 0.053992f
C112 two_stage_opamp_dummy_magic_0.VD3.n6 GNDA 0.053537f
C113 two_stage_opamp_dummy_magic_0.VD3.n7 GNDA 0.100747f
C114 two_stage_opamp_dummy_magic_0.VD3.n8 GNDA 0.300245f
C115 two_stage_opamp_dummy_magic_0.VD3.t36 GNDA 0.448159f
C116 two_stage_opamp_dummy_magic_0.VD3.t0 GNDA 0.25876f
C117 two_stage_opamp_dummy_magic_0.VD3.t6 GNDA 0.25876f
C118 two_stage_opamp_dummy_magic_0.VD3.t14 GNDA 0.25876f
C119 two_stage_opamp_dummy_magic_0.VD3.t10 GNDA 0.25876f
C120 two_stage_opamp_dummy_magic_0.VD3.t16 GNDA 0.19407f
C121 two_stage_opamp_dummy_magic_0.VD3.n9 GNDA 0.12938f
C122 two_stage_opamp_dummy_magic_0.VD3.t18 GNDA 0.19407f
C123 two_stage_opamp_dummy_magic_0.VD3.t2 GNDA 0.25876f
C124 two_stage_opamp_dummy_magic_0.VD3.t8 GNDA 0.25876f
C125 two_stage_opamp_dummy_magic_0.VD3.t4 GNDA 0.25876f
C126 two_stage_opamp_dummy_magic_0.VD3.t12 GNDA 0.25876f
C127 two_stage_opamp_dummy_magic_0.VD3.t33 GNDA 0.448159f
C128 two_stage_opamp_dummy_magic_0.VD3.n10 GNDA 0.300245f
C129 two_stage_opamp_dummy_magic_0.VD3.n11 GNDA 0.073371f
C130 two_stage_opamp_dummy_magic_0.VD3.n12 GNDA 0.108171f
C131 two_stage_opamp_dummy_magic_0.VD3.t30 GNDA 0.026025f
C132 two_stage_opamp_dummy_magic_0.VD3.t22 GNDA 0.026025f
C133 two_stage_opamp_dummy_magic_0.VD3.n13 GNDA 0.090509f
C134 two_stage_opamp_dummy_magic_0.VD3.t24 GNDA 0.026025f
C135 two_stage_opamp_dummy_magic_0.VD3.t28 GNDA 0.026025f
C136 two_stage_opamp_dummy_magic_0.VD3.n14 GNDA 0.090188f
C137 two_stage_opamp_dummy_magic_0.VD3.n15 GNDA 0.170266f
C138 two_stage_opamp_dummy_magic_0.VD3.t26 GNDA 0.026025f
C139 two_stage_opamp_dummy_magic_0.VD3.t29 GNDA 0.026025f
C140 two_stage_opamp_dummy_magic_0.VD3.n16 GNDA 0.090188f
C141 two_stage_opamp_dummy_magic_0.VD3.n17 GNDA 0.088268f
C142 two_stage_opamp_dummy_magic_0.VD3.t20 GNDA 0.026025f
C143 two_stage_opamp_dummy_magic_0.VD3.t21 GNDA 0.026025f
C144 two_stage_opamp_dummy_magic_0.VD3.n18 GNDA 0.090188f
C145 two_stage_opamp_dummy_magic_0.VD3.n19 GNDA 0.088268f
C146 two_stage_opamp_dummy_magic_0.VD3.t25 GNDA 0.026025f
C147 two_stage_opamp_dummy_magic_0.VD3.t23 GNDA 0.026025f
C148 two_stage_opamp_dummy_magic_0.VD3.n20 GNDA 0.090188f
C149 two_stage_opamp_dummy_magic_0.VD3.n21 GNDA 0.088268f
C150 two_stage_opamp_dummy_magic_0.VD3.t27 GNDA 0.026025f
C151 two_stage_opamp_dummy_magic_0.VD3.t31 GNDA 0.026025f
C152 two_stage_opamp_dummy_magic_0.VD3.n22 GNDA 0.090188f
C153 two_stage_opamp_dummy_magic_0.VD3.n23 GNDA 0.169329f
C154 two_stage_opamp_dummy_magic_0.VD3.t1 GNDA 0.026025f
C155 two_stage_opamp_dummy_magic_0.VD3.t7 GNDA 0.026025f
C156 two_stage_opamp_dummy_magic_0.VD3.n24 GNDA 0.090188f
C157 two_stage_opamp_dummy_magic_0.VD3.n25 GNDA 0.163355f
C158 two_stage_opamp_dummy_magic_0.VD3.t15 GNDA 0.026025f
C159 two_stage_opamp_dummy_magic_0.VD3.t11 GNDA 0.026025f
C160 two_stage_opamp_dummy_magic_0.VD3.n26 GNDA 0.090188f
C161 two_stage_opamp_dummy_magic_0.VD3.n27 GNDA 0.088268f
C162 two_stage_opamp_dummy_magic_0.VD3.t5 GNDA 0.026025f
C163 two_stage_opamp_dummy_magic_0.VD3.t13 GNDA 0.026025f
C164 two_stage_opamp_dummy_magic_0.VD3.n28 GNDA 0.090509f
C165 two_stage_opamp_dummy_magic_0.VD3.t3 GNDA 0.026025f
C166 two_stage_opamp_dummy_magic_0.VD3.t9 GNDA 0.026025f
C167 two_stage_opamp_dummy_magic_0.VD3.n29 GNDA 0.090188f
C168 two_stage_opamp_dummy_magic_0.VD3.n30 GNDA 0.170266f
C169 two_stage_opamp_dummy_magic_0.VD3.n31 GNDA 0.023794f
C170 two_stage_opamp_dummy_magic_0.VD3.n32 GNDA 0.069277f
C171 two_stage_opamp_dummy_magic_0.VD3.n33 GNDA 0.08832f
C172 two_stage_opamp_dummy_magic_0.VD3.t19 GNDA 0.026025f
C173 two_stage_opamp_dummy_magic_0.err_amp_out.n0 GNDA 0.018848f
C174 two_stage_opamp_dummy_magic_0.err_amp_out.n1 GNDA 0.018642f
C175 two_stage_opamp_dummy_magic_0.err_amp_out.n2 GNDA 0.371454f
C176 two_stage_opamp_dummy_magic_0.err_amp_out.n3 GNDA 0.018642f
C177 two_stage_opamp_dummy_magic_0.err_amp_out.n4 GNDA 0.020813f
C178 two_stage_opamp_dummy_magic_0.err_amp_out.t12 GNDA 0.074665f
C179 two_stage_opamp_dummy_magic_0.err_amp_out.n5 GNDA 0.022234f
C180 two_stage_opamp_dummy_magic_0.err_amp_out.n6 GNDA 1.11353f
C181 two_stage_opamp_dummy_magic_0.err_amp_out.n7 GNDA 0.022234f
C182 two_stage_opamp_dummy_magic_0.err_amp_out.n8 GNDA 0.195309f
C183 two_stage_opamp_dummy_magic_0.err_amp_out.n9 GNDA 0.190271f
C184 bgr_0.START_UP.t0 GNDA 1.06745f
C185 bgr_0.START_UP.t1 GNDA 0.02806f
C186 bgr_0.START_UP.n0 GNDA 0.714928f
C187 bgr_0.START_UP.t2 GNDA 0.026778f
C188 bgr_0.START_UP.t4 GNDA 0.026778f
C189 bgr_0.START_UP.n1 GNDA 0.097147f
C190 bgr_0.START_UP.t3 GNDA 0.026778f
C191 bgr_0.START_UP.t5 GNDA 0.026778f
C192 bgr_0.START_UP.n2 GNDA 0.08937f
C193 bgr_0.START_UP.n3 GNDA 0.462855f
C194 bgr_0.START_UP.t7 GNDA 0.010062f
C195 bgr_0.START_UP.t6 GNDA 0.010062f
C196 bgr_0.START_UP.n4 GNDA 0.028407f
C197 bgr_0.START_UP.n5 GNDA 0.260836f
C198 VIN-.t6 GNDA 0.050911f
C199 VIN-.t5 GNDA 0.03359f
C200 VIN-.t0 GNDA 0.04147f
C201 VIN-.n0 GNDA 0.05959f
C202 VIN-.n1 GNDA 0.281971f
C203 VIN-.t3 GNDA 0.033038f
C204 VIN-.t9 GNDA 0.041485f
C205 VIN-.n2 GNDA 0.065237f
C206 VIN-.n3 GNDA 0.201948f
C207 VIN-.t8 GNDA 0.050345f
C208 VIN-.n4 GNDA 0.237498f
C209 VIN-.t7 GNDA 0.050694f
C210 VIN-.n5 GNDA 0.181582f
C211 VIN-.t2 GNDA 0.03359f
C212 VIN-.t1 GNDA 0.04147f
C213 VIN-.n6 GNDA 0.05959f
C214 VIN-.n7 GNDA 0.150425f
C215 VIN-.t4 GNDA 0.033038f
C216 VIN-.t10 GNDA 0.041485f
C217 VIN-.n8 GNDA 0.065237f
C218 VIN-.n9 GNDA 0.178598f
C219 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 GNDA 0.020333f
C220 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 GNDA 0.020333f
C221 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 GNDA 0.073906f
C222 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 GNDA 0.020333f
C223 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 GNDA 0.020333f
C224 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 GNDA 0.061415f
C225 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 GNDA 1.19789f
C226 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 GNDA 0.253162f
C227 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 GNDA 0.061f
C228 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 GNDA 0.061f
C229 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 GNDA 0.252259f
C230 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 GNDA 0.061f
C231 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 GNDA 0.061f
C232 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 GNDA 0.251291f
C233 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 GNDA 0.348416f
C234 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 GNDA 0.061f
C235 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 GNDA 0.061f
C236 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 GNDA 0.251291f
C237 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 GNDA 0.181808f
C238 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 GNDA 0.061f
C239 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 GNDA 0.061f
C240 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 GNDA 0.251291f
C241 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 GNDA 0.181808f
C242 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 GNDA 0.061f
C243 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 GNDA 0.061f
C244 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 GNDA 0.251291f
C245 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 GNDA 0.267294f
C246 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 GNDA 1.54748f
C247 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n13 GNDA 1.8279f
C248 bgr_0.V_CMFB_S4 GNDA 0.010167f
C249 two_stage_opamp_dummy_magic_0.V_source.t9 GNDA 0.024498f
C250 two_stage_opamp_dummy_magic_0.V_source.t31 GNDA 0.024498f
C251 two_stage_opamp_dummy_magic_0.V_source.t38 GNDA 0.024498f
C252 two_stage_opamp_dummy_magic_0.V_source.n0 GNDA 0.097805f
C253 two_stage_opamp_dummy_magic_0.V_source.t19 GNDA 0.024498f
C254 two_stage_opamp_dummy_magic_0.V_source.t13 GNDA 0.024498f
C255 two_stage_opamp_dummy_magic_0.V_source.n1 GNDA 0.097268f
C256 two_stage_opamp_dummy_magic_0.V_source.n2 GNDA 0.169458f
C257 two_stage_opamp_dummy_magic_0.V_source.t6 GNDA 0.024498f
C258 two_stage_opamp_dummy_magic_0.V_source.t12 GNDA 0.024498f
C259 two_stage_opamp_dummy_magic_0.V_source.n3 GNDA 0.09772f
C260 two_stage_opamp_dummy_magic_0.V_source.t8 GNDA 0.024498f
C261 two_stage_opamp_dummy_magic_0.V_source.t16 GNDA 0.024498f
C262 two_stage_opamp_dummy_magic_0.V_source.n4 GNDA 0.097268f
C263 two_stage_opamp_dummy_magic_0.V_source.n5 GNDA 0.166602f
C264 two_stage_opamp_dummy_magic_0.V_source.t10 GNDA 0.024498f
C265 two_stage_opamp_dummy_magic_0.V_source.t18 GNDA 0.024498f
C266 two_stage_opamp_dummy_magic_0.V_source.n6 GNDA 0.097268f
C267 two_stage_opamp_dummy_magic_0.V_source.n7 GNDA 0.086957f
C268 two_stage_opamp_dummy_magic_0.V_source.t23 GNDA 0.102648f
C269 two_stage_opamp_dummy_magic_0.V_source.t14 GNDA 0.024498f
C270 two_stage_opamp_dummy_magic_0.V_source.t4 GNDA 0.024498f
C271 two_stage_opamp_dummy_magic_0.V_source.n8 GNDA 0.09453f
C272 two_stage_opamp_dummy_magic_0.V_source.n9 GNDA 0.675932f
C273 two_stage_opamp_dummy_magic_0.V_source.n10 GNDA 0.029398f
C274 two_stage_opamp_dummy_magic_0.V_source.t11 GNDA 0.024498f
C275 two_stage_opamp_dummy_magic_0.V_source.t3 GNDA 0.024498f
C276 two_stage_opamp_dummy_magic_0.V_source.n11 GNDA 0.097268f
C277 two_stage_opamp_dummy_magic_0.V_source.n12 GNDA 0.086957f
C278 two_stage_opamp_dummy_magic_0.V_source.t15 GNDA 0.024498f
C279 two_stage_opamp_dummy_magic_0.V_source.t5 GNDA 0.024498f
C280 two_stage_opamp_dummy_magic_0.V_source.n13 GNDA 0.097268f
C281 two_stage_opamp_dummy_magic_0.V_source.n14 GNDA 0.086957f
C282 two_stage_opamp_dummy_magic_0.V_source.t17 GNDA 0.024498f
C283 two_stage_opamp_dummy_magic_0.V_source.t7 GNDA 0.024498f
C284 two_stage_opamp_dummy_magic_0.V_source.n15 GNDA 0.097268f
C285 two_stage_opamp_dummy_magic_0.V_source.n16 GNDA 0.086957f
C286 two_stage_opamp_dummy_magic_0.V_source.n17 GNDA 0.029398f
C287 two_stage_opamp_dummy_magic_0.V_source.t34 GNDA 0.014699f
C288 two_stage_opamp_dummy_magic_0.V_source.t28 GNDA 0.014699f
C289 two_stage_opamp_dummy_magic_0.V_source.n18 GNDA 0.049939f
C290 two_stage_opamp_dummy_magic_0.V_source.t21 GNDA 0.014699f
C291 two_stage_opamp_dummy_magic_0.V_source.t25 GNDA 0.014699f
C292 two_stage_opamp_dummy_magic_0.V_source.n19 GNDA 0.052807f
C293 two_stage_opamp_dummy_magic_0.V_source.t22 GNDA 0.014699f
C294 two_stage_opamp_dummy_magic_0.V_source.t30 GNDA 0.014699f
C295 two_stage_opamp_dummy_magic_0.V_source.n20 GNDA 0.0524f
C296 two_stage_opamp_dummy_magic_0.V_source.n21 GNDA 0.177206f
C297 two_stage_opamp_dummy_magic_0.V_source.t36 GNDA 0.014699f
C298 two_stage_opamp_dummy_magic_0.V_source.t1 GNDA 0.014699f
C299 two_stage_opamp_dummy_magic_0.V_source.n22 GNDA 0.0524f
C300 two_stage_opamp_dummy_magic_0.V_source.n23 GNDA 0.092237f
C301 two_stage_opamp_dummy_magic_0.V_source.t32 GNDA 0.014699f
C302 two_stage_opamp_dummy_magic_0.V_source.t27 GNDA 0.014699f
C303 two_stage_opamp_dummy_magic_0.V_source.n24 GNDA 0.0524f
C304 two_stage_opamp_dummy_magic_0.V_source.n25 GNDA 0.091747f
C305 two_stage_opamp_dummy_magic_0.V_source.t33 GNDA 0.014699f
C306 two_stage_opamp_dummy_magic_0.V_source.t39 GNDA 0.014699f
C307 two_stage_opamp_dummy_magic_0.V_source.n26 GNDA 0.052785f
C308 two_stage_opamp_dummy_magic_0.V_source.t29 GNDA 0.014699f
C309 two_stage_opamp_dummy_magic_0.V_source.t40 GNDA 0.014699f
C310 two_stage_opamp_dummy_magic_0.V_source.n27 GNDA 0.0524f
C311 two_stage_opamp_dummy_magic_0.V_source.n28 GNDA 0.175465f
C312 two_stage_opamp_dummy_magic_0.V_source.t26 GNDA 0.014699f
C313 two_stage_opamp_dummy_magic_0.V_source.t2 GNDA 0.014699f
C314 two_stage_opamp_dummy_magic_0.V_source.n29 GNDA 0.0524f
C315 two_stage_opamp_dummy_magic_0.V_source.n30 GNDA 0.092237f
C316 two_stage_opamp_dummy_magic_0.V_source.t0 GNDA 0.014699f
C317 two_stage_opamp_dummy_magic_0.V_source.t24 GNDA 0.014699f
C318 two_stage_opamp_dummy_magic_0.V_source.n31 GNDA 0.0524f
C319 two_stage_opamp_dummy_magic_0.V_source.n32 GNDA 0.092237f
C320 two_stage_opamp_dummy_magic_0.V_source.t35 GNDA 0.014699f
C321 two_stage_opamp_dummy_magic_0.V_source.t37 GNDA 0.014699f
C322 two_stage_opamp_dummy_magic_0.V_source.n33 GNDA 0.0524f
C323 two_stage_opamp_dummy_magic_0.V_source.n34 GNDA 0.140743f
C324 two_stage_opamp_dummy_magic_0.V_source.n35 GNDA 0.077414f
C325 two_stage_opamp_dummy_magic_0.V_source.n36 GNDA 0.082836f
C326 two_stage_opamp_dummy_magic_0.V_source.n37 GNDA 0.082155f
C327 two_stage_opamp_dummy_magic_0.V_source.n38 GNDA 0.09453f
C328 two_stage_opamp_dummy_magic_0.V_source.t20 GNDA 0.024498f
C329 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 GNDA 0.016041f
C330 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 GNDA 0.016041f
C331 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 GNDA 0.040208f
C332 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 GNDA 0.016041f
C333 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 GNDA 0.016041f
C334 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 GNDA 0.039996f
C335 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 GNDA 0.355484f
C336 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 GNDA 0.016041f
C337 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 GNDA 0.016041f
C338 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 GNDA 0.032081f
C339 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 GNDA 0.059661f
C340 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 GNDA 0.205433f
C341 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 GNDA 0.032081f
C342 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 GNDA 0.032081f
C343 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 GNDA 0.094125f
C344 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 GNDA 0.032081f
C345 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 GNDA 0.032081f
C346 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 GNDA 0.093697f
C347 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 GNDA 0.323873f
C348 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 GNDA 0.032081f
C349 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 GNDA 0.032081f
C350 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 GNDA 0.093697f
C351 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 GNDA 0.167764f
C352 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 GNDA 0.032081f
C353 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 GNDA 0.032081f
C354 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 GNDA 0.093697f
C355 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 GNDA 0.167764f
C356 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 GNDA 0.032081f
C357 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 GNDA 0.032081f
C358 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 GNDA 0.093697f
C359 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 GNDA 0.245609f
C360 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 GNDA 1.4546f
C361 bgr_0.V_CMFB_S1 GNDA 0.921551f
C362 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA 0.240411f
C363 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA 0.240438f
C364 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA 0.225686f
C365 two_stage_opamp_dummy_magic_0.V_tot.n0 GNDA 1.16969f
C366 two_stage_opamp_dummy_magic_0.V_tot.t11 GNDA 0.011798f
C367 two_stage_opamp_dummy_magic_0.V_tot.t5 GNDA 0.011798f
C368 two_stage_opamp_dummy_magic_0.V_tot.n1 GNDA 0.053113f
C369 two_stage_opamp_dummy_magic_0.V_tot.t12 GNDA 0.011798f
C370 two_stage_opamp_dummy_magic_0.V_tot.t8 GNDA 0.011798f
C371 two_stage_opamp_dummy_magic_0.V_tot.n2 GNDA 0.052149f
C372 two_stage_opamp_dummy_magic_0.V_tot.n3 GNDA 0.289549f
C373 two_stage_opamp_dummy_magic_0.V_tot.t4 GNDA 0.027075f
C374 two_stage_opamp_dummy_magic_0.V_tot.n4 GNDA 0.152118f
C375 two_stage_opamp_dummy_magic_0.V_tot.t6 GNDA 0.027256f
C376 two_stage_opamp_dummy_magic_0.V_tot.t9 GNDA 0.012231f
C377 two_stage_opamp_dummy_magic_0.V_tot.t10 GNDA 0.012231f
C378 two_stage_opamp_dummy_magic_0.V_tot.n5 GNDA 0.044381f
C379 two_stage_opamp_dummy_magic_0.V_tot.n6 GNDA 0.259533f
C380 two_stage_opamp_dummy_magic_0.V_tot.t7 GNDA 0.011798f
C381 two_stage_opamp_dummy_magic_0.V_tot.t13 GNDA 0.011798f
C382 two_stage_opamp_dummy_magic_0.V_tot.n7 GNDA 0.052149f
C383 two_stage_opamp_dummy_magic_0.V_tot.n8 GNDA 0.191378f
C384 two_stage_opamp_dummy_magic_0.V_tot.n9 GNDA 0.206537f
C385 two_stage_opamp_dummy_magic_0.V_tot.n10 GNDA 1.88795f
C386 two_stage_opamp_dummy_magic_0.V_tot.n11 GNDA 1.15965f
C387 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA 0.225686f
C388 two_stage_opamp_dummy_magic_0.V_err_p.n0 GNDA 0.021118f
C389 two_stage_opamp_dummy_magic_0.V_err_p.n1 GNDA 0.020212f
C390 two_stage_opamp_dummy_magic_0.V_err_p.n2 GNDA 0.020262f
C391 two_stage_opamp_dummy_magic_0.V_err_p.n3 GNDA 0.021093f
C392 two_stage_opamp_dummy_magic_0.V_err_p.n4 GNDA 0.020966f
C393 two_stage_opamp_dummy_magic_0.V_err_p.n5 GNDA 0.297859f
C394 two_stage_opamp_dummy_magic_0.V_err_p.n6 GNDA 0.020966f
C395 two_stage_opamp_dummy_magic_0.V_err_p.n7 GNDA 0.155369f
C396 two_stage_opamp_dummy_magic_0.V_err_p.n8 GNDA 0.020966f
C397 two_stage_opamp_dummy_magic_0.V_err_p.n9 GNDA 0.189616f
C398 two_stage_opamp_dummy_magic_0.V_err_p.n10 GNDA 0.160506f
C399 two_stage_opamp_dummy_magic_0.V_err_p.n11 GNDA 0.14076f
C400 two_stage_opamp_dummy_magic_0.V_err_p.n12 GNDA 0.241198f
C401 two_stage_opamp_dummy_magic_0.V_err_p.n13 GNDA 0.021118f
C402 two_stage_opamp_dummy_magic_0.V_err_p.n14 GNDA 0.020826f
C403 two_stage_opamp_dummy_magic_0.V_err_p.n15 GNDA 0.326026f
C404 two_stage_opamp_dummy_magic_0.V_err_p.n16 GNDA 0.020826f
C405 two_stage_opamp_dummy_magic_0.V_err_p.n17 GNDA 0.179554f
C406 two_stage_opamp_dummy_magic_0.V_err_p.n18 GNDA 0.179554f
C407 two_stage_opamp_dummy_magic_0.V_err_p.n19 GNDA 0.020826f
C408 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 GNDA 0.019818f
C409 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 GNDA 0.019818f
C410 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 GNDA 0.072035f
C411 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 GNDA 0.019818f
C412 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 GNDA 0.019818f
C413 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 GNDA 0.05986f
C414 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 GNDA 1.16756f
C415 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 GNDA 0.246752f
C416 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 GNDA 0.059456f
C417 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 GNDA 0.059456f
C418 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 GNDA 0.245873f
C419 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 GNDA 0.059456f
C420 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 GNDA 0.059456f
C421 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 GNDA 0.244929f
C422 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 GNDA 0.339595f
C423 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 GNDA 0.059456f
C424 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 GNDA 0.059456f
C425 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 GNDA 0.244929f
C426 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 GNDA 0.177206f
C427 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA 0.059456f
C428 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 GNDA 0.059456f
C429 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 GNDA 0.244929f
C430 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 GNDA 0.177206f
C431 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA 0.059456f
C432 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 GNDA 0.059456f
C433 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 GNDA 0.244929f
C434 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 GNDA 0.260527f
C435 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 GNDA 1.5083f
C436 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n13 GNDA 1.78163f
C437 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 GNDA 0.21829f
C438 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 GNDA 0.593397f
C439 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 GNDA 0.544212f
C440 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 GNDA 0.544212f
C441 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 GNDA 0.645895f
C442 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 GNDA 0.341156f
C443 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 GNDA 0.215911f
C444 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 GNDA 0.199536f
C445 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 GNDA 1.1506f
C446 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 GNDA 0.544212f
C447 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 GNDA 0.544212f
C448 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 GNDA 0.645895f
C449 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 GNDA 0.341156f
C450 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 GNDA 0.215911f
C451 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 GNDA 0.593397f
C452 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 GNDA 0.199536f
C453 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 GNDA 1.14462f
C454 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 GNDA 0.217852f
C455 bgr_0.Vin-.n0 GNDA 0.069747f
C456 bgr_0.Vin-.n1 GNDA 0.316148f
C457 bgr_0.Vin-.t7 GNDA 0.027101f
C458 bgr_0.Vin-.t5 GNDA 0.027101f
C459 bgr_0.Vin-.n2 GNDA 0.094346f
C460 bgr_0.Vin-.t4 GNDA 0.027101f
C461 bgr_0.Vin-.t6 GNDA 0.027101f
C462 bgr_0.Vin-.n3 GNDA 0.090091f
C463 bgr_0.Vin-.n4 GNDA 0.386489f
C464 bgr_0.Vin-.n5 GNDA 0.027681f
C465 bgr_0.Vin-.n6 GNDA 0.366254f
C466 bgr_0.Vin-.t12 GNDA 0.022346f
C467 bgr_0.Vin-.n7 GNDA 0.026209f
C468 bgr_0.Vin-.n8 GNDA 0.021455f
C469 bgr_0.Vin-.n9 GNDA 0.021455f
C470 bgr_0.Vin-.n10 GNDA 0.036491f
C471 bgr_0.Vin-.n11 GNDA 0.497932f
C472 bgr_0.Vin-.t0 GNDA 0.117924f
C473 bgr_0.Vin-.n12 GNDA 0.655831f
C474 bgr_0.Vin-.n13 GNDA 1.07297f
C475 bgr_0.Vin-.n14 GNDA 0.471323f
C476 bgr_0.Vin-.t3 GNDA 0.261631f
C477 bgr_0.Vin-.n15 GNDA 0.069875f
C478 bgr_0.Vin-.n16 GNDA 0.119593f
C479 bgr_0.Vin-.n17 GNDA 0.07053f
C480 bgr_0.Vin-.n18 GNDA 0.579028f
C481 bgr_0.Vin-.n19 GNDA 0.358216f
C482 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter GNDA 0.086538f
C483 bgr_0.V_mir2.t12 GNDA 0.03537f
C484 bgr_0.V_mir2.t3 GNDA 0.017685f
C485 bgr_0.V_mir2.t1 GNDA 0.017685f
C486 bgr_0.V_mir2.n0 GNDA 0.046242f
C487 bgr_0.V_mir2.t2 GNDA 0.075466f
C488 bgr_0.V_mir2.t4 GNDA 0.017685f
C489 bgr_0.V_mir2.t0 GNDA 0.017685f
C490 bgr_0.V_mir2.n1 GNDA 0.050199f
C491 bgr_0.V_mir2.n2 GNDA 0.827814f
C492 bgr_0.V_mir2.n3 GNDA 0.268286f
C493 bgr_0.V_mir2.t9 GNDA 0.042444f
C494 bgr_0.V_mir2.t17 GNDA 0.042444f
C495 bgr_0.V_mir2.t20 GNDA 0.06851f
C496 bgr_0.V_mir2.n4 GNDA 0.076506f
C497 bgr_0.V_mir2.n5 GNDA 0.052264f
C498 bgr_0.V_mir2.t5 GNDA 0.053881f
C499 bgr_0.V_mir2.n6 GNDA 0.081315f
C500 bgr_0.V_mir2.t10 GNDA 0.03537f
C501 bgr_0.V_mir2.t6 GNDA 0.03537f
C502 bgr_0.V_mir2.n7 GNDA 0.08097f
C503 bgr_0.V_mir2.n8 GNDA 0.201563f
C504 bgr_0.V_mir2.t7 GNDA 0.042444f
C505 bgr_0.V_mir2.t18 GNDA 0.042444f
C506 bgr_0.V_mir2.t22 GNDA 0.06851f
C507 bgr_0.V_mir2.n9 GNDA 0.076506f
C508 bgr_0.V_mir2.n10 GNDA 0.052264f
C509 bgr_0.V_mir2.t13 GNDA 0.053881f
C510 bgr_0.V_mir2.n11 GNDA 0.081315f
C511 bgr_0.V_mir2.t8 GNDA 0.03537f
C512 bgr_0.V_mir2.t14 GNDA 0.03537f
C513 bgr_0.V_mir2.n12 GNDA 0.08097f
C514 bgr_0.V_mir2.n13 GNDA 0.203577f
C515 bgr_0.V_mir2.n14 GNDA 0.699157f
C516 bgr_0.V_mir2.n15 GNDA 0.09373f
C517 bgr_0.V_mir2.t11 GNDA 0.042444f
C518 bgr_0.V_mir2.t19 GNDA 0.042444f
C519 bgr_0.V_mir2.t21 GNDA 0.06851f
C520 bgr_0.V_mir2.n16 GNDA 0.076506f
C521 bgr_0.V_mir2.n17 GNDA 0.052264f
C522 bgr_0.V_mir2.t15 GNDA 0.053881f
C523 bgr_0.V_mir2.n18 GNDA 0.081315f
C524 bgr_0.V_mir2.n19 GNDA 0.156007f
C525 bgr_0.V_mir2.n20 GNDA 0.08097f
C526 bgr_0.V_mir2.t16 GNDA 0.03537f
C527 bgr_0.cap_res1.t12 GNDA 0.331712f
C528 bgr_0.cap_res1.t19 GNDA 0.349187f
C529 bgr_0.cap_res1.t16 GNDA 0.350452f
C530 bgr_0.cap_res1.t5 GNDA 0.331712f
C531 bgr_0.cap_res1.t15 GNDA 0.349187f
C532 bgr_0.cap_res1.t9 GNDA 0.350452f
C533 bgr_0.cap_res1.t11 GNDA 0.331712f
C534 bgr_0.cap_res1.t18 GNDA 0.349187f
C535 bgr_0.cap_res1.t14 GNDA 0.350452f
C536 bgr_0.cap_res1.t4 GNDA 0.331712f
C537 bgr_0.cap_res1.t13 GNDA 0.349187f
C538 bgr_0.cap_res1.t7 GNDA 0.350452f
C539 bgr_0.cap_res1.t20 GNDA 0.331712f
C540 bgr_0.cap_res1.t6 GNDA 0.349187f
C541 bgr_0.cap_res1.t1 GNDA 0.350452f
C542 bgr_0.cap_res1.n0 GNDA 0.23406f
C543 bgr_0.cap_res1.t17 GNDA 0.186395f
C544 bgr_0.cap_res1.n1 GNDA 0.253961f
C545 bgr_0.cap_res1.t2 GNDA 0.186395f
C546 bgr_0.cap_res1.n2 GNDA 0.253961f
C547 bgr_0.cap_res1.t8 GNDA 0.186395f
C548 bgr_0.cap_res1.n3 GNDA 0.253961f
C549 bgr_0.cap_res1.t3 GNDA 0.186395f
C550 bgr_0.cap_res1.n4 GNDA 0.253961f
C551 bgr_0.cap_res1.t10 GNDA 0.363549f
C552 bgr_0.cap_res1.t0 GNDA 0.08421f
C553 two_stage_opamp_dummy_magic_0.cap_res_X.t90 GNDA 0.344645f
C554 two_stage_opamp_dummy_magic_0.cap_res_X.t127 GNDA 0.345894f
C555 two_stage_opamp_dummy_magic_0.cap_res_X.t49 GNDA 0.344645f
C556 two_stage_opamp_dummy_magic_0.cap_res_X.t88 GNDA 0.347347f
C557 two_stage_opamp_dummy_magic_0.cap_res_X.t67 GNDA 0.37779f
C558 two_stage_opamp_dummy_magic_0.cap_res_X.t130 GNDA 0.344645f
C559 two_stage_opamp_dummy_magic_0.cap_res_X.t27 GNDA 0.345894f
C560 two_stage_opamp_dummy_magic_0.cap_res_X.t81 GNDA 0.344645f
C561 two_stage_opamp_dummy_magic_0.cap_res_X.t42 GNDA 0.345894f
C562 two_stage_opamp_dummy_magic_0.cap_res_X.t95 GNDA 0.344645f
C563 two_stage_opamp_dummy_magic_0.cap_res_X.t134 GNDA 0.345894f
C564 two_stage_opamp_dummy_magic_0.cap_res_X.t45 GNDA 0.344645f
C565 two_stage_opamp_dummy_magic_0.cap_res_X.t9 GNDA 0.345894f
C566 two_stage_opamp_dummy_magic_0.cap_res_X.t43 GNDA 0.344645f
C567 two_stage_opamp_dummy_magic_0.cap_res_X.t79 GNDA 0.345894f
C568 two_stage_opamp_dummy_magic_0.cap_res_X.t58 GNDA 0.344645f
C569 two_stage_opamp_dummy_magic_0.cap_res_X.t25 GNDA 0.345894f
C570 two_stage_opamp_dummy_magic_0.cap_res_X.t83 GNDA 0.344645f
C571 two_stage_opamp_dummy_magic_0.cap_res_X.t118 GNDA 0.345894f
C572 two_stage_opamp_dummy_magic_0.cap_res_X.t102 GNDA 0.344645f
C573 two_stage_opamp_dummy_magic_0.cap_res_X.t65 GNDA 0.345894f
C574 two_stage_opamp_dummy_magic_0.cap_res_X.t48 GNDA 0.344645f
C575 two_stage_opamp_dummy_magic_0.cap_res_X.t86 GNDA 0.345894f
C576 two_stage_opamp_dummy_magic_0.cap_res_X.t66 GNDA 0.344645f
C577 two_stage_opamp_dummy_magic_0.cap_res_X.t31 GNDA 0.345894f
C578 two_stage_opamp_dummy_magic_0.cap_res_X.t89 GNDA 0.344645f
C579 two_stage_opamp_dummy_magic_0.cap_res_X.t124 GNDA 0.345894f
C580 two_stage_opamp_dummy_magic_0.cap_res_X.t105 GNDA 0.344645f
C581 two_stage_opamp_dummy_magic_0.cap_res_X.t69 GNDA 0.345894f
C582 two_stage_opamp_dummy_magic_0.cap_res_X.t128 GNDA 0.344645f
C583 two_stage_opamp_dummy_magic_0.cap_res_X.t22 GNDA 0.345894f
C584 two_stage_opamp_dummy_magic_0.cap_res_X.t4 GNDA 0.344645f
C585 two_stage_opamp_dummy_magic_0.cap_res_X.t109 GNDA 0.345894f
C586 two_stage_opamp_dummy_magic_0.cap_res_X.t94 GNDA 0.344645f
C587 two_stage_opamp_dummy_magic_0.cap_res_X.t129 GNDA 0.345894f
C588 two_stage_opamp_dummy_magic_0.cap_res_X.t111 GNDA 0.344645f
C589 two_stage_opamp_dummy_magic_0.cap_res_X.t76 GNDA 0.345894f
C590 two_stage_opamp_dummy_magic_0.cap_res_X.t135 GNDA 0.344645f
C591 two_stage_opamp_dummy_magic_0.cap_res_X.t28 GNDA 0.345894f
C592 two_stage_opamp_dummy_magic_0.cap_res_X.t11 GNDA 0.344645f
C593 two_stage_opamp_dummy_magic_0.cap_res_X.t117 GNDA 0.345894f
C594 two_stage_opamp_dummy_magic_0.cap_res_X.t34 GNDA 0.344645f
C595 two_stage_opamp_dummy_magic_0.cap_res_X.t68 GNDA 0.345894f
C596 two_stage_opamp_dummy_magic_0.cap_res_X.t50 GNDA 0.344645f
C597 two_stage_opamp_dummy_magic_0.cap_res_X.t16 GNDA 0.345894f
C598 two_stage_opamp_dummy_magic_0.cap_res_X.t73 GNDA 0.344645f
C599 two_stage_opamp_dummy_magic_0.cap_res_X.t108 GNDA 0.345894f
C600 two_stage_opamp_dummy_magic_0.cap_res_X.t91 GNDA 0.344645f
C601 two_stage_opamp_dummy_magic_0.cap_res_X.t54 GNDA 0.345894f
C602 two_stage_opamp_dummy_magic_0.cap_res_X.t36 GNDA 0.344645f
C603 two_stage_opamp_dummy_magic_0.cap_res_X.t74 GNDA 0.345894f
C604 two_stage_opamp_dummy_magic_0.cap_res_X.t53 GNDA 0.344645f
C605 two_stage_opamp_dummy_magic_0.cap_res_X.t20 GNDA 0.345894f
C606 two_stage_opamp_dummy_magic_0.cap_res_X.t78 GNDA 0.344645f
C607 two_stage_opamp_dummy_magic_0.cap_res_X.t116 GNDA 0.345894f
C608 two_stage_opamp_dummy_magic_0.cap_res_X.t97 GNDA 0.344645f
C609 two_stage_opamp_dummy_magic_0.cap_res_X.t57 GNDA 0.345894f
C610 two_stage_opamp_dummy_magic_0.cap_res_X.t120 GNDA 0.344645f
C611 two_stage_opamp_dummy_magic_0.cap_res_X.t15 GNDA 0.345894f
C612 two_stage_opamp_dummy_magic_0.cap_res_X.t137 GNDA 0.344645f
C613 two_stage_opamp_dummy_magic_0.cap_res_X.t100 GNDA 0.345894f
C614 two_stage_opamp_dummy_magic_0.cap_res_X.t85 GNDA 0.344645f
C615 two_stage_opamp_dummy_magic_0.cap_res_X.t119 GNDA 0.345894f
C616 two_stage_opamp_dummy_magic_0.cap_res_X.t84 GNDA 0.344645f
C617 two_stage_opamp_dummy_magic_0.cap_res_X.t8 GNDA 0.361543f
C618 two_stage_opamp_dummy_magic_0.cap_res_X.t41 GNDA 0.344645f
C619 two_stage_opamp_dummy_magic_0.cap_res_X.t99 GNDA 0.185116f
C620 two_stage_opamp_dummy_magic_0.cap_res_X.n0 GNDA 0.19812f
C621 two_stage_opamp_dummy_magic_0.cap_res_X.t93 GNDA 0.344645f
C622 two_stage_opamp_dummy_magic_0.cap_res_X.t60 GNDA 0.185116f
C623 two_stage_opamp_dummy_magic_0.cap_res_X.n1 GNDA 0.196522f
C624 two_stage_opamp_dummy_magic_0.cap_res_X.t3 GNDA 0.344645f
C625 two_stage_opamp_dummy_magic_0.cap_res_X.t26 GNDA 0.185116f
C626 two_stage_opamp_dummy_magic_0.cap_res_X.n2 GNDA 0.196522f
C627 two_stage_opamp_dummy_magic_0.cap_res_X.t51 GNDA 0.344645f
C628 two_stage_opamp_dummy_magic_0.cap_res_X.t133 GNDA 0.185116f
C629 two_stage_opamp_dummy_magic_0.cap_res_X.n3 GNDA 0.196522f
C630 two_stage_opamp_dummy_magic_0.cap_res_X.t14 GNDA 0.344645f
C631 two_stage_opamp_dummy_magic_0.cap_res_X.t82 GNDA 0.185116f
C632 two_stage_opamp_dummy_magic_0.cap_res_X.n4 GNDA 0.196522f
C633 two_stage_opamp_dummy_magic_0.cap_res_X.t61 GNDA 0.344645f
C634 two_stage_opamp_dummy_magic_0.cap_res_X.t44 GNDA 0.185116f
C635 two_stage_opamp_dummy_magic_0.cap_res_X.n5 GNDA 0.196522f
C636 two_stage_opamp_dummy_magic_0.cap_res_X.t115 GNDA 0.344645f
C637 two_stage_opamp_dummy_magic_0.cap_res_X.t13 GNDA 0.185116f
C638 two_stage_opamp_dummy_magic_0.cap_res_X.n6 GNDA 0.196522f
C639 two_stage_opamp_dummy_magic_0.cap_res_X.t71 GNDA 0.344645f
C640 two_stage_opamp_dummy_magic_0.cap_res_X.t103 GNDA 0.185116f
C641 two_stage_opamp_dummy_magic_0.cap_res_X.n7 GNDA 0.196522f
C642 two_stage_opamp_dummy_magic_0.cap_res_X.t123 GNDA 0.344645f
C643 two_stage_opamp_dummy_magic_0.cap_res_X.t63 GNDA 0.185116f
C644 two_stage_opamp_dummy_magic_0.cap_res_X.n8 GNDA 0.196522f
C645 two_stage_opamp_dummy_magic_0.cap_res_X.t40 GNDA 0.344645f
C646 two_stage_opamp_dummy_magic_0.cap_res_X.t132 GNDA 0.345894f
C647 two_stage_opamp_dummy_magic_0.cap_res_X.t33 GNDA 0.166619f
C648 two_stage_opamp_dummy_magic_0.cap_res_X.n9 GNDA 0.214914f
C649 two_stage_opamp_dummy_magic_0.cap_res_X.t30 GNDA 0.18397f
C650 two_stage_opamp_dummy_magic_0.cap_res_X.n10 GNDA 0.23341f
C651 two_stage_opamp_dummy_magic_0.cap_res_X.t64 GNDA 0.18397f
C652 two_stage_opamp_dummy_magic_0.cap_res_X.n11 GNDA 0.250658f
C653 two_stage_opamp_dummy_magic_0.cap_res_X.t24 GNDA 0.18397f
C654 two_stage_opamp_dummy_magic_0.cap_res_X.n12 GNDA 0.250658f
C655 two_stage_opamp_dummy_magic_0.cap_res_X.t126 GNDA 0.18397f
C656 two_stage_opamp_dummy_magic_0.cap_res_X.n13 GNDA 0.250658f
C657 two_stage_opamp_dummy_magic_0.cap_res_X.t19 GNDA 0.18397f
C658 two_stage_opamp_dummy_magic_0.cap_res_X.n14 GNDA 0.250658f
C659 two_stage_opamp_dummy_magic_0.cap_res_X.t122 GNDA 0.18397f
C660 two_stage_opamp_dummy_magic_0.cap_res_X.n15 GNDA 0.250658f
C661 two_stage_opamp_dummy_magic_0.cap_res_X.t80 GNDA 0.18397f
C662 two_stage_opamp_dummy_magic_0.cap_res_X.n16 GNDA 0.250658f
C663 two_stage_opamp_dummy_magic_0.cap_res_X.t37 GNDA 0.18397f
C664 two_stage_opamp_dummy_magic_0.cap_res_X.n17 GNDA 0.250658f
C665 two_stage_opamp_dummy_magic_0.cap_res_X.t75 GNDA 0.18397f
C666 two_stage_opamp_dummy_magic_0.cap_res_X.n18 GNDA 0.250658f
C667 two_stage_opamp_dummy_magic_0.cap_res_X.t35 GNDA 0.18397f
C668 two_stage_opamp_dummy_magic_0.cap_res_X.n19 GNDA 0.250658f
C669 two_stage_opamp_dummy_magic_0.cap_res_X.t138 GNDA 0.18397f
C670 two_stage_opamp_dummy_magic_0.cap_res_X.n20 GNDA 0.250658f
C671 two_stage_opamp_dummy_magic_0.cap_res_X.t29 GNDA 0.18397f
C672 two_stage_opamp_dummy_magic_0.cap_res_X.n21 GNDA 0.250658f
C673 two_stage_opamp_dummy_magic_0.cap_res_X.t131 GNDA 0.18397f
C674 two_stage_opamp_dummy_magic_0.cap_res_X.n22 GNDA 0.250658f
C675 two_stage_opamp_dummy_magic_0.cap_res_X.t110 GNDA 0.18397f
C676 two_stage_opamp_dummy_magic_0.cap_res_X.n23 GNDA 0.250658f
C677 two_stage_opamp_dummy_magic_0.cap_res_X.t5 GNDA 0.18397f
C678 two_stage_opamp_dummy_magic_0.cap_res_X.n24 GNDA 0.250658f
C679 two_stage_opamp_dummy_magic_0.cap_res_X.t106 GNDA 0.18397f
C680 two_stage_opamp_dummy_magic_0.cap_res_X.n25 GNDA 0.23341f
C681 two_stage_opamp_dummy_magic_0.cap_res_X.t104 GNDA 0.343499f
C682 two_stage_opamp_dummy_magic_0.cap_res_X.t2 GNDA 0.166619f
C683 two_stage_opamp_dummy_magic_0.cap_res_X.n26 GNDA 0.216163f
C684 two_stage_opamp_dummy_magic_0.cap_res_X.t1 GNDA 0.343499f
C685 two_stage_opamp_dummy_magic_0.cap_res_X.t38 GNDA 0.166619f
C686 two_stage_opamp_dummy_magic_0.cap_res_X.n27 GNDA 0.216163f
C687 two_stage_opamp_dummy_magic_0.cap_res_X.t121 GNDA 0.343499f
C688 two_stage_opamp_dummy_magic_0.cap_res_X.t113 GNDA 0.344645f
C689 two_stage_opamp_dummy_magic_0.cap_res_X.t21 GNDA 0.363141f
C690 two_stage_opamp_dummy_magic_0.cap_res_X.t56 GNDA 0.363141f
C691 two_stage_opamp_dummy_magic_0.cap_res_X.t18 GNDA 0.185116f
C692 two_stage_opamp_dummy_magic_0.cap_res_X.n28 GNDA 0.216163f
C693 two_stage_opamp_dummy_magic_0.cap_res_X.t125 GNDA 0.343499f
C694 two_stage_opamp_dummy_magic_0.cap_res_X.t62 GNDA 0.344645f
C695 two_stage_opamp_dummy_magic_0.cap_res_X.t23 GNDA 0.185116f
C696 two_stage_opamp_dummy_magic_0.cap_res_X.n29 GNDA 0.197667f
C697 two_stage_opamp_dummy_magic_0.cap_res_X.t7 GNDA 0.343499f
C698 two_stage_opamp_dummy_magic_0.cap_res_X.t87 GNDA 0.344645f
C699 two_stage_opamp_dummy_magic_0.cap_res_X.t46 GNDA 0.185116f
C700 two_stage_opamp_dummy_magic_0.cap_res_X.n30 GNDA 0.216163f
C701 two_stage_opamp_dummy_magic_0.cap_res_X.t107 GNDA 0.343499f
C702 two_stage_opamp_dummy_magic_0.cap_res_X.t47 GNDA 0.344645f
C703 two_stage_opamp_dummy_magic_0.cap_res_X.t10 GNDA 0.185116f
C704 two_stage_opamp_dummy_magic_0.cap_res_X.n31 GNDA 0.216163f
C705 two_stage_opamp_dummy_magic_0.cap_res_X.t70 GNDA 0.343499f
C706 two_stage_opamp_dummy_magic_0.cap_res_X.t12 GNDA 0.344645f
C707 two_stage_opamp_dummy_magic_0.cap_res_X.t112 GNDA 0.185116f
C708 two_stage_opamp_dummy_magic_0.cap_res_X.n32 GNDA 0.216163f
C709 two_stage_opamp_dummy_magic_0.cap_res_X.t32 GNDA 0.343499f
C710 two_stage_opamp_dummy_magic_0.cap_res_X.t92 GNDA 0.344645f
C711 two_stage_opamp_dummy_magic_0.cap_res_X.t77 GNDA 0.363141f
C712 two_stage_opamp_dummy_magic_0.cap_res_X.t114 GNDA 0.363141f
C713 two_stage_opamp_dummy_magic_0.cap_res_X.t72 GNDA 0.185116f
C714 two_stage_opamp_dummy_magic_0.cap_res_X.n33 GNDA 0.216163f
C715 two_stage_opamp_dummy_magic_0.cap_res_X.t52 GNDA 0.343499f
C716 two_stage_opamp_dummy_magic_0.cap_res_X.t39 GNDA 0.344645f
C717 two_stage_opamp_dummy_magic_0.cap_res_X.t101 GNDA 0.363141f
C718 two_stage_opamp_dummy_magic_0.cap_res_X.t136 GNDA 0.363141f
C719 two_stage_opamp_dummy_magic_0.cap_res_X.t96 GNDA 0.185116f
C720 two_stage_opamp_dummy_magic_0.cap_res_X.n34 GNDA 0.216163f
C721 two_stage_opamp_dummy_magic_0.cap_res_X.t17 GNDA 0.343499f
C722 two_stage_opamp_dummy_magic_0.cap_res_X.n35 GNDA 0.216163f
C723 two_stage_opamp_dummy_magic_0.cap_res_X.t55 GNDA 0.185116f
C724 two_stage_opamp_dummy_magic_0.cap_res_X.t98 GNDA 0.363141f
C725 two_stage_opamp_dummy_magic_0.cap_res_X.t59 GNDA 0.363141f
C726 two_stage_opamp_dummy_magic_0.cap_res_X.t6 GNDA 0.764814f
C727 two_stage_opamp_dummy_magic_0.cap_res_X.t0 GNDA 0.3034f
C728 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 GNDA 0.019565f
C729 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 GNDA 0.019565f
C730 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 GNDA 0.01946f
C731 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 GNDA 0.132138f
C732 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 GNDA 0.110991f
C733 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 GNDA 0.015631f
C734 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 GNDA 0.027752f
C735 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 GNDA 0.020809f
C736 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 GNDA 0.020809f
C737 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 GNDA 0.020809f
C738 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 GNDA 0.020809f
C739 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 GNDA 0.020809f
C740 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 GNDA 0.020809f
C741 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 GNDA 0.020809f
C742 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 GNDA 0.020809f
C743 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 GNDA 0.020809f
C744 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 GNDA 0.024288f
C745 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 GNDA 0.022899f
C746 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 GNDA 0.014361f
C747 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 GNDA 0.014361f
C748 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 GNDA 0.014361f
C749 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 GNDA 0.014361f
C750 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 GNDA 0.014361f
C751 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 GNDA 0.014361f
C752 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 GNDA 0.014361f
C753 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 GNDA 0.012833f
C754 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 GNDA 0.020809f
C755 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 GNDA 0.020809f
C756 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 GNDA 0.020809f
C757 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 GNDA 0.020809f
C758 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 GNDA 0.020809f
C759 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 GNDA 0.020809f
C760 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 GNDA 0.020809f
C761 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 GNDA 0.020809f
C762 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 GNDA 0.020809f
C763 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 GNDA 0.024288f
C764 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 GNDA 0.022899f
C765 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 GNDA 0.014361f
C766 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 GNDA 0.014361f
C767 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 GNDA 0.014361f
C768 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 GNDA 0.014361f
C769 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 GNDA 0.014361f
C770 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 GNDA 0.014361f
C771 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 GNDA 0.014361f
C772 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 GNDA 0.012833f
C773 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 GNDA 0.032071f
C774 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 GNDA 0.011723f
C775 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 GNDA 0.011723f
C776 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 GNDA 0.023447f
C777 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 GNDA 0.091435f
C778 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 GNDA 0.011723f
C779 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 GNDA 0.011723f
C780 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 GNDA 0.042043f
C781 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 GNDA 0.734273f
C782 bgr_0.TAIL_CUR_MIR_BIAS GNDA 0.626546f
C783 bgr_0.PFET_GATE_10uA.t28 GNDA 0.025549f
C784 bgr_0.PFET_GATE_10uA.t20 GNDA 0.037767f
C785 bgr_0.PFET_GATE_10uA.n0 GNDA 0.041615f
C786 bgr_0.PFET_GATE_10uA.t15 GNDA 0.025549f
C787 bgr_0.PFET_GATE_10uA.t21 GNDA 0.037767f
C788 bgr_0.PFET_GATE_10uA.n1 GNDA 0.041615f
C789 bgr_0.PFET_GATE_10uA.n2 GNDA 0.050075f
C790 bgr_0.PFET_GATE_10uA.t19 GNDA 0.025549f
C791 bgr_0.PFET_GATE_10uA.t12 GNDA 0.037767f
C792 bgr_0.PFET_GATE_10uA.n3 GNDA 0.041615f
C793 bgr_0.PFET_GATE_10uA.t26 GNDA 0.025549f
C794 bgr_0.PFET_GATE_10uA.t13 GNDA 0.037767f
C795 bgr_0.PFET_GATE_10uA.n4 GNDA 0.041615f
C796 bgr_0.PFET_GATE_10uA.n5 GNDA 0.041749f
C797 bgr_0.PFET_GATE_10uA.t7 GNDA 0.38277f
C798 bgr_0.PFET_GATE_10uA.t0 GNDA 0.026204f
C799 bgr_0.PFET_GATE_10uA.t8 GNDA 0.026204f
C800 bgr_0.PFET_GATE_10uA.n6 GNDA 0.066974f
C801 bgr_0.PFET_GATE_10uA.t2 GNDA 0.026204f
C802 bgr_0.PFET_GATE_10uA.t4 GNDA 0.026204f
C803 bgr_0.PFET_GATE_10uA.n7 GNDA 0.065244f
C804 bgr_0.PFET_GATE_10uA.n8 GNDA 0.638167f
C805 bgr_0.PFET_GATE_10uA.t3 GNDA 0.026204f
C806 bgr_0.PFET_GATE_10uA.t5 GNDA 0.026204f
C807 bgr_0.PFET_GATE_10uA.n9 GNDA 0.065244f
C808 bgr_0.PFET_GATE_10uA.n10 GNDA 0.361874f
C809 bgr_0.PFET_GATE_10uA.n11 GNDA 0.738742f
C810 bgr_0.PFET_GATE_10uA.t9 GNDA 0.026204f
C811 bgr_0.PFET_GATE_10uA.t1 GNDA 0.026204f
C812 bgr_0.PFET_GATE_10uA.n12 GNDA 0.063197f
C813 bgr_0.PFET_GATE_10uA.n13 GNDA 0.337378f
C814 bgr_0.PFET_GATE_10uA.t6 GNDA 0.569585f
C815 bgr_0.PFET_GATE_10uA.t27 GNDA 0.02954f
C816 bgr_0.PFET_GATE_10uA.t14 GNDA 0.02954f
C817 bgr_0.PFET_GATE_10uA.n14 GNDA 0.085401f
C818 bgr_0.PFET_GATE_10uA.n15 GNDA 2.35162f
C819 bgr_0.PFET_GATE_10uA.n16 GNDA 0.945097f
C820 bgr_0.PFET_GATE_10uA.n17 GNDA 0.93005f
C821 bgr_0.PFET_GATE_10uA.t11 GNDA 0.025549f
C822 bgr_0.PFET_GATE_10uA.t25 GNDA 0.025549f
C823 bgr_0.PFET_GATE_10uA.t18 GNDA 0.025549f
C824 bgr_0.PFET_GATE_10uA.t10 GNDA 0.025549f
C825 bgr_0.PFET_GATE_10uA.t24 GNDA 0.025549f
C826 bgr_0.PFET_GATE_10uA.t17 GNDA 0.037767f
C827 bgr_0.PFET_GATE_10uA.n18 GNDA 0.046739f
C828 bgr_0.PFET_GATE_10uA.n19 GNDA 0.03341f
C829 bgr_0.PFET_GATE_10uA.n20 GNDA 0.03341f
C830 bgr_0.PFET_GATE_10uA.n21 GNDA 0.03341f
C831 bgr_0.PFET_GATE_10uA.n22 GNDA 0.028286f
C832 bgr_0.PFET_GATE_10uA.t16 GNDA 0.025549f
C833 bgr_0.PFET_GATE_10uA.t23 GNDA 0.025549f
C834 bgr_0.PFET_GATE_10uA.t22 GNDA 0.025549f
C835 bgr_0.PFET_GATE_10uA.t29 GNDA 0.037767f
C836 bgr_0.PFET_GATE_10uA.n23 GNDA 0.046739f
C837 bgr_0.PFET_GATE_10uA.n24 GNDA 0.03341f
C838 bgr_0.PFET_GATE_10uA.n25 GNDA 0.028286f
C839 bgr_0.PFET_GATE_10uA.n26 GNDA 0.038826f
C840 two_stage_opamp_dummy_magic_0.Vb1.t4 GNDA 0.024583f
C841 two_stage_opamp_dummy_magic_0.Vb1.t5 GNDA 0.024583f
C842 two_stage_opamp_dummy_magic_0.Vb1.n0 GNDA 0.061622f
C843 two_stage_opamp_dummy_magic_0.Vb1.t0 GNDA 0.024583f
C844 two_stage_opamp_dummy_magic_0.Vb1.t3 GNDA 0.024583f
C845 two_stage_opamp_dummy_magic_0.Vb1.n1 GNDA 0.061209f
C846 two_stage_opamp_dummy_magic_0.Vb1.n2 GNDA 0.672131f
C847 two_stage_opamp_dummy_magic_0.Vb1.t2 GNDA 0.112982f
C848 two_stage_opamp_dummy_magic_0.Vb1.t1 GNDA 0.744914f
C849 two_stage_opamp_dummy_magic_0.Vb1.n3 GNDA 1.05377f
C850 two_stage_opamp_dummy_magic_0.Vb1.t7 GNDA 0.037797f
C851 two_stage_opamp_dummy_magic_0.Vb1.t15 GNDA 0.037797f
C852 two_stage_opamp_dummy_magic_0.Vb1.t19 GNDA 0.037797f
C853 two_stage_opamp_dummy_magic_0.Vb1.t8 GNDA 0.037797f
C854 two_stage_opamp_dummy_magic_0.Vb1.t17 GNDA 0.049024f
C855 two_stage_opamp_dummy_magic_0.Vb1.n4 GNDA 0.053304f
C856 two_stage_opamp_dummy_magic_0.Vb1.n5 GNDA 0.035953f
C857 two_stage_opamp_dummy_magic_0.Vb1.n6 GNDA 0.035953f
C858 two_stage_opamp_dummy_magic_0.Vb1.n7 GNDA 0.031146f
C859 two_stage_opamp_dummy_magic_0.Vb1.t10 GNDA 0.037797f
C860 two_stage_opamp_dummy_magic_0.Vb1.t22 GNDA 0.037797f
C861 two_stage_opamp_dummy_magic_0.Vb1.t12 GNDA 0.037797f
C862 two_stage_opamp_dummy_magic_0.Vb1.t24 GNDA 0.037797f
C863 two_stage_opamp_dummy_magic_0.Vb1.t13 GNDA 0.049024f
C864 two_stage_opamp_dummy_magic_0.Vb1.n8 GNDA 0.053304f
C865 two_stage_opamp_dummy_magic_0.Vb1.n9 GNDA 0.035953f
C866 two_stage_opamp_dummy_magic_0.Vb1.n10 GNDA 0.035953f
C867 two_stage_opamp_dummy_magic_0.Vb1.n11 GNDA 0.031146f
C868 two_stage_opamp_dummy_magic_0.Vb1.n12 GNDA 0.045597f
C869 two_stage_opamp_dummy_magic_0.Vb1.t9 GNDA 0.037797f
C870 two_stage_opamp_dummy_magic_0.Vb1.t18 GNDA 0.037797f
C871 two_stage_opamp_dummy_magic_0.Vb1.t23 GNDA 0.037797f
C872 two_stage_opamp_dummy_magic_0.Vb1.t11 GNDA 0.037797f
C873 two_stage_opamp_dummy_magic_0.Vb1.t21 GNDA 0.049024f
C874 two_stage_opamp_dummy_magic_0.Vb1.n13 GNDA 0.053304f
C875 two_stage_opamp_dummy_magic_0.Vb1.n14 GNDA 0.035953f
C876 two_stage_opamp_dummy_magic_0.Vb1.n15 GNDA 0.035953f
C877 two_stage_opamp_dummy_magic_0.Vb1.n16 GNDA 0.031146f
C878 two_stage_opamp_dummy_magic_0.Vb1.t20 GNDA 0.037797f
C879 two_stage_opamp_dummy_magic_0.Vb1.t25 GNDA 0.037797f
C880 two_stage_opamp_dummy_magic_0.Vb1.t14 GNDA 0.037797f
C881 two_stage_opamp_dummy_magic_0.Vb1.t6 GNDA 0.037797f
C882 two_stage_opamp_dummy_magic_0.Vb1.t16 GNDA 0.049024f
C883 two_stage_opamp_dummy_magic_0.Vb1.n17 GNDA 0.053304f
C884 two_stage_opamp_dummy_magic_0.Vb1.n18 GNDA 0.035953f
C885 two_stage_opamp_dummy_magic_0.Vb1.n19 GNDA 0.035953f
C886 two_stage_opamp_dummy_magic_0.Vb1.n20 GNDA 0.031146f
C887 two_stage_opamp_dummy_magic_0.Vb1.n21 GNDA 0.034995f
C888 two_stage_opamp_dummy_magic_0.Vb1.n22 GNDA 0.842245f
C889 two_stage_opamp_dummy_magic_0.Vb1.n23 GNDA 2.21699f
C890 bgr_0.VB1_CUR_BIAS GNDA 1.32895f
C891 VOUT+.t17 GNDA 0.043627f
C892 VOUT+.t8 GNDA 0.043627f
C893 VOUT+.n0 GNDA 0.175348f
C894 VOUT+.t3 GNDA 0.043627f
C895 VOUT+.t7 GNDA 0.043627f
C896 VOUT+.n1 GNDA 0.175025f
C897 VOUT+.n2 GNDA 0.17242f
C898 VOUT+.t2 GNDA 0.043627f
C899 VOUT+.t6 GNDA 0.043627f
C900 VOUT+.n3 GNDA 0.175025f
C901 VOUT+.n4 GNDA 0.088916f
C902 VOUT+.t10 GNDA 0.043627f
C903 VOUT+.t4 GNDA 0.043627f
C904 VOUT+.n5 GNDA 0.175025f
C905 VOUT+.n6 GNDA 0.088916f
C906 VOUT+.t9 GNDA 0.043627f
C907 VOUT+.t18 GNDA 0.043627f
C908 VOUT+.n7 GNDA 0.175348f
C909 VOUT+.n8 GNDA 0.105318f
C910 VOUT+.t11 GNDA 0.043627f
C911 VOUT+.t5 GNDA 0.043627f
C912 VOUT+.n9 GNDA 0.172883f
C913 VOUT+.n10 GNDA 0.213802f
C914 VOUT+.t117 GNDA 0.295799f
C915 VOUT+.t25 GNDA 0.290845f
C916 VOUT+.n11 GNDA 0.195002f
C917 VOUT+.t124 GNDA 0.290845f
C918 VOUT+.n12 GNDA 0.127245f
C919 VOUT+.t72 GNDA 0.295799f
C920 VOUT+.t38 GNDA 0.290845f
C921 VOUT+.n13 GNDA 0.195002f
C922 VOUT+.t127 GNDA 0.290845f
C923 VOUT+.t34 GNDA 0.295178f
C924 VOUT+.t86 GNDA 0.295178f
C925 VOUT+.t42 GNDA 0.295178f
C926 VOUT+.t96 GNDA 0.295178f
C927 VOUT+.t143 GNDA 0.295178f
C928 VOUT+.t106 GNDA 0.295178f
C929 VOUT+.t154 GNDA 0.295178f
C930 VOUT+.t64 GNDA 0.295178f
C931 VOUT+.t116 GNDA 0.295178f
C932 VOUT+.t73 GNDA 0.295178f
C933 VOUT+.t149 GNDA 0.290845f
C934 VOUT+.n14 GNDA 0.195622f
C935 VOUT+.t58 GNDA 0.290845f
C936 VOUT+.n15 GNDA 0.250156f
C937 VOUT+.t97 GNDA 0.290845f
C938 VOUT+.n16 GNDA 0.250156f
C939 VOUT+.t131 GNDA 0.290845f
C940 VOUT+.n17 GNDA 0.250156f
C941 VOUT+.t24 GNDA 0.290845f
C942 VOUT+.n18 GNDA 0.250156f
C943 VOUT+.t75 GNDA 0.290845f
C944 VOUT+.n19 GNDA 0.250156f
C945 VOUT+.t113 GNDA 0.290845f
C946 VOUT+.n20 GNDA 0.250156f
C947 VOUT+.t144 GNDA 0.290845f
C948 VOUT+.n21 GNDA 0.250156f
C949 VOUT+.t54 GNDA 0.290845f
C950 VOUT+.n22 GNDA 0.250156f
C951 VOUT+.t94 GNDA 0.290845f
C952 VOUT+.n23 GNDA 0.250156f
C953 VOUT+.n24 GNDA 0.236312f
C954 VOUT+.t37 GNDA 0.295799f
C955 VOUT+.t142 GNDA 0.290845f
C956 VOUT+.n25 GNDA 0.195002f
C957 VOUT+.t93 GNDA 0.290845f
C958 VOUT+.t20 GNDA 0.295799f
C959 VOUT+.t57 GNDA 0.290845f
C960 VOUT+.n26 GNDA 0.195002f
C961 VOUT+.n27 GNDA 0.236312f
C962 VOUT+.t79 GNDA 0.295799f
C963 VOUT+.t41 GNDA 0.290845f
C964 VOUT+.n28 GNDA 0.195002f
C965 VOUT+.t133 GNDA 0.290845f
C966 VOUT+.t60 GNDA 0.295799f
C967 VOUT+.t100 GNDA 0.290845f
C968 VOUT+.n29 GNDA 0.195002f
C969 VOUT+.n30 GNDA 0.236312f
C970 VOUT+.t121 GNDA 0.295799f
C971 VOUT+.t83 GNDA 0.290845f
C972 VOUT+.n31 GNDA 0.195002f
C973 VOUT+.t31 GNDA 0.290845f
C974 VOUT+.t104 GNDA 0.295799f
C975 VOUT+.t137 GNDA 0.290845f
C976 VOUT+.n32 GNDA 0.195002f
C977 VOUT+.n33 GNDA 0.236312f
C978 VOUT+.t84 GNDA 0.295799f
C979 VOUT+.t49 GNDA 0.290845f
C980 VOUT+.n34 GNDA 0.195002f
C981 VOUT+.t138 GNDA 0.290845f
C982 VOUT+.t66 GNDA 0.295799f
C983 VOUT+.t103 GNDA 0.290845f
C984 VOUT+.n35 GNDA 0.195002f
C985 VOUT+.n36 GNDA 0.236312f
C986 VOUT+.t108 GNDA 0.295799f
C987 VOUT+.t69 GNDA 0.290845f
C988 VOUT+.n37 GNDA 0.195002f
C989 VOUT+.t90 GNDA 0.290845f
C990 VOUT+.n38 GNDA 0.127245f
C991 VOUT+.t67 GNDA 0.295799f
C992 VOUT+.t30 GNDA 0.290845f
C993 VOUT+.n39 GNDA 0.195002f
C994 VOUT+.t51 GNDA 0.290845f
C995 VOUT+.t53 GNDA 0.295178f
C996 VOUT+.t156 GNDA 0.295178f
C997 VOUT+.t44 GNDA 0.295799f
C998 VOUT+.t136 GNDA 0.290845f
C999 VOUT+.n40 GNDA 0.195002f
C1000 VOUT+.t101 GNDA 0.290845f
C1001 VOUT+.n41 GNDA 0.1227f
C1002 VOUT+.t36 GNDA 0.295178f
C1003 VOUT+.t151 GNDA 0.295799f
C1004 VOUT+.t98 GNDA 0.290845f
C1005 VOUT+.n42 GNDA 0.195002f
C1006 VOUT+.t59 GNDA 0.290845f
C1007 VOUT+.n43 GNDA 0.1227f
C1008 VOUT+.t140 GNDA 0.295178f
C1009 VOUT+.t118 GNDA 0.295799f
C1010 VOUT+.t56 GNDA 0.290845f
C1011 VOUT+.n44 GNDA 0.195002f
C1012 VOUT+.t21 GNDA 0.290845f
C1013 VOUT+.n45 GNDA 0.1227f
C1014 VOUT+.t105 GNDA 0.295178f
C1015 VOUT+.t65 GNDA 0.295799f
C1016 VOUT+.t80 GNDA 0.290845f
C1017 VOUT+.n46 GNDA 0.195002f
C1018 VOUT+.t43 GNDA 0.290845f
C1019 VOUT+.n47 GNDA 0.1227f
C1020 VOUT+.t125 GNDA 0.295178f
C1021 VOUT+.t145 GNDA 0.295422f
C1022 VOUT+.t87 GNDA 0.295178f
C1023 VOUT+.t110 GNDA 0.295422f
C1024 VOUT+.t50 GNDA 0.295178f
C1025 VOUT+.t70 GNDA 0.295422f
C1026 VOUT+.t150 GNDA 0.295178f
C1027 VOUT+.t95 GNDA 0.295422f
C1028 VOUT+.t32 GNDA 0.295178f
C1029 VOUT+.t134 GNDA 0.290845f
C1030 VOUT+.n48 GNDA 0.321926f
C1031 VOUT+.t111 GNDA 0.290845f
C1032 VOUT+.n49 GNDA 0.376459f
C1033 VOUT+.t147 GNDA 0.290845f
C1034 VOUT+.n50 GNDA 0.376459f
C1035 VOUT+.t45 GNDA 0.290845f
C1036 VOUT+.n51 GNDA 0.376459f
C1037 VOUT+.t85 GNDA 0.290845f
C1038 VOUT+.n52 GNDA 0.309234f
C1039 VOUT+.t61 GNDA 0.290845f
C1040 VOUT+.n53 GNDA 0.309234f
C1041 VOUT+.t102 GNDA 0.290845f
C1042 VOUT+.n54 GNDA 0.309234f
C1043 VOUT+.t139 GNDA 0.290845f
C1044 VOUT+.n55 GNDA 0.309234f
C1045 VOUT+.t119 GNDA 0.290845f
C1046 VOUT+.n56 GNDA 0.250156f
C1047 VOUT+.t155 GNDA 0.290845f
C1048 VOUT+.n57 GNDA 0.250156f
C1049 VOUT+.n58 GNDA 0.236312f
C1050 VOUT+.t27 GNDA 0.295799f
C1051 VOUT+.t130 GNDA 0.290845f
C1052 VOUT+.n59 GNDA 0.195002f
C1053 VOUT+.t152 GNDA 0.290845f
C1054 VOUT+.t76 GNDA 0.295799f
C1055 VOUT+.t115 GNDA 0.290845f
C1056 VOUT+.n60 GNDA 0.195002f
C1057 VOUT+.n61 GNDA 0.236312f
C1058 VOUT+.t62 GNDA 0.295799f
C1059 VOUT+.t23 GNDA 0.290845f
C1060 VOUT+.n62 GNDA 0.195002f
C1061 VOUT+.t47 GNDA 0.290845f
C1062 VOUT+.t112 GNDA 0.295799f
C1063 VOUT+.t148 GNDA 0.290845f
C1064 VOUT+.n63 GNDA 0.195002f
C1065 VOUT+.n64 GNDA 0.236312f
C1066 VOUT+.t114 GNDA 0.295799f
C1067 VOUT+.t78 GNDA 0.290845f
C1068 VOUT+.n65 GNDA 0.195002f
C1069 VOUT+.t26 GNDA 0.290845f
C1070 VOUT+.t99 GNDA 0.295799f
C1071 VOUT+.t132 GNDA 0.290845f
C1072 VOUT+.n66 GNDA 0.195002f
C1073 VOUT+.n67 GNDA 0.236312f
C1074 VOUT+.t74 GNDA 0.295799f
C1075 VOUT+.t39 GNDA 0.290845f
C1076 VOUT+.n68 GNDA 0.195002f
C1077 VOUT+.t128 GNDA 0.290845f
C1078 VOUT+.t55 GNDA 0.295799f
C1079 VOUT+.t92 GNDA 0.290845f
C1080 VOUT+.n69 GNDA 0.195002f
C1081 VOUT+.n70 GNDA 0.236312f
C1082 VOUT+.t109 GNDA 0.295799f
C1083 VOUT+.t71 GNDA 0.290845f
C1084 VOUT+.n71 GNDA 0.195002f
C1085 VOUT+.t19 GNDA 0.290845f
C1086 VOUT+.t91 GNDA 0.295799f
C1087 VOUT+.t126 GNDA 0.290845f
C1088 VOUT+.n72 GNDA 0.195002f
C1089 VOUT+.n73 GNDA 0.236312f
C1090 VOUT+.t68 GNDA 0.295799f
C1091 VOUT+.t33 GNDA 0.290845f
C1092 VOUT+.n74 GNDA 0.195002f
C1093 VOUT+.t122 GNDA 0.290845f
C1094 VOUT+.t52 GNDA 0.295799f
C1095 VOUT+.t88 GNDA 0.290845f
C1096 VOUT+.n75 GNDA 0.195002f
C1097 VOUT+.n76 GNDA 0.236312f
C1098 VOUT+.t29 GNDA 0.295799f
C1099 VOUT+.t135 GNDA 0.290845f
C1100 VOUT+.n77 GNDA 0.195002f
C1101 VOUT+.t82 GNDA 0.290845f
C1102 VOUT+.t153 GNDA 0.295799f
C1103 VOUT+.t48 GNDA 0.290845f
C1104 VOUT+.n78 GNDA 0.195002f
C1105 VOUT+.n79 GNDA 0.236312f
C1106 VOUT+.t63 GNDA 0.295799f
C1107 VOUT+.t28 GNDA 0.290845f
C1108 VOUT+.n80 GNDA 0.195002f
C1109 VOUT+.t120 GNDA 0.290845f
C1110 VOUT+.t46 GNDA 0.295799f
C1111 VOUT+.t81 GNDA 0.290845f
C1112 VOUT+.n81 GNDA 0.195002f
C1113 VOUT+.n82 GNDA 0.236312f
C1114 VOUT+.t22 GNDA 0.295799f
C1115 VOUT+.t129 GNDA 0.290845f
C1116 VOUT+.n83 GNDA 0.195002f
C1117 VOUT+.t77 GNDA 0.290845f
C1118 VOUT+.t146 GNDA 0.295799f
C1119 VOUT+.t40 GNDA 0.290845f
C1120 VOUT+.n84 GNDA 0.195002f
C1121 VOUT+.n85 GNDA 0.236312f
C1122 VOUT+.t123 GNDA 0.295799f
C1123 VOUT+.t89 GNDA 0.290845f
C1124 VOUT+.n86 GNDA 0.195002f
C1125 VOUT+.t35 GNDA 0.290845f
C1126 VOUT+.n87 GNDA 0.236312f
C1127 VOUT+.t141 GNDA 0.290845f
C1128 VOUT+.n88 GNDA 0.127245f
C1129 VOUT+.t107 GNDA 0.290845f
C1130 VOUT+.n89 GNDA 0.231292f
C1131 VOUT+.n90 GNDA 0.2787f
C1132 VOUT+.t12 GNDA 0.050898f
C1133 VOUT+.t16 GNDA 0.050898f
C1134 VOUT+.n91 GNDA 0.235456f
C1135 VOUT+.t13 GNDA 0.050898f
C1136 VOUT+.t1 GNDA 0.050898f
C1137 VOUT+.n92 GNDA 0.234668f
C1138 VOUT+.n93 GNDA 0.145013f
C1139 VOUT+.t15 GNDA 0.050898f
C1140 VOUT+.t14 GNDA 0.050898f
C1141 VOUT+.n94 GNDA 0.234668f
C1142 VOUT+.n95 GNDA 0.089261f
C1143 VOUT+.t0 GNDA 0.084152f
C1144 VOUT+.n96 GNDA 0.120712f
C1145 two_stage_opamp_dummy_magic_0.X.t16 GNDA 0.024316f
C1146 two_stage_opamp_dummy_magic_0.X.t15 GNDA 0.024316f
C1147 two_stage_opamp_dummy_magic_0.X.n0 GNDA 0.082095f
C1148 two_stage_opamp_dummy_magic_0.X.t19 GNDA 0.024316f
C1149 two_stage_opamp_dummy_magic_0.X.t21 GNDA 0.024316f
C1150 two_stage_opamp_dummy_magic_0.X.n1 GNDA 0.087741f
C1151 two_stage_opamp_dummy_magic_0.X.t0 GNDA 0.024316f
C1152 two_stage_opamp_dummy_magic_0.X.t18 GNDA 0.024316f
C1153 two_stage_opamp_dummy_magic_0.X.n2 GNDA 0.087741f
C1154 two_stage_opamp_dummy_magic_0.X.t22 GNDA 0.024316f
C1155 two_stage_opamp_dummy_magic_0.X.t14 GNDA 0.024316f
C1156 two_stage_opamp_dummy_magic_0.X.n3 GNDA 0.086975f
C1157 two_stage_opamp_dummy_magic_0.X.n4 GNDA 0.32294f
C1158 two_stage_opamp_dummy_magic_0.X.t3 GNDA 0.024316f
C1159 two_stage_opamp_dummy_magic_0.X.t20 GNDA 0.024316f
C1160 two_stage_opamp_dummy_magic_0.X.n5 GNDA 0.086975f
C1161 two_stage_opamp_dummy_magic_0.X.n6 GNDA 0.167527f
C1162 two_stage_opamp_dummy_magic_0.X.t17 GNDA 0.024316f
C1163 two_stage_opamp_dummy_magic_0.X.t23 GNDA 0.024316f
C1164 two_stage_opamp_dummy_magic_0.X.n7 GNDA 0.086975f
C1165 two_stage_opamp_dummy_magic_0.X.n8 GNDA 0.167527f
C1166 two_stage_opamp_dummy_magic_0.X.n9 GNDA 0.204045f
C1167 two_stage_opamp_dummy_magic_0.X.n10 GNDA 0.164936f
C1168 two_stage_opamp_dummy_magic_0.X.t1 GNDA 0.79195f
C1169 two_stage_opamp_dummy_magic_0.X.t36 GNDA 0.106988f
C1170 two_stage_opamp_dummy_magic_0.X.t49 GNDA 0.106988f
C1171 two_stage_opamp_dummy_magic_0.X.t34 GNDA 0.11395f
C1172 two_stage_opamp_dummy_magic_0.X.n11 GNDA 0.0903f
C1173 two_stage_opamp_dummy_magic_0.X.n12 GNDA 0.048273f
C1174 two_stage_opamp_dummy_magic_0.X.t51 GNDA 0.106988f
C1175 two_stage_opamp_dummy_magic_0.X.t39 GNDA 0.106988f
C1176 two_stage_opamp_dummy_magic_0.X.t26 GNDA 0.106988f
C1177 two_stage_opamp_dummy_magic_0.X.t44 GNDA 0.106988f
C1178 two_stage_opamp_dummy_magic_0.X.t25 GNDA 0.106988f
C1179 two_stage_opamp_dummy_magic_0.X.t43 GNDA 0.106988f
C1180 two_stage_opamp_dummy_magic_0.X.t29 GNDA 0.11395f
C1181 two_stage_opamp_dummy_magic_0.X.n13 GNDA 0.0903f
C1182 two_stage_opamp_dummy_magic_0.X.n14 GNDA 0.051063f
C1183 two_stage_opamp_dummy_magic_0.X.n15 GNDA 0.051063f
C1184 two_stage_opamp_dummy_magic_0.X.n16 GNDA 0.051063f
C1185 two_stage_opamp_dummy_magic_0.X.n17 GNDA 0.051063f
C1186 two_stage_opamp_dummy_magic_0.X.n18 GNDA 0.048273f
C1187 two_stage_opamp_dummy_magic_0.X.n19 GNDA 0.026157f
C1188 two_stage_opamp_dummy_magic_0.X.n20 GNDA 0.941428f
C1189 two_stage_opamp_dummy_magic_0.X.t7 GNDA 0.056736f
C1190 two_stage_opamp_dummy_magic_0.X.t2 GNDA 0.056736f
C1191 two_stage_opamp_dummy_magic_0.X.n21 GNDA 0.197316f
C1192 two_stage_opamp_dummy_magic_0.X.t5 GNDA 0.056736f
C1193 two_stage_opamp_dummy_magic_0.X.t8 GNDA 0.056736f
C1194 two_stage_opamp_dummy_magic_0.X.n22 GNDA 0.196617f
C1195 two_stage_opamp_dummy_magic_0.X.n23 GNDA 0.371194f
C1196 two_stage_opamp_dummy_magic_0.X.t10 GNDA 0.056736f
C1197 two_stage_opamp_dummy_magic_0.X.t11 GNDA 0.056736f
C1198 two_stage_opamp_dummy_magic_0.X.n24 GNDA 0.196617f
C1199 two_stage_opamp_dummy_magic_0.X.n25 GNDA 0.19243f
C1200 two_stage_opamp_dummy_magic_0.X.t6 GNDA 0.056736f
C1201 two_stage_opamp_dummy_magic_0.X.t4 GNDA 0.056736f
C1202 two_stage_opamp_dummy_magic_0.X.n26 GNDA 0.196617f
C1203 two_stage_opamp_dummy_magic_0.X.n27 GNDA 0.19243f
C1204 two_stage_opamp_dummy_magic_0.X.t9 GNDA 0.056736f
C1205 two_stage_opamp_dummy_magic_0.X.t13 GNDA 0.056736f
C1206 two_stage_opamp_dummy_magic_0.X.n28 GNDA 0.196617f
C1207 two_stage_opamp_dummy_magic_0.X.n29 GNDA 0.226591f
C1208 two_stage_opamp_dummy_magic_0.X.t24 GNDA 0.056736f
C1209 two_stage_opamp_dummy_magic_0.X.t12 GNDA 0.056736f
C1210 two_stage_opamp_dummy_magic_0.X.n30 GNDA 0.192544f
C1211 two_stage_opamp_dummy_magic_0.X.n31 GNDA 0.384076f
C1212 two_stage_opamp_dummy_magic_0.X.t53 GNDA 0.034042f
C1213 two_stage_opamp_dummy_magic_0.X.t42 GNDA 0.034042f
C1214 two_stage_opamp_dummy_magic_0.X.t54 GNDA 0.034042f
C1215 two_stage_opamp_dummy_magic_0.X.t38 GNDA 0.034042f
C1216 two_stage_opamp_dummy_magic_0.X.t50 GNDA 0.034042f
C1217 two_stage_opamp_dummy_magic_0.X.t35 GNDA 0.034042f
C1218 two_stage_opamp_dummy_magic_0.X.t48 GNDA 0.034042f
C1219 two_stage_opamp_dummy_magic_0.X.t33 GNDA 0.041336f
C1220 two_stage_opamp_dummy_magic_0.X.n32 GNDA 0.041336f
C1221 two_stage_opamp_dummy_magic_0.X.n33 GNDA 0.026747f
C1222 two_stage_opamp_dummy_magic_0.X.n34 GNDA 0.026747f
C1223 two_stage_opamp_dummy_magic_0.X.n35 GNDA 0.026747f
C1224 two_stage_opamp_dummy_magic_0.X.n36 GNDA 0.026747f
C1225 two_stage_opamp_dummy_magic_0.X.n37 GNDA 0.026747f
C1226 two_stage_opamp_dummy_magic_0.X.n38 GNDA 0.023958f
C1227 two_stage_opamp_dummy_magic_0.X.t41 GNDA 0.034042f
C1228 two_stage_opamp_dummy_magic_0.X.t28 GNDA 0.041336f
C1229 two_stage_opamp_dummy_magic_0.X.n39 GNDA 0.038547f
C1230 two_stage_opamp_dummy_magic_0.X.n40 GNDA 0.023563f
C1231 two_stage_opamp_dummy_magic_0.X.t30 GNDA 0.052278f
C1232 two_stage_opamp_dummy_magic_0.X.t47 GNDA 0.052278f
C1233 two_stage_opamp_dummy_magic_0.X.t31 GNDA 0.052278f
C1234 two_stage_opamp_dummy_magic_0.X.t45 GNDA 0.052278f
C1235 two_stage_opamp_dummy_magic_0.X.t27 GNDA 0.052278f
C1236 two_stage_opamp_dummy_magic_0.X.t40 GNDA 0.052278f
C1237 two_stage_opamp_dummy_magic_0.X.t52 GNDA 0.052278f
C1238 two_stage_opamp_dummy_magic_0.X.t37 GNDA 0.059432f
C1239 two_stage_opamp_dummy_magic_0.X.n41 GNDA 0.053635f
C1240 two_stage_opamp_dummy_magic_0.X.n42 GNDA 0.032826f
C1241 two_stage_opamp_dummy_magic_0.X.n43 GNDA 0.032826f
C1242 two_stage_opamp_dummy_magic_0.X.n44 GNDA 0.032826f
C1243 two_stage_opamp_dummy_magic_0.X.n45 GNDA 0.032826f
C1244 two_stage_opamp_dummy_magic_0.X.n46 GNDA 0.032826f
C1245 two_stage_opamp_dummy_magic_0.X.n47 GNDA 0.030036f
C1246 two_stage_opamp_dummy_magic_0.X.t46 GNDA 0.052278f
C1247 two_stage_opamp_dummy_magic_0.X.t32 GNDA 0.059432f
C1248 two_stage_opamp_dummy_magic_0.X.n48 GNDA 0.050846f
C1249 two_stage_opamp_dummy_magic_0.X.n49 GNDA 0.023513f
C1250 two_stage_opamp_dummy_magic_0.X.n50 GNDA 0.253421f
C1251 two_stage_opamp_dummy_magic_0.X.n51 GNDA 0.527686f
C1252 two_stage_opamp_dummy_magic_0.X.n52 GNDA 0.246145f
C1253 two_stage_opamp_dummy_magic_0.X.n53 GNDA 0.104986f
C1254 two_stage_opamp_dummy_magic_0.VD4.t15 GNDA 0.026025f
C1255 two_stage_opamp_dummy_magic_0.VD4.t19 GNDA 0.026025f
C1256 two_stage_opamp_dummy_magic_0.VD4.n0 GNDA 0.090508f
C1257 two_stage_opamp_dummy_magic_0.VD4.t23 GNDA 0.026025f
C1258 two_stage_opamp_dummy_magic_0.VD4.t7 GNDA 0.026025f
C1259 two_stage_opamp_dummy_magic_0.VD4.n1 GNDA 0.090188f
C1260 two_stage_opamp_dummy_magic_0.VD4.n2 GNDA 0.170266f
C1261 two_stage_opamp_dummy_magic_0.VD4.n3 GNDA 0.073371f
C1262 two_stage_opamp_dummy_magic_0.VD4.n4 GNDA 0.100747f
C1263 two_stage_opamp_dummy_magic_0.VD4.t2 GNDA 0.128386f
C1264 two_stage_opamp_dummy_magic_0.VD4.t0 GNDA 0.045318f
C1265 two_stage_opamp_dummy_magic_0.VD4.n5 GNDA 0.083755f
C1266 two_stage_opamp_dummy_magic_0.VD4.n6 GNDA 0.053992f
C1267 two_stage_opamp_dummy_magic_0.VD4.t5 GNDA 0.128386f
C1268 two_stage_opamp_dummy_magic_0.VD4.t3 GNDA 0.045318f
C1269 two_stage_opamp_dummy_magic_0.VD4.n7 GNDA 0.083755f
C1270 two_stage_opamp_dummy_magic_0.VD4.n8 GNDA 0.053992f
C1271 two_stage_opamp_dummy_magic_0.VD4.n9 GNDA 0.053537f
C1272 two_stage_opamp_dummy_magic_0.VD4.n10 GNDA 0.100747f
C1273 two_stage_opamp_dummy_magic_0.VD4.n11 GNDA 0.300245f
C1274 two_stage_opamp_dummy_magic_0.VD4.t4 GNDA 0.448159f
C1275 two_stage_opamp_dummy_magic_0.VD4.t14 GNDA 0.25876f
C1276 two_stage_opamp_dummy_magic_0.VD4.t18 GNDA 0.25876f
C1277 two_stage_opamp_dummy_magic_0.VD4.t22 GNDA 0.25876f
C1278 two_stage_opamp_dummy_magic_0.VD4.t6 GNDA 0.25876f
C1279 two_stage_opamp_dummy_magic_0.VD4.t10 GNDA 0.19407f
C1280 two_stage_opamp_dummy_magic_0.VD4.n12 GNDA 0.12938f
C1281 two_stage_opamp_dummy_magic_0.VD4.t12 GNDA 0.19407f
C1282 two_stage_opamp_dummy_magic_0.VD4.t16 GNDA 0.25876f
C1283 two_stage_opamp_dummy_magic_0.VD4.t20 GNDA 0.25876f
C1284 two_stage_opamp_dummy_magic_0.VD4.t24 GNDA 0.25876f
C1285 two_stage_opamp_dummy_magic_0.VD4.t8 GNDA 0.25876f
C1286 two_stage_opamp_dummy_magic_0.VD4.t1 GNDA 0.448159f
C1287 two_stage_opamp_dummy_magic_0.VD4.n13 GNDA 0.300245f
C1288 two_stage_opamp_dummy_magic_0.VD4.n14 GNDA 0.073371f
C1289 two_stage_opamp_dummy_magic_0.VD4.n15 GNDA 0.108171f
C1290 two_stage_opamp_dummy_magic_0.VD4.t11 GNDA 0.026025f
C1291 two_stage_opamp_dummy_magic_0.VD4.t13 GNDA 0.026025f
C1292 two_stage_opamp_dummy_magic_0.VD4.n16 GNDA 0.08832f
C1293 two_stage_opamp_dummy_magic_0.VD4.n17 GNDA 0.069277f
C1294 two_stage_opamp_dummy_magic_0.VD4.n18 GNDA 0.023794f
C1295 two_stage_opamp_dummy_magic_0.VD4.t17 GNDA 0.026025f
C1296 two_stage_opamp_dummy_magic_0.VD4.t21 GNDA 0.026025f
C1297 two_stage_opamp_dummy_magic_0.VD4.n19 GNDA 0.090188f
C1298 two_stage_opamp_dummy_magic_0.VD4.n20 GNDA 0.088268f
C1299 two_stage_opamp_dummy_magic_0.VD4.t25 GNDA 0.026025f
C1300 two_stage_opamp_dummy_magic_0.VD4.t9 GNDA 0.026025f
C1301 two_stage_opamp_dummy_magic_0.VD4.n21 GNDA 0.090188f
C1302 two_stage_opamp_dummy_magic_0.VD4.n22 GNDA 0.115584f
C1303 two_stage_opamp_dummy_magic_0.VD4.t34 GNDA 0.026025f
C1304 two_stage_opamp_dummy_magic_0.VD4.t37 GNDA 0.026025f
C1305 two_stage_opamp_dummy_magic_0.VD4.n23 GNDA 0.090509f
C1306 two_stage_opamp_dummy_magic_0.VD4.t30 GNDA 0.026025f
C1307 two_stage_opamp_dummy_magic_0.VD4.t32 GNDA 0.026025f
C1308 two_stage_opamp_dummy_magic_0.VD4.n24 GNDA 0.090188f
C1309 two_stage_opamp_dummy_magic_0.VD4.n25 GNDA 0.170266f
C1310 two_stage_opamp_dummy_magic_0.VD4.t26 GNDA 0.026025f
C1311 two_stage_opamp_dummy_magic_0.VD4.t28 GNDA 0.026025f
C1312 two_stage_opamp_dummy_magic_0.VD4.n26 GNDA 0.090188f
C1313 two_stage_opamp_dummy_magic_0.VD4.n27 GNDA 0.088268f
C1314 two_stage_opamp_dummy_magic_0.VD4.t33 GNDA 0.026025f
C1315 two_stage_opamp_dummy_magic_0.VD4.t35 GNDA 0.026025f
C1316 two_stage_opamp_dummy_magic_0.VD4.n28 GNDA 0.090188f
C1317 two_stage_opamp_dummy_magic_0.VD4.n29 GNDA 0.088268f
C1318 two_stage_opamp_dummy_magic_0.VD4.t29 GNDA 0.026025f
C1319 two_stage_opamp_dummy_magic_0.VD4.t31 GNDA 0.026025f
C1320 two_stage_opamp_dummy_magic_0.VD4.n30 GNDA 0.090188f
C1321 two_stage_opamp_dummy_magic_0.VD4.n31 GNDA 0.088268f
C1322 two_stage_opamp_dummy_magic_0.VD4.t36 GNDA 0.026025f
C1323 two_stage_opamp_dummy_magic_0.VD4.t27 GNDA 0.026025f
C1324 two_stage_opamp_dummy_magic_0.VD4.n32 GNDA 0.090188f
C1325 two_stage_opamp_dummy_magic_0.VD4.n33 GNDA 0.13596f
C1326 two_stage_opamp_dummy_magic_0.Vb2.n0 GNDA 0.010675f
C1327 two_stage_opamp_dummy_magic_0.Vb2.t0 GNDA 0.015714f
C1328 two_stage_opamp_dummy_magic_0.Vb2.n1 GNDA 0.067122f
C1329 two_stage_opamp_dummy_magic_0.Vb2.t20 GNDA 0.040575f
C1330 two_stage_opamp_dummy_magic_0.Vb2.t23 GNDA 0.040575f
C1331 two_stage_opamp_dummy_magic_0.Vb2.t21 GNDA 0.040575f
C1332 two_stage_opamp_dummy_magic_0.Vb2.t26 GNDA 0.040575f
C1333 two_stage_opamp_dummy_magic_0.Vb2.t31 GNDA 0.046824f
C1334 two_stage_opamp_dummy_magic_0.Vb2.n2 GNDA 0.038016f
C1335 two_stage_opamp_dummy_magic_0.Vb2.n3 GNDA 0.023362f
C1336 two_stage_opamp_dummy_magic_0.Vb2.n4 GNDA 0.023362f
C1337 two_stage_opamp_dummy_magic_0.Vb2.n5 GNDA 0.021875f
C1338 two_stage_opamp_dummy_magic_0.Vb2.t17 GNDA 0.040575f
C1339 two_stage_opamp_dummy_magic_0.Vb2.t30 GNDA 0.040575f
C1340 two_stage_opamp_dummy_magic_0.Vb2.t25 GNDA 0.040575f
C1341 two_stage_opamp_dummy_magic_0.Vb2.t27 GNDA 0.040575f
C1342 two_stage_opamp_dummy_magic_0.Vb2.t22 GNDA 0.046824f
C1343 two_stage_opamp_dummy_magic_0.Vb2.n6 GNDA 0.038016f
C1344 two_stage_opamp_dummy_magic_0.Vb2.n7 GNDA 0.023362f
C1345 two_stage_opamp_dummy_magic_0.Vb2.n8 GNDA 0.023362f
C1346 two_stage_opamp_dummy_magic_0.Vb2.n9 GNDA 0.021875f
C1347 two_stage_opamp_dummy_magic_0.Vb2.n10 GNDA 0.014849f
C1348 two_stage_opamp_dummy_magic_0.Vb2.t24 GNDA 0.040575f
C1349 two_stage_opamp_dummy_magic_0.Vb2.t29 GNDA 0.040575f
C1350 two_stage_opamp_dummy_magic_0.Vb2.t12 GNDA 0.040575f
C1351 two_stage_opamp_dummy_magic_0.Vb2.t14 GNDA 0.040575f
C1352 two_stage_opamp_dummy_magic_0.Vb2.t16 GNDA 0.046824f
C1353 two_stage_opamp_dummy_magic_0.Vb2.n11 GNDA 0.038016f
C1354 two_stage_opamp_dummy_magic_0.Vb2.n12 GNDA 0.023362f
C1355 two_stage_opamp_dummy_magic_0.Vb2.n13 GNDA 0.023362f
C1356 two_stage_opamp_dummy_magic_0.Vb2.n14 GNDA 0.021875f
C1357 two_stage_opamp_dummy_magic_0.Vb2.t18 GNDA 0.040575f
C1358 two_stage_opamp_dummy_magic_0.Vb2.t15 GNDA 0.040575f
C1359 two_stage_opamp_dummy_magic_0.Vb2.t13 GNDA 0.040575f
C1360 two_stage_opamp_dummy_magic_0.Vb2.t11 GNDA 0.040575f
C1361 two_stage_opamp_dummy_magic_0.Vb2.t28 GNDA 0.046824f
C1362 two_stage_opamp_dummy_magic_0.Vb2.n15 GNDA 0.038016f
C1363 two_stage_opamp_dummy_magic_0.Vb2.n16 GNDA 0.023362f
C1364 two_stage_opamp_dummy_magic_0.Vb2.n17 GNDA 0.023362f
C1365 two_stage_opamp_dummy_magic_0.Vb2.n18 GNDA 0.021875f
C1366 two_stage_opamp_dummy_magic_0.Vb2.n19 GNDA 0.014426f
C1367 two_stage_opamp_dummy_magic_0.Vb2.n20 GNDA 0.329391f
C1368 two_stage_opamp_dummy_magic_0.Vb2.n21 GNDA 0.247076f
C1369 two_stage_opamp_dummy_magic_0.Vb2.t19 GNDA 0.048957f
C1370 two_stage_opamp_dummy_magic_0.Vb2.n22 GNDA 0.684913f
C1371 two_stage_opamp_dummy_magic_0.Vb2.n23 GNDA 0.027105f
C1372 two_stage_opamp_dummy_magic_0.Vb2.n24 GNDA 0.747282f
C1373 two_stage_opamp_dummy_magic_0.Vb2.n25 GNDA 0.027105f
C1374 two_stage_opamp_dummy_magic_0.Vb2.n26 GNDA 0.190117f
C1375 two_stage_opamp_dummy_magic_0.Vb2.n27 GNDA 0.027926f
C1376 two_stage_opamp_dummy_magic_0.Vb2.n28 GNDA 0.281868f
C1377 two_stage_opamp_dummy_magic_0.Vb2.n29 GNDA 0.027105f
C1378 bgr_0.cap_res2.t6 GNDA 0.358376f
C1379 bgr_0.cap_res2.t12 GNDA 0.359675f
C1380 bgr_0.cap_res2.t14 GNDA 0.340442f
C1381 bgr_0.cap_res2.t0 GNDA 0.358376f
C1382 bgr_0.cap_res2.t5 GNDA 0.359675f
C1383 bgr_0.cap_res2.t8 GNDA 0.340442f
C1384 bgr_0.cap_res2.t4 GNDA 0.358376f
C1385 bgr_0.cap_res2.t10 GNDA 0.359675f
C1386 bgr_0.cap_res2.t13 GNDA 0.340442f
C1387 bgr_0.cap_res2.t19 GNDA 0.358376f
C1388 bgr_0.cap_res2.t3 GNDA 0.359675f
C1389 bgr_0.cap_res2.t7 GNDA 0.340442f
C1390 bgr_0.cap_res2.t15 GNDA 0.358376f
C1391 bgr_0.cap_res2.t18 GNDA 0.359675f
C1392 bgr_0.cap_res2.t1 GNDA 0.340442f
C1393 bgr_0.cap_res2.n0 GNDA 0.24022f
C1394 bgr_0.cap_res2.t2 GNDA 0.1913f
C1395 bgr_0.cap_res2.n1 GNDA 0.260644f
C1396 bgr_0.cap_res2.t9 GNDA 0.1913f
C1397 bgr_0.cap_res2.n2 GNDA 0.260644f
C1398 bgr_0.cap_res2.t16 GNDA 0.1913f
C1399 bgr_0.cap_res2.n3 GNDA 0.260644f
C1400 bgr_0.cap_res2.t11 GNDA 0.1913f
C1401 bgr_0.cap_res2.n4 GNDA 0.260644f
C1402 bgr_0.cap_res2.t17 GNDA 0.373116f
C1403 bgr_0.cap_res2.t20 GNDA 0.086426f
C1404 bgr_0.1st_Vout_2.n0 GNDA 0.720636f
C1405 bgr_0.1st_Vout_2.n1 GNDA 0.319289f
C1406 bgr_0.1st_Vout_2.n2 GNDA 1.80961f
C1407 bgr_0.1st_Vout_2.n3 GNDA 0.132034f
C1408 bgr_0.1st_Vout_2.n4 GNDA 1.84352f
C1409 bgr_0.1st_Vout_2.t33 GNDA 0.02189f
C1410 bgr_0.1st_Vout_2.t28 GNDA 0.364819f
C1411 bgr_0.1st_Vout_2.t17 GNDA 0.371033f
C1412 bgr_0.1st_Vout_2.t12 GNDA 0.364819f
C1413 bgr_0.1st_Vout_2.t32 GNDA 0.364819f
C1414 bgr_0.1st_Vout_2.t35 GNDA 0.371033f
C1415 bgr_0.1st_Vout_2.t11 GNDA 0.371033f
C1416 bgr_0.1st_Vout_2.t31 GNDA 0.364819f
C1417 bgr_0.1st_Vout_2.t23 GNDA 0.364819f
C1418 bgr_0.1st_Vout_2.t26 GNDA 0.371033f
C1419 bgr_0.1st_Vout_2.t30 GNDA 0.371033f
C1420 bgr_0.1st_Vout_2.t22 GNDA 0.364819f
C1421 bgr_0.1st_Vout_2.t15 GNDA 0.364819f
C1422 bgr_0.1st_Vout_2.t19 GNDA 0.371033f
C1423 bgr_0.1st_Vout_2.t36 GNDA 0.371033f
C1424 bgr_0.1st_Vout_2.t29 GNDA 0.364819f
C1425 bgr_0.1st_Vout_2.t21 GNDA 0.364819f
C1426 bgr_0.1st_Vout_2.t25 GNDA 0.371033f
C1427 bgr_0.1st_Vout_2.t18 GNDA 0.371033f
C1428 bgr_0.1st_Vout_2.t14 GNDA 0.364819f
C1429 bgr_0.1st_Vout_2.t20 GNDA 0.364819f
C1430 bgr_0.1st_Vout_2.t34 GNDA 0.023833f
C1431 bgr_0.1st_Vout_2.n5 GNDA 0.022991f
C1432 bgr_0.1st_Vout_2.t27 GNDA 0.013894f
C1433 bgr_0.1st_Vout_2.t16 GNDA 0.013894f
C1434 bgr_0.1st_Vout_2.n6 GNDA 0.030909f
C1435 bgr_0.1st_Vout_2.n7 GNDA 0.013175f
C1436 bgr_0.1st_Vout_2.t8 GNDA 0.01921f
C1437 bgr_0.1st_Vout_2.n8 GNDA 0.199276f
C1438 bgr_0.1st_Vout_2.n9 GNDA 0.01192f
C1439 bgr_0.1st_Vout_2.n10 GNDA 0.022038f
C1440 bgr_0.1st_Vout_2.t24 GNDA 0.013894f
C1441 bgr_0.1st_Vout_2.t13 GNDA 0.013894f
C1442 bgr_0.1st_Vout_2.n11 GNDA 0.030909f
C1443 bgr_0.1st_Vout_2.n12 GNDA 0.174923f
C1444 bgr_0.1st_Vout_2.n13 GNDA 0.022991f
C1445 two_stage_opamp_dummy_magic_0.V_err_gate.n0 GNDA 1.01381f
C1446 two_stage_opamp_dummy_magic_0.V_err_gate.n1 GNDA 2.13029f
C1447 two_stage_opamp_dummy_magic_0.V_err_gate.t8 GNDA 0.028502f
C1448 two_stage_opamp_dummy_magic_0.V_err_gate.t9 GNDA 0.028502f
C1449 two_stage_opamp_dummy_magic_0.V_err_gate.n2 GNDA 0.433389f
C1450 two_stage_opamp_dummy_magic_0.V_err_gate.t13 GNDA 0.014251f
C1451 two_stage_opamp_dummy_magic_0.V_err_gate.t10 GNDA 0.014251f
C1452 two_stage_opamp_dummy_magic_0.V_err_gate.n3 GNDA 0.033264f
C1453 two_stage_opamp_dummy_magic_0.V_err_gate.t3 GNDA 0.014251f
C1454 two_stage_opamp_dummy_magic_0.V_err_gate.t0 GNDA 0.014251f
C1455 two_stage_opamp_dummy_magic_0.V_err_gate.n4 GNDA 0.033049f
C1456 two_stage_opamp_dummy_magic_0.V_err_gate.t7 GNDA 0.014251f
C1457 two_stage_opamp_dummy_magic_0.V_err_gate.t5 GNDA 0.014251f
C1458 two_stage_opamp_dummy_magic_0.V_err_gate.n5 GNDA 0.033049f
C1459 two_stage_opamp_dummy_magic_0.V_err_gate.t23 GNDA 0.011757f
C1460 two_stage_opamp_dummy_magic_0.V_err_gate.t32 GNDA 0.011757f
C1461 two_stage_opamp_dummy_magic_0.V_err_gate.t21 GNDA 0.011757f
C1462 two_stage_opamp_dummy_magic_0.V_err_gate.t30 GNDA 0.011757f
C1463 two_stage_opamp_dummy_magic_0.V_err_gate.t16 GNDA 0.011757f
C1464 two_stage_opamp_dummy_magic_0.V_err_gate.t25 GNDA 0.011757f
C1465 two_stage_opamp_dummy_magic_0.V_err_gate.t18 GNDA 0.011757f
C1466 two_stage_opamp_dummy_magic_0.V_err_gate.t28 GNDA 0.011757f
C1467 two_stage_opamp_dummy_magic_0.V_err_gate.t15 GNDA 0.011757f
C1468 two_stage_opamp_dummy_magic_0.V_err_gate.t24 GNDA 0.011757f
C1469 two_stage_opamp_dummy_magic_0.V_err_gate.t33 GNDA 0.011757f
C1470 two_stage_opamp_dummy_magic_0.V_err_gate.t22 GNDA 0.011757f
C1471 two_stage_opamp_dummy_magic_0.V_err_gate.t31 GNDA 0.011757f
C1472 two_stage_opamp_dummy_magic_0.V_err_gate.t19 GNDA 0.011757f
C1473 two_stage_opamp_dummy_magic_0.V_err_gate.t26 GNDA 0.011757f
C1474 two_stage_opamp_dummy_magic_0.V_err_gate.t20 GNDA 0.011757f
C1475 two_stage_opamp_dummy_magic_0.V_err_gate.t29 GNDA 0.025473f
C1476 two_stage_opamp_dummy_magic_0.V_err_gate.n6 GNDA 0.039724f
C1477 two_stage_opamp_dummy_magic_0.V_err_gate.n7 GNDA 0.030995f
C1478 two_stage_opamp_dummy_magic_0.V_err_gate.n8 GNDA 0.030995f
C1479 two_stage_opamp_dummy_magic_0.V_err_gate.n9 GNDA 0.030995f
C1480 two_stage_opamp_dummy_magic_0.V_err_gate.n10 GNDA 0.030995f
C1481 two_stage_opamp_dummy_magic_0.V_err_gate.n11 GNDA 0.030995f
C1482 two_stage_opamp_dummy_magic_0.V_err_gate.n12 GNDA 0.030995f
C1483 two_stage_opamp_dummy_magic_0.V_err_gate.n13 GNDA 0.030995f
C1484 two_stage_opamp_dummy_magic_0.V_err_gate.n14 GNDA 0.030995f
C1485 two_stage_opamp_dummy_magic_0.V_err_gate.n15 GNDA 0.030995f
C1486 two_stage_opamp_dummy_magic_0.V_err_gate.n16 GNDA 0.030995f
C1487 two_stage_opamp_dummy_magic_0.V_err_gate.n17 GNDA 0.030995f
C1488 two_stage_opamp_dummy_magic_0.V_err_gate.n18 GNDA 0.030995f
C1489 two_stage_opamp_dummy_magic_0.V_err_gate.n19 GNDA 0.030995f
C1490 two_stage_opamp_dummy_magic_0.V_err_gate.n20 GNDA 0.030995f
C1491 two_stage_opamp_dummy_magic_0.V_err_gate.n21 GNDA 0.026524f
C1492 two_stage_opamp_dummy_magic_0.V_err_gate.t14 GNDA 0.011757f
C1493 two_stage_opamp_dummy_magic_0.V_err_gate.t27 GNDA 0.011757f
C1494 two_stage_opamp_dummy_magic_0.V_err_gate.t17 GNDA 0.025473f
C1495 two_stage_opamp_dummy_magic_0.V_err_gate.n22 GNDA 0.039724f
C1496 two_stage_opamp_dummy_magic_0.V_err_gate.n23 GNDA 0.026524f
C1497 two_stage_opamp_dummy_magic_0.V_err_gate.n24 GNDA 0.043031f
C1498 two_stage_opamp_dummy_magic_0.V_err_gate.t2 GNDA 0.014251f
C1499 two_stage_opamp_dummy_magic_0.V_err_gate.t4 GNDA 0.014251f
C1500 two_stage_opamp_dummy_magic_0.V_err_gate.n25 GNDA 0.028502f
C1501 two_stage_opamp_dummy_magic_0.V_err_gate.n26 GNDA 0.0849f
C1502 two_stage_opamp_dummy_magic_0.V_err_gate.t6 GNDA 0.014251f
C1503 two_stage_opamp_dummy_magic_0.V_err_gate.t12 GNDA 0.014251f
C1504 two_stage_opamp_dummy_magic_0.V_err_gate.n27 GNDA 0.033049f
C1505 two_stage_opamp_dummy_magic_0.V_err_gate.t11 GNDA 0.014251f
C1506 two_stage_opamp_dummy_magic_0.V_err_gate.t1 GNDA 0.014251f
C1507 two_stage_opamp_dummy_magic_0.V_err_gate.n28 GNDA 0.032803f
C1508 bgr_0.1st_Vout_1.n0 GNDA 0.629216f
C1509 bgr_0.1st_Vout_1.n1 GNDA 0.276014f
C1510 bgr_0.1st_Vout_1.n2 GNDA 1.1368f
C1511 bgr_0.1st_Vout_1.n3 GNDA 1.05961f
C1512 bgr_0.1st_Vout_1.n4 GNDA 1.04144f
C1513 bgr_0.1st_Vout_1.t11 GNDA 0.418685f
C1514 bgr_0.1st_Vout_1.t15 GNDA 0.411673f
C1515 bgr_0.1st_Vout_1.t29 GNDA 0.418685f
C1516 bgr_0.1st_Vout_1.t35 GNDA 0.411673f
C1517 bgr_0.1st_Vout_1.t31 GNDA 0.418685f
C1518 bgr_0.1st_Vout_1.t34 GNDA 0.411673f
C1519 bgr_0.1st_Vout_1.t20 GNDA 0.418685f
C1520 bgr_0.1st_Vout_1.t28 GNDA 0.411673f
C1521 bgr_0.1st_Vout_1.t24 GNDA 0.418685f
C1522 bgr_0.1st_Vout_1.t27 GNDA 0.411673f
C1523 bgr_0.1st_Vout_1.t14 GNDA 0.418685f
C1524 bgr_0.1st_Vout_1.t19 GNDA 0.411673f
C1525 bgr_0.1st_Vout_1.t30 GNDA 0.418685f
C1526 bgr_0.1st_Vout_1.t33 GNDA 0.411673f
C1527 bgr_0.1st_Vout_1.t18 GNDA 0.418685f
C1528 bgr_0.1st_Vout_1.t26 GNDA 0.411673f
C1529 bgr_0.1st_Vout_1.t23 GNDA 0.418685f
C1530 bgr_0.1st_Vout_1.t25 GNDA 0.411673f
C1531 bgr_0.1st_Vout_1.t17 GNDA 0.411673f
C1532 bgr_0.1st_Vout_1.t12 GNDA 0.411673f
C1533 bgr_0.1st_Vout_1.t21 GNDA 0.026894f
C1534 bgr_0.1st_Vout_1.n5 GNDA 0.835652f
C1535 bgr_0.1st_Vout_1.t0 GNDA 0.010292f
C1536 bgr_0.1st_Vout_1.t3 GNDA 0.010292f
C1537 bgr_0.1st_Vout_1.n6 GNDA 0.025944f
C1538 bgr_0.1st_Vout_1.n7 GNDA 0.122259f
C1539 bgr_0.1st_Vout_1.t36 GNDA 0.015678f
C1540 bgr_0.1st_Vout_1.t16 GNDA 0.015678f
C1541 bgr_0.1st_Vout_1.n8 GNDA 0.034878f
C1542 bgr_0.1st_Vout_1.n9 GNDA 0.096376f
C1543 bgr_0.1st_Vout_1.t8 GNDA 0.021677f
C1544 bgr_0.1st_Vout_1.n10 GNDA 0.014867f
C1545 bgr_0.1st_Vout_1.n11 GNDA 0.224869f
C1546 bgr_0.1st_Vout_1.n12 GNDA 0.013451f
C1547 bgr_0.1st_Vout_1.n13 GNDA 0.057048f
C1548 bgr_0.1st_Vout_1.t5 GNDA 0.010292f
C1549 bgr_0.1st_Vout_1.t1 GNDA 0.010292f
C1550 bgr_0.1st_Vout_1.n14 GNDA 0.024868f
C1551 bgr_0.1st_Vout_1.n15 GNDA 0.091944f
C1552 bgr_0.1st_Vout_1.n16 GNDA 0.045284f
C1553 bgr_0.1st_Vout_1.t32 GNDA 0.015678f
C1554 bgr_0.1st_Vout_1.t22 GNDA 0.015678f
C1555 bgr_0.1st_Vout_1.n17 GNDA 0.034878f
C1556 bgr_0.1st_Vout_1.n18 GNDA 0.096376f
C1557 bgr_0.1st_Vout_1.t4 GNDA 0.010292f
C1558 bgr_0.1st_Vout_1.t2 GNDA 0.010292f
C1559 bgr_0.1st_Vout_1.n19 GNDA 0.025944f
C1560 bgr_0.1st_Vout_1.n20 GNDA 0.122259f
C1561 bgr_0.1st_Vout_1.t13 GNDA 0.024608f
C1562 bgr_0.V_mir1.t9 GNDA 0.03537f
C1563 bgr_0.V_mir1.t2 GNDA 0.053881f
C1564 bgr_0.V_mir1.t6 GNDA 0.042444f
C1565 bgr_0.V_mir1.t18 GNDA 0.042444f
C1566 bgr_0.V_mir1.t20 GNDA 0.06851f
C1567 bgr_0.V_mir1.n0 GNDA 0.076506f
C1568 bgr_0.V_mir1.n1 GNDA 0.052264f
C1569 bgr_0.V_mir1.n2 GNDA 0.081315f
C1570 bgr_0.V_mir1.t3 GNDA 0.03537f
C1571 bgr_0.V_mir1.t7 GNDA 0.03537f
C1572 bgr_0.V_mir1.n3 GNDA 0.08097f
C1573 bgr_0.V_mir1.n4 GNDA 0.201563f
C1574 bgr_0.V_mir1.t16 GNDA 0.017685f
C1575 bgr_0.V_mir1.t1 GNDA 0.017685f
C1576 bgr_0.V_mir1.n5 GNDA 0.046242f
C1577 bgr_0.V_mir1.t14 GNDA 0.075466f
C1578 bgr_0.V_mir1.t0 GNDA 0.017685f
C1579 bgr_0.V_mir1.t15 GNDA 0.017685f
C1580 bgr_0.V_mir1.n6 GNDA 0.050199f
C1581 bgr_0.V_mir1.n7 GNDA 0.827814f
C1582 bgr_0.V_mir1.n8 GNDA 0.268286f
C1583 bgr_0.V_mir1.t4 GNDA 0.053881f
C1584 bgr_0.V_mir1.t10 GNDA 0.042444f
C1585 bgr_0.V_mir1.t17 GNDA 0.042444f
C1586 bgr_0.V_mir1.t21 GNDA 0.06851f
C1587 bgr_0.V_mir1.n9 GNDA 0.076506f
C1588 bgr_0.V_mir1.n10 GNDA 0.052264f
C1589 bgr_0.V_mir1.n11 GNDA 0.081315f
C1590 bgr_0.V_mir1.t5 GNDA 0.03537f
C1591 bgr_0.V_mir1.t11 GNDA 0.03537f
C1592 bgr_0.V_mir1.n12 GNDA 0.08097f
C1593 bgr_0.V_mir1.n13 GNDA 0.156007f
C1594 bgr_0.V_mir1.n14 GNDA 0.09373f
C1595 bgr_0.V_mir1.n15 GNDA 0.699157f
C1596 bgr_0.V_mir1.t8 GNDA 0.053881f
C1597 bgr_0.V_mir1.t12 GNDA 0.042444f
C1598 bgr_0.V_mir1.t22 GNDA 0.042444f
C1599 bgr_0.V_mir1.t19 GNDA 0.06851f
C1600 bgr_0.V_mir1.n16 GNDA 0.076506f
C1601 bgr_0.V_mir1.n17 GNDA 0.052264f
C1602 bgr_0.V_mir1.n18 GNDA 0.081315f
C1603 bgr_0.V_mir1.n19 GNDA 0.203577f
C1604 bgr_0.V_mir1.n20 GNDA 0.08097f
C1605 bgr_0.V_mir1.t13 GNDA 0.03537f
C1606 bgr_0.Vin+.t1 GNDA 0.173951f
C1607 bgr_0.Vin+.t7 GNDA 0.010696f
C1608 bgr_0.Vin+.t8 GNDA 0.025367f
C1609 bgr_0.Vin+.t9 GNDA 0.01649f
C1610 bgr_0.Vin+.n0 GNDA 0.054406f
C1611 bgr_0.Vin+.t6 GNDA 0.01649f
C1612 bgr_0.Vin+.n1 GNDA 0.042338f
C1613 bgr_0.Vin+.t10 GNDA 0.01649f
C1614 bgr_0.Vin+.n2 GNDA 0.042909f
C1615 bgr_0.Vin+.n3 GNDA 0.130793f
C1616 bgr_0.Vin+.t4 GNDA 0.05348f
C1617 bgr_0.Vin+.t3 GNDA 0.05348f
C1618 bgr_0.Vin+.n4 GNDA 0.176679f
C1619 bgr_0.Vin+.n5 GNDA 1.27851f
C1620 bgr_0.Vin+.t2 GNDA 0.05348f
C1621 bgr_0.Vin+.t5 GNDA 0.05348f
C1622 bgr_0.Vin+.n6 GNDA 0.176679f
C1623 bgr_0.Vin+.n7 GNDA 1.06525f
C1624 bgr_0.Vin+.n8 GNDA 1.7265f
C1625 bgr_0.Vin+.t0 GNDA 0.232527f
C1626 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 GNDA 0.016041f
C1627 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 GNDA 0.016041f
C1628 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 GNDA 0.040225f
C1629 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 GNDA 0.016041f
C1630 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 GNDA 0.016041f
C1631 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 GNDA 0.040013f
C1632 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 GNDA 0.355706f
C1633 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 GNDA 0.016041f
C1634 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 GNDA 0.016041f
C1635 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 GNDA 0.032081f
C1636 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 GNDA 0.059636f
C1637 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 GNDA 0.205433f
C1638 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 GNDA 0.032081f
C1639 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 GNDA 0.032081f
C1640 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 GNDA 0.094125f
C1641 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 GNDA 0.032081f
C1642 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 GNDA 0.032081f
C1643 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 GNDA 0.093697f
C1644 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 GNDA 0.323873f
C1645 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 GNDA 0.032081f
C1646 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 GNDA 0.032081f
C1647 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 GNDA 0.093697f
C1648 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 GNDA 0.167764f
C1649 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 GNDA 0.032081f
C1650 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 GNDA 0.032081f
C1651 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 GNDA 0.093697f
C1652 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 GNDA 0.167764f
C1653 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 GNDA 0.032081f
C1654 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 GNDA 0.032081f
C1655 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 GNDA 0.093697f
C1656 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 GNDA 0.245609f
C1657 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 GNDA 1.4546f
C1658 bgr_0.V_CMFB_S3 GNDA 0.92132f
C1659 two_stage_opamp_dummy_magic_0.Y.t9 GNDA 0.023873f
C1660 two_stage_opamp_dummy_magic_0.Y.t22 GNDA 0.023873f
C1661 two_stage_opamp_dummy_magic_0.Y.n0 GNDA 0.080602f
C1662 two_stage_opamp_dummy_magic_0.Y.t18 GNDA 0.023873f
C1663 two_stage_opamp_dummy_magic_0.Y.t7 GNDA 0.023873f
C1664 two_stage_opamp_dummy_magic_0.Y.n1 GNDA 0.086146f
C1665 two_stage_opamp_dummy_magic_0.Y.t4 GNDA 0.023873f
C1666 two_stage_opamp_dummy_magic_0.Y.t3 GNDA 0.023873f
C1667 two_stage_opamp_dummy_magic_0.Y.n2 GNDA 0.085394f
C1668 two_stage_opamp_dummy_magic_0.Y.n3 GNDA 0.317069f
C1669 two_stage_opamp_dummy_magic_0.Y.t24 GNDA 0.023873f
C1670 two_stage_opamp_dummy_magic_0.Y.t6 GNDA 0.023873f
C1671 two_stage_opamp_dummy_magic_0.Y.n4 GNDA 0.085394f
C1672 two_stage_opamp_dummy_magic_0.Y.n5 GNDA 0.164481f
C1673 two_stage_opamp_dummy_magic_0.Y.t5 GNDA 0.023873f
C1674 two_stage_opamp_dummy_magic_0.Y.t15 GNDA 0.023873f
C1675 two_stage_opamp_dummy_magic_0.Y.n6 GNDA 0.085394f
C1676 two_stage_opamp_dummy_magic_0.Y.n7 GNDA 0.164481f
C1677 two_stage_opamp_dummy_magic_0.Y.t14 GNDA 0.023873f
C1678 two_stage_opamp_dummy_magic_0.Y.t19 GNDA 0.023873f
C1679 two_stage_opamp_dummy_magic_0.Y.n8 GNDA 0.086146f
C1680 two_stage_opamp_dummy_magic_0.Y.n9 GNDA 0.200335f
C1681 two_stage_opamp_dummy_magic_0.Y.n10 GNDA 0.250257f
C1682 two_stage_opamp_dummy_magic_0.Y.t17 GNDA 0.055705f
C1683 two_stage_opamp_dummy_magic_0.Y.t16 GNDA 0.055705f
C1684 two_stage_opamp_dummy_magic_0.Y.n11 GNDA 0.193729f
C1685 two_stage_opamp_dummy_magic_0.Y.t2 GNDA 0.055705f
C1686 two_stage_opamp_dummy_magic_0.Y.t0 GNDA 0.055705f
C1687 two_stage_opamp_dummy_magic_0.Y.n12 GNDA 0.193042f
C1688 two_stage_opamp_dummy_magic_0.Y.n13 GNDA 0.364444f
C1689 two_stage_opamp_dummy_magic_0.Y.t13 GNDA 0.055705f
C1690 two_stage_opamp_dummy_magic_0.Y.t23 GNDA 0.055705f
C1691 two_stage_opamp_dummy_magic_0.Y.n14 GNDA 0.193042f
C1692 two_stage_opamp_dummy_magic_0.Y.n15 GNDA 0.188932f
C1693 two_stage_opamp_dummy_magic_0.Y.t10 GNDA 0.055705f
C1694 two_stage_opamp_dummy_magic_0.Y.t12 GNDA 0.055705f
C1695 two_stage_opamp_dummy_magic_0.Y.n16 GNDA 0.193042f
C1696 two_stage_opamp_dummy_magic_0.Y.n17 GNDA 0.188932f
C1697 two_stage_opamp_dummy_magic_0.Y.t11 GNDA 0.055705f
C1698 two_stage_opamp_dummy_magic_0.Y.t20 GNDA 0.055705f
C1699 two_stage_opamp_dummy_magic_0.Y.n18 GNDA 0.193042f
C1700 two_stage_opamp_dummy_magic_0.Y.n19 GNDA 0.222471f
C1701 two_stage_opamp_dummy_magic_0.Y.t21 GNDA 0.055705f
C1702 two_stage_opamp_dummy_magic_0.Y.t8 GNDA 0.055705f
C1703 two_stage_opamp_dummy_magic_0.Y.n20 GNDA 0.189043f
C1704 two_stage_opamp_dummy_magic_0.Y.n21 GNDA 0.376251f
C1705 two_stage_opamp_dummy_magic_0.Y.t52 GNDA 0.033423f
C1706 two_stage_opamp_dummy_magic_0.Y.t38 GNDA 0.040585f
C1707 two_stage_opamp_dummy_magic_0.Y.n22 GNDA 0.037846f
C1708 two_stage_opamp_dummy_magic_0.Y.t42 GNDA 0.033423f
C1709 two_stage_opamp_dummy_magic_0.Y.t25 GNDA 0.033423f
C1710 two_stage_opamp_dummy_magic_0.Y.t30 GNDA 0.033423f
C1711 two_stage_opamp_dummy_magic_0.Y.t47 GNDA 0.033423f
C1712 two_stage_opamp_dummy_magic_0.Y.t33 GNDA 0.033423f
C1713 two_stage_opamp_dummy_magic_0.Y.t49 GNDA 0.033423f
C1714 two_stage_opamp_dummy_magic_0.Y.t37 GNDA 0.033423f
C1715 two_stage_opamp_dummy_magic_0.Y.t29 GNDA 0.040585f
C1716 two_stage_opamp_dummy_magic_0.Y.n23 GNDA 0.040585f
C1717 two_stage_opamp_dummy_magic_0.Y.n24 GNDA 0.026261f
C1718 two_stage_opamp_dummy_magic_0.Y.n25 GNDA 0.026261f
C1719 two_stage_opamp_dummy_magic_0.Y.n26 GNDA 0.026261f
C1720 two_stage_opamp_dummy_magic_0.Y.n27 GNDA 0.026261f
C1721 two_stage_opamp_dummy_magic_0.Y.n28 GNDA 0.026261f
C1722 two_stage_opamp_dummy_magic_0.Y.n29 GNDA 0.023522f
C1723 two_stage_opamp_dummy_magic_0.Y.n30 GNDA 0.023134f
C1724 two_stage_opamp_dummy_magic_0.Y.t27 GNDA 0.051328f
C1725 two_stage_opamp_dummy_magic_0.Y.t45 GNDA 0.058351f
C1726 two_stage_opamp_dummy_magic_0.Y.n31 GNDA 0.049922f
C1727 two_stage_opamp_dummy_magic_0.Y.t46 GNDA 0.051328f
C1728 two_stage_opamp_dummy_magic_0.Y.t28 GNDA 0.051328f
C1729 two_stage_opamp_dummy_magic_0.Y.t36 GNDA 0.051328f
C1730 two_stage_opamp_dummy_magic_0.Y.t51 GNDA 0.051328f
C1731 two_stage_opamp_dummy_magic_0.Y.t41 GNDA 0.051328f
C1732 two_stage_opamp_dummy_magic_0.Y.t54 GNDA 0.051328f
C1733 two_stage_opamp_dummy_magic_0.Y.t44 GNDA 0.051328f
C1734 two_stage_opamp_dummy_magic_0.Y.t34 GNDA 0.058351f
C1735 two_stage_opamp_dummy_magic_0.Y.n32 GNDA 0.05266f
C1736 two_stage_opamp_dummy_magic_0.Y.n33 GNDA 0.032229f
C1737 two_stage_opamp_dummy_magic_0.Y.n34 GNDA 0.032229f
C1738 two_stage_opamp_dummy_magic_0.Y.n35 GNDA 0.032229f
C1739 two_stage_opamp_dummy_magic_0.Y.n36 GNDA 0.032229f
C1740 two_stage_opamp_dummy_magic_0.Y.n37 GNDA 0.032229f
C1741 two_stage_opamp_dummy_magic_0.Y.n38 GNDA 0.02949f
C1742 two_stage_opamp_dummy_magic_0.Y.n39 GNDA 0.023086f
C1743 two_stage_opamp_dummy_magic_0.Y.n40 GNDA 0.249706f
C1744 two_stage_opamp_dummy_magic_0.Y.n41 GNDA 0.51804f
C1745 two_stage_opamp_dummy_magic_0.Y.n42 GNDA 0.261996f
C1746 two_stage_opamp_dummy_magic_0.Y.t35 GNDA 0.105043f
C1747 two_stage_opamp_dummy_magic_0.Y.t48 GNDA 0.105043f
C1748 two_stage_opamp_dummy_magic_0.Y.t32 GNDA 0.105043f
C1749 two_stage_opamp_dummy_magic_0.Y.t26 GNDA 0.105043f
C1750 two_stage_opamp_dummy_magic_0.Y.t43 GNDA 0.105043f
C1751 two_stage_opamp_dummy_magic_0.Y.t53 GNDA 0.105043f
C1752 two_stage_opamp_dummy_magic_0.Y.t40 GNDA 0.111878f
C1753 two_stage_opamp_dummy_magic_0.Y.n43 GNDA 0.088659f
C1754 two_stage_opamp_dummy_magic_0.Y.n44 GNDA 0.050134f
C1755 two_stage_opamp_dummy_magic_0.Y.n45 GNDA 0.050134f
C1756 two_stage_opamp_dummy_magic_0.Y.n46 GNDA 0.050134f
C1757 two_stage_opamp_dummy_magic_0.Y.n47 GNDA 0.050134f
C1758 two_stage_opamp_dummy_magic_0.Y.n48 GNDA 0.047395f
C1759 two_stage_opamp_dummy_magic_0.Y.t50 GNDA 0.105043f
C1760 two_stage_opamp_dummy_magic_0.Y.t39 GNDA 0.105043f
C1761 two_stage_opamp_dummy_magic_0.Y.t31 GNDA 0.111878f
C1762 two_stage_opamp_dummy_magic_0.Y.n49 GNDA 0.088659f
C1763 two_stage_opamp_dummy_magic_0.Y.n50 GNDA 0.047395f
C1764 two_stage_opamp_dummy_magic_0.Y.n51 GNDA 0.025681f
C1765 two_stage_opamp_dummy_magic_0.Y.n52 GNDA 0.925108f
C1766 two_stage_opamp_dummy_magic_0.Y.t1 GNDA 0.777549f
C1767 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 GNDA 0.034707f
C1768 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 GNDA 0.010902f
C1769 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 GNDA 0.020344f
C1770 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 GNDA 0.04857f
C1771 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 GNDA 0.303701f
C1772 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 GNDA 0.010902f
C1773 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 GNDA 0.020344f
C1774 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 GNDA 0.04857f
C1775 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 GNDA 0.280548f
C1776 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 GNDA 0.034375f
C1777 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 GNDA 0.273171f
C1778 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 GNDA 0.010902f
C1779 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 GNDA 0.020344f
C1780 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 GNDA 0.04857f
C1781 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 GNDA 0.16963f
C1782 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 GNDA 0.010902f
C1783 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 GNDA 0.020344f
C1784 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 GNDA 0.04857f
C1785 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 GNDA 0.215581f
C1786 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 GNDA 0.380652f
C1787 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 GNDA 0.059389f
C1788 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 GNDA 0.022208f
C1789 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 GNDA 0.069655f
C1790 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 GNDA 0.022208f
C1791 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 GNDA 0.05702f
C1792 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 GNDA 0.022208f
C1793 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 GNDA 0.05702f
C1794 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 GNDA 0.022208f
C1795 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 GNDA 0.099349f
C1796 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 GNDA 1.98565f
C1797 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 GNDA 0.072025f
C1798 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 GNDA 0.072025f
C1799 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 GNDA 0.253667f
C1800 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 GNDA 0.072025f
C1801 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 GNDA 0.072025f
C1802 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 GNDA 0.241356f
C1803 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 GNDA 1.12793f
C1804 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 GNDA 0.072025f
C1805 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 GNDA 0.072025f
C1806 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 GNDA 0.241356f
C1807 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 GNDA 0.806559f
C1808 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 GNDA 1.65703f
C1809 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 GNDA 0.343499f
C1810 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 GNDA 0.344645f
C1811 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 GNDA 0.185116f
C1812 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 GNDA 0.197667f
C1813 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 GNDA 0.343499f
C1814 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 GNDA 0.344645f
C1815 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 GNDA 0.185116f
C1816 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 GNDA 0.216163f
C1817 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 GNDA 0.343499f
C1818 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 GNDA 0.344645f
C1819 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 GNDA 0.185116f
C1820 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 GNDA 0.216163f
C1821 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 GNDA 0.343499f
C1822 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 GNDA 0.344645f
C1823 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 GNDA 0.185116f
C1824 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 GNDA 0.216163f
C1825 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 GNDA 0.343499f
C1826 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 GNDA 0.344645f
C1827 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 GNDA 0.363141f
C1828 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 GNDA 0.363141f
C1829 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 GNDA 0.185116f
C1830 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 GNDA 0.216163f
C1831 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 GNDA 0.343499f
C1832 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 GNDA 0.344645f
C1833 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 GNDA 0.363141f
C1834 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 GNDA 0.363141f
C1835 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 GNDA 0.185116f
C1836 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 GNDA 0.216163f
C1837 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 GNDA 0.344645f
C1838 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 GNDA 0.345894f
C1839 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 GNDA 0.344645f
C1840 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 GNDA 0.347347f
C1841 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 GNDA 0.377789f
C1842 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 GNDA 0.344645f
C1843 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 GNDA 0.345894f
C1844 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 GNDA 0.344645f
C1845 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 GNDA 0.345894f
C1846 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 GNDA 0.344645f
C1847 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 GNDA 0.345894f
C1848 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 GNDA 0.344645f
C1849 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 GNDA 0.345894f
C1850 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 GNDA 0.344645f
C1851 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 GNDA 0.345894f
C1852 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 GNDA 0.344645f
C1853 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 GNDA 0.345894f
C1854 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 GNDA 0.344645f
C1855 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 GNDA 0.345894f
C1856 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 GNDA 0.344645f
C1857 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 GNDA 0.345894f
C1858 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 GNDA 0.344645f
C1859 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 GNDA 0.345894f
C1860 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 GNDA 0.344645f
C1861 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 GNDA 0.345894f
C1862 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 GNDA 0.344645f
C1863 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 GNDA 0.345894f
C1864 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 GNDA 0.344645f
C1865 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 GNDA 0.345894f
C1866 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 GNDA 0.344645f
C1867 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 GNDA 0.345894f
C1868 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 GNDA 0.344645f
C1869 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 GNDA 0.345894f
C1870 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 GNDA 0.344645f
C1871 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 GNDA 0.345894f
C1872 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 GNDA 0.344645f
C1873 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 GNDA 0.345894f
C1874 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 GNDA 0.344645f
C1875 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 GNDA 0.345894f
C1876 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 GNDA 0.344645f
C1877 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 GNDA 0.345894f
C1878 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 GNDA 0.344645f
C1879 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 GNDA 0.345894f
C1880 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 GNDA 0.344645f
C1881 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 GNDA 0.345894f
C1882 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 GNDA 0.344645f
C1883 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 GNDA 0.345894f
C1884 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 GNDA 0.344645f
C1885 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 GNDA 0.345894f
C1886 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 GNDA 0.344645f
C1887 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 GNDA 0.345894f
C1888 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 GNDA 0.344645f
C1889 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 GNDA 0.345894f
C1890 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 GNDA 0.344645f
C1891 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 GNDA 0.345894f
C1892 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 GNDA 0.344645f
C1893 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 GNDA 0.345894f
C1894 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 GNDA 0.344645f
C1895 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 GNDA 0.345894f
C1896 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 GNDA 0.344645f
C1897 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 GNDA 0.345894f
C1898 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 GNDA 0.344645f
C1899 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 GNDA 0.361543f
C1900 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 GNDA 0.344645f
C1901 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 GNDA 0.185116f
C1902 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 GNDA 0.19812f
C1903 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 GNDA 0.344645f
C1904 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 GNDA 0.185116f
C1905 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 GNDA 0.196521f
C1906 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 GNDA 0.344645f
C1907 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 GNDA 0.185116f
C1908 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 GNDA 0.196521f
C1909 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 GNDA 0.344645f
C1910 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 GNDA 0.185116f
C1911 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 GNDA 0.196521f
C1912 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 GNDA 0.344645f
C1913 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 GNDA 0.185116f
C1914 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 GNDA 0.196521f
C1915 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 GNDA 0.344645f
C1916 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 GNDA 0.185116f
C1917 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 GNDA 0.196521f
C1918 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 GNDA 0.344645f
C1919 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 GNDA 0.185116f
C1920 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 GNDA 0.196521f
C1921 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 GNDA 0.344645f
C1922 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 GNDA 0.185116f
C1923 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 GNDA 0.196521f
C1924 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 GNDA 0.344645f
C1925 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 GNDA 0.185116f
C1926 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 GNDA 0.196521f
C1927 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 GNDA 0.344645f
C1928 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 GNDA 0.345894f
C1929 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 GNDA 0.344645f
C1930 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 GNDA 0.345894f
C1931 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 GNDA 0.166619f
C1932 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 GNDA 0.214914f
C1933 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 GNDA 0.18397f
C1934 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 GNDA 0.23341f
C1935 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 GNDA 0.18397f
C1936 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 GNDA 0.250658f
C1937 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 GNDA 0.18397f
C1938 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 GNDA 0.250658f
C1939 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 GNDA 0.18397f
C1940 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 GNDA 0.250658f
C1941 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 GNDA 0.18397f
C1942 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 GNDA 0.250658f
C1943 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 GNDA 0.18397f
C1944 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 GNDA 0.250658f
C1945 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 GNDA 0.18397f
C1946 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 GNDA 0.250658f
C1947 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 GNDA 0.18397f
C1948 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 GNDA 0.250658f
C1949 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 GNDA 0.18397f
C1950 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 GNDA 0.250658f
C1951 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 GNDA 0.18397f
C1952 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 GNDA 0.250658f
C1953 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 GNDA 0.18397f
C1954 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 GNDA 0.250658f
C1955 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 GNDA 0.18397f
C1956 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 GNDA 0.250658f
C1957 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 GNDA 0.18397f
C1958 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 GNDA 0.250658f
C1959 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 GNDA 0.18397f
C1960 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 GNDA 0.250658f
C1961 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 GNDA 0.18397f
C1962 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 GNDA 0.250658f
C1963 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 GNDA 0.18397f
C1964 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 GNDA 0.23341f
C1965 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 GNDA 0.343499f
C1966 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 GNDA 0.166619f
C1967 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 GNDA 0.216163f
C1968 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 GNDA 0.343499f
C1969 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 GNDA 0.166619f
C1970 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 GNDA 0.216163f
C1971 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 GNDA 0.343499f
C1972 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 GNDA 0.344645f
C1973 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 GNDA 0.363141f
C1974 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 GNDA 0.363141f
C1975 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 GNDA 0.185116f
C1976 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 GNDA 0.216163f
C1977 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 GNDA 0.343499f
C1978 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 GNDA 0.216163f
C1979 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 GNDA 0.185116f
C1980 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 GNDA 0.363141f
C1981 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 GNDA 0.363141f
C1982 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 GNDA 0.434494f
C1983 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 GNDA 0.297192f
C1984 VOUT-.t13 GNDA 0.050898f
C1985 VOUT-.t3 GNDA 0.050898f
C1986 VOUT-.n0 GNDA 0.235456f
C1987 VOUT-.t11 GNDA 0.050898f
C1988 VOUT-.t16 GNDA 0.050898f
C1989 VOUT-.n1 GNDA 0.234668f
C1990 VOUT-.n2 GNDA 0.145013f
C1991 VOUT-.t17 GNDA 0.050898f
C1992 VOUT-.t12 GNDA 0.050898f
C1993 VOUT-.n3 GNDA 0.234668f
C1994 VOUT-.n4 GNDA 0.090715f
C1995 VOUT-.t18 GNDA 0.084152f
C1996 VOUT-.n5 GNDA 0.120712f
C1997 VOUT-.t14 GNDA 0.043627f
C1998 VOUT-.t6 GNDA 0.043627f
C1999 VOUT-.n6 GNDA 0.175348f
C2000 VOUT-.t8 GNDA 0.043627f
C2001 VOUT-.t15 GNDA 0.043627f
C2002 VOUT-.n7 GNDA 0.175348f
C2003 VOUT-.t1 GNDA 0.043627f
C2004 VOUT-.t10 GNDA 0.043627f
C2005 VOUT-.n8 GNDA 0.175025f
C2006 VOUT-.n9 GNDA 0.172421f
C2007 VOUT-.t7 GNDA 0.043627f
C2008 VOUT-.t0 GNDA 0.043627f
C2009 VOUT-.n10 GNDA 0.175025f
C2010 VOUT-.n11 GNDA 0.088916f
C2011 VOUT-.t5 GNDA 0.043627f
C2012 VOUT-.t4 GNDA 0.043627f
C2013 VOUT-.n12 GNDA 0.175025f
C2014 VOUT-.n13 GNDA 0.088916f
C2015 VOUT-.n14 GNDA 0.105317f
C2016 VOUT-.t2 GNDA 0.043627f
C2017 VOUT-.t9 GNDA 0.043627f
C2018 VOUT-.n15 GNDA 0.172883f
C2019 VOUT-.n16 GNDA 0.213802f
C2020 VOUT-.t101 GNDA 0.290845f
C2021 VOUT-.t108 GNDA 0.295799f
C2022 VOUT-.t149 GNDA 0.290845f
C2023 VOUT-.n17 GNDA 0.195002f
C2024 VOUT-.n18 GNDA 0.127245f
C2025 VOUT-.t48 GNDA 0.295178f
C2026 VOUT-.t92 GNDA 0.295178f
C2027 VOUT-.t42 GNDA 0.295178f
C2028 VOUT-.t130 GNDA 0.295178f
C2029 VOUT-.t84 GNDA 0.295178f
C2030 VOUT-.t125 GNDA 0.295178f
C2031 VOUT-.t74 GNDA 0.295178f
C2032 VOUT-.t23 GNDA 0.295178f
C2033 VOUT-.t64 GNDA 0.295178f
C2034 VOUT-.t150 GNDA 0.295178f
C2035 VOUT-.t88 GNDA 0.290845f
C2036 VOUT-.n19 GNDA 0.195622f
C2037 VOUT-.t51 GNDA 0.290845f
C2038 VOUT-.n20 GNDA 0.250156f
C2039 VOUT-.t137 GNDA 0.290845f
C2040 VOUT-.n21 GNDA 0.250156f
C2041 VOUT-.t106 GNDA 0.290845f
C2042 VOUT-.n22 GNDA 0.250156f
C2043 VOUT-.t75 GNDA 0.290845f
C2044 VOUT-.n23 GNDA 0.250156f
C2045 VOUT-.t25 GNDA 0.290845f
C2046 VOUT-.n24 GNDA 0.250156f
C2047 VOUT-.t128 GNDA 0.290845f
C2048 VOUT-.n25 GNDA 0.250156f
C2049 VOUT-.t90 GNDA 0.290845f
C2050 VOUT-.n26 GNDA 0.250156f
C2051 VOUT-.t54 GNDA 0.290845f
C2052 VOUT-.n27 GNDA 0.250156f
C2053 VOUT-.t140 GNDA 0.290845f
C2054 VOUT-.n28 GNDA 0.250156f
C2055 VOUT-.t110 GNDA 0.290845f
C2056 VOUT-.t28 GNDA 0.295799f
C2057 VOUT-.t79 GNDA 0.290845f
C2058 VOUT-.n29 GNDA 0.195002f
C2059 VOUT-.n30 GNDA 0.236312f
C2060 VOUT-.t24 GNDA 0.295799f
C2061 VOUT-.t113 GNDA 0.290845f
C2062 VOUT-.n31 GNDA 0.195002f
C2063 VOUT-.t78 GNDA 0.290845f
C2064 VOUT-.t129 GNDA 0.295799f
C2065 VOUT-.t38 GNDA 0.290845f
C2066 VOUT-.n32 GNDA 0.195002f
C2067 VOUT-.n33 GNDA 0.236312f
C2068 VOUT-.t61 GNDA 0.295799f
C2069 VOUT-.t147 GNDA 0.290845f
C2070 VOUT-.n34 GNDA 0.195002f
C2071 VOUT-.t117 GNDA 0.290845f
C2072 VOUT-.t32 GNDA 0.295799f
C2073 VOUT-.t83 GNDA 0.290845f
C2074 VOUT-.n35 GNDA 0.195002f
C2075 VOUT-.n36 GNDA 0.236312f
C2076 VOUT-.t100 GNDA 0.295799f
C2077 VOUT-.t47 GNDA 0.290845f
C2078 VOUT-.n37 GNDA 0.195002f
C2079 VOUT-.t153 GNDA 0.290845f
C2080 VOUT-.t71 GNDA 0.295799f
C2081 VOUT-.t123 GNDA 0.290845f
C2082 VOUT-.n38 GNDA 0.195002f
C2083 VOUT-.n39 GNDA 0.236312f
C2084 VOUT-.t69 GNDA 0.295799f
C2085 VOUT-.t154 GNDA 0.290845f
C2086 VOUT-.n40 GNDA 0.195002f
C2087 VOUT-.t124 GNDA 0.290845f
C2088 VOUT-.t35 GNDA 0.295799f
C2089 VOUT-.t86 GNDA 0.290845f
C2090 VOUT-.n41 GNDA 0.195002f
C2091 VOUT-.n42 GNDA 0.236312f
C2092 VOUT-.t96 GNDA 0.290845f
C2093 VOUT-.t85 GNDA 0.295799f
C2094 VOUT-.t57 GNDA 0.290845f
C2095 VOUT-.n43 GNDA 0.195002f
C2096 VOUT-.n44 GNDA 0.127245f
C2097 VOUT-.t132 GNDA 0.295178f
C2098 VOUT-.t115 GNDA 0.295178f
C2099 VOUT-.t131 GNDA 0.295799f
C2100 VOUT-.t104 GNDA 0.290845f
C2101 VOUT-.n45 GNDA 0.195002f
C2102 VOUT-.t73 GNDA 0.290845f
C2103 VOUT-.n46 GNDA 0.1227f
C2104 VOUT-.t146 GNDA 0.295178f
C2105 VOUT-.t31 GNDA 0.295799f
C2106 VOUT-.t138 GNDA 0.290845f
C2107 VOUT-.n47 GNDA 0.195002f
C2108 VOUT-.t107 GNDA 0.290845f
C2109 VOUT-.n48 GNDA 0.1227f
C2110 VOUT-.t46 GNDA 0.295178f
C2111 VOUT-.t62 GNDA 0.295799f
C2112 VOUT-.t41 GNDA 0.290845f
C2113 VOUT-.n49 GNDA 0.195002f
C2114 VOUT-.t143 GNDA 0.290845f
C2115 VOUT-.n50 GNDA 0.1227f
C2116 VOUT-.t87 GNDA 0.295178f
C2117 VOUT-.t114 GNDA 0.295799f
C2118 VOUT-.t21 GNDA 0.290845f
C2119 VOUT-.n51 GNDA 0.195002f
C2120 VOUT-.t126 GNDA 0.290845f
C2121 VOUT-.n52 GNDA 0.1227f
C2122 VOUT-.t65 GNDA 0.295178f
C2123 VOUT-.t26 GNDA 0.295422f
C2124 VOUT-.t102 GNDA 0.295178f
C2125 VOUT-.t59 GNDA 0.295422f
C2126 VOUT-.t134 GNDA 0.295178f
C2127 VOUT-.t37 GNDA 0.295422f
C2128 VOUT-.t120 GNDA 0.295178f
C2129 VOUT-.t81 GNDA 0.295422f
C2130 VOUT-.t155 GNDA 0.295178f
C2131 VOUT-.t119 GNDA 0.290845f
C2132 VOUT-.n53 GNDA 0.321926f
C2133 VOUT-.t82 GNDA 0.290845f
C2134 VOUT-.n54 GNDA 0.376459f
C2135 VOUT-.t97 GNDA 0.290845f
C2136 VOUT-.n55 GNDA 0.376459f
C2137 VOUT-.t63 GNDA 0.290845f
C2138 VOUT-.n56 GNDA 0.376459f
C2139 VOUT-.t27 GNDA 0.290845f
C2140 VOUT-.n57 GNDA 0.309234f
C2141 VOUT-.t45 GNDA 0.290845f
C2142 VOUT-.n58 GNDA 0.309234f
C2143 VOUT-.t144 GNDA 0.290845f
C2144 VOUT-.n59 GNDA 0.309234f
C2145 VOUT-.t112 GNDA 0.290845f
C2146 VOUT-.n60 GNDA 0.309234f
C2147 VOUT-.t76 GNDA 0.290845f
C2148 VOUT-.n61 GNDA 0.250156f
C2149 VOUT-.t93 GNDA 0.290845f
C2150 VOUT-.n62 GNDA 0.250156f
C2151 VOUT-.t56 GNDA 0.290845f
C2152 VOUT-.t40 GNDA 0.295799f
C2153 VOUT-.t19 GNDA 0.290845f
C2154 VOUT-.n63 GNDA 0.195002f
C2155 VOUT-.n64 GNDA 0.236312f
C2156 VOUT-.t34 GNDA 0.295799f
C2157 VOUT-.t52 GNDA 0.290845f
C2158 VOUT-.n65 GNDA 0.195002f
C2159 VOUT-.t156 GNDA 0.290845f
C2160 VOUT-.t136 GNDA 0.295799f
C2161 VOUT-.t121 GNDA 0.290845f
C2162 VOUT-.n66 GNDA 0.195002f
C2163 VOUT-.n67 GNDA 0.236312f
C2164 VOUT-.t70 GNDA 0.295799f
C2165 VOUT-.t89 GNDA 0.290845f
C2166 VOUT-.n68 GNDA 0.195002f
C2167 VOUT-.t50 GNDA 0.290845f
C2168 VOUT-.t36 GNDA 0.295799f
C2169 VOUT-.t151 GNDA 0.290845f
C2170 VOUT-.n69 GNDA 0.195002f
C2171 VOUT-.n70 GNDA 0.236312f
C2172 VOUT-.t95 GNDA 0.295799f
C2173 VOUT-.t43 GNDA 0.290845f
C2174 VOUT-.n71 GNDA 0.195002f
C2175 VOUT-.t145 GNDA 0.290845f
C2176 VOUT-.t66 GNDA 0.295799f
C2177 VOUT-.t118 GNDA 0.290845f
C2178 VOUT-.n72 GNDA 0.195002f
C2179 VOUT-.n73 GNDA 0.236312f
C2180 VOUT-.t55 GNDA 0.295799f
C2181 VOUT-.t141 GNDA 0.290845f
C2182 VOUT-.n74 GNDA 0.195002f
C2183 VOUT-.t111 GNDA 0.290845f
C2184 VOUT-.t29 GNDA 0.295799f
C2185 VOUT-.t80 GNDA 0.290845f
C2186 VOUT-.n75 GNDA 0.195002f
C2187 VOUT-.n76 GNDA 0.236312f
C2188 VOUT-.t91 GNDA 0.295799f
C2189 VOUT-.t39 GNDA 0.290845f
C2190 VOUT-.n77 GNDA 0.195002f
C2191 VOUT-.t139 GNDA 0.290845f
C2192 VOUT-.t58 GNDA 0.295799f
C2193 VOUT-.t109 GNDA 0.290845f
C2194 VOUT-.n78 GNDA 0.195002f
C2195 VOUT-.n79 GNDA 0.236312f
C2196 VOUT-.t49 GNDA 0.295799f
C2197 VOUT-.t135 GNDA 0.290845f
C2198 VOUT-.n80 GNDA 0.195002f
C2199 VOUT-.t103 GNDA 0.290845f
C2200 VOUT-.t20 GNDA 0.295799f
C2201 VOUT-.t72 GNDA 0.290845f
C2202 VOUT-.n81 GNDA 0.195002f
C2203 VOUT-.n82 GNDA 0.236312f
C2204 VOUT-.t148 GNDA 0.295799f
C2205 VOUT-.t99 GNDA 0.290845f
C2206 VOUT-.n83 GNDA 0.195002f
C2207 VOUT-.t68 GNDA 0.290845f
C2208 VOUT-.t122 GNDA 0.295799f
C2209 VOUT-.t33 GNDA 0.290845f
C2210 VOUT-.n84 GNDA 0.195002f
C2211 VOUT-.n85 GNDA 0.236312f
C2212 VOUT-.t44 GNDA 0.295799f
C2213 VOUT-.t133 GNDA 0.290845f
C2214 VOUT-.n86 GNDA 0.195002f
C2215 VOUT-.t98 GNDA 0.290845f
C2216 VOUT-.t152 GNDA 0.295799f
C2217 VOUT-.t67 GNDA 0.290845f
C2218 VOUT-.n87 GNDA 0.195002f
C2219 VOUT-.n88 GNDA 0.236312f
C2220 VOUT-.t142 GNDA 0.295799f
C2221 VOUT-.t94 GNDA 0.290845f
C2222 VOUT-.n89 GNDA 0.195002f
C2223 VOUT-.t60 GNDA 0.290845f
C2224 VOUT-.t116 GNDA 0.295799f
C2225 VOUT-.t30 GNDA 0.290845f
C2226 VOUT-.n90 GNDA 0.195002f
C2227 VOUT-.n91 GNDA 0.236312f
C2228 VOUT-.t77 GNDA 0.295799f
C2229 VOUT-.t127 GNDA 0.290845f
C2230 VOUT-.n92 GNDA 0.195002f
C2231 VOUT-.t22 GNDA 0.290845f
C2232 VOUT-.n93 GNDA 0.236312f
C2233 VOUT-.t53 GNDA 0.290845f
C2234 VOUT-.n94 GNDA 0.127245f
C2235 VOUT-.t105 GNDA 0.290845f
C2236 VOUT-.n95 GNDA 0.231292f
C2237 VOUT-.n96 GNDA 0.2787f
C2238 two_stage_opamp_dummy_magic_0.VD2.t20 GNDA 0.013877f
C2239 two_stage_opamp_dummy_magic_0.VD2.t11 GNDA 0.013877f
C2240 two_stage_opamp_dummy_magic_0.VD2.t8 GNDA 0.013877f
C2241 two_stage_opamp_dummy_magic_0.VD2.n0 GNDA 0.048872f
C2242 two_stage_opamp_dummy_magic_0.VD2.t1 GNDA 0.013877f
C2243 two_stage_opamp_dummy_magic_0.VD2.t17 GNDA 0.013877f
C2244 two_stage_opamp_dummy_magic_0.VD2.n1 GNDA 0.047884f
C2245 two_stage_opamp_dummy_magic_0.VD2.n2 GNDA 0.193373f
C2246 two_stage_opamp_dummy_magic_0.VD2.t13 GNDA 0.013877f
C2247 two_stage_opamp_dummy_magic_0.VD2.t15 GNDA 0.013877f
C2248 two_stage_opamp_dummy_magic_0.VD2.n3 GNDA 0.047884f
C2249 two_stage_opamp_dummy_magic_0.VD2.n4 GNDA 0.140662f
C2250 two_stage_opamp_dummy_magic_0.VD2.t3 GNDA 0.013877f
C2251 two_stage_opamp_dummy_magic_0.VD2.t21 GNDA 0.013877f
C2252 two_stage_opamp_dummy_magic_0.VD2.n5 GNDA 0.04687f
C2253 two_stage_opamp_dummy_magic_0.VD2.t7 GNDA 0.013877f
C2254 two_stage_opamp_dummy_magic_0.VD2.t4 GNDA 0.013877f
C2255 two_stage_opamp_dummy_magic_0.VD2.n6 GNDA 0.050131f
C2256 two_stage_opamp_dummy_magic_0.VD2.t19 GNDA 0.013877f
C2257 two_stage_opamp_dummy_magic_0.VD2.t10 GNDA 0.013877f
C2258 two_stage_opamp_dummy_magic_0.VD2.n7 GNDA 0.050131f
C2259 two_stage_opamp_dummy_magic_0.VD2.t12 GNDA 0.013877f
C2260 two_stage_opamp_dummy_magic_0.VD2.t9 GNDA 0.013877f
C2261 two_stage_opamp_dummy_magic_0.VD2.n8 GNDA 0.04969f
C2262 two_stage_opamp_dummy_magic_0.VD2.n9 GNDA 0.186051f
C2263 two_stage_opamp_dummy_magic_0.VD2.t6 GNDA 0.013877f
C2264 two_stage_opamp_dummy_magic_0.VD2.t5 GNDA 0.013877f
C2265 two_stage_opamp_dummy_magic_0.VD2.n10 GNDA 0.04969f
C2266 two_stage_opamp_dummy_magic_0.VD2.n11 GNDA 0.096484f
C2267 two_stage_opamp_dummy_magic_0.VD2.n12 GNDA 0.117322f
C2268 two_stage_opamp_dummy_magic_0.VD2.n13 GNDA 0.081264f
C2269 two_stage_opamp_dummy_magic_0.VD2.t18 GNDA 0.013877f
C2270 two_stage_opamp_dummy_magic_0.VD2.t0 GNDA 0.013877f
C2271 two_stage_opamp_dummy_magic_0.VD2.n14 GNDA 0.045463f
C2272 two_stage_opamp_dummy_magic_0.VD2.n15 GNDA 0.069533f
C2273 two_stage_opamp_dummy_magic_0.VD2.n16 GNDA 0.083264f
C2274 two_stage_opamp_dummy_magic_0.VD2.t2 GNDA 0.013877f
C2275 two_stage_opamp_dummy_magic_0.VD2.t14 GNDA 0.013877f
C2276 two_stage_opamp_dummy_magic_0.VD2.n17 GNDA 0.047884f
C2277 two_stage_opamp_dummy_magic_0.VD2.n18 GNDA 0.193373f
C2278 two_stage_opamp_dummy_magic_0.VD2.n19 GNDA 0.048872f
C2279 two_stage_opamp_dummy_magic_0.VD2.t16 GNDA 0.013877f
C2280 bgr_0.V_TOP.t24 GNDA 0.107607f
C2281 bgr_0.V_TOP.t33 GNDA 0.107607f
C2282 bgr_0.V_TOP.t39 GNDA 0.107607f
C2283 bgr_0.V_TOP.t16 GNDA 0.107607f
C2284 bgr_0.V_TOP.t15 GNDA 0.107607f
C2285 bgr_0.V_TOP.t28 GNDA 0.107607f
C2286 bgr_0.V_TOP.t38 GNDA 0.107607f
C2287 bgr_0.V_TOP.t14 GNDA 0.107607f
C2288 bgr_0.V_TOP.t27 GNDA 0.107607f
C2289 bgr_0.V_TOP.t26 GNDA 0.107607f
C2290 bgr_0.V_TOP.t37 GNDA 0.107607f
C2291 bgr_0.V_TOP.t46 GNDA 0.107607f
C2292 bgr_0.V_TOP.t18 GNDA 0.107607f
C2293 bgr_0.V_TOP.t30 GNDA 0.107607f
C2294 bgr_0.V_TOP.t29 GNDA 0.140668f
C2295 bgr_0.V_TOP.n0 GNDA 0.078644f
C2296 bgr_0.V_TOP.n1 GNDA 0.05739f
C2297 bgr_0.V_TOP.n2 GNDA 0.05739f
C2298 bgr_0.V_TOP.n3 GNDA 0.05739f
C2299 bgr_0.V_TOP.n4 GNDA 0.05739f
C2300 bgr_0.V_TOP.n5 GNDA 0.053518f
C2301 bgr_0.V_TOP.t9 GNDA 0.138382f
C2302 bgr_0.V_TOP.t40 GNDA 0.40993f
C2303 bgr_0.V_TOP.t31 GNDA 0.416912f
C2304 bgr_0.V_TOP.t35 GNDA 0.40993f
C2305 bgr_0.V_TOP.n6 GNDA 0.274845f
C2306 bgr_0.V_TOP.t32 GNDA 0.40993f
C2307 bgr_0.V_TOP.t22 GNDA 0.416912f
C2308 bgr_0.V_TOP.n7 GNDA 0.351706f
C2309 bgr_0.V_TOP.t20 GNDA 0.416912f
C2310 bgr_0.V_TOP.t25 GNDA 0.40993f
C2311 bgr_0.V_TOP.n8 GNDA 0.274845f
C2312 bgr_0.V_TOP.t21 GNDA 0.40993f
C2313 bgr_0.V_TOP.t45 GNDA 0.416912f
C2314 bgr_0.V_TOP.n9 GNDA 0.428568f
C2315 bgr_0.V_TOP.t42 GNDA 0.416912f
C2316 bgr_0.V_TOP.t49 GNDA 0.40993f
C2317 bgr_0.V_TOP.n10 GNDA 0.274845f
C2318 bgr_0.V_TOP.t44 GNDA 0.40993f
C2319 bgr_0.V_TOP.t36 GNDA 0.416912f
C2320 bgr_0.V_TOP.n11 GNDA 0.428568f
C2321 bgr_0.V_TOP.t17 GNDA 0.416912f
C2322 bgr_0.V_TOP.t23 GNDA 0.40993f
C2323 bgr_0.V_TOP.n12 GNDA 0.274845f
C2324 bgr_0.V_TOP.t19 GNDA 0.40993f
C2325 bgr_0.V_TOP.t43 GNDA 0.416912f
C2326 bgr_0.V_TOP.n13 GNDA 0.428568f
C2327 bgr_0.V_TOP.t34 GNDA 0.416912f
C2328 bgr_0.V_TOP.t41 GNDA 0.40993f
C2329 bgr_0.V_TOP.n14 GNDA 0.351706f
C2330 bgr_0.V_TOP.t47 GNDA 0.40993f
C2331 bgr_0.V_TOP.n15 GNDA 0.179344f
C2332 bgr_0.V_TOP.n16 GNDA 0.613759f
C2333 bgr_0.V_TOP.t2 GNDA 0.115319f
C2334 bgr_0.V_TOP.n17 GNDA 0.816567f
C2335 bgr_0.V_TOP.t10 GNDA 0.010248f
C2336 bgr_0.V_TOP.t7 GNDA 0.010248f
C2337 bgr_0.V_TOP.n18 GNDA 0.025517f
C2338 bgr_0.V_TOP.n19 GNDA 0.46747f
C2339 bgr_0.V_TOP.t5 GNDA 0.010248f
C2340 bgr_0.V_TOP.t1 GNDA 0.010248f
C2341 bgr_0.V_TOP.n20 GNDA 0.024716f
C2342 bgr_0.V_TOP.t12 GNDA 0.010248f
C2343 bgr_0.V_TOP.t4 GNDA 0.010248f
C2344 bgr_0.V_TOP.n21 GNDA 0.025689f
C2345 bgr_0.V_TOP.t3 GNDA 0.010248f
C2346 bgr_0.V_TOP.t13 GNDA 0.010248f
C2347 bgr_0.V_TOP.n22 GNDA 0.025517f
C2348 bgr_0.V_TOP.n23 GNDA 0.236477f
C2349 bgr_0.V_TOP.n24 GNDA 0.143648f
C2350 bgr_0.V_TOP.n25 GNDA 0.081986f
C2351 bgr_0.V_TOP.t6 GNDA 0.010248f
C2352 bgr_0.V_TOP.t8 GNDA 0.010248f
C2353 bgr_0.V_TOP.n26 GNDA 0.025517f
C2354 bgr_0.V_TOP.n27 GNDA 0.141529f
C2355 bgr_0.V_TOP.t0 GNDA 0.010248f
C2356 bgr_0.V_TOP.t11 GNDA 0.010248f
C2357 bgr_0.V_TOP.n28 GNDA 0.025517f
C2358 bgr_0.V_TOP.n29 GNDA 0.140184f
C2359 bgr_0.V_TOP.n30 GNDA 0.308147f
C2360 bgr_0.V_TOP.n31 GNDA 0.021684f
C2361 bgr_0.V_TOP.n32 GNDA 0.053518f
C2362 bgr_0.V_TOP.n33 GNDA 0.05739f
C2363 bgr_0.V_TOP.n34 GNDA 0.05739f
C2364 bgr_0.V_TOP.n35 GNDA 0.05739f
C2365 bgr_0.V_TOP.n36 GNDA 0.05739f
C2366 bgr_0.V_TOP.n37 GNDA 0.05739f
C2367 bgr_0.V_TOP.n38 GNDA 0.05739f
C2368 bgr_0.V_TOP.n39 GNDA 0.053518f
C2369 bgr_0.V_TOP.t48 GNDA 0.124001f
C2370 VDDA.t3 GNDA 0.019167f
C2371 VDDA.t316 GNDA 0.019167f
C2372 VDDA.n0 GNDA 0.079263f
C2373 VDDA.t215 GNDA 0.019167f
C2374 VDDA.t71 GNDA 0.019167f
C2375 VDDA.n1 GNDA 0.078959f
C2376 VDDA.n2 GNDA 0.109472f
C2377 VDDA.t8 GNDA 0.019167f
C2378 VDDA.t81 GNDA 0.019167f
C2379 VDDA.n3 GNDA 0.078959f
C2380 VDDA.n4 GNDA 0.057124f
C2381 VDDA.t94 GNDA 0.019167f
C2382 VDDA.t113 GNDA 0.019167f
C2383 VDDA.n5 GNDA 0.078959f
C2384 VDDA.n6 GNDA 0.057124f
C2385 VDDA.t59 GNDA 0.019167f
C2386 VDDA.t126 GNDA 0.019167f
C2387 VDDA.n7 GNDA 0.078959f
C2388 VDDA.n8 GNDA 0.057124f
C2389 VDDA.t314 GNDA 0.019167f
C2390 VDDA.t72 GNDA 0.019167f
C2391 VDDA.n9 GNDA 0.078959f
C2392 VDDA.n10 GNDA 0.135749f
C2393 VDDA.n11 GNDA 0.061892f
C2394 VDDA.n12 GNDA 0.165234f
C2395 VDDA.t323 GNDA 0.012038f
C2396 VDDA.n13 GNDA 0.025615f
C2397 VDDA.t426 GNDA 0.012038f
C2398 VDDA.n14 GNDA 0.025615f
C2399 VDDA.n15 GNDA 0.037192f
C2400 VDDA.n16 GNDA 0.062513f
C2401 VDDA.n17 GNDA 0.166598f
C2402 VDDA.t384 GNDA 0.012038f
C2403 VDDA.n18 GNDA 0.025615f
C2404 VDDA.t360 GNDA 0.012038f
C2405 VDDA.n19 GNDA 0.025615f
C2406 VDDA.n20 GNDA 0.03466f
C2407 VDDA.n21 GNDA 0.043024f
C2408 VDDA.n22 GNDA 0.166598f
C2409 VDDA.t359 GNDA 0.162068f
C2410 VDDA.t147 GNDA 0.100146f
C2411 VDDA.t68 GNDA 0.100146f
C2412 VDDA.t13 GNDA 0.100146f
C2413 VDDA.t117 GNDA 0.100146f
C2414 VDDA.t121 GNDA 0.075109f
C2415 VDDA.t383 GNDA 0.162068f
C2416 VDDA.t33 GNDA 0.100146f
C2417 VDDA.t120 GNDA 0.100146f
C2418 VDDA.t455 GNDA 0.100146f
C2419 VDDA.t197 GNDA 0.100146f
C2420 VDDA.t35 GNDA 0.075109f
C2421 VDDA.n23 GNDA 0.063133f
C2422 VDDA.n24 GNDA 0.050073f
C2423 VDDA.n25 GNDA 0.063133f
C2424 VDDA.n26 GNDA 0.042167f
C2425 VDDA.n27 GNDA 0.034117f
C2426 VDDA.n28 GNDA 0.079326f
C2427 VDDA.n29 GNDA 0.079326f
C2428 VDDA.n30 GNDA 0.165234f
C2429 VDDA.t425 GNDA 0.1588f
C2430 VDDA.t146 GNDA 0.098389f
C2431 VDDA.t112 GNDA 0.098389f
C2432 VDDA.t433 GNDA 0.098389f
C2433 VDDA.t119 GNDA 0.098389f
C2434 VDDA.t122 GNDA 0.073792f
C2435 VDDA.t322 GNDA 0.1588f
C2436 VDDA.t450 GNDA 0.098389f
C2437 VDDA.t118 GNDA 0.098389f
C2438 VDDA.t148 GNDA 0.098389f
C2439 VDDA.t34 GNDA 0.098389f
C2440 VDDA.t251 GNDA 0.073792f
C2441 VDDA.n31 GNDA 0.063133f
C2442 VDDA.n32 GNDA 0.049194f
C2443 VDDA.n33 GNDA 0.063133f
C2444 VDDA.n34 GNDA 0.041966f
C2445 VDDA.n35 GNDA 0.034117f
C2446 VDDA.n36 GNDA 0.066047f
C2447 VDDA.n37 GNDA 0.19628f
C2448 VDDA.t80 GNDA 0.038333f
C2449 VDDA.t20 GNDA 0.038333f
C2450 VDDA.n38 GNDA 0.153788f
C2451 VDDA.n39 GNDA 0.078128f
C2452 VDDA.t329 GNDA 0.038187f
C2453 VDDA.n40 GNDA 0.077493f
C2454 VDDA.n41 GNDA 0.051708f
C2455 VDDA.n42 GNDA 0.072986f
C2456 VDDA.t363 GNDA 0.04241f
C2457 VDDA.t361 GNDA 0.018572f
C2458 VDDA.n43 GNDA 0.067275f
C2459 VDDA.n44 GNDA 0.039604f
C2460 VDDA.t335 GNDA 0.04241f
C2461 VDDA.t333 GNDA 0.018572f
C2462 VDDA.n45 GNDA 0.067275f
C2463 VDDA.n46 GNDA 0.039604f
C2464 VDDA.n47 GNDA 0.042167f
C2465 VDDA.n48 GNDA 0.072986f
C2466 VDDA.n49 GNDA 0.210995f
C2467 VDDA.t334 GNDA 0.261311f
C2468 VDDA.t238 GNDA 0.151097f
C2469 VDDA.t18 GNDA 0.151097f
C2470 VDDA.t216 GNDA 0.151097f
C2471 VDDA.t96 GNDA 0.151097f
C2472 VDDA.t149 GNDA 0.113323f
C2473 VDDA.n50 GNDA 0.075549f
C2474 VDDA.t127 GNDA 0.113323f
C2475 VDDA.t56 GNDA 0.151097f
C2476 VDDA.t125 GNDA 0.151097f
C2477 VDDA.t114 GNDA 0.151097f
C2478 VDDA.t95 GNDA 0.151097f
C2479 VDDA.t362 GNDA 0.261311f
C2480 VDDA.n51 GNDA 0.210995f
C2481 VDDA.n52 GNDA 0.051708f
C2482 VDDA.n53 GNDA 0.097848f
C2483 VDDA.t354 GNDA 0.038187f
C2484 VDDA.t218 GNDA 0.038333f
C2485 VDDA.t58 GNDA 0.038333f
C2486 VDDA.n54 GNDA 0.153788f
C2487 VDDA.n55 GNDA 0.078128f
C2488 VDDA.t55 GNDA 0.038333f
C2489 VDDA.t124 GNDA 0.038333f
C2490 VDDA.n56 GNDA 0.153788f
C2491 VDDA.n57 GNDA 0.078128f
C2492 VDDA.t5 GNDA 0.038333f
C2493 VDDA.t7 GNDA 0.038333f
C2494 VDDA.n58 GNDA 0.153788f
C2495 VDDA.n59 GNDA 0.078128f
C2496 VDDA.t240 GNDA 0.038333f
C2497 VDDA.t151 GNDA 0.038333f
C2498 VDDA.n60 GNDA 0.153788f
C2499 VDDA.n61 GNDA 0.164176f
C2500 VDDA.n62 GNDA 0.123956f
C2501 VDDA.t352 GNDA 0.046334f
C2502 VDDA.n63 GNDA 0.088651f
C2503 VDDA.n64 GNDA 0.051792f
C2504 VDDA.n65 GNDA 0.341097f
C2505 VDDA.n66 GNDA 0.341097f
C2506 VDDA.t328 GNDA 0.526859f
C2507 VDDA.t79 GNDA 0.291653f
C2508 VDDA.t19 GNDA 0.291653f
C2509 VDDA.t217 GNDA 0.291653f
C2510 VDDA.t57 GNDA 0.291653f
C2511 VDDA.t54 GNDA 0.21874f
C2512 VDDA.n67 GNDA 0.077493f
C2513 VDDA.n68 GNDA 0.099326f
C2514 VDDA.n69 GNDA 0.099326f
C2515 VDDA.t353 GNDA 0.526859f
C2516 VDDA.t150 GNDA 0.291653f
C2517 VDDA.t239 GNDA 0.291653f
C2518 VDDA.t6 GNDA 0.291653f
C2519 VDDA.t4 GNDA 0.291653f
C2520 VDDA.t123 GNDA 0.21874f
C2521 VDDA.n70 GNDA 0.145826f
C2522 VDDA.n71 GNDA 0.098679f
C2523 VDDA.n72 GNDA 0.066964f
C2524 VDDA.n73 GNDA 0.051792f
C2525 VDDA.t327 GNDA 0.046334f
C2526 VDDA.n74 GNDA 0.088651f
C2527 VDDA.n75 GNDA 0.123636f
C2528 VDDA.n76 GNDA 0.110006f
C2529 VDDA.n77 GNDA 0.093597f
C2530 VDDA.t289 GNDA 0.022361f
C2531 VDDA.t297 GNDA 0.022361f
C2532 VDDA.n78 GNDA 0.077767f
C2533 VDDA.t309 GNDA 0.022361f
C2534 VDDA.t303 GNDA 0.022361f
C2535 VDDA.n79 GNDA 0.077492f
C2536 VDDA.n80 GNDA 0.146297f
C2537 VDDA.t295 GNDA 0.022361f
C2538 VDDA.t307 GNDA 0.022361f
C2539 VDDA.n81 GNDA 0.077767f
C2540 VDDA.t277 GNDA 0.022361f
C2541 VDDA.t299 GNDA 0.022361f
C2542 VDDA.n82 GNDA 0.077492f
C2543 VDDA.n83 GNDA 0.146297f
C2544 VDDA.n84 GNDA 0.020444f
C2545 VDDA.n85 GNDA 0.06366f
C2546 VDDA.n86 GNDA 0.086565f
C2547 VDDA.t420 GNDA 0.110312f
C2548 VDDA.t418 GNDA 0.038938f
C2549 VDDA.n87 GNDA 0.071965f
C2550 VDDA.n88 GNDA 0.046392f
C2551 VDDA.t369 GNDA 0.110312f
C2552 VDDA.t367 GNDA 0.038938f
C2553 VDDA.n89 GNDA 0.071965f
C2554 VDDA.n90 GNDA 0.046392f
C2555 VDDA.n91 GNDA 0.046f
C2556 VDDA.n92 GNDA 0.086565f
C2557 VDDA.n93 GNDA 0.257978f
C2558 VDDA.t368 GNDA 0.385069f
C2559 VDDA.t288 GNDA 0.222333f
C2560 VDDA.t296 GNDA 0.222333f
C2561 VDDA.t308 GNDA 0.222333f
C2562 VDDA.t302 GNDA 0.222333f
C2563 VDDA.t312 GNDA 0.16675f
C2564 VDDA.n94 GNDA 0.111167f
C2565 VDDA.t272 GNDA 0.16675f
C2566 VDDA.t276 GNDA 0.222333f
C2567 VDDA.t298 GNDA 0.222333f
C2568 VDDA.t294 GNDA 0.222333f
C2569 VDDA.t306 GNDA 0.222333f
C2570 VDDA.t419 GNDA 0.385069f
C2571 VDDA.n95 GNDA 0.257978f
C2572 VDDA.n96 GNDA 0.06366f
C2573 VDDA.n97 GNDA 0.08912f
C2574 VDDA.t313 GNDA 0.022361f
C2575 VDDA.t273 GNDA 0.022361f
C2576 VDDA.n98 GNDA 0.072907f
C2577 VDDA.n99 GNDA 0.04976f
C2578 VDDA.n100 GNDA 0.041588f
C2579 VDDA.t315 GNDA 0.019167f
C2580 VDDA.t87 GNDA 0.019167f
C2581 VDDA.n101 GNDA 0.079263f
C2582 VDDA.t243 GNDA 0.019167f
C2583 VDDA.t456 GNDA 0.019167f
C2584 VDDA.n102 GNDA 0.078959f
C2585 VDDA.n103 GNDA 0.109472f
C2586 VDDA.t241 GNDA 0.019167f
C2587 VDDA.t88 GNDA 0.019167f
C2588 VDDA.n104 GNDA 0.078959f
C2589 VDDA.n105 GNDA 0.057124f
C2590 VDDA.t25 GNDA 0.019167f
C2591 VDDA.t231 GNDA 0.019167f
C2592 VDDA.n106 GNDA 0.078959f
C2593 VDDA.n107 GNDA 0.057124f
C2594 VDDA.t86 GNDA 0.019167f
C2595 VDDA.t439 GNDA 0.019167f
C2596 VDDA.n108 GNDA 0.078959f
C2597 VDDA.n109 GNDA 0.057124f
C2598 VDDA.t438 GNDA 0.019167f
C2599 VDDA.t317 GNDA 0.019167f
C2600 VDDA.n110 GNDA 0.078959f
C2601 VDDA.n111 GNDA 0.164553f
C2602 VDDA.t466 GNDA 0.038333f
C2603 VDDA.t203 GNDA 0.038333f
C2604 VDDA.n112 GNDA 0.153788f
C2605 VDDA.n113 GNDA 0.078128f
C2606 VDDA.t375 GNDA 0.038187f
C2607 VDDA.n114 GNDA 0.051708f
C2608 VDDA.n115 GNDA 0.072986f
C2609 VDDA.t381 GNDA 0.04241f
C2610 VDDA.t379 GNDA 0.018572f
C2611 VDDA.n116 GNDA 0.067275f
C2612 VDDA.n117 GNDA 0.039604f
C2613 VDDA.t357 GNDA 0.04241f
C2614 VDDA.t355 GNDA 0.018572f
C2615 VDDA.n118 GNDA 0.067275f
C2616 VDDA.n119 GNDA 0.039604f
C2617 VDDA.n120 GNDA 0.042167f
C2618 VDDA.n121 GNDA 0.072986f
C2619 VDDA.n122 GNDA 0.210995f
C2620 VDDA.t356 GNDA 0.261311f
C2621 VDDA.t156 GNDA 0.151097f
C2622 VDDA.t0 GNDA 0.151097f
C2623 VDDA.t444 GNDA 0.151097f
C2624 VDDA.t26 GNDA 0.151097f
C2625 VDDA.t230 GNDA 0.113323f
C2626 VDDA.n123 GNDA 0.075549f
C2627 VDDA.t206 GNDA 0.113323f
C2628 VDDA.t242 GNDA 0.151097f
C2629 VDDA.t190 GNDA 0.151097f
C2630 VDDA.t445 GNDA 0.151097f
C2631 VDDA.t187 GNDA 0.151097f
C2632 VDDA.t380 GNDA 0.261311f
C2633 VDDA.n124 GNDA 0.210995f
C2634 VDDA.n125 GNDA 0.051708f
C2635 VDDA.n126 GNDA 0.097848f
C2636 VDDA.n127 GNDA 0.066964f
C2637 VDDA.n128 GNDA 0.099326f
C2638 VDDA.n129 GNDA 0.099326f
C2639 VDDA.n130 GNDA 0.098679f
C2640 VDDA.t348 GNDA 0.038187f
C2641 VDDA.t205 GNDA 0.038333f
C2642 VDDA.t24 GNDA 0.038333f
C2643 VDDA.n131 GNDA 0.153788f
C2644 VDDA.n132 GNDA 0.078128f
C2645 VDDA.t189 GNDA 0.038333f
C2646 VDDA.t229 GNDA 0.038333f
C2647 VDDA.n133 GNDA 0.153788f
C2648 VDDA.n134 GNDA 0.078128f
C2649 VDDA.t160 GNDA 0.038333f
C2650 VDDA.t235 GNDA 0.038333f
C2651 VDDA.n135 GNDA 0.153788f
C2652 VDDA.n136 GNDA 0.078128f
C2653 VDDA.t452 GNDA 0.038333f
C2654 VDDA.t233 GNDA 0.038333f
C2655 VDDA.n137 GNDA 0.153788f
C2656 VDDA.n138 GNDA 0.164176f
C2657 VDDA.n139 GNDA 0.123956f
C2658 VDDA.t346 GNDA 0.046334f
C2659 VDDA.n140 GNDA 0.088651f
C2660 VDDA.n141 GNDA 0.051792f
C2661 VDDA.n142 GNDA 0.077493f
C2662 VDDA.n143 GNDA 0.341097f
C2663 VDDA.t347 GNDA 0.526859f
C2664 VDDA.t451 GNDA 0.291653f
C2665 VDDA.t232 GNDA 0.291653f
C2666 VDDA.t159 GNDA 0.291653f
C2667 VDDA.t234 GNDA 0.291653f
C2668 VDDA.t188 GNDA 0.21874f
C2669 VDDA.n144 GNDA 0.145826f
C2670 VDDA.t228 GNDA 0.21874f
C2671 VDDA.t204 GNDA 0.291653f
C2672 VDDA.t23 GNDA 0.291653f
C2673 VDDA.t465 GNDA 0.291653f
C2674 VDDA.t202 GNDA 0.291653f
C2675 VDDA.t374 GNDA 0.526859f
C2676 VDDA.n145 GNDA 0.341097f
C2677 VDDA.n146 GNDA 0.077493f
C2678 VDDA.n147 GNDA 0.051792f
C2679 VDDA.t373 GNDA 0.046334f
C2680 VDDA.n148 GNDA 0.088651f
C2681 VDDA.n149 GNDA 0.123636f
C2682 VDDA.n150 GNDA 0.094353f
C2683 VDDA.n152 GNDA 0.048918f
C2684 VDDA.n153 GNDA 0.060687f
C2685 VDDA.n155 GNDA 0.048918f
C2686 VDDA.n157 GNDA 0.048918f
C2687 VDDA.n159 GNDA 0.048918f
C2688 VDDA.n161 GNDA 0.048918f
C2689 VDDA.n163 GNDA 0.048918f
C2690 VDDA.n165 GNDA 0.048918f
C2691 VDDA.n167 GNDA 0.048918f
C2692 VDDA.n169 GNDA 0.048918f
C2693 VDDA.n171 GNDA 0.08005f
C2694 VDDA.t405 GNDA 0.01164f
C2695 VDDA.n172 GNDA 0.017283f
C2696 VDDA.n173 GNDA 0.015292f
C2697 VDDA.n174 GNDA 0.052229f
C2698 VDDA.n175 GNDA 0.200561f
C2699 VDDA.n176 GNDA 0.200561f
C2700 VDDA.t413 GNDA 0.1588f
C2701 VDDA.t40 GNDA 0.098389f
C2702 VDDA.t105 GNDA 0.098389f
C2703 VDDA.t175 GNDA 0.098389f
C2704 VDDA.t103 GNDA 0.098389f
C2705 VDDA.t169 GNDA 0.098389f
C2706 VDDA.t179 GNDA 0.098389f
C2707 VDDA.t62 GNDA 0.098389f
C2708 VDDA.t185 GNDA 0.098389f
C2709 VDDA.t14 GNDA 0.098389f
C2710 VDDA.t49 GNDA 0.073792f
C2711 VDDA.t404 GNDA 0.1588f
C2712 VDDA.t99 GNDA 0.098389f
C2713 VDDA.t47 GNDA 0.098389f
C2714 VDDA.t181 GNDA 0.098389f
C2715 VDDA.t183 GNDA 0.098389f
C2716 VDDA.t171 GNDA 0.098389f
C2717 VDDA.t177 GNDA 0.098389f
C2718 VDDA.t42 GNDA 0.098389f
C2719 VDDA.t16 GNDA 0.098389f
C2720 VDDA.t173 GNDA 0.098389f
C2721 VDDA.t101 GNDA 0.073792f
C2722 VDDA.n177 GNDA 0.060687f
C2723 VDDA.n178 GNDA 0.098084f
C2724 VDDA.n179 GNDA 0.098084f
C2725 VDDA.n180 GNDA 0.049194f
C2726 VDDA.n181 GNDA 0.098084f
C2727 VDDA.n182 GNDA 0.077306f
C2728 VDDA.n183 GNDA 0.052229f
C2729 VDDA.n184 GNDA 0.015292f
C2730 VDDA.t414 GNDA 0.01164f
C2731 VDDA.n185 GNDA 0.016862f
C2732 VDDA.n186 GNDA 0.060623f
C2733 VDDA.n187 GNDA 0.047278f
C2734 VDDA.n188 GNDA 0.243658f
C2735 VDDA.n189 GNDA 0.23184f
C2736 VDDA.t279 GNDA 0.022361f
C2737 VDDA.t285 GNDA 0.022361f
C2738 VDDA.n190 GNDA 0.077767f
C2739 VDDA.t291 GNDA 0.022361f
C2740 VDDA.t301 GNDA 0.022361f
C2741 VDDA.n191 GNDA 0.077492f
C2742 VDDA.n192 GNDA 0.146297f
C2743 VDDA.t293 GNDA 0.022361f
C2744 VDDA.t305 GNDA 0.022361f
C2745 VDDA.n193 GNDA 0.077767f
C2746 VDDA.t281 GNDA 0.022361f
C2747 VDDA.t287 GNDA 0.022361f
C2748 VDDA.n194 GNDA 0.077492f
C2749 VDDA.n195 GNDA 0.146297f
C2750 VDDA.n196 GNDA 0.020444f
C2751 VDDA.n197 GNDA 0.06366f
C2752 VDDA.n198 GNDA 0.086565f
C2753 VDDA.t399 GNDA 0.110312f
C2754 VDDA.t397 GNDA 0.038938f
C2755 VDDA.n199 GNDA 0.071965f
C2756 VDDA.n200 GNDA 0.046392f
C2757 VDDA.t366 GNDA 0.110312f
C2758 VDDA.t364 GNDA 0.038938f
C2759 VDDA.n201 GNDA 0.071965f
C2760 VDDA.n202 GNDA 0.046392f
C2761 VDDA.n203 GNDA 0.046f
C2762 VDDA.n204 GNDA 0.086565f
C2763 VDDA.n205 GNDA 0.257978f
C2764 VDDA.t365 GNDA 0.385069f
C2765 VDDA.t278 GNDA 0.222333f
C2766 VDDA.t284 GNDA 0.222333f
C2767 VDDA.t290 GNDA 0.222333f
C2768 VDDA.t300 GNDA 0.222333f
C2769 VDDA.t310 GNDA 0.16675f
C2770 VDDA.n206 GNDA 0.111167f
C2771 VDDA.t274 GNDA 0.16675f
C2772 VDDA.t280 GNDA 0.222333f
C2773 VDDA.t286 GNDA 0.222333f
C2774 VDDA.t292 GNDA 0.222333f
C2775 VDDA.t304 GNDA 0.222333f
C2776 VDDA.t398 GNDA 0.385069f
C2777 VDDA.n207 GNDA 0.257978f
C2778 VDDA.n208 GNDA 0.06366f
C2779 VDDA.n209 GNDA 0.08912f
C2780 VDDA.t311 GNDA 0.022361f
C2781 VDDA.t275 GNDA 0.022361f
C2782 VDDA.n210 GNDA 0.072907f
C2783 VDDA.n211 GNDA 0.04976f
C2784 VDDA.n212 GNDA 0.041802f
C2785 VDDA.n213 GNDA 0.200657f
C2786 VDDA.n214 GNDA 0.078583f
C2787 VDDA.n216 GNDA 0.06216f
C2788 VDDA.n217 GNDA 0.0115f
C2789 VDDA.n218 GNDA 0.03397f
C2790 VDDA.n219 GNDA 0.03397f
C2791 VDDA.n220 GNDA 0.034637f
C2792 VDDA.n221 GNDA 0.088266f
C2793 VDDA.n222 GNDA 0.0115f
C2794 VDDA.n223 GNDA 0.052059f
C2795 VDDA.n224 GNDA 0.052059f
C2796 VDDA.n225 GNDA 0.054659f
C2797 VDDA.t283 GNDA 0.022681f
C2798 VDDA.n226 GNDA 0.080893f
C2799 VDDA.t341 GNDA 0.103479f
C2800 VDDA.n227 GNDA 0.050777f
C2801 VDDA.n228 GNDA 0.04732f
C2802 VDDA.t339 GNDA 0.037553f
C2803 VDDA.n229 GNDA 0.040428f
C2804 VDDA.n230 GNDA 0.030544f
C2805 VDDA.n231 GNDA 0.045903f
C2806 VDDA.n232 GNDA 0.308645f
C2807 VDDA.t340 GNDA 0.284429f
C2808 VDDA.n233 GNDA 0.094236f
C2809 VDDA.n234 GNDA 0.023559f
C2810 VDDA.t282 GNDA 0.131931f
C2811 VDDA.t395 GNDA 0.312107f
C2812 VDDA.n235 GNDA 0.307488f
C2813 VDDA.n236 GNDA 0.047538f
C2814 VDDA.n237 GNDA 0.030206f
C2815 VDDA.t394 GNDA 0.039408f
C2816 VDDA.n238 GNDA 0.040428f
C2817 VDDA.t396 GNDA 0.080799f
C2818 VDDA.n239 GNDA 0.054478f
C2819 VDDA.n240 GNDA 0.109416f
C2820 VDDA.n241 GNDA 0.072496f
C2821 VDDA.t332 GNDA 0.014173f
C2822 VDDA.n242 GNDA 0.016004f
C2823 VDDA.t330 GNDA 0.012265f
C2824 VDDA.n243 GNDA 0.016125f
C2825 VDDA.n244 GNDA 0.020424f
C2826 VDDA.n245 GNDA 0.028661f
C2827 VDDA.n246 GNDA 0.152876f
C2828 VDDA.t331 GNDA 0.169321f
C2829 VDDA.t115 GNDA 0.115f
C2830 VDDA.t343 GNDA 0.169321f
C2831 VDDA.n247 GNDA 0.152876f
C2832 VDDA.n248 GNDA 0.028661f
C2833 VDDA.n249 GNDA 0.020424f
C2834 VDDA.t342 GNDA 0.012265f
C2835 VDDA.n250 GNDA 0.016125f
C2836 VDDA.t345 GNDA 0.014173f
C2837 VDDA.n251 GNDA 0.017899f
C2838 VDDA.n252 GNDA 0.070792f
C2839 VDDA.n253 GNDA 0.207133f
C2840 VDDA.n254 GNDA 3.59973f
C2841 VDDA.t463 GNDA 0.357139f
C2842 VDDA.t210 GNDA 0.358433f
C2843 VDDA.t135 GNDA 0.339267f
C2844 VDDA.t111 GNDA 0.357139f
C2845 VDDA.t46 GNDA 0.358433f
C2846 VDDA.t52 GNDA 0.339267f
C2847 VDDA.t51 GNDA 0.357139f
C2848 VDDA.t91 GNDA 0.358433f
C2849 VDDA.t128 GNDA 0.339267f
C2850 VDDA.t78 GNDA 0.357139f
C2851 VDDA.t143 GNDA 0.358433f
C2852 VDDA.t207 GNDA 0.339267f
C2853 VDDA.t139 GNDA 0.357139f
C2854 VDDA.t136 GNDA 0.358433f
C2855 VDDA.t45 GNDA 0.339267f
C2856 VDDA.n255 GNDA 0.239391f
C2857 VDDA.t140 GNDA 0.190639f
C2858 VDDA.n256 GNDA 0.259745f
C2859 VDDA.t44 GNDA 0.190639f
C2860 VDDA.n257 GNDA 0.259745f
C2861 VDDA.t53 GNDA 0.190639f
C2862 VDDA.n258 GNDA 0.259745f
C2863 VDDA.t77 GNDA 0.190639f
C2864 VDDA.n259 GNDA 0.259745f
C2865 VDDA.t464 GNDA 0.333969f
C2866 VDDA.n260 GNDA 3.09101f
C2867 VDDA.t469 GNDA 0.706319f
C2868 VDDA.t470 GNDA 0.752801f
C2869 VDDA.t471 GNDA 0.752801f
C2870 VDDA.t472 GNDA 0.721867f
C2871 VDDA.n261 GNDA 0.504605f
C2872 VDDA.n262 GNDA 0.244984f
C2873 VDDA.n263 GNDA 0.358238f
C2874 VDDA.n264 GNDA 0.661249f
C2875 VDDA.n265 GNDA 0.020444f
C2876 VDDA.n266 GNDA 0.015474f
C2877 VDDA.n267 GNDA 0.015474f
C2878 VDDA.n268 GNDA 0.045221f
C2879 VDDA.n269 GNDA 0.020444f
C2880 VDDA.t393 GNDA 0.024f
C2881 VDDA.t391 GNDA 0.015815f
C2882 VDDA.n270 GNDA 0.03765f
C2883 VDDA.n271 GNDA 0.053572f
C2884 VDDA.n272 GNDA 0.100713f
C2885 VDDA.n273 GNDA 0.100713f
C2886 VDDA.t408 GNDA 0.024f
C2887 VDDA.t406 GNDA 0.015815f
C2888 VDDA.n274 GNDA 0.03765f
C2889 VDDA.n275 GNDA 0.076667f
C2890 VDDA.n276 GNDA 0.053572f
C2891 VDDA.n277 GNDA 0.020444f
C2892 VDDA.n278 GNDA 0.015474f
C2893 VDDA.n279 GNDA 0.016179f
C2894 VDDA.n280 GNDA 0.016069f
C2895 VDDA.n281 GNDA 0.124918f
C2896 VDDA.n282 GNDA 0.016069f
C2897 VDDA.n283 GNDA 0.06507f
C2898 VDDA.n284 GNDA 0.016069f
C2899 VDDA.n285 GNDA 0.06507f
C2900 VDDA.n286 GNDA 0.015474f
C2901 VDDA.n287 GNDA 0.062844f
C2902 VDDA.n288 GNDA 0.100713f
C2903 VDDA.t378 GNDA 0.024f
C2904 VDDA.t376 GNDA 0.015815f
C2905 VDDA.n289 GNDA 0.03765f
C2906 VDDA.n290 GNDA 0.053572f
C2907 VDDA.t338 GNDA 0.024f
C2908 VDDA.t336 GNDA 0.015815f
C2909 VDDA.n291 GNDA 0.03765f
C2910 VDDA.n292 GNDA 0.053572f
C2911 VDDA.n293 GNDA 0.076667f
C2912 VDDA.n294 GNDA 0.100713f
C2913 VDDA.n295 GNDA 0.218978f
C2914 VDDA.t337 GNDA 0.199726f
C2915 VDDA.t256 GNDA 0.1265f
C2916 VDDA.t64 GNDA 0.1265f
C2917 VDDA.t60 GNDA 0.1265f
C2918 VDDA.t260 GNDA 0.1265f
C2919 VDDA.t268 GNDA 0.1265f
C2920 VDDA.t252 GNDA 0.1265f
C2921 VDDA.t157 GNDA 0.1265f
C2922 VDDA.t36 GNDA 0.1265f
C2923 VDDA.t21 GNDA 0.094875f
C2924 VDDA.n296 GNDA 0.06325f
C2925 VDDA.t270 GNDA 0.094875f
C2926 VDDA.t264 GNDA 0.1265f
C2927 VDDA.t254 GNDA 0.1265f
C2928 VDDA.t258 GNDA 0.1265f
C2929 VDDA.t442 GNDA 0.1265f
C2930 VDDA.t436 GNDA 0.1265f
C2931 VDDA.t266 GNDA 0.1265f
C2932 VDDA.t262 GNDA 0.1265f
C2933 VDDA.t82 GNDA 0.1265f
C2934 VDDA.t377 GNDA 0.199726f
C2935 VDDA.n297 GNDA 0.218978f
C2936 VDDA.n298 GNDA 0.062844f
C2937 VDDA.n299 GNDA 0.107057f
C2938 VDDA.n300 GNDA 0.045221f
C2939 VDDA.n301 GNDA 0.020444f
C2940 VDDA.n302 GNDA 0.016069f
C2941 VDDA.n303 GNDA 0.06507f
C2942 VDDA.n304 GNDA 0.016069f
C2943 VDDA.n305 GNDA 0.06507f
C2944 VDDA.n306 GNDA 0.016069f
C2945 VDDA.n307 GNDA 0.06507f
C2946 VDDA.n308 GNDA 0.016069f
C2947 VDDA.n309 GNDA 0.093181f
C2948 VDDA.n310 GNDA 0.020444f
C2949 VDDA.n311 GNDA 0.015474f
C2950 VDDA.n312 GNDA 0.015474f
C2951 VDDA.n313 GNDA 0.045221f
C2952 VDDA.n314 GNDA 0.020444f
C2953 VDDA.n315 GNDA 0.015474f
C2954 VDDA.n316 GNDA 0.020444f
C2955 VDDA.n317 GNDA 0.015474f
C2956 VDDA.n318 GNDA 0.045221f
C2957 VDDA.n319 GNDA 0.020444f
C2958 VDDA.n320 GNDA 0.020444f
C2959 VDDA.n321 GNDA 0.045221f
C2960 VDDA.n322 GNDA 0.020444f
C2961 VDDA.n323 GNDA 0.020444f
C2962 VDDA.n324 GNDA 0.015474f
C2963 VDDA.n325 GNDA 0.045221f
C2964 VDDA.n326 GNDA 0.020444f
C2965 VDDA.n327 GNDA 0.020444f
C2966 VDDA.n328 GNDA 0.045221f
C2967 VDDA.n329 GNDA 0.020444f
C2968 VDDA.n330 GNDA 0.015474f
C2969 VDDA.n331 GNDA 0.045221f
C2970 VDDA.n332 GNDA 0.020444f
C2971 VDDA.n333 GNDA 0.048556f
C2972 VDDA.n334 GNDA 0.045221f
C2973 VDDA.n335 GNDA 0.033379f
C2974 VDDA.n336 GNDA 0.031882f
C2975 VDDA.n337 GNDA 0.218978f
C2976 VDDA.t407 GNDA 0.199726f
C2977 VDDA.t200 GNDA 0.1265f
C2978 VDDA.t38 GNDA 0.1265f
C2979 VDDA.t236 GNDA 0.1265f
C2980 VDDA.t69 GNDA 0.1265f
C2981 VDDA.t11 GNDA 0.1265f
C2982 VDDA.t191 GNDA 0.1265f
C2983 VDDA.t459 GNDA 0.1265f
C2984 VDDA.t434 GNDA 0.1265f
C2985 VDDA.t154 GNDA 0.094875f
C2986 VDDA.n338 GNDA 0.06325f
C2987 VDDA.t198 GNDA 0.094875f
C2988 VDDA.t84 GNDA 0.1265f
C2989 VDDA.t27 GNDA 0.1265f
C2990 VDDA.t225 GNDA 0.1265f
C2991 VDDA.t73 GNDA 0.1265f
C2992 VDDA.t97 GNDA 0.1265f
C2993 VDDA.t9 GNDA 0.1265f
C2994 VDDA.t249 GNDA 0.1265f
C2995 VDDA.t66 GNDA 0.1265f
C2996 VDDA.t392 GNDA 0.199726f
C2997 VDDA.n339 GNDA 0.218978f
C2998 VDDA.n340 GNDA 0.031882f
C2999 VDDA.n341 GNDA 0.033379f
C3000 VDDA.n342 GNDA 0.045221f
C3001 VDDA.n343 GNDA 0.104353f
C3002 VDDA.n344 GNDA 0.219564f
C3003 VDDA.t142 GNDA 0.019167f
C3004 VDDA.t90 GNDA 0.019167f
C3005 VDDA.n345 GNDA 0.063321f
C3006 VDDA.n346 GNDA 0.081707f
C3007 VDDA.t320 GNDA 0.058738f
C3008 VDDA.n347 GNDA 0.1035f
C3009 VDDA.n348 GNDA 0.14109f
C3010 VDDA.n349 GNDA 0.14109f
C3011 VDDA.n350 GNDA 0.140442f
C3012 VDDA.t372 GNDA 0.058738f
C3013 VDDA.t370 GNDA 0.091394f
C3014 VDDA.t402 GNDA 0.024f
C3015 VDDA.t400 GNDA 0.012112f
C3016 VDDA.n351 GNDA 0.037839f
C3017 VDDA.n352 GNDA 0.021819f
C3018 VDDA.n353 GNDA 0.038777f
C3019 VDDA.t432 GNDA 0.024f
C3020 VDDA.t430 GNDA 0.012112f
C3021 VDDA.n354 GNDA 0.037839f
C3022 VDDA.n355 GNDA 0.038777f
C3023 VDDA.n356 GNDA 0.038777f
C3024 VDDA.n357 GNDA 0.031817f
C3025 VDDA.n358 GNDA 0.152894f
C3026 VDDA.t401 GNDA 0.191981f
C3027 VDDA.t248 GNDA 0.086969f
C3028 VDDA.n359 GNDA 0.057979f
C3029 VDDA.t227 GNDA 0.086969f
C3030 VDDA.t431 GNDA 0.194813f
C3031 VDDA.n360 GNDA 0.160605f
C3032 VDDA.n361 GNDA 0.031817f
C3033 VDDA.n362 GNDA 0.021819f
C3034 VDDA.n363 GNDA 0.030653f
C3035 VDDA.t462 GNDA 0.019167f
C3036 VDDA.t134 GNDA 0.019167f
C3037 VDDA.n364 GNDA 0.063321f
C3038 VDDA.n365 GNDA 0.081707f
C3039 VDDA.t108 GNDA 0.019167f
C3040 VDDA.t110 GNDA 0.019167f
C3041 VDDA.n366 GNDA 0.063321f
C3042 VDDA.n367 GNDA 0.081707f
C3043 VDDA.t132 GNDA 0.019167f
C3044 VDDA.t166 GNDA 0.019167f
C3045 VDDA.n368 GNDA 0.063321f
C3046 VDDA.n369 GNDA 0.081707f
C3047 VDDA.t164 GNDA 0.019167f
C3048 VDDA.t468 GNDA 0.019167f
C3049 VDDA.n370 GNDA 0.063321f
C3050 VDDA.n371 GNDA 0.081707f
C3051 VDDA.t130 GNDA 0.019167f
C3052 VDDA.t145 GNDA 0.019167f
C3053 VDDA.n372 GNDA 0.063321f
C3054 VDDA.n373 GNDA 0.081707f
C3055 VDDA.t76 GNDA 0.019167f
C3056 VDDA.t209 GNDA 0.019167f
C3057 VDDA.n374 GNDA 0.063321f
C3058 VDDA.n375 GNDA 0.081707f
C3059 VDDA.t168 GNDA 0.019167f
C3060 VDDA.t138 GNDA 0.019167f
C3061 VDDA.n376 GNDA 0.063321f
C3062 VDDA.n377 GNDA 0.081707f
C3063 VDDA.n378 GNDA 0.090214f
C3064 VDDA.n379 GNDA 0.109076f
C3065 VDDA.n380 GNDA 0.073523f
C3066 VDDA.n381 GNDA 0.089766f
C3067 VDDA.n382 GNDA 0.330743f
C3068 VDDA.t371 GNDA 0.426769f
C3069 VDDA.t167 GNDA 0.307625f
C3070 VDDA.t137 GNDA 0.307625f
C3071 VDDA.t75 GNDA 0.307625f
C3072 VDDA.t208 GNDA 0.307625f
C3073 VDDA.t129 GNDA 0.307625f
C3074 VDDA.t144 GNDA 0.307625f
C3075 VDDA.t163 GNDA 0.307625f
C3076 VDDA.t467 GNDA 0.230719f
C3077 VDDA.n383 GNDA 0.153813f
C3078 VDDA.t131 GNDA 0.230719f
C3079 VDDA.t165 GNDA 0.307625f
C3080 VDDA.t107 GNDA 0.307625f
C3081 VDDA.t109 GNDA 0.307625f
C3082 VDDA.t461 GNDA 0.307625f
C3083 VDDA.t133 GNDA 0.307625f
C3084 VDDA.t141 GNDA 0.307625f
C3085 VDDA.t89 GNDA 0.307625f
C3086 VDDA.t319 GNDA 0.426769f
C3087 VDDA.n384 GNDA 0.330743f
C3088 VDDA.n385 GNDA 0.089766f
C3089 VDDA.n386 GNDA 0.073523f
C3090 VDDA.t318 GNDA 0.091394f
C3091 VDDA.n387 GNDA 0.109076f
C3092 VDDA.n388 GNDA 0.05007f
C3093 VDDA.n389 GNDA 0.01543f
C3094 VDDA.t390 GNDA 0.024178f
C3095 VDDA.t388 GNDA 0.011798f
C3096 VDDA.n390 GNDA 0.036218f
C3097 VDDA.n391 GNDA 0.021719f
C3098 VDDA.n392 GNDA 0.038777f
C3099 VDDA.t387 GNDA 0.024178f
C3100 VDDA.t385 GNDA 0.011798f
C3101 VDDA.n393 GNDA 0.036218f
C3102 VDDA.n394 GNDA 0.038777f
C3103 VDDA.n395 GNDA 0.038777f
C3104 VDDA.n396 GNDA 0.031817f
C3105 VDDA.n397 GNDA 0.152894f
C3106 VDDA.t389 GNDA 0.191981f
C3107 VDDA.t446 GNDA 0.086969f
C3108 VDDA.n398 GNDA 0.057979f
C3109 VDDA.t31 GNDA 0.086969f
C3110 VDDA.t386 GNDA 0.191981f
C3111 VDDA.n399 GNDA 0.152894f
C3112 VDDA.n400 GNDA 0.031817f
C3113 VDDA.n401 GNDA 0.021719f
C3114 VDDA.n402 GNDA 0.022817f
C3115 VDDA.n403 GNDA 0.042709f
C3116 VDDA.n404 GNDA 0.132392f
C3117 VDDA.n405 GNDA 0.17326f
C3118 VDDA.n406 GNDA 0.015937f
C3119 VDDA.n407 GNDA 0.056257f
C3120 VDDA.t423 GNDA 0.025214f
C3121 VDDA.n408 GNDA 0.021083f
C3122 VDDA.n409 GNDA 0.045635f
C3123 VDDA.n410 GNDA 0.045635f
C3124 VDDA.n411 GNDA 0.045635f
C3125 VDDA.t351 GNDA 0.025214f
C3126 VDDA.t349 GNDA 0.012582f
C3127 VDDA.n412 GNDA 0.015908f
C3128 VDDA.n413 GNDA 0.056287f
C3129 VDDA.t411 GNDA 0.024062f
C3130 VDDA.n414 GNDA 0.042167f
C3131 VDDA.n415 GNDA 0.066433f
C3132 VDDA.n416 GNDA 0.066433f
C3133 VDDA.n417 GNDA 0.066433f
C3134 VDDA.t429 GNDA 0.024062f
C3135 VDDA.t427 GNDA 0.012582f
C3136 VDDA.n418 GNDA 0.015944f
C3137 VDDA.n419 GNDA 0.056251f
C3138 VDDA.t326 GNDA 0.025224f
C3139 VDDA.n420 GNDA 0.021083f
C3140 VDDA.n421 GNDA 0.045635f
C3141 VDDA.n422 GNDA 0.045635f
C3142 VDDA.n423 GNDA 0.045635f
C3143 VDDA.t417 GNDA 0.025224f
C3144 VDDA.t415 GNDA 0.012582f
C3145 VDDA.n424 GNDA 0.015944f
C3146 VDDA.n425 GNDA 0.076989f
C3147 VDDA.n426 GNDA 0.043199f
C3148 VDDA.n427 GNDA 0.02578f
C3149 VDDA.n428 GNDA 0.035416f
C3150 VDDA.n429 GNDA 0.161347f
C3151 VDDA.t416 GNDA 0.195358f
C3152 VDDA.t244 GNDA 0.117715f
C3153 VDDA.t453 GNDA 0.088287f
C3154 VDDA.n430 GNDA 0.058858f
C3155 VDDA.t1 GNDA 0.088287f
C3156 VDDA.t448 GNDA 0.117715f
C3157 VDDA.t325 GNDA 0.195358f
C3158 VDDA.n431 GNDA 0.161347f
C3159 VDDA.n432 GNDA 0.035416f
C3160 VDDA.n433 GNDA 0.02578f
C3161 VDDA.t324 GNDA 0.012981f
C3162 VDDA.n434 GNDA 0.042753f
C3163 VDDA.n435 GNDA 0.038833f
C3164 VDDA.n436 GNDA 0.015908f
C3165 VDDA.n437 GNDA 0.056287f
C3166 VDDA.n438 GNDA 0.015908f
C3167 VDDA.n439 GNDA 0.056287f
C3168 VDDA.n440 GNDA 0.015908f
C3169 VDDA.n441 GNDA 0.056287f
C3170 VDDA.n442 GNDA 0.015908f
C3171 VDDA.n443 GNDA 0.056287f
C3172 VDDA.n444 GNDA 0.038833f
C3173 VDDA.n445 GNDA 0.043516f
C3174 VDDA.n446 GNDA 0.039836f
C3175 VDDA.n447 GNDA 0.049648f
C3176 VDDA.n448 GNDA 0.189811f
C3177 VDDA.t428 GNDA 0.195358f
C3178 VDDA.t440 GNDA 0.117715f
C3179 VDDA.t219 GNDA 0.117715f
C3180 VDDA.t213 GNDA 0.117715f
C3181 VDDA.t92 GNDA 0.117715f
C3182 VDDA.t29 GNDA 0.117715f
C3183 VDDA.t195 GNDA 0.088287f
C3184 VDDA.n449 GNDA 0.058858f
C3185 VDDA.t221 GNDA 0.088287f
C3186 VDDA.t193 GNDA 0.117715f
C3187 VDDA.t457 GNDA 0.117715f
C3188 VDDA.t152 GNDA 0.117715f
C3189 VDDA.t410 GNDA 0.195358f
C3190 VDDA.n450 GNDA 0.175621f
C3191 VDDA.n451 GNDA 0.042553f
C3192 VDDA.n452 GNDA 0.032808f
C3193 VDDA.t409 GNDA 0.012582f
C3194 VDDA.n453 GNDA 0.043516f
C3195 VDDA.n454 GNDA 0.038833f
C3196 VDDA.n455 GNDA 0.015937f
C3197 VDDA.n456 GNDA 0.056257f
C3198 VDDA.n457 GNDA 0.038833f
C3199 VDDA.n458 GNDA 0.042364f
C3200 VDDA.n459 GNDA 0.02578f
C3201 VDDA.n460 GNDA 0.034927f
C3202 VDDA.n461 GNDA 0.159603f
C3203 VDDA.t350 GNDA 0.191981f
C3204 VDDA.t246 GNDA 0.115958f
C3205 VDDA.t211 GNDA 0.079062f
C3206 VDDA.n462 GNDA 0.02899f
C3207 VDDA.n463 GNDA 0.036896f
C3208 VDDA.t161 GNDA 0.086969f
C3209 VDDA.t223 GNDA 0.115958f
C3210 VDDA.t422 GNDA 0.191981f
C3211 VDDA.n464 GNDA 0.160581f
C3212 VDDA.n465 GNDA 0.035905f
C3213 VDDA.n466 GNDA 0.02578f
C3214 VDDA.t421 GNDA 0.012582f
C3215 VDDA.n467 GNDA 0.042364f
C3216 VDDA.n468 GNDA 0.129197f
C3217 VDDA.n469 GNDA 0.150831f
C3218 VDDA.n470 GNDA 0.480271f
C3219 two_stage_opamp_dummy_magic_0.Vb3.t5 GNDA 0.012871f
C3220 two_stage_opamp_dummy_magic_0.Vb3.t3 GNDA 0.012871f
C3221 two_stage_opamp_dummy_magic_0.Vb3.n0 GNDA 0.041459f
C3222 two_stage_opamp_dummy_magic_0.Vb3.t7 GNDA 0.012871f
C3223 two_stage_opamp_dummy_magic_0.Vb3.t0 GNDA 0.012871f
C3224 two_stage_opamp_dummy_magic_0.Vb3.n1 GNDA 0.04146f
C3225 two_stage_opamp_dummy_magic_0.Vb3.n2 GNDA 0.228564f
C3226 two_stage_opamp_dummy_magic_0.Vb3.t4 GNDA 0.012871f
C3227 two_stage_opamp_dummy_magic_0.Vb3.t6 GNDA 0.012871f
C3228 two_stage_opamp_dummy_magic_0.Vb3.n3 GNDA 0.038876f
C3229 two_stage_opamp_dummy_magic_0.Vb3.n4 GNDA 0.692281f
C3230 two_stage_opamp_dummy_magic_0.Vb3.t2 GNDA 0.046336f
C3231 two_stage_opamp_dummy_magic_0.Vb3.t1 GNDA 0.046336f
C3232 two_stage_opamp_dummy_magic_0.Vb3.n5 GNDA 0.167927f
C3233 two_stage_opamp_dummy_magic_0.Vb3.t22 GNDA 0.079878f
C3234 two_stage_opamp_dummy_magic_0.Vb3.t8 GNDA 0.063713f
C3235 two_stage_opamp_dummy_magic_0.Vb3.t13 GNDA 0.063713f
C3236 two_stage_opamp_dummy_magic_0.Vb3.t10 GNDA 0.063713f
C3237 two_stage_opamp_dummy_magic_0.Vb3.t16 GNDA 0.063713f
C3238 two_stage_opamp_dummy_magic_0.Vb3.t20 GNDA 0.073524f
C3239 two_stage_opamp_dummy_magic_0.Vb3.n6 GNDA 0.059693f
C3240 two_stage_opamp_dummy_magic_0.Vb3.n7 GNDA 0.036683f
C3241 two_stage_opamp_dummy_magic_0.Vb3.n8 GNDA 0.036683f
C3242 two_stage_opamp_dummy_magic_0.Vb3.n9 GNDA 0.034349f
C3243 two_stage_opamp_dummy_magic_0.Vb3.t28 GNDA 0.063713f
C3244 two_stage_opamp_dummy_magic_0.Vb3.t26 GNDA 0.063713f
C3245 two_stage_opamp_dummy_magic_0.Vb3.t15 GNDA 0.063713f
C3246 two_stage_opamp_dummy_magic_0.Vb3.t17 GNDA 0.063713f
C3247 two_stage_opamp_dummy_magic_0.Vb3.t11 GNDA 0.073524f
C3248 two_stage_opamp_dummy_magic_0.Vb3.n10 GNDA 0.059693f
C3249 two_stage_opamp_dummy_magic_0.Vb3.n11 GNDA 0.036683f
C3250 two_stage_opamp_dummy_magic_0.Vb3.n12 GNDA 0.036683f
C3251 two_stage_opamp_dummy_magic_0.Vb3.n13 GNDA 0.034349f
C3252 two_stage_opamp_dummy_magic_0.Vb3.n14 GNDA 0.035386f
C3253 two_stage_opamp_dummy_magic_0.Vb3.t9 GNDA 0.063713f
C3254 two_stage_opamp_dummy_magic_0.Vb3.t14 GNDA 0.063713f
C3255 two_stage_opamp_dummy_magic_0.Vb3.t19 GNDA 0.063713f
C3256 two_stage_opamp_dummy_magic_0.Vb3.t23 GNDA 0.063713f
C3257 two_stage_opamp_dummy_magic_0.Vb3.t25 GNDA 0.073524f
C3258 two_stage_opamp_dummy_magic_0.Vb3.n15 GNDA 0.059693f
C3259 two_stage_opamp_dummy_magic_0.Vb3.n16 GNDA 0.036683f
C3260 two_stage_opamp_dummy_magic_0.Vb3.n17 GNDA 0.036683f
C3261 two_stage_opamp_dummy_magic_0.Vb3.n18 GNDA 0.034349f
C3262 two_stage_opamp_dummy_magic_0.Vb3.t27 GNDA 0.063713f
C3263 two_stage_opamp_dummy_magic_0.Vb3.t24 GNDA 0.063713f
C3264 two_stage_opamp_dummy_magic_0.Vb3.t21 GNDA 0.063713f
C3265 two_stage_opamp_dummy_magic_0.Vb3.t18 GNDA 0.063713f
C3266 two_stage_opamp_dummy_magic_0.Vb3.t12 GNDA 0.073524f
C3267 two_stage_opamp_dummy_magic_0.Vb3.n19 GNDA 0.059693f
C3268 two_stage_opamp_dummy_magic_0.Vb3.n20 GNDA 0.036683f
C3269 two_stage_opamp_dummy_magic_0.Vb3.n21 GNDA 0.036683f
C3270 two_stage_opamp_dummy_magic_0.Vb3.n22 GNDA 0.034349f
C3271 two_stage_opamp_dummy_magic_0.Vb3.n23 GNDA 0.03722f
C3272 two_stage_opamp_dummy_magic_0.Vb3.n24 GNDA 1.01054f
C3273 two_stage_opamp_dummy_magic_0.Vb3.n25 GNDA 0.247796f
C3274 two_stage_opamp_dummy_magic_0.Vb3.n26 GNDA 0.80646f
C3275 bgr_0.VB3_CUR_BIAS GNDA 1.31912f
C3276 bgr_0.NFET_GATE_10uA.t0 GNDA 0.01496f
C3277 bgr_0.NFET_GATE_10uA.t2 GNDA 0.01496f
C3278 bgr_0.NFET_GATE_10uA.n0 GNDA 0.042091f
C3279 bgr_0.NFET_GATE_10uA.t18 GNDA 0.014586f
C3280 bgr_0.NFET_GATE_10uA.t6 GNDA 0.014586f
C3281 bgr_0.NFET_GATE_10uA.t14 GNDA 0.014586f
C3282 bgr_0.NFET_GATE_10uA.t19 GNDA 0.014586f
C3283 bgr_0.NFET_GATE_10uA.t5 GNDA 0.014586f
C3284 bgr_0.NFET_GATE_10uA.t13 GNDA 0.014586f
C3285 bgr_0.NFET_GATE_10uA.t12 GNDA 0.021563f
C3286 bgr_0.NFET_GATE_10uA.n1 GNDA 0.026685f
C3287 bgr_0.NFET_GATE_10uA.n2 GNDA 0.019075f
C3288 bgr_0.NFET_GATE_10uA.n3 GNDA 0.016149f
C3289 bgr_0.NFET_GATE_10uA.t15 GNDA 0.014586f
C3290 bgr_0.NFET_GATE_10uA.t8 GNDA 0.014586f
C3291 bgr_0.NFET_GATE_10uA.t21 GNDA 0.014586f
C3292 bgr_0.NFET_GATE_10uA.t16 GNDA 0.021563f
C3293 bgr_0.NFET_GATE_10uA.n4 GNDA 0.026685f
C3294 bgr_0.NFET_GATE_10uA.n5 GNDA 0.019075f
C3295 bgr_0.NFET_GATE_10uA.n6 GNDA 0.016149f
C3296 bgr_0.NFET_GATE_10uA.t20 GNDA 0.014586f
C3297 bgr_0.NFET_GATE_10uA.t7 GNDA 0.021563f
C3298 bgr_0.NFET_GATE_10uA.n7 GNDA 0.02376f
C3299 bgr_0.NFET_GATE_10uA.n8 GNDA 0.026114f
C3300 bgr_0.NFET_GATE_10uA.t11 GNDA 0.014586f
C3301 bgr_0.NFET_GATE_10uA.t22 GNDA 0.021563f
C3302 bgr_0.NFET_GATE_10uA.n9 GNDA 0.02376f
C3303 bgr_0.NFET_GATE_10uA.t9 GNDA 0.014586f
C3304 bgr_0.NFET_GATE_10uA.t17 GNDA 0.014586f
C3305 bgr_0.NFET_GATE_10uA.t23 GNDA 0.014586f
C3306 bgr_0.NFET_GATE_10uA.t10 GNDA 0.021563f
C3307 bgr_0.NFET_GATE_10uA.n10 GNDA 0.026685f
C3308 bgr_0.NFET_GATE_10uA.n11 GNDA 0.019075f
C3309 bgr_0.NFET_GATE_10uA.n12 GNDA 0.016149f
C3310 bgr_0.NFET_GATE_10uA.n13 GNDA 0.026114f
C3311 bgr_0.NFET_GATE_10uA.n14 GNDA 0.605807f
C3312 bgr_0.NFET_GATE_10uA.n15 GNDA 0.022264f
C3313 bgr_0.NFET_GATE_10uA.n16 GNDA 0.016149f
C3314 bgr_0.NFET_GATE_10uA.n17 GNDA 0.019075f
C3315 bgr_0.NFET_GATE_10uA.n18 GNDA 0.026685f
C3316 bgr_0.NFET_GATE_10uA.t1 GNDA 0.034164f
C3317 bgr_0.NFET_GATE_10uA.n19 GNDA 0.327308f
C3318 bgr_0.NFET_GATE_10uA.t3 GNDA 0.01496f
C3319 bgr_0.NFET_GATE_10uA.t4 GNDA 0.01496f
C3320 bgr_0.NFET_GATE_10uA.n20 GNDA 0.088541f
.ends

