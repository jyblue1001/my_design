magic
tech sky130A
timestamp 1751975008
<< metal1 >>
rect 2960 6685 3000 6690
rect 2960 6655 2965 6685
rect 2995 6655 3000 6685
rect 2960 6650 3000 6655
rect 3030 6685 3070 6690
rect 3030 6655 3035 6685
rect 3065 6655 3070 6685
rect 6060 6685 6100 6690
rect 6060 6655 6065 6685
rect 6095 6655 6100 6685
rect 3030 6650 3070 6655
rect 2915 6580 2955 6585
rect 2915 6550 2920 6580
rect 2950 6550 2955 6580
rect 2915 6545 2955 6550
rect 2925 2710 2945 6545
rect 2970 2520 2990 6650
rect 3280 6525 3300 6650
rect 3400 6645 3440 6650
rect 3400 6615 3405 6645
rect 3435 6615 3440 6645
rect 3400 6610 3440 6615
rect 3270 6520 3310 6525
rect 3270 6490 3275 6520
rect 3305 6490 3310 6520
rect 3270 6485 3310 6490
rect 3555 6480 3575 6655
rect 4010 6645 4050 6650
rect 4010 6615 4015 6645
rect 4045 6615 4050 6645
rect 4010 6610 4050 6615
rect 3545 6475 3585 6480
rect 3545 6445 3550 6475
rect 3580 6445 3585 6475
rect 3545 6440 3585 6445
rect 3975 6475 4005 6480
rect 3975 6440 4005 6445
rect 3985 2790 4005 6440
rect 4020 3365 4040 6610
rect 4340 6585 4360 6655
rect 4330 6580 4370 6585
rect 4330 6550 4335 6580
rect 4365 6550 4370 6580
rect 4330 6545 4370 6550
rect 5085 5495 5105 6655
rect 5730 6585 5750 6655
rect 6060 6650 6100 6655
rect 6700 6685 6740 6690
rect 6700 6655 6705 6685
rect 6735 6655 6740 6685
rect 7020 6685 7060 6690
rect 7020 6655 7025 6685
rect 7055 6655 7060 6685
rect 6700 6650 6740 6655
rect 5720 6580 5760 6585
rect 5720 6550 5725 6580
rect 5755 6550 5760 6580
rect 5720 6545 5760 6550
rect 5375 6520 5415 6525
rect 5375 6490 5380 6520
rect 5410 6490 5415 6520
rect 5375 6485 5415 6490
rect 5065 5490 5105 5495
rect 4770 5470 4810 5475
rect 4770 5440 4775 5470
rect 4805 5440 4810 5470
rect 5065 5460 5070 5490
rect 5100 5460 5105 5490
rect 5065 5455 5105 5460
rect 4770 5435 4810 5440
rect 4780 4805 4800 5435
rect 5385 4950 5405 6485
rect 5375 4945 5415 4950
rect 5375 4915 5380 4945
rect 5410 4915 5415 4945
rect 5375 4910 5415 4915
rect 4770 4800 4810 4805
rect 4770 4770 4775 4800
rect 4805 4770 4810 4800
rect 4770 4765 4810 4770
rect 5025 4800 5065 4805
rect 5025 4770 5030 4800
rect 5060 4770 5065 4800
rect 5025 4765 5065 4770
rect 5035 4075 5055 4765
rect 5025 4070 5065 4075
rect 5025 4040 5030 4070
rect 5060 4040 5065 4070
rect 5025 4035 5065 4040
rect 5970 4070 6010 4075
rect 5970 4040 5975 4070
rect 6005 4040 6010 4070
rect 5970 4035 6010 4040
rect 4995 3665 5035 3670
rect 4995 3635 5000 3665
rect 5030 3635 5035 3665
rect 4995 3630 5035 3635
rect 4020 3360 4060 3365
rect 4020 3330 4025 3360
rect 4055 3330 4060 3360
rect 4020 3325 4060 3330
rect 5005 3305 5025 3630
rect 4995 3300 5035 3305
rect 4995 3270 5000 3300
rect 5030 3270 5035 3300
rect 4995 3265 5035 3270
rect 5980 2410 6000 4035
rect 6070 3670 6090 6650
rect 6785 5090 6805 6655
rect 7020 6650 7060 6655
rect 7090 6685 7130 6690
rect 7090 6655 7095 6685
rect 7125 6655 7130 6685
rect 7090 6650 7130 6655
rect 6410 5085 6450 5090
rect 6410 5055 6415 5085
rect 6445 5055 6450 5085
rect 6410 5050 6450 5055
rect 6775 5085 6815 5090
rect 6775 5055 6780 5085
rect 6810 5055 6815 5085
rect 6775 5050 6815 5055
rect 6420 4850 6440 5050
rect 6410 4845 6450 4850
rect 6410 4815 6415 4845
rect 6445 4815 6450 4845
rect 6410 4810 6450 4815
rect 6060 3665 6100 3670
rect 6060 3635 6065 3665
rect 6095 3635 6100 3665
rect 6060 3630 6100 3635
rect 7100 2520 7120 6650
rect 7135 6580 7175 6585
rect 7135 6550 7140 6580
rect 7170 6550 7175 6580
rect 7135 6545 7175 6550
rect 7145 2710 7165 6545
rect 5970 2405 6010 2410
rect 5970 2375 5975 2405
rect 6005 2375 6010 2405
rect 5970 2370 6010 2375
rect 2440 1790 2480 1830
rect 7610 1790 7650 1830
<< via1 >>
rect 2965 6655 2995 6685
rect 3035 6655 3065 6685
rect 6065 6655 6095 6685
rect 2920 6550 2950 6580
rect 3405 6615 3435 6645
rect 3275 6490 3305 6520
rect 4015 6615 4045 6645
rect 3550 6445 3580 6475
rect 3975 6445 4005 6475
rect 4335 6550 4365 6580
rect 6705 6655 6735 6685
rect 7025 6655 7055 6685
rect 5725 6550 5755 6580
rect 5380 6490 5410 6520
rect 4775 5440 4805 5470
rect 5070 5460 5100 5490
rect 5380 4915 5410 4945
rect 4775 4770 4805 4800
rect 5030 4770 5060 4800
rect 5030 4040 5060 4070
rect 5975 4040 6005 4070
rect 5000 3635 5030 3665
rect 4025 3330 4055 3360
rect 5000 3270 5030 3300
rect 7095 6655 7125 6685
rect 6415 5055 6445 5085
rect 6780 5055 6810 5085
rect 6415 4815 6445 4845
rect 6065 3635 6095 3665
rect 7140 6550 7170 6580
rect 5975 2375 6005 2405
<< metal2 >>
rect 2960 6685 3000 6690
rect 2960 6655 2965 6685
rect 2995 6680 3000 6685
rect 3030 6685 3070 6690
rect 3030 6680 3035 6685
rect 2995 6660 3035 6680
rect 2995 6655 3000 6660
rect 2960 6650 3000 6655
rect 3030 6655 3035 6660
rect 3065 6655 3070 6685
rect 3030 6650 3070 6655
rect 6060 6685 6100 6690
rect 6060 6655 6065 6685
rect 6095 6680 6100 6685
rect 6700 6685 6740 6690
rect 6700 6680 6705 6685
rect 6095 6660 6705 6680
rect 6095 6655 6100 6660
rect 6060 6650 6100 6655
rect 6700 6655 6705 6660
rect 6735 6655 6740 6685
rect 6700 6650 6740 6655
rect 7020 6685 7060 6690
rect 7020 6655 7025 6685
rect 7055 6680 7060 6685
rect 7090 6685 7130 6690
rect 7090 6680 7095 6685
rect 7055 6660 7095 6680
rect 7055 6655 7060 6660
rect 7020 6650 7060 6655
rect 7090 6655 7095 6660
rect 7125 6655 7130 6685
rect 7090 6650 7130 6655
rect 3400 6645 3440 6650
rect 3400 6615 3405 6645
rect 3435 6640 3440 6645
rect 4010 6645 4050 6650
rect 4010 6640 4015 6645
rect 3435 6620 4015 6640
rect 3435 6615 3440 6620
rect 3400 6610 3440 6615
rect 4010 6615 4015 6620
rect 4045 6615 4050 6645
rect 4010 6610 4050 6615
rect 2915 6580 2955 6585
rect 2915 6550 2920 6580
rect 2950 6575 2955 6580
rect 4330 6580 4370 6585
rect 4330 6575 4335 6580
rect 2950 6555 4335 6575
rect 2950 6550 2955 6555
rect 2915 6545 2955 6550
rect 4330 6550 4335 6555
rect 4365 6550 4370 6580
rect 4330 6545 4370 6550
rect 5720 6580 5760 6585
rect 5720 6550 5725 6580
rect 5755 6575 5760 6580
rect 7135 6580 7175 6585
rect 7135 6575 7140 6580
rect 5755 6555 7140 6575
rect 5755 6550 5760 6555
rect 5720 6545 5760 6550
rect 7135 6550 7140 6555
rect 7170 6550 7175 6580
rect 7135 6545 7175 6550
rect 3270 6520 3310 6525
rect 3270 6490 3275 6520
rect 3305 6515 3310 6520
rect 5375 6520 5415 6525
rect 5375 6515 5380 6520
rect 3305 6495 5380 6515
rect 3305 6490 3310 6495
rect 3270 6485 3310 6490
rect 5375 6490 5380 6495
rect 5410 6490 5415 6520
rect 5375 6485 5415 6490
rect 3545 6475 3585 6480
rect 3545 6445 3550 6475
rect 3580 6470 3585 6475
rect 3975 6475 4005 6480
rect 3580 6450 3975 6470
rect 3580 6445 3585 6450
rect 3545 6440 3585 6445
rect 3975 6440 4005 6445
rect 5065 5490 5105 5495
rect 5065 5475 5070 5490
rect 4770 5470 5070 5475
rect 4770 5440 4775 5470
rect 4805 5460 5070 5470
rect 5100 5460 5105 5490
rect 4805 5455 5105 5460
rect 4805 5440 4810 5455
rect 4770 5435 4810 5440
rect 6410 5085 6450 5090
rect 6410 5055 6415 5085
rect 6445 5080 6450 5085
rect 6775 5085 6815 5090
rect 6775 5080 6780 5085
rect 6445 5060 6780 5080
rect 6445 5055 6450 5060
rect 6410 5050 6450 5055
rect 6775 5055 6780 5060
rect 6810 5055 6815 5085
rect 6775 5050 6815 5055
rect 5375 4945 5415 4950
rect 5375 4915 5380 4945
rect 5410 4915 5415 4945
rect 5375 4910 5415 4915
rect 6410 4845 6450 4850
rect 6410 4840 6415 4845
rect 5750 4820 6415 4840
rect 6410 4815 6415 4820
rect 6445 4815 6450 4845
rect 6410 4810 6450 4815
rect 4770 4800 4810 4805
rect 4770 4770 4775 4800
rect 4805 4795 4810 4800
rect 5025 4800 5065 4805
rect 5025 4795 5030 4800
rect 4805 4775 5030 4795
rect 4805 4770 4810 4775
rect 4770 4765 4810 4770
rect 5025 4770 5030 4775
rect 5060 4770 5065 4800
rect 5025 4765 5065 4770
rect 5025 4070 5065 4075
rect 5025 4040 5030 4070
rect 5060 4065 5065 4070
rect 5970 4070 6010 4075
rect 5970 4065 5975 4070
rect 5060 4045 5975 4065
rect 5060 4040 5065 4045
rect 5025 4035 5065 4040
rect 5970 4040 5975 4045
rect 6005 4040 6010 4070
rect 5970 4035 6010 4040
rect 4995 3665 5035 3670
rect 4995 3635 5000 3665
rect 5030 3660 5035 3665
rect 6060 3665 6100 3670
rect 6060 3660 6065 3665
rect 5030 3640 6065 3660
rect 5030 3635 5035 3640
rect 4995 3630 5035 3635
rect 6060 3635 6065 3640
rect 6095 3635 6100 3665
rect 6060 3630 6100 3635
rect 4020 3360 4060 3365
rect 4020 3330 4025 3360
rect 4055 3355 4060 3360
rect 4055 3335 4100 3355
rect 4055 3330 4060 3335
rect 4020 3325 4060 3330
rect 4995 3300 5035 3305
rect 4995 3295 5000 3300
rect 4860 3275 5000 3295
rect 4995 3270 5000 3275
rect 5030 3270 5035 3300
rect 4995 3265 5035 3270
rect 5970 2405 6010 2410
rect 5970 2400 5975 2405
rect 5125 2380 5975 2400
rect 5970 2375 5975 2380
rect 6005 2375 6010 2405
rect 5970 2370 6010 2375
rect 4090 2290 4105 2310
rect 4090 2070 4105 2090
rect 2440 1790 2480 1830
rect 7610 1790 7650 1830
<< metal4 >>
rect 3475 14415 3525 14465
rect 940 6700 990 6750
rect 975 0 1025 50
use bgr  bgr_0
timestamp 1751960357
transform -1 0 22845 0 -1 8250
box 15505 -6295 20095 1600
use two_stage_opamp_dummy_magic  two_stage_opamp_dummy_magic_0
timestamp 1751965702
transform 1 0 -51855 0 1 555
box 51855 -555 61545 6195
<< labels >>
flabel metal4 965 6750 965 6750 1 FreeSans 800 0 0 400 VDDA
port 1 n
flabel metal4 1000 0 1000 0 5 FreeSans 800 0 0 -400 GNDA
port 2 s
flabel metal2 4090 2300 4090 2300 7 FreeSans 400 0 -200 0 VIN-
port 6 w
flabel metal2 4090 2080 4090 2080 7 FreeSans 400 0 -200 0 VIN+
port 5 w
flabel metal2 2460 1790 2460 1790 5 FreeSans 400 0 0 -200 VOUT-
port 4 s
flabel metal2 7630 1790 7630 1790 5 FreeSans 400 0 0 -200 VOUT+
port 3 s
flabel metal4 3500 14415 3500 14415 5 FreeSans 800 0 0 -400 GNDA
port 2 s
<< end >>
