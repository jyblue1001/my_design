** sch_path: /foss/designs/my_design/projects/ASU/EEE572/schematic/tb_buck_converter.sch
**.subckt tb_buck_converter
V1 net2 net4 25
R48 net3 net4 1 m=1
D1 net4 net1 D1N914 area=1
L1 net3 net1 30u m=1
C1 net5 net4 250u m=1
R1 net3 net5 0.05 m=1
V2 net6 GND pulse(0 1.8 0ns 1ns 1ns 24ns 50ns)
S1 net2 net1 net6 GND SW1
**** begin user architecture code



.options method=gear
.options wnflag=1
.options savecurrents


.model D1N914 D(Is=168.1E-21 N=1 Rs=.1 Ikf=0 Xti=3 Eg=1.11 Cjo=4p M=.3333 + Vj=.75 Fc=.5 Bv=100 Ibv=100u Tt=11.54n)


.control
  save all
  * dc V1 0.0 2.0 0.005
  tran 1ps 1us
  remzerovec
  write tb_buck_converter.raw
  set appendwrite

.endc




**** end user architecture code
**.ends
.GLOBAL GND
**** begin user architecture code
.MODEL SW1 SW( VT=0.9 VH=0.01 RON=0.01 ROFF=10G )
**** end user architecture code
.end
