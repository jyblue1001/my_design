magic
tech sky130A
timestamp 1754032204
<< nwell >>
rect 56025 4510 56365 4900
rect 56495 4510 56835 4730
rect 56965 4510 57305 4900
rect 57435 4510 57775 4900
rect 54780 3395 55665 3785
rect 55945 3395 56825 3785
rect 56975 3395 57855 3785
rect 58350 3395 59230 3785
rect 54680 2285 55500 2925
rect 56450 2640 57350 2930
rect 58380 2285 59200 2925
rect 58875 2280 59015 2285
rect 54680 1410 55500 1650
rect 58380 1410 59200 1650
<< nmos >>
rect 56810 2065 56825 2315
rect 56865 2065 56880 2315
rect 56920 2065 56935 2315
rect 56975 2065 56990 2315
rect 56070 1495 56085 1645
rect 56125 1495 56140 1645
rect 56180 1495 56195 1645
rect 56235 1495 56250 1645
rect 56290 1495 56305 1645
rect 56345 1495 56360 1645
rect 56400 1495 56415 1645
rect 56455 1495 56470 1645
rect 56510 1495 56525 1645
rect 56565 1495 56580 1645
rect 56620 1495 56635 1645
rect 56675 1495 56690 1645
rect 57110 1495 57125 1645
rect 57165 1495 57180 1645
rect 57220 1495 57235 1645
rect 57275 1495 57290 1645
rect 57330 1495 57345 1645
rect 57385 1495 57400 1645
rect 57440 1495 57455 1645
rect 57495 1495 57510 1645
rect 57550 1495 57565 1645
rect 57605 1495 57620 1645
rect 57660 1495 57675 1645
rect 57715 1495 57730 1645
rect 54780 890 54795 1190
rect 54835 890 54850 1190
rect 54890 890 54905 1190
rect 54945 890 54960 1190
rect 55000 890 55015 1190
rect 55055 890 55070 1190
rect 55110 890 55125 1190
rect 55165 890 55180 1190
rect 55220 890 55235 1190
rect 55275 890 55290 1190
rect 55330 890 55345 1190
rect 55385 890 55400 1190
rect 56070 820 56085 970
rect 56125 820 56140 970
rect 56180 820 56195 970
rect 56235 820 56250 970
rect 56290 820 56305 970
rect 56345 820 56360 970
rect 56400 820 56415 970
rect 56455 820 56470 970
rect 56510 820 56525 970
rect 56565 820 56580 970
rect 56620 820 56635 970
rect 56675 820 56690 970
rect 56810 820 56825 970
rect 56865 820 56880 970
rect 56920 820 56935 970
rect 56975 820 56990 970
rect 57110 820 57125 970
rect 57165 820 57180 970
rect 57220 820 57235 970
rect 57275 820 57290 970
rect 57330 820 57345 970
rect 57385 820 57400 970
rect 57440 820 57455 970
rect 57495 820 57510 970
rect 57550 820 57565 970
rect 57605 820 57620 970
rect 57660 820 57675 970
rect 57715 820 57730 970
rect 58480 890 58495 1190
rect 58535 890 58550 1190
rect 58590 890 58605 1190
rect 58645 890 58660 1190
rect 58700 890 58715 1190
rect 58755 890 58770 1190
rect 58810 890 58825 1190
rect 58865 890 58880 1190
rect 58920 890 58935 1190
rect 58975 890 58990 1190
rect 59030 890 59045 1190
rect 59085 890 59100 1190
rect 54790 -520 54850 180
rect 54890 -520 54950 180
rect 54990 -520 55050 180
rect 55090 -520 55150 180
rect 55190 -520 55250 180
rect 55290 -520 55350 180
rect 56260 80 56275 330
rect 56315 80 56330 330
rect 56370 80 56385 330
rect 56425 80 56440 330
rect 56480 80 56495 330
rect 56535 80 56550 330
rect 56590 80 56605 330
rect 56645 80 56660 330
rect 56700 80 56715 330
rect 56755 80 56770 330
rect 56810 80 56825 330
rect 56865 80 56880 330
rect 56920 80 56935 330
rect 56975 80 56990 330
rect 57030 80 57045 330
rect 57085 80 57100 330
rect 57140 80 57155 330
rect 57195 80 57210 330
rect 57250 80 57265 330
rect 57305 80 57320 330
rect 57360 80 57375 330
rect 57415 80 57430 330
rect 57470 80 57485 330
rect 56470 -475 56485 -325
rect 56525 -475 56540 -325
rect 56580 -475 56595 -325
rect 56635 -475 56650 -325
rect 56690 -475 56705 -325
rect 56745 -475 56760 -325
rect 56910 -475 57210 -325
rect 58370 -520 58430 180
rect 58470 -520 58530 180
rect 58570 -520 58630 180
rect 58670 -520 58730 180
rect 58770 -520 58830 180
rect 58870 -520 58930 180
<< pmos >>
rect 56125 4530 56145 4880
rect 56185 4530 56205 4880
rect 56245 4530 56265 4880
rect 56595 4530 56615 4710
rect 56655 4530 56675 4710
rect 56715 4530 56735 4710
rect 57065 4530 57085 4880
rect 57125 4530 57145 4880
rect 57185 4530 57205 4880
rect 57535 4530 57555 4880
rect 57595 4530 57615 4880
rect 57655 4530 57675 4880
rect 54880 3415 54900 3765
rect 54940 3415 54960 3765
rect 55000 3415 55020 3765
rect 55060 3415 55080 3765
rect 55120 3415 55140 3765
rect 55180 3415 55200 3765
rect 55240 3415 55260 3765
rect 55300 3415 55320 3765
rect 55360 3415 55380 3765
rect 55420 3415 55440 3765
rect 55480 3415 55500 3765
rect 55540 3415 55560 3765
rect 56045 3415 56065 3765
rect 56105 3415 56125 3765
rect 56165 3415 56185 3765
rect 56225 3415 56245 3765
rect 56285 3415 56305 3765
rect 56345 3415 56365 3765
rect 56405 3415 56425 3765
rect 56465 3415 56485 3765
rect 56525 3415 56545 3765
rect 56585 3415 56605 3765
rect 56645 3415 56665 3765
rect 56705 3415 56725 3765
rect 57075 3415 57095 3765
rect 57135 3415 57155 3765
rect 57195 3415 57215 3765
rect 57255 3415 57275 3765
rect 57315 3415 57335 3765
rect 57375 3415 57395 3765
rect 57435 3415 57455 3765
rect 57495 3415 57515 3765
rect 57555 3415 57575 3765
rect 57615 3415 57635 3765
rect 57675 3415 57695 3765
rect 57735 3415 57755 3765
rect 58450 3415 58470 3765
rect 58510 3415 58530 3765
rect 58570 3415 58590 3765
rect 58630 3415 58650 3765
rect 58690 3415 58710 3765
rect 58750 3415 58770 3765
rect 58810 3415 58830 3765
rect 58870 3415 58890 3765
rect 58930 3415 58950 3765
rect 58990 3415 59010 3765
rect 59050 3415 59070 3765
rect 59110 3415 59130 3765
rect 54780 2305 54795 2905
rect 54835 2305 54850 2905
rect 54890 2305 54905 2905
rect 54945 2305 54960 2905
rect 55000 2305 55015 2905
rect 55055 2305 55070 2905
rect 55110 2305 55125 2905
rect 55165 2305 55180 2905
rect 55220 2305 55235 2905
rect 55275 2305 55290 2905
rect 55330 2305 55345 2905
rect 55385 2305 55400 2905
rect 56550 2660 56565 2910
rect 56605 2660 56620 2910
rect 56660 2660 56675 2910
rect 56715 2660 56730 2910
rect 56770 2660 56785 2910
rect 56825 2660 56840 2910
rect 56960 2660 56975 2910
rect 57015 2660 57030 2910
rect 57070 2660 57085 2910
rect 57125 2660 57140 2910
rect 57180 2660 57195 2910
rect 57235 2660 57250 2910
rect 58480 2305 58495 2905
rect 58535 2305 58550 2905
rect 58590 2305 58605 2905
rect 58645 2305 58660 2905
rect 58700 2305 58715 2905
rect 58755 2305 58770 2905
rect 58810 2305 58825 2905
rect 58865 2305 58880 2905
rect 58920 2305 58935 2905
rect 58975 2305 58990 2905
rect 59030 2305 59045 2905
rect 59085 2305 59100 2905
rect 54780 1430 54795 1630
rect 54835 1430 54850 1630
rect 54890 1430 54905 1630
rect 54945 1430 54960 1630
rect 55000 1430 55015 1630
rect 55055 1430 55070 1630
rect 55110 1430 55125 1630
rect 55165 1430 55180 1630
rect 55220 1430 55235 1630
rect 55275 1430 55290 1630
rect 55330 1430 55345 1630
rect 55385 1430 55400 1630
rect 58480 1430 58495 1630
rect 58535 1430 58550 1630
rect 58590 1430 58605 1630
rect 58645 1430 58660 1630
rect 58700 1430 58715 1630
rect 58755 1430 58770 1630
rect 58810 1430 58825 1630
rect 58865 1430 58880 1630
rect 58920 1430 58935 1630
rect 58975 1430 58990 1630
rect 59030 1430 59045 1630
rect 59085 1430 59100 1630
<< ndiff >>
rect 56770 2300 56810 2315
rect 56770 2080 56780 2300
rect 56800 2080 56810 2300
rect 56770 2065 56810 2080
rect 56825 2300 56865 2315
rect 56825 2080 56835 2300
rect 56855 2080 56865 2300
rect 56825 2065 56865 2080
rect 56880 2300 56920 2315
rect 56880 2080 56890 2300
rect 56910 2080 56920 2300
rect 56880 2065 56920 2080
rect 56935 2300 56975 2315
rect 56935 2080 56945 2300
rect 56965 2080 56975 2300
rect 56935 2065 56975 2080
rect 56990 2300 57030 2315
rect 56990 2080 57000 2300
rect 57020 2080 57030 2300
rect 56990 2065 57030 2080
rect 56030 1630 56070 1645
rect 56030 1510 56040 1630
rect 56060 1510 56070 1630
rect 56030 1495 56070 1510
rect 56085 1630 56125 1645
rect 56085 1510 56095 1630
rect 56115 1510 56125 1630
rect 56085 1495 56125 1510
rect 56140 1630 56180 1645
rect 56140 1510 56150 1630
rect 56170 1510 56180 1630
rect 56140 1495 56180 1510
rect 56195 1630 56235 1645
rect 56195 1510 56205 1630
rect 56225 1510 56235 1630
rect 56195 1495 56235 1510
rect 56250 1630 56290 1645
rect 56250 1510 56260 1630
rect 56280 1510 56290 1630
rect 56250 1495 56290 1510
rect 56305 1630 56345 1645
rect 56305 1510 56315 1630
rect 56335 1510 56345 1630
rect 56305 1495 56345 1510
rect 56360 1630 56400 1645
rect 56360 1510 56370 1630
rect 56390 1510 56400 1630
rect 56360 1495 56400 1510
rect 56415 1630 56455 1645
rect 56415 1510 56425 1630
rect 56445 1510 56455 1630
rect 56415 1495 56455 1510
rect 56470 1630 56510 1645
rect 56470 1510 56480 1630
rect 56500 1510 56510 1630
rect 56470 1495 56510 1510
rect 56525 1630 56565 1645
rect 56525 1510 56535 1630
rect 56555 1510 56565 1630
rect 56525 1495 56565 1510
rect 56580 1630 56620 1645
rect 56580 1510 56590 1630
rect 56610 1510 56620 1630
rect 56580 1495 56620 1510
rect 56635 1630 56675 1645
rect 56635 1510 56645 1630
rect 56665 1510 56675 1630
rect 56635 1495 56675 1510
rect 56690 1630 56730 1645
rect 56690 1510 56700 1630
rect 56720 1510 56730 1630
rect 56690 1495 56730 1510
rect 57070 1630 57110 1645
rect 57070 1510 57080 1630
rect 57100 1510 57110 1630
rect 57070 1495 57110 1510
rect 57125 1630 57165 1645
rect 57125 1510 57135 1630
rect 57155 1510 57165 1630
rect 57125 1495 57165 1510
rect 57180 1630 57220 1645
rect 57180 1510 57190 1630
rect 57210 1510 57220 1630
rect 57180 1495 57220 1510
rect 57235 1630 57275 1645
rect 57235 1510 57245 1630
rect 57265 1510 57275 1630
rect 57235 1495 57275 1510
rect 57290 1630 57330 1645
rect 57290 1510 57300 1630
rect 57320 1510 57330 1630
rect 57290 1495 57330 1510
rect 57345 1630 57385 1645
rect 57345 1510 57355 1630
rect 57375 1510 57385 1630
rect 57345 1495 57385 1510
rect 57400 1630 57440 1645
rect 57400 1510 57410 1630
rect 57430 1510 57440 1630
rect 57400 1495 57440 1510
rect 57455 1630 57495 1645
rect 57455 1510 57465 1630
rect 57485 1510 57495 1630
rect 57455 1495 57495 1510
rect 57510 1630 57550 1645
rect 57510 1510 57520 1630
rect 57540 1510 57550 1630
rect 57510 1495 57550 1510
rect 57565 1630 57605 1645
rect 57565 1510 57575 1630
rect 57595 1510 57605 1630
rect 57565 1495 57605 1510
rect 57620 1630 57660 1645
rect 57620 1510 57630 1630
rect 57650 1510 57660 1630
rect 57620 1495 57660 1510
rect 57675 1630 57715 1645
rect 57675 1510 57685 1630
rect 57705 1510 57715 1630
rect 57675 1495 57715 1510
rect 57730 1630 57770 1645
rect 57730 1510 57740 1630
rect 57760 1510 57770 1630
rect 57730 1495 57770 1510
rect 54740 1175 54780 1190
rect 54740 905 54750 1175
rect 54770 905 54780 1175
rect 54740 890 54780 905
rect 54795 1175 54835 1190
rect 54795 905 54805 1175
rect 54825 905 54835 1175
rect 54795 890 54835 905
rect 54850 1175 54890 1190
rect 54850 905 54860 1175
rect 54880 905 54890 1175
rect 54850 890 54890 905
rect 54905 1175 54945 1190
rect 54905 905 54915 1175
rect 54935 905 54945 1175
rect 54905 890 54945 905
rect 54960 1175 55000 1190
rect 54960 905 54970 1175
rect 54990 905 55000 1175
rect 54960 890 55000 905
rect 55015 1175 55055 1190
rect 55015 905 55025 1175
rect 55045 905 55055 1175
rect 55015 890 55055 905
rect 55070 1175 55110 1190
rect 55070 905 55080 1175
rect 55100 905 55110 1175
rect 55070 890 55110 905
rect 55125 1175 55165 1190
rect 55125 905 55135 1175
rect 55155 905 55165 1175
rect 55125 890 55165 905
rect 55180 1175 55220 1190
rect 55180 905 55190 1175
rect 55210 905 55220 1175
rect 55180 890 55220 905
rect 55235 1175 55275 1190
rect 55235 905 55245 1175
rect 55265 905 55275 1175
rect 55235 890 55275 905
rect 55290 1175 55330 1190
rect 55290 905 55300 1175
rect 55320 905 55330 1175
rect 55290 890 55330 905
rect 55345 1175 55385 1190
rect 55345 905 55355 1175
rect 55375 905 55385 1175
rect 55345 890 55385 905
rect 55400 1175 55440 1190
rect 55400 905 55410 1175
rect 55430 905 55440 1175
rect 58440 1175 58480 1190
rect 55400 890 55440 905
rect 56030 955 56070 970
rect 56030 835 56040 955
rect 56060 835 56070 955
rect 56030 820 56070 835
rect 56085 955 56125 970
rect 56085 835 56095 955
rect 56115 835 56125 955
rect 56085 820 56125 835
rect 56140 955 56180 970
rect 56140 835 56150 955
rect 56170 835 56180 955
rect 56140 820 56180 835
rect 56195 955 56235 970
rect 56195 835 56205 955
rect 56225 835 56235 955
rect 56195 820 56235 835
rect 56250 955 56290 970
rect 56250 835 56260 955
rect 56280 835 56290 955
rect 56250 820 56290 835
rect 56305 955 56345 970
rect 56305 835 56315 955
rect 56335 835 56345 955
rect 56305 820 56345 835
rect 56360 955 56400 970
rect 56360 835 56370 955
rect 56390 835 56400 955
rect 56360 820 56400 835
rect 56415 955 56455 970
rect 56415 835 56425 955
rect 56445 835 56455 955
rect 56415 820 56455 835
rect 56470 955 56510 970
rect 56470 835 56480 955
rect 56500 835 56510 955
rect 56470 820 56510 835
rect 56525 955 56565 970
rect 56525 835 56535 955
rect 56555 835 56565 955
rect 56525 820 56565 835
rect 56580 955 56620 970
rect 56580 835 56590 955
rect 56610 835 56620 955
rect 56580 820 56620 835
rect 56635 955 56675 970
rect 56635 835 56645 955
rect 56665 835 56675 955
rect 56635 820 56675 835
rect 56690 955 56730 970
rect 56770 955 56810 970
rect 56690 835 56700 955
rect 56720 835 56730 955
rect 56770 835 56780 955
rect 56800 835 56810 955
rect 56690 820 56730 835
rect 56770 820 56810 835
rect 56825 955 56865 970
rect 56825 835 56835 955
rect 56855 835 56865 955
rect 56825 820 56865 835
rect 56880 955 56920 970
rect 56880 835 56890 955
rect 56910 835 56920 955
rect 56880 820 56920 835
rect 56935 955 56975 970
rect 56935 835 56945 955
rect 56965 835 56975 955
rect 56935 820 56975 835
rect 56990 955 57030 970
rect 57070 955 57110 970
rect 56990 835 57000 955
rect 57020 835 57030 955
rect 57070 835 57080 955
rect 57100 835 57110 955
rect 56990 820 57030 835
rect 57070 820 57110 835
rect 57125 955 57165 970
rect 57125 835 57135 955
rect 57155 835 57165 955
rect 57125 820 57165 835
rect 57180 955 57220 970
rect 57180 835 57190 955
rect 57210 835 57220 955
rect 57180 820 57220 835
rect 57235 955 57275 970
rect 57235 835 57245 955
rect 57265 835 57275 955
rect 57235 820 57275 835
rect 57290 955 57330 970
rect 57290 835 57300 955
rect 57320 835 57330 955
rect 57290 820 57330 835
rect 57345 955 57385 970
rect 57345 835 57355 955
rect 57375 835 57385 955
rect 57345 820 57385 835
rect 57400 955 57440 970
rect 57400 835 57410 955
rect 57430 835 57440 955
rect 57400 820 57440 835
rect 57455 955 57495 970
rect 57455 835 57465 955
rect 57485 835 57495 955
rect 57455 820 57495 835
rect 57510 955 57550 970
rect 57510 835 57520 955
rect 57540 835 57550 955
rect 57510 820 57550 835
rect 57565 955 57605 970
rect 57565 835 57575 955
rect 57595 835 57605 955
rect 57565 820 57605 835
rect 57620 955 57660 970
rect 57620 835 57630 955
rect 57650 835 57660 955
rect 57620 820 57660 835
rect 57675 955 57715 970
rect 57675 835 57685 955
rect 57705 835 57715 955
rect 57675 820 57715 835
rect 57730 955 57770 970
rect 57730 835 57740 955
rect 57760 835 57770 955
rect 58440 905 58450 1175
rect 58470 905 58480 1175
rect 58440 890 58480 905
rect 58495 1175 58535 1190
rect 58495 905 58505 1175
rect 58525 905 58535 1175
rect 58495 890 58535 905
rect 58550 1175 58590 1190
rect 58550 905 58560 1175
rect 58580 905 58590 1175
rect 58550 890 58590 905
rect 58605 1175 58645 1190
rect 58605 905 58615 1175
rect 58635 905 58645 1175
rect 58605 890 58645 905
rect 58660 1175 58700 1190
rect 58660 905 58670 1175
rect 58690 905 58700 1175
rect 58660 890 58700 905
rect 58715 1175 58755 1190
rect 58715 905 58725 1175
rect 58745 905 58755 1175
rect 58715 890 58755 905
rect 58770 1175 58810 1190
rect 58770 905 58780 1175
rect 58800 905 58810 1175
rect 58770 890 58810 905
rect 58825 1175 58865 1190
rect 58825 905 58835 1175
rect 58855 905 58865 1175
rect 58825 890 58865 905
rect 58880 1175 58920 1190
rect 58880 905 58890 1175
rect 58910 905 58920 1175
rect 58880 890 58920 905
rect 58935 1175 58975 1190
rect 58935 905 58945 1175
rect 58965 905 58975 1175
rect 58935 890 58975 905
rect 58990 1175 59030 1190
rect 58990 905 59000 1175
rect 59020 905 59030 1175
rect 58990 890 59030 905
rect 59045 1175 59085 1190
rect 59045 905 59055 1175
rect 59075 905 59085 1175
rect 59045 890 59085 905
rect 59100 1175 59140 1190
rect 59100 905 59110 1175
rect 59130 905 59140 1175
rect 59100 890 59140 905
rect 57730 820 57770 835
rect 56220 315 56260 330
rect 54750 165 54790 180
rect 54750 -505 54760 165
rect 54780 -505 54790 165
rect 54750 -520 54790 -505
rect 54850 165 54890 180
rect 54850 -505 54860 165
rect 54880 -505 54890 165
rect 54850 -520 54890 -505
rect 54950 165 54990 180
rect 54950 -505 54960 165
rect 54980 -505 54990 165
rect 54950 -520 54990 -505
rect 55050 165 55090 180
rect 55050 -505 55060 165
rect 55080 -505 55090 165
rect 55050 -520 55090 -505
rect 55150 165 55190 180
rect 55150 -505 55160 165
rect 55180 -505 55190 165
rect 55150 -520 55190 -505
rect 55250 165 55290 180
rect 55250 -505 55260 165
rect 55280 -505 55290 165
rect 55250 -520 55290 -505
rect 55350 165 55390 180
rect 55350 -505 55360 165
rect 55380 -505 55390 165
rect 56220 95 56230 315
rect 56250 95 56260 315
rect 56220 80 56260 95
rect 56275 315 56315 330
rect 56275 95 56285 315
rect 56305 95 56315 315
rect 56275 80 56315 95
rect 56330 315 56370 330
rect 56330 95 56340 315
rect 56360 95 56370 315
rect 56330 80 56370 95
rect 56385 315 56425 330
rect 56385 95 56395 315
rect 56415 95 56425 315
rect 56385 80 56425 95
rect 56440 315 56480 330
rect 56440 95 56450 315
rect 56470 95 56480 315
rect 56440 80 56480 95
rect 56495 315 56535 330
rect 56495 95 56505 315
rect 56525 95 56535 315
rect 56495 80 56535 95
rect 56550 315 56590 330
rect 56550 95 56560 315
rect 56580 95 56590 315
rect 56550 80 56590 95
rect 56605 315 56645 330
rect 56605 95 56615 315
rect 56635 95 56645 315
rect 56605 80 56645 95
rect 56660 315 56700 330
rect 56660 95 56670 315
rect 56690 95 56700 315
rect 56660 80 56700 95
rect 56715 315 56755 330
rect 56715 95 56725 315
rect 56745 95 56755 315
rect 56715 80 56755 95
rect 56770 315 56810 330
rect 56770 95 56780 315
rect 56800 95 56810 315
rect 56770 80 56810 95
rect 56825 315 56865 330
rect 56825 95 56835 315
rect 56855 95 56865 315
rect 56825 80 56865 95
rect 56880 315 56920 330
rect 56880 95 56890 315
rect 56910 95 56920 315
rect 56880 80 56920 95
rect 56935 315 56975 330
rect 56935 95 56945 315
rect 56965 95 56975 315
rect 56935 80 56975 95
rect 56990 315 57030 330
rect 56990 95 57000 315
rect 57020 95 57030 315
rect 56990 80 57030 95
rect 57045 315 57085 330
rect 57045 95 57055 315
rect 57075 95 57085 315
rect 57045 80 57085 95
rect 57100 315 57140 330
rect 57100 95 57110 315
rect 57130 95 57140 315
rect 57100 80 57140 95
rect 57155 315 57195 330
rect 57155 95 57165 315
rect 57185 95 57195 315
rect 57155 80 57195 95
rect 57210 315 57250 330
rect 57210 95 57220 315
rect 57240 95 57250 315
rect 57210 80 57250 95
rect 57265 315 57305 330
rect 57265 95 57275 315
rect 57295 95 57305 315
rect 57265 80 57305 95
rect 57320 315 57360 330
rect 57320 95 57330 315
rect 57350 95 57360 315
rect 57320 80 57360 95
rect 57375 315 57415 330
rect 57375 95 57385 315
rect 57405 95 57415 315
rect 57375 80 57415 95
rect 57430 315 57470 330
rect 57430 95 57440 315
rect 57460 95 57470 315
rect 57430 80 57470 95
rect 57485 315 57525 330
rect 57485 95 57495 315
rect 57515 95 57525 315
rect 57485 80 57525 95
rect 58330 165 58370 180
rect 56430 -340 56470 -325
rect 56430 -460 56440 -340
rect 56460 -460 56470 -340
rect 56430 -475 56470 -460
rect 56485 -340 56525 -325
rect 56485 -460 56495 -340
rect 56515 -460 56525 -340
rect 56485 -475 56525 -460
rect 56540 -340 56580 -325
rect 56540 -460 56550 -340
rect 56570 -460 56580 -340
rect 56540 -475 56580 -460
rect 56595 -340 56635 -325
rect 56595 -460 56605 -340
rect 56625 -460 56635 -340
rect 56595 -475 56635 -460
rect 56650 -340 56690 -325
rect 56650 -460 56660 -340
rect 56680 -460 56690 -340
rect 56650 -475 56690 -460
rect 56705 -340 56745 -325
rect 56705 -460 56715 -340
rect 56735 -460 56745 -340
rect 56705 -475 56745 -460
rect 56760 -340 56800 -325
rect 56760 -460 56770 -340
rect 56790 -460 56800 -340
rect 56760 -475 56800 -460
rect 56870 -340 56910 -325
rect 56870 -460 56880 -340
rect 56900 -460 56910 -340
rect 56870 -475 56910 -460
rect 57210 -340 57250 -325
rect 57210 -460 57220 -340
rect 57240 -460 57250 -340
rect 57210 -475 57250 -460
rect 55350 -520 55390 -505
rect 58330 -505 58340 165
rect 58360 -505 58370 165
rect 58330 -520 58370 -505
rect 58430 165 58470 180
rect 58430 -505 58440 165
rect 58460 -505 58470 165
rect 58430 -520 58470 -505
rect 58530 165 58570 180
rect 58530 -505 58540 165
rect 58560 -505 58570 165
rect 58530 -520 58570 -505
rect 58630 165 58670 180
rect 58630 -505 58640 165
rect 58660 -505 58670 165
rect 58630 -520 58670 -505
rect 58730 165 58770 180
rect 58730 -505 58740 165
rect 58760 -505 58770 165
rect 58730 -520 58770 -505
rect 58830 165 58870 180
rect 58830 -505 58840 165
rect 58860 -505 58870 165
rect 58830 -520 58870 -505
rect 58930 165 58970 180
rect 58930 -505 58940 165
rect 58960 -505 58970 165
rect 58930 -520 58970 -505
<< pdiff >>
rect 56085 4865 56125 4880
rect 56085 4545 56095 4865
rect 56115 4545 56125 4865
rect 56085 4530 56125 4545
rect 56145 4865 56185 4880
rect 56145 4545 56155 4865
rect 56175 4545 56185 4865
rect 56145 4530 56185 4545
rect 56205 4865 56245 4880
rect 56205 4545 56215 4865
rect 56235 4545 56245 4865
rect 56205 4530 56245 4545
rect 56265 4865 56305 4880
rect 56265 4545 56275 4865
rect 56295 4545 56305 4865
rect 57025 4865 57065 4880
rect 56265 4530 56305 4545
rect 56555 4695 56595 4710
rect 56555 4545 56565 4695
rect 56585 4545 56595 4695
rect 56555 4530 56595 4545
rect 56615 4695 56655 4710
rect 56615 4545 56625 4695
rect 56645 4545 56655 4695
rect 56615 4530 56655 4545
rect 56675 4695 56715 4710
rect 56675 4545 56685 4695
rect 56705 4545 56715 4695
rect 56675 4530 56715 4545
rect 56735 4695 56775 4710
rect 56735 4545 56745 4695
rect 56765 4545 56775 4695
rect 56735 4530 56775 4545
rect 57025 4545 57035 4865
rect 57055 4545 57065 4865
rect 57025 4530 57065 4545
rect 57085 4865 57125 4880
rect 57085 4545 57095 4865
rect 57115 4545 57125 4865
rect 57085 4530 57125 4545
rect 57145 4865 57185 4880
rect 57145 4545 57155 4865
rect 57175 4545 57185 4865
rect 57145 4530 57185 4545
rect 57205 4865 57245 4880
rect 57205 4545 57215 4865
rect 57235 4545 57245 4865
rect 57205 4530 57245 4545
rect 57495 4865 57535 4880
rect 57495 4545 57505 4865
rect 57525 4545 57535 4865
rect 57495 4530 57535 4545
rect 57555 4865 57595 4880
rect 57555 4545 57565 4865
rect 57585 4545 57595 4865
rect 57555 4530 57595 4545
rect 57615 4865 57655 4880
rect 57615 4545 57625 4865
rect 57645 4545 57655 4865
rect 57615 4530 57655 4545
rect 57675 4865 57715 4880
rect 57675 4545 57685 4865
rect 57705 4545 57715 4865
rect 57675 4530 57715 4545
rect 54840 3750 54880 3765
rect 54840 3430 54850 3750
rect 54870 3430 54880 3750
rect 54840 3415 54880 3430
rect 54900 3750 54940 3765
rect 54900 3430 54910 3750
rect 54930 3430 54940 3750
rect 54900 3415 54940 3430
rect 54960 3750 55000 3765
rect 54960 3430 54970 3750
rect 54990 3430 55000 3750
rect 54960 3415 55000 3430
rect 55020 3750 55060 3765
rect 55020 3430 55030 3750
rect 55050 3430 55060 3750
rect 55020 3415 55060 3430
rect 55080 3750 55120 3765
rect 55080 3430 55090 3750
rect 55110 3430 55120 3750
rect 55080 3415 55120 3430
rect 55140 3750 55180 3765
rect 55140 3430 55150 3750
rect 55170 3430 55180 3750
rect 55140 3415 55180 3430
rect 55200 3750 55240 3765
rect 55200 3430 55210 3750
rect 55230 3430 55240 3750
rect 55200 3415 55240 3430
rect 55260 3750 55300 3765
rect 55260 3430 55270 3750
rect 55290 3430 55300 3750
rect 55260 3415 55300 3430
rect 55320 3750 55360 3765
rect 55320 3430 55330 3750
rect 55350 3430 55360 3750
rect 55320 3415 55360 3430
rect 55380 3750 55420 3765
rect 55380 3430 55390 3750
rect 55410 3430 55420 3750
rect 55380 3415 55420 3430
rect 55440 3750 55480 3765
rect 55440 3430 55450 3750
rect 55470 3430 55480 3750
rect 55440 3415 55480 3430
rect 55500 3750 55540 3765
rect 55500 3430 55510 3750
rect 55530 3430 55540 3750
rect 55500 3415 55540 3430
rect 55560 3750 55600 3765
rect 55560 3430 55570 3750
rect 55590 3430 55600 3750
rect 55560 3415 55600 3430
rect 56005 3750 56045 3765
rect 56005 3430 56015 3750
rect 56035 3430 56045 3750
rect 56005 3415 56045 3430
rect 56065 3750 56105 3765
rect 56065 3430 56075 3750
rect 56095 3430 56105 3750
rect 56065 3415 56105 3430
rect 56125 3750 56165 3765
rect 56125 3430 56135 3750
rect 56155 3430 56165 3750
rect 56125 3415 56165 3430
rect 56185 3750 56225 3765
rect 56185 3430 56195 3750
rect 56215 3430 56225 3750
rect 56185 3415 56225 3430
rect 56245 3750 56285 3765
rect 56245 3430 56255 3750
rect 56275 3430 56285 3750
rect 56245 3415 56285 3430
rect 56305 3750 56345 3765
rect 56305 3430 56315 3750
rect 56335 3430 56345 3750
rect 56305 3415 56345 3430
rect 56365 3750 56405 3765
rect 56365 3430 56375 3750
rect 56395 3430 56405 3750
rect 56365 3415 56405 3430
rect 56425 3750 56465 3765
rect 56425 3430 56435 3750
rect 56455 3430 56465 3750
rect 56425 3415 56465 3430
rect 56485 3750 56525 3765
rect 56485 3430 56495 3750
rect 56515 3430 56525 3750
rect 56485 3415 56525 3430
rect 56545 3750 56585 3765
rect 56545 3430 56555 3750
rect 56575 3430 56585 3750
rect 56545 3415 56585 3430
rect 56605 3750 56645 3765
rect 56605 3430 56615 3750
rect 56635 3430 56645 3750
rect 56605 3415 56645 3430
rect 56665 3750 56705 3765
rect 56665 3430 56675 3750
rect 56695 3430 56705 3750
rect 56665 3415 56705 3430
rect 56725 3750 56765 3765
rect 56725 3430 56735 3750
rect 56755 3430 56765 3750
rect 56725 3415 56765 3430
rect 57035 3750 57075 3765
rect 57035 3430 57045 3750
rect 57065 3430 57075 3750
rect 57035 3415 57075 3430
rect 57095 3750 57135 3765
rect 57095 3430 57105 3750
rect 57125 3430 57135 3750
rect 57095 3415 57135 3430
rect 57155 3750 57195 3765
rect 57155 3430 57165 3750
rect 57185 3430 57195 3750
rect 57155 3415 57195 3430
rect 57215 3750 57255 3765
rect 57215 3430 57225 3750
rect 57245 3430 57255 3750
rect 57215 3415 57255 3430
rect 57275 3750 57315 3765
rect 57275 3430 57285 3750
rect 57305 3430 57315 3750
rect 57275 3415 57315 3430
rect 57335 3750 57375 3765
rect 57335 3430 57345 3750
rect 57365 3430 57375 3750
rect 57335 3415 57375 3430
rect 57395 3750 57435 3765
rect 57395 3430 57405 3750
rect 57425 3430 57435 3750
rect 57395 3415 57435 3430
rect 57455 3750 57495 3765
rect 57455 3430 57465 3750
rect 57485 3430 57495 3750
rect 57455 3415 57495 3430
rect 57515 3750 57555 3765
rect 57515 3430 57525 3750
rect 57545 3430 57555 3750
rect 57515 3415 57555 3430
rect 57575 3750 57615 3765
rect 57575 3430 57585 3750
rect 57605 3430 57615 3750
rect 57575 3415 57615 3430
rect 57635 3750 57675 3765
rect 57635 3430 57645 3750
rect 57665 3430 57675 3750
rect 57635 3415 57675 3430
rect 57695 3750 57735 3765
rect 57695 3430 57705 3750
rect 57725 3430 57735 3750
rect 57695 3415 57735 3430
rect 57755 3750 57795 3765
rect 57755 3430 57765 3750
rect 57785 3430 57795 3750
rect 57755 3415 57795 3430
rect 58410 3750 58450 3765
rect 58410 3430 58420 3750
rect 58440 3430 58450 3750
rect 58410 3415 58450 3430
rect 58470 3750 58510 3765
rect 58470 3430 58480 3750
rect 58500 3430 58510 3750
rect 58470 3415 58510 3430
rect 58530 3750 58570 3765
rect 58530 3430 58540 3750
rect 58560 3430 58570 3750
rect 58530 3415 58570 3430
rect 58590 3750 58630 3765
rect 58590 3430 58600 3750
rect 58620 3430 58630 3750
rect 58590 3415 58630 3430
rect 58650 3750 58690 3765
rect 58650 3430 58660 3750
rect 58680 3430 58690 3750
rect 58650 3415 58690 3430
rect 58710 3750 58750 3765
rect 58710 3430 58720 3750
rect 58740 3430 58750 3750
rect 58710 3415 58750 3430
rect 58770 3750 58810 3765
rect 58770 3430 58780 3750
rect 58800 3430 58810 3750
rect 58770 3415 58810 3430
rect 58830 3750 58870 3765
rect 58830 3430 58840 3750
rect 58860 3430 58870 3750
rect 58830 3415 58870 3430
rect 58890 3750 58930 3765
rect 58890 3430 58900 3750
rect 58920 3430 58930 3750
rect 58890 3415 58930 3430
rect 58950 3750 58990 3765
rect 58950 3430 58960 3750
rect 58980 3430 58990 3750
rect 58950 3415 58990 3430
rect 59010 3750 59050 3765
rect 59010 3430 59020 3750
rect 59040 3430 59050 3750
rect 59010 3415 59050 3430
rect 59070 3750 59110 3765
rect 59070 3430 59080 3750
rect 59100 3430 59110 3750
rect 59070 3415 59110 3430
rect 59130 3750 59170 3765
rect 59130 3430 59140 3750
rect 59160 3430 59170 3750
rect 59130 3415 59170 3430
rect 54740 2890 54780 2905
rect 54740 2320 54750 2890
rect 54770 2320 54780 2890
rect 54740 2305 54780 2320
rect 54795 2890 54835 2905
rect 54795 2320 54805 2890
rect 54825 2320 54835 2890
rect 54795 2305 54835 2320
rect 54850 2890 54890 2905
rect 54850 2320 54860 2890
rect 54880 2320 54890 2890
rect 54850 2305 54890 2320
rect 54905 2890 54945 2905
rect 54905 2320 54915 2890
rect 54935 2320 54945 2890
rect 54905 2305 54945 2320
rect 54960 2890 55000 2905
rect 54960 2320 54970 2890
rect 54990 2320 55000 2890
rect 54960 2305 55000 2320
rect 55015 2890 55055 2905
rect 55015 2320 55025 2890
rect 55045 2320 55055 2890
rect 55015 2305 55055 2320
rect 55070 2890 55110 2905
rect 55070 2320 55080 2890
rect 55100 2320 55110 2890
rect 55070 2305 55110 2320
rect 55125 2890 55165 2905
rect 55125 2320 55135 2890
rect 55155 2320 55165 2890
rect 55125 2305 55165 2320
rect 55180 2890 55220 2905
rect 55180 2320 55190 2890
rect 55210 2320 55220 2890
rect 55180 2305 55220 2320
rect 55235 2890 55275 2905
rect 55235 2320 55245 2890
rect 55265 2320 55275 2890
rect 55235 2305 55275 2320
rect 55290 2890 55330 2905
rect 55290 2320 55300 2890
rect 55320 2320 55330 2890
rect 55290 2305 55330 2320
rect 55345 2890 55385 2905
rect 55345 2320 55355 2890
rect 55375 2320 55385 2890
rect 55345 2305 55385 2320
rect 55400 2890 55440 2905
rect 55400 2320 55410 2890
rect 55430 2320 55440 2890
rect 56510 2895 56550 2910
rect 56510 2875 56520 2895
rect 56540 2875 56550 2895
rect 56510 2845 56550 2875
rect 56510 2825 56520 2845
rect 56540 2825 56550 2845
rect 56510 2795 56550 2825
rect 56510 2775 56520 2795
rect 56540 2775 56550 2795
rect 56510 2745 56550 2775
rect 56510 2725 56520 2745
rect 56540 2725 56550 2745
rect 56510 2695 56550 2725
rect 56510 2675 56520 2695
rect 56540 2675 56550 2695
rect 56510 2660 56550 2675
rect 56565 2895 56605 2910
rect 56565 2875 56575 2895
rect 56595 2875 56605 2895
rect 56565 2845 56605 2875
rect 56565 2825 56575 2845
rect 56595 2825 56605 2845
rect 56565 2795 56605 2825
rect 56565 2775 56575 2795
rect 56595 2775 56605 2795
rect 56565 2745 56605 2775
rect 56565 2725 56575 2745
rect 56595 2725 56605 2745
rect 56565 2695 56605 2725
rect 56565 2675 56575 2695
rect 56595 2675 56605 2695
rect 56565 2660 56605 2675
rect 56620 2895 56660 2910
rect 56620 2875 56630 2895
rect 56650 2875 56660 2895
rect 56620 2845 56660 2875
rect 56620 2825 56630 2845
rect 56650 2825 56660 2845
rect 56620 2795 56660 2825
rect 56620 2775 56630 2795
rect 56650 2775 56660 2795
rect 56620 2745 56660 2775
rect 56620 2725 56630 2745
rect 56650 2725 56660 2745
rect 56620 2695 56660 2725
rect 56620 2675 56630 2695
rect 56650 2675 56660 2695
rect 56620 2660 56660 2675
rect 56675 2895 56715 2910
rect 56675 2875 56685 2895
rect 56705 2875 56715 2895
rect 56675 2845 56715 2875
rect 56675 2825 56685 2845
rect 56705 2825 56715 2845
rect 56675 2795 56715 2825
rect 56675 2775 56685 2795
rect 56705 2775 56715 2795
rect 56675 2745 56715 2775
rect 56675 2725 56685 2745
rect 56705 2725 56715 2745
rect 56675 2695 56715 2725
rect 56675 2675 56685 2695
rect 56705 2675 56715 2695
rect 56675 2660 56715 2675
rect 56730 2895 56770 2910
rect 56730 2875 56740 2895
rect 56760 2875 56770 2895
rect 56730 2845 56770 2875
rect 56730 2825 56740 2845
rect 56760 2825 56770 2845
rect 56730 2795 56770 2825
rect 56730 2775 56740 2795
rect 56760 2775 56770 2795
rect 56730 2745 56770 2775
rect 56730 2725 56740 2745
rect 56760 2725 56770 2745
rect 56730 2695 56770 2725
rect 56730 2675 56740 2695
rect 56760 2675 56770 2695
rect 56730 2660 56770 2675
rect 56785 2895 56825 2910
rect 56785 2875 56795 2895
rect 56815 2875 56825 2895
rect 56785 2845 56825 2875
rect 56785 2825 56795 2845
rect 56815 2825 56825 2845
rect 56785 2795 56825 2825
rect 56785 2775 56795 2795
rect 56815 2775 56825 2795
rect 56785 2745 56825 2775
rect 56785 2725 56795 2745
rect 56815 2725 56825 2745
rect 56785 2695 56825 2725
rect 56785 2675 56795 2695
rect 56815 2675 56825 2695
rect 56785 2660 56825 2675
rect 56840 2895 56880 2910
rect 56920 2895 56960 2910
rect 56840 2875 56850 2895
rect 56870 2875 56880 2895
rect 56920 2875 56930 2895
rect 56950 2875 56960 2895
rect 56840 2845 56880 2875
rect 56920 2845 56960 2875
rect 56840 2825 56850 2845
rect 56870 2825 56880 2845
rect 56920 2825 56930 2845
rect 56950 2825 56960 2845
rect 56840 2795 56880 2825
rect 56920 2795 56960 2825
rect 56840 2775 56850 2795
rect 56870 2775 56880 2795
rect 56920 2775 56930 2795
rect 56950 2775 56960 2795
rect 56840 2745 56880 2775
rect 56920 2745 56960 2775
rect 56840 2725 56850 2745
rect 56870 2725 56880 2745
rect 56920 2725 56930 2745
rect 56950 2725 56960 2745
rect 56840 2695 56880 2725
rect 56920 2695 56960 2725
rect 56840 2675 56850 2695
rect 56870 2675 56880 2695
rect 56920 2675 56930 2695
rect 56950 2675 56960 2695
rect 56840 2660 56880 2675
rect 56920 2660 56960 2675
rect 56975 2895 57015 2910
rect 56975 2875 56985 2895
rect 57005 2875 57015 2895
rect 56975 2845 57015 2875
rect 56975 2825 56985 2845
rect 57005 2825 57015 2845
rect 56975 2795 57015 2825
rect 56975 2775 56985 2795
rect 57005 2775 57015 2795
rect 56975 2745 57015 2775
rect 56975 2725 56985 2745
rect 57005 2725 57015 2745
rect 56975 2695 57015 2725
rect 56975 2675 56985 2695
rect 57005 2675 57015 2695
rect 56975 2660 57015 2675
rect 57030 2895 57070 2910
rect 57030 2875 57040 2895
rect 57060 2875 57070 2895
rect 57030 2845 57070 2875
rect 57030 2825 57040 2845
rect 57060 2825 57070 2845
rect 57030 2795 57070 2825
rect 57030 2775 57040 2795
rect 57060 2775 57070 2795
rect 57030 2745 57070 2775
rect 57030 2725 57040 2745
rect 57060 2725 57070 2745
rect 57030 2695 57070 2725
rect 57030 2675 57040 2695
rect 57060 2675 57070 2695
rect 57030 2660 57070 2675
rect 57085 2895 57125 2910
rect 57085 2875 57095 2895
rect 57115 2875 57125 2895
rect 57085 2845 57125 2875
rect 57085 2825 57095 2845
rect 57115 2825 57125 2845
rect 57085 2795 57125 2825
rect 57085 2775 57095 2795
rect 57115 2775 57125 2795
rect 57085 2745 57125 2775
rect 57085 2725 57095 2745
rect 57115 2725 57125 2745
rect 57085 2695 57125 2725
rect 57085 2675 57095 2695
rect 57115 2675 57125 2695
rect 57085 2660 57125 2675
rect 57140 2895 57180 2910
rect 57140 2875 57150 2895
rect 57170 2875 57180 2895
rect 57140 2845 57180 2875
rect 57140 2825 57150 2845
rect 57170 2825 57180 2845
rect 57140 2795 57180 2825
rect 57140 2775 57150 2795
rect 57170 2775 57180 2795
rect 57140 2745 57180 2775
rect 57140 2725 57150 2745
rect 57170 2725 57180 2745
rect 57140 2695 57180 2725
rect 57140 2675 57150 2695
rect 57170 2675 57180 2695
rect 57140 2660 57180 2675
rect 57195 2895 57235 2910
rect 57195 2875 57205 2895
rect 57225 2875 57235 2895
rect 57195 2845 57235 2875
rect 57195 2825 57205 2845
rect 57225 2825 57235 2845
rect 57195 2795 57235 2825
rect 57195 2775 57205 2795
rect 57225 2775 57235 2795
rect 57195 2745 57235 2775
rect 57195 2725 57205 2745
rect 57225 2725 57235 2745
rect 57195 2695 57235 2725
rect 57195 2675 57205 2695
rect 57225 2675 57235 2695
rect 57195 2660 57235 2675
rect 57250 2895 57290 2910
rect 57250 2875 57260 2895
rect 57280 2875 57290 2895
rect 57250 2845 57290 2875
rect 57250 2825 57260 2845
rect 57280 2825 57290 2845
rect 57250 2795 57290 2825
rect 57250 2775 57260 2795
rect 57280 2775 57290 2795
rect 57250 2745 57290 2775
rect 57250 2725 57260 2745
rect 57280 2725 57290 2745
rect 57250 2695 57290 2725
rect 57250 2675 57260 2695
rect 57280 2675 57290 2695
rect 57250 2660 57290 2675
rect 58440 2890 58480 2905
rect 55400 2305 55440 2320
rect 58440 2320 58450 2890
rect 58470 2320 58480 2890
rect 58440 2305 58480 2320
rect 58495 2890 58535 2905
rect 58495 2320 58505 2890
rect 58525 2320 58535 2890
rect 58495 2305 58535 2320
rect 58550 2890 58590 2905
rect 58550 2320 58560 2890
rect 58580 2320 58590 2890
rect 58550 2305 58590 2320
rect 58605 2890 58645 2905
rect 58605 2320 58615 2890
rect 58635 2320 58645 2890
rect 58605 2305 58645 2320
rect 58660 2890 58700 2905
rect 58660 2320 58670 2890
rect 58690 2320 58700 2890
rect 58660 2305 58700 2320
rect 58715 2890 58755 2905
rect 58715 2320 58725 2890
rect 58745 2320 58755 2890
rect 58715 2305 58755 2320
rect 58770 2890 58810 2905
rect 58770 2320 58780 2890
rect 58800 2320 58810 2890
rect 58770 2305 58810 2320
rect 58825 2890 58865 2905
rect 58825 2320 58835 2890
rect 58855 2320 58865 2890
rect 58825 2305 58865 2320
rect 58880 2890 58920 2905
rect 58880 2320 58890 2890
rect 58910 2320 58920 2890
rect 58880 2305 58920 2320
rect 58935 2890 58975 2905
rect 58935 2320 58945 2890
rect 58965 2320 58975 2890
rect 58935 2305 58975 2320
rect 58990 2890 59030 2905
rect 58990 2320 59000 2890
rect 59020 2320 59030 2890
rect 58990 2305 59030 2320
rect 59045 2890 59085 2905
rect 59045 2320 59055 2890
rect 59075 2320 59085 2890
rect 59045 2305 59085 2320
rect 59100 2890 59140 2905
rect 59100 2320 59110 2890
rect 59130 2320 59140 2890
rect 59100 2305 59140 2320
rect 54740 1615 54780 1630
rect 54740 1445 54750 1615
rect 54770 1445 54780 1615
rect 54740 1430 54780 1445
rect 54795 1615 54835 1630
rect 54795 1445 54805 1615
rect 54825 1445 54835 1615
rect 54795 1430 54835 1445
rect 54850 1615 54890 1630
rect 54850 1445 54860 1615
rect 54880 1445 54890 1615
rect 54850 1430 54890 1445
rect 54905 1615 54945 1630
rect 54905 1445 54915 1615
rect 54935 1445 54945 1615
rect 54905 1430 54945 1445
rect 54960 1615 55000 1630
rect 54960 1445 54970 1615
rect 54990 1445 55000 1615
rect 54960 1430 55000 1445
rect 55015 1615 55055 1630
rect 55015 1445 55025 1615
rect 55045 1445 55055 1615
rect 55015 1430 55055 1445
rect 55070 1615 55110 1630
rect 55070 1445 55080 1615
rect 55100 1445 55110 1615
rect 55070 1430 55110 1445
rect 55125 1615 55165 1630
rect 55125 1445 55135 1615
rect 55155 1445 55165 1615
rect 55125 1430 55165 1445
rect 55180 1615 55220 1630
rect 55180 1445 55190 1615
rect 55210 1445 55220 1615
rect 55180 1430 55220 1445
rect 55235 1615 55275 1630
rect 55235 1445 55245 1615
rect 55265 1445 55275 1615
rect 55235 1430 55275 1445
rect 55290 1615 55330 1630
rect 55290 1445 55300 1615
rect 55320 1445 55330 1615
rect 55290 1430 55330 1445
rect 55345 1615 55385 1630
rect 55345 1445 55355 1615
rect 55375 1445 55385 1615
rect 55345 1430 55385 1445
rect 55400 1615 55440 1630
rect 55400 1445 55410 1615
rect 55430 1445 55440 1615
rect 58440 1615 58480 1630
rect 55400 1430 55440 1445
rect 58440 1445 58450 1615
rect 58470 1445 58480 1615
rect 58440 1430 58480 1445
rect 58495 1615 58535 1630
rect 58495 1445 58505 1615
rect 58525 1445 58535 1615
rect 58495 1430 58535 1445
rect 58550 1615 58590 1630
rect 58550 1445 58560 1615
rect 58580 1445 58590 1615
rect 58550 1430 58590 1445
rect 58605 1615 58645 1630
rect 58605 1445 58615 1615
rect 58635 1445 58645 1615
rect 58605 1430 58645 1445
rect 58660 1615 58700 1630
rect 58660 1445 58670 1615
rect 58690 1445 58700 1615
rect 58660 1430 58700 1445
rect 58715 1615 58755 1630
rect 58715 1445 58725 1615
rect 58745 1445 58755 1615
rect 58715 1430 58755 1445
rect 58770 1615 58810 1630
rect 58770 1445 58780 1615
rect 58800 1445 58810 1615
rect 58770 1430 58810 1445
rect 58825 1615 58865 1630
rect 58825 1445 58835 1615
rect 58855 1445 58865 1615
rect 58825 1430 58865 1445
rect 58880 1615 58920 1630
rect 58880 1445 58890 1615
rect 58910 1445 58920 1615
rect 58880 1430 58920 1445
rect 58935 1615 58975 1630
rect 58935 1445 58945 1615
rect 58965 1445 58975 1615
rect 58935 1430 58975 1445
rect 58990 1615 59030 1630
rect 58990 1445 59000 1615
rect 59020 1445 59030 1615
rect 58990 1430 59030 1445
rect 59045 1615 59085 1630
rect 59045 1445 59055 1615
rect 59075 1445 59085 1615
rect 59045 1430 59085 1445
rect 59100 1615 59140 1630
rect 59100 1445 59110 1615
rect 59130 1445 59140 1615
rect 59100 1430 59140 1445
<< ndiffc >>
rect 56780 2080 56800 2300
rect 56835 2080 56855 2300
rect 56890 2080 56910 2300
rect 56945 2080 56965 2300
rect 57000 2080 57020 2300
rect 56040 1510 56060 1630
rect 56095 1510 56115 1630
rect 56150 1510 56170 1630
rect 56205 1510 56225 1630
rect 56260 1510 56280 1630
rect 56315 1510 56335 1630
rect 56370 1510 56390 1630
rect 56425 1510 56445 1630
rect 56480 1510 56500 1630
rect 56535 1510 56555 1630
rect 56590 1510 56610 1630
rect 56645 1510 56665 1630
rect 56700 1510 56720 1630
rect 57080 1510 57100 1630
rect 57135 1510 57155 1630
rect 57190 1510 57210 1630
rect 57245 1510 57265 1630
rect 57300 1510 57320 1630
rect 57355 1510 57375 1630
rect 57410 1510 57430 1630
rect 57465 1510 57485 1630
rect 57520 1510 57540 1630
rect 57575 1510 57595 1630
rect 57630 1510 57650 1630
rect 57685 1510 57705 1630
rect 57740 1510 57760 1630
rect 54750 905 54770 1175
rect 54805 905 54825 1175
rect 54860 905 54880 1175
rect 54915 905 54935 1175
rect 54970 905 54990 1175
rect 55025 905 55045 1175
rect 55080 905 55100 1175
rect 55135 905 55155 1175
rect 55190 905 55210 1175
rect 55245 905 55265 1175
rect 55300 905 55320 1175
rect 55355 905 55375 1175
rect 55410 905 55430 1175
rect 56040 835 56060 955
rect 56095 835 56115 955
rect 56150 835 56170 955
rect 56205 835 56225 955
rect 56260 835 56280 955
rect 56315 835 56335 955
rect 56370 835 56390 955
rect 56425 835 56445 955
rect 56480 835 56500 955
rect 56535 835 56555 955
rect 56590 835 56610 955
rect 56645 835 56665 955
rect 56700 835 56720 955
rect 56780 835 56800 955
rect 56835 835 56855 955
rect 56890 835 56910 955
rect 56945 835 56965 955
rect 57000 835 57020 955
rect 57080 835 57100 955
rect 57135 835 57155 955
rect 57190 835 57210 955
rect 57245 835 57265 955
rect 57300 835 57320 955
rect 57355 835 57375 955
rect 57410 835 57430 955
rect 57465 835 57485 955
rect 57520 835 57540 955
rect 57575 835 57595 955
rect 57630 835 57650 955
rect 57685 835 57705 955
rect 57740 835 57760 955
rect 58450 905 58470 1175
rect 58505 905 58525 1175
rect 58560 905 58580 1175
rect 58615 905 58635 1175
rect 58670 905 58690 1175
rect 58725 905 58745 1175
rect 58780 905 58800 1175
rect 58835 905 58855 1175
rect 58890 905 58910 1175
rect 58945 905 58965 1175
rect 59000 905 59020 1175
rect 59055 905 59075 1175
rect 59110 905 59130 1175
rect 54760 -505 54780 165
rect 54860 -505 54880 165
rect 54960 -505 54980 165
rect 55060 -505 55080 165
rect 55160 -505 55180 165
rect 55260 -505 55280 165
rect 55360 -505 55380 165
rect 56230 95 56250 315
rect 56285 95 56305 315
rect 56340 95 56360 315
rect 56395 95 56415 315
rect 56450 95 56470 315
rect 56505 95 56525 315
rect 56560 95 56580 315
rect 56615 95 56635 315
rect 56670 95 56690 315
rect 56725 95 56745 315
rect 56780 95 56800 315
rect 56835 95 56855 315
rect 56890 95 56910 315
rect 56945 95 56965 315
rect 57000 95 57020 315
rect 57055 95 57075 315
rect 57110 95 57130 315
rect 57165 95 57185 315
rect 57220 95 57240 315
rect 57275 95 57295 315
rect 57330 95 57350 315
rect 57385 95 57405 315
rect 57440 95 57460 315
rect 57495 95 57515 315
rect 56440 -460 56460 -340
rect 56495 -460 56515 -340
rect 56550 -460 56570 -340
rect 56605 -460 56625 -340
rect 56660 -460 56680 -340
rect 56715 -460 56735 -340
rect 56770 -460 56790 -340
rect 56880 -460 56900 -340
rect 57220 -460 57240 -340
rect 58340 -505 58360 165
rect 58440 -505 58460 165
rect 58540 -505 58560 165
rect 58640 -505 58660 165
rect 58740 -505 58760 165
rect 58840 -505 58860 165
rect 58940 -505 58960 165
<< pdiffc >>
rect 56095 4545 56115 4865
rect 56155 4545 56175 4865
rect 56215 4545 56235 4865
rect 56275 4545 56295 4865
rect 56565 4545 56585 4695
rect 56625 4545 56645 4695
rect 56685 4545 56705 4695
rect 56745 4545 56765 4695
rect 57035 4545 57055 4865
rect 57095 4545 57115 4865
rect 57155 4545 57175 4865
rect 57215 4545 57235 4865
rect 57505 4545 57525 4865
rect 57565 4545 57585 4865
rect 57625 4545 57645 4865
rect 57685 4545 57705 4865
rect 54850 3430 54870 3750
rect 54910 3430 54930 3750
rect 54970 3430 54990 3750
rect 55030 3430 55050 3750
rect 55090 3430 55110 3750
rect 55150 3430 55170 3750
rect 55210 3430 55230 3750
rect 55270 3430 55290 3750
rect 55330 3430 55350 3750
rect 55390 3430 55410 3750
rect 55450 3430 55470 3750
rect 55510 3430 55530 3750
rect 55570 3430 55590 3750
rect 56015 3430 56035 3750
rect 56075 3430 56095 3750
rect 56135 3430 56155 3750
rect 56195 3430 56215 3750
rect 56255 3430 56275 3750
rect 56315 3430 56335 3750
rect 56375 3430 56395 3750
rect 56435 3430 56455 3750
rect 56495 3430 56515 3750
rect 56555 3430 56575 3750
rect 56615 3430 56635 3750
rect 56675 3430 56695 3750
rect 56735 3430 56755 3750
rect 57045 3430 57065 3750
rect 57105 3430 57125 3750
rect 57165 3430 57185 3750
rect 57225 3430 57245 3750
rect 57285 3430 57305 3750
rect 57345 3430 57365 3750
rect 57405 3430 57425 3750
rect 57465 3430 57485 3750
rect 57525 3430 57545 3750
rect 57585 3430 57605 3750
rect 57645 3430 57665 3750
rect 57705 3430 57725 3750
rect 57765 3430 57785 3750
rect 58420 3430 58440 3750
rect 58480 3430 58500 3750
rect 58540 3430 58560 3750
rect 58600 3430 58620 3750
rect 58660 3430 58680 3750
rect 58720 3430 58740 3750
rect 58780 3430 58800 3750
rect 58840 3430 58860 3750
rect 58900 3430 58920 3750
rect 58960 3430 58980 3750
rect 59020 3430 59040 3750
rect 59080 3430 59100 3750
rect 59140 3430 59160 3750
rect 54750 2320 54770 2890
rect 54805 2320 54825 2890
rect 54860 2320 54880 2890
rect 54915 2320 54935 2890
rect 54970 2320 54990 2890
rect 55025 2320 55045 2890
rect 55080 2320 55100 2890
rect 55135 2320 55155 2890
rect 55190 2320 55210 2890
rect 55245 2320 55265 2890
rect 55300 2320 55320 2890
rect 55355 2320 55375 2890
rect 55410 2320 55430 2890
rect 56520 2875 56540 2895
rect 56520 2825 56540 2845
rect 56520 2775 56540 2795
rect 56520 2725 56540 2745
rect 56520 2675 56540 2695
rect 56575 2875 56595 2895
rect 56575 2825 56595 2845
rect 56575 2775 56595 2795
rect 56575 2725 56595 2745
rect 56575 2675 56595 2695
rect 56630 2875 56650 2895
rect 56630 2825 56650 2845
rect 56630 2775 56650 2795
rect 56630 2725 56650 2745
rect 56630 2675 56650 2695
rect 56685 2875 56705 2895
rect 56685 2825 56705 2845
rect 56685 2775 56705 2795
rect 56685 2725 56705 2745
rect 56685 2675 56705 2695
rect 56740 2875 56760 2895
rect 56740 2825 56760 2845
rect 56740 2775 56760 2795
rect 56740 2725 56760 2745
rect 56740 2675 56760 2695
rect 56795 2875 56815 2895
rect 56795 2825 56815 2845
rect 56795 2775 56815 2795
rect 56795 2725 56815 2745
rect 56795 2675 56815 2695
rect 56850 2875 56870 2895
rect 56930 2875 56950 2895
rect 56850 2825 56870 2845
rect 56930 2825 56950 2845
rect 56850 2775 56870 2795
rect 56930 2775 56950 2795
rect 56850 2725 56870 2745
rect 56930 2725 56950 2745
rect 56850 2675 56870 2695
rect 56930 2675 56950 2695
rect 56985 2875 57005 2895
rect 56985 2825 57005 2845
rect 56985 2775 57005 2795
rect 56985 2725 57005 2745
rect 56985 2675 57005 2695
rect 57040 2875 57060 2895
rect 57040 2825 57060 2845
rect 57040 2775 57060 2795
rect 57040 2725 57060 2745
rect 57040 2675 57060 2695
rect 57095 2875 57115 2895
rect 57095 2825 57115 2845
rect 57095 2775 57115 2795
rect 57095 2725 57115 2745
rect 57095 2675 57115 2695
rect 57150 2875 57170 2895
rect 57150 2825 57170 2845
rect 57150 2775 57170 2795
rect 57150 2725 57170 2745
rect 57150 2675 57170 2695
rect 57205 2875 57225 2895
rect 57205 2825 57225 2845
rect 57205 2775 57225 2795
rect 57205 2725 57225 2745
rect 57205 2675 57225 2695
rect 57260 2875 57280 2895
rect 57260 2825 57280 2845
rect 57260 2775 57280 2795
rect 57260 2725 57280 2745
rect 57260 2675 57280 2695
rect 58450 2320 58470 2890
rect 58505 2320 58525 2890
rect 58560 2320 58580 2890
rect 58615 2320 58635 2890
rect 58670 2320 58690 2890
rect 58725 2320 58745 2890
rect 58780 2320 58800 2890
rect 58835 2320 58855 2890
rect 58890 2320 58910 2890
rect 58945 2320 58965 2890
rect 59000 2320 59020 2890
rect 59055 2320 59075 2890
rect 59110 2320 59130 2890
rect 54750 1445 54770 1615
rect 54805 1445 54825 1615
rect 54860 1445 54880 1615
rect 54915 1445 54935 1615
rect 54970 1445 54990 1615
rect 55025 1445 55045 1615
rect 55080 1445 55100 1615
rect 55135 1445 55155 1615
rect 55190 1445 55210 1615
rect 55245 1445 55265 1615
rect 55300 1445 55320 1615
rect 55355 1445 55375 1615
rect 55410 1445 55430 1615
rect 58450 1445 58470 1615
rect 58505 1445 58525 1615
rect 58560 1445 58580 1615
rect 58615 1445 58635 1615
rect 58670 1445 58690 1615
rect 58725 1445 58745 1615
rect 58780 1445 58800 1615
rect 58835 1445 58855 1615
rect 58890 1445 58910 1615
rect 58945 1445 58965 1615
rect 59000 1445 59020 1615
rect 59055 1445 59075 1615
rect 59110 1445 59130 1615
<< psubdiff >>
rect 56730 2300 56770 2315
rect 56730 2080 56740 2300
rect 56760 2080 56770 2300
rect 56730 2065 56770 2080
rect 57030 2300 57070 2315
rect 57030 2080 57040 2300
rect 57060 2080 57070 2300
rect 57030 2065 57070 2080
rect 55990 1630 56030 1645
rect 55990 1510 56000 1630
rect 56020 1510 56030 1630
rect 55990 1495 56030 1510
rect 56730 1630 56770 1645
rect 56730 1510 56740 1630
rect 56760 1510 56770 1630
rect 56730 1495 56770 1510
rect 57030 1630 57070 1645
rect 57030 1510 57040 1630
rect 57060 1510 57070 1630
rect 57030 1495 57070 1510
rect 57770 1630 57810 1645
rect 57770 1510 57780 1630
rect 57800 1510 57810 1630
rect 57770 1495 57810 1510
rect 54700 1175 54740 1190
rect 54700 905 54710 1175
rect 54730 905 54740 1175
rect 54700 890 54740 905
rect 55440 1175 55480 1190
rect 55440 905 55450 1175
rect 55470 905 55480 1175
rect 58400 1175 58440 1190
rect 55440 890 55480 905
rect 55990 955 56030 970
rect 55990 835 56000 955
rect 56020 835 56030 955
rect 55990 820 56030 835
rect 56730 955 56770 970
rect 56730 835 56740 955
rect 56760 835 56770 955
rect 56730 820 56770 835
rect 57030 955 57070 970
rect 57030 835 57040 955
rect 57060 835 57070 955
rect 57030 820 57070 835
rect 57770 955 57810 970
rect 57770 835 57780 955
rect 57800 835 57810 955
rect 58400 905 58410 1175
rect 58430 905 58440 1175
rect 58400 890 58440 905
rect 59140 1175 59180 1190
rect 59140 905 59150 1175
rect 59170 905 59180 1175
rect 59140 890 59180 905
rect 57770 820 57810 835
rect 56180 315 56220 330
rect 54710 165 54750 180
rect 54710 -505 54720 165
rect 54740 -505 54750 165
rect 54710 -520 54750 -505
rect 55390 165 55430 180
rect 55390 -505 55400 165
rect 55420 -505 55430 165
rect 56180 95 56190 315
rect 56210 95 56220 315
rect 56180 80 56220 95
rect 57525 315 57565 330
rect 57525 95 57535 315
rect 57555 95 57565 315
rect 57525 80 57565 95
rect 58290 165 58330 180
rect 56390 -340 56430 -325
rect 56390 -460 56400 -340
rect 56420 -460 56430 -340
rect 56390 -475 56430 -460
rect 56800 -340 56840 -325
rect 56800 -460 56810 -340
rect 56830 -460 56840 -340
rect 56800 -475 56840 -460
rect 55390 -520 55430 -505
rect 58290 -505 58300 165
rect 58320 -505 58330 165
rect 58290 -520 58330 -505
rect 58970 165 59010 180
rect 58970 -505 58980 165
rect 59000 -505 59010 165
rect 58970 -520 59010 -505
<< nsubdiff >>
rect 56045 4865 56085 4880
rect 56045 4545 56055 4865
rect 56075 4545 56085 4865
rect 56045 4530 56085 4545
rect 56305 4865 56345 4880
rect 56305 4545 56315 4865
rect 56335 4545 56345 4865
rect 56985 4865 57025 4880
rect 56305 4530 56345 4545
rect 56515 4695 56555 4710
rect 56515 4545 56525 4695
rect 56545 4545 56555 4695
rect 56515 4530 56555 4545
rect 56775 4695 56815 4710
rect 56775 4545 56785 4695
rect 56805 4545 56815 4695
rect 56775 4530 56815 4545
rect 56985 4545 56995 4865
rect 57015 4545 57025 4865
rect 56985 4530 57025 4545
rect 57245 4865 57285 4880
rect 57245 4545 57255 4865
rect 57275 4545 57285 4865
rect 57245 4530 57285 4545
rect 57455 4865 57495 4880
rect 57455 4545 57465 4865
rect 57485 4545 57495 4865
rect 57455 4530 57495 4545
rect 57715 4865 57755 4880
rect 57715 4545 57725 4865
rect 57745 4545 57755 4865
rect 57715 4530 57755 4545
rect 54800 3750 54840 3765
rect 54800 3430 54810 3750
rect 54830 3430 54840 3750
rect 54800 3415 54840 3430
rect 55600 3750 55640 3765
rect 55600 3430 55610 3750
rect 55630 3430 55640 3750
rect 55600 3415 55640 3430
rect 55965 3750 56005 3765
rect 55965 3430 55975 3750
rect 55995 3430 56005 3750
rect 55965 3415 56005 3430
rect 56765 3750 56805 3765
rect 56765 3430 56775 3750
rect 56795 3430 56805 3750
rect 56765 3415 56805 3430
rect 56995 3750 57035 3765
rect 56995 3430 57005 3750
rect 57025 3430 57035 3750
rect 56995 3415 57035 3430
rect 57795 3750 57835 3765
rect 57795 3430 57805 3750
rect 57825 3430 57835 3750
rect 57795 3415 57835 3430
rect 58370 3750 58410 3765
rect 58370 3430 58380 3750
rect 58400 3430 58410 3750
rect 58370 3415 58410 3430
rect 59170 3750 59210 3765
rect 59170 3430 59180 3750
rect 59200 3430 59210 3750
rect 59170 3415 59210 3430
rect 54700 2890 54740 2905
rect 54700 2320 54710 2890
rect 54730 2320 54740 2890
rect 54700 2305 54740 2320
rect 55440 2890 55480 2905
rect 55440 2320 55450 2890
rect 55470 2320 55480 2890
rect 56470 2895 56510 2910
rect 56470 2875 56480 2895
rect 56500 2875 56510 2895
rect 56470 2845 56510 2875
rect 56470 2825 56480 2845
rect 56500 2825 56510 2845
rect 56470 2795 56510 2825
rect 56470 2775 56480 2795
rect 56500 2775 56510 2795
rect 56470 2745 56510 2775
rect 56470 2725 56480 2745
rect 56500 2725 56510 2745
rect 56470 2695 56510 2725
rect 56470 2675 56480 2695
rect 56500 2675 56510 2695
rect 56470 2660 56510 2675
rect 56880 2895 56920 2910
rect 56880 2875 56890 2895
rect 56910 2875 56920 2895
rect 56880 2845 56920 2875
rect 56880 2825 56890 2845
rect 56910 2825 56920 2845
rect 56880 2795 56920 2825
rect 56880 2775 56890 2795
rect 56910 2775 56920 2795
rect 56880 2745 56920 2775
rect 56880 2725 56890 2745
rect 56910 2725 56920 2745
rect 56880 2695 56920 2725
rect 56880 2675 56890 2695
rect 56910 2675 56920 2695
rect 56880 2660 56920 2675
rect 57290 2895 57330 2910
rect 57290 2875 57300 2895
rect 57320 2875 57330 2895
rect 57290 2845 57330 2875
rect 57290 2825 57300 2845
rect 57320 2825 57330 2845
rect 57290 2795 57330 2825
rect 57290 2775 57300 2795
rect 57320 2775 57330 2795
rect 57290 2745 57330 2775
rect 57290 2725 57300 2745
rect 57320 2725 57330 2745
rect 57290 2695 57330 2725
rect 57290 2675 57300 2695
rect 57320 2675 57330 2695
rect 57290 2660 57330 2675
rect 58400 2890 58440 2905
rect 55440 2305 55480 2320
rect 58400 2320 58410 2890
rect 58430 2320 58440 2890
rect 58400 2305 58440 2320
rect 59140 2890 59180 2905
rect 59140 2320 59150 2890
rect 59170 2320 59180 2890
rect 59140 2305 59180 2320
rect 54700 1615 54740 1630
rect 54700 1445 54710 1615
rect 54730 1445 54740 1615
rect 54700 1430 54740 1445
rect 55440 1615 55480 1630
rect 55440 1445 55450 1615
rect 55470 1445 55480 1615
rect 58400 1615 58440 1630
rect 55440 1430 55480 1445
rect 58400 1445 58410 1615
rect 58430 1445 58440 1615
rect 58400 1430 58440 1445
rect 59140 1615 59180 1630
rect 59140 1445 59150 1615
rect 59170 1445 59180 1615
rect 59140 1430 59180 1445
<< psubdiffcont >>
rect 56740 2080 56760 2300
rect 57040 2080 57060 2300
rect 56000 1510 56020 1630
rect 56740 1510 56760 1630
rect 57040 1510 57060 1630
rect 57780 1510 57800 1630
rect 54710 905 54730 1175
rect 55450 905 55470 1175
rect 56000 835 56020 955
rect 56740 835 56760 955
rect 57040 835 57060 955
rect 57780 835 57800 955
rect 58410 905 58430 1175
rect 59150 905 59170 1175
rect 54720 -505 54740 165
rect 55400 -505 55420 165
rect 56190 95 56210 315
rect 57535 95 57555 315
rect 56400 -460 56420 -340
rect 56810 -460 56830 -340
rect 58300 -505 58320 165
rect 58980 -505 59000 165
<< nsubdiffcont >>
rect 56055 4545 56075 4865
rect 56315 4545 56335 4865
rect 56525 4545 56545 4695
rect 56785 4545 56805 4695
rect 56995 4545 57015 4865
rect 57255 4545 57275 4865
rect 57465 4545 57485 4865
rect 57725 4545 57745 4865
rect 54810 3430 54830 3750
rect 55610 3430 55630 3750
rect 55975 3430 55995 3750
rect 56775 3430 56795 3750
rect 57005 3430 57025 3750
rect 57805 3430 57825 3750
rect 58380 3430 58400 3750
rect 59180 3430 59200 3750
rect 54710 2320 54730 2890
rect 55450 2320 55470 2890
rect 56480 2875 56500 2895
rect 56480 2825 56500 2845
rect 56480 2775 56500 2795
rect 56480 2725 56500 2745
rect 56480 2675 56500 2695
rect 56890 2875 56910 2895
rect 56890 2825 56910 2845
rect 56890 2775 56910 2795
rect 56890 2725 56910 2745
rect 56890 2675 56910 2695
rect 57300 2875 57320 2895
rect 57300 2825 57320 2845
rect 57300 2775 57320 2795
rect 57300 2725 57320 2745
rect 57300 2675 57320 2695
rect 58410 2320 58430 2890
rect 59150 2320 59170 2890
rect 54710 1445 54730 1615
rect 55450 1445 55470 1615
rect 58410 1445 58430 1615
rect 59150 1445 59170 1615
<< poly >>
rect 56085 4925 56125 4935
rect 56085 4905 56095 4925
rect 56115 4910 56125 4925
rect 56265 4925 56305 4935
rect 56265 4910 56275 4925
rect 56115 4905 56145 4910
rect 56085 4895 56145 4905
rect 56245 4905 56275 4910
rect 56295 4905 56305 4925
rect 56245 4895 56305 4905
rect 57025 4925 57065 4935
rect 57025 4905 57035 4925
rect 57055 4910 57065 4925
rect 57205 4925 57245 4935
rect 57205 4910 57215 4925
rect 57055 4905 57085 4910
rect 57025 4895 57085 4905
rect 57185 4905 57215 4910
rect 57235 4905 57245 4925
rect 57185 4895 57245 4905
rect 57495 4925 57535 4935
rect 57495 4905 57505 4925
rect 57525 4910 57535 4925
rect 57675 4925 57715 4935
rect 57675 4910 57685 4925
rect 57525 4905 57555 4910
rect 57495 4895 57555 4905
rect 57655 4905 57685 4910
rect 57705 4905 57715 4925
rect 57655 4895 57715 4905
rect 56125 4880 56145 4895
rect 56185 4880 56205 4895
rect 56245 4880 56265 4895
rect 57065 4880 57085 4895
rect 57125 4880 57145 4895
rect 57185 4880 57205 4895
rect 57535 4880 57555 4895
rect 57595 4880 57615 4895
rect 57655 4880 57675 4895
rect 56555 4755 56595 4765
rect 56555 4735 56565 4755
rect 56585 4740 56595 4755
rect 56735 4755 56775 4765
rect 56735 4740 56745 4755
rect 56585 4735 56615 4740
rect 56555 4725 56615 4735
rect 56715 4735 56745 4740
rect 56765 4735 56775 4755
rect 56715 4725 56775 4735
rect 56595 4710 56615 4725
rect 56655 4710 56675 4725
rect 56715 4710 56735 4725
rect 56125 4515 56145 4530
rect 56185 4485 56205 4530
rect 56245 4515 56265 4530
rect 56595 4515 56615 4530
rect 56655 4485 56675 4530
rect 56715 4515 56735 4530
rect 57065 4515 57085 4530
rect 56150 4475 56205 4485
rect 56150 4455 56160 4475
rect 56180 4455 56205 4475
rect 56150 4445 56205 4455
rect 56630 4475 56675 4485
rect 56630 4455 56635 4475
rect 56655 4470 56675 4475
rect 57125 4485 57145 4530
rect 57185 4515 57205 4530
rect 57535 4515 57555 4530
rect 57125 4475 57170 4485
rect 57595 4475 57615 4530
rect 57655 4515 57675 4530
rect 57125 4470 57145 4475
rect 56655 4455 56660 4470
rect 56630 4445 56660 4455
rect 57140 4455 57145 4470
rect 57165 4455 57170 4475
rect 57140 4445 57170 4455
rect 57576 4465 57615 4475
rect 57576 4445 57581 4465
rect 57601 4460 57615 4465
rect 57601 4445 57606 4460
rect 57576 4435 57606 4445
rect 54880 3765 54900 3780
rect 54940 3765 54960 3780
rect 55000 3765 55020 3780
rect 55060 3765 55080 3780
rect 55120 3765 55140 3780
rect 55180 3765 55200 3780
rect 55240 3765 55260 3780
rect 55300 3765 55320 3780
rect 55360 3765 55380 3780
rect 55420 3765 55440 3780
rect 55480 3765 55500 3780
rect 55540 3765 55560 3780
rect 56045 3765 56065 3780
rect 56105 3765 56125 3780
rect 56165 3765 56185 3780
rect 56225 3765 56245 3780
rect 56285 3765 56305 3780
rect 56345 3765 56365 3780
rect 56405 3765 56425 3780
rect 56465 3765 56485 3780
rect 56525 3765 56545 3780
rect 56585 3765 56605 3780
rect 56645 3765 56665 3780
rect 56705 3765 56725 3780
rect 57075 3765 57095 3780
rect 57135 3765 57155 3780
rect 57195 3765 57215 3780
rect 57255 3765 57275 3780
rect 57315 3765 57335 3780
rect 57375 3765 57395 3780
rect 57435 3765 57455 3780
rect 57495 3765 57515 3780
rect 57555 3765 57575 3780
rect 57615 3765 57635 3780
rect 57675 3765 57695 3780
rect 57735 3765 57755 3780
rect 58450 3765 58470 3780
rect 58510 3765 58530 3780
rect 58570 3765 58590 3780
rect 58630 3765 58650 3780
rect 58690 3765 58710 3780
rect 58750 3765 58770 3780
rect 58810 3765 58830 3780
rect 58870 3765 58890 3780
rect 58930 3765 58950 3780
rect 58990 3765 59010 3780
rect 59050 3765 59070 3780
rect 59110 3765 59130 3780
rect 54880 3400 54900 3415
rect 54845 3390 54900 3400
rect 54940 3405 54960 3415
rect 55000 3405 55020 3415
rect 55060 3405 55080 3415
rect 55120 3405 55140 3415
rect 55180 3405 55200 3415
rect 55240 3405 55260 3415
rect 55300 3405 55320 3415
rect 55360 3405 55380 3415
rect 55420 3405 55440 3415
rect 55480 3405 55500 3415
rect 54940 3390 55500 3405
rect 55540 3400 55560 3415
rect 56045 3400 56065 3415
rect 55540 3390 55595 3400
rect 54845 3370 54850 3390
rect 54870 3385 54900 3390
rect 54870 3370 54875 3385
rect 54845 3360 54875 3370
rect 55205 3370 55210 3390
rect 55230 3370 55235 3390
rect 55540 3385 55570 3390
rect 55205 3360 55235 3370
rect 55565 3370 55570 3385
rect 55590 3370 55595 3390
rect 55565 3360 55595 3370
rect 56010 3390 56065 3400
rect 56105 3405 56125 3415
rect 56165 3405 56185 3415
rect 56225 3405 56245 3415
rect 56285 3405 56305 3415
rect 56345 3405 56365 3415
rect 56405 3405 56425 3415
rect 56465 3405 56485 3415
rect 56525 3405 56545 3415
rect 56585 3405 56605 3415
rect 56645 3405 56665 3415
rect 56105 3390 56665 3405
rect 56705 3400 56725 3415
rect 57075 3400 57095 3415
rect 56705 3390 56760 3400
rect 56010 3370 56015 3390
rect 56035 3385 56065 3390
rect 56035 3370 56040 3385
rect 56010 3360 56040 3370
rect 56370 3370 56375 3390
rect 56395 3370 56400 3390
rect 56705 3385 56735 3390
rect 56370 3360 56400 3370
rect 56730 3370 56735 3385
rect 56755 3370 56760 3390
rect 56730 3360 56760 3370
rect 57040 3390 57095 3400
rect 57135 3405 57155 3415
rect 57195 3405 57215 3415
rect 57255 3405 57275 3415
rect 57315 3405 57335 3415
rect 57375 3405 57395 3415
rect 57435 3405 57455 3415
rect 57495 3405 57515 3415
rect 57555 3405 57575 3415
rect 57615 3405 57635 3415
rect 57675 3405 57695 3415
rect 57135 3390 57695 3405
rect 57735 3400 57755 3415
rect 58450 3400 58470 3415
rect 57735 3390 57790 3400
rect 57040 3370 57045 3390
rect 57065 3385 57095 3390
rect 57065 3370 57070 3385
rect 57040 3360 57070 3370
rect 57400 3370 57405 3390
rect 57425 3370 57430 3390
rect 57735 3385 57765 3390
rect 57400 3360 57430 3370
rect 57760 3370 57765 3385
rect 57785 3370 57790 3390
rect 57760 3360 57790 3370
rect 58415 3390 58470 3400
rect 58510 3405 58530 3415
rect 58570 3405 58590 3415
rect 58630 3405 58650 3415
rect 58690 3405 58710 3415
rect 58750 3405 58770 3415
rect 58810 3405 58830 3415
rect 58870 3405 58890 3415
rect 58930 3405 58950 3415
rect 58990 3405 59010 3415
rect 59050 3405 59070 3415
rect 58510 3390 59070 3405
rect 59110 3400 59130 3415
rect 59110 3390 59165 3400
rect 58415 3370 58420 3390
rect 58440 3385 58470 3390
rect 58440 3370 58445 3385
rect 58415 3360 58445 3370
rect 58775 3370 58780 3390
rect 58800 3370 58805 3390
rect 59110 3385 59140 3390
rect 58775 3360 58805 3370
rect 59135 3370 59140 3385
rect 59160 3370 59165 3390
rect 59135 3360 59165 3370
rect 55210 3290 55230 3360
rect 56375 3335 56395 3360
rect 57405 3335 57425 3360
rect 56365 3325 56405 3335
rect 56365 3305 56375 3325
rect 56395 3305 56405 3325
rect 56365 3295 56405 3305
rect 57395 3325 57435 3335
rect 57395 3305 57405 3325
rect 57425 3305 57435 3325
rect 57395 3295 57435 3305
rect 58780 3290 58800 3360
rect 55200 3280 55240 3290
rect 55200 3260 55210 3280
rect 55230 3260 55240 3280
rect 55200 3250 55240 3260
rect 58770 3280 58810 3290
rect 58770 3260 58780 3280
rect 58800 3260 58810 3280
rect 58770 3250 58810 3260
rect 56510 3010 56550 3020
rect 56510 2990 56520 3010
rect 56540 2995 56550 3010
rect 56840 3010 56880 3020
rect 56840 2995 56850 3010
rect 56540 2990 56565 2995
rect 56510 2980 56565 2990
rect 54745 2950 54775 2960
rect 54745 2930 54750 2950
rect 54770 2935 54775 2950
rect 55405 2950 55435 2960
rect 55405 2935 55410 2950
rect 54770 2930 54795 2935
rect 54745 2920 54795 2930
rect 55385 2930 55410 2935
rect 55430 2930 55435 2950
rect 55385 2920 55435 2930
rect 54780 2905 54795 2920
rect 54835 2905 54850 2920
rect 54890 2905 54905 2920
rect 54945 2905 54960 2920
rect 55000 2905 55015 2920
rect 55055 2905 55070 2920
rect 55110 2905 55125 2920
rect 55165 2905 55180 2920
rect 55220 2905 55235 2920
rect 55275 2905 55290 2920
rect 55330 2905 55345 2920
rect 55385 2905 55400 2920
rect 56550 2910 56565 2980
rect 56825 2990 56850 2995
rect 56870 2990 56880 3010
rect 56825 2980 56880 2990
rect 56920 3010 56960 3020
rect 56920 2990 56930 3010
rect 56950 2995 56960 3010
rect 57250 3010 57290 3020
rect 57250 2995 57260 3010
rect 56950 2990 56975 2995
rect 56920 2980 56975 2990
rect 56605 2910 56620 2925
rect 56660 2910 56675 2925
rect 56715 2910 56730 2925
rect 56770 2910 56785 2925
rect 56825 2910 56840 2980
rect 56960 2910 56975 2980
rect 57235 2990 57260 2995
rect 57280 2990 57290 3010
rect 57235 2980 57290 2990
rect 57015 2910 57030 2925
rect 57070 2910 57085 2925
rect 57125 2910 57140 2925
rect 57180 2910 57195 2925
rect 57235 2910 57250 2980
rect 58445 2950 58475 2960
rect 58445 2930 58450 2950
rect 58470 2935 58475 2950
rect 59105 2950 59135 2960
rect 59105 2935 59110 2950
rect 58470 2930 58495 2935
rect 58445 2920 58495 2930
rect 59085 2930 59110 2935
rect 59130 2930 59135 2950
rect 59085 2920 59135 2930
rect 58480 2905 58495 2920
rect 58535 2905 58550 2920
rect 58590 2905 58605 2920
rect 58645 2905 58660 2920
rect 58700 2905 58715 2920
rect 58755 2905 58770 2920
rect 58810 2905 58825 2920
rect 58865 2905 58880 2920
rect 58920 2905 58935 2920
rect 58975 2905 58990 2920
rect 59030 2905 59045 2920
rect 59085 2905 59100 2920
rect 56550 2645 56565 2660
rect 56605 2645 56620 2660
rect 56660 2650 56675 2660
rect 56715 2650 56730 2660
rect 56605 2635 56637 2645
rect 56660 2635 56730 2650
rect 56770 2645 56785 2660
rect 56825 2645 56840 2660
rect 56960 2645 56975 2660
rect 57015 2645 57030 2660
rect 57070 2650 57085 2660
rect 57125 2650 57140 2660
rect 56753 2635 56785 2645
rect 57015 2635 57047 2645
rect 57070 2635 57140 2650
rect 57180 2645 57195 2660
rect 57235 2645 57250 2660
rect 57163 2635 57195 2645
rect 56607 2615 56612 2635
rect 56632 2615 56637 2635
rect 56607 2605 56637 2615
rect 56675 2615 56685 2635
rect 56705 2615 56715 2635
rect 56675 2605 56715 2615
rect 56753 2615 56758 2635
rect 56778 2615 56783 2635
rect 56753 2605 56783 2615
rect 57017 2615 57022 2635
rect 57042 2615 57047 2635
rect 57017 2605 57047 2615
rect 57085 2615 57095 2635
rect 57115 2615 57125 2635
rect 57085 2605 57125 2615
rect 57163 2615 57168 2635
rect 57188 2615 57193 2635
rect 57163 2605 57193 2615
rect 56850 2360 56890 2370
rect 56850 2340 56860 2360
rect 56880 2340 56890 2360
rect 56850 2330 56935 2340
rect 56810 2315 56825 2330
rect 56865 2325 56935 2330
rect 56865 2315 56880 2325
rect 56920 2315 56935 2325
rect 56975 2315 56990 2330
rect 54780 2290 54795 2305
rect 54835 2295 54850 2305
rect 54890 2295 54905 2305
rect 54945 2295 54960 2305
rect 55000 2295 55015 2305
rect 55055 2295 55070 2305
rect 55110 2295 55125 2305
rect 55165 2295 55180 2305
rect 55220 2295 55235 2305
rect 55275 2295 55290 2305
rect 55330 2295 55345 2305
rect 54835 2280 55345 2295
rect 55385 2290 55400 2305
rect 55075 2260 55080 2280
rect 55100 2260 55105 2280
rect 55075 2225 55105 2260
rect 55070 2215 55110 2225
rect 55070 2195 55080 2215
rect 55100 2195 55110 2215
rect 55070 2175 55110 2195
rect 55070 2155 55080 2175
rect 55100 2155 55110 2175
rect 55070 2135 55110 2155
rect 55070 2115 55080 2135
rect 55100 2115 55110 2135
rect 55070 2105 55110 2115
rect 58480 2290 58495 2305
rect 58535 2295 58550 2305
rect 58590 2295 58605 2305
rect 58645 2295 58660 2305
rect 58700 2295 58715 2305
rect 58755 2295 58770 2305
rect 58810 2295 58825 2305
rect 58865 2295 58880 2305
rect 58920 2295 58935 2305
rect 58975 2295 58990 2305
rect 59030 2295 59045 2305
rect 58535 2280 59045 2295
rect 59085 2290 59100 2305
rect 58775 2260 58780 2280
rect 58800 2260 58805 2280
rect 58775 2225 58805 2260
rect 58770 2215 58810 2225
rect 58770 2195 58780 2215
rect 58800 2195 58810 2215
rect 58770 2175 58810 2195
rect 58770 2155 58780 2175
rect 58800 2155 58810 2175
rect 58770 2135 58810 2155
rect 58770 2115 58780 2135
rect 58800 2115 58810 2135
rect 58770 2105 58810 2115
rect 56810 2050 56825 2065
rect 56865 2050 56880 2065
rect 56920 2050 56935 2065
rect 56975 2050 56990 2065
rect 56770 2040 56825 2050
rect 56770 2020 56780 2040
rect 56800 2035 56825 2040
rect 56975 2040 57030 2050
rect 56975 2035 57000 2040
rect 56800 2020 56810 2035
rect 56770 2010 56810 2020
rect 56990 2020 57000 2035
rect 57020 2020 57030 2040
rect 56990 2010 57030 2020
rect 55995 1730 56025 1740
rect 55995 1710 56000 1730
rect 56020 1715 56025 1730
rect 56690 1730 56720 1740
rect 56690 1715 56695 1730
rect 56020 1710 56140 1715
rect 55995 1700 56140 1710
rect 54745 1675 54775 1685
rect 54745 1655 54750 1675
rect 54770 1660 54775 1675
rect 55405 1675 55435 1685
rect 55405 1660 55410 1675
rect 54770 1655 54795 1660
rect 54745 1645 54795 1655
rect 55385 1655 55410 1660
rect 55430 1655 55435 1675
rect 56125 1670 56140 1700
rect 56620 1710 56695 1715
rect 56715 1710 56720 1730
rect 56620 1700 56720 1710
rect 57080 1730 57110 1740
rect 57080 1710 57085 1730
rect 57105 1715 57110 1730
rect 57105 1710 57180 1715
rect 57080 1700 57180 1710
rect 56620 1670 56635 1700
rect 55385 1645 55435 1655
rect 56070 1645 56085 1660
rect 56125 1655 56635 1670
rect 57165 1670 57180 1700
rect 58445 1675 58475 1685
rect 56125 1645 56140 1655
rect 56180 1645 56195 1655
rect 56235 1645 56250 1655
rect 56290 1645 56305 1655
rect 56345 1645 56360 1655
rect 56400 1645 56415 1655
rect 56455 1645 56470 1655
rect 56510 1645 56525 1655
rect 56565 1645 56580 1655
rect 56620 1645 56635 1655
rect 56675 1645 56690 1660
rect 57110 1645 57125 1660
rect 57165 1655 57675 1670
rect 57165 1645 57180 1655
rect 57220 1645 57235 1655
rect 57275 1645 57290 1655
rect 57330 1645 57345 1655
rect 57385 1645 57400 1655
rect 57440 1645 57455 1655
rect 57495 1645 57510 1655
rect 57550 1645 57565 1655
rect 57605 1645 57620 1655
rect 57660 1645 57675 1655
rect 57715 1645 57730 1660
rect 58445 1655 58450 1675
rect 58470 1660 58475 1675
rect 59105 1675 59135 1685
rect 59105 1660 59110 1675
rect 58470 1655 58495 1660
rect 58445 1645 58495 1655
rect 59085 1655 59110 1660
rect 59130 1655 59135 1675
rect 59085 1645 59135 1655
rect 54780 1630 54795 1645
rect 54835 1630 54850 1645
rect 54890 1630 54905 1645
rect 54945 1630 54960 1645
rect 55000 1630 55015 1645
rect 55055 1630 55070 1645
rect 55110 1630 55125 1645
rect 55165 1630 55180 1645
rect 55220 1630 55235 1645
rect 55275 1630 55290 1645
rect 55330 1630 55345 1645
rect 55385 1630 55400 1645
rect 58480 1630 58495 1645
rect 58535 1630 58550 1645
rect 58590 1630 58605 1645
rect 58645 1630 58660 1645
rect 58700 1630 58715 1645
rect 58755 1630 58770 1645
rect 58810 1630 58825 1645
rect 58865 1630 58880 1645
rect 58920 1630 58935 1645
rect 58975 1630 58990 1645
rect 59030 1630 59045 1645
rect 59085 1630 59100 1645
rect 56070 1480 56085 1495
rect 56125 1480 56140 1495
rect 56180 1480 56195 1495
rect 56235 1480 56250 1495
rect 56290 1480 56305 1495
rect 56345 1480 56360 1495
rect 56400 1480 56415 1495
rect 56455 1480 56470 1495
rect 56510 1480 56525 1495
rect 56565 1480 56580 1495
rect 56620 1480 56635 1495
rect 56675 1480 56690 1495
rect 57110 1480 57125 1495
rect 57165 1480 57180 1495
rect 57220 1480 57235 1495
rect 57275 1480 57290 1495
rect 57330 1480 57345 1495
rect 57385 1480 57400 1495
rect 57440 1480 57455 1495
rect 57495 1480 57510 1495
rect 57550 1480 57565 1495
rect 57605 1480 57620 1495
rect 57660 1480 57675 1495
rect 57715 1480 57730 1495
rect 56035 1470 56085 1480
rect 56035 1450 56040 1470
rect 56060 1465 56085 1470
rect 56675 1470 56725 1480
rect 56675 1465 56700 1470
rect 56060 1450 56065 1465
rect 56035 1440 56065 1450
rect 56695 1450 56700 1465
rect 56720 1450 56725 1470
rect 56695 1440 56725 1450
rect 57075 1470 57125 1480
rect 57075 1450 57080 1470
rect 57100 1465 57125 1470
rect 57715 1470 57765 1480
rect 57715 1465 57740 1470
rect 57100 1450 57105 1465
rect 57075 1440 57105 1450
rect 57735 1450 57740 1465
rect 57760 1450 57765 1470
rect 57735 1440 57765 1450
rect 54780 1415 54795 1430
rect 54835 1420 54850 1430
rect 54890 1420 54905 1430
rect 54945 1420 54960 1430
rect 55000 1420 55015 1430
rect 55055 1420 55070 1430
rect 55110 1420 55125 1430
rect 55165 1420 55180 1430
rect 55220 1420 55235 1430
rect 55275 1420 55290 1430
rect 55330 1420 55345 1430
rect 54835 1405 55345 1420
rect 55385 1415 55400 1430
rect 58480 1415 58495 1430
rect 58535 1420 58550 1430
rect 58590 1420 58605 1430
rect 58645 1420 58660 1430
rect 58700 1420 58715 1430
rect 58755 1420 58770 1430
rect 58810 1420 58825 1430
rect 58865 1420 58880 1430
rect 58920 1420 58935 1430
rect 58975 1420 58990 1430
rect 59030 1420 59045 1430
rect 58535 1405 59045 1420
rect 59085 1415 59100 1430
rect 55240 1385 55245 1405
rect 55265 1385 55270 1405
rect 55240 1375 55270 1385
rect 58610 1385 58615 1405
rect 58635 1385 58640 1405
rect 58610 1375 58640 1385
rect 55245 1350 55265 1375
rect 58615 1350 58635 1375
rect 55235 1340 55275 1350
rect 55235 1320 55245 1340
rect 55265 1320 55275 1340
rect 55235 1300 55275 1320
rect 55235 1280 55245 1300
rect 55265 1280 55275 1300
rect 55235 1270 55275 1280
rect 58605 1340 58645 1350
rect 58605 1320 58615 1340
rect 58635 1320 58645 1340
rect 58605 1300 58645 1320
rect 58605 1280 58615 1300
rect 58635 1280 58645 1300
rect 58605 1270 58645 1280
rect 55245 1245 55265 1270
rect 58615 1245 58635 1270
rect 55240 1235 55270 1245
rect 55240 1215 55245 1235
rect 55265 1215 55270 1235
rect 58610 1235 58640 1245
rect 58610 1215 58615 1235
rect 58635 1215 58640 1235
rect 54780 1190 54795 1205
rect 54835 1200 55345 1215
rect 54835 1190 54850 1200
rect 54890 1190 54905 1200
rect 54945 1190 54960 1200
rect 55000 1190 55015 1200
rect 55055 1190 55070 1200
rect 55110 1190 55125 1200
rect 55165 1190 55180 1200
rect 55220 1190 55235 1200
rect 55275 1190 55290 1200
rect 55330 1190 55345 1200
rect 55385 1190 55400 1205
rect 58480 1190 58495 1205
rect 58535 1200 59045 1215
rect 58535 1190 58550 1200
rect 58590 1190 58605 1200
rect 58645 1190 58660 1200
rect 58700 1190 58715 1200
rect 58755 1190 58770 1200
rect 58810 1190 58825 1200
rect 58865 1190 58880 1200
rect 58920 1190 58935 1200
rect 58975 1190 58990 1200
rect 59030 1190 59045 1200
rect 59085 1190 59100 1205
rect 56690 1050 56720 1060
rect 56040 1040 56070 1050
rect 56040 1020 56045 1040
rect 56065 1025 56070 1040
rect 56690 1035 56695 1050
rect 56620 1030 56695 1035
rect 56715 1030 56720 1050
rect 56065 1020 56140 1025
rect 56040 1010 56140 1020
rect 56125 995 56140 1010
rect 56620 1020 56720 1030
rect 56840 1050 56870 1060
rect 56840 1030 56845 1050
rect 56865 1035 56870 1050
rect 56930 1050 56960 1060
rect 56930 1035 56935 1050
rect 56865 1030 56880 1035
rect 56840 1020 56880 1030
rect 56620 995 56635 1020
rect 56070 970 56085 985
rect 56125 980 56635 995
rect 56125 970 56140 980
rect 56180 970 56195 980
rect 56235 970 56250 980
rect 56290 970 56305 980
rect 56345 970 56360 980
rect 56400 970 56415 980
rect 56455 970 56470 980
rect 56510 970 56525 980
rect 56565 970 56580 980
rect 56620 970 56635 980
rect 56675 970 56690 985
rect 56810 970 56825 985
rect 56865 970 56880 1020
rect 56920 1030 56935 1035
rect 56955 1030 56960 1050
rect 56920 1020 56960 1030
rect 57080 1050 57110 1060
rect 57080 1030 57085 1050
rect 57105 1035 57110 1050
rect 57730 1040 57760 1050
rect 57105 1030 57180 1035
rect 57080 1020 57180 1030
rect 57730 1025 57735 1040
rect 56920 970 56935 1020
rect 57165 995 57180 1020
rect 57660 1020 57735 1025
rect 57755 1020 57760 1040
rect 57660 1010 57760 1020
rect 57660 995 57675 1010
rect 56975 970 56990 985
rect 57110 970 57125 985
rect 57165 980 57675 995
rect 57165 970 57180 980
rect 57220 970 57235 980
rect 57275 970 57290 980
rect 57330 970 57345 980
rect 57385 970 57400 980
rect 57440 970 57455 980
rect 57495 970 57510 980
rect 57550 970 57565 980
rect 57605 970 57620 980
rect 57660 970 57675 980
rect 57715 970 57730 985
rect 54780 875 54795 890
rect 54835 875 54850 890
rect 54890 875 54905 890
rect 54945 875 54960 890
rect 55000 875 55015 890
rect 55055 875 55070 890
rect 55110 875 55125 890
rect 55165 875 55180 890
rect 55220 875 55235 890
rect 55275 875 55290 890
rect 55330 875 55345 890
rect 55385 875 55400 890
rect 54745 865 54795 875
rect 54745 845 54750 865
rect 54770 860 54795 865
rect 55385 865 55435 875
rect 55385 860 55410 865
rect 54770 845 54775 860
rect 54745 830 54775 845
rect 55405 845 55410 860
rect 55430 845 55435 865
rect 55405 830 55435 845
rect 58480 875 58495 890
rect 58535 875 58550 890
rect 58590 875 58605 890
rect 58645 875 58660 890
rect 58700 875 58715 890
rect 58755 875 58770 890
rect 58810 875 58825 890
rect 58865 875 58880 890
rect 58920 875 58935 890
rect 58975 875 58990 890
rect 59030 875 59045 890
rect 59085 875 59100 890
rect 58445 865 58495 875
rect 58445 845 58450 865
rect 58470 860 58495 865
rect 59085 865 59135 875
rect 59085 860 59110 865
rect 58470 845 58475 860
rect 58445 830 58475 845
rect 59105 845 59110 860
rect 59130 845 59135 865
rect 59105 835 59135 845
rect 56070 805 56085 820
rect 56125 805 56140 820
rect 56180 805 56195 820
rect 56235 805 56250 820
rect 56290 805 56305 820
rect 56345 805 56360 820
rect 56400 805 56415 820
rect 56455 805 56470 820
rect 56510 805 56525 820
rect 56565 805 56580 820
rect 56620 805 56635 820
rect 56675 805 56690 820
rect 56810 805 56825 820
rect 56865 805 56880 820
rect 56920 805 56935 820
rect 56975 805 56990 820
rect 57110 805 57125 820
rect 57165 805 57180 820
rect 57220 805 57235 820
rect 57275 805 57290 820
rect 57330 805 57345 820
rect 57385 805 57400 820
rect 57440 805 57455 820
rect 57495 805 57510 820
rect 57550 805 57565 820
rect 57605 805 57620 820
rect 57660 805 57675 820
rect 57715 805 57730 820
rect 56035 795 56085 805
rect 56035 775 56040 795
rect 56060 790 56085 795
rect 56675 795 56825 805
rect 56675 790 56740 795
rect 56060 775 56065 790
rect 56035 765 56065 775
rect 56735 775 56740 790
rect 56760 790 56825 795
rect 56975 795 57125 805
rect 56975 790 57040 795
rect 56760 775 56765 790
rect 56735 765 56765 775
rect 57035 775 57040 790
rect 57060 790 57125 795
rect 57715 795 57765 805
rect 57715 790 57740 795
rect 57060 775 57065 790
rect 57035 765 57065 775
rect 57735 775 57740 790
rect 57760 775 57765 795
rect 57735 765 57765 775
rect 55100 505 55140 515
rect 55100 485 55110 505
rect 55130 485 55140 505
rect 55100 475 55140 485
rect 58580 505 58620 515
rect 58580 485 58590 505
rect 58610 485 58620 505
rect 58580 475 58620 485
rect 55110 205 55130 475
rect 56825 375 56865 385
rect 56825 355 56835 375
rect 56855 355 56865 375
rect 56935 375 56975 385
rect 56935 355 56945 375
rect 56965 355 56975 375
rect 56260 330 56275 345
rect 56315 340 57375 355
rect 56315 330 56330 340
rect 56370 330 56385 340
rect 56425 330 56440 340
rect 56480 330 56495 340
rect 56535 330 56550 340
rect 56590 330 56605 340
rect 56645 330 56660 340
rect 56700 330 56715 340
rect 56755 330 56770 340
rect 56810 330 56825 340
rect 56865 330 56880 340
rect 56920 330 56935 340
rect 56975 330 56990 340
rect 57030 330 57045 340
rect 57085 330 57100 340
rect 57140 330 57155 340
rect 57195 330 57210 340
rect 57250 330 57265 340
rect 57305 330 57320 340
rect 57360 330 57375 340
rect 57415 330 57430 345
rect 57470 330 57485 345
rect 54790 180 54850 195
rect 54890 190 55250 205
rect 54890 180 54950 190
rect 54990 180 55050 190
rect 55090 180 55150 190
rect 55190 180 55250 190
rect 55290 180 55350 195
rect 58590 205 58610 475
rect 58370 180 58430 195
rect 58470 190 58830 205
rect 58470 180 58530 190
rect 58570 180 58630 190
rect 58670 180 58730 190
rect 58770 180 58830 190
rect 58870 180 58930 195
rect 56260 65 56275 80
rect 56315 65 56330 80
rect 56370 65 56385 80
rect 56425 65 56440 80
rect 56480 65 56495 80
rect 56535 65 56550 80
rect 56590 65 56605 80
rect 56645 65 56660 80
rect 56700 65 56715 80
rect 56755 65 56770 80
rect 56810 65 56825 80
rect 56865 65 56880 80
rect 56920 65 56935 80
rect 56975 65 56990 80
rect 57030 65 57045 80
rect 57085 65 57100 80
rect 57140 65 57155 80
rect 57195 65 57210 80
rect 57250 65 57265 80
rect 57305 65 57320 80
rect 57360 65 57375 80
rect 56220 55 56275 65
rect 56220 35 56230 55
rect 56250 50 56275 55
rect 56250 35 56260 50
rect 56220 25 56260 35
rect 57415 -35 57430 80
rect 57470 65 57485 80
rect 57470 55 57525 65
rect 57470 50 57495 55
rect 57485 35 57495 50
rect 57515 35 57525 55
rect 57485 25 57525 35
rect 57415 -45 57455 -35
rect 57415 -65 57425 -45
rect 57445 -65 57455 -45
rect 57415 -75 57455 -65
rect 56595 -280 56635 -270
rect 56595 -300 56605 -280
rect 56625 -300 56635 -280
rect 57040 -280 57080 -270
rect 57040 -300 57050 -280
rect 57070 -300 57080 -280
rect 56470 -325 56485 -310
rect 56525 -315 56705 -300
rect 57040 -310 57080 -300
rect 56525 -325 56540 -315
rect 56580 -325 56595 -315
rect 56635 -325 56650 -315
rect 56690 -325 56705 -315
rect 56745 -325 56760 -310
rect 56910 -325 57210 -310
rect 56470 -490 56485 -475
rect 56525 -490 56540 -475
rect 56580 -490 56595 -475
rect 56635 -490 56650 -475
rect 56690 -490 56705 -475
rect 56745 -490 56760 -475
rect 56910 -490 57210 -475
rect 56435 -500 56485 -490
rect 56435 -520 56440 -500
rect 56460 -505 56485 -500
rect 56745 -500 56795 -490
rect 56745 -505 56770 -500
rect 56460 -520 56465 -505
rect 54790 -535 54850 -520
rect 54890 -535 54950 -520
rect 54990 -535 55050 -520
rect 55090 -535 55150 -520
rect 55190 -535 55250 -520
rect 55290 -535 55350 -520
rect 56435 -530 56465 -520
rect 56765 -520 56770 -505
rect 56790 -520 56795 -500
rect 56765 -530 56795 -520
rect 58370 -535 58430 -520
rect 58470 -535 58530 -520
rect 58570 -535 58630 -520
rect 58670 -535 58730 -520
rect 58770 -535 58830 -520
rect 58870 -535 58930 -520
rect 54755 -545 54850 -535
rect 54755 -565 54760 -545
rect 54780 -550 54850 -545
rect 55290 -545 55385 -535
rect 55290 -550 55360 -545
rect 54780 -565 54785 -550
rect 54755 -575 54785 -565
rect 55355 -565 55360 -550
rect 55380 -565 55385 -545
rect 55355 -575 55385 -565
rect 58335 -545 58430 -535
rect 58335 -565 58340 -545
rect 58360 -550 58430 -545
rect 58870 -545 58965 -535
rect 58870 -550 58940 -545
rect 58360 -565 58365 -550
rect 58335 -575 58365 -565
rect 58935 -565 58940 -550
rect 58960 -565 58965 -545
rect 58935 -575 58965 -565
<< polycont >>
rect 56095 4905 56115 4925
rect 56275 4905 56295 4925
rect 57035 4905 57055 4925
rect 57215 4905 57235 4925
rect 57505 4905 57525 4925
rect 57685 4905 57705 4925
rect 56565 4735 56585 4755
rect 56745 4735 56765 4755
rect 56160 4455 56180 4475
rect 56635 4455 56655 4475
rect 57145 4455 57165 4475
rect 57581 4445 57601 4465
rect 54850 3370 54870 3390
rect 55210 3370 55230 3390
rect 55570 3370 55590 3390
rect 56015 3370 56035 3390
rect 56375 3370 56395 3390
rect 56735 3370 56755 3390
rect 57045 3370 57065 3390
rect 57405 3370 57425 3390
rect 57765 3370 57785 3390
rect 58420 3370 58440 3390
rect 58780 3370 58800 3390
rect 59140 3370 59160 3390
rect 56375 3305 56395 3325
rect 57405 3305 57425 3325
rect 55210 3260 55230 3280
rect 58780 3260 58800 3280
rect 56520 2990 56540 3010
rect 54750 2930 54770 2950
rect 55410 2930 55430 2950
rect 56850 2990 56870 3010
rect 56930 2990 56950 3010
rect 57260 2990 57280 3010
rect 58450 2930 58470 2950
rect 59110 2930 59130 2950
rect 56612 2615 56632 2635
rect 56685 2615 56705 2635
rect 56758 2615 56778 2635
rect 57022 2615 57042 2635
rect 57095 2615 57115 2635
rect 57168 2615 57188 2635
rect 56860 2340 56880 2360
rect 55080 2260 55100 2280
rect 55080 2195 55100 2215
rect 55080 2155 55100 2175
rect 55080 2115 55100 2135
rect 58780 2260 58800 2280
rect 58780 2195 58800 2215
rect 58780 2155 58800 2175
rect 58780 2115 58800 2135
rect 56780 2020 56800 2040
rect 57000 2020 57020 2040
rect 56000 1710 56020 1730
rect 54750 1655 54770 1675
rect 55410 1655 55430 1675
rect 56695 1710 56715 1730
rect 57085 1710 57105 1730
rect 58450 1655 58470 1675
rect 59110 1655 59130 1675
rect 56040 1450 56060 1470
rect 56700 1450 56720 1470
rect 57080 1450 57100 1470
rect 57740 1450 57760 1470
rect 55245 1385 55265 1405
rect 58615 1385 58635 1405
rect 55245 1320 55265 1340
rect 55245 1280 55265 1300
rect 58615 1320 58635 1340
rect 58615 1280 58635 1300
rect 55245 1215 55265 1235
rect 58615 1215 58635 1235
rect 56045 1020 56065 1040
rect 56695 1030 56715 1050
rect 56845 1030 56865 1050
rect 56935 1030 56955 1050
rect 57085 1030 57105 1050
rect 57735 1020 57755 1040
rect 54750 845 54770 865
rect 55410 845 55430 865
rect 58450 845 58470 865
rect 59110 845 59130 865
rect 56040 775 56060 795
rect 56740 775 56760 795
rect 57040 775 57060 795
rect 57740 775 57760 795
rect 55110 485 55130 505
rect 58590 485 58610 505
rect 56835 355 56855 375
rect 56945 355 56965 375
rect 56230 35 56250 55
rect 57495 35 57515 55
rect 57425 -65 57445 -45
rect 56605 -300 56625 -280
rect 57050 -300 57070 -280
rect 56440 -520 56460 -500
rect 56770 -520 56790 -500
rect 54760 -565 54780 -545
rect 55360 -565 55380 -545
rect 58340 -565 58360 -545
rect 58940 -565 58960 -545
<< xpolycontact >>
rect 54124 2790 54265 3010
rect 54124 2445 54265 2665
rect 59805 2705 59946 2925
rect 59805 2360 59946 2580
rect 54380 1294 54415 1514
rect 54380 915 54415 1135
rect 54440 1294 54475 1514
rect 54440 915 54475 1135
rect 54500 1294 54535 1514
rect 54500 915 54535 1135
rect 54560 1294 54595 1514
rect 59475 1294 59510 1514
rect 54560 915 54595 1135
rect 59475 915 59510 1135
rect 59535 1294 59570 1514
rect 59535 915 59570 1135
rect 59595 1294 59630 1514
rect 59595 915 59630 1135
rect 59655 1294 59690 1514
rect 59655 915 59690 1135
rect 54520 -85 54555 135
rect 54520 -552 54555 -332
rect 54580 -85 54615 135
rect 54580 -552 54615 -332
rect 59455 -85 59490 135
rect 59455 -552 59490 -332
rect 59515 -85 59550 135
rect 59515 -552 59550 -332
<< ppolyres >>
rect 54124 2665 54265 2790
rect 59805 2580 59946 2705
<< xpolyres >>
rect 54380 1135 54415 1294
rect 54440 1135 54475 1294
rect 54500 1135 54535 1294
rect 54560 1135 54595 1294
rect 59475 1135 59510 1294
rect 59535 1135 59570 1294
rect 59595 1135 59630 1294
rect 59655 1135 59690 1294
rect 54520 -332 54555 -85
rect 54580 -332 54615 -85
rect 59455 -332 59490 -85
rect 59515 -332 59550 -85
<< locali >>
rect 56085 4925 56125 4935
rect 56085 4905 56095 4925
rect 56115 4905 56125 4925
rect 56085 4895 56125 4905
rect 56265 4925 56305 4935
rect 56265 4905 56275 4925
rect 56295 4905 56305 4925
rect 56265 4895 56305 4905
rect 57025 4925 57065 4935
rect 57025 4905 57035 4925
rect 57055 4905 57065 4925
rect 57025 4895 57065 4905
rect 57205 4925 57245 4935
rect 57205 4905 57215 4925
rect 57235 4905 57245 4925
rect 57205 4895 57245 4905
rect 57495 4925 57535 4935
rect 57495 4905 57505 4925
rect 57525 4905 57535 4925
rect 57495 4895 57535 4905
rect 57675 4925 57715 4935
rect 57675 4905 57685 4925
rect 57705 4905 57715 4925
rect 57675 4895 57715 4905
rect 56050 4865 56120 4875
rect 56050 4545 56055 4865
rect 56075 4545 56095 4865
rect 56115 4545 56120 4865
rect 56050 4535 56120 4545
rect 56150 4865 56180 4875
rect 56150 4545 56155 4865
rect 56175 4545 56180 4865
rect 56150 4535 56180 4545
rect 56210 4865 56240 4875
rect 56210 4545 56215 4865
rect 56235 4545 56240 4865
rect 56210 4535 56240 4545
rect 56270 4865 56340 4875
rect 56270 4545 56275 4865
rect 56295 4545 56315 4865
rect 56335 4545 56340 4865
rect 56990 4865 57060 4875
rect 56555 4755 56595 4765
rect 56555 4735 56565 4755
rect 56585 4735 56595 4755
rect 56555 4725 56595 4735
rect 56735 4755 56775 4765
rect 56735 4735 56745 4755
rect 56765 4735 56775 4755
rect 56735 4725 56775 4735
rect 56270 4535 56340 4545
rect 56520 4695 56590 4705
rect 56520 4545 56525 4695
rect 56545 4545 56565 4695
rect 56585 4545 56590 4695
rect 56520 4535 56590 4545
rect 56620 4695 56650 4705
rect 56620 4545 56625 4695
rect 56645 4545 56650 4695
rect 56620 4535 56650 4545
rect 56680 4695 56710 4705
rect 56680 4545 56685 4695
rect 56705 4545 56710 4695
rect 56680 4535 56710 4545
rect 56740 4695 56810 4705
rect 56740 4545 56745 4695
rect 56765 4545 56785 4695
rect 56805 4545 56810 4695
rect 56740 4535 56810 4545
rect 56990 4545 56995 4865
rect 57015 4545 57035 4865
rect 57055 4545 57060 4865
rect 56990 4535 57060 4545
rect 57090 4865 57120 4875
rect 57090 4545 57095 4865
rect 57115 4545 57120 4865
rect 57090 4535 57120 4545
rect 57150 4865 57180 4875
rect 57150 4545 57155 4865
rect 57175 4545 57180 4865
rect 57150 4535 57180 4545
rect 57210 4865 57280 4875
rect 57210 4545 57215 4865
rect 57235 4545 57255 4865
rect 57275 4545 57280 4865
rect 57210 4535 57280 4545
rect 57460 4865 57530 4875
rect 57460 4545 57465 4865
rect 57485 4545 57505 4865
rect 57525 4545 57530 4865
rect 57460 4535 57530 4545
rect 57560 4865 57590 4875
rect 57560 4545 57565 4865
rect 57585 4545 57590 4865
rect 57560 4535 57590 4545
rect 57620 4865 57650 4875
rect 57620 4545 57625 4865
rect 57645 4545 57650 4865
rect 57620 4535 57650 4545
rect 57680 4865 57750 4875
rect 57680 4545 57685 4865
rect 57705 4545 57725 4865
rect 57745 4545 57750 4865
rect 57680 4535 57750 4545
rect 56150 4475 56190 4485
rect 56150 4455 56160 4475
rect 56180 4455 56190 4475
rect 56150 4445 56190 4455
rect 56630 4475 56660 4485
rect 56630 4455 56635 4475
rect 56655 4455 56660 4475
rect 56630 4445 56660 4455
rect 57140 4475 57170 4485
rect 57140 4455 57145 4475
rect 57165 4455 57170 4475
rect 57140 4445 57170 4455
rect 57576 4465 57606 4475
rect 57576 4445 57581 4465
rect 57601 4445 57606 4465
rect 57576 4435 57606 4445
rect 54805 3750 54875 3760
rect 54805 3430 54810 3750
rect 54830 3430 54850 3750
rect 54870 3430 54875 3750
rect 54805 3420 54875 3430
rect 54905 3750 54935 3760
rect 54905 3430 54910 3750
rect 54930 3430 54935 3750
rect 54905 3420 54935 3430
rect 54965 3750 54995 3760
rect 54965 3430 54970 3750
rect 54990 3430 54995 3750
rect 54965 3420 54995 3430
rect 55025 3750 55055 3760
rect 55025 3430 55030 3750
rect 55050 3430 55055 3750
rect 55025 3420 55055 3430
rect 55085 3750 55115 3760
rect 55085 3430 55090 3750
rect 55110 3430 55115 3750
rect 55085 3420 55115 3430
rect 55145 3750 55175 3760
rect 55145 3430 55150 3750
rect 55170 3430 55175 3750
rect 55145 3420 55175 3430
rect 55205 3750 55235 3760
rect 55205 3430 55210 3750
rect 55230 3430 55235 3750
rect 55205 3420 55235 3430
rect 55265 3750 55295 3760
rect 55265 3430 55270 3750
rect 55290 3430 55295 3750
rect 55265 3420 55295 3430
rect 55325 3750 55355 3760
rect 55325 3430 55330 3750
rect 55350 3430 55355 3750
rect 55325 3420 55355 3430
rect 55385 3750 55415 3760
rect 55385 3430 55390 3750
rect 55410 3430 55415 3750
rect 55385 3420 55415 3430
rect 55445 3750 55475 3760
rect 55445 3430 55450 3750
rect 55470 3430 55475 3750
rect 55445 3420 55475 3430
rect 55505 3750 55535 3760
rect 55505 3430 55510 3750
rect 55530 3430 55535 3750
rect 55505 3420 55535 3430
rect 55565 3750 55635 3760
rect 55565 3430 55570 3750
rect 55590 3430 55610 3750
rect 55630 3430 55635 3750
rect 55565 3420 55635 3430
rect 55970 3750 56040 3760
rect 55970 3430 55975 3750
rect 55995 3430 56015 3750
rect 56035 3430 56040 3750
rect 55970 3420 56040 3430
rect 56070 3750 56100 3760
rect 56070 3430 56075 3750
rect 56095 3430 56100 3750
rect 56070 3420 56100 3430
rect 56130 3750 56160 3760
rect 56130 3430 56135 3750
rect 56155 3430 56160 3750
rect 56130 3420 56160 3430
rect 56190 3750 56220 3760
rect 56190 3430 56195 3750
rect 56215 3430 56220 3750
rect 56190 3420 56220 3430
rect 56250 3750 56280 3760
rect 56250 3430 56255 3750
rect 56275 3430 56280 3750
rect 56250 3420 56280 3430
rect 56310 3750 56340 3760
rect 56310 3430 56315 3750
rect 56335 3430 56340 3750
rect 56310 3420 56340 3430
rect 56370 3750 56400 3760
rect 56370 3430 56375 3750
rect 56395 3430 56400 3750
rect 56370 3420 56400 3430
rect 56430 3750 56460 3760
rect 56430 3430 56435 3750
rect 56455 3430 56460 3750
rect 56430 3420 56460 3430
rect 56490 3750 56520 3760
rect 56490 3430 56495 3750
rect 56515 3430 56520 3750
rect 56490 3420 56520 3430
rect 56550 3750 56580 3760
rect 56550 3430 56555 3750
rect 56575 3430 56580 3750
rect 56550 3420 56580 3430
rect 56610 3750 56640 3760
rect 56610 3430 56615 3750
rect 56635 3430 56640 3750
rect 56610 3420 56640 3430
rect 56670 3750 56700 3760
rect 56670 3430 56675 3750
rect 56695 3430 56700 3750
rect 56670 3420 56700 3430
rect 56730 3750 56800 3760
rect 56730 3430 56735 3750
rect 56755 3430 56775 3750
rect 56795 3430 56800 3750
rect 56730 3420 56800 3430
rect 57000 3750 57070 3760
rect 57000 3430 57005 3750
rect 57025 3430 57045 3750
rect 57065 3430 57070 3750
rect 57000 3420 57070 3430
rect 57100 3750 57130 3760
rect 57100 3430 57105 3750
rect 57125 3430 57130 3750
rect 57100 3420 57130 3430
rect 57160 3750 57190 3760
rect 57160 3430 57165 3750
rect 57185 3430 57190 3750
rect 57160 3420 57190 3430
rect 57220 3750 57250 3760
rect 57220 3430 57225 3750
rect 57245 3430 57250 3750
rect 57220 3420 57250 3430
rect 57280 3750 57310 3760
rect 57280 3430 57285 3750
rect 57305 3430 57310 3750
rect 57280 3420 57310 3430
rect 57340 3750 57370 3760
rect 57340 3430 57345 3750
rect 57365 3430 57370 3750
rect 57340 3420 57370 3430
rect 57400 3750 57430 3760
rect 57400 3430 57405 3750
rect 57425 3430 57430 3750
rect 57400 3420 57430 3430
rect 57460 3750 57490 3760
rect 57460 3430 57465 3750
rect 57485 3430 57490 3750
rect 57460 3420 57490 3430
rect 57520 3750 57550 3760
rect 57520 3430 57525 3750
rect 57545 3430 57550 3750
rect 57520 3420 57550 3430
rect 57580 3750 57610 3760
rect 57580 3430 57585 3750
rect 57605 3430 57610 3750
rect 57580 3420 57610 3430
rect 57640 3750 57670 3760
rect 57640 3430 57645 3750
rect 57665 3430 57670 3750
rect 57640 3420 57670 3430
rect 57700 3750 57730 3760
rect 57700 3430 57705 3750
rect 57725 3430 57730 3750
rect 57700 3420 57730 3430
rect 57760 3750 57830 3760
rect 57760 3430 57765 3750
rect 57785 3430 57805 3750
rect 57825 3430 57830 3750
rect 57760 3420 57830 3430
rect 58375 3750 58445 3760
rect 58375 3430 58380 3750
rect 58400 3430 58420 3750
rect 58440 3430 58445 3750
rect 58375 3420 58445 3430
rect 58475 3750 58505 3760
rect 58475 3430 58480 3750
rect 58500 3430 58505 3750
rect 58475 3420 58505 3430
rect 58535 3750 58565 3760
rect 58535 3430 58540 3750
rect 58560 3430 58565 3750
rect 58535 3420 58565 3430
rect 58595 3750 58625 3760
rect 58595 3430 58600 3750
rect 58620 3430 58625 3750
rect 58595 3420 58625 3430
rect 58655 3750 58685 3760
rect 58655 3430 58660 3750
rect 58680 3430 58685 3750
rect 58655 3420 58685 3430
rect 58715 3750 58745 3760
rect 58715 3430 58720 3750
rect 58740 3430 58745 3750
rect 58715 3420 58745 3430
rect 58775 3750 58805 3760
rect 58775 3430 58780 3750
rect 58800 3430 58805 3750
rect 58775 3420 58805 3430
rect 58835 3750 58865 3760
rect 58835 3430 58840 3750
rect 58860 3430 58865 3750
rect 58835 3420 58865 3430
rect 58895 3750 58925 3760
rect 58895 3430 58900 3750
rect 58920 3430 58925 3750
rect 58895 3420 58925 3430
rect 58955 3750 58985 3760
rect 58955 3430 58960 3750
rect 58980 3430 58985 3750
rect 58955 3420 58985 3430
rect 59015 3750 59045 3760
rect 59015 3430 59020 3750
rect 59040 3430 59045 3750
rect 59015 3420 59045 3430
rect 59075 3750 59105 3760
rect 59075 3430 59080 3750
rect 59100 3430 59105 3750
rect 59075 3420 59105 3430
rect 59135 3750 59205 3760
rect 59135 3430 59140 3750
rect 59160 3430 59180 3750
rect 59200 3430 59205 3750
rect 59135 3420 59205 3430
rect 54845 3390 54875 3400
rect 54845 3370 54850 3390
rect 54870 3370 54875 3390
rect 54845 3360 54875 3370
rect 55205 3390 55235 3400
rect 55205 3370 55210 3390
rect 55230 3370 55235 3390
rect 55205 3360 55235 3370
rect 55565 3390 55595 3400
rect 55565 3370 55570 3390
rect 55590 3370 55595 3390
rect 55565 3360 55595 3370
rect 56010 3390 56040 3400
rect 56010 3370 56015 3390
rect 56035 3370 56040 3390
rect 56010 3360 56040 3370
rect 56370 3390 56400 3400
rect 56370 3370 56375 3390
rect 56395 3370 56400 3390
rect 56370 3360 56400 3370
rect 56730 3390 56760 3400
rect 56730 3370 56735 3390
rect 56755 3370 56760 3390
rect 56730 3360 56760 3370
rect 57040 3390 57070 3400
rect 57040 3370 57045 3390
rect 57065 3370 57070 3390
rect 57040 3360 57070 3370
rect 57400 3390 57430 3400
rect 57400 3370 57405 3390
rect 57425 3370 57430 3390
rect 57400 3360 57430 3370
rect 57760 3390 57790 3400
rect 57760 3370 57765 3390
rect 57785 3370 57790 3390
rect 57760 3360 57790 3370
rect 58415 3390 58445 3400
rect 58415 3370 58420 3390
rect 58440 3370 58445 3390
rect 58415 3360 58445 3370
rect 58775 3390 58805 3400
rect 58775 3370 58780 3390
rect 58800 3370 58805 3390
rect 58775 3360 58805 3370
rect 59135 3390 59165 3400
rect 59135 3370 59140 3390
rect 59160 3370 59165 3390
rect 59135 3360 59165 3370
rect 56365 3325 56405 3335
rect 56365 3305 56375 3325
rect 56395 3305 56405 3325
rect 56365 3295 56405 3305
rect 57395 3325 57435 3335
rect 57395 3305 57405 3325
rect 57425 3305 57435 3325
rect 57395 3295 57435 3305
rect 55200 3280 55240 3290
rect 55200 3260 55210 3280
rect 55230 3260 55240 3280
rect 55200 3250 55240 3260
rect 58770 3280 58810 3290
rect 58770 3260 58780 3280
rect 58800 3260 58810 3280
rect 58770 3250 58810 3260
rect 54124 3040 54265 3050
rect 54124 3020 54130 3040
rect 54150 3020 54185 3040
rect 54205 3020 54240 3040
rect 54260 3020 54265 3040
rect 54124 3010 54265 3020
rect 56510 3010 56550 3020
rect 56510 2990 56520 3010
rect 56540 2990 56550 3010
rect 56510 2980 56550 2990
rect 56680 3010 56710 3020
rect 56680 2990 56685 3010
rect 56705 2990 56710 3010
rect 56680 2980 56710 2990
rect 56840 3010 56880 3020
rect 56840 2990 56850 3010
rect 56870 2990 56880 3010
rect 56840 2980 56880 2990
rect 56920 3010 56960 3020
rect 56920 2990 56930 3010
rect 56950 2990 56960 3010
rect 56920 2980 56960 2990
rect 57090 3010 57120 3020
rect 57090 2990 57095 3010
rect 57115 2990 57120 3010
rect 57090 2980 57120 2990
rect 57250 3010 57290 3020
rect 57250 2990 57260 3010
rect 57280 2990 57290 3010
rect 57250 2980 57290 2990
rect 54745 2950 54775 2960
rect 54745 2930 54750 2950
rect 54770 2930 54775 2950
rect 54745 2920 54775 2930
rect 55405 2950 55435 2960
rect 55405 2930 55410 2950
rect 55430 2930 55435 2950
rect 55405 2920 55435 2930
rect 56520 2905 56540 2980
rect 56620 2955 56660 2965
rect 56620 2935 56630 2955
rect 56650 2935 56660 2955
rect 56620 2925 56660 2935
rect 56630 2905 56650 2925
rect 56685 2905 56705 2980
rect 56730 2955 56770 2965
rect 56730 2935 56740 2955
rect 56760 2935 56770 2955
rect 56730 2925 56770 2935
rect 56740 2905 56760 2925
rect 56850 2905 56870 2980
rect 56930 2905 56950 2980
rect 57030 2955 57070 2965
rect 57030 2935 57040 2955
rect 57060 2935 57070 2955
rect 57030 2925 57070 2935
rect 57040 2905 57060 2925
rect 57095 2905 57115 2980
rect 57140 2955 57180 2965
rect 57140 2935 57150 2955
rect 57170 2935 57180 2955
rect 57140 2925 57180 2935
rect 57150 2905 57170 2925
rect 57260 2905 57280 2980
rect 58445 2950 58475 2960
rect 58445 2930 58450 2950
rect 58470 2930 58475 2950
rect 58445 2920 58475 2930
rect 59105 2950 59135 2960
rect 59105 2930 59110 2950
rect 59130 2930 59135 2950
rect 59105 2920 59135 2930
rect 59805 2955 59946 2965
rect 59805 2935 59810 2955
rect 59830 2935 59865 2955
rect 59885 2935 59920 2955
rect 59940 2935 59946 2955
rect 59805 2925 59946 2935
rect 54705 2890 54775 2900
rect 54124 2435 54265 2445
rect 54124 2415 54130 2435
rect 54150 2415 54185 2435
rect 54205 2415 54240 2435
rect 54260 2415 54265 2435
rect 54124 2405 54265 2415
rect 54705 2320 54710 2890
rect 54730 2320 54750 2890
rect 54770 2320 54775 2890
rect 54705 2310 54775 2320
rect 54800 2890 54830 2900
rect 54800 2320 54805 2890
rect 54825 2320 54830 2890
rect 54800 2310 54830 2320
rect 54855 2890 54885 2900
rect 54855 2320 54860 2890
rect 54880 2320 54885 2890
rect 54855 2310 54885 2320
rect 54910 2890 54940 2900
rect 54910 2320 54915 2890
rect 54935 2320 54940 2890
rect 54910 2310 54940 2320
rect 54965 2890 54995 2900
rect 54965 2320 54970 2890
rect 54990 2320 54995 2890
rect 54965 2310 54995 2320
rect 55020 2890 55050 2900
rect 55020 2320 55025 2890
rect 55045 2320 55050 2890
rect 55020 2310 55050 2320
rect 55075 2890 55105 2900
rect 55075 2320 55080 2890
rect 55100 2320 55105 2890
rect 55075 2310 55105 2320
rect 55130 2890 55160 2900
rect 55130 2320 55135 2890
rect 55155 2320 55160 2890
rect 55130 2310 55160 2320
rect 55185 2890 55215 2900
rect 55185 2320 55190 2890
rect 55210 2320 55215 2890
rect 55185 2310 55215 2320
rect 55240 2890 55270 2900
rect 55240 2320 55245 2890
rect 55265 2320 55270 2890
rect 55240 2310 55270 2320
rect 55295 2890 55325 2900
rect 55295 2320 55300 2890
rect 55320 2320 55325 2890
rect 55295 2310 55325 2320
rect 55350 2890 55380 2900
rect 55350 2320 55355 2890
rect 55375 2320 55380 2890
rect 55350 2310 55380 2320
rect 55405 2890 55475 2900
rect 55405 2320 55410 2890
rect 55430 2320 55450 2890
rect 55470 2320 55475 2890
rect 56475 2895 56545 2905
rect 56475 2875 56480 2895
rect 56500 2875 56520 2895
rect 56540 2875 56545 2895
rect 56475 2845 56545 2875
rect 56475 2825 56480 2845
rect 56500 2825 56520 2845
rect 56540 2825 56545 2845
rect 56475 2795 56545 2825
rect 56475 2775 56480 2795
rect 56500 2775 56520 2795
rect 56540 2775 56545 2795
rect 56475 2745 56545 2775
rect 56475 2725 56480 2745
rect 56500 2725 56520 2745
rect 56540 2725 56545 2745
rect 56475 2695 56545 2725
rect 56475 2675 56480 2695
rect 56500 2675 56520 2695
rect 56540 2675 56545 2695
rect 56475 2665 56545 2675
rect 56570 2895 56600 2905
rect 56570 2875 56575 2895
rect 56595 2875 56600 2895
rect 56570 2845 56600 2875
rect 56570 2825 56575 2845
rect 56595 2825 56600 2845
rect 56570 2795 56600 2825
rect 56570 2775 56575 2795
rect 56595 2775 56600 2795
rect 56570 2745 56600 2775
rect 56570 2725 56575 2745
rect 56595 2725 56600 2745
rect 56570 2695 56600 2725
rect 56570 2675 56575 2695
rect 56595 2675 56600 2695
rect 56570 2665 56600 2675
rect 56625 2895 56655 2905
rect 56625 2875 56630 2895
rect 56650 2875 56655 2895
rect 56625 2845 56655 2875
rect 56625 2825 56630 2845
rect 56650 2825 56655 2845
rect 56625 2795 56655 2825
rect 56625 2775 56630 2795
rect 56650 2775 56655 2795
rect 56625 2745 56655 2775
rect 56625 2725 56630 2745
rect 56650 2725 56655 2745
rect 56625 2695 56655 2725
rect 56625 2675 56630 2695
rect 56650 2675 56655 2695
rect 56625 2665 56655 2675
rect 56680 2895 56710 2905
rect 56680 2875 56685 2895
rect 56705 2875 56710 2895
rect 56680 2845 56710 2875
rect 56680 2825 56685 2845
rect 56705 2825 56710 2845
rect 56680 2795 56710 2825
rect 56680 2775 56685 2795
rect 56705 2775 56710 2795
rect 56680 2745 56710 2775
rect 56680 2725 56685 2745
rect 56705 2725 56710 2745
rect 56680 2695 56710 2725
rect 56680 2675 56685 2695
rect 56705 2675 56710 2695
rect 56680 2665 56710 2675
rect 56735 2895 56765 2905
rect 56735 2875 56740 2895
rect 56760 2875 56765 2895
rect 56735 2845 56765 2875
rect 56735 2825 56740 2845
rect 56760 2825 56765 2845
rect 56735 2795 56765 2825
rect 56735 2775 56740 2795
rect 56760 2775 56765 2795
rect 56735 2745 56765 2775
rect 56735 2725 56740 2745
rect 56760 2725 56765 2745
rect 56735 2695 56765 2725
rect 56735 2675 56740 2695
rect 56760 2675 56765 2695
rect 56735 2665 56765 2675
rect 56790 2895 56820 2905
rect 56790 2875 56795 2895
rect 56815 2875 56820 2895
rect 56790 2845 56820 2875
rect 56790 2825 56795 2845
rect 56815 2825 56820 2845
rect 56790 2795 56820 2825
rect 56790 2775 56795 2795
rect 56815 2775 56820 2795
rect 56790 2745 56820 2775
rect 56790 2725 56795 2745
rect 56815 2725 56820 2745
rect 56790 2695 56820 2725
rect 56790 2675 56795 2695
rect 56815 2675 56820 2695
rect 56790 2665 56820 2675
rect 56845 2895 56955 2905
rect 56845 2875 56850 2895
rect 56870 2875 56890 2895
rect 56910 2875 56930 2895
rect 56950 2875 56955 2895
rect 56845 2845 56955 2875
rect 56845 2825 56850 2845
rect 56870 2825 56890 2845
rect 56910 2825 56930 2845
rect 56950 2825 56955 2845
rect 56845 2795 56955 2825
rect 56845 2775 56850 2795
rect 56870 2775 56890 2795
rect 56910 2775 56930 2795
rect 56950 2775 56955 2795
rect 56845 2745 56955 2775
rect 56845 2725 56850 2745
rect 56870 2725 56890 2745
rect 56910 2725 56930 2745
rect 56950 2725 56955 2745
rect 56845 2695 56955 2725
rect 56845 2675 56850 2695
rect 56870 2675 56890 2695
rect 56910 2675 56930 2695
rect 56950 2675 56955 2695
rect 56845 2665 56955 2675
rect 56980 2895 57010 2905
rect 56980 2875 56985 2895
rect 57005 2875 57010 2895
rect 56980 2845 57010 2875
rect 56980 2825 56985 2845
rect 57005 2825 57010 2845
rect 56980 2795 57010 2825
rect 56980 2775 56985 2795
rect 57005 2775 57010 2795
rect 56980 2745 57010 2775
rect 56980 2725 56985 2745
rect 57005 2725 57010 2745
rect 56980 2695 57010 2725
rect 56980 2675 56985 2695
rect 57005 2675 57010 2695
rect 56980 2665 57010 2675
rect 57035 2895 57065 2905
rect 57035 2875 57040 2895
rect 57060 2875 57065 2895
rect 57035 2845 57065 2875
rect 57035 2825 57040 2845
rect 57060 2825 57065 2845
rect 57035 2795 57065 2825
rect 57035 2775 57040 2795
rect 57060 2775 57065 2795
rect 57035 2745 57065 2775
rect 57035 2725 57040 2745
rect 57060 2725 57065 2745
rect 57035 2695 57065 2725
rect 57035 2675 57040 2695
rect 57060 2675 57065 2695
rect 57035 2665 57065 2675
rect 57090 2895 57120 2905
rect 57090 2875 57095 2895
rect 57115 2875 57120 2895
rect 57090 2845 57120 2875
rect 57090 2825 57095 2845
rect 57115 2825 57120 2845
rect 57090 2795 57120 2825
rect 57090 2775 57095 2795
rect 57115 2775 57120 2795
rect 57090 2745 57120 2775
rect 57090 2725 57095 2745
rect 57115 2725 57120 2745
rect 57090 2695 57120 2725
rect 57090 2675 57095 2695
rect 57115 2675 57120 2695
rect 57090 2665 57120 2675
rect 57145 2895 57175 2905
rect 57145 2875 57150 2895
rect 57170 2875 57175 2895
rect 57145 2845 57175 2875
rect 57145 2825 57150 2845
rect 57170 2825 57175 2845
rect 57145 2795 57175 2825
rect 57145 2775 57150 2795
rect 57170 2775 57175 2795
rect 57145 2745 57175 2775
rect 57145 2725 57150 2745
rect 57170 2725 57175 2745
rect 57145 2695 57175 2725
rect 57145 2675 57150 2695
rect 57170 2675 57175 2695
rect 57145 2665 57175 2675
rect 57200 2895 57230 2905
rect 57200 2875 57205 2895
rect 57225 2875 57230 2895
rect 57200 2845 57230 2875
rect 57200 2825 57205 2845
rect 57225 2825 57230 2845
rect 57200 2795 57230 2825
rect 57200 2775 57205 2795
rect 57225 2775 57230 2795
rect 57200 2745 57230 2775
rect 57200 2725 57205 2745
rect 57225 2725 57230 2745
rect 57200 2695 57230 2725
rect 57200 2675 57205 2695
rect 57225 2675 57230 2695
rect 57200 2665 57230 2675
rect 57255 2895 57325 2905
rect 57255 2875 57260 2895
rect 57280 2875 57300 2895
rect 57320 2875 57325 2895
rect 57255 2845 57325 2875
rect 57255 2825 57260 2845
rect 57280 2825 57300 2845
rect 57320 2825 57325 2845
rect 57255 2795 57325 2825
rect 57255 2775 57260 2795
rect 57280 2775 57300 2795
rect 57320 2775 57325 2795
rect 57255 2745 57325 2775
rect 57255 2725 57260 2745
rect 57280 2725 57300 2745
rect 57320 2725 57325 2745
rect 57255 2695 57325 2725
rect 57255 2675 57260 2695
rect 57280 2675 57300 2695
rect 57320 2675 57325 2695
rect 57255 2665 57325 2675
rect 58405 2890 58475 2900
rect 56570 2655 56590 2665
rect 56560 2645 56590 2655
rect 56800 2655 56820 2665
rect 56980 2655 57000 2665
rect 56800 2645 56830 2655
rect 56560 2625 56565 2645
rect 56585 2625 56590 2645
rect 56560 2615 56590 2625
rect 56607 2635 56637 2645
rect 56607 2615 56612 2635
rect 56632 2615 56637 2635
rect 56607 2605 56637 2615
rect 56675 2635 56715 2645
rect 56675 2615 56685 2635
rect 56705 2615 56715 2635
rect 56675 2605 56715 2615
rect 56753 2635 56783 2645
rect 56753 2615 56758 2635
rect 56778 2615 56783 2635
rect 56800 2625 56805 2645
rect 56825 2625 56830 2645
rect 56800 2615 56830 2625
rect 56970 2645 57000 2655
rect 57210 2655 57230 2665
rect 57210 2645 57240 2655
rect 56970 2625 56975 2645
rect 56995 2625 57000 2645
rect 56970 2615 57000 2625
rect 57017 2635 57047 2645
rect 57017 2615 57022 2635
rect 57042 2615 57047 2635
rect 56753 2605 56783 2615
rect 57017 2605 57047 2615
rect 57085 2635 57125 2645
rect 57085 2615 57095 2635
rect 57115 2615 57125 2635
rect 57085 2605 57125 2615
rect 57163 2635 57193 2645
rect 57163 2615 57168 2635
rect 57188 2615 57193 2635
rect 57210 2625 57215 2645
rect 57235 2625 57240 2645
rect 57210 2615 57240 2625
rect 57163 2605 57193 2615
rect 56600 2575 56640 2585
rect 56600 2555 56610 2575
rect 56630 2555 56640 2575
rect 56600 2545 56640 2555
rect 57160 2575 57200 2585
rect 57160 2555 57170 2575
rect 57190 2555 57200 2575
rect 57160 2545 57200 2555
rect 56850 2360 56890 2370
rect 56850 2340 56860 2360
rect 56880 2340 56890 2360
rect 56850 2330 56890 2340
rect 56935 2360 56975 2370
rect 56935 2340 56945 2360
rect 56965 2340 56975 2360
rect 56935 2330 56975 2340
rect 55405 2310 55475 2320
rect 58405 2320 58410 2890
rect 58430 2320 58450 2890
rect 58470 2320 58475 2890
rect 58405 2310 58475 2320
rect 58500 2890 58530 2900
rect 58500 2320 58505 2890
rect 58525 2320 58530 2890
rect 58500 2310 58530 2320
rect 58555 2890 58585 2900
rect 58555 2320 58560 2890
rect 58580 2320 58585 2890
rect 58555 2310 58585 2320
rect 58610 2890 58640 2900
rect 58610 2320 58615 2890
rect 58635 2320 58640 2890
rect 58610 2310 58640 2320
rect 58665 2890 58695 2900
rect 58665 2320 58670 2890
rect 58690 2320 58695 2890
rect 58665 2310 58695 2320
rect 58720 2890 58750 2900
rect 58720 2320 58725 2890
rect 58745 2320 58750 2890
rect 58720 2310 58750 2320
rect 58775 2890 58805 2900
rect 58775 2320 58780 2890
rect 58800 2320 58805 2890
rect 58775 2310 58805 2320
rect 58830 2890 58860 2900
rect 58830 2320 58835 2890
rect 58855 2320 58860 2890
rect 58830 2310 58860 2320
rect 58885 2890 58915 2900
rect 58885 2320 58890 2890
rect 58910 2320 58915 2890
rect 58885 2310 58915 2320
rect 58940 2890 58970 2900
rect 58940 2320 58945 2890
rect 58965 2320 58970 2890
rect 58940 2310 58970 2320
rect 58995 2890 59025 2900
rect 58995 2320 59000 2890
rect 59020 2320 59025 2890
rect 58995 2310 59025 2320
rect 59050 2890 59080 2900
rect 59050 2320 59055 2890
rect 59075 2320 59080 2890
rect 59050 2310 59080 2320
rect 59105 2890 59175 2900
rect 59105 2320 59110 2890
rect 59130 2320 59150 2890
rect 59170 2320 59175 2890
rect 59805 2350 59946 2360
rect 59805 2330 59810 2350
rect 59830 2330 59865 2350
rect 59885 2330 59920 2350
rect 59940 2330 59946 2350
rect 59805 2320 59946 2330
rect 59105 2310 59175 2320
rect 56735 2300 56805 2310
rect 55075 2280 55105 2290
rect 55075 2260 55080 2280
rect 55100 2260 55105 2280
rect 55075 2250 55105 2260
rect 55070 2215 55110 2225
rect 55070 2195 55080 2215
rect 55100 2195 55110 2215
rect 55070 2175 55110 2195
rect 55070 2155 55080 2175
rect 55100 2155 55110 2175
rect 55070 2135 55110 2155
rect 55070 2115 55080 2135
rect 55100 2115 55110 2135
rect 55070 2105 55110 2115
rect 56735 2080 56740 2300
rect 56760 2080 56780 2300
rect 56800 2080 56805 2300
rect 56735 2070 56805 2080
rect 56830 2300 56860 2310
rect 56830 2080 56835 2300
rect 56855 2080 56860 2300
rect 56830 2070 56860 2080
rect 56885 2300 56915 2310
rect 56885 2080 56890 2300
rect 56910 2080 56915 2300
rect 56885 2070 56915 2080
rect 56940 2300 56970 2310
rect 56940 2080 56945 2300
rect 56965 2080 56970 2300
rect 56940 2070 56970 2080
rect 56995 2300 57065 2310
rect 56995 2080 57000 2300
rect 57020 2080 57040 2300
rect 57060 2080 57065 2300
rect 58775 2280 58805 2290
rect 58775 2260 58780 2280
rect 58800 2260 58805 2280
rect 58775 2250 58805 2260
rect 58770 2215 58810 2225
rect 58770 2195 58780 2215
rect 58800 2195 58810 2215
rect 58770 2175 58810 2195
rect 58770 2155 58780 2175
rect 58800 2155 58810 2175
rect 58770 2135 58810 2155
rect 58770 2115 58780 2135
rect 58800 2115 58810 2135
rect 58770 2105 58810 2115
rect 56995 2070 57065 2080
rect 56770 2040 56810 2050
rect 56770 2020 56780 2040
rect 56800 2020 56810 2040
rect 56770 2010 56810 2020
rect 56990 2040 57030 2050
rect 56990 2020 57000 2040
rect 57020 2020 57030 2040
rect 56990 2010 57030 2020
rect 55995 1730 56025 1740
rect 55995 1710 56000 1730
rect 56020 1710 56025 1730
rect 55995 1700 56025 1710
rect 56690 1730 56720 1740
rect 56690 1710 56695 1730
rect 56715 1710 56720 1730
rect 56690 1700 56720 1710
rect 57080 1730 57110 1740
rect 57080 1710 57085 1730
rect 57105 1710 57110 1730
rect 57080 1700 57110 1710
rect 54745 1675 54775 1685
rect 54745 1655 54750 1675
rect 54770 1655 54775 1675
rect 54745 1645 54775 1655
rect 55405 1675 55435 1685
rect 55405 1655 55410 1675
rect 55430 1655 55435 1675
rect 55405 1645 55435 1655
rect 58445 1675 58475 1685
rect 58445 1655 58450 1675
rect 58470 1655 58475 1675
rect 58445 1645 58475 1655
rect 59105 1675 59135 1685
rect 59105 1655 59110 1675
rect 59130 1655 59135 1675
rect 59105 1645 59135 1655
rect 55995 1630 56065 1640
rect 54705 1615 54775 1625
rect 54380 1531 54595 1551
rect 54380 1514 54415 1531
rect 54560 1514 54595 1531
rect 54475 1464 54500 1514
rect 54705 1445 54710 1615
rect 54730 1445 54750 1615
rect 54770 1445 54775 1615
rect 54705 1435 54775 1445
rect 54800 1615 54830 1625
rect 54800 1445 54805 1615
rect 54825 1445 54830 1615
rect 54800 1435 54830 1445
rect 54855 1615 54885 1625
rect 54855 1445 54860 1615
rect 54880 1445 54885 1615
rect 54855 1435 54885 1445
rect 54910 1615 54940 1625
rect 54910 1445 54915 1615
rect 54935 1445 54940 1615
rect 54910 1435 54940 1445
rect 54965 1615 54995 1625
rect 54965 1445 54970 1615
rect 54990 1445 54995 1615
rect 54965 1435 54995 1445
rect 55020 1615 55050 1625
rect 55020 1445 55025 1615
rect 55045 1445 55050 1615
rect 55020 1435 55050 1445
rect 55075 1615 55105 1625
rect 55075 1445 55080 1615
rect 55100 1445 55105 1615
rect 55075 1435 55105 1445
rect 55130 1615 55160 1625
rect 55130 1445 55135 1615
rect 55155 1445 55160 1615
rect 55130 1435 55160 1445
rect 55185 1615 55215 1625
rect 55185 1445 55190 1615
rect 55210 1445 55215 1615
rect 55185 1435 55215 1445
rect 55240 1615 55270 1625
rect 55240 1445 55245 1615
rect 55265 1445 55270 1615
rect 55240 1435 55270 1445
rect 55295 1615 55325 1625
rect 55295 1445 55300 1615
rect 55320 1445 55325 1615
rect 55295 1435 55325 1445
rect 55350 1615 55380 1625
rect 55350 1445 55355 1615
rect 55375 1445 55380 1615
rect 55350 1435 55380 1445
rect 55405 1615 55475 1625
rect 55405 1445 55410 1615
rect 55430 1445 55450 1615
rect 55470 1445 55475 1615
rect 55995 1510 56000 1630
rect 56020 1510 56040 1630
rect 56060 1510 56065 1630
rect 55995 1500 56065 1510
rect 56090 1630 56120 1640
rect 56090 1510 56095 1630
rect 56115 1510 56120 1630
rect 56090 1500 56120 1510
rect 56145 1630 56175 1640
rect 56145 1510 56150 1630
rect 56170 1510 56175 1630
rect 56145 1500 56175 1510
rect 56200 1630 56230 1640
rect 56200 1510 56205 1630
rect 56225 1510 56230 1630
rect 56200 1500 56230 1510
rect 56255 1630 56285 1640
rect 56255 1510 56260 1630
rect 56280 1510 56285 1630
rect 56255 1500 56285 1510
rect 56310 1630 56340 1640
rect 56310 1510 56315 1630
rect 56335 1510 56340 1630
rect 56310 1500 56340 1510
rect 56365 1630 56395 1640
rect 56365 1510 56370 1630
rect 56390 1510 56395 1630
rect 56365 1500 56395 1510
rect 56420 1630 56450 1640
rect 56420 1510 56425 1630
rect 56445 1510 56450 1630
rect 56420 1500 56450 1510
rect 56475 1630 56505 1640
rect 56475 1510 56480 1630
rect 56500 1510 56505 1630
rect 56475 1500 56505 1510
rect 56530 1630 56560 1640
rect 56530 1510 56535 1630
rect 56555 1510 56560 1630
rect 56530 1500 56560 1510
rect 56585 1630 56615 1640
rect 56585 1510 56590 1630
rect 56610 1510 56615 1630
rect 56585 1500 56615 1510
rect 56640 1630 56670 1640
rect 56640 1510 56645 1630
rect 56665 1510 56670 1630
rect 56640 1500 56670 1510
rect 56695 1630 56765 1640
rect 56695 1510 56700 1630
rect 56720 1510 56740 1630
rect 56760 1510 56765 1630
rect 56695 1500 56765 1510
rect 57035 1630 57105 1640
rect 57035 1510 57040 1630
rect 57060 1510 57080 1630
rect 57100 1510 57105 1630
rect 57035 1500 57105 1510
rect 57130 1630 57160 1640
rect 57130 1510 57135 1630
rect 57155 1510 57160 1630
rect 57130 1500 57160 1510
rect 57185 1630 57215 1640
rect 57185 1510 57190 1630
rect 57210 1510 57215 1630
rect 57185 1500 57215 1510
rect 57240 1630 57270 1640
rect 57240 1510 57245 1630
rect 57265 1510 57270 1630
rect 57240 1500 57270 1510
rect 57295 1630 57325 1640
rect 57295 1510 57300 1630
rect 57320 1510 57325 1630
rect 57295 1500 57325 1510
rect 57350 1630 57380 1640
rect 57350 1510 57355 1630
rect 57375 1510 57380 1630
rect 57350 1500 57380 1510
rect 57405 1630 57435 1640
rect 57405 1510 57410 1630
rect 57430 1510 57435 1630
rect 57405 1500 57435 1510
rect 57460 1630 57490 1640
rect 57460 1510 57465 1630
rect 57485 1510 57490 1630
rect 57460 1500 57490 1510
rect 57515 1630 57545 1640
rect 57515 1510 57520 1630
rect 57540 1510 57545 1630
rect 57515 1500 57545 1510
rect 57570 1630 57600 1640
rect 57570 1510 57575 1630
rect 57595 1510 57600 1630
rect 57570 1500 57600 1510
rect 57625 1630 57655 1640
rect 57625 1510 57630 1630
rect 57650 1510 57655 1630
rect 57625 1500 57655 1510
rect 57680 1630 57710 1640
rect 57680 1510 57685 1630
rect 57705 1510 57710 1630
rect 57680 1500 57710 1510
rect 57735 1630 57805 1640
rect 57735 1510 57740 1630
rect 57760 1510 57780 1630
rect 57800 1510 57805 1630
rect 57735 1500 57805 1510
rect 58405 1615 58475 1625
rect 55405 1435 55475 1445
rect 56035 1470 56065 1500
rect 56035 1450 56040 1470
rect 56060 1450 56065 1470
rect 56035 1440 56065 1450
rect 56695 1470 56725 1480
rect 56695 1450 56700 1470
rect 56720 1450 56725 1470
rect 56695 1440 56725 1450
rect 57075 1470 57105 1480
rect 57075 1450 57080 1470
rect 57100 1450 57105 1470
rect 57075 1440 57105 1450
rect 57735 1470 57765 1500
rect 57735 1450 57740 1470
rect 57760 1450 57765 1470
rect 57735 1440 57765 1450
rect 58405 1445 58410 1615
rect 58430 1445 58450 1615
rect 58470 1445 58475 1615
rect 58405 1435 58475 1445
rect 58500 1615 58530 1625
rect 58500 1445 58505 1615
rect 58525 1445 58530 1615
rect 58500 1435 58530 1445
rect 58555 1615 58585 1625
rect 58555 1445 58560 1615
rect 58580 1445 58585 1615
rect 58555 1435 58585 1445
rect 58610 1615 58640 1625
rect 58610 1445 58615 1615
rect 58635 1445 58640 1615
rect 58610 1435 58640 1445
rect 58665 1615 58695 1625
rect 58665 1445 58670 1615
rect 58690 1445 58695 1615
rect 58665 1435 58695 1445
rect 58720 1615 58750 1625
rect 58720 1445 58725 1615
rect 58745 1445 58750 1615
rect 58720 1435 58750 1445
rect 58775 1615 58805 1625
rect 58775 1445 58780 1615
rect 58800 1445 58805 1615
rect 58775 1435 58805 1445
rect 58830 1615 58860 1625
rect 58830 1445 58835 1615
rect 58855 1445 58860 1615
rect 58830 1435 58860 1445
rect 58885 1615 58915 1625
rect 58885 1445 58890 1615
rect 58910 1445 58915 1615
rect 58885 1435 58915 1445
rect 58940 1615 58970 1625
rect 58940 1445 58945 1615
rect 58965 1445 58970 1615
rect 58940 1435 58970 1445
rect 58995 1615 59025 1625
rect 58995 1445 59000 1615
rect 59020 1445 59025 1615
rect 58995 1435 59025 1445
rect 59050 1615 59080 1625
rect 59050 1445 59055 1615
rect 59075 1445 59080 1615
rect 59050 1435 59080 1445
rect 59105 1615 59175 1625
rect 59105 1445 59110 1615
rect 59130 1445 59150 1615
rect 59170 1445 59175 1615
rect 59105 1435 59175 1445
rect 59475 1531 59690 1551
rect 59475 1514 59510 1531
rect 59655 1514 59690 1531
rect 54850 1405 54890 1415
rect 54850 1385 54860 1405
rect 54880 1385 54890 1405
rect 54850 1375 54890 1385
rect 54960 1405 55000 1415
rect 54960 1385 54970 1405
rect 54990 1385 55000 1405
rect 54960 1375 55000 1385
rect 55070 1405 55110 1415
rect 55070 1385 55080 1405
rect 55100 1385 55110 1405
rect 55070 1375 55110 1385
rect 55180 1405 55220 1415
rect 55180 1385 55190 1405
rect 55210 1385 55220 1405
rect 55180 1375 55220 1385
rect 55240 1405 55270 1415
rect 55240 1385 55245 1405
rect 55265 1385 55270 1405
rect 55240 1375 55270 1385
rect 55290 1405 55330 1415
rect 55290 1385 55300 1405
rect 55320 1385 55330 1405
rect 55290 1375 55330 1385
rect 58550 1405 58590 1415
rect 58550 1385 58560 1405
rect 58580 1385 58590 1405
rect 58550 1375 58590 1385
rect 58610 1405 58640 1415
rect 58610 1385 58615 1405
rect 58635 1385 58640 1405
rect 58610 1375 58640 1385
rect 58660 1405 58700 1415
rect 58660 1385 58670 1405
rect 58690 1385 58700 1405
rect 58660 1375 58700 1385
rect 58770 1405 58810 1415
rect 58770 1385 58780 1405
rect 58800 1385 58810 1405
rect 58770 1375 58810 1385
rect 58880 1405 58920 1415
rect 58880 1385 58890 1405
rect 58910 1385 58920 1405
rect 58880 1375 58920 1385
rect 58990 1405 59030 1415
rect 58990 1385 59000 1405
rect 59020 1385 59030 1405
rect 58990 1375 59030 1385
rect 55235 1340 55275 1350
rect 55235 1320 55245 1340
rect 55265 1320 55275 1340
rect 55235 1300 55275 1320
rect 55235 1280 55245 1300
rect 55265 1280 55275 1300
rect 55235 1270 55275 1280
rect 58605 1340 58645 1350
rect 58605 1320 58615 1340
rect 58635 1320 58645 1340
rect 58605 1300 58645 1320
rect 58605 1280 58615 1300
rect 58635 1280 58645 1300
rect 59570 1464 59595 1514
rect 58605 1270 58645 1280
rect 55240 1235 55270 1245
rect 55240 1215 55245 1235
rect 55265 1215 55270 1235
rect 55240 1205 55270 1215
rect 58610 1235 58640 1245
rect 58610 1215 58615 1235
rect 58635 1215 58640 1235
rect 58610 1205 58640 1215
rect 54705 1175 54775 1185
rect 54380 905 54415 915
rect 54380 880 54385 905
rect 54410 880 54415 905
rect 54380 870 54415 880
rect 54440 905 54475 915
rect 54440 880 54445 905
rect 54470 880 54475 905
rect 54440 870 54475 880
rect 54500 905 54535 915
rect 54500 880 54505 905
rect 54530 880 54535 905
rect 54500 870 54535 880
rect 54560 905 54595 915
rect 54560 880 54565 905
rect 54590 880 54595 905
rect 54705 905 54710 1175
rect 54730 905 54750 1175
rect 54770 905 54775 1175
rect 54705 895 54775 905
rect 54800 1175 54830 1185
rect 54800 905 54805 1175
rect 54825 905 54830 1175
rect 54800 895 54830 905
rect 54855 1175 54885 1185
rect 54855 905 54860 1175
rect 54880 905 54885 1175
rect 54855 895 54885 905
rect 54910 1175 54940 1185
rect 54910 905 54915 1175
rect 54935 905 54940 1175
rect 54910 895 54940 905
rect 54965 1175 54995 1185
rect 54965 905 54970 1175
rect 54990 905 54995 1175
rect 54965 895 54995 905
rect 55020 1175 55050 1185
rect 55020 905 55025 1175
rect 55045 905 55050 1175
rect 55020 895 55050 905
rect 55075 1175 55105 1185
rect 55075 905 55080 1175
rect 55100 905 55105 1175
rect 55075 895 55105 905
rect 55130 1175 55160 1185
rect 55130 905 55135 1175
rect 55155 905 55160 1175
rect 55130 895 55160 905
rect 55185 1175 55215 1185
rect 55185 905 55190 1175
rect 55210 905 55215 1175
rect 55185 895 55215 905
rect 55240 1175 55270 1185
rect 55240 905 55245 1175
rect 55265 905 55270 1175
rect 55240 895 55270 905
rect 55295 1175 55325 1185
rect 55295 905 55300 1175
rect 55320 905 55325 1175
rect 55295 895 55325 905
rect 55350 1175 55380 1185
rect 55350 905 55355 1175
rect 55375 905 55380 1175
rect 55350 895 55380 905
rect 55405 1175 55475 1185
rect 55405 905 55410 1175
rect 55430 905 55450 1175
rect 55470 905 55475 1175
rect 58405 1175 58475 1185
rect 56690 1050 56720 1060
rect 56040 1040 56070 1050
rect 56040 1020 56045 1040
rect 56065 1020 56070 1040
rect 56690 1030 56695 1050
rect 56715 1030 56720 1050
rect 56690 1020 56720 1030
rect 56840 1050 56870 1060
rect 56840 1030 56845 1050
rect 56865 1030 56870 1050
rect 56840 1020 56870 1030
rect 56930 1050 56960 1060
rect 56930 1030 56935 1050
rect 56955 1030 56960 1050
rect 56930 1020 56960 1030
rect 57080 1050 57110 1060
rect 57080 1030 57085 1050
rect 57105 1030 57110 1050
rect 57080 1020 57110 1030
rect 57730 1040 57760 1050
rect 57730 1020 57735 1040
rect 57755 1020 57760 1040
rect 56040 1010 56070 1020
rect 57730 1010 57760 1020
rect 55405 895 55475 905
rect 55995 955 56065 965
rect 54560 870 54595 880
rect 54745 865 54775 875
rect 54745 845 54750 865
rect 54770 845 54775 865
rect 54745 830 54775 845
rect 55405 865 55435 875
rect 55405 845 55410 865
rect 55430 845 55435 865
rect 55405 830 55435 845
rect 55995 835 56000 955
rect 56020 835 56040 955
rect 56060 835 56065 955
rect 55995 825 56065 835
rect 56090 955 56120 965
rect 56090 835 56095 955
rect 56115 835 56120 955
rect 56090 825 56120 835
rect 56145 955 56175 965
rect 56145 835 56150 955
rect 56170 835 56175 955
rect 56145 825 56175 835
rect 56200 955 56230 965
rect 56200 835 56205 955
rect 56225 835 56230 955
rect 56200 825 56230 835
rect 56255 955 56285 965
rect 56255 835 56260 955
rect 56280 835 56285 955
rect 56255 825 56285 835
rect 56310 955 56340 965
rect 56310 835 56315 955
rect 56335 835 56340 955
rect 56310 825 56340 835
rect 56365 955 56395 965
rect 56365 835 56370 955
rect 56390 835 56395 955
rect 56365 825 56395 835
rect 56420 955 56450 965
rect 56420 835 56425 955
rect 56445 835 56450 955
rect 56420 825 56450 835
rect 56475 955 56505 965
rect 56475 835 56480 955
rect 56500 835 56505 955
rect 56475 825 56505 835
rect 56530 955 56560 965
rect 56530 835 56535 955
rect 56555 835 56560 955
rect 56530 825 56560 835
rect 56585 955 56615 965
rect 56585 835 56590 955
rect 56610 835 56615 955
rect 56585 825 56615 835
rect 56640 955 56670 965
rect 56640 835 56645 955
rect 56665 835 56670 955
rect 56640 825 56670 835
rect 56695 955 56805 965
rect 56695 835 56700 955
rect 56720 835 56740 955
rect 56760 835 56780 955
rect 56800 835 56805 955
rect 56695 825 56805 835
rect 56830 955 56860 965
rect 56830 835 56835 955
rect 56855 835 56860 955
rect 56830 825 56860 835
rect 56885 955 56915 965
rect 56885 835 56890 955
rect 56910 835 56915 955
rect 56885 825 56915 835
rect 56940 955 56970 965
rect 56940 835 56945 955
rect 56965 835 56970 955
rect 56940 825 56970 835
rect 56995 955 57105 965
rect 56995 835 57000 955
rect 57020 835 57040 955
rect 57060 835 57080 955
rect 57100 835 57105 955
rect 56995 825 57105 835
rect 57130 955 57160 965
rect 57130 835 57135 955
rect 57155 835 57160 955
rect 57130 825 57160 835
rect 57185 955 57215 965
rect 57185 835 57190 955
rect 57210 835 57215 955
rect 57185 825 57215 835
rect 57240 955 57270 965
rect 57240 835 57245 955
rect 57265 835 57270 955
rect 57240 825 57270 835
rect 57295 955 57325 965
rect 57295 835 57300 955
rect 57320 835 57325 955
rect 57295 825 57325 835
rect 57350 955 57380 965
rect 57350 835 57355 955
rect 57375 835 57380 955
rect 57350 825 57380 835
rect 57405 955 57435 965
rect 57405 835 57410 955
rect 57430 835 57435 955
rect 57405 825 57435 835
rect 57460 955 57490 965
rect 57460 835 57465 955
rect 57485 835 57490 955
rect 57460 825 57490 835
rect 57515 955 57545 965
rect 57515 835 57520 955
rect 57540 835 57545 955
rect 57515 825 57545 835
rect 57570 955 57600 965
rect 57570 835 57575 955
rect 57595 835 57600 955
rect 57570 825 57600 835
rect 57625 955 57655 965
rect 57625 835 57630 955
rect 57650 835 57655 955
rect 57625 825 57655 835
rect 57680 955 57710 965
rect 57680 835 57685 955
rect 57705 835 57710 955
rect 57680 825 57710 835
rect 57735 955 57805 965
rect 57735 835 57740 955
rect 57760 835 57780 955
rect 57800 835 57805 955
rect 58405 905 58410 1175
rect 58430 905 58450 1175
rect 58470 905 58475 1175
rect 58405 895 58475 905
rect 58500 1175 58530 1185
rect 58500 905 58505 1175
rect 58525 905 58530 1175
rect 58500 895 58530 905
rect 58555 1175 58585 1185
rect 58555 905 58560 1175
rect 58580 905 58585 1175
rect 58555 895 58585 905
rect 58610 1175 58640 1185
rect 58610 905 58615 1175
rect 58635 905 58640 1175
rect 58610 895 58640 905
rect 58665 1175 58695 1185
rect 58665 905 58670 1175
rect 58690 905 58695 1175
rect 58665 895 58695 905
rect 58720 1175 58750 1185
rect 58720 905 58725 1175
rect 58745 905 58750 1175
rect 58720 895 58750 905
rect 58775 1175 58805 1185
rect 58775 905 58780 1175
rect 58800 905 58805 1175
rect 58775 895 58805 905
rect 58830 1175 58860 1185
rect 58830 905 58835 1175
rect 58855 905 58860 1175
rect 58830 895 58860 905
rect 58885 1175 58915 1185
rect 58885 905 58890 1175
rect 58910 905 58915 1175
rect 58885 895 58915 905
rect 58940 1175 58970 1185
rect 58940 905 58945 1175
rect 58965 905 58970 1175
rect 58940 895 58970 905
rect 58995 1175 59025 1185
rect 58995 905 59000 1175
rect 59020 905 59025 1175
rect 58995 895 59025 905
rect 59050 1175 59080 1185
rect 59050 905 59055 1175
rect 59075 905 59080 1175
rect 59050 895 59080 905
rect 59105 1175 59175 1185
rect 59105 905 59110 1175
rect 59130 905 59150 1175
rect 59170 905 59175 1175
rect 59105 895 59175 905
rect 59475 905 59510 915
rect 59475 880 59480 905
rect 59505 880 59510 905
rect 57735 825 57805 835
rect 58445 865 58475 875
rect 58445 845 58450 865
rect 58470 845 58475 865
rect 58445 830 58475 845
rect 59105 865 59135 875
rect 59475 870 59510 880
rect 59535 905 59570 915
rect 59535 880 59540 905
rect 59565 880 59570 905
rect 59535 870 59570 880
rect 59595 905 59630 915
rect 59595 880 59600 905
rect 59625 880 59630 905
rect 59595 870 59630 880
rect 59655 905 59690 915
rect 59655 880 59660 905
rect 59685 880 59690 905
rect 59655 870 59690 880
rect 59105 845 59110 865
rect 59130 845 59135 865
rect 59105 835 59135 845
rect 56040 805 56065 825
rect 56035 795 56065 805
rect 56035 775 56040 795
rect 56060 775 56065 795
rect 56035 765 56065 775
rect 56735 795 56765 805
rect 56735 775 56740 795
rect 56760 775 56765 795
rect 56735 765 56765 775
rect 57035 795 57065 805
rect 57035 775 57040 795
rect 57060 775 57065 795
rect 57035 765 57065 775
rect 57735 795 57765 825
rect 57735 775 57740 795
rect 57760 775 57765 795
rect 57735 765 57765 775
rect 55100 505 55140 515
rect 55100 485 55110 505
rect 55130 485 55140 505
rect 55100 475 55140 485
rect 58580 505 58620 515
rect 58580 485 58590 505
rect 58610 485 58620 505
rect 58580 475 58620 485
rect 56825 375 56865 385
rect 56825 355 56835 375
rect 56855 355 56865 375
rect 56825 345 56865 355
rect 56935 375 56975 385
rect 56935 355 56945 375
rect 56965 355 56975 375
rect 56935 345 56975 355
rect 56185 315 56255 325
rect 54520 170 54555 180
rect 54520 145 54525 170
rect 54550 145 54555 170
rect 54520 135 54555 145
rect 54580 170 54615 180
rect 54580 145 54585 170
rect 54610 145 54615 170
rect 54580 135 54615 145
rect 54715 165 54785 175
rect 54555 -552 54580 -502
rect 54715 -505 54720 165
rect 54740 -505 54760 165
rect 54780 -505 54785 165
rect 54715 -515 54785 -505
rect 54855 165 54885 175
rect 54855 -505 54860 165
rect 54880 -505 54885 165
rect 54855 -515 54885 -505
rect 54955 165 54985 175
rect 54955 -505 54960 165
rect 54980 -505 54985 165
rect 54955 -515 54985 -505
rect 55055 165 55085 175
rect 55055 -505 55060 165
rect 55080 -505 55085 165
rect 55055 -515 55085 -505
rect 55155 165 55185 175
rect 55155 -505 55160 165
rect 55180 -505 55185 165
rect 55155 -515 55185 -505
rect 55255 165 55285 175
rect 55255 -505 55260 165
rect 55280 -505 55285 165
rect 55255 -515 55285 -505
rect 55355 165 55425 175
rect 55355 -505 55360 165
rect 55380 -505 55400 165
rect 55420 -505 55425 165
rect 56185 95 56190 315
rect 56210 95 56230 315
rect 56250 95 56255 315
rect 56185 85 56255 95
rect 56280 315 56310 325
rect 56280 95 56285 315
rect 56305 95 56310 315
rect 56280 85 56310 95
rect 56335 315 56365 325
rect 56335 95 56340 315
rect 56360 95 56365 315
rect 56335 85 56365 95
rect 56390 315 56420 325
rect 56390 95 56395 315
rect 56415 95 56420 315
rect 56390 85 56420 95
rect 56445 315 56475 325
rect 56445 95 56450 315
rect 56470 95 56475 315
rect 56445 85 56475 95
rect 56500 315 56530 325
rect 56500 95 56505 315
rect 56525 95 56530 315
rect 56500 85 56530 95
rect 56555 315 56585 325
rect 56555 95 56560 315
rect 56580 95 56585 315
rect 56555 85 56585 95
rect 56610 315 56640 325
rect 56610 95 56615 315
rect 56635 95 56640 315
rect 56610 85 56640 95
rect 56665 315 56695 325
rect 56665 95 56670 315
rect 56690 95 56695 315
rect 56665 85 56695 95
rect 56720 315 56750 325
rect 56720 95 56725 315
rect 56745 95 56750 315
rect 56720 85 56750 95
rect 56775 315 56805 325
rect 56775 95 56780 315
rect 56800 95 56805 315
rect 56775 85 56805 95
rect 56830 315 56860 325
rect 56830 95 56835 315
rect 56855 95 56860 315
rect 56830 85 56860 95
rect 56885 315 56915 325
rect 56885 95 56890 315
rect 56910 95 56915 315
rect 56885 85 56915 95
rect 56940 315 56970 325
rect 56940 95 56945 315
rect 56965 95 56970 315
rect 56940 85 56970 95
rect 56995 315 57025 325
rect 56995 95 57000 315
rect 57020 95 57025 315
rect 56995 85 57025 95
rect 57050 315 57080 325
rect 57050 95 57055 315
rect 57075 95 57080 315
rect 57050 85 57080 95
rect 57105 315 57135 325
rect 57105 95 57110 315
rect 57130 95 57135 315
rect 57105 85 57135 95
rect 57160 315 57190 325
rect 57160 95 57165 315
rect 57185 95 57190 315
rect 57160 85 57190 95
rect 57215 315 57245 325
rect 57215 95 57220 315
rect 57240 95 57245 315
rect 57215 85 57245 95
rect 57270 315 57300 325
rect 57270 95 57275 315
rect 57295 95 57300 315
rect 57270 85 57300 95
rect 57325 315 57355 325
rect 57325 95 57330 315
rect 57350 95 57355 315
rect 57325 85 57355 95
rect 57380 315 57410 325
rect 57380 95 57385 315
rect 57405 95 57410 315
rect 57380 85 57410 95
rect 57435 315 57465 325
rect 57435 95 57440 315
rect 57460 95 57465 315
rect 57435 85 57465 95
rect 57490 315 57560 325
rect 57490 95 57495 315
rect 57515 95 57535 315
rect 57555 95 57560 315
rect 57490 85 57560 95
rect 58295 165 58365 175
rect 56220 55 56260 65
rect 56220 35 56230 55
rect 56250 35 56260 55
rect 56220 25 56260 35
rect 57485 55 57525 65
rect 57485 35 57495 55
rect 57515 35 57525 55
rect 57485 25 57525 35
rect 57415 -45 57455 -35
rect 57415 -65 57425 -45
rect 57445 -65 57455 -45
rect 57415 -75 57455 -65
rect 56595 -280 56635 -270
rect 56595 -300 56605 -280
rect 56625 -300 56635 -280
rect 56595 -310 56635 -300
rect 57040 -280 57080 -270
rect 57040 -300 57050 -280
rect 57070 -300 57080 -280
rect 57040 -310 57080 -300
rect 56395 -340 56465 -330
rect 56395 -460 56400 -340
rect 56420 -460 56440 -340
rect 56460 -460 56465 -340
rect 56395 -470 56465 -460
rect 56490 -340 56520 -330
rect 56490 -460 56495 -340
rect 56515 -460 56520 -340
rect 56490 -470 56520 -460
rect 56545 -340 56575 -330
rect 56545 -460 56550 -340
rect 56570 -460 56575 -340
rect 56545 -470 56575 -460
rect 56600 -340 56630 -330
rect 56600 -460 56605 -340
rect 56625 -460 56630 -340
rect 56600 -470 56630 -460
rect 56655 -340 56685 -330
rect 56655 -460 56660 -340
rect 56680 -460 56685 -340
rect 56655 -470 56685 -460
rect 56710 -340 56740 -330
rect 56710 -460 56715 -340
rect 56735 -460 56740 -340
rect 56710 -470 56740 -460
rect 56765 -340 56835 -330
rect 56765 -460 56770 -340
rect 56790 -460 56810 -340
rect 56830 -460 56835 -340
rect 56765 -470 56835 -460
rect 56875 -340 56905 -330
rect 56875 -460 56880 -340
rect 56900 -460 56905 -340
rect 56875 -470 56905 -460
rect 57215 -340 57245 -330
rect 57215 -460 57220 -340
rect 57240 -460 57245 -340
rect 57215 -470 57245 -460
rect 55355 -515 55425 -505
rect 56435 -500 56465 -490
rect 56435 -520 56440 -500
rect 56460 -520 56465 -500
rect 56435 -530 56465 -520
rect 56765 -500 56795 -490
rect 56765 -520 56770 -500
rect 56790 -520 56795 -500
rect 58295 -505 58300 165
rect 58320 -505 58340 165
rect 58360 -505 58365 165
rect 58295 -515 58365 -505
rect 58435 165 58465 175
rect 58435 -505 58440 165
rect 58460 -505 58465 165
rect 58435 -515 58465 -505
rect 58535 165 58565 175
rect 58535 -505 58540 165
rect 58560 -505 58565 165
rect 58535 -515 58565 -505
rect 58635 165 58665 175
rect 58635 -505 58640 165
rect 58660 -505 58665 165
rect 58635 -515 58665 -505
rect 58735 165 58765 175
rect 58735 -505 58740 165
rect 58760 -505 58765 165
rect 58735 -515 58765 -505
rect 58835 165 58865 175
rect 58835 -505 58840 165
rect 58860 -505 58865 165
rect 58835 -515 58865 -505
rect 58935 165 59005 175
rect 58935 -505 58940 165
rect 58960 -505 58980 165
rect 59000 -505 59005 165
rect 59455 170 59490 180
rect 59455 145 59460 170
rect 59485 145 59490 170
rect 59455 135 59490 145
rect 59515 170 59550 180
rect 59515 145 59520 170
rect 59545 145 59550 170
rect 59515 135 59550 145
rect 58935 -515 59005 -505
rect 56765 -530 56795 -520
rect 54755 -545 54785 -535
rect 54755 -565 54760 -545
rect 54780 -565 54785 -545
rect 54755 -575 54785 -565
rect 55355 -545 55385 -535
rect 55355 -565 55360 -545
rect 55380 -565 55385 -545
rect 55355 -575 55385 -565
rect 58335 -545 58365 -535
rect 58335 -565 58340 -545
rect 58360 -565 58365 -545
rect 58335 -575 58365 -565
rect 58935 -545 58965 -535
rect 58935 -565 58940 -545
rect 58960 -565 58965 -545
rect 59490 -552 59515 -502
rect 58935 -575 58965 -565
<< viali >>
rect 56095 4905 56115 4925
rect 56275 4905 56295 4925
rect 57035 4905 57055 4925
rect 57215 4905 57235 4925
rect 57505 4905 57525 4925
rect 57685 4905 57705 4925
rect 56095 4545 56115 4865
rect 56155 4545 56175 4865
rect 56215 4545 56235 4865
rect 56275 4545 56295 4865
rect 56565 4735 56585 4755
rect 56745 4735 56765 4755
rect 56565 4545 56585 4695
rect 56625 4545 56645 4695
rect 56685 4545 56705 4695
rect 56745 4545 56765 4695
rect 57035 4545 57055 4865
rect 57095 4545 57115 4865
rect 57155 4545 57175 4865
rect 57215 4545 57235 4865
rect 57505 4545 57525 4865
rect 57565 4545 57585 4865
rect 57625 4545 57645 4865
rect 57685 4545 57705 4865
rect 56160 4455 56180 4475
rect 56635 4455 56655 4475
rect 57145 4455 57165 4475
rect 57581 4445 57601 4465
rect 54850 3430 54870 3750
rect 54910 3430 54930 3750
rect 54970 3430 54990 3750
rect 55030 3430 55050 3750
rect 55090 3430 55110 3750
rect 55150 3430 55170 3750
rect 55210 3430 55230 3750
rect 55270 3430 55290 3750
rect 55330 3430 55350 3750
rect 55390 3430 55410 3750
rect 55450 3430 55470 3750
rect 55510 3430 55530 3750
rect 55570 3430 55590 3750
rect 56015 3430 56035 3750
rect 56075 3430 56095 3750
rect 56135 3430 56155 3750
rect 56195 3430 56215 3750
rect 56255 3430 56275 3750
rect 56315 3430 56335 3750
rect 56375 3430 56395 3750
rect 56435 3430 56455 3750
rect 56495 3430 56515 3750
rect 56555 3430 56575 3750
rect 56615 3430 56635 3750
rect 56675 3430 56695 3750
rect 56735 3430 56755 3750
rect 57045 3430 57065 3750
rect 57105 3430 57125 3750
rect 57165 3430 57185 3750
rect 57225 3430 57245 3750
rect 57285 3430 57305 3750
rect 57345 3430 57365 3750
rect 57405 3430 57425 3750
rect 57465 3430 57485 3750
rect 57525 3430 57545 3750
rect 57585 3430 57605 3750
rect 57645 3430 57665 3750
rect 57705 3430 57725 3750
rect 57765 3430 57785 3750
rect 58420 3430 58440 3750
rect 58480 3430 58500 3750
rect 58540 3430 58560 3750
rect 58600 3430 58620 3750
rect 58660 3430 58680 3750
rect 58720 3430 58740 3750
rect 58780 3430 58800 3750
rect 58840 3430 58860 3750
rect 58900 3430 58920 3750
rect 58960 3430 58980 3750
rect 59020 3430 59040 3750
rect 59080 3430 59100 3750
rect 59140 3430 59160 3750
rect 54850 3370 54870 3390
rect 55570 3370 55590 3390
rect 56015 3370 56035 3390
rect 56735 3370 56755 3390
rect 57045 3370 57065 3390
rect 57765 3370 57785 3390
rect 58420 3370 58440 3390
rect 59140 3370 59160 3390
rect 56375 3305 56395 3325
rect 57405 3305 57425 3325
rect 55210 3260 55230 3280
rect 58780 3260 58800 3280
rect 54130 3020 54150 3040
rect 54185 3020 54205 3040
rect 54240 3020 54260 3040
rect 56520 2990 56540 3010
rect 56685 2990 56705 3010
rect 56850 2990 56870 3010
rect 56930 2990 56950 3010
rect 57095 2990 57115 3010
rect 57260 2990 57280 3010
rect 54750 2930 54770 2950
rect 55410 2930 55430 2950
rect 56630 2935 56650 2955
rect 56740 2935 56760 2955
rect 57040 2935 57060 2955
rect 57150 2935 57170 2955
rect 58450 2930 58470 2950
rect 59110 2930 59130 2950
rect 59810 2935 59830 2955
rect 59865 2935 59885 2955
rect 59920 2935 59940 2955
rect 54130 2415 54150 2435
rect 54185 2415 54205 2435
rect 54240 2415 54260 2435
rect 54750 2320 54770 2890
rect 54805 2320 54825 2890
rect 54860 2320 54880 2890
rect 54915 2320 54935 2890
rect 54970 2320 54990 2890
rect 55025 2320 55045 2890
rect 55080 2320 55100 2890
rect 55135 2320 55155 2890
rect 55190 2320 55210 2890
rect 55245 2320 55265 2890
rect 55300 2320 55320 2890
rect 55355 2320 55375 2890
rect 55410 2320 55430 2890
rect 56565 2625 56585 2645
rect 56612 2615 56632 2635
rect 56685 2615 56705 2635
rect 56758 2615 56778 2635
rect 56805 2625 56825 2645
rect 56975 2625 56995 2645
rect 57022 2615 57042 2635
rect 57095 2615 57115 2635
rect 57168 2615 57188 2635
rect 57215 2625 57235 2645
rect 56610 2555 56630 2575
rect 57170 2555 57190 2575
rect 56860 2340 56880 2360
rect 56945 2340 56965 2360
rect 58450 2320 58470 2890
rect 58505 2320 58525 2890
rect 58560 2320 58580 2890
rect 58615 2320 58635 2890
rect 58670 2320 58690 2890
rect 58725 2320 58745 2890
rect 58780 2320 58800 2890
rect 58835 2320 58855 2890
rect 58890 2320 58910 2890
rect 58945 2320 58965 2890
rect 59000 2320 59020 2890
rect 59055 2320 59075 2890
rect 59110 2320 59130 2890
rect 59810 2330 59830 2350
rect 59865 2330 59885 2350
rect 59920 2330 59940 2350
rect 55080 2195 55100 2215
rect 55080 2155 55100 2175
rect 55080 2115 55100 2135
rect 56780 2080 56800 2300
rect 56835 2080 56855 2300
rect 56890 2080 56910 2300
rect 56945 2080 56965 2300
rect 57000 2080 57020 2300
rect 58780 2195 58800 2215
rect 58780 2155 58800 2175
rect 58780 2115 58800 2135
rect 56780 2020 56800 2040
rect 57000 2020 57020 2040
rect 56000 1710 56020 1730
rect 56695 1710 56715 1730
rect 57085 1710 57105 1730
rect 54750 1655 54770 1675
rect 55410 1655 55430 1675
rect 58450 1655 58470 1675
rect 59110 1655 59130 1675
rect 54750 1445 54770 1615
rect 54805 1445 54825 1615
rect 54860 1445 54880 1615
rect 54915 1445 54935 1615
rect 54970 1445 54990 1615
rect 55025 1445 55045 1615
rect 55080 1445 55100 1615
rect 55135 1445 55155 1615
rect 55190 1445 55210 1615
rect 55245 1445 55265 1615
rect 55300 1445 55320 1615
rect 55355 1445 55375 1615
rect 55410 1445 55430 1615
rect 56040 1510 56060 1630
rect 56095 1510 56115 1630
rect 56150 1510 56170 1630
rect 56205 1510 56225 1630
rect 56260 1510 56280 1630
rect 56315 1510 56335 1630
rect 56370 1510 56390 1630
rect 56425 1510 56445 1630
rect 56480 1510 56500 1630
rect 56535 1510 56555 1630
rect 56590 1510 56610 1630
rect 56645 1510 56665 1630
rect 56700 1510 56720 1630
rect 57080 1510 57100 1630
rect 57135 1510 57155 1630
rect 57190 1510 57210 1630
rect 57245 1510 57265 1630
rect 57300 1510 57320 1630
rect 57355 1510 57375 1630
rect 57410 1510 57430 1630
rect 57465 1510 57485 1630
rect 57520 1510 57540 1630
rect 57575 1510 57595 1630
rect 57630 1510 57650 1630
rect 57685 1510 57705 1630
rect 57740 1510 57760 1630
rect 56040 1450 56060 1470
rect 56700 1450 56720 1470
rect 57080 1450 57100 1470
rect 57740 1450 57760 1470
rect 58450 1445 58470 1615
rect 58505 1445 58525 1615
rect 58560 1445 58580 1615
rect 58615 1445 58635 1615
rect 58670 1445 58690 1615
rect 58725 1445 58745 1615
rect 58780 1445 58800 1615
rect 58835 1445 58855 1615
rect 58890 1445 58910 1615
rect 58945 1445 58965 1615
rect 59000 1445 59020 1615
rect 59055 1445 59075 1615
rect 59110 1445 59130 1615
rect 54860 1385 54880 1405
rect 54970 1385 54990 1405
rect 55080 1385 55100 1405
rect 55190 1385 55210 1405
rect 55300 1385 55320 1405
rect 58560 1385 58580 1405
rect 58670 1385 58690 1405
rect 58780 1385 58800 1405
rect 58890 1385 58910 1405
rect 59000 1385 59020 1405
rect 55245 1320 55265 1340
rect 55245 1280 55265 1300
rect 58615 1320 58635 1340
rect 58615 1280 58635 1300
rect 54385 880 54410 905
rect 54445 880 54470 905
rect 54505 880 54530 905
rect 54565 880 54590 905
rect 54750 905 54770 1175
rect 54805 905 54825 1175
rect 54860 905 54880 1175
rect 54915 905 54935 1175
rect 54970 905 54990 1175
rect 55025 905 55045 1175
rect 55080 905 55100 1175
rect 55135 905 55155 1175
rect 55190 905 55210 1175
rect 55245 905 55265 1175
rect 55300 905 55320 1175
rect 55355 905 55375 1175
rect 55410 905 55430 1175
rect 56045 1020 56065 1040
rect 56695 1030 56715 1050
rect 56845 1030 56865 1050
rect 56935 1030 56955 1050
rect 57085 1030 57105 1050
rect 57735 1020 57755 1040
rect 54750 845 54770 865
rect 55410 845 55430 865
rect 56040 835 56060 955
rect 56095 835 56115 955
rect 56150 835 56170 955
rect 56205 835 56225 955
rect 56260 835 56280 955
rect 56315 835 56335 955
rect 56370 835 56390 955
rect 56425 835 56445 955
rect 56480 835 56500 955
rect 56535 835 56555 955
rect 56590 835 56610 955
rect 56645 835 56665 955
rect 56700 835 56720 955
rect 56780 835 56800 955
rect 56835 835 56855 955
rect 56890 835 56910 955
rect 56945 835 56965 955
rect 57000 835 57020 955
rect 57080 835 57100 955
rect 57135 835 57155 955
rect 57190 835 57210 955
rect 57245 835 57265 955
rect 57300 835 57320 955
rect 57355 835 57375 955
rect 57410 835 57430 955
rect 57465 835 57485 955
rect 57520 835 57540 955
rect 57575 835 57595 955
rect 57630 835 57650 955
rect 57685 835 57705 955
rect 57740 835 57760 955
rect 58450 905 58470 1175
rect 58505 905 58525 1175
rect 58560 905 58580 1175
rect 58615 905 58635 1175
rect 58670 905 58690 1175
rect 58725 905 58745 1175
rect 58780 905 58800 1175
rect 58835 905 58855 1175
rect 58890 905 58910 1175
rect 58945 905 58965 1175
rect 59000 905 59020 1175
rect 59055 905 59075 1175
rect 59110 905 59130 1175
rect 59480 880 59505 905
rect 58450 845 58470 865
rect 59540 880 59565 905
rect 59600 880 59625 905
rect 59660 880 59685 905
rect 59110 845 59130 865
rect 56040 775 56060 795
rect 56740 775 56760 795
rect 57040 775 57060 795
rect 57740 775 57760 795
rect 55110 485 55130 505
rect 58590 485 58610 505
rect 56835 355 56855 375
rect 56945 355 56965 375
rect 54525 145 54550 170
rect 54585 145 54610 170
rect 54760 -505 54780 165
rect 54860 -505 54880 165
rect 54960 -505 54980 165
rect 55060 -505 55080 165
rect 55160 -505 55180 165
rect 55260 -505 55280 165
rect 55360 -505 55380 165
rect 56230 95 56250 315
rect 56285 95 56305 315
rect 56340 95 56360 315
rect 56395 95 56415 315
rect 56450 95 56470 315
rect 56505 95 56525 315
rect 56560 95 56580 315
rect 56615 95 56635 315
rect 56670 95 56690 315
rect 56725 95 56745 315
rect 56780 95 56800 315
rect 56835 95 56855 315
rect 56890 95 56910 315
rect 56945 95 56965 315
rect 57000 95 57020 315
rect 57055 95 57075 315
rect 57110 95 57130 315
rect 57165 95 57185 315
rect 57220 95 57240 315
rect 57275 95 57295 315
rect 57330 95 57350 315
rect 57385 95 57405 315
rect 57440 95 57460 315
rect 57495 95 57515 315
rect 56230 35 56250 55
rect 57495 35 57515 55
rect 57425 -65 57445 -45
rect 56605 -300 56625 -280
rect 57050 -300 57070 -280
rect 56440 -460 56460 -340
rect 56495 -460 56515 -340
rect 56550 -460 56570 -340
rect 56605 -460 56625 -340
rect 56660 -460 56680 -340
rect 56715 -460 56735 -340
rect 56770 -460 56790 -340
rect 56880 -460 56900 -340
rect 57220 -460 57240 -340
rect 56440 -520 56460 -500
rect 56770 -520 56790 -500
rect 58340 -505 58360 165
rect 58440 -505 58460 165
rect 58540 -505 58560 165
rect 58640 -505 58660 165
rect 58740 -505 58760 165
rect 58840 -505 58860 165
rect 58940 -505 58960 165
rect 59460 145 59485 170
rect 59520 145 59545 170
rect 54760 -565 54780 -545
rect 55360 -565 55380 -545
rect 58340 -565 58360 -545
rect 58940 -565 58960 -545
<< metal1 >>
rect 52290 4320 52410 6460
rect 52290 4290 52295 4320
rect 52325 4290 52335 4320
rect 52365 4290 52375 4320
rect 52405 4290 52410 4320
rect 52290 4280 52410 4290
rect 52290 4250 52295 4280
rect 52325 4250 52335 4280
rect 52365 4250 52375 4280
rect 52405 4250 52410 4280
rect 52290 4240 52410 4250
rect 52290 4210 52295 4240
rect 52325 4210 52335 4240
rect 52365 4210 52375 4240
rect 52405 4210 52410 4240
rect 52290 4205 52410 4210
rect 52640 4320 52760 6460
rect 52640 4290 52645 4320
rect 52675 4290 52685 4320
rect 52715 4290 52725 4320
rect 52755 4290 52760 4320
rect 52640 4280 52760 4290
rect 52640 4250 52645 4280
rect 52675 4250 52685 4280
rect 52715 4250 52725 4280
rect 52755 4250 52760 4280
rect 52640 4240 52760 4250
rect 52640 4210 52645 4240
rect 52675 4210 52685 4240
rect 52715 4210 52725 4240
rect 52755 4210 52760 4240
rect 52640 4205 52760 4210
rect 52990 4320 53110 6460
rect 52990 4290 52995 4320
rect 53025 4290 53035 4320
rect 53065 4290 53075 4320
rect 53105 4290 53110 4320
rect 52990 4280 53110 4290
rect 52990 4250 52995 4280
rect 53025 4250 53035 4280
rect 53065 4250 53075 4280
rect 53105 4250 53110 4280
rect 52990 4240 53110 4250
rect 52990 4210 52995 4240
rect 53025 4210 53035 4240
rect 53065 4210 53075 4240
rect 53105 4210 53110 4240
rect 52990 4205 53110 4210
rect 53690 4090 53810 6460
rect 54040 4325 54160 6460
rect 56205 5065 56245 5070
rect 56205 5035 56210 5065
rect 56240 5035 56245 5065
rect 56085 4930 56125 4935
rect 56085 4900 56090 4930
rect 56120 4900 56125 4930
rect 56085 4895 56125 4900
rect 56205 4930 56245 5035
rect 56675 5065 56715 5070
rect 56675 5035 56680 5065
rect 56710 5035 56715 5065
rect 56675 5030 56715 5035
rect 57085 5065 57125 5070
rect 57085 5035 57090 5065
rect 57120 5035 57125 5065
rect 57085 5030 57125 5035
rect 57555 5065 57595 5070
rect 57555 5035 57560 5065
rect 57590 5035 57595 5065
rect 56205 4900 56210 4930
rect 56240 4900 56245 4930
rect 56205 4895 56245 4900
rect 56265 4930 56305 4935
rect 56265 4900 56270 4930
rect 56300 4900 56305 4930
rect 56265 4895 56305 4900
rect 56090 4865 56120 4895
rect 56090 4545 56095 4865
rect 56115 4545 56120 4865
rect 56090 4535 56120 4545
rect 56150 4865 56180 4875
rect 56150 4545 56155 4865
rect 56175 4545 56180 4865
rect 56150 4485 56180 4545
rect 56210 4865 56240 4895
rect 56210 4545 56215 4865
rect 56235 4545 56240 4865
rect 56210 4530 56240 4545
rect 56270 4865 56300 4895
rect 56270 4545 56275 4865
rect 56295 4545 56300 4865
rect 56555 4840 56595 4845
rect 56555 4810 56560 4840
rect 56590 4810 56595 4840
rect 56555 4800 56595 4810
rect 56555 4770 56560 4800
rect 56590 4770 56595 4800
rect 56555 4760 56595 4770
rect 56555 4730 56560 4760
rect 56590 4730 56595 4760
rect 56555 4725 56595 4730
rect 56615 4840 56655 4845
rect 56615 4810 56620 4840
rect 56650 4810 56655 4840
rect 56615 4800 56655 4810
rect 56615 4770 56620 4800
rect 56650 4770 56655 4800
rect 56615 4760 56655 4770
rect 56615 4730 56620 4760
rect 56650 4730 56655 4760
rect 56615 4725 56655 4730
rect 56270 4535 56300 4545
rect 56560 4695 56590 4725
rect 56560 4545 56565 4695
rect 56585 4545 56590 4695
rect 56560 4535 56590 4545
rect 56620 4695 56650 4725
rect 56620 4545 56625 4695
rect 56645 4545 56650 4695
rect 56620 4535 56650 4545
rect 56680 4695 56710 5030
rect 56880 5010 56920 5015
rect 56880 4980 56885 5010
rect 56915 4980 56920 5010
rect 56880 4970 56920 4980
rect 56880 4940 56885 4970
rect 56915 4940 56920 4970
rect 56880 4930 56920 4940
rect 56880 4900 56885 4930
rect 56915 4900 56920 4930
rect 56735 4840 56775 4845
rect 56735 4810 56740 4840
rect 56770 4810 56775 4840
rect 56735 4800 56775 4810
rect 56735 4770 56740 4800
rect 56770 4770 56775 4800
rect 56735 4760 56775 4770
rect 56735 4730 56740 4760
rect 56770 4730 56775 4760
rect 56735 4725 56775 4730
rect 56880 4840 56920 4900
rect 57025 5010 57065 5015
rect 57025 4980 57030 5010
rect 57060 4980 57065 5010
rect 57025 4970 57065 4980
rect 57025 4940 57030 4970
rect 57060 4940 57065 4970
rect 57025 4930 57065 4940
rect 57025 4900 57030 4930
rect 57060 4900 57065 4930
rect 57025 4895 57065 4900
rect 56880 4810 56885 4840
rect 56915 4810 56920 4840
rect 56880 4800 56920 4810
rect 56880 4770 56885 4800
rect 56915 4770 56920 4800
rect 56880 4760 56920 4770
rect 56880 4730 56885 4760
rect 56915 4730 56920 4760
rect 56680 4545 56685 4695
rect 56705 4545 56710 4695
rect 56680 4530 56710 4545
rect 56740 4695 56770 4725
rect 56740 4545 56745 4695
rect 56765 4545 56770 4695
rect 56740 4535 56770 4545
rect 56205 4525 56245 4530
rect 56205 4495 56210 4525
rect 56240 4495 56245 4525
rect 56205 4490 56245 4495
rect 56675 4525 56715 4530
rect 56675 4495 56680 4525
rect 56710 4495 56715 4525
rect 56675 4490 56715 4495
rect 56150 4480 56190 4485
rect 56150 4450 56155 4480
rect 56185 4450 56190 4480
rect 56150 4445 56190 4450
rect 56630 4480 56660 4485
rect 56630 4445 56660 4450
rect 56825 4480 56865 4485
rect 56825 4450 56830 4480
rect 56860 4450 56865 4480
rect 56825 4445 56865 4450
rect 53960 4320 54160 4325
rect 53960 4290 53965 4320
rect 53995 4290 54005 4320
rect 54035 4290 54045 4320
rect 54075 4290 54160 4320
rect 53960 4280 54160 4290
rect 53960 4250 53965 4280
rect 53995 4250 54005 4280
rect 54035 4250 54045 4280
rect 54075 4250 54160 4280
rect 53960 4240 54160 4250
rect 53960 4210 53965 4240
rect 53995 4210 54005 4240
rect 54035 4210 54045 4240
rect 54075 4210 54160 4240
rect 53960 4205 54160 4210
rect 54310 4320 54430 4325
rect 54310 4290 54315 4320
rect 54345 4290 54355 4320
rect 54385 4290 54395 4320
rect 54425 4290 54430 4320
rect 54310 4280 54430 4290
rect 54310 4250 54315 4280
rect 54345 4250 54355 4280
rect 54385 4250 54395 4280
rect 54425 4250 54430 4280
rect 54310 4240 54430 4250
rect 54310 4210 54315 4240
rect 54345 4210 54355 4240
rect 54385 4210 54395 4240
rect 54425 4210 54430 4240
rect 54310 4205 54430 4210
rect 54840 4320 54880 4325
rect 54840 4290 54845 4320
rect 54875 4290 54880 4320
rect 54840 4280 54880 4290
rect 54840 4250 54845 4280
rect 54875 4250 54880 4280
rect 54840 4240 54880 4250
rect 54840 4210 54845 4240
rect 54875 4210 54880 4240
rect 54080 4090 54160 4205
rect 54840 3800 54880 4210
rect 55200 4320 55240 4325
rect 55200 4290 55205 4320
rect 55235 4290 55240 4320
rect 55200 4280 55240 4290
rect 55200 4250 55205 4280
rect 55235 4250 55240 4280
rect 55200 4240 55240 4250
rect 55200 4210 55205 4240
rect 55235 4210 55240 4240
rect 54900 3935 55180 3940
rect 54900 3905 54905 3935
rect 54935 3905 54945 3935
rect 54975 3905 54985 3935
rect 55015 3905 55025 3935
rect 55055 3905 55065 3935
rect 55095 3905 55105 3935
rect 55135 3905 55145 3935
rect 55175 3905 55180 3935
rect 54900 3895 55180 3905
rect 54900 3865 54905 3895
rect 54935 3865 54945 3895
rect 54975 3865 54985 3895
rect 55015 3865 55025 3895
rect 55055 3865 55065 3895
rect 55095 3865 55105 3895
rect 55135 3865 55145 3895
rect 55175 3865 55180 3895
rect 54900 3855 55180 3865
rect 54900 3825 54905 3855
rect 54935 3825 54945 3855
rect 54975 3825 54985 3855
rect 55015 3825 55025 3855
rect 55055 3825 55065 3855
rect 55095 3825 55105 3855
rect 55135 3825 55145 3855
rect 55175 3825 55180 3855
rect 54900 3820 55180 3825
rect 54840 3770 54845 3800
rect 54875 3770 54880 3800
rect 54840 3765 54880 3770
rect 54845 3750 54875 3765
rect 54845 3430 54850 3750
rect 54870 3430 54875 3750
rect 54845 3390 54875 3430
rect 54905 3750 54935 3820
rect 54960 3800 55000 3805
rect 54960 3770 54965 3800
rect 54995 3770 55000 3800
rect 54960 3765 55000 3770
rect 54905 3430 54910 3750
rect 54930 3430 54935 3750
rect 54905 3415 54935 3430
rect 54965 3750 54995 3765
rect 54965 3430 54970 3750
rect 54990 3430 54995 3750
rect 54965 3420 54995 3430
rect 55025 3750 55055 3820
rect 55080 3800 55120 3805
rect 55080 3770 55085 3800
rect 55115 3770 55120 3800
rect 55080 3765 55120 3770
rect 55025 3430 55030 3750
rect 55050 3430 55055 3750
rect 55025 3415 55055 3430
rect 55085 3750 55115 3765
rect 55085 3430 55090 3750
rect 55110 3430 55115 3750
rect 55085 3420 55115 3430
rect 55145 3750 55175 3820
rect 55200 3800 55240 4210
rect 55560 4320 55600 4325
rect 55560 4290 55565 4320
rect 55595 4290 55600 4320
rect 55560 4280 55600 4290
rect 55560 4250 55565 4280
rect 55595 4250 55600 4280
rect 55560 4240 55600 4250
rect 55560 4210 55565 4240
rect 55595 4210 55600 4240
rect 55260 3935 55540 3940
rect 55260 3905 55265 3935
rect 55295 3905 55305 3935
rect 55335 3905 55345 3935
rect 55375 3905 55385 3935
rect 55415 3905 55425 3935
rect 55455 3905 55465 3935
rect 55495 3905 55505 3935
rect 55535 3905 55540 3935
rect 55260 3895 55540 3905
rect 55260 3865 55265 3895
rect 55295 3865 55305 3895
rect 55335 3865 55345 3895
rect 55375 3865 55385 3895
rect 55415 3865 55425 3895
rect 55455 3865 55465 3895
rect 55495 3865 55505 3895
rect 55535 3865 55540 3895
rect 55260 3855 55540 3865
rect 55260 3825 55265 3855
rect 55295 3825 55305 3855
rect 55335 3825 55345 3855
rect 55375 3825 55385 3855
rect 55415 3825 55425 3855
rect 55455 3825 55465 3855
rect 55495 3825 55505 3855
rect 55535 3825 55540 3855
rect 55260 3820 55540 3825
rect 55200 3770 55205 3800
rect 55235 3770 55240 3800
rect 55200 3765 55240 3770
rect 55145 3430 55150 3750
rect 55170 3430 55175 3750
rect 55145 3415 55175 3430
rect 55205 3750 55235 3765
rect 55205 3430 55210 3750
rect 55230 3430 55235 3750
rect 55205 3420 55235 3430
rect 55265 3750 55295 3820
rect 55320 3800 55360 3805
rect 55320 3770 55325 3800
rect 55355 3770 55360 3800
rect 55320 3765 55360 3770
rect 55265 3430 55270 3750
rect 55290 3430 55295 3750
rect 55265 3415 55295 3430
rect 55325 3750 55355 3765
rect 55325 3430 55330 3750
rect 55350 3430 55355 3750
rect 55325 3420 55355 3430
rect 55385 3750 55415 3820
rect 55440 3800 55480 3805
rect 55440 3770 55445 3800
rect 55475 3770 55480 3800
rect 55440 3765 55480 3770
rect 55385 3430 55390 3750
rect 55410 3430 55415 3750
rect 55385 3415 55415 3430
rect 55445 3750 55475 3765
rect 55445 3430 55450 3750
rect 55470 3430 55475 3750
rect 55445 3420 55475 3430
rect 55505 3750 55535 3820
rect 55560 3800 55600 4210
rect 55560 3770 55565 3800
rect 55595 3770 55600 3800
rect 55560 3765 55600 3770
rect 55660 4320 55780 4325
rect 55660 4290 55665 4320
rect 55695 4290 55705 4320
rect 55735 4290 55745 4320
rect 55775 4290 55780 4320
rect 55660 4280 55780 4290
rect 55660 4250 55665 4280
rect 55695 4250 55705 4280
rect 55735 4250 55745 4280
rect 55775 4250 55780 4280
rect 55660 4240 55780 4250
rect 55660 4210 55665 4240
rect 55695 4210 55705 4240
rect 55735 4210 55745 4240
rect 55775 4210 55780 4240
rect 55505 3430 55510 3750
rect 55530 3430 55535 3750
rect 55505 3415 55535 3430
rect 55565 3750 55595 3765
rect 55565 3430 55570 3750
rect 55590 3430 55595 3750
rect 54845 3370 54850 3390
rect 54870 3370 54875 3390
rect 54900 3410 54940 3415
rect 54900 3380 54905 3410
rect 54935 3380 54940 3410
rect 54900 3375 54940 3380
rect 55020 3410 55060 3415
rect 55020 3380 55025 3410
rect 55055 3380 55060 3410
rect 55020 3375 55060 3380
rect 55140 3410 55180 3415
rect 55140 3380 55145 3410
rect 55175 3380 55180 3410
rect 55140 3375 55180 3380
rect 55260 3410 55300 3415
rect 55260 3380 55265 3410
rect 55295 3380 55300 3410
rect 55260 3375 55300 3380
rect 55380 3410 55420 3415
rect 55380 3380 55385 3410
rect 55415 3380 55420 3410
rect 55380 3375 55420 3380
rect 55500 3410 55540 3415
rect 55500 3380 55505 3410
rect 55535 3380 55540 3410
rect 55500 3375 55540 3380
rect 55565 3390 55595 3430
rect 54845 3360 54875 3370
rect 55565 3370 55570 3390
rect 55590 3370 55595 3390
rect 55565 3360 55595 3370
rect 55200 3285 55240 3290
rect 55200 3255 55205 3285
rect 55235 3255 55240 3285
rect 55200 3250 55240 3255
rect 55520 3240 55640 3245
rect 55520 3210 55525 3240
rect 55555 3210 55565 3240
rect 55595 3210 55605 3240
rect 55635 3210 55640 3240
rect 55520 3200 55640 3210
rect 55520 3170 55525 3200
rect 55555 3170 55565 3200
rect 55595 3170 55605 3200
rect 55635 3170 55640 3200
rect 55520 3160 55640 3170
rect 55520 3130 55525 3160
rect 55555 3130 55565 3160
rect 55595 3130 55605 3160
rect 55635 3130 55640 3160
rect 54175 3125 54215 3130
rect 54175 3095 54180 3125
rect 54210 3095 54215 3125
rect 54175 3090 54215 3095
rect 54740 3105 54780 3110
rect 54185 3050 54205 3090
rect 54740 3075 54745 3105
rect 54775 3075 54780 3105
rect 54740 3065 54780 3075
rect 54124 3040 54265 3050
rect 54124 3020 54130 3040
rect 54150 3020 54185 3040
rect 54205 3020 54240 3040
rect 54260 3020 54265 3040
rect 54124 3010 54265 3020
rect 54740 3035 54745 3065
rect 54775 3035 54780 3065
rect 54740 3025 54780 3035
rect 54740 2995 54745 3025
rect 54775 2995 54780 3025
rect 54740 2990 54780 2995
rect 54850 3105 54890 3110
rect 54850 3075 54855 3105
rect 54885 3075 54890 3105
rect 54850 3065 54890 3075
rect 54850 3035 54855 3065
rect 54885 3035 54890 3065
rect 54850 3025 54890 3035
rect 54850 2995 54855 3025
rect 54885 2995 54890 3025
rect 54850 2990 54890 2995
rect 54960 3105 55000 3110
rect 54960 3075 54965 3105
rect 54995 3075 55000 3105
rect 54960 3065 55000 3075
rect 54960 3035 54965 3065
rect 54995 3035 55000 3065
rect 54960 3025 55000 3035
rect 54960 2995 54965 3025
rect 54995 2995 55000 3025
rect 54960 2990 55000 2995
rect 55070 3105 55110 3110
rect 55070 3075 55075 3105
rect 55105 3075 55110 3105
rect 55070 3065 55110 3075
rect 55070 3035 55075 3065
rect 55105 3035 55110 3065
rect 55070 3025 55110 3035
rect 55070 2995 55075 3025
rect 55105 2995 55110 3025
rect 55070 2990 55110 2995
rect 55180 3105 55220 3110
rect 55180 3075 55185 3105
rect 55215 3075 55220 3105
rect 55180 3065 55220 3075
rect 55180 3035 55185 3065
rect 55215 3035 55220 3065
rect 55180 3025 55220 3035
rect 55180 2995 55185 3025
rect 55215 2995 55220 3025
rect 55180 2990 55220 2995
rect 55290 3105 55330 3110
rect 55290 3075 55295 3105
rect 55325 3075 55330 3105
rect 55290 3065 55330 3075
rect 55290 3035 55295 3065
rect 55325 3035 55330 3065
rect 55290 3025 55330 3035
rect 55290 2995 55295 3025
rect 55325 2995 55330 3025
rect 55290 2990 55330 2995
rect 55400 3105 55440 3110
rect 55400 3075 55405 3105
rect 55435 3075 55440 3105
rect 55400 3065 55440 3075
rect 55400 3035 55405 3065
rect 55435 3035 55440 3065
rect 55400 3025 55440 3035
rect 55400 2995 55405 3025
rect 55435 2995 55440 3025
rect 55400 2990 55440 2995
rect 54745 2950 54775 2990
rect 54745 2930 54750 2950
rect 54770 2930 54775 2950
rect 54745 2890 54775 2930
rect 54795 2940 54835 2945
rect 54795 2910 54800 2940
rect 54830 2910 54835 2940
rect 54795 2905 54835 2910
rect 54124 2435 54265 2445
rect 54124 2415 54130 2435
rect 54150 2415 54185 2435
rect 54205 2415 54240 2435
rect 54260 2415 54265 2435
rect 54124 2405 54265 2415
rect 54135 2220 54255 2405
rect 54745 2320 54750 2890
rect 54770 2320 54775 2890
rect 54745 2310 54775 2320
rect 54800 2890 54830 2905
rect 54800 2320 54805 2890
rect 54825 2320 54830 2890
rect 54800 2305 54830 2320
rect 54855 2890 54885 2990
rect 54905 2940 54945 2945
rect 54905 2910 54910 2940
rect 54940 2910 54945 2940
rect 54905 2905 54945 2910
rect 54855 2320 54860 2890
rect 54880 2320 54885 2890
rect 54855 2310 54885 2320
rect 54910 2890 54940 2905
rect 54910 2320 54915 2890
rect 54935 2320 54940 2890
rect 54910 2305 54940 2320
rect 54965 2890 54995 2990
rect 55015 2940 55055 2945
rect 55015 2910 55020 2940
rect 55050 2910 55055 2940
rect 55015 2905 55055 2910
rect 54965 2320 54970 2890
rect 54990 2320 54995 2890
rect 54965 2310 54995 2320
rect 55020 2890 55050 2905
rect 55020 2320 55025 2890
rect 55045 2320 55050 2890
rect 55020 2305 55050 2320
rect 55075 2890 55105 2990
rect 55125 2940 55165 2945
rect 55125 2910 55130 2940
rect 55160 2910 55165 2940
rect 55125 2905 55165 2910
rect 55075 2320 55080 2890
rect 55100 2320 55105 2890
rect 55075 2310 55105 2320
rect 55130 2890 55160 2905
rect 55130 2320 55135 2890
rect 55155 2320 55160 2890
rect 55130 2305 55160 2320
rect 55185 2890 55215 2990
rect 55235 2940 55275 2945
rect 55235 2910 55240 2940
rect 55270 2910 55275 2940
rect 55235 2905 55275 2910
rect 55185 2320 55190 2890
rect 55210 2320 55215 2890
rect 55185 2310 55215 2320
rect 55240 2890 55270 2905
rect 55240 2320 55245 2890
rect 55265 2320 55270 2890
rect 55240 2305 55270 2320
rect 55295 2890 55325 2990
rect 55405 2950 55435 2990
rect 55345 2940 55385 2945
rect 55345 2910 55350 2940
rect 55380 2910 55385 2940
rect 55345 2905 55385 2910
rect 55405 2930 55410 2950
rect 55430 2930 55435 2950
rect 55295 2320 55300 2890
rect 55320 2320 55325 2890
rect 55295 2310 55325 2320
rect 55350 2890 55380 2905
rect 55350 2320 55355 2890
rect 55375 2320 55380 2890
rect 55350 2305 55380 2320
rect 55405 2890 55435 2930
rect 55405 2320 55410 2890
rect 55430 2320 55435 2890
rect 55405 2310 55435 2320
rect 54135 2190 54140 2220
rect 54170 2190 54180 2220
rect 54210 2190 54220 2220
rect 54250 2190 54255 2220
rect 54135 2180 54255 2190
rect 54135 2150 54140 2180
rect 54170 2150 54180 2180
rect 54210 2150 54220 2180
rect 54250 2150 54255 2180
rect 54135 2140 54255 2150
rect 54135 2110 54140 2140
rect 54170 2110 54180 2140
rect 54210 2110 54220 2140
rect 54250 2110 54255 2140
rect 54135 2105 54255 2110
rect 54795 2300 54835 2305
rect 54795 2270 54800 2300
rect 54830 2270 54835 2300
rect 54795 2075 54835 2270
rect 54905 2300 54945 2305
rect 54905 2270 54910 2300
rect 54940 2270 54945 2300
rect 54905 2075 54945 2270
rect 55015 2300 55055 2305
rect 55015 2270 55020 2300
rect 55050 2270 55055 2300
rect 55015 2075 55055 2270
rect 55125 2300 55165 2305
rect 55125 2270 55130 2300
rect 55160 2270 55165 2300
rect 55070 2220 55110 2225
rect 55070 2190 55075 2220
rect 55105 2190 55110 2220
rect 55070 2180 55110 2190
rect 55070 2150 55075 2180
rect 55105 2150 55110 2180
rect 55070 2140 55110 2150
rect 55070 2110 55075 2140
rect 55105 2110 55110 2140
rect 55070 2105 55110 2110
rect 55125 2075 55165 2270
rect 55235 2300 55275 2305
rect 55235 2270 55240 2300
rect 55270 2270 55275 2300
rect 55235 2075 55275 2270
rect 55345 2300 55385 2305
rect 55345 2270 55350 2300
rect 55380 2270 55385 2300
rect 55345 2075 55385 2270
rect 54105 2070 54355 2075
rect 54105 2040 54110 2070
rect 54140 2040 54150 2070
rect 54180 2040 54195 2070
rect 54225 2040 54235 2070
rect 54265 2040 54280 2070
rect 54310 2040 54320 2070
rect 54350 2040 54355 2070
rect 54105 2030 54355 2040
rect 54105 2000 54110 2030
rect 54140 2000 54150 2030
rect 54180 2000 54195 2030
rect 54225 2000 54235 2030
rect 54265 2000 54280 2030
rect 54310 2000 54320 2030
rect 54350 2000 54355 2030
rect 54105 1990 54355 2000
rect 54105 1960 54110 1990
rect 54140 1960 54150 1990
rect 54180 1960 54195 1990
rect 54225 1960 54235 1990
rect 54265 1960 54280 1990
rect 54310 1960 54320 1990
rect 54350 1960 54355 1990
rect 53960 1800 54080 1805
rect 53960 1770 53965 1800
rect 53995 1770 54005 1800
rect 54035 1770 54045 1800
rect 54075 1770 54080 1800
rect 53960 1760 54080 1770
rect 53960 1730 53965 1760
rect 53995 1730 54005 1760
rect 54035 1730 54045 1760
rect 54075 1730 54080 1760
rect 53960 1720 54080 1730
rect 53960 1690 53965 1720
rect 53995 1690 54005 1720
rect 54035 1690 54045 1720
rect 54075 1690 54080 1720
rect 53960 690 54080 1690
rect 53960 660 53965 690
rect 53995 660 54005 690
rect 54035 660 54045 690
rect 54075 660 54080 690
rect 53960 650 54080 660
rect 53960 620 53965 650
rect 53995 620 54005 650
rect 54035 620 54045 650
rect 54075 620 54080 650
rect 53960 610 54080 620
rect 53960 580 53965 610
rect 53995 580 54005 610
rect 54035 580 54045 610
rect 54075 580 54080 610
rect 52290 -580 52410 -575
rect 52290 -610 52295 -580
rect 52325 -610 52335 -580
rect 52365 -610 52375 -580
rect 52405 -610 52410 -580
rect 52290 -620 52410 -610
rect 52290 -650 52295 -620
rect 52325 -650 52335 -620
rect 52365 -650 52375 -620
rect 52405 -650 52410 -620
rect 52290 -660 52410 -650
rect 52290 -690 52295 -660
rect 52325 -690 52335 -660
rect 52365 -690 52375 -660
rect 52405 -690 52410 -660
rect 52290 -1500 52410 -690
rect 52640 -580 52760 -575
rect 52640 -610 52645 -580
rect 52675 -610 52685 -580
rect 52715 -610 52725 -580
rect 52755 -610 52760 -580
rect 52640 -620 52760 -610
rect 52640 -650 52645 -620
rect 52675 -650 52685 -620
rect 52715 -650 52725 -620
rect 52755 -650 52760 -620
rect 52640 -660 52760 -650
rect 52640 -690 52645 -660
rect 52675 -690 52685 -660
rect 52715 -690 52725 -660
rect 52755 -690 52760 -660
rect 52640 -1500 52760 -690
rect 52990 -580 53110 -575
rect 52990 -610 52995 -580
rect 53025 -610 53035 -580
rect 53065 -610 53075 -580
rect 53105 -610 53110 -580
rect 52990 -620 53110 -610
rect 52990 -650 52995 -620
rect 53025 -650 53035 -620
rect 53065 -650 53075 -620
rect 53105 -650 53110 -620
rect 52990 -660 53110 -650
rect 52990 -690 52995 -660
rect 53025 -690 53035 -660
rect 53065 -690 53075 -660
rect 53105 -690 53110 -660
rect 52990 -1500 53110 -690
rect 53340 -580 53460 -575
rect 53340 -610 53345 -580
rect 53375 -610 53385 -580
rect 53415 -610 53425 -580
rect 53455 -610 53460 -580
rect 53340 -620 53460 -610
rect 53340 -650 53345 -620
rect 53375 -650 53385 -620
rect 53415 -650 53425 -620
rect 53455 -650 53460 -620
rect 53340 -660 53460 -650
rect 53340 -690 53345 -660
rect 53375 -690 53385 -660
rect 53415 -690 53425 -660
rect 53455 -690 53460 -660
rect 53340 -1500 53460 -690
rect 53960 -580 54080 580
rect 54105 1360 54355 1960
rect 54795 2070 55385 2075
rect 54795 2040 54800 2070
rect 54830 2040 54855 2070
rect 54885 2040 54910 2070
rect 54940 2040 54965 2070
rect 54995 2040 55020 2070
rect 55050 2040 55075 2070
rect 55105 2040 55130 2070
rect 55160 2040 55185 2070
rect 55215 2040 55240 2070
rect 55270 2040 55295 2070
rect 55325 2040 55350 2070
rect 55380 2040 55385 2070
rect 54795 2030 55385 2040
rect 54795 2000 54800 2030
rect 54830 2000 54855 2030
rect 54885 2000 54910 2030
rect 54940 2000 54965 2030
rect 54995 2000 55020 2030
rect 55050 2000 55075 2030
rect 55105 2000 55130 2030
rect 55160 2000 55185 2030
rect 55215 2000 55240 2030
rect 55270 2000 55295 2030
rect 55325 2000 55350 2030
rect 55380 2000 55385 2030
rect 54795 1990 55385 2000
rect 54795 1960 54800 1990
rect 54830 1960 54855 1990
rect 54885 1960 54910 1990
rect 54940 1960 54965 1990
rect 54995 1960 55020 1990
rect 55050 1960 55075 1990
rect 55105 1960 55130 1990
rect 55160 1960 55185 1990
rect 55215 1960 55240 1990
rect 55270 1960 55295 1990
rect 55325 1960 55350 1990
rect 55380 1960 55385 1990
rect 54795 1955 55385 1960
rect 55520 2220 55640 3130
rect 55520 2190 55525 2220
rect 55555 2190 55565 2220
rect 55595 2190 55605 2220
rect 55635 2190 55640 2220
rect 55520 2180 55640 2190
rect 55520 2150 55525 2180
rect 55555 2150 55565 2180
rect 55595 2150 55605 2180
rect 55635 2150 55640 2180
rect 55520 2140 55640 2150
rect 55520 2110 55525 2140
rect 55555 2110 55565 2140
rect 55595 2110 55605 2140
rect 55635 2110 55640 2140
rect 54740 1935 54780 1940
rect 54740 1905 54745 1935
rect 54775 1905 54780 1935
rect 54740 1895 54780 1905
rect 54740 1865 54745 1895
rect 54775 1865 54780 1895
rect 54740 1855 54780 1865
rect 54740 1825 54745 1855
rect 54775 1825 54780 1855
rect 54740 1820 54780 1825
rect 55400 1935 55440 1940
rect 55400 1905 55405 1935
rect 55435 1905 55440 1935
rect 55400 1895 55440 1905
rect 55400 1865 55405 1895
rect 55435 1865 55440 1895
rect 55400 1855 55440 1865
rect 55400 1825 55405 1855
rect 55435 1825 55440 1855
rect 55400 1820 55440 1825
rect 54745 1675 54775 1820
rect 54795 1800 54835 1805
rect 54795 1770 54800 1800
rect 54830 1770 54835 1800
rect 54795 1760 54835 1770
rect 54795 1730 54800 1760
rect 54830 1730 54835 1760
rect 54795 1720 54835 1730
rect 54795 1690 54800 1720
rect 54830 1690 54835 1720
rect 54795 1685 54835 1690
rect 54905 1800 54945 1805
rect 54905 1770 54910 1800
rect 54940 1770 54945 1800
rect 54905 1760 54945 1770
rect 54905 1730 54910 1760
rect 54940 1730 54945 1760
rect 54905 1720 54945 1730
rect 54905 1690 54910 1720
rect 54940 1690 54945 1720
rect 54905 1685 54945 1690
rect 55015 1800 55055 1805
rect 55015 1770 55020 1800
rect 55050 1770 55055 1800
rect 55015 1760 55055 1770
rect 55015 1730 55020 1760
rect 55050 1730 55055 1760
rect 55015 1720 55055 1730
rect 55015 1690 55020 1720
rect 55050 1690 55055 1720
rect 55015 1685 55055 1690
rect 55125 1800 55165 1805
rect 55125 1770 55130 1800
rect 55160 1770 55165 1800
rect 55125 1760 55165 1770
rect 55125 1730 55130 1760
rect 55160 1730 55165 1760
rect 55125 1720 55165 1730
rect 55125 1690 55130 1720
rect 55160 1690 55165 1720
rect 55125 1685 55165 1690
rect 55235 1800 55275 1805
rect 55235 1770 55240 1800
rect 55270 1770 55275 1800
rect 55235 1760 55275 1770
rect 55235 1730 55240 1760
rect 55270 1730 55275 1760
rect 55235 1720 55275 1730
rect 55235 1690 55240 1720
rect 55270 1690 55275 1720
rect 55235 1685 55275 1690
rect 55345 1800 55385 1805
rect 55345 1770 55350 1800
rect 55380 1770 55385 1800
rect 55345 1760 55385 1770
rect 55345 1730 55350 1760
rect 55380 1730 55385 1760
rect 55345 1720 55385 1730
rect 55345 1690 55350 1720
rect 55380 1690 55385 1720
rect 55345 1685 55385 1690
rect 54745 1655 54750 1675
rect 54770 1655 54775 1675
rect 54745 1615 54775 1655
rect 54745 1445 54750 1615
rect 54770 1445 54775 1615
rect 54745 1435 54775 1445
rect 54800 1615 54830 1685
rect 54850 1665 54890 1670
rect 54850 1635 54855 1665
rect 54885 1635 54890 1665
rect 54850 1630 54890 1635
rect 54800 1445 54805 1615
rect 54825 1445 54830 1615
rect 54800 1435 54830 1445
rect 54855 1615 54885 1630
rect 54855 1445 54860 1615
rect 54880 1445 54885 1615
rect 54855 1415 54885 1445
rect 54910 1615 54940 1685
rect 54960 1665 55000 1670
rect 54960 1635 54965 1665
rect 54995 1635 55000 1665
rect 54960 1630 55000 1635
rect 54910 1445 54915 1615
rect 54935 1445 54940 1615
rect 54910 1435 54940 1445
rect 54965 1615 54995 1630
rect 54965 1445 54970 1615
rect 54990 1445 54995 1615
rect 54965 1415 54995 1445
rect 55020 1615 55050 1685
rect 55070 1665 55110 1670
rect 55070 1635 55075 1665
rect 55105 1635 55110 1665
rect 55070 1630 55110 1635
rect 55020 1445 55025 1615
rect 55045 1445 55050 1615
rect 55020 1435 55050 1445
rect 55075 1615 55105 1630
rect 55075 1445 55080 1615
rect 55100 1445 55105 1615
rect 55075 1415 55105 1445
rect 55130 1615 55160 1685
rect 55180 1665 55220 1670
rect 55180 1635 55185 1665
rect 55215 1635 55220 1665
rect 55180 1630 55220 1635
rect 55130 1445 55135 1615
rect 55155 1445 55160 1615
rect 55130 1435 55160 1445
rect 55185 1615 55215 1630
rect 55185 1445 55190 1615
rect 55210 1445 55215 1615
rect 55185 1415 55215 1445
rect 55240 1615 55270 1685
rect 55290 1665 55330 1670
rect 55290 1635 55295 1665
rect 55325 1635 55330 1665
rect 55290 1630 55330 1635
rect 55240 1445 55245 1615
rect 55265 1445 55270 1615
rect 55240 1435 55270 1445
rect 55295 1615 55325 1630
rect 55295 1445 55300 1615
rect 55320 1445 55325 1615
rect 55295 1415 55325 1445
rect 55350 1615 55380 1685
rect 55350 1445 55355 1615
rect 55375 1445 55380 1615
rect 55350 1435 55380 1445
rect 55405 1675 55435 1820
rect 55405 1655 55410 1675
rect 55430 1655 55435 1675
rect 55405 1615 55435 1655
rect 55405 1445 55410 1615
rect 55430 1445 55435 1615
rect 55405 1435 55435 1445
rect 54600 1410 54640 1415
rect 54600 1380 54605 1410
rect 54635 1380 54640 1410
rect 54600 1375 54640 1380
rect 54850 1410 54890 1415
rect 54850 1380 54855 1410
rect 54885 1380 54890 1410
rect 54850 1375 54890 1380
rect 54960 1410 55000 1415
rect 54960 1380 54965 1410
rect 54995 1380 55000 1410
rect 54960 1375 55000 1380
rect 55070 1410 55110 1415
rect 55070 1380 55075 1410
rect 55105 1380 55110 1410
rect 55070 1375 55110 1380
rect 55180 1410 55220 1415
rect 55180 1380 55185 1410
rect 55215 1380 55220 1410
rect 55180 1375 55220 1380
rect 55290 1410 55330 1415
rect 55290 1380 55295 1410
rect 55325 1380 55330 1410
rect 55290 1375 55330 1380
rect 54105 1330 54115 1360
rect 54145 1330 54165 1360
rect 54195 1330 54215 1360
rect 54245 1330 54265 1360
rect 54295 1330 54315 1360
rect 54345 1330 54355 1360
rect 54105 1310 54355 1330
rect 54105 1280 54115 1310
rect 54145 1280 54165 1310
rect 54195 1280 54215 1310
rect 54245 1280 54265 1310
rect 54295 1280 54315 1310
rect 54345 1280 54355 1310
rect 54105 1260 54355 1280
rect 54105 1230 54115 1260
rect 54145 1230 54165 1260
rect 54195 1230 54215 1260
rect 54245 1230 54265 1260
rect 54295 1230 54315 1260
rect 54345 1230 54355 1260
rect 54105 310 54355 1230
rect 54380 910 54415 916
rect 54380 870 54415 875
rect 54440 910 54475 915
rect 54440 870 54475 875
rect 54500 910 54535 915
rect 54500 870 54535 875
rect 54560 910 54595 915
rect 54560 870 54595 875
rect 54390 560 54410 870
rect 54510 840 54530 870
rect 54610 840 54630 1375
rect 55235 1345 55275 1350
rect 55235 1315 55240 1345
rect 55270 1315 55275 1345
rect 55235 1305 55275 1315
rect 55235 1275 55240 1305
rect 55270 1275 55275 1305
rect 55235 1270 55275 1275
rect 55520 1345 55640 2110
rect 55520 1315 55525 1345
rect 55555 1315 55565 1345
rect 55595 1315 55605 1345
rect 55635 1315 55640 1345
rect 55520 1305 55640 1315
rect 55520 1275 55525 1305
rect 55555 1275 55565 1305
rect 55595 1275 55605 1305
rect 55635 1275 55640 1305
rect 55520 1270 55640 1275
rect 55660 3105 55780 4210
rect 56005 3935 56765 3940
rect 56005 3905 56010 3935
rect 56040 3905 56050 3935
rect 56080 3905 56090 3935
rect 56120 3905 56130 3935
rect 56160 3905 56170 3935
rect 56200 3905 56210 3935
rect 56240 3905 56250 3935
rect 56280 3905 56290 3935
rect 56320 3905 56330 3935
rect 56360 3905 56370 3935
rect 56400 3905 56410 3935
rect 56440 3905 56450 3935
rect 56480 3905 56490 3935
rect 56520 3905 56530 3935
rect 56560 3905 56570 3935
rect 56600 3905 56610 3935
rect 56640 3905 56650 3935
rect 56680 3905 56690 3935
rect 56720 3905 56730 3935
rect 56760 3905 56765 3935
rect 56005 3895 56765 3905
rect 56005 3865 56010 3895
rect 56040 3865 56050 3895
rect 56080 3865 56090 3895
rect 56120 3865 56130 3895
rect 56160 3865 56170 3895
rect 56200 3865 56210 3895
rect 56240 3865 56250 3895
rect 56280 3865 56290 3895
rect 56320 3865 56330 3895
rect 56360 3865 56370 3895
rect 56400 3865 56410 3895
rect 56440 3865 56450 3895
rect 56480 3865 56490 3895
rect 56520 3865 56530 3895
rect 56560 3865 56570 3895
rect 56600 3865 56610 3895
rect 56640 3865 56650 3895
rect 56680 3865 56690 3895
rect 56720 3865 56730 3895
rect 56760 3865 56765 3895
rect 56005 3855 56765 3865
rect 56005 3825 56010 3855
rect 56040 3825 56050 3855
rect 56080 3825 56090 3855
rect 56120 3825 56130 3855
rect 56160 3825 56170 3855
rect 56200 3825 56210 3855
rect 56240 3825 56250 3855
rect 56280 3825 56290 3855
rect 56320 3825 56330 3855
rect 56360 3825 56370 3855
rect 56400 3825 56410 3855
rect 56440 3825 56450 3855
rect 56480 3825 56490 3855
rect 56520 3825 56530 3855
rect 56560 3825 56570 3855
rect 56600 3825 56610 3855
rect 56640 3825 56650 3855
rect 56680 3825 56690 3855
rect 56720 3825 56730 3855
rect 56760 3825 56765 3855
rect 56005 3820 56765 3825
rect 56010 3750 56040 3820
rect 56065 3800 56105 3805
rect 56065 3770 56070 3800
rect 56100 3770 56105 3800
rect 56065 3765 56105 3770
rect 56010 3430 56015 3750
rect 56035 3430 56040 3750
rect 56010 3390 56040 3430
rect 56070 3750 56100 3765
rect 56070 3430 56075 3750
rect 56095 3430 56100 3750
rect 56070 3415 56100 3430
rect 56130 3750 56160 3820
rect 56185 3800 56225 3805
rect 56185 3770 56190 3800
rect 56220 3770 56225 3800
rect 56185 3765 56225 3770
rect 56130 3430 56135 3750
rect 56155 3430 56160 3750
rect 56130 3420 56160 3430
rect 56190 3750 56220 3765
rect 56190 3430 56195 3750
rect 56215 3430 56220 3750
rect 56190 3415 56220 3430
rect 56250 3750 56280 3820
rect 56305 3800 56345 3805
rect 56305 3770 56310 3800
rect 56340 3770 56345 3800
rect 56305 3765 56345 3770
rect 56250 3430 56255 3750
rect 56275 3430 56280 3750
rect 56250 3420 56280 3430
rect 56310 3750 56340 3765
rect 56310 3430 56315 3750
rect 56335 3430 56340 3750
rect 56310 3415 56340 3430
rect 56370 3750 56400 3820
rect 56425 3800 56465 3805
rect 56425 3770 56430 3800
rect 56460 3770 56465 3800
rect 56425 3765 56465 3770
rect 56370 3430 56375 3750
rect 56395 3430 56400 3750
rect 56370 3420 56400 3430
rect 56430 3750 56460 3765
rect 56430 3430 56435 3750
rect 56455 3430 56460 3750
rect 56430 3415 56460 3430
rect 56490 3750 56520 3820
rect 56545 3800 56585 3805
rect 56545 3770 56550 3800
rect 56580 3770 56585 3800
rect 56545 3765 56585 3770
rect 56490 3430 56495 3750
rect 56515 3430 56520 3750
rect 56490 3420 56520 3430
rect 56550 3750 56580 3765
rect 56550 3430 56555 3750
rect 56575 3430 56580 3750
rect 56550 3415 56580 3430
rect 56610 3750 56640 3820
rect 56665 3800 56705 3805
rect 56665 3770 56670 3800
rect 56700 3770 56705 3800
rect 56665 3765 56705 3770
rect 56610 3430 56615 3750
rect 56635 3430 56640 3750
rect 56610 3420 56640 3430
rect 56670 3750 56700 3765
rect 56670 3430 56675 3750
rect 56695 3430 56700 3750
rect 56670 3415 56700 3430
rect 56730 3750 56760 3820
rect 56730 3430 56735 3750
rect 56755 3430 56760 3750
rect 56010 3370 56015 3390
rect 56035 3370 56040 3390
rect 56010 3360 56040 3370
rect 56065 3410 56105 3415
rect 56065 3380 56070 3410
rect 56100 3380 56105 3410
rect 56065 3245 56105 3380
rect 56185 3410 56225 3415
rect 56185 3380 56190 3410
rect 56220 3380 56225 3410
rect 56185 3245 56225 3380
rect 56305 3410 56345 3415
rect 56305 3380 56310 3410
rect 56340 3380 56345 3410
rect 56305 3245 56345 3380
rect 56425 3410 56465 3415
rect 56425 3380 56430 3410
rect 56460 3380 56465 3410
rect 56365 3330 56405 3335
rect 56365 3300 56370 3330
rect 56400 3300 56405 3330
rect 56365 3295 56405 3300
rect 56425 3245 56465 3380
rect 56545 3410 56585 3415
rect 56545 3380 56550 3410
rect 56580 3380 56585 3410
rect 56545 3245 56585 3380
rect 56665 3410 56705 3415
rect 56665 3380 56670 3410
rect 56700 3380 56705 3410
rect 56665 3245 56705 3380
rect 56730 3390 56760 3430
rect 56730 3370 56735 3390
rect 56755 3370 56760 3390
rect 56730 3360 56760 3370
rect 56845 3335 56865 4445
rect 56880 4320 56920 4730
rect 57030 4865 57060 4895
rect 57030 4545 57035 4865
rect 57055 4545 57060 4865
rect 57030 4535 57060 4545
rect 57090 4865 57120 5030
rect 57145 5010 57185 5015
rect 57145 4980 57150 5010
rect 57180 4980 57185 5010
rect 57145 4970 57185 4980
rect 57145 4940 57150 4970
rect 57180 4940 57185 4970
rect 57145 4930 57185 4940
rect 57145 4900 57150 4930
rect 57180 4900 57185 4930
rect 57145 4895 57185 4900
rect 57205 5010 57245 5015
rect 57205 4980 57210 5010
rect 57240 4980 57245 5010
rect 57205 4970 57245 4980
rect 57205 4940 57210 4970
rect 57240 4940 57245 4970
rect 57205 4930 57245 4940
rect 57205 4900 57210 4930
rect 57240 4900 57245 4930
rect 57205 4895 57245 4900
rect 57495 4930 57535 4935
rect 57495 4900 57500 4930
rect 57530 4900 57535 4930
rect 57495 4895 57535 4900
rect 57555 4930 57595 5035
rect 57555 4900 57560 4930
rect 57590 4900 57595 4930
rect 57555 4895 57595 4900
rect 57675 4930 57715 4935
rect 57675 4900 57680 4930
rect 57710 4900 57715 4930
rect 57675 4895 57715 4900
rect 57090 4545 57095 4865
rect 57115 4545 57120 4865
rect 57090 4530 57120 4545
rect 57150 4865 57180 4895
rect 57150 4545 57155 4865
rect 57175 4545 57180 4865
rect 57150 4535 57180 4545
rect 57210 4865 57240 4895
rect 57210 4545 57215 4865
rect 57235 4545 57240 4865
rect 57210 4535 57240 4545
rect 57500 4865 57530 4895
rect 57500 4545 57505 4865
rect 57525 4545 57530 4865
rect 57500 4535 57530 4545
rect 57560 4865 57590 4895
rect 57560 4545 57565 4865
rect 57585 4545 57590 4865
rect 57560 4530 57590 4545
rect 57620 4865 57650 4875
rect 57620 4545 57625 4865
rect 57645 4545 57650 4865
rect 57085 4525 57125 4530
rect 57085 4495 57090 4525
rect 57120 4495 57125 4525
rect 57085 4490 57125 4495
rect 57555 4525 57595 4530
rect 57555 4495 57560 4525
rect 57590 4495 57595 4525
rect 57555 4490 57595 4495
rect 57140 4475 57170 4485
rect 57140 4455 57145 4475
rect 57165 4455 57170 4475
rect 56880 4290 56885 4320
rect 56915 4290 56920 4320
rect 56880 4280 56920 4290
rect 56880 4250 56885 4280
rect 56915 4250 56920 4280
rect 56880 4240 56920 4250
rect 56880 4210 56885 4240
rect 56915 4210 56920 4240
rect 56880 4205 56920 4210
rect 56935 4425 56975 4430
rect 56935 4395 56940 4425
rect 56970 4395 56975 4425
rect 57140 4420 57170 4455
rect 57576 4470 57606 4475
rect 57576 4435 57606 4440
rect 57620 4420 57650 4545
rect 57680 4865 57710 4895
rect 57680 4545 57685 4865
rect 57705 4545 57710 4865
rect 57680 4535 57710 4545
rect 56935 4390 56975 4395
rect 57135 4415 57175 4420
rect 56835 3330 56875 3335
rect 56835 3300 56840 3330
rect 56870 3300 56875 3330
rect 56835 3295 56875 3300
rect 56935 3290 56955 4390
rect 57135 4385 57140 4415
rect 57170 4385 57175 4415
rect 57135 4380 57175 4385
rect 57615 4415 57655 4420
rect 57615 4385 57620 4415
rect 57650 4385 57655 4415
rect 57615 4380 57655 4385
rect 58100 4320 58220 4325
rect 58100 4290 58105 4320
rect 58135 4290 58145 4320
rect 58175 4290 58185 4320
rect 58215 4290 58220 4320
rect 58100 4280 58220 4290
rect 58100 4250 58105 4280
rect 58135 4250 58145 4280
rect 58175 4250 58185 4280
rect 58215 4250 58220 4280
rect 58100 4240 58220 4250
rect 58100 4210 58105 4240
rect 58135 4210 58145 4240
rect 58175 4210 58185 4240
rect 58215 4210 58220 4240
rect 57035 3935 57795 3940
rect 57035 3905 57040 3935
rect 57070 3905 57080 3935
rect 57110 3905 57120 3935
rect 57150 3905 57160 3935
rect 57190 3905 57200 3935
rect 57230 3905 57240 3935
rect 57270 3905 57280 3935
rect 57310 3905 57320 3935
rect 57350 3905 57360 3935
rect 57390 3905 57400 3935
rect 57430 3905 57440 3935
rect 57470 3905 57480 3935
rect 57510 3905 57520 3935
rect 57550 3905 57560 3935
rect 57590 3905 57600 3935
rect 57630 3905 57640 3935
rect 57670 3905 57680 3935
rect 57710 3905 57720 3935
rect 57750 3905 57760 3935
rect 57790 3905 57795 3935
rect 57035 3895 57795 3905
rect 57035 3865 57040 3895
rect 57070 3865 57080 3895
rect 57110 3865 57120 3895
rect 57150 3865 57160 3895
rect 57190 3865 57200 3895
rect 57230 3865 57240 3895
rect 57270 3865 57280 3895
rect 57310 3865 57320 3895
rect 57350 3865 57360 3895
rect 57390 3865 57400 3895
rect 57430 3865 57440 3895
rect 57470 3865 57480 3895
rect 57510 3865 57520 3895
rect 57550 3865 57560 3895
rect 57590 3865 57600 3895
rect 57630 3865 57640 3895
rect 57670 3865 57680 3895
rect 57710 3865 57720 3895
rect 57750 3865 57760 3895
rect 57790 3865 57795 3895
rect 57035 3855 57795 3865
rect 57035 3825 57040 3855
rect 57070 3825 57080 3855
rect 57110 3825 57120 3855
rect 57150 3825 57160 3855
rect 57190 3825 57200 3855
rect 57230 3825 57240 3855
rect 57270 3825 57280 3855
rect 57310 3825 57320 3855
rect 57350 3825 57360 3855
rect 57390 3825 57400 3855
rect 57430 3825 57440 3855
rect 57470 3825 57480 3855
rect 57510 3825 57520 3855
rect 57550 3825 57560 3855
rect 57590 3825 57600 3855
rect 57630 3825 57640 3855
rect 57670 3825 57680 3855
rect 57710 3825 57720 3855
rect 57750 3825 57760 3855
rect 57790 3825 57795 3855
rect 57035 3820 57795 3825
rect 57040 3750 57070 3820
rect 57095 3800 57135 3805
rect 57095 3770 57100 3800
rect 57130 3770 57135 3800
rect 57095 3765 57135 3770
rect 57040 3430 57045 3750
rect 57065 3430 57070 3750
rect 57040 3390 57070 3430
rect 57100 3750 57130 3765
rect 57100 3430 57105 3750
rect 57125 3430 57130 3750
rect 57100 3415 57130 3430
rect 57160 3750 57190 3820
rect 57215 3800 57255 3805
rect 57215 3770 57220 3800
rect 57250 3770 57255 3800
rect 57215 3765 57255 3770
rect 57160 3430 57165 3750
rect 57185 3430 57190 3750
rect 57160 3420 57190 3430
rect 57220 3750 57250 3765
rect 57220 3430 57225 3750
rect 57245 3430 57250 3750
rect 57220 3415 57250 3430
rect 57280 3750 57310 3820
rect 57335 3800 57375 3805
rect 57335 3770 57340 3800
rect 57370 3770 57375 3800
rect 57335 3765 57375 3770
rect 57280 3430 57285 3750
rect 57305 3430 57310 3750
rect 57280 3420 57310 3430
rect 57340 3750 57370 3765
rect 57340 3430 57345 3750
rect 57365 3430 57370 3750
rect 57340 3415 57370 3430
rect 57400 3750 57430 3820
rect 57455 3800 57495 3805
rect 57455 3770 57460 3800
rect 57490 3770 57495 3800
rect 57455 3765 57495 3770
rect 57400 3430 57405 3750
rect 57425 3430 57430 3750
rect 57400 3420 57430 3430
rect 57460 3750 57490 3765
rect 57460 3430 57465 3750
rect 57485 3430 57490 3750
rect 57460 3415 57490 3430
rect 57520 3750 57550 3820
rect 57575 3800 57615 3805
rect 57575 3770 57580 3800
rect 57610 3770 57615 3800
rect 57575 3765 57615 3770
rect 57520 3430 57525 3750
rect 57545 3430 57550 3750
rect 57520 3420 57550 3430
rect 57580 3750 57610 3765
rect 57580 3430 57585 3750
rect 57605 3430 57610 3750
rect 57580 3415 57610 3430
rect 57640 3750 57670 3820
rect 57695 3800 57735 3805
rect 57695 3770 57700 3800
rect 57730 3770 57735 3800
rect 57695 3765 57735 3770
rect 57640 3430 57645 3750
rect 57665 3430 57670 3750
rect 57640 3420 57670 3430
rect 57700 3750 57730 3765
rect 57700 3430 57705 3750
rect 57725 3430 57730 3750
rect 57700 3415 57730 3430
rect 57760 3750 57790 3820
rect 57760 3430 57765 3750
rect 57785 3430 57790 3750
rect 57040 3370 57045 3390
rect 57065 3370 57070 3390
rect 57040 3360 57070 3370
rect 57095 3410 57135 3415
rect 57095 3380 57100 3410
rect 57130 3380 57135 3410
rect 56925 3285 56965 3290
rect 56925 3255 56930 3285
rect 56960 3255 56965 3285
rect 56925 3250 56965 3255
rect 56065 3240 56705 3245
rect 56065 3210 56070 3240
rect 56100 3210 56110 3240
rect 56140 3210 56150 3240
rect 56180 3210 56190 3240
rect 56220 3210 56230 3240
rect 56260 3210 56270 3240
rect 56300 3210 56310 3240
rect 56340 3210 56350 3240
rect 56380 3210 56390 3240
rect 56420 3210 56430 3240
rect 56460 3210 56470 3240
rect 56500 3210 56510 3240
rect 56540 3210 56550 3240
rect 56580 3210 56590 3240
rect 56620 3210 56630 3240
rect 56660 3210 56670 3240
rect 56700 3210 56705 3240
rect 56065 3200 56705 3210
rect 56065 3170 56070 3200
rect 56100 3170 56110 3200
rect 56140 3170 56150 3200
rect 56180 3170 56190 3200
rect 56220 3170 56230 3200
rect 56260 3170 56270 3200
rect 56300 3170 56310 3200
rect 56340 3170 56350 3200
rect 56380 3170 56390 3200
rect 56420 3170 56430 3200
rect 56460 3170 56470 3200
rect 56500 3170 56510 3200
rect 56540 3170 56550 3200
rect 56580 3170 56590 3200
rect 56620 3170 56630 3200
rect 56660 3170 56670 3200
rect 56700 3170 56705 3200
rect 56065 3160 56705 3170
rect 56065 3130 56070 3160
rect 56100 3130 56110 3160
rect 56140 3130 56150 3160
rect 56180 3130 56190 3160
rect 56220 3130 56230 3160
rect 56260 3130 56270 3160
rect 56300 3130 56310 3160
rect 56340 3130 56350 3160
rect 56380 3130 56390 3160
rect 56420 3130 56430 3160
rect 56460 3130 56470 3160
rect 56500 3130 56510 3160
rect 56540 3130 56550 3160
rect 56580 3130 56590 3160
rect 56620 3130 56630 3160
rect 56660 3130 56670 3160
rect 56700 3130 56705 3160
rect 56065 3125 56705 3130
rect 57095 3245 57135 3380
rect 57215 3410 57255 3415
rect 57215 3380 57220 3410
rect 57250 3380 57255 3410
rect 57215 3245 57255 3380
rect 57335 3410 57375 3415
rect 57335 3380 57340 3410
rect 57370 3380 57375 3410
rect 57335 3245 57375 3380
rect 57455 3410 57495 3415
rect 57455 3380 57460 3410
rect 57490 3380 57495 3410
rect 57395 3330 57435 3335
rect 57395 3300 57400 3330
rect 57430 3300 57435 3330
rect 57395 3295 57435 3300
rect 57455 3245 57495 3380
rect 57575 3410 57615 3415
rect 57575 3380 57580 3410
rect 57610 3380 57615 3410
rect 57575 3245 57615 3380
rect 57695 3410 57735 3415
rect 57695 3380 57700 3410
rect 57730 3380 57735 3410
rect 57695 3245 57735 3380
rect 57760 3390 57790 3430
rect 57760 3370 57765 3390
rect 57785 3370 57790 3390
rect 57760 3360 57790 3370
rect 57095 3240 57735 3245
rect 57095 3210 57100 3240
rect 57130 3210 57140 3240
rect 57170 3210 57180 3240
rect 57210 3210 57220 3240
rect 57250 3210 57260 3240
rect 57290 3210 57300 3240
rect 57330 3210 57340 3240
rect 57370 3210 57380 3240
rect 57410 3210 57420 3240
rect 57450 3210 57460 3240
rect 57490 3210 57500 3240
rect 57530 3210 57540 3240
rect 57570 3210 57580 3240
rect 57610 3210 57620 3240
rect 57650 3210 57660 3240
rect 57690 3210 57700 3240
rect 57730 3210 57735 3240
rect 57095 3200 57735 3210
rect 57095 3170 57100 3200
rect 57130 3170 57140 3200
rect 57170 3170 57180 3200
rect 57210 3170 57220 3200
rect 57250 3170 57260 3200
rect 57290 3170 57300 3200
rect 57330 3170 57340 3200
rect 57370 3170 57380 3200
rect 57410 3170 57420 3200
rect 57450 3170 57460 3200
rect 57490 3170 57500 3200
rect 57530 3170 57540 3200
rect 57570 3170 57580 3200
rect 57610 3170 57620 3200
rect 57650 3170 57660 3200
rect 57690 3170 57700 3200
rect 57730 3170 57735 3200
rect 57095 3160 57735 3170
rect 57095 3130 57100 3160
rect 57130 3130 57140 3160
rect 57170 3130 57180 3160
rect 57210 3130 57220 3160
rect 57250 3130 57260 3160
rect 57290 3130 57300 3160
rect 57330 3130 57340 3160
rect 57370 3130 57380 3160
rect 57410 3130 57420 3160
rect 57450 3130 57460 3160
rect 57490 3130 57500 3160
rect 57530 3130 57540 3160
rect 57570 3130 57580 3160
rect 57610 3130 57620 3160
rect 57650 3130 57660 3160
rect 57690 3130 57700 3160
rect 57730 3130 57735 3160
rect 57095 3125 57735 3130
rect 55660 3075 55665 3105
rect 55695 3075 55705 3105
rect 55735 3075 55745 3105
rect 55775 3075 55780 3105
rect 58100 3105 58220 4210
rect 58410 4320 58450 4325
rect 58410 4290 58415 4320
rect 58445 4290 58450 4320
rect 58410 4280 58450 4290
rect 58410 4250 58415 4280
rect 58445 4250 58450 4280
rect 58410 4240 58450 4250
rect 58410 4210 58415 4240
rect 58445 4210 58450 4240
rect 58410 3800 58450 4210
rect 58770 4320 58810 4325
rect 58770 4290 58775 4320
rect 58805 4290 58810 4320
rect 58770 4280 58810 4290
rect 58770 4250 58775 4280
rect 58805 4250 58810 4280
rect 58770 4240 58810 4250
rect 58770 4210 58775 4240
rect 58805 4210 58810 4240
rect 58470 3935 58750 3940
rect 58470 3905 58475 3935
rect 58505 3905 58515 3935
rect 58545 3905 58555 3935
rect 58585 3905 58595 3935
rect 58625 3905 58635 3935
rect 58665 3905 58675 3935
rect 58705 3905 58715 3935
rect 58745 3905 58750 3935
rect 58470 3895 58750 3905
rect 58470 3865 58475 3895
rect 58505 3865 58515 3895
rect 58545 3865 58555 3895
rect 58585 3865 58595 3895
rect 58625 3865 58635 3895
rect 58665 3865 58675 3895
rect 58705 3865 58715 3895
rect 58745 3865 58750 3895
rect 58470 3855 58750 3865
rect 58470 3825 58475 3855
rect 58505 3825 58515 3855
rect 58545 3825 58555 3855
rect 58585 3825 58595 3855
rect 58625 3825 58635 3855
rect 58665 3825 58675 3855
rect 58705 3825 58715 3855
rect 58745 3825 58750 3855
rect 58470 3820 58750 3825
rect 58410 3770 58415 3800
rect 58445 3770 58450 3800
rect 58410 3765 58450 3770
rect 58415 3750 58445 3765
rect 58415 3430 58420 3750
rect 58440 3430 58445 3750
rect 58415 3390 58445 3430
rect 58475 3750 58505 3820
rect 58530 3800 58570 3805
rect 58530 3770 58535 3800
rect 58565 3770 58570 3800
rect 58530 3765 58570 3770
rect 58475 3430 58480 3750
rect 58500 3430 58505 3750
rect 58475 3415 58505 3430
rect 58535 3750 58565 3765
rect 58535 3430 58540 3750
rect 58560 3430 58565 3750
rect 58535 3420 58565 3430
rect 58595 3750 58625 3820
rect 58650 3800 58690 3805
rect 58650 3770 58655 3800
rect 58685 3770 58690 3800
rect 58650 3765 58690 3770
rect 58595 3430 58600 3750
rect 58620 3430 58625 3750
rect 58595 3415 58625 3430
rect 58655 3750 58685 3765
rect 58655 3430 58660 3750
rect 58680 3430 58685 3750
rect 58655 3420 58685 3430
rect 58715 3750 58745 3820
rect 58770 3800 58810 4210
rect 59130 4320 59170 4325
rect 59130 4290 59135 4320
rect 59165 4290 59170 4320
rect 59130 4280 59170 4290
rect 59130 4250 59135 4280
rect 59165 4250 59170 4280
rect 59130 4240 59170 4250
rect 59130 4210 59135 4240
rect 59165 4210 59170 4240
rect 58830 3935 59110 3940
rect 58830 3905 58835 3935
rect 58865 3905 58875 3935
rect 58905 3905 58915 3935
rect 58945 3905 58955 3935
rect 58985 3905 58995 3935
rect 59025 3905 59035 3935
rect 59065 3905 59075 3935
rect 59105 3905 59110 3935
rect 58830 3895 59110 3905
rect 58830 3865 58835 3895
rect 58865 3865 58875 3895
rect 58905 3865 58915 3895
rect 58945 3865 58955 3895
rect 58985 3865 58995 3895
rect 59025 3865 59035 3895
rect 59065 3865 59075 3895
rect 59105 3865 59110 3895
rect 58830 3855 59110 3865
rect 58830 3825 58835 3855
rect 58865 3825 58875 3855
rect 58905 3825 58915 3855
rect 58945 3825 58955 3855
rect 58985 3825 58995 3855
rect 59025 3825 59035 3855
rect 59065 3825 59075 3855
rect 59105 3825 59110 3855
rect 58830 3820 59110 3825
rect 58770 3770 58775 3800
rect 58805 3770 58810 3800
rect 58770 3765 58810 3770
rect 58715 3430 58720 3750
rect 58740 3430 58745 3750
rect 58715 3415 58745 3430
rect 58775 3750 58805 3765
rect 58775 3430 58780 3750
rect 58800 3430 58805 3750
rect 58775 3420 58805 3430
rect 58835 3750 58865 3820
rect 58890 3800 58930 3805
rect 58890 3770 58895 3800
rect 58925 3770 58930 3800
rect 58890 3765 58930 3770
rect 58835 3430 58840 3750
rect 58860 3430 58865 3750
rect 58835 3415 58865 3430
rect 58895 3750 58925 3765
rect 58895 3430 58900 3750
rect 58920 3430 58925 3750
rect 58895 3420 58925 3430
rect 58955 3750 58985 3820
rect 59010 3800 59050 3805
rect 59010 3770 59015 3800
rect 59045 3770 59050 3800
rect 59010 3765 59050 3770
rect 58955 3430 58960 3750
rect 58980 3430 58985 3750
rect 58955 3415 58985 3430
rect 59015 3750 59045 3765
rect 59015 3430 59020 3750
rect 59040 3430 59045 3750
rect 59015 3420 59045 3430
rect 59075 3750 59105 3820
rect 59130 3800 59170 4210
rect 59640 4320 59760 6460
rect 59640 4290 59645 4320
rect 59675 4290 59685 4320
rect 59715 4290 59725 4320
rect 59755 4290 59760 4320
rect 59640 4280 59760 4290
rect 59640 4250 59645 4280
rect 59675 4250 59685 4280
rect 59715 4250 59725 4280
rect 59755 4250 59760 4280
rect 59640 4240 59760 4250
rect 59640 4210 59645 4240
rect 59675 4210 59685 4240
rect 59715 4210 59725 4240
rect 59755 4210 59760 4240
rect 59640 4205 59760 4210
rect 59990 4320 60110 6460
rect 59990 4290 59995 4320
rect 60025 4290 60035 4320
rect 60065 4290 60075 4320
rect 60105 4290 60110 4320
rect 59990 4280 60110 4290
rect 59990 4250 59995 4280
rect 60025 4250 60035 4280
rect 60065 4250 60075 4280
rect 60105 4250 60110 4280
rect 59990 4240 60110 4250
rect 59990 4210 59995 4240
rect 60025 4210 60035 4240
rect 60065 4210 60075 4240
rect 60105 4210 60110 4240
rect 59990 4205 60110 4210
rect 60690 4320 60810 6460
rect 60690 4290 60695 4320
rect 60725 4290 60735 4320
rect 60765 4290 60775 4320
rect 60805 4290 60810 4320
rect 60690 4280 60810 4290
rect 60690 4250 60695 4280
rect 60725 4250 60735 4280
rect 60765 4250 60775 4280
rect 60805 4250 60810 4280
rect 60690 4240 60810 4250
rect 60690 4210 60695 4240
rect 60725 4210 60735 4240
rect 60765 4210 60775 4240
rect 60805 4210 60810 4240
rect 60690 4205 60810 4210
rect 61040 4320 61160 6460
rect 61040 4290 61045 4320
rect 61075 4290 61085 4320
rect 61115 4290 61125 4320
rect 61155 4290 61160 4320
rect 61040 4280 61160 4290
rect 61040 4250 61045 4280
rect 61075 4250 61085 4280
rect 61115 4250 61125 4280
rect 61155 4250 61160 4280
rect 61040 4240 61160 4250
rect 61040 4210 61045 4240
rect 61075 4210 61085 4240
rect 61115 4210 61125 4240
rect 61155 4210 61160 4240
rect 61040 4205 61160 4210
rect 61390 4320 61510 6460
rect 61390 4290 61395 4320
rect 61425 4290 61435 4320
rect 61465 4290 61475 4320
rect 61505 4290 61510 4320
rect 61390 4280 61510 4290
rect 61390 4250 61395 4280
rect 61425 4250 61435 4280
rect 61465 4250 61475 4280
rect 61505 4250 61510 4280
rect 61390 4240 61510 4250
rect 61390 4210 61395 4240
rect 61425 4210 61435 4240
rect 61465 4210 61475 4240
rect 61505 4210 61510 4240
rect 61390 4205 61510 4210
rect 59130 3770 59135 3800
rect 59165 3770 59170 3800
rect 59130 3765 59170 3770
rect 59075 3430 59080 3750
rect 59100 3430 59105 3750
rect 59075 3415 59105 3430
rect 59135 3750 59165 3765
rect 59135 3430 59140 3750
rect 59160 3430 59165 3750
rect 58415 3370 58420 3390
rect 58440 3370 58445 3390
rect 58470 3410 58510 3415
rect 58470 3380 58475 3410
rect 58505 3380 58510 3410
rect 58470 3375 58510 3380
rect 58590 3410 58630 3415
rect 58590 3380 58595 3410
rect 58625 3380 58630 3410
rect 58590 3375 58630 3380
rect 58710 3410 58750 3415
rect 58710 3380 58715 3410
rect 58745 3380 58750 3410
rect 58710 3375 58750 3380
rect 58830 3410 58870 3415
rect 58830 3380 58835 3410
rect 58865 3380 58870 3410
rect 58830 3375 58870 3380
rect 58950 3410 58990 3415
rect 58950 3380 58955 3410
rect 58985 3380 58990 3410
rect 58950 3375 58990 3380
rect 59070 3410 59110 3415
rect 59070 3380 59075 3410
rect 59105 3380 59110 3410
rect 59070 3375 59110 3380
rect 59135 3390 59165 3430
rect 58415 3360 58445 3370
rect 59135 3370 59140 3390
rect 59160 3370 59165 3390
rect 59135 3360 59165 3370
rect 58770 3285 58810 3290
rect 58770 3255 58775 3285
rect 58805 3255 58810 3285
rect 58770 3250 58810 3255
rect 55660 3065 55780 3075
rect 55660 3035 55665 3065
rect 55695 3035 55705 3065
rect 55735 3035 55745 3065
rect 55775 3035 55780 3065
rect 55660 3025 55780 3035
rect 55660 2995 55665 3025
rect 55695 2995 55705 3025
rect 55735 2995 55745 3025
rect 55775 2995 55780 3025
rect 55660 1935 55780 2995
rect 56510 3095 56550 3100
rect 56510 3065 56515 3095
rect 56545 3065 56550 3095
rect 56510 3055 56550 3065
rect 56510 3025 56515 3055
rect 56545 3025 56550 3055
rect 56510 3015 56550 3025
rect 56510 2985 56515 3015
rect 56545 2985 56550 3015
rect 56510 2980 56550 2985
rect 56680 3095 56710 3100
rect 56680 3055 56710 3065
rect 56680 3015 56710 3025
rect 56680 2980 56710 2985
rect 56840 3095 56880 3100
rect 56840 3065 56845 3095
rect 56875 3065 56880 3095
rect 56840 3055 56880 3065
rect 56840 3025 56845 3055
rect 56875 3025 56880 3055
rect 56840 3015 56880 3025
rect 56840 2985 56845 3015
rect 56875 2985 56880 3015
rect 56840 2980 56880 2985
rect 56920 3095 56960 3100
rect 56920 3065 56925 3095
rect 56955 3065 56960 3095
rect 56920 3055 56960 3065
rect 56920 3025 56925 3055
rect 56955 3025 56960 3055
rect 56920 3015 56960 3025
rect 56920 2985 56925 3015
rect 56955 2985 56960 3015
rect 56920 2980 56960 2985
rect 57090 3095 57120 3100
rect 57090 3055 57120 3065
rect 57090 3015 57120 3025
rect 57090 2980 57120 2985
rect 57250 3095 57290 3100
rect 57250 3065 57255 3095
rect 57285 3065 57290 3095
rect 57250 3055 57290 3065
rect 57250 3025 57255 3055
rect 57285 3025 57290 3055
rect 57250 3015 57290 3025
rect 57250 2985 57255 3015
rect 57285 2985 57290 3015
rect 57250 2980 57290 2985
rect 58100 3075 58105 3105
rect 58135 3075 58145 3105
rect 58175 3075 58185 3105
rect 58215 3075 58220 3105
rect 58100 3065 58220 3075
rect 58100 3035 58105 3065
rect 58135 3035 58145 3065
rect 58175 3035 58185 3065
rect 58215 3035 58220 3065
rect 58100 3025 58220 3035
rect 58100 2995 58105 3025
rect 58135 2995 58145 3025
rect 58175 2995 58185 3025
rect 58215 2995 58220 3025
rect 56620 2960 56660 2965
rect 56620 2930 56625 2960
rect 56655 2930 56660 2960
rect 56620 2925 56660 2930
rect 56730 2960 56770 2965
rect 56730 2930 56735 2960
rect 56765 2930 56770 2960
rect 56730 2925 56770 2930
rect 57030 2960 57070 2965
rect 57030 2930 57035 2960
rect 57065 2930 57070 2960
rect 57030 2925 57070 2930
rect 57140 2960 57180 2965
rect 57140 2930 57145 2960
rect 57175 2930 57180 2960
rect 57140 2925 57180 2930
rect 56560 2650 56590 2655
rect 56800 2650 56830 2655
rect 56560 2615 56590 2620
rect 56607 2635 56637 2645
rect 56607 2615 56612 2635
rect 56632 2615 56637 2635
rect 56607 2605 56637 2615
rect 56675 2640 56715 2645
rect 56675 2610 56680 2640
rect 56710 2610 56715 2640
rect 56675 2605 56715 2610
rect 56753 2635 56783 2645
rect 56753 2615 56758 2635
rect 56778 2615 56783 2635
rect 56800 2615 56830 2620
rect 56970 2645 57000 2655
rect 57210 2645 57240 2655
rect 56970 2625 56975 2645
rect 56995 2625 57000 2645
rect 56970 2615 57000 2625
rect 57017 2635 57047 2645
rect 57017 2615 57022 2635
rect 57042 2615 57047 2635
rect 56753 2605 56783 2615
rect 56610 2585 56630 2605
rect 56600 2580 56640 2585
rect 56600 2550 56605 2580
rect 56635 2550 56640 2580
rect 56600 2545 56640 2550
rect 56760 2535 56780 2605
rect 55940 2530 55980 2535
rect 55940 2500 55945 2530
rect 55975 2500 55980 2530
rect 55940 2495 55980 2500
rect 56745 2530 56785 2535
rect 56745 2500 56750 2530
rect 56780 2500 56785 2530
rect 56745 2495 56785 2500
rect 55660 1905 55665 1935
rect 55695 1905 55705 1935
rect 55735 1905 55745 1935
rect 55775 1905 55780 1935
rect 55660 1895 55780 1905
rect 55660 1865 55665 1895
rect 55695 1865 55705 1895
rect 55735 1865 55745 1895
rect 55775 1865 55780 1895
rect 55660 1855 55780 1865
rect 55660 1825 55665 1855
rect 55695 1825 55705 1855
rect 55735 1825 55745 1855
rect 55775 1825 55780 1855
rect 54645 1225 54685 1230
rect 54645 1195 54650 1225
rect 54680 1195 54685 1225
rect 54645 1190 54685 1195
rect 54850 1225 54890 1230
rect 54850 1195 54855 1225
rect 54885 1195 54890 1225
rect 54850 1190 54890 1195
rect 54960 1225 55000 1230
rect 54960 1195 54965 1225
rect 54995 1195 55000 1225
rect 54960 1190 55000 1195
rect 55070 1225 55110 1230
rect 55070 1195 55075 1225
rect 55105 1195 55110 1225
rect 55070 1190 55110 1195
rect 55180 1225 55220 1230
rect 55180 1195 55185 1225
rect 55215 1195 55220 1225
rect 55180 1190 55220 1195
rect 55290 1225 55330 1230
rect 55290 1195 55295 1225
rect 55325 1195 55330 1225
rect 55290 1190 55330 1195
rect 54655 910 54675 1190
rect 54745 1175 54775 1185
rect 54645 905 54685 910
rect 54645 875 54650 905
rect 54680 875 54685 905
rect 54645 870 54685 875
rect 54745 905 54750 1175
rect 54770 905 54775 1175
rect 54745 865 54775 905
rect 54745 845 54750 865
rect 54770 845 54775 865
rect 54500 835 54540 840
rect 54500 805 54505 835
rect 54535 805 54540 835
rect 54500 800 54540 805
rect 54600 835 54640 840
rect 54600 805 54605 835
rect 54635 805 54640 835
rect 54600 800 54640 805
rect 54745 695 54775 845
rect 54800 1175 54830 1185
rect 54800 905 54805 1175
rect 54825 905 54830 1175
rect 54800 830 54830 905
rect 54855 1175 54885 1190
rect 54855 905 54860 1175
rect 54880 905 54885 1175
rect 54855 890 54885 905
rect 54910 1175 54940 1185
rect 54910 905 54915 1175
rect 54935 905 54940 1175
rect 54850 885 54890 890
rect 54850 855 54855 885
rect 54885 855 54890 885
rect 54850 850 54890 855
rect 54910 830 54940 905
rect 54965 1175 54995 1190
rect 54965 905 54970 1175
rect 54990 905 54995 1175
rect 54965 890 54995 905
rect 55020 1175 55050 1185
rect 55020 905 55025 1175
rect 55045 905 55050 1175
rect 54960 885 55000 890
rect 54960 855 54965 885
rect 54995 855 55000 885
rect 54960 850 55000 855
rect 55020 830 55050 905
rect 55075 1175 55105 1190
rect 55075 905 55080 1175
rect 55100 905 55105 1175
rect 55075 890 55105 905
rect 55130 1175 55160 1185
rect 55130 905 55135 1175
rect 55155 905 55160 1175
rect 55070 885 55110 890
rect 55070 855 55075 885
rect 55105 855 55110 885
rect 55070 850 55110 855
rect 55130 830 55160 905
rect 55185 1175 55215 1190
rect 55185 905 55190 1175
rect 55210 905 55215 1175
rect 55185 890 55215 905
rect 55240 1175 55270 1185
rect 55240 905 55245 1175
rect 55265 905 55270 1175
rect 55180 885 55220 890
rect 55180 855 55185 885
rect 55215 855 55220 885
rect 55180 850 55220 855
rect 55240 830 55270 905
rect 55295 1175 55325 1190
rect 55295 905 55300 1175
rect 55320 905 55325 1175
rect 55295 890 55325 905
rect 55350 1175 55380 1185
rect 55350 905 55355 1175
rect 55375 905 55380 1175
rect 55290 885 55330 890
rect 55290 855 55295 885
rect 55325 855 55330 885
rect 55290 850 55330 855
rect 55350 830 55380 905
rect 55405 1175 55435 1185
rect 55405 905 55410 1175
rect 55430 905 55435 1175
rect 55405 865 55435 905
rect 55405 845 55410 865
rect 55430 845 55435 865
rect 54795 825 54835 830
rect 54795 795 54800 825
rect 54830 795 54835 825
rect 54795 785 54835 795
rect 54795 755 54800 785
rect 54830 755 54835 785
rect 54795 745 54835 755
rect 54795 715 54800 745
rect 54830 715 54835 745
rect 54795 710 54835 715
rect 54905 825 54945 830
rect 54905 795 54910 825
rect 54940 795 54945 825
rect 54905 785 54945 795
rect 54905 755 54910 785
rect 54940 755 54945 785
rect 54905 745 54945 755
rect 54905 715 54910 745
rect 54940 715 54945 745
rect 54905 710 54945 715
rect 55015 825 55055 830
rect 55015 795 55020 825
rect 55050 795 55055 825
rect 55015 785 55055 795
rect 55015 755 55020 785
rect 55050 755 55055 785
rect 55015 745 55055 755
rect 55015 715 55020 745
rect 55050 715 55055 745
rect 55015 710 55055 715
rect 55125 825 55165 830
rect 55125 795 55130 825
rect 55160 795 55165 825
rect 55125 785 55165 795
rect 55125 755 55130 785
rect 55160 755 55165 785
rect 55125 745 55165 755
rect 55125 715 55130 745
rect 55160 715 55165 745
rect 55125 710 55165 715
rect 55235 825 55275 830
rect 55235 795 55240 825
rect 55270 795 55275 825
rect 55235 785 55275 795
rect 55235 755 55240 785
rect 55270 755 55275 785
rect 55235 745 55275 755
rect 55235 715 55240 745
rect 55270 715 55275 745
rect 55235 710 55275 715
rect 55345 825 55385 830
rect 55345 795 55350 825
rect 55380 795 55385 825
rect 55345 785 55385 795
rect 55345 755 55350 785
rect 55380 755 55385 785
rect 55345 745 55385 755
rect 55345 715 55350 745
rect 55380 715 55385 745
rect 55345 710 55385 715
rect 55405 695 55435 845
rect 55660 825 55780 1825
rect 55895 1735 55935 1740
rect 55895 1705 55900 1735
rect 55930 1705 55935 1735
rect 55895 1700 55935 1705
rect 55660 795 55665 825
rect 55695 795 55705 825
rect 55735 795 55745 825
rect 55775 795 55780 825
rect 55660 785 55780 795
rect 55660 755 55665 785
rect 55695 755 55705 785
rect 55735 755 55745 785
rect 55775 755 55780 785
rect 55660 745 55780 755
rect 55660 715 55665 745
rect 55695 715 55705 745
rect 55735 715 55745 745
rect 55775 715 55780 745
rect 55660 710 55780 715
rect 55795 1235 55875 1240
rect 55795 1205 55800 1235
rect 55830 1205 55840 1235
rect 55870 1205 55875 1235
rect 55795 1195 55875 1205
rect 55795 1165 55800 1195
rect 55830 1165 55840 1195
rect 55870 1165 55875 1195
rect 55795 1155 55875 1165
rect 55795 1125 55800 1155
rect 55830 1125 55840 1155
rect 55870 1125 55875 1155
rect 54740 690 54780 695
rect 54740 660 54745 690
rect 54775 660 54780 690
rect 54740 650 54780 660
rect 54740 620 54745 650
rect 54775 620 54780 650
rect 54740 610 54780 620
rect 54740 580 54745 610
rect 54775 580 54780 610
rect 54740 575 54780 580
rect 55400 690 55440 695
rect 55400 660 55405 690
rect 55435 660 55440 690
rect 55400 650 55440 660
rect 55400 620 55405 650
rect 55435 620 55440 650
rect 55400 610 55440 620
rect 55400 580 55405 610
rect 55435 580 55440 610
rect 55400 575 55440 580
rect 54380 555 54420 560
rect 54380 525 54385 555
rect 54415 525 54420 555
rect 54380 520 54420 525
rect 54515 510 54555 515
rect 54515 480 54520 510
rect 54550 480 54555 510
rect 54515 475 54555 480
rect 55100 510 55140 515
rect 55100 480 55105 510
rect 55135 480 55140 510
rect 55100 475 55140 480
rect 54105 280 54110 310
rect 54140 280 54150 310
rect 54180 280 54195 310
rect 54225 280 54235 310
rect 54265 280 54280 310
rect 54310 280 54320 310
rect 54350 280 54355 310
rect 54105 270 54355 280
rect 54105 240 54110 270
rect 54140 240 54150 270
rect 54180 240 54195 270
rect 54225 240 54235 270
rect 54265 240 54280 270
rect 54310 240 54320 270
rect 54350 240 54355 270
rect 54105 230 54355 240
rect 54105 200 54110 230
rect 54140 200 54150 230
rect 54180 200 54195 230
rect 54225 200 54235 230
rect 54265 200 54280 230
rect 54310 200 54320 230
rect 54350 200 54355 230
rect 54105 195 54355 200
rect 54525 180 54545 475
rect 54580 310 54620 315
rect 54580 280 54585 310
rect 54615 280 54620 310
rect 54580 270 54620 280
rect 54580 240 54585 270
rect 54615 240 54620 270
rect 54580 230 54620 240
rect 54580 200 54585 230
rect 54615 200 54620 230
rect 54580 195 54620 200
rect 54850 310 55290 315
rect 54850 280 54855 310
rect 54885 280 54895 310
rect 54925 280 54935 310
rect 54965 280 54975 310
rect 55005 280 55015 310
rect 55045 280 55055 310
rect 55085 280 55095 310
rect 55125 280 55135 310
rect 55165 280 55175 310
rect 55205 280 55215 310
rect 55245 280 55255 310
rect 55285 280 55290 310
rect 54850 270 55290 280
rect 54850 240 54855 270
rect 54885 240 54895 270
rect 54925 240 54935 270
rect 54965 240 54975 270
rect 55005 240 55015 270
rect 55045 240 55055 270
rect 55085 240 55095 270
rect 55125 240 55135 270
rect 55165 240 55175 270
rect 55205 240 55215 270
rect 55245 240 55255 270
rect 55285 240 55290 270
rect 54850 230 55290 240
rect 54850 200 54855 230
rect 54885 200 54895 230
rect 54925 200 54935 230
rect 54965 200 54975 230
rect 55005 200 55015 230
rect 55045 200 55055 230
rect 55085 200 55095 230
rect 55125 200 55135 230
rect 55165 200 55175 230
rect 55205 200 55215 230
rect 55245 200 55255 230
rect 55285 200 55290 230
rect 54850 195 55290 200
rect 54520 175 54555 180
rect 54520 135 54555 140
rect 54580 175 54615 195
rect 54580 135 54615 140
rect 54755 165 54785 175
rect 54755 -505 54760 165
rect 54780 -505 54785 165
rect 54755 -545 54785 -505
rect 54855 165 54885 195
rect 54855 -505 54860 165
rect 54880 -505 54885 165
rect 54855 -520 54885 -505
rect 54955 165 54985 175
rect 54955 -505 54960 165
rect 54980 -505 54985 165
rect 54755 -565 54760 -545
rect 54780 -565 54785 -545
rect 54850 -525 54890 -520
rect 54850 -555 54855 -525
rect 54885 -555 54890 -525
rect 54850 -560 54890 -555
rect 54755 -575 54785 -565
rect 54955 -575 54985 -505
rect 55055 165 55085 195
rect 55055 -505 55060 165
rect 55080 -505 55085 165
rect 55055 -520 55085 -505
rect 55155 165 55185 175
rect 55155 -505 55160 165
rect 55180 -505 55185 165
rect 55050 -525 55090 -520
rect 55050 -555 55055 -525
rect 55085 -555 55090 -525
rect 55050 -560 55090 -555
rect 55155 -575 55185 -505
rect 55255 165 55285 195
rect 55255 -505 55260 165
rect 55280 -505 55285 165
rect 55255 -520 55285 -505
rect 55355 165 55385 175
rect 55355 -505 55360 165
rect 55380 -505 55385 165
rect 55795 -95 55875 1125
rect 55795 -125 55800 -95
rect 55830 -125 55840 -95
rect 55870 -125 55875 -95
rect 55795 -135 55875 -125
rect 55795 -165 55800 -135
rect 55830 -165 55840 -135
rect 55870 -165 55875 -135
rect 55795 -175 55875 -165
rect 55795 -205 55800 -175
rect 55830 -205 55840 -175
rect 55870 -205 55875 -175
rect 55795 -210 55875 -205
rect 55905 -270 55925 1700
rect 55950 560 55970 2495
rect 56970 2480 56990 2615
rect 57017 2605 57047 2615
rect 57085 2640 57125 2645
rect 57085 2610 57090 2640
rect 57120 2610 57125 2640
rect 57085 2605 57125 2610
rect 57163 2635 57193 2645
rect 57163 2615 57168 2635
rect 57188 2615 57193 2635
rect 57210 2625 57215 2645
rect 57235 2625 57240 2645
rect 57210 2615 57240 2625
rect 57163 2605 57193 2615
rect 57020 2535 57040 2605
rect 57170 2585 57190 2605
rect 57160 2580 57200 2585
rect 57160 2550 57165 2580
rect 57195 2550 57200 2580
rect 57160 2545 57200 2550
rect 57015 2530 57055 2535
rect 57015 2500 57020 2530
rect 57050 2500 57055 2530
rect 57015 2495 57055 2500
rect 56850 2475 56890 2480
rect 56850 2445 56855 2475
rect 56885 2445 56890 2475
rect 56850 2440 56890 2445
rect 56960 2475 57000 2480
rect 56960 2445 56965 2475
rect 56995 2445 57000 2475
rect 56960 2440 57000 2445
rect 56860 2370 56880 2440
rect 57220 2425 57240 2615
rect 57820 2530 57860 2535
rect 57820 2500 57825 2530
rect 57855 2500 57860 2530
rect 57820 2495 57860 2500
rect 56935 2420 56975 2425
rect 56935 2390 56940 2420
rect 56970 2390 56975 2420
rect 56935 2385 56975 2390
rect 57210 2420 57250 2425
rect 57210 2390 57215 2420
rect 57245 2390 57250 2420
rect 57210 2385 57250 2390
rect 56945 2370 56965 2385
rect 56830 2365 56890 2370
rect 56830 2335 56855 2365
rect 56885 2335 56890 2365
rect 56830 2330 56890 2335
rect 56935 2360 56975 2370
rect 56935 2340 56945 2360
rect 56965 2340 56975 2360
rect 56935 2330 56975 2340
rect 56775 2300 56805 2310
rect 56085 2220 56675 2225
rect 56085 2190 56090 2220
rect 56120 2190 56145 2220
rect 56175 2190 56200 2220
rect 56230 2190 56255 2220
rect 56285 2190 56310 2220
rect 56340 2190 56365 2220
rect 56395 2190 56420 2220
rect 56450 2190 56475 2220
rect 56505 2190 56530 2220
rect 56560 2190 56585 2220
rect 56615 2190 56640 2220
rect 56670 2190 56675 2220
rect 56085 2180 56675 2190
rect 56085 2150 56090 2180
rect 56120 2150 56145 2180
rect 56175 2150 56200 2180
rect 56230 2150 56255 2180
rect 56285 2150 56310 2180
rect 56340 2150 56365 2180
rect 56395 2150 56420 2180
rect 56450 2150 56475 2180
rect 56505 2150 56530 2180
rect 56560 2150 56585 2180
rect 56615 2150 56640 2180
rect 56670 2150 56675 2180
rect 56085 2140 56675 2150
rect 56085 2110 56090 2140
rect 56120 2110 56145 2140
rect 56175 2110 56200 2140
rect 56230 2110 56255 2140
rect 56285 2110 56310 2140
rect 56340 2110 56365 2140
rect 56395 2110 56420 2140
rect 56450 2110 56475 2140
rect 56505 2110 56530 2140
rect 56560 2110 56585 2140
rect 56615 2110 56640 2140
rect 56670 2110 56675 2140
rect 56085 2105 56675 2110
rect 55995 1735 56025 1740
rect 55995 1700 56025 1705
rect 56085 1680 56125 2105
rect 56140 1725 56180 1730
rect 56140 1695 56145 1725
rect 56175 1695 56180 1725
rect 56140 1690 56180 1695
rect 56085 1650 56090 1680
rect 56120 1650 56125 1680
rect 56085 1645 56125 1650
rect 56030 1630 56065 1640
rect 56030 1510 56040 1630
rect 56060 1510 56065 1630
rect 56030 1500 56065 1510
rect 56035 1495 56065 1500
rect 56090 1630 56120 1645
rect 56090 1510 56095 1630
rect 56115 1510 56120 1630
rect 56035 1470 56065 1480
rect 56035 1450 56040 1470
rect 56060 1450 56065 1470
rect 56090 1450 56120 1510
rect 56145 1630 56175 1690
rect 56195 1680 56235 2105
rect 56250 1725 56290 1730
rect 56250 1695 56255 1725
rect 56285 1695 56290 1725
rect 56250 1690 56290 1695
rect 56195 1650 56200 1680
rect 56230 1650 56235 1680
rect 56195 1645 56235 1650
rect 56145 1510 56150 1630
rect 56170 1510 56175 1630
rect 56145 1495 56175 1510
rect 56200 1630 56230 1645
rect 56200 1510 56205 1630
rect 56225 1510 56230 1630
rect 56140 1490 56180 1495
rect 56140 1460 56145 1490
rect 56175 1460 56180 1490
rect 56140 1455 56180 1460
rect 56035 1395 56065 1450
rect 56085 1445 56125 1450
rect 56085 1415 56090 1445
rect 56120 1415 56125 1445
rect 56085 1410 56125 1415
rect 56030 1390 56070 1395
rect 56030 1360 56035 1390
rect 56065 1360 56070 1390
rect 56030 1350 56070 1360
rect 56030 1320 56035 1350
rect 56065 1320 56070 1350
rect 56030 1310 56070 1320
rect 56030 1280 56035 1310
rect 56065 1280 56070 1310
rect 56030 1275 56070 1280
rect 56145 1065 56175 1455
rect 56200 1450 56230 1510
rect 56255 1630 56285 1690
rect 56305 1680 56345 2105
rect 56360 1725 56400 1730
rect 56360 1695 56365 1725
rect 56395 1695 56400 1725
rect 56360 1690 56400 1695
rect 56305 1650 56310 1680
rect 56340 1650 56345 1680
rect 56305 1645 56345 1650
rect 56255 1510 56260 1630
rect 56280 1510 56285 1630
rect 56255 1495 56285 1510
rect 56310 1630 56340 1645
rect 56310 1510 56315 1630
rect 56335 1510 56340 1630
rect 56250 1490 56290 1495
rect 56250 1460 56255 1490
rect 56285 1460 56290 1490
rect 56250 1455 56290 1460
rect 56195 1445 56235 1450
rect 56195 1415 56200 1445
rect 56230 1415 56235 1445
rect 56195 1410 56235 1415
rect 56085 1055 56125 1060
rect 56040 1045 56070 1050
rect 56085 1025 56090 1055
rect 56120 1025 56125 1055
rect 56255 1065 56285 1455
rect 56310 1450 56340 1510
rect 56365 1630 56395 1690
rect 56415 1680 56455 2105
rect 56470 1725 56510 1730
rect 56470 1695 56475 1725
rect 56505 1695 56510 1725
rect 56470 1690 56510 1695
rect 56415 1650 56420 1680
rect 56450 1650 56455 1680
rect 56415 1645 56455 1650
rect 56365 1510 56370 1630
rect 56390 1510 56395 1630
rect 56365 1495 56395 1510
rect 56420 1630 56450 1645
rect 56420 1510 56425 1630
rect 56445 1510 56450 1630
rect 56360 1490 56400 1495
rect 56360 1460 56365 1490
rect 56395 1460 56400 1490
rect 56360 1455 56400 1460
rect 56305 1445 56345 1450
rect 56305 1415 56310 1445
rect 56340 1415 56345 1445
rect 56305 1410 56345 1415
rect 56145 1030 56175 1035
rect 56195 1055 56235 1060
rect 56085 1020 56125 1025
rect 56195 1025 56200 1055
rect 56230 1025 56235 1055
rect 56365 1065 56395 1455
rect 56420 1450 56450 1510
rect 56475 1630 56505 1690
rect 56525 1680 56565 2105
rect 56580 1725 56620 1730
rect 56580 1695 56585 1725
rect 56615 1695 56620 1725
rect 56580 1690 56620 1695
rect 56525 1650 56530 1680
rect 56560 1650 56565 1680
rect 56525 1645 56565 1650
rect 56475 1510 56480 1630
rect 56500 1510 56505 1630
rect 56475 1495 56505 1510
rect 56530 1630 56560 1645
rect 56530 1510 56535 1630
rect 56555 1510 56560 1630
rect 56470 1490 56510 1495
rect 56470 1460 56475 1490
rect 56505 1460 56510 1490
rect 56470 1455 56510 1460
rect 56415 1445 56455 1450
rect 56415 1415 56420 1445
rect 56450 1415 56455 1445
rect 56415 1410 56455 1415
rect 56255 1030 56285 1035
rect 56305 1055 56345 1060
rect 56195 1020 56235 1025
rect 56305 1025 56310 1055
rect 56340 1025 56345 1055
rect 56475 1065 56505 1455
rect 56530 1450 56560 1510
rect 56585 1630 56615 1690
rect 56635 1680 56675 2105
rect 56775 2080 56780 2300
rect 56800 2080 56805 2300
rect 56775 2050 56805 2080
rect 56830 2300 56860 2330
rect 56830 2080 56835 2300
rect 56855 2080 56860 2300
rect 56830 2070 56860 2080
rect 56885 2300 56915 2310
rect 56885 2080 56890 2300
rect 56910 2080 56915 2300
rect 56885 2050 56915 2080
rect 56940 2300 56970 2330
rect 56940 2080 56945 2300
rect 56965 2080 56970 2300
rect 56940 2070 56970 2080
rect 56995 2300 57025 2310
rect 56995 2080 57000 2300
rect 57020 2080 57025 2300
rect 56995 2050 57025 2080
rect 57125 2220 57715 2225
rect 57125 2190 57130 2220
rect 57160 2190 57185 2220
rect 57215 2190 57240 2220
rect 57270 2190 57295 2220
rect 57325 2190 57350 2220
rect 57380 2190 57405 2220
rect 57435 2190 57460 2220
rect 57490 2190 57515 2220
rect 57545 2190 57570 2220
rect 57600 2190 57625 2220
rect 57655 2190 57680 2220
rect 57710 2190 57715 2220
rect 57125 2180 57715 2190
rect 57125 2150 57130 2180
rect 57160 2150 57185 2180
rect 57215 2150 57240 2180
rect 57270 2150 57295 2180
rect 57325 2150 57350 2180
rect 57380 2150 57405 2180
rect 57435 2150 57460 2180
rect 57490 2150 57515 2180
rect 57545 2150 57570 2180
rect 57600 2150 57625 2180
rect 57655 2150 57680 2180
rect 57710 2150 57715 2180
rect 57125 2140 57715 2150
rect 57125 2110 57130 2140
rect 57160 2110 57185 2140
rect 57215 2110 57240 2140
rect 57270 2110 57295 2140
rect 57325 2110 57350 2140
rect 57380 2110 57405 2140
rect 57435 2110 57460 2140
rect 57490 2110 57515 2140
rect 57545 2110 57570 2140
rect 57600 2110 57625 2140
rect 57655 2110 57680 2140
rect 57710 2110 57715 2140
rect 57125 2105 57715 2110
rect 56770 2045 56810 2050
rect 56770 2015 56775 2045
rect 56805 2015 56810 2045
rect 56770 2005 56810 2015
rect 56770 1975 56775 2005
rect 56805 1975 56810 2005
rect 56770 1965 56810 1975
rect 56770 1935 56775 1965
rect 56805 1935 56810 1965
rect 56770 1930 56810 1935
rect 56880 2045 56920 2050
rect 56880 2015 56885 2045
rect 56915 2015 56920 2045
rect 56880 2005 56920 2015
rect 56880 1975 56885 2005
rect 56915 1975 56920 2005
rect 56880 1965 56920 1975
rect 56880 1935 56885 1965
rect 56915 1935 56920 1965
rect 56880 1930 56920 1935
rect 56990 2045 57030 2050
rect 56990 2015 56995 2045
rect 57025 2015 57030 2045
rect 56990 2005 57030 2015
rect 56990 1975 56995 2005
rect 57025 1975 57030 2005
rect 56990 1965 57030 1975
rect 56990 1935 56995 1965
rect 57025 1935 57030 1965
rect 56990 1930 57030 1935
rect 56690 1735 56720 1740
rect 56690 1700 56720 1705
rect 57080 1735 57110 1740
rect 57080 1700 57110 1705
rect 56635 1650 56640 1680
rect 56670 1650 56675 1680
rect 56635 1645 56675 1650
rect 57125 1680 57165 2105
rect 57180 1725 57220 1730
rect 57180 1695 57185 1725
rect 57215 1695 57220 1725
rect 57180 1690 57220 1695
rect 57125 1650 57130 1680
rect 57160 1650 57165 1680
rect 57125 1645 57165 1650
rect 56585 1510 56590 1630
rect 56610 1510 56615 1630
rect 56585 1495 56615 1510
rect 56640 1630 56670 1645
rect 56640 1510 56645 1630
rect 56665 1510 56670 1630
rect 56580 1490 56620 1495
rect 56580 1460 56585 1490
rect 56615 1460 56620 1490
rect 56580 1455 56620 1460
rect 56525 1445 56565 1450
rect 56525 1415 56530 1445
rect 56560 1415 56565 1445
rect 56525 1410 56565 1415
rect 56365 1030 56395 1035
rect 56415 1055 56455 1060
rect 56305 1020 56345 1025
rect 56415 1025 56420 1055
rect 56450 1025 56455 1055
rect 56585 1065 56615 1455
rect 56640 1450 56670 1510
rect 56695 1630 56765 1640
rect 56695 1510 56700 1630
rect 56720 1510 56765 1630
rect 56695 1500 56765 1510
rect 57035 1630 57105 1640
rect 57035 1510 57080 1630
rect 57100 1510 57105 1630
rect 57035 1500 57105 1510
rect 56695 1470 56725 1500
rect 56695 1450 56700 1470
rect 56720 1450 56725 1470
rect 56635 1445 56675 1450
rect 56635 1415 56640 1445
rect 56670 1415 56675 1445
rect 56635 1410 56675 1415
rect 56695 1395 56725 1450
rect 57075 1470 57105 1500
rect 57075 1450 57080 1470
rect 57100 1450 57105 1470
rect 57130 1630 57160 1645
rect 57130 1510 57135 1630
rect 57155 1510 57160 1630
rect 57130 1450 57160 1510
rect 57185 1630 57215 1690
rect 57235 1680 57275 2105
rect 57290 1725 57330 1730
rect 57290 1695 57295 1725
rect 57325 1695 57330 1725
rect 57290 1690 57330 1695
rect 57235 1650 57240 1680
rect 57270 1650 57275 1680
rect 57235 1645 57275 1650
rect 57185 1510 57190 1630
rect 57210 1510 57215 1630
rect 57185 1495 57215 1510
rect 57240 1630 57270 1645
rect 57240 1510 57245 1630
rect 57265 1510 57270 1630
rect 57180 1490 57220 1495
rect 57180 1460 57185 1490
rect 57215 1460 57220 1490
rect 57180 1455 57220 1460
rect 57075 1395 57105 1450
rect 57125 1445 57165 1450
rect 57125 1415 57130 1445
rect 57160 1415 57165 1445
rect 57125 1410 57165 1415
rect 56690 1390 56730 1395
rect 56690 1360 56695 1390
rect 56725 1360 56730 1390
rect 56690 1350 56730 1360
rect 56690 1320 56695 1350
rect 56725 1320 56730 1350
rect 56690 1310 56730 1320
rect 56690 1280 56695 1310
rect 56725 1280 56730 1310
rect 56690 1275 56730 1280
rect 57070 1390 57110 1395
rect 57070 1360 57075 1390
rect 57105 1360 57110 1390
rect 57070 1350 57110 1360
rect 57070 1320 57075 1350
rect 57105 1320 57110 1350
rect 57070 1310 57110 1320
rect 57070 1280 57075 1310
rect 57105 1280 57110 1310
rect 57070 1275 57110 1280
rect 56880 1235 56920 1240
rect 56880 1205 56885 1235
rect 56915 1205 56920 1235
rect 56880 1195 56920 1205
rect 56880 1165 56885 1195
rect 56915 1165 56920 1195
rect 56880 1155 56920 1165
rect 56880 1125 56885 1155
rect 56915 1125 56920 1155
rect 56880 1120 56920 1125
rect 56475 1030 56505 1035
rect 56525 1055 56565 1060
rect 56415 1020 56455 1025
rect 56525 1025 56530 1055
rect 56560 1025 56565 1055
rect 56585 1030 56615 1035
rect 56635 1055 56675 1060
rect 56525 1020 56565 1025
rect 56635 1025 56640 1055
rect 56670 1025 56675 1055
rect 56635 1020 56675 1025
rect 56690 1055 56720 1060
rect 56690 1020 56720 1025
rect 56840 1055 56870 1060
rect 56840 1020 56870 1025
rect 56040 1010 56070 1015
rect 56035 955 56065 965
rect 56035 835 56040 955
rect 56060 835 56065 955
rect 56035 825 56065 835
rect 56090 955 56120 1020
rect 56140 1010 56180 1015
rect 56140 980 56145 1010
rect 56175 980 56180 1010
rect 56140 975 56180 980
rect 56090 835 56095 955
rect 56115 835 56120 955
rect 56090 820 56120 835
rect 56145 955 56175 975
rect 56145 835 56150 955
rect 56170 835 56175 955
rect 56085 815 56125 820
rect 56035 795 56065 805
rect 56035 775 56040 795
rect 56060 775 56065 795
rect 56085 785 56090 815
rect 56120 785 56125 815
rect 56085 780 56125 785
rect 56035 765 56065 775
rect 56040 695 56060 765
rect 56145 750 56175 835
rect 56200 955 56230 1020
rect 56250 1010 56290 1015
rect 56250 980 56255 1010
rect 56285 980 56290 1010
rect 56250 975 56290 980
rect 56200 835 56205 955
rect 56225 835 56230 955
rect 56200 820 56230 835
rect 56255 955 56285 975
rect 56255 835 56260 955
rect 56280 835 56285 955
rect 56195 815 56235 820
rect 56195 785 56200 815
rect 56230 785 56235 815
rect 56195 780 56235 785
rect 56255 750 56285 835
rect 56310 955 56340 1020
rect 56360 1010 56400 1015
rect 56360 980 56365 1010
rect 56395 980 56400 1010
rect 56360 975 56400 980
rect 56310 835 56315 955
rect 56335 835 56340 955
rect 56310 820 56340 835
rect 56365 955 56395 975
rect 56365 835 56370 955
rect 56390 835 56395 955
rect 56305 815 56345 820
rect 56305 785 56310 815
rect 56340 785 56345 815
rect 56305 780 56345 785
rect 56365 750 56395 835
rect 56420 955 56450 1020
rect 56470 1010 56510 1015
rect 56470 980 56475 1010
rect 56505 980 56510 1010
rect 56470 975 56510 980
rect 56420 835 56425 955
rect 56445 835 56450 955
rect 56420 820 56450 835
rect 56475 955 56505 975
rect 56475 835 56480 955
rect 56500 835 56505 955
rect 56415 815 56455 820
rect 56415 785 56420 815
rect 56450 785 56455 815
rect 56415 780 56455 785
rect 56475 750 56505 835
rect 56530 955 56560 1020
rect 56580 1010 56620 1015
rect 56580 980 56585 1010
rect 56615 980 56620 1010
rect 56580 975 56620 980
rect 56530 835 56535 955
rect 56555 835 56560 955
rect 56530 820 56560 835
rect 56585 955 56615 975
rect 56585 835 56590 955
rect 56610 835 56615 955
rect 56525 815 56565 820
rect 56525 785 56530 815
rect 56560 785 56565 815
rect 56525 780 56565 785
rect 56585 750 56615 835
rect 56640 955 56670 1020
rect 56640 835 56645 955
rect 56665 835 56670 955
rect 56640 820 56670 835
rect 56695 955 56805 965
rect 56695 835 56700 955
rect 56720 835 56780 955
rect 56800 835 56805 955
rect 56695 825 56805 835
rect 56830 955 56860 965
rect 56830 835 56835 955
rect 56855 835 56860 955
rect 56635 815 56675 820
rect 56635 785 56640 815
rect 56670 785 56675 815
rect 56740 805 56760 825
rect 56830 820 56860 835
rect 56885 955 56915 1120
rect 57185 1065 57215 1455
rect 57240 1450 57270 1510
rect 57295 1630 57325 1690
rect 57345 1680 57385 2105
rect 57400 1725 57440 1730
rect 57400 1695 57405 1725
rect 57435 1695 57440 1725
rect 57400 1690 57440 1695
rect 57345 1650 57350 1680
rect 57380 1650 57385 1680
rect 57345 1645 57385 1650
rect 57295 1510 57300 1630
rect 57320 1510 57325 1630
rect 57295 1495 57325 1510
rect 57350 1630 57380 1645
rect 57350 1510 57355 1630
rect 57375 1510 57380 1630
rect 57290 1490 57330 1495
rect 57290 1460 57295 1490
rect 57325 1460 57330 1490
rect 57290 1455 57330 1460
rect 57235 1445 57275 1450
rect 57235 1415 57240 1445
rect 57270 1415 57275 1445
rect 57235 1410 57275 1415
rect 56930 1055 56960 1060
rect 56930 1020 56960 1025
rect 57080 1055 57110 1060
rect 57080 1020 57110 1025
rect 57125 1055 57165 1060
rect 57125 1025 57130 1055
rect 57160 1025 57165 1055
rect 57295 1065 57325 1455
rect 57350 1450 57380 1510
rect 57405 1630 57435 1690
rect 57455 1680 57495 2105
rect 57510 1725 57550 1730
rect 57510 1695 57515 1725
rect 57545 1695 57550 1725
rect 57510 1690 57550 1695
rect 57455 1650 57460 1680
rect 57490 1650 57495 1680
rect 57455 1645 57495 1650
rect 57405 1510 57410 1630
rect 57430 1510 57435 1630
rect 57405 1495 57435 1510
rect 57460 1630 57490 1645
rect 57460 1510 57465 1630
rect 57485 1510 57490 1630
rect 57400 1490 57440 1495
rect 57400 1460 57405 1490
rect 57435 1460 57440 1490
rect 57400 1455 57440 1460
rect 57345 1445 57385 1450
rect 57345 1415 57350 1445
rect 57380 1415 57385 1445
rect 57345 1410 57385 1415
rect 57185 1030 57215 1035
rect 57235 1055 57275 1060
rect 57125 1020 57165 1025
rect 57235 1025 57240 1055
rect 57270 1025 57275 1055
rect 57405 1065 57435 1455
rect 57460 1450 57490 1510
rect 57515 1630 57545 1690
rect 57565 1680 57605 2105
rect 57620 1725 57660 1730
rect 57620 1695 57625 1725
rect 57655 1695 57660 1725
rect 57620 1690 57660 1695
rect 57565 1650 57570 1680
rect 57600 1650 57605 1680
rect 57565 1645 57605 1650
rect 57515 1510 57520 1630
rect 57540 1510 57545 1630
rect 57515 1495 57545 1510
rect 57570 1630 57600 1645
rect 57570 1510 57575 1630
rect 57595 1510 57600 1630
rect 57510 1490 57550 1495
rect 57510 1460 57515 1490
rect 57545 1460 57550 1490
rect 57510 1455 57550 1460
rect 57455 1445 57495 1450
rect 57455 1415 57460 1445
rect 57490 1415 57495 1445
rect 57455 1410 57495 1415
rect 57295 1030 57325 1035
rect 57345 1055 57385 1060
rect 57235 1020 57275 1025
rect 57345 1025 57350 1055
rect 57380 1025 57385 1055
rect 57515 1065 57545 1455
rect 57570 1450 57600 1510
rect 57625 1630 57655 1690
rect 57675 1680 57715 2105
rect 57675 1650 57680 1680
rect 57710 1650 57715 1680
rect 57675 1645 57715 1650
rect 57625 1510 57630 1630
rect 57650 1510 57655 1630
rect 57625 1495 57655 1510
rect 57680 1630 57710 1645
rect 57680 1510 57685 1630
rect 57705 1510 57710 1630
rect 57620 1490 57660 1495
rect 57620 1460 57625 1490
rect 57655 1460 57660 1490
rect 57620 1455 57660 1460
rect 57565 1445 57605 1450
rect 57565 1415 57570 1445
rect 57600 1415 57605 1445
rect 57565 1410 57605 1415
rect 57405 1030 57435 1035
rect 57455 1055 57495 1060
rect 57345 1020 57385 1025
rect 57455 1025 57460 1055
rect 57490 1025 57495 1055
rect 57625 1065 57655 1455
rect 57680 1450 57710 1510
rect 57735 1630 57765 1640
rect 57735 1510 57740 1630
rect 57760 1510 57765 1630
rect 57735 1500 57765 1510
rect 57735 1470 57765 1480
rect 57735 1450 57740 1470
rect 57760 1450 57765 1470
rect 57675 1445 57715 1450
rect 57675 1415 57680 1445
rect 57710 1415 57715 1445
rect 57675 1410 57715 1415
rect 57735 1395 57765 1450
rect 57730 1390 57770 1395
rect 57730 1360 57735 1390
rect 57765 1360 57770 1390
rect 57730 1350 57770 1360
rect 57730 1320 57735 1350
rect 57765 1320 57770 1350
rect 57730 1310 57770 1320
rect 57730 1280 57735 1310
rect 57765 1280 57770 1310
rect 57730 1275 57770 1280
rect 57515 1030 57545 1035
rect 57565 1055 57605 1060
rect 57455 1020 57495 1025
rect 57565 1025 57570 1055
rect 57600 1025 57605 1055
rect 57625 1030 57655 1035
rect 57675 1055 57715 1060
rect 57565 1020 57605 1025
rect 57675 1025 57680 1055
rect 57710 1025 57715 1055
rect 57675 1020 57715 1025
rect 57730 1045 57760 1050
rect 56885 835 56890 955
rect 56910 835 56915 955
rect 56885 825 56915 835
rect 56940 955 56970 965
rect 56940 835 56945 955
rect 56965 835 56970 955
rect 56940 820 56970 835
rect 56995 955 57105 965
rect 56995 835 57000 955
rect 57020 835 57080 955
rect 57100 835 57105 955
rect 56995 825 57105 835
rect 57130 955 57160 1020
rect 57180 1010 57220 1015
rect 57180 980 57185 1010
rect 57215 980 57220 1010
rect 57180 975 57220 980
rect 57130 835 57135 955
rect 57155 835 57160 955
rect 56825 815 56865 820
rect 56635 780 56675 785
rect 56735 795 56765 805
rect 56735 775 56740 795
rect 56760 775 56765 795
rect 56735 765 56765 775
rect 56825 785 56830 815
rect 56860 785 56865 815
rect 56140 745 56180 750
rect 56140 715 56145 745
rect 56175 715 56180 745
rect 56140 710 56180 715
rect 56250 745 56290 750
rect 56250 715 56255 745
rect 56285 715 56290 745
rect 56250 710 56290 715
rect 56360 745 56400 750
rect 56360 715 56365 745
rect 56395 715 56400 745
rect 56360 710 56400 715
rect 56440 745 56700 750
rect 56440 715 56475 745
rect 56505 715 56585 745
rect 56615 715 56700 745
rect 56030 690 56070 695
rect 56030 660 56035 690
rect 56065 660 56070 690
rect 56030 650 56070 660
rect 56030 620 56035 650
rect 56065 620 56070 650
rect 56030 610 56070 620
rect 56030 580 56035 610
rect 56065 580 56070 610
rect 56030 575 56070 580
rect 55940 555 55980 560
rect 55940 525 55945 555
rect 55975 525 55980 555
rect 55940 520 55980 525
rect 56440 390 56700 715
rect 56740 695 56760 765
rect 56730 690 56770 695
rect 56730 660 56735 690
rect 56765 660 56770 690
rect 56730 650 56770 660
rect 56730 620 56735 650
rect 56765 620 56770 650
rect 56730 610 56770 620
rect 56730 580 56735 610
rect 56765 580 56770 610
rect 56730 575 56770 580
rect 56440 360 56445 390
rect 56475 360 56555 390
rect 56585 360 56665 390
rect 56695 360 56700 390
rect 56440 355 56700 360
rect 56770 390 56810 395
rect 56770 360 56775 390
rect 56805 360 56810 390
rect 56770 355 56810 360
rect 56825 375 56865 785
rect 56935 815 56975 820
rect 56935 785 56940 815
rect 56970 785 56975 815
rect 57040 805 57060 825
rect 57130 820 57160 835
rect 57185 955 57215 975
rect 57185 835 57190 955
rect 57210 835 57215 955
rect 57125 815 57165 820
rect 56825 355 56835 375
rect 56855 355 56865 375
rect 56880 390 56920 395
rect 56880 360 56885 390
rect 56915 360 56920 390
rect 56880 355 56920 360
rect 56935 375 56975 785
rect 57035 795 57065 805
rect 57035 775 57040 795
rect 57060 775 57065 795
rect 57125 785 57130 815
rect 57160 785 57165 815
rect 57125 780 57165 785
rect 57035 765 57065 775
rect 57040 695 57060 765
rect 57185 750 57215 835
rect 57240 955 57270 1020
rect 57290 1010 57330 1015
rect 57290 980 57295 1010
rect 57325 980 57330 1010
rect 57290 975 57330 980
rect 57240 835 57245 955
rect 57265 835 57270 955
rect 57240 820 57270 835
rect 57295 955 57325 975
rect 57295 835 57300 955
rect 57320 835 57325 955
rect 57235 815 57275 820
rect 57235 785 57240 815
rect 57270 785 57275 815
rect 57235 780 57275 785
rect 57295 750 57325 835
rect 57350 955 57380 1020
rect 57400 1010 57440 1015
rect 57400 980 57405 1010
rect 57435 980 57440 1010
rect 57400 975 57440 980
rect 57350 835 57355 955
rect 57375 835 57380 955
rect 57350 820 57380 835
rect 57405 955 57435 975
rect 57405 835 57410 955
rect 57430 835 57435 955
rect 57345 815 57385 820
rect 57345 785 57350 815
rect 57380 785 57385 815
rect 57345 780 57385 785
rect 57405 750 57435 835
rect 57460 955 57490 1020
rect 57510 1010 57550 1015
rect 57510 980 57515 1010
rect 57545 980 57550 1010
rect 57510 975 57550 980
rect 57460 835 57465 955
rect 57485 835 57490 955
rect 57460 820 57490 835
rect 57515 955 57545 975
rect 57515 835 57520 955
rect 57540 835 57545 955
rect 57455 815 57495 820
rect 57455 785 57460 815
rect 57490 785 57495 815
rect 57455 780 57495 785
rect 57515 750 57545 835
rect 57570 955 57600 1020
rect 57620 1010 57660 1015
rect 57620 980 57625 1010
rect 57655 980 57660 1010
rect 57620 975 57660 980
rect 57570 835 57575 955
rect 57595 835 57600 955
rect 57570 820 57600 835
rect 57625 955 57655 975
rect 57625 835 57630 955
rect 57650 835 57655 955
rect 57565 815 57605 820
rect 57565 785 57570 815
rect 57600 785 57605 815
rect 57565 780 57605 785
rect 57625 750 57655 835
rect 57680 955 57710 1020
rect 57730 1010 57760 1015
rect 57680 835 57685 955
rect 57705 835 57710 955
rect 57680 820 57710 835
rect 57735 955 57765 965
rect 57735 835 57740 955
rect 57760 835 57765 955
rect 57735 825 57765 835
rect 57675 815 57715 820
rect 57675 785 57680 815
rect 57710 785 57715 815
rect 57675 780 57715 785
rect 57735 795 57765 805
rect 57735 775 57740 795
rect 57760 775 57765 795
rect 57735 765 57765 775
rect 57100 745 57360 750
rect 57100 715 57185 745
rect 57215 715 57295 745
rect 57325 715 57360 745
rect 57030 690 57070 695
rect 57030 660 57035 690
rect 57065 660 57070 690
rect 57030 650 57070 660
rect 57030 620 57035 650
rect 57065 620 57070 650
rect 57030 610 57070 620
rect 57030 580 57035 610
rect 57065 580 57070 610
rect 57030 575 57070 580
rect 56935 355 56945 375
rect 56965 355 56975 375
rect 56990 390 57030 395
rect 56990 360 56995 390
rect 57025 360 57030 390
rect 56990 355 57030 360
rect 57100 390 57360 715
rect 57400 745 57440 750
rect 57400 715 57405 745
rect 57435 715 57440 745
rect 57400 710 57440 715
rect 57510 745 57550 750
rect 57510 715 57515 745
rect 57545 715 57550 745
rect 57510 710 57550 715
rect 57620 745 57660 750
rect 57620 715 57625 745
rect 57655 715 57660 745
rect 57620 710 57660 715
rect 57740 695 57760 765
rect 57730 690 57770 695
rect 57730 660 57735 690
rect 57765 660 57770 690
rect 57730 650 57770 660
rect 57730 620 57735 650
rect 57765 620 57770 650
rect 57730 610 57770 620
rect 57730 580 57735 610
rect 57765 580 57770 610
rect 57730 575 57770 580
rect 57830 560 57850 2495
rect 57865 2420 57905 2425
rect 57865 2390 57870 2420
rect 57900 2390 57905 2420
rect 57865 2385 57905 2390
rect 57820 555 57860 560
rect 57820 525 57825 555
rect 57855 525 57860 555
rect 57820 520 57860 525
rect 57100 360 57105 390
rect 57135 360 57215 390
rect 57245 360 57325 390
rect 57355 360 57360 390
rect 57100 355 57360 360
rect 57430 390 57470 395
rect 57430 360 57435 390
rect 57465 360 57470 390
rect 57430 355 57470 360
rect 56185 315 56255 325
rect 56185 95 56230 315
rect 56250 95 56255 315
rect 56185 85 56255 95
rect 56225 65 56255 85
rect 56280 315 56310 325
rect 56280 95 56285 315
rect 56305 95 56310 315
rect 56280 65 56310 95
rect 56335 315 56365 325
rect 56335 95 56340 315
rect 56360 95 56365 315
rect 56220 60 56260 65
rect 56220 30 56225 60
rect 56255 30 56260 60
rect 55895 -275 55935 -270
rect 55895 -305 55900 -275
rect 55930 -305 55935 -275
rect 55895 -310 55935 -305
rect 55250 -525 55290 -520
rect 55250 -555 55255 -525
rect 55285 -555 55290 -525
rect 55250 -560 55290 -555
rect 55355 -545 55385 -505
rect 55355 -565 55360 -545
rect 55380 -565 55385 -545
rect 55355 -575 55385 -565
rect 56220 -575 56260 30
rect 56275 60 56315 65
rect 56275 30 56280 60
rect 56310 30 56315 60
rect 56275 25 56315 30
rect 56335 -90 56365 95
rect 56390 315 56420 325
rect 56390 95 56395 315
rect 56415 95 56420 315
rect 56390 65 56420 95
rect 56445 315 56475 355
rect 56445 95 56450 315
rect 56470 95 56475 315
rect 56385 60 56425 65
rect 56385 30 56390 60
rect 56420 30 56425 60
rect 56385 25 56425 30
rect 56445 20 56475 95
rect 56500 315 56530 325
rect 56500 95 56505 315
rect 56525 95 56530 315
rect 56500 65 56530 95
rect 56555 315 56585 355
rect 56555 95 56560 315
rect 56580 95 56585 315
rect 56495 60 56535 65
rect 56495 30 56500 60
rect 56530 30 56535 60
rect 56495 25 56535 30
rect 56555 20 56585 95
rect 56610 315 56640 325
rect 56610 95 56615 315
rect 56635 95 56640 315
rect 56610 65 56640 95
rect 56665 315 56695 355
rect 56665 95 56670 315
rect 56690 95 56695 315
rect 56605 60 56645 65
rect 56605 30 56610 60
rect 56640 30 56645 60
rect 56605 25 56645 30
rect 56665 20 56695 95
rect 56720 315 56750 325
rect 56720 95 56725 315
rect 56745 95 56750 315
rect 56720 65 56750 95
rect 56775 315 56805 355
rect 56825 345 56865 355
rect 56775 95 56780 315
rect 56800 95 56805 315
rect 56715 60 56755 65
rect 56715 30 56720 60
rect 56750 30 56755 60
rect 56715 25 56755 30
rect 56775 20 56805 95
rect 56830 315 56860 325
rect 56830 95 56835 315
rect 56855 95 56860 315
rect 56830 65 56860 95
rect 56885 315 56915 355
rect 56935 345 56975 355
rect 56885 95 56890 315
rect 56910 95 56915 315
rect 56825 60 56865 65
rect 56825 30 56830 60
rect 56860 30 56865 60
rect 56825 25 56865 30
rect 56885 20 56915 95
rect 56940 315 56970 325
rect 56940 95 56945 315
rect 56965 95 56970 315
rect 56940 65 56970 95
rect 56995 315 57025 355
rect 56995 95 57000 315
rect 57020 95 57025 315
rect 56935 60 56975 65
rect 56935 30 56940 60
rect 56970 30 56975 60
rect 56935 25 56975 30
rect 56995 20 57025 95
rect 57050 315 57080 325
rect 57050 95 57055 315
rect 57075 95 57080 315
rect 57050 65 57080 95
rect 57105 315 57135 355
rect 57105 95 57110 315
rect 57130 95 57135 315
rect 57045 60 57085 65
rect 57045 30 57050 60
rect 57080 30 57085 60
rect 57045 25 57085 30
rect 57105 20 57135 95
rect 57160 315 57190 325
rect 57160 95 57165 315
rect 57185 95 57190 315
rect 57160 65 57190 95
rect 57215 315 57245 355
rect 57215 95 57220 315
rect 57240 95 57245 315
rect 57155 60 57195 65
rect 57155 30 57160 60
rect 57190 30 57195 60
rect 57155 25 57195 30
rect 57215 20 57245 95
rect 57270 315 57300 325
rect 57270 95 57275 315
rect 57295 95 57300 315
rect 57270 65 57300 95
rect 57325 315 57355 355
rect 57325 95 57330 315
rect 57350 95 57355 315
rect 57265 60 57305 65
rect 57265 30 57270 60
rect 57300 30 57305 60
rect 57265 25 57305 30
rect 57325 20 57355 95
rect 57380 315 57410 325
rect 57380 95 57385 315
rect 57405 95 57410 315
rect 57380 65 57410 95
rect 57435 315 57465 355
rect 57435 95 57440 315
rect 57460 95 57465 315
rect 57375 60 57415 65
rect 57375 30 57380 60
rect 57410 30 57415 60
rect 57375 25 57415 30
rect 57435 20 57465 95
rect 57490 315 57520 325
rect 57490 95 57495 315
rect 57515 95 57520 315
rect 57490 65 57520 95
rect 57485 60 57525 65
rect 57485 30 57490 60
rect 57520 30 57525 60
rect 56440 15 56480 20
rect 56440 -15 56445 15
rect 56475 -15 56480 15
rect 56440 -20 56480 -15
rect 56550 15 56590 20
rect 56550 -15 56555 15
rect 56585 -15 56590 15
rect 56550 -20 56590 -15
rect 56660 15 56700 20
rect 56660 -15 56665 15
rect 56695 -15 56700 15
rect 56660 -20 56700 -15
rect 56770 15 56810 20
rect 56770 -15 56775 15
rect 56805 -15 56810 15
rect 56770 -20 56810 -15
rect 56880 15 56920 20
rect 56880 -15 56885 15
rect 56915 -15 56920 15
rect 56880 -20 56920 -15
rect 56990 15 57030 20
rect 56990 -15 56995 15
rect 57025 -15 57030 15
rect 56990 -20 57030 -15
rect 57100 15 57140 20
rect 57100 -15 57105 15
rect 57135 -15 57140 15
rect 57100 -20 57140 -15
rect 57210 15 57250 20
rect 57210 -15 57215 15
rect 57245 -15 57250 15
rect 57210 -20 57250 -15
rect 57320 15 57360 20
rect 57320 -15 57325 15
rect 57355 -15 57360 15
rect 57320 -20 57360 -15
rect 57430 15 57470 20
rect 57430 -15 57435 15
rect 57465 -15 57470 15
rect 57430 -20 57470 -15
rect 56330 -95 56370 -90
rect 56330 -125 56335 -95
rect 56365 -125 56370 -95
rect 56330 -135 56370 -125
rect 56330 -165 56335 -135
rect 56365 -165 56370 -135
rect 56330 -175 56370 -165
rect 56330 -205 56335 -175
rect 56365 -205 56370 -175
rect 56330 -210 56370 -205
rect 56540 -230 56580 -225
rect 56540 -260 56545 -230
rect 56575 -260 56580 -230
rect 56540 -265 56580 -260
rect 56650 -230 56690 -225
rect 56650 -260 56655 -230
rect 56685 -260 56690 -230
rect 56650 -265 56690 -260
rect 56870 -230 56910 -225
rect 56870 -260 56875 -230
rect 56905 -260 56910 -230
rect 56870 -265 56910 -260
rect 56485 -275 56525 -270
rect 56485 -305 56490 -275
rect 56520 -305 56525 -275
rect 56485 -310 56525 -305
rect 56395 -340 56465 -330
rect 56395 -460 56440 -340
rect 56460 -460 56465 -340
rect 56395 -470 56465 -460
rect 56435 -500 56465 -470
rect 56435 -520 56440 -500
rect 56460 -520 56465 -500
rect 56490 -340 56520 -310
rect 56490 -460 56495 -340
rect 56515 -460 56520 -340
rect 56490 -520 56520 -460
rect 56545 -340 56575 -265
rect 56595 -275 56635 -270
rect 56595 -305 56600 -275
rect 56630 -305 56635 -275
rect 56595 -310 56635 -305
rect 56545 -460 56550 -340
rect 56570 -460 56575 -340
rect 56545 -475 56575 -460
rect 56600 -340 56630 -310
rect 56600 -460 56605 -340
rect 56625 -460 56630 -340
rect 56540 -480 56580 -475
rect 56540 -510 56545 -480
rect 56575 -510 56580 -480
rect 56540 -515 56580 -510
rect 56600 -520 56630 -460
rect 56655 -340 56685 -265
rect 56705 -275 56745 -270
rect 56705 -305 56710 -275
rect 56740 -305 56745 -275
rect 56705 -310 56745 -305
rect 56655 -460 56660 -340
rect 56680 -460 56685 -340
rect 56655 -475 56685 -460
rect 56710 -340 56740 -310
rect 56710 -460 56715 -340
rect 56735 -460 56740 -340
rect 56650 -480 56690 -475
rect 56650 -510 56655 -480
rect 56685 -510 56690 -480
rect 56650 -515 56690 -510
rect 56710 -520 56740 -460
rect 56765 -340 56835 -330
rect 56765 -460 56770 -340
rect 56790 -460 56835 -340
rect 56765 -470 56835 -460
rect 56875 -340 56905 -265
rect 57040 -275 57080 -270
rect 57040 -305 57045 -275
rect 57075 -305 57080 -275
rect 57040 -310 57080 -305
rect 56875 -460 56880 -340
rect 56900 -460 56905 -340
rect 56765 -500 56795 -470
rect 56875 -475 56905 -460
rect 57215 -340 57245 -20
rect 57415 -40 57455 -35
rect 57415 -70 57420 -40
rect 57450 -70 57455 -40
rect 57415 -75 57455 -70
rect 57215 -460 57220 -340
rect 57240 -460 57245 -340
rect 57215 -470 57245 -460
rect 56765 -520 56770 -500
rect 56790 -520 56795 -500
rect 56870 -480 56910 -475
rect 56870 -510 56875 -480
rect 56905 -510 56910 -480
rect 56870 -515 56910 -510
rect 56435 -575 56465 -520
rect 56485 -525 56525 -520
rect 56485 -555 56490 -525
rect 56520 -555 56525 -525
rect 56485 -560 56525 -555
rect 56595 -525 56635 -520
rect 56595 -555 56600 -525
rect 56630 -555 56635 -525
rect 56595 -560 56635 -555
rect 56705 -525 56745 -520
rect 56705 -555 56710 -525
rect 56740 -555 56745 -525
rect 56705 -560 56745 -555
rect 56765 -575 56795 -520
rect 53960 -610 53965 -580
rect 53995 -610 54005 -580
rect 54035 -610 54045 -580
rect 54075 -610 54080 -580
rect 53960 -620 54080 -610
rect 53960 -650 53965 -620
rect 53995 -650 54005 -620
rect 54035 -650 54045 -620
rect 54075 -650 54080 -620
rect 53960 -660 54080 -650
rect 53960 -690 53965 -660
rect 53995 -690 54005 -660
rect 54035 -690 54045 -660
rect 54075 -690 54080 -660
rect 53960 -695 54080 -690
rect 54390 -580 54510 -575
rect 54390 -610 54395 -580
rect 54425 -610 54435 -580
rect 54465 -610 54475 -580
rect 54505 -610 54510 -580
rect 54390 -620 54510 -610
rect 54390 -650 54395 -620
rect 54425 -650 54435 -620
rect 54465 -650 54475 -620
rect 54505 -650 54510 -620
rect 54390 -660 54510 -650
rect 54390 -690 54395 -660
rect 54425 -690 54435 -660
rect 54465 -690 54475 -660
rect 54505 -690 54510 -660
rect 53690 -1500 53810 -695
rect 54040 -1500 54160 -695
rect 54390 -1500 54510 -690
rect 54740 -580 54860 -575
rect 54740 -610 54745 -580
rect 54775 -610 54785 -580
rect 54815 -610 54825 -580
rect 54855 -610 54860 -580
rect 54740 -620 54860 -610
rect 54740 -650 54745 -620
rect 54775 -650 54785 -620
rect 54815 -650 54825 -620
rect 54855 -650 54860 -620
rect 54740 -660 54860 -650
rect 54740 -690 54745 -660
rect 54775 -690 54785 -660
rect 54815 -690 54825 -660
rect 54855 -690 54860 -660
rect 54740 -1500 54860 -690
rect 55030 -580 55070 -575
rect 55030 -610 55035 -580
rect 55065 -610 55070 -580
rect 55030 -620 55070 -610
rect 55030 -650 55035 -620
rect 55065 -650 55070 -620
rect 55030 -660 55070 -650
rect 55030 -690 55035 -660
rect 55065 -690 55070 -660
rect 55030 -695 55070 -690
rect 55090 -580 55210 -575
rect 55090 -610 55095 -580
rect 55125 -610 55135 -580
rect 55165 -610 55175 -580
rect 55205 -610 55210 -580
rect 55090 -620 55210 -610
rect 55090 -650 55095 -620
rect 55125 -650 55135 -620
rect 55165 -650 55175 -620
rect 55205 -650 55210 -620
rect 55090 -660 55210 -650
rect 55090 -690 55095 -660
rect 55125 -690 55135 -660
rect 55165 -690 55175 -660
rect 55205 -690 55210 -660
rect 55090 -1500 55210 -690
rect 55230 -580 55270 -575
rect 55230 -610 55235 -580
rect 55265 -610 55270 -580
rect 55230 -620 55270 -610
rect 55230 -650 55235 -620
rect 55265 -650 55270 -620
rect 55230 -660 55270 -650
rect 55230 -690 55235 -660
rect 55265 -690 55270 -660
rect 55230 -695 55270 -690
rect 55440 -580 55560 -575
rect 55440 -610 55445 -580
rect 55475 -610 55485 -580
rect 55515 -610 55525 -580
rect 55555 -610 55560 -580
rect 55440 -620 55560 -610
rect 55440 -650 55445 -620
rect 55475 -650 55485 -620
rect 55515 -650 55525 -620
rect 55555 -650 55560 -620
rect 55440 -660 55560 -650
rect 55440 -690 55445 -660
rect 55475 -690 55485 -660
rect 55515 -690 55525 -660
rect 55555 -690 55560 -660
rect 55440 -1500 55560 -690
rect 55790 -580 55910 -575
rect 55790 -610 55795 -580
rect 55825 -610 55835 -580
rect 55865 -610 55875 -580
rect 55905 -610 55910 -580
rect 55790 -620 55910 -610
rect 55790 -650 55795 -620
rect 55825 -650 55835 -620
rect 55865 -650 55875 -620
rect 55905 -650 55910 -620
rect 55790 -660 55910 -650
rect 55790 -690 55795 -660
rect 55825 -690 55835 -660
rect 55865 -690 55875 -660
rect 55905 -690 55910 -660
rect 55790 -1500 55910 -690
rect 56140 -580 56260 -575
rect 56140 -610 56145 -580
rect 56175 -610 56185 -580
rect 56215 -610 56225 -580
rect 56255 -610 56260 -580
rect 56140 -620 56260 -610
rect 56140 -650 56145 -620
rect 56175 -650 56185 -620
rect 56215 -650 56225 -620
rect 56255 -650 56260 -620
rect 56140 -660 56260 -650
rect 56140 -690 56145 -660
rect 56175 -690 56185 -660
rect 56215 -690 56225 -660
rect 56255 -690 56260 -660
rect 56140 -1500 56260 -690
rect 56430 -580 56470 -575
rect 56430 -610 56435 -580
rect 56465 -610 56470 -580
rect 56430 -620 56470 -610
rect 56430 -650 56435 -620
rect 56465 -650 56470 -620
rect 56430 -660 56470 -650
rect 56430 -690 56435 -660
rect 56465 -690 56470 -660
rect 56430 -695 56470 -690
rect 56490 -580 56610 -575
rect 56490 -610 56495 -580
rect 56525 -610 56535 -580
rect 56565 -610 56575 -580
rect 56605 -610 56610 -580
rect 56490 -620 56610 -610
rect 56490 -650 56495 -620
rect 56525 -650 56535 -620
rect 56565 -650 56575 -620
rect 56605 -650 56610 -620
rect 56490 -660 56610 -650
rect 56490 -690 56495 -660
rect 56525 -690 56535 -660
rect 56565 -690 56575 -660
rect 56605 -690 56610 -660
rect 56490 -1500 56610 -690
rect 56760 -580 56800 -575
rect 56760 -610 56765 -580
rect 56795 -610 56800 -580
rect 56760 -620 56800 -610
rect 56760 -650 56765 -620
rect 56795 -650 56800 -620
rect 56760 -660 56800 -650
rect 56760 -690 56765 -660
rect 56795 -690 56800 -660
rect 56760 -695 56800 -690
rect 56840 -580 56960 -575
rect 56840 -610 56845 -580
rect 56875 -610 56885 -580
rect 56915 -610 56925 -580
rect 56955 -610 56960 -580
rect 56840 -620 56960 -610
rect 56840 -650 56845 -620
rect 56875 -650 56885 -620
rect 56915 -650 56925 -620
rect 56955 -650 56960 -620
rect 56840 -660 56960 -650
rect 56840 -690 56845 -660
rect 56875 -690 56885 -660
rect 56915 -690 56925 -660
rect 56955 -690 56960 -660
rect 56840 -1500 56960 -690
rect 57190 -580 57310 -575
rect 57190 -610 57195 -580
rect 57225 -610 57235 -580
rect 57265 -610 57275 -580
rect 57305 -610 57310 -580
rect 57190 -620 57310 -610
rect 57190 -650 57195 -620
rect 57225 -650 57235 -620
rect 57265 -650 57275 -620
rect 57305 -650 57310 -620
rect 57190 -660 57310 -650
rect 57190 -690 57195 -660
rect 57225 -690 57235 -660
rect 57265 -690 57275 -660
rect 57305 -690 57310 -660
rect 57190 -1500 57310 -690
rect 57485 -580 57525 30
rect 57875 -35 57895 2385
rect 57920 2045 58040 2050
rect 57920 2015 57925 2045
rect 57955 2015 57965 2045
rect 57995 2015 58005 2045
rect 58035 2015 58040 2045
rect 57920 2005 58040 2015
rect 57920 1975 57925 2005
rect 57955 1975 57965 2005
rect 57995 1975 58005 2005
rect 58035 1975 58040 2005
rect 57920 1965 58040 1975
rect 57920 1935 57925 1965
rect 57955 1935 57965 1965
rect 57995 1935 58005 1965
rect 58035 1935 58040 1965
rect 57920 1800 58040 1935
rect 57920 1770 57925 1800
rect 57955 1770 57965 1800
rect 57995 1770 58005 1800
rect 58035 1770 58040 1800
rect 57920 1760 58040 1770
rect 57920 1730 57925 1760
rect 57955 1730 57965 1760
rect 57995 1730 58005 1760
rect 58035 1730 58040 1760
rect 57920 1720 58040 1730
rect 57920 1690 57925 1720
rect 57955 1690 57965 1720
rect 57995 1690 58005 1720
rect 58035 1690 58040 1720
rect 57920 1390 58040 1690
rect 57920 1360 57925 1390
rect 57955 1360 57965 1390
rect 57995 1360 58005 1390
rect 58035 1360 58040 1390
rect 57920 1350 58040 1360
rect 57920 1320 57925 1350
rect 57955 1320 57965 1350
rect 57995 1320 58005 1350
rect 58035 1320 58040 1350
rect 57920 1310 58040 1320
rect 57920 1280 57925 1310
rect 57955 1280 57965 1310
rect 57995 1280 58005 1310
rect 58035 1280 58040 1310
rect 57920 1275 58040 1280
rect 58100 1935 58220 2995
rect 58100 1905 58105 1935
rect 58135 1905 58145 1935
rect 58175 1905 58185 1935
rect 58215 1905 58220 1935
rect 58100 1895 58220 1905
rect 58100 1865 58105 1895
rect 58135 1865 58145 1895
rect 58175 1865 58185 1895
rect 58215 1865 58220 1895
rect 58100 1855 58220 1865
rect 58100 1825 58105 1855
rect 58135 1825 58145 1855
rect 58175 1825 58185 1855
rect 58215 1825 58220 1855
rect 57920 1235 58040 1240
rect 57920 1205 57925 1235
rect 57955 1205 57965 1235
rect 57995 1205 58005 1235
rect 58035 1205 58040 1235
rect 57920 1195 58040 1205
rect 57920 1165 57925 1195
rect 57955 1165 57965 1195
rect 57995 1165 58005 1195
rect 58035 1165 58040 1195
rect 57920 1155 58040 1165
rect 57920 1125 57925 1155
rect 57955 1125 57965 1155
rect 57995 1125 58005 1155
rect 58035 1125 58040 1155
rect 57865 -40 57905 -35
rect 57865 -70 57870 -40
rect 57900 -70 57905 -40
rect 57865 -75 57905 -70
rect 57920 -95 58040 1125
rect 58100 830 58220 1825
rect 58240 3240 58360 3245
rect 58240 3210 58245 3240
rect 58275 3210 58285 3240
rect 58315 3210 58325 3240
rect 58355 3210 58360 3240
rect 58240 3200 58360 3210
rect 58240 3170 58245 3200
rect 58275 3170 58285 3200
rect 58315 3170 58325 3200
rect 58355 3170 58360 3200
rect 58240 3160 58360 3170
rect 58240 3130 58245 3160
rect 58275 3130 58285 3160
rect 58315 3130 58325 3160
rect 58355 3130 58360 3160
rect 58240 2220 58360 3130
rect 59855 3125 59895 3130
rect 58440 3105 58480 3110
rect 58440 3075 58445 3105
rect 58475 3075 58480 3105
rect 58440 3065 58480 3075
rect 58440 3035 58445 3065
rect 58475 3035 58480 3065
rect 58440 3025 58480 3035
rect 58440 2995 58445 3025
rect 58475 2995 58480 3025
rect 58440 2990 58480 2995
rect 58550 3105 58590 3110
rect 58550 3075 58555 3105
rect 58585 3075 58590 3105
rect 58550 3065 58590 3075
rect 58550 3035 58555 3065
rect 58585 3035 58590 3065
rect 58550 3025 58590 3035
rect 58550 2995 58555 3025
rect 58585 2995 58590 3025
rect 58550 2990 58590 2995
rect 58660 3105 58700 3110
rect 58660 3075 58665 3105
rect 58695 3075 58700 3105
rect 58660 3065 58700 3075
rect 58660 3035 58665 3065
rect 58695 3035 58700 3065
rect 58660 3025 58700 3035
rect 58660 2995 58665 3025
rect 58695 2995 58700 3025
rect 58660 2990 58700 2995
rect 58770 3105 58810 3110
rect 58770 3075 58775 3105
rect 58805 3075 58810 3105
rect 58770 3065 58810 3075
rect 58770 3035 58775 3065
rect 58805 3035 58810 3065
rect 58770 3025 58810 3035
rect 58770 2995 58775 3025
rect 58805 2995 58810 3025
rect 58770 2990 58810 2995
rect 58880 3105 58920 3110
rect 58880 3075 58885 3105
rect 58915 3075 58920 3105
rect 58880 3065 58920 3075
rect 58880 3035 58885 3065
rect 58915 3035 58920 3065
rect 58880 3025 58920 3035
rect 58880 2995 58885 3025
rect 58915 2995 58920 3025
rect 58880 2990 58920 2995
rect 58990 3105 59030 3110
rect 58990 3075 58995 3105
rect 59025 3075 59030 3105
rect 58990 3065 59030 3075
rect 58990 3035 58995 3065
rect 59025 3035 59030 3065
rect 58990 3025 59030 3035
rect 58990 2995 58995 3025
rect 59025 2995 59030 3025
rect 58990 2990 59030 2995
rect 59100 3105 59140 3110
rect 59100 3075 59105 3105
rect 59135 3075 59140 3105
rect 59855 3095 59860 3125
rect 59890 3095 59895 3125
rect 59855 3090 59895 3095
rect 59100 3065 59140 3075
rect 59100 3035 59105 3065
rect 59135 3035 59140 3065
rect 59100 3025 59140 3035
rect 59100 2995 59105 3025
rect 59135 2995 59140 3025
rect 59100 2990 59140 2995
rect 58445 2950 58475 2990
rect 58445 2930 58450 2950
rect 58470 2930 58475 2950
rect 58445 2890 58475 2930
rect 58495 2940 58535 2945
rect 58495 2910 58500 2940
rect 58530 2910 58535 2940
rect 58495 2905 58535 2910
rect 58445 2320 58450 2890
rect 58470 2320 58475 2890
rect 58445 2310 58475 2320
rect 58500 2890 58530 2905
rect 58500 2320 58505 2890
rect 58525 2320 58530 2890
rect 58500 2305 58530 2320
rect 58555 2890 58585 2990
rect 58605 2940 58645 2945
rect 58605 2910 58610 2940
rect 58640 2910 58645 2940
rect 58605 2905 58645 2910
rect 58555 2320 58560 2890
rect 58580 2320 58585 2890
rect 58555 2310 58585 2320
rect 58610 2890 58640 2905
rect 58610 2320 58615 2890
rect 58635 2320 58640 2890
rect 58610 2305 58640 2320
rect 58665 2890 58695 2990
rect 58715 2940 58755 2945
rect 58715 2910 58720 2940
rect 58750 2910 58755 2940
rect 58715 2905 58755 2910
rect 58665 2320 58670 2890
rect 58690 2320 58695 2890
rect 58665 2310 58695 2320
rect 58720 2890 58750 2905
rect 58720 2320 58725 2890
rect 58745 2320 58750 2890
rect 58720 2305 58750 2320
rect 58775 2890 58805 2990
rect 58825 2940 58865 2945
rect 58825 2910 58830 2940
rect 58860 2910 58865 2940
rect 58825 2905 58865 2910
rect 58775 2320 58780 2890
rect 58800 2320 58805 2890
rect 58775 2310 58805 2320
rect 58830 2890 58860 2905
rect 58830 2320 58835 2890
rect 58855 2320 58860 2890
rect 58830 2305 58860 2320
rect 58885 2890 58915 2990
rect 58935 2940 58975 2945
rect 58935 2910 58940 2940
rect 58970 2910 58975 2940
rect 58935 2905 58975 2910
rect 58885 2320 58890 2890
rect 58910 2320 58915 2890
rect 58885 2310 58915 2320
rect 58940 2890 58970 2905
rect 58940 2320 58945 2890
rect 58965 2320 58970 2890
rect 58940 2305 58970 2320
rect 58995 2890 59025 2990
rect 59105 2950 59135 2990
rect 59865 2965 59885 3090
rect 59045 2940 59085 2945
rect 59045 2910 59050 2940
rect 59080 2910 59085 2940
rect 59045 2905 59085 2910
rect 59105 2930 59110 2950
rect 59130 2930 59135 2950
rect 58995 2320 59000 2890
rect 59020 2320 59025 2890
rect 58995 2310 59025 2320
rect 59050 2890 59080 2905
rect 59050 2320 59055 2890
rect 59075 2320 59080 2890
rect 59050 2305 59080 2320
rect 59105 2890 59135 2930
rect 59805 2955 59946 2965
rect 59805 2935 59810 2955
rect 59830 2935 59865 2955
rect 59885 2935 59920 2955
rect 59940 2935 59946 2955
rect 59805 2925 59946 2935
rect 59105 2320 59110 2890
rect 59130 2320 59135 2890
rect 59805 2350 59946 2360
rect 59805 2330 59810 2350
rect 59830 2330 59865 2350
rect 59885 2330 59920 2350
rect 59940 2330 59946 2350
rect 59805 2320 59946 2330
rect 59105 2310 59135 2320
rect 58240 2190 58245 2220
rect 58275 2190 58285 2220
rect 58315 2190 58325 2220
rect 58355 2190 58360 2220
rect 58240 2180 58360 2190
rect 58240 2150 58245 2180
rect 58275 2150 58285 2180
rect 58315 2150 58325 2180
rect 58355 2150 58360 2180
rect 58240 2140 58360 2150
rect 58240 2110 58245 2140
rect 58275 2110 58285 2140
rect 58315 2110 58325 2140
rect 58355 2110 58360 2140
rect 58240 1345 58360 2110
rect 58495 2300 58535 2305
rect 58495 2270 58500 2300
rect 58530 2270 58535 2300
rect 58495 2075 58535 2270
rect 58605 2300 58645 2305
rect 58605 2270 58610 2300
rect 58640 2270 58645 2300
rect 58605 2075 58645 2270
rect 58715 2300 58755 2305
rect 58715 2270 58720 2300
rect 58750 2270 58755 2300
rect 58715 2075 58755 2270
rect 58825 2300 58865 2305
rect 58825 2270 58830 2300
rect 58860 2270 58865 2300
rect 58770 2220 58810 2225
rect 58770 2190 58775 2220
rect 58805 2190 58810 2220
rect 58770 2180 58810 2190
rect 58770 2150 58775 2180
rect 58805 2150 58810 2180
rect 58770 2140 58810 2150
rect 58770 2110 58775 2140
rect 58805 2110 58810 2140
rect 58770 2105 58810 2110
rect 58825 2075 58865 2270
rect 58935 2300 58975 2305
rect 58935 2270 58940 2300
rect 58970 2270 58975 2300
rect 58935 2075 58975 2270
rect 59045 2300 59085 2305
rect 59045 2270 59050 2300
rect 59080 2270 59085 2300
rect 59045 2075 59085 2270
rect 59815 2220 59935 2320
rect 59815 2190 59820 2220
rect 59850 2190 59860 2220
rect 59890 2190 59900 2220
rect 59930 2190 59935 2220
rect 59815 2180 59935 2190
rect 59815 2150 59820 2180
rect 59850 2150 59860 2180
rect 59890 2150 59900 2180
rect 59930 2150 59935 2180
rect 59815 2140 59935 2150
rect 59815 2110 59820 2140
rect 59850 2110 59860 2140
rect 59890 2110 59900 2140
rect 59930 2110 59935 2140
rect 59815 2105 59935 2110
rect 58495 2070 59085 2075
rect 58495 2040 58500 2070
rect 58530 2040 58555 2070
rect 58585 2040 58610 2070
rect 58640 2040 58665 2070
rect 58695 2040 58720 2070
rect 58750 2040 58775 2070
rect 58805 2040 58830 2070
rect 58860 2040 58885 2070
rect 58915 2040 58940 2070
rect 58970 2040 58995 2070
rect 59025 2040 59050 2070
rect 59080 2040 59085 2070
rect 58495 2030 59085 2040
rect 58495 2000 58500 2030
rect 58530 2000 58555 2030
rect 58585 2000 58610 2030
rect 58640 2000 58665 2030
rect 58695 2000 58720 2030
rect 58750 2000 58775 2030
rect 58805 2000 58830 2030
rect 58860 2000 58885 2030
rect 58915 2000 58940 2030
rect 58970 2000 58995 2030
rect 59025 2000 59050 2030
rect 59080 2000 59085 2030
rect 58495 1990 59085 2000
rect 58495 1960 58500 1990
rect 58530 1960 58555 1990
rect 58585 1960 58610 1990
rect 58640 1960 58665 1990
rect 58695 1960 58720 1990
rect 58750 1960 58775 1990
rect 58805 1960 58830 1990
rect 58860 1960 58885 1990
rect 58915 1960 58940 1990
rect 58970 1960 58995 1990
rect 59025 1960 59050 1990
rect 59080 1960 59085 1990
rect 58495 1955 59085 1960
rect 59715 2070 59965 2075
rect 59715 2040 59720 2070
rect 59750 2040 59760 2070
rect 59790 2040 59805 2070
rect 59835 2040 59845 2070
rect 59875 2040 59890 2070
rect 59920 2040 59930 2070
rect 59960 2040 59965 2070
rect 59715 2030 59965 2040
rect 59715 2000 59720 2030
rect 59750 2000 59760 2030
rect 59790 2000 59805 2030
rect 59835 2000 59845 2030
rect 59875 2000 59890 2030
rect 59920 2000 59930 2030
rect 59960 2000 59965 2030
rect 59715 1990 59965 2000
rect 59715 1960 59720 1990
rect 59750 1960 59760 1990
rect 59790 1960 59805 1990
rect 59835 1960 59845 1990
rect 59875 1960 59890 1990
rect 59920 1960 59930 1990
rect 59960 1960 59965 1990
rect 58440 1935 58480 1940
rect 58440 1905 58445 1935
rect 58475 1905 58480 1935
rect 58440 1895 58480 1905
rect 58440 1865 58445 1895
rect 58475 1865 58480 1895
rect 58440 1855 58480 1865
rect 58440 1825 58445 1855
rect 58475 1825 58480 1855
rect 58440 1820 58480 1825
rect 59100 1935 59140 1940
rect 59100 1905 59105 1935
rect 59135 1905 59140 1935
rect 59100 1895 59140 1905
rect 59100 1865 59105 1895
rect 59135 1865 59140 1895
rect 59100 1855 59140 1865
rect 59100 1825 59105 1855
rect 59135 1825 59140 1855
rect 59100 1820 59140 1825
rect 58445 1675 58475 1820
rect 58495 1800 58535 1805
rect 58495 1770 58500 1800
rect 58530 1770 58535 1800
rect 58495 1760 58535 1770
rect 58495 1730 58500 1760
rect 58530 1730 58535 1760
rect 58495 1720 58535 1730
rect 58495 1690 58500 1720
rect 58530 1690 58535 1720
rect 58495 1685 58535 1690
rect 58605 1800 58645 1805
rect 58605 1770 58610 1800
rect 58640 1770 58645 1800
rect 58605 1760 58645 1770
rect 58605 1730 58610 1760
rect 58640 1730 58645 1760
rect 58605 1720 58645 1730
rect 58605 1690 58610 1720
rect 58640 1690 58645 1720
rect 58605 1685 58645 1690
rect 58715 1800 58755 1805
rect 58715 1770 58720 1800
rect 58750 1770 58755 1800
rect 58715 1760 58755 1770
rect 58715 1730 58720 1760
rect 58750 1730 58755 1760
rect 58715 1720 58755 1730
rect 58715 1690 58720 1720
rect 58750 1690 58755 1720
rect 58715 1685 58755 1690
rect 58825 1800 58865 1805
rect 58825 1770 58830 1800
rect 58860 1770 58865 1800
rect 58825 1760 58865 1770
rect 58825 1730 58830 1760
rect 58860 1730 58865 1760
rect 58825 1720 58865 1730
rect 58825 1690 58830 1720
rect 58860 1690 58865 1720
rect 58825 1685 58865 1690
rect 58935 1800 58975 1805
rect 58935 1770 58940 1800
rect 58970 1770 58975 1800
rect 58935 1760 58975 1770
rect 58935 1730 58940 1760
rect 58970 1730 58975 1760
rect 58935 1720 58975 1730
rect 58935 1690 58940 1720
rect 58970 1690 58975 1720
rect 58935 1685 58975 1690
rect 59045 1800 59085 1805
rect 59045 1770 59050 1800
rect 59080 1770 59085 1800
rect 59045 1760 59085 1770
rect 59045 1730 59050 1760
rect 59080 1730 59085 1760
rect 59045 1720 59085 1730
rect 59045 1690 59050 1720
rect 59080 1690 59085 1720
rect 59045 1685 59085 1690
rect 58445 1655 58450 1675
rect 58470 1655 58475 1675
rect 58445 1615 58475 1655
rect 58445 1445 58450 1615
rect 58470 1445 58475 1615
rect 58445 1435 58475 1445
rect 58500 1615 58530 1685
rect 58550 1665 58590 1670
rect 58550 1635 58555 1665
rect 58585 1635 58590 1665
rect 58550 1630 58590 1635
rect 58500 1445 58505 1615
rect 58525 1445 58530 1615
rect 58500 1435 58530 1445
rect 58555 1615 58585 1630
rect 58555 1445 58560 1615
rect 58580 1445 58585 1615
rect 58555 1415 58585 1445
rect 58610 1615 58640 1685
rect 58660 1665 58700 1670
rect 58660 1635 58665 1665
rect 58695 1635 58700 1665
rect 58660 1630 58700 1635
rect 58610 1445 58615 1615
rect 58635 1445 58640 1615
rect 58610 1435 58640 1445
rect 58665 1615 58695 1630
rect 58665 1445 58670 1615
rect 58690 1445 58695 1615
rect 58665 1415 58695 1445
rect 58720 1615 58750 1685
rect 58770 1665 58810 1670
rect 58770 1635 58775 1665
rect 58805 1635 58810 1665
rect 58770 1630 58810 1635
rect 58720 1445 58725 1615
rect 58745 1445 58750 1615
rect 58720 1435 58750 1445
rect 58775 1615 58805 1630
rect 58775 1445 58780 1615
rect 58800 1445 58805 1615
rect 58775 1415 58805 1445
rect 58830 1615 58860 1685
rect 58880 1665 58920 1670
rect 58880 1635 58885 1665
rect 58915 1635 58920 1665
rect 58880 1630 58920 1635
rect 58830 1445 58835 1615
rect 58855 1445 58860 1615
rect 58830 1435 58860 1445
rect 58885 1615 58915 1630
rect 58885 1445 58890 1615
rect 58910 1445 58915 1615
rect 58885 1415 58915 1445
rect 58940 1615 58970 1685
rect 58990 1665 59030 1670
rect 58990 1635 58995 1665
rect 59025 1635 59030 1665
rect 58990 1630 59030 1635
rect 58940 1445 58945 1615
rect 58965 1445 58970 1615
rect 58940 1435 58970 1445
rect 58995 1615 59025 1630
rect 58995 1445 59000 1615
rect 59020 1445 59025 1615
rect 58995 1415 59025 1445
rect 59050 1615 59080 1685
rect 59050 1445 59055 1615
rect 59075 1445 59080 1615
rect 59050 1435 59080 1445
rect 59105 1675 59135 1820
rect 59105 1655 59110 1675
rect 59130 1655 59135 1675
rect 59105 1615 59135 1655
rect 59105 1445 59110 1615
rect 59130 1445 59135 1615
rect 59105 1435 59135 1445
rect 59715 1435 59965 1960
rect 58550 1410 58590 1415
rect 58550 1380 58555 1410
rect 58585 1380 58590 1410
rect 58550 1375 58590 1380
rect 58660 1410 58700 1415
rect 58660 1380 58665 1410
rect 58695 1380 58700 1410
rect 58660 1375 58700 1380
rect 58770 1410 58810 1415
rect 58770 1380 58775 1410
rect 58805 1380 58810 1410
rect 58770 1375 58810 1380
rect 58880 1410 58920 1415
rect 58880 1380 58885 1410
rect 58915 1380 58920 1410
rect 58880 1375 58920 1380
rect 58990 1410 59030 1415
rect 58990 1380 58995 1410
rect 59025 1380 59030 1410
rect 58990 1375 59030 1380
rect 59430 1410 59470 1415
rect 59430 1380 59435 1410
rect 59465 1380 59470 1410
rect 59430 1375 59470 1380
rect 59715 1405 59725 1435
rect 59755 1405 59775 1435
rect 59805 1405 59825 1435
rect 59855 1405 59875 1435
rect 59905 1405 59925 1435
rect 59955 1405 59965 1435
rect 59715 1385 59965 1405
rect 58240 1315 58245 1345
rect 58275 1315 58285 1345
rect 58315 1315 58325 1345
rect 58355 1315 58360 1345
rect 58240 1305 58360 1315
rect 58240 1275 58245 1305
rect 58275 1275 58285 1305
rect 58315 1275 58325 1305
rect 58355 1275 58360 1305
rect 58240 1270 58360 1275
rect 58605 1345 58645 1350
rect 58605 1315 58610 1345
rect 58640 1315 58645 1345
rect 58605 1305 58645 1315
rect 58605 1275 58610 1305
rect 58640 1275 58645 1305
rect 58605 1270 58645 1275
rect 58550 1225 58590 1230
rect 58550 1195 58555 1225
rect 58585 1195 58590 1225
rect 58550 1190 58590 1195
rect 58660 1225 58700 1230
rect 58660 1195 58665 1225
rect 58695 1195 58700 1225
rect 58660 1190 58700 1195
rect 58770 1225 58810 1230
rect 58770 1195 58775 1225
rect 58805 1195 58810 1225
rect 58770 1190 58810 1195
rect 58880 1225 58920 1230
rect 58880 1195 58885 1225
rect 58915 1195 58920 1225
rect 58880 1190 58920 1195
rect 58990 1225 59030 1230
rect 58990 1195 58995 1225
rect 59025 1195 59030 1225
rect 58990 1190 59030 1195
rect 59195 1225 59235 1230
rect 59195 1195 59200 1225
rect 59230 1195 59235 1225
rect 59195 1190 59235 1195
rect 58100 800 58105 830
rect 58135 800 58145 830
rect 58175 800 58185 830
rect 58215 800 58220 830
rect 58100 790 58220 800
rect 58100 760 58105 790
rect 58135 760 58145 790
rect 58175 760 58185 790
rect 58215 760 58220 790
rect 58100 750 58220 760
rect 58100 720 58105 750
rect 58135 720 58145 750
rect 58175 720 58185 750
rect 58215 720 58220 750
rect 58100 715 58220 720
rect 58445 1175 58475 1185
rect 58445 905 58450 1175
rect 58470 905 58475 1175
rect 58445 865 58475 905
rect 58445 845 58450 865
rect 58470 845 58475 865
rect 58445 695 58475 845
rect 58500 1175 58530 1185
rect 58500 905 58505 1175
rect 58525 905 58530 1175
rect 58500 835 58530 905
rect 58555 1175 58585 1190
rect 58555 905 58560 1175
rect 58580 905 58585 1175
rect 58555 890 58585 905
rect 58610 1175 58640 1185
rect 58610 905 58615 1175
rect 58635 905 58640 1175
rect 58550 885 58590 890
rect 58550 855 58555 885
rect 58585 855 58590 885
rect 58550 850 58590 855
rect 58610 835 58640 905
rect 58665 1175 58695 1190
rect 58665 905 58670 1175
rect 58690 905 58695 1175
rect 58665 890 58695 905
rect 58720 1175 58750 1185
rect 58720 905 58725 1175
rect 58745 905 58750 1175
rect 58660 885 58700 890
rect 58660 855 58665 885
rect 58695 855 58700 885
rect 58660 850 58700 855
rect 58720 835 58750 905
rect 58775 1175 58805 1190
rect 58775 905 58780 1175
rect 58800 905 58805 1175
rect 58775 890 58805 905
rect 58830 1175 58860 1185
rect 58830 905 58835 1175
rect 58855 905 58860 1175
rect 58770 885 58810 890
rect 58770 855 58775 885
rect 58805 855 58810 885
rect 58770 850 58810 855
rect 58830 835 58860 905
rect 58885 1175 58915 1190
rect 58885 905 58890 1175
rect 58910 905 58915 1175
rect 58885 890 58915 905
rect 58940 1175 58970 1185
rect 58940 905 58945 1175
rect 58965 905 58970 1175
rect 58880 885 58920 890
rect 58880 855 58885 885
rect 58915 855 58920 885
rect 58880 850 58920 855
rect 58940 835 58970 905
rect 58995 1175 59025 1190
rect 58995 905 59000 1175
rect 59020 905 59025 1175
rect 58995 890 59025 905
rect 59050 1175 59080 1185
rect 59050 905 59055 1175
rect 59075 905 59080 1175
rect 58990 885 59030 890
rect 58990 855 58995 885
rect 59025 855 59030 885
rect 58990 850 59030 855
rect 59050 835 59080 905
rect 59105 1175 59135 1185
rect 59105 905 59110 1175
rect 59130 905 59135 1175
rect 59205 910 59225 1190
rect 59105 865 59135 905
rect 59195 905 59235 910
rect 59195 875 59200 905
rect 59230 875 59235 905
rect 59195 870 59235 875
rect 59105 845 59110 865
rect 59130 845 59135 865
rect 58495 830 58535 835
rect 58495 800 58500 830
rect 58530 800 58535 830
rect 58495 790 58535 800
rect 58495 760 58500 790
rect 58530 760 58535 790
rect 58495 750 58535 760
rect 58495 720 58500 750
rect 58530 720 58535 750
rect 58495 715 58535 720
rect 58605 830 58645 835
rect 58605 800 58610 830
rect 58640 800 58645 830
rect 58605 790 58645 800
rect 58605 760 58610 790
rect 58640 760 58645 790
rect 58605 750 58645 760
rect 58605 720 58610 750
rect 58640 720 58645 750
rect 58605 715 58645 720
rect 58715 830 58755 835
rect 58715 800 58720 830
rect 58750 800 58755 830
rect 58715 790 58755 800
rect 58715 760 58720 790
rect 58750 760 58755 790
rect 58715 750 58755 760
rect 58715 720 58720 750
rect 58750 720 58755 750
rect 58715 715 58755 720
rect 58825 830 58865 835
rect 58825 800 58830 830
rect 58860 800 58865 830
rect 58825 790 58865 800
rect 58825 760 58830 790
rect 58860 760 58865 790
rect 58825 750 58865 760
rect 58825 720 58830 750
rect 58860 720 58865 750
rect 58825 715 58865 720
rect 58935 830 58975 835
rect 58935 800 58940 830
rect 58970 800 58975 830
rect 58935 790 58975 800
rect 58935 760 58940 790
rect 58970 760 58975 790
rect 58935 750 58975 760
rect 58935 720 58940 750
rect 58970 720 58975 750
rect 58935 715 58975 720
rect 59045 830 59085 835
rect 59045 800 59050 830
rect 59080 800 59085 830
rect 59045 790 59085 800
rect 59045 760 59050 790
rect 59080 760 59085 790
rect 59045 750 59085 760
rect 59045 720 59050 750
rect 59080 720 59085 750
rect 59045 715 59085 720
rect 59105 695 59135 845
rect 59440 840 59460 1375
rect 59715 1355 59725 1385
rect 59755 1355 59775 1385
rect 59805 1355 59825 1385
rect 59855 1355 59875 1385
rect 59905 1355 59925 1385
rect 59955 1355 59965 1385
rect 59715 1335 59965 1355
rect 59715 1305 59725 1335
rect 59755 1305 59775 1335
rect 59805 1305 59825 1335
rect 59855 1305 59875 1335
rect 59905 1305 59925 1335
rect 59955 1305 59965 1335
rect 59475 910 59510 915
rect 59475 870 59510 875
rect 59535 910 59570 915
rect 59535 870 59570 875
rect 59595 910 59630 915
rect 59595 870 59630 875
rect 59655 910 59690 916
rect 59655 870 59690 875
rect 59540 840 59560 870
rect 59430 835 59470 840
rect 59430 805 59435 835
rect 59465 805 59470 835
rect 59430 800 59470 805
rect 59530 835 59570 840
rect 59530 805 59535 835
rect 59565 805 59570 835
rect 59530 800 59570 805
rect 58440 690 58480 695
rect 58440 660 58445 690
rect 58475 660 58480 690
rect 58440 650 58480 660
rect 58440 620 58445 650
rect 58475 620 58480 650
rect 58440 610 58480 620
rect 58440 580 58445 610
rect 58475 580 58480 610
rect 58440 575 58480 580
rect 59100 690 59140 695
rect 59100 660 59105 690
rect 59135 660 59140 690
rect 59100 650 59140 660
rect 59100 620 59105 650
rect 59135 620 59140 650
rect 59100 610 59140 620
rect 59100 580 59105 610
rect 59135 580 59140 610
rect 59100 575 59140 580
rect 59660 560 59680 870
rect 59650 555 59690 560
rect 59650 525 59655 555
rect 59685 525 59690 555
rect 59650 520 59690 525
rect 58580 510 58620 515
rect 58580 480 58585 510
rect 58615 480 58620 510
rect 58580 475 58620 480
rect 59515 510 59555 515
rect 59515 480 59520 510
rect 59550 480 59555 510
rect 59515 475 59555 480
rect 58430 310 58870 315
rect 58430 280 58435 310
rect 58465 280 58475 310
rect 58505 280 58515 310
rect 58545 280 58555 310
rect 58585 280 58595 310
rect 58625 280 58635 310
rect 58665 280 58675 310
rect 58705 280 58715 310
rect 58745 280 58755 310
rect 58785 280 58795 310
rect 58825 280 58835 310
rect 58865 280 58870 310
rect 58430 270 58870 280
rect 58430 240 58435 270
rect 58465 240 58475 270
rect 58505 240 58515 270
rect 58545 240 58555 270
rect 58585 240 58595 270
rect 58625 240 58635 270
rect 58665 240 58675 270
rect 58705 240 58715 270
rect 58745 240 58755 270
rect 58785 240 58795 270
rect 58825 240 58835 270
rect 58865 240 58870 270
rect 58430 230 58870 240
rect 58430 200 58435 230
rect 58465 200 58475 230
rect 58505 200 58515 230
rect 58545 200 58555 230
rect 58585 200 58595 230
rect 58625 200 58635 230
rect 58665 200 58675 230
rect 58705 200 58715 230
rect 58745 200 58755 230
rect 58785 200 58795 230
rect 58825 200 58835 230
rect 58865 200 58870 230
rect 58430 195 58870 200
rect 59450 310 59490 315
rect 59450 280 59455 310
rect 59485 280 59490 310
rect 59450 270 59490 280
rect 59450 240 59455 270
rect 59485 240 59490 270
rect 59450 230 59490 240
rect 59450 200 59455 230
rect 59485 200 59490 230
rect 59450 195 59490 200
rect 57920 -125 57925 -95
rect 57955 -125 57965 -95
rect 57995 -125 58005 -95
rect 58035 -125 58040 -95
rect 57920 -135 58040 -125
rect 57920 -165 57925 -135
rect 57955 -165 57965 -135
rect 57995 -165 58005 -135
rect 58035 -165 58040 -135
rect 57920 -175 58040 -165
rect 57920 -205 57925 -175
rect 57955 -205 57965 -175
rect 57995 -205 58005 -175
rect 58035 -205 58040 -175
rect 57920 -210 58040 -205
rect 58335 165 58365 175
rect 58335 -505 58340 165
rect 58360 -505 58365 165
rect 58335 -545 58365 -505
rect 58435 165 58465 195
rect 58435 -505 58440 165
rect 58460 -505 58465 165
rect 58435 -520 58465 -505
rect 58535 165 58565 175
rect 58535 -505 58540 165
rect 58560 -505 58565 165
rect 58335 -565 58340 -545
rect 58360 -565 58365 -545
rect 58430 -525 58470 -520
rect 58430 -555 58435 -525
rect 58465 -555 58470 -525
rect 58430 -560 58470 -555
rect 58335 -575 58365 -565
rect 58535 -575 58565 -505
rect 58635 165 58665 195
rect 58635 -505 58640 165
rect 58660 -505 58665 165
rect 58635 -520 58665 -505
rect 58735 165 58765 175
rect 58735 -505 58740 165
rect 58760 -505 58765 165
rect 58630 -525 58670 -520
rect 58630 -555 58635 -525
rect 58665 -555 58670 -525
rect 58630 -560 58670 -555
rect 58735 -575 58765 -505
rect 58835 165 58865 195
rect 59455 175 59490 195
rect 59525 180 59545 475
rect 59715 310 59965 1305
rect 59715 280 59720 310
rect 59750 280 59760 310
rect 59790 280 59805 310
rect 59835 280 59845 310
rect 59875 280 59890 310
rect 59920 280 59930 310
rect 59960 280 59965 310
rect 59715 270 59965 280
rect 59715 240 59720 270
rect 59750 240 59760 270
rect 59790 240 59805 270
rect 59835 240 59845 270
rect 59875 240 59890 270
rect 59920 240 59930 270
rect 59960 240 59965 270
rect 59715 230 59965 240
rect 59715 200 59720 230
rect 59750 200 59760 230
rect 59790 200 59805 230
rect 59835 200 59845 230
rect 59875 200 59890 230
rect 59920 200 59930 230
rect 59960 200 59965 230
rect 59715 195 59965 200
rect 59990 1800 60110 1805
rect 59990 1770 59995 1800
rect 60025 1770 60035 1800
rect 60065 1770 60075 1800
rect 60105 1770 60110 1800
rect 59990 1760 60110 1770
rect 59990 1730 59995 1760
rect 60025 1730 60035 1760
rect 60065 1730 60075 1760
rect 60105 1730 60110 1760
rect 59990 1720 60110 1730
rect 59990 1690 59995 1720
rect 60025 1690 60035 1720
rect 60065 1690 60075 1720
rect 60105 1690 60110 1720
rect 59990 690 60110 1690
rect 59990 660 59995 690
rect 60025 660 60035 690
rect 60065 660 60075 690
rect 60105 660 60110 690
rect 59990 650 60110 660
rect 59990 620 59995 650
rect 60025 620 60035 650
rect 60065 620 60075 650
rect 60105 620 60110 650
rect 59990 610 60110 620
rect 59990 580 59995 610
rect 60025 580 60035 610
rect 60065 580 60075 610
rect 60105 580 60110 610
rect 58835 -505 58840 165
rect 58860 -505 58865 165
rect 58835 -520 58865 -505
rect 58935 165 58965 175
rect 58935 -505 58940 165
rect 58960 -505 58965 165
rect 59455 135 59490 140
rect 59515 175 59550 180
rect 59515 135 59550 140
rect 58830 -525 58870 -520
rect 58830 -555 58835 -525
rect 58865 -555 58870 -525
rect 58830 -560 58870 -555
rect 58935 -545 58965 -505
rect 58935 -565 58940 -545
rect 58960 -565 58965 -545
rect 58935 -575 58965 -565
rect 57485 -610 57490 -580
rect 57520 -610 57525 -580
rect 57485 -620 57525 -610
rect 57485 -650 57490 -620
rect 57520 -650 57525 -620
rect 57485 -660 57525 -650
rect 57485 -690 57490 -660
rect 57520 -690 57525 -660
rect 57485 -695 57525 -690
rect 57540 -580 57660 -575
rect 57540 -610 57545 -580
rect 57575 -610 57585 -580
rect 57615 -610 57625 -580
rect 57655 -610 57660 -580
rect 57540 -620 57660 -610
rect 57540 -650 57545 -620
rect 57575 -650 57585 -620
rect 57615 -650 57625 -620
rect 57655 -650 57660 -620
rect 57540 -660 57660 -650
rect 57540 -690 57545 -660
rect 57575 -690 57585 -660
rect 57615 -690 57625 -660
rect 57655 -690 57660 -660
rect 57540 -1500 57660 -690
rect 57890 -580 58010 -575
rect 57890 -610 57895 -580
rect 57925 -610 57935 -580
rect 57965 -610 57975 -580
rect 58005 -610 58010 -580
rect 57890 -620 58010 -610
rect 57890 -650 57895 -620
rect 57925 -650 57935 -620
rect 57965 -650 57975 -620
rect 58005 -650 58010 -620
rect 57890 -660 58010 -650
rect 57890 -690 57895 -660
rect 57925 -690 57935 -660
rect 57965 -690 57975 -660
rect 58005 -690 58010 -660
rect 57890 -1500 58010 -690
rect 58240 -580 58365 -575
rect 58240 -610 58245 -580
rect 58275 -610 58285 -580
rect 58315 -610 58325 -580
rect 58355 -610 58365 -580
rect 58240 -620 58365 -610
rect 58240 -650 58245 -620
rect 58275 -650 58285 -620
rect 58315 -650 58325 -620
rect 58355 -650 58365 -620
rect 58240 -660 58365 -650
rect 58240 -690 58245 -660
rect 58275 -690 58285 -660
rect 58315 -690 58325 -660
rect 58355 -690 58365 -660
rect 58240 -695 58365 -690
rect 58530 -580 58570 -575
rect 58530 -610 58535 -580
rect 58565 -610 58570 -580
rect 58530 -620 58570 -610
rect 58530 -650 58535 -620
rect 58565 -650 58570 -620
rect 58530 -660 58570 -650
rect 58530 -690 58535 -660
rect 58565 -690 58570 -660
rect 58530 -695 58570 -690
rect 58590 -580 58710 -575
rect 58590 -610 58595 -580
rect 58625 -610 58635 -580
rect 58665 -610 58675 -580
rect 58705 -610 58710 -580
rect 58590 -620 58710 -610
rect 58590 -650 58595 -620
rect 58625 -650 58635 -620
rect 58665 -650 58675 -620
rect 58705 -650 58710 -620
rect 58590 -660 58710 -650
rect 58590 -690 58595 -660
rect 58625 -690 58635 -660
rect 58665 -690 58675 -660
rect 58705 -690 58710 -660
rect 58240 -1500 58360 -695
rect 58590 -1500 58710 -690
rect 58730 -580 58770 -575
rect 58730 -610 58735 -580
rect 58765 -610 58770 -580
rect 58730 -620 58770 -610
rect 58730 -650 58735 -620
rect 58765 -650 58770 -620
rect 58730 -660 58770 -650
rect 58730 -690 58735 -660
rect 58765 -690 58770 -660
rect 58730 -695 58770 -690
rect 58935 -580 59060 -575
rect 58935 -610 58945 -580
rect 58975 -610 58985 -580
rect 59015 -610 59025 -580
rect 59055 -610 59060 -580
rect 58935 -620 59060 -610
rect 58935 -650 58945 -620
rect 58975 -650 58985 -620
rect 59015 -650 59025 -620
rect 59055 -650 59060 -620
rect 58935 -660 59060 -650
rect 58935 -690 58945 -660
rect 58975 -690 58985 -660
rect 59015 -690 59025 -660
rect 59055 -690 59060 -660
rect 58935 -695 59060 -690
rect 58940 -1500 59060 -695
rect 59290 -580 59410 -575
rect 59290 -610 59295 -580
rect 59325 -610 59335 -580
rect 59365 -610 59375 -580
rect 59405 -610 59410 -580
rect 59290 -620 59410 -610
rect 59290 -650 59295 -620
rect 59325 -650 59335 -620
rect 59365 -650 59375 -620
rect 59405 -650 59410 -620
rect 59290 -660 59410 -650
rect 59290 -690 59295 -660
rect 59325 -690 59335 -660
rect 59365 -690 59375 -660
rect 59405 -690 59410 -660
rect 59290 -1500 59410 -690
rect 59640 -580 59760 -575
rect 59640 -610 59645 -580
rect 59675 -610 59685 -580
rect 59715 -610 59725 -580
rect 59755 -610 59760 -580
rect 59640 -620 59760 -610
rect 59640 -650 59645 -620
rect 59675 -650 59685 -620
rect 59715 -650 59725 -620
rect 59755 -650 59760 -620
rect 59640 -660 59760 -650
rect 59640 -690 59645 -660
rect 59675 -690 59685 -660
rect 59715 -690 59725 -660
rect 59755 -690 59760 -660
rect 59640 -1500 59760 -690
rect 59990 -580 60110 580
rect 59990 -610 59995 -580
rect 60025 -610 60035 -580
rect 60065 -610 60075 -580
rect 60105 -610 60110 -580
rect 59990 -620 60110 -610
rect 59990 -650 59995 -620
rect 60025 -650 60035 -620
rect 60065 -650 60075 -620
rect 60105 -650 60110 -620
rect 59990 -660 60110 -650
rect 59990 -690 59995 -660
rect 60025 -690 60035 -660
rect 60065 -690 60075 -660
rect 60105 -690 60110 -660
rect 59990 -1500 60110 -690
rect 60340 -580 60460 -575
rect 60340 -610 60345 -580
rect 60375 -610 60385 -580
rect 60415 -610 60425 -580
rect 60455 -610 60460 -580
rect 60340 -620 60460 -610
rect 60340 -650 60345 -620
rect 60375 -650 60385 -620
rect 60415 -650 60425 -620
rect 60455 -650 60460 -620
rect 60340 -660 60460 -650
rect 60340 -690 60345 -660
rect 60375 -690 60385 -660
rect 60415 -690 60425 -660
rect 60455 -690 60460 -660
rect 60340 -1500 60460 -690
rect 60690 -580 60810 -575
rect 60690 -610 60695 -580
rect 60725 -610 60735 -580
rect 60765 -610 60775 -580
rect 60805 -610 60810 -580
rect 60690 -620 60810 -610
rect 60690 -650 60695 -620
rect 60725 -650 60735 -620
rect 60765 -650 60775 -620
rect 60805 -650 60810 -620
rect 60690 -660 60810 -650
rect 60690 -690 60695 -660
rect 60725 -690 60735 -660
rect 60765 -690 60775 -660
rect 60805 -690 60810 -660
rect 60690 -1500 60810 -690
rect 61040 -580 61160 -575
rect 61040 -610 61045 -580
rect 61075 -610 61085 -580
rect 61115 -610 61125 -580
rect 61155 -610 61160 -580
rect 61040 -620 61160 -610
rect 61040 -650 61045 -620
rect 61075 -650 61085 -620
rect 61115 -650 61125 -620
rect 61155 -650 61160 -620
rect 61040 -660 61160 -650
rect 61040 -690 61045 -660
rect 61075 -690 61085 -660
rect 61115 -690 61125 -660
rect 61155 -690 61160 -660
rect 61040 -1500 61160 -690
rect 61390 -580 61510 -575
rect 61390 -610 61395 -580
rect 61425 -610 61435 -580
rect 61465 -610 61475 -580
rect 61505 -610 61510 -580
rect 61390 -620 61510 -610
rect 61390 -650 61395 -620
rect 61425 -650 61435 -620
rect 61465 -650 61475 -620
rect 61505 -650 61510 -620
rect 61390 -660 61510 -650
rect 61390 -690 61395 -660
rect 61425 -690 61435 -660
rect 61465 -690 61475 -660
rect 61505 -690 61510 -660
rect 61390 -1500 61510 -690
<< via1 >>
rect 52295 4290 52325 4320
rect 52335 4290 52365 4320
rect 52375 4290 52405 4320
rect 52295 4250 52325 4280
rect 52335 4250 52365 4280
rect 52375 4250 52405 4280
rect 52295 4210 52325 4240
rect 52335 4210 52365 4240
rect 52375 4210 52405 4240
rect 52645 4290 52675 4320
rect 52685 4290 52715 4320
rect 52725 4290 52755 4320
rect 52645 4250 52675 4280
rect 52685 4250 52715 4280
rect 52725 4250 52755 4280
rect 52645 4210 52675 4240
rect 52685 4210 52715 4240
rect 52725 4210 52755 4240
rect 52995 4290 53025 4320
rect 53035 4290 53065 4320
rect 53075 4290 53105 4320
rect 52995 4250 53025 4280
rect 53035 4250 53065 4280
rect 53075 4250 53105 4280
rect 52995 4210 53025 4240
rect 53035 4210 53065 4240
rect 53075 4210 53105 4240
rect 56210 5035 56240 5065
rect 56090 4925 56120 4930
rect 56090 4905 56095 4925
rect 56095 4905 56115 4925
rect 56115 4905 56120 4925
rect 56090 4900 56120 4905
rect 56680 5035 56710 5065
rect 57090 5035 57120 5065
rect 57560 5035 57590 5065
rect 56210 4900 56240 4930
rect 56270 4925 56300 4930
rect 56270 4905 56275 4925
rect 56275 4905 56295 4925
rect 56295 4905 56300 4925
rect 56270 4900 56300 4905
rect 56560 4810 56590 4840
rect 56560 4770 56590 4800
rect 56560 4755 56590 4760
rect 56560 4735 56565 4755
rect 56565 4735 56585 4755
rect 56585 4735 56590 4755
rect 56560 4730 56590 4735
rect 56620 4810 56650 4840
rect 56620 4770 56650 4800
rect 56620 4730 56650 4760
rect 56885 4980 56915 5010
rect 56885 4940 56915 4970
rect 56885 4900 56915 4930
rect 56740 4810 56770 4840
rect 56740 4770 56770 4800
rect 56740 4755 56770 4760
rect 56740 4735 56745 4755
rect 56745 4735 56765 4755
rect 56765 4735 56770 4755
rect 56740 4730 56770 4735
rect 57030 4980 57060 5010
rect 57030 4940 57060 4970
rect 57030 4925 57060 4930
rect 57030 4905 57035 4925
rect 57035 4905 57055 4925
rect 57055 4905 57060 4925
rect 57030 4900 57060 4905
rect 56885 4810 56915 4840
rect 56885 4770 56915 4800
rect 56885 4730 56915 4760
rect 56210 4495 56240 4525
rect 56680 4495 56710 4525
rect 56155 4475 56185 4480
rect 56155 4455 56160 4475
rect 56160 4455 56180 4475
rect 56180 4455 56185 4475
rect 56155 4450 56185 4455
rect 56630 4475 56660 4480
rect 56630 4455 56635 4475
rect 56635 4455 56655 4475
rect 56655 4455 56660 4475
rect 56630 4450 56660 4455
rect 56830 4450 56860 4480
rect 53965 4290 53995 4320
rect 54005 4290 54035 4320
rect 54045 4290 54075 4320
rect 53965 4250 53995 4280
rect 54005 4250 54035 4280
rect 54045 4250 54075 4280
rect 53965 4210 53995 4240
rect 54005 4210 54035 4240
rect 54045 4210 54075 4240
rect 54315 4290 54345 4320
rect 54355 4290 54385 4320
rect 54395 4290 54425 4320
rect 54315 4250 54345 4280
rect 54355 4250 54385 4280
rect 54395 4250 54425 4280
rect 54315 4210 54345 4240
rect 54355 4210 54385 4240
rect 54395 4210 54425 4240
rect 54845 4290 54875 4320
rect 54845 4250 54875 4280
rect 54845 4210 54875 4240
rect 55205 4290 55235 4320
rect 55205 4250 55235 4280
rect 55205 4210 55235 4240
rect 54905 3905 54935 3935
rect 54945 3905 54975 3935
rect 54985 3905 55015 3935
rect 55025 3905 55055 3935
rect 55065 3905 55095 3935
rect 55105 3905 55135 3935
rect 55145 3905 55175 3935
rect 54905 3865 54935 3895
rect 54945 3865 54975 3895
rect 54985 3865 55015 3895
rect 55025 3865 55055 3895
rect 55065 3865 55095 3895
rect 55105 3865 55135 3895
rect 55145 3865 55175 3895
rect 54905 3825 54935 3855
rect 54945 3825 54975 3855
rect 54985 3825 55015 3855
rect 55025 3825 55055 3855
rect 55065 3825 55095 3855
rect 55105 3825 55135 3855
rect 55145 3825 55175 3855
rect 54845 3770 54875 3800
rect 54965 3770 54995 3800
rect 55085 3770 55115 3800
rect 55565 4290 55595 4320
rect 55565 4250 55595 4280
rect 55565 4210 55595 4240
rect 55265 3905 55295 3935
rect 55305 3905 55335 3935
rect 55345 3905 55375 3935
rect 55385 3905 55415 3935
rect 55425 3905 55455 3935
rect 55465 3905 55495 3935
rect 55505 3905 55535 3935
rect 55265 3865 55295 3895
rect 55305 3865 55335 3895
rect 55345 3865 55375 3895
rect 55385 3865 55415 3895
rect 55425 3865 55455 3895
rect 55465 3865 55495 3895
rect 55505 3865 55535 3895
rect 55265 3825 55295 3855
rect 55305 3825 55335 3855
rect 55345 3825 55375 3855
rect 55385 3825 55415 3855
rect 55425 3825 55455 3855
rect 55465 3825 55495 3855
rect 55505 3825 55535 3855
rect 55205 3770 55235 3800
rect 55325 3770 55355 3800
rect 55445 3770 55475 3800
rect 55565 3770 55595 3800
rect 55665 4290 55695 4320
rect 55705 4290 55735 4320
rect 55745 4290 55775 4320
rect 55665 4250 55695 4280
rect 55705 4250 55735 4280
rect 55745 4250 55775 4280
rect 55665 4210 55695 4240
rect 55705 4210 55735 4240
rect 55745 4210 55775 4240
rect 54905 3380 54935 3410
rect 55025 3380 55055 3410
rect 55145 3380 55175 3410
rect 55265 3380 55295 3410
rect 55385 3380 55415 3410
rect 55505 3380 55535 3410
rect 55205 3280 55235 3285
rect 55205 3260 55210 3280
rect 55210 3260 55230 3280
rect 55230 3260 55235 3280
rect 55205 3255 55235 3260
rect 55525 3210 55555 3240
rect 55565 3210 55595 3240
rect 55605 3210 55635 3240
rect 55525 3170 55555 3200
rect 55565 3170 55595 3200
rect 55605 3170 55635 3200
rect 55525 3130 55555 3160
rect 55565 3130 55595 3160
rect 55605 3130 55635 3160
rect 54180 3095 54210 3125
rect 54745 3075 54775 3105
rect 54745 3035 54775 3065
rect 54745 2995 54775 3025
rect 54855 3075 54885 3105
rect 54855 3035 54885 3065
rect 54855 2995 54885 3025
rect 54965 3075 54995 3105
rect 54965 3035 54995 3065
rect 54965 2995 54995 3025
rect 55075 3075 55105 3105
rect 55075 3035 55105 3065
rect 55075 2995 55105 3025
rect 55185 3075 55215 3105
rect 55185 3035 55215 3065
rect 55185 2995 55215 3025
rect 55295 3075 55325 3105
rect 55295 3035 55325 3065
rect 55295 2995 55325 3025
rect 55405 3075 55435 3105
rect 55405 3035 55435 3065
rect 55405 2995 55435 3025
rect 54800 2910 54830 2940
rect 54910 2910 54940 2940
rect 55020 2910 55050 2940
rect 55130 2910 55160 2940
rect 55240 2910 55270 2940
rect 55350 2910 55380 2940
rect 54140 2190 54170 2220
rect 54180 2190 54210 2220
rect 54220 2190 54250 2220
rect 54140 2150 54170 2180
rect 54180 2150 54210 2180
rect 54220 2150 54250 2180
rect 54140 2110 54170 2140
rect 54180 2110 54210 2140
rect 54220 2110 54250 2140
rect 54800 2270 54830 2300
rect 54910 2270 54940 2300
rect 55020 2270 55050 2300
rect 55130 2270 55160 2300
rect 55075 2215 55105 2220
rect 55075 2195 55080 2215
rect 55080 2195 55100 2215
rect 55100 2195 55105 2215
rect 55075 2190 55105 2195
rect 55075 2175 55105 2180
rect 55075 2155 55080 2175
rect 55080 2155 55100 2175
rect 55100 2155 55105 2175
rect 55075 2150 55105 2155
rect 55075 2135 55105 2140
rect 55075 2115 55080 2135
rect 55080 2115 55100 2135
rect 55100 2115 55105 2135
rect 55075 2110 55105 2115
rect 55240 2270 55270 2300
rect 55350 2270 55380 2300
rect 54110 2040 54140 2070
rect 54150 2040 54180 2070
rect 54195 2040 54225 2070
rect 54235 2040 54265 2070
rect 54280 2040 54310 2070
rect 54320 2040 54350 2070
rect 54110 2000 54140 2030
rect 54150 2000 54180 2030
rect 54195 2000 54225 2030
rect 54235 2000 54265 2030
rect 54280 2000 54310 2030
rect 54320 2000 54350 2030
rect 54110 1960 54140 1990
rect 54150 1960 54180 1990
rect 54195 1960 54225 1990
rect 54235 1960 54265 1990
rect 54280 1960 54310 1990
rect 54320 1960 54350 1990
rect 53965 1770 53995 1800
rect 54005 1770 54035 1800
rect 54045 1770 54075 1800
rect 53965 1730 53995 1760
rect 54005 1730 54035 1760
rect 54045 1730 54075 1760
rect 53965 1690 53995 1720
rect 54005 1690 54035 1720
rect 54045 1690 54075 1720
rect 53965 660 53995 690
rect 54005 660 54035 690
rect 54045 660 54075 690
rect 53965 620 53995 650
rect 54005 620 54035 650
rect 54045 620 54075 650
rect 53965 580 53995 610
rect 54005 580 54035 610
rect 54045 580 54075 610
rect 52295 -610 52325 -580
rect 52335 -610 52365 -580
rect 52375 -610 52405 -580
rect 52295 -650 52325 -620
rect 52335 -650 52365 -620
rect 52375 -650 52405 -620
rect 52295 -690 52325 -660
rect 52335 -690 52365 -660
rect 52375 -690 52405 -660
rect 52645 -610 52675 -580
rect 52685 -610 52715 -580
rect 52725 -610 52755 -580
rect 52645 -650 52675 -620
rect 52685 -650 52715 -620
rect 52725 -650 52755 -620
rect 52645 -690 52675 -660
rect 52685 -690 52715 -660
rect 52725 -690 52755 -660
rect 52995 -610 53025 -580
rect 53035 -610 53065 -580
rect 53075 -610 53105 -580
rect 52995 -650 53025 -620
rect 53035 -650 53065 -620
rect 53075 -650 53105 -620
rect 52995 -690 53025 -660
rect 53035 -690 53065 -660
rect 53075 -690 53105 -660
rect 53345 -610 53375 -580
rect 53385 -610 53415 -580
rect 53425 -610 53455 -580
rect 53345 -650 53375 -620
rect 53385 -650 53415 -620
rect 53425 -650 53455 -620
rect 53345 -690 53375 -660
rect 53385 -690 53415 -660
rect 53425 -690 53455 -660
rect 54800 2040 54830 2070
rect 54855 2040 54885 2070
rect 54910 2040 54940 2070
rect 54965 2040 54995 2070
rect 55020 2040 55050 2070
rect 55075 2040 55105 2070
rect 55130 2040 55160 2070
rect 55185 2040 55215 2070
rect 55240 2040 55270 2070
rect 55295 2040 55325 2070
rect 55350 2040 55380 2070
rect 54800 2000 54830 2030
rect 54855 2000 54885 2030
rect 54910 2000 54940 2030
rect 54965 2000 54995 2030
rect 55020 2000 55050 2030
rect 55075 2000 55105 2030
rect 55130 2000 55160 2030
rect 55185 2000 55215 2030
rect 55240 2000 55270 2030
rect 55295 2000 55325 2030
rect 55350 2000 55380 2030
rect 54800 1960 54830 1990
rect 54855 1960 54885 1990
rect 54910 1960 54940 1990
rect 54965 1960 54995 1990
rect 55020 1960 55050 1990
rect 55075 1960 55105 1990
rect 55130 1960 55160 1990
rect 55185 1960 55215 1990
rect 55240 1960 55270 1990
rect 55295 1960 55325 1990
rect 55350 1960 55380 1990
rect 55525 2190 55555 2220
rect 55565 2190 55595 2220
rect 55605 2190 55635 2220
rect 55525 2150 55555 2180
rect 55565 2150 55595 2180
rect 55605 2150 55635 2180
rect 55525 2110 55555 2140
rect 55565 2110 55595 2140
rect 55605 2110 55635 2140
rect 54745 1905 54775 1935
rect 54745 1865 54775 1895
rect 54745 1825 54775 1855
rect 55405 1905 55435 1935
rect 55405 1865 55435 1895
rect 55405 1825 55435 1855
rect 54800 1770 54830 1800
rect 54800 1730 54830 1760
rect 54800 1690 54830 1720
rect 54910 1770 54940 1800
rect 54910 1730 54940 1760
rect 54910 1690 54940 1720
rect 55020 1770 55050 1800
rect 55020 1730 55050 1760
rect 55020 1690 55050 1720
rect 55130 1770 55160 1800
rect 55130 1730 55160 1760
rect 55130 1690 55160 1720
rect 55240 1770 55270 1800
rect 55240 1730 55270 1760
rect 55240 1690 55270 1720
rect 55350 1770 55380 1800
rect 55350 1730 55380 1760
rect 55350 1690 55380 1720
rect 54855 1635 54885 1665
rect 54965 1635 54995 1665
rect 55075 1635 55105 1665
rect 55185 1635 55215 1665
rect 55295 1635 55325 1665
rect 54605 1380 54635 1410
rect 54855 1405 54885 1410
rect 54855 1385 54860 1405
rect 54860 1385 54880 1405
rect 54880 1385 54885 1405
rect 54855 1380 54885 1385
rect 54965 1405 54995 1410
rect 54965 1385 54970 1405
rect 54970 1385 54990 1405
rect 54990 1385 54995 1405
rect 54965 1380 54995 1385
rect 55075 1405 55105 1410
rect 55075 1385 55080 1405
rect 55080 1385 55100 1405
rect 55100 1385 55105 1405
rect 55075 1380 55105 1385
rect 55185 1405 55215 1410
rect 55185 1385 55190 1405
rect 55190 1385 55210 1405
rect 55210 1385 55215 1405
rect 55185 1380 55215 1385
rect 55295 1405 55325 1410
rect 55295 1385 55300 1405
rect 55300 1385 55320 1405
rect 55320 1385 55325 1405
rect 55295 1380 55325 1385
rect 54115 1330 54145 1360
rect 54165 1330 54195 1360
rect 54215 1330 54245 1360
rect 54265 1330 54295 1360
rect 54315 1330 54345 1360
rect 54115 1280 54145 1310
rect 54165 1280 54195 1310
rect 54215 1280 54245 1310
rect 54265 1280 54295 1310
rect 54315 1280 54345 1310
rect 54115 1230 54145 1260
rect 54165 1230 54195 1260
rect 54215 1230 54245 1260
rect 54265 1230 54295 1260
rect 54315 1230 54345 1260
rect 54380 905 54415 910
rect 54380 880 54385 905
rect 54385 880 54410 905
rect 54410 880 54415 905
rect 54380 875 54415 880
rect 54440 905 54475 910
rect 54440 880 54445 905
rect 54445 880 54470 905
rect 54470 880 54475 905
rect 54440 875 54475 880
rect 54500 905 54535 910
rect 54500 880 54505 905
rect 54505 880 54530 905
rect 54530 880 54535 905
rect 54500 875 54535 880
rect 54560 905 54595 910
rect 54560 880 54565 905
rect 54565 880 54590 905
rect 54590 880 54595 905
rect 54560 875 54595 880
rect 55240 1340 55270 1345
rect 55240 1320 55245 1340
rect 55245 1320 55265 1340
rect 55265 1320 55270 1340
rect 55240 1315 55270 1320
rect 55240 1300 55270 1305
rect 55240 1280 55245 1300
rect 55245 1280 55265 1300
rect 55265 1280 55270 1300
rect 55240 1275 55270 1280
rect 55525 1315 55555 1345
rect 55565 1315 55595 1345
rect 55605 1315 55635 1345
rect 55525 1275 55555 1305
rect 55565 1275 55595 1305
rect 55605 1275 55635 1305
rect 56010 3905 56040 3935
rect 56050 3905 56080 3935
rect 56090 3905 56120 3935
rect 56130 3905 56160 3935
rect 56170 3905 56200 3935
rect 56210 3905 56240 3935
rect 56250 3905 56280 3935
rect 56290 3905 56320 3935
rect 56330 3905 56360 3935
rect 56370 3905 56400 3935
rect 56410 3905 56440 3935
rect 56450 3905 56480 3935
rect 56490 3905 56520 3935
rect 56530 3905 56560 3935
rect 56570 3905 56600 3935
rect 56610 3905 56640 3935
rect 56650 3905 56680 3935
rect 56690 3905 56720 3935
rect 56730 3905 56760 3935
rect 56010 3865 56040 3895
rect 56050 3865 56080 3895
rect 56090 3865 56120 3895
rect 56130 3865 56160 3895
rect 56170 3865 56200 3895
rect 56210 3865 56240 3895
rect 56250 3865 56280 3895
rect 56290 3865 56320 3895
rect 56330 3865 56360 3895
rect 56370 3865 56400 3895
rect 56410 3865 56440 3895
rect 56450 3865 56480 3895
rect 56490 3865 56520 3895
rect 56530 3865 56560 3895
rect 56570 3865 56600 3895
rect 56610 3865 56640 3895
rect 56650 3865 56680 3895
rect 56690 3865 56720 3895
rect 56730 3865 56760 3895
rect 56010 3825 56040 3855
rect 56050 3825 56080 3855
rect 56090 3825 56120 3855
rect 56130 3825 56160 3855
rect 56170 3825 56200 3855
rect 56210 3825 56240 3855
rect 56250 3825 56280 3855
rect 56290 3825 56320 3855
rect 56330 3825 56360 3855
rect 56370 3825 56400 3855
rect 56410 3825 56440 3855
rect 56450 3825 56480 3855
rect 56490 3825 56520 3855
rect 56530 3825 56560 3855
rect 56570 3825 56600 3855
rect 56610 3825 56640 3855
rect 56650 3825 56680 3855
rect 56690 3825 56720 3855
rect 56730 3825 56760 3855
rect 56070 3770 56100 3800
rect 56190 3770 56220 3800
rect 56310 3770 56340 3800
rect 56430 3770 56460 3800
rect 56550 3770 56580 3800
rect 56670 3770 56700 3800
rect 56070 3380 56100 3410
rect 56190 3380 56220 3410
rect 56310 3380 56340 3410
rect 56430 3380 56460 3410
rect 56370 3325 56400 3330
rect 56370 3305 56375 3325
rect 56375 3305 56395 3325
rect 56395 3305 56400 3325
rect 56370 3300 56400 3305
rect 56550 3380 56580 3410
rect 56670 3380 56700 3410
rect 57150 4980 57180 5010
rect 57150 4940 57180 4970
rect 57150 4900 57180 4930
rect 57210 4980 57240 5010
rect 57210 4940 57240 4970
rect 57210 4925 57240 4930
rect 57210 4905 57215 4925
rect 57215 4905 57235 4925
rect 57235 4905 57240 4925
rect 57210 4900 57240 4905
rect 57500 4925 57530 4930
rect 57500 4905 57505 4925
rect 57505 4905 57525 4925
rect 57525 4905 57530 4925
rect 57500 4900 57530 4905
rect 57560 4900 57590 4930
rect 57680 4925 57710 4930
rect 57680 4905 57685 4925
rect 57685 4905 57705 4925
rect 57705 4905 57710 4925
rect 57680 4900 57710 4905
rect 57090 4495 57120 4525
rect 57560 4495 57590 4525
rect 56885 4290 56915 4320
rect 56885 4250 56915 4280
rect 56885 4210 56915 4240
rect 56940 4395 56970 4425
rect 57576 4465 57606 4470
rect 57576 4445 57581 4465
rect 57581 4445 57601 4465
rect 57601 4445 57606 4465
rect 57576 4440 57606 4445
rect 56840 3300 56870 3330
rect 57140 4385 57170 4415
rect 57620 4385 57650 4415
rect 58105 4290 58135 4320
rect 58145 4290 58175 4320
rect 58185 4290 58215 4320
rect 58105 4250 58135 4280
rect 58145 4250 58175 4280
rect 58185 4250 58215 4280
rect 58105 4210 58135 4240
rect 58145 4210 58175 4240
rect 58185 4210 58215 4240
rect 57040 3905 57070 3935
rect 57080 3905 57110 3935
rect 57120 3905 57150 3935
rect 57160 3905 57190 3935
rect 57200 3905 57230 3935
rect 57240 3905 57270 3935
rect 57280 3905 57310 3935
rect 57320 3905 57350 3935
rect 57360 3905 57390 3935
rect 57400 3905 57430 3935
rect 57440 3905 57470 3935
rect 57480 3905 57510 3935
rect 57520 3905 57550 3935
rect 57560 3905 57590 3935
rect 57600 3905 57630 3935
rect 57640 3905 57670 3935
rect 57680 3905 57710 3935
rect 57720 3905 57750 3935
rect 57760 3905 57790 3935
rect 57040 3865 57070 3895
rect 57080 3865 57110 3895
rect 57120 3865 57150 3895
rect 57160 3865 57190 3895
rect 57200 3865 57230 3895
rect 57240 3865 57270 3895
rect 57280 3865 57310 3895
rect 57320 3865 57350 3895
rect 57360 3865 57390 3895
rect 57400 3865 57430 3895
rect 57440 3865 57470 3895
rect 57480 3865 57510 3895
rect 57520 3865 57550 3895
rect 57560 3865 57590 3895
rect 57600 3865 57630 3895
rect 57640 3865 57670 3895
rect 57680 3865 57710 3895
rect 57720 3865 57750 3895
rect 57760 3865 57790 3895
rect 57040 3825 57070 3855
rect 57080 3825 57110 3855
rect 57120 3825 57150 3855
rect 57160 3825 57190 3855
rect 57200 3825 57230 3855
rect 57240 3825 57270 3855
rect 57280 3825 57310 3855
rect 57320 3825 57350 3855
rect 57360 3825 57390 3855
rect 57400 3825 57430 3855
rect 57440 3825 57470 3855
rect 57480 3825 57510 3855
rect 57520 3825 57550 3855
rect 57560 3825 57590 3855
rect 57600 3825 57630 3855
rect 57640 3825 57670 3855
rect 57680 3825 57710 3855
rect 57720 3825 57750 3855
rect 57760 3825 57790 3855
rect 57100 3770 57130 3800
rect 57220 3770 57250 3800
rect 57340 3770 57370 3800
rect 57460 3770 57490 3800
rect 57580 3770 57610 3800
rect 57700 3770 57730 3800
rect 57100 3380 57130 3410
rect 56930 3255 56960 3285
rect 56070 3210 56100 3240
rect 56110 3210 56140 3240
rect 56150 3210 56180 3240
rect 56190 3210 56220 3240
rect 56230 3210 56260 3240
rect 56270 3210 56300 3240
rect 56310 3210 56340 3240
rect 56350 3210 56380 3240
rect 56390 3210 56420 3240
rect 56430 3210 56460 3240
rect 56470 3210 56500 3240
rect 56510 3210 56540 3240
rect 56550 3210 56580 3240
rect 56590 3210 56620 3240
rect 56630 3210 56660 3240
rect 56670 3210 56700 3240
rect 56070 3170 56100 3200
rect 56110 3170 56140 3200
rect 56150 3170 56180 3200
rect 56190 3170 56220 3200
rect 56230 3170 56260 3200
rect 56270 3170 56300 3200
rect 56310 3170 56340 3200
rect 56350 3170 56380 3200
rect 56390 3170 56420 3200
rect 56430 3170 56460 3200
rect 56470 3170 56500 3200
rect 56510 3170 56540 3200
rect 56550 3170 56580 3200
rect 56590 3170 56620 3200
rect 56630 3170 56660 3200
rect 56670 3170 56700 3200
rect 56070 3130 56100 3160
rect 56110 3130 56140 3160
rect 56150 3130 56180 3160
rect 56190 3130 56220 3160
rect 56230 3130 56260 3160
rect 56270 3130 56300 3160
rect 56310 3130 56340 3160
rect 56350 3130 56380 3160
rect 56390 3130 56420 3160
rect 56430 3130 56460 3160
rect 56470 3130 56500 3160
rect 56510 3130 56540 3160
rect 56550 3130 56580 3160
rect 56590 3130 56620 3160
rect 56630 3130 56660 3160
rect 56670 3130 56700 3160
rect 57220 3380 57250 3410
rect 57340 3380 57370 3410
rect 57460 3380 57490 3410
rect 57400 3325 57430 3330
rect 57400 3305 57405 3325
rect 57405 3305 57425 3325
rect 57425 3305 57430 3325
rect 57400 3300 57430 3305
rect 57580 3380 57610 3410
rect 57700 3380 57730 3410
rect 57100 3210 57130 3240
rect 57140 3210 57170 3240
rect 57180 3210 57210 3240
rect 57220 3210 57250 3240
rect 57260 3210 57290 3240
rect 57300 3210 57330 3240
rect 57340 3210 57370 3240
rect 57380 3210 57410 3240
rect 57420 3210 57450 3240
rect 57460 3210 57490 3240
rect 57500 3210 57530 3240
rect 57540 3210 57570 3240
rect 57580 3210 57610 3240
rect 57620 3210 57650 3240
rect 57660 3210 57690 3240
rect 57700 3210 57730 3240
rect 57100 3170 57130 3200
rect 57140 3170 57170 3200
rect 57180 3170 57210 3200
rect 57220 3170 57250 3200
rect 57260 3170 57290 3200
rect 57300 3170 57330 3200
rect 57340 3170 57370 3200
rect 57380 3170 57410 3200
rect 57420 3170 57450 3200
rect 57460 3170 57490 3200
rect 57500 3170 57530 3200
rect 57540 3170 57570 3200
rect 57580 3170 57610 3200
rect 57620 3170 57650 3200
rect 57660 3170 57690 3200
rect 57700 3170 57730 3200
rect 57100 3130 57130 3160
rect 57140 3130 57170 3160
rect 57180 3130 57210 3160
rect 57220 3130 57250 3160
rect 57260 3130 57290 3160
rect 57300 3130 57330 3160
rect 57340 3130 57370 3160
rect 57380 3130 57410 3160
rect 57420 3130 57450 3160
rect 57460 3130 57490 3160
rect 57500 3130 57530 3160
rect 57540 3130 57570 3160
rect 57580 3130 57610 3160
rect 57620 3130 57650 3160
rect 57660 3130 57690 3160
rect 57700 3130 57730 3160
rect 55665 3075 55695 3105
rect 55705 3075 55735 3105
rect 55745 3075 55775 3105
rect 58415 4290 58445 4320
rect 58415 4250 58445 4280
rect 58415 4210 58445 4240
rect 58775 4290 58805 4320
rect 58775 4250 58805 4280
rect 58775 4210 58805 4240
rect 58475 3905 58505 3935
rect 58515 3905 58545 3935
rect 58555 3905 58585 3935
rect 58595 3905 58625 3935
rect 58635 3905 58665 3935
rect 58675 3905 58705 3935
rect 58715 3905 58745 3935
rect 58475 3865 58505 3895
rect 58515 3865 58545 3895
rect 58555 3865 58585 3895
rect 58595 3865 58625 3895
rect 58635 3865 58665 3895
rect 58675 3865 58705 3895
rect 58715 3865 58745 3895
rect 58475 3825 58505 3855
rect 58515 3825 58545 3855
rect 58555 3825 58585 3855
rect 58595 3825 58625 3855
rect 58635 3825 58665 3855
rect 58675 3825 58705 3855
rect 58715 3825 58745 3855
rect 58415 3770 58445 3800
rect 58535 3770 58565 3800
rect 58655 3770 58685 3800
rect 59135 4290 59165 4320
rect 59135 4250 59165 4280
rect 59135 4210 59165 4240
rect 58835 3905 58865 3935
rect 58875 3905 58905 3935
rect 58915 3905 58945 3935
rect 58955 3905 58985 3935
rect 58995 3905 59025 3935
rect 59035 3905 59065 3935
rect 59075 3905 59105 3935
rect 58835 3865 58865 3895
rect 58875 3865 58905 3895
rect 58915 3865 58945 3895
rect 58955 3865 58985 3895
rect 58995 3865 59025 3895
rect 59035 3865 59065 3895
rect 59075 3865 59105 3895
rect 58835 3825 58865 3855
rect 58875 3825 58905 3855
rect 58915 3825 58945 3855
rect 58955 3825 58985 3855
rect 58995 3825 59025 3855
rect 59035 3825 59065 3855
rect 59075 3825 59105 3855
rect 58775 3770 58805 3800
rect 58895 3770 58925 3800
rect 59015 3770 59045 3800
rect 59645 4290 59675 4320
rect 59685 4290 59715 4320
rect 59725 4290 59755 4320
rect 59645 4250 59675 4280
rect 59685 4250 59715 4280
rect 59725 4250 59755 4280
rect 59645 4210 59675 4240
rect 59685 4210 59715 4240
rect 59725 4210 59755 4240
rect 59995 4290 60025 4320
rect 60035 4290 60065 4320
rect 60075 4290 60105 4320
rect 59995 4250 60025 4280
rect 60035 4250 60065 4280
rect 60075 4250 60105 4280
rect 59995 4210 60025 4240
rect 60035 4210 60065 4240
rect 60075 4210 60105 4240
rect 60695 4290 60725 4320
rect 60735 4290 60765 4320
rect 60775 4290 60805 4320
rect 60695 4250 60725 4280
rect 60735 4250 60765 4280
rect 60775 4250 60805 4280
rect 60695 4210 60725 4240
rect 60735 4210 60765 4240
rect 60775 4210 60805 4240
rect 61045 4290 61075 4320
rect 61085 4290 61115 4320
rect 61125 4290 61155 4320
rect 61045 4250 61075 4280
rect 61085 4250 61115 4280
rect 61125 4250 61155 4280
rect 61045 4210 61075 4240
rect 61085 4210 61115 4240
rect 61125 4210 61155 4240
rect 61395 4290 61425 4320
rect 61435 4290 61465 4320
rect 61475 4290 61505 4320
rect 61395 4250 61425 4280
rect 61435 4250 61465 4280
rect 61475 4250 61505 4280
rect 61395 4210 61425 4240
rect 61435 4210 61465 4240
rect 61475 4210 61505 4240
rect 59135 3770 59165 3800
rect 58475 3380 58505 3410
rect 58595 3380 58625 3410
rect 58715 3380 58745 3410
rect 58835 3380 58865 3410
rect 58955 3380 58985 3410
rect 59075 3380 59105 3410
rect 58775 3280 58805 3285
rect 58775 3260 58780 3280
rect 58780 3260 58800 3280
rect 58800 3260 58805 3280
rect 58775 3255 58805 3260
rect 55665 3035 55695 3065
rect 55705 3035 55735 3065
rect 55745 3035 55775 3065
rect 55665 2995 55695 3025
rect 55705 2995 55735 3025
rect 55745 2995 55775 3025
rect 56515 3065 56545 3095
rect 56515 3025 56545 3055
rect 56515 3010 56545 3015
rect 56515 2990 56520 3010
rect 56520 2990 56540 3010
rect 56540 2990 56545 3010
rect 56515 2985 56545 2990
rect 56680 3065 56710 3095
rect 56680 3025 56710 3055
rect 56680 3010 56710 3015
rect 56680 2990 56685 3010
rect 56685 2990 56705 3010
rect 56705 2990 56710 3010
rect 56680 2985 56710 2990
rect 56845 3065 56875 3095
rect 56845 3025 56875 3055
rect 56845 3010 56875 3015
rect 56845 2990 56850 3010
rect 56850 2990 56870 3010
rect 56870 2990 56875 3010
rect 56845 2985 56875 2990
rect 56925 3065 56955 3095
rect 56925 3025 56955 3055
rect 56925 3010 56955 3015
rect 56925 2990 56930 3010
rect 56930 2990 56950 3010
rect 56950 2990 56955 3010
rect 56925 2985 56955 2990
rect 57090 3065 57120 3095
rect 57090 3025 57120 3055
rect 57090 3010 57120 3015
rect 57090 2990 57095 3010
rect 57095 2990 57115 3010
rect 57115 2990 57120 3010
rect 57090 2985 57120 2990
rect 57255 3065 57285 3095
rect 57255 3025 57285 3055
rect 57255 3010 57285 3015
rect 57255 2990 57260 3010
rect 57260 2990 57280 3010
rect 57280 2990 57285 3010
rect 57255 2985 57285 2990
rect 58105 3075 58135 3105
rect 58145 3075 58175 3105
rect 58185 3075 58215 3105
rect 58105 3035 58135 3065
rect 58145 3035 58175 3065
rect 58185 3035 58215 3065
rect 58105 2995 58135 3025
rect 58145 2995 58175 3025
rect 58185 2995 58215 3025
rect 56625 2955 56655 2960
rect 56625 2935 56630 2955
rect 56630 2935 56650 2955
rect 56650 2935 56655 2955
rect 56625 2930 56655 2935
rect 56735 2955 56765 2960
rect 56735 2935 56740 2955
rect 56740 2935 56760 2955
rect 56760 2935 56765 2955
rect 56735 2930 56765 2935
rect 57035 2955 57065 2960
rect 57035 2935 57040 2955
rect 57040 2935 57060 2955
rect 57060 2935 57065 2955
rect 57035 2930 57065 2935
rect 57145 2955 57175 2960
rect 57145 2935 57150 2955
rect 57150 2935 57170 2955
rect 57170 2935 57175 2955
rect 57145 2930 57175 2935
rect 56560 2645 56590 2650
rect 56800 2645 56830 2650
rect 56560 2625 56565 2645
rect 56565 2625 56585 2645
rect 56585 2625 56590 2645
rect 56560 2620 56590 2625
rect 56680 2635 56710 2640
rect 56680 2615 56685 2635
rect 56685 2615 56705 2635
rect 56705 2615 56710 2635
rect 56680 2610 56710 2615
rect 56800 2625 56805 2645
rect 56805 2625 56825 2645
rect 56825 2625 56830 2645
rect 56800 2620 56830 2625
rect 56605 2575 56635 2580
rect 56605 2555 56610 2575
rect 56610 2555 56630 2575
rect 56630 2555 56635 2575
rect 56605 2550 56635 2555
rect 55945 2500 55975 2530
rect 56750 2500 56780 2530
rect 55665 1905 55695 1935
rect 55705 1905 55735 1935
rect 55745 1905 55775 1935
rect 55665 1865 55695 1895
rect 55705 1865 55735 1895
rect 55745 1865 55775 1895
rect 55665 1825 55695 1855
rect 55705 1825 55735 1855
rect 55745 1825 55775 1855
rect 54650 1195 54680 1225
rect 54855 1195 54885 1225
rect 54965 1195 54995 1225
rect 55075 1195 55105 1225
rect 55185 1195 55215 1225
rect 55295 1195 55325 1225
rect 54650 875 54680 905
rect 54505 805 54535 835
rect 54605 805 54635 835
rect 54855 855 54885 885
rect 54965 855 54995 885
rect 55075 855 55105 885
rect 55185 855 55215 885
rect 55295 855 55325 885
rect 54800 795 54830 825
rect 54800 755 54830 785
rect 54800 715 54830 745
rect 54910 795 54940 825
rect 54910 755 54940 785
rect 54910 715 54940 745
rect 55020 795 55050 825
rect 55020 755 55050 785
rect 55020 715 55050 745
rect 55130 795 55160 825
rect 55130 755 55160 785
rect 55130 715 55160 745
rect 55240 795 55270 825
rect 55240 755 55270 785
rect 55240 715 55270 745
rect 55350 795 55380 825
rect 55350 755 55380 785
rect 55350 715 55380 745
rect 55900 1705 55930 1735
rect 55665 795 55695 825
rect 55705 795 55735 825
rect 55745 795 55775 825
rect 55665 755 55695 785
rect 55705 755 55735 785
rect 55745 755 55775 785
rect 55665 715 55695 745
rect 55705 715 55735 745
rect 55745 715 55775 745
rect 55800 1205 55830 1235
rect 55840 1205 55870 1235
rect 55800 1165 55830 1195
rect 55840 1165 55870 1195
rect 55800 1125 55830 1155
rect 55840 1125 55870 1155
rect 54745 660 54775 690
rect 54745 620 54775 650
rect 54745 580 54775 610
rect 55405 660 55435 690
rect 55405 620 55435 650
rect 55405 580 55435 610
rect 54385 525 54415 555
rect 54520 480 54550 510
rect 55105 505 55135 510
rect 55105 485 55110 505
rect 55110 485 55130 505
rect 55130 485 55135 505
rect 55105 480 55135 485
rect 54110 280 54140 310
rect 54150 280 54180 310
rect 54195 280 54225 310
rect 54235 280 54265 310
rect 54280 280 54310 310
rect 54320 280 54350 310
rect 54110 240 54140 270
rect 54150 240 54180 270
rect 54195 240 54225 270
rect 54235 240 54265 270
rect 54280 240 54310 270
rect 54320 240 54350 270
rect 54110 200 54140 230
rect 54150 200 54180 230
rect 54195 200 54225 230
rect 54235 200 54265 230
rect 54280 200 54310 230
rect 54320 200 54350 230
rect 54585 280 54615 310
rect 54585 240 54615 270
rect 54585 200 54615 230
rect 54855 280 54885 310
rect 54895 280 54925 310
rect 54935 280 54965 310
rect 54975 280 55005 310
rect 55015 280 55045 310
rect 55055 280 55085 310
rect 55095 280 55125 310
rect 55135 280 55165 310
rect 55175 280 55205 310
rect 55215 280 55245 310
rect 55255 280 55285 310
rect 54855 240 54885 270
rect 54895 240 54925 270
rect 54935 240 54965 270
rect 54975 240 55005 270
rect 55015 240 55045 270
rect 55055 240 55085 270
rect 55095 240 55125 270
rect 55135 240 55165 270
rect 55175 240 55205 270
rect 55215 240 55245 270
rect 55255 240 55285 270
rect 54855 200 54885 230
rect 54895 200 54925 230
rect 54935 200 54965 230
rect 54975 200 55005 230
rect 55015 200 55045 230
rect 55055 200 55085 230
rect 55095 200 55125 230
rect 55135 200 55165 230
rect 55175 200 55205 230
rect 55215 200 55245 230
rect 55255 200 55285 230
rect 54520 170 54555 175
rect 54520 145 54525 170
rect 54525 145 54550 170
rect 54550 145 54555 170
rect 54520 140 54555 145
rect 54580 170 54615 175
rect 54580 145 54585 170
rect 54585 145 54610 170
rect 54610 145 54615 170
rect 54580 140 54615 145
rect 54855 -555 54885 -525
rect 55055 -555 55085 -525
rect 55800 -125 55830 -95
rect 55840 -125 55870 -95
rect 55800 -165 55830 -135
rect 55840 -165 55870 -135
rect 55800 -205 55830 -175
rect 55840 -205 55870 -175
rect 57090 2635 57120 2640
rect 57090 2615 57095 2635
rect 57095 2615 57115 2635
rect 57115 2615 57120 2635
rect 57090 2610 57120 2615
rect 57165 2575 57195 2580
rect 57165 2555 57170 2575
rect 57170 2555 57190 2575
rect 57190 2555 57195 2575
rect 57165 2550 57195 2555
rect 57020 2500 57050 2530
rect 56855 2445 56885 2475
rect 56965 2445 56995 2475
rect 57825 2500 57855 2530
rect 56940 2390 56970 2420
rect 57215 2390 57245 2420
rect 56855 2360 56885 2365
rect 56855 2340 56860 2360
rect 56860 2340 56880 2360
rect 56880 2340 56885 2360
rect 56855 2335 56885 2340
rect 56090 2190 56120 2220
rect 56145 2190 56175 2220
rect 56200 2190 56230 2220
rect 56255 2190 56285 2220
rect 56310 2190 56340 2220
rect 56365 2190 56395 2220
rect 56420 2190 56450 2220
rect 56475 2190 56505 2220
rect 56530 2190 56560 2220
rect 56585 2190 56615 2220
rect 56640 2190 56670 2220
rect 56090 2150 56120 2180
rect 56145 2150 56175 2180
rect 56200 2150 56230 2180
rect 56255 2150 56285 2180
rect 56310 2150 56340 2180
rect 56365 2150 56395 2180
rect 56420 2150 56450 2180
rect 56475 2150 56505 2180
rect 56530 2150 56560 2180
rect 56585 2150 56615 2180
rect 56640 2150 56670 2180
rect 56090 2110 56120 2140
rect 56145 2110 56175 2140
rect 56200 2110 56230 2140
rect 56255 2110 56285 2140
rect 56310 2110 56340 2140
rect 56365 2110 56395 2140
rect 56420 2110 56450 2140
rect 56475 2110 56505 2140
rect 56530 2110 56560 2140
rect 56585 2110 56615 2140
rect 56640 2110 56670 2140
rect 55995 1730 56025 1735
rect 55995 1710 56000 1730
rect 56000 1710 56020 1730
rect 56020 1710 56025 1730
rect 55995 1705 56025 1710
rect 56145 1695 56175 1725
rect 56090 1650 56120 1680
rect 56255 1695 56285 1725
rect 56200 1650 56230 1680
rect 56145 1460 56175 1490
rect 56090 1415 56120 1445
rect 56035 1360 56065 1390
rect 56035 1320 56065 1350
rect 56035 1280 56065 1310
rect 56365 1695 56395 1725
rect 56310 1650 56340 1680
rect 56255 1460 56285 1490
rect 56200 1415 56230 1445
rect 56040 1040 56070 1045
rect 56040 1020 56045 1040
rect 56045 1020 56065 1040
rect 56065 1020 56070 1040
rect 56090 1025 56120 1055
rect 56145 1035 56175 1065
rect 56475 1695 56505 1725
rect 56420 1650 56450 1680
rect 56365 1460 56395 1490
rect 56310 1415 56340 1445
rect 56200 1025 56230 1055
rect 56255 1035 56285 1065
rect 56585 1695 56615 1725
rect 56530 1650 56560 1680
rect 56475 1460 56505 1490
rect 56420 1415 56450 1445
rect 56310 1025 56340 1055
rect 56365 1035 56395 1065
rect 57130 2190 57160 2220
rect 57185 2190 57215 2220
rect 57240 2190 57270 2220
rect 57295 2190 57325 2220
rect 57350 2190 57380 2220
rect 57405 2190 57435 2220
rect 57460 2190 57490 2220
rect 57515 2190 57545 2220
rect 57570 2190 57600 2220
rect 57625 2190 57655 2220
rect 57680 2190 57710 2220
rect 57130 2150 57160 2180
rect 57185 2150 57215 2180
rect 57240 2150 57270 2180
rect 57295 2150 57325 2180
rect 57350 2150 57380 2180
rect 57405 2150 57435 2180
rect 57460 2150 57490 2180
rect 57515 2150 57545 2180
rect 57570 2150 57600 2180
rect 57625 2150 57655 2180
rect 57680 2150 57710 2180
rect 57130 2110 57160 2140
rect 57185 2110 57215 2140
rect 57240 2110 57270 2140
rect 57295 2110 57325 2140
rect 57350 2110 57380 2140
rect 57405 2110 57435 2140
rect 57460 2110 57490 2140
rect 57515 2110 57545 2140
rect 57570 2110 57600 2140
rect 57625 2110 57655 2140
rect 57680 2110 57710 2140
rect 56775 2040 56805 2045
rect 56775 2020 56780 2040
rect 56780 2020 56800 2040
rect 56800 2020 56805 2040
rect 56775 2015 56805 2020
rect 56775 1975 56805 2005
rect 56775 1935 56805 1965
rect 56885 2015 56915 2045
rect 56885 1975 56915 2005
rect 56885 1935 56915 1965
rect 56995 2040 57025 2045
rect 56995 2020 57000 2040
rect 57000 2020 57020 2040
rect 57020 2020 57025 2040
rect 56995 2015 57025 2020
rect 56995 1975 57025 2005
rect 56995 1935 57025 1965
rect 56690 1730 56720 1735
rect 56690 1710 56695 1730
rect 56695 1710 56715 1730
rect 56715 1710 56720 1730
rect 56690 1705 56720 1710
rect 57080 1730 57110 1735
rect 57080 1710 57085 1730
rect 57085 1710 57105 1730
rect 57105 1710 57110 1730
rect 57080 1705 57110 1710
rect 56640 1650 56670 1680
rect 57185 1695 57215 1725
rect 57130 1650 57160 1680
rect 56585 1460 56615 1490
rect 56530 1415 56560 1445
rect 56420 1025 56450 1055
rect 56475 1035 56505 1065
rect 56640 1415 56670 1445
rect 57295 1695 57325 1725
rect 57240 1650 57270 1680
rect 57185 1460 57215 1490
rect 57130 1415 57160 1445
rect 56695 1360 56725 1390
rect 56695 1320 56725 1350
rect 56695 1280 56725 1310
rect 57075 1360 57105 1390
rect 57075 1320 57105 1350
rect 57075 1280 57105 1310
rect 56885 1205 56915 1235
rect 56885 1165 56915 1195
rect 56885 1125 56915 1155
rect 56530 1025 56560 1055
rect 56585 1035 56615 1065
rect 56640 1025 56670 1055
rect 56690 1050 56720 1055
rect 56690 1030 56695 1050
rect 56695 1030 56715 1050
rect 56715 1030 56720 1050
rect 56690 1025 56720 1030
rect 56840 1050 56870 1055
rect 56840 1030 56845 1050
rect 56845 1030 56865 1050
rect 56865 1030 56870 1050
rect 56840 1025 56870 1030
rect 56040 1015 56070 1020
rect 56145 980 56175 1010
rect 56090 785 56120 815
rect 56255 980 56285 1010
rect 56200 785 56230 815
rect 56365 980 56395 1010
rect 56310 785 56340 815
rect 56475 980 56505 1010
rect 56420 785 56450 815
rect 56585 980 56615 1010
rect 56530 785 56560 815
rect 56640 785 56670 815
rect 57405 1695 57435 1725
rect 57350 1650 57380 1680
rect 57295 1460 57325 1490
rect 57240 1415 57270 1445
rect 56930 1050 56960 1055
rect 56930 1030 56935 1050
rect 56935 1030 56955 1050
rect 56955 1030 56960 1050
rect 56930 1025 56960 1030
rect 57080 1050 57110 1055
rect 57080 1030 57085 1050
rect 57085 1030 57105 1050
rect 57105 1030 57110 1050
rect 57080 1025 57110 1030
rect 57130 1025 57160 1055
rect 57185 1035 57215 1065
rect 57515 1695 57545 1725
rect 57460 1650 57490 1680
rect 57405 1460 57435 1490
rect 57350 1415 57380 1445
rect 57240 1025 57270 1055
rect 57295 1035 57325 1065
rect 57625 1695 57655 1725
rect 57570 1650 57600 1680
rect 57515 1460 57545 1490
rect 57460 1415 57490 1445
rect 57350 1025 57380 1055
rect 57405 1035 57435 1065
rect 57680 1650 57710 1680
rect 57625 1460 57655 1490
rect 57570 1415 57600 1445
rect 57460 1025 57490 1055
rect 57515 1035 57545 1065
rect 57680 1415 57710 1445
rect 57735 1360 57765 1390
rect 57735 1320 57765 1350
rect 57735 1280 57765 1310
rect 57570 1025 57600 1055
rect 57625 1035 57655 1065
rect 57680 1025 57710 1055
rect 57730 1040 57760 1045
rect 57730 1020 57735 1040
rect 57735 1020 57755 1040
rect 57755 1020 57760 1040
rect 57185 980 57215 1010
rect 56830 785 56860 815
rect 56145 715 56175 745
rect 56255 715 56285 745
rect 56365 715 56395 745
rect 56475 715 56505 745
rect 56585 715 56615 745
rect 56035 660 56065 690
rect 56035 620 56065 650
rect 56035 580 56065 610
rect 55945 525 55975 555
rect 56735 660 56765 690
rect 56735 620 56765 650
rect 56735 580 56765 610
rect 56445 360 56475 390
rect 56555 360 56585 390
rect 56665 360 56695 390
rect 56775 360 56805 390
rect 56940 785 56970 815
rect 56885 360 56915 390
rect 57130 785 57160 815
rect 57295 980 57325 1010
rect 57240 785 57270 815
rect 57405 980 57435 1010
rect 57350 785 57380 815
rect 57515 980 57545 1010
rect 57460 785 57490 815
rect 57625 980 57655 1010
rect 57570 785 57600 815
rect 57730 1015 57760 1020
rect 57680 785 57710 815
rect 57185 715 57215 745
rect 57295 715 57325 745
rect 57035 660 57065 690
rect 57035 620 57065 650
rect 57035 580 57065 610
rect 56995 360 57025 390
rect 57405 715 57435 745
rect 57515 715 57545 745
rect 57625 715 57655 745
rect 57735 660 57765 690
rect 57735 620 57765 650
rect 57735 580 57765 610
rect 57870 2390 57900 2420
rect 57825 525 57855 555
rect 57105 360 57135 390
rect 57215 360 57245 390
rect 57325 360 57355 390
rect 57435 360 57465 390
rect 56225 55 56255 60
rect 56225 35 56230 55
rect 56230 35 56250 55
rect 56250 35 56255 55
rect 56225 30 56255 35
rect 55900 -305 55930 -275
rect 55255 -555 55285 -525
rect 56280 30 56310 60
rect 56390 30 56420 60
rect 56500 30 56530 60
rect 56610 30 56640 60
rect 56720 30 56750 60
rect 56830 30 56860 60
rect 56940 30 56970 60
rect 57050 30 57080 60
rect 57160 30 57190 60
rect 57270 30 57300 60
rect 57380 30 57410 60
rect 57490 55 57520 60
rect 57490 35 57495 55
rect 57495 35 57515 55
rect 57515 35 57520 55
rect 57490 30 57520 35
rect 56445 -15 56475 15
rect 56555 -15 56585 15
rect 56665 -15 56695 15
rect 56775 -15 56805 15
rect 56885 -15 56915 15
rect 56995 -15 57025 15
rect 57105 -15 57135 15
rect 57215 -15 57245 15
rect 57325 -15 57355 15
rect 57435 -15 57465 15
rect 56335 -125 56365 -95
rect 56335 -165 56365 -135
rect 56335 -205 56365 -175
rect 56545 -260 56575 -230
rect 56655 -260 56685 -230
rect 56875 -260 56905 -230
rect 56490 -305 56520 -275
rect 56600 -280 56630 -275
rect 56600 -300 56605 -280
rect 56605 -300 56625 -280
rect 56625 -300 56630 -280
rect 56600 -305 56630 -300
rect 56545 -510 56575 -480
rect 56710 -305 56740 -275
rect 56655 -510 56685 -480
rect 57045 -280 57075 -275
rect 57045 -300 57050 -280
rect 57050 -300 57070 -280
rect 57070 -300 57075 -280
rect 57045 -305 57075 -300
rect 57420 -45 57450 -40
rect 57420 -65 57425 -45
rect 57425 -65 57445 -45
rect 57445 -65 57450 -45
rect 57420 -70 57450 -65
rect 56875 -510 56905 -480
rect 56490 -555 56520 -525
rect 56600 -555 56630 -525
rect 56710 -555 56740 -525
rect 53965 -610 53995 -580
rect 54005 -610 54035 -580
rect 54045 -610 54075 -580
rect 53965 -650 53995 -620
rect 54005 -650 54035 -620
rect 54045 -650 54075 -620
rect 53965 -690 53995 -660
rect 54005 -690 54035 -660
rect 54045 -690 54075 -660
rect 54395 -610 54425 -580
rect 54435 -610 54465 -580
rect 54475 -610 54505 -580
rect 54395 -650 54425 -620
rect 54435 -650 54465 -620
rect 54475 -650 54505 -620
rect 54395 -690 54425 -660
rect 54435 -690 54465 -660
rect 54475 -690 54505 -660
rect 54745 -610 54775 -580
rect 54785 -610 54815 -580
rect 54825 -610 54855 -580
rect 54745 -650 54775 -620
rect 54785 -650 54815 -620
rect 54825 -650 54855 -620
rect 54745 -690 54775 -660
rect 54785 -690 54815 -660
rect 54825 -690 54855 -660
rect 55035 -610 55065 -580
rect 55035 -650 55065 -620
rect 55035 -690 55065 -660
rect 55095 -610 55125 -580
rect 55135 -610 55165 -580
rect 55175 -610 55205 -580
rect 55095 -650 55125 -620
rect 55135 -650 55165 -620
rect 55175 -650 55205 -620
rect 55095 -690 55125 -660
rect 55135 -690 55165 -660
rect 55175 -690 55205 -660
rect 55235 -610 55265 -580
rect 55235 -650 55265 -620
rect 55235 -690 55265 -660
rect 55445 -610 55475 -580
rect 55485 -610 55515 -580
rect 55525 -610 55555 -580
rect 55445 -650 55475 -620
rect 55485 -650 55515 -620
rect 55525 -650 55555 -620
rect 55445 -690 55475 -660
rect 55485 -690 55515 -660
rect 55525 -690 55555 -660
rect 55795 -610 55825 -580
rect 55835 -610 55865 -580
rect 55875 -610 55905 -580
rect 55795 -650 55825 -620
rect 55835 -650 55865 -620
rect 55875 -650 55905 -620
rect 55795 -690 55825 -660
rect 55835 -690 55865 -660
rect 55875 -690 55905 -660
rect 56145 -610 56175 -580
rect 56185 -610 56215 -580
rect 56225 -610 56255 -580
rect 56145 -650 56175 -620
rect 56185 -650 56215 -620
rect 56225 -650 56255 -620
rect 56145 -690 56175 -660
rect 56185 -690 56215 -660
rect 56225 -690 56255 -660
rect 56435 -610 56465 -580
rect 56435 -650 56465 -620
rect 56435 -690 56465 -660
rect 56495 -610 56525 -580
rect 56535 -610 56565 -580
rect 56575 -610 56605 -580
rect 56495 -650 56525 -620
rect 56535 -650 56565 -620
rect 56575 -650 56605 -620
rect 56495 -690 56525 -660
rect 56535 -690 56565 -660
rect 56575 -690 56605 -660
rect 56765 -610 56795 -580
rect 56765 -650 56795 -620
rect 56765 -690 56795 -660
rect 56845 -610 56875 -580
rect 56885 -610 56915 -580
rect 56925 -610 56955 -580
rect 56845 -650 56875 -620
rect 56885 -650 56915 -620
rect 56925 -650 56955 -620
rect 56845 -690 56875 -660
rect 56885 -690 56915 -660
rect 56925 -690 56955 -660
rect 57195 -610 57225 -580
rect 57235 -610 57265 -580
rect 57275 -610 57305 -580
rect 57195 -650 57225 -620
rect 57235 -650 57265 -620
rect 57275 -650 57305 -620
rect 57195 -690 57225 -660
rect 57235 -690 57265 -660
rect 57275 -690 57305 -660
rect 57925 2015 57955 2045
rect 57965 2015 57995 2045
rect 58005 2015 58035 2045
rect 57925 1975 57955 2005
rect 57965 1975 57995 2005
rect 58005 1975 58035 2005
rect 57925 1935 57955 1965
rect 57965 1935 57995 1965
rect 58005 1935 58035 1965
rect 57925 1770 57955 1800
rect 57965 1770 57995 1800
rect 58005 1770 58035 1800
rect 57925 1730 57955 1760
rect 57965 1730 57995 1760
rect 58005 1730 58035 1760
rect 57925 1690 57955 1720
rect 57965 1690 57995 1720
rect 58005 1690 58035 1720
rect 57925 1360 57955 1390
rect 57965 1360 57995 1390
rect 58005 1360 58035 1390
rect 57925 1320 57955 1350
rect 57965 1320 57995 1350
rect 58005 1320 58035 1350
rect 57925 1280 57955 1310
rect 57965 1280 57995 1310
rect 58005 1280 58035 1310
rect 58105 1905 58135 1935
rect 58145 1905 58175 1935
rect 58185 1905 58215 1935
rect 58105 1865 58135 1895
rect 58145 1865 58175 1895
rect 58185 1865 58215 1895
rect 58105 1825 58135 1855
rect 58145 1825 58175 1855
rect 58185 1825 58215 1855
rect 57925 1205 57955 1235
rect 57965 1205 57995 1235
rect 58005 1205 58035 1235
rect 57925 1165 57955 1195
rect 57965 1165 57995 1195
rect 58005 1165 58035 1195
rect 57925 1125 57955 1155
rect 57965 1125 57995 1155
rect 58005 1125 58035 1155
rect 57870 -70 57900 -40
rect 58245 3210 58275 3240
rect 58285 3210 58315 3240
rect 58325 3210 58355 3240
rect 58245 3170 58275 3200
rect 58285 3170 58315 3200
rect 58325 3170 58355 3200
rect 58245 3130 58275 3160
rect 58285 3130 58315 3160
rect 58325 3130 58355 3160
rect 58445 3075 58475 3105
rect 58445 3035 58475 3065
rect 58445 2995 58475 3025
rect 58555 3075 58585 3105
rect 58555 3035 58585 3065
rect 58555 2995 58585 3025
rect 58665 3075 58695 3105
rect 58665 3035 58695 3065
rect 58665 2995 58695 3025
rect 58775 3075 58805 3105
rect 58775 3035 58805 3065
rect 58775 2995 58805 3025
rect 58885 3075 58915 3105
rect 58885 3035 58915 3065
rect 58885 2995 58915 3025
rect 58995 3075 59025 3105
rect 58995 3035 59025 3065
rect 58995 2995 59025 3025
rect 59105 3075 59135 3105
rect 59860 3095 59890 3125
rect 59105 3035 59135 3065
rect 59105 2995 59135 3025
rect 58500 2910 58530 2940
rect 58610 2910 58640 2940
rect 58720 2910 58750 2940
rect 58830 2910 58860 2940
rect 58940 2910 58970 2940
rect 59050 2910 59080 2940
rect 58245 2190 58275 2220
rect 58285 2190 58315 2220
rect 58325 2190 58355 2220
rect 58245 2150 58275 2180
rect 58285 2150 58315 2180
rect 58325 2150 58355 2180
rect 58245 2110 58275 2140
rect 58285 2110 58315 2140
rect 58325 2110 58355 2140
rect 58500 2270 58530 2300
rect 58610 2270 58640 2300
rect 58720 2270 58750 2300
rect 58830 2270 58860 2300
rect 58775 2215 58805 2220
rect 58775 2195 58780 2215
rect 58780 2195 58800 2215
rect 58800 2195 58805 2215
rect 58775 2190 58805 2195
rect 58775 2175 58805 2180
rect 58775 2155 58780 2175
rect 58780 2155 58800 2175
rect 58800 2155 58805 2175
rect 58775 2150 58805 2155
rect 58775 2135 58805 2140
rect 58775 2115 58780 2135
rect 58780 2115 58800 2135
rect 58800 2115 58805 2135
rect 58775 2110 58805 2115
rect 58940 2270 58970 2300
rect 59050 2270 59080 2300
rect 59820 2190 59850 2220
rect 59860 2190 59890 2220
rect 59900 2190 59930 2220
rect 59820 2150 59850 2180
rect 59860 2150 59890 2180
rect 59900 2150 59930 2180
rect 59820 2110 59850 2140
rect 59860 2110 59890 2140
rect 59900 2110 59930 2140
rect 58500 2040 58530 2070
rect 58555 2040 58585 2070
rect 58610 2040 58640 2070
rect 58665 2040 58695 2070
rect 58720 2040 58750 2070
rect 58775 2040 58805 2070
rect 58830 2040 58860 2070
rect 58885 2040 58915 2070
rect 58940 2040 58970 2070
rect 58995 2040 59025 2070
rect 59050 2040 59080 2070
rect 58500 2000 58530 2030
rect 58555 2000 58585 2030
rect 58610 2000 58640 2030
rect 58665 2000 58695 2030
rect 58720 2000 58750 2030
rect 58775 2000 58805 2030
rect 58830 2000 58860 2030
rect 58885 2000 58915 2030
rect 58940 2000 58970 2030
rect 58995 2000 59025 2030
rect 59050 2000 59080 2030
rect 58500 1960 58530 1990
rect 58555 1960 58585 1990
rect 58610 1960 58640 1990
rect 58665 1960 58695 1990
rect 58720 1960 58750 1990
rect 58775 1960 58805 1990
rect 58830 1960 58860 1990
rect 58885 1960 58915 1990
rect 58940 1960 58970 1990
rect 58995 1960 59025 1990
rect 59050 1960 59080 1990
rect 59720 2040 59750 2070
rect 59760 2040 59790 2070
rect 59805 2040 59835 2070
rect 59845 2040 59875 2070
rect 59890 2040 59920 2070
rect 59930 2040 59960 2070
rect 59720 2000 59750 2030
rect 59760 2000 59790 2030
rect 59805 2000 59835 2030
rect 59845 2000 59875 2030
rect 59890 2000 59920 2030
rect 59930 2000 59960 2030
rect 59720 1960 59750 1990
rect 59760 1960 59790 1990
rect 59805 1960 59835 1990
rect 59845 1960 59875 1990
rect 59890 1960 59920 1990
rect 59930 1960 59960 1990
rect 58445 1905 58475 1935
rect 58445 1865 58475 1895
rect 58445 1825 58475 1855
rect 59105 1905 59135 1935
rect 59105 1865 59135 1895
rect 59105 1825 59135 1855
rect 58500 1770 58530 1800
rect 58500 1730 58530 1760
rect 58500 1690 58530 1720
rect 58610 1770 58640 1800
rect 58610 1730 58640 1760
rect 58610 1690 58640 1720
rect 58720 1770 58750 1800
rect 58720 1730 58750 1760
rect 58720 1690 58750 1720
rect 58830 1770 58860 1800
rect 58830 1730 58860 1760
rect 58830 1690 58860 1720
rect 58940 1770 58970 1800
rect 58940 1730 58970 1760
rect 58940 1690 58970 1720
rect 59050 1770 59080 1800
rect 59050 1730 59080 1760
rect 59050 1690 59080 1720
rect 58555 1635 58585 1665
rect 58665 1635 58695 1665
rect 58775 1635 58805 1665
rect 58885 1635 58915 1665
rect 58995 1635 59025 1665
rect 58555 1405 58585 1410
rect 58555 1385 58560 1405
rect 58560 1385 58580 1405
rect 58580 1385 58585 1405
rect 58555 1380 58585 1385
rect 58665 1405 58695 1410
rect 58665 1385 58670 1405
rect 58670 1385 58690 1405
rect 58690 1385 58695 1405
rect 58665 1380 58695 1385
rect 58775 1405 58805 1410
rect 58775 1385 58780 1405
rect 58780 1385 58800 1405
rect 58800 1385 58805 1405
rect 58775 1380 58805 1385
rect 58885 1405 58915 1410
rect 58885 1385 58890 1405
rect 58890 1385 58910 1405
rect 58910 1385 58915 1405
rect 58885 1380 58915 1385
rect 58995 1405 59025 1410
rect 58995 1385 59000 1405
rect 59000 1385 59020 1405
rect 59020 1385 59025 1405
rect 58995 1380 59025 1385
rect 59435 1380 59465 1410
rect 59725 1405 59755 1435
rect 59775 1405 59805 1435
rect 59825 1405 59855 1435
rect 59875 1405 59905 1435
rect 59925 1405 59955 1435
rect 58245 1315 58275 1345
rect 58285 1315 58315 1345
rect 58325 1315 58355 1345
rect 58245 1275 58275 1305
rect 58285 1275 58315 1305
rect 58325 1275 58355 1305
rect 58610 1340 58640 1345
rect 58610 1320 58615 1340
rect 58615 1320 58635 1340
rect 58635 1320 58640 1340
rect 58610 1315 58640 1320
rect 58610 1300 58640 1305
rect 58610 1280 58615 1300
rect 58615 1280 58635 1300
rect 58635 1280 58640 1300
rect 58610 1275 58640 1280
rect 58555 1195 58585 1225
rect 58665 1195 58695 1225
rect 58775 1195 58805 1225
rect 58885 1195 58915 1225
rect 58995 1195 59025 1225
rect 59200 1195 59230 1225
rect 58105 800 58135 830
rect 58145 800 58175 830
rect 58185 800 58215 830
rect 58105 760 58135 790
rect 58145 760 58175 790
rect 58185 760 58215 790
rect 58105 720 58135 750
rect 58145 720 58175 750
rect 58185 720 58215 750
rect 58555 855 58585 885
rect 58665 855 58695 885
rect 58775 855 58805 885
rect 58885 855 58915 885
rect 58995 855 59025 885
rect 59200 875 59230 905
rect 58500 800 58530 830
rect 58500 760 58530 790
rect 58500 720 58530 750
rect 58610 800 58640 830
rect 58610 760 58640 790
rect 58610 720 58640 750
rect 58720 800 58750 830
rect 58720 760 58750 790
rect 58720 720 58750 750
rect 58830 800 58860 830
rect 58830 760 58860 790
rect 58830 720 58860 750
rect 58940 800 58970 830
rect 58940 760 58970 790
rect 58940 720 58970 750
rect 59050 800 59080 830
rect 59050 760 59080 790
rect 59050 720 59080 750
rect 59725 1355 59755 1385
rect 59775 1355 59805 1385
rect 59825 1355 59855 1385
rect 59875 1355 59905 1385
rect 59925 1355 59955 1385
rect 59725 1305 59755 1335
rect 59775 1305 59805 1335
rect 59825 1305 59855 1335
rect 59875 1305 59905 1335
rect 59925 1305 59955 1335
rect 59475 905 59510 910
rect 59475 880 59480 905
rect 59480 880 59505 905
rect 59505 880 59510 905
rect 59475 875 59510 880
rect 59535 905 59570 910
rect 59535 880 59540 905
rect 59540 880 59565 905
rect 59565 880 59570 905
rect 59535 875 59570 880
rect 59595 905 59630 910
rect 59595 880 59600 905
rect 59600 880 59625 905
rect 59625 880 59630 905
rect 59595 875 59630 880
rect 59655 905 59690 910
rect 59655 880 59660 905
rect 59660 880 59685 905
rect 59685 880 59690 905
rect 59655 875 59690 880
rect 59435 805 59465 835
rect 59535 805 59565 835
rect 58445 660 58475 690
rect 58445 620 58475 650
rect 58445 580 58475 610
rect 59105 660 59135 690
rect 59105 620 59135 650
rect 59105 580 59135 610
rect 59655 525 59685 555
rect 58585 505 58615 510
rect 58585 485 58590 505
rect 58590 485 58610 505
rect 58610 485 58615 505
rect 58585 480 58615 485
rect 59520 480 59550 510
rect 58435 280 58465 310
rect 58475 280 58505 310
rect 58515 280 58545 310
rect 58555 280 58585 310
rect 58595 280 58625 310
rect 58635 280 58665 310
rect 58675 280 58705 310
rect 58715 280 58745 310
rect 58755 280 58785 310
rect 58795 280 58825 310
rect 58835 280 58865 310
rect 58435 240 58465 270
rect 58475 240 58505 270
rect 58515 240 58545 270
rect 58555 240 58585 270
rect 58595 240 58625 270
rect 58635 240 58665 270
rect 58675 240 58705 270
rect 58715 240 58745 270
rect 58755 240 58785 270
rect 58795 240 58825 270
rect 58835 240 58865 270
rect 58435 200 58465 230
rect 58475 200 58505 230
rect 58515 200 58545 230
rect 58555 200 58585 230
rect 58595 200 58625 230
rect 58635 200 58665 230
rect 58675 200 58705 230
rect 58715 200 58745 230
rect 58755 200 58785 230
rect 58795 200 58825 230
rect 58835 200 58865 230
rect 59455 280 59485 310
rect 59455 240 59485 270
rect 59455 200 59485 230
rect 57925 -125 57955 -95
rect 57965 -125 57995 -95
rect 58005 -125 58035 -95
rect 57925 -165 57955 -135
rect 57965 -165 57995 -135
rect 58005 -165 58035 -135
rect 57925 -205 57955 -175
rect 57965 -205 57995 -175
rect 58005 -205 58035 -175
rect 58435 -555 58465 -525
rect 58635 -555 58665 -525
rect 59720 280 59750 310
rect 59760 280 59790 310
rect 59805 280 59835 310
rect 59845 280 59875 310
rect 59890 280 59920 310
rect 59930 280 59960 310
rect 59720 240 59750 270
rect 59760 240 59790 270
rect 59805 240 59835 270
rect 59845 240 59875 270
rect 59890 240 59920 270
rect 59930 240 59960 270
rect 59720 200 59750 230
rect 59760 200 59790 230
rect 59805 200 59835 230
rect 59845 200 59875 230
rect 59890 200 59920 230
rect 59930 200 59960 230
rect 59995 1770 60025 1800
rect 60035 1770 60065 1800
rect 60075 1770 60105 1800
rect 59995 1730 60025 1760
rect 60035 1730 60065 1760
rect 60075 1730 60105 1760
rect 59995 1690 60025 1720
rect 60035 1690 60065 1720
rect 60075 1690 60105 1720
rect 59995 660 60025 690
rect 60035 660 60065 690
rect 60075 660 60105 690
rect 59995 620 60025 650
rect 60035 620 60065 650
rect 60075 620 60105 650
rect 59995 580 60025 610
rect 60035 580 60065 610
rect 60075 580 60105 610
rect 59455 170 59490 175
rect 59455 145 59460 170
rect 59460 145 59485 170
rect 59485 145 59490 170
rect 59455 140 59490 145
rect 59515 170 59550 175
rect 59515 145 59520 170
rect 59520 145 59545 170
rect 59545 145 59550 170
rect 59515 140 59550 145
rect 58835 -555 58865 -525
rect 57490 -610 57520 -580
rect 57490 -650 57520 -620
rect 57490 -690 57520 -660
rect 57545 -610 57575 -580
rect 57585 -610 57615 -580
rect 57625 -610 57655 -580
rect 57545 -650 57575 -620
rect 57585 -650 57615 -620
rect 57625 -650 57655 -620
rect 57545 -690 57575 -660
rect 57585 -690 57615 -660
rect 57625 -690 57655 -660
rect 57895 -610 57925 -580
rect 57935 -610 57965 -580
rect 57975 -610 58005 -580
rect 57895 -650 57925 -620
rect 57935 -650 57965 -620
rect 57975 -650 58005 -620
rect 57895 -690 57925 -660
rect 57935 -690 57965 -660
rect 57975 -690 58005 -660
rect 58245 -610 58275 -580
rect 58285 -610 58315 -580
rect 58325 -610 58355 -580
rect 58245 -650 58275 -620
rect 58285 -650 58315 -620
rect 58325 -650 58355 -620
rect 58245 -690 58275 -660
rect 58285 -690 58315 -660
rect 58325 -690 58355 -660
rect 58535 -610 58565 -580
rect 58535 -650 58565 -620
rect 58535 -690 58565 -660
rect 58595 -610 58625 -580
rect 58635 -610 58665 -580
rect 58675 -610 58705 -580
rect 58595 -650 58625 -620
rect 58635 -650 58665 -620
rect 58675 -650 58705 -620
rect 58595 -690 58625 -660
rect 58635 -690 58665 -660
rect 58675 -690 58705 -660
rect 58735 -610 58765 -580
rect 58735 -650 58765 -620
rect 58735 -690 58765 -660
rect 58945 -610 58975 -580
rect 58985 -610 59015 -580
rect 59025 -610 59055 -580
rect 58945 -650 58975 -620
rect 58985 -650 59015 -620
rect 59025 -650 59055 -620
rect 58945 -690 58975 -660
rect 58985 -690 59015 -660
rect 59025 -690 59055 -660
rect 59295 -610 59325 -580
rect 59335 -610 59365 -580
rect 59375 -610 59405 -580
rect 59295 -650 59325 -620
rect 59335 -650 59365 -620
rect 59375 -650 59405 -620
rect 59295 -690 59325 -660
rect 59335 -690 59365 -660
rect 59375 -690 59405 -660
rect 59645 -610 59675 -580
rect 59685 -610 59715 -580
rect 59725 -610 59755 -580
rect 59645 -650 59675 -620
rect 59685 -650 59715 -620
rect 59725 -650 59755 -620
rect 59645 -690 59675 -660
rect 59685 -690 59715 -660
rect 59725 -690 59755 -660
rect 59995 -610 60025 -580
rect 60035 -610 60065 -580
rect 60075 -610 60105 -580
rect 59995 -650 60025 -620
rect 60035 -650 60065 -620
rect 60075 -650 60105 -620
rect 59995 -690 60025 -660
rect 60035 -690 60065 -660
rect 60075 -690 60105 -660
rect 60345 -610 60375 -580
rect 60385 -610 60415 -580
rect 60425 -610 60455 -580
rect 60345 -650 60375 -620
rect 60385 -650 60415 -620
rect 60425 -650 60455 -620
rect 60345 -690 60375 -660
rect 60385 -690 60415 -660
rect 60425 -690 60455 -660
rect 60695 -610 60725 -580
rect 60735 -610 60765 -580
rect 60775 -610 60805 -580
rect 60695 -650 60725 -620
rect 60735 -650 60765 -620
rect 60775 -650 60805 -620
rect 60695 -690 60725 -660
rect 60735 -690 60765 -660
rect 60775 -690 60805 -660
rect 61045 -610 61075 -580
rect 61085 -610 61115 -580
rect 61125 -610 61155 -580
rect 61045 -650 61075 -620
rect 61085 -650 61115 -620
rect 61125 -650 61155 -620
rect 61045 -690 61075 -660
rect 61085 -690 61115 -660
rect 61125 -690 61155 -660
rect 61395 -610 61425 -580
rect 61435 -610 61465 -580
rect 61475 -610 61505 -580
rect 61395 -650 61425 -620
rect 61435 -650 61465 -620
rect 61475 -650 61505 -620
rect 61395 -690 61425 -660
rect 61435 -690 61465 -660
rect 61475 -690 61505 -660
<< metal2 >>
rect 56205 5065 56245 5070
rect 56205 5035 56210 5065
rect 56240 5060 56245 5065
rect 56675 5065 56715 5070
rect 56675 5060 56680 5065
rect 56240 5040 56680 5060
rect 56240 5035 56245 5040
rect 56205 5030 56245 5035
rect 56675 5035 56680 5040
rect 56710 5035 56715 5065
rect 56675 5030 56715 5035
rect 57085 5065 57125 5070
rect 57085 5035 57090 5065
rect 57120 5060 57125 5065
rect 57555 5065 57595 5070
rect 57555 5060 57560 5065
rect 57120 5040 57560 5060
rect 57120 5035 57125 5040
rect 57085 5030 57125 5035
rect 57555 5035 57560 5040
rect 57590 5035 57595 5065
rect 57555 5030 57595 5035
rect 56880 5010 57245 5015
rect 56880 4980 56885 5010
rect 56915 4980 57030 5010
rect 57060 4980 57150 5010
rect 57180 4980 57210 5010
rect 57240 4980 57245 5010
rect 56880 4970 57245 4980
rect 56880 4940 56885 4970
rect 56915 4940 57030 4970
rect 57060 4940 57150 4970
rect 57180 4940 57210 4970
rect 57240 4940 57245 4970
rect 56085 4930 56125 4935
rect 56085 4900 56090 4930
rect 56120 4925 56125 4930
rect 56205 4930 56245 4935
rect 56205 4925 56210 4930
rect 56120 4905 56210 4925
rect 56120 4900 56125 4905
rect 56085 4895 56125 4900
rect 56205 4900 56210 4905
rect 56240 4925 56245 4930
rect 56265 4930 56305 4935
rect 56265 4925 56270 4930
rect 56240 4905 56270 4925
rect 56240 4900 56245 4905
rect 56205 4895 56245 4900
rect 56265 4900 56270 4905
rect 56300 4900 56305 4930
rect 56265 4895 56305 4900
rect 56880 4930 57245 4940
rect 56880 4900 56885 4930
rect 56915 4900 57030 4930
rect 57060 4900 57150 4930
rect 57180 4900 57210 4930
rect 57240 4900 57245 4930
rect 56880 4895 57245 4900
rect 57495 4930 57535 4935
rect 57495 4900 57500 4930
rect 57530 4925 57535 4930
rect 57555 4930 57595 4935
rect 57555 4925 57560 4930
rect 57530 4905 57560 4925
rect 57530 4900 57535 4905
rect 57495 4895 57535 4900
rect 57555 4900 57560 4905
rect 57590 4925 57595 4930
rect 57675 4930 57715 4935
rect 57675 4925 57680 4930
rect 57590 4905 57680 4925
rect 57590 4900 57595 4905
rect 57555 4895 57595 4900
rect 57675 4900 57680 4905
rect 57710 4900 57715 4930
rect 57675 4895 57715 4900
rect 56555 4840 56920 4845
rect 56555 4810 56560 4840
rect 56590 4810 56620 4840
rect 56650 4810 56740 4840
rect 56770 4810 56885 4840
rect 56915 4810 56920 4840
rect 56555 4800 56920 4810
rect 56555 4770 56560 4800
rect 56590 4770 56620 4800
rect 56650 4770 56740 4800
rect 56770 4770 56885 4800
rect 56915 4770 56920 4800
rect 56555 4760 56920 4770
rect 56555 4730 56560 4760
rect 56590 4730 56620 4760
rect 56650 4730 56740 4760
rect 56770 4730 56885 4760
rect 56915 4730 56920 4760
rect 56555 4725 56920 4730
rect 56205 4525 56245 4530
rect 56205 4495 56210 4525
rect 56240 4520 56245 4525
rect 56675 4525 56715 4530
rect 56675 4520 56680 4525
rect 56240 4500 56680 4520
rect 56240 4495 56245 4500
rect 56205 4490 56245 4495
rect 56675 4495 56680 4500
rect 56710 4495 56715 4525
rect 56675 4490 56715 4495
rect 57085 4525 57125 4530
rect 57085 4495 57090 4525
rect 57120 4520 57125 4525
rect 57555 4525 57595 4530
rect 57555 4520 57560 4525
rect 57120 4500 57560 4520
rect 57120 4495 57125 4500
rect 57085 4490 57125 4495
rect 57555 4495 57560 4500
rect 57590 4495 57595 4525
rect 57555 4490 57595 4495
rect 56150 4480 56190 4485
rect 56150 4450 56155 4480
rect 56185 4475 56190 4480
rect 56630 4480 56660 4485
rect 56185 4455 56630 4475
rect 56185 4450 56190 4455
rect 56150 4445 56190 4450
rect 56825 4480 56865 4485
rect 56825 4475 56830 4480
rect 56660 4455 56830 4475
rect 56630 4445 56660 4450
rect 56825 4450 56830 4455
rect 56860 4475 56865 4480
rect 56860 4470 57606 4475
rect 56860 4455 57576 4470
rect 56860 4450 56865 4455
rect 56825 4445 56865 4450
rect 57576 4435 57606 4440
rect 56935 4425 56975 4430
rect 56935 4395 56940 4425
rect 56970 4410 56975 4425
rect 57135 4415 57175 4420
rect 57135 4410 57140 4415
rect 56970 4395 57140 4410
rect 56935 4390 57140 4395
rect 57135 4385 57140 4390
rect 57170 4410 57175 4415
rect 57615 4415 57655 4420
rect 57615 4410 57620 4415
rect 57170 4390 57620 4410
rect 57170 4385 57175 4390
rect 57135 4380 57175 4385
rect 57615 4385 57620 4390
rect 57650 4385 57655 4415
rect 57615 4380 57655 4385
rect 52290 4320 61510 4325
rect 52290 4290 52295 4320
rect 52325 4290 52335 4320
rect 52365 4290 52375 4320
rect 52405 4290 52645 4320
rect 52675 4290 52685 4320
rect 52715 4290 52725 4320
rect 52755 4290 52995 4320
rect 53025 4290 53035 4320
rect 53065 4290 53075 4320
rect 53105 4290 53965 4320
rect 53995 4290 54005 4320
rect 54035 4290 54045 4320
rect 54075 4290 54315 4320
rect 54345 4290 54355 4320
rect 54385 4290 54395 4320
rect 54425 4290 54845 4320
rect 54875 4290 55205 4320
rect 55235 4290 55565 4320
rect 55595 4290 55665 4320
rect 55695 4290 55705 4320
rect 55735 4290 55745 4320
rect 55775 4290 56885 4320
rect 56915 4290 58105 4320
rect 58135 4290 58145 4320
rect 58175 4290 58185 4320
rect 58215 4290 58415 4320
rect 58445 4290 58775 4320
rect 58805 4290 59135 4320
rect 59165 4290 59645 4320
rect 59675 4290 59685 4320
rect 59715 4290 59725 4320
rect 59755 4290 59995 4320
rect 60025 4290 60035 4320
rect 60065 4290 60075 4320
rect 60105 4290 60695 4320
rect 60725 4290 60735 4320
rect 60765 4290 60775 4320
rect 60805 4290 61045 4320
rect 61075 4290 61085 4320
rect 61115 4290 61125 4320
rect 61155 4290 61395 4320
rect 61425 4290 61435 4320
rect 61465 4290 61475 4320
rect 61505 4290 61510 4320
rect 52290 4280 61510 4290
rect 52290 4250 52295 4280
rect 52325 4250 52335 4280
rect 52365 4250 52375 4280
rect 52405 4250 52645 4280
rect 52675 4250 52685 4280
rect 52715 4250 52725 4280
rect 52755 4250 52995 4280
rect 53025 4250 53035 4280
rect 53065 4250 53075 4280
rect 53105 4250 53965 4280
rect 53995 4250 54005 4280
rect 54035 4250 54045 4280
rect 54075 4250 54315 4280
rect 54345 4250 54355 4280
rect 54385 4250 54395 4280
rect 54425 4250 54845 4280
rect 54875 4250 55205 4280
rect 55235 4250 55565 4280
rect 55595 4250 55665 4280
rect 55695 4250 55705 4280
rect 55735 4250 55745 4280
rect 55775 4250 56885 4280
rect 56915 4250 58105 4280
rect 58135 4250 58145 4280
rect 58175 4250 58185 4280
rect 58215 4250 58415 4280
rect 58445 4250 58775 4280
rect 58805 4250 59135 4280
rect 59165 4250 59645 4280
rect 59675 4250 59685 4280
rect 59715 4250 59725 4280
rect 59755 4250 59995 4280
rect 60025 4250 60035 4280
rect 60065 4250 60075 4280
rect 60105 4250 60695 4280
rect 60725 4250 60735 4280
rect 60765 4250 60775 4280
rect 60805 4250 61045 4280
rect 61075 4250 61085 4280
rect 61115 4250 61125 4280
rect 61155 4250 61395 4280
rect 61425 4250 61435 4280
rect 61465 4250 61475 4280
rect 61505 4250 61510 4280
rect 52290 4240 61510 4250
rect 52290 4210 52295 4240
rect 52325 4210 52335 4240
rect 52365 4210 52375 4240
rect 52405 4210 52645 4240
rect 52675 4210 52685 4240
rect 52715 4210 52725 4240
rect 52755 4210 52995 4240
rect 53025 4210 53035 4240
rect 53065 4210 53075 4240
rect 53105 4210 53965 4240
rect 53995 4210 54005 4240
rect 54035 4210 54045 4240
rect 54075 4210 54315 4240
rect 54345 4210 54355 4240
rect 54385 4210 54395 4240
rect 54425 4210 54845 4240
rect 54875 4210 55205 4240
rect 55235 4210 55565 4240
rect 55595 4210 55665 4240
rect 55695 4210 55705 4240
rect 55735 4210 55745 4240
rect 55775 4210 56885 4240
rect 56915 4210 58105 4240
rect 58135 4210 58145 4240
rect 58175 4210 58185 4240
rect 58215 4210 58415 4240
rect 58445 4210 58775 4240
rect 58805 4210 59135 4240
rect 59165 4210 59645 4240
rect 59675 4210 59685 4240
rect 59715 4210 59725 4240
rect 59755 4210 59995 4240
rect 60025 4210 60035 4240
rect 60065 4210 60075 4240
rect 60105 4210 60695 4240
rect 60725 4210 60735 4240
rect 60765 4210 60775 4240
rect 60805 4210 61045 4240
rect 61075 4210 61085 4240
rect 61115 4210 61125 4240
rect 61155 4210 61395 4240
rect 61425 4210 61435 4240
rect 61465 4210 61475 4240
rect 61505 4210 61510 4240
rect 52290 4205 61510 4210
rect 54900 3935 56765 3940
rect 54900 3905 54905 3935
rect 54935 3905 54945 3935
rect 54975 3905 54985 3935
rect 55015 3905 55025 3935
rect 55055 3905 55065 3935
rect 55095 3905 55105 3935
rect 55135 3905 55145 3935
rect 55175 3905 55265 3935
rect 55295 3905 55305 3935
rect 55335 3905 55345 3935
rect 55375 3905 55385 3935
rect 55415 3905 55425 3935
rect 55455 3905 55465 3935
rect 55495 3905 55505 3935
rect 55535 3905 56010 3935
rect 56040 3905 56050 3935
rect 56080 3905 56090 3935
rect 56120 3905 56130 3935
rect 56160 3905 56170 3935
rect 56200 3905 56210 3935
rect 56240 3905 56250 3935
rect 56280 3905 56290 3935
rect 56320 3905 56330 3935
rect 56360 3905 56370 3935
rect 56400 3905 56410 3935
rect 56440 3905 56450 3935
rect 56480 3905 56490 3935
rect 56520 3905 56530 3935
rect 56560 3905 56570 3935
rect 56600 3905 56610 3935
rect 56640 3905 56650 3935
rect 56680 3905 56690 3935
rect 56720 3905 56730 3935
rect 56760 3905 56765 3935
rect 54900 3895 56765 3905
rect 54900 3865 54905 3895
rect 54935 3865 54945 3895
rect 54975 3865 54985 3895
rect 55015 3865 55025 3895
rect 55055 3865 55065 3895
rect 55095 3865 55105 3895
rect 55135 3865 55145 3895
rect 55175 3865 55265 3895
rect 55295 3865 55305 3895
rect 55335 3865 55345 3895
rect 55375 3865 55385 3895
rect 55415 3865 55425 3895
rect 55455 3865 55465 3895
rect 55495 3865 55505 3895
rect 55535 3865 56010 3895
rect 56040 3865 56050 3895
rect 56080 3865 56090 3895
rect 56120 3865 56130 3895
rect 56160 3865 56170 3895
rect 56200 3865 56210 3895
rect 56240 3865 56250 3895
rect 56280 3865 56290 3895
rect 56320 3865 56330 3895
rect 56360 3865 56370 3895
rect 56400 3865 56410 3895
rect 56440 3865 56450 3895
rect 56480 3865 56490 3895
rect 56520 3865 56530 3895
rect 56560 3865 56570 3895
rect 56600 3865 56610 3895
rect 56640 3865 56650 3895
rect 56680 3865 56690 3895
rect 56720 3865 56730 3895
rect 56760 3865 56765 3895
rect 54900 3855 56765 3865
rect 54900 3825 54905 3855
rect 54935 3825 54945 3855
rect 54975 3825 54985 3855
rect 55015 3825 55025 3855
rect 55055 3825 55065 3855
rect 55095 3825 55105 3855
rect 55135 3825 55145 3855
rect 55175 3825 55265 3855
rect 55295 3825 55305 3855
rect 55335 3825 55345 3855
rect 55375 3825 55385 3855
rect 55415 3825 55425 3855
rect 55455 3825 55465 3855
rect 55495 3825 55505 3855
rect 55535 3825 56010 3855
rect 56040 3825 56050 3855
rect 56080 3825 56090 3855
rect 56120 3825 56130 3855
rect 56160 3825 56170 3855
rect 56200 3825 56210 3855
rect 56240 3825 56250 3855
rect 56280 3825 56290 3855
rect 56320 3825 56330 3855
rect 56360 3825 56370 3855
rect 56400 3825 56410 3855
rect 56440 3825 56450 3855
rect 56480 3825 56490 3855
rect 56520 3825 56530 3855
rect 56560 3825 56570 3855
rect 56600 3825 56610 3855
rect 56640 3825 56650 3855
rect 56680 3825 56690 3855
rect 56720 3825 56730 3855
rect 56760 3825 56765 3855
rect 54900 3820 56765 3825
rect 57035 3935 59110 3940
rect 57035 3905 57040 3935
rect 57070 3905 57080 3935
rect 57110 3905 57120 3935
rect 57150 3905 57160 3935
rect 57190 3905 57200 3935
rect 57230 3905 57240 3935
rect 57270 3905 57280 3935
rect 57310 3905 57320 3935
rect 57350 3905 57360 3935
rect 57390 3905 57400 3935
rect 57430 3905 57440 3935
rect 57470 3905 57480 3935
rect 57510 3905 57520 3935
rect 57550 3905 57560 3935
rect 57590 3905 57600 3935
rect 57630 3905 57640 3935
rect 57670 3905 57680 3935
rect 57710 3905 57720 3935
rect 57750 3905 57760 3935
rect 57790 3905 58475 3935
rect 58505 3905 58515 3935
rect 58545 3905 58555 3935
rect 58585 3905 58595 3935
rect 58625 3905 58635 3935
rect 58665 3905 58675 3935
rect 58705 3905 58715 3935
rect 58745 3905 58835 3935
rect 58865 3905 58875 3935
rect 58905 3905 58915 3935
rect 58945 3905 58955 3935
rect 58985 3905 58995 3935
rect 59025 3905 59035 3935
rect 59065 3905 59075 3935
rect 59105 3905 59110 3935
rect 57035 3895 59110 3905
rect 57035 3865 57040 3895
rect 57070 3865 57080 3895
rect 57110 3865 57120 3895
rect 57150 3865 57160 3895
rect 57190 3865 57200 3895
rect 57230 3865 57240 3895
rect 57270 3865 57280 3895
rect 57310 3865 57320 3895
rect 57350 3865 57360 3895
rect 57390 3865 57400 3895
rect 57430 3865 57440 3895
rect 57470 3865 57480 3895
rect 57510 3865 57520 3895
rect 57550 3865 57560 3895
rect 57590 3865 57600 3895
rect 57630 3865 57640 3895
rect 57670 3865 57680 3895
rect 57710 3865 57720 3895
rect 57750 3865 57760 3895
rect 57790 3865 58475 3895
rect 58505 3865 58515 3895
rect 58545 3865 58555 3895
rect 58585 3865 58595 3895
rect 58625 3865 58635 3895
rect 58665 3865 58675 3895
rect 58705 3865 58715 3895
rect 58745 3865 58835 3895
rect 58865 3865 58875 3895
rect 58905 3865 58915 3895
rect 58945 3865 58955 3895
rect 58985 3865 58995 3895
rect 59025 3865 59035 3895
rect 59065 3865 59075 3895
rect 59105 3865 59110 3895
rect 57035 3855 59110 3865
rect 57035 3825 57040 3855
rect 57070 3825 57080 3855
rect 57110 3825 57120 3855
rect 57150 3825 57160 3855
rect 57190 3825 57200 3855
rect 57230 3825 57240 3855
rect 57270 3825 57280 3855
rect 57310 3825 57320 3855
rect 57350 3825 57360 3855
rect 57390 3825 57400 3855
rect 57430 3825 57440 3855
rect 57470 3825 57480 3855
rect 57510 3825 57520 3855
rect 57550 3825 57560 3855
rect 57590 3825 57600 3855
rect 57630 3825 57640 3855
rect 57670 3825 57680 3855
rect 57710 3825 57720 3855
rect 57750 3825 57760 3855
rect 57790 3825 58475 3855
rect 58505 3825 58515 3855
rect 58545 3825 58555 3855
rect 58585 3825 58595 3855
rect 58625 3825 58635 3855
rect 58665 3825 58675 3855
rect 58705 3825 58715 3855
rect 58745 3825 58835 3855
rect 58865 3825 58875 3855
rect 58905 3825 58915 3855
rect 58945 3825 58955 3855
rect 58985 3825 58995 3855
rect 59025 3825 59035 3855
rect 59065 3825 59075 3855
rect 59105 3825 59110 3855
rect 57035 3820 59110 3825
rect 54840 3800 54880 3805
rect 54840 3770 54845 3800
rect 54875 3795 54880 3800
rect 54960 3800 55000 3805
rect 54960 3795 54965 3800
rect 54875 3775 54965 3795
rect 54875 3770 54880 3775
rect 54840 3765 54880 3770
rect 54960 3770 54965 3775
rect 54995 3795 55000 3800
rect 55080 3800 55120 3805
rect 55080 3795 55085 3800
rect 54995 3775 55085 3795
rect 54995 3770 55000 3775
rect 54960 3765 55000 3770
rect 55080 3770 55085 3775
rect 55115 3795 55120 3800
rect 55200 3800 55240 3805
rect 55200 3795 55205 3800
rect 55115 3775 55205 3795
rect 55115 3770 55120 3775
rect 55080 3765 55120 3770
rect 55200 3770 55205 3775
rect 55235 3795 55240 3800
rect 55320 3800 55360 3805
rect 55320 3795 55325 3800
rect 55235 3775 55325 3795
rect 55235 3770 55240 3775
rect 55200 3765 55240 3770
rect 55320 3770 55325 3775
rect 55355 3795 55360 3800
rect 55440 3800 55480 3805
rect 55440 3795 55445 3800
rect 55355 3775 55445 3795
rect 55355 3770 55360 3775
rect 55320 3765 55360 3770
rect 55440 3770 55445 3775
rect 55475 3795 55480 3800
rect 55560 3800 55600 3805
rect 55560 3795 55565 3800
rect 55475 3775 55565 3795
rect 55475 3770 55480 3775
rect 55440 3765 55480 3770
rect 55560 3770 55565 3775
rect 55595 3770 55600 3800
rect 55560 3765 55600 3770
rect 56065 3800 56105 3805
rect 56065 3770 56070 3800
rect 56100 3795 56105 3800
rect 56185 3800 56225 3805
rect 56185 3795 56190 3800
rect 56100 3775 56190 3795
rect 56100 3770 56105 3775
rect 56065 3765 56105 3770
rect 56185 3770 56190 3775
rect 56220 3795 56225 3800
rect 56305 3800 56345 3805
rect 56305 3795 56310 3800
rect 56220 3775 56310 3795
rect 56220 3770 56225 3775
rect 56185 3765 56225 3770
rect 56305 3770 56310 3775
rect 56340 3795 56345 3800
rect 56425 3800 56465 3805
rect 56425 3795 56430 3800
rect 56340 3775 56430 3795
rect 56340 3770 56345 3775
rect 56305 3765 56345 3770
rect 56425 3770 56430 3775
rect 56460 3795 56465 3800
rect 56545 3800 56585 3805
rect 56545 3795 56550 3800
rect 56460 3775 56550 3795
rect 56460 3770 56465 3775
rect 56425 3765 56465 3770
rect 56545 3770 56550 3775
rect 56580 3795 56585 3800
rect 56665 3800 56705 3805
rect 56665 3795 56670 3800
rect 56580 3775 56670 3795
rect 56580 3770 56585 3775
rect 56545 3765 56585 3770
rect 56665 3770 56670 3775
rect 56700 3770 56705 3800
rect 56665 3765 56705 3770
rect 57095 3800 57135 3805
rect 57095 3770 57100 3800
rect 57130 3795 57135 3800
rect 57215 3800 57255 3805
rect 57215 3795 57220 3800
rect 57130 3775 57220 3795
rect 57130 3770 57135 3775
rect 57095 3765 57135 3770
rect 57215 3770 57220 3775
rect 57250 3795 57255 3800
rect 57335 3800 57375 3805
rect 57335 3795 57340 3800
rect 57250 3775 57340 3795
rect 57250 3770 57255 3775
rect 57215 3765 57255 3770
rect 57335 3770 57340 3775
rect 57370 3795 57375 3800
rect 57455 3800 57495 3805
rect 57455 3795 57460 3800
rect 57370 3775 57460 3795
rect 57370 3770 57375 3775
rect 57335 3765 57375 3770
rect 57455 3770 57460 3775
rect 57490 3795 57495 3800
rect 57575 3800 57615 3805
rect 57575 3795 57580 3800
rect 57490 3775 57580 3795
rect 57490 3770 57495 3775
rect 57455 3765 57495 3770
rect 57575 3770 57580 3775
rect 57610 3795 57615 3800
rect 57695 3800 57735 3805
rect 57695 3795 57700 3800
rect 57610 3775 57700 3795
rect 57610 3770 57615 3775
rect 57575 3765 57615 3770
rect 57695 3770 57700 3775
rect 57730 3770 57735 3800
rect 57695 3765 57735 3770
rect 58410 3800 58450 3805
rect 58410 3770 58415 3800
rect 58445 3795 58450 3800
rect 58530 3800 58570 3805
rect 58530 3795 58535 3800
rect 58445 3775 58535 3795
rect 58445 3770 58450 3775
rect 58410 3765 58450 3770
rect 58530 3770 58535 3775
rect 58565 3795 58570 3800
rect 58650 3800 58690 3805
rect 58650 3795 58655 3800
rect 58565 3775 58655 3795
rect 58565 3770 58570 3775
rect 58530 3765 58570 3770
rect 58650 3770 58655 3775
rect 58685 3795 58690 3800
rect 58770 3800 58810 3805
rect 58770 3795 58775 3800
rect 58685 3775 58775 3795
rect 58685 3770 58690 3775
rect 58650 3765 58690 3770
rect 58770 3770 58775 3775
rect 58805 3795 58810 3800
rect 58890 3800 58930 3805
rect 58890 3795 58895 3800
rect 58805 3775 58895 3795
rect 58805 3770 58810 3775
rect 58770 3765 58810 3770
rect 58890 3770 58895 3775
rect 58925 3795 58930 3800
rect 59010 3800 59050 3805
rect 59010 3795 59015 3800
rect 58925 3775 59015 3795
rect 58925 3770 58930 3775
rect 58890 3765 58930 3770
rect 59010 3770 59015 3775
rect 59045 3795 59050 3800
rect 59130 3800 59170 3805
rect 59130 3795 59135 3800
rect 59045 3775 59135 3795
rect 59045 3770 59050 3775
rect 59010 3765 59050 3770
rect 59130 3770 59135 3775
rect 59165 3770 59170 3800
rect 59130 3765 59170 3770
rect 54900 3410 54940 3415
rect 54900 3380 54905 3410
rect 54935 3405 54940 3410
rect 55020 3410 55060 3415
rect 55020 3405 55025 3410
rect 54935 3385 55025 3405
rect 54935 3380 54940 3385
rect 54900 3375 54940 3380
rect 55020 3380 55025 3385
rect 55055 3405 55060 3410
rect 55140 3410 55180 3415
rect 55140 3405 55145 3410
rect 55055 3385 55145 3405
rect 55055 3380 55060 3385
rect 55020 3375 55060 3380
rect 55140 3380 55145 3385
rect 55175 3405 55180 3410
rect 55260 3410 55300 3415
rect 55260 3405 55265 3410
rect 55175 3385 55265 3405
rect 55175 3380 55180 3385
rect 55140 3375 55180 3380
rect 55260 3380 55265 3385
rect 55295 3405 55300 3410
rect 55380 3410 55420 3415
rect 55380 3405 55385 3410
rect 55295 3385 55385 3405
rect 55295 3380 55300 3385
rect 55260 3375 55300 3380
rect 55380 3380 55385 3385
rect 55415 3405 55420 3410
rect 55500 3410 55540 3415
rect 55500 3405 55505 3410
rect 55415 3385 55505 3405
rect 55415 3380 55420 3385
rect 55380 3375 55420 3380
rect 55500 3380 55505 3385
rect 55535 3380 55540 3410
rect 55500 3375 55540 3380
rect 56065 3410 56105 3415
rect 56065 3380 56070 3410
rect 56100 3405 56105 3410
rect 56185 3410 56225 3415
rect 56185 3405 56190 3410
rect 56100 3385 56190 3405
rect 56100 3380 56105 3385
rect 56065 3375 56105 3380
rect 56185 3380 56190 3385
rect 56220 3405 56225 3410
rect 56305 3410 56345 3415
rect 56305 3405 56310 3410
rect 56220 3385 56310 3405
rect 56220 3380 56225 3385
rect 56185 3375 56225 3380
rect 56305 3380 56310 3385
rect 56340 3405 56345 3410
rect 56425 3410 56465 3415
rect 56425 3405 56430 3410
rect 56340 3385 56430 3405
rect 56340 3380 56345 3385
rect 56305 3375 56345 3380
rect 56425 3380 56430 3385
rect 56460 3405 56465 3410
rect 56545 3410 56585 3415
rect 56545 3405 56550 3410
rect 56460 3385 56550 3405
rect 56460 3380 56465 3385
rect 56425 3375 56465 3380
rect 56545 3380 56550 3385
rect 56580 3405 56585 3410
rect 56665 3410 56705 3415
rect 56665 3405 56670 3410
rect 56580 3385 56670 3405
rect 56580 3380 56585 3385
rect 56545 3375 56585 3380
rect 56665 3380 56670 3385
rect 56700 3380 56705 3410
rect 56665 3375 56705 3380
rect 57095 3410 57135 3415
rect 57095 3380 57100 3410
rect 57130 3405 57135 3410
rect 57215 3410 57255 3415
rect 57215 3405 57220 3410
rect 57130 3385 57220 3405
rect 57130 3380 57135 3385
rect 57095 3375 57135 3380
rect 57215 3380 57220 3385
rect 57250 3405 57255 3410
rect 57335 3410 57375 3415
rect 57335 3405 57340 3410
rect 57250 3385 57340 3405
rect 57250 3380 57255 3385
rect 57215 3375 57255 3380
rect 57335 3380 57340 3385
rect 57370 3405 57375 3410
rect 57455 3410 57495 3415
rect 57455 3405 57460 3410
rect 57370 3385 57460 3405
rect 57370 3380 57375 3385
rect 57335 3375 57375 3380
rect 57455 3380 57460 3385
rect 57490 3405 57495 3410
rect 57575 3410 57615 3415
rect 57575 3405 57580 3410
rect 57490 3385 57580 3405
rect 57490 3380 57495 3385
rect 57455 3375 57495 3380
rect 57575 3380 57580 3385
rect 57610 3405 57615 3410
rect 57695 3410 57735 3415
rect 57695 3405 57700 3410
rect 57610 3385 57700 3405
rect 57610 3380 57615 3385
rect 57575 3375 57615 3380
rect 57695 3380 57700 3385
rect 57730 3380 57735 3410
rect 57695 3375 57735 3380
rect 58470 3410 58510 3415
rect 58470 3380 58475 3410
rect 58505 3405 58510 3410
rect 58590 3410 58630 3415
rect 58590 3405 58595 3410
rect 58505 3385 58595 3405
rect 58505 3380 58510 3385
rect 58470 3375 58510 3380
rect 58590 3380 58595 3385
rect 58625 3405 58630 3410
rect 58710 3410 58750 3415
rect 58710 3405 58715 3410
rect 58625 3385 58715 3405
rect 58625 3380 58630 3385
rect 58590 3375 58630 3380
rect 58710 3380 58715 3385
rect 58745 3405 58750 3410
rect 58830 3410 58870 3415
rect 58830 3405 58835 3410
rect 58745 3385 58835 3405
rect 58745 3380 58750 3385
rect 58710 3375 58750 3380
rect 58830 3380 58835 3385
rect 58865 3405 58870 3410
rect 58950 3410 58990 3415
rect 58950 3405 58955 3410
rect 58865 3385 58955 3405
rect 58865 3380 58870 3385
rect 58830 3375 58870 3380
rect 58950 3380 58955 3385
rect 58985 3405 58990 3410
rect 59070 3410 59110 3415
rect 59070 3405 59075 3410
rect 58985 3385 59075 3405
rect 58985 3380 58990 3385
rect 58950 3375 58990 3380
rect 59070 3380 59075 3385
rect 59105 3380 59110 3410
rect 59070 3375 59110 3380
rect 56365 3330 56405 3335
rect 56365 3300 56370 3330
rect 56400 3325 56405 3330
rect 56835 3330 56875 3335
rect 56835 3325 56840 3330
rect 56400 3305 56840 3325
rect 56400 3300 56405 3305
rect 56365 3295 56405 3300
rect 56835 3300 56840 3305
rect 56870 3325 56875 3330
rect 57395 3330 57435 3335
rect 57395 3325 57400 3330
rect 56870 3305 57400 3325
rect 56870 3300 56875 3305
rect 56835 3295 56875 3300
rect 57395 3300 57400 3305
rect 57430 3300 57435 3330
rect 57395 3295 57435 3300
rect 55200 3285 55240 3290
rect 55200 3255 55205 3285
rect 55235 3280 55240 3285
rect 56925 3285 56965 3290
rect 56925 3280 56930 3285
rect 55235 3260 56930 3280
rect 55235 3255 55240 3260
rect 55200 3250 55240 3255
rect 56925 3255 56930 3260
rect 56960 3280 56965 3285
rect 58770 3285 58810 3290
rect 58770 3280 58775 3285
rect 56960 3260 58775 3280
rect 56960 3255 56965 3260
rect 56925 3250 56965 3255
rect 58770 3255 58775 3260
rect 58805 3255 58810 3285
rect 58770 3250 58810 3255
rect 55520 3240 56705 3245
rect 55520 3210 55525 3240
rect 55555 3210 55565 3240
rect 55595 3210 55605 3240
rect 55635 3210 56070 3240
rect 56100 3210 56110 3240
rect 56140 3210 56150 3240
rect 56180 3210 56190 3240
rect 56220 3210 56230 3240
rect 56260 3210 56270 3240
rect 56300 3210 56310 3240
rect 56340 3210 56350 3240
rect 56380 3210 56390 3240
rect 56420 3210 56430 3240
rect 56460 3210 56470 3240
rect 56500 3210 56510 3240
rect 56540 3210 56550 3240
rect 56580 3210 56590 3240
rect 56620 3210 56630 3240
rect 56660 3210 56670 3240
rect 56700 3210 56705 3240
rect 55520 3200 56705 3210
rect 55520 3170 55525 3200
rect 55555 3170 55565 3200
rect 55595 3170 55605 3200
rect 55635 3170 56070 3200
rect 56100 3170 56110 3200
rect 56140 3170 56150 3200
rect 56180 3170 56190 3200
rect 56220 3170 56230 3200
rect 56260 3170 56270 3200
rect 56300 3170 56310 3200
rect 56340 3170 56350 3200
rect 56380 3170 56390 3200
rect 56420 3170 56430 3200
rect 56460 3170 56470 3200
rect 56500 3170 56510 3200
rect 56540 3170 56550 3200
rect 56580 3170 56590 3200
rect 56620 3170 56630 3200
rect 56660 3170 56670 3200
rect 56700 3170 56705 3200
rect 55520 3160 56705 3170
rect 55520 3130 55525 3160
rect 55555 3130 55565 3160
rect 55595 3130 55605 3160
rect 55635 3130 56070 3160
rect 56100 3130 56110 3160
rect 56140 3130 56150 3160
rect 56180 3130 56190 3160
rect 56220 3130 56230 3160
rect 56260 3130 56270 3160
rect 56300 3130 56310 3160
rect 56340 3130 56350 3160
rect 56380 3130 56390 3160
rect 56420 3130 56430 3160
rect 56460 3130 56470 3160
rect 56500 3130 56510 3160
rect 56540 3130 56550 3160
rect 56580 3130 56590 3160
rect 56620 3130 56630 3160
rect 56660 3130 56670 3160
rect 56700 3130 56705 3160
rect 54175 3125 54215 3130
rect 55520 3125 56705 3130
rect 57095 3240 58360 3245
rect 57095 3210 57100 3240
rect 57130 3210 57140 3240
rect 57170 3210 57180 3240
rect 57210 3210 57220 3240
rect 57250 3210 57260 3240
rect 57290 3210 57300 3240
rect 57330 3210 57340 3240
rect 57370 3210 57380 3240
rect 57410 3210 57420 3240
rect 57450 3210 57460 3240
rect 57490 3210 57500 3240
rect 57530 3210 57540 3240
rect 57570 3210 57580 3240
rect 57610 3210 57620 3240
rect 57650 3210 57660 3240
rect 57690 3210 57700 3240
rect 57730 3210 58245 3240
rect 58275 3210 58285 3240
rect 58315 3210 58325 3240
rect 58355 3210 58360 3240
rect 57095 3200 58360 3210
rect 57095 3170 57100 3200
rect 57130 3170 57140 3200
rect 57170 3170 57180 3200
rect 57210 3170 57220 3200
rect 57250 3170 57260 3200
rect 57290 3170 57300 3200
rect 57330 3170 57340 3200
rect 57370 3170 57380 3200
rect 57410 3170 57420 3200
rect 57450 3170 57460 3200
rect 57490 3170 57500 3200
rect 57530 3170 57540 3200
rect 57570 3170 57580 3200
rect 57610 3170 57620 3200
rect 57650 3170 57660 3200
rect 57690 3170 57700 3200
rect 57730 3170 58245 3200
rect 58275 3170 58285 3200
rect 58315 3170 58325 3200
rect 58355 3170 58360 3200
rect 57095 3160 58360 3170
rect 57095 3130 57100 3160
rect 57130 3130 57140 3160
rect 57170 3130 57180 3160
rect 57210 3130 57220 3160
rect 57250 3130 57260 3160
rect 57290 3130 57300 3160
rect 57330 3130 57340 3160
rect 57370 3130 57380 3160
rect 57410 3130 57420 3160
rect 57450 3130 57460 3160
rect 57490 3130 57500 3160
rect 57530 3130 57540 3160
rect 57570 3130 57580 3160
rect 57610 3130 57620 3160
rect 57650 3130 57660 3160
rect 57690 3130 57700 3160
rect 57730 3130 58245 3160
rect 58275 3130 58285 3160
rect 58315 3130 58325 3160
rect 58355 3130 58360 3160
rect 57095 3125 58360 3130
rect 59855 3125 59895 3130
rect 54175 3095 54180 3125
rect 54210 3095 54215 3125
rect 54175 3090 54215 3095
rect 54740 3105 55780 3110
rect 54740 3075 54745 3105
rect 54775 3075 54855 3105
rect 54885 3075 54965 3105
rect 54995 3075 55075 3105
rect 55105 3075 55185 3105
rect 55215 3075 55295 3105
rect 55325 3075 55405 3105
rect 55435 3075 55665 3105
rect 55695 3075 55705 3105
rect 55735 3075 55745 3105
rect 55775 3075 55780 3105
rect 57290 3105 59140 3110
rect 57290 3100 58105 3105
rect 54740 3065 55780 3075
rect 54740 3035 54745 3065
rect 54775 3035 54855 3065
rect 54885 3035 54965 3065
rect 54995 3035 55075 3065
rect 55105 3035 55185 3065
rect 55215 3035 55295 3065
rect 55325 3035 55405 3065
rect 55435 3035 55665 3065
rect 55695 3035 55705 3065
rect 55735 3035 55745 3065
rect 55775 3035 55780 3065
rect 54740 3025 55780 3035
rect 54740 2995 54745 3025
rect 54775 2995 54855 3025
rect 54885 2995 54965 3025
rect 54995 2995 55075 3025
rect 55105 2995 55185 3025
rect 55215 2995 55295 3025
rect 55325 2995 55405 3025
rect 55435 2995 55665 3025
rect 55695 2995 55705 3025
rect 55735 2995 55745 3025
rect 55775 2995 55780 3025
rect 54740 2990 55780 2995
rect 56510 3095 58105 3100
rect 56510 3065 56515 3095
rect 56545 3065 56680 3095
rect 56710 3065 56845 3095
rect 56875 3065 56925 3095
rect 56955 3065 57090 3095
rect 57120 3065 57255 3095
rect 57285 3075 58105 3095
rect 58135 3075 58145 3105
rect 58175 3075 58185 3105
rect 58215 3075 58445 3105
rect 58475 3075 58555 3105
rect 58585 3075 58665 3105
rect 58695 3075 58775 3105
rect 58805 3075 58885 3105
rect 58915 3075 58995 3105
rect 59025 3075 59105 3105
rect 59135 3075 59140 3105
rect 59855 3095 59860 3125
rect 59890 3095 59895 3125
rect 59855 3090 59895 3095
rect 57285 3065 59140 3075
rect 56510 3055 58105 3065
rect 56510 3025 56515 3055
rect 56545 3025 56680 3055
rect 56710 3025 56845 3055
rect 56875 3025 56925 3055
rect 56955 3025 57090 3055
rect 57120 3025 57255 3055
rect 57285 3035 58105 3055
rect 58135 3035 58145 3065
rect 58175 3035 58185 3065
rect 58215 3035 58445 3065
rect 58475 3035 58555 3065
rect 58585 3035 58665 3065
rect 58695 3035 58775 3065
rect 58805 3035 58885 3065
rect 58915 3035 58995 3065
rect 59025 3035 59105 3065
rect 59135 3035 59140 3065
rect 57285 3025 59140 3035
rect 56510 3015 58105 3025
rect 56510 2985 56515 3015
rect 56545 2985 56680 3015
rect 56710 2985 56845 3015
rect 56875 2985 56925 3015
rect 56955 2985 57090 3015
rect 57120 2985 57255 3015
rect 57285 2995 58105 3015
rect 58135 2995 58145 3025
rect 58175 2995 58185 3025
rect 58215 2995 58445 3025
rect 58475 2995 58555 3025
rect 58585 2995 58665 3025
rect 58695 2995 58775 3025
rect 58805 2995 58885 3025
rect 58915 2995 58995 3025
rect 59025 2995 59105 3025
rect 59135 2995 59140 3025
rect 57285 2990 59140 2995
rect 57285 2985 57290 2990
rect 56510 2980 57290 2985
rect 56620 2960 56660 2965
rect 54795 2940 54835 2945
rect 54795 2910 54800 2940
rect 54830 2935 54835 2940
rect 54905 2940 54945 2945
rect 54905 2935 54910 2940
rect 54830 2915 54910 2935
rect 54830 2910 54835 2915
rect 54795 2905 54835 2910
rect 54905 2910 54910 2915
rect 54940 2935 54945 2940
rect 55015 2940 55055 2945
rect 55015 2935 55020 2940
rect 54940 2915 55020 2935
rect 54940 2910 54945 2915
rect 54905 2905 54945 2910
rect 55015 2910 55020 2915
rect 55050 2935 55055 2940
rect 55125 2940 55165 2945
rect 55125 2935 55130 2940
rect 55050 2915 55130 2935
rect 55050 2910 55055 2915
rect 55015 2905 55055 2910
rect 55125 2910 55130 2915
rect 55160 2935 55165 2940
rect 55235 2940 55275 2945
rect 55235 2935 55240 2940
rect 55160 2915 55240 2935
rect 55160 2910 55165 2915
rect 55125 2905 55165 2910
rect 55235 2910 55240 2915
rect 55270 2935 55275 2940
rect 55345 2940 55385 2945
rect 55345 2935 55350 2940
rect 55270 2915 55350 2935
rect 55270 2910 55275 2915
rect 55235 2905 55275 2910
rect 55345 2910 55350 2915
rect 55380 2910 55385 2940
rect 56620 2930 56625 2960
rect 56655 2955 56660 2960
rect 56730 2960 56770 2965
rect 56730 2955 56735 2960
rect 56655 2935 56735 2955
rect 56655 2930 56660 2935
rect 56620 2925 56660 2930
rect 56730 2930 56735 2935
rect 56765 2930 56770 2960
rect 56730 2925 56770 2930
rect 57030 2960 57070 2965
rect 57030 2930 57035 2960
rect 57065 2955 57070 2960
rect 57140 2960 57180 2965
rect 57140 2955 57145 2960
rect 57065 2935 57145 2955
rect 57065 2930 57070 2935
rect 57030 2925 57070 2930
rect 57140 2930 57145 2935
rect 57175 2930 57180 2960
rect 57140 2925 57180 2930
rect 58495 2940 58535 2945
rect 55345 2905 55385 2910
rect 58495 2910 58500 2940
rect 58530 2935 58535 2940
rect 58605 2940 58645 2945
rect 58605 2935 58610 2940
rect 58530 2915 58610 2935
rect 58530 2910 58535 2915
rect 58495 2905 58535 2910
rect 58605 2910 58610 2915
rect 58640 2935 58645 2940
rect 58715 2940 58755 2945
rect 58715 2935 58720 2940
rect 58640 2915 58720 2935
rect 58640 2910 58645 2915
rect 58605 2905 58645 2910
rect 58715 2910 58720 2915
rect 58750 2935 58755 2940
rect 58825 2940 58865 2945
rect 58825 2935 58830 2940
rect 58750 2915 58830 2935
rect 58750 2910 58755 2915
rect 58715 2905 58755 2910
rect 58825 2910 58830 2915
rect 58860 2935 58865 2940
rect 58935 2940 58975 2945
rect 58935 2935 58940 2940
rect 58860 2915 58940 2935
rect 58860 2910 58865 2915
rect 58825 2905 58865 2910
rect 58935 2910 58940 2915
rect 58970 2935 58975 2940
rect 59045 2940 59085 2945
rect 59045 2935 59050 2940
rect 58970 2915 59050 2935
rect 58970 2910 58975 2915
rect 58935 2905 58975 2910
rect 59045 2910 59050 2915
rect 59080 2910 59085 2940
rect 59045 2905 59085 2910
rect 56560 2650 56590 2655
rect 56800 2650 56830 2655
rect 56675 2640 56715 2645
rect 56675 2635 56680 2640
rect 56590 2620 56680 2635
rect 56560 2615 56680 2620
rect 56675 2610 56680 2615
rect 56710 2635 56715 2640
rect 56710 2620 56800 2635
rect 57085 2640 57125 2645
rect 57085 2635 57090 2640
rect 56830 2620 57090 2635
rect 56710 2615 57090 2620
rect 56710 2610 56715 2615
rect 56675 2605 56715 2610
rect 57085 2610 57090 2615
rect 57120 2635 57125 2640
rect 57120 2615 57130 2635
rect 57120 2610 57125 2615
rect 57085 2605 57125 2610
rect 56600 2580 56640 2585
rect 56600 2575 56605 2580
rect 56365 2555 56605 2575
rect 56600 2550 56605 2555
rect 56635 2575 56640 2580
rect 57160 2580 57200 2585
rect 57160 2575 57165 2580
rect 56635 2555 57165 2575
rect 56635 2550 56640 2555
rect 56600 2545 56640 2550
rect 57160 2550 57165 2555
rect 57195 2550 57200 2580
rect 57160 2545 57200 2550
rect 55940 2530 55980 2535
rect 55940 2500 55945 2530
rect 55975 2525 55980 2530
rect 56745 2530 56785 2535
rect 56745 2525 56750 2530
rect 55975 2505 56750 2525
rect 55975 2500 55980 2505
rect 55940 2495 55980 2500
rect 56745 2500 56750 2505
rect 56780 2525 56785 2530
rect 57015 2530 57055 2535
rect 57015 2525 57020 2530
rect 56780 2505 57020 2525
rect 56780 2500 56785 2505
rect 56745 2495 56785 2500
rect 57015 2500 57020 2505
rect 57050 2525 57055 2530
rect 57820 2530 57860 2535
rect 57820 2525 57825 2530
rect 57050 2505 57825 2525
rect 57050 2500 57055 2505
rect 57015 2495 57055 2500
rect 57820 2500 57825 2505
rect 57855 2500 57860 2530
rect 57820 2495 57860 2500
rect 56850 2475 56890 2480
rect 56850 2445 56855 2475
rect 56885 2470 56890 2475
rect 56960 2475 57000 2480
rect 56960 2470 56965 2475
rect 56885 2450 56965 2470
rect 56885 2445 56890 2450
rect 56850 2440 56890 2445
rect 56960 2445 56965 2450
rect 56995 2445 57000 2475
rect 56960 2440 57000 2445
rect 56935 2420 56975 2425
rect 56935 2390 56940 2420
rect 56970 2415 56975 2420
rect 57210 2420 57250 2425
rect 57210 2415 57215 2420
rect 56970 2395 57215 2415
rect 56970 2390 56975 2395
rect 56935 2385 56975 2390
rect 57210 2390 57215 2395
rect 57245 2415 57250 2420
rect 57865 2420 57905 2425
rect 57865 2415 57870 2420
rect 57245 2395 57870 2415
rect 57245 2390 57250 2395
rect 57210 2385 57250 2390
rect 57865 2390 57870 2395
rect 57900 2390 57905 2420
rect 57865 2385 57905 2390
rect 56850 2365 56890 2370
rect 56850 2335 56855 2365
rect 56885 2335 56890 2365
rect 56850 2330 56890 2335
rect 54795 2300 54835 2305
rect 54795 2270 54800 2300
rect 54830 2295 54835 2300
rect 54905 2300 54945 2305
rect 54905 2295 54910 2300
rect 54830 2275 54910 2295
rect 54830 2270 54835 2275
rect 54795 2265 54835 2270
rect 54905 2270 54910 2275
rect 54940 2295 54945 2300
rect 55015 2300 55055 2305
rect 55015 2295 55020 2300
rect 54940 2275 55020 2295
rect 54940 2270 54945 2275
rect 54905 2265 54945 2270
rect 55015 2270 55020 2275
rect 55050 2295 55055 2300
rect 55125 2300 55165 2305
rect 55125 2295 55130 2300
rect 55050 2275 55130 2295
rect 55050 2270 55055 2275
rect 55015 2265 55055 2270
rect 55125 2270 55130 2275
rect 55160 2295 55165 2300
rect 55235 2300 55275 2305
rect 55235 2295 55240 2300
rect 55160 2275 55240 2295
rect 55160 2270 55165 2275
rect 55125 2265 55165 2270
rect 55235 2270 55240 2275
rect 55270 2295 55275 2300
rect 55345 2300 55385 2305
rect 55345 2295 55350 2300
rect 55270 2275 55350 2295
rect 55270 2270 55275 2275
rect 55235 2265 55275 2270
rect 55345 2270 55350 2275
rect 55380 2270 55385 2300
rect 55345 2265 55385 2270
rect 58495 2300 58535 2305
rect 58495 2270 58500 2300
rect 58530 2295 58535 2300
rect 58605 2300 58645 2305
rect 58605 2295 58610 2300
rect 58530 2275 58610 2295
rect 58530 2270 58535 2275
rect 58495 2265 58535 2270
rect 58605 2270 58610 2275
rect 58640 2295 58645 2300
rect 58715 2300 58755 2305
rect 58715 2295 58720 2300
rect 58640 2275 58720 2295
rect 58640 2270 58645 2275
rect 58605 2265 58645 2270
rect 58715 2270 58720 2275
rect 58750 2295 58755 2300
rect 58825 2300 58865 2305
rect 58825 2295 58830 2300
rect 58750 2275 58830 2295
rect 58750 2270 58755 2275
rect 58715 2265 58755 2270
rect 58825 2270 58830 2275
rect 58860 2295 58865 2300
rect 58935 2300 58975 2305
rect 58935 2295 58940 2300
rect 58860 2275 58940 2295
rect 58860 2270 58865 2275
rect 58825 2265 58865 2270
rect 58935 2270 58940 2275
rect 58970 2295 58975 2300
rect 59045 2300 59085 2305
rect 59045 2295 59050 2300
rect 58970 2275 59050 2295
rect 58970 2270 58975 2275
rect 58935 2265 58975 2270
rect 59045 2270 59050 2275
rect 59080 2270 59085 2300
rect 59045 2265 59085 2270
rect 54135 2220 56675 2225
rect 54135 2190 54140 2220
rect 54170 2190 54180 2220
rect 54210 2190 54220 2220
rect 54250 2190 55075 2220
rect 55105 2190 55525 2220
rect 55555 2190 55565 2220
rect 55595 2190 55605 2220
rect 55635 2190 56090 2220
rect 56120 2190 56145 2220
rect 56175 2190 56200 2220
rect 56230 2190 56255 2220
rect 56285 2190 56310 2220
rect 56340 2190 56365 2220
rect 56395 2190 56420 2220
rect 56450 2190 56475 2220
rect 56505 2190 56530 2220
rect 56560 2190 56585 2220
rect 56615 2190 56640 2220
rect 56670 2190 56675 2220
rect 54135 2180 56675 2190
rect 54135 2150 54140 2180
rect 54170 2150 54180 2180
rect 54210 2150 54220 2180
rect 54250 2150 55075 2180
rect 55105 2150 55525 2180
rect 55555 2150 55565 2180
rect 55595 2150 55605 2180
rect 55635 2150 56090 2180
rect 56120 2150 56145 2180
rect 56175 2150 56200 2180
rect 56230 2150 56255 2180
rect 56285 2150 56310 2180
rect 56340 2150 56365 2180
rect 56395 2150 56420 2180
rect 56450 2150 56475 2180
rect 56505 2150 56530 2180
rect 56560 2150 56585 2180
rect 56615 2150 56640 2180
rect 56670 2150 56675 2180
rect 54135 2140 56675 2150
rect 54135 2110 54140 2140
rect 54170 2110 54180 2140
rect 54210 2110 54220 2140
rect 54250 2110 55075 2140
rect 55105 2110 55525 2140
rect 55555 2110 55565 2140
rect 55595 2110 55605 2140
rect 55635 2110 56090 2140
rect 56120 2110 56145 2140
rect 56175 2110 56200 2140
rect 56230 2110 56255 2140
rect 56285 2110 56310 2140
rect 56340 2110 56365 2140
rect 56395 2110 56420 2140
rect 56450 2110 56475 2140
rect 56505 2110 56530 2140
rect 56560 2110 56585 2140
rect 56615 2110 56640 2140
rect 56670 2110 56675 2140
rect 54135 2105 56675 2110
rect 57125 2220 59935 2225
rect 57125 2190 57130 2220
rect 57160 2190 57185 2220
rect 57215 2190 57240 2220
rect 57270 2190 57295 2220
rect 57325 2190 57350 2220
rect 57380 2190 57405 2220
rect 57435 2190 57460 2220
rect 57490 2190 57515 2220
rect 57545 2190 57570 2220
rect 57600 2190 57625 2220
rect 57655 2190 57680 2220
rect 57710 2190 58245 2220
rect 58275 2190 58285 2220
rect 58315 2190 58325 2220
rect 58355 2190 58775 2220
rect 58805 2190 59820 2220
rect 59850 2190 59860 2220
rect 59890 2190 59900 2220
rect 59930 2190 59935 2220
rect 57125 2180 59935 2190
rect 57125 2150 57130 2180
rect 57160 2150 57185 2180
rect 57215 2150 57240 2180
rect 57270 2150 57295 2180
rect 57325 2150 57350 2180
rect 57380 2150 57405 2180
rect 57435 2150 57460 2180
rect 57490 2150 57515 2180
rect 57545 2150 57570 2180
rect 57600 2150 57625 2180
rect 57655 2150 57680 2180
rect 57710 2150 58245 2180
rect 58275 2150 58285 2180
rect 58315 2150 58325 2180
rect 58355 2150 58775 2180
rect 58805 2150 59820 2180
rect 59850 2150 59860 2180
rect 59890 2150 59900 2180
rect 59930 2150 59935 2180
rect 57125 2140 59935 2150
rect 57125 2110 57130 2140
rect 57160 2110 57185 2140
rect 57215 2110 57240 2140
rect 57270 2110 57295 2140
rect 57325 2110 57350 2140
rect 57380 2110 57405 2140
rect 57435 2110 57460 2140
rect 57490 2110 57515 2140
rect 57545 2110 57570 2140
rect 57600 2110 57625 2140
rect 57655 2110 57680 2140
rect 57710 2110 58245 2140
rect 58275 2110 58285 2140
rect 58315 2110 58325 2140
rect 58355 2110 58775 2140
rect 58805 2110 59820 2140
rect 59850 2110 59860 2140
rect 59890 2110 59900 2140
rect 59930 2110 59935 2140
rect 57125 2105 59935 2110
rect 54105 2070 55385 2075
rect 54105 2040 54110 2070
rect 54140 2040 54150 2070
rect 54180 2040 54195 2070
rect 54225 2040 54235 2070
rect 54265 2040 54280 2070
rect 54310 2040 54320 2070
rect 54350 2040 54800 2070
rect 54830 2040 54855 2070
rect 54885 2040 54910 2070
rect 54940 2040 54965 2070
rect 54995 2040 55020 2070
rect 55050 2040 55075 2070
rect 55105 2040 55130 2070
rect 55160 2040 55185 2070
rect 55215 2040 55240 2070
rect 55270 2040 55295 2070
rect 55325 2040 55350 2070
rect 55380 2040 55385 2070
rect 58495 2070 59965 2075
rect 54105 2030 55385 2040
rect 54105 2000 54110 2030
rect 54140 2000 54150 2030
rect 54180 2000 54195 2030
rect 54225 2000 54235 2030
rect 54265 2000 54280 2030
rect 54310 2000 54320 2030
rect 54350 2000 54800 2030
rect 54830 2000 54855 2030
rect 54885 2000 54910 2030
rect 54940 2000 54965 2030
rect 54995 2000 55020 2030
rect 55050 2000 55075 2030
rect 55105 2000 55130 2030
rect 55160 2000 55185 2030
rect 55215 2000 55240 2030
rect 55270 2000 55295 2030
rect 55325 2000 55350 2030
rect 55380 2000 55385 2030
rect 54105 1990 55385 2000
rect 54105 1960 54110 1990
rect 54140 1960 54150 1990
rect 54180 1960 54195 1990
rect 54225 1960 54235 1990
rect 54265 1960 54280 1990
rect 54310 1960 54320 1990
rect 54350 1960 54800 1990
rect 54830 1960 54855 1990
rect 54885 1960 54910 1990
rect 54940 1960 54965 1990
rect 54995 1960 55020 1990
rect 55050 1960 55075 1990
rect 55105 1960 55130 1990
rect 55160 1960 55185 1990
rect 55215 1960 55240 1990
rect 55270 1960 55295 1990
rect 55325 1960 55350 1990
rect 55380 1960 55385 1990
rect 54105 1955 55385 1960
rect 56770 2045 58040 2050
rect 56770 2015 56775 2045
rect 56805 2015 56885 2045
rect 56915 2015 56995 2045
rect 57025 2015 57925 2045
rect 57955 2015 57965 2045
rect 57995 2015 58005 2045
rect 58035 2015 58040 2045
rect 56770 2005 58040 2015
rect 56770 1975 56775 2005
rect 56805 1975 56885 2005
rect 56915 1975 56995 2005
rect 57025 1975 57925 2005
rect 57955 1975 57965 2005
rect 57995 1975 58005 2005
rect 58035 1975 58040 2005
rect 56770 1965 58040 1975
rect 54740 1935 55780 1940
rect 54740 1905 54745 1935
rect 54775 1905 55405 1935
rect 55435 1905 55665 1935
rect 55695 1905 55705 1935
rect 55735 1905 55745 1935
rect 55775 1905 55780 1935
rect 56770 1935 56775 1965
rect 56805 1935 56885 1965
rect 56915 1935 56995 1965
rect 57025 1935 57925 1965
rect 57955 1935 57965 1965
rect 57995 1935 58005 1965
rect 58035 1935 58040 1965
rect 58495 2040 58500 2070
rect 58530 2040 58555 2070
rect 58585 2040 58610 2070
rect 58640 2040 58665 2070
rect 58695 2040 58720 2070
rect 58750 2040 58775 2070
rect 58805 2040 58830 2070
rect 58860 2040 58885 2070
rect 58915 2040 58940 2070
rect 58970 2040 58995 2070
rect 59025 2040 59050 2070
rect 59080 2040 59720 2070
rect 59750 2040 59760 2070
rect 59790 2040 59805 2070
rect 59835 2040 59845 2070
rect 59875 2040 59890 2070
rect 59920 2040 59930 2070
rect 59960 2040 59965 2070
rect 58495 2030 59965 2040
rect 58495 2000 58500 2030
rect 58530 2000 58555 2030
rect 58585 2000 58610 2030
rect 58640 2000 58665 2030
rect 58695 2000 58720 2030
rect 58750 2000 58775 2030
rect 58805 2000 58830 2030
rect 58860 2000 58885 2030
rect 58915 2000 58940 2030
rect 58970 2000 58995 2030
rect 59025 2000 59050 2030
rect 59080 2000 59720 2030
rect 59750 2000 59760 2030
rect 59790 2000 59805 2030
rect 59835 2000 59845 2030
rect 59875 2000 59890 2030
rect 59920 2000 59930 2030
rect 59960 2000 59965 2030
rect 58495 1990 59965 2000
rect 58495 1960 58500 1990
rect 58530 1960 58555 1990
rect 58585 1960 58610 1990
rect 58640 1960 58665 1990
rect 58695 1960 58720 1990
rect 58750 1960 58775 1990
rect 58805 1960 58830 1990
rect 58860 1960 58885 1990
rect 58915 1960 58940 1990
rect 58970 1960 58995 1990
rect 59025 1960 59050 1990
rect 59080 1960 59720 1990
rect 59750 1960 59760 1990
rect 59790 1960 59805 1990
rect 59835 1960 59845 1990
rect 59875 1960 59890 1990
rect 59920 1960 59930 1990
rect 59960 1960 59965 1990
rect 58495 1955 59965 1960
rect 56770 1930 58040 1935
rect 58100 1935 59140 1940
rect 54740 1895 55780 1905
rect 54740 1865 54745 1895
rect 54775 1865 55405 1895
rect 55435 1865 55665 1895
rect 55695 1865 55705 1895
rect 55735 1865 55745 1895
rect 55775 1865 55780 1895
rect 54740 1855 55780 1865
rect 54740 1825 54745 1855
rect 54775 1825 55405 1855
rect 55435 1825 55665 1855
rect 55695 1825 55705 1855
rect 55735 1825 55745 1855
rect 55775 1825 55780 1855
rect 54740 1820 55780 1825
rect 58100 1905 58105 1935
rect 58135 1905 58145 1935
rect 58175 1905 58185 1935
rect 58215 1905 58445 1935
rect 58475 1905 59105 1935
rect 59135 1905 59140 1935
rect 58100 1895 59140 1905
rect 58100 1865 58105 1895
rect 58135 1865 58145 1895
rect 58175 1865 58185 1895
rect 58215 1865 58445 1895
rect 58475 1865 59105 1895
rect 59135 1865 59140 1895
rect 58100 1855 59140 1865
rect 58100 1825 58105 1855
rect 58135 1825 58145 1855
rect 58175 1825 58185 1855
rect 58215 1825 58445 1855
rect 58475 1825 59105 1855
rect 59135 1825 59140 1855
rect 58100 1820 59140 1825
rect 53960 1800 55385 1805
rect 53960 1770 53965 1800
rect 53995 1770 54005 1800
rect 54035 1770 54045 1800
rect 54075 1770 54800 1800
rect 54830 1770 54910 1800
rect 54940 1770 55020 1800
rect 55050 1770 55130 1800
rect 55160 1770 55240 1800
rect 55270 1770 55350 1800
rect 55380 1770 55385 1800
rect 53960 1760 55385 1770
rect 53960 1730 53965 1760
rect 53995 1730 54005 1760
rect 54035 1730 54045 1760
rect 54075 1730 54800 1760
rect 54830 1730 54910 1760
rect 54940 1730 55020 1760
rect 55050 1730 55130 1760
rect 55160 1730 55240 1760
rect 55270 1730 55350 1760
rect 55380 1730 55385 1760
rect 57920 1800 60110 1805
rect 57920 1770 57925 1800
rect 57955 1770 57965 1800
rect 57995 1770 58005 1800
rect 58035 1770 58500 1800
rect 58530 1770 58610 1800
rect 58640 1770 58720 1800
rect 58750 1770 58830 1800
rect 58860 1770 58940 1800
rect 58970 1770 59050 1800
rect 59080 1770 59995 1800
rect 60025 1770 60035 1800
rect 60065 1770 60075 1800
rect 60105 1770 60110 1800
rect 57920 1760 60110 1770
rect 53960 1720 55385 1730
rect 53960 1690 53965 1720
rect 53995 1690 54005 1720
rect 54035 1690 54045 1720
rect 54075 1690 54800 1720
rect 54830 1690 54910 1720
rect 54940 1690 55020 1720
rect 55050 1690 55130 1720
rect 55160 1690 55240 1720
rect 55270 1690 55350 1720
rect 55380 1690 55385 1720
rect 55895 1735 55935 1740
rect 55895 1705 55900 1735
rect 55930 1730 55935 1735
rect 55995 1735 56025 1740
rect 55930 1710 55995 1730
rect 55930 1705 55935 1710
rect 55895 1700 55935 1705
rect 56690 1735 56720 1740
rect 55995 1700 56025 1705
rect 56140 1725 56180 1730
rect 56140 1695 56145 1725
rect 56175 1720 56180 1725
rect 56250 1725 56290 1730
rect 56250 1720 56255 1725
rect 56175 1700 56255 1720
rect 56175 1695 56180 1700
rect 56140 1690 56180 1695
rect 56250 1695 56255 1700
rect 56285 1720 56290 1725
rect 56360 1725 56400 1730
rect 56360 1720 56365 1725
rect 56285 1700 56365 1720
rect 56285 1695 56290 1700
rect 56250 1690 56290 1695
rect 56360 1695 56365 1700
rect 56395 1720 56400 1725
rect 56470 1725 56510 1730
rect 56470 1720 56475 1725
rect 56395 1700 56475 1720
rect 56395 1695 56400 1700
rect 56360 1690 56400 1695
rect 56470 1695 56475 1700
rect 56505 1720 56510 1725
rect 56580 1725 56620 1730
rect 56580 1720 56585 1725
rect 56505 1700 56585 1720
rect 56505 1695 56510 1700
rect 56470 1690 56510 1695
rect 56580 1695 56585 1700
rect 56615 1695 56620 1725
rect 57080 1735 57110 1740
rect 56720 1710 57080 1730
rect 56690 1700 56720 1705
rect 57920 1730 57925 1760
rect 57955 1730 57965 1760
rect 57995 1730 58005 1760
rect 58035 1730 58500 1760
rect 58530 1730 58610 1760
rect 58640 1730 58720 1760
rect 58750 1730 58830 1760
rect 58860 1730 58940 1760
rect 58970 1730 59050 1760
rect 59080 1730 59995 1760
rect 60025 1730 60035 1760
rect 60065 1730 60075 1760
rect 60105 1730 60110 1760
rect 57080 1700 57110 1705
rect 57180 1725 57220 1730
rect 56580 1690 56620 1695
rect 57180 1695 57185 1725
rect 57215 1720 57220 1725
rect 57290 1725 57330 1730
rect 57290 1720 57295 1725
rect 57215 1700 57295 1720
rect 57215 1695 57220 1700
rect 57180 1690 57220 1695
rect 57290 1695 57295 1700
rect 57325 1720 57330 1725
rect 57400 1725 57440 1730
rect 57400 1720 57405 1725
rect 57325 1700 57405 1720
rect 57325 1695 57330 1700
rect 57290 1690 57330 1695
rect 57400 1695 57405 1700
rect 57435 1720 57440 1725
rect 57510 1725 57550 1730
rect 57510 1720 57515 1725
rect 57435 1700 57515 1720
rect 57435 1695 57440 1700
rect 57400 1690 57440 1695
rect 57510 1695 57515 1700
rect 57545 1720 57550 1725
rect 57620 1725 57660 1730
rect 57620 1720 57625 1725
rect 57545 1700 57625 1720
rect 57545 1695 57550 1700
rect 57510 1690 57550 1695
rect 57620 1695 57625 1700
rect 57655 1695 57660 1725
rect 57620 1690 57660 1695
rect 57920 1720 60110 1730
rect 57920 1690 57925 1720
rect 57955 1690 57965 1720
rect 57995 1690 58005 1720
rect 58035 1690 58500 1720
rect 58530 1690 58610 1720
rect 58640 1690 58720 1720
rect 58750 1690 58830 1720
rect 58860 1690 58940 1720
rect 58970 1690 59050 1720
rect 59080 1690 59995 1720
rect 60025 1690 60035 1720
rect 60065 1690 60075 1720
rect 60105 1690 60110 1720
rect 53960 1685 55385 1690
rect 57920 1685 60110 1690
rect 54745 1680 54775 1685
rect 56085 1680 56125 1685
rect 54850 1665 54890 1670
rect 54850 1635 54855 1665
rect 54885 1660 54890 1665
rect 54960 1665 55000 1670
rect 54960 1660 54965 1665
rect 54885 1640 54965 1660
rect 54885 1635 54890 1640
rect 54850 1630 54890 1635
rect 54960 1635 54965 1640
rect 54995 1660 55000 1665
rect 55070 1665 55110 1670
rect 55070 1660 55075 1665
rect 54995 1640 55075 1660
rect 54995 1635 55000 1640
rect 54960 1630 55000 1635
rect 55070 1635 55075 1640
rect 55105 1660 55110 1665
rect 55180 1665 55220 1670
rect 55180 1660 55185 1665
rect 55105 1640 55185 1660
rect 55105 1635 55110 1640
rect 55070 1630 55110 1635
rect 55180 1635 55185 1640
rect 55215 1660 55220 1665
rect 55290 1665 55330 1670
rect 55290 1660 55295 1665
rect 55215 1640 55295 1660
rect 55215 1635 55220 1640
rect 55180 1630 55220 1635
rect 55290 1635 55295 1640
rect 55325 1635 55330 1665
rect 56085 1650 56090 1680
rect 56120 1675 56125 1680
rect 56195 1680 56235 1685
rect 56195 1675 56200 1680
rect 56120 1655 56200 1675
rect 56120 1650 56125 1655
rect 56085 1645 56125 1650
rect 56195 1650 56200 1655
rect 56230 1675 56235 1680
rect 56305 1680 56345 1685
rect 56305 1675 56310 1680
rect 56230 1655 56310 1675
rect 56230 1650 56235 1655
rect 56195 1645 56235 1650
rect 56305 1650 56310 1655
rect 56340 1675 56345 1680
rect 56415 1680 56455 1685
rect 56415 1675 56420 1680
rect 56340 1655 56420 1675
rect 56340 1650 56345 1655
rect 56305 1645 56345 1650
rect 56415 1650 56420 1655
rect 56450 1675 56455 1680
rect 56525 1680 56565 1685
rect 56525 1675 56530 1680
rect 56450 1655 56530 1675
rect 56450 1650 56455 1655
rect 56415 1645 56455 1650
rect 56525 1650 56530 1655
rect 56560 1675 56565 1680
rect 56635 1680 56675 1685
rect 56635 1675 56640 1680
rect 56560 1655 56640 1675
rect 56560 1650 56565 1655
rect 56525 1645 56565 1650
rect 56635 1650 56640 1655
rect 56670 1650 56675 1680
rect 56635 1645 56675 1650
rect 57125 1680 57165 1685
rect 57125 1650 57130 1680
rect 57160 1675 57165 1680
rect 57235 1680 57275 1685
rect 57235 1675 57240 1680
rect 57160 1655 57240 1675
rect 57160 1650 57165 1655
rect 57125 1645 57165 1650
rect 57235 1650 57240 1655
rect 57270 1675 57275 1680
rect 57345 1680 57385 1685
rect 57345 1675 57350 1680
rect 57270 1655 57350 1675
rect 57270 1650 57275 1655
rect 57235 1645 57275 1650
rect 57345 1650 57350 1655
rect 57380 1675 57385 1680
rect 57455 1680 57495 1685
rect 57455 1675 57460 1680
rect 57380 1655 57460 1675
rect 57380 1650 57385 1655
rect 57345 1645 57385 1650
rect 57455 1650 57460 1655
rect 57490 1675 57495 1680
rect 57565 1680 57605 1685
rect 57565 1675 57570 1680
rect 57490 1655 57570 1675
rect 57490 1650 57495 1655
rect 57455 1645 57495 1650
rect 57565 1650 57570 1655
rect 57600 1675 57605 1680
rect 57675 1680 57715 1685
rect 58445 1680 58475 1685
rect 59105 1680 59135 1685
rect 57675 1675 57680 1680
rect 57600 1655 57680 1675
rect 57600 1650 57605 1655
rect 57565 1645 57605 1650
rect 57675 1650 57680 1655
rect 57710 1650 57715 1680
rect 57675 1645 57715 1650
rect 58550 1665 58590 1670
rect 55290 1630 55330 1635
rect 58550 1635 58555 1665
rect 58585 1660 58590 1665
rect 58660 1665 58700 1670
rect 58660 1660 58665 1665
rect 58585 1640 58665 1660
rect 58585 1635 58590 1640
rect 58550 1630 58590 1635
rect 58660 1635 58665 1640
rect 58695 1660 58700 1665
rect 58770 1665 58810 1670
rect 58770 1660 58775 1665
rect 58695 1640 58775 1660
rect 58695 1635 58700 1640
rect 58660 1630 58700 1635
rect 58770 1635 58775 1640
rect 58805 1660 58810 1665
rect 58880 1665 58920 1670
rect 58880 1660 58885 1665
rect 58805 1640 58885 1660
rect 58805 1635 58810 1640
rect 58770 1630 58810 1635
rect 58880 1635 58885 1640
rect 58915 1660 58920 1665
rect 58990 1665 59030 1670
rect 58990 1660 58995 1665
rect 58915 1640 58995 1660
rect 58915 1635 58920 1640
rect 58880 1630 58920 1635
rect 58990 1635 58995 1640
rect 59025 1635 59030 1665
rect 58990 1630 59030 1635
rect 56140 1490 56180 1495
rect 56140 1460 56145 1490
rect 56175 1485 56180 1490
rect 56250 1490 56290 1495
rect 56250 1485 56255 1490
rect 56175 1465 56255 1485
rect 56175 1460 56180 1465
rect 56140 1455 56180 1460
rect 56250 1460 56255 1465
rect 56285 1485 56290 1490
rect 56360 1490 56400 1495
rect 56360 1485 56365 1490
rect 56285 1465 56365 1485
rect 56285 1460 56290 1465
rect 56250 1455 56290 1460
rect 56360 1460 56365 1465
rect 56395 1485 56400 1490
rect 56470 1490 56510 1495
rect 56470 1485 56475 1490
rect 56395 1465 56475 1485
rect 56395 1460 56400 1465
rect 56360 1455 56400 1460
rect 56470 1460 56475 1465
rect 56505 1485 56510 1490
rect 56580 1490 56620 1495
rect 56580 1485 56585 1490
rect 56505 1465 56585 1485
rect 56505 1460 56510 1465
rect 56470 1455 56510 1460
rect 56580 1460 56585 1465
rect 56615 1460 56620 1490
rect 56580 1455 56620 1460
rect 57180 1490 57220 1495
rect 57180 1460 57185 1490
rect 57215 1485 57220 1490
rect 57290 1490 57330 1495
rect 57290 1485 57295 1490
rect 57215 1465 57295 1485
rect 57215 1460 57220 1465
rect 57180 1455 57220 1460
rect 57290 1460 57295 1465
rect 57325 1485 57330 1490
rect 57400 1490 57440 1495
rect 57400 1485 57405 1490
rect 57325 1465 57405 1485
rect 57325 1460 57330 1465
rect 57290 1455 57330 1460
rect 57400 1460 57405 1465
rect 57435 1485 57440 1490
rect 57510 1490 57550 1495
rect 57510 1485 57515 1490
rect 57435 1465 57515 1485
rect 57435 1460 57440 1465
rect 57400 1455 57440 1460
rect 57510 1460 57515 1465
rect 57545 1485 57550 1490
rect 57620 1490 57660 1495
rect 57620 1485 57625 1490
rect 57545 1465 57625 1485
rect 57545 1460 57550 1465
rect 57510 1455 57550 1460
rect 57620 1460 57625 1465
rect 57655 1460 57660 1490
rect 57620 1455 57660 1460
rect 56085 1445 56125 1450
rect 56085 1415 56090 1445
rect 56120 1440 56125 1445
rect 56195 1445 56235 1450
rect 56195 1440 56200 1445
rect 56120 1420 56200 1440
rect 56120 1415 56125 1420
rect 54600 1410 54640 1415
rect 54600 1380 54605 1410
rect 54635 1405 54640 1410
rect 54850 1410 54890 1415
rect 54850 1405 54855 1410
rect 54635 1385 54855 1405
rect 54635 1380 54640 1385
rect 54600 1375 54640 1380
rect 54850 1380 54855 1385
rect 54885 1405 54890 1410
rect 54960 1410 55000 1415
rect 54960 1405 54965 1410
rect 54885 1385 54965 1405
rect 54885 1380 54890 1385
rect 54850 1375 54890 1380
rect 54960 1380 54965 1385
rect 54995 1405 55000 1410
rect 55070 1410 55110 1415
rect 55070 1405 55075 1410
rect 54995 1385 55075 1405
rect 54995 1380 55000 1385
rect 54960 1375 55000 1380
rect 55070 1380 55075 1385
rect 55105 1405 55110 1410
rect 55180 1410 55220 1415
rect 55180 1405 55185 1410
rect 55105 1385 55185 1405
rect 55105 1380 55110 1385
rect 55070 1375 55110 1380
rect 55180 1380 55185 1385
rect 55215 1405 55220 1410
rect 55290 1410 55330 1415
rect 56085 1410 56125 1415
rect 56195 1415 56200 1420
rect 56230 1440 56235 1445
rect 56305 1445 56345 1450
rect 56305 1440 56310 1445
rect 56230 1420 56310 1440
rect 56230 1415 56235 1420
rect 56195 1410 56235 1415
rect 56305 1415 56310 1420
rect 56340 1440 56345 1445
rect 56415 1445 56455 1450
rect 56415 1440 56420 1445
rect 56340 1420 56420 1440
rect 56340 1415 56345 1420
rect 56305 1410 56345 1415
rect 56415 1415 56420 1420
rect 56450 1440 56455 1445
rect 56525 1445 56565 1450
rect 56525 1440 56530 1445
rect 56450 1420 56530 1440
rect 56450 1415 56455 1420
rect 56415 1410 56455 1415
rect 56525 1415 56530 1420
rect 56560 1440 56565 1445
rect 56635 1445 56675 1450
rect 56635 1440 56640 1445
rect 56560 1420 56640 1440
rect 56560 1415 56565 1420
rect 56525 1410 56565 1415
rect 56635 1415 56640 1420
rect 56670 1415 56675 1445
rect 56635 1410 56675 1415
rect 57125 1445 57165 1450
rect 57125 1415 57130 1445
rect 57160 1440 57165 1445
rect 57235 1445 57275 1450
rect 57235 1440 57240 1445
rect 57160 1420 57240 1440
rect 57160 1415 57165 1420
rect 57125 1410 57165 1415
rect 57235 1415 57240 1420
rect 57270 1440 57275 1445
rect 57345 1445 57385 1450
rect 57345 1440 57350 1445
rect 57270 1420 57350 1440
rect 57270 1415 57275 1420
rect 57235 1410 57275 1415
rect 57345 1415 57350 1420
rect 57380 1440 57385 1445
rect 57455 1445 57495 1450
rect 57455 1440 57460 1445
rect 57380 1420 57460 1440
rect 57380 1415 57385 1420
rect 57345 1410 57385 1415
rect 57455 1415 57460 1420
rect 57490 1440 57495 1445
rect 57565 1445 57605 1450
rect 57565 1440 57570 1445
rect 57490 1420 57570 1440
rect 57490 1415 57495 1420
rect 57455 1410 57495 1415
rect 57565 1415 57570 1420
rect 57600 1440 57605 1445
rect 57675 1445 57715 1450
rect 57675 1440 57680 1445
rect 57600 1420 57680 1440
rect 57600 1415 57605 1420
rect 57565 1410 57605 1415
rect 57675 1415 57680 1420
rect 57710 1415 57715 1445
rect 59715 1435 59965 1445
rect 57675 1410 57715 1415
rect 58550 1410 58590 1415
rect 55290 1405 55295 1410
rect 55215 1385 55295 1405
rect 55215 1380 55220 1385
rect 55180 1375 55220 1380
rect 55290 1380 55295 1385
rect 55325 1380 55330 1410
rect 55290 1375 55330 1380
rect 56030 1390 58040 1395
rect 54105 1360 54355 1370
rect 54105 1330 54115 1360
rect 54145 1330 54165 1360
rect 54195 1330 54215 1360
rect 54245 1330 54265 1360
rect 54295 1330 54315 1360
rect 54345 1330 54355 1360
rect 56030 1360 56035 1390
rect 56065 1360 56695 1390
rect 56725 1360 57075 1390
rect 57105 1360 57735 1390
rect 57765 1360 57925 1390
rect 57955 1360 57965 1390
rect 57995 1360 58005 1390
rect 58035 1360 58040 1390
rect 58550 1380 58555 1410
rect 58585 1405 58590 1410
rect 58660 1410 58700 1415
rect 58660 1405 58665 1410
rect 58585 1385 58665 1405
rect 58585 1380 58590 1385
rect 58550 1375 58590 1380
rect 58660 1380 58665 1385
rect 58695 1405 58700 1410
rect 58770 1410 58810 1415
rect 58770 1405 58775 1410
rect 58695 1385 58775 1405
rect 58695 1380 58700 1385
rect 58660 1375 58700 1380
rect 58770 1380 58775 1385
rect 58805 1405 58810 1410
rect 58880 1410 58920 1415
rect 58880 1405 58885 1410
rect 58805 1385 58885 1405
rect 58805 1380 58810 1385
rect 58770 1375 58810 1380
rect 58880 1380 58885 1385
rect 58915 1405 58920 1410
rect 58990 1410 59030 1415
rect 58990 1405 58995 1410
rect 58915 1385 58995 1405
rect 58915 1380 58920 1385
rect 58880 1375 58920 1380
rect 58990 1380 58995 1385
rect 59025 1405 59030 1410
rect 59430 1410 59470 1415
rect 59430 1405 59435 1410
rect 59025 1385 59435 1405
rect 59025 1380 59030 1385
rect 58990 1375 59030 1380
rect 59430 1380 59435 1385
rect 59465 1380 59470 1410
rect 59430 1375 59470 1380
rect 59715 1405 59725 1435
rect 59755 1405 59775 1435
rect 59805 1405 59825 1435
rect 59855 1405 59875 1435
rect 59905 1405 59925 1435
rect 59955 1405 59965 1435
rect 59715 1385 59965 1405
rect 56030 1350 58040 1360
rect 59715 1355 59725 1385
rect 59755 1355 59775 1385
rect 59805 1355 59825 1385
rect 59855 1355 59875 1385
rect 59905 1355 59925 1385
rect 59955 1355 59965 1385
rect 54105 1310 54355 1330
rect 54105 1280 54115 1310
rect 54145 1280 54165 1310
rect 54195 1280 54215 1310
rect 54245 1280 54265 1310
rect 54295 1280 54315 1310
rect 54345 1280 54355 1310
rect 54105 1260 54355 1280
rect 55235 1345 55640 1350
rect 55235 1315 55240 1345
rect 55270 1315 55525 1345
rect 55555 1315 55565 1345
rect 55595 1315 55605 1345
rect 55635 1315 55640 1345
rect 55235 1305 55640 1315
rect 55235 1275 55240 1305
rect 55270 1275 55525 1305
rect 55555 1275 55565 1305
rect 55595 1275 55605 1305
rect 55635 1275 55640 1305
rect 56030 1320 56035 1350
rect 56065 1320 56695 1350
rect 56725 1320 57075 1350
rect 57105 1320 57735 1350
rect 57765 1320 57925 1350
rect 57955 1320 57965 1350
rect 57995 1320 58005 1350
rect 58035 1320 58040 1350
rect 56030 1310 58040 1320
rect 56030 1280 56035 1310
rect 56065 1280 56695 1310
rect 56725 1280 57075 1310
rect 57105 1280 57735 1310
rect 57765 1280 57925 1310
rect 57955 1280 57965 1310
rect 57995 1280 58005 1310
rect 58035 1280 58040 1310
rect 56030 1275 58040 1280
rect 58240 1345 58645 1350
rect 58240 1315 58245 1345
rect 58275 1315 58285 1345
rect 58315 1315 58325 1345
rect 58355 1315 58610 1345
rect 58640 1315 58645 1345
rect 58240 1305 58645 1315
rect 58240 1275 58245 1305
rect 58275 1275 58285 1305
rect 58315 1275 58325 1305
rect 58355 1275 58610 1305
rect 58640 1275 58645 1305
rect 59715 1335 59965 1355
rect 59715 1305 59725 1335
rect 59755 1305 59775 1335
rect 59805 1305 59825 1335
rect 59855 1305 59875 1335
rect 59905 1305 59925 1335
rect 59955 1305 59965 1335
rect 59715 1295 59965 1305
rect 55235 1270 55640 1275
rect 58240 1270 58645 1275
rect 54105 1230 54115 1260
rect 54145 1230 54165 1260
rect 54195 1230 54215 1260
rect 54245 1230 54265 1260
rect 54295 1230 54315 1260
rect 54345 1230 54355 1260
rect 55795 1235 58040 1240
rect 54105 1220 54355 1230
rect 54645 1225 54685 1230
rect 54645 1195 54650 1225
rect 54680 1220 54685 1225
rect 54850 1225 54890 1230
rect 54850 1220 54855 1225
rect 54680 1200 54855 1220
rect 54680 1195 54685 1200
rect 54645 1190 54685 1195
rect 54850 1195 54855 1200
rect 54885 1220 54890 1225
rect 54960 1225 55000 1230
rect 54960 1220 54965 1225
rect 54885 1200 54965 1220
rect 54885 1195 54890 1200
rect 54850 1190 54890 1195
rect 54960 1195 54965 1200
rect 54995 1220 55000 1225
rect 55070 1225 55110 1230
rect 55070 1220 55075 1225
rect 54995 1200 55075 1220
rect 54995 1195 55000 1200
rect 54960 1190 55000 1195
rect 55070 1195 55075 1200
rect 55105 1220 55110 1225
rect 55180 1225 55220 1230
rect 55180 1220 55185 1225
rect 55105 1200 55185 1220
rect 55105 1195 55110 1200
rect 55070 1190 55110 1195
rect 55180 1195 55185 1200
rect 55215 1220 55220 1225
rect 55290 1225 55330 1230
rect 55290 1220 55295 1225
rect 55215 1200 55295 1220
rect 55215 1195 55220 1200
rect 55180 1190 55220 1195
rect 55290 1195 55295 1200
rect 55325 1195 55330 1225
rect 55290 1190 55330 1195
rect 55795 1205 55800 1235
rect 55830 1205 55840 1235
rect 55870 1205 56885 1235
rect 56915 1205 57925 1235
rect 57955 1205 57965 1235
rect 57995 1205 58005 1235
rect 58035 1205 58040 1235
rect 55795 1195 58040 1205
rect 55795 1165 55800 1195
rect 55830 1165 55840 1195
rect 55870 1165 56885 1195
rect 56915 1165 57925 1195
rect 57955 1165 57965 1195
rect 57995 1165 58005 1195
rect 58035 1165 58040 1195
rect 58550 1225 58590 1230
rect 58550 1195 58555 1225
rect 58585 1220 58590 1225
rect 58660 1225 58700 1230
rect 58660 1220 58665 1225
rect 58585 1200 58665 1220
rect 58585 1195 58590 1200
rect 58550 1190 58590 1195
rect 58660 1195 58665 1200
rect 58695 1220 58700 1225
rect 58770 1225 58810 1230
rect 58770 1220 58775 1225
rect 58695 1200 58775 1220
rect 58695 1195 58700 1200
rect 58660 1190 58700 1195
rect 58770 1195 58775 1200
rect 58805 1220 58810 1225
rect 58880 1225 58920 1230
rect 58880 1220 58885 1225
rect 58805 1200 58885 1220
rect 58805 1195 58810 1200
rect 58770 1190 58810 1195
rect 58880 1195 58885 1200
rect 58915 1220 58920 1225
rect 58990 1225 59030 1230
rect 58990 1220 58995 1225
rect 58915 1200 58995 1220
rect 58915 1195 58920 1200
rect 58880 1190 58920 1195
rect 58990 1195 58995 1200
rect 59025 1220 59030 1225
rect 59195 1225 59235 1230
rect 59195 1220 59200 1225
rect 59025 1200 59200 1220
rect 59025 1195 59030 1200
rect 58990 1190 59030 1195
rect 59195 1195 59200 1200
rect 59230 1195 59235 1225
rect 59195 1190 59235 1195
rect 55795 1155 58040 1165
rect 55795 1125 55800 1155
rect 55830 1125 55840 1155
rect 55870 1125 56885 1155
rect 56915 1125 57925 1155
rect 57955 1125 57965 1155
rect 57995 1125 58005 1155
rect 58035 1125 58040 1155
rect 55795 1120 58040 1125
rect 56145 1065 56175 1070
rect 56085 1055 56125 1060
rect 56040 1045 56070 1050
rect 56030 1020 56040 1040
rect 56085 1025 56090 1055
rect 56120 1050 56125 1055
rect 56120 1035 56145 1050
rect 56255 1065 56285 1070
rect 56195 1055 56235 1060
rect 56195 1050 56200 1055
rect 56175 1035 56200 1050
rect 56120 1030 56200 1035
rect 56120 1025 56125 1030
rect 56085 1020 56125 1025
rect 56195 1025 56200 1030
rect 56230 1050 56235 1055
rect 56230 1035 56255 1050
rect 56365 1065 56395 1070
rect 56305 1055 56345 1060
rect 56305 1050 56310 1055
rect 56285 1035 56310 1050
rect 56230 1030 56310 1035
rect 56230 1025 56235 1030
rect 56195 1020 56235 1025
rect 56305 1025 56310 1030
rect 56340 1050 56345 1055
rect 56340 1035 56365 1050
rect 56475 1065 56505 1070
rect 56415 1055 56455 1060
rect 56415 1050 56420 1055
rect 56395 1035 56420 1050
rect 56340 1030 56420 1035
rect 56340 1025 56345 1030
rect 56305 1020 56345 1025
rect 56415 1025 56420 1030
rect 56450 1050 56455 1055
rect 56450 1035 56475 1050
rect 56585 1065 56615 1070
rect 56525 1055 56565 1060
rect 56525 1050 56530 1055
rect 56505 1035 56530 1050
rect 56450 1030 56530 1035
rect 56450 1025 56455 1030
rect 56415 1020 56455 1025
rect 56525 1025 56530 1030
rect 56560 1050 56565 1055
rect 56560 1035 56585 1050
rect 57185 1065 57215 1070
rect 56635 1055 56675 1060
rect 56635 1050 56640 1055
rect 56615 1035 56640 1050
rect 56560 1030 56640 1035
rect 56560 1025 56565 1030
rect 56525 1020 56565 1025
rect 56635 1025 56640 1030
rect 56670 1025 56675 1055
rect 56635 1020 56675 1025
rect 56690 1055 56720 1060
rect 56840 1055 56870 1060
rect 56720 1030 56840 1050
rect 56690 1020 56720 1025
rect 56840 1020 56870 1025
rect 56930 1055 56960 1060
rect 57080 1055 57110 1060
rect 56960 1030 57080 1050
rect 56930 1020 56960 1025
rect 57080 1020 57110 1025
rect 57125 1055 57165 1060
rect 57125 1025 57130 1055
rect 57160 1050 57165 1055
rect 57160 1035 57185 1050
rect 57295 1065 57325 1070
rect 57235 1055 57275 1060
rect 57235 1050 57240 1055
rect 57215 1035 57240 1050
rect 57160 1030 57240 1035
rect 57160 1025 57165 1030
rect 57125 1020 57165 1025
rect 57235 1025 57240 1030
rect 57270 1050 57275 1055
rect 57270 1035 57295 1050
rect 57405 1065 57435 1070
rect 57345 1055 57385 1060
rect 57345 1050 57350 1055
rect 57325 1035 57350 1050
rect 57270 1030 57350 1035
rect 57270 1025 57275 1030
rect 57235 1020 57275 1025
rect 57345 1025 57350 1030
rect 57380 1050 57385 1055
rect 57380 1035 57405 1050
rect 57515 1065 57545 1070
rect 57455 1055 57495 1060
rect 57455 1050 57460 1055
rect 57435 1035 57460 1050
rect 57380 1030 57460 1035
rect 57380 1025 57385 1030
rect 57345 1020 57385 1025
rect 57455 1025 57460 1030
rect 57490 1050 57495 1055
rect 57490 1035 57515 1050
rect 57625 1065 57655 1070
rect 57565 1055 57605 1060
rect 57565 1050 57570 1055
rect 57545 1035 57570 1050
rect 57490 1030 57570 1035
rect 57490 1025 57495 1030
rect 57455 1020 57495 1025
rect 57565 1025 57570 1030
rect 57600 1050 57605 1055
rect 57600 1035 57625 1050
rect 57675 1055 57715 1060
rect 57675 1050 57680 1055
rect 57655 1035 57680 1050
rect 57600 1030 57680 1035
rect 57600 1025 57605 1030
rect 57565 1020 57605 1025
rect 57675 1025 57680 1030
rect 57710 1025 57715 1055
rect 57675 1020 57715 1025
rect 57730 1045 57760 1050
rect 57760 1020 57770 1040
rect 56040 1010 56070 1015
rect 56140 1010 56180 1015
rect 56140 980 56145 1010
rect 56175 1005 56180 1010
rect 56250 1010 56290 1015
rect 56250 1005 56255 1010
rect 56175 985 56255 1005
rect 56175 980 56180 985
rect 56140 975 56180 980
rect 56250 980 56255 985
rect 56285 1005 56290 1010
rect 56360 1010 56400 1015
rect 56360 1005 56365 1010
rect 56285 985 56365 1005
rect 56285 980 56290 985
rect 56250 975 56290 980
rect 56360 980 56365 985
rect 56395 1005 56400 1010
rect 56470 1010 56510 1015
rect 56470 1005 56475 1010
rect 56395 985 56475 1005
rect 56395 980 56400 985
rect 56360 975 56400 980
rect 56470 980 56475 985
rect 56505 1005 56510 1010
rect 56580 1010 56620 1015
rect 56580 1005 56585 1010
rect 56505 985 56585 1005
rect 56505 980 56510 985
rect 56470 975 56510 980
rect 56580 980 56585 985
rect 56615 1005 56620 1010
rect 57180 1010 57220 1015
rect 57180 1005 57185 1010
rect 56615 985 57185 1005
rect 56615 980 56620 985
rect 56580 975 56620 980
rect 57180 980 57185 985
rect 57215 1005 57220 1010
rect 57290 1010 57330 1015
rect 57290 1005 57295 1010
rect 57215 985 57295 1005
rect 57215 980 57220 985
rect 57180 975 57220 980
rect 57290 980 57295 985
rect 57325 1005 57330 1010
rect 57400 1010 57440 1015
rect 57400 1005 57405 1010
rect 57325 985 57405 1005
rect 57325 980 57330 985
rect 57290 975 57330 980
rect 57400 980 57405 985
rect 57435 1005 57440 1010
rect 57510 1010 57550 1015
rect 57510 1005 57515 1010
rect 57435 985 57515 1005
rect 57435 980 57440 985
rect 57400 975 57440 980
rect 57510 980 57515 985
rect 57545 1005 57550 1010
rect 57620 1010 57660 1015
rect 57730 1010 57760 1015
rect 57620 1005 57625 1010
rect 57545 985 57625 1005
rect 57545 980 57550 985
rect 57510 975 57550 980
rect 57620 980 57625 985
rect 57655 980 57660 1010
rect 57620 975 57660 980
rect 54380 915 54415 916
rect 59655 915 59690 916
rect 54380 910 54475 915
rect 54415 875 54440 910
rect 54380 870 54475 875
rect 54500 910 54535 915
rect 54500 870 54535 875
rect 54560 910 54595 915
rect 59475 910 59510 915
rect 54645 905 54685 910
rect 54645 900 54650 905
rect 54595 880 54650 900
rect 54560 870 54595 875
rect 54645 875 54650 880
rect 54680 875 54685 905
rect 59195 905 59235 910
rect 54645 870 54685 875
rect 54850 885 54890 890
rect 54850 855 54855 885
rect 54885 880 54890 885
rect 54960 885 55000 890
rect 54960 880 54965 885
rect 54885 860 54965 880
rect 54885 855 54890 860
rect 54850 850 54890 855
rect 54960 855 54965 860
rect 54995 880 55000 885
rect 55070 885 55110 890
rect 55070 880 55075 885
rect 54995 860 55075 880
rect 54995 855 55000 860
rect 54960 850 55000 855
rect 55070 855 55075 860
rect 55105 880 55110 885
rect 55180 885 55220 890
rect 55180 880 55185 885
rect 55105 860 55185 880
rect 55105 855 55110 860
rect 55070 850 55110 855
rect 55180 855 55185 860
rect 55215 880 55220 885
rect 55290 885 55330 890
rect 55290 880 55295 885
rect 55215 860 55295 880
rect 55215 855 55220 860
rect 55180 850 55220 855
rect 55290 855 55295 860
rect 55325 855 55330 885
rect 55290 850 55330 855
rect 58550 885 58590 890
rect 58550 855 58555 885
rect 58585 880 58590 885
rect 58660 885 58700 890
rect 58660 880 58665 885
rect 58585 860 58665 880
rect 58585 855 58590 860
rect 58550 850 58590 855
rect 58660 855 58665 860
rect 58695 880 58700 885
rect 58770 885 58810 890
rect 58770 880 58775 885
rect 58695 860 58775 880
rect 58695 855 58700 860
rect 58660 850 58700 855
rect 58770 855 58775 860
rect 58805 880 58810 885
rect 58880 885 58920 890
rect 58880 880 58885 885
rect 58805 860 58885 880
rect 58805 855 58810 860
rect 58770 850 58810 855
rect 58880 855 58885 860
rect 58915 880 58920 885
rect 58990 885 59030 890
rect 58990 880 58995 885
rect 58915 860 58995 880
rect 58915 855 58920 860
rect 58880 850 58920 855
rect 58990 855 58995 860
rect 59025 855 59030 885
rect 59195 875 59200 905
rect 59230 900 59235 905
rect 59230 880 59475 900
rect 59230 875 59235 880
rect 59195 870 59235 875
rect 59475 870 59510 875
rect 59535 910 59570 915
rect 59535 870 59570 875
rect 59595 910 59690 915
rect 59630 875 59655 910
rect 59595 870 59690 875
rect 58990 850 59030 855
rect 54500 835 54540 840
rect 54500 805 54505 835
rect 54535 825 54540 835
rect 54600 835 54640 840
rect 59430 835 59470 840
rect 54600 825 54605 835
rect 54535 810 54605 825
rect 54535 805 54540 810
rect 54500 800 54540 805
rect 54600 805 54605 810
rect 54635 805 54640 835
rect 58100 830 59085 835
rect 54600 800 54640 805
rect 54795 825 55780 830
rect 54795 795 54800 825
rect 54830 795 54910 825
rect 54940 795 55020 825
rect 55050 795 55130 825
rect 55160 795 55240 825
rect 55270 795 55350 825
rect 55380 795 55665 825
rect 55695 795 55705 825
rect 55735 795 55745 825
rect 55775 795 55780 825
rect 54795 785 55780 795
rect 54795 755 54800 785
rect 54830 755 54910 785
rect 54940 755 55020 785
rect 55050 755 55130 785
rect 55160 755 55240 785
rect 55270 755 55350 785
rect 55380 755 55665 785
rect 55695 755 55705 785
rect 55735 755 55745 785
rect 55775 755 55780 785
rect 56085 815 56125 820
rect 56085 785 56090 815
rect 56120 810 56125 815
rect 56195 815 56235 820
rect 56195 810 56200 815
rect 56120 790 56200 810
rect 56120 785 56125 790
rect 56085 780 56125 785
rect 56195 785 56200 790
rect 56230 810 56235 815
rect 56305 815 56345 820
rect 56305 810 56310 815
rect 56230 790 56310 810
rect 56230 785 56235 790
rect 56195 780 56235 785
rect 56305 785 56310 790
rect 56340 810 56345 815
rect 56415 815 56455 820
rect 56415 810 56420 815
rect 56340 790 56420 810
rect 56340 785 56345 790
rect 56305 780 56345 785
rect 56415 785 56420 790
rect 56450 810 56455 815
rect 56525 815 56565 820
rect 56525 810 56530 815
rect 56450 790 56530 810
rect 56450 785 56455 790
rect 56415 780 56455 785
rect 56525 785 56530 790
rect 56560 810 56565 815
rect 56635 815 56675 820
rect 56635 810 56640 815
rect 56560 790 56640 810
rect 56560 785 56565 790
rect 56525 780 56565 785
rect 56635 785 56640 790
rect 56670 785 56675 815
rect 56635 780 56675 785
rect 56825 815 56865 820
rect 56825 785 56830 815
rect 56860 810 56865 815
rect 56935 815 56975 820
rect 56935 810 56940 815
rect 56860 790 56940 810
rect 56860 785 56865 790
rect 56825 780 56865 785
rect 56935 785 56940 790
rect 56970 785 56975 815
rect 56935 780 56975 785
rect 57125 815 57165 820
rect 57125 785 57130 815
rect 57160 810 57165 815
rect 57235 815 57275 820
rect 57235 810 57240 815
rect 57160 790 57240 810
rect 57160 785 57165 790
rect 57125 780 57165 785
rect 57235 785 57240 790
rect 57270 810 57275 815
rect 57345 815 57385 820
rect 57345 810 57350 815
rect 57270 790 57350 810
rect 57270 785 57275 790
rect 57235 780 57275 785
rect 57345 785 57350 790
rect 57380 810 57385 815
rect 57455 815 57495 820
rect 57455 810 57460 815
rect 57380 790 57460 810
rect 57380 785 57385 790
rect 57345 780 57385 785
rect 57455 785 57460 790
rect 57490 810 57495 815
rect 57565 815 57605 820
rect 57565 810 57570 815
rect 57490 790 57570 810
rect 57490 785 57495 790
rect 57455 780 57495 785
rect 57565 785 57570 790
rect 57600 810 57605 815
rect 57675 815 57715 820
rect 57675 810 57680 815
rect 57600 790 57680 810
rect 57600 785 57605 790
rect 57565 780 57605 785
rect 57675 785 57680 790
rect 57710 785 57715 815
rect 57675 780 57715 785
rect 58100 800 58105 830
rect 58135 800 58145 830
rect 58175 800 58185 830
rect 58215 800 58500 830
rect 58530 800 58610 830
rect 58640 800 58720 830
rect 58750 800 58830 830
rect 58860 800 58940 830
rect 58970 800 59050 830
rect 59080 800 59085 830
rect 59430 805 59435 835
rect 59465 830 59470 835
rect 59530 835 59570 840
rect 59530 830 59535 835
rect 59465 810 59535 830
rect 59465 805 59470 810
rect 59430 800 59470 805
rect 59530 805 59535 810
rect 59565 805 59570 835
rect 59530 800 59570 805
rect 58100 790 59085 800
rect 54795 745 55780 755
rect 58100 760 58105 790
rect 58135 760 58145 790
rect 58175 760 58185 790
rect 58215 760 58500 790
rect 58530 760 58610 790
rect 58640 760 58720 790
rect 58750 760 58830 790
rect 58860 760 58940 790
rect 58970 760 59050 790
rect 59080 760 59085 790
rect 58100 750 59085 760
rect 54795 715 54800 745
rect 54830 715 54910 745
rect 54940 715 55020 745
rect 55050 715 55130 745
rect 55160 715 55240 745
rect 55270 715 55350 745
rect 55380 715 55665 745
rect 55695 715 55705 745
rect 55735 715 55745 745
rect 55775 715 55780 745
rect 54795 710 55780 715
rect 56140 745 57660 750
rect 56140 715 56145 745
rect 56175 715 56255 745
rect 56285 715 56365 745
rect 56395 715 56475 745
rect 56505 715 56585 745
rect 56615 715 57185 745
rect 57215 715 57295 745
rect 57325 715 57405 745
rect 57435 715 57515 745
rect 57545 715 57625 745
rect 57655 715 57660 745
rect 58100 720 58105 750
rect 58135 720 58145 750
rect 58175 720 58185 750
rect 58215 720 58500 750
rect 58530 720 58610 750
rect 58640 720 58720 750
rect 58750 720 58830 750
rect 58860 720 58940 750
rect 58970 720 59050 750
rect 59080 720 59085 750
rect 58100 715 59085 720
rect 56140 710 57660 715
rect 53960 690 60110 695
rect 53960 660 53965 690
rect 53995 660 54005 690
rect 54035 660 54045 690
rect 54075 660 54745 690
rect 54775 660 55405 690
rect 55435 660 56035 690
rect 56065 660 56735 690
rect 56765 660 57035 690
rect 57065 660 57735 690
rect 57765 660 58445 690
rect 58475 660 59105 690
rect 59135 660 59995 690
rect 60025 660 60035 690
rect 60065 660 60075 690
rect 60105 660 60110 690
rect 53960 650 60110 660
rect 53960 620 53965 650
rect 53995 620 54005 650
rect 54035 620 54045 650
rect 54075 620 54745 650
rect 54775 620 55405 650
rect 55435 620 56035 650
rect 56065 620 56735 650
rect 56765 620 57035 650
rect 57065 620 57735 650
rect 57765 620 58445 650
rect 58475 620 59105 650
rect 59135 620 59995 650
rect 60025 620 60035 650
rect 60065 620 60075 650
rect 60105 620 60110 650
rect 53960 610 60110 620
rect 53960 580 53965 610
rect 53995 580 54005 610
rect 54035 580 54045 610
rect 54075 580 54745 610
rect 54775 580 55405 610
rect 55435 580 56035 610
rect 56065 580 56735 610
rect 56765 580 57035 610
rect 57065 580 57735 610
rect 57765 580 58445 610
rect 58475 580 59105 610
rect 59135 580 59995 610
rect 60025 580 60035 610
rect 60065 580 60075 610
rect 60105 580 60110 610
rect 53960 575 60110 580
rect 54380 555 54420 560
rect 54380 525 54385 555
rect 54415 550 54420 555
rect 55940 555 55980 560
rect 55940 550 55945 555
rect 54415 530 55945 550
rect 54415 525 54420 530
rect 54380 520 54420 525
rect 55940 525 55945 530
rect 55975 525 55980 555
rect 55940 520 55980 525
rect 57820 555 57860 560
rect 57820 525 57825 555
rect 57855 550 57860 555
rect 59650 555 59690 560
rect 59650 550 59655 555
rect 57855 530 59655 550
rect 57855 525 57860 530
rect 57820 520 57860 525
rect 59650 525 59655 530
rect 59685 525 59690 555
rect 59650 520 59690 525
rect 54515 510 54555 515
rect 54515 480 54520 510
rect 54550 505 54555 510
rect 55100 510 55140 515
rect 55100 505 55105 510
rect 54550 485 55105 505
rect 54550 480 54555 485
rect 54515 475 54555 480
rect 55100 480 55105 485
rect 55135 505 55140 510
rect 58580 510 58620 515
rect 58580 505 58585 510
rect 55135 485 58585 505
rect 55135 480 55140 485
rect 55100 475 55140 480
rect 58580 480 58585 485
rect 58615 505 58620 510
rect 59515 510 59555 515
rect 59515 505 59520 510
rect 58615 485 59520 505
rect 58615 480 58620 485
rect 58580 475 58620 480
rect 59515 480 59520 485
rect 59550 480 59555 510
rect 59515 475 59555 480
rect 56440 390 57470 395
rect 56440 360 56445 390
rect 56475 360 56555 390
rect 56585 360 56665 390
rect 56695 360 56775 390
rect 56805 360 56885 390
rect 56915 360 56995 390
rect 57025 360 57105 390
rect 57135 360 57215 390
rect 57245 360 57325 390
rect 57355 360 57435 390
rect 57465 360 57470 390
rect 56440 355 57470 360
rect 54105 310 55290 315
rect 54105 280 54110 310
rect 54140 280 54150 310
rect 54180 280 54195 310
rect 54225 280 54235 310
rect 54265 280 54280 310
rect 54310 280 54320 310
rect 54350 280 54585 310
rect 54615 280 54855 310
rect 54885 280 54895 310
rect 54925 280 54935 310
rect 54965 280 54975 310
rect 55005 280 55015 310
rect 55045 280 55055 310
rect 55085 280 55095 310
rect 55125 280 55135 310
rect 55165 280 55175 310
rect 55205 280 55215 310
rect 55245 280 55255 310
rect 55285 280 55290 310
rect 54105 270 55290 280
rect 54105 240 54110 270
rect 54140 240 54150 270
rect 54180 240 54195 270
rect 54225 240 54235 270
rect 54265 240 54280 270
rect 54310 240 54320 270
rect 54350 240 54585 270
rect 54615 240 54855 270
rect 54885 240 54895 270
rect 54925 240 54935 270
rect 54965 240 54975 270
rect 55005 240 55015 270
rect 55045 240 55055 270
rect 55085 240 55095 270
rect 55125 240 55135 270
rect 55165 240 55175 270
rect 55205 240 55215 270
rect 55245 240 55255 270
rect 55285 240 55290 270
rect 54105 230 55290 240
rect 54105 200 54110 230
rect 54140 200 54150 230
rect 54180 200 54195 230
rect 54225 200 54235 230
rect 54265 200 54280 230
rect 54310 200 54320 230
rect 54350 200 54585 230
rect 54615 200 54855 230
rect 54885 200 54895 230
rect 54925 200 54935 230
rect 54965 200 54975 230
rect 55005 200 55015 230
rect 55045 200 55055 230
rect 55085 200 55095 230
rect 55125 200 55135 230
rect 55165 200 55175 230
rect 55205 200 55215 230
rect 55245 200 55255 230
rect 55285 200 55290 230
rect 54105 195 55290 200
rect 58430 310 59965 315
rect 58430 280 58435 310
rect 58465 280 58475 310
rect 58505 280 58515 310
rect 58545 280 58555 310
rect 58585 280 58595 310
rect 58625 280 58635 310
rect 58665 280 58675 310
rect 58705 280 58715 310
rect 58745 280 58755 310
rect 58785 280 58795 310
rect 58825 280 58835 310
rect 58865 280 59455 310
rect 59485 280 59720 310
rect 59750 280 59760 310
rect 59790 280 59805 310
rect 59835 280 59845 310
rect 59875 280 59890 310
rect 59920 280 59930 310
rect 59960 280 59965 310
rect 58430 270 59965 280
rect 58430 240 58435 270
rect 58465 240 58475 270
rect 58505 240 58515 270
rect 58545 240 58555 270
rect 58585 240 58595 270
rect 58625 240 58635 270
rect 58665 240 58675 270
rect 58705 240 58715 270
rect 58745 240 58755 270
rect 58785 240 58795 270
rect 58825 240 58835 270
rect 58865 240 59455 270
rect 59485 240 59720 270
rect 59750 240 59760 270
rect 59790 240 59805 270
rect 59835 240 59845 270
rect 59875 240 59890 270
rect 59920 240 59930 270
rect 59960 240 59965 270
rect 58430 230 59965 240
rect 58430 200 58435 230
rect 58465 200 58475 230
rect 58505 200 58515 230
rect 58545 200 58555 230
rect 58585 200 58595 230
rect 58625 200 58635 230
rect 58665 200 58675 230
rect 58705 200 58715 230
rect 58745 200 58755 230
rect 58785 200 58795 230
rect 58825 200 58835 230
rect 58865 200 59455 230
rect 59485 200 59720 230
rect 59750 200 59760 230
rect 59790 200 59805 230
rect 59835 200 59845 230
rect 59875 200 59890 230
rect 59920 200 59930 230
rect 59960 200 59965 230
rect 58430 195 59965 200
rect 54520 175 54555 180
rect 54520 135 54555 140
rect 54580 175 54615 180
rect 54580 135 54615 140
rect 59455 175 59490 180
rect 59455 135 59490 140
rect 59515 175 59550 180
rect 59515 135 59550 140
rect 56220 60 56260 65
rect 56220 30 56225 60
rect 56255 55 56260 60
rect 56275 60 56315 65
rect 56275 55 56280 60
rect 56255 35 56280 55
rect 56255 30 56260 35
rect 56220 25 56260 30
rect 56275 30 56280 35
rect 56310 55 56315 60
rect 56385 60 56425 65
rect 56385 55 56390 60
rect 56310 35 56390 55
rect 56310 30 56315 35
rect 56275 25 56315 30
rect 56385 30 56390 35
rect 56420 55 56425 60
rect 56495 60 56535 65
rect 56495 55 56500 60
rect 56420 35 56500 55
rect 56420 30 56425 35
rect 56385 25 56425 30
rect 56495 30 56500 35
rect 56530 55 56535 60
rect 56605 60 56645 65
rect 56605 55 56610 60
rect 56530 35 56610 55
rect 56530 30 56535 35
rect 56495 25 56535 30
rect 56605 30 56610 35
rect 56640 55 56645 60
rect 56715 60 56755 65
rect 56715 55 56720 60
rect 56640 35 56720 55
rect 56640 30 56645 35
rect 56605 25 56645 30
rect 56715 30 56720 35
rect 56750 55 56755 60
rect 56825 60 56865 65
rect 56825 55 56830 60
rect 56750 35 56830 55
rect 56750 30 56755 35
rect 56715 25 56755 30
rect 56825 30 56830 35
rect 56860 55 56865 60
rect 56935 60 56975 65
rect 56935 55 56940 60
rect 56860 35 56940 55
rect 56860 30 56865 35
rect 56825 25 56865 30
rect 56935 30 56940 35
rect 56970 55 56975 60
rect 57045 60 57085 65
rect 57045 55 57050 60
rect 56970 35 57050 55
rect 56970 30 56975 35
rect 56935 25 56975 30
rect 57045 30 57050 35
rect 57080 55 57085 60
rect 57155 60 57195 65
rect 57155 55 57160 60
rect 57080 35 57160 55
rect 57080 30 57085 35
rect 57045 25 57085 30
rect 57155 30 57160 35
rect 57190 55 57195 60
rect 57265 60 57305 65
rect 57265 55 57270 60
rect 57190 35 57270 55
rect 57190 30 57195 35
rect 57155 25 57195 30
rect 57265 30 57270 35
rect 57300 55 57305 60
rect 57375 60 57415 65
rect 57375 55 57380 60
rect 57300 35 57380 55
rect 57300 30 57305 35
rect 57265 25 57305 30
rect 57375 30 57380 35
rect 57410 55 57415 60
rect 57485 60 57525 65
rect 57485 55 57490 60
rect 57410 35 57490 55
rect 57410 30 57415 35
rect 57375 25 57415 30
rect 57485 30 57490 35
rect 57520 30 57525 60
rect 57485 25 57525 30
rect 56440 15 56480 20
rect 56440 -15 56445 15
rect 56475 10 56480 15
rect 56550 15 56590 20
rect 56550 10 56555 15
rect 56475 -10 56555 10
rect 56475 -15 56480 -10
rect 56440 -20 56480 -15
rect 56550 -15 56555 -10
rect 56585 10 56590 15
rect 56660 15 56700 20
rect 56660 10 56665 15
rect 56585 -10 56665 10
rect 56585 -15 56590 -10
rect 56550 -20 56590 -15
rect 56660 -15 56665 -10
rect 56695 10 56700 15
rect 56770 15 56810 20
rect 56770 10 56775 15
rect 56695 -10 56775 10
rect 56695 -15 56700 -10
rect 56660 -20 56700 -15
rect 56770 -15 56775 -10
rect 56805 10 56810 15
rect 56880 15 56920 20
rect 56880 10 56885 15
rect 56805 -10 56885 10
rect 56805 -15 56810 -10
rect 56770 -20 56810 -15
rect 56880 -15 56885 -10
rect 56915 10 56920 15
rect 56990 15 57030 20
rect 56990 10 56995 15
rect 56915 -10 56995 10
rect 56915 -15 56920 -10
rect 56880 -20 56920 -15
rect 56990 -15 56995 -10
rect 57025 10 57030 15
rect 57100 15 57140 20
rect 57100 10 57105 15
rect 57025 -10 57105 10
rect 57025 -15 57030 -10
rect 56990 -20 57030 -15
rect 57100 -15 57105 -10
rect 57135 10 57140 15
rect 57210 15 57250 20
rect 57210 10 57215 15
rect 57135 -10 57215 10
rect 57135 -15 57140 -10
rect 57100 -20 57140 -15
rect 57210 -15 57215 -10
rect 57245 10 57250 15
rect 57320 15 57360 20
rect 57320 10 57325 15
rect 57245 -10 57325 10
rect 57245 -15 57250 -10
rect 57210 -20 57250 -15
rect 57320 -15 57325 -10
rect 57355 10 57360 15
rect 57430 15 57470 20
rect 57430 10 57435 15
rect 57355 -10 57435 10
rect 57355 -15 57360 -10
rect 57320 -20 57360 -15
rect 57430 -15 57435 -10
rect 57465 -15 57470 15
rect 57430 -20 57470 -15
rect 57415 -40 57455 -35
rect 57415 -70 57420 -40
rect 57450 -45 57455 -40
rect 57865 -40 57905 -35
rect 57865 -45 57870 -40
rect 57450 -65 57870 -45
rect 57450 -70 57455 -65
rect 57415 -75 57455 -70
rect 57865 -70 57870 -65
rect 57900 -70 57905 -40
rect 57865 -75 57905 -70
rect 55795 -95 58040 -90
rect 55795 -125 55800 -95
rect 55830 -125 55840 -95
rect 55870 -125 56335 -95
rect 56365 -125 57925 -95
rect 57955 -125 57965 -95
rect 57995 -125 58005 -95
rect 58035 -125 58040 -95
rect 55795 -135 58040 -125
rect 55795 -165 55800 -135
rect 55830 -165 55840 -135
rect 55870 -165 56335 -135
rect 56365 -165 57925 -135
rect 57955 -165 57965 -135
rect 57995 -165 58005 -135
rect 58035 -165 58040 -135
rect 55795 -175 58040 -165
rect 55795 -205 55800 -175
rect 55830 -205 55840 -175
rect 55870 -205 56335 -175
rect 56365 -205 57925 -175
rect 57955 -205 57965 -175
rect 57995 -205 58005 -175
rect 58035 -205 58040 -175
rect 55795 -210 58040 -205
rect 56540 -230 56580 -225
rect 56540 -260 56545 -230
rect 56575 -235 56580 -230
rect 56650 -230 56690 -225
rect 56650 -235 56655 -230
rect 56575 -255 56655 -235
rect 56575 -260 56580 -255
rect 56540 -265 56580 -260
rect 56650 -260 56655 -255
rect 56685 -235 56690 -230
rect 56870 -230 56910 -225
rect 56870 -235 56875 -230
rect 56685 -255 56875 -235
rect 56685 -260 56690 -255
rect 56650 -265 56690 -260
rect 56870 -260 56875 -255
rect 56905 -260 56910 -230
rect 56870 -265 56910 -260
rect 55895 -275 55935 -270
rect 55895 -305 55900 -275
rect 55930 -280 55935 -275
rect 56485 -275 56525 -270
rect 56485 -280 56490 -275
rect 55930 -300 56490 -280
rect 55930 -305 55935 -300
rect 55895 -310 55935 -305
rect 56485 -305 56490 -300
rect 56520 -280 56525 -275
rect 56595 -275 56635 -270
rect 56595 -280 56600 -275
rect 56520 -300 56600 -280
rect 56520 -305 56525 -300
rect 56485 -310 56525 -305
rect 56595 -305 56600 -300
rect 56630 -280 56635 -275
rect 56705 -275 56745 -270
rect 56705 -280 56710 -275
rect 56630 -300 56710 -280
rect 56630 -305 56635 -300
rect 56595 -310 56635 -305
rect 56705 -305 56710 -300
rect 56740 -280 56745 -275
rect 57040 -275 57080 -270
rect 57040 -280 57045 -275
rect 56740 -300 57045 -280
rect 56740 -305 56745 -300
rect 56705 -310 56745 -305
rect 57040 -305 57045 -300
rect 57075 -305 57080 -275
rect 57040 -310 57080 -305
rect 56540 -480 56580 -475
rect 56540 -510 56545 -480
rect 56575 -485 56580 -480
rect 56650 -480 56690 -475
rect 56650 -485 56655 -480
rect 56575 -505 56655 -485
rect 56575 -510 56580 -505
rect 56540 -515 56580 -510
rect 56650 -510 56655 -505
rect 56685 -485 56690 -480
rect 56870 -480 56910 -475
rect 56870 -485 56875 -480
rect 56685 -505 56875 -485
rect 56685 -510 56690 -505
rect 56650 -515 56690 -510
rect 56870 -510 56875 -505
rect 56905 -510 56910 -480
rect 56870 -515 56910 -510
rect 54850 -525 55290 -520
rect 54850 -555 54855 -525
rect 54885 -555 55055 -525
rect 55085 -555 55255 -525
rect 55285 -555 55290 -525
rect 54850 -560 55290 -555
rect 56485 -525 56525 -520
rect 56485 -555 56490 -525
rect 56520 -530 56525 -525
rect 56595 -525 56635 -520
rect 56595 -530 56600 -525
rect 56520 -550 56600 -530
rect 56520 -555 56525 -550
rect 56485 -560 56525 -555
rect 56595 -555 56600 -550
rect 56630 -530 56635 -525
rect 56705 -525 56745 -520
rect 56705 -530 56710 -525
rect 56630 -550 56710 -530
rect 56630 -555 56635 -550
rect 56595 -560 56635 -555
rect 56705 -555 56710 -550
rect 56740 -555 56745 -525
rect 56705 -560 56745 -555
rect 58430 -525 58870 -520
rect 58430 -555 58435 -525
rect 58465 -555 58635 -525
rect 58665 -555 58835 -525
rect 58865 -555 58870 -525
rect 58430 -560 58870 -555
rect 52290 -580 61510 -575
rect 52290 -610 52295 -580
rect 52325 -610 52335 -580
rect 52365 -610 52375 -580
rect 52405 -610 52645 -580
rect 52675 -610 52685 -580
rect 52715 -610 52725 -580
rect 52755 -610 52995 -580
rect 53025 -610 53035 -580
rect 53065 -610 53075 -580
rect 53105 -610 53345 -580
rect 53375 -610 53385 -580
rect 53415 -610 53425 -580
rect 53455 -610 53965 -580
rect 53995 -610 54005 -580
rect 54035 -610 54045 -580
rect 54075 -610 54395 -580
rect 54425 -610 54435 -580
rect 54465 -610 54475 -580
rect 54505 -610 54745 -580
rect 54775 -610 54785 -580
rect 54815 -610 54825 -580
rect 54855 -610 55035 -580
rect 55065 -610 55095 -580
rect 55125 -610 55135 -580
rect 55165 -610 55175 -580
rect 55205 -610 55235 -580
rect 55265 -610 55445 -580
rect 55475 -610 55485 -580
rect 55515 -610 55525 -580
rect 55555 -610 55795 -580
rect 55825 -610 55835 -580
rect 55865 -610 55875 -580
rect 55905 -610 56145 -580
rect 56175 -610 56185 -580
rect 56215 -610 56225 -580
rect 56255 -610 56435 -580
rect 56465 -610 56495 -580
rect 56525 -610 56535 -580
rect 56565 -610 56575 -580
rect 56605 -610 56765 -580
rect 56795 -610 56845 -580
rect 56875 -610 56885 -580
rect 56915 -610 56925 -580
rect 56955 -610 57195 -580
rect 57225 -610 57235 -580
rect 57265 -610 57275 -580
rect 57305 -610 57490 -580
rect 57520 -610 57545 -580
rect 57575 -610 57585 -580
rect 57615 -610 57625 -580
rect 57655 -610 57895 -580
rect 57925 -610 57935 -580
rect 57965 -610 57975 -580
rect 58005 -610 58245 -580
rect 58275 -610 58285 -580
rect 58315 -610 58325 -580
rect 58355 -610 58535 -580
rect 58565 -610 58595 -580
rect 58625 -610 58635 -580
rect 58665 -610 58675 -580
rect 58705 -610 58735 -580
rect 58765 -610 58945 -580
rect 58975 -610 58985 -580
rect 59015 -610 59025 -580
rect 59055 -610 59295 -580
rect 59325 -610 59335 -580
rect 59365 -610 59375 -580
rect 59405 -610 59645 -580
rect 59675 -610 59685 -580
rect 59715 -610 59725 -580
rect 59755 -610 59995 -580
rect 60025 -610 60035 -580
rect 60065 -610 60075 -580
rect 60105 -610 60345 -580
rect 60375 -610 60385 -580
rect 60415 -610 60425 -580
rect 60455 -610 60695 -580
rect 60725 -610 60735 -580
rect 60765 -610 60775 -580
rect 60805 -610 61045 -580
rect 61075 -610 61085 -580
rect 61115 -610 61125 -580
rect 61155 -610 61395 -580
rect 61425 -610 61435 -580
rect 61465 -610 61475 -580
rect 61505 -610 61510 -580
rect 52290 -620 61510 -610
rect 52290 -650 52295 -620
rect 52325 -650 52335 -620
rect 52365 -650 52375 -620
rect 52405 -650 52645 -620
rect 52675 -650 52685 -620
rect 52715 -650 52725 -620
rect 52755 -650 52995 -620
rect 53025 -650 53035 -620
rect 53065 -650 53075 -620
rect 53105 -650 53345 -620
rect 53375 -650 53385 -620
rect 53415 -650 53425 -620
rect 53455 -650 53965 -620
rect 53995 -650 54005 -620
rect 54035 -650 54045 -620
rect 54075 -650 54395 -620
rect 54425 -650 54435 -620
rect 54465 -650 54475 -620
rect 54505 -650 54745 -620
rect 54775 -650 54785 -620
rect 54815 -650 54825 -620
rect 54855 -650 55035 -620
rect 55065 -650 55095 -620
rect 55125 -650 55135 -620
rect 55165 -650 55175 -620
rect 55205 -650 55235 -620
rect 55265 -650 55445 -620
rect 55475 -650 55485 -620
rect 55515 -650 55525 -620
rect 55555 -650 55795 -620
rect 55825 -650 55835 -620
rect 55865 -650 55875 -620
rect 55905 -650 56145 -620
rect 56175 -650 56185 -620
rect 56215 -650 56225 -620
rect 56255 -650 56435 -620
rect 56465 -650 56495 -620
rect 56525 -650 56535 -620
rect 56565 -650 56575 -620
rect 56605 -650 56765 -620
rect 56795 -650 56845 -620
rect 56875 -650 56885 -620
rect 56915 -650 56925 -620
rect 56955 -650 57195 -620
rect 57225 -650 57235 -620
rect 57265 -650 57275 -620
rect 57305 -650 57490 -620
rect 57520 -650 57545 -620
rect 57575 -650 57585 -620
rect 57615 -650 57625 -620
rect 57655 -650 57895 -620
rect 57925 -650 57935 -620
rect 57965 -650 57975 -620
rect 58005 -650 58245 -620
rect 58275 -650 58285 -620
rect 58315 -650 58325 -620
rect 58355 -650 58535 -620
rect 58565 -650 58595 -620
rect 58625 -650 58635 -620
rect 58665 -650 58675 -620
rect 58705 -650 58735 -620
rect 58765 -650 58945 -620
rect 58975 -650 58985 -620
rect 59015 -650 59025 -620
rect 59055 -650 59295 -620
rect 59325 -650 59335 -620
rect 59365 -650 59375 -620
rect 59405 -650 59645 -620
rect 59675 -650 59685 -620
rect 59715 -650 59725 -620
rect 59755 -650 59995 -620
rect 60025 -650 60035 -620
rect 60065 -650 60075 -620
rect 60105 -650 60345 -620
rect 60375 -650 60385 -620
rect 60415 -650 60425 -620
rect 60455 -650 60695 -620
rect 60725 -650 60735 -620
rect 60765 -650 60775 -620
rect 60805 -650 61045 -620
rect 61075 -650 61085 -620
rect 61115 -650 61125 -620
rect 61155 -650 61395 -620
rect 61425 -650 61435 -620
rect 61465 -650 61475 -620
rect 61505 -650 61510 -620
rect 52290 -660 61510 -650
rect 52290 -690 52295 -660
rect 52325 -690 52335 -660
rect 52365 -690 52375 -660
rect 52405 -690 52645 -660
rect 52675 -690 52685 -660
rect 52715 -690 52725 -660
rect 52755 -690 52995 -660
rect 53025 -690 53035 -660
rect 53065 -690 53075 -660
rect 53105 -690 53345 -660
rect 53375 -690 53385 -660
rect 53415 -690 53425 -660
rect 53455 -690 53965 -660
rect 53995 -690 54005 -660
rect 54035 -690 54045 -660
rect 54075 -690 54395 -660
rect 54425 -690 54435 -660
rect 54465 -690 54475 -660
rect 54505 -690 54745 -660
rect 54775 -690 54785 -660
rect 54815 -690 54825 -660
rect 54855 -690 55035 -660
rect 55065 -690 55095 -660
rect 55125 -690 55135 -660
rect 55165 -690 55175 -660
rect 55205 -690 55235 -660
rect 55265 -690 55445 -660
rect 55475 -690 55485 -660
rect 55515 -690 55525 -660
rect 55555 -690 55795 -660
rect 55825 -690 55835 -660
rect 55865 -690 55875 -660
rect 55905 -690 56145 -660
rect 56175 -690 56185 -660
rect 56215 -690 56225 -660
rect 56255 -690 56435 -660
rect 56465 -690 56495 -660
rect 56525 -690 56535 -660
rect 56565 -690 56575 -660
rect 56605 -690 56765 -660
rect 56795 -690 56845 -660
rect 56875 -690 56885 -660
rect 56915 -690 56925 -660
rect 56955 -690 57195 -660
rect 57225 -690 57235 -660
rect 57265 -690 57275 -660
rect 57305 -690 57490 -660
rect 57520 -690 57545 -660
rect 57575 -690 57585 -660
rect 57615 -690 57625 -660
rect 57655 -690 57895 -660
rect 57925 -690 57935 -660
rect 57965 -690 57975 -660
rect 58005 -690 58245 -660
rect 58275 -690 58285 -660
rect 58315 -690 58325 -660
rect 58355 -690 58535 -660
rect 58565 -690 58595 -660
rect 58625 -690 58635 -660
rect 58665 -690 58675 -660
rect 58705 -690 58735 -660
rect 58765 -690 58945 -660
rect 58975 -690 58985 -660
rect 59015 -690 59025 -660
rect 59055 -690 59295 -660
rect 59325 -690 59335 -660
rect 59365 -690 59375 -660
rect 59405 -690 59645 -660
rect 59675 -690 59685 -660
rect 59715 -690 59725 -660
rect 59755 -690 59995 -660
rect 60025 -690 60035 -660
rect 60065 -690 60075 -660
rect 60105 -690 60345 -660
rect 60375 -690 60385 -660
rect 60415 -690 60425 -660
rect 60455 -690 60695 -660
rect 60725 -690 60735 -660
rect 60765 -690 60775 -660
rect 60805 -690 61045 -660
rect 61075 -690 61085 -660
rect 61115 -690 61125 -660
rect 61155 -690 61395 -660
rect 61425 -690 61435 -660
rect 61465 -690 61475 -660
rect 61505 -690 61510 -660
rect 52290 -695 61510 -690
<< via2 >>
rect 54180 3095 54210 3125
rect 59860 3095 59890 3125
rect 54115 1330 54145 1360
rect 54165 1330 54195 1360
rect 54215 1330 54245 1360
rect 54265 1330 54295 1360
rect 54315 1330 54345 1360
rect 59725 1405 59755 1435
rect 59775 1405 59805 1435
rect 59825 1405 59855 1435
rect 59875 1405 59905 1435
rect 59925 1405 59955 1435
rect 59725 1355 59755 1385
rect 59775 1355 59805 1385
rect 59825 1355 59855 1385
rect 59875 1355 59905 1385
rect 59925 1355 59955 1385
rect 54115 1280 54145 1310
rect 54165 1280 54195 1310
rect 54215 1280 54245 1310
rect 54265 1280 54295 1310
rect 54315 1280 54345 1310
rect 59725 1305 59755 1335
rect 59775 1305 59805 1335
rect 59825 1305 59855 1335
rect 59875 1305 59905 1335
rect 59925 1305 59955 1335
rect 54115 1230 54145 1260
rect 54165 1230 54195 1260
rect 54215 1230 54245 1260
rect 54265 1230 54295 1260
rect 54315 1230 54345 1260
<< metal3 >>
rect 52060 6220 52290 6305
rect 52410 6220 52640 6305
rect 52760 6220 52990 6305
rect 52060 6170 52990 6220
rect 52060 6075 52290 6170
rect 52410 6075 52640 6170
rect 52760 6075 52990 6170
rect 53110 6075 53340 6305
rect 53460 6075 53690 6305
rect 53810 6075 54040 6305
rect 54160 6075 54390 6305
rect 54510 6075 54740 6305
rect 54860 6075 55090 6305
rect 55210 6075 55440 6305
rect 55560 6075 55790 6305
rect 55910 6075 56140 6305
rect 56260 6075 56490 6305
rect 56610 6075 56840 6305
rect 56960 6075 57190 6305
rect 57310 6075 57540 6305
rect 57660 6075 57890 6305
rect 58010 6075 58240 6305
rect 58360 6075 58590 6305
rect 58710 6075 58940 6305
rect 59060 6075 59290 6305
rect 59410 6075 59640 6305
rect 59760 6075 59990 6305
rect 60110 6075 60340 6305
rect 60460 6075 60690 6305
rect 60810 6220 61040 6305
rect 61160 6220 61390 6305
rect 61510 6220 61740 6305
rect 60810 6170 61740 6220
rect 60810 6075 61040 6170
rect 61160 6075 61390 6170
rect 61510 6075 61740 6170
rect 52850 5955 52900 6075
rect 53200 5955 53250 6075
rect 53550 5955 53600 6075
rect 53900 5955 53950 6075
rect 54250 5955 54300 6075
rect 54600 5955 54650 6075
rect 54950 5955 55000 6075
rect 55300 5955 55350 6075
rect 55650 5955 55700 6075
rect 56000 5955 56050 6075
rect 56350 5955 56400 6075
rect 56700 5955 56750 6075
rect 57050 5955 57100 6075
rect 57400 5955 57450 6075
rect 57750 5955 57800 6075
rect 58100 5955 58150 6075
rect 58450 5955 58500 6075
rect 58800 5955 58850 6075
rect 59150 5955 59200 6075
rect 59500 5955 59550 6075
rect 59850 5955 59900 6075
rect 60200 5955 60250 6075
rect 60550 5955 60600 6075
rect 60900 5955 60950 6075
rect 52060 5870 52290 5955
rect 52410 5870 52640 5955
rect 52760 5870 52990 5955
rect 53110 5870 53340 5955
rect 53460 5870 53690 5955
rect 53810 5870 54040 5955
rect 54160 5870 54390 5955
rect 54510 5870 54740 5955
rect 54860 5870 55090 5955
rect 55210 5870 55440 5955
rect 55560 5870 55790 5955
rect 55910 5870 56140 5955
rect 56260 5870 56490 5955
rect 56610 5870 56840 5955
rect 52060 5820 56840 5870
rect 52060 5725 52290 5820
rect 52410 5725 52640 5820
rect 52760 5725 52990 5820
rect 53110 5725 53340 5820
rect 53460 5725 53690 5820
rect 53810 5725 54040 5820
rect 54160 5725 54390 5820
rect 54510 5725 54740 5820
rect 54860 5725 55090 5820
rect 55210 5725 55440 5820
rect 55560 5725 55790 5820
rect 55910 5725 56140 5820
rect 56260 5725 56490 5820
rect 56610 5725 56840 5820
rect 56960 5870 57190 5955
rect 57310 5870 57540 5955
rect 57660 5870 57890 5955
rect 58010 5870 58240 5955
rect 58360 5870 58590 5955
rect 58710 5870 58940 5955
rect 59060 5870 59290 5955
rect 59410 5870 59640 5955
rect 59760 5870 59990 5955
rect 60110 5870 60340 5955
rect 60460 5870 60690 5955
rect 60810 5870 61040 5955
rect 61160 5870 61390 5955
rect 61510 5870 61740 5955
rect 56960 5820 61740 5870
rect 56960 5725 57190 5820
rect 57310 5725 57540 5820
rect 57660 5725 57890 5820
rect 58010 5725 58240 5820
rect 58360 5725 58590 5820
rect 58710 5725 58940 5820
rect 59060 5725 59290 5820
rect 59410 5725 59640 5820
rect 59760 5725 59990 5820
rect 60110 5725 60340 5820
rect 60460 5725 60690 5820
rect 60810 5725 61040 5820
rect 61160 5725 61390 5820
rect 61510 5725 61740 5820
rect 52850 5605 52900 5725
rect 53900 5605 53950 5725
rect 54250 5605 54300 5725
rect 54600 5605 54650 5725
rect 54950 5605 55000 5725
rect 55300 5605 55350 5725
rect 55650 5605 55700 5725
rect 56000 5605 56050 5725
rect 56350 5605 56400 5725
rect 56700 5605 56750 5725
rect 57050 5605 57100 5725
rect 57400 5605 57450 5725
rect 57750 5605 57800 5725
rect 58100 5605 58150 5725
rect 58450 5605 58500 5725
rect 58800 5605 58850 5725
rect 59150 5605 59200 5725
rect 59500 5605 59550 5725
rect 59850 5605 59900 5725
rect 60900 5605 60950 5725
rect 52060 5520 52290 5605
rect 52410 5520 52640 5605
rect 52760 5520 52990 5605
rect 53110 5520 53340 5605
rect 53460 5520 53690 5605
rect 52060 5470 53690 5520
rect 52060 5375 52290 5470
rect 52410 5375 52640 5470
rect 52760 5375 52990 5470
rect 53110 5375 53340 5470
rect 53460 5375 53690 5470
rect 53810 5375 54040 5605
rect 54160 5375 54390 5605
rect 54510 5375 54740 5605
rect 54860 5375 55090 5605
rect 55210 5375 55440 5605
rect 55560 5375 55790 5605
rect 55910 5375 56140 5605
rect 56260 5375 56490 5605
rect 56610 5375 56840 5605
rect 56960 5375 57190 5605
rect 57310 5375 57540 5605
rect 57660 5375 57890 5605
rect 58010 5375 58240 5605
rect 58360 5375 58590 5605
rect 58710 5375 58940 5605
rect 59060 5375 59290 5605
rect 59410 5375 59640 5605
rect 59760 5375 59990 5605
rect 60110 5520 60340 5605
rect 60460 5520 60690 5605
rect 60810 5520 61040 5605
rect 61160 5520 61390 5605
rect 61510 5520 61740 5605
rect 60110 5470 61740 5520
rect 60110 5375 60340 5470
rect 60460 5375 60690 5470
rect 60810 5375 61040 5470
rect 61160 5375 61390 5470
rect 61510 5375 61740 5470
rect 52850 5255 52900 5375
rect 53900 5255 53950 5375
rect 54250 5255 54300 5375
rect 54600 5255 54650 5375
rect 59150 5255 59200 5375
rect 59500 5255 59550 5375
rect 59850 5255 59900 5375
rect 60900 5255 60950 5375
rect 52060 5170 52290 5255
rect 52410 5170 52640 5255
rect 52760 5170 52990 5255
rect 53110 5170 53340 5255
rect 53460 5170 53690 5255
rect 52060 5120 53690 5170
rect 52060 5025 52290 5120
rect 52410 5025 52640 5120
rect 52760 5025 52990 5120
rect 53110 5025 53340 5120
rect 53460 5025 53690 5120
rect 53810 5025 54040 5255
rect 54160 5025 54390 5255
rect 54510 5025 54740 5255
rect 59060 5025 59290 5255
rect 59410 5025 59640 5255
rect 59760 5025 59990 5255
rect 60110 5170 60340 5255
rect 60460 5170 60690 5255
rect 60810 5170 61040 5255
rect 61160 5170 61390 5255
rect 61510 5170 61740 5255
rect 60110 5120 61740 5170
rect 60110 5025 60340 5120
rect 60460 5025 60690 5120
rect 60810 5025 61040 5120
rect 61160 5025 61390 5120
rect 61510 5025 61740 5120
rect 52850 4905 52900 5025
rect 52060 4820 52290 4905
rect 52410 4820 52640 4905
rect 52760 4820 52990 4905
rect 53110 4820 53340 4905
rect 53460 4820 53690 4905
rect 52060 4770 53690 4820
rect 52060 4675 52290 4770
rect 52410 4675 52640 4770
rect 52760 4675 52990 4770
rect 53110 4675 53340 4770
rect 53460 4675 53690 4770
rect 52850 4555 52900 4675
rect 52060 4470 52290 4555
rect 52410 4470 52640 4555
rect 52760 4470 52990 4555
rect 53110 4470 53340 4555
rect 53460 4470 53690 4555
rect 52060 4420 53690 4470
rect 52060 4325 52290 4420
rect 52410 4325 52640 4420
rect 52760 4325 52990 4420
rect 53110 4325 53340 4420
rect 53460 4325 53690 4420
rect 52850 4205 52900 4325
rect 52060 4120 52290 4205
rect 52410 4120 52640 4205
rect 52760 4120 52990 4205
rect 53110 4120 53340 4205
rect 53460 4120 53690 4205
rect 52060 4070 53690 4120
rect 53905 4090 53945 5025
rect 52060 3975 52290 4070
rect 52410 3975 52640 4070
rect 52760 3975 52990 4070
rect 53110 3975 53340 4070
rect 53460 3975 53690 4070
rect 52850 3855 52900 3975
rect 52060 3770 52290 3855
rect 52410 3770 52640 3855
rect 52760 3770 52990 3855
rect 53110 3770 53340 3855
rect 53460 3770 53690 3855
rect 52060 3720 53690 3770
rect 52060 3625 52290 3720
rect 52410 3625 52640 3720
rect 52760 3625 52990 3720
rect 53110 3625 53340 3720
rect 53460 3625 53690 3720
rect 52850 3505 52900 3625
rect 52060 3420 52290 3505
rect 52410 3420 52640 3505
rect 52760 3420 52990 3505
rect 53110 3420 53340 3505
rect 53460 3420 53690 3505
rect 52060 3370 53690 3420
rect 52060 3275 52290 3370
rect 52410 3275 52640 3370
rect 52760 3275 52990 3370
rect 53110 3275 53340 3370
rect 53460 3275 53690 3370
rect 52850 3155 52900 3275
rect 52060 3070 52290 3155
rect 52410 3070 52640 3155
rect 52760 3070 52990 3155
rect 53110 3070 53340 3155
rect 53460 3070 53690 3155
rect 54175 3125 54215 4325
rect 54175 3095 54180 3125
rect 54210 3095 54215 3125
rect 54175 3090 54215 3095
rect 59855 3125 59895 5025
rect 60900 4905 60950 5025
rect 60110 4820 60340 4905
rect 60460 4820 60690 4905
rect 60810 4820 61040 4905
rect 61160 4820 61390 4905
rect 61510 4820 61740 4905
rect 60110 4770 61740 4820
rect 60110 4675 60340 4770
rect 60460 4675 60690 4770
rect 60810 4675 61040 4770
rect 61160 4675 61390 4770
rect 61510 4675 61740 4770
rect 60900 4555 60950 4675
rect 60110 4470 60340 4555
rect 60460 4470 60690 4555
rect 60810 4470 61040 4555
rect 61160 4470 61390 4555
rect 61510 4470 61740 4555
rect 60110 4420 61740 4470
rect 60110 4325 60340 4420
rect 60460 4325 60690 4420
rect 60810 4325 61040 4420
rect 61160 4325 61390 4420
rect 61510 4325 61740 4420
rect 60900 4205 60950 4325
rect 60110 4120 60340 4205
rect 60460 4120 60690 4205
rect 60810 4120 61040 4205
rect 61160 4120 61390 4205
rect 61510 4120 61740 4205
rect 60110 4070 61740 4120
rect 60110 3975 60340 4070
rect 60460 3975 60690 4070
rect 60810 3975 61040 4070
rect 61160 3975 61390 4070
rect 61510 3975 61740 4070
rect 60900 3855 60950 3975
rect 60110 3770 60340 3855
rect 60460 3770 60690 3855
rect 60810 3770 61040 3855
rect 61160 3770 61390 3855
rect 61510 3770 61740 3855
rect 60110 3720 61740 3770
rect 60110 3625 60340 3720
rect 60460 3625 60690 3720
rect 60810 3625 61040 3720
rect 61160 3625 61390 3720
rect 61510 3625 61740 3720
rect 60900 3505 60950 3625
rect 60110 3420 60340 3505
rect 60460 3420 60690 3505
rect 60810 3420 61040 3505
rect 61160 3420 61390 3505
rect 61510 3420 61740 3505
rect 60110 3370 61740 3420
rect 60110 3275 60340 3370
rect 60460 3275 60690 3370
rect 60810 3275 61040 3370
rect 61160 3275 61390 3370
rect 61510 3275 61740 3370
rect 60900 3155 60950 3275
rect 59855 3095 59860 3125
rect 59890 3095 59895 3125
rect 59855 3090 59895 3095
rect 52060 3020 53690 3070
rect 52060 2925 52290 3020
rect 52410 2925 52640 3020
rect 52760 2925 52990 3020
rect 53110 2925 53340 3020
rect 53460 2925 53690 3020
rect 60110 3070 60340 3155
rect 60460 3070 60690 3155
rect 60810 3070 61040 3155
rect 61160 3070 61390 3155
rect 61510 3070 61740 3155
rect 60110 3020 61740 3070
rect 60110 2925 60340 3020
rect 60460 2925 60690 3020
rect 60810 2925 61040 3020
rect 61160 2925 61390 3020
rect 61510 2925 61740 3020
rect 52850 2805 52900 2925
rect 60900 2805 60950 2925
rect 52060 2720 52290 2805
rect 52410 2720 52640 2805
rect 52760 2720 52990 2805
rect 53110 2720 53340 2805
rect 53460 2720 53690 2805
rect 52060 2670 53690 2720
rect 52060 2575 52290 2670
rect 52410 2575 52640 2670
rect 52760 2575 52990 2670
rect 53110 2575 53340 2670
rect 53460 2575 53690 2670
rect 60110 2720 60340 2805
rect 60460 2720 60690 2805
rect 60810 2720 61040 2805
rect 61160 2720 61390 2805
rect 61510 2720 61740 2805
rect 60110 2670 61740 2720
rect 60110 2575 60340 2670
rect 60460 2575 60690 2670
rect 60810 2575 61040 2670
rect 61160 2575 61390 2670
rect 61510 2575 61740 2670
rect 52850 2455 52900 2575
rect 60900 2455 60950 2575
rect 52060 2370 52290 2455
rect 52410 2370 52640 2455
rect 52760 2370 52990 2455
rect 53110 2370 53340 2455
rect 53460 2370 53690 2455
rect 52060 2320 53690 2370
rect 52060 2225 52290 2320
rect 52410 2225 52640 2320
rect 52760 2225 52990 2320
rect 53110 2225 53340 2320
rect 53460 2225 53690 2320
rect 60110 2370 60340 2455
rect 60460 2370 60690 2455
rect 60810 2370 61040 2455
rect 61160 2370 61390 2455
rect 61510 2370 61740 2455
rect 60110 2320 61740 2370
rect 60110 2225 60340 2320
rect 60460 2225 60690 2320
rect 60810 2225 61040 2320
rect 61160 2225 61390 2320
rect 61510 2225 61740 2320
rect 52850 2105 52900 2225
rect 60900 2105 60950 2225
rect 52060 2020 52290 2105
rect 52410 2020 52640 2105
rect 52760 2020 52990 2105
rect 53110 2020 53340 2105
rect 53460 2020 53690 2105
rect 52060 1970 53690 2020
rect 52060 1875 52290 1970
rect 52410 1875 52640 1970
rect 52760 1875 52990 1970
rect 53110 1875 53340 1970
rect 53460 1875 53690 1970
rect 60110 2020 60340 2105
rect 60460 2020 60690 2105
rect 60810 2020 61040 2105
rect 61160 2020 61390 2105
rect 61510 2020 61740 2105
rect 60110 1970 61740 2020
rect 60110 1875 60340 1970
rect 60460 1875 60690 1970
rect 60810 1875 61040 1970
rect 61160 1875 61390 1970
rect 61510 1875 61740 1970
rect 52850 1755 52900 1875
rect 60900 1755 60950 1875
rect 52060 1670 52290 1755
rect 52410 1670 52640 1755
rect 52760 1670 52990 1755
rect 53110 1670 53340 1755
rect 53460 1670 53690 1755
rect 52060 1620 53690 1670
rect 52060 1525 52290 1620
rect 52410 1525 52640 1620
rect 52760 1525 52990 1620
rect 53110 1525 53340 1620
rect 53460 1525 53690 1620
rect 60110 1670 60340 1755
rect 60460 1670 60690 1755
rect 60810 1670 61040 1755
rect 61160 1670 61390 1755
rect 61510 1670 61740 1755
rect 60110 1620 61740 1670
rect 60110 1525 60340 1620
rect 60460 1525 60690 1620
rect 60810 1525 61040 1620
rect 61160 1525 61390 1620
rect 61510 1525 61740 1620
rect 52850 1405 52900 1525
rect 59715 1440 59965 1445
rect 52060 1320 52290 1405
rect 52410 1320 52640 1405
rect 52760 1320 52990 1405
rect 53110 1320 53340 1405
rect 53460 1320 53690 1405
rect 59715 1400 59720 1440
rect 59760 1400 59770 1440
rect 59810 1400 59820 1440
rect 59860 1400 59870 1440
rect 59910 1400 59920 1440
rect 59960 1400 59965 1440
rect 60900 1405 60950 1525
rect 59715 1390 59965 1400
rect 52060 1270 53690 1320
rect 52060 1175 52290 1270
rect 52410 1175 52640 1270
rect 52760 1175 52990 1270
rect 53110 1175 53340 1270
rect 53460 1175 53690 1270
rect 54105 1365 54355 1370
rect 54105 1325 54110 1365
rect 54150 1325 54160 1365
rect 54200 1325 54210 1365
rect 54250 1325 54260 1365
rect 54300 1325 54310 1365
rect 54350 1325 54355 1365
rect 54105 1315 54355 1325
rect 54105 1275 54110 1315
rect 54150 1275 54160 1315
rect 54200 1275 54210 1315
rect 54250 1275 54260 1315
rect 54300 1275 54310 1315
rect 54350 1275 54355 1315
rect 59715 1350 59720 1390
rect 59760 1350 59770 1390
rect 59810 1350 59820 1390
rect 59860 1350 59870 1390
rect 59910 1350 59920 1390
rect 59960 1350 59965 1390
rect 59715 1340 59965 1350
rect 59715 1300 59720 1340
rect 59760 1300 59770 1340
rect 59810 1300 59820 1340
rect 59860 1300 59870 1340
rect 59910 1300 59920 1340
rect 59960 1300 59965 1340
rect 59715 1295 59965 1300
rect 60110 1320 60340 1405
rect 60460 1320 60690 1405
rect 60810 1320 61040 1405
rect 61160 1320 61390 1405
rect 61510 1320 61740 1405
rect 54105 1265 54355 1275
rect 54105 1225 54110 1265
rect 54150 1225 54160 1265
rect 54200 1225 54210 1265
rect 54250 1225 54260 1265
rect 54300 1225 54310 1265
rect 54350 1225 54355 1265
rect 54105 1220 54355 1225
rect 60110 1270 61740 1320
rect 60110 1175 60340 1270
rect 60460 1175 60690 1270
rect 60810 1175 61040 1270
rect 61160 1175 61390 1270
rect 61510 1175 61740 1270
rect 52850 1055 52900 1175
rect 60900 1055 60950 1175
rect 52060 970 52290 1055
rect 52410 970 52640 1055
rect 52760 970 52990 1055
rect 53110 970 53340 1055
rect 53460 970 53690 1055
rect 52060 920 53690 970
rect 52060 825 52290 920
rect 52410 825 52640 920
rect 52760 825 52990 920
rect 53110 825 53340 920
rect 53460 825 53690 920
rect 60110 970 60340 1055
rect 60460 970 60690 1055
rect 60810 970 61040 1055
rect 61160 970 61390 1055
rect 61510 970 61740 1055
rect 60110 920 61740 970
rect 60110 825 60340 920
rect 60460 825 60690 920
rect 60810 825 61040 920
rect 61160 825 61390 920
rect 61510 825 61740 920
rect 52850 705 52900 825
rect 60900 705 60950 825
rect 52060 620 52290 705
rect 52410 620 52640 705
rect 52760 620 52990 705
rect 53110 620 53340 705
rect 53460 620 53690 705
rect 52060 570 53690 620
rect 52060 475 52290 570
rect 52410 475 52640 570
rect 52760 475 52990 570
rect 53110 475 53340 570
rect 53460 475 53690 570
rect 60110 620 60340 705
rect 60460 620 60690 705
rect 60810 620 61040 705
rect 61160 620 61390 705
rect 61510 620 61740 705
rect 60110 570 61740 620
rect 60110 475 60340 570
rect 60460 475 60690 570
rect 60810 475 61040 570
rect 61160 475 61390 570
rect 61510 475 61740 570
rect 52850 355 52900 475
rect 60900 355 60950 475
rect 52060 270 52290 355
rect 52410 270 52640 355
rect 52760 270 52990 355
rect 53110 270 53340 355
rect 53460 270 53690 355
rect 52060 220 53690 270
rect 52060 125 52290 220
rect 52410 125 52640 220
rect 52760 125 52990 220
rect 53110 125 53340 220
rect 53460 125 53690 220
rect 60110 270 60340 355
rect 60460 270 60690 355
rect 60810 270 61040 355
rect 61160 270 61390 355
rect 61510 270 61740 355
rect 60110 220 61740 270
rect 60110 125 60340 220
rect 60460 125 60690 220
rect 60810 125 61040 220
rect 61160 125 61390 220
rect 61510 125 61740 220
rect 52850 5 52900 125
rect 60900 5 60950 125
rect 52060 -80 52290 5
rect 52410 -80 52640 5
rect 52760 -80 52990 5
rect 53110 -80 53340 5
rect 53460 -80 53690 5
rect 52060 -130 53690 -80
rect 52060 -225 52290 -130
rect 52410 -225 52640 -130
rect 52760 -225 52990 -130
rect 53110 -225 53340 -130
rect 53460 -225 53690 -130
rect 60110 -80 60340 5
rect 60460 -80 60690 5
rect 60810 -80 61040 5
rect 61160 -80 61390 5
rect 61510 -80 61740 5
rect 60110 -130 61740 -80
rect 60110 -225 60340 -130
rect 60460 -225 60690 -130
rect 60810 -225 61040 -130
rect 61160 -225 61390 -130
rect 61510 -225 61740 -130
rect 52850 -345 52900 -225
rect 60900 -345 60950 -225
rect 52060 -430 52290 -345
rect 52410 -430 52640 -345
rect 52760 -430 52990 -345
rect 53110 -430 53340 -345
rect 53460 -430 53690 -345
rect 52060 -480 53690 -430
rect 52060 -575 52290 -480
rect 52410 -575 52640 -480
rect 52760 -575 52990 -480
rect 53110 -575 53340 -480
rect 53460 -575 53690 -480
rect 60110 -430 60340 -345
rect 60460 -430 60690 -345
rect 60810 -430 61040 -345
rect 61160 -430 61390 -345
rect 61510 -430 61740 -345
rect 60110 -480 61740 -430
rect 60110 -575 60340 -480
rect 60460 -575 60690 -480
rect 60810 -575 61040 -480
rect 61160 -575 61390 -480
rect 61510 -575 61740 -480
rect 52850 -695 52900 -575
rect 60900 -695 60950 -575
rect 52060 -780 52290 -695
rect 52410 -780 52640 -695
rect 52760 -780 52990 -695
rect 53110 -780 53340 -695
rect 53460 -780 53690 -695
rect 53810 -780 54040 -695
rect 54160 -780 54390 -695
rect 54510 -780 54740 -695
rect 54860 -780 55090 -695
rect 55210 -780 55440 -695
rect 55560 -780 55790 -695
rect 55910 -780 56140 -695
rect 56260 -780 56490 -695
rect 56610 -780 56840 -695
rect 52060 -830 56840 -780
rect 52060 -925 52290 -830
rect 52410 -925 52640 -830
rect 52760 -925 52990 -830
rect 53110 -925 53340 -830
rect 53460 -925 53690 -830
rect 53810 -925 54040 -830
rect 54160 -925 54390 -830
rect 54510 -925 54740 -830
rect 54860 -925 55090 -830
rect 55210 -925 55440 -830
rect 55560 -925 55790 -830
rect 55910 -925 56140 -830
rect 56260 -925 56490 -830
rect 56610 -925 56840 -830
rect 56960 -780 57190 -695
rect 57310 -780 57540 -695
rect 57660 -780 57890 -695
rect 58010 -780 58240 -695
rect 58360 -780 58590 -695
rect 58710 -780 58940 -695
rect 59060 -780 59290 -695
rect 59410 -780 59640 -695
rect 59760 -780 59990 -695
rect 60110 -780 60340 -695
rect 60460 -780 60690 -695
rect 60810 -780 61040 -695
rect 61160 -780 61390 -695
rect 61510 -780 61740 -695
rect 56960 -830 61740 -780
rect 56960 -925 57190 -830
rect 57310 -925 57540 -830
rect 57660 -925 57890 -830
rect 58010 -925 58240 -830
rect 58360 -925 58590 -830
rect 58710 -925 58940 -830
rect 59060 -925 59290 -830
rect 59410 -925 59640 -830
rect 59760 -925 59990 -830
rect 60110 -925 60340 -830
rect 60460 -925 60690 -830
rect 60810 -925 61040 -830
rect 61160 -925 61390 -830
rect 61510 -925 61740 -830
rect 52850 -1045 52900 -925
rect 53200 -1045 53250 -925
rect 53550 -1045 53600 -925
rect 53900 -1045 53950 -925
rect 54250 -1045 54300 -925
rect 54600 -1045 54650 -925
rect 54950 -1045 55000 -925
rect 55300 -1045 55350 -925
rect 55650 -1045 55700 -925
rect 56000 -1045 56050 -925
rect 56350 -1045 56400 -925
rect 56700 -1045 56750 -925
rect 57050 -1045 57100 -925
rect 57400 -1045 57450 -925
rect 57750 -1045 57800 -925
rect 58100 -1045 58150 -925
rect 58450 -1045 58500 -925
rect 58800 -1045 58850 -925
rect 59150 -1045 59200 -925
rect 59500 -1045 59550 -925
rect 59850 -1045 59900 -925
rect 60200 -1045 60250 -925
rect 60550 -1045 60600 -925
rect 60900 -1045 60950 -925
rect 52060 -1130 52290 -1045
rect 52410 -1130 52640 -1045
rect 52760 -1130 52990 -1045
rect 52060 -1180 52990 -1130
rect 52060 -1275 52290 -1180
rect 52410 -1275 52640 -1180
rect 52760 -1275 52990 -1180
rect 53110 -1275 53340 -1045
rect 53460 -1275 53690 -1045
rect 53810 -1275 54040 -1045
rect 54160 -1275 54390 -1045
rect 54510 -1275 54740 -1045
rect 54860 -1275 55090 -1045
rect 55210 -1275 55440 -1045
rect 55560 -1275 55790 -1045
rect 55910 -1275 56140 -1045
rect 56260 -1275 56490 -1045
rect 56610 -1275 56840 -1045
rect 56960 -1275 57190 -1045
rect 57310 -1275 57540 -1045
rect 57660 -1275 57890 -1045
rect 58010 -1275 58240 -1045
rect 58360 -1275 58590 -1045
rect 58710 -1275 58940 -1045
rect 59060 -1275 59290 -1045
rect 59410 -1275 59640 -1045
rect 59760 -1275 59990 -1045
rect 60110 -1275 60340 -1045
rect 60460 -1275 60690 -1045
rect 60810 -1130 61040 -1045
rect 61160 -1130 61390 -1045
rect 61510 -1130 61740 -1045
rect 60810 -1180 61740 -1130
rect 60810 -1275 61040 -1180
rect 61160 -1275 61390 -1180
rect 61510 -1275 61740 -1180
<< via3 >>
rect 59720 1435 59760 1440
rect 59720 1405 59725 1435
rect 59725 1405 59755 1435
rect 59755 1405 59760 1435
rect 59720 1400 59760 1405
rect 59770 1435 59810 1440
rect 59770 1405 59775 1435
rect 59775 1405 59805 1435
rect 59805 1405 59810 1435
rect 59770 1400 59810 1405
rect 59820 1435 59860 1440
rect 59820 1405 59825 1435
rect 59825 1405 59855 1435
rect 59855 1405 59860 1435
rect 59820 1400 59860 1405
rect 59870 1435 59910 1440
rect 59870 1405 59875 1435
rect 59875 1405 59905 1435
rect 59905 1405 59910 1435
rect 59870 1400 59910 1405
rect 59920 1435 59960 1440
rect 59920 1405 59925 1435
rect 59925 1405 59955 1435
rect 59955 1405 59960 1435
rect 59920 1400 59960 1405
rect 54110 1360 54150 1365
rect 54110 1330 54115 1360
rect 54115 1330 54145 1360
rect 54145 1330 54150 1360
rect 54110 1325 54150 1330
rect 54160 1360 54200 1365
rect 54160 1330 54165 1360
rect 54165 1330 54195 1360
rect 54195 1330 54200 1360
rect 54160 1325 54200 1330
rect 54210 1360 54250 1365
rect 54210 1330 54215 1360
rect 54215 1330 54245 1360
rect 54245 1330 54250 1360
rect 54210 1325 54250 1330
rect 54260 1360 54300 1365
rect 54260 1330 54265 1360
rect 54265 1330 54295 1360
rect 54295 1330 54300 1360
rect 54260 1325 54300 1330
rect 54310 1360 54350 1365
rect 54310 1330 54315 1360
rect 54315 1330 54345 1360
rect 54345 1330 54350 1360
rect 54310 1325 54350 1330
rect 54110 1310 54150 1315
rect 54110 1280 54115 1310
rect 54115 1280 54145 1310
rect 54145 1280 54150 1310
rect 54110 1275 54150 1280
rect 54160 1310 54200 1315
rect 54160 1280 54165 1310
rect 54165 1280 54195 1310
rect 54195 1280 54200 1310
rect 54160 1275 54200 1280
rect 54210 1310 54250 1315
rect 54210 1280 54215 1310
rect 54215 1280 54245 1310
rect 54245 1280 54250 1310
rect 54210 1275 54250 1280
rect 54260 1310 54300 1315
rect 54260 1280 54265 1310
rect 54265 1280 54295 1310
rect 54295 1280 54300 1310
rect 54260 1275 54300 1280
rect 54310 1310 54350 1315
rect 54310 1280 54315 1310
rect 54315 1280 54345 1310
rect 54345 1280 54350 1310
rect 54310 1275 54350 1280
rect 59720 1385 59760 1390
rect 59720 1355 59725 1385
rect 59725 1355 59755 1385
rect 59755 1355 59760 1385
rect 59720 1350 59760 1355
rect 59770 1385 59810 1390
rect 59770 1355 59775 1385
rect 59775 1355 59805 1385
rect 59805 1355 59810 1385
rect 59770 1350 59810 1355
rect 59820 1385 59860 1390
rect 59820 1355 59825 1385
rect 59825 1355 59855 1385
rect 59855 1355 59860 1385
rect 59820 1350 59860 1355
rect 59870 1385 59910 1390
rect 59870 1355 59875 1385
rect 59875 1355 59905 1385
rect 59905 1355 59910 1385
rect 59870 1350 59910 1355
rect 59920 1385 59960 1390
rect 59920 1355 59925 1385
rect 59925 1355 59955 1385
rect 59955 1355 59960 1385
rect 59920 1350 59960 1355
rect 59720 1335 59760 1340
rect 59720 1305 59725 1335
rect 59725 1305 59755 1335
rect 59755 1305 59760 1335
rect 59720 1300 59760 1305
rect 59770 1335 59810 1340
rect 59770 1305 59775 1335
rect 59775 1305 59805 1335
rect 59805 1305 59810 1335
rect 59770 1300 59810 1305
rect 59820 1335 59860 1340
rect 59820 1305 59825 1335
rect 59825 1305 59855 1335
rect 59855 1305 59860 1335
rect 59820 1300 59860 1305
rect 59870 1335 59910 1340
rect 59870 1305 59875 1335
rect 59875 1305 59905 1335
rect 59905 1305 59910 1335
rect 59870 1300 59910 1305
rect 59920 1335 59960 1340
rect 59920 1305 59925 1335
rect 59925 1305 59955 1335
rect 59955 1305 59960 1335
rect 59920 1300 59960 1305
rect 54110 1260 54150 1265
rect 54110 1230 54115 1260
rect 54115 1230 54145 1260
rect 54145 1230 54150 1260
rect 54110 1225 54150 1230
rect 54160 1260 54200 1265
rect 54160 1230 54165 1260
rect 54165 1230 54195 1260
rect 54195 1230 54200 1260
rect 54160 1225 54200 1230
rect 54210 1260 54250 1265
rect 54210 1230 54215 1260
rect 54215 1230 54245 1260
rect 54245 1230 54250 1260
rect 54210 1225 54250 1230
rect 54260 1260 54300 1265
rect 54260 1230 54265 1260
rect 54265 1230 54295 1260
rect 54295 1230 54300 1260
rect 54260 1225 54300 1230
rect 54310 1260 54350 1265
rect 54310 1230 54315 1260
rect 54315 1230 54345 1260
rect 54345 1230 54350 1260
rect 54310 1225 54350 1230
<< mimcap >>
rect 52075 6215 52275 6290
rect 52075 6175 52155 6215
rect 52195 6175 52275 6215
rect 52075 6090 52275 6175
rect 52425 6215 52625 6290
rect 52425 6175 52505 6215
rect 52545 6175 52625 6215
rect 52425 6090 52625 6175
rect 52775 6215 52975 6290
rect 52775 6175 52855 6215
rect 52895 6175 52975 6215
rect 52775 6090 52975 6175
rect 53125 6215 53325 6290
rect 53125 6175 53205 6215
rect 53245 6175 53325 6215
rect 53125 6090 53325 6175
rect 53475 6215 53675 6290
rect 53475 6175 53555 6215
rect 53595 6175 53675 6215
rect 53475 6090 53675 6175
rect 53825 6215 54025 6290
rect 53825 6175 53905 6215
rect 53945 6175 54025 6215
rect 53825 6090 54025 6175
rect 54175 6215 54375 6290
rect 54175 6175 54255 6215
rect 54295 6175 54375 6215
rect 54175 6090 54375 6175
rect 54525 6215 54725 6290
rect 54525 6175 54605 6215
rect 54645 6175 54725 6215
rect 54525 6090 54725 6175
rect 54875 6215 55075 6290
rect 54875 6175 54955 6215
rect 54995 6175 55075 6215
rect 54875 6090 55075 6175
rect 55225 6215 55425 6290
rect 55225 6175 55305 6215
rect 55345 6175 55425 6215
rect 55225 6090 55425 6175
rect 55575 6215 55775 6290
rect 55575 6175 55655 6215
rect 55695 6175 55775 6215
rect 55575 6090 55775 6175
rect 55925 6215 56125 6290
rect 55925 6175 56005 6215
rect 56045 6175 56125 6215
rect 55925 6090 56125 6175
rect 56275 6215 56475 6290
rect 56275 6175 56355 6215
rect 56395 6175 56475 6215
rect 56275 6090 56475 6175
rect 56625 6215 56825 6290
rect 56625 6175 56705 6215
rect 56745 6175 56825 6215
rect 56625 6090 56825 6175
rect 56975 6215 57175 6290
rect 56975 6175 57055 6215
rect 57095 6175 57175 6215
rect 56975 6090 57175 6175
rect 57325 6215 57525 6290
rect 57325 6175 57405 6215
rect 57445 6175 57525 6215
rect 57325 6090 57525 6175
rect 57675 6215 57875 6290
rect 57675 6175 57755 6215
rect 57795 6175 57875 6215
rect 57675 6090 57875 6175
rect 58025 6215 58225 6290
rect 58025 6175 58105 6215
rect 58145 6175 58225 6215
rect 58025 6090 58225 6175
rect 58375 6215 58575 6290
rect 58375 6175 58455 6215
rect 58495 6175 58575 6215
rect 58375 6090 58575 6175
rect 58725 6215 58925 6290
rect 58725 6175 58805 6215
rect 58845 6175 58925 6215
rect 58725 6090 58925 6175
rect 59075 6215 59275 6290
rect 59075 6175 59155 6215
rect 59195 6175 59275 6215
rect 59075 6090 59275 6175
rect 59425 6215 59625 6290
rect 59425 6175 59505 6215
rect 59545 6175 59625 6215
rect 59425 6090 59625 6175
rect 59775 6215 59975 6290
rect 59775 6175 59855 6215
rect 59895 6175 59975 6215
rect 59775 6090 59975 6175
rect 60125 6215 60325 6290
rect 60125 6175 60205 6215
rect 60245 6175 60325 6215
rect 60125 6090 60325 6175
rect 60475 6215 60675 6290
rect 60475 6175 60555 6215
rect 60595 6175 60675 6215
rect 60475 6090 60675 6175
rect 60825 6215 61025 6290
rect 60825 6175 60905 6215
rect 60945 6175 61025 6215
rect 60825 6090 61025 6175
rect 61175 6215 61375 6290
rect 61175 6175 61255 6215
rect 61295 6175 61375 6215
rect 61175 6090 61375 6175
rect 61525 6215 61725 6290
rect 61525 6175 61605 6215
rect 61645 6175 61725 6215
rect 61525 6090 61725 6175
rect 52075 5865 52275 5940
rect 52075 5825 52155 5865
rect 52195 5825 52275 5865
rect 52075 5740 52275 5825
rect 52425 5865 52625 5940
rect 52425 5825 52505 5865
rect 52545 5825 52625 5865
rect 52425 5740 52625 5825
rect 52775 5865 52975 5940
rect 52775 5825 52855 5865
rect 52895 5825 52975 5865
rect 52775 5740 52975 5825
rect 53125 5865 53325 5940
rect 53125 5825 53205 5865
rect 53245 5825 53325 5865
rect 53125 5740 53325 5825
rect 53475 5865 53675 5940
rect 53475 5825 53555 5865
rect 53595 5825 53675 5865
rect 53475 5740 53675 5825
rect 53825 5865 54025 5940
rect 53825 5825 53905 5865
rect 53945 5825 54025 5865
rect 53825 5740 54025 5825
rect 54175 5865 54375 5940
rect 54175 5825 54255 5865
rect 54295 5825 54375 5865
rect 54175 5740 54375 5825
rect 54525 5865 54725 5940
rect 54525 5825 54605 5865
rect 54645 5825 54725 5865
rect 54525 5740 54725 5825
rect 54875 5865 55075 5940
rect 54875 5825 54955 5865
rect 54995 5825 55075 5865
rect 54875 5740 55075 5825
rect 55225 5865 55425 5940
rect 55225 5825 55305 5865
rect 55345 5825 55425 5865
rect 55225 5740 55425 5825
rect 55575 5865 55775 5940
rect 55575 5825 55655 5865
rect 55695 5825 55775 5865
rect 55575 5740 55775 5825
rect 55925 5865 56125 5940
rect 55925 5825 56005 5865
rect 56045 5825 56125 5865
rect 55925 5740 56125 5825
rect 56275 5865 56475 5940
rect 56275 5825 56355 5865
rect 56395 5825 56475 5865
rect 56275 5740 56475 5825
rect 56625 5865 56825 5940
rect 56625 5825 56705 5865
rect 56745 5825 56825 5865
rect 56625 5740 56825 5825
rect 56975 5865 57175 5940
rect 56975 5825 57055 5865
rect 57095 5825 57175 5865
rect 56975 5740 57175 5825
rect 57325 5865 57525 5940
rect 57325 5825 57405 5865
rect 57445 5825 57525 5865
rect 57325 5740 57525 5825
rect 57675 5865 57875 5940
rect 57675 5825 57755 5865
rect 57795 5825 57875 5865
rect 57675 5740 57875 5825
rect 58025 5865 58225 5940
rect 58025 5825 58105 5865
rect 58145 5825 58225 5865
rect 58025 5740 58225 5825
rect 58375 5865 58575 5940
rect 58375 5825 58455 5865
rect 58495 5825 58575 5865
rect 58375 5740 58575 5825
rect 58725 5865 58925 5940
rect 58725 5825 58805 5865
rect 58845 5825 58925 5865
rect 58725 5740 58925 5825
rect 59075 5865 59275 5940
rect 59075 5825 59155 5865
rect 59195 5825 59275 5865
rect 59075 5740 59275 5825
rect 59425 5865 59625 5940
rect 59425 5825 59505 5865
rect 59545 5825 59625 5865
rect 59425 5740 59625 5825
rect 59775 5865 59975 5940
rect 59775 5825 59855 5865
rect 59895 5825 59975 5865
rect 59775 5740 59975 5825
rect 60125 5865 60325 5940
rect 60125 5825 60205 5865
rect 60245 5825 60325 5865
rect 60125 5740 60325 5825
rect 60475 5865 60675 5940
rect 60475 5825 60555 5865
rect 60595 5825 60675 5865
rect 60475 5740 60675 5825
rect 60825 5865 61025 5940
rect 60825 5825 60905 5865
rect 60945 5825 61025 5865
rect 60825 5740 61025 5825
rect 61175 5865 61375 5940
rect 61175 5825 61255 5865
rect 61295 5825 61375 5865
rect 61175 5740 61375 5825
rect 61525 5865 61725 5940
rect 61525 5825 61605 5865
rect 61645 5825 61725 5865
rect 61525 5740 61725 5825
rect 52075 5515 52275 5590
rect 52075 5475 52155 5515
rect 52195 5475 52275 5515
rect 52075 5390 52275 5475
rect 52425 5515 52625 5590
rect 52425 5475 52505 5515
rect 52545 5475 52625 5515
rect 52425 5390 52625 5475
rect 52775 5515 52975 5590
rect 52775 5475 52855 5515
rect 52895 5475 52975 5515
rect 52775 5390 52975 5475
rect 53125 5515 53325 5590
rect 53125 5475 53205 5515
rect 53245 5475 53325 5515
rect 53125 5390 53325 5475
rect 53475 5515 53675 5590
rect 53475 5475 53555 5515
rect 53595 5475 53675 5515
rect 53475 5390 53675 5475
rect 53825 5515 54025 5590
rect 53825 5475 53905 5515
rect 53945 5475 54025 5515
rect 53825 5390 54025 5475
rect 54175 5515 54375 5590
rect 54175 5475 54255 5515
rect 54295 5475 54375 5515
rect 54175 5390 54375 5475
rect 54525 5515 54725 5590
rect 54525 5475 54605 5515
rect 54645 5475 54725 5515
rect 54525 5390 54725 5475
rect 54875 5515 55075 5590
rect 54875 5475 54955 5515
rect 54995 5475 55075 5515
rect 54875 5390 55075 5475
rect 55225 5505 55425 5590
rect 55225 5465 55305 5505
rect 55345 5465 55425 5505
rect 55225 5390 55425 5465
rect 55575 5505 55775 5590
rect 55575 5465 55655 5505
rect 55695 5465 55775 5505
rect 55575 5390 55775 5465
rect 55925 5505 56125 5590
rect 55925 5465 56005 5505
rect 56045 5465 56125 5505
rect 55925 5390 56125 5465
rect 56275 5505 56475 5590
rect 56275 5465 56355 5505
rect 56395 5465 56475 5505
rect 56275 5390 56475 5465
rect 56625 5505 56825 5590
rect 56625 5465 56705 5505
rect 56745 5465 56825 5505
rect 56625 5390 56825 5465
rect 56975 5505 57175 5590
rect 56975 5465 57055 5505
rect 57095 5465 57175 5505
rect 56975 5390 57175 5465
rect 57325 5505 57525 5590
rect 57325 5465 57405 5505
rect 57445 5465 57525 5505
rect 57325 5390 57525 5465
rect 57675 5505 57875 5590
rect 57675 5465 57755 5505
rect 57795 5465 57875 5505
rect 57675 5390 57875 5465
rect 58025 5505 58225 5590
rect 58025 5465 58105 5505
rect 58145 5465 58225 5505
rect 58025 5390 58225 5465
rect 58375 5505 58575 5590
rect 58375 5465 58455 5505
rect 58495 5465 58575 5505
rect 58375 5390 58575 5465
rect 58725 5515 58925 5590
rect 58725 5475 58805 5515
rect 58845 5475 58925 5515
rect 58725 5390 58925 5475
rect 59075 5515 59275 5590
rect 59075 5475 59155 5515
rect 59195 5475 59275 5515
rect 59075 5390 59275 5475
rect 59425 5515 59625 5590
rect 59425 5475 59505 5515
rect 59545 5475 59625 5515
rect 59425 5390 59625 5475
rect 59775 5515 59975 5590
rect 59775 5475 59855 5515
rect 59895 5475 59975 5515
rect 59775 5390 59975 5475
rect 60125 5515 60325 5590
rect 60125 5475 60205 5515
rect 60245 5475 60325 5515
rect 60125 5390 60325 5475
rect 60475 5515 60675 5590
rect 60475 5475 60555 5515
rect 60595 5475 60675 5515
rect 60475 5390 60675 5475
rect 60825 5515 61025 5590
rect 60825 5475 60905 5515
rect 60945 5475 61025 5515
rect 60825 5390 61025 5475
rect 61175 5515 61375 5590
rect 61175 5475 61255 5515
rect 61295 5475 61375 5515
rect 61175 5390 61375 5475
rect 61525 5515 61725 5590
rect 61525 5475 61605 5515
rect 61645 5475 61725 5515
rect 61525 5390 61725 5475
rect 52075 5165 52275 5240
rect 52075 5125 52155 5165
rect 52195 5125 52275 5165
rect 52075 5040 52275 5125
rect 52425 5165 52625 5240
rect 52425 5125 52505 5165
rect 52545 5125 52625 5165
rect 52425 5040 52625 5125
rect 52775 5165 52975 5240
rect 52775 5125 52855 5165
rect 52895 5125 52975 5165
rect 52775 5040 52975 5125
rect 53125 5165 53325 5240
rect 53125 5125 53205 5165
rect 53245 5125 53325 5165
rect 53125 5040 53325 5125
rect 53475 5165 53675 5240
rect 53475 5125 53555 5165
rect 53595 5125 53675 5165
rect 53475 5040 53675 5125
rect 53825 5165 54025 5240
rect 53825 5125 53905 5165
rect 53945 5125 54025 5165
rect 53825 5040 54025 5125
rect 54175 5165 54375 5240
rect 54175 5125 54255 5165
rect 54295 5125 54375 5165
rect 54175 5040 54375 5125
rect 54525 5165 54725 5240
rect 54525 5125 54605 5165
rect 54645 5125 54725 5165
rect 54525 5040 54725 5125
rect 59075 5165 59275 5240
rect 59075 5125 59155 5165
rect 59195 5125 59275 5165
rect 59075 5040 59275 5125
rect 59425 5165 59625 5240
rect 59425 5125 59505 5165
rect 59545 5125 59625 5165
rect 59425 5040 59625 5125
rect 59775 5165 59975 5240
rect 59775 5125 59855 5165
rect 59895 5125 59975 5165
rect 59775 5040 59975 5125
rect 60125 5165 60325 5240
rect 60125 5125 60205 5165
rect 60245 5125 60325 5165
rect 60125 5040 60325 5125
rect 60475 5165 60675 5240
rect 60475 5125 60555 5165
rect 60595 5125 60675 5165
rect 60475 5040 60675 5125
rect 60825 5165 61025 5240
rect 60825 5125 60905 5165
rect 60945 5125 61025 5165
rect 60825 5040 61025 5125
rect 61175 5165 61375 5240
rect 61175 5125 61255 5165
rect 61295 5125 61375 5165
rect 61175 5040 61375 5125
rect 61525 5165 61725 5240
rect 61525 5125 61605 5165
rect 61645 5125 61725 5165
rect 61525 5040 61725 5125
rect 52075 4815 52275 4890
rect 52075 4775 52155 4815
rect 52195 4775 52275 4815
rect 52075 4690 52275 4775
rect 52425 4815 52625 4890
rect 52425 4775 52505 4815
rect 52545 4775 52625 4815
rect 52425 4690 52625 4775
rect 52775 4815 52975 4890
rect 52775 4775 52855 4815
rect 52895 4775 52975 4815
rect 52775 4690 52975 4775
rect 53125 4815 53325 4890
rect 53125 4775 53205 4815
rect 53245 4775 53325 4815
rect 53125 4690 53325 4775
rect 53475 4815 53675 4890
rect 53475 4775 53555 4815
rect 53595 4775 53675 4815
rect 53475 4690 53675 4775
rect 60125 4815 60325 4890
rect 60125 4775 60205 4815
rect 60245 4775 60325 4815
rect 60125 4690 60325 4775
rect 60475 4815 60675 4890
rect 60475 4775 60555 4815
rect 60595 4775 60675 4815
rect 60475 4690 60675 4775
rect 60825 4815 61025 4890
rect 60825 4775 60905 4815
rect 60945 4775 61025 4815
rect 60825 4690 61025 4775
rect 61175 4815 61375 4890
rect 61175 4775 61255 4815
rect 61295 4775 61375 4815
rect 61175 4690 61375 4775
rect 61525 4815 61725 4890
rect 61525 4775 61605 4815
rect 61645 4775 61725 4815
rect 61525 4690 61725 4775
rect 52075 4465 52275 4540
rect 52075 4425 52155 4465
rect 52195 4425 52275 4465
rect 52075 4340 52275 4425
rect 52425 4465 52625 4540
rect 52425 4425 52505 4465
rect 52545 4425 52625 4465
rect 52425 4340 52625 4425
rect 52775 4465 52975 4540
rect 52775 4425 52855 4465
rect 52895 4425 52975 4465
rect 52775 4340 52975 4425
rect 53125 4465 53325 4540
rect 53125 4425 53205 4465
rect 53245 4425 53325 4465
rect 53125 4340 53325 4425
rect 53475 4465 53675 4540
rect 53475 4425 53555 4465
rect 53595 4425 53675 4465
rect 53475 4340 53675 4425
rect 60125 4465 60325 4540
rect 60125 4425 60205 4465
rect 60245 4425 60325 4465
rect 60125 4340 60325 4425
rect 60475 4465 60675 4540
rect 60475 4425 60555 4465
rect 60595 4425 60675 4465
rect 60475 4340 60675 4425
rect 60825 4465 61025 4540
rect 60825 4425 60905 4465
rect 60945 4425 61025 4465
rect 60825 4340 61025 4425
rect 61175 4465 61375 4540
rect 61175 4425 61255 4465
rect 61295 4425 61375 4465
rect 61175 4340 61375 4425
rect 61525 4465 61725 4540
rect 61525 4425 61605 4465
rect 61645 4425 61725 4465
rect 61525 4340 61725 4425
rect 52075 4115 52275 4190
rect 52075 4075 52155 4115
rect 52195 4075 52275 4115
rect 52075 3990 52275 4075
rect 52425 4115 52625 4190
rect 52425 4075 52505 4115
rect 52545 4075 52625 4115
rect 52425 3990 52625 4075
rect 52775 4115 52975 4190
rect 52775 4075 52855 4115
rect 52895 4075 52975 4115
rect 52775 3990 52975 4075
rect 53125 4115 53325 4190
rect 53125 4075 53205 4115
rect 53245 4075 53325 4115
rect 53125 3990 53325 4075
rect 53475 4115 53675 4190
rect 53475 4075 53555 4115
rect 53595 4075 53675 4115
rect 53475 3990 53675 4075
rect 60125 4115 60325 4190
rect 60125 4075 60205 4115
rect 60245 4075 60325 4115
rect 60125 3990 60325 4075
rect 60475 4115 60675 4190
rect 60475 4075 60555 4115
rect 60595 4075 60675 4115
rect 60475 3990 60675 4075
rect 60825 4115 61025 4190
rect 60825 4075 60905 4115
rect 60945 4075 61025 4115
rect 60825 3990 61025 4075
rect 61175 4115 61375 4190
rect 61175 4075 61255 4115
rect 61295 4075 61375 4115
rect 61175 3990 61375 4075
rect 61525 4115 61725 4190
rect 61525 4075 61605 4115
rect 61645 4075 61725 4115
rect 61525 3990 61725 4075
rect 52075 3765 52275 3840
rect 52075 3725 52155 3765
rect 52195 3725 52275 3765
rect 52075 3640 52275 3725
rect 52425 3765 52625 3840
rect 52425 3725 52505 3765
rect 52545 3725 52625 3765
rect 52425 3640 52625 3725
rect 52775 3765 52975 3840
rect 52775 3725 52855 3765
rect 52895 3725 52975 3765
rect 52775 3640 52975 3725
rect 53125 3765 53325 3840
rect 53125 3725 53205 3765
rect 53245 3725 53325 3765
rect 53125 3640 53325 3725
rect 53475 3765 53675 3840
rect 53475 3725 53555 3765
rect 53595 3725 53675 3765
rect 53475 3640 53675 3725
rect 60125 3765 60325 3840
rect 60125 3725 60205 3765
rect 60245 3725 60325 3765
rect 60125 3640 60325 3725
rect 60475 3765 60675 3840
rect 60475 3725 60555 3765
rect 60595 3725 60675 3765
rect 60475 3640 60675 3725
rect 60825 3765 61025 3840
rect 60825 3725 60905 3765
rect 60945 3725 61025 3765
rect 60825 3640 61025 3725
rect 61175 3765 61375 3840
rect 61175 3725 61255 3765
rect 61295 3725 61375 3765
rect 61175 3640 61375 3725
rect 61525 3765 61725 3840
rect 61525 3725 61605 3765
rect 61645 3725 61725 3765
rect 61525 3640 61725 3725
rect 52075 3415 52275 3490
rect 52075 3375 52155 3415
rect 52195 3375 52275 3415
rect 52075 3290 52275 3375
rect 52425 3415 52625 3490
rect 52425 3375 52505 3415
rect 52545 3375 52625 3415
rect 52425 3290 52625 3375
rect 52775 3415 52975 3490
rect 52775 3375 52855 3415
rect 52895 3375 52975 3415
rect 52775 3290 52975 3375
rect 53125 3415 53325 3490
rect 53125 3375 53205 3415
rect 53245 3375 53325 3415
rect 53125 3290 53325 3375
rect 53475 3415 53675 3490
rect 53475 3375 53555 3415
rect 53595 3375 53675 3415
rect 53475 3290 53675 3375
rect 60125 3415 60325 3490
rect 60125 3375 60205 3415
rect 60245 3375 60325 3415
rect 60125 3290 60325 3375
rect 60475 3415 60675 3490
rect 60475 3375 60555 3415
rect 60595 3375 60675 3415
rect 60475 3290 60675 3375
rect 60825 3415 61025 3490
rect 60825 3375 60905 3415
rect 60945 3375 61025 3415
rect 60825 3290 61025 3375
rect 61175 3415 61375 3490
rect 61175 3375 61255 3415
rect 61295 3375 61375 3415
rect 61175 3290 61375 3375
rect 61525 3415 61725 3490
rect 61525 3375 61605 3415
rect 61645 3375 61725 3415
rect 61525 3290 61725 3375
rect 52075 3065 52275 3140
rect 52075 3025 52155 3065
rect 52195 3025 52275 3065
rect 52075 2940 52275 3025
rect 52425 3065 52625 3140
rect 52425 3025 52505 3065
rect 52545 3025 52625 3065
rect 52425 2940 52625 3025
rect 52775 3065 52975 3140
rect 52775 3025 52855 3065
rect 52895 3025 52975 3065
rect 52775 2940 52975 3025
rect 53125 3065 53325 3140
rect 53125 3025 53205 3065
rect 53245 3025 53325 3065
rect 53125 2940 53325 3025
rect 53475 3065 53675 3140
rect 53475 3025 53555 3065
rect 53595 3025 53675 3065
rect 53475 2940 53675 3025
rect 60125 3065 60325 3140
rect 60125 3025 60205 3065
rect 60245 3025 60325 3065
rect 60125 2940 60325 3025
rect 60475 3065 60675 3140
rect 60475 3025 60555 3065
rect 60595 3025 60675 3065
rect 60475 2940 60675 3025
rect 60825 3065 61025 3140
rect 60825 3025 60905 3065
rect 60945 3025 61025 3065
rect 60825 2940 61025 3025
rect 61175 3065 61375 3140
rect 61175 3025 61255 3065
rect 61295 3025 61375 3065
rect 61175 2940 61375 3025
rect 61525 3065 61725 3140
rect 61525 3025 61605 3065
rect 61645 3025 61725 3065
rect 61525 2940 61725 3025
rect 52075 2715 52275 2790
rect 52075 2675 52155 2715
rect 52195 2675 52275 2715
rect 52075 2590 52275 2675
rect 52425 2715 52625 2790
rect 52425 2675 52505 2715
rect 52545 2675 52625 2715
rect 52425 2590 52625 2675
rect 52775 2715 52975 2790
rect 52775 2675 52855 2715
rect 52895 2675 52975 2715
rect 52775 2590 52975 2675
rect 53125 2715 53325 2790
rect 53125 2675 53205 2715
rect 53245 2675 53325 2715
rect 53125 2590 53325 2675
rect 53475 2715 53675 2790
rect 53475 2675 53555 2715
rect 53595 2675 53675 2715
rect 53475 2590 53675 2675
rect 60125 2715 60325 2790
rect 60125 2675 60205 2715
rect 60245 2675 60325 2715
rect 60125 2590 60325 2675
rect 60475 2715 60675 2790
rect 60475 2675 60555 2715
rect 60595 2675 60675 2715
rect 60475 2590 60675 2675
rect 60825 2715 61025 2790
rect 60825 2675 60905 2715
rect 60945 2675 61025 2715
rect 60825 2590 61025 2675
rect 61175 2715 61375 2790
rect 61175 2675 61255 2715
rect 61295 2675 61375 2715
rect 61175 2590 61375 2675
rect 61525 2715 61725 2790
rect 61525 2675 61605 2715
rect 61645 2675 61725 2715
rect 61525 2590 61725 2675
rect 52075 2365 52275 2440
rect 52075 2325 52155 2365
rect 52195 2325 52275 2365
rect 52075 2240 52275 2325
rect 52425 2365 52625 2440
rect 52425 2325 52505 2365
rect 52545 2325 52625 2365
rect 52425 2240 52625 2325
rect 52775 2365 52975 2440
rect 52775 2325 52855 2365
rect 52895 2325 52975 2365
rect 52775 2240 52975 2325
rect 53125 2365 53325 2440
rect 53125 2325 53205 2365
rect 53245 2325 53325 2365
rect 53125 2240 53325 2325
rect 53475 2365 53675 2440
rect 53475 2325 53555 2365
rect 53595 2325 53675 2365
rect 53475 2240 53675 2325
rect 60125 2365 60325 2440
rect 60125 2325 60205 2365
rect 60245 2325 60325 2365
rect 60125 2240 60325 2325
rect 60475 2365 60675 2440
rect 60475 2325 60555 2365
rect 60595 2325 60675 2365
rect 60475 2240 60675 2325
rect 60825 2365 61025 2440
rect 60825 2325 60905 2365
rect 60945 2325 61025 2365
rect 60825 2240 61025 2325
rect 61175 2365 61375 2440
rect 61175 2325 61255 2365
rect 61295 2325 61375 2365
rect 61175 2240 61375 2325
rect 61525 2365 61725 2440
rect 61525 2325 61605 2365
rect 61645 2325 61725 2365
rect 61525 2240 61725 2325
rect 52075 2015 52275 2090
rect 52075 1975 52155 2015
rect 52195 1975 52275 2015
rect 52075 1890 52275 1975
rect 52425 2015 52625 2090
rect 52425 1975 52505 2015
rect 52545 1975 52625 2015
rect 52425 1890 52625 1975
rect 52775 2015 52975 2090
rect 52775 1975 52855 2015
rect 52895 1975 52975 2015
rect 52775 1890 52975 1975
rect 53125 2015 53325 2090
rect 53125 1975 53205 2015
rect 53245 1975 53325 2015
rect 53125 1890 53325 1975
rect 53475 2015 53675 2090
rect 53475 1975 53555 2015
rect 53595 1975 53675 2015
rect 53475 1890 53675 1975
rect 60125 2015 60325 2090
rect 60125 1975 60205 2015
rect 60245 1975 60325 2015
rect 60125 1890 60325 1975
rect 60475 2015 60675 2090
rect 60475 1975 60555 2015
rect 60595 1975 60675 2015
rect 60475 1890 60675 1975
rect 60825 2015 61025 2090
rect 60825 1975 60905 2015
rect 60945 1975 61025 2015
rect 60825 1890 61025 1975
rect 61175 2015 61375 2090
rect 61175 1975 61255 2015
rect 61295 1975 61375 2015
rect 61175 1890 61375 1975
rect 61525 2015 61725 2090
rect 61525 1975 61605 2015
rect 61645 1975 61725 2015
rect 61525 1890 61725 1975
rect 52075 1665 52275 1740
rect 52075 1625 52155 1665
rect 52195 1625 52275 1665
rect 52075 1540 52275 1625
rect 52425 1665 52625 1740
rect 52425 1625 52505 1665
rect 52545 1625 52625 1665
rect 52425 1540 52625 1625
rect 52775 1665 52975 1740
rect 52775 1625 52855 1665
rect 52895 1625 52975 1665
rect 52775 1540 52975 1625
rect 53125 1665 53325 1740
rect 53125 1625 53205 1665
rect 53245 1625 53325 1665
rect 53125 1540 53325 1625
rect 53475 1665 53675 1740
rect 53475 1625 53555 1665
rect 53595 1625 53675 1665
rect 53475 1540 53675 1625
rect 60125 1665 60325 1740
rect 60125 1625 60205 1665
rect 60245 1625 60325 1665
rect 60125 1540 60325 1625
rect 60475 1665 60675 1740
rect 60475 1625 60555 1665
rect 60595 1625 60675 1665
rect 60475 1540 60675 1625
rect 60825 1665 61025 1740
rect 60825 1625 60905 1665
rect 60945 1625 61025 1665
rect 60825 1540 61025 1625
rect 61175 1665 61375 1740
rect 61175 1625 61255 1665
rect 61295 1625 61375 1665
rect 61175 1540 61375 1625
rect 61525 1665 61725 1740
rect 61525 1625 61605 1665
rect 61645 1625 61725 1665
rect 61525 1540 61725 1625
rect 52075 1315 52275 1390
rect 52075 1275 52155 1315
rect 52195 1275 52275 1315
rect 52075 1190 52275 1275
rect 52425 1315 52625 1390
rect 52425 1275 52505 1315
rect 52545 1275 52625 1315
rect 52425 1190 52625 1275
rect 52775 1315 52975 1390
rect 52775 1275 52855 1315
rect 52895 1275 52975 1315
rect 52775 1190 52975 1275
rect 53125 1315 53325 1390
rect 53125 1275 53205 1315
rect 53245 1275 53325 1315
rect 53125 1190 53325 1275
rect 53475 1315 53675 1390
rect 53475 1275 53555 1315
rect 53595 1275 53675 1315
rect 53475 1190 53675 1275
rect 60125 1315 60325 1390
rect 60125 1275 60205 1315
rect 60245 1275 60325 1315
rect 60125 1190 60325 1275
rect 60475 1315 60675 1390
rect 60475 1275 60555 1315
rect 60595 1275 60675 1315
rect 60475 1190 60675 1275
rect 60825 1315 61025 1390
rect 60825 1275 60905 1315
rect 60945 1275 61025 1315
rect 60825 1190 61025 1275
rect 61175 1315 61375 1390
rect 61175 1275 61255 1315
rect 61295 1275 61375 1315
rect 61175 1190 61375 1275
rect 61525 1315 61725 1390
rect 61525 1275 61605 1315
rect 61645 1275 61725 1315
rect 61525 1190 61725 1275
rect 52075 965 52275 1040
rect 52075 925 52155 965
rect 52195 925 52275 965
rect 52075 840 52275 925
rect 52425 965 52625 1040
rect 52425 925 52505 965
rect 52545 925 52625 965
rect 52425 840 52625 925
rect 52775 965 52975 1040
rect 52775 925 52855 965
rect 52895 925 52975 965
rect 52775 840 52975 925
rect 53125 965 53325 1040
rect 53125 925 53205 965
rect 53245 925 53325 965
rect 53125 840 53325 925
rect 53475 965 53675 1040
rect 53475 925 53555 965
rect 53595 925 53675 965
rect 53475 840 53675 925
rect 60125 965 60325 1040
rect 60125 925 60205 965
rect 60245 925 60325 965
rect 60125 840 60325 925
rect 60475 965 60675 1040
rect 60475 925 60555 965
rect 60595 925 60675 965
rect 60475 840 60675 925
rect 60825 965 61025 1040
rect 60825 925 60905 965
rect 60945 925 61025 965
rect 60825 840 61025 925
rect 61175 965 61375 1040
rect 61175 925 61255 965
rect 61295 925 61375 965
rect 61175 840 61375 925
rect 61525 965 61725 1040
rect 61525 925 61605 965
rect 61645 925 61725 965
rect 61525 840 61725 925
rect 52075 615 52275 690
rect 52075 575 52155 615
rect 52195 575 52275 615
rect 52075 490 52275 575
rect 52425 615 52625 690
rect 52425 575 52505 615
rect 52545 575 52625 615
rect 52425 490 52625 575
rect 52775 615 52975 690
rect 52775 575 52855 615
rect 52895 575 52975 615
rect 52775 490 52975 575
rect 53125 615 53325 690
rect 53125 575 53205 615
rect 53245 575 53325 615
rect 53125 490 53325 575
rect 53475 615 53675 690
rect 53475 575 53555 615
rect 53595 575 53675 615
rect 53475 490 53675 575
rect 60125 615 60325 690
rect 60125 575 60205 615
rect 60245 575 60325 615
rect 60125 490 60325 575
rect 60475 615 60675 690
rect 60475 575 60555 615
rect 60595 575 60675 615
rect 60475 490 60675 575
rect 60825 615 61025 690
rect 60825 575 60905 615
rect 60945 575 61025 615
rect 60825 490 61025 575
rect 61175 615 61375 690
rect 61175 575 61255 615
rect 61295 575 61375 615
rect 61175 490 61375 575
rect 61525 615 61725 690
rect 61525 575 61605 615
rect 61645 575 61725 615
rect 61525 490 61725 575
rect 52075 265 52275 340
rect 52075 225 52155 265
rect 52195 225 52275 265
rect 52075 140 52275 225
rect 52425 265 52625 340
rect 52425 225 52505 265
rect 52545 225 52625 265
rect 52425 140 52625 225
rect 52775 265 52975 340
rect 52775 225 52855 265
rect 52895 225 52975 265
rect 52775 140 52975 225
rect 53125 265 53325 340
rect 53125 225 53205 265
rect 53245 225 53325 265
rect 53125 140 53325 225
rect 53475 265 53675 340
rect 53475 225 53555 265
rect 53595 225 53675 265
rect 53475 140 53675 225
rect 60125 265 60325 340
rect 60125 225 60205 265
rect 60245 225 60325 265
rect 60125 140 60325 225
rect 60475 265 60675 340
rect 60475 225 60555 265
rect 60595 225 60675 265
rect 60475 140 60675 225
rect 60825 265 61025 340
rect 60825 225 60905 265
rect 60945 225 61025 265
rect 60825 140 61025 225
rect 61175 265 61375 340
rect 61175 225 61255 265
rect 61295 225 61375 265
rect 61175 140 61375 225
rect 61525 265 61725 340
rect 61525 225 61605 265
rect 61645 225 61725 265
rect 61525 140 61725 225
rect 52075 -85 52275 -10
rect 52075 -125 52155 -85
rect 52195 -125 52275 -85
rect 52075 -210 52275 -125
rect 52425 -85 52625 -10
rect 52425 -125 52505 -85
rect 52545 -125 52625 -85
rect 52425 -210 52625 -125
rect 52775 -85 52975 -10
rect 52775 -125 52855 -85
rect 52895 -125 52975 -85
rect 52775 -210 52975 -125
rect 53125 -85 53325 -10
rect 53125 -125 53205 -85
rect 53245 -125 53325 -85
rect 53125 -210 53325 -125
rect 53475 -85 53675 -10
rect 53475 -125 53555 -85
rect 53595 -125 53675 -85
rect 53475 -210 53675 -125
rect 60125 -85 60325 -10
rect 60125 -125 60205 -85
rect 60245 -125 60325 -85
rect 60125 -210 60325 -125
rect 60475 -85 60675 -10
rect 60475 -125 60555 -85
rect 60595 -125 60675 -85
rect 60475 -210 60675 -125
rect 60825 -85 61025 -10
rect 60825 -125 60905 -85
rect 60945 -125 61025 -85
rect 60825 -210 61025 -125
rect 61175 -85 61375 -10
rect 61175 -125 61255 -85
rect 61295 -125 61375 -85
rect 61175 -210 61375 -125
rect 61525 -85 61725 -10
rect 61525 -125 61605 -85
rect 61645 -125 61725 -85
rect 61525 -210 61725 -125
rect 52075 -435 52275 -360
rect 52075 -475 52155 -435
rect 52195 -475 52275 -435
rect 52075 -560 52275 -475
rect 52425 -435 52625 -360
rect 52425 -475 52505 -435
rect 52545 -475 52625 -435
rect 52425 -560 52625 -475
rect 52775 -435 52975 -360
rect 52775 -475 52855 -435
rect 52895 -475 52975 -435
rect 52775 -560 52975 -475
rect 53125 -435 53325 -360
rect 53125 -475 53205 -435
rect 53245 -475 53325 -435
rect 53125 -560 53325 -475
rect 53475 -435 53675 -360
rect 53475 -475 53555 -435
rect 53595 -475 53675 -435
rect 53475 -560 53675 -475
rect 60125 -435 60325 -360
rect 60125 -475 60205 -435
rect 60245 -475 60325 -435
rect 60125 -560 60325 -475
rect 60475 -435 60675 -360
rect 60475 -475 60555 -435
rect 60595 -475 60675 -435
rect 60475 -560 60675 -475
rect 60825 -435 61025 -360
rect 60825 -475 60905 -435
rect 60945 -475 61025 -435
rect 60825 -560 61025 -475
rect 61175 -435 61375 -360
rect 61175 -475 61255 -435
rect 61295 -475 61375 -435
rect 61175 -560 61375 -475
rect 61525 -435 61725 -360
rect 61525 -475 61605 -435
rect 61645 -475 61725 -435
rect 61525 -560 61725 -475
rect 52075 -785 52275 -710
rect 52075 -825 52155 -785
rect 52195 -825 52275 -785
rect 52075 -910 52275 -825
rect 52425 -785 52625 -710
rect 52425 -825 52505 -785
rect 52545 -825 52625 -785
rect 52425 -910 52625 -825
rect 52775 -785 52975 -710
rect 52775 -825 52855 -785
rect 52895 -825 52975 -785
rect 52775 -910 52975 -825
rect 53125 -785 53325 -710
rect 53125 -825 53205 -785
rect 53245 -825 53325 -785
rect 53125 -910 53325 -825
rect 53475 -785 53675 -710
rect 53475 -825 53555 -785
rect 53595 -825 53675 -785
rect 53475 -910 53675 -825
rect 53825 -785 54025 -710
rect 53825 -825 53905 -785
rect 53945 -825 54025 -785
rect 53825 -910 54025 -825
rect 54175 -785 54375 -710
rect 54175 -825 54255 -785
rect 54295 -825 54375 -785
rect 54175 -910 54375 -825
rect 54525 -785 54725 -710
rect 54525 -825 54605 -785
rect 54645 -825 54725 -785
rect 54525 -910 54725 -825
rect 54875 -785 55075 -710
rect 54875 -825 54955 -785
rect 54995 -825 55075 -785
rect 54875 -910 55075 -825
rect 55225 -785 55425 -710
rect 55225 -825 55305 -785
rect 55345 -825 55425 -785
rect 55225 -910 55425 -825
rect 55575 -785 55775 -710
rect 55575 -825 55655 -785
rect 55695 -825 55775 -785
rect 55575 -910 55775 -825
rect 55925 -785 56125 -710
rect 55925 -825 56005 -785
rect 56045 -825 56125 -785
rect 55925 -910 56125 -825
rect 56275 -785 56475 -710
rect 56275 -825 56355 -785
rect 56395 -825 56475 -785
rect 56275 -910 56475 -825
rect 56625 -785 56825 -710
rect 56625 -825 56705 -785
rect 56745 -825 56825 -785
rect 56625 -910 56825 -825
rect 56975 -785 57175 -710
rect 56975 -825 57055 -785
rect 57095 -825 57175 -785
rect 56975 -910 57175 -825
rect 57325 -785 57525 -710
rect 57325 -825 57405 -785
rect 57445 -825 57525 -785
rect 57325 -910 57525 -825
rect 57675 -785 57875 -710
rect 57675 -825 57755 -785
rect 57795 -825 57875 -785
rect 57675 -910 57875 -825
rect 58025 -785 58225 -710
rect 58025 -825 58105 -785
rect 58145 -825 58225 -785
rect 58025 -910 58225 -825
rect 58375 -785 58575 -710
rect 58375 -825 58455 -785
rect 58495 -825 58575 -785
rect 58375 -910 58575 -825
rect 58725 -785 58925 -710
rect 58725 -825 58805 -785
rect 58845 -825 58925 -785
rect 58725 -910 58925 -825
rect 59075 -785 59275 -710
rect 59075 -825 59155 -785
rect 59195 -825 59275 -785
rect 59075 -910 59275 -825
rect 59425 -785 59625 -710
rect 59425 -825 59505 -785
rect 59545 -825 59625 -785
rect 59425 -910 59625 -825
rect 59775 -785 59975 -710
rect 59775 -825 59855 -785
rect 59895 -825 59975 -785
rect 59775 -910 59975 -825
rect 60125 -785 60325 -710
rect 60125 -825 60205 -785
rect 60245 -825 60325 -785
rect 60125 -910 60325 -825
rect 60475 -785 60675 -710
rect 60475 -825 60555 -785
rect 60595 -825 60675 -785
rect 60475 -910 60675 -825
rect 60825 -785 61025 -710
rect 60825 -825 60905 -785
rect 60945 -825 61025 -785
rect 60825 -910 61025 -825
rect 61175 -785 61375 -710
rect 61175 -825 61255 -785
rect 61295 -825 61375 -785
rect 61175 -910 61375 -825
rect 61525 -785 61725 -710
rect 61525 -825 61605 -785
rect 61645 -825 61725 -785
rect 61525 -910 61725 -825
rect 52075 -1135 52275 -1060
rect 52075 -1175 52155 -1135
rect 52195 -1175 52275 -1135
rect 52075 -1260 52275 -1175
rect 52425 -1135 52625 -1060
rect 52425 -1175 52505 -1135
rect 52545 -1175 52625 -1135
rect 52425 -1260 52625 -1175
rect 52775 -1135 52975 -1060
rect 52775 -1175 52855 -1135
rect 52895 -1175 52975 -1135
rect 52775 -1260 52975 -1175
rect 53125 -1135 53325 -1060
rect 53125 -1175 53205 -1135
rect 53245 -1175 53325 -1135
rect 53125 -1260 53325 -1175
rect 53475 -1135 53675 -1060
rect 53475 -1175 53555 -1135
rect 53595 -1175 53675 -1135
rect 53475 -1260 53675 -1175
rect 53825 -1135 54025 -1060
rect 53825 -1175 53905 -1135
rect 53945 -1175 54025 -1135
rect 53825 -1260 54025 -1175
rect 54175 -1135 54375 -1060
rect 54175 -1175 54255 -1135
rect 54295 -1175 54375 -1135
rect 54175 -1260 54375 -1175
rect 54525 -1135 54725 -1060
rect 54525 -1175 54605 -1135
rect 54645 -1175 54725 -1135
rect 54525 -1260 54725 -1175
rect 54875 -1135 55075 -1060
rect 54875 -1175 54955 -1135
rect 54995 -1175 55075 -1135
rect 54875 -1260 55075 -1175
rect 55225 -1135 55425 -1060
rect 55225 -1175 55305 -1135
rect 55345 -1175 55425 -1135
rect 55225 -1260 55425 -1175
rect 55575 -1135 55775 -1060
rect 55575 -1175 55655 -1135
rect 55695 -1175 55775 -1135
rect 55575 -1260 55775 -1175
rect 55925 -1135 56125 -1060
rect 55925 -1175 56005 -1135
rect 56045 -1175 56125 -1135
rect 55925 -1260 56125 -1175
rect 56275 -1135 56475 -1060
rect 56275 -1175 56355 -1135
rect 56395 -1175 56475 -1135
rect 56275 -1260 56475 -1175
rect 56625 -1135 56825 -1060
rect 56625 -1175 56705 -1135
rect 56745 -1175 56825 -1135
rect 56625 -1260 56825 -1175
rect 56975 -1135 57175 -1060
rect 56975 -1175 57055 -1135
rect 57095 -1175 57175 -1135
rect 56975 -1260 57175 -1175
rect 57325 -1135 57525 -1060
rect 57325 -1175 57405 -1135
rect 57445 -1175 57525 -1135
rect 57325 -1260 57525 -1175
rect 57675 -1135 57875 -1060
rect 57675 -1175 57755 -1135
rect 57795 -1175 57875 -1135
rect 57675 -1260 57875 -1175
rect 58025 -1135 58225 -1060
rect 58025 -1175 58105 -1135
rect 58145 -1175 58225 -1135
rect 58025 -1260 58225 -1175
rect 58375 -1135 58575 -1060
rect 58375 -1175 58455 -1135
rect 58495 -1175 58575 -1135
rect 58375 -1260 58575 -1175
rect 58725 -1135 58925 -1060
rect 58725 -1175 58805 -1135
rect 58845 -1175 58925 -1135
rect 58725 -1260 58925 -1175
rect 59075 -1135 59275 -1060
rect 59075 -1175 59155 -1135
rect 59195 -1175 59275 -1135
rect 59075 -1260 59275 -1175
rect 59425 -1135 59625 -1060
rect 59425 -1175 59505 -1135
rect 59545 -1175 59625 -1135
rect 59425 -1260 59625 -1175
rect 59775 -1135 59975 -1060
rect 59775 -1175 59855 -1135
rect 59895 -1175 59975 -1135
rect 59775 -1260 59975 -1175
rect 60125 -1135 60325 -1060
rect 60125 -1175 60205 -1135
rect 60245 -1175 60325 -1135
rect 60125 -1260 60325 -1175
rect 60475 -1135 60675 -1060
rect 60475 -1175 60555 -1135
rect 60595 -1175 60675 -1135
rect 60475 -1260 60675 -1175
rect 60825 -1135 61025 -1060
rect 60825 -1175 60905 -1135
rect 60945 -1175 61025 -1135
rect 60825 -1260 61025 -1175
rect 61175 -1135 61375 -1060
rect 61175 -1175 61255 -1135
rect 61295 -1175 61375 -1135
rect 61175 -1260 61375 -1175
rect 61525 -1135 61725 -1060
rect 61525 -1175 61605 -1135
rect 61645 -1175 61725 -1135
rect 61525 -1260 61725 -1175
<< mimcapcontact >>
rect 52155 6175 52195 6215
rect 52505 6175 52545 6215
rect 52855 6175 52895 6215
rect 53205 6175 53245 6215
rect 53555 6175 53595 6215
rect 53905 6175 53945 6215
rect 54255 6175 54295 6215
rect 54605 6175 54645 6215
rect 54955 6175 54995 6215
rect 55305 6175 55345 6215
rect 55655 6175 55695 6215
rect 56005 6175 56045 6215
rect 56355 6175 56395 6215
rect 56705 6175 56745 6215
rect 57055 6175 57095 6215
rect 57405 6175 57445 6215
rect 57755 6175 57795 6215
rect 58105 6175 58145 6215
rect 58455 6175 58495 6215
rect 58805 6175 58845 6215
rect 59155 6175 59195 6215
rect 59505 6175 59545 6215
rect 59855 6175 59895 6215
rect 60205 6175 60245 6215
rect 60555 6175 60595 6215
rect 60905 6175 60945 6215
rect 61255 6175 61295 6215
rect 61605 6175 61645 6215
rect 52155 5825 52195 5865
rect 52505 5825 52545 5865
rect 52855 5825 52895 5865
rect 53205 5825 53245 5865
rect 53555 5825 53595 5865
rect 53905 5825 53945 5865
rect 54255 5825 54295 5865
rect 54605 5825 54645 5865
rect 54955 5825 54995 5865
rect 55305 5825 55345 5865
rect 55655 5825 55695 5865
rect 56005 5825 56045 5865
rect 56355 5825 56395 5865
rect 56705 5825 56745 5865
rect 57055 5825 57095 5865
rect 57405 5825 57445 5865
rect 57755 5825 57795 5865
rect 58105 5825 58145 5865
rect 58455 5825 58495 5865
rect 58805 5825 58845 5865
rect 59155 5825 59195 5865
rect 59505 5825 59545 5865
rect 59855 5825 59895 5865
rect 60205 5825 60245 5865
rect 60555 5825 60595 5865
rect 60905 5825 60945 5865
rect 61255 5825 61295 5865
rect 61605 5825 61645 5865
rect 52155 5475 52195 5515
rect 52505 5475 52545 5515
rect 52855 5475 52895 5515
rect 53205 5475 53245 5515
rect 53555 5475 53595 5515
rect 53905 5475 53945 5515
rect 54255 5475 54295 5515
rect 54605 5475 54645 5515
rect 54955 5475 54995 5515
rect 55305 5465 55345 5505
rect 55655 5465 55695 5505
rect 56005 5465 56045 5505
rect 56355 5465 56395 5505
rect 56705 5465 56745 5505
rect 57055 5465 57095 5505
rect 57405 5465 57445 5505
rect 57755 5465 57795 5505
rect 58105 5465 58145 5505
rect 58455 5465 58495 5505
rect 58805 5475 58845 5515
rect 59155 5475 59195 5515
rect 59505 5475 59545 5515
rect 59855 5475 59895 5515
rect 60205 5475 60245 5515
rect 60555 5475 60595 5515
rect 60905 5475 60945 5515
rect 61255 5475 61295 5515
rect 61605 5475 61645 5515
rect 52155 5125 52195 5165
rect 52505 5125 52545 5165
rect 52855 5125 52895 5165
rect 53205 5125 53245 5165
rect 53555 5125 53595 5165
rect 53905 5125 53945 5165
rect 54255 5125 54295 5165
rect 54605 5125 54645 5165
rect 59155 5125 59195 5165
rect 59505 5125 59545 5165
rect 59855 5125 59895 5165
rect 60205 5125 60245 5165
rect 60555 5125 60595 5165
rect 60905 5125 60945 5165
rect 61255 5125 61295 5165
rect 61605 5125 61645 5165
rect 52155 4775 52195 4815
rect 52505 4775 52545 4815
rect 52855 4775 52895 4815
rect 53205 4775 53245 4815
rect 53555 4775 53595 4815
rect 60205 4775 60245 4815
rect 60555 4775 60595 4815
rect 60905 4775 60945 4815
rect 61255 4775 61295 4815
rect 61605 4775 61645 4815
rect 52155 4425 52195 4465
rect 52505 4425 52545 4465
rect 52855 4425 52895 4465
rect 53205 4425 53245 4465
rect 53555 4425 53595 4465
rect 60205 4425 60245 4465
rect 60555 4425 60595 4465
rect 60905 4425 60945 4465
rect 61255 4425 61295 4465
rect 61605 4425 61645 4465
rect 52155 4075 52195 4115
rect 52505 4075 52545 4115
rect 52855 4075 52895 4115
rect 53205 4075 53245 4115
rect 53555 4075 53595 4115
rect 60205 4075 60245 4115
rect 60555 4075 60595 4115
rect 60905 4075 60945 4115
rect 61255 4075 61295 4115
rect 61605 4075 61645 4115
rect 52155 3725 52195 3765
rect 52505 3725 52545 3765
rect 52855 3725 52895 3765
rect 53205 3725 53245 3765
rect 53555 3725 53595 3765
rect 60205 3725 60245 3765
rect 60555 3725 60595 3765
rect 60905 3725 60945 3765
rect 61255 3725 61295 3765
rect 61605 3725 61645 3765
rect 52155 3375 52195 3415
rect 52505 3375 52545 3415
rect 52855 3375 52895 3415
rect 53205 3375 53245 3415
rect 53555 3375 53595 3415
rect 60205 3375 60245 3415
rect 60555 3375 60595 3415
rect 60905 3375 60945 3415
rect 61255 3375 61295 3415
rect 61605 3375 61645 3415
rect 52155 3025 52195 3065
rect 52505 3025 52545 3065
rect 52855 3025 52895 3065
rect 53205 3025 53245 3065
rect 53555 3025 53595 3065
rect 60205 3025 60245 3065
rect 60555 3025 60595 3065
rect 60905 3025 60945 3065
rect 61255 3025 61295 3065
rect 61605 3025 61645 3065
rect 52155 2675 52195 2715
rect 52505 2675 52545 2715
rect 52855 2675 52895 2715
rect 53205 2675 53245 2715
rect 53555 2675 53595 2715
rect 60205 2675 60245 2715
rect 60555 2675 60595 2715
rect 60905 2675 60945 2715
rect 61255 2675 61295 2715
rect 61605 2675 61645 2715
rect 52155 2325 52195 2365
rect 52505 2325 52545 2365
rect 52855 2325 52895 2365
rect 53205 2325 53245 2365
rect 53555 2325 53595 2365
rect 60205 2325 60245 2365
rect 60555 2325 60595 2365
rect 60905 2325 60945 2365
rect 61255 2325 61295 2365
rect 61605 2325 61645 2365
rect 52155 1975 52195 2015
rect 52505 1975 52545 2015
rect 52855 1975 52895 2015
rect 53205 1975 53245 2015
rect 53555 1975 53595 2015
rect 60205 1975 60245 2015
rect 60555 1975 60595 2015
rect 60905 1975 60945 2015
rect 61255 1975 61295 2015
rect 61605 1975 61645 2015
rect 52155 1625 52195 1665
rect 52505 1625 52545 1665
rect 52855 1625 52895 1665
rect 53205 1625 53245 1665
rect 53555 1625 53595 1665
rect 60205 1625 60245 1665
rect 60555 1625 60595 1665
rect 60905 1625 60945 1665
rect 61255 1625 61295 1665
rect 61605 1625 61645 1665
rect 52155 1275 52195 1315
rect 52505 1275 52545 1315
rect 52855 1275 52895 1315
rect 53205 1275 53245 1315
rect 53555 1275 53595 1315
rect 60205 1275 60245 1315
rect 60555 1275 60595 1315
rect 60905 1275 60945 1315
rect 61255 1275 61295 1315
rect 61605 1275 61645 1315
rect 52155 925 52195 965
rect 52505 925 52545 965
rect 52855 925 52895 965
rect 53205 925 53245 965
rect 53555 925 53595 965
rect 60205 925 60245 965
rect 60555 925 60595 965
rect 60905 925 60945 965
rect 61255 925 61295 965
rect 61605 925 61645 965
rect 52155 575 52195 615
rect 52505 575 52545 615
rect 52855 575 52895 615
rect 53205 575 53245 615
rect 53555 575 53595 615
rect 60205 575 60245 615
rect 60555 575 60595 615
rect 60905 575 60945 615
rect 61255 575 61295 615
rect 61605 575 61645 615
rect 52155 225 52195 265
rect 52505 225 52545 265
rect 52855 225 52895 265
rect 53205 225 53245 265
rect 53555 225 53595 265
rect 60205 225 60245 265
rect 60555 225 60595 265
rect 60905 225 60945 265
rect 61255 225 61295 265
rect 61605 225 61645 265
rect 52155 -125 52195 -85
rect 52505 -125 52545 -85
rect 52855 -125 52895 -85
rect 53205 -125 53245 -85
rect 53555 -125 53595 -85
rect 60205 -125 60245 -85
rect 60555 -125 60595 -85
rect 60905 -125 60945 -85
rect 61255 -125 61295 -85
rect 61605 -125 61645 -85
rect 52155 -475 52195 -435
rect 52505 -475 52545 -435
rect 52855 -475 52895 -435
rect 53205 -475 53245 -435
rect 53555 -475 53595 -435
rect 60205 -475 60245 -435
rect 60555 -475 60595 -435
rect 60905 -475 60945 -435
rect 61255 -475 61295 -435
rect 61605 -475 61645 -435
rect 52155 -825 52195 -785
rect 52505 -825 52545 -785
rect 52855 -825 52895 -785
rect 53205 -825 53245 -785
rect 53555 -825 53595 -785
rect 53905 -825 53945 -785
rect 54255 -825 54295 -785
rect 54605 -825 54645 -785
rect 54955 -825 54995 -785
rect 55305 -825 55345 -785
rect 55655 -825 55695 -785
rect 56005 -825 56045 -785
rect 56355 -825 56395 -785
rect 56705 -825 56745 -785
rect 57055 -825 57095 -785
rect 57405 -825 57445 -785
rect 57755 -825 57795 -785
rect 58105 -825 58145 -785
rect 58455 -825 58495 -785
rect 58805 -825 58845 -785
rect 59155 -825 59195 -785
rect 59505 -825 59545 -785
rect 59855 -825 59895 -785
rect 60205 -825 60245 -785
rect 60555 -825 60595 -785
rect 60905 -825 60945 -785
rect 61255 -825 61295 -785
rect 61605 -825 61645 -785
rect 52155 -1175 52195 -1135
rect 52505 -1175 52545 -1135
rect 52855 -1175 52895 -1135
rect 53205 -1175 53245 -1135
rect 53555 -1175 53595 -1135
rect 53905 -1175 53945 -1135
rect 54255 -1175 54295 -1135
rect 54605 -1175 54645 -1135
rect 54955 -1175 54995 -1135
rect 55305 -1175 55345 -1135
rect 55655 -1175 55695 -1135
rect 56005 -1175 56045 -1135
rect 56355 -1175 56395 -1135
rect 56705 -1175 56745 -1135
rect 57055 -1175 57095 -1135
rect 57405 -1175 57445 -1135
rect 57755 -1175 57795 -1135
rect 58105 -1175 58145 -1135
rect 58455 -1175 58495 -1135
rect 58805 -1175 58845 -1135
rect 59155 -1175 59195 -1135
rect 59505 -1175 59545 -1135
rect 59855 -1175 59895 -1135
rect 60205 -1175 60245 -1135
rect 60555 -1175 60595 -1135
rect 60905 -1175 60945 -1135
rect 61255 -1175 61295 -1135
rect 61605 -1175 61645 -1135
<< metal4 >>
rect 52150 6215 52900 6220
rect 52150 6175 52155 6215
rect 52195 6175 52505 6215
rect 52545 6175 52855 6215
rect 52895 6175 52900 6215
rect 52150 6170 52900 6175
rect 52850 5870 52900 6170
rect 53200 6215 53250 6220
rect 53200 6175 53205 6215
rect 53245 6175 53250 6215
rect 53200 5870 53250 6175
rect 53550 6215 53600 6220
rect 53550 6175 53555 6215
rect 53595 6175 53600 6215
rect 53550 5870 53600 6175
rect 53900 6215 53950 6220
rect 53900 6175 53905 6215
rect 53945 6175 53950 6215
rect 53900 5870 53950 6175
rect 54250 6215 54300 6220
rect 54250 6175 54255 6215
rect 54295 6175 54300 6215
rect 54250 5870 54300 6175
rect 54600 6215 54650 6220
rect 54600 6175 54605 6215
rect 54645 6175 54650 6215
rect 54600 5870 54650 6175
rect 54950 6215 55000 6220
rect 54950 6175 54955 6215
rect 54995 6175 55000 6215
rect 54950 5870 55000 6175
rect 55300 6215 55350 6220
rect 55300 6175 55305 6215
rect 55345 6175 55350 6215
rect 55300 5870 55350 6175
rect 55650 6215 55700 6220
rect 55650 6175 55655 6215
rect 55695 6175 55700 6215
rect 55650 5870 55700 6175
rect 56000 6215 56050 6220
rect 56000 6175 56005 6215
rect 56045 6175 56050 6215
rect 56000 5870 56050 6175
rect 56350 6215 56400 6220
rect 56350 6175 56355 6215
rect 56395 6175 56400 6215
rect 56350 5870 56400 6175
rect 56700 6215 56750 6220
rect 56700 6175 56705 6215
rect 56745 6175 56750 6215
rect 56700 5870 56750 6175
rect 52150 5865 56750 5870
rect 52150 5825 52155 5865
rect 52195 5825 52505 5865
rect 52545 5825 52855 5865
rect 52895 5825 53205 5865
rect 53245 5825 53555 5865
rect 53595 5825 53905 5865
rect 53945 5825 54255 5865
rect 54295 5825 54605 5865
rect 54645 5825 54955 5865
rect 54995 5825 55305 5865
rect 55345 5825 55655 5865
rect 55695 5825 56005 5865
rect 56045 5825 56355 5865
rect 56395 5825 56705 5865
rect 56745 5825 56750 5865
rect 52150 5820 56750 5825
rect 52850 5520 52900 5820
rect 52150 5515 53600 5520
rect 52150 5475 52155 5515
rect 52195 5475 52505 5515
rect 52545 5475 52855 5515
rect 52895 5475 53205 5515
rect 53245 5475 53555 5515
rect 53595 5475 53600 5515
rect 52150 5470 53600 5475
rect 53900 5515 53950 5820
rect 53900 5475 53905 5515
rect 53945 5475 53950 5515
rect 52850 5170 52900 5470
rect 52150 5165 53600 5170
rect 52150 5125 52155 5165
rect 52195 5125 52505 5165
rect 52545 5125 52855 5165
rect 52895 5125 53205 5165
rect 53245 5125 53555 5165
rect 53595 5125 53600 5165
rect 52150 5120 53600 5125
rect 53900 5165 53950 5475
rect 53900 5125 53905 5165
rect 53945 5125 53950 5165
rect 53900 5120 53950 5125
rect 54250 5515 54300 5820
rect 54250 5475 54255 5515
rect 54295 5475 54300 5515
rect 54250 5165 54300 5475
rect 54250 5125 54255 5165
rect 54295 5125 54300 5165
rect 54250 5120 54300 5125
rect 54600 5515 54650 5820
rect 54600 5475 54605 5515
rect 54645 5475 54650 5515
rect 54600 5165 54650 5475
rect 54950 5515 55000 5820
rect 54950 5475 54955 5515
rect 54995 5475 55000 5515
rect 54950 5470 55000 5475
rect 55300 5505 55350 5820
rect 55300 5465 55305 5505
rect 55345 5465 55350 5505
rect 55300 5460 55350 5465
rect 55650 5505 55700 5820
rect 55650 5465 55655 5505
rect 55695 5465 55700 5505
rect 55650 5460 55700 5465
rect 56000 5505 56050 5820
rect 56000 5465 56005 5505
rect 56045 5465 56050 5505
rect 56000 5460 56050 5465
rect 56350 5505 56400 5820
rect 56350 5465 56355 5505
rect 56395 5465 56400 5505
rect 56350 5460 56400 5465
rect 56700 5505 56750 5820
rect 56700 5465 56705 5505
rect 56745 5465 56750 5505
rect 56700 5460 56750 5465
rect 57050 6215 57100 6220
rect 57050 6175 57055 6215
rect 57095 6175 57100 6215
rect 57050 5870 57100 6175
rect 57400 6215 57450 6220
rect 57400 6175 57405 6215
rect 57445 6175 57450 6215
rect 57400 5870 57450 6175
rect 57750 6215 57800 6220
rect 57750 6175 57755 6215
rect 57795 6175 57800 6215
rect 57750 5870 57800 6175
rect 58100 6215 58150 6220
rect 58100 6175 58105 6215
rect 58145 6175 58150 6215
rect 58100 5870 58150 6175
rect 58450 6215 58500 6220
rect 58450 6175 58455 6215
rect 58495 6175 58500 6215
rect 58450 5870 58500 6175
rect 58800 6215 58850 6220
rect 58800 6175 58805 6215
rect 58845 6175 58850 6215
rect 58800 5870 58850 6175
rect 59150 6215 59200 6220
rect 59150 6175 59155 6215
rect 59195 6175 59200 6215
rect 59150 5870 59200 6175
rect 59500 6215 59550 6220
rect 59500 6175 59505 6215
rect 59545 6175 59550 6215
rect 59500 5870 59550 6175
rect 59850 6215 59900 6220
rect 59850 6175 59855 6215
rect 59895 6175 59900 6215
rect 59850 5870 59900 6175
rect 60200 6215 60250 6220
rect 60200 6175 60205 6215
rect 60245 6175 60250 6215
rect 60200 5870 60250 6175
rect 60550 6215 60600 6220
rect 60550 6175 60555 6215
rect 60595 6175 60600 6215
rect 60550 5870 60600 6175
rect 60900 6215 61650 6220
rect 60900 6175 60905 6215
rect 60945 6175 61255 6215
rect 61295 6175 61605 6215
rect 61645 6175 61650 6215
rect 60900 6170 61650 6175
rect 60900 5870 60950 6170
rect 57050 5865 61650 5870
rect 57050 5825 57055 5865
rect 57095 5825 57405 5865
rect 57445 5825 57755 5865
rect 57795 5825 58105 5865
rect 58145 5825 58455 5865
rect 58495 5825 58805 5865
rect 58845 5825 59155 5865
rect 59195 5825 59505 5865
rect 59545 5825 59855 5865
rect 59895 5825 60205 5865
rect 60245 5825 60555 5865
rect 60595 5825 60905 5865
rect 60945 5825 61255 5865
rect 61295 5825 61605 5865
rect 61645 5825 61650 5865
rect 57050 5820 61650 5825
rect 57050 5505 57100 5820
rect 57050 5465 57055 5505
rect 57095 5465 57100 5505
rect 57050 5460 57100 5465
rect 57400 5505 57450 5820
rect 57400 5465 57405 5505
rect 57445 5465 57450 5505
rect 57400 5460 57450 5465
rect 57750 5505 57800 5820
rect 57750 5465 57755 5505
rect 57795 5465 57800 5505
rect 57750 5460 57800 5465
rect 58100 5505 58150 5820
rect 58100 5465 58105 5505
rect 58145 5465 58150 5505
rect 58100 5460 58150 5465
rect 58450 5505 58500 5820
rect 58450 5465 58455 5505
rect 58495 5465 58500 5505
rect 58800 5515 58850 5820
rect 58800 5475 58805 5515
rect 58845 5475 58850 5515
rect 58800 5470 58850 5475
rect 59150 5515 59200 5820
rect 59150 5475 59155 5515
rect 59195 5475 59200 5515
rect 58450 5460 58500 5465
rect 54600 5125 54605 5165
rect 54645 5125 54650 5165
rect 54600 5120 54650 5125
rect 59150 5165 59200 5475
rect 59150 5125 59155 5165
rect 59195 5125 59200 5165
rect 59150 5120 59200 5125
rect 59500 5515 59550 5820
rect 59500 5475 59505 5515
rect 59545 5475 59550 5515
rect 59500 5165 59550 5475
rect 59500 5125 59505 5165
rect 59545 5125 59550 5165
rect 59500 5120 59550 5125
rect 59850 5515 59900 5820
rect 60900 5520 60950 5820
rect 59850 5475 59855 5515
rect 59895 5475 59900 5515
rect 59850 5165 59900 5475
rect 60200 5515 61650 5520
rect 60200 5475 60205 5515
rect 60245 5475 60555 5515
rect 60595 5475 60905 5515
rect 60945 5475 61255 5515
rect 61295 5475 61605 5515
rect 61645 5475 61650 5515
rect 60200 5470 61650 5475
rect 60900 5170 60950 5470
rect 59850 5125 59855 5165
rect 59895 5125 59900 5165
rect 59850 5120 59900 5125
rect 60200 5165 61650 5170
rect 60200 5125 60205 5165
rect 60245 5125 60555 5165
rect 60595 5125 60905 5165
rect 60945 5125 61255 5165
rect 61295 5125 61605 5165
rect 61645 5125 61650 5165
rect 60200 5120 61650 5125
rect 52850 4820 52900 5120
rect 60900 4820 60950 5120
rect 52150 4815 53600 4820
rect 52150 4775 52155 4815
rect 52195 4775 52505 4815
rect 52545 4775 52855 4815
rect 52895 4775 53205 4815
rect 53245 4775 53555 4815
rect 53595 4775 53600 4815
rect 52150 4770 53600 4775
rect 60200 4815 61650 4820
rect 60200 4775 60205 4815
rect 60245 4775 60555 4815
rect 60595 4775 60905 4815
rect 60945 4775 61255 4815
rect 61295 4775 61605 4815
rect 61645 4775 61650 4815
rect 60200 4770 61650 4775
rect 52850 4470 52900 4770
rect 60900 4470 60950 4770
rect 52150 4465 53600 4470
rect 52150 4425 52155 4465
rect 52195 4425 52505 4465
rect 52545 4425 52855 4465
rect 52895 4425 53205 4465
rect 53245 4425 53555 4465
rect 53595 4425 53600 4465
rect 52150 4420 53600 4425
rect 60200 4465 61650 4470
rect 60200 4425 60205 4465
rect 60245 4425 60555 4465
rect 60595 4425 60905 4465
rect 60945 4425 61255 4465
rect 61295 4425 61605 4465
rect 61645 4425 61650 4465
rect 60200 4420 61650 4425
rect 52850 4120 52900 4420
rect 60900 4120 60950 4420
rect 52150 4115 53600 4120
rect 52150 4075 52155 4115
rect 52195 4075 52505 4115
rect 52545 4075 52855 4115
rect 52895 4075 53205 4115
rect 53245 4075 53555 4115
rect 53595 4075 53600 4115
rect 52150 4070 53600 4075
rect 60200 4115 61650 4120
rect 60200 4075 60205 4115
rect 60245 4075 60555 4115
rect 60595 4075 60905 4115
rect 60945 4075 61255 4115
rect 61295 4075 61605 4115
rect 61645 4075 61650 4115
rect 60200 4070 61650 4075
rect 52850 3770 52900 4070
rect 60900 3770 60950 4070
rect 52150 3765 53600 3770
rect 52150 3725 52155 3765
rect 52195 3725 52505 3765
rect 52545 3725 52855 3765
rect 52895 3725 53205 3765
rect 53245 3725 53555 3765
rect 53595 3725 53600 3765
rect 52150 3720 53600 3725
rect 60200 3765 61650 3770
rect 60200 3725 60205 3765
rect 60245 3725 60555 3765
rect 60595 3725 60905 3765
rect 60945 3725 61255 3765
rect 61295 3725 61605 3765
rect 61645 3725 61650 3765
rect 60200 3720 61650 3725
rect 52850 3420 52900 3720
rect 60900 3420 60950 3720
rect 52150 3415 53600 3420
rect 52150 3375 52155 3415
rect 52195 3375 52505 3415
rect 52545 3375 52855 3415
rect 52895 3375 53205 3415
rect 53245 3375 53555 3415
rect 53595 3375 53600 3415
rect 52150 3370 53600 3375
rect 60200 3415 61650 3420
rect 60200 3375 60205 3415
rect 60245 3375 60555 3415
rect 60595 3375 60905 3415
rect 60945 3375 61255 3415
rect 61295 3375 61605 3415
rect 61645 3375 61650 3415
rect 60200 3370 61650 3375
rect 52850 3070 52900 3370
rect 60900 3070 60950 3370
rect 52150 3065 53600 3070
rect 52150 3025 52155 3065
rect 52195 3025 52505 3065
rect 52545 3025 52855 3065
rect 52895 3025 53205 3065
rect 53245 3025 53555 3065
rect 53595 3025 53600 3065
rect 52150 3020 53600 3025
rect 60200 3065 61650 3070
rect 60200 3025 60205 3065
rect 60245 3025 60555 3065
rect 60595 3025 60905 3065
rect 60945 3025 61255 3065
rect 61295 3025 61605 3065
rect 61645 3025 61650 3065
rect 60200 3020 61650 3025
rect 52850 2720 52900 3020
rect 60900 2720 60950 3020
rect 52150 2715 53600 2720
rect 52150 2675 52155 2715
rect 52195 2675 52505 2715
rect 52545 2675 52855 2715
rect 52895 2675 53205 2715
rect 53245 2675 53555 2715
rect 53595 2675 53600 2715
rect 52150 2670 53600 2675
rect 60200 2715 61650 2720
rect 60200 2675 60205 2715
rect 60245 2675 60555 2715
rect 60595 2675 60905 2715
rect 60945 2675 61255 2715
rect 61295 2675 61605 2715
rect 61645 2675 61650 2715
rect 60200 2670 61650 2675
rect 52850 2370 52900 2670
rect 60900 2370 60950 2670
rect 52150 2365 53600 2370
rect 52150 2325 52155 2365
rect 52195 2325 52505 2365
rect 52545 2325 52855 2365
rect 52895 2325 53205 2365
rect 53245 2325 53555 2365
rect 53595 2325 53600 2365
rect 52150 2320 53600 2325
rect 60200 2365 61650 2370
rect 60200 2325 60205 2365
rect 60245 2325 60555 2365
rect 60595 2325 60905 2365
rect 60945 2325 61255 2365
rect 61295 2325 61605 2365
rect 61645 2325 61650 2365
rect 60200 2320 61650 2325
rect 52850 2020 52900 2320
rect 60900 2020 60950 2320
rect 52150 2015 53600 2020
rect 52150 1975 52155 2015
rect 52195 1975 52505 2015
rect 52545 1975 52855 2015
rect 52895 1975 53205 2015
rect 53245 1975 53555 2015
rect 53595 1975 53600 2015
rect 52150 1970 53600 1975
rect 60200 2015 61650 2020
rect 60200 1975 60205 2015
rect 60245 1975 60555 2015
rect 60595 1975 60905 2015
rect 60945 1975 61255 2015
rect 61295 1975 61605 2015
rect 61645 1975 61650 2015
rect 60200 1970 61650 1975
rect 52850 1670 52900 1970
rect 60900 1670 60950 1970
rect 52150 1665 53600 1670
rect 52150 1625 52155 1665
rect 52195 1625 52505 1665
rect 52545 1625 52855 1665
rect 52895 1625 53205 1665
rect 53245 1625 53555 1665
rect 53595 1625 53600 1665
rect 52150 1620 53600 1625
rect 60200 1665 61650 1670
rect 60200 1625 60205 1665
rect 60245 1625 60555 1665
rect 60595 1625 60905 1665
rect 60945 1625 61255 1665
rect 61295 1625 61605 1665
rect 61645 1625 61650 1665
rect 60200 1620 61650 1625
rect 52850 1320 52900 1620
rect 59715 1440 60110 1445
rect 59715 1400 59720 1440
rect 59760 1400 59770 1440
rect 59810 1400 59820 1440
rect 59860 1400 59870 1440
rect 59910 1400 59920 1440
rect 59960 1400 60110 1440
rect 59715 1390 60110 1400
rect 53550 1365 54355 1370
rect 53550 1325 54110 1365
rect 54150 1325 54160 1365
rect 54200 1325 54210 1365
rect 54250 1325 54260 1365
rect 54300 1325 54310 1365
rect 54350 1325 54355 1365
rect 53550 1320 54355 1325
rect 52150 1315 54355 1320
rect 52150 1275 52155 1315
rect 52195 1275 52505 1315
rect 52545 1275 52855 1315
rect 52895 1275 53205 1315
rect 53245 1275 53555 1315
rect 53595 1275 54110 1315
rect 54150 1275 54160 1315
rect 54200 1275 54210 1315
rect 54250 1275 54260 1315
rect 54300 1275 54310 1315
rect 54350 1275 54355 1315
rect 59715 1350 59720 1390
rect 59760 1350 59770 1390
rect 59810 1350 59820 1390
rect 59860 1350 59870 1390
rect 59910 1350 59920 1390
rect 59960 1370 60110 1390
rect 59960 1350 60255 1370
rect 59715 1340 60255 1350
rect 59715 1300 59720 1340
rect 59760 1300 59770 1340
rect 59810 1300 59820 1340
rect 59860 1300 59870 1340
rect 59910 1300 59920 1340
rect 59960 1320 60255 1340
rect 60900 1320 60950 1620
rect 59960 1315 61650 1320
rect 59960 1300 60205 1315
rect 59715 1295 60205 1300
rect 52150 1270 54355 1275
rect 52850 970 52900 1270
rect 53550 1265 54355 1270
rect 53550 1225 54110 1265
rect 54150 1225 54160 1265
rect 54200 1225 54210 1265
rect 54250 1225 54260 1265
rect 54300 1225 54310 1265
rect 54350 1225 54355 1265
rect 53550 1220 54355 1225
rect 60110 1275 60205 1295
rect 60245 1275 60555 1315
rect 60595 1275 60905 1315
rect 60945 1275 61255 1315
rect 61295 1275 61605 1315
rect 61645 1275 61650 1315
rect 60110 1270 61650 1275
rect 60110 1220 60255 1270
rect 60900 970 60950 1270
rect 52150 965 53600 970
rect 52150 925 52155 965
rect 52195 925 52505 965
rect 52545 925 52855 965
rect 52895 925 53205 965
rect 53245 925 53555 965
rect 53595 925 53600 965
rect 52150 920 53600 925
rect 60200 965 61650 970
rect 60200 925 60205 965
rect 60245 925 60555 965
rect 60595 925 60905 965
rect 60945 925 61255 965
rect 61295 925 61605 965
rect 61645 925 61650 965
rect 60200 920 61650 925
rect 52850 620 52900 920
rect 60900 620 60950 920
rect 52150 615 53600 620
rect 52150 575 52155 615
rect 52195 575 52505 615
rect 52545 575 52855 615
rect 52895 575 53205 615
rect 53245 575 53555 615
rect 53595 575 53600 615
rect 52150 570 53600 575
rect 60200 615 61650 620
rect 60200 575 60205 615
rect 60245 575 60555 615
rect 60595 575 60905 615
rect 60945 575 61255 615
rect 61295 575 61605 615
rect 61645 575 61650 615
rect 60200 570 61650 575
rect 52850 270 52900 570
rect 60900 270 60950 570
rect 52150 265 53600 270
rect 52150 225 52155 265
rect 52195 225 52505 265
rect 52545 225 52855 265
rect 52895 225 53205 265
rect 53245 225 53555 265
rect 53595 225 53600 265
rect 52150 220 53600 225
rect 60200 265 61650 270
rect 60200 225 60205 265
rect 60245 225 60555 265
rect 60595 225 60905 265
rect 60945 225 61255 265
rect 61295 225 61605 265
rect 61645 225 61650 265
rect 60200 220 61650 225
rect 52850 -80 52900 220
rect 60900 -80 60950 220
rect 52150 -85 53600 -80
rect 52150 -125 52155 -85
rect 52195 -125 52505 -85
rect 52545 -125 52855 -85
rect 52895 -125 53205 -85
rect 53245 -125 53555 -85
rect 53595 -125 53600 -85
rect 52150 -130 53600 -125
rect 60200 -85 61650 -80
rect 60200 -125 60205 -85
rect 60245 -125 60555 -85
rect 60595 -125 60905 -85
rect 60945 -125 61255 -85
rect 61295 -125 61605 -85
rect 61645 -125 61650 -85
rect 60200 -130 61650 -125
rect 52850 -430 52900 -130
rect 60900 -430 60950 -130
rect 52150 -435 53600 -430
rect 52150 -475 52155 -435
rect 52195 -475 52505 -435
rect 52545 -475 52855 -435
rect 52895 -475 53205 -435
rect 53245 -475 53555 -435
rect 53595 -475 53600 -435
rect 52150 -480 53600 -475
rect 60200 -435 61650 -430
rect 60200 -475 60205 -435
rect 60245 -475 60555 -435
rect 60595 -475 60905 -435
rect 60945 -475 61255 -435
rect 61295 -475 61605 -435
rect 61645 -475 61650 -435
rect 60200 -480 61650 -475
rect 52850 -780 52900 -480
rect 60900 -780 60950 -480
rect 52150 -785 56750 -780
rect 52150 -825 52155 -785
rect 52195 -825 52505 -785
rect 52545 -825 52855 -785
rect 52895 -825 53205 -785
rect 53245 -825 53555 -785
rect 53595 -825 53905 -785
rect 53945 -825 54255 -785
rect 54295 -825 54605 -785
rect 54645 -825 54955 -785
rect 54995 -825 55305 -785
rect 55345 -825 55655 -785
rect 55695 -825 56005 -785
rect 56045 -825 56355 -785
rect 56395 -825 56705 -785
rect 56745 -825 56750 -785
rect 52150 -830 56750 -825
rect 52850 -1130 52900 -830
rect 52150 -1135 52900 -1130
rect 52150 -1175 52155 -1135
rect 52195 -1175 52505 -1135
rect 52545 -1175 52855 -1135
rect 52895 -1175 52900 -1135
rect 52150 -1180 52900 -1175
rect 53200 -1135 53250 -830
rect 53200 -1175 53205 -1135
rect 53245 -1175 53250 -1135
rect 53200 -1180 53250 -1175
rect 53550 -1135 53600 -830
rect 53550 -1175 53555 -1135
rect 53595 -1175 53600 -1135
rect 53550 -1180 53600 -1175
rect 53900 -1135 53950 -830
rect 53900 -1175 53905 -1135
rect 53945 -1175 53950 -1135
rect 53900 -1180 53950 -1175
rect 54250 -1135 54300 -830
rect 54250 -1175 54255 -1135
rect 54295 -1175 54300 -1135
rect 54250 -1180 54300 -1175
rect 54600 -1135 54650 -830
rect 54600 -1175 54605 -1135
rect 54645 -1175 54650 -1135
rect 54600 -1180 54650 -1175
rect 54950 -1135 55000 -830
rect 54950 -1175 54955 -1135
rect 54995 -1175 55000 -1135
rect 54950 -1180 55000 -1175
rect 55300 -1135 55350 -830
rect 55300 -1175 55305 -1135
rect 55345 -1175 55350 -1135
rect 55300 -1180 55350 -1175
rect 55650 -1135 55700 -830
rect 55650 -1175 55655 -1135
rect 55695 -1175 55700 -1135
rect 55650 -1180 55700 -1175
rect 56000 -1135 56050 -830
rect 56000 -1175 56005 -1135
rect 56045 -1175 56050 -1135
rect 56000 -1180 56050 -1175
rect 56350 -1135 56400 -830
rect 56350 -1175 56355 -1135
rect 56395 -1175 56400 -1135
rect 56350 -1180 56400 -1175
rect 56700 -1135 56750 -830
rect 56700 -1175 56705 -1135
rect 56745 -1175 56750 -1135
rect 56700 -1180 56750 -1175
rect 57050 -785 61650 -780
rect 57050 -825 57055 -785
rect 57095 -825 57405 -785
rect 57445 -825 57755 -785
rect 57795 -825 58105 -785
rect 58145 -825 58455 -785
rect 58495 -825 58805 -785
rect 58845 -825 59155 -785
rect 59195 -825 59505 -785
rect 59545 -825 59855 -785
rect 59895 -825 60205 -785
rect 60245 -825 60555 -785
rect 60595 -825 60905 -785
rect 60945 -825 61255 -785
rect 61295 -825 61605 -785
rect 61645 -825 61650 -785
rect 57050 -830 61650 -825
rect 57050 -1135 57100 -830
rect 57050 -1175 57055 -1135
rect 57095 -1175 57100 -1135
rect 57050 -1180 57100 -1175
rect 57400 -1135 57450 -830
rect 57400 -1175 57405 -1135
rect 57445 -1175 57450 -1135
rect 57400 -1180 57450 -1175
rect 57750 -1135 57800 -830
rect 57750 -1175 57755 -1135
rect 57795 -1175 57800 -1135
rect 57750 -1180 57800 -1175
rect 58100 -1135 58150 -830
rect 58100 -1175 58105 -1135
rect 58145 -1175 58150 -1135
rect 58100 -1180 58150 -1175
rect 58450 -1135 58500 -830
rect 58450 -1175 58455 -1135
rect 58495 -1175 58500 -1135
rect 58450 -1180 58500 -1175
rect 58800 -1135 58850 -830
rect 58800 -1175 58805 -1135
rect 58845 -1175 58850 -1135
rect 58800 -1180 58850 -1175
rect 59150 -1135 59200 -830
rect 59150 -1175 59155 -1135
rect 59195 -1175 59200 -1135
rect 59150 -1180 59200 -1175
rect 59500 -1135 59550 -830
rect 59500 -1175 59505 -1135
rect 59545 -1175 59550 -1135
rect 59500 -1180 59550 -1175
rect 59850 -1135 59900 -830
rect 59850 -1175 59855 -1135
rect 59895 -1175 59900 -1135
rect 59850 -1180 59900 -1175
rect 60200 -1135 60250 -830
rect 60200 -1175 60205 -1135
rect 60245 -1175 60250 -1135
rect 60200 -1180 60250 -1175
rect 60550 -1135 60600 -830
rect 60550 -1175 60555 -1135
rect 60595 -1175 60600 -1135
rect 60550 -1180 60600 -1175
rect 60900 -1130 60950 -830
rect 60900 -1135 61650 -1130
rect 60900 -1175 60905 -1135
rect 60945 -1175 61255 -1135
rect 61295 -1175 61605 -1135
rect 61645 -1175 61650 -1135
rect 60900 -1180 61650 -1175
<< labels >>
flabel metal2 57365 5060 57365 5060 1 FreeSans 240 0 0 80 Vb2_Vb3
flabel metal2 56455 5060 56455 5060 1 FreeSans 240 0 0 80 Vb2_2
flabel metal2 57000 3260 57000 3260 5 FreeSans 200 0 0 -80 Vb3
port 4 s
flabel metal1 56855 3295 56855 3295 5 FreeSans 200 0 0 -80 Vb2
port 5 s
flabel metal2 57950 3820 57950 3820 5 FreeSans 240 0 0 -80 VD3
flabel metal2 55865 3820 55865 3820 5 FreeSans 240 0 0 -80 VD4
flabel metal1 57220 515 57220 515 3 FreeSans 240 0 80 0 V_source
flabel metal2 57720 485 57720 485 5 FreeSans 200 0 0 -80 V_b_2nd_stage
flabel metal2 56800 -235 56800 -235 1 FreeSans 240 0 0 80 Vb1_2
flabel metal2 56460 -90 56460 -90 1 FreeSans 240 0 0 80 V_p_mir
flabel metal1 56945 405 56945 405 7 FreeSans 240 0 -80 0 V_tail_gate
port 11 w
flabel metal2 57770 1030 57770 1030 3 FreeSans 240 0 80 0 VIN-
flabel metal2 56030 1030 56030 1030 7 FreeSans 240 0 -80 0 VIN+
flabel metal1 57430 1075 57430 1075 3 FreeSans 240 0 80 0 VD1
flabel metal1 56370 1075 56370 1075 7 FreeSans 240 0 -80 0 VD2
flabel metal2 56900 1710 56900 1710 5 FreeSans 240 0 0 -80 Vb1
flabel metal3 59895 3185 59895 3185 3 FreeSans 240 0 80 0 cap_res_X
flabel metal1 59860 195 59860 195 5 FreeSans 240 0 0 -80 VOUT-
port 9 s
flabel metal1 59450 1415 59450 1415 1 FreeSans 240 0 0 80 V_CMFB_S1
port 2 n
flabel metal1 59215 1230 59215 1230 1 FreeSans 240 0 0 80 V_CMFB_S2
port 7 n
flabel metal2 57455 2215 57455 2215 7 FreeSans 240 0 -80 0 X
flabel metal2 57525 2415 57525 2415 1 FreeSans 240 0 0 80 err_amp_out
flabel metal2 57000 2460 57000 2460 3 FreeSans 240 0 80 0 err_amp_mir
flabel metal2 57125 2625 57125 2625 3 FreeSans 240 0 80 0 V_err_gate
port 13 e
flabel metal2 56365 2565 56365 2565 7 FreeSans 240 0 -80 0 V_err_amp_ref
port 12 w
flabel metal1 56620 2945 56620 2945 7 FreeSans 240 0 -80 0 V_err_mir_p
flabel metal2 57180 2945 57180 2945 3 FreeSans 240 0 80 0 V_err_p
flabel metal2 57580 2525 57580 2525 1 FreeSans 240 0 0 160 V_tot
flabel metal1 56345 2205 56345 2205 3 FreeSans 240 0 80 0 Y
flabel metal3 54175 3185 54175 3185 7 FreeSans 240 0 -80 0 cap_res_Y
flabel metal2 54210 195 54210 195 5 FreeSans 240 0 0 -80 VOUT+
port 10 s
flabel metal2 54665 1230 54665 1230 1 FreeSans 240 0 0 80 V_CMFB_S4
port 8 n
flabel metal2 54620 1415 54620 1415 1 FreeSans 240 0 0 80 V_CMFB_S3
port 3 n
<< end >>
