magic
tech sky130A
timestamp 1739794596
<< nwell >>
rect 10240 2215 10730 3105
<< nmos >>
rect 10150 1605 10210 2005
rect 10360 1605 10420 2005
rect 10550 1605 10610 2005
<< pmos >>
rect 10360 2285 10420 3085
rect 10550 2285 10610 3085
<< ndiff >>
rect 10100 1990 10150 2005
rect 10100 1970 10115 1990
rect 10135 1970 10150 1990
rect 10100 1940 10150 1970
rect 10100 1920 10115 1940
rect 10135 1920 10150 1940
rect 10100 1890 10150 1920
rect 10100 1870 10115 1890
rect 10135 1870 10150 1890
rect 10100 1840 10150 1870
rect 10100 1820 10115 1840
rect 10135 1820 10150 1840
rect 10100 1790 10150 1820
rect 10100 1770 10115 1790
rect 10135 1770 10150 1790
rect 10100 1740 10150 1770
rect 10100 1720 10115 1740
rect 10135 1720 10150 1740
rect 10100 1690 10150 1720
rect 10100 1670 10115 1690
rect 10135 1670 10150 1690
rect 10100 1640 10150 1670
rect 10100 1620 10115 1640
rect 10135 1620 10150 1640
rect 10100 1605 10150 1620
rect 10210 1990 10260 2005
rect 10310 1990 10360 2005
rect 10210 1970 10225 1990
rect 10245 1970 10260 1990
rect 10310 1970 10325 1990
rect 10345 1970 10360 1990
rect 10210 1940 10260 1970
rect 10310 1940 10360 1970
rect 10210 1920 10225 1940
rect 10245 1920 10260 1940
rect 10310 1920 10325 1940
rect 10345 1920 10360 1940
rect 10210 1890 10260 1920
rect 10310 1890 10360 1920
rect 10210 1870 10225 1890
rect 10245 1870 10260 1890
rect 10310 1870 10325 1890
rect 10345 1870 10360 1890
rect 10210 1840 10260 1870
rect 10310 1840 10360 1870
rect 10210 1820 10225 1840
rect 10245 1820 10260 1840
rect 10310 1820 10325 1840
rect 10345 1820 10360 1840
rect 10210 1790 10260 1820
rect 10310 1790 10360 1820
rect 10210 1770 10225 1790
rect 10245 1770 10260 1790
rect 10310 1770 10325 1790
rect 10345 1770 10360 1790
rect 10210 1740 10260 1770
rect 10310 1740 10360 1770
rect 10210 1720 10225 1740
rect 10245 1720 10260 1740
rect 10310 1720 10325 1740
rect 10345 1720 10360 1740
rect 10210 1690 10260 1720
rect 10310 1690 10360 1720
rect 10210 1670 10225 1690
rect 10245 1670 10260 1690
rect 10310 1670 10325 1690
rect 10345 1670 10360 1690
rect 10210 1640 10260 1670
rect 10310 1640 10360 1670
rect 10210 1620 10225 1640
rect 10245 1620 10260 1640
rect 10310 1620 10325 1640
rect 10345 1620 10360 1640
rect 10210 1605 10260 1620
rect 10310 1605 10360 1620
rect 10420 1990 10470 2005
rect 10420 1970 10435 1990
rect 10455 1970 10470 1990
rect 10420 1940 10470 1970
rect 10420 1920 10435 1940
rect 10455 1920 10470 1940
rect 10420 1890 10470 1920
rect 10420 1870 10435 1890
rect 10455 1870 10470 1890
rect 10420 1840 10470 1870
rect 10420 1820 10435 1840
rect 10455 1820 10470 1840
rect 10420 1790 10470 1820
rect 10420 1770 10435 1790
rect 10455 1770 10470 1790
rect 10420 1740 10470 1770
rect 10420 1720 10435 1740
rect 10455 1720 10470 1740
rect 10420 1690 10470 1720
rect 10420 1670 10435 1690
rect 10455 1670 10470 1690
rect 10420 1640 10470 1670
rect 10420 1620 10435 1640
rect 10455 1620 10470 1640
rect 10420 1605 10470 1620
rect 10500 1990 10550 2005
rect 10500 1970 10515 1990
rect 10535 1970 10550 1990
rect 10500 1940 10550 1970
rect 10500 1920 10515 1940
rect 10535 1920 10550 1940
rect 10500 1890 10550 1920
rect 10500 1870 10515 1890
rect 10535 1870 10550 1890
rect 10500 1840 10550 1870
rect 10500 1820 10515 1840
rect 10535 1820 10550 1840
rect 10500 1790 10550 1820
rect 10500 1770 10515 1790
rect 10535 1770 10550 1790
rect 10500 1740 10550 1770
rect 10500 1720 10515 1740
rect 10535 1720 10550 1740
rect 10500 1690 10550 1720
rect 10500 1670 10515 1690
rect 10535 1670 10550 1690
rect 10500 1640 10550 1670
rect 10500 1620 10515 1640
rect 10535 1620 10550 1640
rect 10500 1605 10550 1620
rect 10610 1990 10660 2005
rect 10610 1970 10625 1990
rect 10645 1970 10660 1990
rect 10610 1940 10660 1970
rect 10610 1920 10625 1940
rect 10645 1920 10660 1940
rect 10610 1890 10660 1920
rect 10610 1870 10625 1890
rect 10645 1870 10660 1890
rect 10610 1840 10660 1870
rect 10610 1820 10625 1840
rect 10645 1820 10660 1840
rect 10610 1790 10660 1820
rect 10610 1770 10625 1790
rect 10645 1770 10660 1790
rect 10610 1740 10660 1770
rect 10610 1720 10625 1740
rect 10645 1720 10660 1740
rect 10610 1690 10660 1720
rect 10610 1670 10625 1690
rect 10645 1670 10660 1690
rect 10610 1640 10660 1670
rect 10610 1620 10625 1640
rect 10645 1620 10660 1640
rect 10610 1605 10660 1620
<< pdiff >>
rect 10310 3070 10360 3085
rect 10310 3050 10325 3070
rect 10345 3050 10360 3070
rect 10310 3020 10360 3050
rect 10310 3000 10325 3020
rect 10345 3000 10360 3020
rect 10310 2970 10360 3000
rect 10310 2950 10325 2970
rect 10345 2950 10360 2970
rect 10310 2920 10360 2950
rect 10310 2900 10325 2920
rect 10345 2900 10360 2920
rect 10310 2870 10360 2900
rect 10310 2850 10325 2870
rect 10345 2850 10360 2870
rect 10310 2820 10360 2850
rect 10310 2800 10325 2820
rect 10345 2800 10360 2820
rect 10310 2770 10360 2800
rect 10310 2750 10325 2770
rect 10345 2750 10360 2770
rect 10310 2720 10360 2750
rect 10310 2700 10325 2720
rect 10345 2700 10360 2720
rect 10310 2670 10360 2700
rect 10310 2650 10325 2670
rect 10345 2650 10360 2670
rect 10310 2620 10360 2650
rect 10310 2600 10325 2620
rect 10345 2600 10360 2620
rect 10310 2570 10360 2600
rect 10310 2550 10325 2570
rect 10345 2550 10360 2570
rect 10310 2520 10360 2550
rect 10310 2500 10325 2520
rect 10345 2500 10360 2520
rect 10310 2470 10360 2500
rect 10310 2450 10325 2470
rect 10345 2450 10360 2470
rect 10310 2420 10360 2450
rect 10310 2400 10325 2420
rect 10345 2400 10360 2420
rect 10310 2370 10360 2400
rect 10310 2350 10325 2370
rect 10345 2350 10360 2370
rect 10310 2320 10360 2350
rect 10310 2300 10325 2320
rect 10345 2300 10360 2320
rect 10310 2285 10360 2300
rect 10420 3070 10465 3085
rect 10420 3050 10435 3070
rect 10455 3050 10465 3070
rect 10420 3020 10465 3050
rect 10420 3000 10435 3020
rect 10455 3000 10465 3020
rect 10420 2970 10465 3000
rect 10420 2950 10435 2970
rect 10455 2950 10465 2970
rect 10420 2920 10465 2950
rect 10420 2900 10435 2920
rect 10455 2900 10465 2920
rect 10420 2870 10465 2900
rect 10420 2850 10435 2870
rect 10455 2850 10465 2870
rect 10420 2820 10465 2850
rect 10420 2800 10435 2820
rect 10455 2800 10465 2820
rect 10420 2770 10465 2800
rect 10420 2750 10435 2770
rect 10455 2750 10465 2770
rect 10420 2720 10465 2750
rect 10420 2700 10435 2720
rect 10455 2700 10465 2720
rect 10420 2670 10465 2700
rect 10420 2650 10435 2670
rect 10455 2650 10465 2670
rect 10420 2620 10465 2650
rect 10420 2600 10435 2620
rect 10455 2600 10465 2620
rect 10420 2570 10465 2600
rect 10420 2550 10435 2570
rect 10455 2550 10465 2570
rect 10420 2520 10465 2550
rect 10420 2500 10435 2520
rect 10455 2500 10465 2520
rect 10420 2470 10465 2500
rect 10420 2450 10435 2470
rect 10455 2450 10465 2470
rect 10420 2420 10465 2450
rect 10420 2400 10435 2420
rect 10455 2400 10465 2420
rect 10420 2370 10465 2400
rect 10420 2350 10435 2370
rect 10455 2350 10465 2370
rect 10420 2320 10465 2350
rect 10420 2300 10435 2320
rect 10455 2300 10465 2320
rect 10420 2285 10465 2300
rect 10500 3070 10550 3085
rect 10500 3050 10515 3070
rect 10535 3050 10550 3070
rect 10500 3020 10550 3050
rect 10500 3000 10515 3020
rect 10535 3000 10550 3020
rect 10500 2970 10550 3000
rect 10500 2950 10515 2970
rect 10535 2950 10550 2970
rect 10500 2920 10550 2950
rect 10500 2900 10515 2920
rect 10535 2900 10550 2920
rect 10500 2870 10550 2900
rect 10500 2850 10515 2870
rect 10535 2850 10550 2870
rect 10500 2820 10550 2850
rect 10500 2800 10515 2820
rect 10535 2800 10550 2820
rect 10500 2770 10550 2800
rect 10500 2750 10515 2770
rect 10535 2750 10550 2770
rect 10500 2720 10550 2750
rect 10500 2700 10515 2720
rect 10535 2700 10550 2720
rect 10500 2670 10550 2700
rect 10500 2650 10515 2670
rect 10535 2650 10550 2670
rect 10500 2620 10550 2650
rect 10500 2600 10515 2620
rect 10535 2600 10550 2620
rect 10500 2570 10550 2600
rect 10500 2550 10515 2570
rect 10535 2550 10550 2570
rect 10500 2520 10550 2550
rect 10500 2500 10515 2520
rect 10535 2500 10550 2520
rect 10500 2470 10550 2500
rect 10500 2450 10515 2470
rect 10535 2450 10550 2470
rect 10500 2420 10550 2450
rect 10500 2400 10515 2420
rect 10535 2400 10550 2420
rect 10500 2370 10550 2400
rect 10500 2350 10515 2370
rect 10535 2350 10550 2370
rect 10500 2320 10550 2350
rect 10500 2300 10515 2320
rect 10535 2300 10550 2320
rect 10500 2285 10550 2300
rect 10610 3070 10660 3085
rect 10610 3050 10625 3070
rect 10645 3050 10660 3070
rect 10610 3020 10660 3050
rect 10610 3000 10625 3020
rect 10645 3000 10660 3020
rect 10610 2970 10660 3000
rect 10610 2950 10625 2970
rect 10645 2950 10660 2970
rect 10610 2920 10660 2950
rect 10610 2900 10625 2920
rect 10645 2900 10660 2920
rect 10610 2870 10660 2900
rect 10610 2850 10625 2870
rect 10645 2850 10660 2870
rect 10610 2820 10660 2850
rect 10610 2800 10625 2820
rect 10645 2800 10660 2820
rect 10610 2770 10660 2800
rect 10610 2750 10625 2770
rect 10645 2750 10660 2770
rect 10610 2720 10660 2750
rect 10610 2700 10625 2720
rect 10645 2700 10660 2720
rect 10610 2670 10660 2700
rect 10610 2650 10625 2670
rect 10645 2650 10660 2670
rect 10610 2620 10660 2650
rect 10610 2600 10625 2620
rect 10645 2600 10660 2620
rect 10610 2570 10660 2600
rect 10610 2550 10625 2570
rect 10645 2550 10660 2570
rect 10610 2520 10660 2550
rect 10610 2500 10625 2520
rect 10645 2500 10660 2520
rect 10610 2470 10660 2500
rect 10610 2450 10625 2470
rect 10645 2450 10660 2470
rect 10610 2420 10660 2450
rect 10610 2400 10625 2420
rect 10645 2400 10660 2420
rect 10610 2370 10660 2400
rect 10610 2350 10625 2370
rect 10645 2350 10660 2370
rect 10610 2320 10660 2350
rect 10610 2300 10625 2320
rect 10645 2300 10660 2320
rect 10610 2285 10660 2300
<< ndiffc >>
rect 10115 1970 10135 1990
rect 10115 1920 10135 1940
rect 10115 1870 10135 1890
rect 10115 1820 10135 1840
rect 10115 1770 10135 1790
rect 10115 1720 10135 1740
rect 10115 1670 10135 1690
rect 10115 1620 10135 1640
rect 10225 1970 10245 1990
rect 10325 1970 10345 1990
rect 10225 1920 10245 1940
rect 10325 1920 10345 1940
rect 10225 1870 10245 1890
rect 10325 1870 10345 1890
rect 10225 1820 10245 1840
rect 10325 1820 10345 1840
rect 10225 1770 10245 1790
rect 10325 1770 10345 1790
rect 10225 1720 10245 1740
rect 10325 1720 10345 1740
rect 10225 1670 10245 1690
rect 10325 1670 10345 1690
rect 10225 1620 10245 1640
rect 10325 1620 10345 1640
rect 10435 1970 10455 1990
rect 10435 1920 10455 1940
rect 10435 1870 10455 1890
rect 10435 1820 10455 1840
rect 10435 1770 10455 1790
rect 10435 1720 10455 1740
rect 10435 1670 10455 1690
rect 10435 1620 10455 1640
rect 10515 1970 10535 1990
rect 10515 1920 10535 1940
rect 10515 1870 10535 1890
rect 10515 1820 10535 1840
rect 10515 1770 10535 1790
rect 10515 1720 10535 1740
rect 10515 1670 10535 1690
rect 10515 1620 10535 1640
rect 10625 1970 10645 1990
rect 10625 1920 10645 1940
rect 10625 1870 10645 1890
rect 10625 1820 10645 1840
rect 10625 1770 10645 1790
rect 10625 1720 10645 1740
rect 10625 1670 10645 1690
rect 10625 1620 10645 1640
<< pdiffc >>
rect 10325 3050 10345 3070
rect 10325 3000 10345 3020
rect 10325 2950 10345 2970
rect 10325 2900 10345 2920
rect 10325 2850 10345 2870
rect 10325 2800 10345 2820
rect 10325 2750 10345 2770
rect 10325 2700 10345 2720
rect 10325 2650 10345 2670
rect 10325 2600 10345 2620
rect 10325 2550 10345 2570
rect 10325 2500 10345 2520
rect 10325 2450 10345 2470
rect 10325 2400 10345 2420
rect 10325 2350 10345 2370
rect 10325 2300 10345 2320
rect 10435 3050 10455 3070
rect 10435 3000 10455 3020
rect 10435 2950 10455 2970
rect 10435 2900 10455 2920
rect 10435 2850 10455 2870
rect 10435 2800 10455 2820
rect 10435 2750 10455 2770
rect 10435 2700 10455 2720
rect 10435 2650 10455 2670
rect 10435 2600 10455 2620
rect 10435 2550 10455 2570
rect 10435 2500 10455 2520
rect 10435 2450 10455 2470
rect 10435 2400 10455 2420
rect 10435 2350 10455 2370
rect 10435 2300 10455 2320
rect 10515 3050 10535 3070
rect 10515 3000 10535 3020
rect 10515 2950 10535 2970
rect 10515 2900 10535 2920
rect 10515 2850 10535 2870
rect 10515 2800 10535 2820
rect 10515 2750 10535 2770
rect 10515 2700 10535 2720
rect 10515 2650 10535 2670
rect 10515 2600 10535 2620
rect 10515 2550 10535 2570
rect 10515 2500 10535 2520
rect 10515 2450 10535 2470
rect 10515 2400 10535 2420
rect 10515 2350 10535 2370
rect 10515 2300 10535 2320
rect 10625 3050 10645 3070
rect 10625 3000 10645 3020
rect 10625 2950 10645 2970
rect 10625 2900 10645 2920
rect 10625 2850 10645 2870
rect 10625 2800 10645 2820
rect 10625 2750 10645 2770
rect 10625 2700 10645 2720
rect 10625 2650 10645 2670
rect 10625 2600 10645 2620
rect 10625 2550 10645 2570
rect 10625 2500 10645 2520
rect 10625 2450 10645 2470
rect 10625 2400 10645 2420
rect 10625 2350 10645 2370
rect 10625 2300 10645 2320
<< psubdiff >>
rect 10260 1990 10310 2005
rect 10260 1970 10275 1990
rect 10295 1970 10310 1990
rect 10260 1940 10310 1970
rect 10260 1920 10275 1940
rect 10295 1920 10310 1940
rect 10260 1890 10310 1920
rect 10260 1870 10275 1890
rect 10295 1870 10310 1890
rect 10260 1840 10310 1870
rect 10260 1820 10275 1840
rect 10295 1820 10310 1840
rect 10260 1790 10310 1820
rect 10260 1770 10275 1790
rect 10295 1770 10310 1790
rect 10260 1740 10310 1770
rect 10260 1720 10275 1740
rect 10295 1720 10310 1740
rect 10260 1690 10310 1720
rect 10260 1670 10275 1690
rect 10295 1670 10310 1690
rect 10260 1640 10310 1670
rect 10260 1620 10275 1640
rect 10295 1620 10310 1640
rect 10260 1605 10310 1620
rect 10660 1990 10710 2005
rect 10660 1970 10675 1990
rect 10695 1970 10710 1990
rect 10660 1940 10710 1970
rect 10660 1920 10675 1940
rect 10695 1920 10710 1940
rect 10660 1890 10710 1920
rect 10660 1870 10675 1890
rect 10695 1870 10710 1890
rect 10660 1840 10710 1870
rect 10660 1820 10675 1840
rect 10695 1820 10710 1840
rect 10660 1790 10710 1820
rect 10660 1770 10675 1790
rect 10695 1770 10710 1790
rect 10660 1740 10710 1770
rect 10660 1720 10675 1740
rect 10695 1720 10710 1740
rect 10660 1690 10710 1720
rect 10660 1670 10675 1690
rect 10695 1670 10710 1690
rect 10660 1640 10710 1670
rect 10660 1620 10675 1640
rect 10695 1620 10710 1640
rect 10660 1605 10710 1620
<< nsubdiff >>
rect 10260 3070 10310 3085
rect 10260 3050 10275 3070
rect 10295 3050 10310 3070
rect 10260 3020 10310 3050
rect 10260 3000 10275 3020
rect 10295 3000 10310 3020
rect 10260 2970 10310 3000
rect 10260 2950 10275 2970
rect 10295 2950 10310 2970
rect 10260 2920 10310 2950
rect 10260 2900 10275 2920
rect 10295 2900 10310 2920
rect 10260 2870 10310 2900
rect 10260 2850 10275 2870
rect 10295 2850 10310 2870
rect 10260 2820 10310 2850
rect 10260 2800 10275 2820
rect 10295 2800 10310 2820
rect 10260 2770 10310 2800
rect 10260 2750 10275 2770
rect 10295 2750 10310 2770
rect 10260 2720 10310 2750
rect 10260 2700 10275 2720
rect 10295 2700 10310 2720
rect 10260 2670 10310 2700
rect 10260 2650 10275 2670
rect 10295 2650 10310 2670
rect 10260 2620 10310 2650
rect 10260 2600 10275 2620
rect 10295 2600 10310 2620
rect 10260 2570 10310 2600
rect 10260 2550 10275 2570
rect 10295 2550 10310 2570
rect 10260 2520 10310 2550
rect 10260 2500 10275 2520
rect 10295 2500 10310 2520
rect 10260 2470 10310 2500
rect 10260 2450 10275 2470
rect 10295 2450 10310 2470
rect 10260 2420 10310 2450
rect 10260 2400 10275 2420
rect 10295 2400 10310 2420
rect 10260 2370 10310 2400
rect 10260 2350 10275 2370
rect 10295 2350 10310 2370
rect 10260 2320 10310 2350
rect 10260 2300 10275 2320
rect 10295 2300 10310 2320
rect 10260 2285 10310 2300
rect 10660 3070 10710 3085
rect 10660 3050 10675 3070
rect 10695 3050 10710 3070
rect 10660 3020 10710 3050
rect 10660 3000 10675 3020
rect 10695 3000 10710 3020
rect 10660 2970 10710 3000
rect 10660 2950 10675 2970
rect 10695 2950 10710 2970
rect 10660 2920 10710 2950
rect 10660 2900 10675 2920
rect 10695 2900 10710 2920
rect 10660 2870 10710 2900
rect 10660 2850 10675 2870
rect 10695 2850 10710 2870
rect 10660 2820 10710 2850
rect 10660 2800 10675 2820
rect 10695 2800 10710 2820
rect 10660 2770 10710 2800
rect 10660 2750 10675 2770
rect 10695 2750 10710 2770
rect 10660 2720 10710 2750
rect 10660 2700 10675 2720
rect 10695 2700 10710 2720
rect 10660 2670 10710 2700
rect 10660 2650 10675 2670
rect 10695 2650 10710 2670
rect 10660 2620 10710 2650
rect 10660 2600 10675 2620
rect 10695 2600 10710 2620
rect 10660 2570 10710 2600
rect 10660 2550 10675 2570
rect 10695 2550 10710 2570
rect 10660 2520 10710 2550
rect 10660 2500 10675 2520
rect 10695 2500 10710 2520
rect 10660 2470 10710 2500
rect 10660 2450 10675 2470
rect 10695 2450 10710 2470
rect 10660 2420 10710 2450
rect 10660 2400 10675 2420
rect 10695 2400 10710 2420
rect 10660 2370 10710 2400
rect 10660 2350 10675 2370
rect 10695 2350 10710 2370
rect 10660 2320 10710 2350
rect 10660 2300 10675 2320
rect 10695 2300 10710 2320
rect 10660 2285 10710 2300
<< psubdiffcont >>
rect 10275 1970 10295 1990
rect 10275 1920 10295 1940
rect 10275 1870 10295 1890
rect 10275 1820 10295 1840
rect 10275 1770 10295 1790
rect 10275 1720 10295 1740
rect 10275 1670 10295 1690
rect 10275 1620 10295 1640
rect 10675 1970 10695 1990
rect 10675 1920 10695 1940
rect 10675 1870 10695 1890
rect 10675 1820 10695 1840
rect 10675 1770 10695 1790
rect 10675 1720 10695 1740
rect 10675 1670 10695 1690
rect 10675 1620 10695 1640
<< nsubdiffcont >>
rect 10275 3050 10295 3070
rect 10275 3000 10295 3020
rect 10275 2950 10295 2970
rect 10275 2900 10295 2920
rect 10275 2850 10295 2870
rect 10275 2800 10295 2820
rect 10275 2750 10295 2770
rect 10275 2700 10295 2720
rect 10275 2650 10295 2670
rect 10275 2600 10295 2620
rect 10275 2550 10295 2570
rect 10275 2500 10295 2520
rect 10275 2450 10295 2470
rect 10275 2400 10295 2420
rect 10275 2350 10295 2370
rect 10275 2300 10295 2320
rect 10675 3050 10695 3070
rect 10675 3000 10695 3020
rect 10675 2950 10695 2970
rect 10675 2900 10695 2920
rect 10675 2850 10695 2870
rect 10675 2800 10695 2820
rect 10675 2750 10695 2770
rect 10675 2700 10695 2720
rect 10675 2650 10695 2670
rect 10675 2600 10695 2620
rect 10675 2550 10695 2570
rect 10675 2500 10695 2520
rect 10675 2450 10695 2470
rect 10675 2400 10695 2420
rect 10675 2350 10695 2370
rect 10675 2300 10695 2320
<< poly >>
rect 10360 3085 10420 3100
rect 10550 3085 10610 3100
rect 10360 2255 10420 2285
rect 10550 2255 10610 2285
rect 10570 2245 10610 2255
rect 10570 2225 10580 2245
rect 10600 2225 10610 2245
rect 10570 2215 10610 2225
rect 10105 2065 10145 2075
rect 10105 2045 10115 2065
rect 10135 2045 10145 2065
rect 10105 2035 10145 2045
rect 10570 2065 10610 2075
rect 10570 2045 10580 2065
rect 10600 2045 10610 2065
rect 10570 2035 10610 2045
rect 10100 2015 10210 2035
rect 10150 2005 10210 2015
rect 10360 2005 10420 2030
rect 10550 2005 10610 2035
rect 10150 1565 10210 1605
rect 10360 1565 10420 1605
rect 10550 1590 10610 1605
rect 10150 1550 10420 1565
<< polycont >>
rect 10580 2225 10600 2245
rect 10115 2045 10135 2065
rect 10580 2045 10600 2065
<< locali >>
rect 10890 3285 10945 3295
rect 10890 3250 10900 3285
rect 10935 3250 10945 3285
rect 10890 3240 10945 3250
rect 10030 3165 10060 3185
rect 10080 3165 10110 3185
rect 10130 3165 10160 3185
rect 10180 3165 10210 3185
rect 10230 3165 10260 3185
rect 10280 3165 10310 3185
rect 10330 3165 10360 3185
rect 10380 3165 10410 3185
rect 10430 3165 10460 3185
rect 10480 3165 10510 3185
rect 10530 3165 10560 3185
rect 10580 3165 10610 3185
rect 10630 3165 10660 3185
rect 10315 3080 10355 3165
rect 10615 3080 10655 3165
rect 10265 3070 10355 3080
rect 10265 3050 10275 3070
rect 10295 3050 10325 3070
rect 10345 3050 10355 3070
rect 10265 3020 10355 3050
rect 10265 3000 10275 3020
rect 10295 3000 10325 3020
rect 10345 3000 10355 3020
rect 10265 2970 10355 3000
rect 10265 2950 10275 2970
rect 10295 2950 10325 2970
rect 10345 2950 10355 2970
rect 10265 2920 10355 2950
rect 10265 2900 10275 2920
rect 10295 2900 10325 2920
rect 10345 2900 10355 2920
rect 10265 2870 10355 2900
rect 10265 2850 10275 2870
rect 10295 2850 10325 2870
rect 10345 2850 10355 2870
rect 10265 2820 10355 2850
rect 10265 2800 10275 2820
rect 10295 2800 10325 2820
rect 10345 2800 10355 2820
rect 10265 2770 10355 2800
rect 10265 2750 10275 2770
rect 10295 2750 10325 2770
rect 10345 2750 10355 2770
rect 10265 2720 10355 2750
rect 10265 2700 10275 2720
rect 10295 2700 10325 2720
rect 10345 2700 10355 2720
rect 10265 2670 10355 2700
rect 10265 2650 10275 2670
rect 10295 2650 10325 2670
rect 10345 2650 10355 2670
rect 10265 2620 10355 2650
rect 10265 2600 10275 2620
rect 10295 2600 10325 2620
rect 10345 2600 10355 2620
rect 10265 2570 10355 2600
rect 10265 2550 10275 2570
rect 10295 2550 10325 2570
rect 10345 2550 10355 2570
rect 10265 2520 10355 2550
rect 10265 2500 10275 2520
rect 10295 2500 10325 2520
rect 10345 2500 10355 2520
rect 10265 2470 10355 2500
rect 10265 2450 10275 2470
rect 10295 2450 10325 2470
rect 10345 2450 10355 2470
rect 10265 2420 10355 2450
rect 10265 2400 10275 2420
rect 10295 2400 10325 2420
rect 10345 2400 10355 2420
rect 10265 2370 10355 2400
rect 10265 2350 10275 2370
rect 10295 2350 10325 2370
rect 10345 2350 10355 2370
rect 10265 2320 10355 2350
rect 10265 2300 10275 2320
rect 10295 2300 10325 2320
rect 10345 2300 10355 2320
rect 10265 2290 10355 2300
rect 10425 3070 10465 3080
rect 10425 3050 10435 3070
rect 10455 3050 10465 3070
rect 10425 3020 10465 3050
rect 10425 3000 10435 3020
rect 10455 3000 10465 3020
rect 10425 2970 10465 3000
rect 10425 2950 10435 2970
rect 10455 2950 10465 2970
rect 10425 2920 10465 2950
rect 10425 2900 10435 2920
rect 10455 2900 10465 2920
rect 10425 2870 10465 2900
rect 10425 2850 10435 2870
rect 10455 2850 10465 2870
rect 10425 2820 10465 2850
rect 10425 2800 10435 2820
rect 10455 2800 10465 2820
rect 10425 2770 10465 2800
rect 10425 2750 10435 2770
rect 10455 2750 10465 2770
rect 10425 2720 10465 2750
rect 10425 2700 10435 2720
rect 10455 2700 10465 2720
rect 10425 2670 10465 2700
rect 10425 2650 10435 2670
rect 10455 2650 10465 2670
rect 10425 2620 10465 2650
rect 10425 2600 10435 2620
rect 10455 2600 10465 2620
rect 10425 2570 10465 2600
rect 10425 2550 10435 2570
rect 10455 2550 10465 2570
rect 10425 2520 10465 2550
rect 10425 2500 10435 2520
rect 10455 2500 10465 2520
rect 10425 2470 10465 2500
rect 10425 2450 10435 2470
rect 10455 2450 10465 2470
rect 10425 2420 10465 2450
rect 10425 2400 10435 2420
rect 10455 2400 10465 2420
rect 10425 2370 10465 2400
rect 10425 2350 10435 2370
rect 10455 2350 10465 2370
rect 10425 2320 10465 2350
rect 10425 2300 10435 2320
rect 10455 2300 10465 2320
rect 9985 2065 10145 2075
rect 9985 2055 10115 2065
rect 10105 2045 10115 2055
rect 10135 2045 10145 2065
rect 10105 1990 10145 2045
rect 10105 1970 10115 1990
rect 10135 1970 10145 1990
rect 10105 1940 10145 1970
rect 10105 1920 10115 1940
rect 10135 1920 10145 1940
rect 10105 1890 10145 1920
rect 10105 1870 10115 1890
rect 10135 1870 10145 1890
rect 10105 1840 10145 1870
rect 10105 1820 10115 1840
rect 10135 1820 10145 1840
rect 10105 1790 10145 1820
rect 10105 1770 10115 1790
rect 10135 1770 10145 1790
rect 10105 1740 10145 1770
rect 10105 1720 10115 1740
rect 10135 1720 10145 1740
rect 10105 1690 10145 1720
rect 10105 1670 10115 1690
rect 10135 1670 10145 1690
rect 10105 1640 10145 1670
rect 10105 1620 10115 1640
rect 10135 1620 10145 1640
rect 10105 1610 10145 1620
rect 10215 1990 10355 2000
rect 10215 1970 10225 1990
rect 10245 1970 10275 1990
rect 10295 1970 10325 1990
rect 10345 1970 10355 1990
rect 10215 1940 10355 1970
rect 10215 1920 10225 1940
rect 10245 1920 10275 1940
rect 10295 1920 10325 1940
rect 10345 1920 10355 1940
rect 10215 1890 10355 1920
rect 10215 1870 10225 1890
rect 10245 1870 10275 1890
rect 10295 1870 10325 1890
rect 10345 1870 10355 1890
rect 10215 1840 10355 1870
rect 10215 1820 10225 1840
rect 10245 1820 10275 1840
rect 10295 1820 10325 1840
rect 10345 1820 10355 1840
rect 10215 1790 10355 1820
rect 10215 1770 10225 1790
rect 10245 1770 10275 1790
rect 10295 1770 10325 1790
rect 10345 1770 10355 1790
rect 10215 1740 10355 1770
rect 10215 1720 10225 1740
rect 10245 1720 10275 1740
rect 10295 1720 10325 1740
rect 10345 1720 10355 1740
rect 10215 1690 10355 1720
rect 10215 1670 10225 1690
rect 10245 1670 10275 1690
rect 10295 1670 10325 1690
rect 10345 1670 10355 1690
rect 10215 1640 10355 1670
rect 10215 1620 10225 1640
rect 10245 1620 10275 1640
rect 10295 1620 10325 1640
rect 10345 1620 10355 1640
rect 10215 1610 10355 1620
rect 10425 1990 10465 2300
rect 10425 1970 10435 1990
rect 10455 1970 10465 1990
rect 10425 1940 10465 1970
rect 10425 1920 10435 1940
rect 10455 1920 10465 1940
rect 10425 1890 10465 1920
rect 10425 1870 10435 1890
rect 10455 1870 10465 1890
rect 10425 1840 10465 1870
rect 10425 1820 10435 1840
rect 10455 1820 10465 1840
rect 10425 1790 10465 1820
rect 10425 1770 10435 1790
rect 10455 1770 10465 1790
rect 10425 1740 10465 1770
rect 10425 1720 10435 1740
rect 10455 1720 10465 1740
rect 10425 1690 10465 1720
rect 10425 1670 10435 1690
rect 10455 1670 10465 1690
rect 10425 1640 10465 1670
rect 10425 1620 10435 1640
rect 10455 1620 10465 1640
rect 10425 1610 10465 1620
rect 10505 3070 10545 3080
rect 10505 3050 10515 3070
rect 10535 3050 10545 3070
rect 10505 3020 10545 3050
rect 10505 3000 10515 3020
rect 10535 3000 10545 3020
rect 10505 2970 10545 3000
rect 10505 2950 10515 2970
rect 10535 2950 10545 2970
rect 10505 2920 10545 2950
rect 10505 2900 10515 2920
rect 10535 2900 10545 2920
rect 10505 2870 10545 2900
rect 10505 2850 10515 2870
rect 10535 2850 10545 2870
rect 10505 2820 10545 2850
rect 10505 2800 10515 2820
rect 10535 2800 10545 2820
rect 10505 2770 10545 2800
rect 10505 2750 10515 2770
rect 10535 2750 10545 2770
rect 10505 2720 10545 2750
rect 10505 2700 10515 2720
rect 10535 2700 10545 2720
rect 10505 2670 10545 2700
rect 10505 2650 10515 2670
rect 10535 2650 10545 2670
rect 10505 2620 10545 2650
rect 10505 2600 10515 2620
rect 10535 2600 10545 2620
rect 10505 2570 10545 2600
rect 10505 2550 10515 2570
rect 10535 2550 10545 2570
rect 10505 2520 10545 2550
rect 10505 2500 10515 2520
rect 10535 2500 10545 2520
rect 10505 2470 10545 2500
rect 10505 2450 10515 2470
rect 10535 2450 10545 2470
rect 10505 2420 10545 2450
rect 10505 2400 10515 2420
rect 10535 2400 10545 2420
rect 10505 2370 10545 2400
rect 10505 2350 10515 2370
rect 10535 2350 10545 2370
rect 10505 2320 10545 2350
rect 10505 2300 10515 2320
rect 10535 2300 10545 2320
rect 10505 2170 10545 2300
rect 10615 3070 10705 3080
rect 10615 3050 10625 3070
rect 10645 3050 10675 3070
rect 10695 3050 10705 3070
rect 10615 3020 10705 3050
rect 10615 3000 10625 3020
rect 10645 3000 10675 3020
rect 10695 3000 10705 3020
rect 10615 2970 10705 3000
rect 10615 2950 10625 2970
rect 10645 2950 10675 2970
rect 10695 2950 10705 2970
rect 10615 2920 10705 2950
rect 10615 2900 10625 2920
rect 10645 2900 10675 2920
rect 10695 2900 10705 2920
rect 10615 2870 10705 2900
rect 10615 2850 10625 2870
rect 10645 2850 10675 2870
rect 10695 2850 10705 2870
rect 10615 2820 10705 2850
rect 10615 2800 10625 2820
rect 10645 2800 10675 2820
rect 10695 2800 10705 2820
rect 10615 2770 10705 2800
rect 10615 2750 10625 2770
rect 10645 2750 10675 2770
rect 10695 2750 10705 2770
rect 10615 2720 10705 2750
rect 10615 2700 10625 2720
rect 10645 2700 10675 2720
rect 10695 2700 10705 2720
rect 10615 2670 10705 2700
rect 10615 2650 10625 2670
rect 10645 2650 10675 2670
rect 10695 2650 10705 2670
rect 10615 2620 10705 2650
rect 10615 2600 10625 2620
rect 10645 2600 10675 2620
rect 10695 2600 10705 2620
rect 10615 2570 10705 2600
rect 10615 2550 10625 2570
rect 10645 2550 10675 2570
rect 10695 2550 10705 2570
rect 10615 2520 10705 2550
rect 10615 2500 10625 2520
rect 10645 2500 10675 2520
rect 10695 2500 10705 2520
rect 10615 2470 10705 2500
rect 10615 2450 10625 2470
rect 10645 2450 10675 2470
rect 10695 2450 10705 2470
rect 10615 2420 10705 2450
rect 10615 2400 10625 2420
rect 10645 2400 10675 2420
rect 10695 2400 10705 2420
rect 10615 2370 10705 2400
rect 10615 2350 10625 2370
rect 10645 2350 10675 2370
rect 10695 2350 10705 2370
rect 10615 2320 10705 2350
rect 10615 2300 10625 2320
rect 10645 2300 10675 2320
rect 10695 2300 10705 2320
rect 10615 2290 10705 2300
rect 10905 2260 10960 2270
rect 10905 2255 10915 2260
rect 10570 2245 10915 2255
rect 10570 2225 10580 2245
rect 10600 2225 10915 2245
rect 10950 2225 10960 2260
rect 10570 2215 10960 2225
rect 10505 2130 10860 2170
rect 10505 1990 10545 2130
rect 10570 2065 10960 2075
rect 10570 2045 10580 2065
rect 10600 2045 10915 2065
rect 10570 2035 10915 2045
rect 10905 2030 10915 2035
rect 10950 2030 10960 2065
rect 10905 2020 10960 2030
rect 10505 1970 10515 1990
rect 10535 1970 10545 1990
rect 10505 1940 10545 1970
rect 10505 1920 10515 1940
rect 10535 1920 10545 1940
rect 10505 1890 10545 1920
rect 10505 1870 10515 1890
rect 10535 1870 10545 1890
rect 10505 1840 10545 1870
rect 10505 1820 10515 1840
rect 10535 1820 10545 1840
rect 10505 1790 10545 1820
rect 10505 1770 10515 1790
rect 10535 1770 10545 1790
rect 10505 1740 10545 1770
rect 10505 1720 10515 1740
rect 10535 1720 10545 1740
rect 10505 1690 10545 1720
rect 10505 1670 10515 1690
rect 10535 1670 10545 1690
rect 10505 1640 10545 1670
rect 10505 1620 10515 1640
rect 10535 1620 10545 1640
rect 10505 1610 10545 1620
rect 10615 1990 10705 2000
rect 10615 1970 10625 1990
rect 10645 1970 10675 1990
rect 10695 1970 10705 1990
rect 10615 1940 10705 1970
rect 10615 1920 10625 1940
rect 10645 1920 10675 1940
rect 10695 1920 10705 1940
rect 10615 1890 10705 1920
rect 10615 1870 10625 1890
rect 10645 1870 10675 1890
rect 10695 1870 10705 1890
rect 10615 1840 10705 1870
rect 10615 1820 10625 1840
rect 10645 1820 10675 1840
rect 10695 1820 10705 1840
rect 10615 1790 10705 1820
rect 10615 1770 10625 1790
rect 10645 1770 10675 1790
rect 10695 1770 10705 1790
rect 10615 1740 10705 1770
rect 10615 1720 10625 1740
rect 10645 1720 10675 1740
rect 10695 1720 10705 1740
rect 10615 1690 10705 1720
rect 10615 1670 10625 1690
rect 10645 1670 10675 1690
rect 10695 1670 10705 1690
rect 10615 1640 10705 1670
rect 10615 1620 10625 1640
rect 10645 1620 10675 1640
rect 10695 1620 10705 1640
rect 10615 1610 10705 1620
rect 10265 1535 10305 1610
rect 10615 1535 10655 1610
rect 10045 1515 10075 1535
rect 10095 1515 10125 1535
rect 10145 1515 10175 1535
rect 10195 1515 10225 1535
rect 10245 1515 10275 1535
rect 10295 1515 10325 1535
rect 10345 1515 10375 1535
rect 10395 1515 10425 1535
rect 10445 1515 10475 1535
rect 10495 1515 10525 1535
rect 10545 1515 10575 1535
rect 10595 1515 10625 1535
rect 10645 1515 10660 1535
rect 10890 1400 10945 1410
rect 10890 1365 10900 1400
rect 10935 1365 10945 1400
rect 10890 1355 10945 1365
<< viali >>
rect 10900 3250 10935 3285
rect 10060 3165 10080 3185
rect 10110 3165 10130 3185
rect 10160 3165 10180 3185
rect 10210 3165 10230 3185
rect 10260 3165 10280 3185
rect 10310 3165 10330 3185
rect 10360 3165 10380 3185
rect 10410 3165 10430 3185
rect 10460 3165 10480 3185
rect 10510 3165 10530 3185
rect 10560 3165 10580 3185
rect 10610 3165 10630 3185
rect 10915 2225 10950 2260
rect 10915 2030 10950 2065
rect 10075 1515 10095 1535
rect 10125 1515 10145 1535
rect 10175 1515 10195 1535
rect 10225 1515 10245 1535
rect 10275 1515 10295 1535
rect 10325 1515 10345 1535
rect 10375 1515 10395 1535
rect 10425 1515 10445 1535
rect 10475 1515 10495 1535
rect 10525 1515 10545 1535
rect 10575 1515 10595 1535
rect 10625 1515 10645 1535
rect 10900 1365 10935 1400
<< metal1 >>
rect 9985 3285 10945 3295
rect 9985 3250 10900 3285
rect 10935 3250 10945 3285
rect 9985 3240 10945 3250
rect 10030 3185 10660 3195
rect 10030 3165 10060 3185
rect 10080 3165 10110 3185
rect 10130 3165 10160 3185
rect 10180 3165 10210 3185
rect 10230 3165 10260 3185
rect 10280 3165 10310 3185
rect 10330 3165 10360 3185
rect 10380 3165 10410 3185
rect 10430 3165 10460 3185
rect 10480 3165 10510 3185
rect 10530 3165 10560 3185
rect 10580 3165 10610 3185
rect 10630 3165 10660 3185
rect 10030 3155 10660 3165
rect 10905 2260 10960 2270
rect 10905 2225 10915 2260
rect 10950 2225 10960 2260
rect 10905 2215 10960 2225
rect 10905 2065 10960 2075
rect 10905 2030 10915 2065
rect 10950 2030 10960 2065
rect 10905 2020 10960 2030
rect 10045 1535 10660 1545
rect 10045 1515 10075 1535
rect 10095 1515 10125 1535
rect 10145 1515 10175 1535
rect 10195 1515 10225 1535
rect 10245 1515 10275 1535
rect 10295 1515 10325 1535
rect 10345 1515 10375 1535
rect 10395 1515 10425 1535
rect 10445 1515 10475 1535
rect 10495 1515 10525 1535
rect 10545 1515 10575 1535
rect 10595 1515 10625 1535
rect 10645 1515 10660 1535
rect 10045 1505 10660 1515
rect 9995 1400 10945 1410
rect 9995 1365 10900 1400
rect 10935 1365 10945 1400
rect 9995 1355 10945 1365
<< via1 >>
rect 10900 3250 10935 3285
rect 10915 2225 10950 2260
rect 10915 2030 10950 2065
rect 10900 1365 10935 1400
<< metal2 >>
rect 10890 3285 10945 3295
rect 10890 3250 10900 3285
rect 10935 3250 10945 3285
rect 10890 3240 10945 3250
rect 10905 2260 10960 2270
rect 10905 2225 10915 2260
rect 10950 2225 10960 2260
rect 10905 2215 10960 2225
rect 10905 2065 10960 2075
rect 10905 2030 10915 2065
rect 10950 2030 10960 2065
rect 10905 2020 10960 2030
rect 10890 1400 10945 1410
rect 10890 1365 10900 1400
rect 10935 1365 10945 1400
rect 10890 1355 10945 1365
<< via2 >>
rect 10900 3250 10935 3285
rect 10915 2225 10950 2260
rect 10915 2030 10950 2065
rect 10900 1365 10935 1400
<< metal3 >>
rect 10890 3285 10945 3295
rect 10890 3250 10900 3285
rect 10935 3250 10945 3285
rect 10890 3050 10945 3250
rect 10890 2390 11795 3050
rect 10905 2260 10960 2270
rect 10905 2225 10915 2260
rect 10950 2225 10960 2260
rect 10905 2215 10960 2225
rect 10905 2065 10960 2075
rect 10905 2030 10915 2065
rect 10950 2030 10960 2065
rect 10905 2020 10960 2030
rect 10890 1610 11230 1900
rect 10890 1400 10945 1610
rect 10890 1365 10900 1400
rect 10935 1365 10945 1400
rect 10890 1355 10945 1365
<< via3 >>
rect 10915 2225 10950 2260
rect 10915 2030 10950 2065
<< mimcap >>
rect 10905 2450 11780 3035
rect 10905 2415 10915 2450
rect 10950 2415 11780 2450
rect 10905 2405 11780 2415
rect 10905 1875 11215 1885
rect 10905 1840 10915 1875
rect 10950 1840 11215 1875
rect 10905 1625 11215 1840
<< mimcapcontact >>
rect 10915 2415 10950 2450
rect 10915 1840 10950 1875
<< metal4 >>
rect 10905 2450 10960 2460
rect 10905 2415 10915 2450
rect 10950 2415 10960 2450
rect 10905 2260 10960 2415
rect 10905 2225 10915 2260
rect 10950 2225 10960 2260
rect 10905 2215 10960 2225
rect 10905 2065 10960 2075
rect 10905 2030 10915 2065
rect 10950 2030 10960 2065
rect 10905 1875 10960 2030
rect 10905 1840 10915 1875
rect 10950 1840 10960 1875
rect 10905 1830 10960 1840
<< labels >>
flabel locali 10545 2105 10545 2105 3 FreeSans 400 0 160 0 vout
port 4 e
flabel poly 10610 2270 10610 2270 3 FreeSans 400 0 200 0 UP_input
port 8 e
flabel locali 10465 2150 10465 2150 3 FreeSans 400 0 200 0 x
port 3 e
flabel poly 10610 2020 10610 2020 3 FreeSans 400 0 200 0 DOWN_input
port 9 e
flabel poly 10360 2255 10360 2255 7 FreeSans 400 0 -200 0 opamp_out
port 10 w
flabel metal1 9995 1380 9995 1380 7 FreeSans 400 0 -200 0 DOWN
port 6 w
flabel metal1 10045 1525 10045 1525 7 FreeSans 400 0 -200 0 GNDA
port 2 w
flabel metal1 10030 3175 10030 3175 7 FreeSans 400 0 -200 0 VDDA
port 1 w
flabel metal1 9985 3265 9985 3265 7 FreeSans 400 0 -200 0 UP_b
port 5 w
flabel locali 9985 2065 9985 2065 7 FreeSans 400 0 -200 0 I_IN
port 7 w
<< end >>
