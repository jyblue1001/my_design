* PEX produced on Mon Feb 17 06:03:56 PM CET 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from pfd_cp_magic_3.ext - technology: sky130A

.subckt pfd_cp_magic V_OUT VDDA GNDA F_REF F_VCO I_IN
X0 a_6400_6270.t4 a_6400_6270.t3 GNDA.t92 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X1 VDDA.t108 opamp_cell_4_0.n_left.t6 opamp_cell_4_0.n_right.t3 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X2 VDDA.t116 opamp_cell_4_0.n_right.t5 pfd_8_0.opamp_out.t8 VDDA.t115 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X3 GNDA.t138 a_6380_5710.t2 a_6380_5710.t3 GNDA.t137 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X4 a_6500_6300.t4 a_6500_6300.t2 a_6500_6300.t3 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X5 pfd_8_0.DOWN_b.t0 VDDA.t129 pfd_8_0.DOWN_PFD_b.t2 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X6 a_870_1400.t0 pfd_8_0.QA_b.t3 VDDA.t71 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X7 a_6500_6300.t12 a_6400_6270.t9 GNDA.t90 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X8 a_6150_5090.t4 opamp_cell_4_0.p_bias.t9 VDDA.t11 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X9 pfd_8_0.DOWN.t0 pfd_8_0.DOWN_b.t2 VDDA.t122 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X10 V_OUT.t3 pfd_8_0.UP_input.t3 VDDA.t90 VDDA.t89 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X11 opamp_cell_4_0.p_bias.t7 opamp_cell_4_0.p_bias.t6 VDDA.t94 VDDA.t93 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X12 a_6150_5090.t12 V_OUT.t6 a_6380_5710.t5 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X13 VDDA.t69 VDDA.t66 VDDA.t68 VDDA.t67 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X14 a_2350_1400.t1 pfd_8_0.before_Reset.t3 GNDA.t27 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X15 pfd_8_0.DOWN.t1 pfd_8_0.DOWN_b.t3 GNDA.t74 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X16 GNDA.t134 GNDA.t131 GNDA.t133 GNDA.t132 sky130_fd_pr__nfet_01v8 ad=0.625 pd=3.5 as=0 ps=0 w=1.25 l=0.5
X17 a_n30_1400.t1 F_REF.t0 VDDA.t28 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X18 pfd_8_0.opamp_out.t3 a_6670_5090.t5 GNDA.t29 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X19 GNDA.t13 pfd_8_0.QA.t3 pfd_8_0.QA_b.t0 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X20 GNDA.t88 a_6400_6270.t10 a_6500_6300.t11 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X21 pfd_8_0.DOWN_input.t0 pfd_8_0.DOWN_b.t4 I_IN.t0 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X22 pfd_8_0.opamp_out.t7 opamp_cell_4_0.n_right.t6 VDDA.t114 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X23 a_1910_2020.t0 pfd_8_0.QB.t3 GNDA.t61 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X24 a_6500_6300.t1 a_6500_6300.t0 a_6500_6300.t1 GNDA.t143 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X25 pfd_8_0.UP.t0 pfd_8_0.UP_PFD_b.t2 VDDA.t100 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X26 pfd_8_0.UP_input.t2 pfd_8_0.UP.t2 pfd_8_0.opamp_out.t9 GNDA.t152 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X27 pfd_8_0.QA.t1 pfd_8_0.QA_b.t4 GNDA.t69 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X28 pfd_8_0.opamp_out.t10 a_9540_3974.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X29 pfd_8_0.DOWN_input.t2 pfd_8_0.DOWN.t3 I_IN.t1 GNDA.t70 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X30 a_1390_1400.t1 pfd_8_0.E.t3 pfd_8_0.E_b.t1 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X31 a_870_640.t1 pfd_8_0.QB_b.t3 VDDA.t128 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X32 VDDA.t65 VDDA.t63 VDDA.t65 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X33 VDDA.t15 a_2530_190.t2 a_2200_190.t0 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X34 GNDA.t130 GNDA.t127 GNDA.t129 GNDA.t128 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X35 pfd_8_0.DOWN_input.t1 pfd_8_0.DOWN_b.t5 GNDA.t39 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X36 GNDA.t48 a_2530_190.t3 a_2200_190.t1 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X37 pfd_8_0.F.t1 pfd_8_0.QB_b.t4 GNDA.t54 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X38 pfd_8_0.UP_b.t2 pfd_8_0.UP.t3 GNDA.t52 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X39 GNDA.t46 pfd_8_0.E_b.t3 pfd_8_0.E.t0 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X40 a_1390_640.t0 pfd_8_0.F.t3 pfd_8_0.F_b.t0 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X41 VDDA.t62 VDDA.t59 VDDA.t61 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X42 a_2350_1400.t0 pfd_8_0.before_Reset.t4 VDDA.t22 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X43 pfd_8_0.F_b.t1 pfd_8_0.F.t4 GNDA.t56 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X44 VDDA.t35 pfd_8_0.F.t5 a_490_640.t0 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X45 pfd_8_0.QA_b.t1 pfd_8_0.QA.t4 a_n30_1400.t0 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X46 GNDA.t126 GNDA.t124 GNDA.t126 GNDA.t125 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X47 opamp_cell_4_0.n_right.t1 opamp_cell_4_0.VIN+.t6 a_6500_6300.t6 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X48 VDDA.t58 VDDA.t56 VDDA.t58 VDDA.t57 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X49 GNDA.t151 pfd_8_0.F.t6 pfd_8_0.QB.t2 GNDA.t150 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X50 pfd_8_0.before_Reset.t0 pfd_8_0.QB.t4 VDDA.t4 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.805 ps=5 w=2 l=0.15
X51 GNDA.t123 GNDA.t121 GNDA.t123 GNDA.t122 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0 ps=0 w=1.25 l=0.5
X52 a_6150_5090.t10 a_6150_5090.t9 a_6150_5090.t10 VDDA.t78 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X53 opamp_cell_4_0.n_right.t4 opamp_cell_4_0.n_left.t7 VDDA.t106 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X54 pfd_8_0.UP_input.t0 pfd_8_0.UP_b.t3 pfd_8_0.opamp_out.t2 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X55 a_490_1400.t1 pfd_8_0.QA_b.t5 pfd_8_0.QA.t0 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X56 a_6380_5710.t1 a_6380_5710.t0 GNDA.t17 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X57 GNDA.t23 pfd_8_0.Reset.t2 pfd_8_0.E_b.t0 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X58 opamp_cell_4_0.p_bias.t5 opamp_cell_4_0.p_bias.t4 VDDA.t96 VDDA.t95 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X59 opamp_cell_4_0.VIN+.t3 pfd_8_0.opamp_out.t11 VDDA.t80 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X60 a_2530_190.t1 a_2350_1400.t2 GNDA.t32 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X61 VDDA.t55 VDDA.t53 VDDA.t55 VDDA.t54 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X62 a_6150_5090.t3 opamp_cell_4_0.p_bias.t10 VDDA.t121 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X63 a_6380_5710.t4 V_OUT.t7 a_6150_5090.t11 VDDA.t91 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X64 GNDA.t86 a_6400_6270.t1 a_6400_6270.t2 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X65 pfd_8_0.E.t2 pfd_8_0.E_b.t4 a_870_1400.t1 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X66 a_6500_6300.t8 V_OUT.t8 opamp_cell_4_0.n_left.t1 GNDA.t72 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X67 pfd_8_0.UP_b.t1 pfd_8_0.UP.t4 VDDA.t32 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X68 GNDA.t84 a_6400_6270.t7 a_6400_6270.t8 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X69 VDDA.t52 VDDA.t50 VDDA.t51 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0 ps=0 w=2.5 l=0.5
X70 VDDA.t98 a_1870_190.t2 pfd_8_0.Reset.t1 VDDA.t97 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X71 VDDA.t76 pfd_8_0.opamp_out.t12 opamp_cell_4_0.VIN+.t2 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X72 VDDA.t104 opamp_cell_4_0.n_left.t4 opamp_cell_4_0.n_left.t5 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X73 VDDA.t88 pfd_8_0.UP_input.t4 V_OUT.t2 VDDA.t87 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X74 GNDA.t82 a_6400_6270.t11 a_6500_6300.t10 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X75 VDDA.t73 opamp_cell_4_0.p_bias.t11 a_6150_5090.t2 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X76 V_OUT.t5 pfd_8_0.DOWN_input.t3 GNDA.t63 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X77 GNDA.t120 GNDA.t117 GNDA.t119 GNDA.t118 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X78 GNDA.t41 a_1870_190.t3 pfd_8_0.Reset.t0 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X79 pfd_8_0.opamp_out.t0 a_6670_5090.t6 GNDA.t7 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X80 opamp_cell_4_0.n_right.t2 a_9540_3974.t1 GNDA.t57 sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X81 GNDA.t116 GNDA.t114 GNDA.t116 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X82 a_6150_5090.t8 a_6150_5090.t6 a_6150_5090.t7 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X83 a_6500_6300.t9 a_6400_6270.t12 GNDA.t80 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X84 opamp_cell_4_0.VIN+.t1 pfd_8_0.opamp_out.t13 VDDA.t126 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X85 pfd_8_0.before_Reset.t2 pfd_8_0.QA.t5 a_1910_2020.t1 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X86 pfd_8_0.opamp_out.t6 opamp_cell_4_0.n_right.t7 VDDA.t112 VDDA.t111 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X87 GNDA.t113 GNDA.t111 GNDA.t113 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X88 pfd_8_0.UP_PFD_b.t1 pfd_8_0.QA.t6 GNDA.t11 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X89 opamp_cell_4_0.p_bias.t8 a_6400_6270.t0 GNDA.t35 sky130_fd_pr__res_xhigh_po_5p73 l=1
X90 a_6400_6270.t6 a_6400_6270.t5 GNDA.t78 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X91 opamp_cell_4_0.n_left.t0 V_OUT.t9 a_6500_6300.t7 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X92 GNDA.t110 GNDA.t108 GNDA.t110 GNDA.t109 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X93 GNDA.t154 pfd_8_0.E.t4 pfd_8_0.QA.t2 GNDA.t153 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X94 pfd_8_0.F.t0 pfd_8_0.F_b.t3 a_870_640.t0 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X95 VDDA.t7 pfd_8_0.Reset.t3 a_1390_1400.t0 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X96 GNDA.t107 GNDA.t105 GNDA.t107 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X97 GNDA.t104 GNDA.t101 GNDA.t103 GNDA.t102 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X98 pfd_8_0.UP_input.t5 pfd_8_0.UP_b.t0 sky130_fd_pr__cap_mim_m3_1 l=6.3 w=7
X99 a_2530_190.t0 a_2350_1400.t3 VDDA.t119 VDDA.t118 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X100 VDDA.t49 VDDA.t47 VDDA.t49 VDDA.t48 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X101 a_9540_6900.t1 a_6670_5090.t1 GNDA.t24 sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X102 opamp_cell_4_0.n_left.t3 opamp_cell_4_0.n_left.t2 VDDA.t102 VDDA.t101 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X103 GNDA.t100 GNDA.t97 GNDA.t99 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X104 GNDA.t67 pfd_8_0.F_b.t4 pfd_8_0.F.t2 GNDA.t66 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X105 GNDA.t59 pfd_8_0.DOWN_input.t4 V_OUT.t4 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X106 pfd_8_0.QB_b.t0 pfd_8_0.QB.t5 a_n30_640.t0 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X107 VDDA.t30 pfd_8_0.opamp_out.t14 opamp_cell_4_0.VIN+.t0 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X108 VDDA.t46 VDDA.t43 VDDA.t45 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X109 pfd_8_0.opamp_out.t15 a_9540_6900.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X110 VDDA.t74 pfd_8_0.Reset.t4 a_1390_640.t1 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X111 GNDA.t76 I_IN.t6 opamp_cell_4_0.VIN+.t5 GNDA.t75 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X112 pfd_8_0.UP_input.t1 pfd_8_0.UP.t5 VDDA.t124 VDDA.t123 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X113 GNDA.t147 a_6380_5710.t6 a_6670_5090.t3 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X114 GNDA.t5 pfd_8_0.QB.t6 pfd_8_0.QB_b.t1 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X115 GNDA.t1 I_IN.t4 I_IN.t5 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X116 GNDA.t21 pfd_8_0.Reset.t5 pfd_8_0.F_b.t2 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X117 GNDA.t9 a_6670_5090.t7 pfd_8_0.opamp_out.t1 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X118 a_6150_5090.t5 opamp_cell_4_0.VIN+.t7 a_6670_5090.t4 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X119 VDDA.t42 VDDA.t39 VDDA.t41 VDDA.t40 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X120 pfd_8_0.E.t1 pfd_8_0.QA_b.t6 GNDA.t37 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X121 VDDA.t110 opamp_cell_4_0.n_right.t8 pfd_8_0.opamp_out.t5 VDDA.t109 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X122 VDDA.t38 VDDA.t36 VDDA.t38 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0 ps=0 w=2.5 l=0.5
X123 VDDA.t13 pfd_8_0.QA.t7 pfd_8_0.before_Reset.t1 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X124 opamp_cell_4_0.VIN+.t4 I_IN.t7 GNDA.t136 GNDA.t135 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X125 a_n30_640.t1 F_VCO.t0 VDDA.t117 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X126 pfd_8_0.UP_PFD_b.t0 pfd_8_0.QA.t8 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X127 VDDA.t127 pfd_8_0.E.t5 a_490_1400.t0 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X128 I_IN.t3 I_IN.t2 GNDA.t140 GNDA.t139 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X129 VDDA.t24 a_2200_190.t2 a_1870_190.t0 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X130 V_OUT.t1 pfd_8_0.UP_input.t6 VDDA.t86 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X131 pfd_8_0.QA_b.t2 F_REF.t1 GNDA.t43 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X132 a_6670_5090.t2 a_6380_5710.t7 GNDA.t145 GNDA.t144 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X133 pfd_8_0.QB_b.t2 F_VCO.t1 GNDA.t65 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X134 a_490_640.t1 pfd_8_0.QB_b.t5 pfd_8_0.QB.t0 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X135 GNDA.t50 a_2200_190.t3 a_1870_190.t1 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X136 VDDA.t9 opamp_cell_4_0.p_bias.t2 opamp_cell_4_0.p_bias.t3 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X137 pfd_8_0.DOWN_input.t5 pfd_8_0.DOWN.t2 sky130_fd_pr__cap_mim_m3_1 l=2.6 w=3.8
X138 pfd_8_0.QB.t1 pfd_8_0.QB_b.t6 GNDA.t149 GNDA.t148 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X139 pfd_8_0.DOWN_PFD_b.t1 pfd_8_0.QB.t7 VDDA.t2 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X140 a_6670_5090.t0 opamp_cell_4_0.VIN+.t8 a_6150_5090.t0 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X141 pfd_8_0.UP.t1 pfd_8_0.UP_PFD_b.t3 GNDA.t15 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X142 VDDA.t82 opamp_cell_4_0.p_bias.t0 opamp_cell_4_0.p_bias.t1 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X143 a_6500_6300.t5 opamp_cell_4_0.VIN+.t9 opamp_cell_4_0.n_right.t0 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X144 GNDA.t34 a_6670_5090.t8 pfd_8_0.opamp_out.t4 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X145 pfd_8_0.DOWN_PFD_b.t0 pfd_8_0.QB.t8 GNDA.t3 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X146 VDDA.t84 pfd_8_0.UP_input.t7 V_OUT.t0 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X147 pfd_8_0.E_b.t2 pfd_8_0.E.t6 GNDA.t142 GNDA.t141 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X148 VDDA.t19 opamp_cell_4_0.p_bias.t12 a_6150_5090.t1 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X149 GNDA.t96 GNDA.t93 GNDA.t95 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X150 pfd_8_0.DOWN_b.t1 GNDA.t155 pfd_8_0.DOWN_PFD_b.t3 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
R0 a_6400_6270.n4 a_6400_6270.t12 317.317
R1 a_6400_6270.n2 a_6400_6270.t11 317.317
R2 a_6400_6270.n5 a_6400_6270.n4 257.067
R3 a_6400_6270.n3 a_6400_6270.n2 257.067
R4 a_6400_6270.n10 a_6400_6270.n9 257.067
R5 a_6400_6270.t0 a_6400_6270.n12 194.478
R6 a_6400_6270.n8 a_6400_6270.n7 152
R7 a_6400_6270.n12 a_6400_6270.n11 152
R8 a_6400_6270.n1 a_6400_6270.n0 120.981
R9 a_6400_6270.n7 a_6400_6270.n6 117.781
R10 a_6400_6270.n7 a_6400_6270.n1 108.8
R11 a_6400_6270.n8 a_6400_6270.n5 85.6894
R12 a_6400_6270.n11 a_6400_6270.n3 85.6894
R13 a_6400_6270.n11 a_6400_6270.n10 85.6894
R14 a_6400_6270.n9 a_6400_6270.n8 85.6894
R15 a_6400_6270.n4 a_6400_6270.t10 60.2505
R16 a_6400_6270.n5 a_6400_6270.t5 60.2505
R17 a_6400_6270.n2 a_6400_6270.t9 60.2505
R18 a_6400_6270.n3 a_6400_6270.t7 60.2505
R19 a_6400_6270.n10 a_6400_6270.t3 60.2505
R20 a_6400_6270.n9 a_6400_6270.t1 60.2505
R21 a_6400_6270.n6 a_6400_6270.t2 24.0005
R22 a_6400_6270.n6 a_6400_6270.t6 24.0005
R23 a_6400_6270.n0 a_6400_6270.t8 24.0005
R24 a_6400_6270.n0 a_6400_6270.t4 24.0005
R25 a_6400_6270.n12 a_6400_6270.n1 3.2005
R26 GNDA.n392 GNDA.n391 19798.9
R27 GNDA.t57 GNDA.n242 6651.75
R28 GNDA.t38 GNDA.n135 5107.62
R29 GNDA.n243 GNDA.t57 3567.2
R30 GNDA.t55 GNDA.t66 2577.14
R31 GNDA.t148 GNDA.t4 2577.14
R32 GNDA.t44 GNDA.t2 2451.43
R33 GNDA.t73 GNDA.t70 1822.86
R34 GNDA.t40 GNDA.n395 1665.71
R35 GNDA.n398 GNDA.n23 1634.29
R36 GNDA.t70 GNDA.n137 1414.29
R37 GNDA.n138 GNDA.t44 1414.29
R38 GNDA.t152 GNDA.n307 1397.16
R39 GNDA.t47 GNDA.n397 1225.71
R40 GNDA.t49 GNDA.n396 1225.71
R41 GNDA.n257 GNDA.n256 1186
R42 GNDA.n58 GNDA.n50 1186
R43 GNDA.n252 GNDA.n251 1186
R44 GNDA.n247 GNDA.n246 1186
R45 GNDA.n137 GNDA.t38 1037.14
R46 GNDA.n138 GNDA.t73 1037.14
R47 GNDA.t2 GNDA.n23 1037.14
R48 GNDA.n398 GNDA.t47 848.572
R49 GNDA.n397 GNDA.t49 848.572
R50 GNDA.n396 GNDA.t40 848.572
R51 GNDA.n395 GNDA.t20 848.572
R52 GNDA.t53 GNDA.n394 848.572
R53 GNDA.n394 GNDA.t150 848.572
R54 GNDA.t64 GNDA.n392 848.572
R55 GNDA.t58 GNDA.t115 733.333
R56 GNDA.t62 GNDA.t58 733.333
R57 GNDA.t102 GNDA.t62 733.333
R58 GNDA.t75 GNDA.t112 733.333
R59 GNDA.t135 GNDA.t75 733.333
R60 GNDA.t98 GNDA.t135 733.333
R61 GNDA.t0 GNDA.t106 733.333
R62 GNDA.t139 GNDA.t0 733.333
R63 GNDA.t94 GNDA.t139 733.333
R64 GNDA.n242 GNDA.t115 700
R65 GNDA.n215 GNDA.t102 700
R66 GNDA.n215 GNDA.t112 700
R67 GNDA.n194 GNDA.t98 700
R68 GNDA.n194 GNDA.t106 700
R69 GNDA.n135 GNDA.t94 700
R70 GNDA.t20 GNDA.t55 691.429
R71 GNDA.t66 GNDA.t53 691.429
R72 GNDA.t150 GNDA.t148 691.429
R73 GNDA.t4 GNDA.t64 691.429
R74 GNDA.n193 GNDA.n192 669.307
R75 GNDA.n196 GNDA.n195 669.307
R76 GNDA.n214 GNDA.n213 669.307
R77 GNDA.n217 GNDA.n216 669.307
R78 GNDA.n241 GNDA.n240 669.307
R79 GNDA.n235 GNDA.n77 669.307
R80 GNDA.n356 GNDA.n355 585.003
R81 GNDA.n394 GNDA.n393 585.003
R82 GNDA.n391 GNDA.n390 585.001
R83 GNDA.n358 GNDA.n357 585.001
R84 GNDA.n353 GNDA.n352 585.001
R85 GNDA.n309 GNDA.n308 585.001
R86 GNDA.n311 GNDA.n310 585.001
R87 GNDA.n137 GNDA.n136 585.001
R88 GNDA.n139 GNDA.n138 585.001
R89 GNDA.n145 GNDA.n23 585.001
R90 GNDA.n399 GNDA.n398 585.001
R91 GNDA.n397 GNDA.n19 585.001
R92 GNDA.n396 GNDA.n16 585.001
R93 GNDA.n395 GNDA.n13 585.001
R94 GNDA.n392 GNDA.n2 585.001
R95 GNDA.n315 GNDA.n314 585.001
R96 GNDA.n313 GNDA.n47 585.001
R97 GNDA.n312 GNDA.n44 585.001
R98 GNDA.n255 GNDA.n254 585.001
R99 GNDA.n307 GNDA.n306 585.001
R100 GNDA.n239 GNDA.n78 585
R101 GNDA.n237 GNDA.n236 585
R102 GNDA.n93 GNDA.n89 585
R103 GNDA.n91 GNDA.n88 585
R104 GNDA.n110 GNDA.n106 585
R105 GNDA.n108 GNDA.n105 585
R106 GNDA.n134 GNDA.n133 585
R107 GNDA.n135 GNDA.n134 585
R108 GNDA.n132 GNDA.n125 585
R109 GNDA.n130 GNDA.n129 585
R110 GNDA.n128 GNDA.n124 585
R111 GNDA.n135 GNDA.n124 585
R112 GNDA.n143 GNDA.t155 566.966
R113 GNDA.n243 GNDA.t24 340.536
R114 GNDA.n107 GNDA.t105 336.329
R115 GNDA.n107 GNDA.t97 336.329
R116 GNDA.n90 GNDA.t111 336.329
R117 GNDA.n90 GNDA.t101 336.329
R118 GNDA.n255 GNDA.t143 333.075
R119 GNDA.n127 GNDA.t93 320.7
R120 GNDA.n234 GNDA.t114 320.7
R121 GNDA.n244 GNDA.t108 304.634
R122 GNDA.n258 GNDA.t127 304.634
R123 GNDA.n59 GNDA.t117 304.634
R124 GNDA.n250 GNDA.t124 304.634
R125 GNDA.t141 GNDA.t45 296.906
R126 GNDA.t68 GNDA.t12 296.906
R127 GNDA.n253 GNDA.t121 292.584
R128 GNDA.n305 GNDA.t131 292.584
R129 GNDA.t91 GNDA.n252 290.373
R130 GNDA.t109 GNDA.n247 281.832
R131 GNDA.n256 GNDA.t128 281.832
R132 GNDA.t30 GNDA.t91 264.752
R133 GNDA.t132 GNDA.n50 256.212
R134 GNDA.n242 GNDA.n241 250.349
R135 GNDA.n242 GNDA.n77 250.349
R136 GNDA.n215 GNDA.n214 250.349
R137 GNDA.n216 GNDA.n215 250.349
R138 GNDA.n194 GNDA.n193 250.349
R139 GNDA.n195 GNDA.n194 250.349
R140 GNDA.n135 GNDA.n123 250.349
R141 GNDA.n246 GNDA.t110 245
R142 GNDA.n257 GNDA.t130 245
R143 GNDA.n58 GNDA.t120 245
R144 GNDA.n251 GNDA.t126 245
R145 GNDA.t85 GNDA.t125 230.59
R146 GNDA.t8 GNDA.t109 222.05
R147 GNDA.t6 GNDA.t8 222.05
R148 GNDA.t33 GNDA.t6 222.05
R149 GNDA.t28 GNDA.t33 222.05
R150 GNDA.t128 GNDA.t28 222.05
R151 GNDA.n256 GNDA.n255 222.05
R152 GNDA.t25 GNDA.t72 222.05
R153 GNDA.t146 GNDA.t144 222.05
R154 GNDA.t16 GNDA.t118 222.05
R155 GNDA.t122 GNDA.t19 213.51
R156 GNDA.t87 GNDA.t137 213.51
R157 GNDA.t51 GNDA.t152 210.007
R158 GNDA.n312 GNDA.t31 206.387
R159 GNDA.n260 GNDA.n74 204.201
R160 GNDA.n61 GNDA.n56 204.201
R161 GNDA.n60 GNDA.n57 204.201
R162 GNDA.n249 GNDA.n248 204.201
R163 GNDA.n259 GNDA.n76 204.201
R164 GNDA.n245 GNDA.n75 204.201
R165 GNDA.n3 GNDA.t5 198.058
R166 GNDA.n440 GNDA.t149 198.058
R167 GNDA.n428 GNDA.t67 198.058
R168 GNDA.n11 GNDA.t56 198.058
R169 GNDA.n384 GNDA.t13 198.058
R170 GNDA.n26 GNDA.t69 198.058
R171 GNDA.n370 GNDA.t46 198.058
R172 GNDA.n365 GNDA.t142 198.058
R173 GNDA.n106 GNDA.n105 197
R174 GNDA.n89 GNDA.n88 197
R175 GNDA.n236 GNDA.n78 197
R176 GNDA.n134 GNDA.n125 197
R177 GNDA.n129 GNDA.n124 197
R178 GNDA.t89 GNDA.t71 196.429
R179 GNDA.n192 GNDA.n104 185
R180 GNDA.n196 GNDA.n104 185
R181 GNDA.n213 GNDA.n87 185
R182 GNDA.n217 GNDA.n87 185
R183 GNDA.n240 GNDA.n79 185
R184 GNDA.n235 GNDA.n79 185
R185 GNDA.n133 GNDA.n126 185
R186 GNDA.n128 GNDA.n126 185
R187 GNDA.n314 GNDA.t14 170.179
R188 GNDA.n313 GNDA.t10 170.179
R189 GNDA.n192 GNDA.n107 166.63
R190 GNDA.n213 GNDA.n90 166.63
R191 GNDA.n247 GNDA.n243 153.727
R192 GNDA.t71 GNDA.t83 145.186
R193 GNDA.n311 GNDA.t26 141.212
R194 GNDA.n309 GNDA.t18 141.212
R195 GNDA.n254 GNDA.t123 134.501
R196 GNDA.n306 GNDA.t134 134.501
R197 GNDA.n7 GNDA.t151 130.713
R198 GNDA.n390 GNDA.t43 130.001
R199 GNDA.n358 GNDA.t23 130.001
R200 GNDA.n352 GNDA.t61 130.001
R201 GNDA.n308 GNDA.t27 130.001
R202 GNDA.n310 GNDA.t32 130.001
R203 GNDA.n2 GNDA.t65 130.001
R204 GNDA.n13 GNDA.t21 130.001
R205 GNDA.n16 GNDA.t41 130.001
R206 GNDA.n19 GNDA.t50 130.001
R207 GNDA.n399 GNDA.t48 130.001
R208 GNDA.n354 GNDA.t37 130.001
R209 GNDA.n28 GNDA.t154 130.001
R210 GNDA.n8 GNDA.t54 130.001
R211 GNDA.t19 GNDA.t81 128.107
R212 GNDA.t137 GNDA.t79 128.107
R213 GNDA.n44 GNDA.t11 122.501
R214 GNDA.n47 GNDA.t15 122.501
R215 GNDA.n315 GNDA.t52 122.501
R216 GNDA.n145 GNDA.t3 122.501
R217 GNDA.n139 GNDA.t74 122.501
R218 GNDA.n136 GNDA.t39 122.501
R219 GNDA.n314 GNDA.t51 112.246
R220 GNDA.t14 GNDA.n313 112.246
R221 GNDA.t10 GNDA.n312 112.246
R222 GNDA.t125 GNDA.t77 111.025
R223 GNDA.t77 GNDA.t146 111.025
R224 GNDA.n357 GNDA.n353 101.382
R225 GNDA.n265 GNDA.n72 97.8707
R226 GNDA.n272 GNDA.n69 97.8707
R227 GNDA.n279 GNDA.n66 97.8707
R228 GNDA.n286 GNDA.n63 97.8707
R229 GNDA.n294 GNDA.n54 97.8707
R230 GNDA.t31 GNDA.n311 97.7622
R231 GNDA.t26 GNDA.n309 97.7622
R232 GNDA.n353 GNDA.t60 97.7622
R233 GNDA.n357 GNDA.t22 97.7622
R234 GNDA.t36 GNDA.n356 97.7622
R235 GNDA.n356 GNDA.t153 97.7622
R236 GNDA.n391 GNDA.t42 97.7622
R237 GNDA.t81 GNDA.t25 93.9446
R238 GNDA.n224 GNDA.n223 92.2612
R239 GNDA.n232 GNDA.n231 92.2612
R240 GNDA.n210 GNDA.n209 92.2612
R241 GNDA.n203 GNDA.n99 92.2612
R242 GNDA.n189 GNDA.n188 92.2612
R243 GNDA.n182 GNDA.n117 92.2612
R244 GNDA.n109 GNDA.n104 91.3721
R245 GNDA.n191 GNDA.n190 91.3721
R246 GNDA.n190 GNDA.n103 91.3721
R247 GNDA.n92 GNDA.n87 91.3721
R248 GNDA.n212 GNDA.n211 91.3721
R249 GNDA.n211 GNDA.n86 91.3721
R250 GNDA.n238 GNDA.n79 90.7567
R251 GNDA.n131 GNDA.n126 90.7567
R252 GNDA.n307 GNDA.n50 85.4042
R253 GNDA.n241 GNDA.n78 84.306
R254 GNDA.n236 GNDA.n77 84.306
R255 GNDA.n214 GNDA.n89 84.306
R256 GNDA.n216 GNDA.n88 84.306
R257 GNDA.n193 GNDA.n106 84.306
R258 GNDA.n195 GNDA.n105 84.306
R259 GNDA.n125 GNDA.n123 84.306
R260 GNDA.n129 GNDA.n123 84.306
R261 GNDA.n249 GNDA.n61 83.2005
R262 GNDA.n61 GNDA.n60 83.2005
R263 GNDA.t18 GNDA.t60 79.6582
R264 GNDA.t22 GNDA.t141 79.6582
R265 GNDA.t45 GNDA.t36 79.6582
R266 GNDA.t153 GNDA.t68 79.6582
R267 GNDA.t12 GNDA.t42 79.6582
R268 GNDA.t83 GNDA.t30 76.8638
R269 GNDA.n260 GNDA.n75 66.5605
R270 GNDA.n260 GNDA.n259 66.5605
R271 GNDA.n261 GNDA.n260 65.9634
R272 GNDA.n390 GNDA.n389 60.29
R273 GNDA.n359 GNDA.n358 60.29
R274 GNDA.n352 GNDA.n351 60.29
R275 GNDA.n308 GNDA.n38 60.29
R276 GNDA.n310 GNDA.n40 60.29
R277 GNDA.n400 GNDA.n399 60.29
R278 GNDA.n407 GNDA.n19 60.29
R279 GNDA.n413 GNDA.n16 60.29
R280 GNDA.n420 GNDA.n13 60.29
R281 GNDA.n448 GNDA.n2 60.29
R282 GNDA.n74 GNDA.t7 60.0005
R283 GNDA.n74 GNDA.t34 60.0005
R284 GNDA.n56 GNDA.t145 60.0005
R285 GNDA.n56 GNDA.t138 60.0005
R286 GNDA.n57 GNDA.t17 60.0005
R287 GNDA.n57 GNDA.t119 60.0005
R288 GNDA.n248 GNDA.t126 60.0005
R289 GNDA.n248 GNDA.t147 60.0005
R290 GNDA.n76 GNDA.t29 60.0005
R291 GNDA.n76 GNDA.t129 60.0005
R292 GNDA.t110 GNDA.n245 60.0005
R293 GNDA.n245 GNDA.t9 60.0005
R294 GNDA.n329 GNDA.n44 59.5478
R295 GNDA.n322 GNDA.n47 59.5478
R296 GNDA.n316 GNDA.n315 59.5478
R297 GNDA.n164 GNDA.n139 58.9809
R298 GNDA.n152 GNDA.n145 58.9809
R299 GNDA.n136 GNDA.n119 58.9809
R300 GNDA.n376 GNDA.n28 54.4005
R301 GNDA.n354 GNDA.n29 54.4005
R302 GNDA.n433 GNDA.n8 54.4005
R303 GNDA.n435 GNDA.n7 54.4005
R304 GNDA.t35 GNDA.t16 52.9508
R305 GNDA.n252 GNDA.t85 51.2427
R306 GNDA.n290 GNDA.n61 41.6005
R307 GNDA.n177 GNDA.n176 41.3005
R308 GNDA.t79 GNDA.t35 40.9943
R309 GNDA.n262 GNDA.n261 39.4985
R310 GNDA.n389 GNDA.n0 33.0991
R311 GNDA.n449 GNDA.n448 33.0991
R312 GNDA.n224 GNDA.n222 32.0005
R313 GNDA.n222 GNDA.n83 32.0005
R314 GNDA.n230 GNDA.n229 32.0005
R315 GNDA.n229 GNDA.n81 32.0005
R316 GNDA.n225 GNDA.n81 32.0005
R317 GNDA.n94 GNDA.n85 32.0005
R318 GNDA.n208 GNDA.n97 32.0005
R319 GNDA.n204 GNDA.n97 32.0005
R320 GNDA.n204 GNDA.n203 32.0005
R321 GNDA.n202 GNDA.n100 32.0005
R322 GNDA.n198 GNDA.n100 32.0005
R323 GNDA.n197 GNDA.n102 32.0005
R324 GNDA.n111 GNDA.n102 32.0005
R325 GNDA.n187 GNDA.n115 32.0005
R326 GNDA.n183 GNDA.n115 32.0005
R327 GNDA.n181 GNDA.n118 32.0005
R328 GNDA.n262 GNDA.n71 32.0005
R329 GNDA.n267 GNDA.n71 32.0005
R330 GNDA.n268 GNDA.n267 32.0005
R331 GNDA.n269 GNDA.n268 32.0005
R332 GNDA.n269 GNDA.n68 32.0005
R333 GNDA.n274 GNDA.n68 32.0005
R334 GNDA.n275 GNDA.n274 32.0005
R335 GNDA.n276 GNDA.n275 32.0005
R336 GNDA.n276 GNDA.n65 32.0005
R337 GNDA.n281 GNDA.n65 32.0005
R338 GNDA.n282 GNDA.n281 32.0005
R339 GNDA.n283 GNDA.n282 32.0005
R340 GNDA.n283 GNDA.n62 32.0005
R341 GNDA.n288 GNDA.n62 32.0005
R342 GNDA.n289 GNDA.n288 32.0005
R343 GNDA.n291 GNDA.n53 32.0005
R344 GNDA.n296 GNDA.n53 32.0005
R345 GNDA.n297 GNDA.n296 32.0005
R346 GNDA.n302 GNDA.n297 32.0005
R347 GNDA.n302 GNDA.n301 32.0005
R348 GNDA.n301 GNDA.n300 32.0005
R349 GNDA.n316 GNDA.n48 32.0005
R350 GNDA.n320 GNDA.n48 32.0005
R351 GNDA.n321 GNDA.n320 32.0005
R352 GNDA.n323 GNDA.n45 32.0005
R353 GNDA.n327 GNDA.n45 32.0005
R354 GNDA.n328 GNDA.n327 32.0005
R355 GNDA.n330 GNDA.n42 32.0005
R356 GNDA.n334 GNDA.n42 32.0005
R357 GNDA.n335 GNDA.n334 32.0005
R358 GNDA.n336 GNDA.n335 32.0005
R359 GNDA.n340 GNDA.n339 32.0005
R360 GNDA.n341 GNDA.n340 32.0005
R361 GNDA.n345 GNDA.n344 32.0005
R362 GNDA.n346 GNDA.n345 32.0005
R363 GNDA.n346 GNDA.n36 32.0005
R364 GNDA.n350 GNDA.n35 32.0005
R365 GNDA.n360 GNDA.n35 32.0005
R366 GNDA.n364 GNDA.n33 32.0005
R367 GNDA.n365 GNDA.n364 32.0005
R368 GNDA.n366 GNDA.n365 32.0005
R369 GNDA.n366 GNDA.n31 32.0005
R370 GNDA.n370 GNDA.n31 32.0005
R371 GNDA.n371 GNDA.n370 32.0005
R372 GNDA.n372 GNDA.n371 32.0005
R373 GNDA.n378 GNDA.n377 32.0005
R374 GNDA.n378 GNDA.n26 32.0005
R375 GNDA.n382 GNDA.n26 32.0005
R376 GNDA.n383 GNDA.n382 32.0005
R377 GNDA.n384 GNDA.n383 32.0005
R378 GNDA.n384 GNDA.n24 32.0005
R379 GNDA.n388 GNDA.n24 32.0005
R380 GNDA.n172 GNDA.n171 32.0005
R381 GNDA.n171 GNDA.n170 32.0005
R382 GNDA.n170 GNDA.n121 32.0005
R383 GNDA.n166 GNDA.n121 32.0005
R384 GNDA.n166 GNDA.n165 32.0005
R385 GNDA.n165 GNDA.n164 32.0005
R386 GNDA.n164 GNDA.n140 32.0005
R387 GNDA.n160 GNDA.n140 32.0005
R388 GNDA.n160 GNDA.n159 32.0005
R389 GNDA.n159 GNDA.n158 32.0005
R390 GNDA.n158 GNDA.n142 32.0005
R391 GNDA.n154 GNDA.n142 32.0005
R392 GNDA.n154 GNDA.n153 32.0005
R393 GNDA.n151 GNDA.n146 32.0005
R394 GNDA.n147 GNDA.n146 32.0005
R395 GNDA.n147 GNDA.n22 32.0005
R396 GNDA.n401 GNDA.n22 32.0005
R397 GNDA.n405 GNDA.n20 32.0005
R398 GNDA.n406 GNDA.n405 32.0005
R399 GNDA.n408 GNDA.n17 32.0005
R400 GNDA.n412 GNDA.n17 32.0005
R401 GNDA.n415 GNDA.n414 32.0005
R402 GNDA.n415 GNDA.n14 32.0005
R403 GNDA.n419 GNDA.n14 32.0005
R404 GNDA.n422 GNDA.n421 32.0005
R405 GNDA.n422 GNDA.n11 32.0005
R406 GNDA.n426 GNDA.n11 32.0005
R407 GNDA.n427 GNDA.n426 32.0005
R408 GNDA.n428 GNDA.n427 32.0005
R409 GNDA.n428 GNDA.n9 32.0005
R410 GNDA.n432 GNDA.n9 32.0005
R411 GNDA.n436 GNDA.n5 32.0005
R412 GNDA.n440 GNDA.n5 32.0005
R413 GNDA.n441 GNDA.n440 32.0005
R414 GNDA.n442 GNDA.n441 32.0005
R415 GNDA.n442 GNDA.n3 32.0005
R416 GNDA.n446 GNDA.n3 32.0005
R417 GNDA.n447 GNDA.n446 32.0005
R418 GNDA.n197 GNDA.n196 29.0291
R419 GNDA.n218 GNDA.n217 29.0291
R420 GNDA.n322 GNDA.n321 28.8005
R421 GNDA.n339 GNDA.n40 28.8005
R422 GNDA.n258 GNDA.n257 27.2005
R423 GNDA.n246 GNDA.n244 27.2005
R424 GNDA.t72 GNDA.t89 25.6216
R425 GNDA.t118 GNDA.t132 25.6216
R426 GNDA.n218 GNDA.n85 25.6005
R427 GNDA.n188 GNDA.n187 25.6005
R428 GNDA.n183 GNDA.n182 25.6005
R429 GNDA.n59 GNDA.n58 25.6005
R430 GNDA.n251 GNDA.n250 25.6005
R431 GNDA.n291 GNDA.n290 25.6005
R432 GNDA.n300 GNDA 25.6005
R433 GNDA.n329 GNDA.n328 25.6005
R434 GNDA.n351 GNDA.n36 25.6005
R435 GNDA.n360 GNDA.n359 25.6005
R436 GNDA.n375 GNDA.n29 25.6005
R437 GNDA.n376 GNDA.n375 25.6005
R438 GNDA.n172 GNDA.n119 25.6005
R439 GNDA.n153 GNDA.n152 25.6005
R440 GNDA.n400 GNDA.n20 25.6005
R441 GNDA.n413 GNDA.n412 25.6005
R442 GNDA.n420 GNDA.n419 25.6005
R443 GNDA.n434 GNDA.n433 25.6005
R444 GNDA.n254 GNDA.n253 24.8279
R445 GNDA.n306 GNDA.n305 24.8279
R446 GNDA.t123 GNDA.n72 24.0005
R447 GNDA.n72 GNDA.t82 24.0005
R448 GNDA.n69 GNDA.t90 24.0005
R449 GNDA.n69 GNDA.t84 24.0005
R450 GNDA.n66 GNDA.t92 24.0005
R451 GNDA.n66 GNDA.t86 24.0005
R452 GNDA.n63 GNDA.t78 24.0005
R453 GNDA.n63 GNDA.t88 24.0005
R454 GNDA.n54 GNDA.t80 24.0005
R455 GNDA.n54 GNDA.t133 24.0005
R456 GNDA.n435 GNDA.n434 22.4005
R457 GNDA.n234 GNDA.n233 20.9665
R458 GNDA.n209 GNDA.n94 19.2005
R459 GNDA.n209 GNDA.n208 19.2005
R460 GNDA.n344 GNDA.n38 19.2005
R461 GNDA.n407 GNDA.n406 16.0005
R462 GNDA.n408 GNDA.n407 16.0005
R463 GNDA.n298 GNDA 15.7005
R464 GNDA.n235 GNDA.n234 15.6449
R465 GNDA.n128 GNDA.n127 15.6449
R466 GNDA.n223 GNDA.t63 15.0005
R467 GNDA.n223 GNDA.t103 15.0005
R468 GNDA.n231 GNDA.t116 15.0005
R469 GNDA.n231 GNDA.t59 15.0005
R470 GNDA.t113 GNDA.n210 15.0005
R471 GNDA.n210 GNDA.t76 15.0005
R472 GNDA.n99 GNDA.t136 15.0005
R473 GNDA.n99 GNDA.t99 15.0005
R474 GNDA.t107 GNDA.n189 15.0005
R475 GNDA.n189 GNDA.t1 15.0005
R476 GNDA.n117 GNDA.t140 15.0005
R477 GNDA.n117 GNDA.t95 15.0005
R478 GNDA.n190 GNDA.t107 15.0005
R479 GNDA.n104 GNDA.t100 15.0005
R480 GNDA.n211 GNDA.t113 15.0005
R481 GNDA.n87 GNDA.t104 15.0005
R482 GNDA.t116 GNDA.n79 15.0005
R483 GNDA.n126 GNDA.t96 15.0005
R484 GNDA.n127 GNDA.n118 14.4005
R485 GNDA.n259 GNDA.n258 14.0805
R486 GNDA.n244 GNDA.n75 14.0805
R487 GNDA.n174 GNDA.n119 13.9181
R488 GNDA.n298 GNDA.n49 13.506
R489 GNDA.n317 GNDA.n49 12.8163
R490 GNDA.n218 GNDA.n83 12.8005
R491 GNDA.n232 GNDA.n230 12.8005
R492 GNDA.n188 GNDA.n111 12.8005
R493 GNDA.n182 GNDA.n181 12.8005
R494 GNDA.n60 GNDA.n59 12.8005
R495 GNDA.n250 GNDA.n249 12.8005
R496 GNDA.n341 GNDA.n38 12.8005
R497 GNDA GNDA.n0 12.7806
R498 GNDA GNDA.n449 11.8829
R499 GNDA.n176 GNDA.n175 11.8187
R500 GNDA.n175 GNDA.n174 11.8152
R501 GNDA.n436 GNDA.n435 9.6005
R502 GNDA.n253 GNDA.n73 9.58175
R503 GNDA.n305 GNDA.n304 9.58175
R504 GNDA.n263 GNDA.n262 9.3005
R505 GNDA.n264 GNDA.n71 9.3005
R506 GNDA.n267 GNDA.n266 9.3005
R507 GNDA.n268 GNDA.n70 9.3005
R508 GNDA.n270 GNDA.n269 9.3005
R509 GNDA.n271 GNDA.n68 9.3005
R510 GNDA.n274 GNDA.n273 9.3005
R511 GNDA.n275 GNDA.n67 9.3005
R512 GNDA.n277 GNDA.n276 9.3005
R513 GNDA.n278 GNDA.n65 9.3005
R514 GNDA.n281 GNDA.n280 9.3005
R515 GNDA.n282 GNDA.n64 9.3005
R516 GNDA.n284 GNDA.n283 9.3005
R517 GNDA.n285 GNDA.n62 9.3005
R518 GNDA.n288 GNDA.n287 9.3005
R519 GNDA.n289 GNDA.n55 9.3005
R520 GNDA.n292 GNDA.n291 9.3005
R521 GNDA.n293 GNDA.n53 9.3005
R522 GNDA.n296 GNDA.n295 9.3005
R523 GNDA.n297 GNDA.n51 9.3005
R524 GNDA.n303 GNDA.n302 9.3005
R525 GNDA.n301 GNDA.n52 9.3005
R526 GNDA.n300 GNDA.n299 9.3005
R527 GNDA.n318 GNDA.n48 9.3005
R528 GNDA.n320 GNDA.n319 9.3005
R529 GNDA.n321 GNDA.n46 9.3005
R530 GNDA.n324 GNDA.n323 9.3005
R531 GNDA.n325 GNDA.n45 9.3005
R532 GNDA.n327 GNDA.n326 9.3005
R533 GNDA.n328 GNDA.n43 9.3005
R534 GNDA.n331 GNDA.n330 9.3005
R535 GNDA.n332 GNDA.n42 9.3005
R536 GNDA.n334 GNDA.n333 9.3005
R537 GNDA.n335 GNDA.n41 9.3005
R538 GNDA.n337 GNDA.n336 9.3005
R539 GNDA.n339 GNDA.n338 9.3005
R540 GNDA.n340 GNDA.n39 9.3005
R541 GNDA.n342 GNDA.n341 9.3005
R542 GNDA.n344 GNDA.n343 9.3005
R543 GNDA.n345 GNDA.n37 9.3005
R544 GNDA.n347 GNDA.n346 9.3005
R545 GNDA.n348 GNDA.n36 9.3005
R546 GNDA.n350 GNDA.n349 9.3005
R547 GNDA.n35 GNDA.n34 9.3005
R548 GNDA.n361 GNDA.n360 9.3005
R549 GNDA.n362 GNDA.n33 9.3005
R550 GNDA.n364 GNDA.n363 9.3005
R551 GNDA.n365 GNDA.n32 9.3005
R552 GNDA.n367 GNDA.n366 9.3005
R553 GNDA.n368 GNDA.n31 9.3005
R554 GNDA.n370 GNDA.n369 9.3005
R555 GNDA.n371 GNDA.n30 9.3005
R556 GNDA.n373 GNDA.n372 9.3005
R557 GNDA.n375 GNDA.n374 9.3005
R558 GNDA.n377 GNDA.n27 9.3005
R559 GNDA.n379 GNDA.n378 9.3005
R560 GNDA.n380 GNDA.n26 9.3005
R561 GNDA.n382 GNDA.n381 9.3005
R562 GNDA.n383 GNDA.n25 9.3005
R563 GNDA.n385 GNDA.n384 9.3005
R564 GNDA.n386 GNDA.n24 9.3005
R565 GNDA.n388 GNDA.n387 9.3005
R566 GNDA.n178 GNDA.n177 9.3005
R567 GNDA.n179 GNDA.n118 9.3005
R568 GNDA.n181 GNDA.n180 9.3005
R569 GNDA.n182 GNDA.n116 9.3005
R570 GNDA.n184 GNDA.n183 9.3005
R571 GNDA.n185 GNDA.n115 9.3005
R572 GNDA.n187 GNDA.n186 9.3005
R573 GNDA.n188 GNDA.n114 9.3005
R574 GNDA.n113 GNDA.n111 9.3005
R575 GNDA.n112 GNDA.n102 9.3005
R576 GNDA.n197 GNDA.n101 9.3005
R577 GNDA.n230 GNDA.n80 9.3005
R578 GNDA.n229 GNDA.n228 9.3005
R579 GNDA.n227 GNDA.n81 9.3005
R580 GNDA.n226 GNDA.n225 9.3005
R581 GNDA.n224 GNDA.n82 9.3005
R582 GNDA.n222 GNDA.n221 9.3005
R583 GNDA.n220 GNDA.n83 9.3005
R584 GNDA.n219 GNDA.n218 9.3005
R585 GNDA.n85 GNDA.n84 9.3005
R586 GNDA.n95 GNDA.n94 9.3005
R587 GNDA.n209 GNDA.n96 9.3005
R588 GNDA.n208 GNDA.n207 9.3005
R589 GNDA.n206 GNDA.n97 9.3005
R590 GNDA.n205 GNDA.n204 9.3005
R591 GNDA.n203 GNDA.n98 9.3005
R592 GNDA.n202 GNDA.n201 9.3005
R593 GNDA.n200 GNDA.n100 9.3005
R594 GNDA.n199 GNDA.n198 9.3005
R595 GNDA.n173 GNDA.n172 9.3005
R596 GNDA.n171 GNDA.n120 9.3005
R597 GNDA.n170 GNDA.n169 9.3005
R598 GNDA.n168 GNDA.n121 9.3005
R599 GNDA.n167 GNDA.n166 9.3005
R600 GNDA.n165 GNDA.n122 9.3005
R601 GNDA.n164 GNDA.n163 9.3005
R602 GNDA.n162 GNDA.n140 9.3005
R603 GNDA.n161 GNDA.n160 9.3005
R604 GNDA.n159 GNDA.n141 9.3005
R605 GNDA.n158 GNDA.n157 9.3005
R606 GNDA.n156 GNDA.n142 9.3005
R607 GNDA.n155 GNDA.n154 9.3005
R608 GNDA.n153 GNDA.n144 9.3005
R609 GNDA.n151 GNDA.n150 9.3005
R610 GNDA.n149 GNDA.n146 9.3005
R611 GNDA.n148 GNDA.n147 9.3005
R612 GNDA.n22 GNDA.n21 9.3005
R613 GNDA.n402 GNDA.n401 9.3005
R614 GNDA.n403 GNDA.n20 9.3005
R615 GNDA.n405 GNDA.n404 9.3005
R616 GNDA.n406 GNDA.n18 9.3005
R617 GNDA.n409 GNDA.n408 9.3005
R618 GNDA.n410 GNDA.n17 9.3005
R619 GNDA.n412 GNDA.n411 9.3005
R620 GNDA.n414 GNDA.n15 9.3005
R621 GNDA.n416 GNDA.n415 9.3005
R622 GNDA.n417 GNDA.n14 9.3005
R623 GNDA.n419 GNDA.n418 9.3005
R624 GNDA.n421 GNDA.n12 9.3005
R625 GNDA.n423 GNDA.n422 9.3005
R626 GNDA.n424 GNDA.n11 9.3005
R627 GNDA.n426 GNDA.n425 9.3005
R628 GNDA.n427 GNDA.n10 9.3005
R629 GNDA.n429 GNDA.n428 9.3005
R630 GNDA.n430 GNDA.n9 9.3005
R631 GNDA.n432 GNDA.n431 9.3005
R632 GNDA.n434 GNDA.n6 9.3005
R633 GNDA.n437 GNDA.n436 9.3005
R634 GNDA.n438 GNDA.n5 9.3005
R635 GNDA.n440 GNDA.n439 9.3005
R636 GNDA.n441 GNDA.n4 9.3005
R637 GNDA.n443 GNDA.n442 9.3005
R638 GNDA.n444 GNDA.n3 9.3005
R639 GNDA.n446 GNDA.n445 9.3005
R640 GNDA.n447 GNDA.n1 9.3005
R641 GNDA.t143 GNDA.t122 8.54087
R642 GNDA.t144 GNDA.t87 8.54087
R643 GNDA.n317 GNDA.n316 7.49888
R644 GNDA.n240 GNDA.n239 7.11161
R645 GNDA.n237 GNDA.n235 7.11161
R646 GNDA.n133 GNDA.n132 7.11161
R647 GNDA.n130 GNDA.n128 7.11161
R648 GNDA.n233 GNDA.n232 6.69883
R649 GNDA.n225 GNDA.n224 6.4005
R650 GNDA.n203 GNDA.n202 6.4005
R651 GNDA.n198 GNDA.n197 6.4005
R652 GNDA.n290 GNDA.n289 6.4005
R653 GNDA.n330 GNDA.n329 6.4005
R654 GNDA.n351 GNDA.n350 6.4005
R655 GNDA.n359 GNDA.n33 6.4005
R656 GNDA.n372 GNDA.n29 6.4005
R657 GNDA.n377 GNDA.n376 6.4005
R658 GNDA.n389 GNDA.n388 6.4005
R659 GNDA.n152 GNDA.n151 6.4005
R660 GNDA.n401 GNDA.n400 6.4005
R661 GNDA.n414 GNDA.n413 6.4005
R662 GNDA.n421 GNDA.n420 6.4005
R663 GNDA.n433 GNDA.n432 6.4005
R664 GNDA.n448 GNDA.n447 6.4005
R665 GNDA.n177 GNDA.n118 6.4005
R666 GNDA.n355 GNDA.n354 5.68939
R667 GNDA.n355 GNDA.n28 5.68939
R668 GNDA.n393 GNDA.n8 5.68939
R669 GNDA.n393 GNDA.n7 4.97828
R670 GNDA.n239 GNDA.n238 3.48951
R671 GNDA.n238 GNDA.n237 3.48951
R672 GNDA.n132 GNDA.n131 3.48951
R673 GNDA.n131 GNDA.n130 3.48951
R674 GNDA.n323 GNDA.n322 3.2005
R675 GNDA.n336 GNDA.n40 3.2005
R676 GNDA.n191 GNDA.n110 2.25882
R677 GNDA.n110 GNDA.n109 2.25882
R678 GNDA.n196 GNDA.n103 2.25882
R679 GNDA.n109 GNDA.n108 2.25882
R680 GNDA.n192 GNDA.n191 2.25882
R681 GNDA.n108 GNDA.n103 2.25882
R682 GNDA.n212 GNDA.n93 2.25882
R683 GNDA.n93 GNDA.n92 2.25882
R684 GNDA.n217 GNDA.n86 2.25882
R685 GNDA.n92 GNDA.n91 2.25882
R686 GNDA.n213 GNDA.n212 2.25882
R687 GNDA.n91 GNDA.n86 2.25882
R688 GNDA.n175 GNDA.n49 1.0063
R689 GNDA.n233 GNDA.n80 0.703977
R690 GNDA.n318 GNDA.n317 0.193977
R691 GNDA.n387 GNDA.n0 0.193881
R692 GNDA.n449 GNDA.n1 0.193881
R693 GNDA.n174 GNDA.n173 0.193695
R694 GNDA.n299 GNDA.n298 0.188
R695 GNDA.n264 GNDA.n263 0.15675
R696 GNDA.n266 GNDA.n70 0.15675
R697 GNDA.n270 GNDA.n70 0.15675
R698 GNDA.n271 GNDA.n270 0.15675
R699 GNDA.n273 GNDA.n67 0.15675
R700 GNDA.n277 GNDA.n67 0.15675
R701 GNDA.n278 GNDA.n277 0.15675
R702 GNDA.n280 GNDA.n64 0.15675
R703 GNDA.n284 GNDA.n64 0.15675
R704 GNDA.n285 GNDA.n284 0.15675
R705 GNDA.n287 GNDA.n55 0.15675
R706 GNDA.n292 GNDA.n55 0.15675
R707 GNDA.n293 GNDA.n292 0.15675
R708 GNDA.n295 GNDA.n51 0.15675
R709 GNDA.n303 GNDA.n52 0.15675
R710 GNDA.n299 GNDA.n52 0.15675
R711 GNDA.n319 GNDA.n318 0.15675
R712 GNDA.n319 GNDA.n46 0.15675
R713 GNDA.n324 GNDA.n46 0.15675
R714 GNDA.n325 GNDA.n324 0.15675
R715 GNDA.n326 GNDA.n325 0.15675
R716 GNDA.n326 GNDA.n43 0.15675
R717 GNDA.n331 GNDA.n43 0.15675
R718 GNDA.n332 GNDA.n331 0.15675
R719 GNDA.n333 GNDA.n332 0.15675
R720 GNDA.n333 GNDA.n41 0.15675
R721 GNDA.n337 GNDA.n41 0.15675
R722 GNDA.n338 GNDA.n337 0.15675
R723 GNDA.n338 GNDA.n39 0.15675
R724 GNDA.n342 GNDA.n39 0.15675
R725 GNDA.n343 GNDA.n342 0.15675
R726 GNDA.n343 GNDA.n37 0.15675
R727 GNDA.n347 GNDA.n37 0.15675
R728 GNDA.n348 GNDA.n347 0.15675
R729 GNDA.n349 GNDA.n348 0.15675
R730 GNDA.n349 GNDA.n34 0.15675
R731 GNDA.n361 GNDA.n34 0.15675
R732 GNDA.n362 GNDA.n361 0.15675
R733 GNDA.n363 GNDA.n362 0.15675
R734 GNDA.n363 GNDA.n32 0.15675
R735 GNDA.n367 GNDA.n32 0.15675
R736 GNDA.n368 GNDA.n367 0.15675
R737 GNDA.n369 GNDA.n368 0.15675
R738 GNDA.n369 GNDA.n30 0.15675
R739 GNDA.n373 GNDA.n30 0.15675
R740 GNDA.n374 GNDA.n373 0.15675
R741 GNDA.n374 GNDA.n27 0.15675
R742 GNDA.n379 GNDA.n27 0.15675
R743 GNDA.n380 GNDA.n379 0.15675
R744 GNDA.n381 GNDA.n380 0.15675
R745 GNDA.n381 GNDA.n25 0.15675
R746 GNDA.n385 GNDA.n25 0.15675
R747 GNDA.n386 GNDA.n385 0.15675
R748 GNDA.n387 GNDA.n386 0.15675
R749 GNDA.n228 GNDA.n80 0.15675
R750 GNDA.n228 GNDA.n227 0.15675
R751 GNDA.n227 GNDA.n226 0.15675
R752 GNDA.n226 GNDA.n82 0.15675
R753 GNDA.n221 GNDA.n82 0.15675
R754 GNDA.n221 GNDA.n220 0.15675
R755 GNDA.n220 GNDA.n219 0.15675
R756 GNDA.n219 GNDA.n84 0.15675
R757 GNDA.n95 GNDA.n84 0.15675
R758 GNDA.n96 GNDA.n95 0.15675
R759 GNDA.n207 GNDA.n96 0.15675
R760 GNDA.n207 GNDA.n206 0.15675
R761 GNDA.n206 GNDA.n205 0.15675
R762 GNDA.n205 GNDA.n98 0.15675
R763 GNDA.n201 GNDA.n98 0.15675
R764 GNDA.n201 GNDA.n200 0.15675
R765 GNDA.n200 GNDA.n199 0.15675
R766 GNDA.n199 GNDA.n101 0.15675
R767 GNDA.n112 GNDA.n101 0.15675
R768 GNDA.n113 GNDA.n112 0.15675
R769 GNDA.n114 GNDA.n113 0.15675
R770 GNDA.n186 GNDA.n114 0.15675
R771 GNDA.n186 GNDA.n185 0.15675
R772 GNDA.n185 GNDA.n184 0.15675
R773 GNDA.n184 GNDA.n116 0.15675
R774 GNDA.n180 GNDA.n116 0.15675
R775 GNDA.n180 GNDA.n179 0.15675
R776 GNDA.n179 GNDA.n178 0.15675
R777 GNDA.n173 GNDA.n120 0.15675
R778 GNDA.n169 GNDA.n120 0.15675
R779 GNDA.n169 GNDA.n168 0.15675
R780 GNDA.n168 GNDA.n167 0.15675
R781 GNDA.n167 GNDA.n122 0.15675
R782 GNDA.n163 GNDA.n122 0.15675
R783 GNDA.n163 GNDA.n162 0.15675
R784 GNDA.n162 GNDA.n161 0.15675
R785 GNDA.n161 GNDA.n141 0.15675
R786 GNDA.n157 GNDA.n156 0.15675
R787 GNDA.n156 GNDA.n155 0.15675
R788 GNDA.n155 GNDA.n144 0.15675
R789 GNDA.n150 GNDA.n144 0.15675
R790 GNDA.n150 GNDA.n149 0.15675
R791 GNDA.n149 GNDA.n148 0.15675
R792 GNDA.n148 GNDA.n21 0.15675
R793 GNDA.n402 GNDA.n21 0.15675
R794 GNDA.n403 GNDA.n402 0.15675
R795 GNDA.n404 GNDA.n403 0.15675
R796 GNDA.n404 GNDA.n18 0.15675
R797 GNDA.n409 GNDA.n18 0.15675
R798 GNDA.n410 GNDA.n409 0.15675
R799 GNDA.n411 GNDA.n410 0.15675
R800 GNDA.n411 GNDA.n15 0.15675
R801 GNDA.n416 GNDA.n15 0.15675
R802 GNDA.n417 GNDA.n416 0.15675
R803 GNDA.n418 GNDA.n417 0.15675
R804 GNDA.n418 GNDA.n12 0.15675
R805 GNDA.n423 GNDA.n12 0.15675
R806 GNDA.n424 GNDA.n423 0.15675
R807 GNDA.n425 GNDA.n424 0.15675
R808 GNDA.n425 GNDA.n10 0.15675
R809 GNDA.n429 GNDA.n10 0.15675
R810 GNDA.n430 GNDA.n429 0.15675
R811 GNDA.n431 GNDA.n430 0.15675
R812 GNDA.n431 GNDA.n6 0.15675
R813 GNDA.n437 GNDA.n6 0.15675
R814 GNDA.n438 GNDA.n437 0.15675
R815 GNDA.n439 GNDA.n438 0.15675
R816 GNDA.n439 GNDA.n4 0.15675
R817 GNDA.n443 GNDA.n4 0.15675
R818 GNDA.n444 GNDA.n443 0.15675
R819 GNDA.n445 GNDA.n444 0.15675
R820 GNDA.n445 GNDA.n1 0.15675
R821 GNDA.n261 GNDA.n73 0.131895
R822 GNDA.n178 GNDA 0.1255
R823 GNDA.n143 GNDA.n141 0.109875
R824 GNDA.n265 GNDA.n264 0.09425
R825 GNDA.n272 GNDA.n271 0.09425
R826 GNDA.n279 GNDA.n278 0.09425
R827 GNDA.n286 GNDA.n285 0.09425
R828 GNDA.n294 GNDA.n293 0.09425
R829 GNDA.n304 GNDA.n51 0.09425
R830 GNDA.n263 GNDA.n73 0.063
R831 GNDA.n266 GNDA.n265 0.063
R832 GNDA.n273 GNDA.n272 0.063
R833 GNDA.n280 GNDA.n279 0.063
R834 GNDA.n287 GNDA.n286 0.063
R835 GNDA.n295 GNDA.n294 0.063
R836 GNDA.n304 GNDA.n303 0.063
R837 GNDA.n176 GNDA 0.063
R838 GNDA.n157 GNDA.n143 0.047375
R839 opamp_cell_4_0.n_left.n1 opamp_cell_4_0.n_left.t6 401.668
R840 opamp_cell_4_0.n_left.n5 opamp_cell_4_0.n_left.n4 325.248
R841 opamp_cell_4_0.n_left.n4 opamp_cell_4_0.n_left.n0 313
R842 opamp_cell_4_0.n_left.n3 opamp_cell_4_0.n_left.t2 252.248
R843 opamp_cell_4_0.n_left.n2 opamp_cell_4_0.n_left.n1 208.868
R844 opamp_cell_4_0.n_left.n2 opamp_cell_4_0.n_left.t4 192.8
R845 opamp_cell_4_0.n_left.n1 opamp_cell_4_0.n_left.t7 192.8
R846 opamp_cell_4_0.n_left.n4 opamp_cell_4_0.n_left.n3 152
R847 opamp_cell_4_0.n_left.n0 opamp_cell_4_0.n_left.t1 60.0005
R848 opamp_cell_4_0.n_left.n0 opamp_cell_4_0.n_left.t0 60.0005
R849 opamp_cell_4_0.n_left.n3 opamp_cell_4_0.n_left.n2 59.4472
R850 opamp_cell_4_0.n_left.n5 opamp_cell_4_0.n_left.t5 49.2505
R851 opamp_cell_4_0.n_left.t3 opamp_cell_4_0.n_left.n5 49.2505
R852 opamp_cell_4_0.n_right.t2 opamp_cell_4_0.n_right.n6 1010.36
R853 opamp_cell_4_0.n_right.n3 opamp_cell_4_0.n_right.n2 416.101
R854 opamp_cell_4_0.n_right.n2 opamp_cell_4_0.n_right.n1 354.048
R855 opamp_cell_4_0.n_right.n3 opamp_cell_4_0.n_right.t6 289.2
R856 opamp_cell_4_0.n_right.n4 opamp_cell_4_0.n_right.t5 289.2
R857 opamp_cell_4_0.n_right.n5 opamp_cell_4_0.n_right.t7 289.2
R858 opamp_cell_4_0.n_right.n6 opamp_cell_4_0.n_right.t8 289.2
R859 opamp_cell_4_0.n_right.n2 opamp_cell_4_0.n_right.n0 284.2
R860 opamp_cell_4_0.n_right.n6 opamp_cell_4_0.n_right.n5 208.868
R861 opamp_cell_4_0.n_right.n5 opamp_cell_4_0.n_right.n4 208.868
R862 opamp_cell_4_0.n_right.n4 opamp_cell_4_0.n_right.n3 208.868
R863 opamp_cell_4_0.n_right.n0 opamp_cell_4_0.n_right.t0 60.0005
R864 opamp_cell_4_0.n_right.n0 opamp_cell_4_0.n_right.t1 60.0005
R865 opamp_cell_4_0.n_right.n1 opamp_cell_4_0.n_right.t3 49.2505
R866 opamp_cell_4_0.n_right.n1 opamp_cell_4_0.n_right.t4 49.2505
R867 VDDA.n164 VDDA.n130 3803.21
R868 VDDA.n261 VDDA.t123 2266.27
R869 VDDA.n441 VDDA.n433 831.25
R870 VDDA.n436 VDDA.n435 831.25
R871 VDDA.n452 VDDA.n444 831.25
R872 VDDA.n447 VDDA.n446 831.25
R873 VDDA.n151 VDDA.n150 585
R874 VDDA.n263 VDDA.n60 585
R875 VDDA.n256 VDDA.n60 585
R876 VDDA.n200 VDDA.n199 585
R877 VDDA.n199 VDDA.n198 585
R878 VDDA.n362 VDDA.n357 585
R879 VDDA.n357 VDDA.n48 585
R880 VDDA.n291 VDDA.n55 585
R881 VDDA.n286 VDDA.n55 585
R882 VDDA.n348 VDDA.n343 585
R883 VDDA.n343 VDDA.n45 585
R884 VDDA.n328 VDDA.n42 585
R885 VDDA.n328 VDDA.n327 585
R886 VDDA.n339 VDDA.n334 585
R887 VDDA.n334 VDDA.n41 585
R888 VDDA.n434 VDDA.n433 585
R889 VDDA.n438 VDDA.n436 585
R890 VDDA.n445 VDDA.n444 585
R891 VDDA.n449 VDDA.n447 585
R892 VDDA.n366 VDDA.n50 585
R893 VDDA.n351 VDDA.n50 585
R894 VDDA.n253 VDDA.n246 585
R895 VDDA.n169 VDDA.n168 585
R896 VDDA.n169 VDDA.n125 585
R897 VDDA.n440 VDDA.t128 465.079
R898 VDDA.t128 VDDA.n439 465.079
R899 VDDA.n451 VDDA.t71 465.079
R900 VDDA.t71 VDDA.n450 465.079
R901 VDDA.n313 VDDA.t119 464.281
R902 VDDA.t119 VDDA.n312 464.281
R903 VDDA.n29 VDDA.t22 464.281
R904 VDDA.t22 VDDA.n26 464.281
R905 VDDA.n474 VDDA.t4 464.281
R906 VDDA.t4 VDDA.n18 464.281
R907 VDDA.t74 VDDA.n457 464.281
R908 VDDA.n458 VDDA.t74 464.281
R909 VDDA.n468 VDDA.t7 464.281
R910 VDDA.t7 VDDA.n467 464.281
R911 VDDA.t117 VDDA.n417 464.281
R912 VDDA.n418 VDDA.t117 464.281
R913 VDDA.n428 VDDA.t28 464.281
R914 VDDA.t28 VDDA.n427 464.281
R915 VDDA.n408 VDDA.t98 464.281
R916 VDDA.t98 VDDA.n407 464.281
R917 VDDA.t24 VDDA.n301 464.281
R918 VDDA.n302 VDDA.t24 464.281
R919 VDDA.t15 VDDA.n317 464.281
R920 VDDA.n318 VDDA.t15 464.281
R921 VDDA.n371 VDDA.t129 415.336
R922 VDDA.n157 VDDA.t47 384.967
R923 VDDA.n161 VDDA.t59 384.967
R924 VDDA.n205 VDDA.t66 384.967
R925 VDDA.n133 VDDA.t63 384.967
R926 VDDA.n150 VDDA.t36 374.878
R927 VDDA.n245 VDDA.t50 352.834
R928 VDDA.t49 VDDA.n130 341.991
R929 VDDA.n134 VDDA.t65 341.752
R930 VDDA.n162 VDDA.t62 341.752
R931 VDDA.n204 VDDA.t69 341.752
R932 VDDA.n197 VDDA.t56 336.329
R933 VDDA.n197 VDDA.t39 336.329
R934 VDDA.n126 VDDA.t53 320.7
R935 VDDA.n264 VDDA.t43 320.7
R936 VDDA.n158 VDDA.n156 315.647
R937 VDDA.n207 VDDA.n81 315.647
R938 VDDA.n132 VDDA.n82 315.647
R939 VDDA.n206 VDDA.n83 315.647
R940 VDDA.n159 VDDA.n138 315.647
R941 VDDA.n160 VDDA.n137 315.647
R942 VDDA.n23 VDDA.t13 315.25
R943 VDDA.t25 VDDA.t16 314.113
R944 VDDA.t33 VDDA.t20 314.113
R945 VDDA.n199 VDDA.n89 291.363
R946 VDDA.n195 VDDA.n87 291.363
R947 VDDA.n196 VDDA.n195 291.363
R948 VDDA.n151 VDDA.n140 290.733
R949 VDDA.n151 VDDA.n141 290.733
R950 VDDA.n257 VDDA.n60 290.733
R951 VDDA.n360 VDDA.n357 290.733
R952 VDDA.n289 VDDA.n55 290.733
R953 VDDA.n346 VDDA.n343 290.733
R954 VDDA.n329 VDDA.n328 290.733
R955 VDDA.n337 VDDA.n334 290.733
R956 VDDA.n352 VDDA.n50 290.733
R957 VDDA.n251 VDDA.n246 290.733
R958 VDDA.n247 VDDA.n246 290.733
R959 VDDA.n169 VDDA.n124 290.733
R960 VDDA.n429 VDDA.n428 243.698
R961 VDDA.n469 VDDA.n468 243.698
R962 VDDA.n475 VDDA.n474 243.698
R963 VDDA.n29 VDDA.n28 243.698
R964 VDDA.n314 VDDA.n313 243.698
R965 VDDA.n407 VDDA.n21 243.698
R966 VDDA.n302 VDDA.n299 243.698
R967 VDDA.n318 VDDA.n297 243.698
R968 VDDA.n458 VDDA.n455 243.698
R969 VDDA.n418 VDDA.n415 243.698
R970 VDDA.n414 VDDA.n1 238.367
R971 VDDA.n453 VDDA.n452 238.367
R972 VDDA.n446 VDDA.n413 238.367
R973 VDDA.n412 VDDA.n13 238.367
R974 VDDA.n478 VDDA.n477 238.367
R975 VDDA.n34 VDDA.n33 238.367
R976 VDDA.n298 VDDA.n38 238.367
R977 VDDA.n422 VDDA.n2 238.367
R978 VDDA.n442 VDDA.n441 238.367
R979 VDDA.n462 VDDA.n14 238.367
R980 VDDA.n410 VDDA.n409 238.367
R981 VDDA.n306 VDDA.n25 238.367
R982 VDDA.n322 VDDA.n37 238.367
R983 VDDA.n435 VDDA.n431 238.367
R984 VDDA.n143 VDDA.n141 233.841
R985 VDDA.n247 VDDA.n63 233.841
R986 VDDA.n254 VDDA.n253 230.308
R987 VDDA.n150 VDDA.n149 230.308
R988 VDDA.n263 VDDA.n262 230.308
R989 VDDA.n260 VDDA.n256 230.308
R990 VDDA.n201 VDDA.n200 230.308
R991 VDDA.n198 VDDA.n84 230.308
R992 VDDA.n340 VDDA.n339 230.308
R993 VDDA.n296 VDDA.n41 230.308
R994 VDDA.n349 VDDA.n348 230.308
R995 VDDA.n295 VDDA.n45 230.308
R996 VDDA.n363 VDDA.n362 230.308
R997 VDDA.n294 VDDA.n48 230.308
R998 VDDA.n292 VDDA.n291 230.308
R999 VDDA.n286 VDDA.n53 230.308
R1000 VDDA.n332 VDDA.n42 230.308
R1001 VDDA.n366 VDDA.n365 230.308
R1002 VDDA.n355 VDDA.n351 230.308
R1003 VDDA.n327 VDDA.n324 230.308
R1004 VDDA.t31 VDDA.t17 222.178
R1005 VDDA.n341 VDDA.n323 199.195
R1006 VDDA.n98 VDDA.n97 196.502
R1007 VDDA.n95 VDDA.n94 196.502
R1008 VDDA.n194 VDDA.n193 196.502
R1009 VDDA.n185 VDDA.n117 196.502
R1010 VDDA.n178 VDDA.n120 196.502
R1011 VDDA.n171 VDDA.n170 196.502
R1012 VDDA.n163 VDDA.n162 185.001
R1013 VDDA.n135 VDDA.n134 185.001
R1014 VDDA.n204 VDDA.n203 185.001
R1015 VDDA.n52 VDDA.n51 185
R1016 VDDA.n354 VDDA.n353 185
R1017 VDDA.n331 VDDA.n330 185
R1018 VDDA.n326 VDDA.n325 185
R1019 VDDA.n321 VDDA.n320 185
R1020 VDDA.n319 VDDA.n316 185
R1021 VDDA.n305 VDDA.n304 185
R1022 VDDA.n303 VDDA.n300 185
R1023 VDDA.n404 VDDA.n22 185
R1024 VDDA.n406 VDDA.n405 185
R1025 VDDA.n461 VDDA.n460 185
R1026 VDDA.n459 VDDA.n456 185
R1027 VDDA.n434 VDDA.n432 185
R1028 VDDA.n438 VDDA.n437 185
R1029 VDDA.n421 VDDA.n420 185
R1030 VDDA.n419 VDDA.n416 185
R1031 VDDA.n290 VDDA.n54 185
R1032 VDDA.n288 VDDA.n287 185
R1033 VDDA.n361 VDDA.n356 185
R1034 VDDA.n359 VDDA.n358 185
R1035 VDDA.n347 VDDA.n342 185
R1036 VDDA.n345 VDDA.n344 185
R1037 VDDA.n338 VDDA.n333 185
R1038 VDDA.n336 VDDA.n335 185
R1039 VDDA.n309 VDDA.n308 185
R1040 VDDA.n311 VDDA.n310 185
R1041 VDDA.n30 VDDA.n27 185
R1042 VDDA.n32 VDDA.n31 185
R1043 VDDA.n473 VDDA.n471 185
R1044 VDDA.n472 VDDA.n19 185
R1045 VDDA.n464 VDDA.n463 185
R1046 VDDA.n466 VDDA.n465 185
R1047 VDDA.n445 VDDA.n443 185
R1048 VDDA.n449 VDDA.n448 185
R1049 VDDA.n424 VDDA.n423 185
R1050 VDDA.n426 VDDA.n425 185
R1051 VDDA.n88 VDDA.n85 185
R1052 VDDA.n91 VDDA.n90 185
R1053 VDDA.n62 VDDA.n61 185
R1054 VDDA.n259 VDDA.n258 185
R1055 VDDA.n148 VDDA.n142 185
R1056 VDDA.n147 VDDA.n146 185
R1057 VDDA.n147 VDDA.n136 185
R1058 VDDA.n145 VDDA.n144 185
R1059 VDDA.n252 VDDA.n65 185
R1060 VDDA.n250 VDDA.n64 185
R1061 VDDA.n255 VDDA.n64 185
R1062 VDDA.n249 VDDA.n248 185
R1063 VDDA.n168 VDDA.n127 185
R1064 VDDA.n164 VDDA.n127 185
R1065 VDDA.n167 VDDA.n166 185
R1066 VDDA.n129 VDDA.n128 185
R1067 VDDA.n131 VDDA.n125 185
R1068 VDDA.n164 VDDA.n131 185
R1069 VDDA.t17 VDDA.n293 172.38
R1070 VDDA.n364 VDDA.t99 172.38
R1071 VDDA.n350 VDDA.t0 172.38
R1072 VDDA.n198 VDDA.n197 166.63
R1073 VDDA.n425 VDDA.n423 150
R1074 VDDA.n448 VDDA.n443 150
R1075 VDDA.n465 VDDA.n463 150
R1076 VDDA.n471 VDDA.n19 150
R1077 VDDA.n32 VDDA.n27 150
R1078 VDDA.n310 VDDA.n308 150
R1079 VDDA.n421 VDDA.n416 150
R1080 VDDA.n437 VDDA.n432 150
R1081 VDDA.n461 VDDA.n456 150
R1082 VDDA.n405 VDDA.n22 150
R1083 VDDA.n305 VDDA.n300 150
R1084 VDDA.n321 VDDA.n316 150
R1085 VDDA.n315 VDDA.n307 137.904
R1086 VDDA.n411 VDDA.n20 137.904
R1087 VDDA.n293 VDDA.t123 126.412
R1088 VDDA.n364 VDDA.t31 126.412
R1089 VDDA.t99 VDDA.n350 126.412
R1090 VDDA.t0 VDDA.n341 126.412
R1091 VDDA.t35 VDDA.n433 123.126
R1092 VDDA.n436 VDDA.t35 123.126
R1093 VDDA.t127 VDDA.n444 123.126
R1094 VDDA.n447 VDDA.t127 123.126
R1095 VDDA.n65 VDDA.n64 120.001
R1096 VDDA.n248 VDDA.n64 120.001
R1097 VDDA.n148 VDDA.n147 120.001
R1098 VDDA.n147 VDDA.n144 120.001
R1099 VDDA.n259 VDDA.n62 120.001
R1100 VDDA.n90 VDDA.n85 120.001
R1101 VDDA.n335 VDDA.n333 120.001
R1102 VDDA.n344 VDDA.n342 120.001
R1103 VDDA.n358 VDDA.n356 120.001
R1104 VDDA.n287 VDDA.n54 120.001
R1105 VDDA.n331 VDDA.n325 120.001
R1106 VDDA.n354 VDDA.n52 120.001
R1107 VDDA.n166 VDDA.n127 120.001
R1108 VDDA.n131 VDDA.n129 120.001
R1109 VDDA.n233 VDDA.n69 119.737
R1110 VDDA.n226 VDDA.n72 119.737
R1111 VDDA.n219 VDDA.n75 119.737
R1112 VDDA.n212 VDDA.n78 119.737
R1113 VDDA.n154 VDDA.n152 119.737
R1114 VDDA.n476 VDDA.n470 107.258
R1115 VDDA.n470 VDDA.t6 103.427
R1116 VDDA.t70 VDDA.n454 103.427
R1117 VDDA.n454 VDDA.t34 103.427
R1118 VDDA.t27 VDDA.n430 103.427
R1119 VDDA.n476 VDDA.t97 95.7666
R1120 VDDA.t118 VDDA.t14 91.936
R1121 VDDA.t21 VDDA.t23 91.936
R1122 VDDA.t3 VDDA.t12 84.2747
R1123 VDDA.t6 VDDA.t25 84.2747
R1124 VDDA.t16 VDDA.t70 84.2747
R1125 VDDA.t34 VDDA.t33 84.2747
R1126 VDDA.t20 VDDA.t27 84.2747
R1127 VDDA.n207 VDDA.n82 83.2005
R1128 VDDA.n207 VDDA.n206 83.2005
R1129 VDDA.n159 VDDA.n158 83.2005
R1130 VDDA.n160 VDDA.n159 83.2005
R1131 VDDA.n365 VDDA.n364 69.8479
R1132 VDDA.n364 VDDA.n355 69.8479
R1133 VDDA.n341 VDDA.n332 69.8479
R1134 VDDA.n341 VDDA.n324 69.8479
R1135 VDDA.n293 VDDA.n292 69.8479
R1136 VDDA.n293 VDDA.n53 69.8479
R1137 VDDA.n364 VDDA.n363 69.8479
R1138 VDDA.n364 VDDA.n294 69.8479
R1139 VDDA.n350 VDDA.n349 69.8479
R1140 VDDA.n350 VDDA.n295 69.8479
R1141 VDDA.n341 VDDA.n340 69.8479
R1142 VDDA.n341 VDDA.n296 69.8479
R1143 VDDA.n202 VDDA.n201 69.8479
R1144 VDDA.n202 VDDA.n84 69.8479
R1145 VDDA.n262 VDDA.n261 69.8479
R1146 VDDA.n261 VDDA.n260 69.8479
R1147 VDDA.n149 VDDA.n136 69.8479
R1148 VDDA.n143 VDDA.n136 69.8479
R1149 VDDA.n255 VDDA.n254 69.8479
R1150 VDDA.n255 VDDA.n63 69.8479
R1151 VDDA.n165 VDDA.n164 69.8479
R1152 VDDA.n159 VDDA.n155 69.3203
R1153 VDDA.n323 VDDA.n322 65.8183
R1154 VDDA.n323 VDDA.n297 65.8183
R1155 VDDA.n307 VDDA.n306 65.8183
R1156 VDDA.n307 VDDA.n299 65.8183
R1157 VDDA.n411 VDDA.n410 65.8183
R1158 VDDA.n411 VDDA.n21 65.8183
R1159 VDDA.n470 VDDA.n462 65.8183
R1160 VDDA.n470 VDDA.n455 65.8183
R1161 VDDA.n454 VDDA.n442 65.8183
R1162 VDDA.n454 VDDA.n431 65.8183
R1163 VDDA.n430 VDDA.n422 65.8183
R1164 VDDA.n430 VDDA.n415 65.8183
R1165 VDDA.n315 VDDA.n314 65.8183
R1166 VDDA.n315 VDDA.n298 65.8183
R1167 VDDA.n28 VDDA.n20 65.8183
R1168 VDDA.n33 VDDA.n20 65.8183
R1169 VDDA.n476 VDDA.n475 65.8183
R1170 VDDA.n477 VDDA.n476 65.8183
R1171 VDDA.n470 VDDA.n469 65.8183
R1172 VDDA.n470 VDDA.n412 65.8183
R1173 VDDA.n454 VDDA.n453 65.8183
R1174 VDDA.n454 VDDA.n413 65.8183
R1175 VDDA.n430 VDDA.n429 65.8183
R1176 VDDA.n430 VDDA.n414 65.8183
R1177 VDDA.n389 VDDA.n38 58.0576
R1178 VDDA.n396 VDDA.n34 58.0576
R1179 VDDA.n479 VDDA.n478 58.0576
R1180 VDDA.n485 VDDA.n14 58.0576
R1181 VDDA.n485 VDDA.n13 58.0576
R1182 VDDA.n513 VDDA.n2 58.0576
R1183 VDDA.n513 VDDA.n1 58.0576
R1184 VDDA.n409 VDDA.n403 58.0576
R1185 VDDA.n397 VDDA.n25 58.0576
R1186 VDDA.n390 VDDA.n37 58.0576
R1187 VDDA.n367 VDDA.n48 57.2449
R1188 VDDA.n286 VDDA.n285 57.2449
R1189 VDDA.n374 VDDA.n45 57.2449
R1190 VDDA.n381 VDDA.n42 57.2449
R1191 VDDA.n381 VDDA.n41 57.2449
R1192 VDDA.n367 VDDA.n366 57.2449
R1193 VDDA.n498 VDDA.n8 54.4005
R1194 VDDA.n498 VDDA.n7 54.4005
R1195 VDDA.n500 VDDA.n7 54.4005
R1196 VDDA.n500 VDDA.n8 54.4005
R1197 VDDA.n416 VDDA.n415 53.3664
R1198 VDDA.n437 VDDA.n431 53.3664
R1199 VDDA.n456 VDDA.n455 53.3664
R1200 VDDA.n322 VDDA.n321 53.3664
R1201 VDDA.n316 VDDA.n297 53.3664
R1202 VDDA.n306 VDDA.n305 53.3664
R1203 VDDA.n300 VDDA.n299 53.3664
R1204 VDDA.n410 VDDA.n22 53.3664
R1205 VDDA.n405 VDDA.n21 53.3664
R1206 VDDA.n462 VDDA.n461 53.3664
R1207 VDDA.n442 VDDA.n432 53.3664
R1208 VDDA.n422 VDDA.n421 53.3664
R1209 VDDA.n314 VDDA.n308 53.3664
R1210 VDDA.n310 VDDA.n298 53.3664
R1211 VDDA.n28 VDDA.n27 53.3664
R1212 VDDA.n33 VDDA.n32 53.3664
R1213 VDDA.n475 VDDA.n471 53.3664
R1214 VDDA.n477 VDDA.n19 53.3664
R1215 VDDA.n469 VDDA.n463 53.3664
R1216 VDDA.n465 VDDA.n412 53.3664
R1217 VDDA.n453 VDDA.n443 53.3664
R1218 VDDA.n448 VDDA.n413 53.3664
R1219 VDDA.n429 VDDA.n423 53.3664
R1220 VDDA.n425 VDDA.n414 53.3664
R1221 VDDA.n156 VDDA.t49 49.2505
R1222 VDDA.n156 VDDA.t110 49.2505
R1223 VDDA.n81 VDDA.t106 49.2505
R1224 VDDA.n81 VDDA.t104 49.2505
R1225 VDDA.t65 VDDA.n132 49.2505
R1226 VDDA.n132 VDDA.t108 49.2505
R1227 VDDA.n83 VDDA.t102 49.2505
R1228 VDDA.n83 VDDA.t68 49.2505
R1229 VDDA.n138 VDDA.t112 49.2505
R1230 VDDA.n138 VDDA.t116 49.2505
R1231 VDDA.n137 VDDA.t114 49.2505
R1232 VDDA.n137 VDDA.t61 49.2505
R1233 VDDA.n248 VDDA.n63 45.3071
R1234 VDDA.n144 VDDA.n143 45.3071
R1235 VDDA.n325 VDDA.n324 45.3071
R1236 VDDA.n355 VDDA.n354 45.3071
R1237 VDDA.n365 VDDA.n52 45.3071
R1238 VDDA.n332 VDDA.n331 45.3071
R1239 VDDA.n292 VDDA.n54 45.3071
R1240 VDDA.n287 VDDA.n53 45.3071
R1241 VDDA.n363 VDDA.n356 45.3071
R1242 VDDA.n358 VDDA.n294 45.3071
R1243 VDDA.n349 VDDA.n342 45.3071
R1244 VDDA.n344 VDDA.n295 45.3071
R1245 VDDA.n340 VDDA.n333 45.3071
R1246 VDDA.n335 VDDA.n296 45.3071
R1247 VDDA.n201 VDDA.n85 45.3071
R1248 VDDA.n90 VDDA.n84 45.3071
R1249 VDDA.n262 VDDA.n62 45.3071
R1250 VDDA.n260 VDDA.n259 45.3071
R1251 VDDA.n149 VDDA.n148 45.3071
R1252 VDDA.n254 VDDA.n65 45.3071
R1253 VDDA.n166 VDDA.n165 45.3071
R1254 VDDA.n165 VDDA.n129 45.3071
R1255 VDDA.n208 VDDA.n207 41.6005
R1256 VDDA.n155 VDDA.n139 39.4988
R1257 VDDA.n271 VDDA.n270 38.1005
R1258 VDDA.t60 VDDA.n163 38.0466
R1259 VDDA.n514 VDDA.n513 34.9005
R1260 VDDA.t8 VDDA.t79 32.2821
R1261 VDDA.n200 VDDA.n86 32.2291
R1262 VDDA.n266 VDDA.n57 32.0005
R1263 VDDA.n270 VDDA.n57 32.0005
R1264 VDDA.n104 VDDA.n103 32.0005
R1265 VDDA.n103 VDDA.n102 32.0005
R1266 VDDA.n110 VDDA.n92 32.0005
R1267 VDDA.n110 VDDA.n109 32.0005
R1268 VDDA.n109 VDDA.n108 32.0005
R1269 VDDA.n192 VDDA.n114 32.0005
R1270 VDDA.n187 VDDA.n186 32.0005
R1271 VDDA.n180 VDDA.n179 32.0005
R1272 VDDA.n180 VDDA.n118 32.0005
R1273 VDDA.n184 VDDA.n118 32.0005
R1274 VDDA.n173 VDDA.n172 32.0005
R1275 VDDA.n173 VDDA.n121 32.0005
R1276 VDDA.n177 VDDA.n121 32.0005
R1277 VDDA.n284 VDDA.n274 32.0005
R1278 VDDA.n280 VDDA.n274 32.0005
R1279 VDDA.n280 VDDA.n279 32.0005
R1280 VDDA.n279 VDDA.n278 32.0005
R1281 VDDA.n278 VDDA.n49 32.0005
R1282 VDDA.n367 VDDA.n49 32.0005
R1283 VDDA.n368 VDDA.n367 32.0005
R1284 VDDA.n368 VDDA.n46 32.0005
R1285 VDDA.n373 VDDA.n46 32.0005
R1286 VDDA.n376 VDDA.n375 32.0005
R1287 VDDA.n376 VDDA.n43 32.0005
R1288 VDDA.n380 VDDA.n43 32.0005
R1289 VDDA.n383 VDDA.n382 32.0005
R1290 VDDA.n383 VDDA.n39 32.0005
R1291 VDDA.n387 VDDA.n39 32.0005
R1292 VDDA.n388 VDDA.n387 32.0005
R1293 VDDA.n391 VDDA.n35 32.0005
R1294 VDDA.n395 VDDA.n35 32.0005
R1295 VDDA.n399 VDDA.n398 32.0005
R1296 VDDA.n480 VDDA.n17 32.0005
R1297 VDDA.n484 VDDA.n15 32.0005
R1298 VDDA.n487 VDDA.n486 32.0005
R1299 VDDA.n487 VDDA.n11 32.0005
R1300 VDDA.n491 VDDA.n11 32.0005
R1301 VDDA.n492 VDDA.n491 32.0005
R1302 VDDA.n493 VDDA.n492 32.0005
R1303 VDDA.n493 VDDA.n9 32.0005
R1304 VDDA.n497 VDDA.n9 32.0005
R1305 VDDA.n501 VDDA.n5 32.0005
R1306 VDDA.n505 VDDA.n5 32.0005
R1307 VDDA.n506 VDDA.n505 32.0005
R1308 VDDA.n507 VDDA.n506 32.0005
R1309 VDDA.n507 VDDA.n3 32.0005
R1310 VDDA.n511 VDDA.n3 32.0005
R1311 VDDA.n512 VDDA.n511 32.0005
R1312 VDDA.n139 VDDA.n80 32.0005
R1313 VDDA.n209 VDDA.n80 32.0005
R1314 VDDA.n214 VDDA.n77 32.0005
R1315 VDDA.n215 VDDA.n214 32.0005
R1316 VDDA.n216 VDDA.n215 32.0005
R1317 VDDA.n216 VDDA.n74 32.0005
R1318 VDDA.n221 VDDA.n74 32.0005
R1319 VDDA.n222 VDDA.n221 32.0005
R1320 VDDA.n223 VDDA.n222 32.0005
R1321 VDDA.n223 VDDA.n71 32.0005
R1322 VDDA.n228 VDDA.n71 32.0005
R1323 VDDA.n229 VDDA.n228 32.0005
R1324 VDDA.n230 VDDA.n229 32.0005
R1325 VDDA.n230 VDDA.n68 32.0005
R1326 VDDA.n235 VDDA.n68 32.0005
R1327 VDDA.n236 VDDA.n235 32.0005
R1328 VDDA.n242 VDDA.n236 32.0005
R1329 VDDA.n242 VDDA.n241 32.0005
R1330 VDDA.n241 VDDA.n240 32.0005
R1331 VDDA.n240 VDDA.n237 32.0005
R1332 VDDA.n162 VDDA.n161 30.754
R1333 VDDA.n205 VDDA.n204 30.754
R1334 VDDA.n134 VDDA.n133 30.186
R1335 VDDA.t48 VDDA.t109 29.9762
R1336 VDDA.t111 VDDA.t115 29.9762
R1337 VDDA.t92 VDDA.t91 29.9762
R1338 VDDA.n157 VDDA.n130 29.9467
R1339 VDDA.t113 VDDA.t85 28.8233
R1340 VDDA.n265 VDDA.n59 28.8005
R1341 VDDA.n104 VDDA.n95 28.8005
R1342 VDDA.n193 VDDA.n192 28.8005
R1343 VDDA.n374 VDDA.n373 28.8005
R1344 VDDA.t29 VDDA.t95 27.6704
R1345 VDDA.t72 VDDA.t5 26.5175
R1346 VDDA.n285 VDDA.n284 25.6005
R1347 VDDA.n381 VDDA.n380 25.6005
R1348 VDDA.n391 VDDA.n390 25.6005
R1349 VDDA.n403 VDDA.n402 25.6005
R1350 VDDA.n479 VDDA.n15 25.6005
R1351 VDDA.n485 VDDA.n484 25.6005
R1352 VDDA.n499 VDDA.n498 25.6005
R1353 VDDA.n500 VDDA.n499 25.6005
R1354 VDDA.n209 VDDA.n208 25.6005
R1355 VDDA.n237 VDDA 25.6005
R1356 VDDA.t83 VDDA.n135 25.3646
R1357 VDDA.n97 VDDA.t126 24.6255
R1358 VDDA.n97 VDDA.t45 24.6255
R1359 VDDA.n94 VDDA.t80 24.6255
R1360 VDDA.n94 VDDA.t76 24.6255
R1361 VDDA.t58 VDDA.n194 24.6255
R1362 VDDA.n194 VDDA.t30 24.6255
R1363 VDDA.n117 VDDA.t90 24.6255
R1364 VDDA.n117 VDDA.t41 24.6255
R1365 VDDA.n120 VDDA.t86 24.6255
R1366 VDDA.n120 VDDA.t84 24.6255
R1367 VDDA.n170 VDDA.t55 24.6255
R1368 VDDA.n170 VDDA.t88 24.6255
R1369 VDDA.t55 VDDA.n169 24.6255
R1370 VDDA.n60 VDDA.t46 24.6255
R1371 VDDA.n195 VDDA.t58 24.6255
R1372 VDDA.n199 VDDA.t42 24.6255
R1373 VDDA.n50 VDDA.t122 24.6255
R1374 VDDA.n357 VDDA.t32 24.6255
R1375 VDDA.n55 VDDA.t124 24.6255
R1376 VDDA.n343 VDDA.t100 24.6255
R1377 VDDA.n328 VDDA.t2 24.6255
R1378 VDDA.n334 VDDA.t1 24.6255
R1379 VDDA.n126 VDDA.n123 24.361
R1380 VDDA.t78 VDDA.t75 24.2117
R1381 VDDA.t44 VDDA.t77 24.2117
R1382 VDDA.n102 VDDA.n98 22.4005
R1383 VDDA.n186 VDDA.n185 22.4005
R1384 VDDA.n187 VDDA.n86 22.4005
R1385 VDDA.n253 VDDA.n245 22.0449
R1386 VDDA.t87 VDDA.t113 21.9058
R1387 VDDA.t40 VDDA.t105 21.9058
R1388 VDDA.t81 VDDA.t103 21.9058
R1389 VDDA.n255 VDDA.t77 21.9058
R1390 VDDA.n202 VDDA.t120 20.7529
R1391 VDDA.t38 VDDA.n151 19.7005
R1392 VDDA.n246 VDDA.t52 19.7005
R1393 VDDA.n69 VDDA.t11 19.7005
R1394 VDDA.n69 VDDA.t51 19.7005
R1395 VDDA.n72 VDDA.t94 19.7005
R1396 VDDA.n72 VDDA.t73 19.7005
R1397 VDDA.n75 VDDA.t96 19.7005
R1398 VDDA.n75 VDDA.t9 19.7005
R1399 VDDA.n78 VDDA.t121 19.7005
R1400 VDDA.n78 VDDA.t82 19.7005
R1401 VDDA.n152 VDDA.t38 19.7005
R1402 VDDA.n152 VDDA.t19 19.7005
R1403 VDDA.t64 VDDA.t18 19.6
R1404 VDDA.n399 VDDA.n23 19.2005
R1405 VDDA.n265 VDDA.n264 17.6005
R1406 VDDA.t109 VDDA.t54 17.2942
R1407 VDDA.n203 VDDA.t8 16.1413
R1408 VDDA.n98 VDDA.n59 16.0005
R1409 VDDA.n114 VDDA.n86 16.0005
R1410 VDDA.n185 VDDA.n184 16.0005
R1411 VDDA.n172 VDDA.n171 16.0005
R1412 VDDA.n398 VDDA.n397 16.0005
R1413 VDDA.n161 VDDA.n160 16.0005
R1414 VDDA.n206 VDDA.n205 16.0005
R1415 VDDA.n133 VDDA.n82 16.0005
R1416 VDDA.n158 VDDA.n157 16.0005
R1417 VDDA VDDA.n56 15.7005
R1418 VDDA.n264 VDDA.n263 15.6449
R1419 VDDA.n168 VDDA.n126 15.6449
R1420 VDDA.t57 VDDA.t101 14.9884
R1421 VDDA.t67 VDDA.t57 14.9884
R1422 VDDA.t5 VDDA.t125 14.9884
R1423 VDDA.n285 VDDA.n273 13.9187
R1424 VDDA.t37 VDDA.t89 13.8355
R1425 VDDA.t79 VDDA.t93 13.8355
R1426 VDDA.n272 VDDA.n56 13.0501
R1427 VDDA.n396 VDDA.n395 12.8005
R1428 VDDA.n402 VDDA.n23 12.8005
R1429 VDDA.t54 VDDA.t111 12.6825
R1430 VDDA.t89 VDDA.t64 12.6825
R1431 VDDA.t93 VDDA.t78 12.6825
R1432 VDDA.n273 VDDA.n272 12.425
R1433 VDDA.n272 VDDA.n271 11.7059
R1434 VDDA.n135 VDDA.t37 11.5296
R1435 VDDA.n323 VDDA.t118 11.4924
R1436 VDDA.t14 VDDA.n315 11.4924
R1437 VDDA.n307 VDDA.t21 11.4924
R1438 VDDA.t23 VDDA.n20 11.4924
R1439 VDDA.t12 VDDA.n411 11.4924
R1440 VDDA.t18 VDDA.t107 10.3767
R1441 VDDA.t10 VDDA.t92 10.3767
R1442 VDDA.n245 VDDA.n244 9.613
R1443 VDDA.n266 VDDA.n265 9.6005
R1444 VDDA.n193 VDDA.n92 9.6005
R1445 VDDA.n108 VDDA.n95 9.6005
R1446 VDDA.n238 VDDA.n237 9.3005
R1447 VDDA.n240 VDDA.n239 9.3005
R1448 VDDA.n241 VDDA.n67 9.3005
R1449 VDDA.n243 VDDA.n242 9.3005
R1450 VDDA.n236 VDDA.n66 9.3005
R1451 VDDA.n235 VDDA.n234 9.3005
R1452 VDDA.n232 VDDA.n68 9.3005
R1453 VDDA.n231 VDDA.n230 9.3005
R1454 VDDA.n229 VDDA.n70 9.3005
R1455 VDDA.n228 VDDA.n227 9.3005
R1456 VDDA.n225 VDDA.n71 9.3005
R1457 VDDA.n224 VDDA.n223 9.3005
R1458 VDDA.n222 VDDA.n73 9.3005
R1459 VDDA.n221 VDDA.n220 9.3005
R1460 VDDA.n218 VDDA.n74 9.3005
R1461 VDDA.n217 VDDA.n216 9.3005
R1462 VDDA.n215 VDDA.n76 9.3005
R1463 VDDA.n214 VDDA.n213 9.3005
R1464 VDDA.n211 VDDA.n77 9.3005
R1465 VDDA.n153 VDDA.n139 9.3005
R1466 VDDA.n80 VDDA.n79 9.3005
R1467 VDDA.n210 VDDA.n209 9.3005
R1468 VDDA.n172 VDDA.n122 9.3005
R1469 VDDA.n174 VDDA.n173 9.3005
R1470 VDDA.n175 VDDA.n121 9.3005
R1471 VDDA.n177 VDDA.n176 9.3005
R1472 VDDA.n179 VDDA.n119 9.3005
R1473 VDDA.n181 VDDA.n180 9.3005
R1474 VDDA.n182 VDDA.n118 9.3005
R1475 VDDA.n184 VDDA.n183 9.3005
R1476 VDDA.n185 VDDA.n116 9.3005
R1477 VDDA.n186 VDDA.n115 9.3005
R1478 VDDA.n188 VDDA.n187 9.3005
R1479 VDDA.n189 VDDA.n86 9.3005
R1480 VDDA.n190 VDDA.n114 9.3005
R1481 VDDA.n192 VDDA.n191 9.3005
R1482 VDDA.n193 VDDA.n113 9.3005
R1483 VDDA.n112 VDDA.n92 9.3005
R1484 VDDA.n111 VDDA.n110 9.3005
R1485 VDDA.n109 VDDA.n93 9.3005
R1486 VDDA.n108 VDDA.n107 9.3005
R1487 VDDA.n106 VDDA.n95 9.3005
R1488 VDDA.n105 VDDA.n104 9.3005
R1489 VDDA.n103 VDDA.n96 9.3005
R1490 VDDA.n102 VDDA.n101 9.3005
R1491 VDDA.n100 VDDA.n98 9.3005
R1492 VDDA.n99 VDDA.n59 9.3005
R1493 VDDA.n265 VDDA.n58 9.3005
R1494 VDDA.n267 VDDA.n266 9.3005
R1495 VDDA.n268 VDDA.n57 9.3005
R1496 VDDA.n270 VDDA.n269 9.3005
R1497 VDDA.n284 VDDA.n283 9.3005
R1498 VDDA.n282 VDDA.n274 9.3005
R1499 VDDA.n281 VDDA.n280 9.3005
R1500 VDDA.n279 VDDA.n275 9.3005
R1501 VDDA.n278 VDDA.n277 9.3005
R1502 VDDA.n276 VDDA.n49 9.3005
R1503 VDDA.n367 VDDA.n47 9.3005
R1504 VDDA.n369 VDDA.n368 9.3005
R1505 VDDA.n370 VDDA.n46 9.3005
R1506 VDDA.n373 VDDA.n372 9.3005
R1507 VDDA.n375 VDDA.n44 9.3005
R1508 VDDA.n377 VDDA.n376 9.3005
R1509 VDDA.n378 VDDA.n43 9.3005
R1510 VDDA.n380 VDDA.n379 9.3005
R1511 VDDA.n382 VDDA.n40 9.3005
R1512 VDDA.n384 VDDA.n383 9.3005
R1513 VDDA.n385 VDDA.n39 9.3005
R1514 VDDA.n387 VDDA.n386 9.3005
R1515 VDDA.n388 VDDA.n36 9.3005
R1516 VDDA.n392 VDDA.n391 9.3005
R1517 VDDA.n393 VDDA.n35 9.3005
R1518 VDDA.n395 VDDA.n394 9.3005
R1519 VDDA.n398 VDDA.n24 9.3005
R1520 VDDA.n400 VDDA.n399 9.3005
R1521 VDDA.n402 VDDA.n401 9.3005
R1522 VDDA.n17 VDDA.n16 9.3005
R1523 VDDA.n481 VDDA.n480 9.3005
R1524 VDDA.n482 VDDA.n15 9.3005
R1525 VDDA.n484 VDDA.n483 9.3005
R1526 VDDA.n486 VDDA.n12 9.3005
R1527 VDDA.n488 VDDA.n487 9.3005
R1528 VDDA.n489 VDDA.n11 9.3005
R1529 VDDA.n491 VDDA.n490 9.3005
R1530 VDDA.n492 VDDA.n10 9.3005
R1531 VDDA.n494 VDDA.n493 9.3005
R1532 VDDA.n495 VDDA.n9 9.3005
R1533 VDDA.n497 VDDA.n496 9.3005
R1534 VDDA.n499 VDDA.n6 9.3005
R1535 VDDA.n502 VDDA.n501 9.3005
R1536 VDDA.n503 VDDA.n5 9.3005
R1537 VDDA.n505 VDDA.n504 9.3005
R1538 VDDA.n506 VDDA.n4 9.3005
R1539 VDDA.n508 VDDA.n507 9.3005
R1540 VDDA.n509 VDDA.n3 9.3005
R1541 VDDA.n511 VDDA.n510 9.3005
R1542 VDDA.n512 VDDA.n0 9.3005
R1543 VDDA.n136 VDDA.t83 9.2238
R1544 VDDA.n311 VDDA.n309 9.14336
R1545 VDDA.n31 VDDA.n30 9.14336
R1546 VDDA.n473 VDDA.n472 9.14336
R1547 VDDA.n460 VDDA.n459 9.14336
R1548 VDDA.n466 VDDA.n464 9.14336
R1549 VDDA.n420 VDDA.n419 9.14336
R1550 VDDA.n426 VDDA.n424 9.14336
R1551 VDDA.n406 VDDA.n404 9.14336
R1552 VDDA.n304 VDDA.n303 9.14336
R1553 VDDA.n320 VDDA.n319 9.14336
R1554 VDDA.t115 VDDA.t87 8.07089
R1555 VDDA.t107 VDDA.t40 8.07089
R1556 VDDA.t101 VDDA.t81 8.07089
R1557 VDDA.t95 VDDA.t67 8.07089
R1558 VDDA.t97 VDDA.t3 7.66179
R1559 VDDA.n150 VDDA.n142 7.11161
R1560 VDDA.n146 VDDA.n145 7.11161
R1561 VDDA.n263 VDDA.n61 7.11161
R1562 VDDA.n258 VDDA.n256 7.11161
R1563 VDDA.n362 VDDA.n361 7.11161
R1564 VDDA.n359 VDDA.n48 7.11161
R1565 VDDA.n291 VDDA.n290 7.11161
R1566 VDDA.n288 VDDA.n286 7.11161
R1567 VDDA.n348 VDDA.n347 7.11161
R1568 VDDA.n345 VDDA.n45 7.11161
R1569 VDDA.n330 VDDA.n42 7.11161
R1570 VDDA.n327 VDDA.n326 7.11161
R1571 VDDA.n339 VDDA.n338 7.11161
R1572 VDDA.n336 VDDA.n41 7.11161
R1573 VDDA.n366 VDDA.n51 7.11161
R1574 VDDA.n353 VDDA.n351 7.11161
R1575 VDDA.n253 VDDA.n252 7.11161
R1576 VDDA.n250 VDDA.n249 7.11161
R1577 VDDA.n168 VDDA.n167 7.11161
R1578 VDDA.n128 VDDA.n125 7.11161
R1579 VDDA.n171 VDDA.n123 6.54033
R1580 VDDA.n382 VDDA.n381 6.4005
R1581 VDDA.n403 VDDA.n17 6.4005
R1582 VDDA.n480 VDDA.n479 6.4005
R1583 VDDA.n486 VDDA.n485 6.4005
R1584 VDDA.n498 VDDA.n497 6.4005
R1585 VDDA.n501 VDDA.n500 6.4005
R1586 VDDA.n513 VDDA.n512 6.4005
R1587 VDDA.n208 VDDA.n77 6.4005
R1588 VDDA.n438 VDDA.n434 5.81868
R1589 VDDA.n449 VDDA.n445 5.81868
R1590 VDDA.t105 VDDA.t120 5.76506
R1591 VDDA.t75 VDDA.t26 5.76506
R1592 VDDA.t91 VDDA.t44 5.76506
R1593 VDDA.n312 VDDA.n38 5.33286
R1594 VDDA.n34 VDDA.n26 5.33286
R1595 VDDA.n478 VDDA.n18 5.33286
R1596 VDDA.n457 VDDA.n14 5.33286
R1597 VDDA.n467 VDDA.n13 5.33286
R1598 VDDA.n417 VDDA.n2 5.33286
R1599 VDDA.n427 VDDA.n1 5.33286
R1600 VDDA.n409 VDDA.n408 5.33286
R1601 VDDA.n301 VDDA.n25 5.33286
R1602 VDDA.n317 VDDA.n37 5.33286
R1603 VDDA.t125 VDDA.t10 4.61215
R1604 VDDA.n313 VDDA.n309 3.75335
R1605 VDDA.n312 VDDA.n311 3.75335
R1606 VDDA.n30 VDDA.n29 3.75335
R1607 VDDA.n31 VDDA.n26 3.75335
R1608 VDDA.n474 VDDA.n473 3.75335
R1609 VDDA.n472 VDDA.n18 3.75335
R1610 VDDA.n460 VDDA.n457 3.75335
R1611 VDDA.n459 VDDA.n458 3.75335
R1612 VDDA.n468 VDDA.n464 3.75335
R1613 VDDA.n467 VDDA.n466 3.75335
R1614 VDDA.n420 VDDA.n417 3.75335
R1615 VDDA.n419 VDDA.n418 3.75335
R1616 VDDA.n428 VDDA.n424 3.75335
R1617 VDDA.n427 VDDA.n426 3.75335
R1618 VDDA.n408 VDDA.n404 3.75335
R1619 VDDA.n407 VDDA.n406 3.75335
R1620 VDDA.n304 VDDA.n301 3.75335
R1621 VDDA.n303 VDDA.n302 3.75335
R1622 VDDA.n320 VDDA.n317 3.75335
R1623 VDDA.n319 VDDA.n318 3.75335
R1624 VDDA.n142 VDDA.n140 3.53508
R1625 VDDA.n145 VDDA.n141 3.53508
R1626 VDDA.n146 VDDA.n140 3.53508
R1627 VDDA.n257 VDDA.n61 3.53508
R1628 VDDA.n258 VDDA.n257 3.53508
R1629 VDDA.n361 VDDA.n360 3.53508
R1630 VDDA.n360 VDDA.n359 3.53508
R1631 VDDA.n290 VDDA.n289 3.53508
R1632 VDDA.n289 VDDA.n288 3.53508
R1633 VDDA.n347 VDDA.n346 3.53508
R1634 VDDA.n346 VDDA.n345 3.53508
R1635 VDDA.n330 VDDA.n329 3.53508
R1636 VDDA.n329 VDDA.n326 3.53508
R1637 VDDA.n338 VDDA.n337 3.53508
R1638 VDDA.n337 VDDA.n336 3.53508
R1639 VDDA.n352 VDDA.n51 3.53508
R1640 VDDA.n353 VDDA.n352 3.53508
R1641 VDDA.n252 VDDA.n251 3.53508
R1642 VDDA.n249 VDDA.n247 3.53508
R1643 VDDA.n251 VDDA.n250 3.53508
R1644 VDDA.n167 VDDA.n124 3.53508
R1645 VDDA.n128 VDDA.n124 3.53508
R1646 VDDA.t103 VDDA.n202 3.45924
R1647 VDDA.t26 VDDA.t72 3.45924
R1648 VDDA.n441 VDDA.n440 3.40194
R1649 VDDA.n439 VDDA.n435 3.40194
R1650 VDDA.n452 VDDA.n451 3.40194
R1651 VDDA.n450 VDDA.n446 3.40194
R1652 VDDA.n179 VDDA.n178 3.2005
R1653 VDDA.n178 VDDA.n177 3.2005
R1654 VDDA.n375 VDDA.n374 3.2005
R1655 VDDA.n389 VDDA.n388 3.2005
R1656 VDDA.n390 VDDA.n389 3.2005
R1657 VDDA.n397 VDDA.n396 3.2005
R1658 VDDA.n440 VDDA.n434 2.39444
R1659 VDDA.n439 VDDA.n438 2.39444
R1660 VDDA.n451 VDDA.n445 2.39444
R1661 VDDA.n450 VDDA.n449 2.39444
R1662 VDDA.n441 VDDA.n8 2.32777
R1663 VDDA.n446 VDDA.n7 2.32777
R1664 VDDA.n163 VDDA.n136 2.30633
R1665 VDDA.n203 VDDA.t29 2.30633
R1666 VDDA.n261 VDDA.n255 2.30633
R1667 VDDA.n88 VDDA.n87 2.27782
R1668 VDDA.n89 VDDA.n88 2.27782
R1669 VDDA.n198 VDDA.n196 2.27782
R1670 VDDA.n91 VDDA.n89 2.27782
R1671 VDDA.n200 VDDA.n87 2.27782
R1672 VDDA.n196 VDDA.n91 2.27782
R1673 VDDA.n164 VDDA.t48 1.15341
R1674 VDDA.t85 VDDA.t60 1.15341
R1675 VDDA.n123 VDDA.n122 0.703395
R1676 VDDA.n283 VDDA.n273 0.194055
R1677 VDDA.n238 VDDA.n56 0.188
R1678 VDDA.n153 VDDA.n79 0.15675
R1679 VDDA.n210 VDDA.n79 0.15675
R1680 VDDA.n211 VDDA.n210 0.15675
R1681 VDDA.n213 VDDA.n76 0.15675
R1682 VDDA.n217 VDDA.n76 0.15675
R1683 VDDA.n218 VDDA.n217 0.15675
R1684 VDDA.n220 VDDA.n73 0.15675
R1685 VDDA.n224 VDDA.n73 0.15675
R1686 VDDA.n225 VDDA.n224 0.15675
R1687 VDDA.n227 VDDA.n70 0.15675
R1688 VDDA.n231 VDDA.n70 0.15675
R1689 VDDA.n232 VDDA.n231 0.15675
R1690 VDDA.n234 VDDA.n66 0.15675
R1691 VDDA.n243 VDDA.n67 0.15675
R1692 VDDA.n239 VDDA.n67 0.15675
R1693 VDDA.n239 VDDA.n238 0.15675
R1694 VDDA.n174 VDDA.n122 0.15675
R1695 VDDA.n175 VDDA.n174 0.15675
R1696 VDDA.n176 VDDA.n175 0.15675
R1697 VDDA.n176 VDDA.n119 0.15675
R1698 VDDA.n181 VDDA.n119 0.15675
R1699 VDDA.n182 VDDA.n181 0.15675
R1700 VDDA.n183 VDDA.n182 0.15675
R1701 VDDA.n183 VDDA.n116 0.15675
R1702 VDDA.n116 VDDA.n115 0.15675
R1703 VDDA.n188 VDDA.n115 0.15675
R1704 VDDA.n189 VDDA.n188 0.15675
R1705 VDDA.n190 VDDA.n189 0.15675
R1706 VDDA.n191 VDDA.n190 0.15675
R1707 VDDA.n191 VDDA.n113 0.15675
R1708 VDDA.n113 VDDA.n112 0.15675
R1709 VDDA.n112 VDDA.n111 0.15675
R1710 VDDA.n111 VDDA.n93 0.15675
R1711 VDDA.n107 VDDA.n93 0.15675
R1712 VDDA.n107 VDDA.n106 0.15675
R1713 VDDA.n106 VDDA.n105 0.15675
R1714 VDDA.n105 VDDA.n96 0.15675
R1715 VDDA.n101 VDDA.n96 0.15675
R1716 VDDA.n101 VDDA.n100 0.15675
R1717 VDDA.n100 VDDA.n99 0.15675
R1718 VDDA.n99 VDDA.n58 0.15675
R1719 VDDA.n267 VDDA.n58 0.15675
R1720 VDDA.n268 VDDA.n267 0.15675
R1721 VDDA.n269 VDDA.n268 0.15675
R1722 VDDA.n283 VDDA.n282 0.15675
R1723 VDDA.n282 VDDA.n281 0.15675
R1724 VDDA.n281 VDDA.n275 0.15675
R1725 VDDA.n277 VDDA.n275 0.15675
R1726 VDDA.n277 VDDA.n276 0.15675
R1727 VDDA.n276 VDDA.n47 0.15675
R1728 VDDA.n369 VDDA.n47 0.15675
R1729 VDDA.n370 VDDA.n369 0.15675
R1730 VDDA.n372 VDDA.n44 0.15675
R1731 VDDA.n377 VDDA.n44 0.15675
R1732 VDDA.n378 VDDA.n377 0.15675
R1733 VDDA.n379 VDDA.n378 0.15675
R1734 VDDA.n379 VDDA.n40 0.15675
R1735 VDDA.n384 VDDA.n40 0.15675
R1736 VDDA.n385 VDDA.n384 0.15675
R1737 VDDA.n386 VDDA.n385 0.15675
R1738 VDDA.n386 VDDA.n36 0.15675
R1739 VDDA.n392 VDDA.n36 0.15675
R1740 VDDA.n393 VDDA.n392 0.15675
R1741 VDDA.n394 VDDA.n393 0.15675
R1742 VDDA.n394 VDDA.n24 0.15675
R1743 VDDA.n400 VDDA.n24 0.15675
R1744 VDDA.n401 VDDA.n400 0.15675
R1745 VDDA.n401 VDDA.n16 0.15675
R1746 VDDA.n481 VDDA.n16 0.15675
R1747 VDDA.n482 VDDA.n481 0.15675
R1748 VDDA.n483 VDDA.n482 0.15675
R1749 VDDA.n483 VDDA.n12 0.15675
R1750 VDDA.n488 VDDA.n12 0.15675
R1751 VDDA.n489 VDDA.n488 0.15675
R1752 VDDA.n490 VDDA.n489 0.15675
R1753 VDDA.n490 VDDA.n10 0.15675
R1754 VDDA.n494 VDDA.n10 0.15675
R1755 VDDA.n495 VDDA.n494 0.15675
R1756 VDDA.n496 VDDA.n495 0.15675
R1757 VDDA.n496 VDDA.n6 0.15675
R1758 VDDA.n502 VDDA.n6 0.15675
R1759 VDDA.n503 VDDA.n502 0.15675
R1760 VDDA.n504 VDDA.n503 0.15675
R1761 VDDA.n504 VDDA.n4 0.15675
R1762 VDDA.n508 VDDA.n4 0.15675
R1763 VDDA.n509 VDDA.n508 0.15675
R1764 VDDA.n510 VDDA.n509 0.15675
R1765 VDDA.n510 VDDA.n0 0.15675
R1766 VDDA.n514 VDDA.n0 0.15675
R1767 VDDA VDDA.n514 0.1255
R1768 VDDA.n269 VDDA 0.122375
R1769 VDDA.n155 VDDA.n154 0.100307
R1770 VDDA.n154 VDDA.n153 0.09425
R1771 VDDA.n213 VDDA.n212 0.09425
R1772 VDDA.n220 VDDA.n219 0.09425
R1773 VDDA.n227 VDDA.n226 0.09425
R1774 VDDA.n234 VDDA.n233 0.09425
R1775 VDDA.n244 VDDA.n243 0.09425
R1776 VDDA.n371 VDDA.n370 0.078625
R1777 VDDA.n372 VDDA.n371 0.078625
R1778 VDDA.n212 VDDA.n211 0.063
R1779 VDDA.n219 VDDA.n218 0.063
R1780 VDDA.n226 VDDA.n225 0.063
R1781 VDDA.n233 VDDA.n232 0.063
R1782 VDDA.n244 VDDA.n66 0.063
R1783 VDDA.n271 VDDA 0.0505
R1784 opamp_cell_4_0.VOUT pfd_8_0.opamp_out.n6 3993.6
R1785 pfd_8_0.opamp_out.n6 pfd_8_0.opamp_out.n4 823.75
R1786 pfd_8_0.opamp_out.n6 pfd_8_0.opamp_out.n5 753.326
R1787 pfd_8_0.opamp_out.n13 pfd_8_0.opamp_out.n12 424.447
R1788 pfd_8_0.opamp_out.n13 pfd_8_0.opamp_out.n11 354.048
R1789 pfd_8_0.opamp_out.n9 pfd_8_0.opamp_out.n8 313
R1790 pfd_8_0.opamp_out.t14 pfd_8_0.opamp_out.n0 297.233
R1791 pfd_8_0.opamp_out.n1 pfd_8_0.opamp_out.t14 297.233
R1792 pfd_8_0.opamp_out.n2 pfd_8_0.opamp_out.t13 297.233
R1793 pfd_8_0.opamp_out.n5 pfd_8_0.opamp_out.t2 281.596
R1794 pfd_8_0.opamp_out.n9 pfd_8_0.opamp_out.n7 242.601
R1795 pfd_8_0.opamp_out.n10 pfd_8_0.opamp_out.n9 220.8
R1796 pfd_8_0.opamp_out.n14 pfd_8_0.opamp_out.n13 220.8
R1797 pfd_8_0.opamp_out.n2 pfd_8_0.opamp_out.n1 216.9
R1798 pfd_8_0.opamp_out.n3 pfd_8_0.opamp_out.n0 216.9
R1799 charge_pump_cell_6_0.opamp_out pfd_8_0.opamp_out.n3 176.733
R1800 pfd_8_0.opamp_out.n5 pfd_8_0.opamp_out.t9 118.666
R1801 pfd_8_0.opamp_out.n1 pfd_8_0.opamp_out.t11 80.3338
R1802 pfd_8_0.opamp_out.t11 pfd_8_0.opamp_out.n0 80.3338
R1803 pfd_8_0.opamp_out.t12 pfd_8_0.opamp_out.n2 80.3338
R1804 pfd_8_0.opamp_out.n3 pfd_8_0.opamp_out.t12 80.3338
R1805 pfd_8_0.opamp_out.n4 pfd_8_0.opamp_out.t13 80.3338
R1806 pfd_8_0.opamp_out.n10 pfd_8_0.opamp_out.t15 70.0829
R1807 pfd_8_0.opamp_out.n15 pfd_8_0.opamp_out.n14 64.0005
R1808 pfd_8_0.opamp_out.n14 pfd_8_0.opamp_out.t10 63.6829
R1809 pfd_8_0.opamp_out.n15 pfd_8_0.opamp_out.n10 60.8005
R1810 pfd_8_0.opamp_out.n7 pfd_8_0.opamp_out.t1 60.0005
R1811 pfd_8_0.opamp_out.n7 pfd_8_0.opamp_out.t0 60.0005
R1812 pfd_8_0.opamp_out.n8 pfd_8_0.opamp_out.t4 60.0005
R1813 pfd_8_0.opamp_out.n8 pfd_8_0.opamp_out.t3 60.0005
R1814 pfd_8_0.opamp_out.n11 pfd_8_0.opamp_out.t5 49.2505
R1815 pfd_8_0.opamp_out.n11 pfd_8_0.opamp_out.t6 49.2505
R1816 pfd_8_0.opamp_out.n12 pfd_8_0.opamp_out.t8 49.2505
R1817 pfd_8_0.opamp_out.n12 pfd_8_0.opamp_out.t7 49.2505
R1818 pfd_8_0.opamp_out.n4 charge_pump_cell_6_0.opamp_out 16.0672
R1819 opamp_cell_4_0.VOUT pfd_8_0.opamp_out.n15 6.4005
R1820 a_6380_5710.n4 a_6380_5710.n0 427.647
R1821 a_6380_5710.n1 a_6380_5710.t6 321.334
R1822 a_6380_5710.n5 a_6380_5710.n4 210.601
R1823 a_6380_5710.n2 a_6380_5710.n1 208.868
R1824 a_6380_5710.n3 a_6380_5710.t0 174.056
R1825 a_6380_5710.n4 a_6380_5710.n3 152
R1826 a_6380_5710.n1 a_6380_5710.t7 112.468
R1827 a_6380_5710.n2 a_6380_5710.t2 112.468
R1828 a_6380_5710.n3 a_6380_5710.n2 61.5894
R1829 a_6380_5710.t3 a_6380_5710.n5 60.0005
R1830 a_6380_5710.n5 a_6380_5710.t1 60.0005
R1831 a_6380_5710.n0 a_6380_5710.t5 49.2505
R1832 a_6380_5710.n0 a_6380_5710.t4 49.2505
R1833 a_6500_6300.n7 a_6500_6300.n5 482.582
R1834 a_6500_6300.n10 a_6500_6300.t2 304.634
R1835 a_6500_6300.n3 a_6500_6300.t0 304.634
R1836 a_6500_6300.t4 a_6500_6300.n10 277.914
R1837 a_6500_6300.n3 a_6500_6300.t1 276.289
R1838 a_6500_6300.n8 a_6500_6300.n1 204.201
R1839 a_6500_6300.n4 a_6500_6300.n2 204.201
R1840 a_6500_6300.n9 a_6500_6300.n0 204.201
R1841 a_6500_6300.n7 a_6500_6300.n6 120.981
R1842 a_6500_6300.n8 a_6500_6300.n4 74.6672
R1843 a_6500_6300.n9 a_6500_6300.n8 74.6672
R1844 a_6500_6300.n1 a_6500_6300.t6 60.0005
R1845 a_6500_6300.n1 a_6500_6300.t8 60.0005
R1846 a_6500_6300.t1 a_6500_6300.n2 60.0005
R1847 a_6500_6300.n2 a_6500_6300.t5 60.0005
R1848 a_6500_6300.n0 a_6500_6300.t7 60.0005
R1849 a_6500_6300.n0 a_6500_6300.t3 60.0005
R1850 a_6500_6300.n8 a_6500_6300.n7 37.763
R1851 a_6500_6300.n5 a_6500_6300.t11 24.0005
R1852 a_6500_6300.n5 a_6500_6300.t9 24.0005
R1853 a_6500_6300.n6 a_6500_6300.t10 24.0005
R1854 a_6500_6300.n6 a_6500_6300.t12 24.0005
R1855 a_6500_6300.n4 a_6500_6300.n3 16.0005
R1856 a_6500_6300.n10 a_6500_6300.n9 16.0005
R1857 pfd_8_0.DOWN_PFD_b.t1 pfd_8_0.DOWN_PFD_b.n1 203.528
R1858 pfd_8_0.DOWN_PFD_b.n0 pfd_8_0.DOWN_PFD_b.t3 203.528
R1859 pfd_8_0.DOWN_PFD_b.n1 pfd_8_0.DOWN_PFD_b.t0 183.935
R1860 pfd_8_0.DOWN_PFD_b.n0 pfd_8_0.DOWN_PFD_b.t2 183.935
R1861 pfd_8_0.DOWN_PFD_b.n1 pfd_8_0.DOWN_PFD_b.n0 83.2005
R1862 pfd_8_0.DOWN_b.n0 pfd_8_0.DOWN_b.t5 1028.27
R1863 pfd_8_0.DOWN_b.n2 pfd_8_0.DOWN_b.n1 569.734
R1864 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.n0 465.933
R1865 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.t3 401.668
R1866 pfd_8_0.DOWN_b.n0 pfd_8_0.DOWN_b.t4 385.601
R1867 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.t2 385.601
R1868 pfd_8_0.DOWN_b.t1 pfd_8_0.DOWN_b.n2 211.847
R1869 pfd_8_0.DOWN_b.n2 pfd_8_0.DOWN_b.t0 173.055
R1870 pfd_8_0.QA_b.t4 pfd_8_0.QA_b.t6 1188.93
R1871 pfd_8_0.QA_b pfd_8_0.QA_b.n2 837.38
R1872 pfd_8_0.QA_b.t6 pfd_8_0.QA_b.t3 835.467
R1873 pfd_8_0.QA_b.n0 pfd_8_0.QA_b.t5 562.333
R1874 pfd_8_0.QA_b pfd_8_0.QA_b.n0 482
R1875 pfd_8_0.QA_b.n2 pfd_8_0.QA_b.n1 247.917
R1876 pfd_8_0.QA_b.n0 pfd_8_0.QA_b.t4 224.934
R1877 pfd_8_0.QA_b.n2 pfd_8_0.QA_b.t1 221.411
R1878 pfd_8_0.QA_b.n1 pfd_8_0.QA_b.t0 24.0005
R1879 pfd_8_0.QA_b.n1 pfd_8_0.QA_b.t2 24.0005
R1880 a_870_1400.t0 a_870_1400.t1 39.4005
R1881 opamp_cell_4_0.p_bias opamp_cell_4_0.p_bias.t8 918.318
R1882 opamp_cell_4_0.p_bias opamp_cell_4_0.p_bias.n11 540.801
R1883 opamp_cell_4_0.p_bias.n8 opamp_cell_4_0.p_bias.t9 377.567
R1884 opamp_cell_4_0.p_bias.n3 opamp_cell_4_0.p_bias.t12 377.567
R1885 opamp_cell_4_0.p_bias.n9 opamp_cell_4_0.p_bias.n8 257.067
R1886 opamp_cell_4_0.p_bias.n7 opamp_cell_4_0.p_bias.n6 257.067
R1887 opamp_cell_4_0.p_bias.n4 opamp_cell_4_0.p_bias.n3 257.067
R1888 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n0 154.321
R1889 opamp_cell_4_0.p_bias.n2 opamp_cell_4_0.p_bias.n1 154.321
R1890 opamp_cell_4_0.p_bias.n5 opamp_cell_4_0.p_bias.n2 152
R1891 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n10 152
R1892 opamp_cell_4_0.p_bias.n8 opamp_cell_4_0.p_bias.t11 120.501
R1893 opamp_cell_4_0.p_bias.n9 opamp_cell_4_0.p_bias.t6 120.501
R1894 opamp_cell_4_0.p_bias.n7 opamp_cell_4_0.p_bias.t2 120.501
R1895 opamp_cell_4_0.p_bias.n6 opamp_cell_4_0.p_bias.t4 120.501
R1896 opamp_cell_4_0.p_bias.n3 opamp_cell_4_0.p_bias.t10 120.501
R1897 opamp_cell_4_0.p_bias.n4 opamp_cell_4_0.p_bias.t0 120.501
R1898 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n2 115.201
R1899 opamp_cell_4_0.p_bias.n10 opamp_cell_4_0.p_bias.n9 85.6894
R1900 opamp_cell_4_0.p_bias.n10 opamp_cell_4_0.p_bias.n7 85.6894
R1901 opamp_cell_4_0.p_bias.n6 opamp_cell_4_0.p_bias.n5 85.6894
R1902 opamp_cell_4_0.p_bias.n5 opamp_cell_4_0.p_bias.n4 85.6894
R1903 opamp_cell_4_0.p_bias.n0 opamp_cell_4_0.p_bias.t3 19.7005
R1904 opamp_cell_4_0.p_bias.n0 opamp_cell_4_0.p_bias.t7 19.7005
R1905 opamp_cell_4_0.p_bias.n1 opamp_cell_4_0.p_bias.t1 19.7005
R1906 opamp_cell_4_0.p_bias.n1 opamp_cell_4_0.p_bias.t5 19.7005
R1907 a_6150_5090.n8 a_6150_5090.n6 522.322
R1908 a_6150_5090.n3 a_6150_5090.t6 384.967
R1909 a_6150_5090.n0 a_6150_5090.t9 384.967
R1910 a_6150_5090.n3 a_6150_5090.t8 379.166
R1911 a_6150_5090.t10 a_6150_5090.n0 376.56
R1912 a_6150_5090.n5 a_6150_5090.n1 315.647
R1913 a_6150_5090.n4 a_6150_5090.n2 315.647
R1914 a_6150_5090.n11 a_6150_5090.n10 314.502
R1915 a_6150_5090.n8 a_6150_5090.n7 160.721
R1916 a_6150_5090.n5 a_6150_5090.n4 83.2005
R1917 a_6150_5090.n1 a_6150_5090.t0 49.2505
R1918 a_6150_5090.n1 a_6150_5090.t12 49.2505
R1919 a_6150_5090.n2 a_6150_5090.t11 49.2505
R1920 a_6150_5090.n2 a_6150_5090.t7 49.2505
R1921 a_6150_5090.t10 a_6150_5090.n11 49.2505
R1922 a_6150_5090.n11 a_6150_5090.t5 49.2505
R1923 a_6150_5090.n10 a_6150_5090.n9 42.6672
R1924 a_6150_5090.n9 a_6150_5090.n8 37.763
R1925 a_6150_5090.n9 a_6150_5090.n5 23.4672
R1926 a_6150_5090.n6 a_6150_5090.t1 19.7005
R1927 a_6150_5090.n6 a_6150_5090.t3 19.7005
R1928 a_6150_5090.n7 a_6150_5090.t2 19.7005
R1929 a_6150_5090.n7 a_6150_5090.t4 19.7005
R1930 a_6150_5090.n4 a_6150_5090.n3 16.0005
R1931 a_6150_5090.n10 a_6150_5090.n0 16.0005
R1932 pfd_8_0.DOWN.t3 pfd_8_0.DOWN.n0 605.311
R1933 charge_pump_cell_6_0.DOWN pfd_8_0.DOWN.t3 398.807
R1934 pfd_8_0.DOWN.n0 pfd_8_0.DOWN.t0 240.327
R1935 pfd_8_0.DOWN.n0 pfd_8_0.DOWN.t1 148.736
R1936 charge_pump_cell_6_0.DOWN pfd_8_0.DOWN.t2 12.0821
R1937 pfd_8_0.UP_input.n1 pfd_8_0.UP_input.t5 326.658
R1938 pfd_8_0.UP_input.n3 pfd_8_0.UP_input.t4 297.233
R1939 pfd_8_0.UP_input.t3 pfd_8_0.UP_input.n4 297.233
R1940 pfd_8_0.UP_input.n2 pfd_8_0.UP_input.n0 257.067
R1941 pfd_8_0.UP_input.t0 pfd_8_0.UP_input.n7 241.928
R1942 pfd_8_0.UP_input.n5 pfd_8_0.UP_input.n0 226.942
R1943 pfd_8_0.UP_input.n2 pfd_8_0.UP_input.n1 226.942
R1944 pfd_8_0.UP_input.n6 pfd_8_0.UP_input.n5 225.417
R1945 pfd_8_0.UP_input.n4 pfd_8_0.UP_input.n3 216.9
R1946 pfd_8_0.UP_input.n6 pfd_8_0.UP_input.t1 209.928
R1947 pfd_8_0.UP_input.n7 pfd_8_0.UP_input.t2 145.536
R1948 pfd_8_0.UP_input.n7 pfd_8_0.UP_input.n6 144
R1949 pfd_8_0.UP_input.n1 pfd_8_0.UP_input.t4 92.3838
R1950 pfd_8_0.UP_input.n5 pfd_8_0.UP_input.t3 92.3838
R1951 pfd_8_0.UP_input.n3 pfd_8_0.UP_input.t6 80.3338
R1952 pfd_8_0.UP_input.t6 pfd_8_0.UP_input.n2 80.3338
R1953 pfd_8_0.UP_input.n4 pfd_8_0.UP_input.t7 80.3338
R1954 pfd_8_0.UP_input.t7 pfd_8_0.UP_input.n0 80.3338
R1955 V_OUT.n2 V_OUT.n1 2008.33
R1956 V_OUT V_OUT.n8 1614.79
R1957 V_OUT V_OUT.n2 618.567
R1958 V_OUT.n0 V_OUT.t6 401.668
R1959 V_OUT.n2 V_OUT.n0 369.534
R1960 V_OUT.n1 V_OUT.t8 321.334
R1961 V_OUT.n5 V_OUT.n4 242.903
R1962 V_OUT.n0 V_OUT.t7 192.8
R1963 V_OUT.n5 V_OUT.n3 172.502
R1964 V_OUT.n8 V_OUT.n7 113.178
R1965 V_OUT.n1 V_OUT.t9 112.468
R1966 V_OUT.n7 V_OUT.n6 106.662
R1967 V_OUT.n3 V_OUT.t2 24.6255
R1968 V_OUT.n3 V_OUT.t1 24.6255
R1969 V_OUT.n4 V_OUT.t0 24.6255
R1970 V_OUT.n4 V_OUT.t3 24.6255
R1971 V_OUT.n7 V_OUT.n5 19.2005
R1972 V_OUT.n6 V_OUT.t4 15.0005
R1973 V_OUT.n6 V_OUT.t5 15.0005
R1974 V_OUT.n8 V_OUT 0.063
R1975 pfd_8_0.before_Reset.n1 pfd_8_0.before_Reset.n0 481.334
R1976 pfd_8_0.before_Reset.n0 pfd_8_0.before_Reset.t4 465.933
R1977 pfd_8_0.before_Reset.n0 pfd_8_0.before_Reset.t3 321.334
R1978 pfd_8_0.before_Reset.n2 pfd_8_0.before_Reset.n1 226.889
R1979 pfd_8_0.before_Reset.n1 pfd_8_0.before_Reset.t2 172.458
R1980 pfd_8_0.before_Reset.n2 pfd_8_0.before_Reset.t1 19.7005
R1981 pfd_8_0.before_Reset.t0 pfd_8_0.before_Reset.n2 19.7005
R1982 a_2350_1400.t0 a_2350_1400.n2 500.086
R1983 a_2350_1400.n1 a_2350_1400.n0 473.334
R1984 a_2350_1400.n0 a_2350_1400.t3 465.933
R1985 a_2350_1400.t0 a_2350_1400.n2 461.389
R1986 a_2350_1400.n0 a_2350_1400.t2 321.334
R1987 a_2350_1400.n1 a_2350_1400.t1 177.577
R1988 a_2350_1400.n2 a_2350_1400.n1 48.3899
R1989 F_REF.n0 F_REF.t0 514.134
R1990 F_REF.n0 F_REF.t1 273.134
R1991 F_REF F_REF.n0 216.9
R1992 a_n30_1400.t0 a_n30_1400.t1 39.4005
R1993 a_6670_5090.t1 a_6670_5090.n6 1112.76
R1994 a_6670_5090.n3 a_6670_5090.n2 416.863
R1995 a_6670_5090.n2 a_6670_5090.n1 366.848
R1996 a_6670_5090.n2 a_6670_5090.n0 271.401
R1997 a_6670_5090.n3 a_6670_5090.t5 208.868
R1998 a_6670_5090.n6 a_6670_5090.t7 208.868
R1999 a_6670_5090.n5 a_6670_5090.t6 208.868
R2000 a_6670_5090.n4 a_6670_5090.t8 208.868
R2001 a_6670_5090.n6 a_6670_5090.n5 208.868
R2002 a_6670_5090.n5 a_6670_5090.n4 208.868
R2003 a_6670_5090.n4 a_6670_5090.n3 193.804
R2004 a_6670_5090.n0 a_6670_5090.t3 60.0005
R2005 a_6670_5090.n0 a_6670_5090.t2 60.0005
R2006 a_6670_5090.n1 a_6670_5090.t4 49.2505
R2007 a_6670_5090.n1 a_6670_5090.t0 49.2505
R2008 pfd_8_0.QA.t5 pfd_8_0.QA.t7 835.467
R2009 pfd_8_0.QA.n2 pfd_8_0.QA.t4 517.347
R2010 pfd_8_0.QA.n0 pfd_8_0.QA.t8 465.933
R2011 pfd_8_0.QA.n1 pfd_8_0.QA.n0 454.031
R2012 pfd_8_0.QA.n1 pfd_8_0.QA.t5 394.267
R2013 pfd_8_0.QA.n0 pfd_8_0.QA.t6 321.334
R2014 pfd_8_0.QA.n4 pfd_8_0.QA.n3 244.715
R2015 pfd_8_0.QA.n2 pfd_8_0.QA.t3 228.148
R2016 pfd_8_0.QA.n4 pfd_8_0.QA.t0 221.411
R2017 pfd_8_0.QA.n5 pfd_8_0.QA.n2 216
R2018 pfd_8_0.QA.n5 pfd_8_0.QA.n4 201.573
R2019 pfd_8_0.QA pfd_8_0.QA.n5 60.8005
R2020 pfd_8_0.QA pfd_8_0.QA.n1 56.1505
R2021 pfd_8_0.QA.n3 pfd_8_0.QA.t2 24.0005
R2022 pfd_8_0.QA.n3 pfd_8_0.QA.t1 24.0005
R2023 I_IN.n2 I_IN.n1 1269.42
R2024 I_IN I_IN.n5 589.356
R2025 I_IN.n2 I_IN.t2 275.325
R2026 I_IN.n4 I_IN.n3 248.4
R2027 I_IN.n5 I_IN.t1 238.892
R2028 I_IN I_IN.n4 214.4
R2029 I_IN.n5 I_IN.t0 161.371
R2030 I_IN.n1 I_IN.t6 151.792
R2031 I_IN.n3 I_IN.t4 140.583
R2032 I_IN.n3 I_IN.t2 140.583
R2033 I_IN.n4 I_IN.n0 98.6614
R2034 I_IN.t4 I_IN.n2 80.3338
R2035 I_IN.n1 I_IN.t7 44.2902
R2036 I_IN.n0 I_IN.t5 15.0005
R2037 I_IN.n0 I_IN.t3 15.0005
R2038 pfd_8_0.DOWN_input pfd_8_0.DOWN_input.n1 539.794
R2039 pfd_8_0.DOWN_input.t3 pfd_8_0.DOWN_input.t4 377.567
R2040 pfd_8_0.DOWN_input.n0 pfd_8_0.DOWN_input.t5 326.658
R2041 pfd_8_0.DOWN_input.n2 pfd_8_0.DOWN_input.t0 229.127
R2042 pfd_8_0.DOWN_input.n1 pfd_8_0.DOWN_input.n0 196.817
R2043 pfd_8_0.DOWN_input.n2 pfd_8_0.DOWN_input.t2 158.335
R2044 pfd_8_0.DOWN_input.n3 pfd_8_0.DOWN_input.t1 158.335
R2045 pfd_8_0.DOWN_input.n3 pfd_8_0.DOWN_input.n2 124.8
R2046 pfd_8_0.DOWN_input.t4 pfd_8_0.DOWN_input.n0 92.3838
R2047 pfd_8_0.DOWN_input.n1 pfd_8_0.DOWN_input.t3 92.3838
R2048 pfd_8_0.DOWN_input pfd_8_0.DOWN_input.n3 6.4005
R2049 pfd_8_0.QB.t4 pfd_8_0.QB.t3 835.467
R2050 pfd_8_0.QB.n1 pfd_8_0.QB.t4 564.496
R2051 pfd_8_0.QB.n2 pfd_8_0.QB.t5 517.347
R2052 pfd_8_0.QB.n0 pfd_8_0.QB.t7 514.134
R2053 pfd_8_0.QB.n1 pfd_8_0.QB.n0 455.219
R2054 pfd_8_0.QB.n5 pfd_8_0.QB.n2 363.2
R2055 pfd_8_0.QB.n0 pfd_8_0.QB.t8 273.134
R2056 pfd_8_0.QB.n4 pfd_8_0.QB.n3 244.716
R2057 pfd_8_0.QB.n2 pfd_8_0.QB.t6 228.148
R2058 pfd_8_0.QB.n4 pfd_8_0.QB.t0 221.411
R2059 pfd_8_0.QB.n5 pfd_8_0.QB.n4 54.3734
R2060 pfd_8_0.QB pfd_8_0.QB.n1 26.7568
R2061 pfd_8_0.QB.n3 pfd_8_0.QB.t2 24.0005
R2062 pfd_8_0.QB.n3 pfd_8_0.QB.t1 24.0005
R2063 pfd_8_0.QB pfd_8_0.QB.n5 6.4005
R2064 a_1910_2020.t0 a_1910_2020.t1 48.0005
R2065 pfd_8_0.UP_PFD_b.n0 pfd_8_0.UP_PFD_b.t2 441.834
R2066 pfd_8_0.UP_PFD_b.n0 pfd_8_0.UP_PFD_b.t3 313.3
R2067 pfd_8_0.UP_PFD_b.n1 pfd_8_0.UP_PFD_b.n0 235.201
R2068 pfd_8_0.UP_PFD_b.t0 pfd_8_0.UP_PFD_b.n1 219.528
R2069 pfd_8_0.UP_PFD_b.n1 pfd_8_0.UP_PFD_b.t1 167.935
R2070 pfd_8_0.UP.n0 pfd_8_0.UP.t5 1205
R2071 pfd_8_0.UP.n2 pfd_8_0.UP.t4 522.168
R2072 pfd_8_0.UP.n1 pfd_8_0.UP.n0 441.834
R2073 pfd_8_0.UP.n3 pfd_8_0.UP.n2 235.201
R2074 pfd_8_0.UP.t0 pfd_8_0.UP.n3 229.127
R2075 pfd_8_0.UP.n1 pfd_8_0.UP.t3 217.905
R2076 pfd_8_0.UP.n0 pfd_8_0.UP.t2 208.868
R2077 pfd_8_0.UP.n3 pfd_8_0.UP.t1 158.335
R2078 pfd_8_0.UP.n2 pfd_8_0.UP.n1 15.063
R2079 a_9540_3974.t1 a_9540_3974.t0 323.964
R2080 pfd_8_0.E.n4 pfd_8_0.E.n0 1319.38
R2081 pfd_8_0.E.n0 pfd_8_0.E.t3 562.333
R2082 pfd_8_0.E.n2 pfd_8_0.E.t5 388.813
R2083 pfd_8_0.E.n2 pfd_8_0.E.t4 356.68
R2084 pfd_8_0.E.n3 pfd_8_0.E.n2 232
R2085 pfd_8_0.E.n0 pfd_8_0.E.t6 224.934
R2086 pfd_8_0.E.t2 pfd_8_0.E.n4 221.411
R2087 pfd_8_0.E.n3 pfd_8_0.E.n1 157.278
R2088 pfd_8_0.E.n4 pfd_8_0.E.n3 90.64
R2089 pfd_8_0.E.n1 pfd_8_0.E.t0 24.0005
R2090 pfd_8_0.E.n1 pfd_8_0.E.t1 24.0005
R2091 pfd_8_0.E_b.n0 pfd_8_0.E_b.t4 517.347
R2092 pfd_8_0.E_b.n2 pfd_8_0.E_b.n0 417.574
R2093 pfd_8_0.E_b.n2 pfd_8_0.E_b.n1 244.716
R2094 pfd_8_0.E_b.n0 pfd_8_0.E_b.t3 228.148
R2095 pfd_8_0.E_b.t1 pfd_8_0.E_b.n2 221.411
R2096 pfd_8_0.E_b.n1 pfd_8_0.E_b.t0 24.0005
R2097 pfd_8_0.E_b.n1 pfd_8_0.E_b.t2 24.0005
R2098 a_1390_1400.t0 a_1390_1400.t1 39.4005
R2099 pfd_8_0.QB_b.t6 pfd_8_0.QB_b.t4 1188.93
R2100 pfd_8_0.QB_b pfd_8_0.QB_b.n2 899.734
R2101 pfd_8_0.QB_b.t4 pfd_8_0.QB_b.t3 835.467
R2102 pfd_8_0.QB_b.n2 pfd_8_0.QB_b.t5 562.333
R2103 pfd_8_0.QB_b pfd_8_0.QB_b.n1 419.647
R2104 pfd_8_0.QB_b.n1 pfd_8_0.QB_b.n0 247.917
R2105 pfd_8_0.QB_b.n2 pfd_8_0.QB_b.t6 224.934
R2106 pfd_8_0.QB_b.n1 pfd_8_0.QB_b.t0 221.411
R2107 pfd_8_0.QB_b.n0 pfd_8_0.QB_b.t1 24.0005
R2108 pfd_8_0.QB_b.n0 pfd_8_0.QB_b.t2 24.0005
R2109 a_870_640.t0 a_870_640.t1 39.4005
R2110 a_2530_190.t0 a_2530_190.n2 500.086
R2111 a_2530_190.n0 a_2530_190.t2 465.933
R2112 a_2530_190.t0 a_2530_190.n2 461.389
R2113 a_2530_190.n1 a_2530_190.n0 392.623
R2114 a_2530_190.n0 a_2530_190.t3 321.334
R2115 a_2530_190.n1 a_2530_190.t1 177.577
R2116 a_2530_190.n2 a_2530_190.n1 48.3899
R2117 a_2200_190.t0 a_2200_190.n2 500.086
R2118 a_2200_190.n1 a_2200_190.n0 473.334
R2119 a_2200_190.n0 a_2200_190.t2 465.933
R2120 a_2200_190.t0 a_2200_190.n2 461.389
R2121 a_2200_190.n0 a_2200_190.t3 321.334
R2122 a_2200_190.n1 a_2200_190.t1 177.577
R2123 a_2200_190.n2 a_2200_190.n1 48.3898
R2124 pfd_8_0.F.n4 pfd_8_0.F.n0 1319.38
R2125 pfd_8_0.F.n0 pfd_8_0.F.t3 562.333
R2126 pfd_8_0.F.n2 pfd_8_0.F.t5 388.813
R2127 pfd_8_0.F.n2 pfd_8_0.F.t6 356.68
R2128 pfd_8_0.F.n3 pfd_8_0.F.n2 232
R2129 pfd_8_0.F.n0 pfd_8_0.F.t4 224.934
R2130 pfd_8_0.F.t0 pfd_8_0.F.n4 221.411
R2131 pfd_8_0.F.n3 pfd_8_0.F.n1 157.278
R2132 pfd_8_0.F.n4 pfd_8_0.F.n3 90.64
R2133 pfd_8_0.F.n1 pfd_8_0.F.t2 24.0005
R2134 pfd_8_0.F.n1 pfd_8_0.F.t1 24.0005
R2135 charge_pump_cell_6_0.UP_b pfd_8_0.UP_b.n1 485.846
R2136 pfd_8_0.UP_b.n1 pfd_8_0.UP_b.n0 409.067
R2137 pfd_8_0.UP_b.n1 pfd_8_0.UP_b.t3 369.534
R2138 pfd_8_0.UP_b.n0 pfd_8_0.UP_b.t1 209.928
R2139 pfd_8_0.UP_b.n0 pfd_8_0.UP_b.t2 177.536
R2140 charge_pump_cell_6_0.UP_b pfd_8_0.UP_b.t0 12.0774
R2141 pfd_8_0.F_b.n0 pfd_8_0.F_b.t3 517.347
R2142 pfd_8_0.F_b.n2 pfd_8_0.F_b.n0 417.574
R2143 pfd_8_0.F_b.n2 pfd_8_0.F_b.n1 244.716
R2144 pfd_8_0.F_b.n0 pfd_8_0.F_b.t4 228.148
R2145 pfd_8_0.F_b.t0 pfd_8_0.F_b.n2 221.411
R2146 pfd_8_0.F_b.n1 pfd_8_0.F_b.t2 24.0005
R2147 pfd_8_0.F_b.n1 pfd_8_0.F_b.t1 24.0005
R2148 a_1390_640.t0 a_1390_640.t1 39.4005
R2149 a_490_640.t0 a_490_640.t1 39.4005
R2150 opamp_cell_4_0.VIN+ opamp_cell_4_0.VIN+.n7 933.13
R2151 opamp_cell_4_0.VIN+.n0 opamp_cell_4_0.VIN+.t8 377.567
R2152 opamp_cell_4_0.VIN+.n1 opamp_cell_4_0.VIN+.t9 297.233
R2153 opamp_cell_4_0.VIN+.n2 opamp_cell_4_0.VIN+.n1 243.44
R2154 opamp_cell_4_0.VIN+.n2 opamp_cell_4_0.VIN+.n0 224.496
R2155 opamp_cell_4_0.VIN+.n0 opamp_cell_4_0.VIN+.t7 216.9
R2156 opamp_cell_4_0.VIN+.n6 opamp_cell_4_0.VIN+.n4 196.262
R2157 opamp_cell_4_0.VIN+.n7 opamp_cell_4_0.VIN+.n3 172.502
R2158 opamp_cell_4_0.VIN+.n6 opamp_cell_4_0.VIN+.n5 172.5
R2159 opamp_cell_4_0.VIN+.n1 opamp_cell_4_0.VIN+.t6 136.567
R2160 opamp_cell_4_0.VIN+.n7 opamp_cell_4_0.VIN+.n6 70.4005
R2161 opamp_cell_4_0.VIN+.n3 opamp_cell_4_0.VIN+.t2 24.6255
R2162 opamp_cell_4_0.VIN+.n3 opamp_cell_4_0.VIN+.t1 24.6255
R2163 opamp_cell_4_0.VIN+.n5 opamp_cell_4_0.VIN+.t0 24.6255
R2164 opamp_cell_4_0.VIN+.n5 opamp_cell_4_0.VIN+.t3 24.6255
R2165 opamp_cell_4_0.VIN+.n4 opamp_cell_4_0.VIN+.t5 15.0005
R2166 opamp_cell_4_0.VIN+.n4 opamp_cell_4_0.VIN+.t4 15.0005
R2167 opamp_cell_4_0.VIN+ opamp_cell_4_0.VIN+.n2 3.438
R2168 a_490_1400.t0 a_490_1400.t1 39.4005
R2169 pfd_8_0.Reset.n1 pfd_8_0.Reset.t3 562.333
R2170 pfd_8_0.Reset.n2 pfd_8_0.Reset.n1 480.45
R2171 pfd_8_0.Reset.n0 pfd_8_0.Reset.t4 417.733
R2172 pfd_8_0.Reset.n0 pfd_8_0.Reset.t5 369.534
R2173 pfd_8_0.Reset.n3 pfd_8_0.Reset.n2 328.733
R2174 pfd_8_0.Reset.t1 pfd_8_0.Reset.n3 288.37
R2175 pfd_8_0.Reset.n1 pfd_8_0.Reset.t2 224.934
R2176 pfd_8_0.Reset.n3 pfd_8_0.Reset.t0 177.577
R2177 pfd_8_0.Reset.n2 pfd_8_0.Reset.n0 176.733
R2178 a_1870_190.t0 a_1870_190.n2 500.086
R2179 a_1870_190.n1 a_1870_190.n0 473.334
R2180 a_1870_190.n0 a_1870_190.t2 465.933
R2181 a_1870_190.t0 a_1870_190.n2 461.389
R2182 a_1870_190.n0 a_1870_190.t3 321.334
R2183 a_1870_190.n1 a_1870_190.t1 177.577
R2184 a_1870_190.n2 a_1870_190.n1 48.3898
R2185 a_9540_6900.t1 a_9540_6900.t0 245.883
R2186 a_n30_640.t0 a_n30_640.t1 39.4005
R2187 F_VCO.n0 F_VCO.t0 514.134
R2188 F_VCO.n0 F_VCO.t1 273.134
R2189 F_VCO F_VCO.n0 216.9
C0 opamp_cell_4_0.p_bias opamp_cell_4_0.VIN+ 0.498662f
C1 I_IN opamp_cell_4_0.VIN+ 0.544835f
C2 VDDA opamp_cell_4_0.VIN+ 1.06587f
C3 pfd_8_0.QB_b pfd_8_0.QB 0.388258f
C4 I_IN pfd_8_0.DOWN_input 0.581394f
C5 VDDA pfd_8_0.DOWN_input 0.168412f
C6 V_OUT opamp_cell_4_0.VIN+ 1.18544f
C7 pfd_8_0.QB_b VDDA 0.511838f
C8 pfd_8_0.DOWN_input V_OUT 0.406052f
C9 pfd_8_0.QB VDDA 2.74984f
C10 F_REF VDDA 0.098433f
C11 VDDA opamp_cell_4_0.p_bias 3.3163f
C12 I_IN VDDA 0.452819f
C13 pfd_8_0.QA_b F_REF 0.027208f
C14 pfd_8_0.QA_b VDDA 0.52066f
C15 opamp_cell_4_0.p_bias V_OUT 0.049138f
C16 F_VCO pfd_8_0.QB_b 0.027208f
C17 pfd_8_0.QA pfd_8_0.QB 0.074487f
C18 pfd_8_0.QA F_REF 0.056f
C19 VDDA V_OUT 1.44907f
C20 pfd_8_0.DOWN_input opamp_cell_4_0.VIN+ 0.132099f
C21 F_VCO pfd_8_0.QB 0.056153f
C22 pfd_8_0.QA VDDA 0.550605f
C23 F_VCO VDDA 0.098386f
C24 pfd_8_0.QA_b pfd_8_0.QA 0.422694f
C25 I_IN GNDA 3.05272f
C26 F_VCO GNDA 0.277756f
C27 F_REF GNDA 0.277756f
C28 V_OUT GNDA 5.87015f
C29 VDDA GNDA 65.92424f
C30 pfd_8_0.DOWN_input GNDA 3.21943f
C31 pfd_8_0.QB_b GNDA 1.06334f
C32 pfd_8_0.QB GNDA 1.3083f
C33 pfd_8_0.QA GNDA 3.10074f
C34 pfd_8_0.QA_b GNDA 1.05138f
C35 opamp_cell_4_0.VIN+ GNDA 2.71146f
C36 opamp_cell_4_0.p_bias GNDA 3.153184f
C37 pfd_8_0.QB.t7 GNDA 0.066708f
C38 pfd_8_0.QB.t8 GNDA 0.031333f
C39 pfd_8_0.QB.n0 GNDA 0.096363f
C40 pfd_8_0.QB.t3 GNDA 0.066708f
C41 pfd_8_0.QB.t4 GNDA 0.100569f
C42 pfd_8_0.QB.n1 GNDA 1.20598f
C43 pfd_8_0.QB.t5 GNDA 0.067367f
C44 pfd_8_0.QB.t6 GNDA 0.029539f
C45 pfd_8_0.QB.n2 GNDA 0.170164f
C46 pfd_8_0.QB.t0 GNDA 0.14186f
C47 pfd_8_0.QB.t2 GNDA 0.026953f
C48 pfd_8_0.QB.t1 GNDA 0.026953f
C49 pfd_8_0.QB.n3 GNDA 0.143916f
C50 pfd_8_0.QB.n4 GNDA 0.255686f
C51 pfd_8_0.QB.n5 GNDA 0.218372f
C52 pfd_8_0.UP_input.t2 GNDA 0.019943f
C53 pfd_8_0.UP_input.t1 GNDA 0.043912f
C54 pfd_8_0.UP_input.n0 GNDA 0.022544f
C55 pfd_8_0.UP_input.t7 GNDA 0.024945f
C56 pfd_8_0.UP_input.t4 GNDA 0.042895f
C57 pfd_8_0.UP_input.t5 GNDA 1.97861f
C58 pfd_8_0.UP_input.n1 GNDA 0.043722f
C59 pfd_8_0.UP_input.n2 GNDA 0.022544f
C60 pfd_8_0.UP_input.t6 GNDA 0.024945f
C61 pfd_8_0.UP_input.n3 GNDA 0.030069f
C62 pfd_8_0.UP_input.n4 GNDA 0.030069f
C63 pfd_8_0.UP_input.t3 GNDA 0.042895f
C64 pfd_8_0.UP_input.n5 GNDA 0.039471f
C65 pfd_8_0.UP_input.n6 GNDA 0.22578f
C66 pfd_8_0.UP_input.n7 GNDA 0.059297f
C67 pfd_8_0.UP_input.t0 GNDA 0.048355f
C68 a_6150_5090.t9 GNDA 0.030769f
C69 a_6150_5090.n0 GNDA 0.124795f
C70 a_6150_5090.t5 GNDA 0.020325f
C71 a_6150_5090.t0 GNDA 0.020325f
C72 a_6150_5090.t12 GNDA 0.020325f
C73 a_6150_5090.n1 GNDA 0.044943f
C74 a_6150_5090.t11 GNDA 0.020325f
C75 a_6150_5090.t7 GNDA 0.020325f
C76 a_6150_5090.n2 GNDA 0.044943f
C77 a_6150_5090.t8 GNDA 0.077457f
C78 a_6150_5090.t6 GNDA 0.030769f
C79 a_6150_5090.n3 GNDA 0.097952f
C80 a_6150_5090.n4 GNDA 0.087903f
C81 a_6150_5090.n5 GNDA 0.089425f
C82 a_6150_5090.t1 GNDA 0.050813f
C83 a_6150_5090.t3 GNDA 0.050813f
C84 a_6150_5090.n6 GNDA 0.295522f
C85 a_6150_5090.t2 GNDA 0.050813f
C86 a_6150_5090.t4 GNDA 0.050813f
C87 a_6150_5090.n7 GNDA 0.144587f
C88 a_6150_5090.n8 GNDA 0.360746f
C89 a_6150_5090.n9 GNDA 0.13437f
C90 a_6150_5090.n10 GNDA 0.085474f
C91 a_6150_5090.n11 GNDA 0.045257f
C92 a_6150_5090.t10 GNDA 0.100208f
C93 opamp_cell_4_0.p_bias.t8 GNDA 1.892f
C94 opamp_cell_4_0.p_bias.t3 GNDA 0.022409f
C95 opamp_cell_4_0.p_bias.t7 GNDA 0.022409f
C96 opamp_cell_4_0.p_bias.n0 GNDA 0.061525f
C97 opamp_cell_4_0.p_bias.t1 GNDA 0.022409f
C98 opamp_cell_4_0.p_bias.t5 GNDA 0.022409f
C99 opamp_cell_4_0.p_bias.n1 GNDA 0.061525f
C100 opamp_cell_4_0.p_bias.n2 GNDA 0.07795f
C101 opamp_cell_4_0.p_bias.t2 GNDA 0.061849f
C102 opamp_cell_4_0.p_bias.t4 GNDA 0.061849f
C103 opamp_cell_4_0.p_bias.t0 GNDA 0.061849f
C104 opamp_cell_4_0.p_bias.t10 GNDA 0.061849f
C105 opamp_cell_4_0.p_bias.t12 GNDA 0.085041f
C106 opamp_cell_4_0.p_bias.n3 GNDA 0.047622f
C107 opamp_cell_4_0.p_bias.n4 GNDA 0.033793f
C108 opamp_cell_4_0.p_bias.n5 GNDA 0.014521f
C109 opamp_cell_4_0.p_bias.n6 GNDA 0.033793f
C110 opamp_cell_4_0.p_bias.n7 GNDA 0.033793f
C111 opamp_cell_4_0.p_bias.t6 GNDA 0.061849f
C112 opamp_cell_4_0.p_bias.t11 GNDA 0.061849f
C113 opamp_cell_4_0.p_bias.t9 GNDA 0.085041f
C114 opamp_cell_4_0.p_bias.n8 GNDA 0.047622f
C115 opamp_cell_4_0.p_bias.n9 GNDA 0.033793f
C116 opamp_cell_4_0.p_bias.n10 GNDA 0.014521f
C117 opamp_cell_4_0.p_bias.n11 GNDA 0.137263f
C118 pfd_8_0.opamp_out.t13 GNDA 0.016624f
C119 pfd_8_0.opamp_out.n0 GNDA 0.012184f
C120 pfd_8_0.opamp_out.t14 GNDA 0.02314f
C121 pfd_8_0.opamp_out.t11 GNDA 0.010108f
C122 pfd_8_0.opamp_out.n1 GNDA 0.012184f
C123 pfd_8_0.opamp_out.n2 GNDA 0.012184f
C124 pfd_8_0.opamp_out.t12 GNDA 0.010108f
C125 pfd_8_0.opamp_out.n4 GNDA 0.01577f
C126 pfd_8_0.opamp_out.t2 GNDA 0.021617f
C127 pfd_8_0.opamp_out.n5 GNDA 0.039426f
C128 pfd_8_0.opamp_out.n6 GNDA 0.150316f
C129 pfd_8_0.opamp_out.t15 GNDA 1.72189f
C130 pfd_8_0.opamp_out.n9 GNDA 0.017323f
C131 pfd_8_0.opamp_out.n10 GNDA 0.014909f
C132 pfd_8_0.opamp_out.t10 GNDA 1.72116f
C133 pfd_8_0.opamp_out.n13 GNDA 0.023291f
C134 pfd_8_0.opamp_out.n14 GNDA 0.015404f
C135 opamp_cell_4_0.VOUT GNDA 0.10585f
C136 VDDA.n1 GNDA 0.010245f
C137 VDDA.n2 GNDA 0.010245f
C138 VDDA.n13 GNDA 0.010245f
C139 VDDA.n14 GNDA 0.010245f
C140 VDDA.n20 GNDA 0.062647f
C141 VDDA.t13 GNDA 0.015729f
C142 VDDA.n23 GNDA 0.017227f
C143 VDDA.n25 GNDA 0.010245f
C144 VDDA.t22 GNDA 0.010929f
C145 VDDA.n29 GNDA 0.010093f
C146 VDDA.n34 GNDA 0.010245f
C147 VDDA.n37 GNDA 0.010245f
C148 VDDA.n38 GNDA 0.010245f
C149 VDDA.n41 GNDA 0.010995f
C150 VDDA.n42 GNDA 0.010995f
C151 VDDA.n45 GNDA 0.010995f
C152 VDDA.n48 GNDA 0.010995f
C153 VDDA.n50 GNDA 0.015545f
C154 VDDA.t123 GNDA 0.339084f
C155 VDDA.n55 GNDA 0.015545f
C156 VDDA.n56 GNDA 0.035604f
C157 VDDA.n60 GNDA 0.015545f
C158 VDDA.t77 GNDA 0.213486f
C159 VDDA.t50 GNDA 0.025667f
C160 VDDA.n69 GNDA 0.013565f
C161 VDDA.n72 GNDA 0.013565f
C162 VDDA.n75 GNDA 0.013565f
C163 VDDA.n78 GNDA 0.013565f
C164 VDDA.n82 GNDA 0.011205f
C165 VDDA.t120 GNDA 0.122755f
C166 VDDA.n88 GNDA 0.014509f
C167 VDDA.n91 GNDA 0.014509f
C168 VDDA.n94 GNDA 0.014982f
C169 VDDA.n95 GNDA 0.021082f
C170 VDDA.n97 GNDA 0.014982f
C171 VDDA.n98 GNDA 0.021082f
C172 VDDA.n117 GNDA 0.014982f
C173 VDDA.n120 GNDA 0.014982f
C174 VDDA.n122 GNDA 0.013328f
C175 VDDA.t53 GNDA 0.025829f
C176 VDDA.n126 GNDA 0.010158f
C177 VDDA.n130 GNDA 0.068227f
C178 VDDA.t105 GNDA 0.128092f
C179 VDDA.t40 GNDA 0.138766f
C180 VDDA.t107 GNDA 0.085395f
C181 VDDA.t18 GNDA 0.138766f
C182 VDDA.t64 GNDA 0.14944f
C183 VDDA.t89 GNDA 0.122755f
C184 VDDA.t37 GNDA 0.117418f
C185 VDDA.t65 GNDA 0.011882f
C186 VDDA.n134 GNDA 0.023158f
C187 VDDA.n135 GNDA 0.176059f
C188 VDDA.t83 GNDA 0.160115f
C189 VDDA.n136 GNDA 0.053372f
C190 VDDA.t36 GNDA 0.026192f
C191 VDDA.n150 GNDA 0.018302f
C192 VDDA.n151 GNDA 0.019431f
C193 VDDA.t38 GNDA 0.012954f
C194 VDDA.n152 GNDA 0.013565f
C195 VDDA.n154 GNDA 0.046819f
C196 VDDA.n155 GNDA 0.046596f
C197 VDDA.t49 GNDA 0.011911f
C198 VDDA.n158 GNDA 0.011205f
C199 VDDA.n159 GNDA 0.016038f
C200 VDDA.n160 GNDA 0.011205f
C201 VDDA.n162 GNDA 0.019491f
C202 VDDA.n163 GNDA 0.192062f
C203 VDDA.t60 GNDA 0.181463f
C204 VDDA.t85 GNDA 0.138766f
C205 VDDA.t113 GNDA 0.234835f
C206 VDDA.t87 GNDA 0.138766f
C207 VDDA.t115 GNDA 0.176126f
C208 VDDA.t111 GNDA 0.197475f
C209 VDDA.t54 GNDA 0.138766f
C210 VDDA.t109 GNDA 0.218824f
C211 VDDA.t48 GNDA 0.144103f
C212 VDDA.n164 GNDA 0.289573f
C213 VDDA.n169 GNDA 0.015545f
C214 VDDA.t55 GNDA 0.010363f
C215 VDDA.n170 GNDA 0.014982f
C216 VDDA.n171 GNDA 0.02135f
C217 VDDA.n178 GNDA 0.020046f
C218 VDDA.n185 GNDA 0.021082f
C219 VDDA.n193 GNDA 0.021082f
C220 VDDA.n194 GNDA 0.014982f
C221 VDDA.t58 GNDA 0.010363f
C222 VDDA.n195 GNDA 0.015545f
C223 VDDA.t39 GNDA 0.024372f
C224 VDDA.t56 GNDA 0.024372f
C225 VDDA.n197 GNDA 0.01098f
C226 VDDA.n198 GNDA 0.018711f
C227 VDDA.n199 GNDA 0.015545f
C228 VDDA.n200 GNDA 0.017627f
C229 VDDA.n202 GNDA 0.11208f
C230 VDDA.t103 GNDA 0.117418f
C231 VDDA.t81 GNDA 0.138766f
C232 VDDA.t101 GNDA 0.106743f
C233 VDDA.t57 GNDA 0.138766f
C234 VDDA.t67 GNDA 0.106743f
C235 VDDA.t95 GNDA 0.165452f
C236 VDDA.t29 GNDA 0.138766f
C237 VDDA.t44 GNDA 0.138766f
C238 VDDA.t91 GNDA 0.165452f
C239 VDDA.t92 GNDA 0.186801f
C240 VDDA.t10 GNDA 0.069383f
C241 VDDA.t125 GNDA 0.090732f
C242 VDDA.t5 GNDA 0.192138f
C243 VDDA.t72 GNDA 0.138766f
C244 VDDA.t26 GNDA 0.042697f
C245 VDDA.t75 GNDA 0.138766f
C246 VDDA.t78 GNDA 0.170789f
C247 VDDA.t93 GNDA 0.122755f
C248 VDDA.t79 GNDA 0.213486f
C249 VDDA.t8 GNDA 0.224161f
C250 VDDA.n203 GNDA 0.090656f
C251 VDDA.n204 GNDA 0.019491f
C252 VDDA.n206 GNDA 0.011205f
C253 VDDA.n207 GNDA 0.01448f
C254 VDDA.n212 GNDA 0.045403f
C255 VDDA.n219 GNDA 0.045403f
C256 VDDA.n226 GNDA 0.045403f
C257 VDDA.n233 GNDA 0.045403f
C258 VDDA.n246 GNDA 0.019431f
C259 VDDA.n255 GNDA 0.11208f
C260 VDDA.n261 GNDA 0.532116f
C261 VDDA.n263 GNDA 0.010431f
C262 VDDA.t43 GNDA 0.025829f
C263 VDDA.n271 GNDA 0.025615f
C264 VDDA.n272 GNDA 0.25605f
C265 VDDA.n273 GNDA 0.044061f
C266 VDDA.n286 GNDA 0.010995f
C267 VDDA.n293 GNDA 0.125294f
C268 VDDA.t17 GNDA 0.165452f
C269 VDDA.t31 GNDA 0.146176f
C270 VDDA.t23 GNDA 0.043371f
C271 VDDA.t21 GNDA 0.043371f
C272 VDDA.t24 GNDA 0.010929f
C273 VDDA.n302 GNDA 0.010093f
C274 VDDA.n307 GNDA 0.062647f
C275 VDDA.t119 GNDA 0.010929f
C276 VDDA.n313 GNDA 0.010093f
C277 VDDA.n315 GNDA 0.062647f
C278 VDDA.t14 GNDA 0.043371f
C279 VDDA.t118 GNDA 0.043371f
C280 VDDA.t15 GNDA 0.010929f
C281 VDDA.n318 GNDA 0.010093f
C282 VDDA.n323 GNDA 0.088348f
C283 VDDA.n328 GNDA 0.015545f
C284 VDDA.n334 GNDA 0.015545f
C285 VDDA.n341 GNDA 0.136538f
C286 VDDA.t0 GNDA 0.125294f
C287 VDDA.n343 GNDA 0.015545f
C288 VDDA.n350 GNDA 0.125294f
C289 VDDA.t99 GNDA 0.125294f
C290 VDDA.n357 GNDA 0.015545f
C291 VDDA.n364 GNDA 0.125294f
C292 VDDA.n366 GNDA 0.010995f
C293 VDDA.n371 GNDA 0.039908f
C294 VDDA.n407 GNDA 0.010093f
C295 VDDA.t98 GNDA 0.010929f
C296 VDDA.n409 GNDA 0.010245f
C297 VDDA.n411 GNDA 0.062647f
C298 VDDA.t12 GNDA 0.040158f
C299 VDDA.t3 GNDA 0.038552f
C300 VDDA.t97 GNDA 0.043371f
C301 VDDA.t117 GNDA 0.010929f
C302 VDDA.n418 GNDA 0.010093f
C303 VDDA.t28 GNDA 0.010929f
C304 VDDA.n428 GNDA 0.010093f
C305 VDDA.n430 GNDA 0.094773f
C306 VDDA.t27 GNDA 0.07871f
C307 VDDA.t20 GNDA 0.167058f
C308 VDDA.t33 GNDA 0.167058f
C309 VDDA.t34 GNDA 0.07871f
C310 VDDA.n434 GNDA 0.0114f
C311 VDDA.n435 GNDA 0.013644f
C312 VDDA.n438 GNDA 0.0114f
C313 VDDA.t128 GNDA 0.010935f
C314 VDDA.n441 GNDA 0.011364f
C315 VDDA.n445 GNDA 0.0114f
C316 VDDA.n446 GNDA 0.011364f
C317 VDDA.n449 GNDA 0.0114f
C318 VDDA.t71 GNDA 0.010935f
C319 VDDA.n452 GNDA 0.013644f
C320 VDDA.n454 GNDA 0.086742f
C321 VDDA.t70 GNDA 0.07871f
C322 VDDA.t16 GNDA 0.167058f
C323 VDDA.t25 GNDA 0.167058f
C324 VDDA.t6 GNDA 0.07871f
C325 VDDA.t74 GNDA 0.010929f
C326 VDDA.n458 GNDA 0.010093f
C327 VDDA.t7 GNDA 0.010929f
C328 VDDA.n468 GNDA 0.010093f
C329 VDDA.n470 GNDA 0.088348f
C330 VDDA.t4 GNDA 0.010875f
C331 VDDA.n474 GNDA 0.010093f
C332 VDDA.n476 GNDA 0.085135f
C333 VDDA.n478 GNDA 0.010051f
.ends

