** sch_path: /foss/designs/my_design/projects/pll/bandgapref/xschem_ngspice/tb_opamp_bandgap.sch
**.subckt tb_opamp_bandgap
VDDA VDDA GND 0.6
Vin1 Vin1 GND 0.3
Vin2 Vin2 GND 0.3 AC 1
x1 VDDA Vout Vin2 Vin1 GND opamp_bandgap2
**** begin user architecture code



.option wnflag=1

* .param VDDGAUSS = agauss(1.8, 0.05, 1)
* .param VDD = VDDGAUSS
* .param VDD = 1.8

* .param TEMPGAUSS = agauss(40, 30, 1)
* .param temp = TEMPGAUSS
.option temp = 26

.control

  save all
   *tran 1u 20m
   ac dec 20 1 1T

  write tb_opamp_bandgap.raw
  set appendwrite

.endc




.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/my_design/projects/pll/bandgapref/xschem_ngspice/opamp_bandgap2.sym # of pins=5
** sym_path: /foss/designs/my_design/projects/pll/bandgapref/xschem_ngspice/opamp_bandgap2.sym
** sch_path: /foss/designs/my_design/projects/pll/bandgapref/xschem_ngspice/opamp_bandgap2.sch
.subckt opamp_bandgap2 VDDA Vout Vin- Vin+ GNDA
*.ipin Vin+
*.opin Vout
*.ipin Vin-
*.ipin GNDA
*.ipin VDDA
XM2 net2 Vin+ net1 GNDA sky130_fd_pr__nfet_01v8 L=0.2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vout Vin- net1 GNDA sky130_fd_pr__nfet_01v8 L=0.2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 net1 net1 GNDA GNDA sky130_fd_pr__nfet_01v8 L=0.2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 net2 net2 VDDA VDDA sky130_fd_pr__pfet_01v8 L=0.2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 Vout net2 VDDA VDDA sky130_fd_pr__pfet_01v8 L=0.2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
