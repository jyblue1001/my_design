magic
tech sky130A
timestamp 1753019372
<< metal1 >>
rect 2950 6685 2990 6690
rect 2950 6655 2955 6685
rect 2985 6655 2990 6685
rect 2950 6650 2990 6655
rect 3030 6685 3070 6690
rect 3030 6655 3035 6685
rect 3065 6655 3070 6685
rect 6045 6685 6085 6690
rect 6045 6655 6050 6685
rect 6080 6655 6085 6685
rect 3030 6650 3070 6655
rect 2905 6580 2945 6585
rect 2905 6550 2910 6580
rect 2940 6550 2945 6580
rect 2905 6545 2945 6550
rect 2915 2760 2935 6545
rect 2960 2455 2980 6650
rect 3280 6525 3300 6650
rect 3400 6645 3440 6650
rect 3400 6615 3405 6645
rect 3435 6615 3440 6645
rect 3400 6610 3440 6615
rect 3270 6520 3310 6525
rect 3270 6490 3275 6520
rect 3305 6490 3310 6520
rect 3270 6485 3310 6490
rect 3555 6480 3575 6655
rect 3955 6645 3995 6650
rect 3955 6615 3960 6645
rect 3990 6615 3995 6645
rect 3955 6610 3995 6615
rect 3545 6475 3585 6480
rect 3545 6445 3550 6475
rect 3580 6445 3585 6475
rect 3545 6440 3585 6445
rect 3965 3410 3985 6610
rect 4340 6585 4360 6655
rect 4330 6580 4370 6585
rect 4330 6550 4335 6580
rect 4365 6550 4370 6580
rect 4330 6545 4370 6550
rect 4025 6475 4065 6480
rect 4025 6445 4030 6475
rect 4060 6445 4065 6475
rect 4025 6440 4065 6445
rect 3955 3405 3995 3410
rect 3955 3375 3960 3405
rect 3990 3375 3995 3405
rect 3955 3370 3995 3375
rect 4035 2920 4055 6440
rect 5085 5465 5105 6655
rect 5730 6585 5750 6655
rect 6045 6650 6085 6655
rect 6700 6685 6740 6690
rect 6700 6655 6705 6685
rect 6735 6655 6740 6685
rect 7020 6685 7060 6690
rect 7020 6655 7025 6685
rect 7055 6655 7060 6685
rect 6700 6650 6740 6655
rect 5720 6580 5760 6585
rect 5720 6550 5725 6580
rect 5755 6550 5760 6580
rect 5720 6545 5760 6550
rect 5375 6520 5415 6525
rect 5375 6490 5380 6520
rect 5410 6490 5415 6520
rect 5375 6485 5415 6490
rect 5075 5460 5115 5465
rect 5075 5430 5080 5460
rect 5110 5430 5115 5460
rect 5075 5425 5115 5430
rect 5385 5420 5405 6485
rect 5375 5415 5415 5420
rect 5375 5385 5380 5415
rect 5410 5385 5415 5415
rect 5375 5380 5415 5385
rect 5495 5415 5535 5420
rect 5495 5385 5500 5415
rect 5530 5385 5535 5415
rect 5495 5380 5535 5385
rect 5505 4805 5525 5380
rect 5495 4800 5535 4805
rect 5495 4770 5500 4800
rect 5530 4770 5535 4800
rect 5495 4765 5535 4770
rect 6055 3730 6075 6650
rect 6105 5460 6145 5465
rect 6105 5430 6110 5460
rect 6140 5430 6145 5460
rect 6785 5440 6805 6655
rect 7020 6650 7060 6655
rect 7100 6685 7140 6690
rect 7100 6655 7105 6685
rect 7135 6655 7140 6685
rect 7100 6650 7140 6655
rect 6105 5425 6145 5430
rect 6425 5435 6465 5440
rect 6045 3725 6085 3730
rect 6045 3695 6050 3725
rect 6080 3695 6085 3725
rect 6045 3690 6085 3695
rect 6115 2920 6135 5425
rect 6425 5405 6430 5435
rect 6460 5405 6465 5435
rect 6425 5400 6465 5405
rect 6775 5435 6815 5440
rect 6775 5405 6780 5435
rect 6810 5405 6815 5435
rect 6775 5400 6815 5405
rect 6435 4870 6455 5400
rect 6425 4865 6465 4870
rect 6425 4835 6430 4865
rect 6460 4835 6465 4865
rect 6425 4830 6465 4835
rect 4025 2915 4065 2920
rect 4025 2885 4030 2915
rect 4060 2885 4065 2915
rect 4025 2880 4065 2885
rect 4970 2915 5010 2920
rect 4970 2885 4975 2915
rect 5005 2885 5010 2915
rect 4970 2880 5010 2885
rect 5025 2915 5065 2920
rect 5025 2885 5030 2915
rect 5060 2885 5065 2915
rect 5025 2880 5065 2885
rect 6105 2915 6145 2920
rect 6105 2885 6110 2915
rect 6140 2885 6145 2915
rect 6105 2880 6145 2885
rect 4980 2830 5000 2880
rect 4970 2825 5010 2830
rect 4970 2795 4975 2825
rect 5005 2795 5010 2825
rect 4970 2790 5010 2795
rect 5035 2400 5055 2880
rect 7110 2455 7130 6650
rect 7145 6580 7185 6585
rect 7145 6550 7150 6580
rect 7180 6550 7185 6580
rect 7145 6545 7185 6550
rect 7155 2760 7175 6545
rect 5025 2395 5065 2400
rect 5025 2365 5030 2395
rect 5060 2365 5065 2395
rect 5025 2360 5065 2365
<< via1 >>
rect 2955 6655 2985 6685
rect 3035 6655 3065 6685
rect 6050 6655 6080 6685
rect 2910 6550 2940 6580
rect 3405 6615 3435 6645
rect 3275 6490 3305 6520
rect 3960 6615 3990 6645
rect 3550 6445 3580 6475
rect 4335 6550 4365 6580
rect 4030 6445 4060 6475
rect 3960 3375 3990 3405
rect 6705 6655 6735 6685
rect 7025 6655 7055 6685
rect 5725 6550 5755 6580
rect 5380 6490 5410 6520
rect 5080 5430 5110 5460
rect 5380 5385 5410 5415
rect 5500 5385 5530 5415
rect 5500 4770 5530 4800
rect 6110 5430 6140 5460
rect 7105 6655 7135 6685
rect 4945 3680 4975 3710
rect 6050 3695 6080 3725
rect 6430 5405 6460 5435
rect 6780 5405 6810 5435
rect 6430 4835 6460 4865
rect 4030 2885 4060 2915
rect 4975 2885 5005 2915
rect 5030 2885 5060 2915
rect 6110 2885 6140 2915
rect 4975 2795 5005 2825
rect 7150 6550 7180 6580
rect 5030 2365 5060 2395
<< metal2 >>
rect 2950 6685 2990 6690
rect 2950 6655 2955 6685
rect 2985 6680 2990 6685
rect 3030 6685 3070 6690
rect 3030 6680 3035 6685
rect 2985 6660 3035 6680
rect 2985 6655 2990 6660
rect 2950 6650 2990 6655
rect 3030 6655 3035 6660
rect 3065 6655 3070 6685
rect 3030 6650 3070 6655
rect 6045 6685 6085 6690
rect 6045 6655 6050 6685
rect 6080 6680 6085 6685
rect 6700 6685 6740 6690
rect 6700 6680 6705 6685
rect 6080 6660 6705 6680
rect 6080 6655 6085 6660
rect 6045 6650 6085 6655
rect 6700 6655 6705 6660
rect 6735 6655 6740 6685
rect 7020 6685 7060 6690
rect 7020 6680 7025 6685
rect 7010 6660 7025 6680
rect 6700 6650 6740 6655
rect 7020 6655 7025 6660
rect 7055 6680 7060 6685
rect 7100 6685 7140 6690
rect 7100 6680 7105 6685
rect 7055 6660 7105 6680
rect 7055 6655 7060 6660
rect 7020 6650 7060 6655
rect 7100 6655 7105 6660
rect 7135 6655 7140 6685
rect 7100 6650 7140 6655
rect 3400 6645 3440 6650
rect 3400 6615 3405 6645
rect 3435 6640 3440 6645
rect 3955 6645 3995 6650
rect 3955 6640 3960 6645
rect 3435 6620 3960 6640
rect 3435 6615 3440 6620
rect 3400 6610 3440 6615
rect 3955 6615 3960 6620
rect 3990 6615 3995 6645
rect 3955 6610 3995 6615
rect 2905 6580 2945 6585
rect 2905 6550 2910 6580
rect 2940 6575 2945 6580
rect 4330 6580 4370 6585
rect 4330 6575 4335 6580
rect 2940 6555 4335 6575
rect 2940 6550 2945 6555
rect 2905 6545 2945 6550
rect 4330 6550 4335 6555
rect 4365 6550 4370 6580
rect 4330 6545 4370 6550
rect 5720 6580 5760 6585
rect 5720 6550 5725 6580
rect 5755 6575 5760 6580
rect 7145 6580 7185 6585
rect 7145 6575 7150 6580
rect 5755 6555 7150 6575
rect 5755 6550 5760 6555
rect 5720 6545 5760 6550
rect 7145 6550 7150 6555
rect 7180 6550 7185 6580
rect 7145 6545 7185 6550
rect 3270 6520 3310 6525
rect 3270 6490 3275 6520
rect 3305 6515 3310 6520
rect 5375 6520 5415 6525
rect 5375 6515 5380 6520
rect 3305 6495 5380 6515
rect 3305 6490 3310 6495
rect 3270 6485 3310 6490
rect 5375 6490 5380 6495
rect 5410 6490 5415 6520
rect 5375 6485 5415 6490
rect 3545 6475 3585 6480
rect 3545 6445 3550 6475
rect 3580 6470 3585 6475
rect 4025 6475 4065 6480
rect 4025 6470 4030 6475
rect 3580 6450 4030 6470
rect 3580 6445 3585 6450
rect 3545 6440 3585 6445
rect 4025 6445 4030 6450
rect 4060 6445 4065 6475
rect 4025 6440 4065 6445
rect 5075 5460 5115 5465
rect 5075 5430 5080 5460
rect 5110 5455 5115 5460
rect 6105 5460 6145 5465
rect 6105 5455 6110 5460
rect 5110 5435 6110 5455
rect 5110 5430 5115 5435
rect 5075 5425 5115 5430
rect 6105 5430 6110 5435
rect 6140 5430 6145 5460
rect 6105 5425 6145 5430
rect 6425 5435 6465 5440
rect 5375 5415 5415 5420
rect 5375 5385 5380 5415
rect 5410 5410 5415 5415
rect 5495 5415 5535 5420
rect 5495 5410 5500 5415
rect 5410 5390 5500 5410
rect 5410 5385 5415 5390
rect 5375 5380 5415 5385
rect 5495 5385 5500 5390
rect 5530 5385 5535 5415
rect 6425 5405 6430 5435
rect 6460 5430 6465 5435
rect 6775 5435 6815 5440
rect 6775 5430 6780 5435
rect 6460 5410 6780 5430
rect 6460 5405 6465 5410
rect 6425 5400 6465 5405
rect 6775 5405 6780 5410
rect 6810 5405 6815 5435
rect 6775 5400 6815 5405
rect 5495 5380 5535 5385
rect 6425 4865 6465 4870
rect 6425 4860 6430 4865
rect 5750 4840 6430 4860
rect 6425 4835 6430 4840
rect 6460 4835 6465 4865
rect 6425 4830 6465 4835
rect 5495 4800 5535 4805
rect 5495 4770 5500 4800
rect 5530 4770 5535 4800
rect 5495 4765 5535 4770
rect 6045 3725 6085 3730
rect 6045 3715 6050 3725
rect 4940 3710 6050 3715
rect 4940 3680 4945 3710
rect 4975 3695 6050 3710
rect 6080 3695 6085 3725
rect 4975 3680 4980 3695
rect 6045 3690 6085 3695
rect 4940 3675 4980 3680
rect 3955 3405 3995 3410
rect 3955 3375 3960 3405
rect 3990 3390 3995 3405
rect 3990 3375 4100 3390
rect 3955 3370 4100 3375
rect 4025 2915 4065 2920
rect 4025 2885 4030 2915
rect 4060 2910 4065 2915
rect 4970 2915 5010 2920
rect 4970 2910 4975 2915
rect 4060 2890 4975 2910
rect 4060 2885 4065 2890
rect 4025 2880 4065 2885
rect 4970 2885 4975 2890
rect 5005 2885 5010 2915
rect 4970 2880 5010 2885
rect 5025 2915 5065 2920
rect 5025 2885 5030 2915
rect 5060 2910 5065 2915
rect 6105 2915 6145 2920
rect 6105 2910 6110 2915
rect 5060 2890 6110 2910
rect 5060 2885 5065 2890
rect 5025 2880 5065 2885
rect 6105 2885 6110 2890
rect 6140 2885 6145 2915
rect 6105 2880 6145 2885
rect 4970 2825 5010 2830
rect 4970 2795 4975 2825
rect 5005 2795 5010 2825
rect 4970 2790 5010 2795
rect 5025 2395 5065 2400
rect 5025 2365 5030 2395
rect 5060 2365 5065 2395
rect 5025 2360 5065 2365
rect 4110 2315 4130 2335
rect 5960 2315 5980 2335
rect 2645 1735 2665 1755
rect 7380 1735 7400 1755
<< metal3 >>
rect 9685 14460 9735 14465
rect 9685 14420 9690 14460
rect 9730 14420 9735 14460
rect 9685 14415 9735 14420
rect 9690 50 9730 14415
rect 9685 45 9735 50
rect 9685 5 9690 45
rect 9730 5 9735 45
rect 9685 0 9735 5
<< via3 >>
rect 9690 14420 9730 14460
rect 9690 5 9730 45
<< metal4 >>
rect 7255 14460 9735 14465
rect 7255 14420 9690 14460
rect 9730 14420 9735 14460
rect 7255 14415 9735 14420
rect 540 6700 590 6750
rect 540 0 590 50
rect 9685 45 9735 50
rect 9685 5 9690 45
rect 9730 5 9735 45
rect 9685 0 9735 5
use bgr_10  bgr_10_0
timestamp 1753013163
transform -1 0 22845 0 -1 8250
box 15505 -6295 20095 1600
use two_stage_opamp_dummy_magic_20  two_stage_opamp_dummy_magic_20_0
timestamp 1753018492
transform 1 0 -51855 0 1 555
box 51855 -555 61545 6195
<< labels >>
flabel metal4 565 0 565 0 5 FreeSans 800 0 0 -320 GNDA
port 2 s
flabel metal4 565 6750 565 6750 1 FreeSans 800 0 0 320 VDDA
port 1 n
flabel metal2 5980 2325 5980 2325 3 FreeSans 800 0 320 0 VIN-
port 6 e
flabel metal2 4110 2325 4110 2325 7 FreeSans 800 0 -320 0 VIN+
port 5 w
flabel metal2 7390 1735 7390 1735 5 FreeSans 800 0 0 -320 VOUT-
port 4 s
flabel metal2 2655 1735 2655 1735 5 FreeSans 800 0 0 -320 VOUT+
port 3 s
<< end >>
