** sch_path: /foss/designs/my_design/projects/pll/charge_pump/magic/pfd_charge_pump_magic_2.sch
**.subckt pfd_charge_pump_magic_2
V1 VDD GND 1.8
V2 F_REF GND pulse(0 1.8 12ns 1ns 1ns 24ns 50ns)
V3 F_VCO GND pulse(0 1.8 12ns 1ns 1ns 24ns 50ns)
I1 GND I_IN 100u
x3 DOWN_input VDD GND UP_input net1 F_REF I_IN F_VCO UP_b DOWN pfd_cp_input_magic
x2 VDD GND x V_OUT UP_b DOWN I_IN UP_input DOWN_input opamp_out charge_pump_magic
x4 VDD V_OUT x opamp_out GND rail_to_rail_opamp_magic
x1 V_OUT GND loop_filter_magic
**** begin user architecture code
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt



.include /foss/designs/my_design/projects/pll/charge_pump/magic/pfd_cp_input_magic.spice
.include /foss/designs/my_design/projects/pll/charge_pump/magic/charge_pump_magic.spice
.include /foss/designs/my_design/projects/pll/charge_pump/magic/rail_to_rail_opamp_magic.spice
.include /foss/designs/my_design/projects/pll/charge_pump/magic/loop_filter_magic.spice

.option method=gear
.option wnflag=1
.option savecurrents

* V_out initial voltage value for the F_VCO delay of 2ns  (leading)
* .ic v(v_out) = 1.8

* V_out initial voltage value for the F_VCO delay of 12ns (lock condition)
.ic v(v_out) = 0.9

* V_out initial voltage value for the F_VCO delay of 22ns (lagging)
* .ic v(v_out) = 0.0

.control
  save v(f_ref) save v(f_vco) save v(i_in) save v(up_pfd) v(down_pfd) v(up_pfd_b) v(down_pfd_b) v(up) v(up_b) v(down) v(down_b) v(x) v(opamp_out) v(up_input) v(down_input) v(down_gate) v(v_out)
  * save all

  * timestep for exact simulation results
  * tran 5ps 0.5us

  * timestep for faster simulation results
  tran 50ps 0.5us

  remzerovec
  write pfd_charge_pump_magic_2.raw
  set appendwrite

.endc



**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
