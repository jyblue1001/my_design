magic
tech sky130A
timestamp 1737881691
<< error_p >>
rect 1175 295 1190 305
<< nmos >>
rect 270 655 320 905
rect 370 655 420 905
rect 470 655 520 905
rect 570 655 620 905
rect 670 655 720 905
rect 770 655 820 905
rect 870 655 920 905
rect 970 655 1020 905
rect 400 485 415 535
rect 465 485 480 535
rect 530 485 545 535
rect 595 485 610 535
rect 660 485 675 535
rect 725 485 740 535
rect 790 485 805 535
rect 855 485 870 535
rect 400 345 415 395
rect 465 345 480 395
rect 530 345 545 395
rect 595 345 610 395
rect 660 345 675 395
rect 725 345 740 395
rect 790 345 805 395
rect 855 345 870 395
rect 1045 390 1060 440
rect 1110 390 1125 440
rect 1175 390 1190 440
rect 1240 390 1255 440
rect 1305 390 1320 440
rect 1370 390 1385 440
rect 1435 390 1450 440
rect 1500 390 1515 440
rect 1310 230 1325 280
rect 1375 230 1390 280
rect 1440 230 1455 280
rect 1505 230 1520 280
rect 305 90 320 140
rect 370 90 385 140
rect 435 90 450 140
rect 500 90 515 140
rect 660 90 675 140
rect 725 90 740 140
rect 790 90 805 140
rect 855 90 870 140
rect 765 -215 815 35
rect 865 -215 915 35
rect 965 -215 1015 35
rect 1065 -215 1115 35
<< ndiff >>
rect 220 890 270 905
rect 220 670 235 890
rect 255 670 270 890
rect 220 655 270 670
rect 320 890 370 905
rect 320 670 335 890
rect 355 670 370 890
rect 320 655 370 670
rect 420 890 470 905
rect 420 670 435 890
rect 455 670 470 890
rect 420 655 470 670
rect 520 890 570 905
rect 520 670 535 890
rect 555 670 570 890
rect 520 655 570 670
rect 620 890 670 905
rect 620 670 635 890
rect 655 670 670 890
rect 620 655 670 670
rect 720 890 770 905
rect 720 670 735 890
rect 755 670 770 890
rect 720 655 770 670
rect 820 890 870 905
rect 820 670 835 890
rect 855 670 870 890
rect 820 655 870 670
rect 920 890 970 905
rect 920 670 935 890
rect 955 670 970 890
rect 920 655 970 670
rect 1020 890 1070 905
rect 1020 670 1035 890
rect 1055 670 1070 890
rect 1020 655 1070 670
rect 350 520 400 535
rect 350 500 365 520
rect 385 500 400 520
rect 350 485 400 500
rect 415 520 465 535
rect 415 500 430 520
rect 450 500 465 520
rect 415 485 465 500
rect 480 520 530 535
rect 480 500 495 520
rect 515 500 530 520
rect 480 485 530 500
rect 545 520 595 535
rect 545 500 560 520
rect 580 500 595 520
rect 545 485 595 500
rect 610 520 660 535
rect 610 500 625 520
rect 645 500 660 520
rect 610 485 660 500
rect 675 520 725 535
rect 675 500 690 520
rect 710 500 725 520
rect 675 485 725 500
rect 740 520 790 535
rect 740 500 755 520
rect 775 500 790 520
rect 740 485 790 500
rect 805 520 855 535
rect 805 500 820 520
rect 840 500 855 520
rect 805 485 855 500
rect 870 520 920 535
rect 870 500 885 520
rect 905 500 920 520
rect 870 485 920 500
rect 995 425 1045 440
rect 995 405 1010 425
rect 1030 405 1045 425
rect 350 380 400 395
rect 350 360 365 380
rect 385 360 400 380
rect 350 345 400 360
rect 415 380 465 395
rect 415 360 430 380
rect 450 360 465 380
rect 415 345 465 360
rect 480 380 530 395
rect 480 360 495 380
rect 515 360 530 380
rect 480 345 530 360
rect 545 380 595 395
rect 545 360 560 380
rect 580 360 595 380
rect 545 345 595 360
rect 610 380 660 395
rect 610 360 625 380
rect 645 360 660 380
rect 610 345 660 360
rect 675 380 725 395
rect 675 360 690 380
rect 710 360 725 380
rect 675 345 725 360
rect 740 380 790 395
rect 740 360 755 380
rect 775 360 790 380
rect 740 345 790 360
rect 805 380 855 395
rect 805 360 820 380
rect 840 360 855 380
rect 805 345 855 360
rect 870 380 920 395
rect 995 390 1045 405
rect 1060 425 1110 440
rect 1060 405 1075 425
rect 1095 405 1110 425
rect 1060 390 1110 405
rect 1125 425 1175 440
rect 1125 405 1140 425
rect 1160 405 1175 425
rect 1125 390 1175 405
rect 1190 425 1240 440
rect 1190 405 1205 425
rect 1225 405 1240 425
rect 1190 390 1240 405
rect 1255 425 1305 440
rect 1255 405 1270 425
rect 1290 405 1305 425
rect 1255 390 1305 405
rect 1320 425 1370 440
rect 1320 405 1335 425
rect 1355 405 1370 425
rect 1320 390 1370 405
rect 1385 425 1435 440
rect 1385 405 1400 425
rect 1420 405 1435 425
rect 1385 390 1435 405
rect 1450 425 1500 440
rect 1450 405 1465 425
rect 1485 405 1500 425
rect 1450 390 1500 405
rect 1515 425 1565 440
rect 1515 405 1530 425
rect 1550 405 1565 425
rect 1515 390 1565 405
rect 870 360 885 380
rect 905 360 920 380
rect 870 345 920 360
rect 1260 265 1310 280
rect 1260 245 1275 265
rect 1295 245 1310 265
rect 1260 230 1310 245
rect 1325 265 1375 280
rect 1325 245 1340 265
rect 1360 245 1375 265
rect 1325 230 1375 245
rect 1390 265 1440 280
rect 1390 245 1405 265
rect 1425 245 1440 265
rect 1390 230 1440 245
rect 1455 265 1505 280
rect 1455 245 1470 265
rect 1490 245 1505 265
rect 1455 230 1505 245
rect 1520 265 1570 280
rect 1520 245 1535 265
rect 1555 245 1570 265
rect 1520 230 1570 245
rect 255 125 305 140
rect 255 105 270 125
rect 290 105 305 125
rect 255 90 305 105
rect 320 125 370 140
rect 320 105 335 125
rect 355 105 370 125
rect 320 90 370 105
rect 385 125 435 140
rect 385 105 400 125
rect 420 105 435 125
rect 385 90 435 105
rect 450 125 500 140
rect 450 105 465 125
rect 485 105 500 125
rect 450 90 500 105
rect 515 125 565 140
rect 515 105 530 125
rect 550 105 565 125
rect 515 90 565 105
rect 610 125 660 140
rect 610 105 625 125
rect 645 105 660 125
rect 610 90 660 105
rect 675 125 725 140
rect 675 105 690 125
rect 710 105 725 125
rect 675 90 725 105
rect 740 125 790 140
rect 740 105 755 125
rect 775 105 790 125
rect 740 90 790 105
rect 805 125 855 140
rect 805 105 820 125
rect 840 105 855 125
rect 805 90 855 105
rect 870 125 920 140
rect 870 105 885 125
rect 905 105 920 125
rect 870 90 920 105
rect 715 20 765 35
rect 715 -200 730 20
rect 750 -200 765 20
rect 715 -215 765 -200
rect 815 20 865 35
rect 815 -200 830 20
rect 850 -200 865 20
rect 815 -215 865 -200
rect 915 20 965 35
rect 915 -200 930 20
rect 950 -200 965 20
rect 915 -215 965 -200
rect 1015 20 1065 35
rect 1015 -200 1030 20
rect 1050 -200 1065 20
rect 1015 -215 1065 -200
rect 1115 20 1165 35
rect 1115 -200 1130 20
rect 1150 -200 1165 20
rect 1115 -215 1165 -200
<< ndiffc >>
rect 235 670 255 890
rect 335 670 355 890
rect 435 670 455 890
rect 535 670 555 890
rect 635 670 655 890
rect 735 670 755 890
rect 835 670 855 890
rect 935 670 955 890
rect 1035 670 1055 890
rect 365 500 385 520
rect 430 500 450 520
rect 495 500 515 520
rect 560 500 580 520
rect 625 500 645 520
rect 690 500 710 520
rect 755 500 775 520
rect 820 500 840 520
rect 885 500 905 520
rect 1010 405 1030 425
rect 365 360 385 380
rect 430 360 450 380
rect 495 360 515 380
rect 560 360 580 380
rect 625 360 645 380
rect 690 360 710 380
rect 755 360 775 380
rect 820 360 840 380
rect 1075 405 1095 425
rect 1140 405 1160 425
rect 1205 405 1225 425
rect 1270 405 1290 425
rect 1335 405 1355 425
rect 1400 405 1420 425
rect 1465 405 1485 425
rect 1530 405 1550 425
rect 885 360 905 380
rect 1275 245 1295 265
rect 1340 245 1360 265
rect 1405 245 1425 265
rect 1470 245 1490 265
rect 1535 245 1555 265
rect 270 105 290 125
rect 335 105 355 125
rect 400 105 420 125
rect 465 105 485 125
rect 530 105 550 125
rect 625 105 645 125
rect 690 105 710 125
rect 755 105 775 125
rect 820 105 840 125
rect 885 105 905 125
rect 730 -200 750 20
rect 830 -200 850 20
rect 930 -200 950 20
rect 1030 -200 1050 20
rect 1130 -200 1150 20
<< poly >>
rect 325 950 365 960
rect 325 935 335 950
rect 270 930 335 935
rect 355 935 365 950
rect 725 950 765 960
rect 725 935 735 950
rect 355 930 735 935
rect 755 935 765 950
rect 755 930 1020 935
rect 270 920 1020 930
rect 270 905 320 920
rect 370 905 420 920
rect 470 905 520 920
rect 570 905 620 920
rect 670 905 720 920
rect 770 905 820 920
rect 870 905 920 920
rect 970 905 1020 920
rect 270 640 320 655
rect 370 640 420 655
rect 470 640 520 655
rect 570 640 620 655
rect 670 640 720 655
rect 770 640 820 655
rect 870 640 920 655
rect 970 640 1020 655
rect 420 580 460 590
rect 420 565 430 580
rect 400 560 430 565
rect 450 565 460 580
rect 680 580 720 590
rect 680 565 690 580
rect 450 560 690 565
rect 710 565 720 580
rect 710 560 870 565
rect 400 550 870 560
rect 400 535 415 550
rect 465 535 480 550
rect 530 535 545 550
rect 595 535 610 550
rect 660 535 675 550
rect 725 535 740 550
rect 790 535 805 550
rect 855 535 870 550
rect 400 470 415 485
rect 465 470 480 485
rect 530 470 545 485
rect 595 470 610 485
rect 660 470 675 485
rect 725 470 740 485
rect 790 470 805 485
rect 855 470 870 485
rect 1215 465 1255 495
rect 980 450 1515 465
rect 1045 440 1060 450
rect 1110 440 1125 450
rect 1175 440 1190 450
rect 1240 440 1255 450
rect 1305 440 1320 450
rect 1370 440 1385 450
rect 1435 440 1450 450
rect 1500 440 1515 450
rect 400 395 415 410
rect 465 395 480 410
rect 530 405 610 420
rect 530 395 545 405
rect 595 395 610 405
rect 660 395 675 410
rect 725 395 740 410
rect 790 405 870 420
rect 790 395 805 405
rect 855 395 870 405
rect 1045 375 1060 390
rect 1110 375 1125 390
rect 1175 375 1190 390
rect 1240 375 1255 390
rect 1305 375 1320 390
rect 1370 375 1385 390
rect 1435 375 1450 390
rect 1500 375 1515 390
rect 400 335 415 345
rect 465 335 480 345
rect 400 320 480 335
rect 530 330 545 345
rect 595 330 610 345
rect 660 335 675 345
rect 725 335 740 345
rect 660 320 740 335
rect 790 330 805 345
rect 855 330 870 345
rect 1190 295 1325 305
rect 550 290 1325 295
rect 550 285 1190 290
rect 550 265 560 285
rect 580 280 810 285
rect 580 265 590 280
rect 550 255 590 265
rect 800 265 810 280
rect 830 280 1190 285
rect 1310 280 1325 290
rect 1375 280 1390 295
rect 1440 280 1455 295
rect 1505 280 1520 295
rect 830 265 840 280
rect 800 255 840 265
rect 1310 215 1325 230
rect 1375 215 1390 230
rect 1440 215 1455 230
rect 1505 215 1520 230
rect 1310 200 1520 215
rect 680 185 720 195
rect 680 170 690 185
rect 660 165 690 170
rect 710 170 720 185
rect 1480 175 1520 200
rect 710 165 870 170
rect 305 140 320 155
rect 370 140 385 155
rect 435 150 515 165
rect 435 140 450 150
rect 500 140 515 150
rect 660 155 870 165
rect 660 140 675 155
rect 725 140 740 155
rect 790 140 805 155
rect 855 140 870 155
rect 305 80 320 90
rect 370 80 385 90
rect 305 65 385 80
rect 435 75 450 90
rect 500 75 515 90
rect 660 75 675 90
rect 725 75 740 90
rect 790 75 805 90
rect 855 75 870 90
rect 765 35 815 50
rect 865 35 915 50
rect 965 35 1015 50
rect 1065 35 1115 50
rect 765 -230 815 -215
rect 865 -230 915 -215
rect 965 -230 1015 -215
rect 1065 -230 1115 -215
rect 765 -240 1115 -230
rect 765 -245 830 -240
rect 820 -260 830 -245
rect 850 -245 1115 -240
rect 850 -260 860 -245
rect 820 -270 860 -260
<< polycont >>
rect 335 930 355 950
rect 735 930 755 950
rect 430 560 450 580
rect 690 560 710 580
rect 560 265 580 285
rect 810 265 830 285
rect 690 165 710 185
rect 830 -260 850 -240
<< xpolycontact >>
rect 1220 880 1255 1100
rect 1220 545 1255 765
rect 170 -270 390 15
rect 440 -270 660 15
rect 1220 -95 1255 125
rect 1220 -400 1255 -180
<< xpolyres >>
rect 1220 765 1255 880
rect 390 -270 440 15
rect 1220 -180 1255 -95
<< locali >>
rect 1585 1290 1625 1300
rect 1235 1270 1625 1290
rect 1235 1100 1255 1270
rect 1585 1260 1625 1270
rect 285 950 365 960
rect 285 940 335 950
rect 225 890 265 900
rect 225 670 235 890
rect 255 670 265 890
rect 225 660 265 670
rect 285 630 305 940
rect 325 930 335 940
rect 355 930 365 950
rect 325 920 365 930
rect 725 950 765 960
rect 725 930 735 950
rect 755 930 765 950
rect 725 920 765 930
rect 335 900 355 920
rect 735 900 755 920
rect 325 890 365 900
rect 325 670 335 890
rect 355 670 365 890
rect 325 660 365 670
rect 425 890 465 900
rect 425 670 435 890
rect 455 670 465 890
rect 425 660 465 670
rect 525 890 565 900
rect 525 670 535 890
rect 555 670 565 890
rect 525 660 565 670
rect 625 890 665 900
rect 625 670 635 890
rect 655 670 665 890
rect 625 660 665 670
rect 725 890 765 900
rect 725 670 735 890
rect 755 670 765 890
rect 725 660 765 670
rect 825 890 865 900
rect 825 670 835 890
rect 855 670 865 890
rect 825 660 865 670
rect 925 890 965 900
rect 925 670 935 890
rect 955 670 965 890
rect 925 660 965 670
rect 1025 890 1065 900
rect 1025 670 1035 890
rect 1055 670 1065 890
rect 1025 660 1065 670
rect 220 610 305 630
rect 535 630 555 660
rect 935 630 955 660
rect 535 610 955 630
rect 220 15 240 610
rect 275 580 720 590
rect 275 570 430 580
rect 275 190 295 570
rect 420 560 430 570
rect 450 570 690 580
rect 450 560 460 570
rect 420 550 460 560
rect 680 560 690 570
rect 710 560 720 580
rect 680 550 720 560
rect 430 530 450 550
rect 690 530 710 550
rect 355 520 395 530
rect 355 500 365 520
rect 385 500 395 520
rect 355 490 395 500
rect 420 520 460 530
rect 420 500 430 520
rect 450 500 460 520
rect 420 490 460 500
rect 485 520 525 530
rect 485 500 495 520
rect 515 500 525 520
rect 485 490 525 500
rect 550 520 590 530
rect 550 500 560 520
rect 580 500 590 520
rect 550 490 590 500
rect 615 520 655 530
rect 615 500 625 520
rect 645 500 655 520
rect 615 490 655 500
rect 680 520 720 530
rect 680 500 690 520
rect 710 500 720 520
rect 680 490 720 500
rect 745 520 785 530
rect 745 500 755 520
rect 775 500 785 520
rect 745 490 785 500
rect 810 520 850 530
rect 810 500 820 520
rect 840 500 850 520
rect 810 490 850 500
rect 875 520 915 530
rect 875 500 885 520
rect 905 500 915 520
rect 875 490 915 500
rect 560 470 580 490
rect 820 470 840 490
rect 315 450 840 470
rect 315 250 335 450
rect 935 430 955 610
rect 1235 495 1255 545
rect 1215 455 1255 495
rect 1585 495 1625 535
rect 365 410 955 430
rect 1000 425 1040 435
rect 365 390 385 410
rect 495 390 515 410
rect 625 390 645 410
rect 755 390 775 410
rect 885 390 905 410
rect 1000 405 1010 425
rect 1030 405 1040 425
rect 1000 395 1040 405
rect 1065 425 1105 435
rect 1065 405 1075 425
rect 1095 405 1105 425
rect 1065 395 1105 405
rect 1130 425 1170 435
rect 1130 405 1140 425
rect 1160 405 1170 425
rect 1130 395 1170 405
rect 1195 425 1235 435
rect 1195 405 1205 425
rect 1225 405 1235 425
rect 1195 395 1235 405
rect 1260 425 1300 435
rect 1260 405 1270 425
rect 1290 405 1300 425
rect 1260 395 1300 405
rect 1325 425 1365 435
rect 1325 405 1335 425
rect 1355 405 1365 425
rect 1325 395 1365 405
rect 1390 425 1430 435
rect 1390 405 1400 425
rect 1420 405 1430 425
rect 1390 395 1430 405
rect 1455 425 1495 435
rect 1455 405 1465 425
rect 1485 405 1495 425
rect 1455 395 1495 405
rect 1520 425 1560 435
rect 1520 405 1530 425
rect 1550 405 1560 425
rect 1520 395 1560 405
rect 355 380 395 390
rect 355 360 365 380
rect 385 360 395 380
rect 355 350 395 360
rect 420 380 460 390
rect 420 360 430 380
rect 450 360 460 380
rect 420 350 460 360
rect 485 380 525 390
rect 485 360 495 380
rect 515 360 525 380
rect 485 350 525 360
rect 550 380 590 390
rect 550 360 560 380
rect 580 360 590 380
rect 550 350 590 360
rect 615 380 655 390
rect 615 360 625 380
rect 645 360 655 380
rect 615 350 655 360
rect 680 380 720 390
rect 680 360 690 380
rect 710 360 720 380
rect 680 350 720 360
rect 745 380 785 390
rect 745 360 755 380
rect 775 360 785 380
rect 745 350 785 360
rect 810 380 850 390
rect 810 360 820 380
rect 840 360 850 380
rect 810 350 850 360
rect 875 380 915 390
rect 875 360 885 380
rect 905 360 915 380
rect 875 350 915 360
rect 1075 370 1095 395
rect 1205 370 1225 395
rect 1335 370 1355 395
rect 1465 370 1485 395
rect 1585 370 1605 495
rect 1075 350 1740 370
rect 315 230 410 250
rect 275 170 355 190
rect 335 135 355 170
rect 390 175 410 230
rect 430 235 450 350
rect 560 295 580 350
rect 550 285 590 295
rect 550 265 560 285
rect 580 265 590 285
rect 550 255 590 265
rect 690 235 710 350
rect 820 295 840 350
rect 800 285 840 295
rect 800 265 810 285
rect 830 265 840 285
rect 1340 295 1740 315
rect 1340 275 1360 295
rect 1470 275 1490 295
rect 800 255 840 265
rect 430 215 710 235
rect 690 195 710 215
rect 680 185 720 195
rect 390 155 485 175
rect 680 165 690 185
rect 710 165 720 185
rect 680 155 720 165
rect 465 135 485 155
rect 690 135 710 155
rect 820 135 840 255
rect 1265 265 1305 275
rect 1265 245 1275 265
rect 1295 245 1305 265
rect 1265 235 1305 245
rect 1330 265 1370 275
rect 1330 245 1340 265
rect 1360 245 1370 265
rect 1330 235 1370 245
rect 1395 265 1435 275
rect 1395 245 1405 265
rect 1425 245 1435 265
rect 1395 235 1435 245
rect 1460 265 1500 275
rect 1460 245 1470 265
rect 1490 245 1500 265
rect 1460 235 1500 245
rect 1525 265 1565 275
rect 1525 245 1535 265
rect 1555 245 1565 265
rect 1525 235 1565 245
rect 1585 235 1605 295
rect 1480 175 1520 215
rect 1585 195 1625 235
rect 1500 170 1520 175
rect 260 125 300 135
rect 260 105 270 125
rect 290 105 300 125
rect 260 95 300 105
rect 325 125 365 135
rect 325 105 335 125
rect 355 105 365 125
rect 325 95 365 105
rect 390 125 430 135
rect 390 105 400 125
rect 420 105 430 125
rect 390 95 430 105
rect 455 125 495 135
rect 455 105 465 125
rect 485 105 495 125
rect 455 95 495 105
rect 520 125 560 135
rect 520 105 530 125
rect 550 105 560 125
rect 520 95 560 105
rect 615 125 655 135
rect 615 105 625 125
rect 645 105 655 125
rect 615 95 655 105
rect 680 125 720 135
rect 680 105 690 125
rect 710 105 720 125
rect 680 95 720 105
rect 745 125 785 135
rect 745 105 755 125
rect 775 105 785 125
rect 745 95 785 105
rect 810 125 850 135
rect 810 105 820 125
rect 840 105 850 125
rect 810 95 850 105
rect 875 125 915 135
rect 1235 125 1255 170
rect 875 105 885 125
rect 905 105 915 125
rect 875 95 915 105
rect 270 70 290 95
rect 400 70 420 95
rect 530 70 550 95
rect 270 50 1050 70
rect 1030 30 1050 50
rect 720 20 760 30
rect 720 -200 730 20
rect 750 -200 760 20
rect 720 -210 760 -200
rect 820 20 860 30
rect 820 -200 830 20
rect 850 -200 860 20
rect 820 -210 860 -200
rect 920 20 960 30
rect 920 -200 930 20
rect 950 -200 960 20
rect 920 -210 960 -200
rect 1020 20 1060 30
rect 1020 -200 1030 20
rect 1050 -200 1060 20
rect 1020 -210 1060 -200
rect 1120 20 1160 30
rect 1120 -200 1130 20
rect 1150 -200 1160 20
rect 1120 -210 1160 -200
rect 830 -230 850 -210
rect 820 -240 860 -230
rect 820 -245 830 -240
rect 660 -260 830 -245
rect 850 -260 860 -240
rect 660 -270 860 -260
rect 1235 -540 1255 -400
rect 1585 -540 1625 -530
rect 1235 -560 1625 -540
rect 1585 -570 1625 -560
<< metal3 >>
rect 1585 1260 2470 1305
rect 1640 475 2470 1260
rect 1640 -530 2470 255
rect 1585 -575 2470 -530
<< mimcap >>
rect 1655 535 2455 1290
rect 1655 500 1665 535
rect 1700 500 2455 535
rect 1655 490 2455 500
rect 1655 230 2455 240
rect 1655 195 1665 230
rect 1700 195 2455 230
rect 1655 -560 2455 195
<< mimcapcontact >>
rect 1665 500 1700 535
rect 1665 195 1700 230
<< metal4 >>
rect 1585 535 1705 540
rect 1585 500 1665 535
rect 1700 500 1705 535
rect 1585 495 1705 500
rect 1585 230 1705 235
rect 1585 195 1665 230
rect 1700 195 1705 230
rect 1585 190 1705 195
<< end >>
