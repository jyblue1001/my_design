* NGSPICE file created from charge_pump_full_5.ext - technology: sky130A

.subckt charge_pump_cell w_17500_3540# a_19460_4470# a_17540_4470# OPAMP_out a_17800_2610#
X0 a_17540_4470# OPAMP_out w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X1 a_17540_4470# OPAMP_out w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X2 a_17540_4470# I_IN a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X3 a_17540_4470# OPAMP_out w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X4 w_17500_3540# a_18890_3120# a_19460_4470# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X5 a_19460_4470# a_18890_3120# w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X6 a_18600_3120# a_18310_3120# a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X7 a_20050_3120# a_19470_3120# a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X8 I_IN I_IN a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X9 a_17800_2610# I_IN a_17540_4470# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X10 w_17500_3540# OPAMP_out a_17540_4470# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X11 a_19470_3120# w_17500_3540# a_19050_3120# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X12 a_19460_4470# a_18890_3120# w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X13 w_17500_3540# a_18890_3120# a_19460_4470# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X14 a_18310_3120# a_18020_3120# w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X15 a_20050_3120# a_19470_3120# I_IN w_17500_3540# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X16 I_IN I_IN a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X17 a_18890_3120# a_18600_3120# sky130_fd_pr__cap_mim_m3_1 l=6 w=4.2
X18 w_17500_3540# DOWN_PFD a_19050_3120# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X19 w_17500_3540# OPAMP_out a_17540_4470# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X20 a_19460_4470# a_18890_3120# w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X21 a_18020_3120# UP_PFD w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X22 a_17800_2610# I_IN I_IN a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X23 a_18890_3120# a_18600_3120# OPAMP_out w_17500_3540# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X24 w_17500_3540# a_18890_3120# a_19460_4470# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X25 a_17800_2610# I_IN I_IN a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X26 a_19760_3120# a_19470_3120# w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X27 a_19460_4470# a_18890_3120# w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X28 a_18310_3120# a_18020_3120# a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X29 a_20050_3120# a_19760_3120# I_IN a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X30 a_17800_2610# DOWN_PFD a_19050_3120# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X31 a_17800_2610# a_20050_3120# a_19460_4470# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X32 a_19460_4470# a_20050_3120# a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X33 w_17500_3540# a_18890_3120# a_19460_4470# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X34 a_18020_3120# UP_PFD a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X35 a_20050_3120# a_19760_3120# sky130_fd_pr__cap_mim_m3_1 l=2.6 w=2.6
X36 a_19460_4470# a_20050_3120# a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X37 a_18890_3120# a_18310_3120# OPAMP_out a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X38 a_19760_3120# a_19470_3120# a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X39 w_17500_3540# OPAMP_out a_17540_4470# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X40 a_17800_2610# a_20050_3120# a_19460_4470# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X41 a_17540_4470# OPAMP_out w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X42 a_18890_3120# a_18310_3120# w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X43 a_18600_3120# a_18310_3120# w_17500_3540# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X44 a_19470_3120# a_17800_2610# a_19050_3120# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X45 a_17540_4470# I_IN a_17800_2610# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X46 w_17500_3540# OPAMP_out a_17540_4470# w_17500_3540# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X47 a_17800_2610# I_IN a_17540_4470# a_17800_2610# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
.ends

.subckt opamp_cell w_8020_4460# a_9460_3850# a_7750_4400# a_8190_3850# a_7320_4730#
X0 w_8020_4460# p_bias p_bias w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=1.25 ps=6 w=2.5 l=0.5
X1 w_8020_4460# n_left n_left w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X2 v_common_n a_7320_4730# n_left a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X3 w_8020_4460# p_bias v_common_p w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X4 w_8020_4460# p_bias p_bias w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X5 n_left a_7320_4730# v_common_n a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X6 a_7760_2448# p_right a_8190_3850# sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X7 a_9460_3850# n_right w_8020_4460# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X8 a_9460_3850# a_10686_2448# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X9 v_common_p a_7320_4730# p_left w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X10 a_9460_3850# p_right a_8190_3850# a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X11 w_8020_4460# n_right a_9460_3850# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X12 p_right p_left a_8190_3850# a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X13 p_left a_7320_4730# v_common_p w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X14 a_8190_3850# p_right a_9460_3850# a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X15 a_8190_3850# p_left p_left a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X16 w_8020_4460# p_bias v_common_p w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X17 v_common_n n_bias a_8190_3850# a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X18 n_bias n_bias a_8190_3850# a_8190_3850# sky130_fd_pr__nfet_01v8 ad=1.25 pd=6 as=0.625 ps=3 w=2.5 l=0.5
X19 v_common_p p_bias w_8020_4460# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X20 n_right a_10686_2448# a_8190_3850# sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X21 p_bias p_bias w_8020_4460# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X22 a_9460_3850# n_right w_8020_4460# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X23 a_9460_3850# a_7760_2448# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X24 v_common_p a_7750_4400# p_right w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X25 a_9460_3850# p_right a_8190_3850# a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X26 n_left n_left w_8020_4460# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X27 w_8020_4460# n_right a_9460_3850# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X28 p_left p_left a_8190_3850# a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X29 v_common_n a_7750_4400# n_right a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X30 p_right a_7750_4400# v_common_p w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X31 w_8020_4460# n_left n_right w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X32 a_8190_3850# p_right a_9460_3850# a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X33 a_8190_3850# p_left p_right a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X34 n_right a_7750_4400# v_common_n a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X35 p_bias n_bias a_8190_3850# sky130_fd_pr__res_xhigh_po_2p85 l=0.51
X36 v_common_p p_bias w_8020_4460# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X37 a_8190_3850# n_bias n_bias a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=1.25 ps=6 w=2.5 l=0.5
X38 p_bias p_bias w_8020_4460# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0.625 ps=3 w=2.5 l=0.5
X39 n_right n_left w_8020_4460# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X40 a_8190_3850# n_bias v_common_n a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
.ends

**.subckt charge_pump_full_5
Xcharge_pump_cell_0 VDDA VOUT a_12100_n1150# charge_pump_cell_0/OPAMP_out GNDA charge_pump_cell
Xopamp_cell_0 VDDA charge_pump_cell_0/OPAMP_out a_12100_n1150# GNDA VOUT opamp_cell
**.ends

