magic
tech sky130A
timestamp 1753679884
<< nwell >>
rect 56025 4545 56365 4935
rect 56495 4545 56835 4765
rect 56965 4545 57305 4935
rect 57435 4545 57775 4935
rect 54860 3670 55745 4060
rect 55945 3670 56825 4060
rect 56975 3670 57855 4060
rect 58055 3670 58940 4060
rect 54760 2645 55580 3285
rect 56215 3185 57585 3275
rect 55970 2875 56790 2965
rect 57010 2875 57830 2965
rect 58220 2645 59040 3285
rect 58715 2640 58855 2645
rect 54760 1945 55580 2185
rect 58220 1945 59040 2185
<< nmos >>
rect 56810 2335 56825 2585
rect 56865 2335 56880 2585
rect 56920 2335 56935 2585
rect 56975 2335 56990 2585
rect 56070 2030 56085 2180
rect 56125 2030 56140 2180
rect 56180 2030 56195 2180
rect 56235 2030 56250 2180
rect 56290 2030 56305 2180
rect 56345 2030 56360 2180
rect 56400 2030 56415 2180
rect 56455 2030 56470 2180
rect 56510 2030 56525 2180
rect 56565 2030 56580 2180
rect 56620 2030 56635 2180
rect 56675 2030 56690 2180
rect 57110 2030 57125 2180
rect 57165 2030 57180 2180
rect 57220 2030 57235 2180
rect 57275 2030 57290 2180
rect 57330 2030 57345 2180
rect 57385 2030 57400 2180
rect 57440 2030 57455 2180
rect 57495 2030 57510 2180
rect 57550 2030 57565 2180
rect 57605 2030 57620 2180
rect 57660 2030 57675 2180
rect 57715 2030 57730 2180
rect 54860 1425 54875 1725
rect 54915 1425 54930 1725
rect 54970 1425 54985 1725
rect 55025 1425 55040 1725
rect 55080 1425 55095 1725
rect 55135 1425 55150 1725
rect 55190 1425 55205 1725
rect 55245 1425 55260 1725
rect 55300 1425 55315 1725
rect 55355 1425 55370 1725
rect 55410 1425 55425 1725
rect 55465 1425 55480 1725
rect 56070 1560 56085 1710
rect 56125 1560 56140 1710
rect 56180 1560 56195 1710
rect 56235 1560 56250 1710
rect 56290 1560 56305 1710
rect 56345 1560 56360 1710
rect 56400 1560 56415 1710
rect 56455 1560 56470 1710
rect 56510 1560 56525 1710
rect 56565 1560 56580 1710
rect 56620 1560 56635 1710
rect 56675 1560 56690 1710
rect 56810 1560 56825 1710
rect 56865 1560 56880 1710
rect 56920 1560 56935 1710
rect 56975 1560 56990 1710
rect 57110 1560 57125 1710
rect 57165 1560 57180 1710
rect 57220 1560 57235 1710
rect 57275 1560 57290 1710
rect 57330 1560 57345 1710
rect 57385 1560 57400 1710
rect 57440 1560 57455 1710
rect 57495 1560 57510 1710
rect 57550 1560 57565 1710
rect 57605 1560 57620 1710
rect 57660 1560 57675 1710
rect 57715 1560 57730 1710
rect 58320 1425 58335 1725
rect 58375 1425 58390 1725
rect 58430 1425 58445 1725
rect 58485 1425 58500 1725
rect 58540 1425 58555 1725
rect 58595 1425 58610 1725
rect 58650 1425 58665 1725
rect 58705 1425 58720 1725
rect 58760 1425 58775 1725
rect 58815 1425 58830 1725
rect 58870 1425 58885 1725
rect 58925 1425 58940 1725
rect 54870 355 54930 1055
rect 54970 355 55030 1055
rect 55070 355 55130 1055
rect 55170 355 55230 1055
rect 55270 355 55330 1055
rect 55370 355 55430 1055
rect 56260 760 56275 1010
rect 56315 760 56330 1010
rect 56370 760 56385 1010
rect 56425 760 56440 1010
rect 56480 760 56495 1010
rect 56535 760 56550 1010
rect 56590 760 56605 1010
rect 56645 760 56660 1010
rect 56700 760 56715 1010
rect 56755 760 56770 1010
rect 56810 760 56825 1010
rect 56865 760 56880 1010
rect 56920 760 56935 1010
rect 56975 760 56990 1010
rect 57030 760 57045 1010
rect 57085 760 57100 1010
rect 57140 760 57155 1010
rect 57195 760 57210 1010
rect 57250 760 57265 1010
rect 57305 760 57320 1010
rect 57360 760 57375 1010
rect 57415 760 57430 1010
rect 57470 760 57485 1010
rect 56470 395 56485 545
rect 56525 395 56540 545
rect 56580 395 56595 545
rect 56635 395 56650 545
rect 56690 395 56705 545
rect 56745 395 56760 545
rect 56910 395 57210 545
rect 58370 355 58430 1055
rect 58470 355 58530 1055
rect 58570 355 58630 1055
rect 58670 355 58730 1055
rect 58770 355 58830 1055
rect 58870 355 58930 1055
<< pmos >>
rect 56125 4565 56145 4915
rect 56185 4565 56205 4915
rect 56245 4565 56265 4915
rect 56595 4565 56615 4745
rect 56655 4565 56675 4745
rect 56715 4565 56735 4745
rect 57065 4565 57085 4915
rect 57125 4565 57145 4915
rect 57185 4565 57205 4915
rect 57535 4565 57555 4915
rect 57595 4565 57615 4915
rect 57655 4565 57675 4915
rect 54960 3690 54980 4040
rect 55020 3690 55040 4040
rect 55080 3690 55100 4040
rect 55140 3690 55160 4040
rect 55200 3690 55220 4040
rect 55260 3690 55280 4040
rect 55320 3690 55340 4040
rect 55380 3690 55400 4040
rect 55440 3690 55460 4040
rect 55500 3690 55520 4040
rect 55560 3690 55580 4040
rect 55620 3690 55640 4040
rect 56045 3690 56065 4040
rect 56105 3690 56125 4040
rect 56165 3690 56185 4040
rect 56225 3690 56245 4040
rect 56285 3690 56305 4040
rect 56345 3690 56365 4040
rect 56405 3690 56425 4040
rect 56465 3690 56485 4040
rect 56525 3690 56545 4040
rect 56585 3690 56605 4040
rect 56645 3690 56665 4040
rect 56705 3690 56725 4040
rect 57075 3690 57095 4040
rect 57135 3690 57155 4040
rect 57195 3690 57215 4040
rect 57255 3690 57275 4040
rect 57315 3690 57335 4040
rect 57375 3690 57395 4040
rect 57435 3690 57455 4040
rect 57495 3690 57515 4040
rect 57555 3690 57575 4040
rect 57615 3690 57635 4040
rect 57675 3690 57695 4040
rect 57735 3690 57755 4040
rect 58160 3690 58180 4040
rect 58220 3690 58240 4040
rect 58280 3690 58300 4040
rect 58340 3690 58360 4040
rect 58400 3690 58420 4040
rect 58460 3690 58480 4040
rect 58520 3690 58540 4040
rect 58580 3690 58600 4040
rect 58640 3690 58660 4040
rect 58700 3690 58720 4040
rect 58760 3690 58780 4040
rect 58820 3690 58840 4040
rect 54860 2665 54875 3265
rect 54915 2665 54930 3265
rect 54970 2665 54985 3265
rect 55025 2665 55040 3265
rect 55080 2665 55095 3265
rect 55135 2665 55150 3265
rect 55190 2665 55205 3265
rect 55245 2665 55260 3265
rect 55300 2665 55315 3265
rect 55355 2665 55370 3265
rect 55410 2665 55425 3265
rect 55465 2665 55480 3265
rect 56315 3205 56330 3255
rect 56370 3205 56385 3255
rect 56425 3205 56440 3255
rect 56480 3205 56495 3255
rect 56535 3205 56550 3255
rect 56590 3205 56605 3255
rect 56645 3205 56660 3255
rect 56700 3205 56715 3255
rect 56755 3205 56770 3255
rect 56810 3205 56825 3255
rect 56865 3205 56880 3255
rect 56920 3205 56935 3255
rect 56975 3205 56990 3255
rect 57030 3205 57045 3255
rect 57085 3205 57100 3255
rect 57140 3205 57155 3255
rect 57195 3205 57210 3255
rect 57250 3205 57265 3255
rect 57305 3205 57320 3255
rect 57360 3205 57375 3255
rect 57415 3205 57430 3255
rect 57470 3205 57485 3255
rect 56070 2895 56085 2945
rect 56125 2895 56140 2945
rect 56180 2895 56195 2945
rect 56235 2895 56250 2945
rect 56290 2895 56305 2945
rect 56345 2895 56360 2945
rect 56400 2895 56415 2945
rect 56455 2895 56470 2945
rect 56510 2895 56525 2945
rect 56565 2895 56580 2945
rect 56620 2895 56635 2945
rect 56675 2895 56690 2945
rect 57110 2895 57125 2945
rect 57165 2895 57180 2945
rect 57220 2895 57235 2945
rect 57275 2895 57290 2945
rect 57330 2895 57345 2945
rect 57385 2895 57400 2945
rect 57440 2895 57455 2945
rect 57495 2895 57510 2945
rect 57550 2895 57565 2945
rect 57605 2895 57620 2945
rect 57660 2895 57675 2945
rect 57715 2895 57730 2945
rect 58320 2665 58335 3265
rect 58375 2665 58390 3265
rect 58430 2665 58445 3265
rect 58485 2665 58500 3265
rect 58540 2665 58555 3265
rect 58595 2665 58610 3265
rect 58650 2665 58665 3265
rect 58705 2665 58720 3265
rect 58760 2665 58775 3265
rect 58815 2665 58830 3265
rect 58870 2665 58885 3265
rect 58925 2665 58940 3265
rect 54860 1965 54875 2165
rect 54915 1965 54930 2165
rect 54970 1965 54985 2165
rect 55025 1965 55040 2165
rect 55080 1965 55095 2165
rect 55135 1965 55150 2165
rect 55190 1965 55205 2165
rect 55245 1965 55260 2165
rect 55300 1965 55315 2165
rect 55355 1965 55370 2165
rect 55410 1965 55425 2165
rect 55465 1965 55480 2165
rect 58320 1965 58335 2165
rect 58375 1965 58390 2165
rect 58430 1965 58445 2165
rect 58485 1965 58500 2165
rect 58540 1965 58555 2165
rect 58595 1965 58610 2165
rect 58650 1965 58665 2165
rect 58705 1965 58720 2165
rect 58760 1965 58775 2165
rect 58815 1965 58830 2165
rect 58870 1965 58885 2165
rect 58925 1965 58940 2165
<< ndiff >>
rect 56770 2570 56810 2585
rect 56770 2350 56780 2570
rect 56800 2350 56810 2570
rect 56770 2335 56810 2350
rect 56825 2570 56865 2585
rect 56825 2350 56835 2570
rect 56855 2350 56865 2570
rect 56825 2335 56865 2350
rect 56880 2570 56920 2585
rect 56880 2350 56890 2570
rect 56910 2350 56920 2570
rect 56880 2335 56920 2350
rect 56935 2570 56975 2585
rect 56935 2350 56945 2570
rect 56965 2350 56975 2570
rect 56935 2335 56975 2350
rect 56990 2570 57030 2585
rect 56990 2350 57000 2570
rect 57020 2350 57030 2570
rect 56990 2335 57030 2350
rect 56030 2165 56070 2180
rect 56030 2045 56040 2165
rect 56060 2045 56070 2165
rect 56030 2030 56070 2045
rect 56085 2165 56125 2180
rect 56085 2045 56095 2165
rect 56115 2045 56125 2165
rect 56085 2030 56125 2045
rect 56140 2165 56180 2180
rect 56140 2045 56150 2165
rect 56170 2045 56180 2165
rect 56140 2030 56180 2045
rect 56195 2165 56235 2180
rect 56195 2045 56205 2165
rect 56225 2045 56235 2165
rect 56195 2030 56235 2045
rect 56250 2165 56290 2180
rect 56250 2045 56260 2165
rect 56280 2045 56290 2165
rect 56250 2030 56290 2045
rect 56305 2165 56345 2180
rect 56305 2045 56315 2165
rect 56335 2045 56345 2165
rect 56305 2030 56345 2045
rect 56360 2165 56400 2180
rect 56360 2045 56370 2165
rect 56390 2045 56400 2165
rect 56360 2030 56400 2045
rect 56415 2165 56455 2180
rect 56415 2045 56425 2165
rect 56445 2045 56455 2165
rect 56415 2030 56455 2045
rect 56470 2165 56510 2180
rect 56470 2045 56480 2165
rect 56500 2045 56510 2165
rect 56470 2030 56510 2045
rect 56525 2165 56565 2180
rect 56525 2045 56535 2165
rect 56555 2045 56565 2165
rect 56525 2030 56565 2045
rect 56580 2165 56620 2180
rect 56580 2045 56590 2165
rect 56610 2045 56620 2165
rect 56580 2030 56620 2045
rect 56635 2165 56675 2180
rect 56635 2045 56645 2165
rect 56665 2045 56675 2165
rect 56635 2030 56675 2045
rect 56690 2165 56730 2180
rect 56690 2045 56700 2165
rect 56720 2045 56730 2165
rect 56690 2030 56730 2045
rect 57070 2165 57110 2180
rect 57070 2045 57080 2165
rect 57100 2045 57110 2165
rect 57070 2030 57110 2045
rect 57125 2165 57165 2180
rect 57125 2045 57135 2165
rect 57155 2045 57165 2165
rect 57125 2030 57165 2045
rect 57180 2165 57220 2180
rect 57180 2045 57190 2165
rect 57210 2045 57220 2165
rect 57180 2030 57220 2045
rect 57235 2165 57275 2180
rect 57235 2045 57245 2165
rect 57265 2045 57275 2165
rect 57235 2030 57275 2045
rect 57290 2165 57330 2180
rect 57290 2045 57300 2165
rect 57320 2045 57330 2165
rect 57290 2030 57330 2045
rect 57345 2165 57385 2180
rect 57345 2045 57355 2165
rect 57375 2045 57385 2165
rect 57345 2030 57385 2045
rect 57400 2165 57440 2180
rect 57400 2045 57410 2165
rect 57430 2045 57440 2165
rect 57400 2030 57440 2045
rect 57455 2165 57495 2180
rect 57455 2045 57465 2165
rect 57485 2045 57495 2165
rect 57455 2030 57495 2045
rect 57510 2165 57550 2180
rect 57510 2045 57520 2165
rect 57540 2045 57550 2165
rect 57510 2030 57550 2045
rect 57565 2165 57605 2180
rect 57565 2045 57575 2165
rect 57595 2045 57605 2165
rect 57565 2030 57605 2045
rect 57620 2165 57660 2180
rect 57620 2045 57630 2165
rect 57650 2045 57660 2165
rect 57620 2030 57660 2045
rect 57675 2165 57715 2180
rect 57675 2045 57685 2165
rect 57705 2045 57715 2165
rect 57675 2030 57715 2045
rect 57730 2165 57770 2180
rect 57730 2045 57740 2165
rect 57760 2045 57770 2165
rect 57730 2030 57770 2045
rect 54820 1710 54860 1725
rect 54820 1440 54830 1710
rect 54850 1440 54860 1710
rect 54820 1425 54860 1440
rect 54875 1710 54915 1725
rect 54875 1440 54885 1710
rect 54905 1440 54915 1710
rect 54875 1425 54915 1440
rect 54930 1710 54970 1725
rect 54930 1440 54940 1710
rect 54960 1440 54970 1710
rect 54930 1425 54970 1440
rect 54985 1710 55025 1725
rect 54985 1440 54995 1710
rect 55015 1440 55025 1710
rect 54985 1425 55025 1440
rect 55040 1710 55080 1725
rect 55040 1440 55050 1710
rect 55070 1440 55080 1710
rect 55040 1425 55080 1440
rect 55095 1710 55135 1725
rect 55095 1440 55105 1710
rect 55125 1440 55135 1710
rect 55095 1425 55135 1440
rect 55150 1710 55190 1725
rect 55150 1440 55160 1710
rect 55180 1440 55190 1710
rect 55150 1425 55190 1440
rect 55205 1710 55245 1725
rect 55205 1440 55215 1710
rect 55235 1440 55245 1710
rect 55205 1425 55245 1440
rect 55260 1710 55300 1725
rect 55260 1440 55270 1710
rect 55290 1440 55300 1710
rect 55260 1425 55300 1440
rect 55315 1710 55355 1725
rect 55315 1440 55325 1710
rect 55345 1440 55355 1710
rect 55315 1425 55355 1440
rect 55370 1710 55410 1725
rect 55370 1440 55380 1710
rect 55400 1440 55410 1710
rect 55370 1425 55410 1440
rect 55425 1710 55465 1725
rect 55425 1440 55435 1710
rect 55455 1440 55465 1710
rect 55425 1425 55465 1440
rect 55480 1710 55520 1725
rect 58280 1710 58320 1725
rect 55480 1440 55490 1710
rect 55510 1440 55520 1710
rect 56030 1695 56070 1710
rect 56030 1575 56040 1695
rect 56060 1575 56070 1695
rect 56030 1560 56070 1575
rect 56085 1695 56125 1710
rect 56085 1575 56095 1695
rect 56115 1575 56125 1695
rect 56085 1560 56125 1575
rect 56140 1695 56180 1710
rect 56140 1575 56150 1695
rect 56170 1575 56180 1695
rect 56140 1560 56180 1575
rect 56195 1695 56235 1710
rect 56195 1575 56205 1695
rect 56225 1575 56235 1695
rect 56195 1560 56235 1575
rect 56250 1695 56290 1710
rect 56250 1575 56260 1695
rect 56280 1575 56290 1695
rect 56250 1560 56290 1575
rect 56305 1695 56345 1710
rect 56305 1575 56315 1695
rect 56335 1575 56345 1695
rect 56305 1560 56345 1575
rect 56360 1695 56400 1710
rect 56360 1575 56370 1695
rect 56390 1575 56400 1695
rect 56360 1560 56400 1575
rect 56415 1695 56455 1710
rect 56415 1575 56425 1695
rect 56445 1575 56455 1695
rect 56415 1560 56455 1575
rect 56470 1695 56510 1710
rect 56470 1575 56480 1695
rect 56500 1575 56510 1695
rect 56470 1560 56510 1575
rect 56525 1695 56565 1710
rect 56525 1575 56535 1695
rect 56555 1575 56565 1695
rect 56525 1560 56565 1575
rect 56580 1695 56620 1710
rect 56580 1575 56590 1695
rect 56610 1575 56620 1695
rect 56580 1560 56620 1575
rect 56635 1695 56675 1710
rect 56635 1575 56645 1695
rect 56665 1575 56675 1695
rect 56635 1560 56675 1575
rect 56690 1695 56730 1710
rect 56770 1695 56810 1710
rect 56690 1575 56700 1695
rect 56720 1575 56730 1695
rect 56770 1575 56780 1695
rect 56800 1575 56810 1695
rect 56690 1560 56730 1575
rect 56770 1560 56810 1575
rect 56825 1695 56865 1710
rect 56825 1575 56835 1695
rect 56855 1575 56865 1695
rect 56825 1560 56865 1575
rect 56880 1695 56920 1710
rect 56880 1575 56890 1695
rect 56910 1575 56920 1695
rect 56880 1560 56920 1575
rect 56935 1695 56975 1710
rect 56935 1575 56945 1695
rect 56965 1575 56975 1695
rect 56935 1560 56975 1575
rect 56990 1695 57030 1710
rect 57070 1695 57110 1710
rect 56990 1575 57000 1695
rect 57020 1575 57030 1695
rect 57070 1575 57080 1695
rect 57100 1575 57110 1695
rect 56990 1560 57030 1575
rect 57070 1560 57110 1575
rect 57125 1695 57165 1710
rect 57125 1575 57135 1695
rect 57155 1575 57165 1695
rect 57125 1560 57165 1575
rect 57180 1695 57220 1710
rect 57180 1575 57190 1695
rect 57210 1575 57220 1695
rect 57180 1560 57220 1575
rect 57235 1695 57275 1710
rect 57235 1575 57245 1695
rect 57265 1575 57275 1695
rect 57235 1560 57275 1575
rect 57290 1695 57330 1710
rect 57290 1575 57300 1695
rect 57320 1575 57330 1695
rect 57290 1560 57330 1575
rect 57345 1695 57385 1710
rect 57345 1575 57355 1695
rect 57375 1575 57385 1695
rect 57345 1560 57385 1575
rect 57400 1695 57440 1710
rect 57400 1575 57410 1695
rect 57430 1575 57440 1695
rect 57400 1560 57440 1575
rect 57455 1695 57495 1710
rect 57455 1575 57465 1695
rect 57485 1575 57495 1695
rect 57455 1560 57495 1575
rect 57510 1695 57550 1710
rect 57510 1575 57520 1695
rect 57540 1575 57550 1695
rect 57510 1560 57550 1575
rect 57565 1695 57605 1710
rect 57565 1575 57575 1695
rect 57595 1575 57605 1695
rect 57565 1560 57605 1575
rect 57620 1695 57660 1710
rect 57620 1575 57630 1695
rect 57650 1575 57660 1695
rect 57620 1560 57660 1575
rect 57675 1695 57715 1710
rect 57675 1575 57685 1695
rect 57705 1575 57715 1695
rect 57675 1560 57715 1575
rect 57730 1695 57770 1710
rect 57730 1575 57740 1695
rect 57760 1575 57770 1695
rect 57730 1560 57770 1575
rect 55480 1425 55520 1440
rect 58280 1440 58290 1710
rect 58310 1440 58320 1710
rect 58280 1425 58320 1440
rect 58335 1710 58375 1725
rect 58335 1440 58345 1710
rect 58365 1440 58375 1710
rect 58335 1425 58375 1440
rect 58390 1710 58430 1725
rect 58390 1440 58400 1710
rect 58420 1440 58430 1710
rect 58390 1425 58430 1440
rect 58445 1710 58485 1725
rect 58445 1440 58455 1710
rect 58475 1440 58485 1710
rect 58445 1425 58485 1440
rect 58500 1710 58540 1725
rect 58500 1440 58510 1710
rect 58530 1440 58540 1710
rect 58500 1425 58540 1440
rect 58555 1710 58595 1725
rect 58555 1440 58565 1710
rect 58585 1440 58595 1710
rect 58555 1425 58595 1440
rect 58610 1710 58650 1725
rect 58610 1440 58620 1710
rect 58640 1440 58650 1710
rect 58610 1425 58650 1440
rect 58665 1710 58705 1725
rect 58665 1440 58675 1710
rect 58695 1440 58705 1710
rect 58665 1425 58705 1440
rect 58720 1710 58760 1725
rect 58720 1440 58730 1710
rect 58750 1440 58760 1710
rect 58720 1425 58760 1440
rect 58775 1710 58815 1725
rect 58775 1440 58785 1710
rect 58805 1440 58815 1710
rect 58775 1425 58815 1440
rect 58830 1710 58870 1725
rect 58830 1440 58840 1710
rect 58860 1440 58870 1710
rect 58830 1425 58870 1440
rect 58885 1710 58925 1725
rect 58885 1440 58895 1710
rect 58915 1440 58925 1710
rect 58885 1425 58925 1440
rect 58940 1710 58980 1725
rect 58940 1440 58950 1710
rect 58970 1440 58980 1710
rect 58940 1425 58980 1440
rect 54830 1040 54870 1055
rect 54830 370 54840 1040
rect 54860 370 54870 1040
rect 54830 355 54870 370
rect 54930 1040 54970 1055
rect 54930 370 54940 1040
rect 54960 370 54970 1040
rect 54930 355 54970 370
rect 55030 1040 55070 1055
rect 55030 370 55040 1040
rect 55060 370 55070 1040
rect 55030 355 55070 370
rect 55130 1040 55170 1055
rect 55130 370 55140 1040
rect 55160 370 55170 1040
rect 55130 355 55170 370
rect 55230 1040 55270 1055
rect 55230 370 55240 1040
rect 55260 370 55270 1040
rect 55230 355 55270 370
rect 55330 1040 55370 1055
rect 55330 370 55340 1040
rect 55360 370 55370 1040
rect 55330 355 55370 370
rect 55430 1040 55470 1055
rect 55430 370 55440 1040
rect 55460 370 55470 1040
rect 58330 1040 58370 1055
rect 56220 995 56260 1010
rect 56220 775 56230 995
rect 56250 775 56260 995
rect 56220 760 56260 775
rect 56275 995 56315 1010
rect 56275 775 56285 995
rect 56305 775 56315 995
rect 56275 760 56315 775
rect 56330 995 56370 1010
rect 56330 775 56340 995
rect 56360 775 56370 995
rect 56330 760 56370 775
rect 56385 995 56425 1010
rect 56385 775 56395 995
rect 56415 775 56425 995
rect 56385 760 56425 775
rect 56440 995 56480 1010
rect 56440 775 56450 995
rect 56470 775 56480 995
rect 56440 760 56480 775
rect 56495 995 56535 1010
rect 56495 775 56505 995
rect 56525 775 56535 995
rect 56495 760 56535 775
rect 56550 995 56590 1010
rect 56550 775 56560 995
rect 56580 775 56590 995
rect 56550 760 56590 775
rect 56605 995 56645 1010
rect 56605 775 56615 995
rect 56635 775 56645 995
rect 56605 760 56645 775
rect 56660 995 56700 1010
rect 56660 775 56670 995
rect 56690 775 56700 995
rect 56660 760 56700 775
rect 56715 995 56755 1010
rect 56715 775 56725 995
rect 56745 775 56755 995
rect 56715 760 56755 775
rect 56770 995 56810 1010
rect 56770 775 56780 995
rect 56800 775 56810 995
rect 56770 760 56810 775
rect 56825 995 56865 1010
rect 56825 775 56835 995
rect 56855 775 56865 995
rect 56825 760 56865 775
rect 56880 995 56920 1010
rect 56880 775 56890 995
rect 56910 775 56920 995
rect 56880 760 56920 775
rect 56935 995 56975 1010
rect 56935 775 56945 995
rect 56965 775 56975 995
rect 56935 760 56975 775
rect 56990 995 57030 1010
rect 56990 775 57000 995
rect 57020 775 57030 995
rect 56990 760 57030 775
rect 57045 995 57085 1010
rect 57045 775 57055 995
rect 57075 775 57085 995
rect 57045 760 57085 775
rect 57100 995 57140 1010
rect 57100 775 57110 995
rect 57130 775 57140 995
rect 57100 760 57140 775
rect 57155 995 57195 1010
rect 57155 775 57165 995
rect 57185 775 57195 995
rect 57155 760 57195 775
rect 57210 995 57250 1010
rect 57210 775 57220 995
rect 57240 775 57250 995
rect 57210 760 57250 775
rect 57265 995 57305 1010
rect 57265 775 57275 995
rect 57295 775 57305 995
rect 57265 760 57305 775
rect 57320 995 57360 1010
rect 57320 775 57330 995
rect 57350 775 57360 995
rect 57320 760 57360 775
rect 57375 995 57415 1010
rect 57375 775 57385 995
rect 57405 775 57415 995
rect 57375 760 57415 775
rect 57430 995 57470 1010
rect 57430 775 57440 995
rect 57460 775 57470 995
rect 57430 760 57470 775
rect 57485 995 57525 1010
rect 57485 775 57495 995
rect 57515 775 57525 995
rect 57485 760 57525 775
rect 56430 530 56470 545
rect 56430 410 56440 530
rect 56460 410 56470 530
rect 56430 395 56470 410
rect 56485 530 56525 545
rect 56485 410 56495 530
rect 56515 410 56525 530
rect 56485 395 56525 410
rect 56540 530 56580 545
rect 56540 410 56550 530
rect 56570 410 56580 530
rect 56540 395 56580 410
rect 56595 530 56635 545
rect 56595 410 56605 530
rect 56625 410 56635 530
rect 56595 395 56635 410
rect 56650 530 56690 545
rect 56650 410 56660 530
rect 56680 410 56690 530
rect 56650 395 56690 410
rect 56705 530 56745 545
rect 56705 410 56715 530
rect 56735 410 56745 530
rect 56705 395 56745 410
rect 56760 530 56800 545
rect 56760 410 56770 530
rect 56790 410 56800 530
rect 56760 395 56800 410
rect 56870 530 56910 545
rect 56870 410 56880 530
rect 56900 410 56910 530
rect 56870 395 56910 410
rect 57210 530 57250 545
rect 57210 410 57220 530
rect 57240 410 57250 530
rect 57210 395 57250 410
rect 55430 355 55470 370
rect 58330 370 58340 1040
rect 58360 370 58370 1040
rect 58330 355 58370 370
rect 58430 1040 58470 1055
rect 58430 370 58440 1040
rect 58460 370 58470 1040
rect 58430 355 58470 370
rect 58530 1040 58570 1055
rect 58530 370 58540 1040
rect 58560 370 58570 1040
rect 58530 355 58570 370
rect 58630 1040 58670 1055
rect 58630 370 58640 1040
rect 58660 370 58670 1040
rect 58630 355 58670 370
rect 58730 1040 58770 1055
rect 58730 370 58740 1040
rect 58760 370 58770 1040
rect 58730 355 58770 370
rect 58830 1040 58870 1055
rect 58830 370 58840 1040
rect 58860 370 58870 1040
rect 58830 355 58870 370
rect 58930 1040 58970 1055
rect 58930 370 58940 1040
rect 58960 370 58970 1040
rect 58930 355 58970 370
<< pdiff >>
rect 56085 4900 56125 4915
rect 56085 4580 56095 4900
rect 56115 4580 56125 4900
rect 56085 4565 56125 4580
rect 56145 4900 56185 4915
rect 56145 4580 56155 4900
rect 56175 4580 56185 4900
rect 56145 4565 56185 4580
rect 56205 4900 56245 4915
rect 56205 4580 56215 4900
rect 56235 4580 56245 4900
rect 56205 4565 56245 4580
rect 56265 4900 56305 4915
rect 56265 4580 56275 4900
rect 56295 4580 56305 4900
rect 57025 4900 57065 4915
rect 56265 4565 56305 4580
rect 56555 4730 56595 4745
rect 56555 4580 56565 4730
rect 56585 4580 56595 4730
rect 56555 4565 56595 4580
rect 56615 4730 56655 4745
rect 56615 4580 56625 4730
rect 56645 4580 56655 4730
rect 56615 4565 56655 4580
rect 56675 4730 56715 4745
rect 56675 4580 56685 4730
rect 56705 4580 56715 4730
rect 56675 4565 56715 4580
rect 56735 4730 56775 4745
rect 56735 4580 56745 4730
rect 56765 4580 56775 4730
rect 56735 4565 56775 4580
rect 57025 4580 57035 4900
rect 57055 4580 57065 4900
rect 57025 4565 57065 4580
rect 57085 4900 57125 4915
rect 57085 4580 57095 4900
rect 57115 4580 57125 4900
rect 57085 4565 57125 4580
rect 57145 4900 57185 4915
rect 57145 4580 57155 4900
rect 57175 4580 57185 4900
rect 57145 4565 57185 4580
rect 57205 4900 57245 4915
rect 57205 4580 57215 4900
rect 57235 4580 57245 4900
rect 57205 4565 57245 4580
rect 57495 4900 57535 4915
rect 57495 4580 57505 4900
rect 57525 4580 57535 4900
rect 57495 4565 57535 4580
rect 57555 4900 57595 4915
rect 57555 4580 57565 4900
rect 57585 4580 57595 4900
rect 57555 4565 57595 4580
rect 57615 4900 57655 4915
rect 57615 4580 57625 4900
rect 57645 4580 57655 4900
rect 57615 4565 57655 4580
rect 57675 4900 57715 4915
rect 57675 4580 57685 4900
rect 57705 4580 57715 4900
rect 57675 4565 57715 4580
rect 54920 4025 54960 4040
rect 54920 3705 54930 4025
rect 54950 3705 54960 4025
rect 54920 3690 54960 3705
rect 54980 4025 55020 4040
rect 54980 3705 54990 4025
rect 55010 3705 55020 4025
rect 54980 3690 55020 3705
rect 55040 4025 55080 4040
rect 55040 3705 55050 4025
rect 55070 3705 55080 4025
rect 55040 3690 55080 3705
rect 55100 4025 55140 4040
rect 55100 3705 55110 4025
rect 55130 3705 55140 4025
rect 55100 3690 55140 3705
rect 55160 4025 55200 4040
rect 55160 3705 55170 4025
rect 55190 3705 55200 4025
rect 55160 3690 55200 3705
rect 55220 4025 55260 4040
rect 55220 3705 55230 4025
rect 55250 3705 55260 4025
rect 55220 3690 55260 3705
rect 55280 4025 55320 4040
rect 55280 3705 55290 4025
rect 55310 3705 55320 4025
rect 55280 3690 55320 3705
rect 55340 4025 55380 4040
rect 55340 3705 55350 4025
rect 55370 3705 55380 4025
rect 55340 3690 55380 3705
rect 55400 4025 55440 4040
rect 55400 3705 55410 4025
rect 55430 3705 55440 4025
rect 55400 3690 55440 3705
rect 55460 4025 55500 4040
rect 55460 3705 55470 4025
rect 55490 3705 55500 4025
rect 55460 3690 55500 3705
rect 55520 4025 55560 4040
rect 55520 3705 55530 4025
rect 55550 3705 55560 4025
rect 55520 3690 55560 3705
rect 55580 4025 55620 4040
rect 55580 3705 55590 4025
rect 55610 3705 55620 4025
rect 55580 3690 55620 3705
rect 55640 4025 55680 4040
rect 55640 3705 55650 4025
rect 55670 3705 55680 4025
rect 55640 3690 55680 3705
rect 56005 4025 56045 4040
rect 56005 3705 56015 4025
rect 56035 3705 56045 4025
rect 56005 3690 56045 3705
rect 56065 4025 56105 4040
rect 56065 3705 56075 4025
rect 56095 3705 56105 4025
rect 56065 3690 56105 3705
rect 56125 4025 56165 4040
rect 56125 3705 56135 4025
rect 56155 3705 56165 4025
rect 56125 3690 56165 3705
rect 56185 4025 56225 4040
rect 56185 3705 56195 4025
rect 56215 3705 56225 4025
rect 56185 3690 56225 3705
rect 56245 4025 56285 4040
rect 56245 3705 56255 4025
rect 56275 3705 56285 4025
rect 56245 3690 56285 3705
rect 56305 4025 56345 4040
rect 56305 3705 56315 4025
rect 56335 3705 56345 4025
rect 56305 3690 56345 3705
rect 56365 4025 56405 4040
rect 56365 3705 56375 4025
rect 56395 3705 56405 4025
rect 56365 3690 56405 3705
rect 56425 4025 56465 4040
rect 56425 3705 56435 4025
rect 56455 3705 56465 4025
rect 56425 3690 56465 3705
rect 56485 4025 56525 4040
rect 56485 3705 56495 4025
rect 56515 3705 56525 4025
rect 56485 3690 56525 3705
rect 56545 4025 56585 4040
rect 56545 3705 56555 4025
rect 56575 3705 56585 4025
rect 56545 3690 56585 3705
rect 56605 4025 56645 4040
rect 56605 3705 56615 4025
rect 56635 3705 56645 4025
rect 56605 3690 56645 3705
rect 56665 4025 56705 4040
rect 56665 3705 56675 4025
rect 56695 3705 56705 4025
rect 56665 3690 56705 3705
rect 56725 4025 56765 4040
rect 56725 3705 56735 4025
rect 56755 3705 56765 4025
rect 56725 3690 56765 3705
rect 57035 4025 57075 4040
rect 57035 3705 57045 4025
rect 57065 3705 57075 4025
rect 57035 3690 57075 3705
rect 57095 4025 57135 4040
rect 57095 3705 57105 4025
rect 57125 3705 57135 4025
rect 57095 3690 57135 3705
rect 57155 4025 57195 4040
rect 57155 3705 57165 4025
rect 57185 3705 57195 4025
rect 57155 3690 57195 3705
rect 57215 4025 57255 4040
rect 57215 3705 57225 4025
rect 57245 3705 57255 4025
rect 57215 3690 57255 3705
rect 57275 4025 57315 4040
rect 57275 3705 57285 4025
rect 57305 3705 57315 4025
rect 57275 3690 57315 3705
rect 57335 4025 57375 4040
rect 57335 3705 57345 4025
rect 57365 3705 57375 4025
rect 57335 3690 57375 3705
rect 57395 4025 57435 4040
rect 57395 3705 57405 4025
rect 57425 3705 57435 4025
rect 57395 3690 57435 3705
rect 57455 4025 57495 4040
rect 57455 3705 57465 4025
rect 57485 3705 57495 4025
rect 57455 3690 57495 3705
rect 57515 4025 57555 4040
rect 57515 3705 57525 4025
rect 57545 3705 57555 4025
rect 57515 3690 57555 3705
rect 57575 4025 57615 4040
rect 57575 3705 57585 4025
rect 57605 3705 57615 4025
rect 57575 3690 57615 3705
rect 57635 4025 57675 4040
rect 57635 3705 57645 4025
rect 57665 3705 57675 4025
rect 57635 3690 57675 3705
rect 57695 4025 57735 4040
rect 57695 3705 57705 4025
rect 57725 3705 57735 4025
rect 57695 3690 57735 3705
rect 57755 4025 57795 4040
rect 57755 3705 57765 4025
rect 57785 3705 57795 4025
rect 57755 3690 57795 3705
rect 58120 4025 58160 4040
rect 58120 3705 58130 4025
rect 58150 3705 58160 4025
rect 58120 3690 58160 3705
rect 58180 4025 58220 4040
rect 58180 3705 58190 4025
rect 58210 3705 58220 4025
rect 58180 3690 58220 3705
rect 58240 4025 58280 4040
rect 58240 3705 58250 4025
rect 58270 3705 58280 4025
rect 58240 3690 58280 3705
rect 58300 4025 58340 4040
rect 58300 3705 58310 4025
rect 58330 3705 58340 4025
rect 58300 3690 58340 3705
rect 58360 4025 58400 4040
rect 58360 3705 58370 4025
rect 58390 3705 58400 4025
rect 58360 3690 58400 3705
rect 58420 4025 58460 4040
rect 58420 3705 58430 4025
rect 58450 3705 58460 4025
rect 58420 3690 58460 3705
rect 58480 4025 58520 4040
rect 58480 3705 58490 4025
rect 58510 3705 58520 4025
rect 58480 3690 58520 3705
rect 58540 4025 58580 4040
rect 58540 3705 58550 4025
rect 58570 3705 58580 4025
rect 58540 3690 58580 3705
rect 58600 4025 58640 4040
rect 58600 3705 58610 4025
rect 58630 3705 58640 4025
rect 58600 3690 58640 3705
rect 58660 4025 58700 4040
rect 58660 3705 58670 4025
rect 58690 3705 58700 4025
rect 58660 3690 58700 3705
rect 58720 4025 58760 4040
rect 58720 3705 58730 4025
rect 58750 3705 58760 4025
rect 58720 3690 58760 3705
rect 58780 4025 58820 4040
rect 58780 3705 58790 4025
rect 58810 3705 58820 4025
rect 58780 3690 58820 3705
rect 58840 4025 58880 4040
rect 58840 3705 58850 4025
rect 58870 3705 58880 4025
rect 58840 3690 58880 3705
rect 54820 3250 54860 3265
rect 54820 2680 54830 3250
rect 54850 2680 54860 3250
rect 54820 2665 54860 2680
rect 54875 3250 54915 3265
rect 54875 2680 54885 3250
rect 54905 2680 54915 3250
rect 54875 2665 54915 2680
rect 54930 3250 54970 3265
rect 54930 2680 54940 3250
rect 54960 2680 54970 3250
rect 54930 2665 54970 2680
rect 54985 3250 55025 3265
rect 54985 2680 54995 3250
rect 55015 2680 55025 3250
rect 54985 2665 55025 2680
rect 55040 3250 55080 3265
rect 55040 2680 55050 3250
rect 55070 2680 55080 3250
rect 55040 2665 55080 2680
rect 55095 3250 55135 3265
rect 55095 2680 55105 3250
rect 55125 2680 55135 3250
rect 55095 2665 55135 2680
rect 55150 3250 55190 3265
rect 55150 2680 55160 3250
rect 55180 2680 55190 3250
rect 55150 2665 55190 2680
rect 55205 3250 55245 3265
rect 55205 2680 55215 3250
rect 55235 2680 55245 3250
rect 55205 2665 55245 2680
rect 55260 3250 55300 3265
rect 55260 2680 55270 3250
rect 55290 2680 55300 3250
rect 55260 2665 55300 2680
rect 55315 3250 55355 3265
rect 55315 2680 55325 3250
rect 55345 2680 55355 3250
rect 55315 2665 55355 2680
rect 55370 3250 55410 3265
rect 55370 2680 55380 3250
rect 55400 2680 55410 3250
rect 55370 2665 55410 2680
rect 55425 3250 55465 3265
rect 55425 2680 55435 3250
rect 55455 2680 55465 3250
rect 55425 2665 55465 2680
rect 55480 3250 55520 3265
rect 55480 2680 55490 3250
rect 55510 2680 55520 3250
rect 56275 3240 56315 3255
rect 56275 3220 56285 3240
rect 56305 3220 56315 3240
rect 56275 3205 56315 3220
rect 56330 3240 56370 3255
rect 56330 3220 56340 3240
rect 56360 3220 56370 3240
rect 56330 3205 56370 3220
rect 56385 3240 56425 3255
rect 56385 3220 56395 3240
rect 56415 3220 56425 3240
rect 56385 3205 56425 3220
rect 56440 3240 56480 3255
rect 56440 3220 56450 3240
rect 56470 3220 56480 3240
rect 56440 3205 56480 3220
rect 56495 3240 56535 3255
rect 56495 3220 56505 3240
rect 56525 3220 56535 3240
rect 56495 3205 56535 3220
rect 56550 3240 56590 3255
rect 56550 3220 56560 3240
rect 56580 3220 56590 3240
rect 56550 3205 56590 3220
rect 56605 3240 56645 3255
rect 56605 3220 56615 3240
rect 56635 3220 56645 3240
rect 56605 3205 56645 3220
rect 56660 3240 56700 3255
rect 56660 3220 56670 3240
rect 56690 3220 56700 3240
rect 56660 3205 56700 3220
rect 56715 3240 56755 3255
rect 56715 3220 56725 3240
rect 56745 3220 56755 3240
rect 56715 3205 56755 3220
rect 56770 3240 56810 3255
rect 56770 3220 56780 3240
rect 56800 3220 56810 3240
rect 56770 3205 56810 3220
rect 56825 3240 56865 3255
rect 56825 3220 56835 3240
rect 56855 3220 56865 3240
rect 56825 3205 56865 3220
rect 56880 3240 56920 3255
rect 56880 3220 56890 3240
rect 56910 3220 56920 3240
rect 56880 3205 56920 3220
rect 56935 3240 56975 3255
rect 56935 3220 56945 3240
rect 56965 3220 56975 3240
rect 56935 3205 56975 3220
rect 56990 3240 57030 3255
rect 56990 3220 57000 3240
rect 57020 3220 57030 3240
rect 56990 3205 57030 3220
rect 57045 3240 57085 3255
rect 57045 3220 57055 3240
rect 57075 3220 57085 3240
rect 57045 3205 57085 3220
rect 57100 3240 57140 3255
rect 57100 3220 57110 3240
rect 57130 3220 57140 3240
rect 57100 3205 57140 3220
rect 57155 3240 57195 3255
rect 57155 3220 57165 3240
rect 57185 3220 57195 3240
rect 57155 3205 57195 3220
rect 57210 3240 57250 3255
rect 57210 3220 57220 3240
rect 57240 3220 57250 3240
rect 57210 3205 57250 3220
rect 57265 3240 57305 3255
rect 57265 3220 57275 3240
rect 57295 3220 57305 3240
rect 57265 3205 57305 3220
rect 57320 3240 57360 3255
rect 57320 3220 57330 3240
rect 57350 3220 57360 3240
rect 57320 3205 57360 3220
rect 57375 3240 57415 3255
rect 57375 3220 57385 3240
rect 57405 3220 57415 3240
rect 57375 3205 57415 3220
rect 57430 3240 57470 3255
rect 57430 3220 57440 3240
rect 57460 3220 57470 3240
rect 57430 3205 57470 3220
rect 57485 3240 57525 3255
rect 57485 3220 57495 3240
rect 57515 3220 57525 3240
rect 57485 3205 57525 3220
rect 58280 3250 58320 3265
rect 56030 2930 56070 2945
rect 56030 2910 56040 2930
rect 56060 2910 56070 2930
rect 56030 2895 56070 2910
rect 56085 2930 56125 2945
rect 56085 2910 56095 2930
rect 56115 2910 56125 2930
rect 56085 2895 56125 2910
rect 56140 2930 56180 2945
rect 56140 2910 56150 2930
rect 56170 2910 56180 2930
rect 56140 2895 56180 2910
rect 56195 2930 56235 2945
rect 56195 2910 56205 2930
rect 56225 2910 56235 2930
rect 56195 2895 56235 2910
rect 56250 2930 56290 2945
rect 56250 2910 56260 2930
rect 56280 2910 56290 2930
rect 56250 2895 56290 2910
rect 56305 2930 56345 2945
rect 56305 2910 56315 2930
rect 56335 2910 56345 2930
rect 56305 2895 56345 2910
rect 56360 2930 56400 2945
rect 56360 2910 56370 2930
rect 56390 2910 56400 2930
rect 56360 2895 56400 2910
rect 56415 2930 56455 2945
rect 56415 2910 56425 2930
rect 56445 2910 56455 2930
rect 56415 2895 56455 2910
rect 56470 2930 56510 2945
rect 56470 2910 56480 2930
rect 56500 2910 56510 2930
rect 56470 2895 56510 2910
rect 56525 2930 56565 2945
rect 56525 2910 56535 2930
rect 56555 2910 56565 2930
rect 56525 2895 56565 2910
rect 56580 2930 56620 2945
rect 56580 2910 56590 2930
rect 56610 2910 56620 2930
rect 56580 2895 56620 2910
rect 56635 2930 56675 2945
rect 56635 2910 56645 2930
rect 56665 2910 56675 2930
rect 56635 2895 56675 2910
rect 56690 2930 56730 2945
rect 56690 2910 56700 2930
rect 56720 2910 56730 2930
rect 56690 2895 56730 2910
rect 57070 2930 57110 2945
rect 57070 2910 57080 2930
rect 57100 2910 57110 2930
rect 57070 2895 57110 2910
rect 57125 2930 57165 2945
rect 57125 2910 57135 2930
rect 57155 2910 57165 2930
rect 57125 2895 57165 2910
rect 57180 2930 57220 2945
rect 57180 2910 57190 2930
rect 57210 2910 57220 2930
rect 57180 2895 57220 2910
rect 57235 2930 57275 2945
rect 57235 2910 57245 2930
rect 57265 2910 57275 2930
rect 57235 2895 57275 2910
rect 57290 2930 57330 2945
rect 57290 2910 57300 2930
rect 57320 2910 57330 2930
rect 57290 2895 57330 2910
rect 57345 2930 57385 2945
rect 57345 2910 57355 2930
rect 57375 2910 57385 2930
rect 57345 2895 57385 2910
rect 57400 2930 57440 2945
rect 57400 2910 57410 2930
rect 57430 2910 57440 2930
rect 57400 2895 57440 2910
rect 57455 2930 57495 2945
rect 57455 2910 57465 2930
rect 57485 2910 57495 2930
rect 57455 2895 57495 2910
rect 57510 2930 57550 2945
rect 57510 2910 57520 2930
rect 57540 2910 57550 2930
rect 57510 2895 57550 2910
rect 57565 2930 57605 2945
rect 57565 2910 57575 2930
rect 57595 2910 57605 2930
rect 57565 2895 57605 2910
rect 57620 2930 57660 2945
rect 57620 2910 57630 2930
rect 57650 2910 57660 2930
rect 57620 2895 57660 2910
rect 57675 2930 57715 2945
rect 57675 2910 57685 2930
rect 57705 2910 57715 2930
rect 57675 2895 57715 2910
rect 57730 2930 57770 2945
rect 57730 2910 57740 2930
rect 57760 2910 57770 2930
rect 57730 2895 57770 2910
rect 55480 2665 55520 2680
rect 58280 2680 58290 3250
rect 58310 2680 58320 3250
rect 58280 2665 58320 2680
rect 58335 3250 58375 3265
rect 58335 2680 58345 3250
rect 58365 2680 58375 3250
rect 58335 2665 58375 2680
rect 58390 3250 58430 3265
rect 58390 2680 58400 3250
rect 58420 2680 58430 3250
rect 58390 2665 58430 2680
rect 58445 3250 58485 3265
rect 58445 2680 58455 3250
rect 58475 2680 58485 3250
rect 58445 2665 58485 2680
rect 58500 3250 58540 3265
rect 58500 2680 58510 3250
rect 58530 2680 58540 3250
rect 58500 2665 58540 2680
rect 58555 3250 58595 3265
rect 58555 2680 58565 3250
rect 58585 2680 58595 3250
rect 58555 2665 58595 2680
rect 58610 3250 58650 3265
rect 58610 2680 58620 3250
rect 58640 2680 58650 3250
rect 58610 2665 58650 2680
rect 58665 3250 58705 3265
rect 58665 2680 58675 3250
rect 58695 2680 58705 3250
rect 58665 2665 58705 2680
rect 58720 3250 58760 3265
rect 58720 2680 58730 3250
rect 58750 2680 58760 3250
rect 58720 2665 58760 2680
rect 58775 3250 58815 3265
rect 58775 2680 58785 3250
rect 58805 2680 58815 3250
rect 58775 2665 58815 2680
rect 58830 3250 58870 3265
rect 58830 2680 58840 3250
rect 58860 2680 58870 3250
rect 58830 2665 58870 2680
rect 58885 3250 58925 3265
rect 58885 2680 58895 3250
rect 58915 2680 58925 3250
rect 58885 2665 58925 2680
rect 58940 3250 58980 3265
rect 58940 2680 58950 3250
rect 58970 2680 58980 3250
rect 58940 2665 58980 2680
rect 54820 2150 54860 2165
rect 54820 1980 54830 2150
rect 54850 1980 54860 2150
rect 54820 1965 54860 1980
rect 54875 2150 54915 2165
rect 54875 1980 54885 2150
rect 54905 1980 54915 2150
rect 54875 1965 54915 1980
rect 54930 2150 54970 2165
rect 54930 1980 54940 2150
rect 54960 1980 54970 2150
rect 54930 1965 54970 1980
rect 54985 2150 55025 2165
rect 54985 1980 54995 2150
rect 55015 1980 55025 2150
rect 54985 1965 55025 1980
rect 55040 2150 55080 2165
rect 55040 1980 55050 2150
rect 55070 1980 55080 2150
rect 55040 1965 55080 1980
rect 55095 2150 55135 2165
rect 55095 1980 55105 2150
rect 55125 1980 55135 2150
rect 55095 1965 55135 1980
rect 55150 2150 55190 2165
rect 55150 1980 55160 2150
rect 55180 1980 55190 2150
rect 55150 1965 55190 1980
rect 55205 2150 55245 2165
rect 55205 1980 55215 2150
rect 55235 1980 55245 2150
rect 55205 1965 55245 1980
rect 55260 2150 55300 2165
rect 55260 1980 55270 2150
rect 55290 1980 55300 2150
rect 55260 1965 55300 1980
rect 55315 2150 55355 2165
rect 55315 1980 55325 2150
rect 55345 1980 55355 2150
rect 55315 1965 55355 1980
rect 55370 2150 55410 2165
rect 55370 1980 55380 2150
rect 55400 1980 55410 2150
rect 55370 1965 55410 1980
rect 55425 2150 55465 2165
rect 55425 1980 55435 2150
rect 55455 1980 55465 2150
rect 55425 1965 55465 1980
rect 55480 2150 55520 2165
rect 55480 1980 55490 2150
rect 55510 1980 55520 2150
rect 58280 2150 58320 2165
rect 55480 1965 55520 1980
rect 58280 1980 58290 2150
rect 58310 1980 58320 2150
rect 58280 1965 58320 1980
rect 58335 2150 58375 2165
rect 58335 1980 58345 2150
rect 58365 1980 58375 2150
rect 58335 1965 58375 1980
rect 58390 2150 58430 2165
rect 58390 1980 58400 2150
rect 58420 1980 58430 2150
rect 58390 1965 58430 1980
rect 58445 2150 58485 2165
rect 58445 1980 58455 2150
rect 58475 1980 58485 2150
rect 58445 1965 58485 1980
rect 58500 2150 58540 2165
rect 58500 1980 58510 2150
rect 58530 1980 58540 2150
rect 58500 1965 58540 1980
rect 58555 2150 58595 2165
rect 58555 1980 58565 2150
rect 58585 1980 58595 2150
rect 58555 1965 58595 1980
rect 58610 2150 58650 2165
rect 58610 1980 58620 2150
rect 58640 1980 58650 2150
rect 58610 1965 58650 1980
rect 58665 2150 58705 2165
rect 58665 1980 58675 2150
rect 58695 1980 58705 2150
rect 58665 1965 58705 1980
rect 58720 2150 58760 2165
rect 58720 1980 58730 2150
rect 58750 1980 58760 2150
rect 58720 1965 58760 1980
rect 58775 2150 58815 2165
rect 58775 1980 58785 2150
rect 58805 1980 58815 2150
rect 58775 1965 58815 1980
rect 58830 2150 58870 2165
rect 58830 1980 58840 2150
rect 58860 1980 58870 2150
rect 58830 1965 58870 1980
rect 58885 2150 58925 2165
rect 58885 1980 58895 2150
rect 58915 1980 58925 2150
rect 58885 1965 58925 1980
rect 58940 2150 58980 2165
rect 58940 1980 58950 2150
rect 58970 1980 58980 2150
rect 58940 1965 58980 1980
<< ndiffc >>
rect 56780 2350 56800 2570
rect 56835 2350 56855 2570
rect 56890 2350 56910 2570
rect 56945 2350 56965 2570
rect 57000 2350 57020 2570
rect 56040 2045 56060 2165
rect 56095 2045 56115 2165
rect 56150 2045 56170 2165
rect 56205 2045 56225 2165
rect 56260 2045 56280 2165
rect 56315 2045 56335 2165
rect 56370 2045 56390 2165
rect 56425 2045 56445 2165
rect 56480 2045 56500 2165
rect 56535 2045 56555 2165
rect 56590 2045 56610 2165
rect 56645 2045 56665 2165
rect 56700 2045 56720 2165
rect 57080 2045 57100 2165
rect 57135 2045 57155 2165
rect 57190 2045 57210 2165
rect 57245 2045 57265 2165
rect 57300 2045 57320 2165
rect 57355 2045 57375 2165
rect 57410 2045 57430 2165
rect 57465 2045 57485 2165
rect 57520 2045 57540 2165
rect 57575 2045 57595 2165
rect 57630 2045 57650 2165
rect 57685 2045 57705 2165
rect 57740 2045 57760 2165
rect 54830 1440 54850 1710
rect 54885 1440 54905 1710
rect 54940 1440 54960 1710
rect 54995 1440 55015 1710
rect 55050 1440 55070 1710
rect 55105 1440 55125 1710
rect 55160 1440 55180 1710
rect 55215 1440 55235 1710
rect 55270 1440 55290 1710
rect 55325 1440 55345 1710
rect 55380 1440 55400 1710
rect 55435 1440 55455 1710
rect 55490 1440 55510 1710
rect 56040 1575 56060 1695
rect 56095 1575 56115 1695
rect 56150 1575 56170 1695
rect 56205 1575 56225 1695
rect 56260 1575 56280 1695
rect 56315 1575 56335 1695
rect 56370 1575 56390 1695
rect 56425 1575 56445 1695
rect 56480 1575 56500 1695
rect 56535 1575 56555 1695
rect 56590 1575 56610 1695
rect 56645 1575 56665 1695
rect 56700 1575 56720 1695
rect 56780 1575 56800 1695
rect 56835 1575 56855 1695
rect 56890 1575 56910 1695
rect 56945 1575 56965 1695
rect 57000 1575 57020 1695
rect 57080 1575 57100 1695
rect 57135 1575 57155 1695
rect 57190 1575 57210 1695
rect 57245 1575 57265 1695
rect 57300 1575 57320 1695
rect 57355 1575 57375 1695
rect 57410 1575 57430 1695
rect 57465 1575 57485 1695
rect 57520 1575 57540 1695
rect 57575 1575 57595 1695
rect 57630 1575 57650 1695
rect 57685 1575 57705 1695
rect 57740 1575 57760 1695
rect 58290 1440 58310 1710
rect 58345 1440 58365 1710
rect 58400 1440 58420 1710
rect 58455 1440 58475 1710
rect 58510 1440 58530 1710
rect 58565 1440 58585 1710
rect 58620 1440 58640 1710
rect 58675 1440 58695 1710
rect 58730 1440 58750 1710
rect 58785 1440 58805 1710
rect 58840 1440 58860 1710
rect 58895 1440 58915 1710
rect 58950 1440 58970 1710
rect 54840 370 54860 1040
rect 54940 370 54960 1040
rect 55040 370 55060 1040
rect 55140 370 55160 1040
rect 55240 370 55260 1040
rect 55340 370 55360 1040
rect 55440 370 55460 1040
rect 56230 775 56250 995
rect 56285 775 56305 995
rect 56340 775 56360 995
rect 56395 775 56415 995
rect 56450 775 56470 995
rect 56505 775 56525 995
rect 56560 775 56580 995
rect 56615 775 56635 995
rect 56670 775 56690 995
rect 56725 775 56745 995
rect 56780 775 56800 995
rect 56835 775 56855 995
rect 56890 775 56910 995
rect 56945 775 56965 995
rect 57000 775 57020 995
rect 57055 775 57075 995
rect 57110 775 57130 995
rect 57165 775 57185 995
rect 57220 775 57240 995
rect 57275 775 57295 995
rect 57330 775 57350 995
rect 57385 775 57405 995
rect 57440 775 57460 995
rect 57495 775 57515 995
rect 56440 410 56460 530
rect 56495 410 56515 530
rect 56550 410 56570 530
rect 56605 410 56625 530
rect 56660 410 56680 530
rect 56715 410 56735 530
rect 56770 410 56790 530
rect 56880 410 56900 530
rect 57220 410 57240 530
rect 58340 370 58360 1040
rect 58440 370 58460 1040
rect 58540 370 58560 1040
rect 58640 370 58660 1040
rect 58740 370 58760 1040
rect 58840 370 58860 1040
rect 58940 370 58960 1040
<< pdiffc >>
rect 56095 4580 56115 4900
rect 56155 4580 56175 4900
rect 56215 4580 56235 4900
rect 56275 4580 56295 4900
rect 56565 4580 56585 4730
rect 56625 4580 56645 4730
rect 56685 4580 56705 4730
rect 56745 4580 56765 4730
rect 57035 4580 57055 4900
rect 57095 4580 57115 4900
rect 57155 4580 57175 4900
rect 57215 4580 57235 4900
rect 57505 4580 57525 4900
rect 57565 4580 57585 4900
rect 57625 4580 57645 4900
rect 57685 4580 57705 4900
rect 54930 3705 54950 4025
rect 54990 3705 55010 4025
rect 55050 3705 55070 4025
rect 55110 3705 55130 4025
rect 55170 3705 55190 4025
rect 55230 3705 55250 4025
rect 55290 3705 55310 4025
rect 55350 3705 55370 4025
rect 55410 3705 55430 4025
rect 55470 3705 55490 4025
rect 55530 3705 55550 4025
rect 55590 3705 55610 4025
rect 55650 3705 55670 4025
rect 56015 3705 56035 4025
rect 56075 3705 56095 4025
rect 56135 3705 56155 4025
rect 56195 3705 56215 4025
rect 56255 3705 56275 4025
rect 56315 3705 56335 4025
rect 56375 3705 56395 4025
rect 56435 3705 56455 4025
rect 56495 3705 56515 4025
rect 56555 3705 56575 4025
rect 56615 3705 56635 4025
rect 56675 3705 56695 4025
rect 56735 3705 56755 4025
rect 57045 3705 57065 4025
rect 57105 3705 57125 4025
rect 57165 3705 57185 4025
rect 57225 3705 57245 4025
rect 57285 3705 57305 4025
rect 57345 3705 57365 4025
rect 57405 3705 57425 4025
rect 57465 3705 57485 4025
rect 57525 3705 57545 4025
rect 57585 3705 57605 4025
rect 57645 3705 57665 4025
rect 57705 3705 57725 4025
rect 57765 3705 57785 4025
rect 58130 3705 58150 4025
rect 58190 3705 58210 4025
rect 58250 3705 58270 4025
rect 58310 3705 58330 4025
rect 58370 3705 58390 4025
rect 58430 3705 58450 4025
rect 58490 3705 58510 4025
rect 58550 3705 58570 4025
rect 58610 3705 58630 4025
rect 58670 3705 58690 4025
rect 58730 3705 58750 4025
rect 58790 3705 58810 4025
rect 58850 3705 58870 4025
rect 54830 2680 54850 3250
rect 54885 2680 54905 3250
rect 54940 2680 54960 3250
rect 54995 2680 55015 3250
rect 55050 2680 55070 3250
rect 55105 2680 55125 3250
rect 55160 2680 55180 3250
rect 55215 2680 55235 3250
rect 55270 2680 55290 3250
rect 55325 2680 55345 3250
rect 55380 2680 55400 3250
rect 55435 2680 55455 3250
rect 55490 2680 55510 3250
rect 56285 3220 56305 3240
rect 56340 3220 56360 3240
rect 56395 3220 56415 3240
rect 56450 3220 56470 3240
rect 56505 3220 56525 3240
rect 56560 3220 56580 3240
rect 56615 3220 56635 3240
rect 56670 3220 56690 3240
rect 56725 3220 56745 3240
rect 56780 3220 56800 3240
rect 56835 3220 56855 3240
rect 56890 3220 56910 3240
rect 56945 3220 56965 3240
rect 57000 3220 57020 3240
rect 57055 3220 57075 3240
rect 57110 3220 57130 3240
rect 57165 3220 57185 3240
rect 57220 3220 57240 3240
rect 57275 3220 57295 3240
rect 57330 3220 57350 3240
rect 57385 3220 57405 3240
rect 57440 3220 57460 3240
rect 57495 3220 57515 3240
rect 56040 2910 56060 2930
rect 56095 2910 56115 2930
rect 56150 2910 56170 2930
rect 56205 2910 56225 2930
rect 56260 2910 56280 2930
rect 56315 2910 56335 2930
rect 56370 2910 56390 2930
rect 56425 2910 56445 2930
rect 56480 2910 56500 2930
rect 56535 2910 56555 2930
rect 56590 2910 56610 2930
rect 56645 2910 56665 2930
rect 56700 2910 56720 2930
rect 57080 2910 57100 2930
rect 57135 2910 57155 2930
rect 57190 2910 57210 2930
rect 57245 2910 57265 2930
rect 57300 2910 57320 2930
rect 57355 2910 57375 2930
rect 57410 2910 57430 2930
rect 57465 2910 57485 2930
rect 57520 2910 57540 2930
rect 57575 2910 57595 2930
rect 57630 2910 57650 2930
rect 57685 2910 57705 2930
rect 57740 2910 57760 2930
rect 58290 2680 58310 3250
rect 58345 2680 58365 3250
rect 58400 2680 58420 3250
rect 58455 2680 58475 3250
rect 58510 2680 58530 3250
rect 58565 2680 58585 3250
rect 58620 2680 58640 3250
rect 58675 2680 58695 3250
rect 58730 2680 58750 3250
rect 58785 2680 58805 3250
rect 58840 2680 58860 3250
rect 58895 2680 58915 3250
rect 58950 2680 58970 3250
rect 54830 1980 54850 2150
rect 54885 1980 54905 2150
rect 54940 1980 54960 2150
rect 54995 1980 55015 2150
rect 55050 1980 55070 2150
rect 55105 1980 55125 2150
rect 55160 1980 55180 2150
rect 55215 1980 55235 2150
rect 55270 1980 55290 2150
rect 55325 1980 55345 2150
rect 55380 1980 55400 2150
rect 55435 1980 55455 2150
rect 55490 1980 55510 2150
rect 58290 1980 58310 2150
rect 58345 1980 58365 2150
rect 58400 1980 58420 2150
rect 58455 1980 58475 2150
rect 58510 1980 58530 2150
rect 58565 1980 58585 2150
rect 58620 1980 58640 2150
rect 58675 1980 58695 2150
rect 58730 1980 58750 2150
rect 58785 1980 58805 2150
rect 58840 1980 58860 2150
rect 58895 1980 58915 2150
rect 58950 1980 58970 2150
<< psubdiff >>
rect 56730 2570 56770 2585
rect 56730 2350 56740 2570
rect 56760 2350 56770 2570
rect 56730 2335 56770 2350
rect 57030 2570 57070 2585
rect 57030 2350 57040 2570
rect 57060 2350 57070 2570
rect 57030 2335 57070 2350
rect 55990 2165 56030 2180
rect 55990 2045 56000 2165
rect 56020 2045 56030 2165
rect 55990 2030 56030 2045
rect 56730 2165 56770 2180
rect 56730 2045 56740 2165
rect 56760 2045 56770 2165
rect 56730 2030 56770 2045
rect 57030 2165 57070 2180
rect 57030 2045 57040 2165
rect 57060 2045 57070 2165
rect 57030 2030 57070 2045
rect 57770 2165 57810 2180
rect 57770 2045 57780 2165
rect 57800 2045 57810 2165
rect 57770 2030 57810 2045
rect 54780 1710 54820 1725
rect 54780 1440 54790 1710
rect 54810 1440 54820 1710
rect 54780 1425 54820 1440
rect 55520 1710 55560 1725
rect 58240 1710 58280 1725
rect 55520 1440 55530 1710
rect 55550 1440 55560 1710
rect 55990 1695 56030 1710
rect 55990 1575 56000 1695
rect 56020 1575 56030 1695
rect 55990 1560 56030 1575
rect 56730 1695 56770 1710
rect 56730 1575 56740 1695
rect 56760 1575 56770 1695
rect 56730 1560 56770 1575
rect 57030 1695 57070 1710
rect 57030 1575 57040 1695
rect 57060 1575 57070 1695
rect 57030 1560 57070 1575
rect 57770 1695 57810 1710
rect 57770 1575 57780 1695
rect 57800 1575 57810 1695
rect 57770 1560 57810 1575
rect 55520 1425 55560 1440
rect 58240 1440 58250 1710
rect 58270 1440 58280 1710
rect 58240 1425 58280 1440
rect 58980 1710 59020 1725
rect 58980 1440 58990 1710
rect 59010 1440 59020 1710
rect 58980 1425 59020 1440
rect 54790 1040 54830 1055
rect 54790 370 54800 1040
rect 54820 370 54830 1040
rect 54790 355 54830 370
rect 55470 1040 55510 1055
rect 55470 370 55480 1040
rect 55500 370 55510 1040
rect 58290 1040 58330 1055
rect 56180 995 56220 1010
rect 56180 775 56190 995
rect 56210 775 56220 995
rect 56180 760 56220 775
rect 57525 995 57565 1010
rect 57525 775 57535 995
rect 57555 775 57565 995
rect 57525 760 57565 775
rect 56390 530 56430 545
rect 56390 410 56400 530
rect 56420 410 56430 530
rect 56390 395 56430 410
rect 56800 530 56840 545
rect 56800 410 56810 530
rect 56830 410 56840 530
rect 56800 395 56840 410
rect 55470 355 55510 370
rect 58290 370 58300 1040
rect 58320 370 58330 1040
rect 58290 355 58330 370
rect 58970 1040 59010 1055
rect 58970 370 58980 1040
rect 59000 370 59010 1040
rect 58970 355 59010 370
<< nsubdiff >>
rect 56045 4900 56085 4915
rect 56045 4580 56055 4900
rect 56075 4580 56085 4900
rect 56045 4565 56085 4580
rect 56305 4900 56345 4915
rect 56305 4580 56315 4900
rect 56335 4580 56345 4900
rect 56985 4900 57025 4915
rect 56305 4565 56345 4580
rect 56515 4730 56555 4745
rect 56515 4580 56525 4730
rect 56545 4580 56555 4730
rect 56515 4565 56555 4580
rect 56775 4730 56815 4745
rect 56775 4580 56785 4730
rect 56805 4580 56815 4730
rect 56775 4565 56815 4580
rect 56985 4580 56995 4900
rect 57015 4580 57025 4900
rect 56985 4565 57025 4580
rect 57245 4900 57285 4915
rect 57245 4580 57255 4900
rect 57275 4580 57285 4900
rect 57245 4565 57285 4580
rect 57455 4900 57495 4915
rect 57455 4580 57465 4900
rect 57485 4580 57495 4900
rect 57455 4565 57495 4580
rect 57715 4900 57755 4915
rect 57715 4580 57725 4900
rect 57745 4580 57755 4900
rect 57715 4565 57755 4580
rect 54880 4025 54920 4040
rect 54880 3705 54890 4025
rect 54910 3705 54920 4025
rect 54880 3690 54920 3705
rect 55680 4025 55720 4040
rect 55680 3705 55690 4025
rect 55710 3705 55720 4025
rect 55680 3690 55720 3705
rect 55965 4025 56005 4040
rect 55965 3705 55975 4025
rect 55995 3705 56005 4025
rect 55965 3690 56005 3705
rect 56765 4025 56805 4040
rect 56765 3705 56775 4025
rect 56795 3705 56805 4025
rect 56765 3690 56805 3705
rect 56995 4025 57035 4040
rect 56995 3705 57005 4025
rect 57025 3705 57035 4025
rect 56995 3690 57035 3705
rect 57795 4025 57835 4040
rect 57795 3705 57805 4025
rect 57825 3705 57835 4025
rect 57795 3690 57835 3705
rect 58080 4025 58120 4040
rect 58080 3705 58090 4025
rect 58110 3705 58120 4025
rect 58080 3690 58120 3705
rect 58880 4025 58920 4040
rect 58880 3705 58890 4025
rect 58910 3705 58920 4025
rect 58880 3690 58920 3705
rect 54780 3250 54820 3265
rect 54780 2680 54790 3250
rect 54810 2680 54820 3250
rect 54780 2665 54820 2680
rect 55520 3250 55560 3265
rect 55520 2680 55530 3250
rect 55550 2680 55560 3250
rect 56235 3240 56275 3255
rect 56235 3220 56245 3240
rect 56265 3220 56275 3240
rect 56235 3205 56275 3220
rect 57525 3240 57565 3255
rect 57525 3220 57535 3240
rect 57555 3220 57565 3240
rect 57525 3205 57565 3220
rect 58240 3250 58280 3265
rect 55990 2930 56030 2945
rect 55990 2910 56000 2930
rect 56020 2910 56030 2930
rect 55990 2895 56030 2910
rect 56730 2930 56770 2945
rect 56730 2910 56740 2930
rect 56760 2910 56770 2930
rect 56730 2895 56770 2910
rect 57030 2930 57070 2945
rect 57030 2910 57040 2930
rect 57060 2910 57070 2930
rect 57030 2895 57070 2910
rect 57770 2930 57810 2945
rect 57770 2910 57780 2930
rect 57800 2910 57810 2930
rect 57770 2895 57810 2910
rect 55520 2665 55560 2680
rect 58240 2680 58250 3250
rect 58270 2680 58280 3250
rect 58240 2665 58280 2680
rect 58980 3250 59020 3265
rect 58980 2680 58990 3250
rect 59010 2680 59020 3250
rect 58980 2665 59020 2680
rect 54780 2150 54820 2165
rect 54780 1980 54790 2150
rect 54810 1980 54820 2150
rect 54780 1965 54820 1980
rect 55520 2150 55560 2165
rect 55520 1980 55530 2150
rect 55550 1980 55560 2150
rect 58240 2150 58280 2165
rect 55520 1965 55560 1980
rect 58240 1980 58250 2150
rect 58270 1980 58280 2150
rect 58240 1965 58280 1980
rect 58980 2150 59020 2165
rect 58980 1980 58990 2150
rect 59010 1980 59020 2150
rect 58980 1965 59020 1980
<< psubdiffcont >>
rect 56740 2350 56760 2570
rect 57040 2350 57060 2570
rect 56000 2045 56020 2165
rect 56740 2045 56760 2165
rect 57040 2045 57060 2165
rect 57780 2045 57800 2165
rect 54790 1440 54810 1710
rect 55530 1440 55550 1710
rect 56000 1575 56020 1695
rect 56740 1575 56760 1695
rect 57040 1575 57060 1695
rect 57780 1575 57800 1695
rect 58250 1440 58270 1710
rect 58990 1440 59010 1710
rect 54800 370 54820 1040
rect 55480 370 55500 1040
rect 56190 775 56210 995
rect 57535 775 57555 995
rect 56400 410 56420 530
rect 56810 410 56830 530
rect 58300 370 58320 1040
rect 58980 370 59000 1040
<< nsubdiffcont >>
rect 56055 4580 56075 4900
rect 56315 4580 56335 4900
rect 56525 4580 56545 4730
rect 56785 4580 56805 4730
rect 56995 4580 57015 4900
rect 57255 4580 57275 4900
rect 57465 4580 57485 4900
rect 57725 4580 57745 4900
rect 54890 3705 54910 4025
rect 55690 3705 55710 4025
rect 55975 3705 55995 4025
rect 56775 3705 56795 4025
rect 57005 3705 57025 4025
rect 57805 3705 57825 4025
rect 58090 3705 58110 4025
rect 58890 3705 58910 4025
rect 54790 2680 54810 3250
rect 55530 2680 55550 3250
rect 56245 3220 56265 3240
rect 57535 3220 57555 3240
rect 56000 2910 56020 2930
rect 56740 2910 56760 2930
rect 57040 2910 57060 2930
rect 57780 2910 57800 2930
rect 58250 2680 58270 3250
rect 58990 2680 59010 3250
rect 54790 1980 54810 2150
rect 55530 1980 55550 2150
rect 58250 1980 58270 2150
rect 58990 1980 59010 2150
<< poly >>
rect 56085 4960 56125 4970
rect 56085 4940 56095 4960
rect 56115 4945 56125 4960
rect 56265 4960 56305 4970
rect 56265 4945 56275 4960
rect 56115 4940 56145 4945
rect 56085 4930 56145 4940
rect 56245 4940 56275 4945
rect 56295 4940 56305 4960
rect 56245 4930 56305 4940
rect 57025 4960 57065 4970
rect 57025 4940 57035 4960
rect 57055 4945 57065 4960
rect 57205 4960 57245 4970
rect 57205 4945 57215 4960
rect 57055 4940 57085 4945
rect 57025 4930 57085 4940
rect 57185 4940 57215 4945
rect 57235 4940 57245 4960
rect 57185 4930 57245 4940
rect 57495 4960 57535 4970
rect 57495 4940 57505 4960
rect 57525 4945 57535 4960
rect 57675 4960 57715 4970
rect 57675 4945 57685 4960
rect 57525 4940 57555 4945
rect 57495 4930 57555 4940
rect 57655 4940 57685 4945
rect 57705 4940 57715 4960
rect 57655 4930 57715 4940
rect 56125 4915 56145 4930
rect 56185 4915 56205 4930
rect 56245 4915 56265 4930
rect 57065 4915 57085 4930
rect 57125 4915 57145 4930
rect 57185 4915 57205 4930
rect 57535 4915 57555 4930
rect 57595 4915 57615 4930
rect 57655 4915 57675 4930
rect 56555 4790 56595 4800
rect 56555 4770 56565 4790
rect 56585 4775 56595 4790
rect 56735 4790 56775 4800
rect 56735 4775 56745 4790
rect 56585 4770 56615 4775
rect 56555 4760 56615 4770
rect 56715 4770 56745 4775
rect 56765 4770 56775 4790
rect 56715 4760 56775 4770
rect 56595 4745 56615 4760
rect 56655 4745 56675 4760
rect 56715 4745 56735 4760
rect 56125 4550 56145 4565
rect 56185 4520 56205 4565
rect 56245 4550 56265 4565
rect 56595 4550 56615 4565
rect 56655 4520 56675 4565
rect 56715 4550 56735 4565
rect 57065 4550 57085 4565
rect 56150 4510 56205 4520
rect 56150 4490 56160 4510
rect 56180 4490 56205 4510
rect 56150 4480 56205 4490
rect 56630 4510 56675 4520
rect 56630 4490 56635 4510
rect 56655 4505 56675 4510
rect 57125 4520 57145 4565
rect 57185 4550 57205 4565
rect 57535 4550 57555 4565
rect 57125 4510 57170 4520
rect 57595 4510 57615 4565
rect 57655 4550 57675 4565
rect 57125 4505 57145 4510
rect 56655 4490 56660 4505
rect 56630 4480 56660 4490
rect 57140 4490 57145 4505
rect 57165 4490 57170 4510
rect 57140 4480 57170 4490
rect 57576 4500 57615 4510
rect 57576 4480 57581 4500
rect 57601 4495 57615 4500
rect 57601 4480 57606 4495
rect 57576 4470 57606 4480
rect 54960 4040 54980 4055
rect 55020 4040 55040 4055
rect 55080 4040 55100 4055
rect 55140 4040 55160 4055
rect 55200 4040 55220 4055
rect 55260 4040 55280 4055
rect 55320 4040 55340 4055
rect 55380 4040 55400 4055
rect 55440 4040 55460 4055
rect 55500 4040 55520 4055
rect 55560 4040 55580 4055
rect 55620 4040 55640 4055
rect 56045 4040 56065 4055
rect 56105 4040 56125 4055
rect 56165 4040 56185 4055
rect 56225 4040 56245 4055
rect 56285 4040 56305 4055
rect 56345 4040 56365 4055
rect 56405 4040 56425 4055
rect 56465 4040 56485 4055
rect 56525 4040 56545 4055
rect 56585 4040 56605 4055
rect 56645 4040 56665 4055
rect 56705 4040 56725 4055
rect 57075 4040 57095 4055
rect 57135 4040 57155 4055
rect 57195 4040 57215 4055
rect 57255 4040 57275 4055
rect 57315 4040 57335 4055
rect 57375 4040 57395 4055
rect 57435 4040 57455 4055
rect 57495 4040 57515 4055
rect 57555 4040 57575 4055
rect 57615 4040 57635 4055
rect 57675 4040 57695 4055
rect 57735 4040 57755 4055
rect 58160 4040 58180 4055
rect 58220 4040 58240 4055
rect 58280 4040 58300 4055
rect 58340 4040 58360 4055
rect 58400 4040 58420 4055
rect 58460 4040 58480 4055
rect 58520 4040 58540 4055
rect 58580 4040 58600 4055
rect 58640 4040 58660 4055
rect 58700 4040 58720 4055
rect 58760 4040 58780 4055
rect 58820 4040 58840 4055
rect 54960 3675 54980 3690
rect 54925 3665 54980 3675
rect 55020 3680 55040 3690
rect 55080 3680 55100 3690
rect 55140 3680 55160 3690
rect 55200 3680 55220 3690
rect 55260 3680 55280 3690
rect 55320 3680 55340 3690
rect 55380 3680 55400 3690
rect 55440 3680 55460 3690
rect 55500 3680 55520 3690
rect 55560 3680 55580 3690
rect 55020 3665 55580 3680
rect 55620 3675 55640 3690
rect 56045 3675 56065 3690
rect 55620 3665 55675 3675
rect 54925 3645 54930 3665
rect 54950 3660 54980 3665
rect 54950 3645 54955 3660
rect 54925 3635 54955 3645
rect 55285 3645 55290 3665
rect 55310 3645 55315 3665
rect 55620 3660 55650 3665
rect 55285 3635 55315 3645
rect 55645 3645 55650 3660
rect 55670 3645 55675 3665
rect 55645 3635 55675 3645
rect 56010 3665 56065 3675
rect 56105 3680 56125 3690
rect 56165 3680 56185 3690
rect 56225 3680 56245 3690
rect 56285 3680 56305 3690
rect 56345 3680 56365 3690
rect 56405 3680 56425 3690
rect 56465 3680 56485 3690
rect 56525 3680 56545 3690
rect 56585 3680 56605 3690
rect 56645 3680 56665 3690
rect 56105 3665 56665 3680
rect 56705 3675 56725 3690
rect 57075 3675 57095 3690
rect 56705 3665 56760 3675
rect 56010 3645 56015 3665
rect 56035 3660 56065 3665
rect 56035 3645 56040 3660
rect 56010 3635 56040 3645
rect 56370 3645 56375 3665
rect 56395 3645 56400 3665
rect 56705 3660 56735 3665
rect 56370 3635 56400 3645
rect 56730 3645 56735 3660
rect 56755 3645 56760 3665
rect 56730 3635 56760 3645
rect 57040 3665 57095 3675
rect 57135 3680 57155 3690
rect 57195 3680 57215 3690
rect 57255 3680 57275 3690
rect 57315 3680 57335 3690
rect 57375 3680 57395 3690
rect 57435 3680 57455 3690
rect 57495 3680 57515 3690
rect 57555 3680 57575 3690
rect 57615 3680 57635 3690
rect 57675 3680 57695 3690
rect 57135 3665 57695 3680
rect 57735 3675 57755 3690
rect 58160 3675 58180 3690
rect 57735 3665 57790 3675
rect 57040 3645 57045 3665
rect 57065 3660 57095 3665
rect 57065 3645 57070 3660
rect 57040 3635 57070 3645
rect 57400 3645 57405 3665
rect 57425 3645 57430 3665
rect 57735 3660 57765 3665
rect 57400 3635 57430 3645
rect 57760 3645 57765 3660
rect 57785 3645 57790 3665
rect 57760 3635 57790 3645
rect 58125 3665 58180 3675
rect 58220 3680 58240 3690
rect 58280 3680 58300 3690
rect 58340 3680 58360 3690
rect 58400 3680 58420 3690
rect 58460 3680 58480 3690
rect 58520 3680 58540 3690
rect 58580 3680 58600 3690
rect 58640 3680 58660 3690
rect 58700 3680 58720 3690
rect 58760 3680 58780 3690
rect 58220 3665 58780 3680
rect 58820 3675 58840 3690
rect 58820 3665 58875 3675
rect 58125 3645 58130 3665
rect 58150 3660 58180 3665
rect 58150 3645 58155 3660
rect 58125 3635 58155 3645
rect 58485 3645 58490 3665
rect 58510 3645 58515 3665
rect 58820 3660 58850 3665
rect 58485 3635 58515 3645
rect 58845 3645 58850 3660
rect 58870 3645 58875 3665
rect 58845 3635 58875 3645
rect 55290 3565 55310 3635
rect 56375 3610 56395 3635
rect 57405 3610 57425 3635
rect 56365 3600 56405 3610
rect 56365 3580 56375 3600
rect 56395 3580 56405 3600
rect 56365 3570 56405 3580
rect 57395 3600 57435 3610
rect 57395 3580 57405 3600
rect 57425 3580 57435 3600
rect 57395 3570 57435 3580
rect 58490 3565 58510 3635
rect 55280 3555 55320 3565
rect 55280 3535 55290 3555
rect 55310 3535 55320 3555
rect 55280 3525 55320 3535
rect 58480 3555 58520 3565
rect 58480 3535 58490 3555
rect 58510 3535 58520 3555
rect 58480 3525 58520 3535
rect 54825 3310 54855 3320
rect 54825 3290 54830 3310
rect 54850 3295 54855 3310
rect 55485 3310 55515 3320
rect 55485 3295 55490 3310
rect 54850 3290 54875 3295
rect 54825 3280 54875 3290
rect 55465 3290 55490 3295
rect 55510 3290 55515 3310
rect 55465 3280 55515 3290
rect 58285 3310 58315 3320
rect 58285 3290 58290 3310
rect 58310 3295 58315 3310
rect 58945 3310 58975 3320
rect 58945 3295 58950 3310
rect 58310 3290 58335 3295
rect 58285 3280 58335 3290
rect 58925 3290 58950 3295
rect 58970 3290 58975 3310
rect 58925 3280 58975 3290
rect 54860 3265 54875 3280
rect 54915 3265 54930 3280
rect 54970 3265 54985 3280
rect 55025 3265 55040 3280
rect 55080 3265 55095 3280
rect 55135 3265 55150 3280
rect 55190 3265 55205 3280
rect 55245 3265 55260 3280
rect 55300 3265 55315 3280
rect 55355 3265 55370 3280
rect 55410 3265 55425 3280
rect 55465 3265 55480 3280
rect 56315 3255 56330 3270
rect 56370 3255 56385 3270
rect 56425 3255 56440 3270
rect 56480 3255 56495 3270
rect 56535 3255 56550 3270
rect 56590 3255 56605 3270
rect 56645 3255 56660 3270
rect 56700 3255 56715 3270
rect 56755 3255 56770 3270
rect 56810 3255 56825 3270
rect 56865 3255 56880 3270
rect 56920 3255 56935 3270
rect 56975 3255 56990 3270
rect 57030 3255 57045 3270
rect 57085 3255 57100 3270
rect 57140 3255 57155 3270
rect 57195 3255 57210 3270
rect 57250 3255 57265 3270
rect 57305 3255 57320 3270
rect 57360 3255 57375 3270
rect 57415 3255 57430 3270
rect 57470 3255 57485 3270
rect 58320 3265 58335 3280
rect 58375 3265 58390 3280
rect 58430 3265 58445 3280
rect 58485 3265 58500 3280
rect 58540 3265 58555 3280
rect 58595 3265 58610 3280
rect 58650 3265 58665 3280
rect 58705 3265 58720 3280
rect 58760 3265 58775 3280
rect 58815 3265 58830 3280
rect 58870 3265 58885 3280
rect 58925 3265 58940 3280
rect 56315 3190 56330 3205
rect 56280 3180 56330 3190
rect 56370 3195 56385 3205
rect 56425 3195 56440 3205
rect 56480 3195 56495 3205
rect 56535 3195 56550 3205
rect 56590 3195 56605 3205
rect 56645 3195 56660 3205
rect 56700 3195 56715 3205
rect 56755 3195 56770 3205
rect 56810 3195 56825 3205
rect 56865 3195 56880 3205
rect 56920 3195 56935 3205
rect 56975 3195 56990 3205
rect 57030 3195 57045 3205
rect 57085 3195 57100 3205
rect 57140 3195 57155 3205
rect 57195 3195 57210 3205
rect 57250 3195 57265 3205
rect 57305 3195 57320 3205
rect 57360 3195 57375 3205
rect 57415 3195 57430 3205
rect 56370 3180 57430 3195
rect 57470 3190 57485 3205
rect 57470 3180 57520 3190
rect 56280 3160 56285 3180
rect 56305 3175 56330 3180
rect 56305 3160 56310 3175
rect 56280 3150 56310 3160
rect 56390 3160 56395 3180
rect 56415 3160 56420 3180
rect 56390 3150 56420 3160
rect 56830 3160 56835 3180
rect 56855 3160 56860 3180
rect 57470 3175 57495 3180
rect 56830 3150 56860 3160
rect 57490 3160 57495 3175
rect 57515 3160 57520 3180
rect 57490 3150 57520 3160
rect 56040 3015 56070 3025
rect 56040 2995 56045 3015
rect 56065 3000 56070 3015
rect 56690 3015 56720 3025
rect 56690 3000 56695 3015
rect 56065 2995 56695 3000
rect 56715 2995 56720 3015
rect 56040 2985 56720 2995
rect 57080 3015 57110 3025
rect 57080 2995 57085 3015
rect 57105 3000 57110 3015
rect 57730 3015 57760 3025
rect 57730 3000 57735 3015
rect 57105 2995 57735 3000
rect 57755 2995 57760 3015
rect 57080 2985 57760 2995
rect 56070 2945 56085 2960
rect 56125 2945 56140 2960
rect 56180 2945 56195 2985
rect 56235 2945 56250 2985
rect 56290 2945 56305 2960
rect 56345 2945 56360 2960
rect 56400 2945 56415 2985
rect 56455 2945 56470 2985
rect 56510 2945 56525 2960
rect 56565 2945 56580 2960
rect 56620 2945 56635 2985
rect 56675 2945 56690 2960
rect 57110 2945 57125 2960
rect 57165 2945 57180 2985
rect 57220 2945 57235 2960
rect 57275 2945 57290 2960
rect 57330 2945 57345 2985
rect 57385 2945 57400 2985
rect 57440 2945 57455 2960
rect 57495 2945 57510 2960
rect 57550 2945 57565 2985
rect 57605 2945 57620 2985
rect 57660 2945 57675 2960
rect 57715 2945 57730 2960
rect 56070 2880 56085 2895
rect 56035 2870 56085 2880
rect 56035 2850 56040 2870
rect 56060 2865 56085 2870
rect 56060 2850 56065 2865
rect 56035 2840 56065 2850
rect 56125 2855 56140 2895
rect 56180 2880 56195 2895
rect 56235 2880 56250 2895
rect 56290 2855 56305 2895
rect 56345 2855 56360 2895
rect 56400 2880 56415 2895
rect 56455 2880 56470 2895
rect 56510 2855 56525 2895
rect 56565 2855 56580 2895
rect 56620 2880 56635 2895
rect 56675 2880 56690 2895
rect 57110 2880 57125 2895
rect 57165 2880 57180 2895
rect 56675 2870 56725 2880
rect 56675 2865 56700 2870
rect 56125 2840 56580 2855
rect 56695 2850 56700 2865
rect 56720 2850 56725 2870
rect 56695 2840 56725 2850
rect 57075 2870 57125 2880
rect 57075 2850 57080 2870
rect 57100 2865 57125 2870
rect 57100 2850 57105 2865
rect 57075 2840 57105 2850
rect 57220 2855 57235 2895
rect 57275 2855 57290 2895
rect 57330 2880 57345 2895
rect 57385 2880 57400 2895
rect 57440 2855 57455 2895
rect 57495 2855 57510 2895
rect 57550 2880 57565 2895
rect 57605 2880 57620 2895
rect 57660 2855 57675 2895
rect 57715 2880 57730 2895
rect 57715 2870 57765 2880
rect 57715 2865 57740 2870
rect 57220 2840 57675 2855
rect 57735 2850 57740 2865
rect 57760 2850 57765 2870
rect 57735 2840 57765 2850
rect 56125 2795 56140 2840
rect 56095 2785 56140 2795
rect 56565 2805 56580 2840
rect 57220 2805 57235 2840
rect 56565 2795 56610 2805
rect 56565 2785 56585 2795
rect 56095 2765 56100 2785
rect 56120 2775 56140 2785
rect 56580 2775 56585 2785
rect 56605 2775 56610 2795
rect 56120 2765 56125 2775
rect 56580 2765 56610 2775
rect 57190 2795 57235 2805
rect 57190 2775 57195 2795
rect 57215 2785 57235 2795
rect 57215 2775 57220 2785
rect 57190 2765 57220 2775
rect 56095 2755 56125 2765
rect 54860 2650 54875 2665
rect 54915 2655 54930 2665
rect 54970 2655 54985 2665
rect 55025 2655 55040 2665
rect 55080 2655 55095 2665
rect 55135 2655 55150 2665
rect 55190 2655 55205 2665
rect 55245 2655 55260 2665
rect 55300 2655 55315 2665
rect 55355 2655 55370 2665
rect 55410 2655 55425 2665
rect 54915 2640 55425 2655
rect 55465 2650 55480 2665
rect 58320 2650 58335 2665
rect 58375 2655 58390 2665
rect 58430 2655 58445 2665
rect 58485 2655 58500 2665
rect 58540 2655 58555 2665
rect 58595 2655 58610 2665
rect 58650 2655 58665 2665
rect 58705 2655 58720 2665
rect 58760 2655 58775 2665
rect 58815 2655 58830 2665
rect 58870 2655 58885 2665
rect 58375 2640 58885 2655
rect 58925 2650 58940 2665
rect 55155 2620 55160 2640
rect 55180 2620 55185 2640
rect 55155 2585 55185 2620
rect 56850 2630 56890 2640
rect 56850 2610 56860 2630
rect 56880 2610 56890 2630
rect 58615 2620 58620 2640
rect 58640 2620 58645 2640
rect 56850 2600 56935 2610
rect 56810 2585 56825 2600
rect 56865 2595 56935 2600
rect 56865 2585 56880 2595
rect 56920 2585 56935 2595
rect 56975 2585 56990 2600
rect 58615 2585 58645 2620
rect 55150 2575 55190 2585
rect 55150 2555 55160 2575
rect 55180 2555 55190 2575
rect 55150 2535 55190 2555
rect 55150 2515 55160 2535
rect 55180 2515 55190 2535
rect 55150 2495 55190 2515
rect 55150 2475 55160 2495
rect 55180 2475 55190 2495
rect 55150 2465 55190 2475
rect 58610 2575 58650 2585
rect 58610 2555 58620 2575
rect 58640 2555 58650 2575
rect 58610 2535 58650 2555
rect 58610 2515 58620 2535
rect 58640 2515 58650 2535
rect 58610 2495 58650 2515
rect 58610 2475 58620 2495
rect 58640 2475 58650 2495
rect 58610 2465 58650 2475
rect 56810 2320 56825 2335
rect 56865 2320 56880 2335
rect 56920 2320 56935 2335
rect 56975 2320 56990 2335
rect 56770 2310 56825 2320
rect 56770 2290 56780 2310
rect 56800 2305 56825 2310
rect 56975 2310 57030 2320
rect 56975 2305 57000 2310
rect 56800 2290 56810 2305
rect 56770 2280 56810 2290
rect 56990 2290 57000 2305
rect 57020 2290 57030 2310
rect 56990 2280 57030 2290
rect 55995 2265 56025 2275
rect 55995 2245 56000 2265
rect 56020 2250 56025 2265
rect 56690 2265 56720 2275
rect 56690 2250 56695 2265
rect 56020 2245 56140 2250
rect 55995 2235 56140 2245
rect 54825 2210 54855 2220
rect 54825 2190 54830 2210
rect 54850 2195 54855 2210
rect 55485 2210 55515 2220
rect 55485 2195 55490 2210
rect 54850 2190 54875 2195
rect 54825 2180 54875 2190
rect 55465 2190 55490 2195
rect 55510 2190 55515 2210
rect 56125 2205 56140 2235
rect 56620 2245 56695 2250
rect 56715 2245 56720 2265
rect 56620 2235 56720 2245
rect 57080 2265 57110 2275
rect 57080 2245 57085 2265
rect 57105 2250 57110 2265
rect 57105 2245 57180 2250
rect 57080 2235 57180 2245
rect 56620 2205 56635 2235
rect 55465 2180 55515 2190
rect 56070 2180 56085 2195
rect 56125 2190 56635 2205
rect 57165 2205 57180 2235
rect 58285 2210 58315 2220
rect 56125 2180 56140 2190
rect 56180 2180 56195 2190
rect 56235 2180 56250 2190
rect 56290 2180 56305 2190
rect 56345 2180 56360 2190
rect 56400 2180 56415 2190
rect 56455 2180 56470 2190
rect 56510 2180 56525 2190
rect 56565 2180 56580 2190
rect 56620 2180 56635 2190
rect 56675 2180 56690 2195
rect 57110 2180 57125 2195
rect 57165 2190 57675 2205
rect 57165 2180 57180 2190
rect 57220 2180 57235 2190
rect 57275 2180 57290 2190
rect 57330 2180 57345 2190
rect 57385 2180 57400 2190
rect 57440 2180 57455 2190
rect 57495 2180 57510 2190
rect 57550 2180 57565 2190
rect 57605 2180 57620 2190
rect 57660 2180 57675 2190
rect 57715 2180 57730 2195
rect 58285 2190 58290 2210
rect 58310 2195 58315 2210
rect 58945 2210 58975 2220
rect 58945 2195 58950 2210
rect 58310 2190 58335 2195
rect 58285 2180 58335 2190
rect 58925 2190 58950 2195
rect 58970 2190 58975 2210
rect 58925 2180 58975 2190
rect 54860 2165 54875 2180
rect 54915 2165 54930 2180
rect 54970 2165 54985 2180
rect 55025 2165 55040 2180
rect 55080 2165 55095 2180
rect 55135 2165 55150 2180
rect 55190 2165 55205 2180
rect 55245 2165 55260 2180
rect 55300 2165 55315 2180
rect 55355 2165 55370 2180
rect 55410 2165 55425 2180
rect 55465 2165 55480 2180
rect 58320 2165 58335 2180
rect 58375 2165 58390 2180
rect 58430 2165 58445 2180
rect 58485 2165 58500 2180
rect 58540 2165 58555 2180
rect 58595 2165 58610 2180
rect 58650 2165 58665 2180
rect 58705 2165 58720 2180
rect 58760 2165 58775 2180
rect 58815 2165 58830 2180
rect 58870 2165 58885 2180
rect 58925 2165 58940 2180
rect 56070 2015 56085 2030
rect 56125 2015 56140 2030
rect 56180 2015 56195 2030
rect 56235 2015 56250 2030
rect 56290 2015 56305 2030
rect 56345 2015 56360 2030
rect 56400 2015 56415 2030
rect 56455 2015 56470 2030
rect 56510 2015 56525 2030
rect 56565 2015 56580 2030
rect 56620 2015 56635 2030
rect 56675 2015 56690 2030
rect 57110 2015 57125 2030
rect 57165 2015 57180 2030
rect 57220 2015 57235 2030
rect 57275 2015 57290 2030
rect 57330 2015 57345 2030
rect 57385 2015 57400 2030
rect 57440 2015 57455 2030
rect 57495 2015 57510 2030
rect 57550 2015 57565 2030
rect 57605 2015 57620 2030
rect 57660 2015 57675 2030
rect 57715 2015 57730 2030
rect 56035 2005 56085 2015
rect 56035 1985 56040 2005
rect 56060 2000 56085 2005
rect 56675 2005 56725 2015
rect 56675 2000 56700 2005
rect 56060 1985 56065 2000
rect 56035 1975 56065 1985
rect 56695 1985 56700 2000
rect 56720 1985 56725 2005
rect 56695 1975 56725 1985
rect 57075 2005 57125 2015
rect 57075 1985 57080 2005
rect 57100 2000 57125 2005
rect 57715 2005 57765 2015
rect 57715 2000 57740 2005
rect 57100 1985 57105 2000
rect 57075 1975 57105 1985
rect 57735 1985 57740 2000
rect 57760 1985 57765 2005
rect 57735 1975 57765 1985
rect 54860 1950 54875 1965
rect 54915 1955 54930 1965
rect 54970 1955 54985 1965
rect 55025 1955 55040 1965
rect 55080 1955 55095 1965
rect 55135 1955 55150 1965
rect 55190 1955 55205 1965
rect 55245 1955 55260 1965
rect 55300 1955 55315 1965
rect 55355 1955 55370 1965
rect 55410 1955 55425 1965
rect 54915 1940 55425 1955
rect 55465 1950 55480 1965
rect 58320 1950 58335 1965
rect 58375 1955 58390 1965
rect 58430 1955 58445 1965
rect 58485 1955 58500 1965
rect 58540 1955 58555 1965
rect 58595 1955 58610 1965
rect 58650 1955 58665 1965
rect 58705 1955 58720 1965
rect 58760 1955 58775 1965
rect 58815 1955 58830 1965
rect 58870 1955 58885 1965
rect 58375 1940 58885 1955
rect 58925 1950 58940 1965
rect 55320 1920 55325 1940
rect 55345 1920 55350 1940
rect 55320 1910 55350 1920
rect 58450 1920 58455 1940
rect 58475 1920 58480 1940
rect 58450 1910 58480 1920
rect 55325 1885 55345 1910
rect 58455 1885 58475 1910
rect 55315 1875 55355 1885
rect 55315 1855 55325 1875
rect 55345 1855 55355 1875
rect 55315 1835 55355 1855
rect 55315 1815 55325 1835
rect 55345 1815 55355 1835
rect 55315 1805 55355 1815
rect 58445 1875 58485 1885
rect 58445 1855 58455 1875
rect 58475 1855 58485 1875
rect 58445 1835 58485 1855
rect 58445 1815 58455 1835
rect 58475 1815 58485 1835
rect 58445 1805 58485 1815
rect 55325 1780 55345 1805
rect 56040 1780 56070 1790
rect 55320 1770 55350 1780
rect 55320 1750 55325 1770
rect 55345 1750 55350 1770
rect 56040 1760 56045 1780
rect 56065 1765 56070 1780
rect 56690 1780 56720 1790
rect 56690 1765 56695 1780
rect 56065 1760 56140 1765
rect 56040 1750 56140 1760
rect 54860 1725 54875 1740
rect 54915 1735 55425 1750
rect 54915 1725 54930 1735
rect 54970 1725 54985 1735
rect 55025 1725 55040 1735
rect 55080 1725 55095 1735
rect 55135 1725 55150 1735
rect 55190 1725 55205 1735
rect 55245 1725 55260 1735
rect 55300 1725 55315 1735
rect 55355 1725 55370 1735
rect 55410 1725 55425 1735
rect 55465 1725 55480 1740
rect 56125 1735 56140 1750
rect 56620 1760 56695 1765
rect 56715 1760 56720 1780
rect 56620 1750 56720 1760
rect 56850 1780 56880 1790
rect 56850 1760 56855 1780
rect 56875 1760 56880 1780
rect 56850 1750 56880 1760
rect 56903 1780 56933 1790
rect 56903 1760 56908 1780
rect 56928 1760 56933 1780
rect 57080 1780 57110 1790
rect 57080 1760 57085 1780
rect 57105 1765 57110 1780
rect 57730 1780 57760 1790
rect 58455 1780 58475 1805
rect 57730 1765 57735 1780
rect 57105 1760 57180 1765
rect 56903 1750 56935 1760
rect 57080 1750 57180 1760
rect 56620 1735 56635 1750
rect 56070 1710 56085 1725
rect 56125 1720 56635 1735
rect 56125 1710 56140 1720
rect 56180 1710 56195 1720
rect 56235 1710 56250 1720
rect 56290 1710 56305 1720
rect 56345 1710 56360 1720
rect 56400 1710 56415 1720
rect 56455 1710 56470 1720
rect 56510 1710 56525 1720
rect 56565 1710 56580 1720
rect 56620 1710 56635 1720
rect 56675 1710 56690 1725
rect 56810 1710 56825 1725
rect 56865 1710 56880 1750
rect 56920 1710 56935 1750
rect 57165 1735 57180 1750
rect 57660 1760 57735 1765
rect 57755 1760 57760 1780
rect 57660 1750 57760 1760
rect 58450 1770 58480 1780
rect 58450 1750 58455 1770
rect 58475 1750 58480 1770
rect 57660 1735 57675 1750
rect 56975 1710 56990 1725
rect 57110 1710 57125 1725
rect 57165 1720 57675 1735
rect 58320 1725 58335 1740
rect 58375 1735 58885 1750
rect 58375 1725 58390 1735
rect 58430 1725 58445 1735
rect 58485 1725 58500 1735
rect 58540 1725 58555 1735
rect 58595 1725 58610 1735
rect 58650 1725 58665 1735
rect 58705 1725 58720 1735
rect 58760 1725 58775 1735
rect 58815 1725 58830 1735
rect 58870 1725 58885 1735
rect 58925 1725 58940 1740
rect 57165 1710 57180 1720
rect 57220 1710 57235 1720
rect 57275 1710 57290 1720
rect 57330 1710 57345 1720
rect 57385 1710 57400 1720
rect 57440 1710 57455 1720
rect 57495 1710 57510 1720
rect 57550 1710 57565 1720
rect 57605 1710 57620 1720
rect 57660 1710 57675 1720
rect 57715 1710 57730 1725
rect 56070 1545 56085 1560
rect 56125 1545 56140 1560
rect 56180 1545 56195 1560
rect 56235 1545 56250 1560
rect 56290 1545 56305 1560
rect 56345 1545 56360 1560
rect 56400 1545 56415 1560
rect 56455 1545 56470 1560
rect 56510 1545 56525 1560
rect 56565 1545 56580 1560
rect 56620 1545 56635 1560
rect 56675 1545 56690 1560
rect 56810 1545 56825 1560
rect 56865 1545 56880 1560
rect 56920 1545 56935 1560
rect 56975 1545 56990 1560
rect 57110 1545 57125 1560
rect 57165 1545 57180 1560
rect 57220 1545 57235 1560
rect 57275 1545 57290 1560
rect 57330 1545 57345 1560
rect 57385 1545 57400 1560
rect 57440 1545 57455 1560
rect 57495 1545 57510 1560
rect 57550 1545 57565 1560
rect 57605 1545 57620 1560
rect 57660 1545 57675 1560
rect 57715 1545 57730 1560
rect 56035 1535 56085 1545
rect 56035 1515 56040 1535
rect 56060 1530 56085 1535
rect 56675 1535 56825 1545
rect 56675 1530 56740 1535
rect 56060 1515 56065 1530
rect 56035 1505 56065 1515
rect 56735 1515 56740 1530
rect 56760 1530 56825 1535
rect 56975 1535 57125 1545
rect 56975 1530 57040 1535
rect 56760 1515 56765 1530
rect 56735 1505 56765 1515
rect 57035 1515 57040 1530
rect 57060 1530 57125 1535
rect 57715 1535 57765 1545
rect 57715 1530 57740 1535
rect 57060 1515 57065 1530
rect 57035 1505 57065 1515
rect 57735 1515 57740 1530
rect 57760 1515 57765 1535
rect 57735 1505 57765 1515
rect 54860 1410 54875 1425
rect 54915 1410 54930 1425
rect 54970 1410 54985 1425
rect 55025 1410 55040 1425
rect 55080 1410 55095 1425
rect 55135 1410 55150 1425
rect 55190 1410 55205 1425
rect 55245 1410 55260 1425
rect 55300 1410 55315 1425
rect 55355 1410 55370 1425
rect 55410 1410 55425 1425
rect 55465 1410 55480 1425
rect 58320 1410 58335 1425
rect 58375 1410 58390 1425
rect 58430 1410 58445 1425
rect 58485 1410 58500 1425
rect 58540 1410 58555 1425
rect 58595 1410 58610 1425
rect 58650 1410 58665 1425
rect 58705 1410 58720 1425
rect 58760 1410 58775 1425
rect 58815 1410 58830 1425
rect 58870 1410 58885 1425
rect 58925 1410 58940 1425
rect 54825 1400 54875 1410
rect 54825 1380 54830 1400
rect 54850 1395 54875 1400
rect 55465 1400 55515 1410
rect 55465 1395 55490 1400
rect 54850 1380 54855 1395
rect 54825 1370 54855 1380
rect 55485 1380 55490 1395
rect 55510 1380 55515 1400
rect 55485 1370 55515 1380
rect 58285 1400 58335 1410
rect 58285 1380 58290 1400
rect 58310 1395 58335 1400
rect 58925 1400 58975 1410
rect 58925 1395 58950 1400
rect 58310 1380 58315 1395
rect 58285 1370 58315 1380
rect 58945 1380 58950 1395
rect 58970 1380 58975 1400
rect 58945 1370 58975 1380
rect 55180 1235 55220 1245
rect 55180 1215 55190 1235
rect 55210 1215 55220 1235
rect 55180 1205 55220 1215
rect 58580 1235 58620 1245
rect 58580 1215 58590 1235
rect 58610 1215 58620 1235
rect 58580 1205 58620 1215
rect 55190 1080 55210 1205
rect 57390 1110 57430 1120
rect 57390 1090 57400 1110
rect 57420 1090 57430 1110
rect 57390 1080 57430 1090
rect 58590 1080 58610 1205
rect 54870 1055 54930 1070
rect 54970 1065 55330 1080
rect 54970 1055 55030 1065
rect 55070 1055 55130 1065
rect 55170 1055 55230 1065
rect 55270 1055 55330 1065
rect 55370 1055 55430 1070
rect 56830 1055 56860 1065
rect 56830 1035 56835 1055
rect 56855 1035 56860 1055
rect 56260 1010 56275 1025
rect 56315 1020 57375 1035
rect 56315 1010 56330 1020
rect 56370 1010 56385 1020
rect 56425 1010 56440 1020
rect 56480 1010 56495 1020
rect 56535 1010 56550 1020
rect 56590 1010 56605 1020
rect 56645 1010 56660 1020
rect 56700 1010 56715 1020
rect 56755 1010 56770 1020
rect 56810 1010 56825 1020
rect 56865 1010 56880 1020
rect 56920 1010 56935 1020
rect 56975 1010 56990 1020
rect 57030 1010 57045 1020
rect 57085 1010 57100 1020
rect 57140 1010 57155 1020
rect 57195 1010 57210 1020
rect 57250 1010 57265 1020
rect 57305 1010 57320 1020
rect 57360 1010 57375 1020
rect 57415 1010 57430 1080
rect 58370 1055 58430 1070
rect 58470 1065 58830 1080
rect 58470 1055 58530 1065
rect 58570 1055 58630 1065
rect 58670 1055 58730 1065
rect 58770 1055 58830 1065
rect 58870 1055 58930 1070
rect 57470 1010 57485 1025
rect 56260 745 56275 760
rect 56315 745 56330 760
rect 56370 745 56385 760
rect 56425 745 56440 760
rect 56480 745 56495 760
rect 56535 745 56550 760
rect 56590 745 56605 760
rect 56645 745 56660 760
rect 56700 745 56715 760
rect 56755 745 56770 760
rect 56810 745 56825 760
rect 56865 745 56880 760
rect 56920 745 56935 760
rect 56975 745 56990 760
rect 57030 745 57045 760
rect 57085 745 57100 760
rect 57140 745 57155 760
rect 57195 745 57210 760
rect 57250 745 57265 760
rect 57305 745 57320 760
rect 57360 745 57375 760
rect 57415 745 57430 760
rect 57470 745 57485 760
rect 56220 735 56275 745
rect 56220 715 56230 735
rect 56250 730 56275 735
rect 57470 735 57525 745
rect 57470 730 57495 735
rect 56250 715 56260 730
rect 56220 705 56260 715
rect 57485 715 57495 730
rect 57515 715 57525 735
rect 57485 705 57525 715
rect 56595 590 56635 600
rect 56595 570 56605 590
rect 56625 570 56635 590
rect 57040 590 57080 600
rect 57040 570 57050 590
rect 57070 570 57080 590
rect 56470 545 56485 560
rect 56525 555 56705 570
rect 57040 560 57080 570
rect 56525 545 56540 555
rect 56580 545 56595 555
rect 56635 545 56650 555
rect 56690 545 56705 555
rect 56745 545 56760 560
rect 56910 545 57210 560
rect 56470 380 56485 395
rect 56525 380 56540 395
rect 56580 380 56595 395
rect 56635 380 56650 395
rect 56690 380 56705 395
rect 56745 380 56760 395
rect 56910 380 57210 395
rect 56435 370 56485 380
rect 54870 340 54930 355
rect 54970 340 55030 355
rect 55070 340 55130 355
rect 55170 340 55230 355
rect 55270 340 55330 355
rect 55370 340 55430 355
rect 56435 350 56440 370
rect 56460 365 56485 370
rect 56745 370 56795 380
rect 56745 365 56770 370
rect 56460 350 56465 365
rect 56435 340 56465 350
rect 56765 350 56770 365
rect 56790 350 56795 370
rect 56765 340 56795 350
rect 58370 340 58430 355
rect 58470 340 58530 355
rect 58570 340 58630 355
rect 58670 340 58730 355
rect 58770 340 58830 355
rect 58870 340 58930 355
rect 54835 330 54930 340
rect 54835 310 54840 330
rect 54860 325 54930 330
rect 55370 330 55465 340
rect 55370 325 55440 330
rect 54860 310 54865 325
rect 54835 300 54865 310
rect 55435 310 55440 325
rect 55460 310 55465 330
rect 55435 300 55465 310
rect 58335 330 58430 340
rect 58335 310 58340 330
rect 58360 325 58430 330
rect 58870 330 58965 340
rect 58870 325 58940 330
rect 58360 310 58365 325
rect 58335 300 58365 310
rect 58935 310 58940 325
rect 58960 310 58965 330
rect 58935 300 58965 310
<< polycont >>
rect 56095 4940 56115 4960
rect 56275 4940 56295 4960
rect 57035 4940 57055 4960
rect 57215 4940 57235 4960
rect 57505 4940 57525 4960
rect 57685 4940 57705 4960
rect 56565 4770 56585 4790
rect 56745 4770 56765 4790
rect 56160 4490 56180 4510
rect 56635 4490 56655 4510
rect 57145 4490 57165 4510
rect 57581 4480 57601 4500
rect 54930 3645 54950 3665
rect 55290 3645 55310 3665
rect 55650 3645 55670 3665
rect 56015 3645 56035 3665
rect 56375 3645 56395 3665
rect 56735 3645 56755 3665
rect 57045 3645 57065 3665
rect 57405 3645 57425 3665
rect 57765 3645 57785 3665
rect 58130 3645 58150 3665
rect 58490 3645 58510 3665
rect 58850 3645 58870 3665
rect 56375 3580 56395 3600
rect 57405 3580 57425 3600
rect 55290 3535 55310 3555
rect 58490 3535 58510 3555
rect 54830 3290 54850 3310
rect 55490 3290 55510 3310
rect 58290 3290 58310 3310
rect 58950 3290 58970 3310
rect 56285 3160 56305 3180
rect 56395 3160 56415 3180
rect 56835 3160 56855 3180
rect 57495 3160 57515 3180
rect 56045 2995 56065 3015
rect 56695 2995 56715 3015
rect 57085 2995 57105 3015
rect 57735 2995 57755 3015
rect 56040 2850 56060 2870
rect 56700 2850 56720 2870
rect 57080 2850 57100 2870
rect 57740 2850 57760 2870
rect 56100 2765 56120 2785
rect 56585 2775 56605 2795
rect 57195 2775 57215 2795
rect 55160 2620 55180 2640
rect 56860 2610 56880 2630
rect 58620 2620 58640 2640
rect 55160 2555 55180 2575
rect 55160 2515 55180 2535
rect 55160 2475 55180 2495
rect 58620 2555 58640 2575
rect 58620 2515 58640 2535
rect 58620 2475 58640 2495
rect 56780 2290 56800 2310
rect 57000 2290 57020 2310
rect 56000 2245 56020 2265
rect 54830 2190 54850 2210
rect 55490 2190 55510 2210
rect 56695 2245 56715 2265
rect 57085 2245 57105 2265
rect 58290 2190 58310 2210
rect 58950 2190 58970 2210
rect 56040 1985 56060 2005
rect 56700 1985 56720 2005
rect 57080 1985 57100 2005
rect 57740 1985 57760 2005
rect 55325 1920 55345 1940
rect 58455 1920 58475 1940
rect 55325 1855 55345 1875
rect 55325 1815 55345 1835
rect 58455 1855 58475 1875
rect 58455 1815 58475 1835
rect 55325 1750 55345 1770
rect 56045 1760 56065 1780
rect 56695 1760 56715 1780
rect 56855 1760 56875 1780
rect 56908 1760 56928 1780
rect 57085 1760 57105 1780
rect 57735 1760 57755 1780
rect 58455 1750 58475 1770
rect 56040 1515 56060 1535
rect 56740 1515 56760 1535
rect 57040 1515 57060 1535
rect 57740 1515 57760 1535
rect 54830 1380 54850 1400
rect 55490 1380 55510 1400
rect 58290 1380 58310 1400
rect 58950 1380 58970 1400
rect 55190 1215 55210 1235
rect 58590 1215 58610 1235
rect 57400 1090 57420 1110
rect 56835 1035 56855 1055
rect 56230 715 56250 735
rect 57495 715 57515 735
rect 56605 570 56625 590
rect 57050 570 57070 590
rect 56440 350 56460 370
rect 56770 350 56790 370
rect 54840 310 54860 330
rect 55440 310 55460 330
rect 58340 310 58360 330
rect 58940 310 58960 330
<< xpolycontact >>
rect 54554 3065 54695 3285
rect 54554 2720 54695 2940
rect 59105 3065 59246 3285
rect 59105 2720 59246 2940
rect 54460 1779 54495 1999
rect 54460 1400 54495 1620
rect 54520 1779 54555 1999
rect 54520 1400 54555 1620
rect 54580 1779 54615 1999
rect 54580 1400 54615 1620
rect 54640 1779 54675 1999
rect 54640 1400 54675 1620
rect 59125 1779 59160 1999
rect 59125 1400 59160 1620
rect 59185 1779 59220 1999
rect 59185 1400 59220 1620
rect 59245 1779 59280 1999
rect 59245 1400 59280 1620
rect 59305 1779 59340 1999
rect 59305 1400 59340 1620
rect 54600 790 54635 1010
rect 54600 323 54635 543
rect 54660 790 54695 1010
rect 54660 323 54695 543
rect 59105 790 59140 1010
rect 59105 323 59140 543
rect 59165 790 59200 1010
rect 59165 323 59200 543
<< ppolyres >>
rect 54554 2940 54695 3065
rect 59105 2940 59246 3065
<< xpolyres >>
rect 54460 1620 54495 1779
rect 54520 1620 54555 1779
rect 54580 1620 54615 1779
rect 54640 1620 54675 1779
rect 59125 1620 59160 1779
rect 59185 1620 59220 1779
rect 59245 1620 59280 1779
rect 59305 1620 59340 1779
rect 54600 543 54635 790
rect 54660 543 54695 790
rect 59105 543 59140 790
rect 59165 543 59200 790
<< locali >>
rect 56085 4960 56125 4970
rect 56085 4940 56095 4960
rect 56115 4940 56125 4960
rect 56085 4930 56125 4940
rect 56265 4960 56305 4970
rect 56265 4940 56275 4960
rect 56295 4940 56305 4960
rect 56265 4930 56305 4940
rect 57025 4960 57065 4970
rect 57025 4940 57035 4960
rect 57055 4940 57065 4960
rect 57025 4930 57065 4940
rect 57205 4960 57245 4970
rect 57205 4940 57215 4960
rect 57235 4940 57245 4960
rect 57205 4930 57245 4940
rect 57495 4960 57535 4970
rect 57495 4940 57505 4960
rect 57525 4940 57535 4960
rect 57495 4930 57535 4940
rect 57675 4960 57715 4970
rect 57675 4940 57685 4960
rect 57705 4940 57715 4960
rect 57675 4930 57715 4940
rect 56050 4900 56120 4910
rect 56050 4580 56055 4900
rect 56075 4580 56095 4900
rect 56115 4580 56120 4900
rect 56050 4570 56120 4580
rect 56150 4900 56180 4910
rect 56150 4580 56155 4900
rect 56175 4580 56180 4900
rect 56150 4570 56180 4580
rect 56210 4900 56240 4910
rect 56210 4580 56215 4900
rect 56235 4580 56240 4900
rect 56210 4570 56240 4580
rect 56270 4900 56340 4910
rect 56270 4580 56275 4900
rect 56295 4580 56315 4900
rect 56335 4580 56340 4900
rect 56990 4900 57060 4910
rect 56555 4790 56595 4800
rect 56555 4770 56565 4790
rect 56585 4770 56595 4790
rect 56555 4760 56595 4770
rect 56735 4790 56775 4800
rect 56735 4770 56745 4790
rect 56765 4770 56775 4790
rect 56735 4760 56775 4770
rect 56270 4570 56340 4580
rect 56520 4730 56590 4740
rect 56520 4580 56525 4730
rect 56545 4580 56565 4730
rect 56585 4580 56590 4730
rect 56520 4570 56590 4580
rect 56620 4730 56650 4740
rect 56620 4580 56625 4730
rect 56645 4580 56650 4730
rect 56620 4570 56650 4580
rect 56680 4730 56710 4740
rect 56680 4580 56685 4730
rect 56705 4580 56710 4730
rect 56680 4570 56710 4580
rect 56740 4730 56810 4740
rect 56740 4580 56745 4730
rect 56765 4580 56785 4730
rect 56805 4580 56810 4730
rect 56740 4570 56810 4580
rect 56990 4580 56995 4900
rect 57015 4580 57035 4900
rect 57055 4580 57060 4900
rect 56990 4570 57060 4580
rect 57090 4900 57120 4910
rect 57090 4580 57095 4900
rect 57115 4580 57120 4900
rect 57090 4570 57120 4580
rect 57150 4900 57180 4910
rect 57150 4580 57155 4900
rect 57175 4580 57180 4900
rect 57150 4570 57180 4580
rect 57210 4900 57280 4910
rect 57210 4580 57215 4900
rect 57235 4580 57255 4900
rect 57275 4580 57280 4900
rect 57210 4570 57280 4580
rect 57460 4900 57530 4910
rect 57460 4580 57465 4900
rect 57485 4580 57505 4900
rect 57525 4580 57530 4900
rect 57460 4570 57530 4580
rect 57560 4900 57590 4910
rect 57560 4580 57565 4900
rect 57585 4580 57590 4900
rect 57560 4570 57590 4580
rect 57620 4900 57650 4910
rect 57620 4580 57625 4900
rect 57645 4580 57650 4900
rect 57620 4570 57650 4580
rect 57680 4900 57750 4910
rect 57680 4580 57685 4900
rect 57705 4580 57725 4900
rect 57745 4580 57750 4900
rect 57680 4570 57750 4580
rect 56150 4510 56190 4520
rect 56150 4490 56160 4510
rect 56180 4490 56190 4510
rect 56150 4480 56190 4490
rect 56630 4510 56660 4520
rect 56630 4490 56635 4510
rect 56655 4490 56660 4510
rect 56630 4480 56660 4490
rect 57140 4510 57170 4520
rect 57140 4490 57145 4510
rect 57165 4490 57170 4510
rect 57140 4480 57170 4490
rect 57576 4500 57606 4510
rect 57576 4480 57581 4500
rect 57601 4480 57606 4500
rect 57576 4470 57606 4480
rect 54885 4025 54955 4035
rect 54885 3705 54890 4025
rect 54910 3705 54930 4025
rect 54950 3705 54955 4025
rect 54885 3695 54955 3705
rect 54985 4025 55015 4035
rect 54985 3705 54990 4025
rect 55010 3705 55015 4025
rect 54985 3695 55015 3705
rect 55045 4025 55075 4035
rect 55045 3705 55050 4025
rect 55070 3705 55075 4025
rect 55045 3695 55075 3705
rect 55105 4025 55135 4035
rect 55105 3705 55110 4025
rect 55130 3705 55135 4025
rect 55105 3695 55135 3705
rect 55165 4025 55195 4035
rect 55165 3705 55170 4025
rect 55190 3705 55195 4025
rect 55165 3695 55195 3705
rect 55225 4025 55255 4035
rect 55225 3705 55230 4025
rect 55250 3705 55255 4025
rect 55225 3695 55255 3705
rect 55285 4025 55315 4035
rect 55285 3705 55290 4025
rect 55310 3705 55315 4025
rect 55285 3695 55315 3705
rect 55345 4025 55375 4035
rect 55345 3705 55350 4025
rect 55370 3705 55375 4025
rect 55345 3695 55375 3705
rect 55405 4025 55435 4035
rect 55405 3705 55410 4025
rect 55430 3705 55435 4025
rect 55405 3695 55435 3705
rect 55465 4025 55495 4035
rect 55465 3705 55470 4025
rect 55490 3705 55495 4025
rect 55465 3695 55495 3705
rect 55525 4025 55555 4035
rect 55525 3705 55530 4025
rect 55550 3705 55555 4025
rect 55525 3695 55555 3705
rect 55585 4025 55615 4035
rect 55585 3705 55590 4025
rect 55610 3705 55615 4025
rect 55585 3695 55615 3705
rect 55645 4025 55715 4035
rect 55645 3705 55650 4025
rect 55670 3705 55690 4025
rect 55710 3705 55715 4025
rect 55645 3695 55715 3705
rect 55970 4025 56040 4035
rect 55970 3705 55975 4025
rect 55995 3705 56015 4025
rect 56035 3705 56040 4025
rect 55970 3695 56040 3705
rect 56070 4025 56100 4035
rect 56070 3705 56075 4025
rect 56095 3705 56100 4025
rect 56070 3695 56100 3705
rect 56130 4025 56160 4035
rect 56130 3705 56135 4025
rect 56155 3705 56160 4025
rect 56130 3695 56160 3705
rect 56190 4025 56220 4035
rect 56190 3705 56195 4025
rect 56215 3705 56220 4025
rect 56190 3695 56220 3705
rect 56250 4025 56280 4035
rect 56250 3705 56255 4025
rect 56275 3705 56280 4025
rect 56250 3695 56280 3705
rect 56310 4025 56340 4035
rect 56310 3705 56315 4025
rect 56335 3705 56340 4025
rect 56310 3695 56340 3705
rect 56370 4025 56400 4035
rect 56370 3705 56375 4025
rect 56395 3705 56400 4025
rect 56370 3695 56400 3705
rect 56430 4025 56460 4035
rect 56430 3705 56435 4025
rect 56455 3705 56460 4025
rect 56430 3695 56460 3705
rect 56490 4025 56520 4035
rect 56490 3705 56495 4025
rect 56515 3705 56520 4025
rect 56490 3695 56520 3705
rect 56550 4025 56580 4035
rect 56550 3705 56555 4025
rect 56575 3705 56580 4025
rect 56550 3695 56580 3705
rect 56610 4025 56640 4035
rect 56610 3705 56615 4025
rect 56635 3705 56640 4025
rect 56610 3695 56640 3705
rect 56670 4025 56700 4035
rect 56670 3705 56675 4025
rect 56695 3705 56700 4025
rect 56670 3695 56700 3705
rect 56730 4025 56800 4035
rect 56730 3705 56735 4025
rect 56755 3705 56775 4025
rect 56795 3705 56800 4025
rect 56730 3695 56800 3705
rect 57000 4025 57070 4035
rect 57000 3705 57005 4025
rect 57025 3705 57045 4025
rect 57065 3705 57070 4025
rect 57000 3695 57070 3705
rect 57100 4025 57130 4035
rect 57100 3705 57105 4025
rect 57125 3705 57130 4025
rect 57100 3695 57130 3705
rect 57160 4025 57190 4035
rect 57160 3705 57165 4025
rect 57185 3705 57190 4025
rect 57160 3695 57190 3705
rect 57220 4025 57250 4035
rect 57220 3705 57225 4025
rect 57245 3705 57250 4025
rect 57220 3695 57250 3705
rect 57280 4025 57310 4035
rect 57280 3705 57285 4025
rect 57305 3705 57310 4025
rect 57280 3695 57310 3705
rect 57340 4025 57370 4035
rect 57340 3705 57345 4025
rect 57365 3705 57370 4025
rect 57340 3695 57370 3705
rect 57400 4025 57430 4035
rect 57400 3705 57405 4025
rect 57425 3705 57430 4025
rect 57400 3695 57430 3705
rect 57460 4025 57490 4035
rect 57460 3705 57465 4025
rect 57485 3705 57490 4025
rect 57460 3695 57490 3705
rect 57520 4025 57550 4035
rect 57520 3705 57525 4025
rect 57545 3705 57550 4025
rect 57520 3695 57550 3705
rect 57580 4025 57610 4035
rect 57580 3705 57585 4025
rect 57605 3705 57610 4025
rect 57580 3695 57610 3705
rect 57640 4025 57670 4035
rect 57640 3705 57645 4025
rect 57665 3705 57670 4025
rect 57640 3695 57670 3705
rect 57700 4025 57730 4035
rect 57700 3705 57705 4025
rect 57725 3705 57730 4025
rect 57700 3695 57730 3705
rect 57760 4025 57830 4035
rect 57760 3705 57765 4025
rect 57785 3705 57805 4025
rect 57825 3705 57830 4025
rect 57760 3695 57830 3705
rect 58085 4025 58155 4035
rect 58085 3705 58090 4025
rect 58110 3705 58130 4025
rect 58150 3705 58155 4025
rect 58085 3695 58155 3705
rect 58185 4025 58215 4035
rect 58185 3705 58190 4025
rect 58210 3705 58215 4025
rect 58185 3695 58215 3705
rect 58245 4025 58275 4035
rect 58245 3705 58250 4025
rect 58270 3705 58275 4025
rect 58245 3695 58275 3705
rect 58305 4025 58335 4035
rect 58305 3705 58310 4025
rect 58330 3705 58335 4025
rect 58305 3695 58335 3705
rect 58365 4025 58395 4035
rect 58365 3705 58370 4025
rect 58390 3705 58395 4025
rect 58365 3695 58395 3705
rect 58425 4025 58455 4035
rect 58425 3705 58430 4025
rect 58450 3705 58455 4025
rect 58425 3695 58455 3705
rect 58485 4025 58515 4035
rect 58485 3705 58490 4025
rect 58510 3705 58515 4025
rect 58485 3695 58515 3705
rect 58545 4025 58575 4035
rect 58545 3705 58550 4025
rect 58570 3705 58575 4025
rect 58545 3695 58575 3705
rect 58605 4025 58635 4035
rect 58605 3705 58610 4025
rect 58630 3705 58635 4025
rect 58605 3695 58635 3705
rect 58665 4025 58695 4035
rect 58665 3705 58670 4025
rect 58690 3705 58695 4025
rect 58665 3695 58695 3705
rect 58725 4025 58755 4035
rect 58725 3705 58730 4025
rect 58750 3705 58755 4025
rect 58725 3695 58755 3705
rect 58785 4025 58815 4035
rect 58785 3705 58790 4025
rect 58810 3705 58815 4025
rect 58785 3695 58815 3705
rect 58845 4025 58915 4035
rect 58845 3705 58850 4025
rect 58870 3705 58890 4025
rect 58910 3705 58915 4025
rect 58845 3695 58915 3705
rect 54925 3665 54955 3675
rect 54925 3645 54930 3665
rect 54950 3645 54955 3665
rect 54925 3635 54955 3645
rect 55285 3665 55315 3675
rect 55285 3645 55290 3665
rect 55310 3645 55315 3665
rect 55285 3635 55315 3645
rect 55645 3665 55675 3675
rect 55645 3645 55650 3665
rect 55670 3645 55675 3665
rect 55645 3635 55675 3645
rect 56010 3665 56040 3675
rect 56010 3645 56015 3665
rect 56035 3645 56040 3665
rect 56010 3635 56040 3645
rect 56370 3665 56400 3675
rect 56370 3645 56375 3665
rect 56395 3645 56400 3665
rect 56370 3635 56400 3645
rect 56730 3665 56760 3675
rect 56730 3645 56735 3665
rect 56755 3645 56760 3665
rect 56730 3635 56760 3645
rect 57040 3665 57070 3675
rect 57040 3645 57045 3665
rect 57065 3645 57070 3665
rect 57040 3635 57070 3645
rect 57400 3665 57430 3675
rect 57400 3645 57405 3665
rect 57425 3645 57430 3665
rect 57400 3635 57430 3645
rect 57760 3665 57790 3675
rect 57760 3645 57765 3665
rect 57785 3645 57790 3665
rect 57760 3635 57790 3645
rect 58125 3665 58155 3675
rect 58125 3645 58130 3665
rect 58150 3645 58155 3665
rect 58125 3635 58155 3645
rect 58485 3665 58515 3675
rect 58485 3645 58490 3665
rect 58510 3645 58515 3665
rect 58485 3635 58515 3645
rect 58845 3665 58875 3675
rect 58845 3645 58850 3665
rect 58870 3645 58875 3665
rect 58845 3635 58875 3645
rect 56365 3600 56405 3610
rect 56365 3580 56375 3600
rect 56395 3580 56405 3600
rect 56365 3570 56405 3580
rect 57395 3600 57435 3610
rect 57395 3580 57405 3600
rect 57425 3580 57435 3600
rect 57395 3570 57435 3580
rect 55280 3555 55320 3565
rect 55280 3535 55290 3555
rect 55310 3535 55320 3555
rect 55280 3525 55320 3535
rect 58480 3555 58520 3565
rect 58480 3535 58490 3555
rect 58510 3535 58520 3555
rect 58480 3525 58520 3535
rect 54554 3315 54695 3325
rect 54554 3295 54560 3315
rect 54580 3295 54615 3315
rect 54635 3295 54670 3315
rect 54690 3295 54695 3315
rect 54554 3285 54695 3295
rect 54825 3310 54855 3320
rect 54825 3290 54830 3310
rect 54850 3290 54855 3310
rect 54825 3280 54855 3290
rect 55485 3310 55515 3320
rect 55485 3290 55490 3310
rect 55510 3290 55515 3310
rect 55485 3280 55515 3290
rect 58285 3310 58315 3320
rect 58285 3290 58290 3310
rect 58310 3290 58315 3310
rect 58285 3280 58315 3290
rect 58945 3310 58975 3320
rect 58945 3290 58950 3310
rect 58970 3290 58975 3310
rect 58945 3280 58975 3290
rect 59105 3315 59246 3325
rect 59105 3295 59110 3315
rect 59130 3295 59165 3315
rect 59185 3295 59220 3315
rect 59240 3295 59246 3315
rect 59105 3285 59246 3295
rect 54785 3250 54855 3260
rect 54554 2710 54695 2720
rect 54554 2690 54560 2710
rect 54580 2690 54615 2710
rect 54635 2690 54670 2710
rect 54690 2690 54695 2710
rect 54554 2680 54695 2690
rect 54785 2680 54790 3250
rect 54810 2680 54830 3250
rect 54850 2680 54855 3250
rect 54785 2670 54855 2680
rect 54880 3250 54910 3260
rect 54880 2680 54885 3250
rect 54905 2680 54910 3250
rect 54880 2670 54910 2680
rect 54935 3250 54965 3260
rect 54935 2680 54940 3250
rect 54960 2680 54965 3250
rect 54935 2670 54965 2680
rect 54990 3250 55020 3260
rect 54990 2680 54995 3250
rect 55015 2680 55020 3250
rect 54990 2670 55020 2680
rect 55045 3250 55075 3260
rect 55045 2680 55050 3250
rect 55070 2680 55075 3250
rect 55045 2670 55075 2680
rect 55100 3250 55130 3260
rect 55100 2680 55105 3250
rect 55125 2680 55130 3250
rect 55100 2670 55130 2680
rect 55155 3250 55185 3260
rect 55155 2680 55160 3250
rect 55180 2680 55185 3250
rect 55155 2670 55185 2680
rect 55210 3250 55240 3260
rect 55210 2680 55215 3250
rect 55235 2680 55240 3250
rect 55210 2670 55240 2680
rect 55265 3250 55295 3260
rect 55265 2680 55270 3250
rect 55290 2680 55295 3250
rect 55265 2670 55295 2680
rect 55320 3250 55350 3260
rect 55320 2680 55325 3250
rect 55345 2680 55350 3250
rect 55320 2670 55350 2680
rect 55375 3250 55405 3260
rect 55375 2680 55380 3250
rect 55400 2680 55405 3250
rect 55375 2670 55405 2680
rect 55430 3250 55460 3260
rect 55430 2680 55435 3250
rect 55455 2680 55460 3250
rect 55430 2670 55460 2680
rect 55485 3250 55555 3260
rect 58245 3250 58315 3260
rect 55485 2680 55490 3250
rect 55510 2680 55530 3250
rect 55550 2680 55555 3250
rect 56240 3240 56310 3250
rect 56240 3220 56245 3240
rect 56265 3220 56285 3240
rect 56305 3220 56310 3240
rect 56240 3210 56310 3220
rect 56335 3240 56365 3250
rect 56335 3220 56340 3240
rect 56360 3220 56365 3240
rect 56335 3210 56365 3220
rect 56390 3240 56420 3250
rect 56390 3220 56395 3240
rect 56415 3220 56420 3240
rect 56390 3210 56420 3220
rect 56445 3240 56475 3250
rect 56445 3220 56450 3240
rect 56470 3220 56475 3240
rect 56445 3210 56475 3220
rect 56500 3240 56530 3250
rect 56500 3220 56505 3240
rect 56525 3220 56530 3240
rect 56500 3210 56530 3220
rect 56555 3240 56585 3250
rect 56555 3220 56560 3240
rect 56580 3220 56585 3240
rect 56555 3210 56585 3220
rect 56610 3240 56640 3250
rect 56610 3220 56615 3240
rect 56635 3220 56640 3240
rect 56610 3210 56640 3220
rect 56665 3240 56695 3250
rect 56665 3220 56670 3240
rect 56690 3220 56695 3240
rect 56665 3210 56695 3220
rect 56720 3240 56750 3250
rect 56720 3220 56725 3240
rect 56745 3220 56750 3240
rect 56720 3210 56750 3220
rect 56775 3240 56805 3250
rect 56775 3220 56780 3240
rect 56800 3220 56805 3240
rect 56775 3210 56805 3220
rect 56830 3240 56860 3250
rect 56830 3220 56835 3240
rect 56855 3220 56860 3240
rect 56830 3210 56860 3220
rect 56885 3240 56915 3250
rect 56885 3220 56890 3240
rect 56910 3220 56915 3240
rect 56885 3210 56915 3220
rect 56940 3240 56970 3250
rect 56940 3220 56945 3240
rect 56965 3220 56970 3240
rect 56940 3210 56970 3220
rect 56995 3240 57025 3250
rect 56995 3220 57000 3240
rect 57020 3220 57025 3240
rect 56995 3210 57025 3220
rect 57050 3240 57080 3250
rect 57050 3220 57055 3240
rect 57075 3220 57080 3240
rect 57050 3210 57080 3220
rect 57105 3240 57135 3250
rect 57105 3220 57110 3240
rect 57130 3220 57135 3240
rect 57105 3210 57135 3220
rect 57160 3240 57190 3250
rect 57160 3220 57165 3240
rect 57185 3220 57190 3240
rect 57160 3210 57190 3220
rect 57215 3240 57245 3250
rect 57215 3220 57220 3240
rect 57240 3220 57245 3240
rect 57215 3210 57245 3220
rect 57270 3240 57300 3250
rect 57270 3220 57275 3240
rect 57295 3220 57300 3240
rect 57270 3210 57300 3220
rect 57325 3240 57355 3250
rect 57325 3220 57330 3240
rect 57350 3220 57355 3240
rect 57325 3210 57355 3220
rect 57380 3240 57410 3250
rect 57380 3220 57385 3240
rect 57405 3220 57410 3240
rect 57380 3210 57410 3220
rect 57435 3240 57465 3250
rect 57435 3220 57440 3240
rect 57460 3220 57465 3240
rect 57435 3210 57465 3220
rect 57490 3240 57560 3250
rect 57490 3220 57495 3240
rect 57515 3220 57535 3240
rect 57555 3220 57560 3240
rect 57490 3210 57560 3220
rect 56280 3180 56310 3190
rect 56280 3160 56285 3180
rect 56305 3160 56310 3180
rect 56280 3150 56310 3160
rect 56390 3180 56420 3190
rect 56390 3160 56395 3180
rect 56415 3160 56420 3180
rect 56390 3150 56420 3160
rect 56830 3180 56860 3190
rect 56830 3160 56835 3180
rect 56855 3160 56860 3180
rect 56830 3150 56860 3160
rect 57490 3180 57520 3190
rect 57490 3160 57495 3180
rect 57515 3160 57520 3180
rect 57490 3150 57520 3160
rect 56040 3015 56070 3025
rect 56040 2995 56045 3015
rect 56065 2995 56070 3015
rect 56040 2985 56070 2995
rect 56690 3015 56720 3025
rect 56690 2995 56695 3015
rect 56715 2995 56720 3015
rect 56690 2985 56720 2995
rect 57080 3015 57110 3025
rect 57080 2995 57085 3015
rect 57105 2995 57110 3015
rect 57080 2985 57110 2995
rect 57730 3015 57760 3025
rect 57730 2995 57735 3015
rect 57755 2995 57760 3015
rect 57730 2985 57760 2995
rect 55995 2930 56065 2940
rect 55995 2910 56000 2930
rect 56020 2910 56040 2930
rect 56060 2910 56065 2930
rect 55995 2900 56065 2910
rect 56090 2930 56120 2940
rect 56090 2910 56095 2930
rect 56115 2910 56120 2930
rect 56090 2900 56120 2910
rect 56145 2930 56175 2940
rect 56145 2910 56150 2930
rect 56170 2910 56175 2930
rect 56145 2900 56175 2910
rect 56200 2930 56230 2940
rect 56200 2910 56205 2930
rect 56225 2910 56230 2930
rect 56200 2900 56230 2910
rect 56255 2930 56285 2940
rect 56255 2910 56260 2930
rect 56280 2910 56285 2930
rect 56255 2900 56285 2910
rect 56310 2930 56340 2940
rect 56310 2910 56315 2930
rect 56335 2910 56340 2930
rect 56310 2900 56340 2910
rect 56365 2930 56395 2940
rect 56365 2910 56370 2930
rect 56390 2910 56395 2930
rect 56365 2900 56395 2910
rect 56420 2930 56450 2940
rect 56420 2910 56425 2930
rect 56445 2910 56450 2930
rect 56420 2900 56450 2910
rect 56475 2930 56505 2940
rect 56475 2910 56480 2930
rect 56500 2910 56505 2930
rect 56475 2900 56505 2910
rect 56530 2930 56560 2940
rect 56530 2910 56535 2930
rect 56555 2910 56560 2930
rect 56530 2900 56560 2910
rect 56585 2930 56615 2940
rect 56585 2910 56590 2930
rect 56610 2910 56615 2930
rect 56585 2900 56615 2910
rect 56640 2930 56670 2940
rect 56640 2910 56645 2930
rect 56665 2910 56670 2930
rect 56640 2900 56670 2910
rect 56695 2930 56765 2940
rect 56695 2910 56700 2930
rect 56720 2910 56740 2930
rect 56760 2910 56765 2930
rect 56695 2900 56765 2910
rect 57035 2930 57105 2940
rect 57035 2910 57040 2930
rect 57060 2910 57080 2930
rect 57100 2910 57105 2930
rect 57035 2900 57105 2910
rect 57130 2930 57160 2940
rect 57130 2910 57135 2930
rect 57155 2910 57160 2930
rect 57130 2900 57160 2910
rect 57185 2930 57215 2940
rect 57185 2910 57190 2930
rect 57210 2910 57215 2930
rect 57185 2900 57215 2910
rect 57240 2930 57270 2940
rect 57240 2910 57245 2930
rect 57265 2910 57270 2930
rect 57240 2900 57270 2910
rect 57295 2930 57325 2940
rect 57295 2910 57300 2930
rect 57320 2910 57325 2930
rect 57295 2900 57325 2910
rect 57350 2930 57380 2940
rect 57350 2910 57355 2930
rect 57375 2910 57380 2930
rect 57350 2900 57380 2910
rect 57405 2930 57435 2940
rect 57405 2910 57410 2930
rect 57430 2910 57435 2930
rect 57405 2900 57435 2910
rect 57460 2930 57490 2940
rect 57460 2910 57465 2930
rect 57485 2910 57490 2930
rect 57460 2900 57490 2910
rect 57515 2930 57545 2940
rect 57515 2910 57520 2930
rect 57540 2910 57545 2930
rect 57515 2900 57545 2910
rect 57570 2930 57600 2940
rect 57570 2910 57575 2930
rect 57595 2910 57600 2930
rect 57570 2900 57600 2910
rect 57625 2930 57655 2940
rect 57625 2910 57630 2930
rect 57650 2910 57655 2930
rect 57625 2900 57655 2910
rect 57680 2930 57710 2940
rect 57680 2910 57685 2930
rect 57705 2910 57710 2930
rect 57680 2900 57710 2910
rect 57735 2930 57805 2940
rect 57735 2910 57740 2930
rect 57760 2910 57780 2930
rect 57800 2910 57805 2930
rect 57735 2900 57805 2910
rect 56035 2870 56065 2880
rect 56035 2850 56040 2870
rect 56060 2850 56065 2870
rect 56035 2840 56065 2850
rect 56695 2870 56725 2880
rect 56695 2850 56700 2870
rect 56720 2850 56725 2870
rect 56695 2840 56725 2850
rect 57075 2870 57105 2880
rect 57075 2850 57080 2870
rect 57100 2850 57105 2870
rect 57075 2840 57105 2850
rect 57735 2870 57765 2880
rect 57735 2850 57740 2870
rect 57760 2850 57765 2870
rect 57735 2840 57765 2850
rect 56580 2795 56610 2805
rect 56095 2785 56125 2795
rect 56095 2765 56100 2785
rect 56120 2765 56125 2785
rect 56580 2775 56585 2795
rect 56605 2775 56610 2795
rect 56580 2765 56610 2775
rect 57190 2795 57220 2805
rect 57190 2775 57195 2795
rect 57215 2775 57220 2795
rect 57190 2765 57220 2775
rect 56095 2755 56125 2765
rect 55485 2670 55555 2680
rect 58245 2680 58250 3250
rect 58270 2680 58290 3250
rect 58310 2680 58315 3250
rect 58245 2670 58315 2680
rect 58340 3250 58370 3260
rect 58340 2680 58345 3250
rect 58365 2680 58370 3250
rect 58340 2670 58370 2680
rect 58395 3250 58425 3260
rect 58395 2680 58400 3250
rect 58420 2680 58425 3250
rect 58395 2670 58425 2680
rect 58450 3250 58480 3260
rect 58450 2680 58455 3250
rect 58475 2680 58480 3250
rect 58450 2670 58480 2680
rect 58505 3250 58535 3260
rect 58505 2680 58510 3250
rect 58530 2680 58535 3250
rect 58505 2670 58535 2680
rect 58560 3250 58590 3260
rect 58560 2680 58565 3250
rect 58585 2680 58590 3250
rect 58560 2670 58590 2680
rect 58615 3250 58645 3260
rect 58615 2680 58620 3250
rect 58640 2680 58645 3250
rect 58615 2670 58645 2680
rect 58670 3250 58700 3260
rect 58670 2680 58675 3250
rect 58695 2680 58700 3250
rect 58670 2670 58700 2680
rect 58725 3250 58755 3260
rect 58725 2680 58730 3250
rect 58750 2680 58755 3250
rect 58725 2670 58755 2680
rect 58780 3250 58810 3260
rect 58780 2680 58785 3250
rect 58805 2680 58810 3250
rect 58780 2670 58810 2680
rect 58835 3250 58865 3260
rect 58835 2680 58840 3250
rect 58860 2680 58865 3250
rect 58835 2670 58865 2680
rect 58890 3250 58920 3260
rect 58890 2680 58895 3250
rect 58915 2680 58920 3250
rect 58890 2670 58920 2680
rect 58945 3250 59015 3260
rect 58945 2680 58950 3250
rect 58970 2680 58990 3250
rect 59010 2680 59015 3250
rect 59105 2710 59246 2720
rect 59105 2690 59110 2710
rect 59130 2690 59165 2710
rect 59185 2690 59220 2710
rect 59240 2690 59246 2710
rect 59105 2680 59246 2690
rect 58945 2670 59015 2680
rect 55155 2640 55185 2650
rect 58615 2640 58645 2650
rect 55155 2620 55160 2640
rect 55180 2620 55185 2640
rect 55155 2610 55185 2620
rect 56850 2630 56890 2640
rect 56850 2610 56860 2630
rect 56880 2610 56890 2630
rect 56850 2600 56890 2610
rect 56935 2630 56975 2640
rect 56935 2610 56945 2630
rect 56965 2610 56975 2630
rect 58615 2620 58620 2640
rect 58640 2620 58645 2640
rect 58615 2610 58645 2620
rect 56935 2600 56975 2610
rect 55150 2575 55190 2585
rect 55150 2555 55160 2575
rect 55180 2555 55190 2575
rect 55150 2535 55190 2555
rect 55150 2515 55160 2535
rect 55180 2515 55190 2535
rect 55150 2495 55190 2515
rect 55150 2475 55160 2495
rect 55180 2475 55190 2495
rect 55150 2465 55190 2475
rect 56735 2570 56805 2580
rect 56735 2350 56740 2570
rect 56760 2350 56780 2570
rect 56800 2350 56805 2570
rect 56735 2340 56805 2350
rect 56830 2570 56860 2580
rect 56830 2350 56835 2570
rect 56855 2350 56860 2570
rect 56830 2340 56860 2350
rect 56885 2570 56915 2580
rect 56885 2350 56890 2570
rect 56910 2350 56915 2570
rect 56885 2340 56915 2350
rect 56940 2570 56970 2580
rect 56940 2350 56945 2570
rect 56965 2350 56970 2570
rect 56940 2340 56970 2350
rect 56995 2570 57065 2580
rect 56995 2350 57000 2570
rect 57020 2350 57040 2570
rect 57060 2350 57065 2570
rect 58610 2575 58650 2585
rect 58610 2555 58620 2575
rect 58640 2555 58650 2575
rect 58610 2535 58650 2555
rect 58610 2515 58620 2535
rect 58640 2515 58650 2535
rect 58610 2495 58650 2515
rect 58610 2475 58620 2495
rect 58640 2475 58650 2495
rect 58610 2465 58650 2475
rect 56995 2340 57065 2350
rect 56770 2310 56810 2320
rect 56770 2290 56780 2310
rect 56800 2290 56810 2310
rect 56770 2280 56810 2290
rect 56990 2310 57030 2320
rect 56990 2290 57000 2310
rect 57020 2290 57030 2310
rect 56990 2280 57030 2290
rect 55995 2265 56025 2275
rect 55995 2245 56000 2265
rect 56020 2245 56025 2265
rect 55995 2235 56025 2245
rect 56690 2265 56720 2275
rect 56690 2245 56695 2265
rect 56715 2245 56720 2265
rect 56690 2235 56720 2245
rect 57080 2265 57110 2275
rect 57080 2245 57085 2265
rect 57105 2245 57110 2265
rect 57080 2235 57110 2245
rect 54825 2210 54855 2220
rect 54825 2190 54830 2210
rect 54850 2190 54855 2210
rect 54825 2180 54855 2190
rect 55485 2210 55515 2220
rect 55485 2190 55490 2210
rect 55510 2190 55515 2210
rect 55485 2180 55515 2190
rect 58285 2210 58315 2220
rect 58285 2190 58290 2210
rect 58310 2190 58315 2210
rect 58285 2180 58315 2190
rect 58945 2210 58975 2220
rect 58945 2190 58950 2210
rect 58970 2190 58975 2210
rect 58945 2180 58975 2190
rect 55995 2165 56065 2175
rect 54785 2150 54855 2160
rect 54460 2016 54675 2036
rect 54460 1999 54495 2016
rect 54640 1999 54675 2016
rect 54555 1949 54580 1999
rect 54785 1980 54790 2150
rect 54810 1980 54830 2150
rect 54850 1980 54855 2150
rect 54785 1970 54855 1980
rect 54880 2150 54910 2160
rect 54880 1980 54885 2150
rect 54905 1980 54910 2150
rect 54880 1970 54910 1980
rect 54935 2150 54965 2160
rect 54935 1980 54940 2150
rect 54960 1980 54965 2150
rect 54935 1970 54965 1980
rect 54990 2150 55020 2160
rect 54990 1980 54995 2150
rect 55015 1980 55020 2150
rect 54990 1970 55020 1980
rect 55045 2150 55075 2160
rect 55045 1980 55050 2150
rect 55070 1980 55075 2150
rect 55045 1970 55075 1980
rect 55100 2150 55130 2160
rect 55100 1980 55105 2150
rect 55125 1980 55130 2150
rect 55100 1970 55130 1980
rect 55155 2150 55185 2160
rect 55155 1980 55160 2150
rect 55180 1980 55185 2150
rect 55155 1970 55185 1980
rect 55210 2150 55240 2160
rect 55210 1980 55215 2150
rect 55235 1980 55240 2150
rect 55210 1970 55240 1980
rect 55265 2150 55295 2160
rect 55265 1980 55270 2150
rect 55290 1980 55295 2150
rect 55265 1970 55295 1980
rect 55320 2150 55350 2160
rect 55320 1980 55325 2150
rect 55345 1980 55350 2150
rect 55320 1970 55350 1980
rect 55375 2150 55405 2160
rect 55375 1980 55380 2150
rect 55400 1980 55405 2150
rect 55375 1970 55405 1980
rect 55430 2150 55460 2160
rect 55430 1980 55435 2150
rect 55455 1980 55460 2150
rect 55430 1970 55460 1980
rect 55485 2150 55555 2160
rect 55485 1980 55490 2150
rect 55510 1980 55530 2150
rect 55550 1980 55555 2150
rect 55995 2045 56000 2165
rect 56020 2045 56040 2165
rect 56060 2045 56065 2165
rect 55995 2035 56065 2045
rect 56090 2165 56120 2175
rect 56090 2045 56095 2165
rect 56115 2045 56120 2165
rect 56090 2035 56120 2045
rect 56145 2165 56175 2175
rect 56145 2045 56150 2165
rect 56170 2045 56175 2165
rect 56145 2035 56175 2045
rect 56200 2165 56230 2175
rect 56200 2045 56205 2165
rect 56225 2045 56230 2165
rect 56200 2035 56230 2045
rect 56255 2165 56285 2175
rect 56255 2045 56260 2165
rect 56280 2045 56285 2165
rect 56255 2035 56285 2045
rect 56310 2165 56340 2175
rect 56310 2045 56315 2165
rect 56335 2045 56340 2165
rect 56310 2035 56340 2045
rect 56365 2165 56395 2175
rect 56365 2045 56370 2165
rect 56390 2045 56395 2165
rect 56365 2035 56395 2045
rect 56420 2165 56450 2175
rect 56420 2045 56425 2165
rect 56445 2045 56450 2165
rect 56420 2035 56450 2045
rect 56475 2165 56505 2175
rect 56475 2045 56480 2165
rect 56500 2045 56505 2165
rect 56475 2035 56505 2045
rect 56530 2165 56560 2175
rect 56530 2045 56535 2165
rect 56555 2045 56560 2165
rect 56530 2035 56560 2045
rect 56585 2165 56615 2175
rect 56585 2045 56590 2165
rect 56610 2045 56615 2165
rect 56585 2035 56615 2045
rect 56640 2165 56670 2175
rect 56640 2045 56645 2165
rect 56665 2045 56670 2165
rect 56640 2035 56670 2045
rect 56695 2165 56765 2175
rect 56695 2045 56700 2165
rect 56720 2045 56740 2165
rect 56760 2045 56765 2165
rect 56695 2035 56765 2045
rect 57035 2165 57105 2175
rect 57035 2045 57040 2165
rect 57060 2045 57080 2165
rect 57100 2045 57105 2165
rect 57035 2035 57105 2045
rect 57130 2165 57160 2175
rect 57130 2045 57135 2165
rect 57155 2045 57160 2165
rect 57130 2035 57160 2045
rect 57185 2165 57215 2175
rect 57185 2045 57190 2165
rect 57210 2045 57215 2165
rect 57185 2035 57215 2045
rect 57240 2165 57270 2175
rect 57240 2045 57245 2165
rect 57265 2045 57270 2165
rect 57240 2035 57270 2045
rect 57295 2165 57325 2175
rect 57295 2045 57300 2165
rect 57320 2045 57325 2165
rect 57295 2035 57325 2045
rect 57350 2165 57380 2175
rect 57350 2045 57355 2165
rect 57375 2045 57380 2165
rect 57350 2035 57380 2045
rect 57405 2165 57435 2175
rect 57405 2045 57410 2165
rect 57430 2045 57435 2165
rect 57405 2035 57435 2045
rect 57460 2165 57490 2175
rect 57460 2045 57465 2165
rect 57485 2045 57490 2165
rect 57460 2035 57490 2045
rect 57515 2165 57545 2175
rect 57515 2045 57520 2165
rect 57540 2045 57545 2165
rect 57515 2035 57545 2045
rect 57570 2165 57600 2175
rect 57570 2045 57575 2165
rect 57595 2045 57600 2165
rect 57570 2035 57600 2045
rect 57625 2165 57655 2175
rect 57625 2045 57630 2165
rect 57650 2045 57655 2165
rect 57625 2035 57655 2045
rect 57680 2165 57710 2175
rect 57680 2045 57685 2165
rect 57705 2045 57710 2165
rect 57680 2035 57710 2045
rect 57735 2165 57805 2175
rect 57735 2045 57740 2165
rect 57760 2045 57780 2165
rect 57800 2045 57805 2165
rect 57735 2035 57805 2045
rect 58245 2150 58315 2160
rect 55485 1970 55555 1980
rect 56035 2005 56065 2035
rect 56035 1985 56040 2005
rect 56060 1985 56065 2005
rect 56035 1975 56065 1985
rect 56695 2005 56725 2015
rect 56695 1985 56700 2005
rect 56720 1985 56725 2005
rect 56695 1975 56725 1985
rect 57075 2005 57105 2015
rect 57075 1985 57080 2005
rect 57100 1985 57105 2005
rect 57075 1975 57105 1985
rect 57735 2005 57765 2035
rect 57735 1985 57740 2005
rect 57760 1985 57765 2005
rect 57735 1975 57765 1985
rect 58245 1980 58250 2150
rect 58270 1980 58290 2150
rect 58310 1980 58315 2150
rect 58245 1970 58315 1980
rect 58340 2150 58370 2160
rect 58340 1980 58345 2150
rect 58365 1980 58370 2150
rect 58340 1970 58370 1980
rect 58395 2150 58425 2160
rect 58395 1980 58400 2150
rect 58420 1980 58425 2150
rect 58395 1970 58425 1980
rect 58450 2150 58480 2160
rect 58450 1980 58455 2150
rect 58475 1980 58480 2150
rect 58450 1970 58480 1980
rect 58505 2150 58535 2160
rect 58505 1980 58510 2150
rect 58530 1980 58535 2150
rect 58505 1970 58535 1980
rect 58560 2150 58590 2160
rect 58560 1980 58565 2150
rect 58585 1980 58590 2150
rect 58560 1970 58590 1980
rect 58615 2150 58645 2160
rect 58615 1980 58620 2150
rect 58640 1980 58645 2150
rect 58615 1970 58645 1980
rect 58670 2150 58700 2160
rect 58670 1980 58675 2150
rect 58695 1980 58700 2150
rect 58670 1970 58700 1980
rect 58725 2150 58755 2160
rect 58725 1980 58730 2150
rect 58750 1980 58755 2150
rect 58725 1970 58755 1980
rect 58780 2150 58810 2160
rect 58780 1980 58785 2150
rect 58805 1980 58810 2150
rect 58780 1970 58810 1980
rect 58835 2150 58865 2160
rect 58835 1980 58840 2150
rect 58860 1980 58865 2150
rect 58835 1970 58865 1980
rect 58890 2150 58920 2160
rect 58890 1980 58895 2150
rect 58915 1980 58920 2150
rect 58890 1970 58920 1980
rect 58945 2150 59015 2160
rect 58945 1980 58950 2150
rect 58970 1980 58990 2150
rect 59010 1980 59015 2150
rect 58945 1970 59015 1980
rect 59125 2016 59340 2036
rect 59125 1999 59160 2016
rect 59305 1999 59340 2016
rect 54930 1940 54970 1950
rect 54930 1920 54940 1940
rect 54960 1920 54970 1940
rect 54930 1910 54970 1920
rect 55040 1940 55080 1950
rect 55040 1920 55050 1940
rect 55070 1920 55080 1940
rect 55040 1910 55080 1920
rect 55150 1940 55190 1950
rect 55150 1920 55160 1940
rect 55180 1920 55190 1940
rect 55150 1910 55190 1920
rect 55260 1940 55300 1950
rect 55260 1920 55270 1940
rect 55290 1920 55300 1940
rect 55260 1910 55300 1920
rect 55320 1940 55350 1950
rect 55320 1920 55325 1940
rect 55345 1920 55350 1940
rect 55320 1910 55350 1920
rect 55370 1940 55410 1950
rect 55370 1920 55380 1940
rect 55400 1920 55410 1940
rect 55370 1910 55410 1920
rect 58390 1940 58430 1950
rect 58390 1920 58400 1940
rect 58420 1920 58430 1940
rect 58390 1910 58430 1920
rect 58450 1940 58480 1950
rect 58450 1920 58455 1940
rect 58475 1920 58480 1940
rect 58450 1910 58480 1920
rect 58500 1940 58540 1950
rect 58500 1920 58510 1940
rect 58530 1920 58540 1940
rect 58500 1910 58540 1920
rect 58610 1940 58650 1950
rect 58610 1920 58620 1940
rect 58640 1920 58650 1940
rect 58610 1910 58650 1920
rect 58720 1940 58760 1950
rect 58720 1920 58730 1940
rect 58750 1920 58760 1940
rect 58720 1910 58760 1920
rect 58830 1940 58870 1950
rect 58830 1920 58840 1940
rect 58860 1920 58870 1940
rect 58830 1910 58870 1920
rect 55315 1875 55355 1885
rect 55315 1855 55325 1875
rect 55345 1855 55355 1875
rect 55315 1835 55355 1855
rect 55315 1815 55325 1835
rect 55345 1815 55355 1835
rect 55315 1805 55355 1815
rect 58445 1875 58485 1885
rect 58445 1855 58455 1875
rect 58475 1855 58485 1875
rect 58445 1835 58485 1855
rect 58445 1815 58455 1835
rect 58475 1815 58485 1835
rect 58445 1805 58485 1815
rect 56040 1780 56070 1790
rect 55320 1770 55350 1780
rect 55320 1750 55325 1770
rect 55345 1750 55350 1770
rect 56040 1760 56045 1780
rect 56065 1760 56070 1780
rect 56040 1750 56070 1760
rect 56690 1780 56720 1790
rect 56690 1760 56695 1780
rect 56715 1760 56720 1780
rect 56690 1750 56720 1760
rect 56850 1780 56880 1790
rect 56850 1760 56855 1780
rect 56875 1760 56880 1780
rect 56850 1750 56880 1760
rect 56903 1780 56933 1790
rect 56903 1760 56908 1780
rect 56928 1760 56933 1780
rect 56903 1750 56933 1760
rect 57080 1780 57110 1790
rect 57080 1760 57085 1780
rect 57105 1760 57110 1780
rect 57080 1750 57110 1760
rect 57730 1780 57760 1790
rect 57730 1760 57735 1780
rect 57755 1760 57760 1780
rect 57730 1750 57760 1760
rect 58450 1770 58480 1780
rect 59220 1949 59245 1999
rect 58450 1750 58455 1770
rect 58475 1750 58480 1770
rect 55320 1740 55350 1750
rect 58450 1740 58480 1750
rect 54785 1710 54855 1720
rect 54460 1390 54495 1400
rect 54460 1365 54465 1390
rect 54490 1365 54495 1390
rect 54460 1355 54495 1365
rect 54520 1390 54555 1400
rect 54520 1365 54525 1390
rect 54550 1365 54555 1390
rect 54520 1355 54555 1365
rect 54580 1390 54615 1400
rect 54580 1365 54585 1390
rect 54610 1365 54615 1390
rect 54580 1355 54615 1365
rect 54785 1440 54790 1710
rect 54810 1440 54830 1710
rect 54850 1440 54855 1710
rect 54785 1430 54855 1440
rect 54880 1710 54910 1720
rect 54880 1440 54885 1710
rect 54905 1440 54910 1710
rect 54880 1430 54910 1440
rect 54935 1710 54965 1720
rect 54935 1440 54940 1710
rect 54960 1440 54965 1710
rect 54935 1430 54965 1440
rect 54990 1710 55020 1720
rect 54990 1440 54995 1710
rect 55015 1440 55020 1710
rect 54990 1430 55020 1440
rect 55045 1710 55075 1720
rect 55045 1440 55050 1710
rect 55070 1440 55075 1710
rect 55045 1430 55075 1440
rect 55100 1710 55130 1720
rect 55100 1440 55105 1710
rect 55125 1440 55130 1710
rect 55100 1430 55130 1440
rect 55155 1710 55185 1720
rect 55155 1440 55160 1710
rect 55180 1440 55185 1710
rect 55155 1430 55185 1440
rect 55210 1710 55240 1720
rect 55210 1440 55215 1710
rect 55235 1440 55240 1710
rect 55210 1430 55240 1440
rect 55265 1710 55295 1720
rect 55265 1440 55270 1710
rect 55290 1440 55295 1710
rect 55265 1430 55295 1440
rect 55320 1710 55350 1720
rect 55320 1440 55325 1710
rect 55345 1440 55350 1710
rect 55320 1430 55350 1440
rect 55375 1710 55405 1720
rect 55375 1440 55380 1710
rect 55400 1440 55405 1710
rect 55375 1430 55405 1440
rect 55430 1710 55460 1720
rect 55430 1440 55435 1710
rect 55455 1440 55460 1710
rect 55430 1430 55460 1440
rect 55485 1710 55555 1720
rect 55485 1440 55490 1710
rect 55510 1440 55530 1710
rect 55550 1440 55555 1710
rect 58245 1710 58315 1720
rect 55995 1695 56065 1705
rect 55995 1575 56000 1695
rect 56020 1575 56040 1695
rect 56060 1575 56065 1695
rect 55995 1565 56065 1575
rect 56090 1695 56120 1705
rect 56090 1575 56095 1695
rect 56115 1575 56120 1695
rect 56090 1565 56120 1575
rect 56145 1695 56175 1705
rect 56145 1575 56150 1695
rect 56170 1575 56175 1695
rect 56145 1565 56175 1575
rect 56200 1695 56230 1705
rect 56200 1575 56205 1695
rect 56225 1575 56230 1695
rect 56200 1565 56230 1575
rect 56255 1695 56285 1705
rect 56255 1575 56260 1695
rect 56280 1575 56285 1695
rect 56255 1565 56285 1575
rect 56310 1695 56340 1705
rect 56310 1575 56315 1695
rect 56335 1575 56340 1695
rect 56310 1565 56340 1575
rect 56365 1695 56395 1705
rect 56365 1575 56370 1695
rect 56390 1575 56395 1695
rect 56365 1565 56395 1575
rect 56420 1695 56450 1705
rect 56420 1575 56425 1695
rect 56445 1575 56450 1695
rect 56420 1565 56450 1575
rect 56475 1695 56505 1705
rect 56475 1575 56480 1695
rect 56500 1575 56505 1695
rect 56475 1565 56505 1575
rect 56530 1695 56560 1705
rect 56530 1575 56535 1695
rect 56555 1575 56560 1695
rect 56530 1565 56560 1575
rect 56585 1695 56615 1705
rect 56585 1575 56590 1695
rect 56610 1575 56615 1695
rect 56585 1565 56615 1575
rect 56640 1695 56670 1705
rect 56640 1575 56645 1695
rect 56665 1575 56670 1695
rect 56640 1565 56670 1575
rect 56695 1695 56805 1705
rect 56695 1575 56700 1695
rect 56720 1575 56740 1695
rect 56760 1575 56780 1695
rect 56800 1575 56805 1695
rect 56695 1565 56805 1575
rect 56830 1695 56860 1705
rect 56830 1575 56835 1695
rect 56855 1575 56860 1695
rect 56830 1565 56860 1575
rect 56885 1695 56915 1705
rect 56885 1575 56890 1695
rect 56910 1575 56915 1695
rect 56885 1565 56915 1575
rect 56940 1695 56970 1705
rect 56940 1575 56945 1695
rect 56965 1575 56970 1695
rect 56940 1565 56970 1575
rect 56995 1695 57105 1705
rect 56995 1575 57000 1695
rect 57020 1575 57040 1695
rect 57060 1575 57080 1695
rect 57100 1575 57105 1695
rect 56995 1565 57105 1575
rect 57130 1695 57160 1705
rect 57130 1575 57135 1695
rect 57155 1575 57160 1695
rect 57130 1565 57160 1575
rect 57185 1695 57215 1705
rect 57185 1575 57190 1695
rect 57210 1575 57215 1695
rect 57185 1565 57215 1575
rect 57240 1695 57270 1705
rect 57240 1575 57245 1695
rect 57265 1575 57270 1695
rect 57240 1565 57270 1575
rect 57295 1695 57325 1705
rect 57295 1575 57300 1695
rect 57320 1575 57325 1695
rect 57295 1565 57325 1575
rect 57350 1695 57380 1705
rect 57350 1575 57355 1695
rect 57375 1575 57380 1695
rect 57350 1565 57380 1575
rect 57405 1695 57435 1705
rect 57405 1575 57410 1695
rect 57430 1575 57435 1695
rect 57405 1565 57435 1575
rect 57460 1695 57490 1705
rect 57460 1575 57465 1695
rect 57485 1575 57490 1695
rect 57460 1565 57490 1575
rect 57515 1695 57545 1705
rect 57515 1575 57520 1695
rect 57540 1575 57545 1695
rect 57515 1565 57545 1575
rect 57570 1695 57600 1705
rect 57570 1575 57575 1695
rect 57595 1575 57600 1695
rect 57570 1565 57600 1575
rect 57625 1695 57655 1705
rect 57625 1575 57630 1695
rect 57650 1575 57655 1695
rect 57625 1565 57655 1575
rect 57680 1695 57710 1705
rect 57680 1575 57685 1695
rect 57705 1575 57710 1695
rect 57680 1565 57710 1575
rect 57735 1695 57805 1705
rect 57735 1575 57740 1695
rect 57760 1575 57780 1695
rect 57800 1575 57805 1695
rect 57735 1565 57805 1575
rect 56040 1545 56065 1565
rect 56035 1535 56065 1545
rect 56035 1515 56040 1535
rect 56060 1515 56065 1535
rect 56035 1505 56065 1515
rect 56735 1535 56765 1545
rect 56735 1515 56740 1535
rect 56760 1515 56765 1535
rect 56735 1505 56765 1515
rect 57035 1535 57065 1545
rect 57035 1515 57040 1535
rect 57060 1515 57065 1535
rect 57035 1505 57065 1515
rect 57735 1535 57765 1565
rect 57735 1515 57740 1535
rect 57760 1515 57765 1535
rect 57735 1505 57765 1515
rect 55485 1430 55555 1440
rect 58245 1440 58250 1710
rect 58270 1440 58290 1710
rect 58310 1440 58315 1710
rect 58245 1430 58315 1440
rect 58340 1710 58370 1720
rect 58340 1440 58345 1710
rect 58365 1440 58370 1710
rect 58340 1430 58370 1440
rect 58395 1710 58425 1720
rect 58395 1440 58400 1710
rect 58420 1440 58425 1710
rect 58395 1430 58425 1440
rect 58450 1710 58480 1720
rect 58450 1440 58455 1710
rect 58475 1440 58480 1710
rect 58450 1430 58480 1440
rect 58505 1710 58535 1720
rect 58505 1440 58510 1710
rect 58530 1440 58535 1710
rect 58505 1430 58535 1440
rect 58560 1710 58590 1720
rect 58560 1440 58565 1710
rect 58585 1440 58590 1710
rect 58560 1430 58590 1440
rect 58615 1710 58645 1720
rect 58615 1440 58620 1710
rect 58640 1440 58645 1710
rect 58615 1430 58645 1440
rect 58670 1710 58700 1720
rect 58670 1440 58675 1710
rect 58695 1440 58700 1710
rect 58670 1430 58700 1440
rect 58725 1710 58755 1720
rect 58725 1440 58730 1710
rect 58750 1440 58755 1710
rect 58725 1430 58755 1440
rect 58780 1710 58810 1720
rect 58780 1440 58785 1710
rect 58805 1440 58810 1710
rect 58780 1430 58810 1440
rect 58835 1710 58865 1720
rect 58835 1440 58840 1710
rect 58860 1440 58865 1710
rect 58835 1430 58865 1440
rect 58890 1710 58920 1720
rect 58890 1440 58895 1710
rect 58915 1440 58920 1710
rect 58890 1430 58920 1440
rect 58945 1710 59015 1720
rect 58945 1440 58950 1710
rect 58970 1440 58990 1710
rect 59010 1440 59015 1710
rect 58945 1430 59015 1440
rect 54640 1390 54675 1400
rect 54640 1365 54645 1390
rect 54670 1365 54675 1390
rect 54825 1400 54855 1410
rect 54825 1380 54830 1400
rect 54850 1380 54855 1400
rect 54825 1370 54855 1380
rect 55485 1400 55515 1410
rect 55485 1380 55490 1400
rect 55510 1380 55515 1400
rect 55485 1370 55515 1380
rect 58285 1400 58315 1410
rect 58285 1380 58290 1400
rect 58310 1380 58315 1400
rect 58285 1370 58315 1380
rect 58945 1400 58975 1410
rect 58945 1380 58950 1400
rect 58970 1380 58975 1400
rect 58945 1370 58975 1380
rect 59125 1390 59160 1400
rect 54640 1355 54675 1365
rect 59125 1365 59130 1390
rect 59155 1365 59160 1390
rect 59125 1355 59160 1365
rect 59185 1390 59220 1400
rect 59185 1365 59190 1390
rect 59215 1365 59220 1390
rect 59185 1355 59220 1365
rect 59245 1390 59280 1400
rect 59245 1365 59250 1390
rect 59275 1365 59280 1390
rect 59245 1355 59280 1365
rect 59305 1390 59340 1400
rect 59305 1365 59310 1390
rect 59335 1365 59340 1390
rect 59305 1355 59340 1365
rect 55180 1235 55220 1245
rect 55180 1215 55190 1235
rect 55210 1215 55220 1235
rect 55180 1205 55220 1215
rect 58580 1235 58620 1245
rect 58580 1215 58590 1235
rect 58610 1215 58620 1235
rect 58580 1205 58620 1215
rect 57390 1110 57430 1120
rect 57390 1090 57400 1110
rect 57420 1090 57430 1110
rect 57390 1080 57430 1090
rect 56830 1055 56860 1065
rect 54600 1045 54635 1055
rect 54600 1020 54605 1045
rect 54630 1020 54635 1045
rect 54600 1010 54635 1020
rect 54660 1045 54695 1055
rect 54660 1020 54665 1045
rect 54690 1020 54695 1045
rect 54660 1010 54695 1020
rect 54795 1040 54865 1050
rect 54635 323 54660 373
rect 54795 370 54800 1040
rect 54820 370 54840 1040
rect 54860 370 54865 1040
rect 54795 360 54865 370
rect 54935 1040 54965 1050
rect 54935 370 54940 1040
rect 54960 370 54965 1040
rect 54935 360 54965 370
rect 55035 1040 55065 1050
rect 55035 370 55040 1040
rect 55060 370 55065 1040
rect 55035 360 55065 370
rect 55135 1040 55165 1050
rect 55135 370 55140 1040
rect 55160 370 55165 1040
rect 55135 360 55165 370
rect 55235 1040 55265 1050
rect 55235 370 55240 1040
rect 55260 370 55265 1040
rect 55235 360 55265 370
rect 55335 1040 55365 1050
rect 55335 370 55340 1040
rect 55360 370 55365 1040
rect 55335 360 55365 370
rect 55435 1040 55505 1050
rect 55435 370 55440 1040
rect 55460 370 55480 1040
rect 55500 370 55505 1040
rect 56830 1035 56835 1055
rect 56855 1035 56860 1055
rect 56830 1025 56860 1035
rect 58295 1040 58365 1050
rect 56185 995 56255 1005
rect 56185 775 56190 995
rect 56210 775 56230 995
rect 56250 775 56255 995
rect 56185 765 56255 775
rect 56280 995 56310 1005
rect 56280 775 56285 995
rect 56305 775 56310 995
rect 56280 765 56310 775
rect 56335 995 56365 1005
rect 56335 775 56340 995
rect 56360 775 56365 995
rect 56335 765 56365 775
rect 56390 995 56420 1005
rect 56390 775 56395 995
rect 56415 775 56420 995
rect 56390 765 56420 775
rect 56445 995 56475 1005
rect 56445 775 56450 995
rect 56470 775 56475 995
rect 56445 765 56475 775
rect 56500 995 56530 1005
rect 56500 775 56505 995
rect 56525 775 56530 995
rect 56500 765 56530 775
rect 56555 995 56585 1005
rect 56555 775 56560 995
rect 56580 775 56585 995
rect 56555 765 56585 775
rect 56610 995 56640 1005
rect 56610 775 56615 995
rect 56635 775 56640 995
rect 56610 765 56640 775
rect 56665 995 56695 1005
rect 56665 775 56670 995
rect 56690 775 56695 995
rect 56665 765 56695 775
rect 56720 995 56750 1005
rect 56720 775 56725 995
rect 56745 775 56750 995
rect 56720 765 56750 775
rect 56775 995 56805 1005
rect 56775 775 56780 995
rect 56800 775 56805 995
rect 56775 765 56805 775
rect 56830 995 56860 1005
rect 56830 775 56835 995
rect 56855 775 56860 995
rect 56830 765 56860 775
rect 56885 995 56915 1005
rect 56885 775 56890 995
rect 56910 775 56915 995
rect 56885 765 56915 775
rect 56940 995 56970 1005
rect 56940 775 56945 995
rect 56965 775 56970 995
rect 56940 765 56970 775
rect 56995 995 57025 1005
rect 56995 775 57000 995
rect 57020 775 57025 995
rect 56995 765 57025 775
rect 57050 995 57080 1005
rect 57050 775 57055 995
rect 57075 775 57080 995
rect 57050 765 57080 775
rect 57105 995 57135 1005
rect 57105 775 57110 995
rect 57130 775 57135 995
rect 57105 765 57135 775
rect 57160 995 57190 1005
rect 57160 775 57165 995
rect 57185 775 57190 995
rect 57160 765 57190 775
rect 57215 995 57245 1005
rect 57215 775 57220 995
rect 57240 775 57245 995
rect 57215 765 57245 775
rect 57270 995 57300 1005
rect 57270 775 57275 995
rect 57295 775 57300 995
rect 57270 765 57300 775
rect 57325 995 57355 1005
rect 57325 775 57330 995
rect 57350 775 57355 995
rect 57325 765 57355 775
rect 57380 995 57410 1005
rect 57380 775 57385 995
rect 57405 775 57410 995
rect 57380 765 57410 775
rect 57435 995 57465 1005
rect 57435 775 57440 995
rect 57460 775 57465 995
rect 57435 765 57465 775
rect 57490 995 57560 1005
rect 57490 775 57495 995
rect 57515 775 57535 995
rect 57555 775 57560 995
rect 57490 765 57560 775
rect 56220 735 56260 745
rect 56220 715 56230 735
rect 56250 715 56260 735
rect 56220 705 56260 715
rect 57485 735 57525 745
rect 57485 715 57495 735
rect 57515 715 57525 735
rect 57485 705 57525 715
rect 56595 590 56635 600
rect 56595 570 56605 590
rect 56625 570 56635 590
rect 56595 560 56635 570
rect 57040 590 57080 600
rect 57040 570 57050 590
rect 57070 570 57080 590
rect 57040 560 57080 570
rect 56395 530 56465 540
rect 56395 410 56400 530
rect 56420 410 56440 530
rect 56460 410 56465 530
rect 56395 400 56465 410
rect 56490 530 56520 540
rect 56490 410 56495 530
rect 56515 410 56520 530
rect 56490 400 56520 410
rect 56545 530 56575 540
rect 56545 410 56550 530
rect 56570 410 56575 530
rect 56545 400 56575 410
rect 56600 530 56630 540
rect 56600 410 56605 530
rect 56625 410 56630 530
rect 56600 400 56630 410
rect 56655 530 56685 540
rect 56655 410 56660 530
rect 56680 410 56685 530
rect 56655 400 56685 410
rect 56710 530 56740 540
rect 56710 410 56715 530
rect 56735 410 56740 530
rect 56710 400 56740 410
rect 56765 530 56835 540
rect 56765 410 56770 530
rect 56790 410 56810 530
rect 56830 410 56835 530
rect 56765 400 56835 410
rect 56875 530 56905 540
rect 56875 410 56880 530
rect 56900 410 56905 530
rect 56875 400 56905 410
rect 57215 530 57245 540
rect 57215 410 57220 530
rect 57240 410 57245 530
rect 57215 400 57245 410
rect 55435 360 55505 370
rect 56435 370 56465 380
rect 56435 350 56440 370
rect 56460 350 56465 370
rect 56435 340 56465 350
rect 56765 370 56795 380
rect 56765 350 56770 370
rect 56790 350 56795 370
rect 58295 370 58300 1040
rect 58320 370 58340 1040
rect 58360 370 58365 1040
rect 58295 360 58365 370
rect 58435 1040 58465 1050
rect 58435 370 58440 1040
rect 58460 370 58465 1040
rect 58435 360 58465 370
rect 58535 1040 58565 1050
rect 58535 370 58540 1040
rect 58560 370 58565 1040
rect 58535 360 58565 370
rect 58635 1040 58665 1050
rect 58635 370 58640 1040
rect 58660 370 58665 1040
rect 58635 360 58665 370
rect 58735 1040 58765 1050
rect 58735 370 58740 1040
rect 58760 370 58765 1040
rect 58735 360 58765 370
rect 58835 1040 58865 1050
rect 58835 370 58840 1040
rect 58860 370 58865 1040
rect 58835 360 58865 370
rect 58935 1040 59005 1050
rect 58935 370 58940 1040
rect 58960 370 58980 1040
rect 59000 370 59005 1040
rect 59105 1045 59140 1055
rect 59105 1020 59110 1045
rect 59135 1020 59140 1045
rect 59105 1010 59140 1020
rect 59165 1045 59200 1055
rect 59165 1020 59170 1045
rect 59195 1020 59200 1045
rect 59165 1010 59200 1020
rect 58935 360 59005 370
rect 56765 340 56795 350
rect 54835 330 54865 340
rect 54835 310 54840 330
rect 54860 310 54865 330
rect 54835 300 54865 310
rect 55435 330 55465 340
rect 55435 310 55440 330
rect 55460 310 55465 330
rect 55435 300 55465 310
rect 58335 330 58365 340
rect 58335 310 58340 330
rect 58360 310 58365 330
rect 58335 300 58365 310
rect 58935 330 58965 340
rect 58935 310 58940 330
rect 58960 310 58965 330
rect 59140 323 59165 373
rect 58935 300 58965 310
<< viali >>
rect 56095 4940 56115 4960
rect 56275 4940 56295 4960
rect 57035 4940 57055 4960
rect 57215 4940 57235 4960
rect 57505 4940 57525 4960
rect 57685 4940 57705 4960
rect 56095 4580 56115 4900
rect 56155 4580 56175 4900
rect 56215 4580 56235 4900
rect 56275 4580 56295 4900
rect 56565 4770 56585 4790
rect 56745 4770 56765 4790
rect 56565 4580 56585 4730
rect 56625 4580 56645 4730
rect 56685 4580 56705 4730
rect 56745 4580 56765 4730
rect 57035 4580 57055 4900
rect 57095 4580 57115 4900
rect 57155 4580 57175 4900
rect 57215 4580 57235 4900
rect 57505 4580 57525 4900
rect 57565 4580 57585 4900
rect 57625 4580 57645 4900
rect 57685 4580 57705 4900
rect 56160 4490 56180 4510
rect 56635 4490 56655 4510
rect 57145 4490 57165 4510
rect 57581 4480 57601 4500
rect 54930 3705 54950 4025
rect 54990 3705 55010 4025
rect 55050 3705 55070 4025
rect 55110 3705 55130 4025
rect 55170 3705 55190 4025
rect 55230 3705 55250 4025
rect 55290 3705 55310 4025
rect 55350 3705 55370 4025
rect 55410 3705 55430 4025
rect 55470 3705 55490 4025
rect 55530 3705 55550 4025
rect 55590 3705 55610 4025
rect 55650 3705 55670 4025
rect 56015 3705 56035 4025
rect 56075 3705 56095 4025
rect 56135 3705 56155 4025
rect 56195 3705 56215 4025
rect 56255 3705 56275 4025
rect 56315 3705 56335 4025
rect 56375 3705 56395 4025
rect 56435 3705 56455 4025
rect 56495 3705 56515 4025
rect 56555 3705 56575 4025
rect 56615 3705 56635 4025
rect 56675 3705 56695 4025
rect 56735 3705 56755 4025
rect 57045 3705 57065 4025
rect 57105 3705 57125 4025
rect 57165 3705 57185 4025
rect 57225 3705 57245 4025
rect 57285 3705 57305 4025
rect 57345 3705 57365 4025
rect 57405 3705 57425 4025
rect 57465 3705 57485 4025
rect 57525 3705 57545 4025
rect 57585 3705 57605 4025
rect 57645 3705 57665 4025
rect 57705 3705 57725 4025
rect 57765 3705 57785 4025
rect 58130 3705 58150 4025
rect 58190 3705 58210 4025
rect 58250 3705 58270 4025
rect 58310 3705 58330 4025
rect 58370 3705 58390 4025
rect 58430 3705 58450 4025
rect 58490 3705 58510 4025
rect 58550 3705 58570 4025
rect 58610 3705 58630 4025
rect 58670 3705 58690 4025
rect 58730 3705 58750 4025
rect 58790 3705 58810 4025
rect 58850 3705 58870 4025
rect 54930 3645 54950 3665
rect 55650 3645 55670 3665
rect 56015 3645 56035 3665
rect 56735 3645 56755 3665
rect 57045 3645 57065 3665
rect 57765 3645 57785 3665
rect 58130 3645 58150 3665
rect 58850 3645 58870 3665
rect 56375 3580 56395 3600
rect 57405 3580 57425 3600
rect 55290 3535 55310 3555
rect 58490 3535 58510 3555
rect 54560 3295 54580 3315
rect 54615 3295 54635 3315
rect 54670 3295 54690 3315
rect 54830 3290 54850 3310
rect 55490 3290 55510 3310
rect 58290 3290 58310 3310
rect 58950 3290 58970 3310
rect 59110 3295 59130 3315
rect 59165 3295 59185 3315
rect 59220 3295 59240 3315
rect 54560 2690 54580 2710
rect 54615 2690 54635 2710
rect 54670 2690 54690 2710
rect 54830 2680 54850 3250
rect 54885 2680 54905 3250
rect 54940 2680 54960 3250
rect 54995 2680 55015 3250
rect 55050 2680 55070 3250
rect 55105 2680 55125 3250
rect 55160 2680 55180 3250
rect 55215 2680 55235 3250
rect 55270 2680 55290 3250
rect 55325 2680 55345 3250
rect 55380 2680 55400 3250
rect 55435 2680 55455 3250
rect 55490 2680 55510 3250
rect 56285 3220 56305 3240
rect 56340 3220 56360 3240
rect 56395 3220 56415 3240
rect 56450 3220 56470 3240
rect 56505 3220 56525 3240
rect 56560 3220 56580 3240
rect 56615 3220 56635 3240
rect 56670 3220 56690 3240
rect 56725 3220 56745 3240
rect 56780 3220 56800 3240
rect 56835 3220 56855 3240
rect 56890 3220 56910 3240
rect 56945 3220 56965 3240
rect 57000 3220 57020 3240
rect 57055 3220 57075 3240
rect 57110 3220 57130 3240
rect 57165 3220 57185 3240
rect 57220 3220 57240 3240
rect 57275 3220 57295 3240
rect 57330 3220 57350 3240
rect 57385 3220 57405 3240
rect 57440 3220 57460 3240
rect 57495 3220 57515 3240
rect 56285 3160 56305 3180
rect 56395 3160 56415 3180
rect 56835 3160 56855 3180
rect 57495 3160 57515 3180
rect 56045 2995 56065 3015
rect 56695 2995 56715 3015
rect 57085 2995 57105 3015
rect 57735 2995 57755 3015
rect 56040 2910 56060 2930
rect 56095 2910 56115 2930
rect 56150 2910 56170 2930
rect 56205 2910 56225 2930
rect 56260 2910 56280 2930
rect 56315 2910 56335 2930
rect 56370 2910 56390 2930
rect 56425 2910 56445 2930
rect 56480 2910 56500 2930
rect 56535 2910 56555 2930
rect 56590 2910 56610 2930
rect 56645 2910 56665 2930
rect 56700 2910 56720 2930
rect 57080 2910 57100 2930
rect 57135 2910 57155 2930
rect 57190 2910 57210 2930
rect 57245 2910 57265 2930
rect 57300 2910 57320 2930
rect 57355 2910 57375 2930
rect 57410 2910 57430 2930
rect 57465 2910 57485 2930
rect 57520 2910 57540 2930
rect 57575 2910 57595 2930
rect 57630 2910 57650 2930
rect 57685 2910 57705 2930
rect 57740 2910 57760 2930
rect 56040 2850 56060 2870
rect 56700 2850 56720 2870
rect 57080 2850 57100 2870
rect 57740 2850 57760 2870
rect 56100 2765 56120 2785
rect 56585 2775 56605 2795
rect 57195 2775 57215 2795
rect 58290 2680 58310 3250
rect 58345 2680 58365 3250
rect 58400 2680 58420 3250
rect 58455 2680 58475 3250
rect 58510 2680 58530 3250
rect 58565 2680 58585 3250
rect 58620 2680 58640 3250
rect 58675 2680 58695 3250
rect 58730 2680 58750 3250
rect 58785 2680 58805 3250
rect 58840 2680 58860 3250
rect 58895 2680 58915 3250
rect 58950 2680 58970 3250
rect 59110 2690 59130 2710
rect 59165 2690 59185 2710
rect 59220 2690 59240 2710
rect 56860 2610 56880 2630
rect 56945 2610 56965 2630
rect 55160 2555 55180 2575
rect 55160 2515 55180 2535
rect 55160 2475 55180 2495
rect 56780 2350 56800 2570
rect 56835 2350 56855 2570
rect 56890 2350 56910 2570
rect 56945 2350 56965 2570
rect 57000 2350 57020 2570
rect 58620 2555 58640 2575
rect 58620 2515 58640 2535
rect 58620 2475 58640 2495
rect 56780 2290 56800 2310
rect 57000 2290 57020 2310
rect 56000 2245 56020 2265
rect 56695 2245 56715 2265
rect 57085 2245 57105 2265
rect 54830 2190 54850 2210
rect 55490 2190 55510 2210
rect 58290 2190 58310 2210
rect 58950 2190 58970 2210
rect 54830 1980 54850 2150
rect 54885 1980 54905 2150
rect 54940 1980 54960 2150
rect 54995 1980 55015 2150
rect 55050 1980 55070 2150
rect 55105 1980 55125 2150
rect 55160 1980 55180 2150
rect 55215 1980 55235 2150
rect 55270 1980 55290 2150
rect 55325 1980 55345 2150
rect 55380 1980 55400 2150
rect 55435 1980 55455 2150
rect 55490 1980 55510 2150
rect 56040 2045 56060 2165
rect 56095 2045 56115 2165
rect 56150 2045 56170 2165
rect 56205 2045 56225 2165
rect 56260 2045 56280 2165
rect 56315 2045 56335 2165
rect 56370 2045 56390 2165
rect 56425 2045 56445 2165
rect 56480 2045 56500 2165
rect 56535 2045 56555 2165
rect 56590 2045 56610 2165
rect 56645 2045 56665 2165
rect 56700 2045 56720 2165
rect 57080 2045 57100 2165
rect 57135 2045 57155 2165
rect 57190 2045 57210 2165
rect 57245 2045 57265 2165
rect 57300 2045 57320 2165
rect 57355 2045 57375 2165
rect 57410 2045 57430 2165
rect 57465 2045 57485 2165
rect 57520 2045 57540 2165
rect 57575 2045 57595 2165
rect 57630 2045 57650 2165
rect 57685 2045 57705 2165
rect 57740 2045 57760 2165
rect 56040 1985 56060 2005
rect 56700 1985 56720 2005
rect 57080 1985 57100 2005
rect 57740 1985 57760 2005
rect 58290 1980 58310 2150
rect 58345 1980 58365 2150
rect 58400 1980 58420 2150
rect 58455 1980 58475 2150
rect 58510 1980 58530 2150
rect 58565 1980 58585 2150
rect 58620 1980 58640 2150
rect 58675 1980 58695 2150
rect 58730 1980 58750 2150
rect 58785 1980 58805 2150
rect 58840 1980 58860 2150
rect 58895 1980 58915 2150
rect 58950 1980 58970 2150
rect 54940 1920 54960 1940
rect 55050 1920 55070 1940
rect 55160 1920 55180 1940
rect 55270 1920 55290 1940
rect 55380 1920 55400 1940
rect 58400 1920 58420 1940
rect 58510 1920 58530 1940
rect 58620 1920 58640 1940
rect 58730 1920 58750 1940
rect 58840 1920 58860 1940
rect 55325 1855 55345 1875
rect 55325 1815 55345 1835
rect 58455 1855 58475 1875
rect 58455 1815 58475 1835
rect 56045 1760 56065 1780
rect 56695 1760 56715 1780
rect 56855 1760 56875 1780
rect 56908 1760 56928 1780
rect 57085 1760 57105 1780
rect 57735 1760 57755 1780
rect 54465 1365 54490 1390
rect 54525 1365 54550 1390
rect 54585 1365 54610 1390
rect 54830 1440 54850 1710
rect 54885 1440 54905 1710
rect 54940 1440 54960 1710
rect 54995 1440 55015 1710
rect 55050 1440 55070 1710
rect 55105 1440 55125 1710
rect 55160 1440 55180 1710
rect 55215 1440 55235 1710
rect 55270 1440 55290 1710
rect 55325 1440 55345 1710
rect 55380 1440 55400 1710
rect 55435 1440 55455 1710
rect 55490 1440 55510 1710
rect 56040 1575 56060 1695
rect 56095 1575 56115 1695
rect 56150 1575 56170 1695
rect 56205 1575 56225 1695
rect 56260 1575 56280 1695
rect 56315 1575 56335 1695
rect 56370 1575 56390 1695
rect 56425 1575 56445 1695
rect 56480 1575 56500 1695
rect 56535 1575 56555 1695
rect 56590 1575 56610 1695
rect 56645 1575 56665 1695
rect 56700 1575 56720 1695
rect 56780 1575 56800 1695
rect 56835 1575 56855 1695
rect 56890 1575 56910 1695
rect 56945 1575 56965 1695
rect 57000 1575 57020 1695
rect 57080 1575 57100 1695
rect 57135 1575 57155 1695
rect 57190 1575 57210 1695
rect 57245 1575 57265 1695
rect 57300 1575 57320 1695
rect 57355 1575 57375 1695
rect 57410 1575 57430 1695
rect 57465 1575 57485 1695
rect 57520 1575 57540 1695
rect 57575 1575 57595 1695
rect 57630 1575 57650 1695
rect 57685 1575 57705 1695
rect 57740 1575 57760 1695
rect 56040 1515 56060 1535
rect 56740 1515 56760 1535
rect 57040 1515 57060 1535
rect 57740 1515 57760 1535
rect 58290 1440 58310 1710
rect 58345 1440 58365 1710
rect 58400 1440 58420 1710
rect 58455 1440 58475 1710
rect 58510 1440 58530 1710
rect 58565 1440 58585 1710
rect 58620 1440 58640 1710
rect 58675 1440 58695 1710
rect 58730 1440 58750 1710
rect 58785 1440 58805 1710
rect 58840 1440 58860 1710
rect 58895 1440 58915 1710
rect 58950 1440 58970 1710
rect 54645 1365 54670 1390
rect 54830 1380 54850 1400
rect 55490 1380 55510 1400
rect 58290 1380 58310 1400
rect 58950 1380 58970 1400
rect 59130 1365 59155 1390
rect 59190 1365 59215 1390
rect 59250 1365 59275 1390
rect 59310 1365 59335 1390
rect 55190 1215 55210 1235
rect 58590 1215 58610 1235
rect 57400 1090 57420 1110
rect 54605 1020 54630 1045
rect 54665 1020 54690 1045
rect 54840 370 54860 1040
rect 54940 370 54960 1040
rect 55040 370 55060 1040
rect 55140 370 55160 1040
rect 55240 370 55260 1040
rect 55340 370 55360 1040
rect 55440 370 55460 1040
rect 56835 1035 56855 1055
rect 56230 775 56250 995
rect 56285 775 56305 995
rect 56340 775 56360 995
rect 56395 775 56415 995
rect 56450 775 56470 995
rect 56505 775 56525 995
rect 56560 775 56580 995
rect 56615 775 56635 995
rect 56670 775 56690 995
rect 56725 775 56745 995
rect 56780 775 56800 995
rect 56835 775 56855 995
rect 56890 775 56910 995
rect 56945 775 56965 995
rect 57000 775 57020 995
rect 57055 775 57075 995
rect 57110 775 57130 995
rect 57165 775 57185 995
rect 57220 775 57240 995
rect 57275 775 57295 995
rect 57330 775 57350 995
rect 57385 775 57405 995
rect 57440 775 57460 995
rect 57495 775 57515 995
rect 56230 715 56250 735
rect 57495 715 57515 735
rect 56605 570 56625 590
rect 57050 570 57070 590
rect 56440 410 56460 530
rect 56495 410 56515 530
rect 56550 410 56570 530
rect 56605 410 56625 530
rect 56660 410 56680 530
rect 56715 410 56735 530
rect 56770 410 56790 530
rect 56880 410 56900 530
rect 57220 410 57240 530
rect 56440 350 56460 370
rect 56770 350 56790 370
rect 58340 370 58360 1040
rect 58440 370 58460 1040
rect 58540 370 58560 1040
rect 58640 370 58660 1040
rect 58740 370 58760 1040
rect 58840 370 58860 1040
rect 58940 370 58960 1040
rect 59110 1020 59135 1045
rect 59170 1020 59195 1045
rect 54840 310 54860 330
rect 55440 310 55460 330
rect 58340 310 58360 330
rect 58940 310 58960 330
<< metal1 >>
rect 52640 4305 52760 6275
rect 52640 4275 52645 4305
rect 52675 4275 52685 4305
rect 52715 4275 52725 4305
rect 52755 4275 52760 4305
rect 52640 4270 52760 4275
rect 52990 4305 53110 6275
rect 52990 4275 52995 4305
rect 53025 4275 53035 4305
rect 53065 4275 53075 4305
rect 53105 4275 53110 4305
rect 52990 4270 53110 4275
rect 53340 4305 53460 6275
rect 53340 4275 53345 4305
rect 53375 4275 53385 4305
rect 53415 4275 53425 4305
rect 53455 4275 53460 4305
rect 53340 4270 53460 4275
rect 53690 4305 53810 6275
rect 53690 4275 53695 4305
rect 53725 4275 53735 4305
rect 53765 4275 53775 4305
rect 53805 4275 53810 4305
rect 53690 4270 53810 4275
rect 54040 4305 54160 6275
rect 54040 4275 54045 4305
rect 54075 4275 54085 4305
rect 54115 4275 54125 4305
rect 54155 4275 54160 4305
rect 54040 4270 54160 4275
rect 54390 4305 54510 6275
rect 54390 4275 54395 4305
rect 54425 4275 54435 4305
rect 54465 4275 54475 4305
rect 54505 4275 54510 4305
rect 54390 4270 54510 4275
rect 54740 4305 54860 6275
rect 54740 4275 54745 4305
rect 54775 4275 54785 4305
rect 54815 4275 54825 4305
rect 54855 4275 54860 4305
rect 54740 4270 54860 4275
rect 55090 4305 55210 6275
rect 55090 4275 55095 4305
rect 55125 4275 55135 4305
rect 55165 4275 55175 4305
rect 55205 4275 55210 4305
rect 55090 4270 55210 4275
rect 55280 4305 55320 4310
rect 55280 4275 55285 4305
rect 55315 4275 55320 4305
rect 54980 4210 55260 4215
rect 54980 4180 54985 4210
rect 55015 4180 55025 4210
rect 55055 4180 55065 4210
rect 55095 4180 55105 4210
rect 55135 4180 55145 4210
rect 55175 4180 55185 4210
rect 55215 4180 55225 4210
rect 55255 4180 55260 4210
rect 54980 4170 55260 4180
rect 54980 4140 54985 4170
rect 55015 4140 55025 4170
rect 55055 4140 55065 4170
rect 55095 4140 55105 4170
rect 55135 4140 55145 4170
rect 55175 4140 55185 4170
rect 55215 4140 55225 4170
rect 55255 4140 55260 4170
rect 54980 4130 55260 4140
rect 54980 4100 54985 4130
rect 55015 4100 55025 4130
rect 55055 4100 55065 4130
rect 55095 4100 55105 4130
rect 55135 4100 55145 4130
rect 55175 4100 55185 4130
rect 55215 4100 55225 4130
rect 55255 4100 55260 4130
rect 54980 4095 55260 4100
rect 54920 4075 54960 4080
rect 54920 4045 54925 4075
rect 54955 4045 54960 4075
rect 54920 4040 54960 4045
rect 54925 4025 54955 4040
rect 54925 3705 54930 4025
rect 54950 3705 54955 4025
rect 54925 3665 54955 3705
rect 54985 4025 55015 4095
rect 55040 4075 55080 4080
rect 55040 4045 55045 4075
rect 55075 4045 55080 4075
rect 55040 4040 55080 4045
rect 54985 3705 54990 4025
rect 55010 3705 55015 4025
rect 54985 3690 55015 3705
rect 55045 4025 55075 4040
rect 55045 3705 55050 4025
rect 55070 3705 55075 4025
rect 55045 3695 55075 3705
rect 55105 4025 55135 4095
rect 55160 4075 55200 4080
rect 55160 4045 55165 4075
rect 55195 4045 55200 4075
rect 55160 4040 55200 4045
rect 55105 3705 55110 4025
rect 55130 3705 55135 4025
rect 55105 3690 55135 3705
rect 55165 4025 55195 4040
rect 55165 3705 55170 4025
rect 55190 3705 55195 4025
rect 55165 3695 55195 3705
rect 55225 4025 55255 4095
rect 55280 4075 55320 4275
rect 55440 4305 55560 6275
rect 55790 4310 55910 6275
rect 56205 5020 56245 5025
rect 56205 4990 56210 5020
rect 56240 4990 56245 5020
rect 56085 4965 56125 4970
rect 56085 4935 56090 4965
rect 56120 4935 56125 4965
rect 56085 4930 56125 4935
rect 56205 4965 56245 4990
rect 56675 5020 56715 5025
rect 56675 4990 56680 5020
rect 56710 4990 56715 5020
rect 56675 4985 56715 4990
rect 56205 4935 56210 4965
rect 56240 4935 56245 4965
rect 56205 4930 56245 4935
rect 56265 4965 56305 4970
rect 56265 4935 56270 4965
rect 56300 4935 56305 4965
rect 56265 4930 56305 4935
rect 56090 4900 56120 4930
rect 56090 4580 56095 4900
rect 56115 4580 56120 4900
rect 56090 4570 56120 4580
rect 56150 4900 56180 4910
rect 56150 4580 56155 4900
rect 56175 4580 56180 4900
rect 56150 4520 56180 4580
rect 56210 4900 56240 4930
rect 56210 4580 56215 4900
rect 56235 4580 56240 4900
rect 56210 4565 56240 4580
rect 56270 4900 56300 4930
rect 56270 4580 56275 4900
rect 56295 4580 56300 4900
rect 56555 4795 56595 4800
rect 56555 4765 56560 4795
rect 56590 4765 56595 4795
rect 56555 4760 56595 4765
rect 56615 4795 56655 4800
rect 56615 4765 56620 4795
rect 56650 4765 56655 4795
rect 56615 4760 56655 4765
rect 56270 4570 56300 4580
rect 56560 4730 56590 4760
rect 56560 4580 56565 4730
rect 56585 4580 56590 4730
rect 56560 4570 56590 4580
rect 56620 4730 56650 4760
rect 56620 4580 56625 4730
rect 56645 4580 56650 4730
rect 56620 4570 56650 4580
rect 56680 4730 56710 4985
rect 56890 4970 56910 6275
rect 57085 5020 57125 5025
rect 57085 4990 57090 5020
rect 57120 4990 57125 5020
rect 57085 4985 57125 4990
rect 57555 5020 57595 5025
rect 57555 4990 57560 5020
rect 57590 4990 57595 5020
rect 56880 4965 56920 4970
rect 56880 4935 56885 4965
rect 56915 4935 56920 4965
rect 56880 4930 56920 4935
rect 57025 4965 57065 4970
rect 57025 4935 57030 4965
rect 57060 4935 57065 4965
rect 57025 4930 57065 4935
rect 56890 4800 56910 4930
rect 57030 4900 57060 4930
rect 56735 4795 56775 4800
rect 56735 4765 56740 4795
rect 56770 4765 56775 4795
rect 56735 4760 56775 4765
rect 56880 4795 56920 4800
rect 56880 4765 56885 4795
rect 56915 4765 56920 4795
rect 56880 4760 56920 4765
rect 56680 4580 56685 4730
rect 56705 4580 56710 4730
rect 56680 4565 56710 4580
rect 56740 4730 56770 4760
rect 56740 4580 56745 4730
rect 56765 4580 56770 4730
rect 56740 4570 56770 4580
rect 56205 4560 56245 4565
rect 56205 4530 56210 4560
rect 56240 4530 56245 4560
rect 56205 4525 56245 4530
rect 56675 4560 56715 4565
rect 56675 4530 56680 4560
rect 56710 4530 56715 4560
rect 56675 4525 56715 4530
rect 56150 4515 56190 4520
rect 56150 4485 56155 4515
rect 56185 4485 56190 4515
rect 56150 4480 56190 4485
rect 56630 4515 56660 4520
rect 56630 4480 56660 4485
rect 56825 4515 56865 4520
rect 56825 4485 56830 4515
rect 56860 4485 56865 4515
rect 56825 4480 56865 4485
rect 55440 4275 55445 4305
rect 55475 4275 55485 4305
rect 55515 4275 55525 4305
rect 55555 4275 55560 4305
rect 55440 4270 55560 4275
rect 55750 4305 55910 4310
rect 55750 4275 55755 4305
rect 55785 4275 55795 4305
rect 55825 4275 55835 4305
rect 55865 4275 55875 4305
rect 55905 4275 55910 4305
rect 55750 4270 55910 4275
rect 55340 4210 55620 4215
rect 55340 4180 55345 4210
rect 55375 4180 55385 4210
rect 55415 4180 55425 4210
rect 55455 4180 55465 4210
rect 55495 4180 55505 4210
rect 55535 4180 55545 4210
rect 55575 4180 55585 4210
rect 55615 4180 55620 4210
rect 55340 4170 55620 4180
rect 55340 4140 55345 4170
rect 55375 4140 55385 4170
rect 55415 4140 55425 4170
rect 55455 4140 55465 4170
rect 55495 4140 55505 4170
rect 55535 4140 55545 4170
rect 55575 4140 55585 4170
rect 55615 4140 55620 4170
rect 55340 4130 55620 4140
rect 55340 4100 55345 4130
rect 55375 4100 55385 4130
rect 55415 4100 55425 4130
rect 55455 4100 55465 4130
rect 55495 4100 55505 4130
rect 55535 4100 55545 4130
rect 55575 4100 55585 4130
rect 55615 4100 55620 4130
rect 55340 4095 55620 4100
rect 55280 4045 55285 4075
rect 55315 4045 55320 4075
rect 55280 4040 55320 4045
rect 55225 3705 55230 4025
rect 55250 3705 55255 4025
rect 55225 3690 55255 3705
rect 55285 4025 55315 4040
rect 55285 3705 55290 4025
rect 55310 3705 55315 4025
rect 55285 3695 55315 3705
rect 55345 4025 55375 4095
rect 55400 4075 55440 4080
rect 55400 4045 55405 4075
rect 55435 4045 55440 4075
rect 55400 4040 55440 4045
rect 55345 3705 55350 4025
rect 55370 3705 55375 4025
rect 55345 3690 55375 3705
rect 55405 4025 55435 4040
rect 55405 3705 55410 4025
rect 55430 3705 55435 4025
rect 55405 3695 55435 3705
rect 55465 4025 55495 4095
rect 55520 4075 55560 4080
rect 55520 4045 55525 4075
rect 55555 4045 55560 4075
rect 55520 4040 55560 4045
rect 55465 3705 55470 4025
rect 55490 3705 55495 4025
rect 55465 3690 55495 3705
rect 55525 4025 55555 4040
rect 55525 3705 55530 4025
rect 55550 3705 55555 4025
rect 55525 3695 55555 3705
rect 55585 4025 55615 4095
rect 55640 4075 55680 4080
rect 55640 4045 55645 4075
rect 55675 4045 55680 4075
rect 55640 4040 55680 4045
rect 55585 3705 55590 4025
rect 55610 3705 55615 4025
rect 55585 3690 55615 3705
rect 55645 4025 55675 4040
rect 55645 3705 55650 4025
rect 55670 3705 55675 4025
rect 54925 3645 54930 3665
rect 54950 3645 54955 3665
rect 54980 3685 55020 3690
rect 54980 3655 54985 3685
rect 55015 3655 55020 3685
rect 54980 3650 55020 3655
rect 55100 3685 55140 3690
rect 55100 3655 55105 3685
rect 55135 3655 55140 3685
rect 55100 3650 55140 3655
rect 55220 3685 55260 3690
rect 55220 3655 55225 3685
rect 55255 3655 55260 3685
rect 55220 3650 55260 3655
rect 55340 3685 55380 3690
rect 55340 3655 55345 3685
rect 55375 3655 55380 3685
rect 55340 3650 55380 3655
rect 55460 3685 55500 3690
rect 55460 3655 55465 3685
rect 55495 3655 55500 3685
rect 55460 3650 55500 3655
rect 55580 3685 55620 3690
rect 55580 3655 55585 3685
rect 55615 3655 55620 3685
rect 55580 3650 55620 3655
rect 55645 3665 55675 3705
rect 54925 3635 54955 3645
rect 55645 3645 55650 3665
rect 55670 3645 55675 3665
rect 55645 3635 55675 3645
rect 55280 3560 55320 3565
rect 55280 3530 55285 3560
rect 55315 3530 55320 3560
rect 55280 3525 55320 3530
rect 55600 3515 55720 3520
rect 55600 3485 55605 3515
rect 55635 3485 55645 3515
rect 55675 3485 55685 3515
rect 55715 3485 55720 3515
rect 55600 3475 55720 3485
rect 55600 3445 55605 3475
rect 55635 3445 55645 3475
rect 55675 3445 55685 3475
rect 55715 3445 55720 3475
rect 55600 3435 55720 3445
rect 55600 3405 55605 3435
rect 55635 3405 55645 3435
rect 55675 3405 55685 3435
rect 55715 3405 55720 3435
rect 54605 3400 54645 3405
rect 54605 3370 54610 3400
rect 54640 3370 54645 3400
rect 54605 3365 54645 3370
rect 54820 3380 54860 3385
rect 54615 3325 54635 3365
rect 54820 3350 54825 3380
rect 54855 3350 54860 3380
rect 54820 3345 54860 3350
rect 54930 3380 54970 3385
rect 54930 3350 54935 3380
rect 54965 3350 54970 3380
rect 54930 3345 54970 3350
rect 55040 3380 55080 3385
rect 55040 3350 55045 3380
rect 55075 3350 55080 3380
rect 55040 3345 55080 3350
rect 55150 3380 55190 3385
rect 55150 3350 55155 3380
rect 55185 3350 55190 3380
rect 55150 3345 55190 3350
rect 55260 3380 55300 3385
rect 55260 3350 55265 3380
rect 55295 3350 55300 3380
rect 55260 3345 55300 3350
rect 55370 3380 55410 3385
rect 55370 3350 55375 3380
rect 55405 3350 55410 3380
rect 55370 3345 55410 3350
rect 55480 3380 55520 3385
rect 55480 3350 55485 3380
rect 55515 3350 55520 3380
rect 55480 3345 55520 3350
rect 54554 3315 54695 3325
rect 54554 3295 54560 3315
rect 54580 3295 54615 3315
rect 54635 3295 54670 3315
rect 54690 3295 54695 3315
rect 54554 3285 54695 3295
rect 54825 3310 54855 3345
rect 54825 3290 54830 3310
rect 54850 3290 54855 3310
rect 54825 3250 54855 3290
rect 54875 3300 54915 3305
rect 54875 3270 54880 3300
rect 54910 3270 54915 3300
rect 54875 3265 54915 3270
rect 54554 2710 54695 2720
rect 54554 2690 54560 2710
rect 54580 2690 54615 2710
rect 54635 2690 54670 2710
rect 54690 2690 54695 2710
rect 54554 2680 54695 2690
rect 54825 2680 54830 3250
rect 54850 2680 54855 3250
rect 54605 2625 54645 2680
rect 54825 2670 54855 2680
rect 54880 3250 54910 3265
rect 54880 2680 54885 3250
rect 54905 2680 54910 3250
rect 54880 2665 54910 2680
rect 54935 3250 54965 3345
rect 54985 3300 55025 3305
rect 54985 3270 54990 3300
rect 55020 3270 55025 3300
rect 54985 3265 55025 3270
rect 54935 2680 54940 3250
rect 54960 2680 54965 3250
rect 54935 2670 54965 2680
rect 54990 3250 55020 3265
rect 54990 2680 54995 3250
rect 55015 2680 55020 3250
rect 54990 2665 55020 2680
rect 55045 3250 55075 3345
rect 55095 3300 55135 3305
rect 55095 3270 55100 3300
rect 55130 3270 55135 3300
rect 55095 3265 55135 3270
rect 55045 2680 55050 3250
rect 55070 2680 55075 3250
rect 55045 2670 55075 2680
rect 55100 3250 55130 3265
rect 55100 2680 55105 3250
rect 55125 2680 55130 3250
rect 55100 2665 55130 2680
rect 55155 3250 55185 3345
rect 55205 3300 55245 3305
rect 55205 3270 55210 3300
rect 55240 3270 55245 3300
rect 55205 3265 55245 3270
rect 55155 2680 55160 3250
rect 55180 2680 55185 3250
rect 55155 2670 55185 2680
rect 55210 3250 55240 3265
rect 55210 2680 55215 3250
rect 55235 2680 55240 3250
rect 55210 2665 55240 2680
rect 55265 3250 55295 3345
rect 55315 3300 55355 3305
rect 55315 3270 55320 3300
rect 55350 3270 55355 3300
rect 55315 3265 55355 3270
rect 55265 2680 55270 3250
rect 55290 2680 55295 3250
rect 55265 2670 55295 2680
rect 55320 3250 55350 3265
rect 55320 2680 55325 3250
rect 55345 2680 55350 3250
rect 55320 2665 55350 2680
rect 55375 3250 55405 3345
rect 55485 3310 55515 3345
rect 55425 3300 55465 3305
rect 55425 3270 55430 3300
rect 55460 3270 55465 3300
rect 55425 3265 55465 3270
rect 55485 3290 55490 3310
rect 55510 3290 55515 3310
rect 55375 2680 55380 3250
rect 55400 2680 55405 3250
rect 55375 2670 55405 2680
rect 55430 3250 55460 3265
rect 55430 2680 55435 3250
rect 55455 2680 55460 3250
rect 55430 2665 55460 2680
rect 55485 3250 55515 3290
rect 55485 2680 55490 3250
rect 55510 2680 55515 3250
rect 55485 2670 55515 2680
rect 54875 2660 54915 2665
rect 54875 2630 54880 2660
rect 54910 2630 54915 2660
rect 54565 2580 54685 2625
rect 54565 2550 54570 2580
rect 54600 2550 54610 2580
rect 54640 2550 54650 2580
rect 54680 2550 54685 2580
rect 54565 2540 54685 2550
rect 54565 2510 54570 2540
rect 54600 2510 54610 2540
rect 54640 2510 54650 2540
rect 54680 2510 54685 2540
rect 54565 2500 54685 2510
rect 54565 2470 54570 2500
rect 54600 2470 54610 2500
rect 54640 2470 54650 2500
rect 54680 2470 54685 2500
rect 54565 2465 54685 2470
rect 54875 2435 54915 2630
rect 54985 2660 55025 2665
rect 54985 2630 54990 2660
rect 55020 2630 55025 2660
rect 54985 2435 55025 2630
rect 55095 2660 55135 2665
rect 55095 2630 55100 2660
rect 55130 2630 55135 2660
rect 55095 2435 55135 2630
rect 55205 2660 55245 2665
rect 55205 2630 55210 2660
rect 55240 2630 55245 2660
rect 55150 2580 55190 2585
rect 55150 2550 55155 2580
rect 55185 2550 55190 2580
rect 55150 2540 55190 2550
rect 55150 2510 55155 2540
rect 55185 2510 55190 2540
rect 55150 2500 55190 2510
rect 55150 2470 55155 2500
rect 55185 2470 55190 2500
rect 55150 2465 55190 2470
rect 55205 2435 55245 2630
rect 55315 2660 55355 2665
rect 55315 2630 55320 2660
rect 55350 2630 55355 2660
rect 55315 2435 55355 2630
rect 55425 2660 55465 2665
rect 55425 2630 55430 2660
rect 55460 2630 55465 2660
rect 55425 2435 55465 2630
rect 54185 2430 54435 2435
rect 54185 2400 54190 2430
rect 54220 2400 54230 2430
rect 54260 2400 54275 2430
rect 54305 2400 54315 2430
rect 54345 2400 54360 2430
rect 54390 2400 54400 2430
rect 54430 2400 54435 2430
rect 54185 2390 54435 2400
rect 54185 2360 54190 2390
rect 54220 2360 54230 2390
rect 54260 2360 54275 2390
rect 54305 2360 54315 2390
rect 54345 2360 54360 2390
rect 54390 2360 54400 2390
rect 54430 2360 54435 2390
rect 54185 2350 54435 2360
rect 54185 2320 54190 2350
rect 54220 2320 54230 2350
rect 54260 2320 54275 2350
rect 54305 2320 54315 2350
rect 54345 2320 54360 2350
rect 54390 2320 54400 2350
rect 54430 2320 54435 2350
rect 54115 2245 54155 2250
rect 54115 2215 54120 2245
rect 54150 2215 54155 2245
rect 54115 2210 54155 2215
rect 54125 50 54145 2210
rect 54185 1710 54435 2320
rect 54875 2430 55465 2435
rect 54875 2400 54880 2430
rect 54910 2400 54935 2430
rect 54965 2400 54990 2430
rect 55020 2400 55045 2430
rect 55075 2400 55100 2430
rect 55130 2400 55155 2430
rect 55185 2400 55210 2430
rect 55240 2400 55265 2430
rect 55295 2400 55320 2430
rect 55350 2400 55375 2430
rect 55405 2400 55430 2430
rect 55460 2400 55465 2430
rect 54875 2390 55465 2400
rect 54875 2360 54880 2390
rect 54910 2360 54935 2390
rect 54965 2360 54990 2390
rect 55020 2360 55045 2390
rect 55075 2360 55100 2390
rect 55130 2360 55155 2390
rect 55185 2360 55210 2390
rect 55240 2360 55265 2390
rect 55295 2360 55320 2390
rect 55350 2360 55375 2390
rect 55405 2360 55430 2390
rect 55460 2360 55465 2390
rect 54875 2350 55465 2360
rect 54875 2320 54880 2350
rect 54910 2320 54935 2350
rect 54965 2320 54990 2350
rect 55020 2320 55045 2350
rect 55075 2320 55100 2350
rect 55130 2320 55155 2350
rect 55185 2320 55210 2350
rect 55240 2320 55265 2350
rect 55295 2320 55320 2350
rect 55350 2320 55375 2350
rect 55405 2320 55430 2350
rect 55460 2320 55465 2350
rect 54875 2315 55465 2320
rect 55600 2580 55720 3405
rect 55760 3400 55780 4270
rect 56005 4210 56765 4215
rect 56005 4180 56010 4210
rect 56040 4180 56050 4210
rect 56080 4180 56090 4210
rect 56120 4180 56130 4210
rect 56160 4180 56170 4210
rect 56200 4180 56210 4210
rect 56240 4180 56250 4210
rect 56280 4180 56290 4210
rect 56320 4180 56330 4210
rect 56360 4180 56370 4210
rect 56400 4180 56410 4210
rect 56440 4180 56450 4210
rect 56480 4180 56490 4210
rect 56520 4180 56530 4210
rect 56560 4180 56570 4210
rect 56600 4180 56610 4210
rect 56640 4180 56650 4210
rect 56680 4180 56690 4210
rect 56720 4180 56730 4210
rect 56760 4180 56765 4210
rect 56005 4170 56765 4180
rect 56005 4140 56010 4170
rect 56040 4140 56050 4170
rect 56080 4140 56090 4170
rect 56120 4140 56130 4170
rect 56160 4140 56170 4170
rect 56200 4140 56210 4170
rect 56240 4140 56250 4170
rect 56280 4140 56290 4170
rect 56320 4140 56330 4170
rect 56360 4140 56370 4170
rect 56400 4140 56410 4170
rect 56440 4140 56450 4170
rect 56480 4140 56490 4170
rect 56520 4140 56530 4170
rect 56560 4140 56570 4170
rect 56600 4140 56610 4170
rect 56640 4140 56650 4170
rect 56680 4140 56690 4170
rect 56720 4140 56730 4170
rect 56760 4140 56765 4170
rect 56005 4130 56765 4140
rect 56005 4100 56010 4130
rect 56040 4100 56050 4130
rect 56080 4100 56090 4130
rect 56120 4100 56130 4130
rect 56160 4100 56170 4130
rect 56200 4100 56210 4130
rect 56240 4100 56250 4130
rect 56280 4100 56290 4130
rect 56320 4100 56330 4130
rect 56360 4100 56370 4130
rect 56400 4100 56410 4130
rect 56440 4100 56450 4130
rect 56480 4100 56490 4130
rect 56520 4100 56530 4130
rect 56560 4100 56570 4130
rect 56600 4100 56610 4130
rect 56640 4100 56650 4130
rect 56680 4100 56690 4130
rect 56720 4100 56730 4130
rect 56760 4100 56765 4130
rect 56005 4095 56765 4100
rect 56010 4025 56040 4095
rect 56065 4075 56105 4080
rect 56065 4045 56070 4075
rect 56100 4045 56105 4075
rect 56065 4040 56105 4045
rect 56010 3705 56015 4025
rect 56035 3705 56040 4025
rect 56010 3665 56040 3705
rect 56070 4025 56100 4040
rect 56070 3705 56075 4025
rect 56095 3705 56100 4025
rect 56070 3690 56100 3705
rect 56130 4025 56160 4095
rect 56185 4075 56225 4080
rect 56185 4045 56190 4075
rect 56220 4045 56225 4075
rect 56185 4040 56225 4045
rect 56130 3705 56135 4025
rect 56155 3705 56160 4025
rect 56130 3695 56160 3705
rect 56190 4025 56220 4040
rect 56190 3705 56195 4025
rect 56215 3705 56220 4025
rect 56190 3690 56220 3705
rect 56250 4025 56280 4095
rect 56305 4075 56345 4080
rect 56305 4045 56310 4075
rect 56340 4045 56345 4075
rect 56305 4040 56345 4045
rect 56250 3705 56255 4025
rect 56275 3705 56280 4025
rect 56250 3695 56280 3705
rect 56310 4025 56340 4040
rect 56310 3705 56315 4025
rect 56335 3705 56340 4025
rect 56310 3690 56340 3705
rect 56370 4025 56400 4095
rect 56425 4075 56465 4080
rect 56425 4045 56430 4075
rect 56460 4045 56465 4075
rect 56425 4040 56465 4045
rect 56370 3705 56375 4025
rect 56395 3705 56400 4025
rect 56370 3695 56400 3705
rect 56430 4025 56460 4040
rect 56430 3705 56435 4025
rect 56455 3705 56460 4025
rect 56430 3690 56460 3705
rect 56490 4025 56520 4095
rect 56545 4075 56585 4080
rect 56545 4045 56550 4075
rect 56580 4045 56585 4075
rect 56545 4040 56585 4045
rect 56490 3705 56495 4025
rect 56515 3705 56520 4025
rect 56490 3695 56520 3705
rect 56550 4025 56580 4040
rect 56550 3705 56555 4025
rect 56575 3705 56580 4025
rect 56550 3690 56580 3705
rect 56610 4025 56640 4095
rect 56665 4075 56705 4080
rect 56665 4045 56670 4075
rect 56700 4045 56705 4075
rect 56665 4040 56705 4045
rect 56610 3705 56615 4025
rect 56635 3705 56640 4025
rect 56610 3695 56640 3705
rect 56670 4025 56700 4040
rect 56670 3705 56675 4025
rect 56695 3705 56700 4025
rect 56670 3690 56700 3705
rect 56730 4025 56760 4095
rect 56730 3705 56735 4025
rect 56755 3705 56760 4025
rect 56010 3645 56015 3665
rect 56035 3645 56040 3665
rect 56010 3635 56040 3645
rect 56065 3685 56105 3690
rect 56065 3655 56070 3685
rect 56100 3655 56105 3685
rect 56065 3520 56105 3655
rect 56185 3685 56225 3690
rect 56185 3655 56190 3685
rect 56220 3655 56225 3685
rect 56185 3520 56225 3655
rect 56305 3685 56345 3690
rect 56305 3655 56310 3685
rect 56340 3655 56345 3685
rect 56305 3520 56345 3655
rect 56425 3685 56465 3690
rect 56425 3655 56430 3685
rect 56460 3655 56465 3685
rect 56365 3605 56405 3610
rect 56365 3575 56370 3605
rect 56400 3575 56405 3605
rect 56365 3570 56405 3575
rect 56425 3520 56465 3655
rect 56545 3685 56585 3690
rect 56545 3655 56550 3685
rect 56580 3655 56585 3685
rect 56545 3520 56585 3655
rect 56665 3685 56705 3690
rect 56665 3655 56670 3685
rect 56700 3655 56705 3685
rect 56665 3520 56705 3655
rect 56730 3665 56760 3705
rect 56730 3645 56735 3665
rect 56755 3645 56760 3665
rect 56730 3635 56760 3645
rect 56845 3610 56865 4480
rect 56890 4310 56910 4760
rect 57030 4580 57035 4900
rect 57055 4580 57060 4900
rect 57030 4570 57060 4580
rect 57090 4900 57120 4985
rect 57145 4965 57185 4970
rect 57145 4935 57150 4965
rect 57180 4935 57185 4965
rect 57145 4930 57185 4935
rect 57205 4965 57245 4970
rect 57205 4935 57210 4965
rect 57240 4935 57245 4965
rect 57205 4930 57245 4935
rect 57495 4965 57535 4970
rect 57495 4935 57500 4965
rect 57530 4935 57535 4965
rect 57495 4930 57535 4935
rect 57555 4965 57595 4990
rect 57555 4935 57560 4965
rect 57590 4935 57595 4965
rect 57555 4930 57595 4935
rect 57675 4965 57715 4970
rect 57675 4935 57680 4965
rect 57710 4935 57715 4965
rect 57675 4930 57715 4935
rect 57090 4580 57095 4900
rect 57115 4580 57120 4900
rect 57090 4565 57120 4580
rect 57150 4900 57180 4930
rect 57150 4580 57155 4900
rect 57175 4580 57180 4900
rect 57150 4570 57180 4580
rect 57210 4900 57240 4930
rect 57210 4580 57215 4900
rect 57235 4580 57240 4900
rect 57210 4570 57240 4580
rect 57500 4900 57530 4930
rect 57500 4580 57505 4900
rect 57525 4580 57530 4900
rect 57500 4570 57530 4580
rect 57560 4900 57590 4930
rect 57560 4580 57565 4900
rect 57585 4580 57590 4900
rect 57560 4565 57590 4580
rect 57620 4900 57650 4910
rect 57620 4580 57625 4900
rect 57645 4580 57650 4900
rect 57085 4560 57125 4565
rect 57085 4530 57090 4560
rect 57120 4530 57125 4560
rect 57085 4525 57125 4530
rect 57555 4560 57595 4565
rect 57555 4530 57560 4560
rect 57590 4530 57595 4560
rect 57555 4525 57595 4530
rect 57140 4510 57170 4520
rect 57140 4490 57145 4510
rect 57165 4490 57170 4510
rect 56935 4460 56975 4465
rect 56935 4430 56940 4460
rect 56970 4430 56975 4460
rect 57140 4455 57170 4490
rect 57576 4505 57606 4510
rect 57576 4470 57606 4475
rect 57620 4455 57650 4580
rect 57680 4900 57710 4930
rect 57680 4580 57685 4900
rect 57705 4580 57710 4900
rect 57680 4570 57710 4580
rect 56935 4425 56975 4430
rect 57135 4450 57175 4455
rect 56880 4305 56920 4310
rect 56880 4275 56885 4305
rect 56915 4275 56920 4305
rect 56880 4270 56920 4275
rect 56835 3605 56875 3610
rect 56835 3575 56840 3605
rect 56870 3575 56875 3605
rect 56835 3570 56875 3575
rect 56935 3565 56955 4425
rect 57135 4420 57140 4450
rect 57170 4420 57175 4450
rect 57135 4415 57175 4420
rect 57615 4450 57655 4455
rect 57615 4420 57620 4450
rect 57650 4420 57655 4450
rect 57615 4415 57655 4420
rect 57890 4310 58010 6275
rect 57890 4305 58050 4310
rect 57890 4275 57895 4305
rect 57925 4275 57935 4305
rect 57965 4275 57975 4305
rect 58005 4275 58015 4305
rect 58045 4275 58050 4305
rect 57890 4270 58050 4275
rect 58240 4305 58360 6275
rect 58240 4275 58245 4305
rect 58275 4275 58285 4305
rect 58315 4275 58325 4305
rect 58355 4275 58360 4305
rect 58240 4270 58360 4275
rect 58480 4305 58520 4310
rect 58480 4275 58485 4305
rect 58515 4275 58520 4305
rect 57035 4210 57795 4215
rect 57035 4180 57040 4210
rect 57070 4180 57080 4210
rect 57110 4180 57120 4210
rect 57150 4180 57160 4210
rect 57190 4180 57200 4210
rect 57230 4180 57240 4210
rect 57270 4180 57280 4210
rect 57310 4180 57320 4210
rect 57350 4180 57360 4210
rect 57390 4180 57400 4210
rect 57430 4180 57440 4210
rect 57470 4180 57480 4210
rect 57510 4180 57520 4210
rect 57550 4180 57560 4210
rect 57590 4180 57600 4210
rect 57630 4180 57640 4210
rect 57670 4180 57680 4210
rect 57710 4180 57720 4210
rect 57750 4180 57760 4210
rect 57790 4180 57795 4210
rect 57035 4170 57795 4180
rect 57035 4140 57040 4170
rect 57070 4140 57080 4170
rect 57110 4140 57120 4170
rect 57150 4140 57160 4170
rect 57190 4140 57200 4170
rect 57230 4140 57240 4170
rect 57270 4140 57280 4170
rect 57310 4140 57320 4170
rect 57350 4140 57360 4170
rect 57390 4140 57400 4170
rect 57430 4140 57440 4170
rect 57470 4140 57480 4170
rect 57510 4140 57520 4170
rect 57550 4140 57560 4170
rect 57590 4140 57600 4170
rect 57630 4140 57640 4170
rect 57670 4140 57680 4170
rect 57710 4140 57720 4170
rect 57750 4140 57760 4170
rect 57790 4140 57795 4170
rect 57035 4130 57795 4140
rect 57035 4100 57040 4130
rect 57070 4100 57080 4130
rect 57110 4100 57120 4130
rect 57150 4100 57160 4130
rect 57190 4100 57200 4130
rect 57230 4100 57240 4130
rect 57270 4100 57280 4130
rect 57310 4100 57320 4130
rect 57350 4100 57360 4130
rect 57390 4100 57400 4130
rect 57430 4100 57440 4130
rect 57470 4100 57480 4130
rect 57510 4100 57520 4130
rect 57550 4100 57560 4130
rect 57590 4100 57600 4130
rect 57630 4100 57640 4130
rect 57670 4100 57680 4130
rect 57710 4100 57720 4130
rect 57750 4100 57760 4130
rect 57790 4100 57795 4130
rect 57035 4095 57795 4100
rect 57040 4025 57070 4095
rect 57095 4075 57135 4080
rect 57095 4045 57100 4075
rect 57130 4045 57135 4075
rect 57095 4040 57135 4045
rect 57040 3705 57045 4025
rect 57065 3705 57070 4025
rect 57040 3665 57070 3705
rect 57100 4025 57130 4040
rect 57100 3705 57105 4025
rect 57125 3705 57130 4025
rect 57100 3690 57130 3705
rect 57160 4025 57190 4095
rect 57215 4075 57255 4080
rect 57215 4045 57220 4075
rect 57250 4045 57255 4075
rect 57215 4040 57255 4045
rect 57160 3705 57165 4025
rect 57185 3705 57190 4025
rect 57160 3695 57190 3705
rect 57220 4025 57250 4040
rect 57220 3705 57225 4025
rect 57245 3705 57250 4025
rect 57220 3690 57250 3705
rect 57280 4025 57310 4095
rect 57335 4075 57375 4080
rect 57335 4045 57340 4075
rect 57370 4045 57375 4075
rect 57335 4040 57375 4045
rect 57280 3705 57285 4025
rect 57305 3705 57310 4025
rect 57280 3695 57310 3705
rect 57340 4025 57370 4040
rect 57340 3705 57345 4025
rect 57365 3705 57370 4025
rect 57340 3690 57370 3705
rect 57400 4025 57430 4095
rect 57455 4075 57495 4080
rect 57455 4045 57460 4075
rect 57490 4045 57495 4075
rect 57455 4040 57495 4045
rect 57400 3705 57405 4025
rect 57425 3705 57430 4025
rect 57400 3695 57430 3705
rect 57460 4025 57490 4040
rect 57460 3705 57465 4025
rect 57485 3705 57490 4025
rect 57460 3690 57490 3705
rect 57520 4025 57550 4095
rect 57575 4075 57615 4080
rect 57575 4045 57580 4075
rect 57610 4045 57615 4075
rect 57575 4040 57615 4045
rect 57520 3705 57525 4025
rect 57545 3705 57550 4025
rect 57520 3695 57550 3705
rect 57580 4025 57610 4040
rect 57580 3705 57585 4025
rect 57605 3705 57610 4025
rect 57580 3690 57610 3705
rect 57640 4025 57670 4095
rect 57695 4075 57735 4080
rect 57695 4045 57700 4075
rect 57730 4045 57735 4075
rect 57695 4040 57735 4045
rect 57640 3705 57645 4025
rect 57665 3705 57670 4025
rect 57640 3695 57670 3705
rect 57700 4025 57730 4040
rect 57700 3705 57705 4025
rect 57725 3705 57730 4025
rect 57700 3690 57730 3705
rect 57760 4025 57790 4095
rect 57760 3705 57765 4025
rect 57785 3705 57790 4025
rect 57040 3645 57045 3665
rect 57065 3645 57070 3665
rect 57040 3635 57070 3645
rect 57095 3685 57135 3690
rect 57095 3655 57100 3685
rect 57130 3655 57135 3685
rect 56925 3560 56965 3565
rect 56925 3530 56930 3560
rect 56960 3530 56965 3560
rect 56925 3525 56965 3530
rect 56065 3515 56705 3520
rect 56065 3485 56070 3515
rect 56100 3485 56110 3515
rect 56140 3485 56150 3515
rect 56180 3485 56190 3515
rect 56220 3485 56230 3515
rect 56260 3485 56270 3515
rect 56300 3485 56310 3515
rect 56340 3485 56350 3515
rect 56380 3485 56390 3515
rect 56420 3485 56430 3515
rect 56460 3485 56470 3515
rect 56500 3485 56510 3515
rect 56540 3485 56550 3515
rect 56580 3485 56590 3515
rect 56620 3485 56630 3515
rect 56660 3485 56670 3515
rect 56700 3485 56705 3515
rect 56065 3475 56705 3485
rect 56065 3445 56070 3475
rect 56100 3445 56110 3475
rect 56140 3445 56150 3475
rect 56180 3445 56190 3475
rect 56220 3445 56230 3475
rect 56260 3445 56270 3475
rect 56300 3445 56310 3475
rect 56340 3445 56350 3475
rect 56380 3445 56390 3475
rect 56420 3445 56430 3475
rect 56460 3445 56470 3475
rect 56500 3445 56510 3475
rect 56540 3445 56550 3475
rect 56580 3445 56590 3475
rect 56620 3445 56630 3475
rect 56660 3445 56670 3475
rect 56700 3445 56705 3475
rect 56065 3435 56705 3445
rect 56065 3405 56070 3435
rect 56100 3405 56110 3435
rect 56140 3405 56150 3435
rect 56180 3405 56190 3435
rect 56220 3405 56230 3435
rect 56260 3405 56270 3435
rect 56300 3405 56310 3435
rect 56340 3405 56350 3435
rect 56380 3405 56390 3435
rect 56420 3405 56430 3435
rect 56460 3405 56470 3435
rect 56500 3405 56510 3435
rect 56540 3405 56550 3435
rect 56580 3405 56590 3435
rect 56620 3405 56630 3435
rect 56660 3405 56670 3435
rect 56700 3405 56705 3435
rect 56065 3400 56705 3405
rect 57095 3520 57135 3655
rect 57215 3685 57255 3690
rect 57215 3655 57220 3685
rect 57250 3655 57255 3685
rect 57215 3520 57255 3655
rect 57335 3685 57375 3690
rect 57335 3655 57340 3685
rect 57370 3655 57375 3685
rect 57335 3520 57375 3655
rect 57455 3685 57495 3690
rect 57455 3655 57460 3685
rect 57490 3655 57495 3685
rect 57395 3605 57435 3610
rect 57395 3575 57400 3605
rect 57430 3575 57435 3605
rect 57395 3570 57435 3575
rect 57455 3520 57495 3655
rect 57575 3685 57615 3690
rect 57575 3655 57580 3685
rect 57610 3655 57615 3685
rect 57575 3520 57615 3655
rect 57695 3685 57735 3690
rect 57695 3655 57700 3685
rect 57730 3655 57735 3685
rect 57695 3520 57735 3655
rect 57760 3665 57790 3705
rect 57760 3645 57765 3665
rect 57785 3645 57790 3665
rect 57760 3635 57790 3645
rect 57095 3515 57735 3520
rect 57095 3485 57100 3515
rect 57130 3485 57140 3515
rect 57170 3485 57180 3515
rect 57210 3485 57220 3515
rect 57250 3485 57260 3515
rect 57290 3485 57300 3515
rect 57330 3485 57340 3515
rect 57370 3485 57380 3515
rect 57410 3485 57420 3515
rect 57450 3485 57460 3515
rect 57490 3485 57500 3515
rect 57530 3485 57540 3515
rect 57570 3485 57580 3515
rect 57610 3485 57620 3515
rect 57650 3485 57660 3515
rect 57690 3485 57700 3515
rect 57730 3485 57735 3515
rect 57095 3475 57735 3485
rect 57095 3445 57100 3475
rect 57130 3445 57140 3475
rect 57170 3445 57180 3475
rect 57210 3445 57220 3475
rect 57250 3445 57260 3475
rect 57290 3445 57300 3475
rect 57330 3445 57340 3475
rect 57370 3445 57380 3475
rect 57410 3445 57420 3475
rect 57450 3445 57460 3475
rect 57490 3445 57500 3475
rect 57530 3445 57540 3475
rect 57570 3445 57580 3475
rect 57610 3445 57620 3475
rect 57650 3445 57660 3475
rect 57690 3445 57700 3475
rect 57730 3445 57735 3475
rect 57095 3435 57735 3445
rect 57095 3405 57100 3435
rect 57130 3405 57140 3435
rect 57170 3405 57180 3435
rect 57210 3405 57220 3435
rect 57250 3405 57260 3435
rect 57290 3405 57300 3435
rect 57330 3405 57340 3435
rect 57370 3405 57380 3435
rect 57410 3405 57420 3435
rect 57450 3405 57460 3435
rect 57490 3405 57500 3435
rect 57530 3405 57540 3435
rect 57570 3405 57580 3435
rect 57610 3405 57620 3435
rect 57650 3405 57660 3435
rect 57690 3405 57700 3435
rect 57730 3405 57735 3435
rect 57095 3400 57735 3405
rect 55765 3385 55785 3400
rect 58020 3385 58040 4270
rect 58180 4210 58460 4215
rect 58180 4180 58185 4210
rect 58215 4180 58225 4210
rect 58255 4180 58265 4210
rect 58295 4180 58305 4210
rect 58335 4180 58345 4210
rect 58375 4180 58385 4210
rect 58415 4180 58425 4210
rect 58455 4180 58460 4210
rect 58180 4170 58460 4180
rect 58180 4140 58185 4170
rect 58215 4140 58225 4170
rect 58255 4140 58265 4170
rect 58295 4140 58305 4170
rect 58335 4140 58345 4170
rect 58375 4140 58385 4170
rect 58415 4140 58425 4170
rect 58455 4140 58460 4170
rect 58180 4130 58460 4140
rect 58180 4100 58185 4130
rect 58215 4100 58225 4130
rect 58255 4100 58265 4130
rect 58295 4100 58305 4130
rect 58335 4100 58345 4130
rect 58375 4100 58385 4130
rect 58415 4100 58425 4130
rect 58455 4100 58460 4130
rect 58180 4095 58460 4100
rect 58120 4075 58160 4080
rect 58120 4045 58125 4075
rect 58155 4045 58160 4075
rect 58120 4040 58160 4045
rect 58125 4025 58155 4040
rect 58125 3705 58130 4025
rect 58150 3705 58155 4025
rect 58125 3665 58155 3705
rect 58185 4025 58215 4095
rect 58240 4075 58280 4080
rect 58240 4045 58245 4075
rect 58275 4045 58280 4075
rect 58240 4040 58280 4045
rect 58185 3705 58190 4025
rect 58210 3705 58215 4025
rect 58185 3690 58215 3705
rect 58245 4025 58275 4040
rect 58245 3705 58250 4025
rect 58270 3705 58275 4025
rect 58245 3695 58275 3705
rect 58305 4025 58335 4095
rect 58360 4075 58400 4080
rect 58360 4045 58365 4075
rect 58395 4045 58400 4075
rect 58360 4040 58400 4045
rect 58305 3705 58310 4025
rect 58330 3705 58335 4025
rect 58305 3690 58335 3705
rect 58365 4025 58395 4040
rect 58365 3705 58370 4025
rect 58390 3705 58395 4025
rect 58365 3695 58395 3705
rect 58425 4025 58455 4095
rect 58480 4075 58520 4275
rect 58590 4305 58710 6275
rect 58590 4275 58595 4305
rect 58625 4275 58635 4305
rect 58665 4275 58675 4305
rect 58705 4275 58710 4305
rect 58590 4270 58710 4275
rect 58940 4305 59060 6275
rect 58940 4275 58945 4305
rect 58975 4275 58985 4305
rect 59015 4275 59025 4305
rect 59055 4275 59060 4305
rect 58940 4270 59060 4275
rect 59290 4305 59410 6275
rect 59290 4275 59295 4305
rect 59325 4275 59335 4305
rect 59365 4275 59375 4305
rect 59405 4275 59410 4305
rect 59290 4270 59410 4275
rect 59640 4305 59760 6275
rect 59640 4275 59645 4305
rect 59675 4275 59685 4305
rect 59715 4275 59725 4305
rect 59755 4275 59760 4305
rect 59640 4270 59760 4275
rect 59990 4305 60110 6275
rect 59990 4275 59995 4305
rect 60025 4275 60035 4305
rect 60065 4275 60075 4305
rect 60105 4275 60110 4305
rect 59990 4270 60110 4275
rect 60340 4305 60460 6275
rect 60340 4275 60345 4305
rect 60375 4275 60385 4305
rect 60415 4275 60425 4305
rect 60455 4275 60460 4305
rect 60340 4270 60460 4275
rect 60690 4305 60810 6275
rect 60690 4275 60695 4305
rect 60725 4275 60735 4305
rect 60765 4275 60775 4305
rect 60805 4275 60810 4305
rect 60690 4270 60810 4275
rect 61040 4305 61160 6275
rect 61040 4275 61045 4305
rect 61075 4275 61085 4305
rect 61115 4275 61125 4305
rect 61155 4275 61160 4305
rect 61040 4270 61160 4275
rect 58540 4210 58820 4215
rect 58540 4180 58545 4210
rect 58575 4180 58585 4210
rect 58615 4180 58625 4210
rect 58655 4180 58665 4210
rect 58695 4180 58705 4210
rect 58735 4180 58745 4210
rect 58775 4180 58785 4210
rect 58815 4180 58820 4210
rect 58540 4170 58820 4180
rect 58540 4140 58545 4170
rect 58575 4140 58585 4170
rect 58615 4140 58625 4170
rect 58655 4140 58665 4170
rect 58695 4140 58705 4170
rect 58735 4140 58745 4170
rect 58775 4140 58785 4170
rect 58815 4140 58820 4170
rect 58540 4130 58820 4140
rect 58540 4100 58545 4130
rect 58575 4100 58585 4130
rect 58615 4100 58625 4130
rect 58655 4100 58665 4130
rect 58695 4100 58705 4130
rect 58735 4100 58745 4130
rect 58775 4100 58785 4130
rect 58815 4100 58820 4130
rect 58540 4095 58820 4100
rect 58480 4045 58485 4075
rect 58515 4045 58520 4075
rect 58480 4040 58520 4045
rect 58425 3705 58430 4025
rect 58450 3705 58455 4025
rect 58425 3690 58455 3705
rect 58485 4025 58515 4040
rect 58485 3705 58490 4025
rect 58510 3705 58515 4025
rect 58485 3695 58515 3705
rect 58545 4025 58575 4095
rect 58600 4075 58640 4080
rect 58600 4045 58605 4075
rect 58635 4045 58640 4075
rect 58600 4040 58640 4045
rect 58545 3705 58550 4025
rect 58570 3705 58575 4025
rect 58545 3690 58575 3705
rect 58605 4025 58635 4040
rect 58605 3705 58610 4025
rect 58630 3705 58635 4025
rect 58605 3695 58635 3705
rect 58665 4025 58695 4095
rect 58720 4075 58760 4080
rect 58720 4045 58725 4075
rect 58755 4045 58760 4075
rect 58720 4040 58760 4045
rect 58665 3705 58670 4025
rect 58690 3705 58695 4025
rect 58665 3690 58695 3705
rect 58725 4025 58755 4040
rect 58725 3705 58730 4025
rect 58750 3705 58755 4025
rect 58725 3695 58755 3705
rect 58785 4025 58815 4095
rect 58840 4075 58880 4080
rect 58840 4045 58845 4075
rect 58875 4045 58880 4075
rect 58840 4040 58880 4045
rect 58785 3705 58790 4025
rect 58810 3705 58815 4025
rect 58785 3690 58815 3705
rect 58845 4025 58875 4040
rect 58845 3705 58850 4025
rect 58870 3705 58875 4025
rect 58125 3645 58130 3665
rect 58150 3645 58155 3665
rect 58180 3685 58220 3690
rect 58180 3655 58185 3685
rect 58215 3655 58220 3685
rect 58180 3650 58220 3655
rect 58300 3685 58340 3690
rect 58300 3655 58305 3685
rect 58335 3655 58340 3685
rect 58300 3650 58340 3655
rect 58420 3685 58460 3690
rect 58420 3655 58425 3685
rect 58455 3655 58460 3685
rect 58420 3650 58460 3655
rect 58540 3685 58580 3690
rect 58540 3655 58545 3685
rect 58575 3655 58580 3685
rect 58540 3650 58580 3655
rect 58660 3685 58700 3690
rect 58660 3655 58665 3685
rect 58695 3655 58700 3685
rect 58660 3650 58700 3655
rect 58780 3685 58820 3690
rect 58780 3655 58785 3685
rect 58815 3655 58820 3685
rect 58780 3650 58820 3655
rect 58845 3665 58875 3705
rect 58125 3635 58155 3645
rect 58845 3645 58850 3665
rect 58870 3645 58875 3665
rect 58845 3635 58875 3645
rect 58480 3560 58520 3565
rect 58480 3530 58485 3560
rect 58515 3530 58520 3560
rect 58480 3525 58520 3530
rect 58080 3515 58200 3520
rect 58080 3485 58085 3515
rect 58115 3485 58125 3515
rect 58155 3485 58165 3515
rect 58195 3485 58200 3515
rect 58080 3475 58200 3485
rect 58080 3445 58085 3475
rect 58115 3445 58125 3475
rect 58155 3445 58165 3475
rect 58195 3445 58200 3475
rect 58080 3435 58200 3445
rect 58080 3405 58085 3435
rect 58115 3405 58125 3435
rect 58155 3405 58165 3435
rect 58195 3405 58200 3435
rect 55750 3380 55790 3385
rect 55750 3350 55755 3380
rect 55785 3350 55790 3380
rect 55750 3345 55790 3350
rect 56275 3380 56315 3385
rect 56275 3350 56280 3380
rect 56310 3350 56315 3380
rect 56275 3345 56315 3350
rect 56385 3380 56425 3385
rect 56385 3350 56390 3380
rect 56420 3350 56425 3380
rect 56385 3345 56425 3350
rect 56495 3380 56535 3385
rect 56495 3350 56500 3380
rect 56530 3350 56535 3380
rect 56495 3345 56535 3350
rect 56605 3380 56645 3385
rect 56605 3350 56610 3380
rect 56640 3350 56645 3380
rect 56605 3345 56645 3350
rect 56715 3380 56755 3385
rect 56715 3350 56720 3380
rect 56750 3350 56755 3380
rect 56715 3345 56755 3350
rect 56825 3380 56865 3385
rect 56825 3350 56830 3380
rect 56860 3350 56865 3380
rect 56825 3345 56865 3350
rect 56935 3380 56975 3385
rect 56935 3350 56940 3380
rect 56970 3350 56975 3380
rect 56935 3345 56975 3350
rect 57045 3380 57085 3385
rect 57045 3350 57050 3380
rect 57080 3350 57085 3380
rect 57045 3345 57085 3350
rect 57155 3380 57195 3385
rect 57155 3350 57160 3380
rect 57190 3350 57195 3380
rect 57155 3345 57195 3350
rect 57265 3380 57305 3385
rect 57265 3350 57270 3380
rect 57300 3350 57305 3380
rect 57265 3345 57305 3350
rect 57375 3380 57415 3385
rect 57375 3350 57380 3380
rect 57410 3350 57415 3380
rect 57375 3345 57415 3350
rect 57485 3380 57525 3385
rect 57485 3350 57490 3380
rect 57520 3350 57525 3380
rect 57485 3345 57525 3350
rect 58010 3380 58050 3385
rect 58010 3350 58015 3380
rect 58045 3350 58050 3380
rect 58010 3345 58050 3350
rect 55760 2750 55780 3345
rect 56280 3240 56310 3345
rect 56330 3335 56370 3340
rect 56330 3305 56335 3335
rect 56365 3305 56370 3335
rect 56330 3300 56370 3305
rect 56280 3220 56285 3240
rect 56305 3220 56310 3240
rect 56280 3180 56310 3220
rect 56335 3240 56365 3300
rect 56335 3220 56340 3240
rect 56360 3220 56365 3240
rect 56335 3205 56365 3220
rect 56390 3240 56420 3345
rect 56440 3290 56480 3295
rect 56440 3260 56445 3290
rect 56475 3260 56480 3290
rect 56440 3255 56480 3260
rect 56390 3220 56395 3240
rect 56415 3220 56420 3240
rect 56390 3210 56420 3220
rect 56445 3240 56475 3255
rect 56445 3220 56450 3240
rect 56470 3220 56475 3240
rect 56280 3160 56285 3180
rect 56305 3160 56310 3180
rect 56330 3200 56370 3205
rect 56330 3170 56335 3200
rect 56365 3170 56370 3200
rect 56330 3165 56370 3170
rect 56390 3180 56420 3190
rect 56280 3150 56310 3160
rect 56390 3160 56395 3180
rect 56415 3160 56420 3180
rect 56390 3150 56420 3160
rect 56445 3135 56475 3220
rect 56500 3240 56530 3345
rect 56550 3335 56590 3340
rect 56550 3305 56555 3335
rect 56585 3305 56590 3335
rect 56550 3300 56590 3305
rect 56500 3220 56505 3240
rect 56525 3220 56530 3240
rect 56500 3210 56530 3220
rect 56555 3240 56585 3300
rect 56555 3220 56560 3240
rect 56580 3220 56585 3240
rect 56555 3205 56585 3220
rect 56610 3240 56640 3345
rect 56660 3290 56700 3295
rect 56660 3260 56665 3290
rect 56695 3260 56700 3290
rect 56660 3255 56700 3260
rect 56610 3220 56615 3240
rect 56635 3220 56640 3240
rect 56610 3210 56640 3220
rect 56665 3240 56695 3255
rect 56665 3220 56670 3240
rect 56690 3220 56695 3240
rect 56550 3200 56590 3205
rect 56550 3170 56555 3200
rect 56585 3170 56590 3200
rect 56550 3165 56590 3170
rect 56665 3135 56695 3220
rect 56720 3240 56750 3345
rect 56770 3335 56810 3340
rect 56770 3305 56775 3335
rect 56805 3305 56810 3335
rect 56770 3300 56810 3305
rect 56720 3220 56725 3240
rect 56745 3220 56750 3240
rect 56720 3210 56750 3220
rect 56775 3240 56805 3300
rect 56775 3220 56780 3240
rect 56800 3220 56805 3240
rect 56775 3205 56805 3220
rect 56830 3240 56860 3345
rect 56880 3290 56920 3295
rect 56880 3260 56885 3290
rect 56915 3260 56920 3290
rect 56880 3255 56920 3260
rect 56830 3220 56835 3240
rect 56855 3220 56860 3240
rect 56830 3210 56860 3220
rect 56885 3240 56915 3255
rect 56885 3220 56890 3240
rect 56910 3220 56915 3240
rect 56770 3200 56810 3205
rect 56770 3170 56775 3200
rect 56805 3170 56810 3200
rect 56770 3165 56810 3170
rect 56830 3180 56860 3190
rect 56830 3160 56835 3180
rect 56855 3160 56860 3180
rect 56830 3150 56860 3160
rect 56440 3130 56490 3135
rect 56440 3100 56445 3130
rect 56475 3100 56490 3130
rect 56440 3095 56490 3100
rect 56660 3130 56700 3135
rect 56660 3100 56665 3130
rect 56695 3100 56700 3130
rect 56660 3095 56700 3100
rect 56470 3030 56490 3095
rect 56140 3025 56180 3030
rect 55940 3020 55980 3025
rect 55940 2990 55945 3020
rect 55975 2990 55980 3020
rect 55940 2985 55980 2990
rect 56040 3020 56070 3025
rect 56140 2995 56145 3025
rect 56175 2995 56180 3025
rect 56140 2990 56180 2995
rect 56250 3025 56290 3030
rect 56250 2995 56255 3025
rect 56285 2995 56290 3025
rect 56250 2990 56290 2995
rect 56360 3025 56400 3030
rect 56360 2995 56365 3025
rect 56395 2995 56400 3025
rect 56360 2990 56400 2995
rect 56470 3025 56510 3030
rect 56470 2995 56475 3025
rect 56505 2995 56510 3025
rect 56470 2990 56510 2995
rect 56580 3025 56620 3030
rect 56580 2995 56585 3025
rect 56615 2995 56620 3025
rect 56580 2990 56620 2995
rect 56690 3020 56720 3025
rect 56040 2985 56070 2990
rect 55750 2745 55790 2750
rect 55750 2715 55755 2745
rect 55785 2715 55790 2745
rect 55750 2710 55790 2715
rect 55600 2550 55605 2580
rect 55635 2550 55645 2580
rect 55675 2550 55685 2580
rect 55715 2550 55720 2580
rect 55600 2540 55720 2550
rect 55600 2510 55605 2540
rect 55635 2510 55645 2540
rect 55675 2510 55685 2540
rect 55715 2510 55720 2540
rect 55600 2500 55720 2510
rect 55600 2470 55605 2500
rect 55635 2470 55645 2500
rect 55675 2470 55685 2500
rect 55715 2470 55720 2500
rect 54820 2290 54860 2295
rect 54820 2260 54825 2290
rect 54855 2260 54860 2290
rect 54820 2255 54860 2260
rect 55480 2290 55520 2295
rect 55480 2260 55485 2290
rect 55515 2260 55520 2290
rect 55480 2255 55520 2260
rect 54825 2210 54855 2255
rect 54875 2245 54915 2250
rect 54875 2215 54880 2245
rect 54910 2215 54915 2245
rect 54875 2210 54915 2215
rect 54985 2245 55025 2250
rect 54985 2215 54990 2245
rect 55020 2215 55025 2245
rect 54985 2210 55025 2215
rect 55095 2245 55135 2250
rect 55095 2215 55100 2245
rect 55130 2215 55135 2245
rect 55095 2210 55135 2215
rect 55205 2245 55245 2250
rect 55205 2215 55210 2245
rect 55240 2215 55245 2245
rect 55205 2210 55245 2215
rect 55315 2245 55355 2250
rect 55315 2215 55320 2245
rect 55350 2215 55355 2245
rect 55315 2210 55355 2215
rect 55425 2245 55465 2250
rect 55425 2215 55430 2245
rect 55460 2215 55465 2245
rect 55425 2210 55465 2215
rect 55485 2210 55515 2255
rect 54825 2190 54830 2210
rect 54850 2190 54855 2210
rect 54825 2150 54855 2190
rect 54825 1980 54830 2150
rect 54850 1980 54855 2150
rect 54825 1970 54855 1980
rect 54880 2150 54910 2210
rect 54930 2200 54970 2205
rect 54930 2170 54935 2200
rect 54965 2170 54970 2200
rect 54930 2165 54970 2170
rect 54880 1980 54885 2150
rect 54905 1980 54910 2150
rect 54880 1970 54910 1980
rect 54935 2150 54965 2165
rect 54935 1980 54940 2150
rect 54960 1980 54965 2150
rect 54935 1950 54965 1980
rect 54990 2150 55020 2210
rect 55040 2200 55080 2205
rect 55040 2170 55045 2200
rect 55075 2170 55080 2200
rect 55040 2165 55080 2170
rect 54990 1980 54995 2150
rect 55015 1980 55020 2150
rect 54990 1970 55020 1980
rect 55045 2150 55075 2165
rect 55045 1980 55050 2150
rect 55070 1980 55075 2150
rect 55045 1950 55075 1980
rect 55100 2150 55130 2210
rect 55150 2200 55190 2205
rect 55150 2170 55155 2200
rect 55185 2170 55190 2200
rect 55150 2165 55190 2170
rect 55100 1980 55105 2150
rect 55125 1980 55130 2150
rect 55100 1970 55130 1980
rect 55155 2150 55185 2165
rect 55155 1980 55160 2150
rect 55180 1980 55185 2150
rect 55155 1950 55185 1980
rect 55210 2150 55240 2210
rect 55260 2200 55300 2205
rect 55260 2170 55265 2200
rect 55295 2170 55300 2200
rect 55260 2165 55300 2170
rect 55210 1980 55215 2150
rect 55235 1980 55240 2150
rect 55210 1970 55240 1980
rect 55265 2150 55295 2165
rect 55265 1980 55270 2150
rect 55290 1980 55295 2150
rect 55265 1950 55295 1980
rect 55320 2150 55350 2210
rect 55370 2200 55410 2205
rect 55370 2170 55375 2200
rect 55405 2170 55410 2200
rect 55370 2165 55410 2170
rect 55320 1980 55325 2150
rect 55345 1980 55350 2150
rect 55320 1970 55350 1980
rect 55375 2150 55405 2165
rect 55375 1980 55380 2150
rect 55400 1980 55405 2150
rect 55375 1950 55405 1980
rect 55430 2150 55460 2210
rect 55430 1980 55435 2150
rect 55455 1980 55460 2150
rect 55430 1970 55460 1980
rect 55485 2190 55490 2210
rect 55510 2190 55515 2210
rect 55485 2150 55515 2190
rect 55485 1980 55490 2150
rect 55510 1980 55515 2150
rect 55485 1970 55515 1980
rect 54680 1945 54720 1950
rect 54680 1915 54685 1945
rect 54715 1915 54720 1945
rect 54680 1910 54720 1915
rect 54930 1945 54970 1950
rect 54930 1915 54935 1945
rect 54965 1915 54970 1945
rect 54930 1910 54970 1915
rect 55040 1945 55080 1950
rect 55040 1915 55045 1945
rect 55075 1915 55080 1945
rect 55040 1910 55080 1915
rect 55150 1945 55190 1950
rect 55150 1915 55155 1945
rect 55185 1915 55190 1945
rect 55150 1910 55190 1915
rect 55260 1945 55300 1950
rect 55260 1915 55265 1945
rect 55295 1915 55300 1945
rect 55260 1910 55300 1915
rect 55370 1945 55410 1950
rect 55370 1915 55375 1945
rect 55405 1915 55410 1945
rect 55370 1910 55410 1915
rect 54185 1680 54195 1710
rect 54225 1680 54245 1710
rect 54275 1680 54295 1710
rect 54325 1680 54345 1710
rect 54375 1680 54395 1710
rect 54425 1680 54435 1710
rect 54185 1660 54435 1680
rect 54185 1630 54195 1660
rect 54225 1630 54245 1660
rect 54275 1630 54295 1660
rect 54325 1630 54345 1660
rect 54375 1630 54395 1660
rect 54425 1630 54435 1660
rect 54185 1610 54435 1630
rect 54185 1580 54195 1610
rect 54225 1580 54245 1610
rect 54275 1580 54295 1610
rect 54325 1580 54345 1610
rect 54375 1580 54395 1610
rect 54425 1580 54435 1610
rect 54185 1185 54435 1580
rect 54460 1395 54495 1401
rect 54460 1355 54495 1360
rect 54520 1395 54555 1400
rect 54520 1355 54555 1360
rect 54580 1395 54615 1400
rect 54580 1355 54615 1360
rect 54640 1395 54675 1400
rect 54640 1355 54675 1360
rect 54470 1290 54490 1355
rect 54590 1340 54610 1355
rect 54690 1340 54710 1910
rect 55315 1880 55355 1885
rect 55315 1850 55320 1880
rect 55350 1850 55355 1880
rect 55315 1840 55355 1850
rect 55315 1810 55320 1840
rect 55350 1810 55355 1840
rect 55315 1805 55355 1810
rect 55600 1880 55720 2470
rect 55760 2295 55780 2710
rect 55750 2290 55790 2295
rect 55750 2260 55755 2290
rect 55785 2260 55790 2290
rect 55750 2255 55790 2260
rect 55895 2270 55935 2275
rect 55600 1850 55605 1880
rect 55635 1850 55645 1880
rect 55675 1850 55685 1880
rect 55715 1850 55720 1880
rect 55600 1840 55720 1850
rect 55600 1810 55605 1840
rect 55635 1810 55645 1840
rect 55675 1810 55685 1840
rect 55715 1810 55720 1840
rect 55600 1805 55720 1810
rect 54725 1760 54765 1765
rect 54725 1730 54730 1760
rect 54760 1730 54765 1760
rect 54725 1725 54765 1730
rect 54930 1760 54970 1765
rect 54930 1730 54935 1760
rect 54965 1730 54970 1760
rect 54930 1725 54970 1730
rect 55040 1760 55080 1765
rect 55040 1730 55045 1760
rect 55075 1730 55080 1760
rect 55040 1725 55080 1730
rect 55150 1760 55190 1765
rect 55150 1730 55155 1760
rect 55185 1730 55190 1760
rect 55150 1725 55190 1730
rect 55260 1760 55300 1765
rect 55260 1730 55265 1760
rect 55295 1730 55300 1760
rect 55260 1725 55300 1730
rect 55370 1760 55410 1765
rect 55370 1730 55375 1760
rect 55405 1730 55410 1760
rect 55370 1725 55410 1730
rect 54735 1395 54755 1725
rect 54825 1710 54855 1720
rect 54825 1440 54830 1710
rect 54850 1440 54855 1710
rect 54825 1400 54855 1440
rect 54725 1390 54765 1395
rect 54725 1360 54730 1390
rect 54760 1360 54765 1390
rect 54725 1355 54765 1360
rect 54825 1380 54830 1400
rect 54850 1380 54855 1400
rect 54880 1710 54910 1720
rect 54880 1440 54885 1710
rect 54905 1440 54910 1710
rect 54880 1380 54910 1440
rect 54935 1710 54965 1725
rect 54935 1440 54940 1710
rect 54960 1440 54965 1710
rect 54935 1425 54965 1440
rect 54990 1710 55020 1720
rect 54990 1440 54995 1710
rect 55015 1440 55020 1710
rect 54930 1420 54970 1425
rect 54930 1390 54935 1420
rect 54965 1390 54970 1420
rect 54930 1385 54970 1390
rect 54990 1380 55020 1440
rect 55045 1710 55075 1725
rect 55045 1440 55050 1710
rect 55070 1440 55075 1710
rect 55045 1425 55075 1440
rect 55100 1710 55130 1720
rect 55100 1440 55105 1710
rect 55125 1440 55130 1710
rect 55040 1420 55080 1425
rect 55040 1390 55045 1420
rect 55075 1390 55080 1420
rect 55040 1385 55080 1390
rect 55100 1380 55130 1440
rect 55155 1710 55185 1725
rect 55155 1440 55160 1710
rect 55180 1440 55185 1710
rect 55155 1425 55185 1440
rect 55210 1710 55240 1720
rect 55210 1440 55215 1710
rect 55235 1440 55240 1710
rect 55150 1420 55190 1425
rect 55150 1390 55155 1420
rect 55185 1390 55190 1420
rect 55150 1385 55190 1390
rect 55210 1380 55240 1440
rect 55265 1710 55295 1725
rect 55265 1440 55270 1710
rect 55290 1440 55295 1710
rect 55265 1425 55295 1440
rect 55320 1710 55350 1720
rect 55320 1440 55325 1710
rect 55345 1440 55350 1710
rect 55260 1420 55300 1425
rect 55260 1390 55265 1420
rect 55295 1390 55300 1420
rect 55260 1385 55300 1390
rect 55320 1380 55350 1440
rect 55375 1710 55405 1725
rect 55375 1440 55380 1710
rect 55400 1440 55405 1710
rect 55375 1425 55405 1440
rect 55430 1710 55460 1720
rect 55430 1440 55435 1710
rect 55455 1440 55460 1710
rect 55370 1420 55410 1425
rect 55370 1390 55375 1420
rect 55405 1390 55410 1420
rect 55370 1385 55410 1390
rect 55430 1380 55460 1440
rect 55485 1710 55515 1720
rect 55485 1440 55490 1710
rect 55510 1440 55515 1710
rect 55485 1400 55515 1440
rect 55485 1380 55490 1400
rect 55510 1380 55515 1400
rect 55760 1380 55780 2255
rect 55895 2240 55900 2270
rect 55930 2240 55935 2270
rect 55895 2235 55935 2240
rect 54580 1335 54620 1340
rect 54580 1305 54585 1335
rect 54615 1305 54620 1335
rect 54580 1300 54620 1305
rect 54680 1335 54720 1340
rect 54825 1335 54855 1380
rect 54875 1375 54915 1380
rect 54875 1345 54880 1375
rect 54910 1345 54915 1375
rect 54875 1340 54915 1345
rect 54985 1375 55025 1380
rect 54985 1345 54990 1375
rect 55020 1345 55025 1375
rect 54985 1340 55025 1345
rect 55095 1375 55135 1380
rect 55095 1345 55100 1375
rect 55130 1345 55135 1375
rect 55095 1340 55135 1345
rect 55205 1375 55245 1380
rect 55205 1345 55210 1375
rect 55240 1345 55245 1375
rect 55205 1340 55245 1345
rect 55315 1375 55355 1380
rect 55315 1345 55320 1375
rect 55350 1345 55355 1375
rect 55315 1340 55355 1345
rect 55425 1375 55465 1380
rect 55425 1345 55430 1375
rect 55460 1345 55465 1375
rect 55425 1340 55465 1345
rect 55485 1335 55515 1380
rect 55750 1375 55790 1380
rect 55750 1345 55755 1375
rect 55785 1345 55790 1375
rect 55750 1340 55790 1345
rect 54680 1305 54685 1335
rect 54715 1305 54720 1335
rect 54680 1300 54720 1305
rect 54820 1330 54860 1335
rect 54820 1300 54825 1330
rect 54855 1300 54860 1330
rect 54820 1295 54860 1300
rect 55480 1330 55520 1335
rect 55480 1300 55485 1330
rect 55515 1300 55520 1330
rect 55480 1295 55520 1300
rect 55830 1330 55870 1335
rect 55830 1300 55835 1330
rect 55865 1300 55870 1330
rect 55830 1295 55870 1300
rect 54460 1285 54500 1290
rect 54460 1255 54465 1285
rect 54495 1255 54500 1285
rect 54460 1250 54500 1255
rect 54595 1240 54635 1245
rect 54595 1210 54600 1240
rect 54630 1210 54635 1240
rect 54595 1205 54635 1210
rect 55180 1240 55220 1245
rect 55180 1210 55185 1240
rect 55215 1210 55220 1240
rect 55180 1205 55220 1210
rect 54185 1155 54190 1185
rect 54220 1155 54230 1185
rect 54260 1155 54275 1185
rect 54305 1155 54315 1185
rect 54345 1155 54360 1185
rect 54390 1155 54400 1185
rect 54430 1155 54435 1185
rect 54185 1145 54435 1155
rect 54185 1115 54190 1145
rect 54220 1115 54230 1145
rect 54260 1115 54275 1145
rect 54305 1115 54315 1145
rect 54345 1115 54360 1145
rect 54390 1115 54400 1145
rect 54430 1115 54435 1145
rect 54185 1105 54435 1115
rect 54185 1075 54190 1105
rect 54220 1075 54230 1105
rect 54260 1075 54275 1105
rect 54305 1075 54315 1105
rect 54345 1075 54360 1105
rect 54390 1075 54400 1105
rect 54430 1075 54435 1105
rect 54185 1070 54435 1075
rect 54605 1055 54625 1205
rect 54660 1185 54700 1190
rect 54660 1155 54665 1185
rect 54695 1155 54700 1185
rect 54660 1145 54700 1155
rect 54660 1115 54665 1145
rect 54695 1115 54700 1145
rect 54660 1105 54700 1115
rect 54660 1075 54665 1105
rect 54695 1075 54700 1105
rect 54660 1070 54700 1075
rect 54930 1185 55370 1190
rect 54930 1155 54935 1185
rect 54965 1155 54975 1185
rect 55005 1155 55015 1185
rect 55045 1155 55055 1185
rect 55085 1155 55095 1185
rect 55125 1155 55135 1185
rect 55165 1155 55175 1185
rect 55205 1155 55215 1185
rect 55245 1155 55255 1185
rect 55285 1155 55295 1185
rect 55325 1155 55335 1185
rect 55365 1155 55370 1185
rect 54930 1145 55370 1155
rect 54930 1115 54935 1145
rect 54965 1115 54975 1145
rect 55005 1115 55015 1145
rect 55045 1115 55055 1145
rect 55085 1115 55095 1145
rect 55125 1115 55135 1145
rect 55165 1115 55175 1145
rect 55205 1115 55215 1145
rect 55245 1115 55255 1145
rect 55285 1115 55295 1145
rect 55325 1115 55335 1145
rect 55365 1115 55370 1145
rect 54930 1105 55370 1115
rect 54930 1075 54935 1105
rect 54965 1075 54975 1105
rect 55005 1075 55015 1105
rect 55045 1075 55055 1105
rect 55085 1075 55095 1105
rect 55125 1075 55135 1105
rect 55165 1075 55175 1105
rect 55205 1075 55215 1105
rect 55245 1075 55255 1105
rect 55285 1075 55295 1105
rect 55325 1075 55335 1105
rect 55365 1075 55370 1105
rect 54930 1070 55370 1075
rect 54600 1050 54635 1055
rect 54600 1010 54635 1015
rect 54660 1050 54695 1070
rect 54660 1010 54695 1015
rect 54835 1040 54865 1050
rect 54835 370 54840 1040
rect 54860 370 54865 1040
rect 54835 330 54865 370
rect 54935 1040 54965 1070
rect 54935 370 54940 1040
rect 54960 370 54965 1040
rect 54935 355 54965 370
rect 55035 1040 55065 1050
rect 55035 370 55040 1040
rect 55060 370 55065 1040
rect 54835 310 54840 330
rect 54860 310 54865 330
rect 54930 350 54970 355
rect 54930 320 54935 350
rect 54965 320 54970 350
rect 54930 315 54970 320
rect 54835 50 54865 310
rect 55035 50 55065 370
rect 55135 1040 55165 1070
rect 55135 370 55140 1040
rect 55160 370 55165 1040
rect 55135 355 55165 370
rect 55235 1040 55265 1050
rect 55235 370 55240 1040
rect 55260 370 55265 1040
rect 55130 350 55170 355
rect 55130 320 55135 350
rect 55165 320 55170 350
rect 55130 315 55170 320
rect 55235 50 55265 370
rect 55335 1040 55365 1070
rect 55335 370 55340 1040
rect 55360 370 55365 1040
rect 55335 355 55365 370
rect 55435 1040 55465 1050
rect 55435 370 55440 1040
rect 55460 370 55465 1040
rect 55840 745 55860 1295
rect 55830 740 55870 745
rect 55830 710 55835 740
rect 55865 710 55870 740
rect 55830 705 55870 710
rect 55330 350 55370 355
rect 55330 320 55335 350
rect 55365 320 55370 350
rect 55330 315 55370 320
rect 55435 330 55465 370
rect 55435 310 55440 330
rect 55460 310 55465 330
rect 55435 50 55465 310
rect 55840 50 55860 705
rect 55905 600 55925 2235
rect 55950 1290 55970 2985
rect 56085 2980 56125 2985
rect 56085 2950 56090 2980
rect 56120 2950 56125 2980
rect 56085 2945 56125 2950
rect 56035 2930 56065 2940
rect 56035 2910 56040 2930
rect 56060 2910 56065 2930
rect 56035 2870 56065 2910
rect 56035 2850 56040 2870
rect 56060 2850 56065 2870
rect 56090 2930 56120 2945
rect 56090 2910 56095 2930
rect 56115 2910 56120 2930
rect 56090 2850 56120 2910
rect 56145 2930 56175 2990
rect 56195 2980 56235 2985
rect 56195 2950 56200 2980
rect 56230 2950 56235 2980
rect 56195 2945 56235 2950
rect 56145 2910 56150 2930
rect 56170 2910 56175 2930
rect 56145 2895 56175 2910
rect 56200 2930 56230 2945
rect 56200 2910 56205 2930
rect 56225 2910 56230 2930
rect 56140 2890 56180 2895
rect 56140 2860 56145 2890
rect 56175 2860 56180 2890
rect 56140 2855 56180 2860
rect 56200 2850 56230 2910
rect 56255 2930 56285 2990
rect 56305 2980 56345 2985
rect 56305 2950 56310 2980
rect 56340 2950 56345 2980
rect 56305 2945 56345 2950
rect 56255 2910 56260 2930
rect 56280 2910 56285 2930
rect 56255 2895 56285 2910
rect 56310 2930 56340 2945
rect 56310 2910 56315 2930
rect 56335 2910 56340 2930
rect 56250 2890 56290 2895
rect 56250 2860 56255 2890
rect 56285 2860 56290 2890
rect 56250 2855 56290 2860
rect 56310 2850 56340 2910
rect 56365 2930 56395 2990
rect 56415 2980 56455 2985
rect 56415 2950 56420 2980
rect 56450 2950 56455 2980
rect 56415 2945 56455 2950
rect 56365 2910 56370 2930
rect 56390 2910 56395 2930
rect 56365 2895 56395 2910
rect 56420 2930 56450 2945
rect 56420 2910 56425 2930
rect 56445 2910 56450 2930
rect 56360 2890 56400 2895
rect 56360 2860 56365 2890
rect 56395 2860 56400 2890
rect 56360 2855 56400 2860
rect 56420 2850 56450 2910
rect 56475 2930 56505 2990
rect 56525 2980 56565 2985
rect 56525 2950 56530 2980
rect 56560 2950 56565 2980
rect 56525 2945 56565 2950
rect 56475 2910 56480 2930
rect 56500 2910 56505 2930
rect 56475 2895 56505 2910
rect 56530 2930 56560 2945
rect 56530 2910 56535 2930
rect 56555 2910 56560 2930
rect 56470 2890 56510 2895
rect 56470 2860 56475 2890
rect 56505 2860 56510 2890
rect 56470 2855 56510 2860
rect 56530 2850 56560 2910
rect 56585 2930 56615 2990
rect 56690 2985 56720 2990
rect 56635 2980 56675 2985
rect 56635 2950 56640 2980
rect 56670 2950 56675 2980
rect 56635 2945 56675 2950
rect 56585 2910 56590 2930
rect 56610 2910 56615 2930
rect 56585 2895 56615 2910
rect 56640 2930 56670 2945
rect 56640 2910 56645 2930
rect 56665 2910 56670 2930
rect 56580 2890 56620 2895
rect 56580 2860 56585 2890
rect 56615 2860 56620 2890
rect 56580 2855 56620 2860
rect 56640 2850 56670 2910
rect 56695 2930 56725 2940
rect 56695 2910 56700 2930
rect 56720 2910 56725 2930
rect 56695 2870 56725 2910
rect 56695 2850 56700 2870
rect 56720 2850 56725 2870
rect 56835 2850 56855 3150
rect 56885 3135 56915 3220
rect 56940 3240 56970 3345
rect 56990 3335 57030 3340
rect 56990 3305 56995 3335
rect 57025 3305 57030 3335
rect 56990 3300 57030 3305
rect 56940 3220 56945 3240
rect 56965 3220 56970 3240
rect 56940 3210 56970 3220
rect 56995 3240 57025 3300
rect 56995 3220 57000 3240
rect 57020 3220 57025 3240
rect 56995 3205 57025 3220
rect 57050 3240 57080 3345
rect 57100 3290 57140 3295
rect 57100 3260 57105 3290
rect 57135 3260 57140 3290
rect 57100 3255 57140 3260
rect 57050 3220 57055 3240
rect 57075 3220 57080 3240
rect 57050 3210 57080 3220
rect 57105 3240 57135 3255
rect 57105 3220 57110 3240
rect 57130 3220 57135 3240
rect 56990 3200 57030 3205
rect 56990 3170 56995 3200
rect 57025 3170 57030 3200
rect 56990 3165 57030 3170
rect 57105 3135 57135 3220
rect 57160 3240 57190 3345
rect 57210 3335 57250 3340
rect 57210 3305 57215 3335
rect 57245 3305 57250 3335
rect 57210 3300 57250 3305
rect 57160 3220 57165 3240
rect 57185 3220 57190 3240
rect 57160 3210 57190 3220
rect 57215 3240 57245 3300
rect 57215 3220 57220 3240
rect 57240 3220 57245 3240
rect 57215 3205 57245 3220
rect 57270 3240 57300 3345
rect 57320 3290 57360 3295
rect 57320 3260 57325 3290
rect 57355 3260 57360 3290
rect 57320 3255 57360 3260
rect 57270 3220 57275 3240
rect 57295 3220 57300 3240
rect 57270 3210 57300 3220
rect 57325 3240 57355 3255
rect 57325 3220 57330 3240
rect 57350 3220 57355 3240
rect 57210 3200 57250 3205
rect 57210 3170 57215 3200
rect 57245 3170 57250 3200
rect 57210 3165 57250 3170
rect 56880 3130 56920 3135
rect 56880 3100 56885 3130
rect 56915 3100 56920 3130
rect 56880 3095 56920 3100
rect 57100 3130 57140 3135
rect 57100 3100 57105 3130
rect 57135 3100 57140 3130
rect 57100 3095 57140 3100
rect 57220 3030 57240 3165
rect 57325 3135 57355 3220
rect 57380 3240 57410 3345
rect 57430 3335 57470 3340
rect 57430 3305 57435 3335
rect 57465 3305 57470 3335
rect 57430 3300 57470 3305
rect 57380 3220 57385 3240
rect 57405 3220 57410 3240
rect 57380 3210 57410 3220
rect 57435 3240 57465 3300
rect 57435 3220 57440 3240
rect 57460 3220 57465 3240
rect 57435 3205 57465 3220
rect 57490 3240 57520 3345
rect 57490 3220 57495 3240
rect 57515 3220 57520 3240
rect 57430 3200 57470 3205
rect 57430 3170 57435 3200
rect 57465 3170 57470 3200
rect 57430 3165 57470 3170
rect 57490 3180 57520 3220
rect 57490 3160 57495 3180
rect 57515 3160 57520 3180
rect 57490 3150 57520 3160
rect 57320 3130 57360 3135
rect 57320 3100 57325 3130
rect 57355 3100 57360 3130
rect 57320 3095 57360 3100
rect 57180 3025 57240 3030
rect 57080 3020 57110 3025
rect 57180 2995 57185 3025
rect 57215 2995 57240 3025
rect 57180 2990 57240 2995
rect 57290 3025 57330 3030
rect 57290 2995 57295 3025
rect 57325 2995 57330 3025
rect 57290 2990 57330 2995
rect 57400 3025 57440 3030
rect 57400 2995 57405 3025
rect 57435 2995 57440 3025
rect 57400 2990 57440 2995
rect 57510 3025 57550 3030
rect 57510 2995 57515 3025
rect 57545 2995 57550 3025
rect 57510 2990 57550 2995
rect 57620 3025 57660 3030
rect 57620 2995 57625 3025
rect 57655 2995 57660 3025
rect 57620 2990 57660 2995
rect 57730 3020 57760 3025
rect 57080 2985 57110 2990
rect 57125 2980 57165 2985
rect 57125 2950 57130 2980
rect 57160 2950 57165 2980
rect 57125 2945 57165 2950
rect 57075 2930 57105 2940
rect 57075 2910 57080 2930
rect 57100 2910 57105 2930
rect 57075 2870 57105 2910
rect 57075 2850 57080 2870
rect 57100 2850 57105 2870
rect 57130 2930 57160 2945
rect 57130 2910 57135 2930
rect 57155 2910 57160 2930
rect 57130 2850 57160 2910
rect 57185 2930 57215 2990
rect 57185 2910 57190 2930
rect 57210 2910 57215 2930
rect 57185 2895 57215 2910
rect 57240 2930 57270 2940
rect 57240 2910 57245 2930
rect 57265 2910 57270 2930
rect 57180 2890 57220 2895
rect 57180 2860 57185 2890
rect 57215 2860 57220 2890
rect 57180 2855 57220 2860
rect 56035 2750 56065 2850
rect 56085 2845 56125 2850
rect 56085 2815 56090 2845
rect 56120 2815 56125 2845
rect 56085 2810 56125 2815
rect 56195 2845 56235 2850
rect 56195 2815 56200 2845
rect 56230 2815 56235 2845
rect 56195 2810 56235 2815
rect 56305 2845 56345 2850
rect 56305 2815 56310 2845
rect 56340 2815 56345 2845
rect 56305 2810 56345 2815
rect 56415 2845 56455 2850
rect 56415 2815 56420 2845
rect 56450 2815 56455 2845
rect 56415 2810 56455 2815
rect 56525 2845 56565 2850
rect 56525 2815 56530 2845
rect 56560 2815 56565 2845
rect 56525 2810 56565 2815
rect 56635 2845 56675 2850
rect 56635 2815 56640 2845
rect 56670 2815 56675 2845
rect 56635 2810 56675 2815
rect 56580 2800 56610 2805
rect 56095 2790 56125 2795
rect 56580 2765 56610 2770
rect 56095 2755 56125 2760
rect 56695 2750 56725 2850
rect 56825 2845 56865 2850
rect 56825 2815 56830 2845
rect 56860 2815 56865 2845
rect 56825 2810 56865 2815
rect 57075 2750 57105 2850
rect 57125 2845 57165 2850
rect 57125 2815 57130 2845
rect 57160 2815 57165 2845
rect 57125 2810 57165 2815
rect 57190 2800 57220 2805
rect 57190 2765 57220 2770
rect 56030 2745 56070 2750
rect 56030 2715 56035 2745
rect 56065 2715 56070 2745
rect 56030 2710 56070 2715
rect 56690 2745 56730 2750
rect 56690 2715 56695 2745
rect 56725 2715 56730 2745
rect 56690 2710 56730 2715
rect 57070 2745 57110 2750
rect 57070 2715 57075 2745
rect 57105 2715 57110 2745
rect 57070 2710 57110 2715
rect 57240 2695 57270 2910
rect 57295 2930 57325 2990
rect 57345 2980 57385 2985
rect 57345 2950 57350 2980
rect 57380 2950 57385 2980
rect 57345 2945 57385 2950
rect 57295 2910 57300 2930
rect 57320 2910 57325 2930
rect 57295 2895 57325 2910
rect 57350 2930 57380 2945
rect 57350 2910 57355 2930
rect 57375 2910 57380 2930
rect 57290 2890 57330 2895
rect 57290 2860 57295 2890
rect 57325 2860 57330 2890
rect 57290 2855 57330 2860
rect 57350 2850 57380 2910
rect 57405 2930 57435 2990
rect 57405 2910 57410 2930
rect 57430 2910 57435 2930
rect 57405 2895 57435 2910
rect 57460 2930 57490 2940
rect 57460 2910 57465 2930
rect 57485 2910 57490 2930
rect 57400 2890 57440 2895
rect 57400 2860 57405 2890
rect 57435 2860 57440 2890
rect 57400 2855 57440 2860
rect 57345 2845 57385 2850
rect 57345 2815 57350 2845
rect 57380 2815 57385 2845
rect 57345 2810 57385 2815
rect 56935 2690 56975 2695
rect 56935 2660 56940 2690
rect 56970 2660 56975 2690
rect 56935 2655 56975 2660
rect 57235 2690 57275 2695
rect 57235 2660 57240 2690
rect 57270 2660 57275 2690
rect 57235 2655 57275 2660
rect 56945 2640 56965 2655
rect 57350 2640 57380 2810
rect 57460 2695 57490 2910
rect 57515 2930 57545 2990
rect 57565 2980 57605 2985
rect 57565 2950 57570 2980
rect 57600 2950 57605 2980
rect 57565 2945 57605 2950
rect 57515 2910 57520 2930
rect 57540 2910 57545 2930
rect 57515 2895 57545 2910
rect 57570 2930 57600 2945
rect 57570 2910 57575 2930
rect 57595 2910 57600 2930
rect 57510 2890 57550 2895
rect 57510 2860 57515 2890
rect 57545 2860 57550 2890
rect 57510 2855 57550 2860
rect 57570 2850 57600 2910
rect 57625 2930 57655 2990
rect 57730 2985 57760 2990
rect 57820 3020 57860 3025
rect 57820 2990 57825 3020
rect 57855 2990 57860 3020
rect 57820 2985 57860 2990
rect 57625 2910 57630 2930
rect 57650 2910 57655 2930
rect 57625 2895 57655 2910
rect 57680 2930 57710 2940
rect 57680 2910 57685 2930
rect 57705 2910 57710 2930
rect 57620 2890 57660 2895
rect 57620 2860 57625 2890
rect 57655 2860 57660 2890
rect 57620 2855 57660 2860
rect 57565 2845 57605 2850
rect 57565 2815 57570 2845
rect 57600 2815 57605 2845
rect 57565 2810 57605 2815
rect 57680 2695 57710 2910
rect 57735 2930 57765 2940
rect 57735 2910 57740 2930
rect 57760 2910 57765 2930
rect 57735 2870 57765 2910
rect 57735 2850 57740 2870
rect 57760 2850 57765 2870
rect 57735 2750 57765 2850
rect 57730 2745 57770 2750
rect 57730 2715 57735 2745
rect 57765 2715 57770 2745
rect 57730 2710 57770 2715
rect 57455 2690 57495 2695
rect 57455 2660 57460 2690
rect 57490 2660 57495 2690
rect 57455 2655 57495 2660
rect 57675 2690 57715 2695
rect 57675 2660 57680 2690
rect 57710 2660 57715 2690
rect 57675 2655 57715 2660
rect 56830 2635 56890 2640
rect 56830 2605 56855 2635
rect 56885 2605 56890 2635
rect 56830 2600 56890 2605
rect 56935 2630 56975 2640
rect 56935 2610 56945 2630
rect 56965 2610 56975 2630
rect 56935 2600 56975 2610
rect 57345 2635 57385 2640
rect 57345 2605 57350 2635
rect 57380 2605 57385 2635
rect 57345 2600 57385 2605
rect 56085 2580 56675 2585
rect 56085 2550 56090 2580
rect 56120 2550 56145 2580
rect 56175 2550 56200 2580
rect 56230 2550 56255 2580
rect 56285 2550 56310 2580
rect 56340 2550 56365 2580
rect 56395 2550 56420 2580
rect 56450 2550 56475 2580
rect 56505 2550 56530 2580
rect 56560 2550 56585 2580
rect 56615 2550 56640 2580
rect 56670 2550 56675 2580
rect 56085 2540 56675 2550
rect 56085 2510 56090 2540
rect 56120 2510 56145 2540
rect 56175 2510 56200 2540
rect 56230 2510 56255 2540
rect 56285 2510 56310 2540
rect 56340 2510 56365 2540
rect 56395 2510 56420 2540
rect 56450 2510 56475 2540
rect 56505 2510 56530 2540
rect 56560 2510 56585 2540
rect 56615 2510 56640 2540
rect 56670 2510 56675 2540
rect 56085 2500 56675 2510
rect 56085 2470 56090 2500
rect 56120 2470 56145 2500
rect 56175 2470 56200 2500
rect 56230 2470 56255 2500
rect 56285 2470 56310 2500
rect 56340 2470 56365 2500
rect 56395 2470 56420 2500
rect 56450 2470 56475 2500
rect 56505 2470 56530 2500
rect 56560 2470 56585 2500
rect 56615 2470 56640 2500
rect 56670 2470 56675 2500
rect 56085 2465 56675 2470
rect 55995 2270 56025 2275
rect 55995 2235 56025 2240
rect 56085 2215 56125 2465
rect 56140 2260 56180 2265
rect 56140 2230 56145 2260
rect 56175 2230 56180 2260
rect 56140 2225 56180 2230
rect 56085 2185 56090 2215
rect 56120 2185 56125 2215
rect 56085 2180 56125 2185
rect 56030 2165 56065 2175
rect 56030 2045 56040 2165
rect 56060 2045 56065 2165
rect 56030 2035 56065 2045
rect 56035 2030 56065 2035
rect 56090 2165 56120 2180
rect 56090 2045 56095 2165
rect 56115 2045 56120 2165
rect 56035 2005 56065 2015
rect 56035 1985 56040 2005
rect 56060 1985 56065 2005
rect 56090 1985 56120 2045
rect 56145 2165 56175 2225
rect 56195 2215 56235 2465
rect 56250 2260 56290 2265
rect 56250 2230 56255 2260
rect 56285 2230 56290 2260
rect 56250 2225 56290 2230
rect 56195 2185 56200 2215
rect 56230 2185 56235 2215
rect 56195 2180 56235 2185
rect 56145 2045 56150 2165
rect 56170 2045 56175 2165
rect 56145 2030 56175 2045
rect 56200 2165 56230 2180
rect 56200 2045 56205 2165
rect 56225 2045 56230 2165
rect 56140 2025 56180 2030
rect 56140 1995 56145 2025
rect 56175 1995 56180 2025
rect 56140 1990 56180 1995
rect 56035 1940 56065 1985
rect 56085 1980 56125 1985
rect 56085 1950 56090 1980
rect 56120 1950 56125 1980
rect 56085 1945 56125 1950
rect 56030 1935 56070 1940
rect 56030 1905 56035 1935
rect 56065 1905 56070 1935
rect 56030 1900 56070 1905
rect 56145 1805 56175 1990
rect 56200 1985 56230 2045
rect 56255 2165 56285 2225
rect 56305 2215 56345 2465
rect 56360 2260 56400 2265
rect 56360 2230 56365 2260
rect 56395 2230 56400 2260
rect 56360 2225 56400 2230
rect 56305 2185 56310 2215
rect 56340 2185 56345 2215
rect 56305 2180 56345 2185
rect 56255 2045 56260 2165
rect 56280 2045 56285 2165
rect 56255 2030 56285 2045
rect 56310 2165 56340 2180
rect 56310 2045 56315 2165
rect 56335 2045 56340 2165
rect 56250 2025 56290 2030
rect 56250 1995 56255 2025
rect 56285 1995 56290 2025
rect 56250 1990 56290 1995
rect 56195 1980 56235 1985
rect 56195 1950 56200 1980
rect 56230 1950 56235 1980
rect 56195 1945 56235 1950
rect 56085 1795 56125 1800
rect 56040 1785 56070 1790
rect 56085 1765 56090 1795
rect 56120 1765 56125 1795
rect 56255 1805 56285 1990
rect 56310 1985 56340 2045
rect 56365 2165 56395 2225
rect 56415 2215 56455 2465
rect 56470 2260 56510 2265
rect 56470 2230 56475 2260
rect 56505 2230 56510 2260
rect 56470 2225 56510 2230
rect 56415 2185 56420 2215
rect 56450 2185 56455 2215
rect 56415 2180 56455 2185
rect 56365 2045 56370 2165
rect 56390 2045 56395 2165
rect 56365 2030 56395 2045
rect 56420 2165 56450 2180
rect 56420 2045 56425 2165
rect 56445 2045 56450 2165
rect 56360 2025 56400 2030
rect 56360 1995 56365 2025
rect 56395 1995 56400 2025
rect 56360 1990 56400 1995
rect 56305 1980 56345 1985
rect 56305 1950 56310 1980
rect 56340 1950 56345 1980
rect 56305 1945 56345 1950
rect 56145 1770 56175 1775
rect 56195 1795 56235 1800
rect 56085 1760 56125 1765
rect 56195 1765 56200 1795
rect 56230 1765 56235 1795
rect 56365 1805 56395 1990
rect 56420 1985 56450 2045
rect 56475 2165 56505 2225
rect 56525 2215 56565 2465
rect 56580 2260 56620 2265
rect 56580 2230 56585 2260
rect 56615 2230 56620 2260
rect 56580 2225 56620 2230
rect 56525 2185 56530 2215
rect 56560 2185 56565 2215
rect 56525 2180 56565 2185
rect 56475 2045 56480 2165
rect 56500 2045 56505 2165
rect 56475 2030 56505 2045
rect 56530 2165 56560 2180
rect 56530 2045 56535 2165
rect 56555 2045 56560 2165
rect 56470 2025 56510 2030
rect 56470 1995 56475 2025
rect 56505 1995 56510 2025
rect 56470 1990 56510 1995
rect 56415 1980 56455 1985
rect 56415 1950 56420 1980
rect 56450 1950 56455 1980
rect 56415 1945 56455 1950
rect 56255 1770 56285 1775
rect 56305 1795 56345 1800
rect 56195 1760 56235 1765
rect 56305 1765 56310 1795
rect 56340 1765 56345 1795
rect 56475 1805 56505 1990
rect 56530 1985 56560 2045
rect 56585 2165 56615 2225
rect 56635 2215 56675 2465
rect 56775 2570 56805 2580
rect 56775 2350 56780 2570
rect 56800 2350 56805 2570
rect 56775 2320 56805 2350
rect 56830 2570 56860 2600
rect 56830 2350 56835 2570
rect 56855 2350 56860 2570
rect 56830 2340 56860 2350
rect 56885 2570 56915 2580
rect 56885 2350 56890 2570
rect 56910 2350 56915 2570
rect 56885 2320 56915 2350
rect 56940 2570 56970 2600
rect 57125 2580 57715 2585
rect 56940 2350 56945 2570
rect 56965 2350 56970 2570
rect 56940 2340 56970 2350
rect 56995 2570 57025 2580
rect 56995 2350 57000 2570
rect 57020 2350 57025 2570
rect 56995 2320 57025 2350
rect 57125 2550 57130 2580
rect 57160 2550 57185 2580
rect 57215 2550 57240 2580
rect 57270 2550 57295 2580
rect 57325 2550 57350 2580
rect 57380 2550 57405 2580
rect 57435 2550 57460 2580
rect 57490 2550 57515 2580
rect 57545 2550 57570 2580
rect 57600 2550 57625 2580
rect 57655 2550 57680 2580
rect 57710 2550 57715 2580
rect 57125 2540 57715 2550
rect 57125 2510 57130 2540
rect 57160 2510 57185 2540
rect 57215 2510 57240 2540
rect 57270 2510 57295 2540
rect 57325 2510 57350 2540
rect 57380 2510 57405 2540
rect 57435 2510 57460 2540
rect 57490 2510 57515 2540
rect 57545 2510 57570 2540
rect 57600 2510 57625 2540
rect 57655 2510 57680 2540
rect 57710 2510 57715 2540
rect 57125 2500 57715 2510
rect 57125 2470 57130 2500
rect 57160 2470 57185 2500
rect 57215 2470 57240 2500
rect 57270 2470 57295 2500
rect 57325 2470 57350 2500
rect 57380 2470 57405 2500
rect 57435 2470 57460 2500
rect 57490 2470 57515 2500
rect 57545 2470 57570 2500
rect 57600 2470 57625 2500
rect 57655 2470 57680 2500
rect 57710 2470 57715 2500
rect 57125 2465 57715 2470
rect 56770 2315 56810 2320
rect 56770 2285 56775 2315
rect 56805 2285 56810 2315
rect 56770 2280 56810 2285
rect 56880 2315 56920 2320
rect 56880 2285 56885 2315
rect 56915 2285 56920 2315
rect 56880 2280 56920 2285
rect 56990 2315 57030 2320
rect 56990 2285 56995 2315
rect 57025 2285 57030 2315
rect 56990 2280 57030 2285
rect 56690 2270 56720 2275
rect 56690 2235 56720 2240
rect 57080 2270 57110 2275
rect 57080 2235 57110 2240
rect 56635 2185 56640 2215
rect 56670 2185 56675 2215
rect 56635 2180 56675 2185
rect 57125 2215 57165 2465
rect 57180 2260 57220 2265
rect 57180 2230 57185 2260
rect 57215 2230 57220 2260
rect 57180 2225 57220 2230
rect 57125 2185 57130 2215
rect 57160 2185 57165 2215
rect 57125 2180 57165 2185
rect 56585 2045 56590 2165
rect 56610 2045 56615 2165
rect 56585 2030 56615 2045
rect 56640 2165 56670 2180
rect 56640 2045 56645 2165
rect 56665 2045 56670 2165
rect 56580 2025 56620 2030
rect 56580 1995 56585 2025
rect 56615 1995 56620 2025
rect 56580 1990 56620 1995
rect 56525 1980 56565 1985
rect 56525 1950 56530 1980
rect 56560 1950 56565 1980
rect 56525 1945 56565 1950
rect 56365 1770 56395 1775
rect 56415 1795 56455 1800
rect 56305 1760 56345 1765
rect 56415 1765 56420 1795
rect 56450 1765 56455 1795
rect 56585 1805 56615 1990
rect 56640 1985 56670 2045
rect 56695 2165 56765 2175
rect 56695 2045 56700 2165
rect 56720 2045 56765 2165
rect 56695 2035 56765 2045
rect 57035 2165 57105 2175
rect 57035 2045 57080 2165
rect 57100 2045 57105 2165
rect 57035 2035 57105 2045
rect 56695 2005 56725 2035
rect 56695 1985 56700 2005
rect 56720 1985 56725 2005
rect 56635 1980 56675 1985
rect 56635 1950 56640 1980
rect 56670 1950 56675 1980
rect 56635 1945 56675 1950
rect 56695 1940 56725 1985
rect 57075 2005 57105 2035
rect 57075 1985 57080 2005
rect 57100 1985 57105 2005
rect 57130 2165 57160 2180
rect 57130 2045 57135 2165
rect 57155 2045 57160 2165
rect 57130 1985 57160 2045
rect 57185 2165 57215 2225
rect 57235 2215 57275 2465
rect 57290 2260 57330 2265
rect 57290 2230 57295 2260
rect 57325 2230 57330 2260
rect 57290 2225 57330 2230
rect 57235 2185 57240 2215
rect 57270 2185 57275 2215
rect 57235 2180 57275 2185
rect 57185 2045 57190 2165
rect 57210 2045 57215 2165
rect 57185 2030 57215 2045
rect 57240 2165 57270 2180
rect 57240 2045 57245 2165
rect 57265 2045 57270 2165
rect 57180 2025 57220 2030
rect 57180 1995 57185 2025
rect 57215 1995 57220 2025
rect 57180 1990 57220 1995
rect 57075 1940 57105 1985
rect 57125 1980 57165 1985
rect 57125 1950 57130 1980
rect 57160 1950 57165 1980
rect 57125 1945 57165 1950
rect 56690 1935 56730 1940
rect 56690 1905 56695 1935
rect 56725 1905 56730 1935
rect 56690 1900 56730 1905
rect 57070 1935 57110 1940
rect 57070 1905 57075 1935
rect 57105 1905 57110 1935
rect 57070 1900 57110 1905
rect 56475 1770 56505 1775
rect 56525 1795 56565 1800
rect 56415 1760 56455 1765
rect 56525 1765 56530 1795
rect 56560 1765 56565 1795
rect 56585 1770 56615 1775
rect 56635 1795 56675 1800
rect 56525 1760 56565 1765
rect 56635 1765 56640 1795
rect 56670 1765 56675 1795
rect 56635 1760 56675 1765
rect 56690 1785 56720 1790
rect 56040 1750 56070 1755
rect 56035 1695 56065 1705
rect 56035 1575 56040 1695
rect 56060 1575 56065 1695
rect 56035 1565 56065 1575
rect 56090 1695 56120 1760
rect 56140 1750 56180 1755
rect 56140 1720 56145 1750
rect 56175 1720 56180 1750
rect 56140 1715 56180 1720
rect 56090 1575 56095 1695
rect 56115 1575 56120 1695
rect 56090 1560 56120 1575
rect 56145 1695 56175 1715
rect 56145 1575 56150 1695
rect 56170 1575 56175 1695
rect 56085 1555 56125 1560
rect 56035 1535 56065 1545
rect 56035 1515 56040 1535
rect 56060 1515 56065 1535
rect 56085 1525 56090 1555
rect 56120 1525 56125 1555
rect 56085 1520 56125 1525
rect 56035 1505 56065 1515
rect 56145 1505 56175 1575
rect 56200 1695 56230 1760
rect 56250 1750 56290 1755
rect 56250 1720 56255 1750
rect 56285 1720 56290 1750
rect 56250 1715 56290 1720
rect 56200 1575 56205 1695
rect 56225 1575 56230 1695
rect 56200 1560 56230 1575
rect 56255 1695 56285 1715
rect 56255 1575 56260 1695
rect 56280 1575 56285 1695
rect 56195 1555 56235 1560
rect 56195 1525 56200 1555
rect 56230 1525 56235 1555
rect 56195 1520 56235 1525
rect 56255 1505 56285 1575
rect 56310 1695 56340 1760
rect 56360 1750 56400 1755
rect 56360 1720 56365 1750
rect 56395 1720 56400 1750
rect 56360 1715 56400 1720
rect 56310 1575 56315 1695
rect 56335 1575 56340 1695
rect 56310 1560 56340 1575
rect 56365 1695 56395 1715
rect 56365 1575 56370 1695
rect 56390 1575 56395 1695
rect 56305 1555 56345 1560
rect 56305 1525 56310 1555
rect 56340 1525 56345 1555
rect 56305 1520 56345 1525
rect 56365 1505 56395 1575
rect 56420 1695 56450 1760
rect 56470 1750 56510 1755
rect 56470 1720 56475 1750
rect 56505 1720 56510 1750
rect 56470 1715 56510 1720
rect 56420 1575 56425 1695
rect 56445 1575 56450 1695
rect 56420 1560 56450 1575
rect 56475 1695 56505 1715
rect 56475 1575 56480 1695
rect 56500 1575 56505 1695
rect 56415 1555 56455 1560
rect 56415 1525 56420 1555
rect 56450 1525 56455 1555
rect 56415 1520 56455 1525
rect 56475 1505 56505 1575
rect 56530 1695 56560 1760
rect 56580 1750 56620 1755
rect 56580 1720 56585 1750
rect 56615 1720 56620 1750
rect 56580 1715 56620 1720
rect 56530 1575 56535 1695
rect 56555 1575 56560 1695
rect 56530 1560 56560 1575
rect 56585 1695 56615 1715
rect 56585 1575 56590 1695
rect 56610 1575 56615 1695
rect 56525 1555 56565 1560
rect 56525 1525 56530 1555
rect 56560 1525 56565 1555
rect 56525 1520 56565 1525
rect 56585 1505 56615 1575
rect 56640 1695 56670 1760
rect 56690 1750 56720 1755
rect 56850 1785 56880 1790
rect 56850 1750 56880 1755
rect 56903 1785 56933 1790
rect 56903 1750 56933 1755
rect 56950 1705 56970 1855
rect 57185 1805 57215 1990
rect 57240 1985 57270 2045
rect 57295 2165 57325 2225
rect 57345 2215 57385 2465
rect 57400 2260 57440 2265
rect 57400 2230 57405 2260
rect 57435 2230 57440 2260
rect 57400 2225 57440 2230
rect 57345 2185 57350 2215
rect 57380 2185 57385 2215
rect 57345 2180 57385 2185
rect 57295 2045 57300 2165
rect 57320 2045 57325 2165
rect 57295 2030 57325 2045
rect 57350 2165 57380 2180
rect 57350 2045 57355 2165
rect 57375 2045 57380 2165
rect 57290 2025 57330 2030
rect 57290 1995 57295 2025
rect 57325 1995 57330 2025
rect 57290 1990 57330 1995
rect 57235 1980 57275 1985
rect 57235 1950 57240 1980
rect 57270 1950 57275 1980
rect 57235 1945 57275 1950
rect 57125 1795 57165 1800
rect 57080 1785 57110 1790
rect 57125 1765 57130 1795
rect 57160 1765 57165 1795
rect 57295 1805 57325 1990
rect 57350 1985 57380 2045
rect 57405 2165 57435 2225
rect 57455 2215 57495 2465
rect 57510 2260 57550 2265
rect 57510 2230 57515 2260
rect 57545 2230 57550 2260
rect 57510 2225 57550 2230
rect 57455 2185 57460 2215
rect 57490 2185 57495 2215
rect 57455 2180 57495 2185
rect 57405 2045 57410 2165
rect 57430 2045 57435 2165
rect 57405 2030 57435 2045
rect 57460 2165 57490 2180
rect 57460 2045 57465 2165
rect 57485 2045 57490 2165
rect 57400 2025 57440 2030
rect 57400 1995 57405 2025
rect 57435 1995 57440 2025
rect 57400 1990 57440 1995
rect 57345 1980 57385 1985
rect 57345 1950 57350 1980
rect 57380 1950 57385 1980
rect 57345 1945 57385 1950
rect 57185 1770 57215 1775
rect 57235 1795 57275 1800
rect 57125 1760 57165 1765
rect 57235 1765 57240 1795
rect 57270 1765 57275 1795
rect 57405 1805 57435 1990
rect 57460 1985 57490 2045
rect 57515 2165 57545 2225
rect 57565 2215 57605 2465
rect 57620 2260 57660 2265
rect 57620 2230 57625 2260
rect 57655 2230 57660 2260
rect 57620 2225 57660 2230
rect 57565 2185 57570 2215
rect 57600 2185 57605 2215
rect 57565 2180 57605 2185
rect 57515 2045 57520 2165
rect 57540 2045 57545 2165
rect 57515 2030 57545 2045
rect 57570 2165 57600 2180
rect 57570 2045 57575 2165
rect 57595 2045 57600 2165
rect 57510 2025 57550 2030
rect 57510 1995 57515 2025
rect 57545 1995 57550 2025
rect 57510 1990 57550 1995
rect 57455 1980 57495 1985
rect 57455 1950 57460 1980
rect 57490 1950 57495 1980
rect 57455 1945 57495 1950
rect 57295 1770 57325 1775
rect 57345 1795 57385 1800
rect 57235 1760 57275 1765
rect 57345 1765 57350 1795
rect 57380 1765 57385 1795
rect 57515 1805 57545 1990
rect 57570 1985 57600 2045
rect 57625 2165 57655 2225
rect 57675 2215 57715 2465
rect 57675 2185 57680 2215
rect 57710 2185 57715 2215
rect 57675 2180 57715 2185
rect 57625 2045 57630 2165
rect 57650 2045 57655 2165
rect 57625 2030 57655 2045
rect 57680 2165 57710 2180
rect 57680 2045 57685 2165
rect 57705 2045 57710 2165
rect 57620 2025 57660 2030
rect 57620 1995 57625 2025
rect 57655 1995 57660 2025
rect 57620 1990 57660 1995
rect 57565 1980 57605 1985
rect 57565 1950 57570 1980
rect 57600 1950 57605 1980
rect 57565 1945 57605 1950
rect 57405 1770 57435 1775
rect 57455 1795 57495 1800
rect 57345 1760 57385 1765
rect 57455 1765 57460 1795
rect 57490 1765 57495 1795
rect 57625 1805 57655 1990
rect 57680 1985 57710 2045
rect 57735 2165 57765 2175
rect 57735 2045 57740 2165
rect 57760 2045 57765 2165
rect 57735 2035 57765 2045
rect 57735 2005 57765 2015
rect 57735 1985 57740 2005
rect 57760 1985 57765 2005
rect 57675 1980 57715 1985
rect 57675 1950 57680 1980
rect 57710 1950 57715 1980
rect 57675 1945 57715 1950
rect 57735 1940 57765 1985
rect 57730 1935 57770 1940
rect 57730 1905 57735 1935
rect 57765 1905 57770 1935
rect 57730 1900 57770 1905
rect 57515 1770 57545 1775
rect 57565 1795 57605 1800
rect 57455 1760 57495 1765
rect 57565 1765 57570 1795
rect 57600 1765 57605 1795
rect 57625 1770 57655 1775
rect 57675 1795 57715 1800
rect 57565 1760 57605 1765
rect 57675 1765 57680 1795
rect 57710 1765 57715 1795
rect 57675 1760 57715 1765
rect 57730 1785 57760 1790
rect 57080 1750 57110 1755
rect 56640 1575 56645 1695
rect 56665 1575 56670 1695
rect 56640 1560 56670 1575
rect 56695 1695 56805 1705
rect 56695 1575 56700 1695
rect 56720 1575 56780 1695
rect 56800 1575 56805 1695
rect 56695 1565 56805 1575
rect 56830 1695 56860 1705
rect 56830 1575 56835 1695
rect 56855 1575 56860 1695
rect 56830 1565 56860 1575
rect 56885 1695 56915 1705
rect 56885 1575 56890 1695
rect 56910 1575 56915 1695
rect 56885 1565 56915 1575
rect 56940 1695 56970 1705
rect 56940 1575 56945 1695
rect 56965 1575 56970 1695
rect 56940 1565 56970 1575
rect 56995 1695 57105 1705
rect 56995 1575 57000 1695
rect 57020 1575 57080 1695
rect 57100 1575 57105 1695
rect 56995 1565 57105 1575
rect 57130 1695 57160 1760
rect 57180 1750 57220 1755
rect 57180 1720 57185 1750
rect 57215 1720 57220 1750
rect 57180 1715 57220 1720
rect 57130 1575 57135 1695
rect 57155 1575 57160 1695
rect 56635 1555 56675 1560
rect 56635 1525 56640 1555
rect 56670 1525 56675 1555
rect 56740 1545 56760 1565
rect 56635 1520 56675 1525
rect 56735 1535 56765 1545
rect 56735 1515 56740 1535
rect 56760 1515 56765 1535
rect 56735 1505 56765 1515
rect 56040 1335 56060 1505
rect 56140 1500 56180 1505
rect 56140 1470 56145 1500
rect 56175 1470 56180 1500
rect 56140 1465 56180 1470
rect 56250 1500 56290 1505
rect 56250 1470 56255 1500
rect 56285 1470 56290 1500
rect 56250 1465 56290 1470
rect 56360 1500 56400 1505
rect 56360 1470 56365 1500
rect 56395 1470 56400 1500
rect 56360 1465 56400 1470
rect 56470 1500 56700 1505
rect 56470 1470 56475 1500
rect 56505 1470 56585 1500
rect 56615 1470 56700 1500
rect 56030 1330 56070 1335
rect 56030 1300 56035 1330
rect 56065 1300 56070 1330
rect 56030 1295 56070 1300
rect 55940 1285 55980 1290
rect 55940 1255 55945 1285
rect 55975 1255 55980 1285
rect 55940 1250 55980 1255
rect 56330 1115 56370 1120
rect 56330 1085 56335 1115
rect 56365 1085 56370 1115
rect 56330 1080 56370 1085
rect 56185 995 56255 1005
rect 56185 775 56230 995
rect 56250 775 56255 995
rect 56185 765 56255 775
rect 56225 745 56255 765
rect 56280 995 56310 1005
rect 56280 775 56285 995
rect 56305 775 56310 995
rect 56280 745 56310 775
rect 56335 995 56365 1080
rect 56470 1065 56700 1470
rect 56740 1335 56760 1505
rect 56835 1425 56855 1565
rect 56825 1420 56865 1425
rect 56825 1390 56830 1420
rect 56860 1390 56865 1420
rect 56825 1385 56865 1390
rect 56730 1330 56770 1335
rect 56730 1300 56735 1330
rect 56765 1300 56770 1330
rect 56730 1295 56770 1300
rect 56835 1065 56855 1385
rect 56890 1120 56910 1565
rect 56945 1425 56965 1565
rect 57040 1545 57060 1565
rect 57130 1560 57160 1575
rect 57185 1695 57215 1715
rect 57185 1575 57190 1695
rect 57210 1575 57215 1695
rect 57125 1555 57165 1560
rect 57035 1535 57065 1545
rect 57035 1515 57040 1535
rect 57060 1515 57065 1535
rect 57125 1525 57130 1555
rect 57160 1525 57165 1555
rect 57125 1520 57165 1525
rect 57035 1505 57065 1515
rect 57185 1505 57215 1575
rect 57240 1695 57270 1760
rect 57290 1750 57330 1755
rect 57290 1720 57295 1750
rect 57325 1720 57330 1750
rect 57290 1715 57330 1720
rect 57240 1575 57245 1695
rect 57265 1575 57270 1695
rect 57240 1560 57270 1575
rect 57295 1695 57325 1715
rect 57295 1575 57300 1695
rect 57320 1575 57325 1695
rect 57235 1555 57275 1560
rect 57235 1525 57240 1555
rect 57270 1525 57275 1555
rect 57235 1520 57275 1525
rect 57295 1505 57325 1575
rect 57350 1695 57380 1760
rect 57400 1750 57440 1755
rect 57400 1720 57405 1750
rect 57435 1720 57440 1750
rect 57400 1715 57440 1720
rect 57350 1575 57355 1695
rect 57375 1575 57380 1695
rect 57350 1560 57380 1575
rect 57405 1695 57435 1715
rect 57405 1575 57410 1695
rect 57430 1575 57435 1695
rect 57345 1555 57385 1560
rect 57345 1525 57350 1555
rect 57380 1525 57385 1555
rect 57345 1520 57385 1525
rect 57405 1505 57435 1575
rect 57460 1695 57490 1760
rect 57510 1750 57550 1755
rect 57510 1720 57515 1750
rect 57545 1720 57550 1750
rect 57510 1715 57550 1720
rect 57460 1575 57465 1695
rect 57485 1575 57490 1695
rect 57460 1560 57490 1575
rect 57515 1695 57545 1715
rect 57515 1575 57520 1695
rect 57540 1575 57545 1695
rect 57455 1555 57495 1560
rect 57455 1525 57460 1555
rect 57490 1525 57495 1555
rect 57455 1520 57495 1525
rect 57515 1505 57545 1575
rect 57570 1695 57600 1760
rect 57620 1750 57660 1755
rect 57620 1720 57625 1750
rect 57655 1720 57660 1750
rect 57620 1715 57660 1720
rect 57570 1575 57575 1695
rect 57595 1575 57600 1695
rect 57570 1560 57600 1575
rect 57625 1695 57655 1715
rect 57625 1575 57630 1695
rect 57650 1575 57655 1695
rect 57565 1555 57605 1560
rect 57565 1525 57570 1555
rect 57600 1525 57605 1555
rect 57565 1520 57605 1525
rect 57625 1505 57655 1575
rect 57680 1695 57710 1760
rect 57730 1750 57760 1755
rect 57680 1575 57685 1695
rect 57705 1575 57710 1695
rect 57680 1560 57710 1575
rect 57735 1695 57765 1705
rect 57735 1575 57740 1695
rect 57760 1575 57765 1695
rect 57735 1565 57765 1575
rect 57675 1555 57715 1560
rect 57675 1525 57680 1555
rect 57710 1525 57715 1555
rect 57675 1520 57715 1525
rect 57735 1535 57765 1545
rect 57735 1515 57740 1535
rect 57760 1515 57765 1535
rect 57735 1505 57765 1515
rect 56935 1420 56975 1425
rect 56935 1390 56940 1420
rect 56970 1390 56975 1420
rect 56935 1385 56975 1390
rect 57040 1335 57060 1505
rect 57100 1500 57330 1505
rect 57100 1470 57185 1500
rect 57215 1470 57295 1500
rect 57325 1470 57330 1500
rect 57030 1330 57070 1335
rect 57030 1300 57035 1330
rect 57065 1300 57070 1330
rect 57030 1295 57070 1300
rect 56880 1115 56920 1120
rect 56880 1085 56885 1115
rect 56915 1085 56920 1115
rect 56880 1080 56920 1085
rect 57100 1065 57330 1470
rect 57400 1500 57440 1505
rect 57400 1470 57405 1500
rect 57435 1470 57440 1500
rect 57400 1465 57440 1470
rect 57510 1500 57550 1505
rect 57510 1470 57515 1500
rect 57545 1470 57550 1500
rect 57510 1465 57550 1470
rect 57620 1500 57660 1505
rect 57620 1470 57625 1500
rect 57655 1470 57660 1500
rect 57620 1465 57660 1470
rect 57740 1335 57760 1505
rect 57730 1330 57770 1335
rect 57730 1300 57735 1330
rect 57765 1300 57770 1330
rect 57730 1295 57770 1300
rect 57830 1290 57850 2985
rect 58020 2750 58040 3345
rect 58010 2745 58050 2750
rect 58010 2715 58015 2745
rect 58045 2715 58050 2745
rect 58010 2710 58050 2715
rect 57865 2690 57905 2695
rect 57865 2660 57870 2690
rect 57900 2660 57905 2690
rect 57865 2655 57905 2660
rect 57820 1285 57860 1290
rect 57820 1255 57825 1285
rect 57855 1255 57860 1285
rect 57820 1250 57860 1255
rect 57875 1120 57895 2655
rect 57930 2315 57970 2320
rect 57930 2285 57935 2315
rect 57965 2285 57970 2315
rect 58020 2295 58040 2710
rect 58080 2580 58200 3405
rect 59155 3400 59195 3405
rect 58280 3380 58320 3385
rect 58280 3350 58285 3380
rect 58315 3350 58320 3380
rect 58280 3345 58320 3350
rect 58390 3380 58430 3385
rect 58390 3350 58395 3380
rect 58425 3350 58430 3380
rect 58390 3345 58430 3350
rect 58500 3380 58540 3385
rect 58500 3350 58505 3380
rect 58535 3350 58540 3380
rect 58500 3345 58540 3350
rect 58610 3380 58650 3385
rect 58610 3350 58615 3380
rect 58645 3350 58650 3380
rect 58610 3345 58650 3350
rect 58720 3380 58760 3385
rect 58720 3350 58725 3380
rect 58755 3350 58760 3380
rect 58720 3345 58760 3350
rect 58830 3380 58870 3385
rect 58830 3350 58835 3380
rect 58865 3350 58870 3380
rect 58830 3345 58870 3350
rect 58940 3380 58980 3385
rect 58940 3350 58945 3380
rect 58975 3350 58980 3380
rect 59155 3370 59160 3400
rect 59190 3370 59195 3400
rect 59155 3365 59195 3370
rect 58940 3345 58980 3350
rect 58285 3310 58315 3345
rect 58285 3290 58290 3310
rect 58310 3290 58315 3310
rect 58285 3250 58315 3290
rect 58335 3300 58375 3305
rect 58335 3270 58340 3300
rect 58370 3270 58375 3300
rect 58335 3265 58375 3270
rect 58285 2680 58290 3250
rect 58310 2680 58315 3250
rect 58285 2670 58315 2680
rect 58340 3250 58370 3265
rect 58340 2680 58345 3250
rect 58365 2680 58370 3250
rect 58340 2665 58370 2680
rect 58395 3250 58425 3345
rect 58445 3300 58485 3305
rect 58445 3270 58450 3300
rect 58480 3270 58485 3300
rect 58445 3265 58485 3270
rect 58395 2680 58400 3250
rect 58420 2680 58425 3250
rect 58395 2670 58425 2680
rect 58450 3250 58480 3265
rect 58450 2680 58455 3250
rect 58475 2680 58480 3250
rect 58450 2665 58480 2680
rect 58505 3250 58535 3345
rect 58555 3300 58595 3305
rect 58555 3270 58560 3300
rect 58590 3270 58595 3300
rect 58555 3265 58595 3270
rect 58505 2680 58510 3250
rect 58530 2680 58535 3250
rect 58505 2670 58535 2680
rect 58560 3250 58590 3265
rect 58560 2680 58565 3250
rect 58585 2680 58590 3250
rect 58560 2665 58590 2680
rect 58615 3250 58645 3345
rect 58665 3300 58705 3305
rect 58665 3270 58670 3300
rect 58700 3270 58705 3300
rect 58665 3265 58705 3270
rect 58615 2680 58620 3250
rect 58640 2680 58645 3250
rect 58615 2670 58645 2680
rect 58670 3250 58700 3265
rect 58670 2680 58675 3250
rect 58695 2680 58700 3250
rect 58670 2665 58700 2680
rect 58725 3250 58755 3345
rect 58775 3300 58815 3305
rect 58775 3270 58780 3300
rect 58810 3270 58815 3300
rect 58775 3265 58815 3270
rect 58725 2680 58730 3250
rect 58750 2680 58755 3250
rect 58725 2670 58755 2680
rect 58780 3250 58810 3265
rect 58780 2680 58785 3250
rect 58805 2680 58810 3250
rect 58780 2665 58810 2680
rect 58835 3250 58865 3345
rect 58945 3310 58975 3345
rect 59165 3325 59185 3365
rect 58885 3300 58925 3305
rect 58885 3270 58890 3300
rect 58920 3270 58925 3300
rect 58885 3265 58925 3270
rect 58945 3290 58950 3310
rect 58970 3290 58975 3310
rect 58835 2680 58840 3250
rect 58860 2680 58865 3250
rect 58835 2670 58865 2680
rect 58890 3250 58920 3265
rect 58890 2680 58895 3250
rect 58915 2680 58920 3250
rect 58890 2665 58920 2680
rect 58945 3250 58975 3290
rect 59105 3315 59246 3325
rect 59105 3295 59110 3315
rect 59130 3295 59165 3315
rect 59185 3295 59220 3315
rect 59240 3295 59246 3315
rect 59105 3285 59246 3295
rect 58945 2680 58950 3250
rect 58970 2680 58975 3250
rect 59105 2710 59246 2720
rect 59105 2690 59110 2710
rect 59130 2690 59165 2710
rect 59185 2690 59220 2710
rect 59240 2690 59246 2710
rect 59105 2680 59246 2690
rect 58945 2670 58975 2680
rect 58080 2550 58085 2580
rect 58115 2550 58125 2580
rect 58155 2550 58165 2580
rect 58195 2550 58200 2580
rect 58080 2540 58200 2550
rect 58080 2510 58085 2540
rect 58115 2510 58125 2540
rect 58155 2510 58165 2540
rect 58195 2510 58200 2540
rect 58080 2500 58200 2510
rect 58080 2470 58085 2500
rect 58115 2470 58125 2500
rect 58155 2470 58165 2500
rect 58195 2470 58200 2500
rect 57930 2280 57970 2285
rect 58010 2290 58050 2295
rect 57940 1940 57960 2280
rect 58010 2260 58015 2290
rect 58045 2260 58050 2290
rect 58010 2255 58050 2260
rect 57930 1935 57970 1940
rect 57930 1905 57935 1935
rect 57965 1905 57970 1935
rect 57930 1900 57970 1905
rect 57940 1335 57960 1900
rect 58020 1380 58040 2255
rect 58080 1880 58200 2470
rect 58335 2660 58375 2665
rect 58335 2630 58340 2660
rect 58370 2630 58375 2660
rect 58335 2435 58375 2630
rect 58445 2660 58485 2665
rect 58445 2630 58450 2660
rect 58480 2630 58485 2660
rect 58445 2435 58485 2630
rect 58555 2660 58595 2665
rect 58555 2630 58560 2660
rect 58590 2630 58595 2660
rect 58555 2435 58595 2630
rect 58665 2660 58705 2665
rect 58665 2630 58670 2660
rect 58700 2630 58705 2660
rect 58610 2580 58650 2585
rect 58610 2550 58615 2580
rect 58645 2550 58650 2580
rect 58610 2540 58650 2550
rect 58610 2510 58615 2540
rect 58645 2510 58650 2540
rect 58610 2500 58650 2510
rect 58610 2470 58615 2500
rect 58645 2470 58650 2500
rect 58610 2465 58650 2470
rect 58665 2435 58705 2630
rect 58775 2660 58815 2665
rect 58775 2630 58780 2660
rect 58810 2630 58815 2660
rect 58775 2435 58815 2630
rect 58885 2660 58925 2665
rect 58885 2630 58890 2660
rect 58920 2630 58925 2660
rect 58885 2435 58925 2630
rect 59115 2580 59235 2680
rect 59115 2550 59120 2580
rect 59150 2550 59160 2580
rect 59190 2550 59200 2580
rect 59230 2550 59235 2580
rect 59115 2540 59235 2550
rect 59115 2510 59120 2540
rect 59150 2510 59160 2540
rect 59190 2510 59200 2540
rect 59230 2510 59235 2540
rect 59115 2500 59235 2510
rect 59115 2470 59120 2500
rect 59150 2470 59160 2500
rect 59190 2470 59200 2500
rect 59230 2470 59235 2500
rect 59115 2465 59235 2470
rect 58335 2430 58925 2435
rect 58335 2400 58340 2430
rect 58370 2400 58395 2430
rect 58425 2400 58450 2430
rect 58480 2400 58505 2430
rect 58535 2400 58560 2430
rect 58590 2400 58615 2430
rect 58645 2400 58670 2430
rect 58700 2400 58725 2430
rect 58755 2400 58780 2430
rect 58810 2400 58835 2430
rect 58865 2400 58890 2430
rect 58920 2400 58925 2430
rect 58335 2390 58925 2400
rect 58335 2360 58340 2390
rect 58370 2360 58395 2390
rect 58425 2360 58450 2390
rect 58480 2360 58505 2390
rect 58535 2360 58560 2390
rect 58590 2360 58615 2390
rect 58645 2360 58670 2390
rect 58700 2360 58725 2390
rect 58755 2360 58780 2390
rect 58810 2360 58835 2390
rect 58865 2360 58890 2390
rect 58920 2360 58925 2390
rect 58335 2350 58925 2360
rect 58335 2320 58340 2350
rect 58370 2320 58395 2350
rect 58425 2320 58450 2350
rect 58480 2320 58505 2350
rect 58535 2320 58560 2350
rect 58590 2320 58615 2350
rect 58645 2320 58670 2350
rect 58700 2320 58725 2350
rect 58755 2320 58780 2350
rect 58810 2320 58835 2350
rect 58865 2320 58890 2350
rect 58920 2320 58925 2350
rect 58335 2315 58925 2320
rect 59365 2430 59615 2435
rect 59365 2400 59370 2430
rect 59400 2400 59410 2430
rect 59440 2400 59455 2430
rect 59485 2400 59495 2430
rect 59525 2400 59540 2430
rect 59570 2400 59580 2430
rect 59610 2400 59615 2430
rect 59365 2390 59615 2400
rect 59365 2360 59370 2390
rect 59400 2360 59410 2390
rect 59440 2360 59455 2390
rect 59485 2360 59495 2390
rect 59525 2360 59540 2390
rect 59570 2360 59580 2390
rect 59610 2360 59615 2390
rect 59365 2350 59615 2360
rect 59365 2320 59370 2350
rect 59400 2320 59410 2350
rect 59440 2320 59455 2350
rect 59485 2320 59495 2350
rect 59525 2320 59540 2350
rect 59570 2320 59580 2350
rect 59610 2320 59615 2350
rect 58280 2290 58320 2295
rect 58280 2260 58285 2290
rect 58315 2260 58320 2290
rect 58280 2255 58320 2260
rect 58940 2290 58980 2295
rect 58940 2260 58945 2290
rect 58975 2260 58980 2290
rect 58940 2255 58980 2260
rect 58285 2210 58315 2255
rect 58335 2245 58375 2250
rect 58335 2215 58340 2245
rect 58370 2215 58375 2245
rect 58335 2210 58375 2215
rect 58445 2245 58485 2250
rect 58445 2215 58450 2245
rect 58480 2215 58485 2245
rect 58445 2210 58485 2215
rect 58555 2245 58595 2250
rect 58555 2215 58560 2245
rect 58590 2215 58595 2245
rect 58555 2210 58595 2215
rect 58665 2245 58705 2250
rect 58665 2215 58670 2245
rect 58700 2215 58705 2245
rect 58665 2210 58705 2215
rect 58775 2245 58815 2250
rect 58775 2215 58780 2245
rect 58810 2215 58815 2245
rect 58775 2210 58815 2215
rect 58885 2245 58925 2250
rect 58885 2215 58890 2245
rect 58920 2215 58925 2245
rect 58885 2210 58925 2215
rect 58945 2210 58975 2255
rect 58285 2190 58290 2210
rect 58310 2190 58315 2210
rect 58285 2150 58315 2190
rect 58285 1980 58290 2150
rect 58310 1980 58315 2150
rect 58285 1970 58315 1980
rect 58340 2150 58370 2210
rect 58390 2200 58430 2205
rect 58390 2170 58395 2200
rect 58425 2170 58430 2200
rect 58390 2165 58430 2170
rect 58340 1980 58345 2150
rect 58365 1980 58370 2150
rect 58340 1970 58370 1980
rect 58395 2150 58425 2165
rect 58395 1980 58400 2150
rect 58420 1980 58425 2150
rect 58395 1950 58425 1980
rect 58450 2150 58480 2210
rect 58500 2200 58540 2205
rect 58500 2170 58505 2200
rect 58535 2170 58540 2200
rect 58500 2165 58540 2170
rect 58450 1980 58455 2150
rect 58475 1980 58480 2150
rect 58450 1970 58480 1980
rect 58505 2150 58535 2165
rect 58505 1980 58510 2150
rect 58530 1980 58535 2150
rect 58505 1950 58535 1980
rect 58560 2150 58590 2210
rect 58610 2200 58650 2205
rect 58610 2170 58615 2200
rect 58645 2170 58650 2200
rect 58610 2165 58650 2170
rect 58560 1980 58565 2150
rect 58585 1980 58590 2150
rect 58560 1970 58590 1980
rect 58615 2150 58645 2165
rect 58615 1980 58620 2150
rect 58640 1980 58645 2150
rect 58615 1950 58645 1980
rect 58670 2150 58700 2210
rect 58720 2200 58760 2205
rect 58720 2170 58725 2200
rect 58755 2170 58760 2200
rect 58720 2165 58760 2170
rect 58670 1980 58675 2150
rect 58695 1980 58700 2150
rect 58670 1970 58700 1980
rect 58725 2150 58755 2165
rect 58725 1980 58730 2150
rect 58750 1980 58755 2150
rect 58725 1950 58755 1980
rect 58780 2150 58810 2210
rect 58830 2200 58870 2205
rect 58830 2170 58835 2200
rect 58865 2170 58870 2200
rect 58830 2165 58870 2170
rect 58780 1980 58785 2150
rect 58805 1980 58810 2150
rect 58780 1970 58810 1980
rect 58835 2150 58865 2165
rect 58835 1980 58840 2150
rect 58860 1980 58865 2150
rect 58835 1950 58865 1980
rect 58890 2150 58920 2210
rect 58890 1980 58895 2150
rect 58915 1980 58920 2150
rect 58890 1970 58920 1980
rect 58945 2190 58950 2210
rect 58970 2190 58975 2210
rect 58945 2150 58975 2190
rect 58945 1980 58950 2150
rect 58970 1980 58975 2150
rect 58945 1970 58975 1980
rect 58390 1945 58430 1950
rect 58390 1915 58395 1945
rect 58425 1915 58430 1945
rect 58390 1910 58430 1915
rect 58500 1945 58540 1950
rect 58500 1915 58505 1945
rect 58535 1915 58540 1945
rect 58500 1910 58540 1915
rect 58610 1945 58650 1950
rect 58610 1915 58615 1945
rect 58645 1915 58650 1945
rect 58610 1910 58650 1915
rect 58720 1945 58760 1950
rect 58720 1915 58725 1945
rect 58755 1915 58760 1945
rect 58720 1910 58760 1915
rect 58830 1945 58870 1950
rect 58830 1915 58835 1945
rect 58865 1915 58870 1945
rect 58830 1910 58870 1915
rect 59080 1945 59120 1950
rect 59080 1915 59085 1945
rect 59115 1915 59120 1945
rect 59080 1910 59120 1915
rect 58080 1850 58085 1880
rect 58115 1850 58125 1880
rect 58155 1850 58165 1880
rect 58195 1850 58200 1880
rect 58080 1840 58200 1850
rect 58080 1810 58085 1840
rect 58115 1810 58125 1840
rect 58155 1810 58165 1840
rect 58195 1810 58200 1840
rect 58080 1805 58200 1810
rect 58445 1880 58485 1885
rect 58445 1850 58450 1880
rect 58480 1850 58485 1880
rect 58445 1840 58485 1850
rect 58445 1810 58450 1840
rect 58480 1810 58485 1840
rect 58445 1805 58485 1810
rect 58390 1760 58430 1765
rect 58390 1730 58395 1760
rect 58425 1730 58430 1760
rect 58390 1725 58430 1730
rect 58500 1760 58540 1765
rect 58500 1730 58505 1760
rect 58535 1730 58540 1760
rect 58500 1725 58540 1730
rect 58610 1760 58650 1765
rect 58610 1730 58615 1760
rect 58645 1730 58650 1760
rect 58610 1725 58650 1730
rect 58720 1760 58760 1765
rect 58720 1730 58725 1760
rect 58755 1730 58760 1760
rect 58720 1725 58760 1730
rect 58830 1760 58870 1765
rect 58830 1730 58835 1760
rect 58865 1730 58870 1760
rect 58830 1725 58870 1730
rect 59035 1760 59075 1765
rect 59035 1730 59040 1760
rect 59070 1730 59075 1760
rect 59035 1725 59075 1730
rect 58285 1710 58315 1720
rect 58285 1440 58290 1710
rect 58310 1440 58315 1710
rect 58285 1400 58315 1440
rect 58285 1380 58290 1400
rect 58310 1380 58315 1400
rect 58340 1710 58370 1720
rect 58340 1440 58345 1710
rect 58365 1440 58370 1710
rect 58340 1380 58370 1440
rect 58395 1710 58425 1725
rect 58395 1440 58400 1710
rect 58420 1440 58425 1710
rect 58395 1425 58425 1440
rect 58450 1710 58480 1720
rect 58450 1440 58455 1710
rect 58475 1440 58480 1710
rect 58390 1420 58430 1425
rect 58390 1390 58395 1420
rect 58425 1390 58430 1420
rect 58390 1385 58430 1390
rect 58450 1380 58480 1440
rect 58505 1710 58535 1725
rect 58505 1440 58510 1710
rect 58530 1440 58535 1710
rect 58505 1425 58535 1440
rect 58560 1710 58590 1720
rect 58560 1440 58565 1710
rect 58585 1440 58590 1710
rect 58500 1420 58540 1425
rect 58500 1390 58505 1420
rect 58535 1390 58540 1420
rect 58500 1385 58540 1390
rect 58560 1380 58590 1440
rect 58615 1710 58645 1725
rect 58615 1440 58620 1710
rect 58640 1440 58645 1710
rect 58615 1425 58645 1440
rect 58670 1710 58700 1720
rect 58670 1440 58675 1710
rect 58695 1440 58700 1710
rect 58610 1420 58650 1425
rect 58610 1390 58615 1420
rect 58645 1390 58650 1420
rect 58610 1385 58650 1390
rect 58670 1380 58700 1440
rect 58725 1710 58755 1725
rect 58725 1440 58730 1710
rect 58750 1440 58755 1710
rect 58725 1425 58755 1440
rect 58780 1710 58810 1720
rect 58780 1440 58785 1710
rect 58805 1440 58810 1710
rect 58720 1420 58760 1425
rect 58720 1390 58725 1420
rect 58755 1390 58760 1420
rect 58720 1385 58760 1390
rect 58780 1380 58810 1440
rect 58835 1710 58865 1725
rect 58835 1440 58840 1710
rect 58860 1440 58865 1710
rect 58835 1425 58865 1440
rect 58890 1710 58920 1720
rect 58890 1440 58895 1710
rect 58915 1440 58920 1710
rect 58830 1420 58870 1425
rect 58830 1390 58835 1420
rect 58865 1390 58870 1420
rect 58830 1385 58870 1390
rect 58890 1380 58920 1440
rect 58945 1710 58975 1720
rect 58945 1440 58950 1710
rect 58970 1440 58975 1710
rect 58945 1400 58975 1440
rect 58945 1380 58950 1400
rect 58970 1380 58975 1400
rect 59045 1395 59065 1725
rect 58010 1375 58050 1380
rect 58010 1345 58015 1375
rect 58045 1345 58050 1375
rect 58010 1340 58050 1345
rect 58285 1335 58315 1380
rect 58335 1375 58375 1380
rect 58335 1345 58340 1375
rect 58370 1345 58375 1375
rect 58335 1340 58375 1345
rect 58445 1375 58485 1380
rect 58445 1345 58450 1375
rect 58480 1345 58485 1375
rect 58445 1340 58485 1345
rect 58555 1375 58595 1380
rect 58555 1345 58560 1375
rect 58590 1345 58595 1375
rect 58555 1340 58595 1345
rect 58665 1375 58705 1380
rect 58665 1345 58670 1375
rect 58700 1345 58705 1375
rect 58665 1340 58705 1345
rect 58775 1375 58815 1380
rect 58775 1345 58780 1375
rect 58810 1345 58815 1375
rect 58775 1340 58815 1345
rect 58885 1375 58925 1380
rect 58885 1345 58890 1375
rect 58920 1345 58925 1375
rect 58885 1340 58925 1345
rect 58945 1335 58975 1380
rect 59035 1390 59075 1395
rect 59035 1360 59040 1390
rect 59070 1360 59075 1390
rect 59035 1355 59075 1360
rect 59090 1340 59110 1910
rect 59365 1710 59615 2320
rect 59645 2245 59685 2250
rect 59645 2215 59650 2245
rect 59680 2215 59685 2245
rect 59645 2210 59685 2215
rect 59365 1680 59375 1710
rect 59405 1680 59425 1710
rect 59455 1680 59475 1710
rect 59505 1680 59525 1710
rect 59555 1680 59575 1710
rect 59605 1680 59615 1710
rect 59365 1660 59615 1680
rect 59365 1630 59375 1660
rect 59405 1630 59425 1660
rect 59455 1630 59475 1660
rect 59505 1630 59525 1660
rect 59555 1630 59575 1660
rect 59605 1630 59615 1660
rect 59365 1610 59615 1630
rect 59365 1580 59375 1610
rect 59405 1580 59425 1610
rect 59455 1580 59475 1610
rect 59505 1580 59525 1610
rect 59555 1580 59575 1610
rect 59605 1580 59615 1610
rect 59125 1395 59160 1400
rect 59125 1355 59160 1360
rect 59185 1395 59220 1400
rect 59185 1355 59220 1360
rect 59245 1395 59280 1400
rect 59245 1355 59280 1360
rect 59305 1395 59340 1401
rect 59305 1355 59340 1360
rect 59190 1340 59210 1355
rect 59080 1335 59120 1340
rect 57930 1330 57970 1335
rect 57930 1300 57935 1330
rect 57965 1300 57970 1330
rect 57930 1295 57970 1300
rect 58280 1330 58320 1335
rect 58280 1300 58285 1330
rect 58315 1300 58320 1330
rect 58280 1295 58320 1300
rect 58940 1330 58980 1335
rect 58940 1300 58945 1330
rect 58975 1300 58980 1330
rect 59080 1305 59085 1335
rect 59115 1305 59120 1335
rect 59080 1300 59120 1305
rect 59180 1335 59220 1340
rect 59180 1305 59185 1335
rect 59215 1305 59220 1335
rect 59180 1300 59220 1305
rect 58940 1295 58980 1300
rect 57390 1115 57430 1120
rect 57390 1085 57395 1115
rect 57425 1085 57430 1115
rect 57390 1080 57430 1085
rect 57865 1115 57905 1120
rect 57865 1085 57870 1115
rect 57900 1085 57905 1115
rect 57865 1080 57905 1085
rect 56440 1060 56700 1065
rect 56440 1030 56445 1060
rect 56475 1030 56555 1060
rect 56585 1030 56665 1060
rect 56695 1030 56700 1060
rect 56440 1025 56700 1030
rect 56770 1060 56810 1065
rect 56770 1030 56775 1060
rect 56805 1030 56810 1060
rect 56770 1025 56810 1030
rect 56830 1055 56860 1065
rect 56830 1035 56835 1055
rect 56855 1035 56860 1055
rect 56830 1025 56860 1035
rect 56880 1060 56920 1065
rect 56880 1030 56885 1060
rect 56915 1030 56920 1060
rect 56880 1025 56920 1030
rect 56990 1060 57030 1065
rect 56990 1030 56995 1060
rect 57025 1030 57030 1060
rect 56990 1025 57030 1030
rect 57100 1060 57360 1065
rect 57100 1030 57105 1060
rect 57135 1030 57215 1060
rect 57245 1030 57325 1060
rect 57355 1030 57360 1060
rect 57100 1025 57360 1030
rect 57430 1060 57470 1065
rect 57430 1030 57435 1060
rect 57465 1030 57470 1060
rect 57430 1025 57470 1030
rect 56335 775 56340 995
rect 56360 775 56365 995
rect 56335 765 56365 775
rect 56390 995 56420 1005
rect 56390 775 56395 995
rect 56415 775 56420 995
rect 56390 745 56420 775
rect 56445 995 56475 1025
rect 56445 775 56450 995
rect 56470 775 56475 995
rect 56220 740 56260 745
rect 56220 710 56225 740
rect 56255 710 56260 740
rect 56220 705 56260 710
rect 56275 740 56315 745
rect 56275 710 56280 740
rect 56310 710 56315 740
rect 56275 705 56315 710
rect 56385 740 56425 745
rect 56385 710 56390 740
rect 56420 710 56425 740
rect 56385 705 56425 710
rect 56445 700 56475 775
rect 56500 995 56530 1005
rect 56500 775 56505 995
rect 56525 775 56530 995
rect 56500 745 56530 775
rect 56555 995 56585 1025
rect 56555 775 56560 995
rect 56580 775 56585 995
rect 56495 740 56535 745
rect 56495 710 56500 740
rect 56530 710 56535 740
rect 56495 705 56535 710
rect 56555 700 56585 775
rect 56610 995 56640 1005
rect 56610 775 56615 995
rect 56635 775 56640 995
rect 56610 745 56640 775
rect 56665 995 56695 1025
rect 56665 775 56670 995
rect 56690 775 56695 995
rect 56605 740 56645 745
rect 56605 710 56610 740
rect 56640 710 56645 740
rect 56605 705 56645 710
rect 56665 700 56695 775
rect 56720 995 56750 1005
rect 56720 775 56725 995
rect 56745 775 56750 995
rect 56720 745 56750 775
rect 56775 995 56805 1025
rect 56775 775 56780 995
rect 56800 775 56805 995
rect 56715 740 56755 745
rect 56715 710 56720 740
rect 56750 710 56755 740
rect 56715 705 56755 710
rect 56775 700 56805 775
rect 56830 995 56860 1005
rect 56830 775 56835 995
rect 56855 775 56860 995
rect 56830 745 56860 775
rect 56885 995 56915 1025
rect 56885 775 56890 995
rect 56910 775 56915 995
rect 56825 740 56865 745
rect 56825 710 56830 740
rect 56860 710 56865 740
rect 56825 705 56865 710
rect 56885 700 56915 775
rect 56940 995 56970 1005
rect 56940 775 56945 995
rect 56965 775 56970 995
rect 56940 745 56970 775
rect 56995 995 57025 1025
rect 56995 775 57000 995
rect 57020 775 57025 995
rect 56935 740 56975 745
rect 56935 710 56940 740
rect 56970 710 56975 740
rect 56935 705 56975 710
rect 56995 700 57025 775
rect 57050 995 57080 1005
rect 57050 775 57055 995
rect 57075 775 57080 995
rect 57050 745 57080 775
rect 57105 995 57135 1025
rect 57105 775 57110 995
rect 57130 775 57135 995
rect 57045 740 57085 745
rect 57045 710 57050 740
rect 57080 710 57085 740
rect 57045 705 57085 710
rect 57105 700 57135 775
rect 57160 995 57190 1005
rect 57160 775 57165 995
rect 57185 775 57190 995
rect 57160 745 57190 775
rect 57215 995 57245 1025
rect 57215 775 57220 995
rect 57240 775 57245 995
rect 57155 740 57195 745
rect 57155 710 57160 740
rect 57190 710 57195 740
rect 57155 705 57195 710
rect 57215 700 57245 775
rect 57270 995 57300 1005
rect 57270 775 57275 995
rect 57295 775 57300 995
rect 57270 745 57300 775
rect 57325 995 57355 1025
rect 57325 775 57330 995
rect 57350 775 57355 995
rect 57265 740 57305 745
rect 57265 710 57270 740
rect 57300 710 57305 740
rect 57265 705 57305 710
rect 57325 700 57355 775
rect 57380 995 57410 1005
rect 57380 775 57385 995
rect 57405 775 57410 995
rect 57380 745 57410 775
rect 57435 995 57465 1025
rect 57435 775 57440 995
rect 57460 775 57465 995
rect 57375 740 57415 745
rect 57375 710 57380 740
rect 57410 710 57415 740
rect 57375 705 57415 710
rect 57435 700 57465 775
rect 57490 995 57520 1005
rect 57490 775 57495 995
rect 57515 775 57520 995
rect 57490 745 57520 775
rect 57940 745 57960 1295
rect 59310 1290 59330 1355
rect 59300 1285 59340 1290
rect 59300 1255 59305 1285
rect 59335 1255 59340 1285
rect 59300 1250 59340 1255
rect 58580 1240 58620 1245
rect 58580 1210 58585 1240
rect 58615 1210 58620 1240
rect 58580 1205 58620 1210
rect 59165 1240 59205 1245
rect 59165 1210 59170 1240
rect 59200 1210 59205 1240
rect 59165 1205 59205 1210
rect 58430 1185 58870 1190
rect 58430 1155 58435 1185
rect 58465 1155 58475 1185
rect 58505 1155 58515 1185
rect 58545 1155 58555 1185
rect 58585 1155 58595 1185
rect 58625 1155 58635 1185
rect 58665 1155 58675 1185
rect 58705 1155 58715 1185
rect 58745 1155 58755 1185
rect 58785 1155 58795 1185
rect 58825 1155 58835 1185
rect 58865 1155 58870 1185
rect 58430 1145 58870 1155
rect 58430 1115 58435 1145
rect 58465 1115 58475 1145
rect 58505 1115 58515 1145
rect 58545 1115 58555 1145
rect 58585 1115 58595 1145
rect 58625 1115 58635 1145
rect 58665 1115 58675 1145
rect 58705 1115 58715 1145
rect 58745 1115 58755 1145
rect 58785 1115 58795 1145
rect 58825 1115 58835 1145
rect 58865 1115 58870 1145
rect 58430 1105 58870 1115
rect 58430 1075 58435 1105
rect 58465 1075 58475 1105
rect 58505 1075 58515 1105
rect 58545 1075 58555 1105
rect 58585 1075 58595 1105
rect 58625 1075 58635 1105
rect 58665 1075 58675 1105
rect 58705 1075 58715 1105
rect 58745 1075 58755 1105
rect 58785 1075 58795 1105
rect 58825 1075 58835 1105
rect 58865 1075 58870 1105
rect 58430 1070 58870 1075
rect 59100 1185 59140 1190
rect 59100 1155 59105 1185
rect 59135 1155 59140 1185
rect 59100 1145 59140 1155
rect 59100 1115 59105 1145
rect 59135 1115 59140 1145
rect 59100 1105 59140 1115
rect 59100 1075 59105 1105
rect 59135 1075 59140 1105
rect 59100 1070 59140 1075
rect 58335 1040 58365 1050
rect 57485 740 57525 745
rect 57485 710 57490 740
rect 57520 710 57525 740
rect 57485 705 57525 710
rect 57930 740 57970 745
rect 57930 710 57935 740
rect 57965 710 57970 740
rect 57930 705 57970 710
rect 56440 695 56480 700
rect 56440 665 56445 695
rect 56475 665 56480 695
rect 56440 660 56480 665
rect 56550 695 56590 700
rect 56550 665 56555 695
rect 56585 665 56590 695
rect 56550 660 56590 665
rect 56660 695 56700 700
rect 56660 665 56665 695
rect 56695 665 56700 695
rect 56660 660 56700 665
rect 56770 695 56810 700
rect 56770 665 56775 695
rect 56805 665 56810 695
rect 56770 660 56810 665
rect 56880 695 56920 700
rect 56880 665 56885 695
rect 56915 665 56920 695
rect 56880 660 56920 665
rect 56990 695 57030 700
rect 56990 665 56995 695
rect 57025 665 57030 695
rect 56990 660 57030 665
rect 57100 695 57140 700
rect 57100 665 57105 695
rect 57135 665 57140 695
rect 57100 660 57140 665
rect 57210 695 57250 700
rect 57210 665 57215 695
rect 57245 665 57250 695
rect 57210 660 57250 665
rect 57320 695 57360 700
rect 57320 665 57325 695
rect 57355 665 57360 695
rect 57320 660 57360 665
rect 57430 695 57470 700
rect 57430 665 57435 695
rect 57465 665 57470 695
rect 57430 660 57470 665
rect 56540 640 56580 645
rect 56540 610 56545 640
rect 56575 610 56580 640
rect 56540 605 56580 610
rect 56650 640 56690 645
rect 56650 610 56655 640
rect 56685 610 56690 640
rect 56650 605 56690 610
rect 56870 640 56910 645
rect 56870 610 56875 640
rect 56905 610 56910 640
rect 56870 605 56910 610
rect 55895 595 55935 600
rect 55895 565 55900 595
rect 55930 565 55935 595
rect 55895 560 55935 565
rect 56485 595 56525 600
rect 56485 565 56490 595
rect 56520 565 56525 595
rect 56485 560 56525 565
rect 56395 530 56465 540
rect 56395 410 56440 530
rect 56460 410 56465 530
rect 56395 400 56465 410
rect 56435 370 56465 400
rect 56435 350 56440 370
rect 56460 350 56465 370
rect 56490 530 56520 560
rect 56490 410 56495 530
rect 56515 410 56520 530
rect 56490 350 56520 410
rect 56545 530 56575 605
rect 56595 595 56635 600
rect 56595 565 56600 595
rect 56630 565 56635 595
rect 56595 560 56635 565
rect 56545 410 56550 530
rect 56570 410 56575 530
rect 56545 395 56575 410
rect 56600 530 56630 560
rect 56600 410 56605 530
rect 56625 410 56630 530
rect 56540 390 56580 395
rect 56540 360 56545 390
rect 56575 360 56580 390
rect 56540 355 56580 360
rect 56600 350 56630 410
rect 56655 530 56685 605
rect 56705 595 56745 600
rect 56705 565 56710 595
rect 56740 565 56745 595
rect 56705 560 56745 565
rect 56655 410 56660 530
rect 56680 410 56685 530
rect 56655 395 56685 410
rect 56710 530 56740 560
rect 56710 410 56715 530
rect 56735 410 56740 530
rect 56650 390 56690 395
rect 56650 360 56655 390
rect 56685 360 56690 390
rect 56650 355 56690 360
rect 56710 350 56740 410
rect 56765 530 56835 540
rect 56765 410 56770 530
rect 56790 410 56835 530
rect 56765 400 56835 410
rect 56875 530 56905 605
rect 57040 595 57080 600
rect 57040 565 57045 595
rect 57075 565 57080 595
rect 57040 560 57080 565
rect 56875 410 56880 530
rect 56900 410 56905 530
rect 56765 370 56795 400
rect 56875 395 56905 410
rect 57215 530 57245 660
rect 57215 410 57220 530
rect 57240 410 57245 530
rect 57215 400 57245 410
rect 56765 350 56770 370
rect 56790 350 56795 370
rect 56870 390 56910 395
rect 56870 360 56875 390
rect 56905 360 56910 390
rect 56870 355 56910 360
rect 56435 50 56465 350
rect 56485 345 56525 350
rect 56485 315 56490 345
rect 56520 315 56525 345
rect 56595 345 56635 350
rect 56595 315 56600 345
rect 56630 315 56635 345
rect 56705 345 56745 350
rect 56705 315 56710 345
rect 56740 315 56745 345
rect 56765 50 56795 350
rect 57940 50 57960 705
rect 58335 370 58340 1040
rect 58360 370 58365 1040
rect 58335 330 58365 370
rect 58435 1040 58465 1070
rect 58435 370 58440 1040
rect 58460 370 58465 1040
rect 58435 355 58465 370
rect 58535 1040 58565 1050
rect 58535 370 58540 1040
rect 58560 370 58565 1040
rect 58335 310 58340 330
rect 58360 310 58365 330
rect 58430 350 58470 355
rect 58430 320 58435 350
rect 58465 320 58470 350
rect 58430 315 58470 320
rect 58335 50 58365 310
rect 58535 50 58565 370
rect 58635 1040 58665 1070
rect 58635 370 58640 1040
rect 58660 370 58665 1040
rect 58635 355 58665 370
rect 58735 1040 58765 1050
rect 58735 370 58740 1040
rect 58760 370 58765 1040
rect 58630 350 58670 355
rect 58630 320 58635 350
rect 58665 320 58670 350
rect 58630 315 58670 320
rect 58735 50 58765 370
rect 58835 1040 58865 1070
rect 59105 1050 59140 1070
rect 59175 1055 59195 1205
rect 59365 1185 59615 1580
rect 59365 1155 59370 1185
rect 59400 1155 59410 1185
rect 59440 1155 59455 1185
rect 59485 1155 59495 1185
rect 59525 1155 59540 1185
rect 59570 1155 59580 1185
rect 59610 1155 59615 1185
rect 59365 1145 59615 1155
rect 59365 1115 59370 1145
rect 59400 1115 59410 1145
rect 59440 1115 59455 1145
rect 59485 1115 59495 1145
rect 59525 1115 59540 1145
rect 59570 1115 59580 1145
rect 59610 1115 59615 1145
rect 59365 1105 59615 1115
rect 59365 1075 59370 1105
rect 59400 1075 59410 1105
rect 59440 1075 59455 1105
rect 59485 1075 59495 1105
rect 59525 1075 59540 1105
rect 59570 1075 59580 1105
rect 59610 1075 59615 1105
rect 59365 1070 59615 1075
rect 58835 370 58840 1040
rect 58860 370 58865 1040
rect 58835 355 58865 370
rect 58935 1040 58965 1050
rect 58935 370 58940 1040
rect 58960 370 58965 1040
rect 59105 1010 59140 1015
rect 59165 1050 59200 1055
rect 59165 1010 59200 1015
rect 58830 350 58870 355
rect 58830 320 58835 350
rect 58865 320 58870 350
rect 58830 315 58870 320
rect 58935 330 58965 370
rect 58935 310 58940 330
rect 58960 310 58965 330
rect 58935 50 58965 310
rect 59655 50 59675 2210
rect 52640 45 52760 50
rect 52640 15 52645 45
rect 52675 15 52685 45
rect 52715 15 52725 45
rect 52755 15 52760 45
rect 52640 -800 52760 15
rect 52990 45 53110 50
rect 52990 15 52995 45
rect 53025 15 53035 45
rect 53065 15 53075 45
rect 53105 15 53110 45
rect 52990 -800 53110 15
rect 53340 45 53460 50
rect 53340 15 53345 45
rect 53375 15 53385 45
rect 53415 15 53425 45
rect 53455 15 53460 45
rect 53340 -800 53460 15
rect 53690 45 53810 50
rect 53690 15 53695 45
rect 53725 15 53735 45
rect 53765 15 53775 45
rect 53805 15 53810 45
rect 53690 -800 53810 15
rect 54040 45 54160 50
rect 54040 15 54045 45
rect 54075 15 54085 45
rect 54115 15 54125 45
rect 54155 15 54160 45
rect 54040 -800 54160 15
rect 54390 45 54510 50
rect 54390 15 54395 45
rect 54425 15 54435 45
rect 54465 15 54475 45
rect 54505 15 54510 45
rect 54390 -800 54510 15
rect 54740 45 54865 50
rect 54740 15 54745 45
rect 54775 15 54785 45
rect 54815 15 54825 45
rect 54855 15 54865 45
rect 54740 10 54865 15
rect 55030 45 55070 50
rect 55030 15 55035 45
rect 55065 15 55070 45
rect 55030 10 55070 15
rect 55090 45 55210 50
rect 55090 15 55095 45
rect 55125 15 55135 45
rect 55165 15 55175 45
rect 55205 15 55210 45
rect 54740 -800 54860 10
rect 55090 -800 55210 15
rect 55230 45 55270 50
rect 55230 15 55235 45
rect 55265 15 55270 45
rect 55230 10 55270 15
rect 55435 45 55560 50
rect 55435 15 55445 45
rect 55475 15 55485 45
rect 55515 15 55525 45
rect 55555 15 55560 45
rect 55435 10 55560 15
rect 55440 -800 55560 10
rect 55790 45 55910 50
rect 55790 15 55795 45
rect 55825 15 55835 45
rect 55865 15 55875 45
rect 55905 15 55910 45
rect 55790 -800 55910 15
rect 56140 45 56260 50
rect 56140 15 56145 45
rect 56175 15 56185 45
rect 56215 15 56225 45
rect 56255 15 56260 45
rect 56140 -800 56260 15
rect 56430 45 56470 50
rect 56430 15 56435 45
rect 56465 15 56470 45
rect 56430 10 56470 15
rect 56490 45 56610 50
rect 56490 15 56495 45
rect 56525 15 56535 45
rect 56565 15 56575 45
rect 56605 15 56610 45
rect 56490 -800 56610 15
rect 56760 45 56800 50
rect 56760 15 56765 45
rect 56795 15 56800 45
rect 56760 10 56800 15
rect 56840 45 56960 50
rect 56840 15 56845 45
rect 56875 15 56885 45
rect 56915 15 56925 45
rect 56955 15 56960 45
rect 56840 -800 56960 15
rect 57190 45 57310 50
rect 57190 15 57195 45
rect 57225 15 57235 45
rect 57265 15 57275 45
rect 57305 15 57310 45
rect 57190 -800 57310 15
rect 57540 45 57660 50
rect 57540 15 57545 45
rect 57575 15 57585 45
rect 57615 15 57625 45
rect 57655 15 57660 45
rect 57540 -800 57660 15
rect 57890 45 58010 50
rect 57890 15 57895 45
rect 57925 15 57935 45
rect 57965 15 57975 45
rect 58005 15 58010 45
rect 57890 -800 58010 15
rect 58240 45 58365 50
rect 58240 15 58245 45
rect 58275 15 58285 45
rect 58315 15 58325 45
rect 58355 15 58365 45
rect 58240 10 58365 15
rect 58530 45 58570 50
rect 58530 15 58535 45
rect 58565 15 58570 45
rect 58530 10 58570 15
rect 58590 45 58710 50
rect 58590 15 58595 45
rect 58625 15 58635 45
rect 58665 15 58675 45
rect 58705 15 58710 45
rect 58240 -800 58360 10
rect 58590 -800 58710 15
rect 58730 45 58770 50
rect 58730 15 58735 45
rect 58765 15 58770 45
rect 58730 10 58770 15
rect 58935 45 59060 50
rect 58935 15 58945 45
rect 58975 15 58985 45
rect 59015 15 59025 45
rect 59055 15 59060 45
rect 58935 10 59060 15
rect 58940 -800 59060 10
rect 59290 45 59410 50
rect 59290 15 59295 45
rect 59325 15 59335 45
rect 59365 15 59375 45
rect 59405 15 59410 45
rect 59290 -800 59410 15
rect 59640 45 59760 50
rect 59640 15 59645 45
rect 59675 15 59685 45
rect 59715 15 59725 45
rect 59755 15 59760 45
rect 59640 -800 59760 15
rect 59990 45 60110 50
rect 59990 15 59995 45
rect 60025 15 60035 45
rect 60065 15 60075 45
rect 60105 15 60110 45
rect 59990 -800 60110 15
rect 60340 45 60460 50
rect 60340 15 60345 45
rect 60375 15 60385 45
rect 60415 15 60425 45
rect 60455 15 60460 45
rect 60340 -800 60460 15
rect 60690 45 60810 50
rect 60690 15 60695 45
rect 60725 15 60735 45
rect 60765 15 60775 45
rect 60805 15 60810 45
rect 60690 -800 60810 15
rect 61040 45 61160 50
rect 61040 15 61045 45
rect 61075 15 61085 45
rect 61115 15 61125 45
rect 61155 15 61160 45
rect 61040 -800 61160 15
<< via1 >>
rect 52645 4275 52675 4305
rect 52685 4275 52715 4305
rect 52725 4275 52755 4305
rect 52995 4275 53025 4305
rect 53035 4275 53065 4305
rect 53075 4275 53105 4305
rect 53345 4275 53375 4305
rect 53385 4275 53415 4305
rect 53425 4275 53455 4305
rect 53695 4275 53725 4305
rect 53735 4275 53765 4305
rect 53775 4275 53805 4305
rect 54045 4275 54075 4305
rect 54085 4275 54115 4305
rect 54125 4275 54155 4305
rect 54395 4275 54425 4305
rect 54435 4275 54465 4305
rect 54475 4275 54505 4305
rect 54745 4275 54775 4305
rect 54785 4275 54815 4305
rect 54825 4275 54855 4305
rect 55095 4275 55125 4305
rect 55135 4275 55165 4305
rect 55175 4275 55205 4305
rect 55285 4275 55315 4305
rect 54985 4180 55015 4210
rect 55025 4180 55055 4210
rect 55065 4180 55095 4210
rect 55105 4180 55135 4210
rect 55145 4180 55175 4210
rect 55185 4180 55215 4210
rect 55225 4180 55255 4210
rect 54985 4140 55015 4170
rect 55025 4140 55055 4170
rect 55065 4140 55095 4170
rect 55105 4140 55135 4170
rect 55145 4140 55175 4170
rect 55185 4140 55215 4170
rect 55225 4140 55255 4170
rect 54985 4100 55015 4130
rect 55025 4100 55055 4130
rect 55065 4100 55095 4130
rect 55105 4100 55135 4130
rect 55145 4100 55175 4130
rect 55185 4100 55215 4130
rect 55225 4100 55255 4130
rect 54925 4045 54955 4075
rect 55045 4045 55075 4075
rect 55165 4045 55195 4075
rect 56210 4990 56240 5020
rect 56090 4960 56120 4965
rect 56090 4940 56095 4960
rect 56095 4940 56115 4960
rect 56115 4940 56120 4960
rect 56090 4935 56120 4940
rect 56680 4990 56710 5020
rect 56210 4935 56240 4965
rect 56270 4960 56300 4965
rect 56270 4940 56275 4960
rect 56275 4940 56295 4960
rect 56295 4940 56300 4960
rect 56270 4935 56300 4940
rect 56560 4790 56590 4795
rect 56560 4770 56565 4790
rect 56565 4770 56585 4790
rect 56585 4770 56590 4790
rect 56560 4765 56590 4770
rect 56620 4765 56650 4795
rect 57090 4990 57120 5020
rect 57560 4990 57590 5020
rect 56885 4935 56915 4965
rect 57030 4960 57060 4965
rect 57030 4940 57035 4960
rect 57035 4940 57055 4960
rect 57055 4940 57060 4960
rect 57030 4935 57060 4940
rect 56740 4790 56770 4795
rect 56740 4770 56745 4790
rect 56745 4770 56765 4790
rect 56765 4770 56770 4790
rect 56740 4765 56770 4770
rect 56885 4765 56915 4795
rect 56210 4530 56240 4560
rect 56680 4530 56710 4560
rect 56155 4510 56185 4515
rect 56155 4490 56160 4510
rect 56160 4490 56180 4510
rect 56180 4490 56185 4510
rect 56155 4485 56185 4490
rect 56630 4510 56660 4515
rect 56630 4490 56635 4510
rect 56635 4490 56655 4510
rect 56655 4490 56660 4510
rect 56630 4485 56660 4490
rect 56830 4485 56860 4515
rect 55445 4275 55475 4305
rect 55485 4275 55515 4305
rect 55525 4275 55555 4305
rect 55755 4275 55785 4305
rect 55795 4275 55825 4305
rect 55835 4275 55865 4305
rect 55875 4275 55905 4305
rect 55345 4180 55375 4210
rect 55385 4180 55415 4210
rect 55425 4180 55455 4210
rect 55465 4180 55495 4210
rect 55505 4180 55535 4210
rect 55545 4180 55575 4210
rect 55585 4180 55615 4210
rect 55345 4140 55375 4170
rect 55385 4140 55415 4170
rect 55425 4140 55455 4170
rect 55465 4140 55495 4170
rect 55505 4140 55535 4170
rect 55545 4140 55575 4170
rect 55585 4140 55615 4170
rect 55345 4100 55375 4130
rect 55385 4100 55415 4130
rect 55425 4100 55455 4130
rect 55465 4100 55495 4130
rect 55505 4100 55535 4130
rect 55545 4100 55575 4130
rect 55585 4100 55615 4130
rect 55285 4045 55315 4075
rect 55405 4045 55435 4075
rect 55525 4045 55555 4075
rect 55645 4045 55675 4075
rect 54985 3655 55015 3685
rect 55105 3655 55135 3685
rect 55225 3655 55255 3685
rect 55345 3655 55375 3685
rect 55465 3655 55495 3685
rect 55585 3655 55615 3685
rect 55285 3555 55315 3560
rect 55285 3535 55290 3555
rect 55290 3535 55310 3555
rect 55310 3535 55315 3555
rect 55285 3530 55315 3535
rect 55605 3485 55635 3515
rect 55645 3485 55675 3515
rect 55685 3485 55715 3515
rect 55605 3445 55635 3475
rect 55645 3445 55675 3475
rect 55685 3445 55715 3475
rect 55605 3405 55635 3435
rect 55645 3405 55675 3435
rect 55685 3405 55715 3435
rect 54610 3370 54640 3400
rect 54825 3350 54855 3380
rect 54935 3350 54965 3380
rect 55045 3350 55075 3380
rect 55155 3350 55185 3380
rect 55265 3350 55295 3380
rect 55375 3350 55405 3380
rect 55485 3350 55515 3380
rect 54880 3270 54910 3300
rect 54990 3270 55020 3300
rect 55100 3270 55130 3300
rect 55210 3270 55240 3300
rect 55320 3270 55350 3300
rect 55430 3270 55460 3300
rect 54880 2630 54910 2660
rect 54570 2550 54600 2580
rect 54610 2550 54640 2580
rect 54650 2550 54680 2580
rect 54570 2510 54600 2540
rect 54610 2510 54640 2540
rect 54650 2510 54680 2540
rect 54570 2470 54600 2500
rect 54610 2470 54640 2500
rect 54650 2470 54680 2500
rect 54990 2630 55020 2660
rect 55100 2630 55130 2660
rect 55210 2630 55240 2660
rect 55155 2575 55185 2580
rect 55155 2555 55160 2575
rect 55160 2555 55180 2575
rect 55180 2555 55185 2575
rect 55155 2550 55185 2555
rect 55155 2535 55185 2540
rect 55155 2515 55160 2535
rect 55160 2515 55180 2535
rect 55180 2515 55185 2535
rect 55155 2510 55185 2515
rect 55155 2495 55185 2500
rect 55155 2475 55160 2495
rect 55160 2475 55180 2495
rect 55180 2475 55185 2495
rect 55155 2470 55185 2475
rect 55320 2630 55350 2660
rect 55430 2630 55460 2660
rect 54190 2400 54220 2430
rect 54230 2400 54260 2430
rect 54275 2400 54305 2430
rect 54315 2400 54345 2430
rect 54360 2400 54390 2430
rect 54400 2400 54430 2430
rect 54190 2360 54220 2390
rect 54230 2360 54260 2390
rect 54275 2360 54305 2390
rect 54315 2360 54345 2390
rect 54360 2360 54390 2390
rect 54400 2360 54430 2390
rect 54190 2320 54220 2350
rect 54230 2320 54260 2350
rect 54275 2320 54305 2350
rect 54315 2320 54345 2350
rect 54360 2320 54390 2350
rect 54400 2320 54430 2350
rect 54120 2215 54150 2245
rect 54880 2400 54910 2430
rect 54935 2400 54965 2430
rect 54990 2400 55020 2430
rect 55045 2400 55075 2430
rect 55100 2400 55130 2430
rect 55155 2400 55185 2430
rect 55210 2400 55240 2430
rect 55265 2400 55295 2430
rect 55320 2400 55350 2430
rect 55375 2400 55405 2430
rect 55430 2400 55460 2430
rect 54880 2360 54910 2390
rect 54935 2360 54965 2390
rect 54990 2360 55020 2390
rect 55045 2360 55075 2390
rect 55100 2360 55130 2390
rect 55155 2360 55185 2390
rect 55210 2360 55240 2390
rect 55265 2360 55295 2390
rect 55320 2360 55350 2390
rect 55375 2360 55405 2390
rect 55430 2360 55460 2390
rect 54880 2320 54910 2350
rect 54935 2320 54965 2350
rect 54990 2320 55020 2350
rect 55045 2320 55075 2350
rect 55100 2320 55130 2350
rect 55155 2320 55185 2350
rect 55210 2320 55240 2350
rect 55265 2320 55295 2350
rect 55320 2320 55350 2350
rect 55375 2320 55405 2350
rect 55430 2320 55460 2350
rect 56010 4180 56040 4210
rect 56050 4180 56080 4210
rect 56090 4180 56120 4210
rect 56130 4180 56160 4210
rect 56170 4180 56200 4210
rect 56210 4180 56240 4210
rect 56250 4180 56280 4210
rect 56290 4180 56320 4210
rect 56330 4180 56360 4210
rect 56370 4180 56400 4210
rect 56410 4180 56440 4210
rect 56450 4180 56480 4210
rect 56490 4180 56520 4210
rect 56530 4180 56560 4210
rect 56570 4180 56600 4210
rect 56610 4180 56640 4210
rect 56650 4180 56680 4210
rect 56690 4180 56720 4210
rect 56730 4180 56760 4210
rect 56010 4140 56040 4170
rect 56050 4140 56080 4170
rect 56090 4140 56120 4170
rect 56130 4140 56160 4170
rect 56170 4140 56200 4170
rect 56210 4140 56240 4170
rect 56250 4140 56280 4170
rect 56290 4140 56320 4170
rect 56330 4140 56360 4170
rect 56370 4140 56400 4170
rect 56410 4140 56440 4170
rect 56450 4140 56480 4170
rect 56490 4140 56520 4170
rect 56530 4140 56560 4170
rect 56570 4140 56600 4170
rect 56610 4140 56640 4170
rect 56650 4140 56680 4170
rect 56690 4140 56720 4170
rect 56730 4140 56760 4170
rect 56010 4100 56040 4130
rect 56050 4100 56080 4130
rect 56090 4100 56120 4130
rect 56130 4100 56160 4130
rect 56170 4100 56200 4130
rect 56210 4100 56240 4130
rect 56250 4100 56280 4130
rect 56290 4100 56320 4130
rect 56330 4100 56360 4130
rect 56370 4100 56400 4130
rect 56410 4100 56440 4130
rect 56450 4100 56480 4130
rect 56490 4100 56520 4130
rect 56530 4100 56560 4130
rect 56570 4100 56600 4130
rect 56610 4100 56640 4130
rect 56650 4100 56680 4130
rect 56690 4100 56720 4130
rect 56730 4100 56760 4130
rect 56070 4045 56100 4075
rect 56190 4045 56220 4075
rect 56310 4045 56340 4075
rect 56430 4045 56460 4075
rect 56550 4045 56580 4075
rect 56670 4045 56700 4075
rect 56070 3655 56100 3685
rect 56190 3655 56220 3685
rect 56310 3655 56340 3685
rect 56430 3655 56460 3685
rect 56370 3600 56400 3605
rect 56370 3580 56375 3600
rect 56375 3580 56395 3600
rect 56395 3580 56400 3600
rect 56370 3575 56400 3580
rect 56550 3655 56580 3685
rect 56670 3655 56700 3685
rect 57150 4935 57180 4965
rect 57210 4960 57240 4965
rect 57210 4940 57215 4960
rect 57215 4940 57235 4960
rect 57235 4940 57240 4960
rect 57210 4935 57240 4940
rect 57500 4960 57530 4965
rect 57500 4940 57505 4960
rect 57505 4940 57525 4960
rect 57525 4940 57530 4960
rect 57500 4935 57530 4940
rect 57560 4935 57590 4965
rect 57680 4960 57710 4965
rect 57680 4940 57685 4960
rect 57685 4940 57705 4960
rect 57705 4940 57710 4960
rect 57680 4935 57710 4940
rect 57090 4530 57120 4560
rect 57560 4530 57590 4560
rect 56940 4430 56970 4460
rect 57576 4500 57606 4505
rect 57576 4480 57581 4500
rect 57581 4480 57601 4500
rect 57601 4480 57606 4500
rect 57576 4475 57606 4480
rect 56885 4275 56915 4305
rect 56840 3575 56870 3605
rect 57140 4420 57170 4450
rect 57620 4420 57650 4450
rect 57895 4275 57925 4305
rect 57935 4275 57965 4305
rect 57975 4275 58005 4305
rect 58015 4275 58045 4305
rect 58245 4275 58275 4305
rect 58285 4275 58315 4305
rect 58325 4275 58355 4305
rect 58485 4275 58515 4305
rect 57040 4180 57070 4210
rect 57080 4180 57110 4210
rect 57120 4180 57150 4210
rect 57160 4180 57190 4210
rect 57200 4180 57230 4210
rect 57240 4180 57270 4210
rect 57280 4180 57310 4210
rect 57320 4180 57350 4210
rect 57360 4180 57390 4210
rect 57400 4180 57430 4210
rect 57440 4180 57470 4210
rect 57480 4180 57510 4210
rect 57520 4180 57550 4210
rect 57560 4180 57590 4210
rect 57600 4180 57630 4210
rect 57640 4180 57670 4210
rect 57680 4180 57710 4210
rect 57720 4180 57750 4210
rect 57760 4180 57790 4210
rect 57040 4140 57070 4170
rect 57080 4140 57110 4170
rect 57120 4140 57150 4170
rect 57160 4140 57190 4170
rect 57200 4140 57230 4170
rect 57240 4140 57270 4170
rect 57280 4140 57310 4170
rect 57320 4140 57350 4170
rect 57360 4140 57390 4170
rect 57400 4140 57430 4170
rect 57440 4140 57470 4170
rect 57480 4140 57510 4170
rect 57520 4140 57550 4170
rect 57560 4140 57590 4170
rect 57600 4140 57630 4170
rect 57640 4140 57670 4170
rect 57680 4140 57710 4170
rect 57720 4140 57750 4170
rect 57760 4140 57790 4170
rect 57040 4100 57070 4130
rect 57080 4100 57110 4130
rect 57120 4100 57150 4130
rect 57160 4100 57190 4130
rect 57200 4100 57230 4130
rect 57240 4100 57270 4130
rect 57280 4100 57310 4130
rect 57320 4100 57350 4130
rect 57360 4100 57390 4130
rect 57400 4100 57430 4130
rect 57440 4100 57470 4130
rect 57480 4100 57510 4130
rect 57520 4100 57550 4130
rect 57560 4100 57590 4130
rect 57600 4100 57630 4130
rect 57640 4100 57670 4130
rect 57680 4100 57710 4130
rect 57720 4100 57750 4130
rect 57760 4100 57790 4130
rect 57100 4045 57130 4075
rect 57220 4045 57250 4075
rect 57340 4045 57370 4075
rect 57460 4045 57490 4075
rect 57580 4045 57610 4075
rect 57700 4045 57730 4075
rect 57100 3655 57130 3685
rect 56930 3530 56960 3560
rect 56070 3485 56100 3515
rect 56110 3485 56140 3515
rect 56150 3485 56180 3515
rect 56190 3485 56220 3515
rect 56230 3485 56260 3515
rect 56270 3485 56300 3515
rect 56310 3485 56340 3515
rect 56350 3485 56380 3515
rect 56390 3485 56420 3515
rect 56430 3485 56460 3515
rect 56470 3485 56500 3515
rect 56510 3485 56540 3515
rect 56550 3485 56580 3515
rect 56590 3485 56620 3515
rect 56630 3485 56660 3515
rect 56670 3485 56700 3515
rect 56070 3445 56100 3475
rect 56110 3445 56140 3475
rect 56150 3445 56180 3475
rect 56190 3445 56220 3475
rect 56230 3445 56260 3475
rect 56270 3445 56300 3475
rect 56310 3445 56340 3475
rect 56350 3445 56380 3475
rect 56390 3445 56420 3475
rect 56430 3445 56460 3475
rect 56470 3445 56500 3475
rect 56510 3445 56540 3475
rect 56550 3445 56580 3475
rect 56590 3445 56620 3475
rect 56630 3445 56660 3475
rect 56670 3445 56700 3475
rect 56070 3405 56100 3435
rect 56110 3405 56140 3435
rect 56150 3405 56180 3435
rect 56190 3405 56220 3435
rect 56230 3405 56260 3435
rect 56270 3405 56300 3435
rect 56310 3405 56340 3435
rect 56350 3405 56380 3435
rect 56390 3405 56420 3435
rect 56430 3405 56460 3435
rect 56470 3405 56500 3435
rect 56510 3405 56540 3435
rect 56550 3405 56580 3435
rect 56590 3405 56620 3435
rect 56630 3405 56660 3435
rect 56670 3405 56700 3435
rect 57220 3655 57250 3685
rect 57340 3655 57370 3685
rect 57460 3655 57490 3685
rect 57400 3600 57430 3605
rect 57400 3580 57405 3600
rect 57405 3580 57425 3600
rect 57425 3580 57430 3600
rect 57400 3575 57430 3580
rect 57580 3655 57610 3685
rect 57700 3655 57730 3685
rect 57100 3485 57130 3515
rect 57140 3485 57170 3515
rect 57180 3485 57210 3515
rect 57220 3485 57250 3515
rect 57260 3485 57290 3515
rect 57300 3485 57330 3515
rect 57340 3485 57370 3515
rect 57380 3485 57410 3515
rect 57420 3485 57450 3515
rect 57460 3485 57490 3515
rect 57500 3485 57530 3515
rect 57540 3485 57570 3515
rect 57580 3485 57610 3515
rect 57620 3485 57650 3515
rect 57660 3485 57690 3515
rect 57700 3485 57730 3515
rect 57100 3445 57130 3475
rect 57140 3445 57170 3475
rect 57180 3445 57210 3475
rect 57220 3445 57250 3475
rect 57260 3445 57290 3475
rect 57300 3445 57330 3475
rect 57340 3445 57370 3475
rect 57380 3445 57410 3475
rect 57420 3445 57450 3475
rect 57460 3445 57490 3475
rect 57500 3445 57530 3475
rect 57540 3445 57570 3475
rect 57580 3445 57610 3475
rect 57620 3445 57650 3475
rect 57660 3445 57690 3475
rect 57700 3445 57730 3475
rect 57100 3405 57130 3435
rect 57140 3405 57170 3435
rect 57180 3405 57210 3435
rect 57220 3405 57250 3435
rect 57260 3405 57290 3435
rect 57300 3405 57330 3435
rect 57340 3405 57370 3435
rect 57380 3405 57410 3435
rect 57420 3405 57450 3435
rect 57460 3405 57490 3435
rect 57500 3405 57530 3435
rect 57540 3405 57570 3435
rect 57580 3405 57610 3435
rect 57620 3405 57650 3435
rect 57660 3405 57690 3435
rect 57700 3405 57730 3435
rect 58185 4180 58215 4210
rect 58225 4180 58255 4210
rect 58265 4180 58295 4210
rect 58305 4180 58335 4210
rect 58345 4180 58375 4210
rect 58385 4180 58415 4210
rect 58425 4180 58455 4210
rect 58185 4140 58215 4170
rect 58225 4140 58255 4170
rect 58265 4140 58295 4170
rect 58305 4140 58335 4170
rect 58345 4140 58375 4170
rect 58385 4140 58415 4170
rect 58425 4140 58455 4170
rect 58185 4100 58215 4130
rect 58225 4100 58255 4130
rect 58265 4100 58295 4130
rect 58305 4100 58335 4130
rect 58345 4100 58375 4130
rect 58385 4100 58415 4130
rect 58425 4100 58455 4130
rect 58125 4045 58155 4075
rect 58245 4045 58275 4075
rect 58365 4045 58395 4075
rect 58595 4275 58625 4305
rect 58635 4275 58665 4305
rect 58675 4275 58705 4305
rect 58945 4275 58975 4305
rect 58985 4275 59015 4305
rect 59025 4275 59055 4305
rect 59295 4275 59325 4305
rect 59335 4275 59365 4305
rect 59375 4275 59405 4305
rect 59645 4275 59675 4305
rect 59685 4275 59715 4305
rect 59725 4275 59755 4305
rect 59995 4275 60025 4305
rect 60035 4275 60065 4305
rect 60075 4275 60105 4305
rect 60345 4275 60375 4305
rect 60385 4275 60415 4305
rect 60425 4275 60455 4305
rect 60695 4275 60725 4305
rect 60735 4275 60765 4305
rect 60775 4275 60805 4305
rect 61045 4275 61075 4305
rect 61085 4275 61115 4305
rect 61125 4275 61155 4305
rect 58545 4180 58575 4210
rect 58585 4180 58615 4210
rect 58625 4180 58655 4210
rect 58665 4180 58695 4210
rect 58705 4180 58735 4210
rect 58745 4180 58775 4210
rect 58785 4180 58815 4210
rect 58545 4140 58575 4170
rect 58585 4140 58615 4170
rect 58625 4140 58655 4170
rect 58665 4140 58695 4170
rect 58705 4140 58735 4170
rect 58745 4140 58775 4170
rect 58785 4140 58815 4170
rect 58545 4100 58575 4130
rect 58585 4100 58615 4130
rect 58625 4100 58655 4130
rect 58665 4100 58695 4130
rect 58705 4100 58735 4130
rect 58745 4100 58775 4130
rect 58785 4100 58815 4130
rect 58485 4045 58515 4075
rect 58605 4045 58635 4075
rect 58725 4045 58755 4075
rect 58845 4045 58875 4075
rect 58185 3655 58215 3685
rect 58305 3655 58335 3685
rect 58425 3655 58455 3685
rect 58545 3655 58575 3685
rect 58665 3655 58695 3685
rect 58785 3655 58815 3685
rect 58485 3555 58515 3560
rect 58485 3535 58490 3555
rect 58490 3535 58510 3555
rect 58510 3535 58515 3555
rect 58485 3530 58515 3535
rect 58085 3485 58115 3515
rect 58125 3485 58155 3515
rect 58165 3485 58195 3515
rect 58085 3445 58115 3475
rect 58125 3445 58155 3475
rect 58165 3445 58195 3475
rect 58085 3405 58115 3435
rect 58125 3405 58155 3435
rect 58165 3405 58195 3435
rect 55755 3350 55785 3380
rect 56280 3350 56310 3380
rect 56390 3350 56420 3380
rect 56500 3350 56530 3380
rect 56610 3350 56640 3380
rect 56720 3350 56750 3380
rect 56830 3350 56860 3380
rect 56940 3350 56970 3380
rect 57050 3350 57080 3380
rect 57160 3350 57190 3380
rect 57270 3350 57300 3380
rect 57380 3350 57410 3380
rect 57490 3350 57520 3380
rect 58015 3350 58045 3380
rect 56335 3305 56365 3335
rect 56445 3260 56475 3290
rect 56335 3170 56365 3200
rect 56555 3305 56585 3335
rect 56665 3260 56695 3290
rect 56555 3170 56585 3200
rect 56775 3305 56805 3335
rect 56885 3260 56915 3290
rect 56775 3170 56805 3200
rect 56445 3100 56475 3130
rect 56665 3100 56695 3130
rect 55945 2990 55975 3020
rect 56040 3015 56070 3020
rect 56040 2995 56045 3015
rect 56045 2995 56065 3015
rect 56065 2995 56070 3015
rect 56040 2990 56070 2995
rect 56145 2995 56175 3025
rect 56255 2995 56285 3025
rect 56365 2995 56395 3025
rect 56475 2995 56505 3025
rect 56585 2995 56615 3025
rect 56690 3015 56720 3020
rect 56690 2995 56695 3015
rect 56695 2995 56715 3015
rect 56715 2995 56720 3015
rect 56690 2990 56720 2995
rect 55755 2715 55785 2745
rect 55605 2550 55635 2580
rect 55645 2550 55675 2580
rect 55685 2550 55715 2580
rect 55605 2510 55635 2540
rect 55645 2510 55675 2540
rect 55685 2510 55715 2540
rect 55605 2470 55635 2500
rect 55645 2470 55675 2500
rect 55685 2470 55715 2500
rect 54825 2260 54855 2290
rect 55485 2260 55515 2290
rect 54880 2215 54910 2245
rect 54990 2215 55020 2245
rect 55100 2215 55130 2245
rect 55210 2215 55240 2245
rect 55320 2215 55350 2245
rect 55430 2215 55460 2245
rect 54935 2170 54965 2200
rect 55045 2170 55075 2200
rect 55155 2170 55185 2200
rect 55265 2170 55295 2200
rect 55375 2170 55405 2200
rect 54685 1915 54715 1945
rect 54935 1940 54965 1945
rect 54935 1920 54940 1940
rect 54940 1920 54960 1940
rect 54960 1920 54965 1940
rect 54935 1915 54965 1920
rect 55045 1940 55075 1945
rect 55045 1920 55050 1940
rect 55050 1920 55070 1940
rect 55070 1920 55075 1940
rect 55045 1915 55075 1920
rect 55155 1940 55185 1945
rect 55155 1920 55160 1940
rect 55160 1920 55180 1940
rect 55180 1920 55185 1940
rect 55155 1915 55185 1920
rect 55265 1940 55295 1945
rect 55265 1920 55270 1940
rect 55270 1920 55290 1940
rect 55290 1920 55295 1940
rect 55265 1915 55295 1920
rect 55375 1940 55405 1945
rect 55375 1920 55380 1940
rect 55380 1920 55400 1940
rect 55400 1920 55405 1940
rect 55375 1915 55405 1920
rect 54195 1680 54225 1710
rect 54245 1680 54275 1710
rect 54295 1680 54325 1710
rect 54345 1680 54375 1710
rect 54395 1680 54425 1710
rect 54195 1630 54225 1660
rect 54245 1630 54275 1660
rect 54295 1630 54325 1660
rect 54345 1630 54375 1660
rect 54395 1630 54425 1660
rect 54195 1580 54225 1610
rect 54245 1580 54275 1610
rect 54295 1580 54325 1610
rect 54345 1580 54375 1610
rect 54395 1580 54425 1610
rect 54460 1390 54495 1395
rect 54460 1365 54465 1390
rect 54465 1365 54490 1390
rect 54490 1365 54495 1390
rect 54460 1360 54495 1365
rect 54520 1390 54555 1395
rect 54520 1365 54525 1390
rect 54525 1365 54550 1390
rect 54550 1365 54555 1390
rect 54520 1360 54555 1365
rect 54580 1390 54615 1395
rect 54580 1365 54585 1390
rect 54585 1365 54610 1390
rect 54610 1365 54615 1390
rect 54580 1360 54615 1365
rect 54640 1390 54675 1395
rect 54640 1365 54645 1390
rect 54645 1365 54670 1390
rect 54670 1365 54675 1390
rect 54640 1360 54675 1365
rect 55320 1875 55350 1880
rect 55320 1855 55325 1875
rect 55325 1855 55345 1875
rect 55345 1855 55350 1875
rect 55320 1850 55350 1855
rect 55320 1835 55350 1840
rect 55320 1815 55325 1835
rect 55325 1815 55345 1835
rect 55345 1815 55350 1835
rect 55320 1810 55350 1815
rect 55755 2260 55785 2290
rect 55605 1850 55635 1880
rect 55645 1850 55675 1880
rect 55685 1850 55715 1880
rect 55605 1810 55635 1840
rect 55645 1810 55675 1840
rect 55685 1810 55715 1840
rect 54730 1730 54760 1760
rect 54935 1730 54965 1760
rect 55045 1730 55075 1760
rect 55155 1730 55185 1760
rect 55265 1730 55295 1760
rect 55375 1730 55405 1760
rect 54730 1360 54760 1390
rect 54935 1390 54965 1420
rect 55045 1390 55075 1420
rect 55155 1390 55185 1420
rect 55265 1390 55295 1420
rect 55375 1390 55405 1420
rect 55900 2240 55930 2270
rect 54585 1305 54615 1335
rect 54880 1345 54910 1375
rect 54990 1345 55020 1375
rect 55100 1345 55130 1375
rect 55210 1345 55240 1375
rect 55320 1345 55350 1375
rect 55430 1345 55460 1375
rect 55755 1345 55785 1375
rect 54685 1305 54715 1335
rect 54825 1300 54855 1330
rect 55485 1300 55515 1330
rect 55835 1300 55865 1330
rect 54465 1255 54495 1285
rect 54600 1210 54630 1240
rect 55185 1235 55215 1240
rect 55185 1215 55190 1235
rect 55190 1215 55210 1235
rect 55210 1215 55215 1235
rect 55185 1210 55215 1215
rect 54190 1155 54220 1185
rect 54230 1155 54260 1185
rect 54275 1155 54305 1185
rect 54315 1155 54345 1185
rect 54360 1155 54390 1185
rect 54400 1155 54430 1185
rect 54190 1115 54220 1145
rect 54230 1115 54260 1145
rect 54275 1115 54305 1145
rect 54315 1115 54345 1145
rect 54360 1115 54390 1145
rect 54400 1115 54430 1145
rect 54190 1075 54220 1105
rect 54230 1075 54260 1105
rect 54275 1075 54305 1105
rect 54315 1075 54345 1105
rect 54360 1075 54390 1105
rect 54400 1075 54430 1105
rect 54665 1155 54695 1185
rect 54665 1115 54695 1145
rect 54665 1075 54695 1105
rect 54935 1155 54965 1185
rect 54975 1155 55005 1185
rect 55015 1155 55045 1185
rect 55055 1155 55085 1185
rect 55095 1155 55125 1185
rect 55135 1155 55165 1185
rect 55175 1155 55205 1185
rect 55215 1155 55245 1185
rect 55255 1155 55285 1185
rect 55295 1155 55325 1185
rect 55335 1155 55365 1185
rect 54935 1115 54965 1145
rect 54975 1115 55005 1145
rect 55015 1115 55045 1145
rect 55055 1115 55085 1145
rect 55095 1115 55125 1145
rect 55135 1115 55165 1145
rect 55175 1115 55205 1145
rect 55215 1115 55245 1145
rect 55255 1115 55285 1145
rect 55295 1115 55325 1145
rect 55335 1115 55365 1145
rect 54935 1075 54965 1105
rect 54975 1075 55005 1105
rect 55015 1075 55045 1105
rect 55055 1075 55085 1105
rect 55095 1075 55125 1105
rect 55135 1075 55165 1105
rect 55175 1075 55205 1105
rect 55215 1075 55245 1105
rect 55255 1075 55285 1105
rect 55295 1075 55325 1105
rect 55335 1075 55365 1105
rect 54600 1045 54635 1050
rect 54600 1020 54605 1045
rect 54605 1020 54630 1045
rect 54630 1020 54635 1045
rect 54600 1015 54635 1020
rect 54660 1045 54695 1050
rect 54660 1020 54665 1045
rect 54665 1020 54690 1045
rect 54690 1020 54695 1045
rect 54660 1015 54695 1020
rect 54935 320 54965 350
rect 55135 320 55165 350
rect 55835 710 55865 740
rect 55335 320 55365 350
rect 56090 2950 56120 2980
rect 56200 2950 56230 2980
rect 56145 2860 56175 2890
rect 56310 2950 56340 2980
rect 56255 2860 56285 2890
rect 56420 2950 56450 2980
rect 56365 2860 56395 2890
rect 56530 2950 56560 2980
rect 56475 2860 56505 2890
rect 56640 2950 56670 2980
rect 56585 2860 56615 2890
rect 56995 3305 57025 3335
rect 57105 3260 57135 3290
rect 56995 3170 57025 3200
rect 57215 3305 57245 3335
rect 57325 3260 57355 3290
rect 57215 3170 57245 3200
rect 56885 3100 56915 3130
rect 57105 3100 57135 3130
rect 57435 3305 57465 3335
rect 57435 3170 57465 3200
rect 57325 3100 57355 3130
rect 57080 3015 57110 3020
rect 57080 2995 57085 3015
rect 57085 2995 57105 3015
rect 57105 2995 57110 3015
rect 57080 2990 57110 2995
rect 57185 2995 57215 3025
rect 57295 2995 57325 3025
rect 57405 2995 57435 3025
rect 57515 2995 57545 3025
rect 57625 2995 57655 3025
rect 57730 3015 57760 3020
rect 57730 2995 57735 3015
rect 57735 2995 57755 3015
rect 57755 2995 57760 3015
rect 57730 2990 57760 2995
rect 57130 2950 57160 2980
rect 57185 2860 57215 2890
rect 56090 2815 56120 2845
rect 56200 2815 56230 2845
rect 56310 2815 56340 2845
rect 56420 2815 56450 2845
rect 56530 2815 56560 2845
rect 56640 2815 56670 2845
rect 56580 2795 56610 2800
rect 56095 2785 56125 2790
rect 56095 2765 56100 2785
rect 56100 2765 56120 2785
rect 56120 2765 56125 2785
rect 56580 2775 56585 2795
rect 56585 2775 56605 2795
rect 56605 2775 56610 2795
rect 56580 2770 56610 2775
rect 56095 2760 56125 2765
rect 56830 2815 56860 2845
rect 57130 2815 57160 2845
rect 57190 2795 57220 2800
rect 57190 2775 57195 2795
rect 57195 2775 57215 2795
rect 57215 2775 57220 2795
rect 57190 2770 57220 2775
rect 56035 2715 56065 2745
rect 56695 2715 56725 2745
rect 57075 2715 57105 2745
rect 57350 2950 57380 2980
rect 57295 2860 57325 2890
rect 57405 2860 57435 2890
rect 57350 2815 57380 2845
rect 56940 2660 56970 2690
rect 57240 2660 57270 2690
rect 57570 2950 57600 2980
rect 57515 2860 57545 2890
rect 57825 2990 57855 3020
rect 57625 2860 57655 2890
rect 57570 2815 57600 2845
rect 57735 2715 57765 2745
rect 57460 2660 57490 2690
rect 57680 2660 57710 2690
rect 56855 2630 56885 2635
rect 56855 2610 56860 2630
rect 56860 2610 56880 2630
rect 56880 2610 56885 2630
rect 56855 2605 56885 2610
rect 57350 2605 57380 2635
rect 56090 2550 56120 2580
rect 56145 2550 56175 2580
rect 56200 2550 56230 2580
rect 56255 2550 56285 2580
rect 56310 2550 56340 2580
rect 56365 2550 56395 2580
rect 56420 2550 56450 2580
rect 56475 2550 56505 2580
rect 56530 2550 56560 2580
rect 56585 2550 56615 2580
rect 56640 2550 56670 2580
rect 56090 2510 56120 2540
rect 56145 2510 56175 2540
rect 56200 2510 56230 2540
rect 56255 2510 56285 2540
rect 56310 2510 56340 2540
rect 56365 2510 56395 2540
rect 56420 2510 56450 2540
rect 56475 2510 56505 2540
rect 56530 2510 56560 2540
rect 56585 2510 56615 2540
rect 56640 2510 56670 2540
rect 56090 2470 56120 2500
rect 56145 2470 56175 2500
rect 56200 2470 56230 2500
rect 56255 2470 56285 2500
rect 56310 2470 56340 2500
rect 56365 2470 56395 2500
rect 56420 2470 56450 2500
rect 56475 2470 56505 2500
rect 56530 2470 56560 2500
rect 56585 2470 56615 2500
rect 56640 2470 56670 2500
rect 55995 2265 56025 2270
rect 55995 2245 56000 2265
rect 56000 2245 56020 2265
rect 56020 2245 56025 2265
rect 55995 2240 56025 2245
rect 56145 2230 56175 2260
rect 56090 2185 56120 2215
rect 56255 2230 56285 2260
rect 56200 2185 56230 2215
rect 56145 1995 56175 2025
rect 56090 1950 56120 1980
rect 56035 1905 56065 1935
rect 56365 2230 56395 2260
rect 56310 2185 56340 2215
rect 56255 1995 56285 2025
rect 56200 1950 56230 1980
rect 56040 1780 56070 1785
rect 56040 1760 56045 1780
rect 56045 1760 56065 1780
rect 56065 1760 56070 1780
rect 56090 1765 56120 1795
rect 56145 1775 56175 1805
rect 56475 2230 56505 2260
rect 56420 2185 56450 2215
rect 56365 1995 56395 2025
rect 56310 1950 56340 1980
rect 56200 1765 56230 1795
rect 56255 1775 56285 1805
rect 56585 2230 56615 2260
rect 56530 2185 56560 2215
rect 56475 1995 56505 2025
rect 56420 1950 56450 1980
rect 56310 1765 56340 1795
rect 56365 1775 56395 1805
rect 57130 2550 57160 2580
rect 57185 2550 57215 2580
rect 57240 2550 57270 2580
rect 57295 2550 57325 2580
rect 57350 2550 57380 2580
rect 57405 2550 57435 2580
rect 57460 2550 57490 2580
rect 57515 2550 57545 2580
rect 57570 2550 57600 2580
rect 57625 2550 57655 2580
rect 57680 2550 57710 2580
rect 57130 2510 57160 2540
rect 57185 2510 57215 2540
rect 57240 2510 57270 2540
rect 57295 2510 57325 2540
rect 57350 2510 57380 2540
rect 57405 2510 57435 2540
rect 57460 2510 57490 2540
rect 57515 2510 57545 2540
rect 57570 2510 57600 2540
rect 57625 2510 57655 2540
rect 57680 2510 57710 2540
rect 57130 2470 57160 2500
rect 57185 2470 57215 2500
rect 57240 2470 57270 2500
rect 57295 2470 57325 2500
rect 57350 2470 57380 2500
rect 57405 2470 57435 2500
rect 57460 2470 57490 2500
rect 57515 2470 57545 2500
rect 57570 2470 57600 2500
rect 57625 2470 57655 2500
rect 57680 2470 57710 2500
rect 56775 2310 56805 2315
rect 56775 2290 56780 2310
rect 56780 2290 56800 2310
rect 56800 2290 56805 2310
rect 56775 2285 56805 2290
rect 56885 2285 56915 2315
rect 56995 2310 57025 2315
rect 56995 2290 57000 2310
rect 57000 2290 57020 2310
rect 57020 2290 57025 2310
rect 56995 2285 57025 2290
rect 56690 2265 56720 2270
rect 56690 2245 56695 2265
rect 56695 2245 56715 2265
rect 56715 2245 56720 2265
rect 56690 2240 56720 2245
rect 57080 2265 57110 2270
rect 57080 2245 57085 2265
rect 57085 2245 57105 2265
rect 57105 2245 57110 2265
rect 57080 2240 57110 2245
rect 56640 2185 56670 2215
rect 57185 2230 57215 2260
rect 57130 2185 57160 2215
rect 56585 1995 56615 2025
rect 56530 1950 56560 1980
rect 56420 1765 56450 1795
rect 56475 1775 56505 1805
rect 56640 1950 56670 1980
rect 57295 2230 57325 2260
rect 57240 2185 57270 2215
rect 57185 1995 57215 2025
rect 57130 1950 57160 1980
rect 56695 1905 56725 1935
rect 57075 1905 57105 1935
rect 56530 1765 56560 1795
rect 56585 1775 56615 1805
rect 56640 1765 56670 1795
rect 56690 1780 56720 1785
rect 56690 1760 56695 1780
rect 56695 1760 56715 1780
rect 56715 1760 56720 1780
rect 56040 1755 56070 1760
rect 56145 1720 56175 1750
rect 56090 1525 56120 1555
rect 56255 1720 56285 1750
rect 56200 1525 56230 1555
rect 56365 1720 56395 1750
rect 56310 1525 56340 1555
rect 56475 1720 56505 1750
rect 56420 1525 56450 1555
rect 56585 1720 56615 1750
rect 56530 1525 56560 1555
rect 56690 1755 56720 1760
rect 56850 1780 56880 1785
rect 56850 1760 56855 1780
rect 56855 1760 56875 1780
rect 56875 1760 56880 1780
rect 56850 1755 56880 1760
rect 56903 1780 56933 1785
rect 56903 1760 56908 1780
rect 56908 1760 56928 1780
rect 56928 1760 56933 1780
rect 56903 1755 56933 1760
rect 57405 2230 57435 2260
rect 57350 2185 57380 2215
rect 57295 1995 57325 2025
rect 57240 1950 57270 1980
rect 57080 1780 57110 1785
rect 57080 1760 57085 1780
rect 57085 1760 57105 1780
rect 57105 1760 57110 1780
rect 57130 1765 57160 1795
rect 57185 1775 57215 1805
rect 57515 2230 57545 2260
rect 57460 2185 57490 2215
rect 57405 1995 57435 2025
rect 57350 1950 57380 1980
rect 57240 1765 57270 1795
rect 57295 1775 57325 1805
rect 57625 2230 57655 2260
rect 57570 2185 57600 2215
rect 57515 1995 57545 2025
rect 57460 1950 57490 1980
rect 57350 1765 57380 1795
rect 57405 1775 57435 1805
rect 57680 2185 57710 2215
rect 57625 1995 57655 2025
rect 57570 1950 57600 1980
rect 57460 1765 57490 1795
rect 57515 1775 57545 1805
rect 57680 1950 57710 1980
rect 57735 1905 57765 1935
rect 57570 1765 57600 1795
rect 57625 1775 57655 1805
rect 57680 1765 57710 1795
rect 57730 1780 57760 1785
rect 57730 1760 57735 1780
rect 57735 1760 57755 1780
rect 57755 1760 57760 1780
rect 57080 1755 57110 1760
rect 57185 1720 57215 1750
rect 56640 1525 56670 1555
rect 56145 1470 56175 1500
rect 56255 1470 56285 1500
rect 56365 1470 56395 1500
rect 56475 1470 56505 1500
rect 56585 1470 56615 1500
rect 56035 1300 56065 1330
rect 55945 1255 55975 1285
rect 56335 1085 56365 1115
rect 56830 1390 56860 1420
rect 56735 1300 56765 1330
rect 57130 1525 57160 1555
rect 57295 1720 57325 1750
rect 57240 1525 57270 1555
rect 57405 1720 57435 1750
rect 57350 1525 57380 1555
rect 57515 1720 57545 1750
rect 57460 1525 57490 1555
rect 57625 1720 57655 1750
rect 57570 1525 57600 1555
rect 57730 1755 57760 1760
rect 57680 1525 57710 1555
rect 56940 1390 56970 1420
rect 57185 1470 57215 1500
rect 57295 1470 57325 1500
rect 57035 1300 57065 1330
rect 56885 1085 56915 1115
rect 57405 1470 57435 1500
rect 57515 1470 57545 1500
rect 57625 1470 57655 1500
rect 57735 1300 57765 1330
rect 58015 2715 58045 2745
rect 57870 2660 57900 2690
rect 57825 1255 57855 1285
rect 57935 2285 57965 2315
rect 58285 3350 58315 3380
rect 58395 3350 58425 3380
rect 58505 3350 58535 3380
rect 58615 3350 58645 3380
rect 58725 3350 58755 3380
rect 58835 3350 58865 3380
rect 58945 3350 58975 3380
rect 59160 3370 59190 3400
rect 58340 3270 58370 3300
rect 58450 3270 58480 3300
rect 58560 3270 58590 3300
rect 58670 3270 58700 3300
rect 58780 3270 58810 3300
rect 58890 3270 58920 3300
rect 58085 2550 58115 2580
rect 58125 2550 58155 2580
rect 58165 2550 58195 2580
rect 58085 2510 58115 2540
rect 58125 2510 58155 2540
rect 58165 2510 58195 2540
rect 58085 2470 58115 2500
rect 58125 2470 58155 2500
rect 58165 2470 58195 2500
rect 58015 2260 58045 2290
rect 57935 1905 57965 1935
rect 58340 2630 58370 2660
rect 58450 2630 58480 2660
rect 58560 2630 58590 2660
rect 58670 2630 58700 2660
rect 58615 2575 58645 2580
rect 58615 2555 58620 2575
rect 58620 2555 58640 2575
rect 58640 2555 58645 2575
rect 58615 2550 58645 2555
rect 58615 2535 58645 2540
rect 58615 2515 58620 2535
rect 58620 2515 58640 2535
rect 58640 2515 58645 2535
rect 58615 2510 58645 2515
rect 58615 2495 58645 2500
rect 58615 2475 58620 2495
rect 58620 2475 58640 2495
rect 58640 2475 58645 2495
rect 58615 2470 58645 2475
rect 58780 2630 58810 2660
rect 58890 2630 58920 2660
rect 59120 2550 59150 2580
rect 59160 2550 59190 2580
rect 59200 2550 59230 2580
rect 59120 2510 59150 2540
rect 59160 2510 59190 2540
rect 59200 2510 59230 2540
rect 59120 2470 59150 2500
rect 59160 2470 59190 2500
rect 59200 2470 59230 2500
rect 58340 2400 58370 2430
rect 58395 2400 58425 2430
rect 58450 2400 58480 2430
rect 58505 2400 58535 2430
rect 58560 2400 58590 2430
rect 58615 2400 58645 2430
rect 58670 2400 58700 2430
rect 58725 2400 58755 2430
rect 58780 2400 58810 2430
rect 58835 2400 58865 2430
rect 58890 2400 58920 2430
rect 58340 2360 58370 2390
rect 58395 2360 58425 2390
rect 58450 2360 58480 2390
rect 58505 2360 58535 2390
rect 58560 2360 58590 2390
rect 58615 2360 58645 2390
rect 58670 2360 58700 2390
rect 58725 2360 58755 2390
rect 58780 2360 58810 2390
rect 58835 2360 58865 2390
rect 58890 2360 58920 2390
rect 58340 2320 58370 2350
rect 58395 2320 58425 2350
rect 58450 2320 58480 2350
rect 58505 2320 58535 2350
rect 58560 2320 58590 2350
rect 58615 2320 58645 2350
rect 58670 2320 58700 2350
rect 58725 2320 58755 2350
rect 58780 2320 58810 2350
rect 58835 2320 58865 2350
rect 58890 2320 58920 2350
rect 59370 2400 59400 2430
rect 59410 2400 59440 2430
rect 59455 2400 59485 2430
rect 59495 2400 59525 2430
rect 59540 2400 59570 2430
rect 59580 2400 59610 2430
rect 59370 2360 59400 2390
rect 59410 2360 59440 2390
rect 59455 2360 59485 2390
rect 59495 2360 59525 2390
rect 59540 2360 59570 2390
rect 59580 2360 59610 2390
rect 59370 2320 59400 2350
rect 59410 2320 59440 2350
rect 59455 2320 59485 2350
rect 59495 2320 59525 2350
rect 59540 2320 59570 2350
rect 59580 2320 59610 2350
rect 58285 2260 58315 2290
rect 58945 2260 58975 2290
rect 58340 2215 58370 2245
rect 58450 2215 58480 2245
rect 58560 2215 58590 2245
rect 58670 2215 58700 2245
rect 58780 2215 58810 2245
rect 58890 2215 58920 2245
rect 58395 2170 58425 2200
rect 58505 2170 58535 2200
rect 58615 2170 58645 2200
rect 58725 2170 58755 2200
rect 58835 2170 58865 2200
rect 58395 1940 58425 1945
rect 58395 1920 58400 1940
rect 58400 1920 58420 1940
rect 58420 1920 58425 1940
rect 58395 1915 58425 1920
rect 58505 1940 58535 1945
rect 58505 1920 58510 1940
rect 58510 1920 58530 1940
rect 58530 1920 58535 1940
rect 58505 1915 58535 1920
rect 58615 1940 58645 1945
rect 58615 1920 58620 1940
rect 58620 1920 58640 1940
rect 58640 1920 58645 1940
rect 58615 1915 58645 1920
rect 58725 1940 58755 1945
rect 58725 1920 58730 1940
rect 58730 1920 58750 1940
rect 58750 1920 58755 1940
rect 58725 1915 58755 1920
rect 58835 1940 58865 1945
rect 58835 1920 58840 1940
rect 58840 1920 58860 1940
rect 58860 1920 58865 1940
rect 58835 1915 58865 1920
rect 59085 1915 59115 1945
rect 58085 1850 58115 1880
rect 58125 1850 58155 1880
rect 58165 1850 58195 1880
rect 58085 1810 58115 1840
rect 58125 1810 58155 1840
rect 58165 1810 58195 1840
rect 58450 1875 58480 1880
rect 58450 1855 58455 1875
rect 58455 1855 58475 1875
rect 58475 1855 58480 1875
rect 58450 1850 58480 1855
rect 58450 1835 58480 1840
rect 58450 1815 58455 1835
rect 58455 1815 58475 1835
rect 58475 1815 58480 1835
rect 58450 1810 58480 1815
rect 58395 1730 58425 1760
rect 58505 1730 58535 1760
rect 58615 1730 58645 1760
rect 58725 1730 58755 1760
rect 58835 1730 58865 1760
rect 59040 1730 59070 1760
rect 58395 1390 58425 1420
rect 58505 1390 58535 1420
rect 58615 1390 58645 1420
rect 58725 1390 58755 1420
rect 58835 1390 58865 1420
rect 58015 1345 58045 1375
rect 58340 1345 58370 1375
rect 58450 1345 58480 1375
rect 58560 1345 58590 1375
rect 58670 1345 58700 1375
rect 58780 1345 58810 1375
rect 58890 1345 58920 1375
rect 59040 1360 59070 1390
rect 59650 2215 59680 2245
rect 59375 1680 59405 1710
rect 59425 1680 59455 1710
rect 59475 1680 59505 1710
rect 59525 1680 59555 1710
rect 59575 1680 59605 1710
rect 59375 1630 59405 1660
rect 59425 1630 59455 1660
rect 59475 1630 59505 1660
rect 59525 1630 59555 1660
rect 59575 1630 59605 1660
rect 59375 1580 59405 1610
rect 59425 1580 59455 1610
rect 59475 1580 59505 1610
rect 59525 1580 59555 1610
rect 59575 1580 59605 1610
rect 59125 1390 59160 1395
rect 59125 1365 59130 1390
rect 59130 1365 59155 1390
rect 59155 1365 59160 1390
rect 59125 1360 59160 1365
rect 59185 1390 59220 1395
rect 59185 1365 59190 1390
rect 59190 1365 59215 1390
rect 59215 1365 59220 1390
rect 59185 1360 59220 1365
rect 59245 1390 59280 1395
rect 59245 1365 59250 1390
rect 59250 1365 59275 1390
rect 59275 1365 59280 1390
rect 59245 1360 59280 1365
rect 59305 1390 59340 1395
rect 59305 1365 59310 1390
rect 59310 1365 59335 1390
rect 59335 1365 59340 1390
rect 59305 1360 59340 1365
rect 57935 1300 57965 1330
rect 58285 1300 58315 1330
rect 58945 1300 58975 1330
rect 59085 1305 59115 1335
rect 59185 1305 59215 1335
rect 57395 1110 57425 1115
rect 57395 1090 57400 1110
rect 57400 1090 57420 1110
rect 57420 1090 57425 1110
rect 57395 1085 57425 1090
rect 57870 1085 57900 1115
rect 56445 1030 56475 1060
rect 56555 1030 56585 1060
rect 56665 1030 56695 1060
rect 56775 1030 56805 1060
rect 56885 1030 56915 1060
rect 56995 1030 57025 1060
rect 57105 1030 57135 1060
rect 57215 1030 57245 1060
rect 57325 1030 57355 1060
rect 57435 1030 57465 1060
rect 56225 735 56255 740
rect 56225 715 56230 735
rect 56230 715 56250 735
rect 56250 715 56255 735
rect 56225 710 56255 715
rect 56280 710 56310 740
rect 56390 710 56420 740
rect 56500 710 56530 740
rect 56610 710 56640 740
rect 56720 710 56750 740
rect 56830 710 56860 740
rect 56940 710 56970 740
rect 57050 710 57080 740
rect 57160 710 57190 740
rect 57270 710 57300 740
rect 57380 710 57410 740
rect 59305 1255 59335 1285
rect 58585 1235 58615 1240
rect 58585 1215 58590 1235
rect 58590 1215 58610 1235
rect 58610 1215 58615 1235
rect 58585 1210 58615 1215
rect 59170 1210 59200 1240
rect 58435 1155 58465 1185
rect 58475 1155 58505 1185
rect 58515 1155 58545 1185
rect 58555 1155 58585 1185
rect 58595 1155 58625 1185
rect 58635 1155 58665 1185
rect 58675 1155 58705 1185
rect 58715 1155 58745 1185
rect 58755 1155 58785 1185
rect 58795 1155 58825 1185
rect 58835 1155 58865 1185
rect 58435 1115 58465 1145
rect 58475 1115 58505 1145
rect 58515 1115 58545 1145
rect 58555 1115 58585 1145
rect 58595 1115 58625 1145
rect 58635 1115 58665 1145
rect 58675 1115 58705 1145
rect 58715 1115 58745 1145
rect 58755 1115 58785 1145
rect 58795 1115 58825 1145
rect 58835 1115 58865 1145
rect 58435 1075 58465 1105
rect 58475 1075 58505 1105
rect 58515 1075 58545 1105
rect 58555 1075 58585 1105
rect 58595 1075 58625 1105
rect 58635 1075 58665 1105
rect 58675 1075 58705 1105
rect 58715 1075 58745 1105
rect 58755 1075 58785 1105
rect 58795 1075 58825 1105
rect 58835 1075 58865 1105
rect 59105 1155 59135 1185
rect 59105 1115 59135 1145
rect 59105 1075 59135 1105
rect 57490 735 57520 740
rect 57490 715 57495 735
rect 57495 715 57515 735
rect 57515 715 57520 735
rect 57490 710 57520 715
rect 57935 710 57965 740
rect 56445 665 56475 695
rect 56555 665 56585 695
rect 56665 665 56695 695
rect 56775 665 56805 695
rect 56885 665 56915 695
rect 56995 665 57025 695
rect 57105 665 57135 695
rect 57215 665 57245 695
rect 57325 665 57355 695
rect 57435 665 57465 695
rect 56545 610 56575 640
rect 56655 610 56685 640
rect 56875 610 56905 640
rect 55900 565 55930 595
rect 56490 565 56520 595
rect 56600 590 56630 595
rect 56600 570 56605 590
rect 56605 570 56625 590
rect 56625 570 56630 590
rect 56600 565 56630 570
rect 56545 360 56575 390
rect 56710 565 56740 595
rect 56655 360 56685 390
rect 57045 590 57075 595
rect 57045 570 57050 590
rect 57050 570 57070 590
rect 57070 570 57075 590
rect 57045 565 57075 570
rect 56875 360 56905 390
rect 56490 315 56520 345
rect 56600 315 56630 345
rect 56710 315 56740 345
rect 58435 320 58465 350
rect 58635 320 58665 350
rect 59370 1155 59400 1185
rect 59410 1155 59440 1185
rect 59455 1155 59485 1185
rect 59495 1155 59525 1185
rect 59540 1155 59570 1185
rect 59580 1155 59610 1185
rect 59370 1115 59400 1145
rect 59410 1115 59440 1145
rect 59455 1115 59485 1145
rect 59495 1115 59525 1145
rect 59540 1115 59570 1145
rect 59580 1115 59610 1145
rect 59370 1075 59400 1105
rect 59410 1075 59440 1105
rect 59455 1075 59485 1105
rect 59495 1075 59525 1105
rect 59540 1075 59570 1105
rect 59580 1075 59610 1105
rect 59105 1045 59140 1050
rect 59105 1020 59110 1045
rect 59110 1020 59135 1045
rect 59135 1020 59140 1045
rect 59105 1015 59140 1020
rect 59165 1045 59200 1050
rect 59165 1020 59170 1045
rect 59170 1020 59195 1045
rect 59195 1020 59200 1045
rect 59165 1015 59200 1020
rect 58835 320 58865 350
rect 52645 15 52675 45
rect 52685 15 52715 45
rect 52725 15 52755 45
rect 52995 15 53025 45
rect 53035 15 53065 45
rect 53075 15 53105 45
rect 53345 15 53375 45
rect 53385 15 53415 45
rect 53425 15 53455 45
rect 53695 15 53725 45
rect 53735 15 53765 45
rect 53775 15 53805 45
rect 54045 15 54075 45
rect 54085 15 54115 45
rect 54125 15 54155 45
rect 54395 15 54425 45
rect 54435 15 54465 45
rect 54475 15 54505 45
rect 54745 15 54775 45
rect 54785 15 54815 45
rect 54825 15 54855 45
rect 55035 15 55065 45
rect 55095 15 55125 45
rect 55135 15 55165 45
rect 55175 15 55205 45
rect 55235 15 55265 45
rect 55445 15 55475 45
rect 55485 15 55515 45
rect 55525 15 55555 45
rect 55795 15 55825 45
rect 55835 15 55865 45
rect 55875 15 55905 45
rect 56145 15 56175 45
rect 56185 15 56215 45
rect 56225 15 56255 45
rect 56435 15 56465 45
rect 56495 15 56525 45
rect 56535 15 56565 45
rect 56575 15 56605 45
rect 56765 15 56795 45
rect 56845 15 56875 45
rect 56885 15 56915 45
rect 56925 15 56955 45
rect 57195 15 57225 45
rect 57235 15 57265 45
rect 57275 15 57305 45
rect 57545 15 57575 45
rect 57585 15 57615 45
rect 57625 15 57655 45
rect 57895 15 57925 45
rect 57935 15 57965 45
rect 57975 15 58005 45
rect 58245 15 58275 45
rect 58285 15 58315 45
rect 58325 15 58355 45
rect 58535 15 58565 45
rect 58595 15 58625 45
rect 58635 15 58665 45
rect 58675 15 58705 45
rect 58735 15 58765 45
rect 58945 15 58975 45
rect 58985 15 59015 45
rect 59025 15 59055 45
rect 59295 15 59325 45
rect 59335 15 59365 45
rect 59375 15 59405 45
rect 59645 15 59675 45
rect 59685 15 59715 45
rect 59725 15 59755 45
rect 59995 15 60025 45
rect 60035 15 60065 45
rect 60075 15 60105 45
rect 60345 15 60375 45
rect 60385 15 60415 45
rect 60425 15 60455 45
rect 60695 15 60725 45
rect 60735 15 60765 45
rect 60775 15 60805 45
rect 61045 15 61075 45
rect 61085 15 61115 45
rect 61125 15 61155 45
<< metal2 >>
rect 56205 5020 56245 5025
rect 56205 4990 56210 5020
rect 56240 5015 56245 5020
rect 56675 5020 56715 5025
rect 56675 5015 56680 5020
rect 56240 4995 56680 5015
rect 56240 4990 56245 4995
rect 56205 4985 56245 4990
rect 56675 4990 56680 4995
rect 56710 4990 56715 5020
rect 56675 4985 56715 4990
rect 57085 5020 57125 5025
rect 57085 4990 57090 5020
rect 57120 5015 57125 5020
rect 57555 5020 57595 5025
rect 57555 5015 57560 5020
rect 57120 4995 57560 5015
rect 57120 4990 57125 4995
rect 57085 4985 57125 4990
rect 57555 4990 57560 4995
rect 57590 4990 57595 5020
rect 57555 4985 57595 4990
rect 56085 4965 56125 4970
rect 56085 4935 56090 4965
rect 56120 4960 56125 4965
rect 56205 4965 56245 4970
rect 56205 4960 56210 4965
rect 56120 4940 56210 4960
rect 56120 4935 56125 4940
rect 56085 4930 56125 4935
rect 56205 4935 56210 4940
rect 56240 4960 56245 4965
rect 56265 4965 56305 4970
rect 56265 4960 56270 4965
rect 56240 4940 56270 4960
rect 56240 4935 56245 4940
rect 56205 4930 56245 4935
rect 56265 4935 56270 4940
rect 56300 4935 56305 4965
rect 56265 4930 56305 4935
rect 56880 4965 56920 4970
rect 56880 4935 56885 4965
rect 56915 4960 56920 4965
rect 57025 4965 57065 4970
rect 57025 4960 57030 4965
rect 56915 4940 57030 4960
rect 56915 4935 56920 4940
rect 56880 4930 56920 4935
rect 57025 4935 57030 4940
rect 57060 4960 57065 4965
rect 57145 4965 57185 4970
rect 57145 4960 57150 4965
rect 57060 4940 57150 4960
rect 57060 4935 57065 4940
rect 57025 4930 57065 4935
rect 57145 4935 57150 4940
rect 57180 4960 57185 4965
rect 57205 4965 57245 4970
rect 57205 4960 57210 4965
rect 57180 4940 57210 4960
rect 57180 4935 57185 4940
rect 57145 4930 57185 4935
rect 57205 4935 57210 4940
rect 57240 4935 57245 4965
rect 57205 4930 57245 4935
rect 57495 4965 57535 4970
rect 57495 4935 57500 4965
rect 57530 4960 57535 4965
rect 57555 4965 57595 4970
rect 57555 4960 57560 4965
rect 57530 4940 57560 4960
rect 57530 4935 57535 4940
rect 57495 4930 57535 4935
rect 57555 4935 57560 4940
rect 57590 4960 57595 4965
rect 57675 4965 57715 4970
rect 57675 4960 57680 4965
rect 57590 4940 57680 4960
rect 57590 4935 57595 4940
rect 57555 4930 57595 4935
rect 57675 4935 57680 4940
rect 57710 4935 57715 4965
rect 57675 4930 57715 4935
rect 56555 4795 56595 4800
rect 56555 4765 56560 4795
rect 56590 4790 56595 4795
rect 56615 4795 56655 4800
rect 56615 4790 56620 4795
rect 56590 4770 56620 4790
rect 56590 4765 56595 4770
rect 56555 4760 56595 4765
rect 56615 4765 56620 4770
rect 56650 4790 56655 4795
rect 56735 4795 56775 4800
rect 56735 4790 56740 4795
rect 56650 4770 56740 4790
rect 56650 4765 56655 4770
rect 56615 4760 56655 4765
rect 56735 4765 56740 4770
rect 56770 4790 56775 4795
rect 56880 4795 56920 4800
rect 56880 4790 56885 4795
rect 56770 4770 56885 4790
rect 56770 4765 56775 4770
rect 56735 4760 56775 4765
rect 56880 4765 56885 4770
rect 56915 4765 56920 4795
rect 56880 4760 56920 4765
rect 56205 4560 56245 4565
rect 56205 4530 56210 4560
rect 56240 4555 56245 4560
rect 56675 4560 56715 4565
rect 56675 4555 56680 4560
rect 56240 4535 56680 4555
rect 56240 4530 56245 4535
rect 56205 4525 56245 4530
rect 56675 4530 56680 4535
rect 56710 4530 56715 4560
rect 56675 4525 56715 4530
rect 57085 4560 57125 4565
rect 57085 4530 57090 4560
rect 57120 4555 57125 4560
rect 57555 4560 57595 4565
rect 57555 4555 57560 4560
rect 57120 4535 57560 4555
rect 57120 4530 57125 4535
rect 57085 4525 57125 4530
rect 57555 4530 57560 4535
rect 57590 4530 57595 4560
rect 57555 4525 57595 4530
rect 56150 4515 56190 4520
rect 56150 4485 56155 4515
rect 56185 4510 56190 4515
rect 56630 4515 56660 4520
rect 56185 4490 56630 4510
rect 56185 4485 56190 4490
rect 56150 4480 56190 4485
rect 56825 4515 56865 4520
rect 56825 4510 56830 4515
rect 56660 4490 56830 4510
rect 56630 4480 56660 4485
rect 56825 4485 56830 4490
rect 56860 4510 56865 4515
rect 56860 4505 57606 4510
rect 56860 4490 57576 4505
rect 56860 4485 56865 4490
rect 56825 4480 56865 4485
rect 57576 4470 57606 4475
rect 56935 4460 56975 4465
rect 56935 4430 56940 4460
rect 56970 4445 56975 4460
rect 57135 4450 57175 4455
rect 57135 4445 57140 4450
rect 56970 4430 57140 4445
rect 56935 4425 57140 4430
rect 57135 4420 57140 4425
rect 57170 4445 57175 4450
rect 57615 4450 57655 4455
rect 57615 4445 57620 4450
rect 57170 4425 57620 4445
rect 57170 4420 57175 4425
rect 57135 4415 57175 4420
rect 57615 4420 57620 4425
rect 57650 4420 57655 4450
rect 57615 4415 57655 4420
rect 52640 4305 61160 4310
rect 52640 4275 52645 4305
rect 52675 4275 52685 4305
rect 52715 4275 52725 4305
rect 52755 4275 52995 4305
rect 53025 4275 53035 4305
rect 53065 4275 53075 4305
rect 53105 4275 53345 4305
rect 53375 4275 53385 4305
rect 53415 4275 53425 4305
rect 53455 4275 53695 4305
rect 53725 4275 53735 4305
rect 53765 4275 53775 4305
rect 53805 4275 54045 4305
rect 54075 4275 54085 4305
rect 54115 4275 54125 4305
rect 54155 4275 54395 4305
rect 54425 4275 54435 4305
rect 54465 4275 54475 4305
rect 54505 4275 54745 4305
rect 54775 4275 54785 4305
rect 54815 4275 54825 4305
rect 54855 4275 55095 4305
rect 55125 4275 55135 4305
rect 55165 4275 55175 4305
rect 55205 4275 55285 4305
rect 55315 4275 55445 4305
rect 55475 4275 55485 4305
rect 55515 4275 55525 4305
rect 55555 4275 55755 4305
rect 55785 4275 55795 4305
rect 55825 4275 55835 4305
rect 55865 4275 55875 4305
rect 55905 4275 56885 4305
rect 56915 4275 57895 4305
rect 57925 4275 57935 4305
rect 57965 4275 57975 4305
rect 58005 4275 58015 4305
rect 58045 4275 58245 4305
rect 58275 4275 58285 4305
rect 58315 4275 58325 4305
rect 58355 4275 58485 4305
rect 58515 4275 58595 4305
rect 58625 4275 58635 4305
rect 58665 4275 58675 4305
rect 58705 4275 58945 4305
rect 58975 4275 58985 4305
rect 59015 4275 59025 4305
rect 59055 4275 59295 4305
rect 59325 4275 59335 4305
rect 59365 4275 59375 4305
rect 59405 4275 59645 4305
rect 59675 4275 59685 4305
rect 59715 4275 59725 4305
rect 59755 4275 59995 4305
rect 60025 4275 60035 4305
rect 60065 4275 60075 4305
rect 60105 4275 60345 4305
rect 60375 4275 60385 4305
rect 60415 4275 60425 4305
rect 60455 4275 60695 4305
rect 60725 4275 60735 4305
rect 60765 4275 60775 4305
rect 60805 4275 61045 4305
rect 61075 4275 61085 4305
rect 61115 4275 61125 4305
rect 61155 4275 61160 4305
rect 52640 4270 61160 4275
rect 54980 4210 56765 4215
rect 54980 4180 54985 4210
rect 55015 4180 55025 4210
rect 55055 4180 55065 4210
rect 55095 4180 55105 4210
rect 55135 4180 55145 4210
rect 55175 4180 55185 4210
rect 55215 4180 55225 4210
rect 55255 4180 55345 4210
rect 55375 4180 55385 4210
rect 55415 4180 55425 4210
rect 55455 4180 55465 4210
rect 55495 4180 55505 4210
rect 55535 4180 55545 4210
rect 55575 4180 55585 4210
rect 55615 4180 56010 4210
rect 56040 4180 56050 4210
rect 56080 4180 56090 4210
rect 56120 4180 56130 4210
rect 56160 4180 56170 4210
rect 56200 4180 56210 4210
rect 56240 4180 56250 4210
rect 56280 4180 56290 4210
rect 56320 4180 56330 4210
rect 56360 4180 56370 4210
rect 56400 4180 56410 4210
rect 56440 4180 56450 4210
rect 56480 4180 56490 4210
rect 56520 4180 56530 4210
rect 56560 4180 56570 4210
rect 56600 4180 56610 4210
rect 56640 4180 56650 4210
rect 56680 4180 56690 4210
rect 56720 4180 56730 4210
rect 56760 4180 56765 4210
rect 54980 4170 56765 4180
rect 54980 4140 54985 4170
rect 55015 4140 55025 4170
rect 55055 4140 55065 4170
rect 55095 4140 55105 4170
rect 55135 4140 55145 4170
rect 55175 4140 55185 4170
rect 55215 4140 55225 4170
rect 55255 4140 55345 4170
rect 55375 4140 55385 4170
rect 55415 4140 55425 4170
rect 55455 4140 55465 4170
rect 55495 4140 55505 4170
rect 55535 4140 55545 4170
rect 55575 4140 55585 4170
rect 55615 4140 56010 4170
rect 56040 4140 56050 4170
rect 56080 4140 56090 4170
rect 56120 4140 56130 4170
rect 56160 4140 56170 4170
rect 56200 4140 56210 4170
rect 56240 4140 56250 4170
rect 56280 4140 56290 4170
rect 56320 4140 56330 4170
rect 56360 4140 56370 4170
rect 56400 4140 56410 4170
rect 56440 4140 56450 4170
rect 56480 4140 56490 4170
rect 56520 4140 56530 4170
rect 56560 4140 56570 4170
rect 56600 4140 56610 4170
rect 56640 4140 56650 4170
rect 56680 4140 56690 4170
rect 56720 4140 56730 4170
rect 56760 4140 56765 4170
rect 54980 4130 56765 4140
rect 54980 4100 54985 4130
rect 55015 4100 55025 4130
rect 55055 4100 55065 4130
rect 55095 4100 55105 4130
rect 55135 4100 55145 4130
rect 55175 4100 55185 4130
rect 55215 4100 55225 4130
rect 55255 4100 55345 4130
rect 55375 4100 55385 4130
rect 55415 4100 55425 4130
rect 55455 4100 55465 4130
rect 55495 4100 55505 4130
rect 55535 4100 55545 4130
rect 55575 4100 55585 4130
rect 55615 4100 56010 4130
rect 56040 4100 56050 4130
rect 56080 4100 56090 4130
rect 56120 4100 56130 4130
rect 56160 4100 56170 4130
rect 56200 4100 56210 4130
rect 56240 4100 56250 4130
rect 56280 4100 56290 4130
rect 56320 4100 56330 4130
rect 56360 4100 56370 4130
rect 56400 4100 56410 4130
rect 56440 4100 56450 4130
rect 56480 4100 56490 4130
rect 56520 4100 56530 4130
rect 56560 4100 56570 4130
rect 56600 4100 56610 4130
rect 56640 4100 56650 4130
rect 56680 4100 56690 4130
rect 56720 4100 56730 4130
rect 56760 4100 56765 4130
rect 54980 4095 56765 4100
rect 57035 4210 58820 4215
rect 57035 4180 57040 4210
rect 57070 4180 57080 4210
rect 57110 4180 57120 4210
rect 57150 4180 57160 4210
rect 57190 4180 57200 4210
rect 57230 4180 57240 4210
rect 57270 4180 57280 4210
rect 57310 4180 57320 4210
rect 57350 4180 57360 4210
rect 57390 4180 57400 4210
rect 57430 4180 57440 4210
rect 57470 4180 57480 4210
rect 57510 4180 57520 4210
rect 57550 4180 57560 4210
rect 57590 4180 57600 4210
rect 57630 4180 57640 4210
rect 57670 4180 57680 4210
rect 57710 4180 57720 4210
rect 57750 4180 57760 4210
rect 57790 4180 58185 4210
rect 58215 4180 58225 4210
rect 58255 4180 58265 4210
rect 58295 4180 58305 4210
rect 58335 4180 58345 4210
rect 58375 4180 58385 4210
rect 58415 4180 58425 4210
rect 58455 4180 58545 4210
rect 58575 4180 58585 4210
rect 58615 4180 58625 4210
rect 58655 4180 58665 4210
rect 58695 4180 58705 4210
rect 58735 4180 58745 4210
rect 58775 4180 58785 4210
rect 58815 4180 58820 4210
rect 57035 4170 58820 4180
rect 57035 4140 57040 4170
rect 57070 4140 57080 4170
rect 57110 4140 57120 4170
rect 57150 4140 57160 4170
rect 57190 4140 57200 4170
rect 57230 4140 57240 4170
rect 57270 4140 57280 4170
rect 57310 4140 57320 4170
rect 57350 4140 57360 4170
rect 57390 4140 57400 4170
rect 57430 4140 57440 4170
rect 57470 4140 57480 4170
rect 57510 4140 57520 4170
rect 57550 4140 57560 4170
rect 57590 4140 57600 4170
rect 57630 4140 57640 4170
rect 57670 4140 57680 4170
rect 57710 4140 57720 4170
rect 57750 4140 57760 4170
rect 57790 4140 58185 4170
rect 58215 4140 58225 4170
rect 58255 4140 58265 4170
rect 58295 4140 58305 4170
rect 58335 4140 58345 4170
rect 58375 4140 58385 4170
rect 58415 4140 58425 4170
rect 58455 4140 58545 4170
rect 58575 4140 58585 4170
rect 58615 4140 58625 4170
rect 58655 4140 58665 4170
rect 58695 4140 58705 4170
rect 58735 4140 58745 4170
rect 58775 4140 58785 4170
rect 58815 4140 58820 4170
rect 57035 4130 58820 4140
rect 57035 4100 57040 4130
rect 57070 4100 57080 4130
rect 57110 4100 57120 4130
rect 57150 4100 57160 4130
rect 57190 4100 57200 4130
rect 57230 4100 57240 4130
rect 57270 4100 57280 4130
rect 57310 4100 57320 4130
rect 57350 4100 57360 4130
rect 57390 4100 57400 4130
rect 57430 4100 57440 4130
rect 57470 4100 57480 4130
rect 57510 4100 57520 4130
rect 57550 4100 57560 4130
rect 57590 4100 57600 4130
rect 57630 4100 57640 4130
rect 57670 4100 57680 4130
rect 57710 4100 57720 4130
rect 57750 4100 57760 4130
rect 57790 4100 58185 4130
rect 58215 4100 58225 4130
rect 58255 4100 58265 4130
rect 58295 4100 58305 4130
rect 58335 4100 58345 4130
rect 58375 4100 58385 4130
rect 58415 4100 58425 4130
rect 58455 4100 58545 4130
rect 58575 4100 58585 4130
rect 58615 4100 58625 4130
rect 58655 4100 58665 4130
rect 58695 4100 58705 4130
rect 58735 4100 58745 4130
rect 58775 4100 58785 4130
rect 58815 4100 58820 4130
rect 57035 4095 58820 4100
rect 54920 4075 54960 4080
rect 54920 4045 54925 4075
rect 54955 4070 54960 4075
rect 55040 4075 55080 4080
rect 55040 4070 55045 4075
rect 54955 4050 55045 4070
rect 54955 4045 54960 4050
rect 54920 4040 54960 4045
rect 55040 4045 55045 4050
rect 55075 4070 55080 4075
rect 55160 4075 55200 4080
rect 55160 4070 55165 4075
rect 55075 4050 55165 4070
rect 55075 4045 55080 4050
rect 55040 4040 55080 4045
rect 55160 4045 55165 4050
rect 55195 4070 55200 4075
rect 55280 4075 55320 4080
rect 55280 4070 55285 4075
rect 55195 4050 55285 4070
rect 55195 4045 55200 4050
rect 55160 4040 55200 4045
rect 55280 4045 55285 4050
rect 55315 4070 55320 4075
rect 55400 4075 55440 4080
rect 55400 4070 55405 4075
rect 55315 4050 55405 4070
rect 55315 4045 55320 4050
rect 55280 4040 55320 4045
rect 55400 4045 55405 4050
rect 55435 4070 55440 4075
rect 55520 4075 55560 4080
rect 55520 4070 55525 4075
rect 55435 4050 55525 4070
rect 55435 4045 55440 4050
rect 55400 4040 55440 4045
rect 55520 4045 55525 4050
rect 55555 4070 55560 4075
rect 55640 4075 55680 4080
rect 55640 4070 55645 4075
rect 55555 4050 55645 4070
rect 55555 4045 55560 4050
rect 55520 4040 55560 4045
rect 55640 4045 55645 4050
rect 55675 4045 55680 4075
rect 55640 4040 55680 4045
rect 56065 4075 56105 4080
rect 56065 4045 56070 4075
rect 56100 4070 56105 4075
rect 56185 4075 56225 4080
rect 56185 4070 56190 4075
rect 56100 4050 56190 4070
rect 56100 4045 56105 4050
rect 56065 4040 56105 4045
rect 56185 4045 56190 4050
rect 56220 4070 56225 4075
rect 56305 4075 56345 4080
rect 56305 4070 56310 4075
rect 56220 4050 56310 4070
rect 56220 4045 56225 4050
rect 56185 4040 56225 4045
rect 56305 4045 56310 4050
rect 56340 4070 56345 4075
rect 56425 4075 56465 4080
rect 56425 4070 56430 4075
rect 56340 4050 56430 4070
rect 56340 4045 56345 4050
rect 56305 4040 56345 4045
rect 56425 4045 56430 4050
rect 56460 4070 56465 4075
rect 56545 4075 56585 4080
rect 56545 4070 56550 4075
rect 56460 4050 56550 4070
rect 56460 4045 56465 4050
rect 56425 4040 56465 4045
rect 56545 4045 56550 4050
rect 56580 4070 56585 4075
rect 56665 4075 56705 4080
rect 56665 4070 56670 4075
rect 56580 4050 56670 4070
rect 56580 4045 56585 4050
rect 56545 4040 56585 4045
rect 56665 4045 56670 4050
rect 56700 4045 56705 4075
rect 56665 4040 56705 4045
rect 57095 4075 57135 4080
rect 57095 4045 57100 4075
rect 57130 4070 57135 4075
rect 57215 4075 57255 4080
rect 57215 4070 57220 4075
rect 57130 4050 57220 4070
rect 57130 4045 57135 4050
rect 57095 4040 57135 4045
rect 57215 4045 57220 4050
rect 57250 4070 57255 4075
rect 57335 4075 57375 4080
rect 57335 4070 57340 4075
rect 57250 4050 57340 4070
rect 57250 4045 57255 4050
rect 57215 4040 57255 4045
rect 57335 4045 57340 4050
rect 57370 4070 57375 4075
rect 57455 4075 57495 4080
rect 57455 4070 57460 4075
rect 57370 4050 57460 4070
rect 57370 4045 57375 4050
rect 57335 4040 57375 4045
rect 57455 4045 57460 4050
rect 57490 4070 57495 4075
rect 57575 4075 57615 4080
rect 57575 4070 57580 4075
rect 57490 4050 57580 4070
rect 57490 4045 57495 4050
rect 57455 4040 57495 4045
rect 57575 4045 57580 4050
rect 57610 4070 57615 4075
rect 57695 4075 57735 4080
rect 57695 4070 57700 4075
rect 57610 4050 57700 4070
rect 57610 4045 57615 4050
rect 57575 4040 57615 4045
rect 57695 4045 57700 4050
rect 57730 4045 57735 4075
rect 57695 4040 57735 4045
rect 58120 4075 58160 4080
rect 58120 4045 58125 4075
rect 58155 4070 58160 4075
rect 58240 4075 58280 4080
rect 58240 4070 58245 4075
rect 58155 4050 58245 4070
rect 58155 4045 58160 4050
rect 58120 4040 58160 4045
rect 58240 4045 58245 4050
rect 58275 4070 58280 4075
rect 58360 4075 58400 4080
rect 58360 4070 58365 4075
rect 58275 4050 58365 4070
rect 58275 4045 58280 4050
rect 58240 4040 58280 4045
rect 58360 4045 58365 4050
rect 58395 4070 58400 4075
rect 58480 4075 58520 4080
rect 58480 4070 58485 4075
rect 58395 4050 58485 4070
rect 58395 4045 58400 4050
rect 58360 4040 58400 4045
rect 58480 4045 58485 4050
rect 58515 4070 58520 4075
rect 58600 4075 58640 4080
rect 58600 4070 58605 4075
rect 58515 4050 58605 4070
rect 58515 4045 58520 4050
rect 58480 4040 58520 4045
rect 58600 4045 58605 4050
rect 58635 4070 58640 4075
rect 58720 4075 58760 4080
rect 58720 4070 58725 4075
rect 58635 4050 58725 4070
rect 58635 4045 58640 4050
rect 58600 4040 58640 4045
rect 58720 4045 58725 4050
rect 58755 4070 58760 4075
rect 58840 4075 58880 4080
rect 58840 4070 58845 4075
rect 58755 4050 58845 4070
rect 58755 4045 58760 4050
rect 58720 4040 58760 4045
rect 58840 4045 58845 4050
rect 58875 4045 58880 4075
rect 58840 4040 58880 4045
rect 54980 3685 55020 3690
rect 54980 3655 54985 3685
rect 55015 3680 55020 3685
rect 55100 3685 55140 3690
rect 55100 3680 55105 3685
rect 55015 3660 55105 3680
rect 55015 3655 55020 3660
rect 54980 3650 55020 3655
rect 55100 3655 55105 3660
rect 55135 3680 55140 3685
rect 55220 3685 55260 3690
rect 55220 3680 55225 3685
rect 55135 3660 55225 3680
rect 55135 3655 55140 3660
rect 55100 3650 55140 3655
rect 55220 3655 55225 3660
rect 55255 3680 55260 3685
rect 55340 3685 55380 3690
rect 55340 3680 55345 3685
rect 55255 3660 55345 3680
rect 55255 3655 55260 3660
rect 55220 3650 55260 3655
rect 55340 3655 55345 3660
rect 55375 3680 55380 3685
rect 55460 3685 55500 3690
rect 55460 3680 55465 3685
rect 55375 3660 55465 3680
rect 55375 3655 55380 3660
rect 55340 3650 55380 3655
rect 55460 3655 55465 3660
rect 55495 3680 55500 3685
rect 55580 3685 55620 3690
rect 55580 3680 55585 3685
rect 55495 3660 55585 3680
rect 55495 3655 55500 3660
rect 55460 3650 55500 3655
rect 55580 3655 55585 3660
rect 55615 3655 55620 3685
rect 55580 3650 55620 3655
rect 56065 3685 56105 3690
rect 56065 3655 56070 3685
rect 56100 3680 56105 3685
rect 56185 3685 56225 3690
rect 56185 3680 56190 3685
rect 56100 3660 56190 3680
rect 56100 3655 56105 3660
rect 56065 3650 56105 3655
rect 56185 3655 56190 3660
rect 56220 3680 56225 3685
rect 56305 3685 56345 3690
rect 56305 3680 56310 3685
rect 56220 3660 56310 3680
rect 56220 3655 56225 3660
rect 56185 3650 56225 3655
rect 56305 3655 56310 3660
rect 56340 3680 56345 3685
rect 56425 3685 56465 3690
rect 56425 3680 56430 3685
rect 56340 3660 56430 3680
rect 56340 3655 56345 3660
rect 56305 3650 56345 3655
rect 56425 3655 56430 3660
rect 56460 3680 56465 3685
rect 56545 3685 56585 3690
rect 56545 3680 56550 3685
rect 56460 3660 56550 3680
rect 56460 3655 56465 3660
rect 56425 3650 56465 3655
rect 56545 3655 56550 3660
rect 56580 3680 56585 3685
rect 56665 3685 56705 3690
rect 56665 3680 56670 3685
rect 56580 3660 56670 3680
rect 56580 3655 56585 3660
rect 56545 3650 56585 3655
rect 56665 3655 56670 3660
rect 56700 3655 56705 3685
rect 56665 3650 56705 3655
rect 57095 3685 57135 3690
rect 57095 3655 57100 3685
rect 57130 3680 57135 3685
rect 57215 3685 57255 3690
rect 57215 3680 57220 3685
rect 57130 3660 57220 3680
rect 57130 3655 57135 3660
rect 57095 3650 57135 3655
rect 57215 3655 57220 3660
rect 57250 3680 57255 3685
rect 57335 3685 57375 3690
rect 57335 3680 57340 3685
rect 57250 3660 57340 3680
rect 57250 3655 57255 3660
rect 57215 3650 57255 3655
rect 57335 3655 57340 3660
rect 57370 3680 57375 3685
rect 57455 3685 57495 3690
rect 57455 3680 57460 3685
rect 57370 3660 57460 3680
rect 57370 3655 57375 3660
rect 57335 3650 57375 3655
rect 57455 3655 57460 3660
rect 57490 3680 57495 3685
rect 57575 3685 57615 3690
rect 57575 3680 57580 3685
rect 57490 3660 57580 3680
rect 57490 3655 57495 3660
rect 57455 3650 57495 3655
rect 57575 3655 57580 3660
rect 57610 3680 57615 3685
rect 57695 3685 57735 3690
rect 57695 3680 57700 3685
rect 57610 3660 57700 3680
rect 57610 3655 57615 3660
rect 57575 3650 57615 3655
rect 57695 3655 57700 3660
rect 57730 3655 57735 3685
rect 57695 3650 57735 3655
rect 58180 3685 58220 3690
rect 58180 3655 58185 3685
rect 58215 3680 58220 3685
rect 58300 3685 58340 3690
rect 58300 3680 58305 3685
rect 58215 3660 58305 3680
rect 58215 3655 58220 3660
rect 58180 3650 58220 3655
rect 58300 3655 58305 3660
rect 58335 3680 58340 3685
rect 58420 3685 58460 3690
rect 58420 3680 58425 3685
rect 58335 3660 58425 3680
rect 58335 3655 58340 3660
rect 58300 3650 58340 3655
rect 58420 3655 58425 3660
rect 58455 3680 58460 3685
rect 58540 3685 58580 3690
rect 58540 3680 58545 3685
rect 58455 3660 58545 3680
rect 58455 3655 58460 3660
rect 58420 3650 58460 3655
rect 58540 3655 58545 3660
rect 58575 3680 58580 3685
rect 58660 3685 58700 3690
rect 58660 3680 58665 3685
rect 58575 3660 58665 3680
rect 58575 3655 58580 3660
rect 58540 3650 58580 3655
rect 58660 3655 58665 3660
rect 58695 3680 58700 3685
rect 58780 3685 58820 3690
rect 58780 3680 58785 3685
rect 58695 3660 58785 3680
rect 58695 3655 58700 3660
rect 58660 3650 58700 3655
rect 58780 3655 58785 3660
rect 58815 3655 58820 3685
rect 58780 3650 58820 3655
rect 56365 3605 56405 3610
rect 56365 3575 56370 3605
rect 56400 3600 56405 3605
rect 56835 3605 56875 3610
rect 56835 3600 56840 3605
rect 56400 3580 56840 3600
rect 56400 3575 56405 3580
rect 56365 3570 56405 3575
rect 56835 3575 56840 3580
rect 56870 3600 56875 3605
rect 57395 3605 57435 3610
rect 57395 3600 57400 3605
rect 56870 3580 57400 3600
rect 56870 3575 56875 3580
rect 56835 3570 56875 3575
rect 57395 3575 57400 3580
rect 57430 3575 57435 3605
rect 57395 3570 57435 3575
rect 55280 3560 55320 3565
rect 55280 3530 55285 3560
rect 55315 3555 55320 3560
rect 56925 3560 56965 3565
rect 56925 3555 56930 3560
rect 55315 3535 56930 3555
rect 55315 3530 55320 3535
rect 55280 3525 55320 3530
rect 56925 3530 56930 3535
rect 56960 3555 56965 3560
rect 58480 3560 58520 3565
rect 58480 3555 58485 3560
rect 56960 3535 58485 3555
rect 56960 3530 56965 3535
rect 56925 3525 56965 3530
rect 58480 3530 58485 3535
rect 58515 3530 58520 3560
rect 58480 3525 58520 3530
rect 55600 3515 56705 3520
rect 55600 3485 55605 3515
rect 55635 3485 55645 3515
rect 55675 3485 55685 3515
rect 55715 3485 56070 3515
rect 56100 3485 56110 3515
rect 56140 3485 56150 3515
rect 56180 3485 56190 3515
rect 56220 3485 56230 3515
rect 56260 3485 56270 3515
rect 56300 3485 56310 3515
rect 56340 3485 56350 3515
rect 56380 3485 56390 3515
rect 56420 3485 56430 3515
rect 56460 3485 56470 3515
rect 56500 3485 56510 3515
rect 56540 3485 56550 3515
rect 56580 3485 56590 3515
rect 56620 3485 56630 3515
rect 56660 3485 56670 3515
rect 56700 3485 56705 3515
rect 55600 3475 56705 3485
rect 55600 3445 55605 3475
rect 55635 3445 55645 3475
rect 55675 3445 55685 3475
rect 55715 3445 56070 3475
rect 56100 3445 56110 3475
rect 56140 3445 56150 3475
rect 56180 3445 56190 3475
rect 56220 3445 56230 3475
rect 56260 3445 56270 3475
rect 56300 3445 56310 3475
rect 56340 3445 56350 3475
rect 56380 3445 56390 3475
rect 56420 3445 56430 3475
rect 56460 3445 56470 3475
rect 56500 3445 56510 3475
rect 56540 3445 56550 3475
rect 56580 3445 56590 3475
rect 56620 3445 56630 3475
rect 56660 3445 56670 3475
rect 56700 3445 56705 3475
rect 55600 3435 56705 3445
rect 55600 3405 55605 3435
rect 55635 3405 55645 3435
rect 55675 3405 55685 3435
rect 55715 3405 56070 3435
rect 56100 3405 56110 3435
rect 56140 3405 56150 3435
rect 56180 3405 56190 3435
rect 56220 3405 56230 3435
rect 56260 3405 56270 3435
rect 56300 3405 56310 3435
rect 56340 3405 56350 3435
rect 56380 3405 56390 3435
rect 56420 3405 56430 3435
rect 56460 3405 56470 3435
rect 56500 3405 56510 3435
rect 56540 3405 56550 3435
rect 56580 3405 56590 3435
rect 56620 3405 56630 3435
rect 56660 3405 56670 3435
rect 56700 3405 56705 3435
rect 54605 3400 54645 3405
rect 55600 3400 56705 3405
rect 57095 3515 58200 3520
rect 57095 3485 57100 3515
rect 57130 3485 57140 3515
rect 57170 3485 57180 3515
rect 57210 3485 57220 3515
rect 57250 3485 57260 3515
rect 57290 3485 57300 3515
rect 57330 3485 57340 3515
rect 57370 3485 57380 3515
rect 57410 3485 57420 3515
rect 57450 3485 57460 3515
rect 57490 3485 57500 3515
rect 57530 3485 57540 3515
rect 57570 3485 57580 3515
rect 57610 3485 57620 3515
rect 57650 3485 57660 3515
rect 57690 3485 57700 3515
rect 57730 3485 58085 3515
rect 58115 3485 58125 3515
rect 58155 3485 58165 3515
rect 58195 3485 58200 3515
rect 57095 3475 58200 3485
rect 57095 3445 57100 3475
rect 57130 3445 57140 3475
rect 57170 3445 57180 3475
rect 57210 3445 57220 3475
rect 57250 3445 57260 3475
rect 57290 3445 57300 3475
rect 57330 3445 57340 3475
rect 57370 3445 57380 3475
rect 57410 3445 57420 3475
rect 57450 3445 57460 3475
rect 57490 3445 57500 3475
rect 57530 3445 57540 3475
rect 57570 3445 57580 3475
rect 57610 3445 57620 3475
rect 57650 3445 57660 3475
rect 57690 3445 57700 3475
rect 57730 3445 58085 3475
rect 58115 3445 58125 3475
rect 58155 3445 58165 3475
rect 58195 3445 58200 3475
rect 57095 3435 58200 3445
rect 57095 3405 57100 3435
rect 57130 3405 57140 3435
rect 57170 3405 57180 3435
rect 57210 3405 57220 3435
rect 57250 3405 57260 3435
rect 57290 3405 57300 3435
rect 57330 3405 57340 3435
rect 57370 3405 57380 3435
rect 57410 3405 57420 3435
rect 57450 3405 57460 3435
rect 57490 3405 57500 3435
rect 57530 3405 57540 3435
rect 57570 3405 57580 3435
rect 57610 3405 57620 3435
rect 57650 3405 57660 3435
rect 57690 3405 57700 3435
rect 57730 3405 58085 3435
rect 58115 3405 58125 3435
rect 58155 3405 58165 3435
rect 58195 3405 58200 3435
rect 57095 3400 58200 3405
rect 59155 3400 59195 3405
rect 54605 3370 54610 3400
rect 54640 3370 54645 3400
rect 54605 3365 54645 3370
rect 54820 3380 54860 3385
rect 54820 3350 54825 3380
rect 54855 3375 54860 3380
rect 54930 3380 54970 3385
rect 54930 3375 54935 3380
rect 54855 3355 54935 3375
rect 54855 3350 54860 3355
rect 54820 3345 54860 3350
rect 54930 3350 54935 3355
rect 54965 3375 54970 3380
rect 55040 3380 55080 3385
rect 55040 3375 55045 3380
rect 54965 3355 55045 3375
rect 54965 3350 54970 3355
rect 54930 3345 54970 3350
rect 55040 3350 55045 3355
rect 55075 3375 55080 3380
rect 55150 3380 55190 3385
rect 55150 3375 55155 3380
rect 55075 3355 55155 3375
rect 55075 3350 55080 3355
rect 55040 3345 55080 3350
rect 55150 3350 55155 3355
rect 55185 3375 55190 3380
rect 55260 3380 55300 3385
rect 55260 3375 55265 3380
rect 55185 3355 55265 3375
rect 55185 3350 55190 3355
rect 55150 3345 55190 3350
rect 55260 3350 55265 3355
rect 55295 3375 55300 3380
rect 55370 3380 55410 3385
rect 55370 3375 55375 3380
rect 55295 3355 55375 3375
rect 55295 3350 55300 3355
rect 55260 3345 55300 3350
rect 55370 3350 55375 3355
rect 55405 3375 55410 3380
rect 55480 3380 55520 3385
rect 55480 3375 55485 3380
rect 55405 3355 55485 3375
rect 55405 3350 55410 3355
rect 55370 3345 55410 3350
rect 55480 3350 55485 3355
rect 55515 3375 55520 3380
rect 55750 3380 55790 3385
rect 55750 3375 55755 3380
rect 55515 3355 55755 3375
rect 55515 3350 55520 3355
rect 55480 3345 55520 3350
rect 55750 3350 55755 3355
rect 55785 3350 55790 3380
rect 55750 3345 55790 3350
rect 56275 3380 56315 3385
rect 56275 3350 56280 3380
rect 56310 3375 56315 3380
rect 56385 3380 56425 3385
rect 56385 3375 56390 3380
rect 56310 3355 56390 3375
rect 56310 3350 56315 3355
rect 56275 3345 56315 3350
rect 56385 3350 56390 3355
rect 56420 3375 56425 3380
rect 56495 3380 56535 3385
rect 56495 3375 56500 3380
rect 56420 3355 56500 3375
rect 56420 3350 56425 3355
rect 56385 3345 56425 3350
rect 56495 3350 56500 3355
rect 56530 3375 56535 3380
rect 56605 3380 56645 3385
rect 56605 3375 56610 3380
rect 56530 3355 56610 3375
rect 56530 3350 56535 3355
rect 56495 3345 56535 3350
rect 56605 3350 56610 3355
rect 56640 3375 56645 3380
rect 56715 3380 56755 3385
rect 56715 3375 56720 3380
rect 56640 3355 56720 3375
rect 56640 3350 56645 3355
rect 56605 3345 56645 3350
rect 56715 3350 56720 3355
rect 56750 3375 56755 3380
rect 56825 3380 56865 3385
rect 56825 3375 56830 3380
rect 56750 3355 56830 3375
rect 56750 3350 56755 3355
rect 56715 3345 56755 3350
rect 56825 3350 56830 3355
rect 56860 3375 56865 3380
rect 56935 3380 56975 3385
rect 56935 3375 56940 3380
rect 56860 3355 56940 3375
rect 56860 3350 56865 3355
rect 56825 3345 56865 3350
rect 56935 3350 56940 3355
rect 56970 3375 56975 3380
rect 57045 3380 57085 3385
rect 57045 3375 57050 3380
rect 56970 3355 57050 3375
rect 56970 3350 56975 3355
rect 56935 3345 56975 3350
rect 57045 3350 57050 3355
rect 57080 3375 57085 3380
rect 57155 3380 57195 3385
rect 57155 3375 57160 3380
rect 57080 3355 57160 3375
rect 57080 3350 57085 3355
rect 57045 3345 57085 3350
rect 57155 3350 57160 3355
rect 57190 3375 57195 3380
rect 57265 3380 57305 3385
rect 57265 3375 57270 3380
rect 57190 3355 57270 3375
rect 57190 3350 57195 3355
rect 57155 3345 57195 3350
rect 57265 3350 57270 3355
rect 57300 3375 57305 3380
rect 57375 3380 57415 3385
rect 57375 3375 57380 3380
rect 57300 3355 57380 3375
rect 57300 3350 57305 3355
rect 57265 3345 57305 3350
rect 57375 3350 57380 3355
rect 57410 3375 57415 3380
rect 57485 3380 57525 3385
rect 57485 3375 57490 3380
rect 57410 3355 57490 3375
rect 57410 3350 57415 3355
rect 57375 3345 57415 3350
rect 57485 3350 57490 3355
rect 57520 3375 57525 3380
rect 58010 3380 58050 3385
rect 58010 3375 58015 3380
rect 57520 3355 58015 3375
rect 57520 3350 57525 3355
rect 57485 3345 57525 3350
rect 58010 3350 58015 3355
rect 58045 3375 58050 3380
rect 58280 3380 58320 3385
rect 58280 3375 58285 3380
rect 58045 3355 58285 3375
rect 58045 3350 58050 3355
rect 58010 3345 58050 3350
rect 58280 3350 58285 3355
rect 58315 3375 58320 3380
rect 58390 3380 58430 3385
rect 58390 3375 58395 3380
rect 58315 3355 58395 3375
rect 58315 3350 58320 3355
rect 58280 3345 58320 3350
rect 58390 3350 58395 3355
rect 58425 3375 58430 3380
rect 58500 3380 58540 3385
rect 58500 3375 58505 3380
rect 58425 3355 58505 3375
rect 58425 3350 58430 3355
rect 58390 3345 58430 3350
rect 58500 3350 58505 3355
rect 58535 3375 58540 3380
rect 58610 3380 58650 3385
rect 58610 3375 58615 3380
rect 58535 3355 58615 3375
rect 58535 3350 58540 3355
rect 58500 3345 58540 3350
rect 58610 3350 58615 3355
rect 58645 3375 58650 3380
rect 58720 3380 58760 3385
rect 58720 3375 58725 3380
rect 58645 3355 58725 3375
rect 58645 3350 58650 3355
rect 58610 3345 58650 3350
rect 58720 3350 58725 3355
rect 58755 3375 58760 3380
rect 58830 3380 58870 3385
rect 58830 3375 58835 3380
rect 58755 3355 58835 3375
rect 58755 3350 58760 3355
rect 58720 3345 58760 3350
rect 58830 3350 58835 3355
rect 58865 3375 58870 3380
rect 58940 3380 58980 3385
rect 58940 3375 58945 3380
rect 58865 3355 58945 3375
rect 58865 3350 58870 3355
rect 58830 3345 58870 3350
rect 58940 3350 58945 3355
rect 58975 3350 58980 3380
rect 59155 3370 59160 3400
rect 59190 3370 59195 3400
rect 59155 3365 59195 3370
rect 58940 3345 58980 3350
rect 56330 3335 56370 3340
rect 56330 3305 56335 3335
rect 56365 3330 56370 3335
rect 56550 3335 56590 3340
rect 56550 3330 56555 3335
rect 56365 3310 56555 3330
rect 56365 3305 56370 3310
rect 54875 3300 54915 3305
rect 54875 3270 54880 3300
rect 54910 3295 54915 3300
rect 54985 3300 55025 3305
rect 54985 3295 54990 3300
rect 54910 3275 54990 3295
rect 54910 3270 54915 3275
rect 54875 3265 54915 3270
rect 54985 3270 54990 3275
rect 55020 3295 55025 3300
rect 55095 3300 55135 3305
rect 55095 3295 55100 3300
rect 55020 3275 55100 3295
rect 55020 3270 55025 3275
rect 54985 3265 55025 3270
rect 55095 3270 55100 3275
rect 55130 3295 55135 3300
rect 55205 3300 55245 3305
rect 55205 3295 55210 3300
rect 55130 3275 55210 3295
rect 55130 3270 55135 3275
rect 55095 3265 55135 3270
rect 55205 3270 55210 3275
rect 55240 3295 55245 3300
rect 55315 3300 55355 3305
rect 55315 3295 55320 3300
rect 55240 3275 55320 3295
rect 55240 3270 55245 3275
rect 55205 3265 55245 3270
rect 55315 3270 55320 3275
rect 55350 3295 55355 3300
rect 55425 3300 55465 3305
rect 56330 3300 56370 3305
rect 56550 3305 56555 3310
rect 56585 3330 56590 3335
rect 56770 3335 56810 3340
rect 56770 3330 56775 3335
rect 56585 3310 56775 3330
rect 56585 3305 56590 3310
rect 56550 3300 56590 3305
rect 56770 3305 56775 3310
rect 56805 3330 56810 3335
rect 56990 3335 57030 3340
rect 56990 3330 56995 3335
rect 56805 3310 56995 3330
rect 56805 3305 56810 3310
rect 56770 3300 56810 3305
rect 56990 3305 56995 3310
rect 57025 3330 57030 3335
rect 57210 3335 57250 3340
rect 57210 3330 57215 3335
rect 57025 3310 57215 3330
rect 57025 3305 57030 3310
rect 56990 3300 57030 3305
rect 57210 3305 57215 3310
rect 57245 3330 57250 3335
rect 57430 3335 57470 3340
rect 57430 3330 57435 3335
rect 57245 3310 57435 3330
rect 57245 3305 57250 3310
rect 57210 3300 57250 3305
rect 57430 3305 57435 3310
rect 57465 3305 57470 3335
rect 57430 3300 57470 3305
rect 58335 3300 58375 3305
rect 55425 3295 55430 3300
rect 55350 3275 55430 3295
rect 55350 3270 55355 3275
rect 55315 3265 55355 3270
rect 55425 3270 55430 3275
rect 55460 3270 55465 3300
rect 55425 3265 55465 3270
rect 56440 3290 56480 3295
rect 56440 3260 56445 3290
rect 56475 3285 56480 3290
rect 56660 3290 56700 3295
rect 56660 3285 56665 3290
rect 56475 3265 56665 3285
rect 56475 3260 56480 3265
rect 56440 3255 56480 3260
rect 56660 3260 56665 3265
rect 56695 3285 56700 3290
rect 56880 3290 56920 3295
rect 56880 3285 56885 3290
rect 56695 3265 56885 3285
rect 56695 3260 56700 3265
rect 56660 3255 56700 3260
rect 56880 3260 56885 3265
rect 56915 3285 56920 3290
rect 57100 3290 57140 3295
rect 57100 3285 57105 3290
rect 56915 3265 57105 3285
rect 56915 3260 56920 3265
rect 56880 3255 56920 3260
rect 57100 3260 57105 3265
rect 57135 3285 57140 3290
rect 57320 3290 57360 3295
rect 57320 3285 57325 3290
rect 57135 3265 57325 3285
rect 57135 3260 57140 3265
rect 57100 3255 57140 3260
rect 57320 3260 57325 3265
rect 57355 3260 57360 3290
rect 58335 3270 58340 3300
rect 58370 3295 58375 3300
rect 58445 3300 58485 3305
rect 58445 3295 58450 3300
rect 58370 3275 58450 3295
rect 58370 3270 58375 3275
rect 58335 3265 58375 3270
rect 58445 3270 58450 3275
rect 58480 3295 58485 3300
rect 58555 3300 58595 3305
rect 58555 3295 58560 3300
rect 58480 3275 58560 3295
rect 58480 3270 58485 3275
rect 58445 3265 58485 3270
rect 58555 3270 58560 3275
rect 58590 3295 58595 3300
rect 58665 3300 58705 3305
rect 58665 3295 58670 3300
rect 58590 3275 58670 3295
rect 58590 3270 58595 3275
rect 58555 3265 58595 3270
rect 58665 3270 58670 3275
rect 58700 3295 58705 3300
rect 58775 3300 58815 3305
rect 58775 3295 58780 3300
rect 58700 3275 58780 3295
rect 58700 3270 58705 3275
rect 58665 3265 58705 3270
rect 58775 3270 58780 3275
rect 58810 3295 58815 3300
rect 58885 3300 58925 3305
rect 58885 3295 58890 3300
rect 58810 3275 58890 3295
rect 58810 3270 58815 3275
rect 58775 3265 58815 3270
rect 58885 3270 58890 3275
rect 58920 3270 58925 3300
rect 58885 3265 58925 3270
rect 57320 3255 57360 3260
rect 56330 3200 56370 3205
rect 56330 3170 56335 3200
rect 56365 3195 56370 3200
rect 56550 3200 56590 3205
rect 56550 3195 56555 3200
rect 56365 3175 56555 3195
rect 56365 3170 56370 3175
rect 56330 3165 56370 3170
rect 56550 3170 56555 3175
rect 56585 3195 56590 3200
rect 56770 3200 56810 3205
rect 56770 3195 56775 3200
rect 56585 3175 56775 3195
rect 56585 3170 56590 3175
rect 56550 3165 56590 3170
rect 56770 3170 56775 3175
rect 56805 3195 56810 3200
rect 56990 3200 57030 3205
rect 56990 3195 56995 3200
rect 56805 3175 56995 3195
rect 56805 3170 56810 3175
rect 56770 3165 56810 3170
rect 56990 3170 56995 3175
rect 57025 3195 57030 3200
rect 57210 3200 57250 3205
rect 57210 3195 57215 3200
rect 57025 3175 57215 3195
rect 57025 3170 57030 3175
rect 56990 3165 57030 3170
rect 57210 3170 57215 3175
rect 57245 3195 57250 3200
rect 57430 3200 57470 3205
rect 57430 3195 57435 3200
rect 57245 3175 57435 3195
rect 57245 3170 57250 3175
rect 57210 3165 57250 3170
rect 57430 3170 57435 3175
rect 57465 3170 57470 3200
rect 57430 3165 57470 3170
rect 56440 3130 56480 3135
rect 56440 3100 56445 3130
rect 56475 3125 56480 3130
rect 56660 3130 56700 3135
rect 56660 3125 56665 3130
rect 56475 3105 56665 3125
rect 56475 3100 56480 3105
rect 56440 3095 56480 3100
rect 56660 3100 56665 3105
rect 56695 3125 56700 3130
rect 56880 3130 56920 3135
rect 56880 3125 56885 3130
rect 56695 3105 56885 3125
rect 56695 3100 56700 3105
rect 56660 3095 56700 3100
rect 56880 3100 56885 3105
rect 56915 3125 56920 3130
rect 57100 3130 57140 3135
rect 57100 3125 57105 3130
rect 56915 3105 57105 3125
rect 56915 3100 56920 3105
rect 56880 3095 56920 3100
rect 57100 3100 57105 3105
rect 57135 3125 57140 3130
rect 57320 3130 57360 3135
rect 57320 3125 57325 3130
rect 57135 3105 57325 3125
rect 57135 3100 57140 3105
rect 57100 3095 57140 3100
rect 57320 3100 57325 3105
rect 57355 3100 57360 3130
rect 57320 3095 57360 3100
rect 56140 3025 56180 3030
rect 55940 3020 55980 3025
rect 55940 2990 55945 3020
rect 55975 3015 55980 3020
rect 56040 3020 56070 3025
rect 55975 2995 56040 3015
rect 55975 2990 55980 2995
rect 55940 2985 55980 2990
rect 56140 2995 56145 3025
rect 56175 3020 56180 3025
rect 56250 3025 56290 3030
rect 56250 3020 56255 3025
rect 56175 3000 56255 3020
rect 56175 2995 56180 3000
rect 56140 2990 56180 2995
rect 56250 2995 56255 3000
rect 56285 3020 56290 3025
rect 56360 3025 56400 3030
rect 56360 3020 56365 3025
rect 56285 3000 56365 3020
rect 56285 2995 56290 3000
rect 56250 2990 56290 2995
rect 56360 2995 56365 3000
rect 56395 3020 56400 3025
rect 56470 3025 56510 3030
rect 56470 3020 56475 3025
rect 56395 3000 56475 3020
rect 56395 2995 56400 3000
rect 56360 2990 56400 2995
rect 56470 2995 56475 3000
rect 56505 3020 56510 3025
rect 56580 3025 56620 3030
rect 57180 3025 57220 3030
rect 56580 3020 56585 3025
rect 56505 3000 56585 3020
rect 56505 2995 56510 3000
rect 56470 2990 56510 2995
rect 56580 2995 56585 3000
rect 56615 2995 56620 3025
rect 56580 2990 56620 2995
rect 56690 3020 56720 3025
rect 57080 3020 57110 3025
rect 56720 2995 57080 3015
rect 56040 2985 56070 2990
rect 56690 2985 56720 2990
rect 57180 2995 57185 3025
rect 57215 3020 57220 3025
rect 57290 3025 57330 3030
rect 57290 3020 57295 3025
rect 57215 3000 57295 3020
rect 57215 2995 57220 3000
rect 57180 2990 57220 2995
rect 57290 2995 57295 3000
rect 57325 3020 57330 3025
rect 57400 3025 57440 3030
rect 57400 3020 57405 3025
rect 57325 3000 57405 3020
rect 57325 2995 57330 3000
rect 57290 2990 57330 2995
rect 57400 2995 57405 3000
rect 57435 3020 57440 3025
rect 57510 3025 57550 3030
rect 57510 3020 57515 3025
rect 57435 3000 57515 3020
rect 57435 2995 57440 3000
rect 57400 2990 57440 2995
rect 57510 2995 57515 3000
rect 57545 3020 57550 3025
rect 57620 3025 57660 3030
rect 57620 3020 57625 3025
rect 57545 3000 57625 3020
rect 57545 2995 57550 3000
rect 57510 2990 57550 2995
rect 57620 2995 57625 3000
rect 57655 2995 57660 3025
rect 57620 2990 57660 2995
rect 57730 3020 57760 3025
rect 57820 3020 57860 3025
rect 57820 3015 57825 3020
rect 57760 2995 57825 3015
rect 57080 2985 57110 2990
rect 57730 2985 57760 2990
rect 57820 2990 57825 2995
rect 57855 2990 57860 3020
rect 57820 2985 57860 2990
rect 56085 2980 56125 2985
rect 56085 2950 56090 2980
rect 56120 2975 56125 2980
rect 56195 2980 56235 2985
rect 56195 2975 56200 2980
rect 56120 2955 56200 2975
rect 56120 2950 56125 2955
rect 56085 2945 56125 2950
rect 56195 2950 56200 2955
rect 56230 2975 56235 2980
rect 56305 2980 56345 2985
rect 56305 2975 56310 2980
rect 56230 2955 56310 2975
rect 56230 2950 56235 2955
rect 56195 2945 56235 2950
rect 56305 2950 56310 2955
rect 56340 2975 56345 2980
rect 56415 2980 56455 2985
rect 56415 2975 56420 2980
rect 56340 2955 56420 2975
rect 56340 2950 56345 2955
rect 56305 2945 56345 2950
rect 56415 2950 56420 2955
rect 56450 2975 56455 2980
rect 56525 2980 56565 2985
rect 56525 2975 56530 2980
rect 56450 2955 56530 2975
rect 56450 2950 56455 2955
rect 56415 2945 56455 2950
rect 56525 2950 56530 2955
rect 56560 2975 56565 2980
rect 56635 2980 56675 2985
rect 56635 2975 56640 2980
rect 56560 2955 56640 2975
rect 56560 2950 56565 2955
rect 56525 2945 56565 2950
rect 56635 2950 56640 2955
rect 56670 2950 56675 2980
rect 56635 2945 56675 2950
rect 57125 2980 57165 2985
rect 57125 2950 57130 2980
rect 57160 2975 57165 2980
rect 57345 2980 57385 2985
rect 57345 2975 57350 2980
rect 57160 2955 57350 2975
rect 57160 2950 57165 2955
rect 57125 2945 57165 2950
rect 57345 2950 57350 2955
rect 57380 2975 57385 2980
rect 57565 2980 57605 2985
rect 57565 2975 57570 2980
rect 57380 2955 57570 2975
rect 57380 2950 57385 2955
rect 57345 2945 57385 2950
rect 57565 2950 57570 2955
rect 57600 2950 57605 2980
rect 57565 2945 57605 2950
rect 56140 2890 56180 2895
rect 56140 2860 56145 2890
rect 56175 2885 56180 2890
rect 56250 2890 56290 2895
rect 56250 2885 56255 2890
rect 56175 2865 56255 2885
rect 56175 2860 56180 2865
rect 56140 2855 56180 2860
rect 56250 2860 56255 2865
rect 56285 2885 56290 2890
rect 56360 2890 56400 2895
rect 56360 2885 56365 2890
rect 56285 2865 56365 2885
rect 56285 2860 56290 2865
rect 56250 2855 56290 2860
rect 56360 2860 56365 2865
rect 56395 2885 56400 2890
rect 56470 2890 56510 2895
rect 56470 2885 56475 2890
rect 56395 2865 56475 2885
rect 56395 2860 56400 2865
rect 56360 2855 56400 2860
rect 56470 2860 56475 2865
rect 56505 2885 56510 2890
rect 56580 2890 56620 2895
rect 56580 2885 56585 2890
rect 56505 2865 56585 2885
rect 56505 2860 56510 2865
rect 56470 2855 56510 2860
rect 56580 2860 56585 2865
rect 56615 2860 56620 2890
rect 56580 2855 56620 2860
rect 57180 2890 57220 2895
rect 57180 2860 57185 2890
rect 57215 2885 57220 2890
rect 57290 2890 57330 2895
rect 57290 2885 57295 2890
rect 57215 2865 57295 2885
rect 57215 2860 57220 2865
rect 57180 2855 57220 2860
rect 57290 2860 57295 2865
rect 57325 2885 57330 2890
rect 57400 2890 57440 2895
rect 57400 2885 57405 2890
rect 57325 2865 57405 2885
rect 57325 2860 57330 2865
rect 57290 2855 57330 2860
rect 57400 2860 57405 2865
rect 57435 2885 57440 2890
rect 57510 2890 57550 2895
rect 57510 2885 57515 2890
rect 57435 2865 57515 2885
rect 57435 2860 57440 2865
rect 57400 2855 57440 2860
rect 57510 2860 57515 2865
rect 57545 2885 57550 2890
rect 57620 2890 57660 2895
rect 57620 2885 57625 2890
rect 57545 2865 57625 2885
rect 57545 2860 57550 2865
rect 57510 2855 57550 2860
rect 57620 2860 57625 2865
rect 57655 2860 57660 2890
rect 57620 2855 57660 2860
rect 56085 2845 56125 2850
rect 56085 2815 56090 2845
rect 56120 2840 56125 2845
rect 56195 2845 56235 2850
rect 56195 2840 56200 2845
rect 56120 2820 56200 2840
rect 56120 2815 56125 2820
rect 56085 2810 56125 2815
rect 56195 2815 56200 2820
rect 56230 2840 56235 2845
rect 56305 2845 56345 2850
rect 56305 2840 56310 2845
rect 56230 2820 56310 2840
rect 56230 2815 56235 2820
rect 56195 2810 56235 2815
rect 56305 2815 56310 2820
rect 56340 2840 56345 2845
rect 56415 2845 56455 2850
rect 56415 2840 56420 2845
rect 56340 2820 56420 2840
rect 56340 2815 56345 2820
rect 56305 2810 56345 2815
rect 56415 2815 56420 2820
rect 56450 2840 56455 2845
rect 56525 2845 56565 2850
rect 56525 2840 56530 2845
rect 56450 2820 56530 2840
rect 56450 2815 56455 2820
rect 56415 2810 56455 2815
rect 56525 2815 56530 2820
rect 56560 2840 56565 2845
rect 56635 2845 56675 2850
rect 56635 2840 56640 2845
rect 56560 2820 56640 2840
rect 56560 2815 56565 2820
rect 56525 2810 56565 2815
rect 56635 2815 56640 2820
rect 56670 2840 56675 2845
rect 56825 2845 56865 2850
rect 56825 2840 56830 2845
rect 56670 2820 56830 2840
rect 56670 2815 56675 2820
rect 56635 2810 56675 2815
rect 56825 2815 56830 2820
rect 56860 2815 56865 2845
rect 56825 2810 56865 2815
rect 57125 2845 57165 2850
rect 57125 2815 57130 2845
rect 57160 2840 57165 2845
rect 57345 2845 57385 2850
rect 57345 2840 57350 2845
rect 57160 2820 57350 2840
rect 57160 2815 57165 2820
rect 57125 2810 57165 2815
rect 57345 2815 57350 2820
rect 57380 2840 57385 2845
rect 57565 2845 57605 2850
rect 57565 2840 57570 2845
rect 57380 2820 57570 2840
rect 57380 2815 57385 2820
rect 57345 2810 57385 2815
rect 57565 2815 57570 2820
rect 57600 2815 57605 2845
rect 57565 2810 57605 2815
rect 56580 2800 56610 2805
rect 56095 2790 56125 2795
rect 55955 2765 56095 2785
rect 57190 2800 57220 2805
rect 56610 2775 57190 2795
rect 56580 2765 56610 2770
rect 57190 2765 57220 2770
rect 56095 2755 56125 2760
rect 55750 2745 55790 2750
rect 55750 2715 55755 2745
rect 55785 2740 55790 2745
rect 56030 2745 56070 2750
rect 56030 2740 56035 2745
rect 55785 2720 56035 2740
rect 55785 2715 55790 2720
rect 55750 2710 55790 2715
rect 56030 2715 56035 2720
rect 56065 2740 56070 2745
rect 56690 2745 56730 2750
rect 56690 2740 56695 2745
rect 56065 2720 56695 2740
rect 56065 2715 56070 2720
rect 56030 2710 56070 2715
rect 56690 2715 56695 2720
rect 56725 2715 56730 2745
rect 56690 2710 56730 2715
rect 57070 2745 57110 2750
rect 57070 2715 57075 2745
rect 57105 2740 57110 2745
rect 57730 2745 57770 2750
rect 57730 2740 57735 2745
rect 57105 2720 57735 2740
rect 57105 2715 57110 2720
rect 57070 2710 57110 2715
rect 57730 2715 57735 2720
rect 57765 2740 57770 2745
rect 58010 2745 58050 2750
rect 58010 2740 58015 2745
rect 57765 2720 58015 2740
rect 57765 2715 57770 2720
rect 57730 2710 57770 2715
rect 58010 2715 58015 2720
rect 58045 2715 58050 2745
rect 58010 2710 58050 2715
rect 56935 2690 56975 2695
rect 54875 2660 54915 2665
rect 54875 2630 54880 2660
rect 54910 2655 54915 2660
rect 54985 2660 55025 2665
rect 54985 2655 54990 2660
rect 54910 2635 54990 2655
rect 54910 2630 54915 2635
rect 54875 2625 54915 2630
rect 54985 2630 54990 2635
rect 55020 2655 55025 2660
rect 55095 2660 55135 2665
rect 55095 2655 55100 2660
rect 55020 2635 55100 2655
rect 55020 2630 55025 2635
rect 54985 2625 55025 2630
rect 55095 2630 55100 2635
rect 55130 2655 55135 2660
rect 55205 2660 55245 2665
rect 55205 2655 55210 2660
rect 55130 2635 55210 2655
rect 55130 2630 55135 2635
rect 55095 2625 55135 2630
rect 55205 2630 55210 2635
rect 55240 2655 55245 2660
rect 55315 2660 55355 2665
rect 55315 2655 55320 2660
rect 55240 2635 55320 2655
rect 55240 2630 55245 2635
rect 55205 2625 55245 2630
rect 55315 2630 55320 2635
rect 55350 2655 55355 2660
rect 55425 2660 55465 2665
rect 55425 2655 55430 2660
rect 55350 2635 55430 2655
rect 55350 2630 55355 2635
rect 55315 2625 55355 2630
rect 55425 2630 55430 2635
rect 55460 2630 55465 2660
rect 56935 2660 56940 2690
rect 56970 2685 56975 2690
rect 57235 2690 57275 2695
rect 57235 2685 57240 2690
rect 56970 2665 57240 2685
rect 56970 2660 56975 2665
rect 56935 2655 56975 2660
rect 57235 2660 57240 2665
rect 57270 2685 57275 2690
rect 57455 2690 57495 2695
rect 57455 2685 57460 2690
rect 57270 2665 57460 2685
rect 57270 2660 57275 2665
rect 57235 2655 57275 2660
rect 57455 2660 57460 2665
rect 57490 2685 57495 2690
rect 57675 2690 57715 2695
rect 57675 2685 57680 2690
rect 57490 2665 57680 2685
rect 57490 2660 57495 2665
rect 57455 2655 57495 2660
rect 57675 2660 57680 2665
rect 57710 2685 57715 2690
rect 57865 2690 57905 2695
rect 57865 2685 57870 2690
rect 57710 2665 57870 2685
rect 57710 2660 57715 2665
rect 57675 2655 57715 2660
rect 57865 2660 57870 2665
rect 57900 2660 57905 2690
rect 57865 2655 57905 2660
rect 58335 2660 58375 2665
rect 55425 2625 55465 2630
rect 56850 2635 56890 2640
rect 56850 2605 56855 2635
rect 56885 2630 56890 2635
rect 57345 2635 57385 2640
rect 57345 2630 57350 2635
rect 56885 2610 57350 2630
rect 56885 2605 56890 2610
rect 56850 2600 56890 2605
rect 57345 2605 57350 2610
rect 57380 2605 57385 2635
rect 58335 2630 58340 2660
rect 58370 2655 58375 2660
rect 58445 2660 58485 2665
rect 58445 2655 58450 2660
rect 58370 2635 58450 2655
rect 58370 2630 58375 2635
rect 58335 2625 58375 2630
rect 58445 2630 58450 2635
rect 58480 2655 58485 2660
rect 58555 2660 58595 2665
rect 58555 2655 58560 2660
rect 58480 2635 58560 2655
rect 58480 2630 58485 2635
rect 58445 2625 58485 2630
rect 58555 2630 58560 2635
rect 58590 2655 58595 2660
rect 58665 2660 58705 2665
rect 58665 2655 58670 2660
rect 58590 2635 58670 2655
rect 58590 2630 58595 2635
rect 58555 2625 58595 2630
rect 58665 2630 58670 2635
rect 58700 2655 58705 2660
rect 58775 2660 58815 2665
rect 58775 2655 58780 2660
rect 58700 2635 58780 2655
rect 58700 2630 58705 2635
rect 58665 2625 58705 2630
rect 58775 2630 58780 2635
rect 58810 2655 58815 2660
rect 58885 2660 58925 2665
rect 58885 2655 58890 2660
rect 58810 2635 58890 2655
rect 58810 2630 58815 2635
rect 58775 2625 58815 2630
rect 58885 2630 58890 2635
rect 58920 2630 58925 2660
rect 58885 2625 58925 2630
rect 57345 2600 57385 2605
rect 54565 2580 56675 2585
rect 54565 2550 54570 2580
rect 54600 2550 54610 2580
rect 54640 2550 54650 2580
rect 54680 2550 55155 2580
rect 55185 2550 55605 2580
rect 55635 2550 55645 2580
rect 55675 2550 55685 2580
rect 55715 2550 56090 2580
rect 56120 2550 56145 2580
rect 56175 2550 56200 2580
rect 56230 2550 56255 2580
rect 56285 2550 56310 2580
rect 56340 2550 56365 2580
rect 56395 2550 56420 2580
rect 56450 2550 56475 2580
rect 56505 2550 56530 2580
rect 56560 2550 56585 2580
rect 56615 2550 56640 2580
rect 56670 2550 56675 2580
rect 54565 2540 56675 2550
rect 54565 2510 54570 2540
rect 54600 2510 54610 2540
rect 54640 2510 54650 2540
rect 54680 2510 55155 2540
rect 55185 2510 55605 2540
rect 55635 2510 55645 2540
rect 55675 2510 55685 2540
rect 55715 2510 56090 2540
rect 56120 2510 56145 2540
rect 56175 2510 56200 2540
rect 56230 2510 56255 2540
rect 56285 2510 56310 2540
rect 56340 2510 56365 2540
rect 56395 2510 56420 2540
rect 56450 2510 56475 2540
rect 56505 2510 56530 2540
rect 56560 2510 56585 2540
rect 56615 2510 56640 2540
rect 56670 2510 56675 2540
rect 54565 2500 56675 2510
rect 54565 2470 54570 2500
rect 54600 2470 54610 2500
rect 54640 2470 54650 2500
rect 54680 2470 55155 2500
rect 55185 2470 55605 2500
rect 55635 2470 55645 2500
rect 55675 2470 55685 2500
rect 55715 2470 56090 2500
rect 56120 2470 56145 2500
rect 56175 2470 56200 2500
rect 56230 2470 56255 2500
rect 56285 2470 56310 2500
rect 56340 2470 56365 2500
rect 56395 2470 56420 2500
rect 56450 2470 56475 2500
rect 56505 2470 56530 2500
rect 56560 2470 56585 2500
rect 56615 2470 56640 2500
rect 56670 2470 56675 2500
rect 54565 2465 56675 2470
rect 57125 2580 59235 2585
rect 57125 2550 57130 2580
rect 57160 2550 57185 2580
rect 57215 2550 57240 2580
rect 57270 2550 57295 2580
rect 57325 2550 57350 2580
rect 57380 2550 57405 2580
rect 57435 2550 57460 2580
rect 57490 2550 57515 2580
rect 57545 2550 57570 2580
rect 57600 2550 57625 2580
rect 57655 2550 57680 2580
rect 57710 2550 58085 2580
rect 58115 2550 58125 2580
rect 58155 2550 58165 2580
rect 58195 2550 58615 2580
rect 58645 2550 59120 2580
rect 59150 2550 59160 2580
rect 59190 2550 59200 2580
rect 59230 2550 59235 2580
rect 57125 2540 59235 2550
rect 57125 2510 57130 2540
rect 57160 2510 57185 2540
rect 57215 2510 57240 2540
rect 57270 2510 57295 2540
rect 57325 2510 57350 2540
rect 57380 2510 57405 2540
rect 57435 2510 57460 2540
rect 57490 2510 57515 2540
rect 57545 2510 57570 2540
rect 57600 2510 57625 2540
rect 57655 2510 57680 2540
rect 57710 2510 58085 2540
rect 58115 2510 58125 2540
rect 58155 2510 58165 2540
rect 58195 2510 58615 2540
rect 58645 2510 59120 2540
rect 59150 2510 59160 2540
rect 59190 2510 59200 2540
rect 59230 2510 59235 2540
rect 57125 2500 59235 2510
rect 57125 2470 57130 2500
rect 57160 2470 57185 2500
rect 57215 2470 57240 2500
rect 57270 2470 57295 2500
rect 57325 2470 57350 2500
rect 57380 2470 57405 2500
rect 57435 2470 57460 2500
rect 57490 2470 57515 2500
rect 57545 2470 57570 2500
rect 57600 2470 57625 2500
rect 57655 2470 57680 2500
rect 57710 2470 58085 2500
rect 58115 2470 58125 2500
rect 58155 2470 58165 2500
rect 58195 2470 58615 2500
rect 58645 2470 59120 2500
rect 59150 2470 59160 2500
rect 59190 2470 59200 2500
rect 59230 2470 59235 2500
rect 57125 2465 59235 2470
rect 54185 2430 55465 2435
rect 54185 2400 54190 2430
rect 54220 2400 54230 2430
rect 54260 2400 54275 2430
rect 54305 2400 54315 2430
rect 54345 2400 54360 2430
rect 54390 2400 54400 2430
rect 54430 2400 54880 2430
rect 54910 2400 54935 2430
rect 54965 2400 54990 2430
rect 55020 2400 55045 2430
rect 55075 2400 55100 2430
rect 55130 2400 55155 2430
rect 55185 2400 55210 2430
rect 55240 2400 55265 2430
rect 55295 2400 55320 2430
rect 55350 2400 55375 2430
rect 55405 2400 55430 2430
rect 55460 2400 55465 2430
rect 54185 2390 55465 2400
rect 54185 2360 54190 2390
rect 54220 2360 54230 2390
rect 54260 2360 54275 2390
rect 54305 2360 54315 2390
rect 54345 2360 54360 2390
rect 54390 2360 54400 2390
rect 54430 2360 54880 2390
rect 54910 2360 54935 2390
rect 54965 2360 54990 2390
rect 55020 2360 55045 2390
rect 55075 2360 55100 2390
rect 55130 2360 55155 2390
rect 55185 2360 55210 2390
rect 55240 2360 55265 2390
rect 55295 2360 55320 2390
rect 55350 2360 55375 2390
rect 55405 2360 55430 2390
rect 55460 2360 55465 2390
rect 54185 2350 55465 2360
rect 54185 2320 54190 2350
rect 54220 2320 54230 2350
rect 54260 2320 54275 2350
rect 54305 2320 54315 2350
rect 54345 2320 54360 2350
rect 54390 2320 54400 2350
rect 54430 2320 54880 2350
rect 54910 2320 54935 2350
rect 54965 2320 54990 2350
rect 55020 2320 55045 2350
rect 55075 2320 55100 2350
rect 55130 2320 55155 2350
rect 55185 2320 55210 2350
rect 55240 2320 55265 2350
rect 55295 2320 55320 2350
rect 55350 2320 55375 2350
rect 55405 2320 55430 2350
rect 55460 2320 55465 2350
rect 58335 2430 59615 2435
rect 58335 2400 58340 2430
rect 58370 2400 58395 2430
rect 58425 2400 58450 2430
rect 58480 2400 58505 2430
rect 58535 2400 58560 2430
rect 58590 2400 58615 2430
rect 58645 2400 58670 2430
rect 58700 2400 58725 2430
rect 58755 2400 58780 2430
rect 58810 2400 58835 2430
rect 58865 2400 58890 2430
rect 58920 2400 59370 2430
rect 59400 2400 59410 2430
rect 59440 2400 59455 2430
rect 59485 2400 59495 2430
rect 59525 2400 59540 2430
rect 59570 2400 59580 2430
rect 59610 2400 59615 2430
rect 58335 2390 59615 2400
rect 58335 2360 58340 2390
rect 58370 2360 58395 2390
rect 58425 2360 58450 2390
rect 58480 2360 58505 2390
rect 58535 2360 58560 2390
rect 58590 2360 58615 2390
rect 58645 2360 58670 2390
rect 58700 2360 58725 2390
rect 58755 2360 58780 2390
rect 58810 2360 58835 2390
rect 58865 2360 58890 2390
rect 58920 2360 59370 2390
rect 59400 2360 59410 2390
rect 59440 2360 59455 2390
rect 59485 2360 59495 2390
rect 59525 2360 59540 2390
rect 59570 2360 59580 2390
rect 59610 2360 59615 2390
rect 58335 2350 59615 2360
rect 58335 2320 58340 2350
rect 58370 2320 58395 2350
rect 58425 2320 58450 2350
rect 58480 2320 58505 2350
rect 58535 2320 58560 2350
rect 58590 2320 58615 2350
rect 58645 2320 58670 2350
rect 58700 2320 58725 2350
rect 58755 2320 58780 2350
rect 58810 2320 58835 2350
rect 58865 2320 58890 2350
rect 58920 2320 59370 2350
rect 59400 2320 59410 2350
rect 59440 2320 59455 2350
rect 59485 2320 59495 2350
rect 59525 2320 59540 2350
rect 59570 2320 59580 2350
rect 59610 2320 59615 2350
rect 54185 2315 55465 2320
rect 56770 2315 56810 2320
rect 54820 2290 54860 2295
rect 54820 2260 54825 2290
rect 54855 2285 54860 2290
rect 55480 2290 55520 2295
rect 55480 2285 55485 2290
rect 54855 2265 55485 2285
rect 54855 2260 54860 2265
rect 54820 2255 54860 2260
rect 55480 2260 55485 2265
rect 55515 2285 55520 2290
rect 55750 2290 55790 2295
rect 55750 2285 55755 2290
rect 55515 2265 55755 2285
rect 55515 2260 55520 2265
rect 55480 2255 55520 2260
rect 55750 2260 55755 2265
rect 55785 2260 55790 2290
rect 56770 2285 56775 2315
rect 56805 2310 56810 2315
rect 56880 2315 56920 2320
rect 56880 2310 56885 2315
rect 56805 2290 56885 2310
rect 56805 2285 56810 2290
rect 56770 2280 56810 2285
rect 56880 2285 56885 2290
rect 56915 2310 56920 2315
rect 56990 2315 57030 2320
rect 56990 2310 56995 2315
rect 56915 2290 56995 2310
rect 56915 2285 56920 2290
rect 56880 2280 56920 2285
rect 56990 2285 56995 2290
rect 57025 2310 57030 2315
rect 57930 2315 57970 2320
rect 58335 2315 59615 2320
rect 57930 2310 57935 2315
rect 57025 2290 57935 2310
rect 57025 2285 57030 2290
rect 56990 2280 57030 2285
rect 57930 2285 57935 2290
rect 57965 2285 57970 2315
rect 57930 2280 57970 2285
rect 58010 2290 58050 2295
rect 55750 2255 55790 2260
rect 55895 2270 55935 2275
rect 54115 2245 54155 2250
rect 54115 2215 54120 2245
rect 54150 2240 54155 2245
rect 54875 2245 54915 2250
rect 54875 2240 54880 2245
rect 54150 2220 54880 2240
rect 54150 2215 54155 2220
rect 54115 2210 54155 2215
rect 54875 2215 54880 2220
rect 54910 2240 54915 2245
rect 54985 2245 55025 2250
rect 54985 2240 54990 2245
rect 54910 2220 54990 2240
rect 54910 2215 54915 2220
rect 54875 2210 54915 2215
rect 54985 2215 54990 2220
rect 55020 2240 55025 2245
rect 55095 2245 55135 2250
rect 55095 2240 55100 2245
rect 55020 2220 55100 2240
rect 55020 2215 55025 2220
rect 54985 2210 55025 2215
rect 55095 2215 55100 2220
rect 55130 2240 55135 2245
rect 55205 2245 55245 2250
rect 55205 2240 55210 2245
rect 55130 2220 55210 2240
rect 55130 2215 55135 2220
rect 55095 2210 55135 2215
rect 55205 2215 55210 2220
rect 55240 2240 55245 2245
rect 55315 2245 55355 2250
rect 55315 2240 55320 2245
rect 55240 2220 55320 2240
rect 55240 2215 55245 2220
rect 55205 2210 55245 2215
rect 55315 2215 55320 2220
rect 55350 2240 55355 2245
rect 55425 2245 55465 2250
rect 55425 2240 55430 2245
rect 55350 2220 55430 2240
rect 55350 2215 55355 2220
rect 55315 2210 55355 2215
rect 55425 2215 55430 2220
rect 55460 2215 55465 2245
rect 55895 2240 55900 2270
rect 55930 2265 55935 2270
rect 55995 2270 56025 2275
rect 55930 2245 55995 2265
rect 55930 2240 55935 2245
rect 55895 2235 55935 2240
rect 56690 2270 56720 2275
rect 55995 2235 56025 2240
rect 56140 2260 56180 2265
rect 56140 2230 56145 2260
rect 56175 2255 56180 2260
rect 56250 2260 56290 2265
rect 56250 2255 56255 2260
rect 56175 2235 56255 2255
rect 56175 2230 56180 2235
rect 56140 2225 56180 2230
rect 56250 2230 56255 2235
rect 56285 2255 56290 2260
rect 56360 2260 56400 2265
rect 56360 2255 56365 2260
rect 56285 2235 56365 2255
rect 56285 2230 56290 2235
rect 56250 2225 56290 2230
rect 56360 2230 56365 2235
rect 56395 2255 56400 2260
rect 56470 2260 56510 2265
rect 56470 2255 56475 2260
rect 56395 2235 56475 2255
rect 56395 2230 56400 2235
rect 56360 2225 56400 2230
rect 56470 2230 56475 2235
rect 56505 2255 56510 2260
rect 56580 2260 56620 2265
rect 56580 2255 56585 2260
rect 56505 2235 56585 2255
rect 56505 2230 56510 2235
rect 56470 2225 56510 2230
rect 56580 2230 56585 2235
rect 56615 2230 56620 2260
rect 56635 2235 56675 2255
rect 57080 2270 57110 2275
rect 56720 2245 57080 2265
rect 56690 2235 56720 2240
rect 57080 2235 57110 2240
rect 57180 2260 57220 2265
rect 56580 2225 56620 2230
rect 57180 2230 57185 2260
rect 57215 2255 57220 2260
rect 57290 2260 57330 2265
rect 57290 2255 57295 2260
rect 57215 2235 57295 2255
rect 57215 2230 57220 2235
rect 57180 2225 57220 2230
rect 57290 2230 57295 2235
rect 57325 2255 57330 2260
rect 57400 2260 57440 2265
rect 57400 2255 57405 2260
rect 57325 2235 57405 2255
rect 57325 2230 57330 2235
rect 57290 2225 57330 2230
rect 57400 2230 57405 2235
rect 57435 2255 57440 2260
rect 57510 2260 57550 2265
rect 57510 2255 57515 2260
rect 57435 2235 57515 2255
rect 57435 2230 57440 2235
rect 57400 2225 57440 2230
rect 57510 2230 57515 2235
rect 57545 2255 57550 2260
rect 57620 2260 57660 2265
rect 57620 2255 57625 2260
rect 57545 2235 57625 2255
rect 57545 2230 57550 2235
rect 57510 2225 57550 2230
rect 57620 2230 57625 2235
rect 57655 2230 57660 2260
rect 58010 2260 58015 2290
rect 58045 2285 58050 2290
rect 58280 2290 58320 2295
rect 58280 2285 58285 2290
rect 58045 2265 58285 2285
rect 58045 2260 58050 2265
rect 58010 2255 58050 2260
rect 58280 2260 58285 2265
rect 58315 2285 58320 2290
rect 58940 2290 58980 2295
rect 58940 2285 58945 2290
rect 58315 2265 58945 2285
rect 58315 2260 58320 2265
rect 58280 2255 58320 2260
rect 58940 2260 58945 2265
rect 58975 2260 58980 2290
rect 58940 2255 58980 2260
rect 57620 2225 57660 2230
rect 58335 2245 58375 2250
rect 55425 2210 55465 2215
rect 56085 2215 56125 2220
rect 54930 2200 54970 2205
rect 54930 2170 54935 2200
rect 54965 2195 54970 2200
rect 55040 2200 55080 2205
rect 55040 2195 55045 2200
rect 54965 2175 55045 2195
rect 54965 2170 54970 2175
rect 54930 2165 54970 2170
rect 55040 2170 55045 2175
rect 55075 2195 55080 2200
rect 55150 2200 55190 2205
rect 55150 2195 55155 2200
rect 55075 2175 55155 2195
rect 55075 2170 55080 2175
rect 55040 2165 55080 2170
rect 55150 2170 55155 2175
rect 55185 2195 55190 2200
rect 55260 2200 55300 2205
rect 55260 2195 55265 2200
rect 55185 2175 55265 2195
rect 55185 2170 55190 2175
rect 55150 2165 55190 2170
rect 55260 2170 55265 2175
rect 55295 2195 55300 2200
rect 55370 2200 55410 2205
rect 55370 2195 55375 2200
rect 55295 2175 55375 2195
rect 55295 2170 55300 2175
rect 55260 2165 55300 2170
rect 55370 2170 55375 2175
rect 55405 2170 55410 2200
rect 56085 2185 56090 2215
rect 56120 2210 56125 2215
rect 56195 2215 56235 2220
rect 56195 2210 56200 2215
rect 56120 2190 56200 2210
rect 56120 2185 56125 2190
rect 56085 2180 56125 2185
rect 56195 2185 56200 2190
rect 56230 2210 56235 2215
rect 56305 2215 56345 2220
rect 56305 2210 56310 2215
rect 56230 2190 56310 2210
rect 56230 2185 56235 2190
rect 56195 2180 56235 2185
rect 56305 2185 56310 2190
rect 56340 2210 56345 2215
rect 56415 2215 56455 2220
rect 56415 2210 56420 2215
rect 56340 2190 56420 2210
rect 56340 2185 56345 2190
rect 56305 2180 56345 2185
rect 56415 2185 56420 2190
rect 56450 2210 56455 2215
rect 56525 2215 56565 2220
rect 56525 2210 56530 2215
rect 56450 2190 56530 2210
rect 56450 2185 56455 2190
rect 56415 2180 56455 2185
rect 56525 2185 56530 2190
rect 56560 2210 56565 2215
rect 56635 2215 56675 2220
rect 56635 2210 56640 2215
rect 56560 2190 56640 2210
rect 56560 2185 56565 2190
rect 56525 2180 56565 2185
rect 56635 2185 56640 2190
rect 56670 2185 56675 2215
rect 56635 2180 56675 2185
rect 57125 2215 57165 2220
rect 57125 2185 57130 2215
rect 57160 2210 57165 2215
rect 57235 2215 57275 2220
rect 57235 2210 57240 2215
rect 57160 2190 57240 2210
rect 57160 2185 57165 2190
rect 57125 2180 57165 2185
rect 57235 2185 57240 2190
rect 57270 2210 57275 2215
rect 57345 2215 57385 2220
rect 57345 2210 57350 2215
rect 57270 2190 57350 2210
rect 57270 2185 57275 2190
rect 57235 2180 57275 2185
rect 57345 2185 57350 2190
rect 57380 2210 57385 2215
rect 57455 2215 57495 2220
rect 57455 2210 57460 2215
rect 57380 2190 57460 2210
rect 57380 2185 57385 2190
rect 57345 2180 57385 2185
rect 57455 2185 57460 2190
rect 57490 2210 57495 2215
rect 57565 2215 57605 2220
rect 57565 2210 57570 2215
rect 57490 2190 57570 2210
rect 57490 2185 57495 2190
rect 57455 2180 57495 2185
rect 57565 2185 57570 2190
rect 57600 2210 57605 2215
rect 57675 2215 57715 2220
rect 57675 2210 57680 2215
rect 57600 2190 57680 2210
rect 57600 2185 57605 2190
rect 57565 2180 57605 2185
rect 57675 2185 57680 2190
rect 57710 2185 57715 2215
rect 58335 2215 58340 2245
rect 58370 2240 58375 2245
rect 58445 2245 58485 2250
rect 58445 2240 58450 2245
rect 58370 2220 58450 2240
rect 58370 2215 58375 2220
rect 58335 2210 58375 2215
rect 58445 2215 58450 2220
rect 58480 2240 58485 2245
rect 58555 2245 58595 2250
rect 58555 2240 58560 2245
rect 58480 2220 58560 2240
rect 58480 2215 58485 2220
rect 58445 2210 58485 2215
rect 58555 2215 58560 2220
rect 58590 2240 58595 2245
rect 58665 2245 58705 2250
rect 58665 2240 58670 2245
rect 58590 2220 58670 2240
rect 58590 2215 58595 2220
rect 58555 2210 58595 2215
rect 58665 2215 58670 2220
rect 58700 2240 58705 2245
rect 58775 2245 58815 2250
rect 58775 2240 58780 2245
rect 58700 2220 58780 2240
rect 58700 2215 58705 2220
rect 58665 2210 58705 2215
rect 58775 2215 58780 2220
rect 58810 2240 58815 2245
rect 58885 2245 58925 2250
rect 58885 2240 58890 2245
rect 58810 2220 58890 2240
rect 58810 2215 58815 2220
rect 58775 2210 58815 2215
rect 58885 2215 58890 2220
rect 58920 2240 58925 2245
rect 59645 2245 59685 2250
rect 59645 2240 59650 2245
rect 58920 2220 59650 2240
rect 58920 2215 58925 2220
rect 58885 2210 58925 2215
rect 59645 2215 59650 2220
rect 59680 2215 59685 2245
rect 59645 2210 59685 2215
rect 57675 2180 57715 2185
rect 58390 2200 58430 2205
rect 55370 2165 55410 2170
rect 58390 2170 58395 2200
rect 58425 2195 58430 2200
rect 58500 2200 58540 2205
rect 58500 2195 58505 2200
rect 58425 2175 58505 2195
rect 58425 2170 58430 2175
rect 58390 2165 58430 2170
rect 58500 2170 58505 2175
rect 58535 2195 58540 2200
rect 58610 2200 58650 2205
rect 58610 2195 58615 2200
rect 58535 2175 58615 2195
rect 58535 2170 58540 2175
rect 58500 2165 58540 2170
rect 58610 2170 58615 2175
rect 58645 2195 58650 2200
rect 58720 2200 58760 2205
rect 58720 2195 58725 2200
rect 58645 2175 58725 2195
rect 58645 2170 58650 2175
rect 58610 2165 58650 2170
rect 58720 2170 58725 2175
rect 58755 2195 58760 2200
rect 58830 2200 58870 2205
rect 58830 2195 58835 2200
rect 58755 2175 58835 2195
rect 58755 2170 58760 2175
rect 58720 2165 58760 2170
rect 58830 2170 58835 2175
rect 58865 2170 58870 2200
rect 58830 2165 58870 2170
rect 56140 2025 56180 2030
rect 56140 1995 56145 2025
rect 56175 2020 56180 2025
rect 56250 2025 56290 2030
rect 56250 2020 56255 2025
rect 56175 2000 56255 2020
rect 56175 1995 56180 2000
rect 56140 1990 56180 1995
rect 56250 1995 56255 2000
rect 56285 2020 56290 2025
rect 56360 2025 56400 2030
rect 56360 2020 56365 2025
rect 56285 2000 56365 2020
rect 56285 1995 56290 2000
rect 56250 1990 56290 1995
rect 56360 1995 56365 2000
rect 56395 2020 56400 2025
rect 56470 2025 56510 2030
rect 56470 2020 56475 2025
rect 56395 2000 56475 2020
rect 56395 1995 56400 2000
rect 56360 1990 56400 1995
rect 56470 1995 56475 2000
rect 56505 2020 56510 2025
rect 56580 2025 56620 2030
rect 56580 2020 56585 2025
rect 56505 2000 56585 2020
rect 56505 1995 56510 2000
rect 56470 1990 56510 1995
rect 56580 1995 56585 2000
rect 56615 1995 56620 2025
rect 56580 1990 56620 1995
rect 57180 2025 57220 2030
rect 57180 1995 57185 2025
rect 57215 2020 57220 2025
rect 57290 2025 57330 2030
rect 57290 2020 57295 2025
rect 57215 2000 57295 2020
rect 57215 1995 57220 2000
rect 57180 1990 57220 1995
rect 57290 1995 57295 2000
rect 57325 2020 57330 2025
rect 57400 2025 57440 2030
rect 57400 2020 57405 2025
rect 57325 2000 57405 2020
rect 57325 1995 57330 2000
rect 57290 1990 57330 1995
rect 57400 1995 57405 2000
rect 57435 2020 57440 2025
rect 57510 2025 57550 2030
rect 57510 2020 57515 2025
rect 57435 2000 57515 2020
rect 57435 1995 57440 2000
rect 57400 1990 57440 1995
rect 57510 1995 57515 2000
rect 57545 2020 57550 2025
rect 57620 2025 57660 2030
rect 57620 2020 57625 2025
rect 57545 2000 57625 2020
rect 57545 1995 57550 2000
rect 57510 1990 57550 1995
rect 57620 1995 57625 2000
rect 57655 1995 57660 2025
rect 57620 1990 57660 1995
rect 56085 1980 56125 1985
rect 56085 1950 56090 1980
rect 56120 1975 56125 1980
rect 56195 1980 56235 1985
rect 56195 1975 56200 1980
rect 56120 1955 56200 1975
rect 56120 1950 56125 1955
rect 54680 1945 54720 1950
rect 54680 1915 54685 1945
rect 54715 1940 54720 1945
rect 54930 1945 54970 1950
rect 54930 1940 54935 1945
rect 54715 1920 54935 1940
rect 54715 1915 54720 1920
rect 54680 1910 54720 1915
rect 54930 1915 54935 1920
rect 54965 1940 54970 1945
rect 55040 1945 55080 1950
rect 55040 1940 55045 1945
rect 54965 1920 55045 1940
rect 54965 1915 54970 1920
rect 54930 1910 54970 1915
rect 55040 1915 55045 1920
rect 55075 1940 55080 1945
rect 55150 1945 55190 1950
rect 55150 1940 55155 1945
rect 55075 1920 55155 1940
rect 55075 1915 55080 1920
rect 55040 1910 55080 1915
rect 55150 1915 55155 1920
rect 55185 1940 55190 1945
rect 55260 1945 55300 1950
rect 55260 1940 55265 1945
rect 55185 1920 55265 1940
rect 55185 1915 55190 1920
rect 55150 1910 55190 1915
rect 55260 1915 55265 1920
rect 55295 1940 55300 1945
rect 55370 1945 55410 1950
rect 56085 1945 56125 1950
rect 56195 1950 56200 1955
rect 56230 1975 56235 1980
rect 56305 1980 56345 1985
rect 56305 1975 56310 1980
rect 56230 1955 56310 1975
rect 56230 1950 56235 1955
rect 56195 1945 56235 1950
rect 56305 1950 56310 1955
rect 56340 1975 56345 1980
rect 56415 1980 56455 1985
rect 56415 1975 56420 1980
rect 56340 1955 56420 1975
rect 56340 1950 56345 1955
rect 56305 1945 56345 1950
rect 56415 1950 56420 1955
rect 56450 1975 56455 1980
rect 56525 1980 56565 1985
rect 56525 1975 56530 1980
rect 56450 1955 56530 1975
rect 56450 1950 56455 1955
rect 56415 1945 56455 1950
rect 56525 1950 56530 1955
rect 56560 1975 56565 1980
rect 56635 1980 56675 1985
rect 56635 1975 56640 1980
rect 56560 1955 56640 1975
rect 56560 1950 56565 1955
rect 56525 1945 56565 1950
rect 56635 1950 56640 1955
rect 56670 1950 56675 1980
rect 56635 1945 56675 1950
rect 57125 1980 57165 1985
rect 57125 1950 57130 1980
rect 57160 1975 57165 1980
rect 57235 1980 57275 1985
rect 57235 1975 57240 1980
rect 57160 1955 57240 1975
rect 57160 1950 57165 1955
rect 57125 1945 57165 1950
rect 57235 1950 57240 1955
rect 57270 1975 57275 1980
rect 57345 1980 57385 1985
rect 57345 1975 57350 1980
rect 57270 1955 57350 1975
rect 57270 1950 57275 1955
rect 57235 1945 57275 1950
rect 57345 1950 57350 1955
rect 57380 1975 57385 1980
rect 57455 1980 57495 1985
rect 57455 1975 57460 1980
rect 57380 1955 57460 1975
rect 57380 1950 57385 1955
rect 57345 1945 57385 1950
rect 57455 1950 57460 1955
rect 57490 1975 57495 1980
rect 57565 1980 57605 1985
rect 57565 1975 57570 1980
rect 57490 1955 57570 1975
rect 57490 1950 57495 1955
rect 57455 1945 57495 1950
rect 57565 1950 57570 1955
rect 57600 1975 57605 1980
rect 57675 1980 57715 1985
rect 57675 1975 57680 1980
rect 57600 1955 57680 1975
rect 57600 1950 57605 1955
rect 57565 1945 57605 1950
rect 57675 1950 57680 1955
rect 57710 1950 57715 1980
rect 57675 1945 57715 1950
rect 58390 1945 58430 1950
rect 55370 1940 55375 1945
rect 55295 1920 55375 1940
rect 55295 1915 55300 1920
rect 55260 1910 55300 1915
rect 55370 1915 55375 1920
rect 55405 1915 55410 1945
rect 55370 1910 55410 1915
rect 56030 1935 56070 1940
rect 56030 1905 56035 1935
rect 56065 1930 56070 1935
rect 56690 1935 56730 1940
rect 56690 1930 56695 1935
rect 56065 1910 56695 1930
rect 56065 1905 56070 1910
rect 56030 1900 56070 1905
rect 56690 1905 56695 1910
rect 56725 1930 56730 1935
rect 57070 1935 57110 1940
rect 57070 1930 57075 1935
rect 56725 1910 57075 1930
rect 56725 1905 56730 1910
rect 56690 1900 56730 1905
rect 57070 1905 57075 1910
rect 57105 1930 57110 1935
rect 57730 1935 57770 1940
rect 57730 1930 57735 1935
rect 57105 1910 57735 1930
rect 57105 1905 57110 1910
rect 57070 1900 57110 1905
rect 57730 1905 57735 1910
rect 57765 1930 57770 1935
rect 57930 1935 57970 1940
rect 57930 1930 57935 1935
rect 57765 1910 57935 1930
rect 57765 1905 57770 1910
rect 57730 1900 57770 1905
rect 57930 1905 57935 1910
rect 57965 1905 57970 1935
rect 58390 1915 58395 1945
rect 58425 1940 58430 1945
rect 58500 1945 58540 1950
rect 58500 1940 58505 1945
rect 58425 1920 58505 1940
rect 58425 1915 58430 1920
rect 58390 1910 58430 1915
rect 58500 1915 58505 1920
rect 58535 1940 58540 1945
rect 58610 1945 58650 1950
rect 58610 1940 58615 1945
rect 58535 1920 58615 1940
rect 58535 1915 58540 1920
rect 58500 1910 58540 1915
rect 58610 1915 58615 1920
rect 58645 1940 58650 1945
rect 58720 1945 58760 1950
rect 58720 1940 58725 1945
rect 58645 1920 58725 1940
rect 58645 1915 58650 1920
rect 58610 1910 58650 1915
rect 58720 1915 58725 1920
rect 58755 1940 58760 1945
rect 58830 1945 58870 1950
rect 58830 1940 58835 1945
rect 58755 1920 58835 1940
rect 58755 1915 58760 1920
rect 58720 1910 58760 1915
rect 58830 1915 58835 1920
rect 58865 1940 58870 1945
rect 59080 1945 59120 1950
rect 59080 1940 59085 1945
rect 58865 1920 59085 1940
rect 58865 1915 58870 1920
rect 58830 1910 58870 1915
rect 59080 1915 59085 1920
rect 59115 1915 59120 1945
rect 59080 1910 59120 1915
rect 57930 1900 57970 1905
rect 55315 1880 55720 1885
rect 55315 1850 55320 1880
rect 55350 1850 55605 1880
rect 55635 1850 55645 1880
rect 55675 1850 55685 1880
rect 55715 1850 55720 1880
rect 55315 1840 55720 1850
rect 55315 1810 55320 1840
rect 55350 1810 55605 1840
rect 55635 1810 55645 1840
rect 55675 1810 55685 1840
rect 55715 1810 55720 1840
rect 58080 1880 58485 1885
rect 58080 1850 58085 1880
rect 58115 1850 58125 1880
rect 58155 1850 58165 1880
rect 58195 1850 58450 1880
rect 58480 1850 58485 1880
rect 58080 1840 58485 1850
rect 58080 1810 58085 1840
rect 58115 1810 58125 1840
rect 58155 1810 58165 1840
rect 58195 1810 58450 1840
rect 58480 1810 58485 1840
rect 55315 1805 55720 1810
rect 56145 1805 56175 1810
rect 56085 1795 56125 1800
rect 56040 1785 56070 1790
rect 54725 1760 54765 1765
rect 54725 1730 54730 1760
rect 54760 1755 54765 1760
rect 54930 1760 54970 1765
rect 54930 1755 54935 1760
rect 54760 1735 54935 1755
rect 54760 1730 54765 1735
rect 54725 1725 54765 1730
rect 54930 1730 54935 1735
rect 54965 1755 54970 1760
rect 55040 1760 55080 1765
rect 55040 1755 55045 1760
rect 54965 1735 55045 1755
rect 54965 1730 54970 1735
rect 54930 1725 54970 1730
rect 55040 1730 55045 1735
rect 55075 1755 55080 1760
rect 55150 1760 55190 1765
rect 55150 1755 55155 1760
rect 55075 1735 55155 1755
rect 55075 1730 55080 1735
rect 55040 1725 55080 1730
rect 55150 1730 55155 1735
rect 55185 1755 55190 1760
rect 55260 1760 55300 1765
rect 55260 1755 55265 1760
rect 55185 1735 55265 1755
rect 55185 1730 55190 1735
rect 55150 1725 55190 1730
rect 55260 1730 55265 1735
rect 55295 1755 55300 1760
rect 55370 1760 55410 1765
rect 56030 1760 56040 1780
rect 55370 1755 55375 1760
rect 55295 1735 55375 1755
rect 55295 1730 55300 1735
rect 55260 1725 55300 1730
rect 55370 1730 55375 1735
rect 55405 1730 55410 1760
rect 56085 1765 56090 1795
rect 56120 1790 56125 1795
rect 56120 1775 56145 1790
rect 56255 1805 56285 1810
rect 56195 1795 56235 1800
rect 56195 1790 56200 1795
rect 56175 1775 56200 1790
rect 56120 1770 56200 1775
rect 56120 1765 56125 1770
rect 56085 1760 56125 1765
rect 56195 1765 56200 1770
rect 56230 1790 56235 1795
rect 56230 1775 56255 1790
rect 56365 1805 56395 1810
rect 56305 1795 56345 1800
rect 56305 1790 56310 1795
rect 56285 1775 56310 1790
rect 56230 1770 56310 1775
rect 56230 1765 56235 1770
rect 56195 1760 56235 1765
rect 56305 1765 56310 1770
rect 56340 1790 56345 1795
rect 56340 1775 56365 1790
rect 56475 1805 56505 1810
rect 56415 1795 56455 1800
rect 56415 1790 56420 1795
rect 56395 1775 56420 1790
rect 56340 1770 56420 1775
rect 56340 1765 56345 1770
rect 56305 1760 56345 1765
rect 56415 1765 56420 1770
rect 56450 1790 56455 1795
rect 56450 1775 56475 1790
rect 56585 1805 56615 1810
rect 56525 1795 56565 1800
rect 56525 1790 56530 1795
rect 56505 1775 56530 1790
rect 56450 1770 56530 1775
rect 56450 1765 56455 1770
rect 56415 1760 56455 1765
rect 56525 1765 56530 1770
rect 56560 1790 56565 1795
rect 56560 1775 56585 1790
rect 57185 1805 57215 1810
rect 56635 1795 56675 1800
rect 56635 1790 56640 1795
rect 56615 1775 56640 1790
rect 56560 1770 56640 1775
rect 56560 1765 56565 1770
rect 56525 1760 56565 1765
rect 56635 1765 56640 1770
rect 56670 1765 56675 1795
rect 57125 1795 57165 1800
rect 56635 1760 56675 1765
rect 56690 1785 56720 1790
rect 56850 1785 56880 1790
rect 56720 1760 56850 1780
rect 56040 1750 56070 1755
rect 56140 1750 56180 1755
rect 55370 1725 55410 1730
rect 56140 1720 56145 1750
rect 56175 1745 56180 1750
rect 56250 1750 56290 1755
rect 56250 1745 56255 1750
rect 56175 1725 56255 1745
rect 56175 1720 56180 1725
rect 54185 1710 54435 1720
rect 56140 1715 56180 1720
rect 56250 1720 56255 1725
rect 56285 1745 56290 1750
rect 56360 1750 56400 1755
rect 56360 1745 56365 1750
rect 56285 1725 56365 1745
rect 56285 1720 56290 1725
rect 56250 1715 56290 1720
rect 56360 1720 56365 1725
rect 56395 1745 56400 1750
rect 56470 1750 56510 1755
rect 56470 1745 56475 1750
rect 56395 1725 56475 1745
rect 56395 1720 56400 1725
rect 56360 1715 56400 1720
rect 56470 1720 56475 1725
rect 56505 1745 56510 1750
rect 56580 1750 56620 1755
rect 56690 1750 56720 1755
rect 56850 1750 56880 1755
rect 56903 1785 56933 1790
rect 57080 1785 57110 1790
rect 56933 1760 57080 1780
rect 56903 1750 56933 1755
rect 57125 1765 57130 1795
rect 57160 1790 57165 1795
rect 57160 1775 57185 1790
rect 57295 1805 57325 1810
rect 57235 1795 57275 1800
rect 57235 1790 57240 1795
rect 57215 1775 57240 1790
rect 57160 1770 57240 1775
rect 57160 1765 57165 1770
rect 57125 1760 57165 1765
rect 57235 1765 57240 1770
rect 57270 1790 57275 1795
rect 57270 1775 57295 1790
rect 57405 1805 57435 1810
rect 57345 1795 57385 1800
rect 57345 1790 57350 1795
rect 57325 1775 57350 1790
rect 57270 1770 57350 1775
rect 57270 1765 57275 1770
rect 57235 1760 57275 1765
rect 57345 1765 57350 1770
rect 57380 1790 57385 1795
rect 57380 1775 57405 1790
rect 57515 1805 57545 1810
rect 57455 1795 57495 1800
rect 57455 1790 57460 1795
rect 57435 1775 57460 1790
rect 57380 1770 57460 1775
rect 57380 1765 57385 1770
rect 57345 1760 57385 1765
rect 57455 1765 57460 1770
rect 57490 1790 57495 1795
rect 57490 1775 57515 1790
rect 57625 1805 57655 1810
rect 58080 1805 58485 1810
rect 57565 1795 57605 1800
rect 57565 1790 57570 1795
rect 57545 1775 57570 1790
rect 57490 1770 57570 1775
rect 57490 1765 57495 1770
rect 57455 1760 57495 1765
rect 57565 1765 57570 1770
rect 57600 1790 57605 1795
rect 57600 1775 57625 1790
rect 57675 1795 57715 1800
rect 57675 1790 57680 1795
rect 57655 1775 57680 1790
rect 57600 1770 57680 1775
rect 57600 1765 57605 1770
rect 57565 1760 57605 1765
rect 57675 1765 57680 1770
rect 57710 1765 57715 1795
rect 57675 1760 57715 1765
rect 57730 1785 57760 1790
rect 57760 1760 57770 1780
rect 58390 1760 58430 1765
rect 57080 1750 57110 1755
rect 57180 1750 57220 1755
rect 56580 1745 56585 1750
rect 56505 1725 56585 1745
rect 56505 1720 56510 1725
rect 56470 1715 56510 1720
rect 56580 1720 56585 1725
rect 56615 1720 56620 1750
rect 56580 1715 56620 1720
rect 57180 1720 57185 1750
rect 57215 1745 57220 1750
rect 57290 1750 57330 1755
rect 57290 1745 57295 1750
rect 57215 1725 57295 1745
rect 57215 1720 57220 1725
rect 57180 1715 57220 1720
rect 57290 1720 57295 1725
rect 57325 1745 57330 1750
rect 57400 1750 57440 1755
rect 57400 1745 57405 1750
rect 57325 1725 57405 1745
rect 57325 1720 57330 1725
rect 57290 1715 57330 1720
rect 57400 1720 57405 1725
rect 57435 1745 57440 1750
rect 57510 1750 57550 1755
rect 57510 1745 57515 1750
rect 57435 1725 57515 1745
rect 57435 1720 57440 1725
rect 57400 1715 57440 1720
rect 57510 1720 57515 1725
rect 57545 1745 57550 1750
rect 57620 1750 57660 1755
rect 57730 1750 57760 1755
rect 57620 1745 57625 1750
rect 57545 1725 57625 1745
rect 57545 1720 57550 1725
rect 57510 1715 57550 1720
rect 57620 1720 57625 1725
rect 57655 1720 57660 1750
rect 58390 1730 58395 1760
rect 58425 1755 58430 1760
rect 58500 1760 58540 1765
rect 58500 1755 58505 1760
rect 58425 1735 58505 1755
rect 58425 1730 58430 1735
rect 58390 1725 58430 1730
rect 58500 1730 58505 1735
rect 58535 1755 58540 1760
rect 58610 1760 58650 1765
rect 58610 1755 58615 1760
rect 58535 1735 58615 1755
rect 58535 1730 58540 1735
rect 58500 1725 58540 1730
rect 58610 1730 58615 1735
rect 58645 1755 58650 1760
rect 58720 1760 58760 1765
rect 58720 1755 58725 1760
rect 58645 1735 58725 1755
rect 58645 1730 58650 1735
rect 58610 1725 58650 1730
rect 58720 1730 58725 1735
rect 58755 1755 58760 1760
rect 58830 1760 58870 1765
rect 58830 1755 58835 1760
rect 58755 1735 58835 1755
rect 58755 1730 58760 1735
rect 58720 1725 58760 1730
rect 58830 1730 58835 1735
rect 58865 1755 58870 1760
rect 59035 1760 59075 1765
rect 59035 1755 59040 1760
rect 58865 1735 59040 1755
rect 58865 1730 58870 1735
rect 58830 1725 58870 1730
rect 59035 1730 59040 1735
rect 59070 1730 59075 1760
rect 59035 1725 59075 1730
rect 57620 1715 57660 1720
rect 54185 1680 54195 1710
rect 54225 1680 54245 1710
rect 54275 1680 54295 1710
rect 54325 1680 54345 1710
rect 54375 1680 54395 1710
rect 54425 1680 54435 1710
rect 54185 1660 54435 1680
rect 54185 1630 54195 1660
rect 54225 1630 54245 1660
rect 54275 1630 54295 1660
rect 54325 1630 54345 1660
rect 54375 1630 54395 1660
rect 54425 1630 54435 1660
rect 54185 1610 54435 1630
rect 54185 1580 54195 1610
rect 54225 1580 54245 1610
rect 54275 1580 54295 1610
rect 54325 1580 54345 1610
rect 54375 1580 54395 1610
rect 54425 1580 54435 1610
rect 54185 1570 54435 1580
rect 59365 1710 59615 1720
rect 59365 1680 59375 1710
rect 59405 1680 59425 1710
rect 59455 1680 59475 1710
rect 59505 1680 59525 1710
rect 59555 1680 59575 1710
rect 59605 1680 59615 1710
rect 59365 1660 59615 1680
rect 59365 1630 59375 1660
rect 59405 1630 59425 1660
rect 59455 1630 59475 1660
rect 59505 1630 59525 1660
rect 59555 1630 59575 1660
rect 59605 1630 59615 1660
rect 59365 1610 59615 1630
rect 59365 1580 59375 1610
rect 59405 1580 59425 1610
rect 59455 1580 59475 1610
rect 59505 1580 59525 1610
rect 59555 1580 59575 1610
rect 59605 1580 59615 1610
rect 59365 1570 59615 1580
rect 56085 1555 56125 1560
rect 56085 1525 56090 1555
rect 56120 1550 56125 1555
rect 56195 1555 56235 1560
rect 56195 1550 56200 1555
rect 56120 1530 56200 1550
rect 56120 1525 56125 1530
rect 56085 1520 56125 1525
rect 56195 1525 56200 1530
rect 56230 1550 56235 1555
rect 56305 1555 56345 1560
rect 56305 1550 56310 1555
rect 56230 1530 56310 1550
rect 56230 1525 56235 1530
rect 56195 1520 56235 1525
rect 56305 1525 56310 1530
rect 56340 1550 56345 1555
rect 56415 1555 56455 1560
rect 56415 1550 56420 1555
rect 56340 1530 56420 1550
rect 56340 1525 56345 1530
rect 56305 1520 56345 1525
rect 56415 1525 56420 1530
rect 56450 1550 56455 1555
rect 56525 1555 56565 1560
rect 56525 1550 56530 1555
rect 56450 1530 56530 1550
rect 56450 1525 56455 1530
rect 56415 1520 56455 1525
rect 56525 1525 56530 1530
rect 56560 1550 56565 1555
rect 56635 1555 56675 1560
rect 56635 1550 56640 1555
rect 56560 1530 56640 1550
rect 56560 1525 56565 1530
rect 56525 1520 56565 1525
rect 56635 1525 56640 1530
rect 56670 1525 56675 1555
rect 56635 1520 56675 1525
rect 57125 1555 57165 1560
rect 57125 1525 57130 1555
rect 57160 1550 57165 1555
rect 57235 1555 57275 1560
rect 57235 1550 57240 1555
rect 57160 1530 57240 1550
rect 57160 1525 57165 1530
rect 57125 1520 57165 1525
rect 57235 1525 57240 1530
rect 57270 1550 57275 1555
rect 57345 1555 57385 1560
rect 57345 1550 57350 1555
rect 57270 1530 57350 1550
rect 57270 1525 57275 1530
rect 57235 1520 57275 1525
rect 57345 1525 57350 1530
rect 57380 1550 57385 1555
rect 57455 1555 57495 1560
rect 57455 1550 57460 1555
rect 57380 1530 57460 1550
rect 57380 1525 57385 1530
rect 57345 1520 57385 1525
rect 57455 1525 57460 1530
rect 57490 1550 57495 1555
rect 57565 1555 57605 1560
rect 57565 1550 57570 1555
rect 57490 1530 57570 1550
rect 57490 1525 57495 1530
rect 57455 1520 57495 1525
rect 57565 1525 57570 1530
rect 57600 1550 57605 1555
rect 57675 1555 57715 1560
rect 57675 1550 57680 1555
rect 57600 1530 57680 1550
rect 57600 1525 57605 1530
rect 57565 1520 57605 1525
rect 57675 1525 57680 1530
rect 57710 1525 57715 1555
rect 57675 1520 57715 1525
rect 56140 1500 56180 1505
rect 56140 1470 56145 1500
rect 56175 1495 56180 1500
rect 56250 1500 56290 1505
rect 56250 1495 56255 1500
rect 56175 1475 56255 1495
rect 56175 1470 56180 1475
rect 56140 1465 56180 1470
rect 56250 1470 56255 1475
rect 56285 1495 56290 1500
rect 56360 1500 56400 1505
rect 56360 1495 56365 1500
rect 56285 1475 56365 1495
rect 56285 1470 56290 1475
rect 56250 1465 56290 1470
rect 56360 1470 56365 1475
rect 56395 1495 56400 1500
rect 56470 1500 56510 1505
rect 56470 1495 56475 1500
rect 56395 1475 56475 1495
rect 56395 1470 56400 1475
rect 56360 1465 56400 1470
rect 56470 1470 56475 1475
rect 56505 1495 56510 1500
rect 56580 1500 56620 1505
rect 56580 1495 56585 1500
rect 56505 1475 56585 1495
rect 56505 1470 56510 1475
rect 56470 1465 56510 1470
rect 56580 1470 56585 1475
rect 56615 1495 56620 1500
rect 57180 1500 57220 1505
rect 57180 1495 57185 1500
rect 56615 1475 57185 1495
rect 56615 1470 56620 1475
rect 56580 1465 56620 1470
rect 57180 1470 57185 1475
rect 57215 1495 57220 1500
rect 57290 1500 57330 1505
rect 57290 1495 57295 1500
rect 57215 1475 57295 1495
rect 57215 1470 57220 1475
rect 57180 1465 57220 1470
rect 57290 1470 57295 1475
rect 57325 1495 57330 1500
rect 57400 1500 57440 1505
rect 57400 1495 57405 1500
rect 57325 1475 57405 1495
rect 57325 1470 57330 1475
rect 57290 1465 57330 1470
rect 57400 1470 57405 1475
rect 57435 1495 57440 1500
rect 57510 1500 57550 1505
rect 57510 1495 57515 1500
rect 57435 1475 57515 1495
rect 57435 1470 57440 1475
rect 57400 1465 57440 1470
rect 57510 1470 57515 1475
rect 57545 1495 57550 1500
rect 57620 1500 57660 1505
rect 57620 1495 57625 1500
rect 57545 1475 57625 1495
rect 57545 1470 57550 1475
rect 57510 1465 57550 1470
rect 57620 1470 57625 1475
rect 57655 1470 57660 1500
rect 57620 1465 57660 1470
rect 54930 1420 54970 1425
rect 54460 1400 54495 1401
rect 54460 1395 54555 1400
rect 54495 1360 54520 1395
rect 54460 1355 54555 1360
rect 54580 1395 54615 1400
rect 54580 1355 54615 1360
rect 54640 1395 54675 1400
rect 54725 1390 54765 1395
rect 54725 1385 54730 1390
rect 54675 1365 54730 1385
rect 54640 1355 54675 1360
rect 54725 1360 54730 1365
rect 54760 1360 54765 1390
rect 54930 1390 54935 1420
rect 54965 1415 54970 1420
rect 55040 1420 55080 1425
rect 55040 1415 55045 1420
rect 54965 1395 55045 1415
rect 54965 1390 54970 1395
rect 54930 1385 54970 1390
rect 55040 1390 55045 1395
rect 55075 1415 55080 1420
rect 55150 1420 55190 1425
rect 55150 1415 55155 1420
rect 55075 1395 55155 1415
rect 55075 1390 55080 1395
rect 55040 1385 55080 1390
rect 55150 1390 55155 1395
rect 55185 1415 55190 1420
rect 55260 1420 55300 1425
rect 55260 1415 55265 1420
rect 55185 1395 55265 1415
rect 55185 1390 55190 1395
rect 55150 1385 55190 1390
rect 55260 1390 55265 1395
rect 55295 1415 55300 1420
rect 55370 1420 55410 1425
rect 55370 1415 55375 1420
rect 55295 1395 55375 1415
rect 55295 1390 55300 1395
rect 55260 1385 55300 1390
rect 55370 1390 55375 1395
rect 55405 1390 55410 1420
rect 55370 1385 55410 1390
rect 56825 1420 56865 1425
rect 56825 1390 56830 1420
rect 56860 1415 56865 1420
rect 56935 1420 56975 1425
rect 56935 1415 56940 1420
rect 56860 1395 56940 1415
rect 56860 1390 56865 1395
rect 56825 1385 56865 1390
rect 56935 1390 56940 1395
rect 56970 1390 56975 1420
rect 56935 1385 56975 1390
rect 58390 1420 58430 1425
rect 58390 1390 58395 1420
rect 58425 1415 58430 1420
rect 58500 1420 58540 1425
rect 58500 1415 58505 1420
rect 58425 1395 58505 1415
rect 58425 1390 58430 1395
rect 58390 1385 58430 1390
rect 58500 1390 58505 1395
rect 58535 1415 58540 1420
rect 58610 1420 58650 1425
rect 58610 1415 58615 1420
rect 58535 1395 58615 1415
rect 58535 1390 58540 1395
rect 58500 1385 58540 1390
rect 58610 1390 58615 1395
rect 58645 1415 58650 1420
rect 58720 1420 58760 1425
rect 58720 1415 58725 1420
rect 58645 1395 58725 1415
rect 58645 1390 58650 1395
rect 58610 1385 58650 1390
rect 58720 1390 58725 1395
rect 58755 1415 58760 1420
rect 58830 1420 58870 1425
rect 58830 1415 58835 1420
rect 58755 1395 58835 1415
rect 58755 1390 58760 1395
rect 58720 1385 58760 1390
rect 58830 1390 58835 1395
rect 58865 1390 58870 1420
rect 59305 1400 59340 1401
rect 59125 1395 59160 1400
rect 58830 1385 58870 1390
rect 59035 1390 59075 1395
rect 54725 1355 54765 1360
rect 54875 1375 54915 1380
rect 54875 1345 54880 1375
rect 54910 1370 54915 1375
rect 54985 1375 55025 1380
rect 54985 1370 54990 1375
rect 54910 1350 54990 1370
rect 54910 1345 54915 1350
rect 54875 1340 54915 1345
rect 54985 1345 54990 1350
rect 55020 1370 55025 1375
rect 55095 1375 55135 1380
rect 55095 1370 55100 1375
rect 55020 1350 55100 1370
rect 55020 1345 55025 1350
rect 54985 1340 55025 1345
rect 55095 1345 55100 1350
rect 55130 1370 55135 1375
rect 55205 1375 55245 1380
rect 55205 1370 55210 1375
rect 55130 1350 55210 1370
rect 55130 1345 55135 1350
rect 55095 1340 55135 1345
rect 55205 1345 55210 1350
rect 55240 1370 55245 1375
rect 55315 1375 55355 1380
rect 55315 1370 55320 1375
rect 55240 1350 55320 1370
rect 55240 1345 55245 1350
rect 55205 1340 55245 1345
rect 55315 1345 55320 1350
rect 55350 1370 55355 1375
rect 55425 1375 55465 1380
rect 55425 1370 55430 1375
rect 55350 1350 55430 1370
rect 55350 1345 55355 1350
rect 55315 1340 55355 1345
rect 55425 1345 55430 1350
rect 55460 1370 55465 1375
rect 55750 1375 55790 1380
rect 55750 1370 55755 1375
rect 55460 1350 55755 1370
rect 55460 1345 55465 1350
rect 55425 1340 55465 1345
rect 55750 1345 55755 1350
rect 55785 1345 55790 1375
rect 55750 1340 55790 1345
rect 58010 1375 58050 1380
rect 58010 1345 58015 1375
rect 58045 1370 58050 1375
rect 58335 1375 58375 1380
rect 58335 1370 58340 1375
rect 58045 1350 58340 1370
rect 58045 1345 58050 1350
rect 58010 1340 58050 1345
rect 58335 1345 58340 1350
rect 58370 1370 58375 1375
rect 58445 1375 58485 1380
rect 58445 1370 58450 1375
rect 58370 1350 58450 1370
rect 58370 1345 58375 1350
rect 58335 1340 58375 1345
rect 58445 1345 58450 1350
rect 58480 1370 58485 1375
rect 58555 1375 58595 1380
rect 58555 1370 58560 1375
rect 58480 1350 58560 1370
rect 58480 1345 58485 1350
rect 58445 1340 58485 1345
rect 58555 1345 58560 1350
rect 58590 1370 58595 1375
rect 58665 1375 58705 1380
rect 58665 1370 58670 1375
rect 58590 1350 58670 1370
rect 58590 1345 58595 1350
rect 58555 1340 58595 1345
rect 58665 1345 58670 1350
rect 58700 1370 58705 1375
rect 58775 1375 58815 1380
rect 58775 1370 58780 1375
rect 58700 1350 58780 1370
rect 58700 1345 58705 1350
rect 58665 1340 58705 1345
rect 58775 1345 58780 1350
rect 58810 1370 58815 1375
rect 58885 1375 58925 1380
rect 58885 1370 58890 1375
rect 58810 1350 58890 1370
rect 58810 1345 58815 1350
rect 58775 1340 58815 1345
rect 58885 1345 58890 1350
rect 58920 1345 58925 1375
rect 59035 1360 59040 1390
rect 59070 1385 59075 1390
rect 59070 1365 59125 1385
rect 59070 1360 59075 1365
rect 59035 1355 59075 1360
rect 59125 1355 59160 1360
rect 59185 1395 59220 1400
rect 59185 1355 59220 1360
rect 59245 1395 59340 1400
rect 59280 1360 59305 1395
rect 59245 1355 59340 1360
rect 58885 1340 58925 1345
rect 54580 1335 54620 1340
rect 54580 1305 54585 1335
rect 54615 1330 54620 1335
rect 54680 1335 54720 1340
rect 59080 1335 59120 1340
rect 54680 1330 54685 1335
rect 54615 1310 54685 1330
rect 54615 1305 54620 1310
rect 54580 1300 54620 1305
rect 54680 1305 54685 1310
rect 54715 1305 54720 1335
rect 54680 1300 54720 1305
rect 54820 1330 54860 1335
rect 54820 1300 54825 1330
rect 54855 1325 54860 1330
rect 55480 1330 55520 1335
rect 55480 1325 55485 1330
rect 54855 1305 55485 1325
rect 54855 1300 54860 1305
rect 54820 1295 54860 1300
rect 55480 1300 55485 1305
rect 55515 1325 55520 1330
rect 55830 1330 55870 1335
rect 55830 1325 55835 1330
rect 55515 1305 55835 1325
rect 55515 1300 55520 1305
rect 55480 1295 55520 1300
rect 55830 1300 55835 1305
rect 55865 1300 55870 1330
rect 55830 1295 55870 1300
rect 56030 1330 56070 1335
rect 56030 1300 56035 1330
rect 56065 1325 56070 1330
rect 56730 1330 56770 1335
rect 56730 1325 56735 1330
rect 56065 1305 56735 1325
rect 56065 1300 56070 1305
rect 56030 1295 56070 1300
rect 56730 1300 56735 1305
rect 56765 1325 56770 1330
rect 57030 1330 57070 1335
rect 57030 1325 57035 1330
rect 56765 1305 57035 1325
rect 56765 1300 56770 1305
rect 56730 1295 56770 1300
rect 57030 1300 57035 1305
rect 57065 1325 57070 1330
rect 57730 1330 57770 1335
rect 57730 1325 57735 1330
rect 57065 1305 57735 1325
rect 57065 1300 57070 1305
rect 57030 1295 57070 1300
rect 57730 1300 57735 1305
rect 57765 1325 57770 1330
rect 57930 1330 57970 1335
rect 57930 1325 57935 1330
rect 57765 1305 57935 1325
rect 57765 1300 57770 1305
rect 57730 1295 57770 1300
rect 57930 1300 57935 1305
rect 57965 1325 57970 1330
rect 58280 1330 58320 1335
rect 58280 1325 58285 1330
rect 57965 1305 58285 1325
rect 57965 1300 57970 1305
rect 57930 1295 57970 1300
rect 58280 1300 58285 1305
rect 58315 1325 58320 1330
rect 58940 1330 58980 1335
rect 58940 1325 58945 1330
rect 58315 1305 58945 1325
rect 58315 1300 58320 1305
rect 58280 1295 58320 1300
rect 58940 1300 58945 1305
rect 58975 1300 58980 1330
rect 59080 1305 59085 1335
rect 59115 1330 59120 1335
rect 59180 1335 59220 1340
rect 59180 1330 59185 1335
rect 59115 1310 59185 1330
rect 59115 1305 59120 1310
rect 59080 1300 59120 1305
rect 59180 1305 59185 1310
rect 59215 1305 59220 1335
rect 59180 1300 59220 1305
rect 58940 1295 58980 1300
rect 54460 1285 54500 1290
rect 54460 1255 54465 1285
rect 54495 1280 54500 1285
rect 55940 1285 55980 1290
rect 55940 1280 55945 1285
rect 54495 1260 55945 1280
rect 54495 1255 54500 1260
rect 54460 1250 54500 1255
rect 55940 1255 55945 1260
rect 55975 1255 55980 1285
rect 55940 1250 55980 1255
rect 57820 1285 57860 1290
rect 57820 1255 57825 1285
rect 57855 1280 57860 1285
rect 59300 1285 59340 1290
rect 59300 1280 59305 1285
rect 57855 1260 59305 1280
rect 57855 1255 57860 1260
rect 57820 1250 57860 1255
rect 59300 1255 59305 1260
rect 59335 1255 59340 1285
rect 59300 1250 59340 1255
rect 54595 1240 54635 1245
rect 54595 1210 54600 1240
rect 54630 1235 54635 1240
rect 55180 1240 55220 1245
rect 55180 1235 55185 1240
rect 54630 1215 55185 1235
rect 54630 1210 54635 1215
rect 54595 1205 54635 1210
rect 55180 1210 55185 1215
rect 55215 1235 55220 1240
rect 58580 1240 58620 1245
rect 58580 1235 58585 1240
rect 55215 1215 58585 1235
rect 55215 1210 55220 1215
rect 55180 1205 55220 1210
rect 58580 1210 58585 1215
rect 58615 1235 58620 1240
rect 59165 1240 59205 1245
rect 59165 1235 59170 1240
rect 58615 1215 59170 1235
rect 58615 1210 58620 1215
rect 58580 1205 58620 1210
rect 59165 1210 59170 1215
rect 59200 1210 59205 1240
rect 59165 1205 59205 1210
rect 54185 1185 55370 1190
rect 54185 1155 54190 1185
rect 54220 1155 54230 1185
rect 54260 1155 54275 1185
rect 54305 1155 54315 1185
rect 54345 1155 54360 1185
rect 54390 1155 54400 1185
rect 54430 1155 54665 1185
rect 54695 1155 54935 1185
rect 54965 1155 54975 1185
rect 55005 1155 55015 1185
rect 55045 1155 55055 1185
rect 55085 1155 55095 1185
rect 55125 1155 55135 1185
rect 55165 1155 55175 1185
rect 55205 1155 55215 1185
rect 55245 1155 55255 1185
rect 55285 1155 55295 1185
rect 55325 1155 55335 1185
rect 55365 1155 55370 1185
rect 54185 1145 55370 1155
rect 54185 1115 54190 1145
rect 54220 1115 54230 1145
rect 54260 1115 54275 1145
rect 54305 1115 54315 1145
rect 54345 1115 54360 1145
rect 54390 1115 54400 1145
rect 54430 1115 54665 1145
rect 54695 1115 54935 1145
rect 54965 1115 54975 1145
rect 55005 1115 55015 1145
rect 55045 1115 55055 1145
rect 55085 1115 55095 1145
rect 55125 1115 55135 1145
rect 55165 1115 55175 1145
rect 55205 1115 55215 1145
rect 55245 1115 55255 1145
rect 55285 1115 55295 1145
rect 55325 1115 55335 1145
rect 55365 1115 55370 1145
rect 58430 1185 59615 1190
rect 58430 1155 58435 1185
rect 58465 1155 58475 1185
rect 58505 1155 58515 1185
rect 58545 1155 58555 1185
rect 58585 1155 58595 1185
rect 58625 1155 58635 1185
rect 58665 1155 58675 1185
rect 58705 1155 58715 1185
rect 58745 1155 58755 1185
rect 58785 1155 58795 1185
rect 58825 1155 58835 1185
rect 58865 1155 59105 1185
rect 59135 1155 59370 1185
rect 59400 1155 59410 1185
rect 59440 1155 59455 1185
rect 59485 1155 59495 1185
rect 59525 1155 59540 1185
rect 59570 1155 59580 1185
rect 59610 1155 59615 1185
rect 58430 1145 59615 1155
rect 54185 1105 55370 1115
rect 54185 1075 54190 1105
rect 54220 1075 54230 1105
rect 54260 1075 54275 1105
rect 54305 1075 54315 1105
rect 54345 1075 54360 1105
rect 54390 1075 54400 1105
rect 54430 1075 54665 1105
rect 54695 1075 54935 1105
rect 54965 1075 54975 1105
rect 55005 1075 55015 1105
rect 55045 1075 55055 1105
rect 55085 1075 55095 1105
rect 55125 1075 55135 1105
rect 55165 1075 55175 1105
rect 55205 1075 55215 1105
rect 55245 1075 55255 1105
rect 55285 1075 55295 1105
rect 55325 1075 55335 1105
rect 55365 1075 55370 1105
rect 56330 1115 56370 1120
rect 56330 1085 56335 1115
rect 56365 1110 56370 1115
rect 56880 1115 56920 1120
rect 56880 1110 56885 1115
rect 56365 1090 56885 1110
rect 56365 1085 56370 1090
rect 56330 1080 56370 1085
rect 56880 1085 56885 1090
rect 56915 1085 56920 1115
rect 56880 1080 56920 1085
rect 57390 1115 57430 1120
rect 57390 1085 57395 1115
rect 57425 1110 57430 1115
rect 57865 1115 57905 1120
rect 57865 1110 57870 1115
rect 57425 1090 57870 1110
rect 57425 1085 57430 1090
rect 57390 1080 57430 1085
rect 57865 1085 57870 1090
rect 57900 1085 57905 1115
rect 57865 1080 57905 1085
rect 58430 1115 58435 1145
rect 58465 1115 58475 1145
rect 58505 1115 58515 1145
rect 58545 1115 58555 1145
rect 58585 1115 58595 1145
rect 58625 1115 58635 1145
rect 58665 1115 58675 1145
rect 58705 1115 58715 1145
rect 58745 1115 58755 1145
rect 58785 1115 58795 1145
rect 58825 1115 58835 1145
rect 58865 1115 59105 1145
rect 59135 1115 59370 1145
rect 59400 1115 59410 1145
rect 59440 1115 59455 1145
rect 59485 1115 59495 1145
rect 59525 1115 59540 1145
rect 59570 1115 59580 1145
rect 59610 1115 59615 1145
rect 58430 1105 59615 1115
rect 54185 1070 55370 1075
rect 58430 1075 58435 1105
rect 58465 1075 58475 1105
rect 58505 1075 58515 1105
rect 58545 1075 58555 1105
rect 58585 1075 58595 1105
rect 58625 1075 58635 1105
rect 58665 1075 58675 1105
rect 58705 1075 58715 1105
rect 58745 1075 58755 1105
rect 58785 1075 58795 1105
rect 58825 1075 58835 1105
rect 58865 1075 59105 1105
rect 59135 1075 59370 1105
rect 59400 1075 59410 1105
rect 59440 1075 59455 1105
rect 59485 1075 59495 1105
rect 59525 1075 59540 1105
rect 59570 1075 59580 1105
rect 59610 1075 59615 1105
rect 58430 1070 59615 1075
rect 56440 1060 56480 1065
rect 54600 1050 54635 1055
rect 54600 1010 54635 1015
rect 54660 1050 54695 1055
rect 56440 1030 56445 1060
rect 56475 1055 56480 1060
rect 56550 1060 56590 1065
rect 56550 1055 56555 1060
rect 56475 1035 56555 1055
rect 56475 1030 56480 1035
rect 56440 1025 56480 1030
rect 56550 1030 56555 1035
rect 56585 1055 56590 1060
rect 56660 1060 56700 1065
rect 56660 1055 56665 1060
rect 56585 1035 56665 1055
rect 56585 1030 56590 1035
rect 56550 1025 56590 1030
rect 56660 1030 56665 1035
rect 56695 1055 56700 1060
rect 56770 1060 56810 1065
rect 56770 1055 56775 1060
rect 56695 1035 56775 1055
rect 56695 1030 56700 1035
rect 56660 1025 56700 1030
rect 56770 1030 56775 1035
rect 56805 1055 56810 1060
rect 56880 1060 56920 1065
rect 56880 1055 56885 1060
rect 56805 1035 56885 1055
rect 56805 1030 56810 1035
rect 56770 1025 56810 1030
rect 56880 1030 56885 1035
rect 56915 1055 56920 1060
rect 56990 1060 57030 1065
rect 56990 1055 56995 1060
rect 56915 1035 56995 1055
rect 56915 1030 56920 1035
rect 56880 1025 56920 1030
rect 56990 1030 56995 1035
rect 57025 1055 57030 1060
rect 57100 1060 57140 1065
rect 57100 1055 57105 1060
rect 57025 1035 57105 1055
rect 57025 1030 57030 1035
rect 56990 1025 57030 1030
rect 57100 1030 57105 1035
rect 57135 1055 57140 1060
rect 57210 1060 57250 1065
rect 57210 1055 57215 1060
rect 57135 1035 57215 1055
rect 57135 1030 57140 1035
rect 57100 1025 57140 1030
rect 57210 1030 57215 1035
rect 57245 1055 57250 1060
rect 57320 1060 57360 1065
rect 57320 1055 57325 1060
rect 57245 1035 57325 1055
rect 57245 1030 57250 1035
rect 57210 1025 57250 1030
rect 57320 1030 57325 1035
rect 57355 1055 57360 1060
rect 57430 1060 57470 1065
rect 57430 1055 57435 1060
rect 57355 1035 57435 1055
rect 57355 1030 57360 1035
rect 57320 1025 57360 1030
rect 57430 1030 57435 1035
rect 57465 1030 57470 1060
rect 57430 1025 57470 1030
rect 59105 1050 59140 1055
rect 54660 1010 54695 1015
rect 59105 1010 59140 1015
rect 59165 1050 59200 1055
rect 59165 1010 59200 1015
rect 55830 740 55870 745
rect 55830 710 55835 740
rect 55865 735 55870 740
rect 56220 740 56260 745
rect 56220 735 56225 740
rect 55865 715 56225 735
rect 55865 710 55870 715
rect 55830 705 55870 710
rect 56220 710 56225 715
rect 56255 735 56260 740
rect 56275 740 56315 745
rect 56275 735 56280 740
rect 56255 715 56280 735
rect 56255 710 56260 715
rect 56220 705 56260 710
rect 56275 710 56280 715
rect 56310 735 56315 740
rect 56385 740 56425 745
rect 56385 735 56390 740
rect 56310 715 56390 735
rect 56310 710 56315 715
rect 56275 705 56315 710
rect 56385 710 56390 715
rect 56420 735 56425 740
rect 56495 740 56535 745
rect 56495 735 56500 740
rect 56420 715 56500 735
rect 56420 710 56425 715
rect 56385 705 56425 710
rect 56495 710 56500 715
rect 56530 735 56535 740
rect 56605 740 56645 745
rect 56605 735 56610 740
rect 56530 715 56610 735
rect 56530 710 56535 715
rect 56495 705 56535 710
rect 56605 710 56610 715
rect 56640 735 56645 740
rect 56715 740 56755 745
rect 56715 735 56720 740
rect 56640 715 56720 735
rect 56640 710 56645 715
rect 56605 705 56645 710
rect 56715 710 56720 715
rect 56750 735 56755 740
rect 56825 740 56865 745
rect 56825 735 56830 740
rect 56750 715 56830 735
rect 56750 710 56755 715
rect 56715 705 56755 710
rect 56825 710 56830 715
rect 56860 735 56865 740
rect 56935 740 56975 745
rect 56935 735 56940 740
rect 56860 715 56940 735
rect 56860 710 56865 715
rect 56825 705 56865 710
rect 56935 710 56940 715
rect 56970 735 56975 740
rect 57045 740 57085 745
rect 57045 735 57050 740
rect 56970 715 57050 735
rect 56970 710 56975 715
rect 56935 705 56975 710
rect 57045 710 57050 715
rect 57080 735 57085 740
rect 57155 740 57195 745
rect 57155 735 57160 740
rect 57080 715 57160 735
rect 57080 710 57085 715
rect 57045 705 57085 710
rect 57155 710 57160 715
rect 57190 735 57195 740
rect 57265 740 57305 745
rect 57265 735 57270 740
rect 57190 715 57270 735
rect 57190 710 57195 715
rect 57155 705 57195 710
rect 57265 710 57270 715
rect 57300 735 57305 740
rect 57375 740 57415 745
rect 57375 735 57380 740
rect 57300 715 57380 735
rect 57300 710 57305 715
rect 57265 705 57305 710
rect 57375 710 57380 715
rect 57410 735 57415 740
rect 57485 740 57525 745
rect 57485 735 57490 740
rect 57410 715 57490 735
rect 57410 710 57415 715
rect 57375 705 57415 710
rect 57485 710 57490 715
rect 57520 735 57525 740
rect 57930 740 57970 745
rect 57930 735 57935 740
rect 57520 715 57935 735
rect 57520 710 57525 715
rect 57485 705 57525 710
rect 57930 710 57935 715
rect 57965 710 57970 740
rect 57930 705 57970 710
rect 56440 695 56480 700
rect 56440 665 56445 695
rect 56475 690 56480 695
rect 56550 695 56590 700
rect 56550 690 56555 695
rect 56475 670 56555 690
rect 56475 665 56480 670
rect 56440 660 56480 665
rect 56550 665 56555 670
rect 56585 690 56590 695
rect 56660 695 56700 700
rect 56660 690 56665 695
rect 56585 670 56665 690
rect 56585 665 56590 670
rect 56550 660 56590 665
rect 56660 665 56665 670
rect 56695 690 56700 695
rect 56770 695 56810 700
rect 56770 690 56775 695
rect 56695 670 56775 690
rect 56695 665 56700 670
rect 56660 660 56700 665
rect 56770 665 56775 670
rect 56805 690 56810 695
rect 56880 695 56920 700
rect 56880 690 56885 695
rect 56805 670 56885 690
rect 56805 665 56810 670
rect 56770 660 56810 665
rect 56880 665 56885 670
rect 56915 690 56920 695
rect 56990 695 57030 700
rect 56990 690 56995 695
rect 56915 670 56995 690
rect 56915 665 56920 670
rect 56880 660 56920 665
rect 56990 665 56995 670
rect 57025 690 57030 695
rect 57100 695 57140 700
rect 57100 690 57105 695
rect 57025 670 57105 690
rect 57025 665 57030 670
rect 56990 660 57030 665
rect 57100 665 57105 670
rect 57135 690 57140 695
rect 57210 695 57250 700
rect 57210 690 57215 695
rect 57135 670 57215 690
rect 57135 665 57140 670
rect 57100 660 57140 665
rect 57210 665 57215 670
rect 57245 690 57250 695
rect 57320 695 57360 700
rect 57320 690 57325 695
rect 57245 670 57325 690
rect 57245 665 57250 670
rect 57210 660 57250 665
rect 57320 665 57325 670
rect 57355 690 57360 695
rect 57430 695 57470 700
rect 57430 690 57435 695
rect 57355 670 57435 690
rect 57355 665 57360 670
rect 57320 660 57360 665
rect 57430 665 57435 670
rect 57465 665 57470 695
rect 57430 660 57470 665
rect 56540 640 56580 645
rect 56540 610 56545 640
rect 56575 635 56580 640
rect 56650 640 56690 645
rect 56650 635 56655 640
rect 56575 615 56655 635
rect 56575 610 56580 615
rect 56540 605 56580 610
rect 56650 610 56655 615
rect 56685 635 56690 640
rect 56870 640 56910 645
rect 56870 635 56875 640
rect 56685 615 56875 635
rect 56685 610 56690 615
rect 56650 605 56690 610
rect 56870 610 56875 615
rect 56905 610 56910 640
rect 56870 605 56910 610
rect 55895 595 55935 600
rect 55895 565 55900 595
rect 55930 590 55935 595
rect 56485 595 56525 600
rect 56485 590 56490 595
rect 55930 570 56490 590
rect 55930 565 55935 570
rect 55895 560 55935 565
rect 56485 565 56490 570
rect 56520 590 56525 595
rect 56595 595 56635 600
rect 56595 590 56600 595
rect 56520 570 56600 590
rect 56520 565 56525 570
rect 56485 560 56525 565
rect 56595 565 56600 570
rect 56630 590 56635 595
rect 56705 595 56745 600
rect 56705 590 56710 595
rect 56630 570 56710 590
rect 56630 565 56635 570
rect 56595 560 56635 565
rect 56705 565 56710 570
rect 56740 590 56745 595
rect 57040 595 57080 600
rect 57040 590 57045 595
rect 56740 570 57045 590
rect 56740 565 56745 570
rect 56705 560 56745 565
rect 57040 565 57045 570
rect 57075 565 57080 595
rect 57040 560 57080 565
rect 56540 390 56580 395
rect 56540 360 56545 390
rect 56575 385 56580 390
rect 56650 390 56690 395
rect 56650 385 56655 390
rect 56575 365 56655 385
rect 56575 360 56580 365
rect 56540 355 56580 360
rect 56650 360 56655 365
rect 56685 385 56690 390
rect 56870 390 56910 395
rect 56870 385 56875 390
rect 56685 365 56875 385
rect 56685 360 56690 365
rect 56650 355 56690 360
rect 56870 360 56875 365
rect 56905 360 56910 390
rect 56870 355 56910 360
rect 54930 350 55370 355
rect 58430 350 58870 355
rect 54930 320 54935 350
rect 54965 320 55135 350
rect 55165 320 55335 350
rect 55365 320 55370 350
rect 54930 315 55370 320
rect 56485 345 56525 350
rect 56485 315 56490 345
rect 56520 340 56525 345
rect 56595 345 56635 350
rect 56595 340 56600 345
rect 56520 320 56600 340
rect 56520 315 56525 320
rect 56595 315 56600 320
rect 56630 340 56635 345
rect 56705 345 56745 350
rect 56705 340 56710 345
rect 56630 320 56710 340
rect 56630 315 56635 320
rect 56705 315 56710 320
rect 56740 315 56745 345
rect 58430 320 58435 350
rect 58465 320 58635 350
rect 58665 320 58835 350
rect 58865 320 58870 350
rect 58430 315 58870 320
rect 52640 45 61160 50
rect 52640 15 52645 45
rect 52675 15 52685 45
rect 52715 15 52725 45
rect 52755 15 52995 45
rect 53025 15 53035 45
rect 53065 15 53075 45
rect 53105 15 53345 45
rect 53375 15 53385 45
rect 53415 15 53425 45
rect 53455 15 53695 45
rect 53725 15 53735 45
rect 53765 15 53775 45
rect 53805 15 54045 45
rect 54075 15 54085 45
rect 54115 15 54125 45
rect 54155 15 54395 45
rect 54425 15 54435 45
rect 54465 15 54475 45
rect 54505 15 54745 45
rect 54775 15 54785 45
rect 54815 15 54825 45
rect 54855 15 55035 45
rect 55065 15 55095 45
rect 55125 15 55135 45
rect 55165 15 55175 45
rect 55205 15 55235 45
rect 55265 15 55445 45
rect 55475 15 55485 45
rect 55515 15 55525 45
rect 55555 15 55795 45
rect 55825 15 55835 45
rect 55865 15 55875 45
rect 55905 15 56145 45
rect 56175 15 56185 45
rect 56215 15 56225 45
rect 56255 15 56435 45
rect 56465 15 56495 45
rect 56525 15 56535 45
rect 56565 15 56575 45
rect 56605 15 56765 45
rect 56795 15 56845 45
rect 56875 15 56885 45
rect 56915 15 56925 45
rect 56955 15 57195 45
rect 57225 15 57235 45
rect 57265 15 57275 45
rect 57305 15 57545 45
rect 57575 15 57585 45
rect 57615 15 57625 45
rect 57655 15 57895 45
rect 57925 15 57935 45
rect 57965 15 57975 45
rect 58005 15 58245 45
rect 58275 15 58285 45
rect 58315 15 58325 45
rect 58355 15 58535 45
rect 58565 15 58595 45
rect 58625 15 58635 45
rect 58665 15 58675 45
rect 58705 15 58735 45
rect 58765 15 58945 45
rect 58975 15 58985 45
rect 59015 15 59025 45
rect 59055 15 59295 45
rect 59325 15 59335 45
rect 59365 15 59375 45
rect 59405 15 59645 45
rect 59675 15 59685 45
rect 59715 15 59725 45
rect 59755 15 59995 45
rect 60025 15 60035 45
rect 60065 15 60075 45
rect 60105 15 60345 45
rect 60375 15 60385 45
rect 60415 15 60425 45
rect 60455 15 60695 45
rect 60725 15 60735 45
rect 60765 15 60775 45
rect 60805 15 61045 45
rect 61075 15 61085 45
rect 61115 15 61125 45
rect 61155 15 61160 45
rect 52640 10 61160 15
<< via2 >>
rect 54610 3370 54640 3400
rect 59160 3370 59190 3400
rect 54195 1680 54225 1710
rect 54245 1680 54275 1710
rect 54295 1680 54325 1710
rect 54345 1680 54375 1710
rect 54395 1680 54425 1710
rect 54195 1630 54225 1660
rect 54245 1630 54275 1660
rect 54295 1630 54325 1660
rect 54345 1630 54375 1660
rect 54395 1630 54425 1660
rect 54195 1580 54225 1610
rect 54245 1580 54275 1610
rect 54295 1580 54325 1610
rect 54345 1580 54375 1610
rect 54395 1580 54425 1610
rect 59375 1680 59405 1710
rect 59425 1680 59455 1710
rect 59475 1680 59505 1710
rect 59525 1680 59555 1710
rect 59575 1680 59605 1710
rect 59375 1630 59405 1660
rect 59425 1630 59455 1660
rect 59475 1630 59505 1660
rect 59525 1630 59555 1660
rect 59575 1630 59605 1660
rect 59375 1580 59405 1610
rect 59425 1580 59455 1610
rect 59475 1580 59505 1610
rect 59525 1580 59555 1610
rect 59575 1580 59605 1610
<< metal3 >>
rect 52410 5870 52640 5955
rect 52760 5870 52990 5955
rect 53110 5870 53340 5955
rect 52410 5820 53340 5870
rect 52410 5725 52640 5820
rect 52760 5725 52990 5820
rect 53110 5725 53340 5820
rect 53460 5725 53690 5955
rect 53810 5725 54040 5955
rect 54160 5725 54390 5955
rect 54510 5725 54740 5955
rect 54860 5725 55090 5955
rect 55210 5725 55440 5955
rect 55560 5725 55790 5955
rect 55910 5725 56140 5955
rect 56260 5725 56490 5955
rect 56610 5725 56840 5955
rect 56960 5725 57190 5955
rect 57310 5725 57540 5955
rect 57660 5725 57890 5955
rect 58010 5725 58240 5955
rect 58360 5725 58590 5955
rect 58710 5725 58940 5955
rect 59060 5725 59290 5955
rect 59410 5725 59640 5955
rect 59760 5725 59990 5955
rect 60110 5725 60340 5955
rect 60460 5870 60690 5955
rect 60810 5870 61040 5955
rect 61160 5870 61390 5955
rect 60460 5820 61390 5870
rect 60460 5725 60690 5820
rect 60810 5725 61040 5820
rect 61160 5725 61390 5820
rect 53200 5605 53250 5725
rect 53550 5605 53600 5725
rect 53900 5605 53950 5725
rect 54250 5605 54300 5725
rect 54600 5605 54650 5725
rect 54950 5605 55000 5725
rect 55300 5605 55350 5725
rect 55650 5605 55700 5725
rect 56000 5605 56050 5725
rect 56350 5605 56400 5725
rect 56700 5605 56750 5725
rect 57050 5605 57100 5725
rect 57400 5605 57450 5725
rect 57750 5605 57800 5725
rect 58100 5605 58150 5725
rect 58450 5605 58500 5725
rect 58800 5605 58850 5725
rect 59150 5605 59200 5725
rect 59500 5605 59550 5725
rect 59850 5605 59900 5725
rect 60200 5605 60250 5725
rect 60550 5605 60600 5725
rect 52410 5520 52640 5605
rect 52760 5520 52990 5605
rect 53110 5520 53340 5605
rect 53460 5520 53690 5605
rect 53810 5520 54040 5605
rect 54160 5520 54390 5605
rect 54510 5520 54740 5605
rect 54860 5520 55090 5605
rect 55210 5520 55440 5605
rect 55560 5520 55790 5605
rect 55910 5520 56140 5605
rect 56260 5520 56490 5605
rect 56610 5520 56840 5605
rect 52410 5470 56840 5520
rect 52410 5375 52640 5470
rect 52760 5375 52990 5470
rect 53110 5375 53340 5470
rect 53460 5375 53690 5470
rect 53810 5375 54040 5470
rect 54160 5375 54390 5470
rect 54510 5375 54740 5470
rect 54860 5375 55090 5470
rect 55210 5375 55440 5470
rect 55560 5375 55790 5470
rect 55910 5375 56140 5470
rect 56260 5375 56490 5470
rect 56610 5375 56840 5470
rect 56960 5520 57190 5605
rect 57310 5520 57540 5605
rect 57660 5520 57890 5605
rect 58010 5520 58240 5605
rect 58360 5520 58590 5605
rect 58710 5520 58940 5605
rect 59060 5520 59290 5605
rect 59410 5520 59640 5605
rect 59760 5520 59990 5605
rect 60110 5520 60340 5605
rect 60460 5520 60690 5605
rect 60810 5520 61040 5605
rect 61160 5520 61390 5605
rect 56960 5470 61390 5520
rect 56960 5375 57190 5470
rect 57310 5375 57540 5470
rect 57660 5375 57890 5470
rect 58010 5375 58240 5470
rect 58360 5375 58590 5470
rect 58710 5375 58940 5470
rect 59060 5375 59290 5470
rect 59410 5375 59640 5470
rect 59760 5375 59990 5470
rect 60110 5375 60340 5470
rect 60460 5375 60690 5470
rect 60810 5375 61040 5470
rect 61160 5375 61390 5470
rect 53200 5255 53250 5375
rect 54250 5255 54300 5375
rect 54600 5255 54650 5375
rect 54950 5255 55000 5375
rect 55300 5255 55350 5375
rect 55650 5255 55700 5375
rect 56000 5255 56050 5375
rect 56350 5255 56400 5375
rect 56700 5255 56750 5375
rect 57050 5255 57100 5375
rect 57400 5255 57450 5375
rect 57750 5255 57800 5375
rect 58100 5255 58150 5375
rect 58450 5255 58500 5375
rect 58800 5255 58850 5375
rect 59150 5255 59200 5375
rect 59500 5255 59550 5375
rect 60550 5255 60600 5375
rect 52410 5170 52640 5255
rect 52760 5170 52990 5255
rect 53110 5170 53340 5255
rect 53460 5170 53690 5255
rect 53810 5170 54040 5255
rect 52410 5120 54040 5170
rect 52410 5025 52640 5120
rect 52760 5025 52990 5120
rect 53110 5025 53340 5120
rect 53460 5025 53690 5120
rect 53810 5025 54040 5120
rect 54160 5025 54390 5255
rect 54510 5025 54740 5255
rect 54860 5025 55090 5255
rect 55210 5025 55440 5255
rect 55560 5025 55790 5255
rect 55910 5025 56140 5255
rect 56260 5025 56490 5255
rect 56610 5025 56840 5255
rect 56960 5025 57190 5255
rect 57310 5025 57540 5255
rect 57660 5025 57890 5255
rect 58010 5025 58240 5255
rect 58360 5025 58590 5255
rect 58710 5025 58940 5255
rect 59060 5025 59290 5255
rect 59410 5025 59640 5255
rect 59760 5170 59990 5255
rect 60110 5170 60340 5255
rect 60460 5170 60690 5255
rect 60810 5170 61040 5255
rect 61160 5170 61390 5255
rect 59760 5120 61390 5170
rect 59760 5025 59990 5120
rect 60110 5025 60340 5120
rect 60460 5025 60690 5120
rect 60810 5025 61040 5120
rect 61160 5025 61390 5120
rect 53200 4905 53250 5025
rect 54250 4905 54300 5025
rect 54600 4905 54650 5025
rect 54950 4905 55000 5025
rect 55300 4905 55350 5025
rect 55650 4905 55700 5025
rect 58100 4905 58150 5025
rect 58450 4905 58500 5025
rect 58800 4905 58850 5025
rect 59150 4905 59200 5025
rect 59500 4905 59550 5025
rect 60550 4905 60600 5025
rect 52410 4820 52640 4905
rect 52760 4820 52990 4905
rect 53110 4820 53340 4905
rect 53460 4820 53690 4905
rect 53810 4820 54040 4905
rect 52410 4770 54040 4820
rect 52410 4675 52640 4770
rect 52760 4675 52990 4770
rect 53110 4675 53340 4770
rect 53460 4675 53690 4770
rect 53810 4675 54040 4770
rect 54160 4675 54390 4905
rect 54510 4675 54740 4905
rect 54860 4675 55090 4905
rect 55210 4675 55440 4905
rect 55560 4675 55790 4905
rect 58010 4675 58240 4905
rect 58360 4675 58590 4905
rect 58710 4675 58940 4905
rect 59060 4675 59290 4905
rect 59410 4675 59640 4905
rect 59760 4820 59990 4905
rect 60110 4820 60340 4905
rect 60460 4820 60690 4905
rect 60810 4820 61040 4905
rect 61160 4820 61390 4905
rect 59760 4770 61390 4820
rect 59760 4675 59990 4770
rect 60110 4675 60340 4770
rect 60460 4675 60690 4770
rect 60810 4675 61040 4770
rect 61160 4675 61390 4770
rect 53200 4555 53250 4675
rect 52410 4470 52640 4555
rect 52760 4470 52990 4555
rect 53110 4470 53340 4555
rect 53460 4470 53690 4555
rect 53810 4470 54040 4555
rect 52410 4420 54040 4470
rect 52410 4325 52640 4420
rect 52760 4325 52990 4420
rect 53110 4325 53340 4420
rect 53460 4325 53690 4420
rect 53810 4325 54040 4420
rect 53200 4205 53250 4325
rect 52410 4120 52640 4205
rect 52760 4120 52990 4205
rect 53110 4120 53340 4205
rect 53460 4120 53690 4205
rect 53810 4120 54040 4205
rect 52410 4070 54040 4120
rect 52410 3975 52640 4070
rect 52760 3975 52990 4070
rect 53110 3975 53340 4070
rect 53460 3975 53690 4070
rect 53810 3975 54040 4070
rect 53200 3855 53250 3975
rect 52410 3770 52640 3855
rect 52760 3770 52990 3855
rect 53110 3770 53340 3855
rect 53460 3770 53690 3855
rect 53810 3770 54040 3855
rect 52410 3720 54040 3770
rect 52410 3625 52640 3720
rect 52760 3625 52990 3720
rect 53110 3625 53340 3720
rect 53460 3625 53690 3720
rect 53810 3625 54040 3720
rect 53200 3505 53250 3625
rect 52410 3420 52640 3505
rect 52760 3420 52990 3505
rect 53110 3420 53340 3505
rect 53460 3420 53690 3505
rect 53810 3420 54040 3505
rect 52410 3370 54040 3420
rect 52410 3275 52640 3370
rect 52760 3275 52990 3370
rect 53110 3275 53340 3370
rect 53460 3275 53690 3370
rect 53810 3275 54040 3370
rect 54605 3400 54645 4675
rect 54605 3370 54610 3400
rect 54640 3370 54645 3400
rect 54605 3365 54645 3370
rect 59155 3400 59195 4675
rect 60550 4555 60600 4675
rect 59760 4470 59990 4555
rect 60110 4470 60340 4555
rect 60460 4470 60690 4555
rect 60810 4470 61040 4555
rect 61160 4470 61390 4555
rect 59760 4420 61390 4470
rect 59760 4325 59990 4420
rect 60110 4325 60340 4420
rect 60460 4325 60690 4420
rect 60810 4325 61040 4420
rect 61160 4325 61390 4420
rect 60550 4205 60600 4325
rect 59760 4120 59990 4205
rect 60110 4120 60340 4205
rect 60460 4120 60690 4205
rect 60810 4120 61040 4205
rect 61160 4120 61390 4205
rect 59760 4070 61390 4120
rect 59760 3975 59990 4070
rect 60110 3975 60340 4070
rect 60460 3975 60690 4070
rect 60810 3975 61040 4070
rect 61160 3975 61390 4070
rect 60550 3855 60600 3975
rect 59760 3770 59990 3855
rect 60110 3770 60340 3855
rect 60460 3770 60690 3855
rect 60810 3770 61040 3855
rect 61160 3770 61390 3855
rect 59760 3720 61390 3770
rect 59760 3625 59990 3720
rect 60110 3625 60340 3720
rect 60460 3625 60690 3720
rect 60810 3625 61040 3720
rect 61160 3625 61390 3720
rect 60550 3505 60600 3625
rect 59155 3370 59160 3400
rect 59190 3370 59195 3400
rect 59155 3365 59195 3370
rect 59760 3420 59990 3505
rect 60110 3420 60340 3505
rect 60460 3420 60690 3505
rect 60810 3420 61040 3505
rect 61160 3420 61390 3505
rect 59760 3370 61390 3420
rect 59760 3275 59990 3370
rect 60110 3275 60340 3370
rect 60460 3275 60690 3370
rect 60810 3275 61040 3370
rect 61160 3275 61390 3370
rect 53200 3155 53250 3275
rect 60550 3155 60600 3275
rect 52410 3070 52640 3155
rect 52760 3070 52990 3155
rect 53110 3070 53340 3155
rect 53460 3070 53690 3155
rect 53810 3070 54040 3155
rect 52410 3020 54040 3070
rect 52410 2925 52640 3020
rect 52760 2925 52990 3020
rect 53110 2925 53340 3020
rect 53460 2925 53690 3020
rect 53810 2925 54040 3020
rect 59760 3070 59990 3155
rect 60110 3070 60340 3155
rect 60460 3070 60690 3155
rect 60810 3070 61040 3155
rect 61160 3070 61390 3155
rect 59760 3020 61390 3070
rect 59760 2925 59990 3020
rect 60110 2925 60340 3020
rect 60460 2925 60690 3020
rect 60810 2925 61040 3020
rect 61160 2925 61390 3020
rect 53200 2805 53250 2925
rect 60550 2805 60600 2925
rect 52410 2720 52640 2805
rect 52760 2720 52990 2805
rect 53110 2720 53340 2805
rect 53460 2720 53690 2805
rect 53810 2720 54040 2805
rect 52410 2670 54040 2720
rect 52410 2575 52640 2670
rect 52760 2575 52990 2670
rect 53110 2575 53340 2670
rect 53460 2575 53690 2670
rect 53810 2575 54040 2670
rect 59760 2720 59990 2805
rect 60110 2720 60340 2805
rect 60460 2720 60690 2805
rect 60810 2720 61040 2805
rect 61160 2720 61390 2805
rect 59760 2670 61390 2720
rect 59760 2575 59990 2670
rect 60110 2575 60340 2670
rect 60460 2575 60690 2670
rect 60810 2575 61040 2670
rect 61160 2575 61390 2670
rect 53200 2455 53250 2575
rect 60550 2455 60600 2575
rect 52410 2370 52640 2455
rect 52760 2370 52990 2455
rect 53110 2370 53340 2455
rect 53460 2370 53690 2455
rect 53810 2370 54040 2455
rect 52410 2320 54040 2370
rect 52410 2225 52640 2320
rect 52760 2225 52990 2320
rect 53110 2225 53340 2320
rect 53460 2225 53690 2320
rect 53810 2225 54040 2320
rect 59760 2370 59990 2455
rect 60110 2370 60340 2455
rect 60460 2370 60690 2455
rect 60810 2370 61040 2455
rect 61160 2370 61390 2455
rect 59760 2320 61390 2370
rect 59760 2225 59990 2320
rect 60110 2225 60340 2320
rect 60460 2225 60690 2320
rect 60810 2225 61040 2320
rect 61160 2225 61390 2320
rect 53200 2105 53250 2225
rect 60550 2105 60600 2225
rect 52410 2020 52640 2105
rect 52760 2020 52990 2105
rect 53110 2020 53340 2105
rect 53460 2020 53690 2105
rect 53810 2020 54040 2105
rect 52410 1970 54040 2020
rect 52410 1875 52640 1970
rect 52760 1875 52990 1970
rect 53110 1875 53340 1970
rect 53460 1875 53690 1970
rect 53810 1875 54040 1970
rect 59760 2020 59990 2105
rect 60110 2020 60340 2105
rect 60460 2020 60690 2105
rect 60810 2020 61040 2105
rect 61160 2020 61390 2105
rect 59760 1970 61390 2020
rect 59760 1875 59990 1970
rect 60110 1875 60340 1970
rect 60460 1875 60690 1970
rect 60810 1875 61040 1970
rect 61160 1875 61390 1970
rect 53200 1755 53250 1875
rect 60550 1755 60600 1875
rect 52410 1670 52640 1755
rect 52760 1670 52990 1755
rect 53110 1670 53340 1755
rect 53460 1670 53690 1755
rect 53810 1670 54040 1755
rect 52410 1620 54040 1670
rect 52410 1525 52640 1620
rect 52760 1525 52990 1620
rect 53110 1525 53340 1620
rect 53460 1525 53690 1620
rect 53810 1525 54040 1620
rect 54185 1715 54435 1720
rect 54185 1675 54190 1715
rect 54230 1675 54240 1715
rect 54280 1675 54290 1715
rect 54330 1675 54340 1715
rect 54380 1675 54390 1715
rect 54430 1675 54435 1715
rect 54185 1665 54435 1675
rect 54185 1625 54190 1665
rect 54230 1625 54240 1665
rect 54280 1625 54290 1665
rect 54330 1625 54340 1665
rect 54380 1625 54390 1665
rect 54430 1625 54435 1665
rect 54185 1615 54435 1625
rect 54185 1575 54190 1615
rect 54230 1575 54240 1615
rect 54280 1575 54290 1615
rect 54330 1575 54340 1615
rect 54380 1575 54390 1615
rect 54430 1575 54435 1615
rect 54185 1570 54435 1575
rect 59365 1715 59615 1720
rect 59365 1675 59370 1715
rect 59410 1675 59420 1715
rect 59460 1675 59470 1715
rect 59510 1675 59520 1715
rect 59560 1675 59570 1715
rect 59610 1675 59615 1715
rect 59365 1665 59615 1675
rect 59365 1625 59370 1665
rect 59410 1625 59420 1665
rect 59460 1625 59470 1665
rect 59510 1625 59520 1665
rect 59560 1625 59570 1665
rect 59610 1625 59615 1665
rect 59365 1615 59615 1625
rect 59365 1575 59370 1615
rect 59410 1575 59420 1615
rect 59460 1575 59470 1615
rect 59510 1575 59520 1615
rect 59560 1575 59570 1615
rect 59610 1575 59615 1615
rect 59365 1570 59615 1575
rect 59760 1670 59990 1755
rect 60110 1670 60340 1755
rect 60460 1670 60690 1755
rect 60810 1670 61040 1755
rect 61160 1670 61390 1755
rect 59760 1620 61390 1670
rect 59760 1525 59990 1620
rect 60110 1525 60340 1620
rect 60460 1525 60690 1620
rect 60810 1525 61040 1620
rect 61160 1525 61390 1620
rect 53200 1405 53250 1525
rect 60550 1405 60600 1525
rect 52410 1320 52640 1405
rect 52760 1320 52990 1405
rect 53110 1320 53340 1405
rect 53460 1320 53690 1405
rect 53810 1320 54040 1405
rect 52410 1270 54040 1320
rect 52410 1175 52640 1270
rect 52760 1175 52990 1270
rect 53110 1175 53340 1270
rect 53460 1175 53690 1270
rect 53810 1175 54040 1270
rect 59760 1320 59990 1405
rect 60110 1320 60340 1405
rect 60460 1320 60690 1405
rect 60810 1320 61040 1405
rect 61160 1320 61390 1405
rect 59760 1270 61390 1320
rect 59760 1175 59990 1270
rect 60110 1175 60340 1270
rect 60460 1175 60690 1270
rect 60810 1175 61040 1270
rect 61160 1175 61390 1270
rect 53200 1055 53250 1175
rect 60550 1055 60600 1175
rect 52410 970 52640 1055
rect 52760 970 52990 1055
rect 53110 970 53340 1055
rect 53460 970 53690 1055
rect 53810 970 54040 1055
rect 52410 920 54040 970
rect 52410 825 52640 920
rect 52760 825 52990 920
rect 53110 825 53340 920
rect 53460 825 53690 920
rect 53810 825 54040 920
rect 59760 970 59990 1055
rect 60110 970 60340 1055
rect 60460 970 60690 1055
rect 60810 970 61040 1055
rect 61160 970 61390 1055
rect 59760 920 61390 970
rect 59760 825 59990 920
rect 60110 825 60340 920
rect 60460 825 60690 920
rect 60810 825 61040 920
rect 61160 825 61390 920
rect 53200 705 53250 825
rect 60550 705 60600 825
rect 52410 620 52640 705
rect 52760 620 52990 705
rect 53110 620 53340 705
rect 53460 620 53690 705
rect 53810 620 54040 705
rect 52410 570 54040 620
rect 52410 475 52640 570
rect 52760 475 52990 570
rect 53110 475 53340 570
rect 53460 475 53690 570
rect 53810 475 54040 570
rect 59760 620 59990 705
rect 60110 620 60340 705
rect 60460 620 60690 705
rect 60810 620 61040 705
rect 61160 620 61390 705
rect 59760 570 61390 620
rect 59760 475 59990 570
rect 60110 475 60340 570
rect 60460 475 60690 570
rect 60810 475 61040 570
rect 61160 475 61390 570
rect 53200 355 53250 475
rect 60550 355 60600 475
rect 52410 270 52640 355
rect 52760 270 52990 355
rect 53110 270 53340 355
rect 53460 270 53690 355
rect 53810 270 54040 355
rect 52410 220 54040 270
rect 52410 125 52640 220
rect 52760 125 52990 220
rect 53110 125 53340 220
rect 53460 125 53690 220
rect 53810 125 54040 220
rect 59760 270 59990 355
rect 60110 270 60340 355
rect 60460 270 60690 355
rect 60810 270 61040 355
rect 61160 270 61390 355
rect 59760 220 61390 270
rect 59760 125 59990 220
rect 60110 125 60340 220
rect 60460 125 60690 220
rect 60810 125 61040 220
rect 61160 125 61390 220
rect 53200 5 53250 125
rect 60550 5 60600 125
rect 52410 -80 52640 5
rect 52760 -80 52990 5
rect 53110 -80 53340 5
rect 53460 -80 53690 5
rect 53810 -80 54040 5
rect 54160 -80 54390 5
rect 54510 -80 54740 5
rect 54860 -80 55090 5
rect 55210 -80 55440 5
rect 55560 -80 55790 5
rect 55910 -80 56140 5
rect 56260 -80 56490 5
rect 56610 -80 56840 5
rect 52410 -130 56840 -80
rect 52410 -225 52640 -130
rect 52760 -225 52990 -130
rect 53110 -225 53340 -130
rect 53460 -225 53690 -130
rect 53810 -225 54040 -130
rect 54160 -225 54390 -130
rect 54510 -225 54740 -130
rect 54860 -225 55090 -130
rect 55210 -225 55440 -130
rect 55560 -225 55790 -130
rect 55910 -225 56140 -130
rect 56260 -225 56490 -130
rect 56610 -225 56840 -130
rect 56960 -80 57190 5
rect 57310 -80 57540 5
rect 57660 -80 57890 5
rect 58010 -80 58240 5
rect 58360 -80 58590 5
rect 58710 -80 58940 5
rect 59060 -80 59290 5
rect 59410 -80 59640 5
rect 59760 -80 59990 5
rect 60110 -80 60340 5
rect 60460 -80 60690 5
rect 60810 -80 61040 5
rect 61160 -80 61390 5
rect 56960 -130 61390 -80
rect 56960 -225 57190 -130
rect 57310 -225 57540 -130
rect 57660 -225 57890 -130
rect 58010 -225 58240 -130
rect 58360 -225 58590 -130
rect 58710 -225 58940 -130
rect 59060 -225 59290 -130
rect 59410 -225 59640 -130
rect 59760 -225 59990 -130
rect 60110 -225 60340 -130
rect 60460 -225 60690 -130
rect 60810 -225 61040 -130
rect 61160 -225 61390 -130
rect 53200 -345 53250 -225
rect 53550 -345 53600 -225
rect 53900 -345 53950 -225
rect 54250 -345 54300 -225
rect 54600 -345 54650 -225
rect 54950 -345 55000 -225
rect 55300 -345 55350 -225
rect 55650 -345 55700 -225
rect 56000 -345 56050 -225
rect 56350 -345 56400 -225
rect 56700 -345 56750 -225
rect 57050 -345 57100 -225
rect 57400 -345 57450 -225
rect 57750 -345 57800 -225
rect 58100 -345 58150 -225
rect 58450 -345 58500 -225
rect 58800 -345 58850 -225
rect 59150 -345 59200 -225
rect 59500 -345 59550 -225
rect 59850 -345 59900 -225
rect 60200 -345 60250 -225
rect 60550 -345 60600 -225
rect 52410 -430 52640 -345
rect 52760 -430 52990 -345
rect 53110 -430 53340 -345
rect 52410 -480 53340 -430
rect 52410 -575 52640 -480
rect 52760 -575 52990 -480
rect 53110 -575 53340 -480
rect 53460 -575 53690 -345
rect 53810 -575 54040 -345
rect 54160 -575 54390 -345
rect 54510 -575 54740 -345
rect 54860 -575 55090 -345
rect 55210 -575 55440 -345
rect 55560 -575 55790 -345
rect 55910 -575 56140 -345
rect 56260 -575 56490 -345
rect 56610 -575 56840 -345
rect 56960 -575 57190 -345
rect 57310 -575 57540 -345
rect 57660 -575 57890 -345
rect 58010 -575 58240 -345
rect 58360 -575 58590 -345
rect 58710 -575 58940 -345
rect 59060 -575 59290 -345
rect 59410 -575 59640 -345
rect 59760 -575 59990 -345
rect 60110 -575 60340 -345
rect 60460 -430 60690 -345
rect 60810 -430 61040 -345
rect 61160 -430 61390 -345
rect 60460 -480 61390 -430
rect 60460 -575 60690 -480
rect 60810 -575 61040 -480
rect 61160 -575 61390 -480
<< via3 >>
rect 54190 1710 54230 1715
rect 54190 1680 54195 1710
rect 54195 1680 54225 1710
rect 54225 1680 54230 1710
rect 54190 1675 54230 1680
rect 54240 1710 54280 1715
rect 54240 1680 54245 1710
rect 54245 1680 54275 1710
rect 54275 1680 54280 1710
rect 54240 1675 54280 1680
rect 54290 1710 54330 1715
rect 54290 1680 54295 1710
rect 54295 1680 54325 1710
rect 54325 1680 54330 1710
rect 54290 1675 54330 1680
rect 54340 1710 54380 1715
rect 54340 1680 54345 1710
rect 54345 1680 54375 1710
rect 54375 1680 54380 1710
rect 54340 1675 54380 1680
rect 54390 1710 54430 1715
rect 54390 1680 54395 1710
rect 54395 1680 54425 1710
rect 54425 1680 54430 1710
rect 54390 1675 54430 1680
rect 54190 1660 54230 1665
rect 54190 1630 54195 1660
rect 54195 1630 54225 1660
rect 54225 1630 54230 1660
rect 54190 1625 54230 1630
rect 54240 1660 54280 1665
rect 54240 1630 54245 1660
rect 54245 1630 54275 1660
rect 54275 1630 54280 1660
rect 54240 1625 54280 1630
rect 54290 1660 54330 1665
rect 54290 1630 54295 1660
rect 54295 1630 54325 1660
rect 54325 1630 54330 1660
rect 54290 1625 54330 1630
rect 54340 1660 54380 1665
rect 54340 1630 54345 1660
rect 54345 1630 54375 1660
rect 54375 1630 54380 1660
rect 54340 1625 54380 1630
rect 54390 1660 54430 1665
rect 54390 1630 54395 1660
rect 54395 1630 54425 1660
rect 54425 1630 54430 1660
rect 54390 1625 54430 1630
rect 54190 1610 54230 1615
rect 54190 1580 54195 1610
rect 54195 1580 54225 1610
rect 54225 1580 54230 1610
rect 54190 1575 54230 1580
rect 54240 1610 54280 1615
rect 54240 1580 54245 1610
rect 54245 1580 54275 1610
rect 54275 1580 54280 1610
rect 54240 1575 54280 1580
rect 54290 1610 54330 1615
rect 54290 1580 54295 1610
rect 54295 1580 54325 1610
rect 54325 1580 54330 1610
rect 54290 1575 54330 1580
rect 54340 1610 54380 1615
rect 54340 1580 54345 1610
rect 54345 1580 54375 1610
rect 54375 1580 54380 1610
rect 54340 1575 54380 1580
rect 54390 1610 54430 1615
rect 54390 1580 54395 1610
rect 54395 1580 54425 1610
rect 54425 1580 54430 1610
rect 54390 1575 54430 1580
rect 59370 1710 59410 1715
rect 59370 1680 59375 1710
rect 59375 1680 59405 1710
rect 59405 1680 59410 1710
rect 59370 1675 59410 1680
rect 59420 1710 59460 1715
rect 59420 1680 59425 1710
rect 59425 1680 59455 1710
rect 59455 1680 59460 1710
rect 59420 1675 59460 1680
rect 59470 1710 59510 1715
rect 59470 1680 59475 1710
rect 59475 1680 59505 1710
rect 59505 1680 59510 1710
rect 59470 1675 59510 1680
rect 59520 1710 59560 1715
rect 59520 1680 59525 1710
rect 59525 1680 59555 1710
rect 59555 1680 59560 1710
rect 59520 1675 59560 1680
rect 59570 1710 59610 1715
rect 59570 1680 59575 1710
rect 59575 1680 59605 1710
rect 59605 1680 59610 1710
rect 59570 1675 59610 1680
rect 59370 1660 59410 1665
rect 59370 1630 59375 1660
rect 59375 1630 59405 1660
rect 59405 1630 59410 1660
rect 59370 1625 59410 1630
rect 59420 1660 59460 1665
rect 59420 1630 59425 1660
rect 59425 1630 59455 1660
rect 59455 1630 59460 1660
rect 59420 1625 59460 1630
rect 59470 1660 59510 1665
rect 59470 1630 59475 1660
rect 59475 1630 59505 1660
rect 59505 1630 59510 1660
rect 59470 1625 59510 1630
rect 59520 1660 59560 1665
rect 59520 1630 59525 1660
rect 59525 1630 59555 1660
rect 59555 1630 59560 1660
rect 59520 1625 59560 1630
rect 59570 1660 59610 1665
rect 59570 1630 59575 1660
rect 59575 1630 59605 1660
rect 59605 1630 59610 1660
rect 59570 1625 59610 1630
rect 59370 1610 59410 1615
rect 59370 1580 59375 1610
rect 59375 1580 59405 1610
rect 59405 1580 59410 1610
rect 59370 1575 59410 1580
rect 59420 1610 59460 1615
rect 59420 1580 59425 1610
rect 59425 1580 59455 1610
rect 59455 1580 59460 1610
rect 59420 1575 59460 1580
rect 59470 1610 59510 1615
rect 59470 1580 59475 1610
rect 59475 1580 59505 1610
rect 59505 1580 59510 1610
rect 59470 1575 59510 1580
rect 59520 1610 59560 1615
rect 59520 1580 59525 1610
rect 59525 1580 59555 1610
rect 59555 1580 59560 1610
rect 59520 1575 59560 1580
rect 59570 1610 59610 1615
rect 59570 1580 59575 1610
rect 59575 1580 59605 1610
rect 59605 1580 59610 1610
rect 59570 1575 59610 1580
<< mimcap >>
rect 52425 5865 52625 5940
rect 52425 5825 52505 5865
rect 52545 5825 52625 5865
rect 52425 5740 52625 5825
rect 52775 5865 52975 5940
rect 52775 5825 52855 5865
rect 52895 5825 52975 5865
rect 52775 5740 52975 5825
rect 53125 5865 53325 5940
rect 53125 5825 53205 5865
rect 53245 5825 53325 5865
rect 53125 5740 53325 5825
rect 53475 5865 53675 5940
rect 53475 5825 53555 5865
rect 53595 5825 53675 5865
rect 53475 5740 53675 5825
rect 53825 5865 54025 5940
rect 53825 5825 53905 5865
rect 53945 5825 54025 5865
rect 53825 5740 54025 5825
rect 54175 5865 54375 5940
rect 54175 5825 54255 5865
rect 54295 5825 54375 5865
rect 54175 5740 54375 5825
rect 54525 5865 54725 5940
rect 54525 5825 54605 5865
rect 54645 5825 54725 5865
rect 54525 5740 54725 5825
rect 54875 5865 55075 5940
rect 54875 5825 54955 5865
rect 54995 5825 55075 5865
rect 54875 5740 55075 5825
rect 55225 5865 55425 5940
rect 55225 5825 55305 5865
rect 55345 5825 55425 5865
rect 55225 5740 55425 5825
rect 55575 5865 55775 5940
rect 55575 5825 55655 5865
rect 55695 5825 55775 5865
rect 55575 5740 55775 5825
rect 55925 5865 56125 5940
rect 55925 5825 56005 5865
rect 56045 5825 56125 5865
rect 55925 5740 56125 5825
rect 56275 5865 56475 5940
rect 56275 5825 56355 5865
rect 56395 5825 56475 5865
rect 56275 5740 56475 5825
rect 56625 5865 56825 5940
rect 56625 5825 56705 5865
rect 56745 5825 56825 5865
rect 56625 5740 56825 5825
rect 56975 5865 57175 5940
rect 56975 5825 57055 5865
rect 57095 5825 57175 5865
rect 56975 5740 57175 5825
rect 57325 5865 57525 5940
rect 57325 5825 57405 5865
rect 57445 5825 57525 5865
rect 57325 5740 57525 5825
rect 57675 5865 57875 5940
rect 57675 5825 57755 5865
rect 57795 5825 57875 5865
rect 57675 5740 57875 5825
rect 58025 5865 58225 5940
rect 58025 5825 58105 5865
rect 58145 5825 58225 5865
rect 58025 5740 58225 5825
rect 58375 5865 58575 5940
rect 58375 5825 58455 5865
rect 58495 5825 58575 5865
rect 58375 5740 58575 5825
rect 58725 5865 58925 5940
rect 58725 5825 58805 5865
rect 58845 5825 58925 5865
rect 58725 5740 58925 5825
rect 59075 5865 59275 5940
rect 59075 5825 59155 5865
rect 59195 5825 59275 5865
rect 59075 5740 59275 5825
rect 59425 5865 59625 5940
rect 59425 5825 59505 5865
rect 59545 5825 59625 5865
rect 59425 5740 59625 5825
rect 59775 5865 59975 5940
rect 59775 5825 59855 5865
rect 59895 5825 59975 5865
rect 59775 5740 59975 5825
rect 60125 5865 60325 5940
rect 60125 5825 60205 5865
rect 60245 5825 60325 5865
rect 60125 5740 60325 5825
rect 60475 5865 60675 5940
rect 60475 5825 60555 5865
rect 60595 5825 60675 5865
rect 60475 5740 60675 5825
rect 60825 5865 61025 5940
rect 60825 5825 60905 5865
rect 60945 5825 61025 5865
rect 60825 5740 61025 5825
rect 61175 5865 61375 5940
rect 61175 5825 61255 5865
rect 61295 5825 61375 5865
rect 61175 5740 61375 5825
rect 52425 5515 52625 5590
rect 52425 5475 52505 5515
rect 52545 5475 52625 5515
rect 52425 5390 52625 5475
rect 52775 5515 52975 5590
rect 52775 5475 52855 5515
rect 52895 5475 52975 5515
rect 52775 5390 52975 5475
rect 53125 5515 53325 5590
rect 53125 5475 53205 5515
rect 53245 5475 53325 5515
rect 53125 5390 53325 5475
rect 53475 5515 53675 5590
rect 53475 5475 53555 5515
rect 53595 5475 53675 5515
rect 53475 5390 53675 5475
rect 53825 5515 54025 5590
rect 53825 5475 53905 5515
rect 53945 5475 54025 5515
rect 53825 5390 54025 5475
rect 54175 5515 54375 5590
rect 54175 5475 54255 5515
rect 54295 5475 54375 5515
rect 54175 5390 54375 5475
rect 54525 5515 54725 5590
rect 54525 5475 54605 5515
rect 54645 5475 54725 5515
rect 54525 5390 54725 5475
rect 54875 5515 55075 5590
rect 54875 5475 54955 5515
rect 54995 5475 55075 5515
rect 54875 5390 55075 5475
rect 55225 5515 55425 5590
rect 55225 5475 55305 5515
rect 55345 5475 55425 5515
rect 55225 5390 55425 5475
rect 55575 5515 55775 5590
rect 55575 5475 55655 5515
rect 55695 5475 55775 5515
rect 55575 5390 55775 5475
rect 55925 5515 56125 5590
rect 55925 5475 56005 5515
rect 56045 5475 56125 5515
rect 55925 5390 56125 5475
rect 56275 5515 56475 5590
rect 56275 5475 56355 5515
rect 56395 5475 56475 5515
rect 56275 5390 56475 5475
rect 56625 5515 56825 5590
rect 56625 5475 56705 5515
rect 56745 5475 56825 5515
rect 56625 5390 56825 5475
rect 56975 5515 57175 5590
rect 56975 5475 57055 5515
rect 57095 5475 57175 5515
rect 56975 5390 57175 5475
rect 57325 5515 57525 5590
rect 57325 5475 57405 5515
rect 57445 5475 57525 5515
rect 57325 5390 57525 5475
rect 57675 5515 57875 5590
rect 57675 5475 57755 5515
rect 57795 5475 57875 5515
rect 57675 5390 57875 5475
rect 58025 5515 58225 5590
rect 58025 5475 58105 5515
rect 58145 5475 58225 5515
rect 58025 5390 58225 5475
rect 58375 5515 58575 5590
rect 58375 5475 58455 5515
rect 58495 5475 58575 5515
rect 58375 5390 58575 5475
rect 58725 5515 58925 5590
rect 58725 5475 58805 5515
rect 58845 5475 58925 5515
rect 58725 5390 58925 5475
rect 59075 5515 59275 5590
rect 59075 5475 59155 5515
rect 59195 5475 59275 5515
rect 59075 5390 59275 5475
rect 59425 5515 59625 5590
rect 59425 5475 59505 5515
rect 59545 5475 59625 5515
rect 59425 5390 59625 5475
rect 59775 5515 59975 5590
rect 59775 5475 59855 5515
rect 59895 5475 59975 5515
rect 59775 5390 59975 5475
rect 60125 5515 60325 5590
rect 60125 5475 60205 5515
rect 60245 5475 60325 5515
rect 60125 5390 60325 5475
rect 60475 5515 60675 5590
rect 60475 5475 60555 5515
rect 60595 5475 60675 5515
rect 60475 5390 60675 5475
rect 60825 5515 61025 5590
rect 60825 5475 60905 5515
rect 60945 5475 61025 5515
rect 60825 5390 61025 5475
rect 61175 5515 61375 5590
rect 61175 5475 61255 5515
rect 61295 5475 61375 5515
rect 61175 5390 61375 5475
rect 52425 5165 52625 5240
rect 52425 5125 52505 5165
rect 52545 5125 52625 5165
rect 52425 5040 52625 5125
rect 52775 5165 52975 5240
rect 52775 5125 52855 5165
rect 52895 5125 52975 5165
rect 52775 5040 52975 5125
rect 53125 5165 53325 5240
rect 53125 5125 53205 5165
rect 53245 5125 53325 5165
rect 53125 5040 53325 5125
rect 53475 5165 53675 5240
rect 53475 5125 53555 5165
rect 53595 5125 53675 5165
rect 53475 5040 53675 5125
rect 53825 5165 54025 5240
rect 53825 5125 53905 5165
rect 53945 5125 54025 5165
rect 53825 5040 54025 5125
rect 54175 5165 54375 5240
rect 54175 5125 54255 5165
rect 54295 5125 54375 5165
rect 54175 5040 54375 5125
rect 54525 5165 54725 5240
rect 54525 5125 54605 5165
rect 54645 5125 54725 5165
rect 54525 5040 54725 5125
rect 54875 5165 55075 5240
rect 54875 5125 54955 5165
rect 54995 5125 55075 5165
rect 54875 5040 55075 5125
rect 55225 5165 55425 5240
rect 55225 5125 55305 5165
rect 55345 5125 55425 5165
rect 55225 5040 55425 5125
rect 55575 5155 55775 5240
rect 55575 5115 55655 5155
rect 55695 5115 55775 5155
rect 55575 5040 55775 5115
rect 55925 5155 56125 5240
rect 55925 5115 56005 5155
rect 56045 5115 56125 5155
rect 55925 5040 56125 5115
rect 56275 5155 56475 5240
rect 56275 5115 56355 5155
rect 56395 5115 56475 5155
rect 56275 5040 56475 5115
rect 56625 5155 56825 5240
rect 56625 5115 56705 5155
rect 56745 5115 56825 5155
rect 56625 5040 56825 5115
rect 56975 5155 57175 5240
rect 56975 5115 57055 5155
rect 57095 5115 57175 5155
rect 56975 5040 57175 5115
rect 57325 5155 57525 5240
rect 57325 5115 57405 5155
rect 57445 5115 57525 5155
rect 57325 5040 57525 5115
rect 57675 5155 57875 5240
rect 57675 5115 57755 5155
rect 57795 5115 57875 5155
rect 57675 5040 57875 5115
rect 58025 5155 58225 5240
rect 58025 5115 58105 5155
rect 58145 5115 58225 5155
rect 58025 5040 58225 5115
rect 58375 5165 58575 5240
rect 58375 5125 58455 5165
rect 58495 5125 58575 5165
rect 58375 5040 58575 5125
rect 58725 5165 58925 5240
rect 58725 5125 58805 5165
rect 58845 5125 58925 5165
rect 58725 5040 58925 5125
rect 59075 5165 59275 5240
rect 59075 5125 59155 5165
rect 59195 5125 59275 5165
rect 59075 5040 59275 5125
rect 59425 5165 59625 5240
rect 59425 5125 59505 5165
rect 59545 5125 59625 5165
rect 59425 5040 59625 5125
rect 59775 5165 59975 5240
rect 59775 5125 59855 5165
rect 59895 5125 59975 5165
rect 59775 5040 59975 5125
rect 60125 5165 60325 5240
rect 60125 5125 60205 5165
rect 60245 5125 60325 5165
rect 60125 5040 60325 5125
rect 60475 5165 60675 5240
rect 60475 5125 60555 5165
rect 60595 5125 60675 5165
rect 60475 5040 60675 5125
rect 60825 5165 61025 5240
rect 60825 5125 60905 5165
rect 60945 5125 61025 5165
rect 60825 5040 61025 5125
rect 61175 5165 61375 5240
rect 61175 5125 61255 5165
rect 61295 5125 61375 5165
rect 61175 5040 61375 5125
rect 52425 4815 52625 4890
rect 52425 4775 52505 4815
rect 52545 4775 52625 4815
rect 52425 4690 52625 4775
rect 52775 4815 52975 4890
rect 52775 4775 52855 4815
rect 52895 4775 52975 4815
rect 52775 4690 52975 4775
rect 53125 4815 53325 4890
rect 53125 4775 53205 4815
rect 53245 4775 53325 4815
rect 53125 4690 53325 4775
rect 53475 4815 53675 4890
rect 53475 4775 53555 4815
rect 53595 4775 53675 4815
rect 53475 4690 53675 4775
rect 53825 4815 54025 4890
rect 53825 4775 53905 4815
rect 53945 4775 54025 4815
rect 53825 4690 54025 4775
rect 54175 4815 54375 4890
rect 54175 4775 54255 4815
rect 54295 4775 54375 4815
rect 54175 4690 54375 4775
rect 54525 4815 54725 4890
rect 54525 4775 54605 4815
rect 54645 4775 54725 4815
rect 54525 4690 54725 4775
rect 54875 4815 55075 4890
rect 54875 4775 54955 4815
rect 54995 4775 55075 4815
rect 54875 4690 55075 4775
rect 55225 4815 55425 4890
rect 55225 4775 55305 4815
rect 55345 4775 55425 4815
rect 55225 4690 55425 4775
rect 55575 4815 55775 4890
rect 55575 4775 55655 4815
rect 55695 4775 55775 4815
rect 55575 4690 55775 4775
rect 58025 4805 58225 4890
rect 58025 4765 58105 4805
rect 58145 4765 58225 4805
rect 58025 4690 58225 4765
rect 58375 4815 58575 4890
rect 58375 4775 58455 4815
rect 58495 4775 58575 4815
rect 58375 4690 58575 4775
rect 58725 4815 58925 4890
rect 58725 4775 58805 4815
rect 58845 4775 58925 4815
rect 58725 4690 58925 4775
rect 59075 4815 59275 4890
rect 59075 4775 59155 4815
rect 59195 4775 59275 4815
rect 59075 4690 59275 4775
rect 59425 4815 59625 4890
rect 59425 4775 59505 4815
rect 59545 4775 59625 4815
rect 59425 4690 59625 4775
rect 59775 4815 59975 4890
rect 59775 4775 59855 4815
rect 59895 4775 59975 4815
rect 59775 4690 59975 4775
rect 60125 4815 60325 4890
rect 60125 4775 60205 4815
rect 60245 4775 60325 4815
rect 60125 4690 60325 4775
rect 60475 4815 60675 4890
rect 60475 4775 60555 4815
rect 60595 4775 60675 4815
rect 60475 4690 60675 4775
rect 60825 4815 61025 4890
rect 60825 4775 60905 4815
rect 60945 4775 61025 4815
rect 60825 4690 61025 4775
rect 61175 4815 61375 4890
rect 61175 4775 61255 4815
rect 61295 4775 61375 4815
rect 61175 4690 61375 4775
rect 52425 4465 52625 4540
rect 52425 4425 52505 4465
rect 52545 4425 52625 4465
rect 52425 4340 52625 4425
rect 52775 4465 52975 4540
rect 52775 4425 52855 4465
rect 52895 4425 52975 4465
rect 52775 4340 52975 4425
rect 53125 4465 53325 4540
rect 53125 4425 53205 4465
rect 53245 4425 53325 4465
rect 53125 4340 53325 4425
rect 53475 4465 53675 4540
rect 53475 4425 53555 4465
rect 53595 4425 53675 4465
rect 53475 4340 53675 4425
rect 53825 4465 54025 4540
rect 53825 4425 53905 4465
rect 53945 4425 54025 4465
rect 53825 4340 54025 4425
rect 59775 4465 59975 4540
rect 59775 4425 59855 4465
rect 59895 4425 59975 4465
rect 59775 4340 59975 4425
rect 60125 4465 60325 4540
rect 60125 4425 60205 4465
rect 60245 4425 60325 4465
rect 60125 4340 60325 4425
rect 60475 4465 60675 4540
rect 60475 4425 60555 4465
rect 60595 4425 60675 4465
rect 60475 4340 60675 4425
rect 60825 4465 61025 4540
rect 60825 4425 60905 4465
rect 60945 4425 61025 4465
rect 60825 4340 61025 4425
rect 61175 4465 61375 4540
rect 61175 4425 61255 4465
rect 61295 4425 61375 4465
rect 61175 4340 61375 4425
rect 52425 4115 52625 4190
rect 52425 4075 52505 4115
rect 52545 4075 52625 4115
rect 52425 3990 52625 4075
rect 52775 4115 52975 4190
rect 52775 4075 52855 4115
rect 52895 4075 52975 4115
rect 52775 3990 52975 4075
rect 53125 4115 53325 4190
rect 53125 4075 53205 4115
rect 53245 4075 53325 4115
rect 53125 3990 53325 4075
rect 53475 4115 53675 4190
rect 53475 4075 53555 4115
rect 53595 4075 53675 4115
rect 53475 3990 53675 4075
rect 53825 4115 54025 4190
rect 53825 4075 53905 4115
rect 53945 4075 54025 4115
rect 53825 3990 54025 4075
rect 59775 4115 59975 4190
rect 59775 4075 59855 4115
rect 59895 4075 59975 4115
rect 59775 3990 59975 4075
rect 60125 4115 60325 4190
rect 60125 4075 60205 4115
rect 60245 4075 60325 4115
rect 60125 3990 60325 4075
rect 60475 4115 60675 4190
rect 60475 4075 60555 4115
rect 60595 4075 60675 4115
rect 60475 3990 60675 4075
rect 60825 4115 61025 4190
rect 60825 4075 60905 4115
rect 60945 4075 61025 4115
rect 60825 3990 61025 4075
rect 61175 4115 61375 4190
rect 61175 4075 61255 4115
rect 61295 4075 61375 4115
rect 61175 3990 61375 4075
rect 52425 3765 52625 3840
rect 52425 3725 52505 3765
rect 52545 3725 52625 3765
rect 52425 3640 52625 3725
rect 52775 3765 52975 3840
rect 52775 3725 52855 3765
rect 52895 3725 52975 3765
rect 52775 3640 52975 3725
rect 53125 3765 53325 3840
rect 53125 3725 53205 3765
rect 53245 3725 53325 3765
rect 53125 3640 53325 3725
rect 53475 3765 53675 3840
rect 53475 3725 53555 3765
rect 53595 3725 53675 3765
rect 53475 3640 53675 3725
rect 53825 3765 54025 3840
rect 53825 3725 53905 3765
rect 53945 3725 54025 3765
rect 53825 3640 54025 3725
rect 59775 3765 59975 3840
rect 59775 3725 59855 3765
rect 59895 3725 59975 3765
rect 59775 3640 59975 3725
rect 60125 3765 60325 3840
rect 60125 3725 60205 3765
rect 60245 3725 60325 3765
rect 60125 3640 60325 3725
rect 60475 3765 60675 3840
rect 60475 3725 60555 3765
rect 60595 3725 60675 3765
rect 60475 3640 60675 3725
rect 60825 3765 61025 3840
rect 60825 3725 60905 3765
rect 60945 3725 61025 3765
rect 60825 3640 61025 3725
rect 61175 3765 61375 3840
rect 61175 3725 61255 3765
rect 61295 3725 61375 3765
rect 61175 3640 61375 3725
rect 52425 3415 52625 3490
rect 52425 3375 52505 3415
rect 52545 3375 52625 3415
rect 52425 3290 52625 3375
rect 52775 3415 52975 3490
rect 52775 3375 52855 3415
rect 52895 3375 52975 3415
rect 52775 3290 52975 3375
rect 53125 3415 53325 3490
rect 53125 3375 53205 3415
rect 53245 3375 53325 3415
rect 53125 3290 53325 3375
rect 53475 3415 53675 3490
rect 53475 3375 53555 3415
rect 53595 3375 53675 3415
rect 53475 3290 53675 3375
rect 53825 3415 54025 3490
rect 53825 3375 53905 3415
rect 53945 3375 54025 3415
rect 53825 3290 54025 3375
rect 59775 3415 59975 3490
rect 59775 3375 59855 3415
rect 59895 3375 59975 3415
rect 59775 3290 59975 3375
rect 60125 3415 60325 3490
rect 60125 3375 60205 3415
rect 60245 3375 60325 3415
rect 60125 3290 60325 3375
rect 60475 3415 60675 3490
rect 60475 3375 60555 3415
rect 60595 3375 60675 3415
rect 60475 3290 60675 3375
rect 60825 3415 61025 3490
rect 60825 3375 60905 3415
rect 60945 3375 61025 3415
rect 60825 3290 61025 3375
rect 61175 3415 61375 3490
rect 61175 3375 61255 3415
rect 61295 3375 61375 3415
rect 61175 3290 61375 3375
rect 52425 3065 52625 3140
rect 52425 3025 52505 3065
rect 52545 3025 52625 3065
rect 52425 2940 52625 3025
rect 52775 3065 52975 3140
rect 52775 3025 52855 3065
rect 52895 3025 52975 3065
rect 52775 2940 52975 3025
rect 53125 3065 53325 3140
rect 53125 3025 53205 3065
rect 53245 3025 53325 3065
rect 53125 2940 53325 3025
rect 53475 3065 53675 3140
rect 53475 3025 53555 3065
rect 53595 3025 53675 3065
rect 53475 2940 53675 3025
rect 53825 3065 54025 3140
rect 53825 3025 53905 3065
rect 53945 3025 54025 3065
rect 53825 2940 54025 3025
rect 59775 3065 59975 3140
rect 59775 3025 59855 3065
rect 59895 3025 59975 3065
rect 59775 2940 59975 3025
rect 60125 3065 60325 3140
rect 60125 3025 60205 3065
rect 60245 3025 60325 3065
rect 60125 2940 60325 3025
rect 60475 3065 60675 3140
rect 60475 3025 60555 3065
rect 60595 3025 60675 3065
rect 60475 2940 60675 3025
rect 60825 3065 61025 3140
rect 60825 3025 60905 3065
rect 60945 3025 61025 3065
rect 60825 2940 61025 3025
rect 61175 3065 61375 3140
rect 61175 3025 61255 3065
rect 61295 3025 61375 3065
rect 61175 2940 61375 3025
rect 52425 2715 52625 2790
rect 52425 2675 52505 2715
rect 52545 2675 52625 2715
rect 52425 2590 52625 2675
rect 52775 2715 52975 2790
rect 52775 2675 52855 2715
rect 52895 2675 52975 2715
rect 52775 2590 52975 2675
rect 53125 2715 53325 2790
rect 53125 2675 53205 2715
rect 53245 2675 53325 2715
rect 53125 2590 53325 2675
rect 53475 2715 53675 2790
rect 53475 2675 53555 2715
rect 53595 2675 53675 2715
rect 53475 2590 53675 2675
rect 53825 2715 54025 2790
rect 53825 2675 53905 2715
rect 53945 2675 54025 2715
rect 53825 2590 54025 2675
rect 59775 2715 59975 2790
rect 59775 2675 59855 2715
rect 59895 2675 59975 2715
rect 59775 2590 59975 2675
rect 60125 2715 60325 2790
rect 60125 2675 60205 2715
rect 60245 2675 60325 2715
rect 60125 2590 60325 2675
rect 60475 2715 60675 2790
rect 60475 2675 60555 2715
rect 60595 2675 60675 2715
rect 60475 2590 60675 2675
rect 60825 2715 61025 2790
rect 60825 2675 60905 2715
rect 60945 2675 61025 2715
rect 60825 2590 61025 2675
rect 61175 2715 61375 2790
rect 61175 2675 61255 2715
rect 61295 2675 61375 2715
rect 61175 2590 61375 2675
rect 52425 2365 52625 2440
rect 52425 2325 52505 2365
rect 52545 2325 52625 2365
rect 52425 2240 52625 2325
rect 52775 2365 52975 2440
rect 52775 2325 52855 2365
rect 52895 2325 52975 2365
rect 52775 2240 52975 2325
rect 53125 2365 53325 2440
rect 53125 2325 53205 2365
rect 53245 2325 53325 2365
rect 53125 2240 53325 2325
rect 53475 2365 53675 2440
rect 53475 2325 53555 2365
rect 53595 2325 53675 2365
rect 53475 2240 53675 2325
rect 53825 2365 54025 2440
rect 53825 2325 53905 2365
rect 53945 2325 54025 2365
rect 53825 2240 54025 2325
rect 59775 2365 59975 2440
rect 59775 2325 59855 2365
rect 59895 2325 59975 2365
rect 59775 2240 59975 2325
rect 60125 2365 60325 2440
rect 60125 2325 60205 2365
rect 60245 2325 60325 2365
rect 60125 2240 60325 2325
rect 60475 2365 60675 2440
rect 60475 2325 60555 2365
rect 60595 2325 60675 2365
rect 60475 2240 60675 2325
rect 60825 2365 61025 2440
rect 60825 2325 60905 2365
rect 60945 2325 61025 2365
rect 60825 2240 61025 2325
rect 61175 2365 61375 2440
rect 61175 2325 61255 2365
rect 61295 2325 61375 2365
rect 61175 2240 61375 2325
rect 52425 2015 52625 2090
rect 52425 1975 52505 2015
rect 52545 1975 52625 2015
rect 52425 1890 52625 1975
rect 52775 2015 52975 2090
rect 52775 1975 52855 2015
rect 52895 1975 52975 2015
rect 52775 1890 52975 1975
rect 53125 2015 53325 2090
rect 53125 1975 53205 2015
rect 53245 1975 53325 2015
rect 53125 1890 53325 1975
rect 53475 2015 53675 2090
rect 53475 1975 53555 2015
rect 53595 1975 53675 2015
rect 53475 1890 53675 1975
rect 53825 2015 54025 2090
rect 53825 1975 53905 2015
rect 53945 1975 54025 2015
rect 53825 1890 54025 1975
rect 59775 2015 59975 2090
rect 59775 1975 59855 2015
rect 59895 1975 59975 2015
rect 59775 1890 59975 1975
rect 60125 2015 60325 2090
rect 60125 1975 60205 2015
rect 60245 1975 60325 2015
rect 60125 1890 60325 1975
rect 60475 2015 60675 2090
rect 60475 1975 60555 2015
rect 60595 1975 60675 2015
rect 60475 1890 60675 1975
rect 60825 2015 61025 2090
rect 60825 1975 60905 2015
rect 60945 1975 61025 2015
rect 60825 1890 61025 1975
rect 61175 2015 61375 2090
rect 61175 1975 61255 2015
rect 61295 1975 61375 2015
rect 61175 1890 61375 1975
rect 52425 1665 52625 1740
rect 52425 1625 52505 1665
rect 52545 1625 52625 1665
rect 52425 1540 52625 1625
rect 52775 1665 52975 1740
rect 52775 1625 52855 1665
rect 52895 1625 52975 1665
rect 52775 1540 52975 1625
rect 53125 1665 53325 1740
rect 53125 1625 53205 1665
rect 53245 1625 53325 1665
rect 53125 1540 53325 1625
rect 53475 1665 53675 1740
rect 53475 1625 53555 1665
rect 53595 1625 53675 1665
rect 53475 1540 53675 1625
rect 53825 1665 54025 1740
rect 53825 1625 53905 1665
rect 53945 1625 54025 1665
rect 53825 1540 54025 1625
rect 59775 1665 59975 1740
rect 59775 1625 59855 1665
rect 59895 1625 59975 1665
rect 59775 1540 59975 1625
rect 60125 1665 60325 1740
rect 60125 1625 60205 1665
rect 60245 1625 60325 1665
rect 60125 1540 60325 1625
rect 60475 1665 60675 1740
rect 60475 1625 60555 1665
rect 60595 1625 60675 1665
rect 60475 1540 60675 1625
rect 60825 1665 61025 1740
rect 60825 1625 60905 1665
rect 60945 1625 61025 1665
rect 60825 1540 61025 1625
rect 61175 1665 61375 1740
rect 61175 1625 61255 1665
rect 61295 1625 61375 1665
rect 61175 1540 61375 1625
rect 52425 1315 52625 1390
rect 52425 1275 52505 1315
rect 52545 1275 52625 1315
rect 52425 1190 52625 1275
rect 52775 1315 52975 1390
rect 52775 1275 52855 1315
rect 52895 1275 52975 1315
rect 52775 1190 52975 1275
rect 53125 1315 53325 1390
rect 53125 1275 53205 1315
rect 53245 1275 53325 1315
rect 53125 1190 53325 1275
rect 53475 1315 53675 1390
rect 53475 1275 53555 1315
rect 53595 1275 53675 1315
rect 53475 1190 53675 1275
rect 53825 1315 54025 1390
rect 53825 1275 53905 1315
rect 53945 1275 54025 1315
rect 53825 1190 54025 1275
rect 59775 1315 59975 1390
rect 59775 1275 59855 1315
rect 59895 1275 59975 1315
rect 59775 1190 59975 1275
rect 60125 1315 60325 1390
rect 60125 1275 60205 1315
rect 60245 1275 60325 1315
rect 60125 1190 60325 1275
rect 60475 1315 60675 1390
rect 60475 1275 60555 1315
rect 60595 1275 60675 1315
rect 60475 1190 60675 1275
rect 60825 1315 61025 1390
rect 60825 1275 60905 1315
rect 60945 1275 61025 1315
rect 60825 1190 61025 1275
rect 61175 1315 61375 1390
rect 61175 1275 61255 1315
rect 61295 1275 61375 1315
rect 61175 1190 61375 1275
rect 52425 965 52625 1040
rect 52425 925 52505 965
rect 52545 925 52625 965
rect 52425 840 52625 925
rect 52775 965 52975 1040
rect 52775 925 52855 965
rect 52895 925 52975 965
rect 52775 840 52975 925
rect 53125 965 53325 1040
rect 53125 925 53205 965
rect 53245 925 53325 965
rect 53125 840 53325 925
rect 53475 965 53675 1040
rect 53475 925 53555 965
rect 53595 925 53675 965
rect 53475 840 53675 925
rect 53825 965 54025 1040
rect 53825 925 53905 965
rect 53945 925 54025 965
rect 53825 840 54025 925
rect 59775 965 59975 1040
rect 59775 925 59855 965
rect 59895 925 59975 965
rect 59775 840 59975 925
rect 60125 965 60325 1040
rect 60125 925 60205 965
rect 60245 925 60325 965
rect 60125 840 60325 925
rect 60475 965 60675 1040
rect 60475 925 60555 965
rect 60595 925 60675 965
rect 60475 840 60675 925
rect 60825 965 61025 1040
rect 60825 925 60905 965
rect 60945 925 61025 965
rect 60825 840 61025 925
rect 61175 965 61375 1040
rect 61175 925 61255 965
rect 61295 925 61375 965
rect 61175 840 61375 925
rect 52425 615 52625 690
rect 52425 575 52505 615
rect 52545 575 52625 615
rect 52425 490 52625 575
rect 52775 615 52975 690
rect 52775 575 52855 615
rect 52895 575 52975 615
rect 52775 490 52975 575
rect 53125 615 53325 690
rect 53125 575 53205 615
rect 53245 575 53325 615
rect 53125 490 53325 575
rect 53475 615 53675 690
rect 53475 575 53555 615
rect 53595 575 53675 615
rect 53475 490 53675 575
rect 53825 615 54025 690
rect 53825 575 53905 615
rect 53945 575 54025 615
rect 53825 490 54025 575
rect 59775 615 59975 690
rect 59775 575 59855 615
rect 59895 575 59975 615
rect 59775 490 59975 575
rect 60125 615 60325 690
rect 60125 575 60205 615
rect 60245 575 60325 615
rect 60125 490 60325 575
rect 60475 615 60675 690
rect 60475 575 60555 615
rect 60595 575 60675 615
rect 60475 490 60675 575
rect 60825 615 61025 690
rect 60825 575 60905 615
rect 60945 575 61025 615
rect 60825 490 61025 575
rect 61175 615 61375 690
rect 61175 575 61255 615
rect 61295 575 61375 615
rect 61175 490 61375 575
rect 52425 265 52625 340
rect 52425 225 52505 265
rect 52545 225 52625 265
rect 52425 140 52625 225
rect 52775 265 52975 340
rect 52775 225 52855 265
rect 52895 225 52975 265
rect 52775 140 52975 225
rect 53125 265 53325 340
rect 53125 225 53205 265
rect 53245 225 53325 265
rect 53125 140 53325 225
rect 53475 265 53675 340
rect 53475 225 53555 265
rect 53595 225 53675 265
rect 53475 140 53675 225
rect 53825 265 54025 340
rect 53825 225 53905 265
rect 53945 225 54025 265
rect 53825 140 54025 225
rect 59775 265 59975 340
rect 59775 225 59855 265
rect 59895 225 59975 265
rect 59775 140 59975 225
rect 60125 265 60325 340
rect 60125 225 60205 265
rect 60245 225 60325 265
rect 60125 140 60325 225
rect 60475 265 60675 340
rect 60475 225 60555 265
rect 60595 225 60675 265
rect 60475 140 60675 225
rect 60825 265 61025 340
rect 60825 225 60905 265
rect 60945 225 61025 265
rect 60825 140 61025 225
rect 61175 265 61375 340
rect 61175 225 61255 265
rect 61295 225 61375 265
rect 61175 140 61375 225
rect 52425 -85 52625 -10
rect 52425 -125 52505 -85
rect 52545 -125 52625 -85
rect 52425 -210 52625 -125
rect 52775 -85 52975 -10
rect 52775 -125 52855 -85
rect 52895 -125 52975 -85
rect 52775 -210 52975 -125
rect 53125 -85 53325 -10
rect 53125 -125 53205 -85
rect 53245 -125 53325 -85
rect 53125 -210 53325 -125
rect 53475 -85 53675 -10
rect 53475 -125 53555 -85
rect 53595 -125 53675 -85
rect 53475 -210 53675 -125
rect 53825 -85 54025 -10
rect 53825 -125 53905 -85
rect 53945 -125 54025 -85
rect 53825 -210 54025 -125
rect 54175 -85 54375 -10
rect 54175 -125 54255 -85
rect 54295 -125 54375 -85
rect 54175 -210 54375 -125
rect 54525 -85 54725 -10
rect 54525 -125 54605 -85
rect 54645 -125 54725 -85
rect 54525 -210 54725 -125
rect 54875 -85 55075 -10
rect 54875 -125 54955 -85
rect 54995 -125 55075 -85
rect 54875 -210 55075 -125
rect 55225 -85 55425 -10
rect 55225 -125 55305 -85
rect 55345 -125 55425 -85
rect 55225 -210 55425 -125
rect 55575 -85 55775 -10
rect 55575 -125 55655 -85
rect 55695 -125 55775 -85
rect 55575 -210 55775 -125
rect 55925 -85 56125 -10
rect 55925 -125 56005 -85
rect 56045 -125 56125 -85
rect 55925 -210 56125 -125
rect 56275 -85 56475 -10
rect 56275 -125 56355 -85
rect 56395 -125 56475 -85
rect 56275 -210 56475 -125
rect 56625 -85 56825 -10
rect 56625 -125 56705 -85
rect 56745 -125 56825 -85
rect 56625 -210 56825 -125
rect 56975 -85 57175 -10
rect 56975 -125 57055 -85
rect 57095 -125 57175 -85
rect 56975 -210 57175 -125
rect 57325 -85 57525 -10
rect 57325 -125 57405 -85
rect 57445 -125 57525 -85
rect 57325 -210 57525 -125
rect 57675 -85 57875 -10
rect 57675 -125 57755 -85
rect 57795 -125 57875 -85
rect 57675 -210 57875 -125
rect 58025 -85 58225 -10
rect 58025 -125 58105 -85
rect 58145 -125 58225 -85
rect 58025 -210 58225 -125
rect 58375 -85 58575 -10
rect 58375 -125 58455 -85
rect 58495 -125 58575 -85
rect 58375 -210 58575 -125
rect 58725 -85 58925 -10
rect 58725 -125 58805 -85
rect 58845 -125 58925 -85
rect 58725 -210 58925 -125
rect 59075 -85 59275 -10
rect 59075 -125 59155 -85
rect 59195 -125 59275 -85
rect 59075 -210 59275 -125
rect 59425 -85 59625 -10
rect 59425 -125 59505 -85
rect 59545 -125 59625 -85
rect 59425 -210 59625 -125
rect 59775 -85 59975 -10
rect 59775 -125 59855 -85
rect 59895 -125 59975 -85
rect 59775 -210 59975 -125
rect 60125 -85 60325 -10
rect 60125 -125 60205 -85
rect 60245 -125 60325 -85
rect 60125 -210 60325 -125
rect 60475 -85 60675 -10
rect 60475 -125 60555 -85
rect 60595 -125 60675 -85
rect 60475 -210 60675 -125
rect 60825 -85 61025 -10
rect 60825 -125 60905 -85
rect 60945 -125 61025 -85
rect 60825 -210 61025 -125
rect 61175 -85 61375 -10
rect 61175 -125 61255 -85
rect 61295 -125 61375 -85
rect 61175 -210 61375 -125
rect 52425 -435 52625 -360
rect 52425 -475 52505 -435
rect 52545 -475 52625 -435
rect 52425 -560 52625 -475
rect 52775 -435 52975 -360
rect 52775 -475 52855 -435
rect 52895 -475 52975 -435
rect 52775 -560 52975 -475
rect 53125 -435 53325 -360
rect 53125 -475 53205 -435
rect 53245 -475 53325 -435
rect 53125 -560 53325 -475
rect 53475 -435 53675 -360
rect 53475 -475 53555 -435
rect 53595 -475 53675 -435
rect 53475 -560 53675 -475
rect 53825 -435 54025 -360
rect 53825 -475 53905 -435
rect 53945 -475 54025 -435
rect 53825 -560 54025 -475
rect 54175 -435 54375 -360
rect 54175 -475 54255 -435
rect 54295 -475 54375 -435
rect 54175 -560 54375 -475
rect 54525 -435 54725 -360
rect 54525 -475 54605 -435
rect 54645 -475 54725 -435
rect 54525 -560 54725 -475
rect 54875 -435 55075 -360
rect 54875 -475 54955 -435
rect 54995 -475 55075 -435
rect 54875 -560 55075 -475
rect 55225 -435 55425 -360
rect 55225 -475 55305 -435
rect 55345 -475 55425 -435
rect 55225 -560 55425 -475
rect 55575 -435 55775 -360
rect 55575 -475 55655 -435
rect 55695 -475 55775 -435
rect 55575 -560 55775 -475
rect 55925 -435 56125 -360
rect 55925 -475 56005 -435
rect 56045 -475 56125 -435
rect 55925 -560 56125 -475
rect 56275 -435 56475 -360
rect 56275 -475 56355 -435
rect 56395 -475 56475 -435
rect 56275 -560 56475 -475
rect 56625 -435 56825 -360
rect 56625 -475 56705 -435
rect 56745 -475 56825 -435
rect 56625 -560 56825 -475
rect 56975 -435 57175 -360
rect 56975 -475 57055 -435
rect 57095 -475 57175 -435
rect 56975 -560 57175 -475
rect 57325 -435 57525 -360
rect 57325 -475 57405 -435
rect 57445 -475 57525 -435
rect 57325 -560 57525 -475
rect 57675 -435 57875 -360
rect 57675 -475 57755 -435
rect 57795 -475 57875 -435
rect 57675 -560 57875 -475
rect 58025 -435 58225 -360
rect 58025 -475 58105 -435
rect 58145 -475 58225 -435
rect 58025 -560 58225 -475
rect 58375 -435 58575 -360
rect 58375 -475 58455 -435
rect 58495 -475 58575 -435
rect 58375 -560 58575 -475
rect 58725 -435 58925 -360
rect 58725 -475 58805 -435
rect 58845 -475 58925 -435
rect 58725 -560 58925 -475
rect 59075 -435 59275 -360
rect 59075 -475 59155 -435
rect 59195 -475 59275 -435
rect 59075 -560 59275 -475
rect 59425 -435 59625 -360
rect 59425 -475 59505 -435
rect 59545 -475 59625 -435
rect 59425 -560 59625 -475
rect 59775 -435 59975 -360
rect 59775 -475 59855 -435
rect 59895 -475 59975 -435
rect 59775 -560 59975 -475
rect 60125 -435 60325 -360
rect 60125 -475 60205 -435
rect 60245 -475 60325 -435
rect 60125 -560 60325 -475
rect 60475 -435 60675 -360
rect 60475 -475 60555 -435
rect 60595 -475 60675 -435
rect 60475 -560 60675 -475
rect 60825 -435 61025 -360
rect 60825 -475 60905 -435
rect 60945 -475 61025 -435
rect 60825 -560 61025 -475
rect 61175 -435 61375 -360
rect 61175 -475 61255 -435
rect 61295 -475 61375 -435
rect 61175 -560 61375 -475
<< mimcapcontact >>
rect 52505 5825 52545 5865
rect 52855 5825 52895 5865
rect 53205 5825 53245 5865
rect 53555 5825 53595 5865
rect 53905 5825 53945 5865
rect 54255 5825 54295 5865
rect 54605 5825 54645 5865
rect 54955 5825 54995 5865
rect 55305 5825 55345 5865
rect 55655 5825 55695 5865
rect 56005 5825 56045 5865
rect 56355 5825 56395 5865
rect 56705 5825 56745 5865
rect 57055 5825 57095 5865
rect 57405 5825 57445 5865
rect 57755 5825 57795 5865
rect 58105 5825 58145 5865
rect 58455 5825 58495 5865
rect 58805 5825 58845 5865
rect 59155 5825 59195 5865
rect 59505 5825 59545 5865
rect 59855 5825 59895 5865
rect 60205 5825 60245 5865
rect 60555 5825 60595 5865
rect 60905 5825 60945 5865
rect 61255 5825 61295 5865
rect 52505 5475 52545 5515
rect 52855 5475 52895 5515
rect 53205 5475 53245 5515
rect 53555 5475 53595 5515
rect 53905 5475 53945 5515
rect 54255 5475 54295 5515
rect 54605 5475 54645 5515
rect 54955 5475 54995 5515
rect 55305 5475 55345 5515
rect 55655 5475 55695 5515
rect 56005 5475 56045 5515
rect 56355 5475 56395 5515
rect 56705 5475 56745 5515
rect 57055 5475 57095 5515
rect 57405 5475 57445 5515
rect 57755 5475 57795 5515
rect 58105 5475 58145 5515
rect 58455 5475 58495 5515
rect 58805 5475 58845 5515
rect 59155 5475 59195 5515
rect 59505 5475 59545 5515
rect 59855 5475 59895 5515
rect 60205 5475 60245 5515
rect 60555 5475 60595 5515
rect 60905 5475 60945 5515
rect 61255 5475 61295 5515
rect 52505 5125 52545 5165
rect 52855 5125 52895 5165
rect 53205 5125 53245 5165
rect 53555 5125 53595 5165
rect 53905 5125 53945 5165
rect 54255 5125 54295 5165
rect 54605 5125 54645 5165
rect 54955 5125 54995 5165
rect 55305 5125 55345 5165
rect 55655 5115 55695 5155
rect 56005 5115 56045 5155
rect 56355 5115 56395 5155
rect 56705 5115 56745 5155
rect 57055 5115 57095 5155
rect 57405 5115 57445 5155
rect 57755 5115 57795 5155
rect 58105 5115 58145 5155
rect 58455 5125 58495 5165
rect 58805 5125 58845 5165
rect 59155 5125 59195 5165
rect 59505 5125 59545 5165
rect 59855 5125 59895 5165
rect 60205 5125 60245 5165
rect 60555 5125 60595 5165
rect 60905 5125 60945 5165
rect 61255 5125 61295 5165
rect 52505 4775 52545 4815
rect 52855 4775 52895 4815
rect 53205 4775 53245 4815
rect 53555 4775 53595 4815
rect 53905 4775 53945 4815
rect 54255 4775 54295 4815
rect 54605 4775 54645 4815
rect 54955 4775 54995 4815
rect 55305 4775 55345 4815
rect 55655 4775 55695 4815
rect 58105 4765 58145 4805
rect 58455 4775 58495 4815
rect 58805 4775 58845 4815
rect 59155 4775 59195 4815
rect 59505 4775 59545 4815
rect 59855 4775 59895 4815
rect 60205 4775 60245 4815
rect 60555 4775 60595 4815
rect 60905 4775 60945 4815
rect 61255 4775 61295 4815
rect 52505 4425 52545 4465
rect 52855 4425 52895 4465
rect 53205 4425 53245 4465
rect 53555 4425 53595 4465
rect 53905 4425 53945 4465
rect 59855 4425 59895 4465
rect 60205 4425 60245 4465
rect 60555 4425 60595 4465
rect 60905 4425 60945 4465
rect 61255 4425 61295 4465
rect 52505 4075 52545 4115
rect 52855 4075 52895 4115
rect 53205 4075 53245 4115
rect 53555 4075 53595 4115
rect 53905 4075 53945 4115
rect 59855 4075 59895 4115
rect 60205 4075 60245 4115
rect 60555 4075 60595 4115
rect 60905 4075 60945 4115
rect 61255 4075 61295 4115
rect 52505 3725 52545 3765
rect 52855 3725 52895 3765
rect 53205 3725 53245 3765
rect 53555 3725 53595 3765
rect 53905 3725 53945 3765
rect 59855 3725 59895 3765
rect 60205 3725 60245 3765
rect 60555 3725 60595 3765
rect 60905 3725 60945 3765
rect 61255 3725 61295 3765
rect 52505 3375 52545 3415
rect 52855 3375 52895 3415
rect 53205 3375 53245 3415
rect 53555 3375 53595 3415
rect 53905 3375 53945 3415
rect 59855 3375 59895 3415
rect 60205 3375 60245 3415
rect 60555 3375 60595 3415
rect 60905 3375 60945 3415
rect 61255 3375 61295 3415
rect 52505 3025 52545 3065
rect 52855 3025 52895 3065
rect 53205 3025 53245 3065
rect 53555 3025 53595 3065
rect 53905 3025 53945 3065
rect 59855 3025 59895 3065
rect 60205 3025 60245 3065
rect 60555 3025 60595 3065
rect 60905 3025 60945 3065
rect 61255 3025 61295 3065
rect 52505 2675 52545 2715
rect 52855 2675 52895 2715
rect 53205 2675 53245 2715
rect 53555 2675 53595 2715
rect 53905 2675 53945 2715
rect 59855 2675 59895 2715
rect 60205 2675 60245 2715
rect 60555 2675 60595 2715
rect 60905 2675 60945 2715
rect 61255 2675 61295 2715
rect 52505 2325 52545 2365
rect 52855 2325 52895 2365
rect 53205 2325 53245 2365
rect 53555 2325 53595 2365
rect 53905 2325 53945 2365
rect 59855 2325 59895 2365
rect 60205 2325 60245 2365
rect 60555 2325 60595 2365
rect 60905 2325 60945 2365
rect 61255 2325 61295 2365
rect 52505 1975 52545 2015
rect 52855 1975 52895 2015
rect 53205 1975 53245 2015
rect 53555 1975 53595 2015
rect 53905 1975 53945 2015
rect 59855 1975 59895 2015
rect 60205 1975 60245 2015
rect 60555 1975 60595 2015
rect 60905 1975 60945 2015
rect 61255 1975 61295 2015
rect 52505 1625 52545 1665
rect 52855 1625 52895 1665
rect 53205 1625 53245 1665
rect 53555 1625 53595 1665
rect 53905 1625 53945 1665
rect 59855 1625 59895 1665
rect 60205 1625 60245 1665
rect 60555 1625 60595 1665
rect 60905 1625 60945 1665
rect 61255 1625 61295 1665
rect 52505 1275 52545 1315
rect 52855 1275 52895 1315
rect 53205 1275 53245 1315
rect 53555 1275 53595 1315
rect 53905 1275 53945 1315
rect 59855 1275 59895 1315
rect 60205 1275 60245 1315
rect 60555 1275 60595 1315
rect 60905 1275 60945 1315
rect 61255 1275 61295 1315
rect 52505 925 52545 965
rect 52855 925 52895 965
rect 53205 925 53245 965
rect 53555 925 53595 965
rect 53905 925 53945 965
rect 59855 925 59895 965
rect 60205 925 60245 965
rect 60555 925 60595 965
rect 60905 925 60945 965
rect 61255 925 61295 965
rect 52505 575 52545 615
rect 52855 575 52895 615
rect 53205 575 53245 615
rect 53555 575 53595 615
rect 53905 575 53945 615
rect 59855 575 59895 615
rect 60205 575 60245 615
rect 60555 575 60595 615
rect 60905 575 60945 615
rect 61255 575 61295 615
rect 52505 225 52545 265
rect 52855 225 52895 265
rect 53205 225 53245 265
rect 53555 225 53595 265
rect 53905 225 53945 265
rect 59855 225 59895 265
rect 60205 225 60245 265
rect 60555 225 60595 265
rect 60905 225 60945 265
rect 61255 225 61295 265
rect 52505 -125 52545 -85
rect 52855 -125 52895 -85
rect 53205 -125 53245 -85
rect 53555 -125 53595 -85
rect 53905 -125 53945 -85
rect 54255 -125 54295 -85
rect 54605 -125 54645 -85
rect 54955 -125 54995 -85
rect 55305 -125 55345 -85
rect 55655 -125 55695 -85
rect 56005 -125 56045 -85
rect 56355 -125 56395 -85
rect 56705 -125 56745 -85
rect 57055 -125 57095 -85
rect 57405 -125 57445 -85
rect 57755 -125 57795 -85
rect 58105 -125 58145 -85
rect 58455 -125 58495 -85
rect 58805 -125 58845 -85
rect 59155 -125 59195 -85
rect 59505 -125 59545 -85
rect 59855 -125 59895 -85
rect 60205 -125 60245 -85
rect 60555 -125 60595 -85
rect 60905 -125 60945 -85
rect 61255 -125 61295 -85
rect 52505 -475 52545 -435
rect 52855 -475 52895 -435
rect 53205 -475 53245 -435
rect 53555 -475 53595 -435
rect 53905 -475 53945 -435
rect 54255 -475 54295 -435
rect 54605 -475 54645 -435
rect 54955 -475 54995 -435
rect 55305 -475 55345 -435
rect 55655 -475 55695 -435
rect 56005 -475 56045 -435
rect 56355 -475 56395 -435
rect 56705 -475 56745 -435
rect 57055 -475 57095 -435
rect 57405 -475 57445 -435
rect 57755 -475 57795 -435
rect 58105 -475 58145 -435
rect 58455 -475 58495 -435
rect 58805 -475 58845 -435
rect 59155 -475 59195 -435
rect 59505 -475 59545 -435
rect 59855 -475 59895 -435
rect 60205 -475 60245 -435
rect 60555 -475 60595 -435
rect 60905 -475 60945 -435
rect 61255 -475 61295 -435
<< metal4 >>
rect 52500 5865 53250 5870
rect 52500 5825 52505 5865
rect 52545 5825 52855 5865
rect 52895 5825 53205 5865
rect 53245 5825 53250 5865
rect 52500 5820 53250 5825
rect 53200 5520 53250 5820
rect 53550 5865 53600 5870
rect 53550 5825 53555 5865
rect 53595 5825 53600 5865
rect 53550 5520 53600 5825
rect 53900 5865 53950 5870
rect 53900 5825 53905 5865
rect 53945 5825 53950 5865
rect 53900 5520 53950 5825
rect 54250 5865 54300 5870
rect 54250 5825 54255 5865
rect 54295 5825 54300 5865
rect 54250 5520 54300 5825
rect 54600 5865 54650 5870
rect 54600 5825 54605 5865
rect 54645 5825 54650 5865
rect 54600 5520 54650 5825
rect 54950 5865 55000 5870
rect 54950 5825 54955 5865
rect 54995 5825 55000 5865
rect 54950 5520 55000 5825
rect 55300 5865 55350 5870
rect 55300 5825 55305 5865
rect 55345 5825 55350 5865
rect 55300 5520 55350 5825
rect 55650 5865 55700 5870
rect 55650 5825 55655 5865
rect 55695 5825 55700 5865
rect 55650 5520 55700 5825
rect 56000 5865 56050 5870
rect 56000 5825 56005 5865
rect 56045 5825 56050 5865
rect 56000 5520 56050 5825
rect 56350 5865 56400 5870
rect 56350 5825 56355 5865
rect 56395 5825 56400 5865
rect 56350 5520 56400 5825
rect 56700 5865 56750 5870
rect 56700 5825 56705 5865
rect 56745 5825 56750 5865
rect 56700 5520 56750 5825
rect 52500 5515 56750 5520
rect 52500 5475 52505 5515
rect 52545 5475 52855 5515
rect 52895 5475 53205 5515
rect 53245 5475 53555 5515
rect 53595 5475 53905 5515
rect 53945 5475 54255 5515
rect 54295 5475 54605 5515
rect 54645 5475 54955 5515
rect 54995 5475 55305 5515
rect 55345 5475 55655 5515
rect 55695 5475 56005 5515
rect 56045 5475 56355 5515
rect 56395 5475 56705 5515
rect 56745 5475 56750 5515
rect 52500 5470 56750 5475
rect 53200 5170 53250 5470
rect 52500 5165 53950 5170
rect 52500 5125 52505 5165
rect 52545 5125 52855 5165
rect 52895 5125 53205 5165
rect 53245 5125 53555 5165
rect 53595 5125 53905 5165
rect 53945 5125 53950 5165
rect 52500 5120 53950 5125
rect 54250 5165 54300 5470
rect 54250 5125 54255 5165
rect 54295 5125 54300 5165
rect 53200 4820 53250 5120
rect 52500 4815 53950 4820
rect 52500 4775 52505 4815
rect 52545 4775 52855 4815
rect 52895 4775 53205 4815
rect 53245 4775 53555 4815
rect 53595 4775 53905 4815
rect 53945 4775 53950 4815
rect 52500 4770 53950 4775
rect 54250 4815 54300 5125
rect 54250 4775 54255 4815
rect 54295 4775 54300 4815
rect 54250 4770 54300 4775
rect 54600 5165 54650 5470
rect 54600 5125 54605 5165
rect 54645 5125 54650 5165
rect 54600 4815 54650 5125
rect 54600 4775 54605 4815
rect 54645 4775 54650 4815
rect 54600 4770 54650 4775
rect 54950 5165 55000 5470
rect 54950 5125 54955 5165
rect 54995 5125 55000 5165
rect 54950 4815 55000 5125
rect 54950 4775 54955 4815
rect 54995 4775 55000 4815
rect 54950 4770 55000 4775
rect 55300 5165 55350 5470
rect 55300 5125 55305 5165
rect 55345 5125 55350 5165
rect 55300 4815 55350 5125
rect 55300 4775 55305 4815
rect 55345 4775 55350 4815
rect 55300 4770 55350 4775
rect 55650 5155 55700 5470
rect 55650 5115 55655 5155
rect 55695 5115 55700 5155
rect 55650 4815 55700 5115
rect 56000 5155 56050 5470
rect 56000 5115 56005 5155
rect 56045 5115 56050 5155
rect 56000 5110 56050 5115
rect 56350 5155 56400 5470
rect 56350 5115 56355 5155
rect 56395 5115 56400 5155
rect 56350 5110 56400 5115
rect 56700 5155 56750 5470
rect 56700 5115 56705 5155
rect 56745 5115 56750 5155
rect 56700 5110 56750 5115
rect 57050 5865 57100 5870
rect 57050 5825 57055 5865
rect 57095 5825 57100 5865
rect 57050 5520 57100 5825
rect 57400 5865 57450 5870
rect 57400 5825 57405 5865
rect 57445 5825 57450 5865
rect 57400 5520 57450 5825
rect 57750 5865 57800 5870
rect 57750 5825 57755 5865
rect 57795 5825 57800 5865
rect 57750 5520 57800 5825
rect 58100 5865 58150 5870
rect 58100 5825 58105 5865
rect 58145 5825 58150 5865
rect 58100 5520 58150 5825
rect 58450 5865 58500 5870
rect 58450 5825 58455 5865
rect 58495 5825 58500 5865
rect 58450 5520 58500 5825
rect 58800 5865 58850 5870
rect 58800 5825 58805 5865
rect 58845 5825 58850 5865
rect 58800 5520 58850 5825
rect 59150 5865 59200 5870
rect 59150 5825 59155 5865
rect 59195 5825 59200 5865
rect 59150 5520 59200 5825
rect 59500 5865 59550 5870
rect 59500 5825 59505 5865
rect 59545 5825 59550 5865
rect 59500 5520 59550 5825
rect 59850 5865 59900 5870
rect 59850 5825 59855 5865
rect 59895 5825 59900 5865
rect 59850 5520 59900 5825
rect 60200 5865 60250 5870
rect 60200 5825 60205 5865
rect 60245 5825 60250 5865
rect 60200 5520 60250 5825
rect 60550 5865 61300 5870
rect 60550 5825 60555 5865
rect 60595 5825 60905 5865
rect 60945 5825 61255 5865
rect 61295 5825 61300 5865
rect 60550 5820 61300 5825
rect 60550 5520 60600 5820
rect 57050 5515 61300 5520
rect 57050 5475 57055 5515
rect 57095 5475 57405 5515
rect 57445 5475 57755 5515
rect 57795 5475 58105 5515
rect 58145 5475 58455 5515
rect 58495 5475 58805 5515
rect 58845 5475 59155 5515
rect 59195 5475 59505 5515
rect 59545 5475 59855 5515
rect 59895 5475 60205 5515
rect 60245 5475 60555 5515
rect 60595 5475 60905 5515
rect 60945 5475 61255 5515
rect 61295 5475 61300 5515
rect 57050 5470 61300 5475
rect 57050 5155 57100 5470
rect 57050 5115 57055 5155
rect 57095 5115 57100 5155
rect 57050 5110 57100 5115
rect 57400 5155 57450 5470
rect 57400 5115 57405 5155
rect 57445 5115 57450 5155
rect 57400 5110 57450 5115
rect 57750 5155 57800 5470
rect 57750 5115 57755 5155
rect 57795 5115 57800 5155
rect 57750 5110 57800 5115
rect 58100 5155 58150 5470
rect 58100 5115 58105 5155
rect 58145 5115 58150 5155
rect 55650 4775 55655 4815
rect 55695 4775 55700 4815
rect 55650 4770 55700 4775
rect 58100 4805 58150 5115
rect 53200 4470 53250 4770
rect 58100 4765 58105 4805
rect 58145 4765 58150 4805
rect 58450 5165 58500 5470
rect 58450 5125 58455 5165
rect 58495 5125 58500 5165
rect 58450 4815 58500 5125
rect 58450 4775 58455 4815
rect 58495 4775 58500 4815
rect 58450 4770 58500 4775
rect 58800 5165 58850 5470
rect 58800 5125 58805 5165
rect 58845 5125 58850 5165
rect 58800 4815 58850 5125
rect 58800 4775 58805 4815
rect 58845 4775 58850 4815
rect 58800 4770 58850 4775
rect 59150 5165 59200 5470
rect 59150 5125 59155 5165
rect 59195 5125 59200 5165
rect 59150 4815 59200 5125
rect 59150 4775 59155 4815
rect 59195 4775 59200 4815
rect 59150 4770 59200 4775
rect 59500 5165 59550 5470
rect 60550 5170 60600 5470
rect 59500 5125 59505 5165
rect 59545 5125 59550 5165
rect 59500 4815 59550 5125
rect 59850 5165 61300 5170
rect 59850 5125 59855 5165
rect 59895 5125 60205 5165
rect 60245 5125 60555 5165
rect 60595 5125 60905 5165
rect 60945 5125 61255 5165
rect 61295 5125 61300 5165
rect 59850 5120 61300 5125
rect 60550 4820 60600 5120
rect 59500 4775 59505 4815
rect 59545 4775 59550 4815
rect 59500 4770 59550 4775
rect 59850 4815 61300 4820
rect 59850 4775 59855 4815
rect 59895 4775 60205 4815
rect 60245 4775 60555 4815
rect 60595 4775 60905 4815
rect 60945 4775 61255 4815
rect 61295 4775 61300 4815
rect 59850 4770 61300 4775
rect 58100 4760 58150 4765
rect 60550 4470 60600 4770
rect 52500 4465 53950 4470
rect 52500 4425 52505 4465
rect 52545 4425 52855 4465
rect 52895 4425 53205 4465
rect 53245 4425 53555 4465
rect 53595 4425 53905 4465
rect 53945 4425 53950 4465
rect 52500 4420 53950 4425
rect 59850 4465 61300 4470
rect 59850 4425 59855 4465
rect 59895 4425 60205 4465
rect 60245 4425 60555 4465
rect 60595 4425 60905 4465
rect 60945 4425 61255 4465
rect 61295 4425 61300 4465
rect 59850 4420 61300 4425
rect 53200 4120 53250 4420
rect 60550 4120 60600 4420
rect 52500 4115 53950 4120
rect 52500 4075 52505 4115
rect 52545 4075 52855 4115
rect 52895 4075 53205 4115
rect 53245 4075 53555 4115
rect 53595 4075 53905 4115
rect 53945 4075 53950 4115
rect 52500 4070 53950 4075
rect 59850 4115 61300 4120
rect 59850 4075 59855 4115
rect 59895 4075 60205 4115
rect 60245 4075 60555 4115
rect 60595 4075 60905 4115
rect 60945 4075 61255 4115
rect 61295 4075 61300 4115
rect 59850 4070 61300 4075
rect 53200 3770 53250 4070
rect 60550 3770 60600 4070
rect 52500 3765 53950 3770
rect 52500 3725 52505 3765
rect 52545 3725 52855 3765
rect 52895 3725 53205 3765
rect 53245 3725 53555 3765
rect 53595 3725 53905 3765
rect 53945 3725 53950 3765
rect 52500 3720 53950 3725
rect 59850 3765 61300 3770
rect 59850 3725 59855 3765
rect 59895 3725 60205 3765
rect 60245 3725 60555 3765
rect 60595 3725 60905 3765
rect 60945 3725 61255 3765
rect 61295 3725 61300 3765
rect 59850 3720 61300 3725
rect 53200 3420 53250 3720
rect 60550 3420 60600 3720
rect 52500 3415 53950 3420
rect 52500 3375 52505 3415
rect 52545 3375 52855 3415
rect 52895 3375 53205 3415
rect 53245 3375 53555 3415
rect 53595 3375 53905 3415
rect 53945 3375 53950 3415
rect 52500 3370 53950 3375
rect 59850 3415 61300 3420
rect 59850 3375 59855 3415
rect 59895 3375 60205 3415
rect 60245 3375 60555 3415
rect 60595 3375 60905 3415
rect 60945 3375 61255 3415
rect 61295 3375 61300 3415
rect 59850 3370 61300 3375
rect 53200 3070 53250 3370
rect 60550 3070 60600 3370
rect 52500 3065 53950 3070
rect 52500 3025 52505 3065
rect 52545 3025 52855 3065
rect 52895 3025 53205 3065
rect 53245 3025 53555 3065
rect 53595 3025 53905 3065
rect 53945 3025 53950 3065
rect 52500 3020 53950 3025
rect 59850 3065 61300 3070
rect 59850 3025 59855 3065
rect 59895 3025 60205 3065
rect 60245 3025 60555 3065
rect 60595 3025 60905 3065
rect 60945 3025 61255 3065
rect 61295 3025 61300 3065
rect 59850 3020 61300 3025
rect 53200 2720 53250 3020
rect 60550 2720 60600 3020
rect 52500 2715 53950 2720
rect 52500 2675 52505 2715
rect 52545 2675 52855 2715
rect 52895 2675 53205 2715
rect 53245 2675 53555 2715
rect 53595 2675 53905 2715
rect 53945 2675 53950 2715
rect 52500 2670 53950 2675
rect 59850 2715 61300 2720
rect 59850 2675 59855 2715
rect 59895 2675 60205 2715
rect 60245 2675 60555 2715
rect 60595 2675 60905 2715
rect 60945 2675 61255 2715
rect 61295 2675 61300 2715
rect 59850 2670 61300 2675
rect 53200 2370 53250 2670
rect 60550 2370 60600 2670
rect 52500 2365 53950 2370
rect 52500 2325 52505 2365
rect 52545 2325 52855 2365
rect 52895 2325 53205 2365
rect 53245 2325 53555 2365
rect 53595 2325 53905 2365
rect 53945 2325 53950 2365
rect 52500 2320 53950 2325
rect 59850 2365 61300 2370
rect 59850 2325 59855 2365
rect 59895 2325 60205 2365
rect 60245 2325 60555 2365
rect 60595 2325 60905 2365
rect 60945 2325 61255 2365
rect 61295 2325 61300 2365
rect 59850 2320 61300 2325
rect 53200 2020 53250 2320
rect 60550 2020 60600 2320
rect 52500 2015 53950 2020
rect 52500 1975 52505 2015
rect 52545 1975 52855 2015
rect 52895 1975 53205 2015
rect 53245 1975 53555 2015
rect 53595 1975 53905 2015
rect 53945 1975 53950 2015
rect 52500 1970 53950 1975
rect 59850 2015 61300 2020
rect 59850 1975 59855 2015
rect 59895 1975 60205 2015
rect 60245 1975 60555 2015
rect 60595 1975 60905 2015
rect 60945 1975 61255 2015
rect 61295 1975 61300 2015
rect 59850 1970 61300 1975
rect 53200 1670 53250 1970
rect 53900 1715 54435 1720
rect 53900 1675 54190 1715
rect 54230 1675 54240 1715
rect 54280 1675 54290 1715
rect 54330 1675 54340 1715
rect 54380 1675 54390 1715
rect 54430 1675 54435 1715
rect 53900 1670 54435 1675
rect 52500 1665 54435 1670
rect 52500 1625 52505 1665
rect 52545 1625 52855 1665
rect 52895 1625 53205 1665
rect 53245 1625 53555 1665
rect 53595 1625 53905 1665
rect 53945 1625 54190 1665
rect 54230 1625 54240 1665
rect 54280 1625 54290 1665
rect 54330 1625 54340 1665
rect 54380 1625 54390 1665
rect 54430 1625 54435 1665
rect 52500 1620 54435 1625
rect 53200 1320 53250 1620
rect 53900 1615 54435 1620
rect 53900 1575 54190 1615
rect 54230 1575 54240 1615
rect 54280 1575 54290 1615
rect 54330 1575 54340 1615
rect 54380 1575 54390 1615
rect 54430 1575 54435 1615
rect 53900 1570 54435 1575
rect 59365 1715 59905 1720
rect 59365 1675 59370 1715
rect 59410 1675 59420 1715
rect 59460 1675 59470 1715
rect 59510 1675 59520 1715
rect 59560 1675 59570 1715
rect 59610 1675 59905 1715
rect 59365 1670 59905 1675
rect 60550 1670 60600 1970
rect 59365 1665 61300 1670
rect 59365 1625 59370 1665
rect 59410 1625 59420 1665
rect 59460 1625 59470 1665
rect 59510 1625 59520 1665
rect 59560 1625 59570 1665
rect 59610 1625 59855 1665
rect 59895 1625 60205 1665
rect 60245 1625 60555 1665
rect 60595 1625 60905 1665
rect 60945 1625 61255 1665
rect 61295 1625 61300 1665
rect 59365 1620 61300 1625
rect 59365 1615 59905 1620
rect 59365 1575 59370 1615
rect 59410 1575 59420 1615
rect 59460 1575 59470 1615
rect 59510 1575 59520 1615
rect 59560 1575 59570 1615
rect 59610 1575 59905 1615
rect 59365 1570 59905 1575
rect 60550 1320 60600 1620
rect 52500 1315 53950 1320
rect 52500 1275 52505 1315
rect 52545 1275 52855 1315
rect 52895 1275 53205 1315
rect 53245 1275 53555 1315
rect 53595 1275 53905 1315
rect 53945 1275 53950 1315
rect 52500 1270 53950 1275
rect 59850 1315 61300 1320
rect 59850 1275 59855 1315
rect 59895 1275 60205 1315
rect 60245 1275 60555 1315
rect 60595 1275 60905 1315
rect 60945 1275 61255 1315
rect 61295 1275 61300 1315
rect 59850 1270 61300 1275
rect 53200 970 53250 1270
rect 60550 970 60600 1270
rect 52500 965 53950 970
rect 52500 925 52505 965
rect 52545 925 52855 965
rect 52895 925 53205 965
rect 53245 925 53555 965
rect 53595 925 53905 965
rect 53945 925 53950 965
rect 52500 920 53950 925
rect 59850 965 61300 970
rect 59850 925 59855 965
rect 59895 925 60205 965
rect 60245 925 60555 965
rect 60595 925 60905 965
rect 60945 925 61255 965
rect 61295 925 61300 965
rect 59850 920 61300 925
rect 53200 620 53250 920
rect 60550 620 60600 920
rect 52500 615 53950 620
rect 52500 575 52505 615
rect 52545 575 52855 615
rect 52895 575 53205 615
rect 53245 575 53555 615
rect 53595 575 53905 615
rect 53945 575 53950 615
rect 52500 570 53950 575
rect 59850 615 61300 620
rect 59850 575 59855 615
rect 59895 575 60205 615
rect 60245 575 60555 615
rect 60595 575 60905 615
rect 60945 575 61255 615
rect 61295 575 61300 615
rect 59850 570 61300 575
rect 53200 270 53250 570
rect 60550 270 60600 570
rect 52500 265 53950 270
rect 52500 225 52505 265
rect 52545 225 52855 265
rect 52895 225 53205 265
rect 53245 225 53555 265
rect 53595 225 53905 265
rect 53945 225 53950 265
rect 52500 220 53950 225
rect 59850 265 61300 270
rect 59850 225 59855 265
rect 59895 225 60205 265
rect 60245 225 60555 265
rect 60595 225 60905 265
rect 60945 225 61255 265
rect 61295 225 61300 265
rect 59850 220 61300 225
rect 53200 -80 53250 220
rect 60550 -80 60600 220
rect 52500 -85 56750 -80
rect 52500 -125 52505 -85
rect 52545 -125 52855 -85
rect 52895 -125 53205 -85
rect 53245 -125 53555 -85
rect 53595 -125 53905 -85
rect 53945 -125 54255 -85
rect 54295 -125 54605 -85
rect 54645 -125 54955 -85
rect 54995 -125 55305 -85
rect 55345 -125 55655 -85
rect 55695 -125 56005 -85
rect 56045 -125 56355 -85
rect 56395 -125 56705 -85
rect 56745 -125 56750 -85
rect 52500 -130 56750 -125
rect 53200 -430 53250 -130
rect 52500 -435 53250 -430
rect 52500 -475 52505 -435
rect 52545 -475 52855 -435
rect 52895 -475 53205 -435
rect 53245 -475 53250 -435
rect 52500 -480 53250 -475
rect 53550 -435 53600 -130
rect 53550 -475 53555 -435
rect 53595 -475 53600 -435
rect 53550 -480 53600 -475
rect 53900 -435 53950 -130
rect 53900 -475 53905 -435
rect 53945 -475 53950 -435
rect 53900 -480 53950 -475
rect 54250 -435 54300 -130
rect 54250 -475 54255 -435
rect 54295 -475 54300 -435
rect 54250 -480 54300 -475
rect 54600 -435 54650 -130
rect 54600 -475 54605 -435
rect 54645 -475 54650 -435
rect 54600 -480 54650 -475
rect 54950 -435 55000 -130
rect 54950 -475 54955 -435
rect 54995 -475 55000 -435
rect 54950 -480 55000 -475
rect 55300 -435 55350 -130
rect 55300 -475 55305 -435
rect 55345 -475 55350 -435
rect 55300 -480 55350 -475
rect 55650 -435 55700 -130
rect 55650 -475 55655 -435
rect 55695 -475 55700 -435
rect 55650 -480 55700 -475
rect 56000 -435 56050 -130
rect 56000 -475 56005 -435
rect 56045 -475 56050 -435
rect 56000 -480 56050 -475
rect 56350 -435 56400 -130
rect 56350 -475 56355 -435
rect 56395 -475 56400 -435
rect 56350 -480 56400 -475
rect 56700 -435 56750 -130
rect 56700 -475 56705 -435
rect 56745 -475 56750 -435
rect 56700 -480 56750 -475
rect 57050 -85 61300 -80
rect 57050 -125 57055 -85
rect 57095 -125 57405 -85
rect 57445 -125 57755 -85
rect 57795 -125 58105 -85
rect 58145 -125 58455 -85
rect 58495 -125 58805 -85
rect 58845 -125 59155 -85
rect 59195 -125 59505 -85
rect 59545 -125 59855 -85
rect 59895 -125 60205 -85
rect 60245 -125 60555 -85
rect 60595 -125 60905 -85
rect 60945 -125 61255 -85
rect 61295 -125 61300 -85
rect 57050 -130 61300 -125
rect 57050 -435 57100 -130
rect 57050 -475 57055 -435
rect 57095 -475 57100 -435
rect 57050 -480 57100 -475
rect 57400 -435 57450 -130
rect 57400 -475 57405 -435
rect 57445 -475 57450 -435
rect 57400 -480 57450 -475
rect 57750 -435 57800 -130
rect 57750 -475 57755 -435
rect 57795 -475 57800 -435
rect 57750 -480 57800 -475
rect 58100 -435 58150 -130
rect 58100 -475 58105 -435
rect 58145 -475 58150 -435
rect 58100 -480 58150 -475
rect 58450 -435 58500 -130
rect 58450 -475 58455 -435
rect 58495 -475 58500 -435
rect 58450 -480 58500 -475
rect 58800 -435 58850 -130
rect 58800 -475 58805 -435
rect 58845 -475 58850 -435
rect 58800 -480 58850 -475
rect 59150 -435 59200 -130
rect 59150 -475 59155 -435
rect 59195 -475 59200 -435
rect 59150 -480 59200 -475
rect 59500 -435 59550 -130
rect 59500 -475 59505 -435
rect 59545 -475 59550 -435
rect 59500 -480 59550 -475
rect 59850 -435 59900 -130
rect 59850 -475 59855 -435
rect 59895 -475 59900 -435
rect 59850 -480 59900 -475
rect 60200 -435 60250 -130
rect 60200 -475 60205 -435
rect 60245 -475 60250 -435
rect 60200 -480 60250 -475
rect 60550 -430 60600 -130
rect 60550 -435 61300 -430
rect 60550 -475 60555 -435
rect 60595 -475 60905 -435
rect 60945 -475 61255 -435
rect 61295 -475 61300 -435
rect 60550 -480 61300 -475
<< labels >>
flabel metal3 59195 3460 59195 3460 3 FreeSans 240 0 80 0 cap_res_X
flabel metal3 54605 3460 54605 3460 7 FreeSans 240 0 -80 0 cap_res_Y
flabel metal1 56370 1880 56370 1880 7 FreeSans 240 0 -80 0 VD2
flabel metal1 57430 1875 57430 1875 3 FreeSans 240 0 80 0 VD1
flabel metal1 56950 1825 56950 1825 7 FreeSans 240 0 -80 0 V_tail_gate
port 11 w
flabel metal2 57605 2830 57605 2830 3 FreeSans 200 0 80 0 err_amp_mir
flabel metal2 56900 3015 56900 3015 1 FreeSans 240 0 0 80 V_tot
flabel metal1 57240 3065 57240 3065 3 FreeSans 200 0 80 0 V_err_p
flabel metal2 57770 1770 57770 1770 3 FreeSans 240 0 80 0 VIN-
flabel metal2 56030 1770 56030 1770 7 FreeSans 240 0 -80 0 VIN+
flabel metal1 56835 3065 56835 3065 7 FreeSans 200 0 -80 0 V_err_gate
port 13 w
flabel metal2 55960 2775 55960 2775 7 FreeSans 200 0 -80 0 V_err_amp_ref
port 12 w
flabel metal2 57000 3535 57000 3535 5 FreeSans 200 0 0 -80 Vb3
port 4 s
flabel metal1 56855 3570 56855 3570 5 FreeSans 200 0 0 -80 Vb2
port 5 s
flabel metal2 57455 2575 57455 2575 7 FreeSans 240 0 -80 0 X
flabel metal1 59510 1070 59510 1070 5 FreeSans 240 0 0 -80 VOUT-
port 9 s
flabel metal1 57220 1235 57220 1235 3 FreeSans 240 0 80 0 V_source
flabel metal2 57720 1215 57720 1215 5 FreeSans 200 0 0 -80 V_b_2nd_stage
flabel metal1 56910 1205 56910 1205 3 FreeSans 200 0 80 0 V_p_mir
flabel metal1 59100 1950 59100 1950 1 FreeSans 240 0 0 80 V_CMFB_S1
port 2 n
flabel metal1 59055 1765 59055 1765 1 FreeSans 240 0 0 80 V_CMFB_S2
port 7 n
flabel metal2 56955 2695 56955 2695 1 FreeSans 240 0 0 80 err_amp_out
flabel metal1 56345 2565 56345 2565 3 FreeSans 240 0 80 0 Y
flabel metal2 56455 5015 56455 5015 1 FreeSans 240 0 0 80 Vb2_2
flabel metal2 57365 5015 57365 5015 1 FreeSans 240 0 0 80 Vb2_Vb3
flabel metal2 57950 4095 57950 4095 5 FreeSans 240 0 0 -80 VD3
flabel metal2 55865 4095 55865 4095 5 FreeSans 240 0 0 -80 VD4
flabel metal2 54290 1070 54290 1070 5 FreeSans 240 0 0 -80 VOUT+
port 10 s
flabel metal2 54700 1950 54700 1950 1 FreeSans 240 0 0 80 V_CMFB_S3
port 3 n
flabel metal2 54745 1765 54745 1765 1 FreeSans 240 0 0 80 V_CMFB_S4
port 8 n
<< end >>
