* NGSPICE file created from vco2_3.ext - technology: sky130A

**.subckt vco2_3 VDDA V_OSC V_CONT GNDA
X0 a_3910_10# a_3870_n240# a_3270_n240# VDDA sky130_fd_pr__pfet_01v8 ad=0.44 pd=3 as=0.44 ps=3 w=1.1 l=0.2
X1 a_4510_n780# VDDA GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X2 a_3310_10# a_2390_720# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X3 a_3910_n780# VDDA GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X4 a_4510_n780# V_OSC a_3870_n240# GNDA sky130_fd_pr__nfet_01v8 ad=0.22 pd=1.9 as=0.22 ps=1.9 w=0.55 l=0.2
X5 a_4510_n780# V_CONT GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X6 a_4510_10# a_2390_720# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X7 a_3910_10# a_2390_720# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X8 a_3910_n780# a_3870_n240# a_3270_n240# GNDA sky130_fd_pr__nfet_01v8 ad=0.22 pd=1.9 as=0.22 ps=1.9 w=0.55 l=0.2
X9 a_3910_n780# V_CONT GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X10 a_3310_10# a_3270_n240# V_OSC VDDA sky130_fd_pr__pfet_01v8 ad=0.44 pd=3 as=0.44 ps=3 w=1.1 l=0.2
X11 GNDA V_CONT a_2390_720# GNDA sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X12 a_3310_10# GNDA VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X13 a_4510_10# GNDA VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X14 a_4510_10# V_OSC a_3870_n240# VDDA sky130_fd_pr__pfet_01v8 ad=0.44 pd=3 as=0.44 ps=3 w=1.1 l=0.2
X15 VDDA a_2390_720# a_2390_720# VDDA sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X16 a_3910_10# GNDA VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X17 a_3310_n780# VDDA GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X18 a_3310_n780# a_3270_n240# V_OSC GNDA sky130_fd_pr__nfet_01v8 ad=0.22 pd=1.9 as=0.22 ps=1.9 w=0.55 l=0.2
X19 a_3310_n780# V_CONT GNDA GNDA sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
.ends

