magic
tech sky130A
timestamp 1749295395
<< error_p >>
rect -2925 -390 -2917 -382
rect -2913 -390 -2905 -382
rect -2933 -398 -2897 -390
rect -2925 -402 -2905 -398
rect -2933 -410 -2897 -402
rect -2925 -418 -2917 -410
rect -2913 -418 -2905 -410
<< nwell >>
rect 2545 1880 5285 2950
<< pwell >>
rect 10955 3550 11100 3580
rect 10490 3230 10710 3293
rect 10820 3230 11100 3550
rect 11220 3175 12580 3575
rect 18455 3550 18600 3580
rect 12890 2940 14140 3240
rect 17990 3230 18210 3293
rect 18320 3230 18600 3550
rect 18720 3175 20080 3575
rect 20390 2940 21640 3240
rect 9680 2520 10930 2620
rect 11220 2495 12580 2895
rect 12890 2520 14140 2620
rect 17180 2520 18430 2620
rect 18720 2495 20080 2895
rect 20390 2520 21640 2620
rect 9680 2020 10930 2170
rect 11275 1980 12525 2130
rect 12890 2020 14140 2170
rect 17180 2020 18430 2170
rect 18775 1980 20025 2130
rect 20390 2020 21640 2170
rect -45 1685 130 1725
rect 20490 1705 20860 1855
rect 3165 1615 3805 1665
rect 4205 1615 4845 1665
rect 11030 1515 11730 1665
rect 11770 1515 12030 1665
rect 12070 1515 12770 1665
rect 18530 1515 19230 1665
rect 19270 1515 19530 1665
rect 19570 1515 20270 1665
rect 2835 1205 3955 1455
rect 4055 1205 5175 1455
rect 20395 1370 20655 1520
rect 20695 1370 20955 1520
rect 2945 975 5065 1075
rect 11205 925 12620 1175
rect 12925 990 14165 1270
rect 18705 975 20120 1225
rect 20545 1030 20805 1180
rect 2995 780 5015 880
rect 9275 -1010 10515 -730
<< nmos >>
rect 10530 3230 10550 3293
rect 10590 3230 10610 3293
rect 10650 3230 10670 3293
rect 10860 3230 10880 3550
rect 10920 3230 10940 3550
rect 10980 3230 11000 3580
rect 11040 3230 11060 3580
rect 11260 3175 11280 3575
rect 11320 3175 11340 3575
rect 11380 3175 11400 3575
rect 11440 3175 11460 3575
rect 11500 3175 11520 3575
rect 11560 3175 11580 3575
rect 11620 3175 11640 3575
rect 11680 3175 11700 3575
rect 11740 3175 11760 3575
rect 11800 3175 11820 3575
rect 11860 3175 11880 3575
rect 11920 3175 11940 3575
rect 11980 3175 12000 3575
rect 12040 3175 12060 3575
rect 12100 3175 12120 3575
rect 12160 3175 12180 3575
rect 12220 3175 12240 3575
rect 12280 3175 12300 3575
rect 12340 3175 12360 3575
rect 12400 3175 12420 3575
rect 12460 3175 12480 3575
rect 12520 3175 12540 3575
rect 12930 2940 12945 3240
rect 12985 2940 13000 3240
rect 13040 2940 13055 3240
rect 13095 2940 13110 3240
rect 13150 2940 13165 3240
rect 13205 2940 13220 3240
rect 13260 2940 13275 3240
rect 13315 2940 13330 3240
rect 13370 2940 13385 3240
rect 13425 2940 13440 3240
rect 13480 2940 13495 3240
rect 13535 2940 13550 3240
rect 13590 2940 13605 3240
rect 13645 2940 13660 3240
rect 13700 2940 13715 3240
rect 13755 2940 13770 3240
rect 13810 2940 13825 3240
rect 13865 2940 13880 3240
rect 13920 2940 13935 3240
rect 13975 2940 13990 3240
rect 14030 2940 14045 3240
rect 14085 2940 14100 3240
rect 18030 3230 18050 3293
rect 18090 3230 18110 3293
rect 18150 3230 18170 3293
rect 18360 3230 18380 3550
rect 18420 3230 18440 3550
rect 18480 3230 18500 3580
rect 18540 3230 18560 3580
rect 18760 3175 18780 3575
rect 18820 3175 18840 3575
rect 18880 3175 18900 3575
rect 18940 3175 18960 3575
rect 19000 3175 19020 3575
rect 19060 3175 19080 3575
rect 19120 3175 19140 3575
rect 19180 3175 19200 3575
rect 19240 3175 19260 3575
rect 19300 3175 19320 3575
rect 19360 3175 19380 3575
rect 19420 3175 19440 3575
rect 19480 3175 19500 3575
rect 19540 3175 19560 3575
rect 19600 3175 19620 3575
rect 19660 3175 19680 3575
rect 19720 3175 19740 3575
rect 19780 3175 19800 3575
rect 19840 3175 19860 3575
rect 19900 3175 19920 3575
rect 19960 3175 19980 3575
rect 20020 3175 20040 3575
rect 9720 2520 9735 2620
rect 9775 2520 9790 2620
rect 9830 2520 9845 2620
rect 9885 2520 9900 2620
rect 9940 2520 9955 2620
rect 9995 2520 10010 2620
rect 10050 2520 10065 2620
rect 10105 2520 10120 2620
rect 10160 2520 10175 2620
rect 10215 2520 10230 2620
rect 10270 2520 10285 2620
rect 10325 2520 10340 2620
rect 10380 2520 10395 2620
rect 10435 2520 10450 2620
rect 10490 2520 10505 2620
rect 10545 2520 10560 2620
rect 10600 2520 10615 2620
rect 10655 2520 10670 2620
rect 10710 2520 10725 2620
rect 10765 2520 10780 2620
rect 10820 2520 10835 2620
rect 10875 2520 10890 2620
rect 11260 2495 11280 2895
rect 11320 2495 11340 2895
rect 11380 2495 11400 2895
rect 11440 2495 11460 2895
rect 11500 2495 11520 2895
rect 11560 2495 11580 2895
rect 11620 2495 11640 2895
rect 11680 2495 11700 2895
rect 11740 2495 11760 2895
rect 11800 2495 11820 2895
rect 11860 2495 11880 2895
rect 11920 2495 11940 2895
rect 11980 2495 12000 2895
rect 12040 2495 12060 2895
rect 12100 2495 12120 2895
rect 12160 2495 12180 2895
rect 12220 2495 12240 2895
rect 12280 2495 12300 2895
rect 12340 2495 12360 2895
rect 12400 2495 12420 2895
rect 12460 2495 12480 2895
rect 12520 2495 12540 2895
rect 20430 2940 20445 3240
rect 20485 2940 20500 3240
rect 20540 2940 20555 3240
rect 20595 2940 20610 3240
rect 20650 2940 20665 3240
rect 20705 2940 20720 3240
rect 20760 2940 20775 3240
rect 20815 2940 20830 3240
rect 20870 2940 20885 3240
rect 20925 2940 20940 3240
rect 20980 2940 20995 3240
rect 21035 2940 21050 3240
rect 21090 2940 21105 3240
rect 21145 2940 21160 3240
rect 21200 2940 21215 3240
rect 21255 2940 21270 3240
rect 21310 2940 21325 3240
rect 21365 2940 21380 3240
rect 21420 2940 21435 3240
rect 21475 2940 21490 3240
rect 21530 2940 21545 3240
rect 21585 2940 21600 3240
rect 12930 2520 12945 2620
rect 12985 2520 13000 2620
rect 13040 2520 13055 2620
rect 13095 2520 13110 2620
rect 13150 2520 13165 2620
rect 13205 2520 13220 2620
rect 13260 2520 13275 2620
rect 13315 2520 13330 2620
rect 13370 2520 13385 2620
rect 13425 2520 13440 2620
rect 13480 2520 13495 2620
rect 13535 2520 13550 2620
rect 13590 2520 13605 2620
rect 13645 2520 13660 2620
rect 13700 2520 13715 2620
rect 13755 2520 13770 2620
rect 13810 2520 13825 2620
rect 13865 2520 13880 2620
rect 13920 2520 13935 2620
rect 13975 2520 13990 2620
rect 14030 2520 14045 2620
rect 14085 2520 14100 2620
rect 17220 2520 17235 2620
rect 17275 2520 17290 2620
rect 17330 2520 17345 2620
rect 17385 2520 17400 2620
rect 17440 2520 17455 2620
rect 17495 2520 17510 2620
rect 17550 2520 17565 2620
rect 17605 2520 17620 2620
rect 17660 2520 17675 2620
rect 17715 2520 17730 2620
rect 17770 2520 17785 2620
rect 17825 2520 17840 2620
rect 17880 2520 17895 2620
rect 17935 2520 17950 2620
rect 17990 2520 18005 2620
rect 18045 2520 18060 2620
rect 18100 2520 18115 2620
rect 18155 2520 18170 2620
rect 18210 2520 18225 2620
rect 18265 2520 18280 2620
rect 18320 2520 18335 2620
rect 18375 2520 18390 2620
rect 18760 2495 18780 2895
rect 18820 2495 18840 2895
rect 18880 2495 18900 2895
rect 18940 2495 18960 2895
rect 19000 2495 19020 2895
rect 19060 2495 19080 2895
rect 19120 2495 19140 2895
rect 19180 2495 19200 2895
rect 19240 2495 19260 2895
rect 19300 2495 19320 2895
rect 19360 2495 19380 2895
rect 19420 2495 19440 2895
rect 19480 2495 19500 2895
rect 19540 2495 19560 2895
rect 19600 2495 19620 2895
rect 19660 2495 19680 2895
rect 19720 2495 19740 2895
rect 19780 2495 19800 2895
rect 19840 2495 19860 2895
rect 19900 2495 19920 2895
rect 19960 2495 19980 2895
rect 20020 2495 20040 2895
rect 20430 2520 20445 2620
rect 20485 2520 20500 2620
rect 20540 2520 20555 2620
rect 20595 2520 20610 2620
rect 20650 2520 20665 2620
rect 20705 2520 20720 2620
rect 20760 2520 20775 2620
rect 20815 2520 20830 2620
rect 20870 2520 20885 2620
rect 20925 2520 20940 2620
rect 20980 2520 20995 2620
rect 21035 2520 21050 2620
rect 21090 2520 21105 2620
rect 21145 2520 21160 2620
rect 21200 2520 21215 2620
rect 21255 2520 21270 2620
rect 21310 2520 21325 2620
rect 21365 2520 21380 2620
rect 21420 2520 21435 2620
rect 21475 2520 21490 2620
rect 21530 2520 21545 2620
rect 21585 2520 21600 2620
rect 9720 2020 9735 2170
rect 9775 2020 9790 2170
rect 9830 2020 9845 2170
rect 9885 2020 9900 2170
rect 9940 2020 9955 2170
rect 9995 2020 10010 2170
rect 10050 2020 10065 2170
rect 10105 2020 10120 2170
rect 10160 2020 10175 2170
rect 10215 2020 10230 2170
rect 10270 2020 10285 2170
rect 10325 2020 10340 2170
rect 10380 2020 10395 2170
rect 10435 2020 10450 2170
rect 10490 2020 10505 2170
rect 10545 2020 10560 2170
rect 10600 2020 10615 2170
rect 10655 2020 10670 2170
rect 10710 2020 10725 2170
rect 10765 2020 10780 2170
rect 10820 2020 10835 2170
rect 10875 2020 10890 2170
rect 11315 1980 11330 2130
rect 11370 1980 11385 2130
rect 11425 1980 11440 2130
rect 11480 1980 11495 2130
rect 11535 1980 11550 2130
rect 11590 1980 11605 2130
rect 11645 1980 11660 2130
rect 11700 1980 11715 2130
rect 11755 1980 11770 2130
rect 11810 1980 11825 2130
rect 11865 1980 11880 2130
rect 11920 1980 11935 2130
rect 11975 1980 11990 2130
rect 12030 1980 12045 2130
rect 12085 1980 12100 2130
rect 12140 1980 12155 2130
rect 12195 1980 12210 2130
rect 12250 1980 12265 2130
rect 12305 1980 12320 2130
rect 12360 1980 12375 2130
rect 12415 1980 12430 2130
rect 12470 1980 12485 2130
rect 12930 2020 12945 2170
rect 12985 2020 13000 2170
rect 13040 2020 13055 2170
rect 13095 2020 13110 2170
rect 13150 2020 13165 2170
rect 13205 2020 13220 2170
rect 13260 2020 13275 2170
rect 13315 2020 13330 2170
rect 13370 2020 13385 2170
rect 13425 2020 13440 2170
rect 13480 2020 13495 2170
rect 13535 2020 13550 2170
rect 13590 2020 13605 2170
rect 13645 2020 13660 2170
rect 13700 2020 13715 2170
rect 13755 2020 13770 2170
rect 13810 2020 13825 2170
rect 13865 2020 13880 2170
rect 13920 2020 13935 2170
rect 13975 2020 13990 2170
rect 14030 2020 14045 2170
rect 14085 2020 14100 2170
rect 17220 2020 17235 2170
rect 17275 2020 17290 2170
rect 17330 2020 17345 2170
rect 17385 2020 17400 2170
rect 17440 2020 17455 2170
rect 17495 2020 17510 2170
rect 17550 2020 17565 2170
rect 17605 2020 17620 2170
rect 17660 2020 17675 2170
rect 17715 2020 17730 2170
rect 17770 2020 17785 2170
rect 17825 2020 17840 2170
rect 17880 2020 17895 2170
rect 17935 2020 17950 2170
rect 17990 2020 18005 2170
rect 18045 2020 18060 2170
rect 18100 2020 18115 2170
rect 18155 2020 18170 2170
rect 18210 2020 18225 2170
rect 18265 2020 18280 2170
rect 18320 2020 18335 2170
rect 18375 2020 18390 2170
rect 18815 1980 18830 2130
rect 18870 1980 18885 2130
rect 18925 1980 18940 2130
rect 18980 1980 18995 2130
rect 19035 1980 19050 2130
rect 19090 1980 19105 2130
rect 19145 1980 19160 2130
rect 19200 1980 19215 2130
rect 19255 1980 19270 2130
rect 19310 1980 19325 2130
rect 19365 1980 19380 2130
rect 19420 1980 19435 2130
rect 19475 1980 19490 2130
rect 19530 1980 19545 2130
rect 19585 1980 19600 2130
rect 19640 1980 19655 2130
rect 19695 1980 19710 2130
rect 19750 1980 19765 2130
rect 19805 1980 19820 2130
rect 19860 1980 19875 2130
rect 19915 1980 19930 2130
rect 19970 1980 19985 2130
rect 20430 2020 20445 2170
rect 20485 2020 20500 2170
rect 20540 2020 20555 2170
rect 20595 2020 20610 2170
rect 20650 2020 20665 2170
rect 20705 2020 20720 2170
rect 20760 2020 20775 2170
rect 20815 2020 20830 2170
rect 20870 2020 20885 2170
rect 20925 2020 20940 2170
rect 20980 2020 20995 2170
rect 21035 2020 21050 2170
rect 21090 2020 21105 2170
rect 21145 2020 21160 2170
rect 21200 2020 21215 2170
rect 21255 2020 21270 2170
rect 21310 2020 21325 2170
rect 21365 2020 21380 2170
rect 21420 2020 21435 2170
rect 21475 2020 21490 2170
rect 21530 2020 21545 2170
rect 21585 2020 21600 2170
rect 20530 1705 20545 1855
rect 20585 1705 20600 1855
rect 20640 1705 20655 1855
rect 20695 1705 20710 1855
rect 20750 1705 20765 1855
rect 20805 1705 20820 1855
rect 3205 1615 3225 1665
rect 3265 1615 3285 1665
rect 3325 1615 3345 1665
rect 3385 1615 3405 1665
rect 3445 1615 3465 1665
rect 3505 1615 3525 1665
rect 3565 1615 3585 1665
rect 3625 1615 3645 1665
rect 3685 1615 3705 1665
rect 3745 1615 3765 1665
rect 4245 1615 4265 1665
rect 4305 1615 4325 1665
rect 4365 1615 4385 1665
rect 4425 1615 4445 1665
rect 4485 1615 4505 1665
rect 4545 1615 4565 1665
rect 4605 1615 4625 1665
rect 4665 1615 4685 1665
rect 4725 1615 4745 1665
rect 4785 1615 4805 1665
rect 11070 1515 11085 1665
rect 11125 1515 11140 1665
rect 11180 1515 11195 1665
rect 11235 1515 11250 1665
rect 11290 1515 11305 1665
rect 11345 1515 11360 1665
rect 11400 1515 11415 1665
rect 11455 1515 11470 1665
rect 11510 1515 11525 1665
rect 11565 1515 11580 1665
rect 11620 1515 11635 1665
rect 11675 1515 11690 1665
rect 11810 1515 11825 1665
rect 11865 1515 11880 1665
rect 11920 1515 11935 1665
rect 11975 1515 11990 1665
rect 12110 1515 12125 1665
rect 12165 1515 12180 1665
rect 12220 1515 12235 1665
rect 12275 1515 12290 1665
rect 12330 1515 12345 1665
rect 12385 1515 12400 1665
rect 12440 1515 12455 1665
rect 12495 1515 12510 1665
rect 12550 1515 12565 1665
rect 12605 1515 12620 1665
rect 12660 1515 12675 1665
rect 12715 1515 12730 1665
rect 18570 1515 18585 1665
rect 18625 1515 18640 1665
rect 18680 1515 18695 1665
rect 18735 1515 18750 1665
rect 18790 1515 18805 1665
rect 18845 1515 18860 1665
rect 18900 1515 18915 1665
rect 18955 1515 18970 1665
rect 19010 1515 19025 1665
rect 19065 1515 19080 1665
rect 19120 1515 19135 1665
rect 19175 1515 19190 1665
rect 19310 1515 19325 1665
rect 19365 1515 19380 1665
rect 19420 1515 19435 1665
rect 19475 1515 19490 1665
rect 19610 1515 19625 1665
rect 19665 1515 19680 1665
rect 19720 1515 19735 1665
rect 19775 1515 19790 1665
rect 19830 1515 19845 1665
rect 19885 1515 19900 1665
rect 19940 1515 19955 1665
rect 19995 1515 20010 1665
rect 20050 1515 20065 1665
rect 20105 1515 20120 1665
rect 20160 1515 20175 1665
rect 20215 1515 20230 1665
rect 2875 1205 3375 1455
rect 3415 1205 3915 1455
rect 4095 1205 4595 1455
rect 4635 1205 5135 1455
rect 20435 1370 20450 1520
rect 20490 1370 20505 1520
rect 20545 1370 20560 1520
rect 20600 1370 20615 1520
rect 20735 1370 20750 1520
rect 20790 1370 20805 1520
rect 20845 1370 20860 1520
rect 20900 1370 20915 1520
rect 2985 975 3985 1075
rect 4025 975 5025 1075
rect 11245 925 11260 1175
rect 11300 925 11315 1175
rect 11355 925 11370 1175
rect 11410 925 11425 1175
rect 11465 925 11480 1175
rect 11520 925 11535 1175
rect 11575 925 11590 1175
rect 11630 925 11645 1175
rect 11685 925 11700 1175
rect 11740 925 11755 1175
rect 11795 925 11810 1175
rect 11850 925 11865 1175
rect 11905 925 11920 1175
rect 11960 925 11975 1175
rect 12015 925 12030 1175
rect 12070 925 12085 1175
rect 12125 925 12140 1175
rect 12180 925 12195 1175
rect 12235 925 12250 1175
rect 12290 925 12305 1175
rect 12345 925 12360 1175
rect 12400 925 12415 1175
rect 12455 925 12470 1175
rect 12510 925 12525 1175
rect 12565 925 12580 1175
rect 12965 990 13025 1270
rect 13065 990 13125 1270
rect 13165 990 13225 1270
rect 13265 990 13325 1270
rect 13365 990 13425 1270
rect 13465 990 13525 1270
rect 13565 990 13625 1270
rect 13665 990 13725 1270
rect 13765 990 13825 1270
rect 13865 990 13925 1270
rect 13965 990 14025 1270
rect 14065 990 14125 1270
rect 18745 975 18760 1225
rect 18800 975 18815 1225
rect 18855 975 18870 1225
rect 18910 975 18925 1225
rect 18965 975 18980 1225
rect 19020 975 19035 1225
rect 19075 975 19090 1225
rect 19130 975 19145 1225
rect 19185 975 19200 1225
rect 19240 975 19255 1225
rect 19295 975 19310 1225
rect 19350 975 19365 1225
rect 19405 975 19420 1225
rect 19460 975 19475 1225
rect 19515 975 19530 1225
rect 19570 975 19585 1225
rect 19625 975 19640 1225
rect 19680 975 19695 1225
rect 19735 975 19750 1225
rect 19790 975 19805 1225
rect 19845 975 19860 1225
rect 19900 975 19915 1225
rect 19955 975 19970 1225
rect 20010 975 20025 1225
rect 20065 975 20080 1225
rect 20585 1030 20600 1180
rect 20640 1030 20655 1180
rect 20695 1030 20710 1180
rect 20750 1030 20765 1180
rect 3035 780 3085 880
rect 3125 780 3175 880
rect 3215 780 3265 880
rect 3305 780 3355 880
rect 3395 780 3445 880
rect 3485 780 3535 880
rect 3575 780 3625 880
rect 3665 780 3715 880
rect 3755 780 3805 880
rect 3845 780 3895 880
rect 3935 780 3985 880
rect 4025 780 4075 880
rect 4115 780 4165 880
rect 4205 780 4255 880
rect 4295 780 4345 880
rect 4385 780 4435 880
rect 4475 780 4525 880
rect 4565 780 4615 880
rect 4655 780 4705 880
rect 4745 780 4795 880
rect 4835 780 4885 880
rect 4925 780 4975 880
rect 9315 -1010 9375 -730
rect 9415 -1010 9475 -730
rect 9515 -1010 9575 -730
rect 9615 -1010 9675 -730
rect 9715 -1010 9775 -730
rect 9815 -1010 9875 -730
rect 9915 -1010 9975 -730
rect 10015 -1010 10075 -730
rect 10115 -1010 10175 -730
rect 10215 -1010 10275 -730
rect 10315 -1010 10375 -730
rect 10415 -1010 10475 -730
<< pmos >>
rect 3035 2830 3085 2930
rect 3125 2830 3175 2930
rect 3215 2830 3265 2930
rect 3305 2830 3355 2930
rect 3395 2830 3445 2930
rect 3485 2830 3535 2930
rect 3575 2830 3625 2930
rect 3665 2830 3715 2930
rect 3755 2830 3805 2930
rect 3845 2830 3895 2930
rect 3935 2830 3985 2930
rect 4025 2830 4075 2930
rect 4115 2830 4165 2930
rect 4205 2830 4255 2930
rect 4295 2830 4345 2930
rect 4385 2830 4435 2930
rect 4475 2830 4525 2930
rect 4565 2830 4615 2930
rect 4655 2830 4705 2930
rect 4745 2830 4795 2930
rect 4835 2830 4885 2930
rect 4925 2830 4975 2930
rect 3215 2400 3265 2700
rect 3305 2400 3355 2700
rect 3395 2400 3445 2700
rect 3485 2400 3535 2700
rect 3575 2400 3625 2700
rect 3665 2400 3715 2700
rect 3755 2400 3805 2700
rect 3845 2400 3895 2700
rect 3935 2400 3985 2700
rect 4025 2400 4075 2700
rect 4115 2400 4165 2700
rect 4205 2400 4255 2700
rect 4295 2400 4345 2700
rect 4385 2400 4435 2700
rect 4475 2400 4525 2700
rect 4565 2400 4615 2700
rect 4655 2400 4705 2700
rect 4745 2400 4795 2700
rect 2605 1900 2620 2000
rect 2660 1900 2675 2000
rect 2785 1900 2805 2000
rect 2845 1900 2865 2000
rect 2905 1900 2925 2000
rect 2965 1900 2985 2000
rect 3025 1900 3045 2000
rect 3085 1900 3105 2000
rect 3145 1900 3165 2000
rect 3205 1900 3225 2000
rect 3265 1900 3285 2000
rect 3325 1900 3345 2000
rect 3385 1900 3405 2000
rect 3445 1900 3465 2000
rect 3505 1900 3525 2000
rect 3565 1900 3585 2000
rect 3625 1900 3645 2000
rect 3685 1900 3705 2000
rect 3745 1900 3765 2000
rect 3805 1900 3825 2000
rect 3865 1900 3885 2000
rect 3925 1900 3945 2000
rect 4065 1900 4085 2000
rect 4125 1900 4145 2000
rect 4185 1900 4205 2000
rect 4245 1900 4265 2000
rect 4305 1900 4325 2000
rect 4365 1900 4385 2000
rect 4425 1900 4445 2000
rect 4485 1900 4505 2000
rect 4545 1900 4565 2000
rect 4605 1900 4625 2000
rect 4665 1900 4685 2000
rect 4725 1900 4745 2000
rect 4785 1900 4805 2000
rect 4845 1900 4865 2000
rect 4905 1900 4925 2000
rect 4965 1900 4985 2000
rect 5025 1900 5045 2000
rect 5085 1900 5105 2000
rect 5145 1900 5165 2000
rect 5205 1900 5225 2000
<< ndiff >>
rect 10955 3550 10980 3580
rect 10820 3515 10860 3550
rect 10820 3495 10830 3515
rect 10850 3495 10860 3515
rect 10820 3465 10860 3495
rect 10820 3445 10830 3465
rect 10850 3445 10860 3465
rect 10820 3415 10860 3445
rect 10820 3395 10830 3415
rect 10850 3395 10860 3415
rect 10820 3365 10860 3395
rect 10820 3345 10830 3365
rect 10850 3345 10860 3365
rect 10820 3315 10860 3345
rect 10820 3295 10830 3315
rect 10850 3295 10860 3315
rect 10490 3265 10530 3293
rect 10490 3245 10500 3265
rect 10520 3245 10530 3265
rect 10490 3230 10530 3245
rect 10550 3270 10590 3293
rect 10550 3250 10560 3270
rect 10580 3250 10590 3270
rect 10550 3230 10590 3250
rect 10610 3270 10650 3293
rect 10610 3250 10620 3270
rect 10640 3250 10650 3270
rect 10610 3230 10650 3250
rect 10670 3265 10710 3293
rect 10670 3245 10680 3265
rect 10700 3245 10710 3265
rect 10670 3230 10710 3245
rect 10820 3265 10860 3295
rect 10820 3245 10830 3265
rect 10850 3245 10860 3265
rect 10820 3230 10860 3245
rect 10880 3515 10920 3550
rect 10880 3495 10890 3515
rect 10910 3495 10920 3515
rect 10880 3465 10920 3495
rect 10880 3445 10890 3465
rect 10910 3445 10920 3465
rect 10880 3415 10920 3445
rect 10880 3395 10890 3415
rect 10910 3395 10920 3415
rect 10880 3365 10920 3395
rect 10880 3345 10890 3365
rect 10910 3345 10920 3365
rect 10880 3315 10920 3345
rect 10880 3295 10890 3315
rect 10910 3295 10920 3315
rect 10880 3265 10920 3295
rect 10880 3245 10890 3265
rect 10910 3245 10920 3265
rect 10880 3230 10920 3245
rect 10940 3515 10980 3550
rect 10940 3495 10950 3515
rect 10970 3495 10980 3515
rect 10940 3465 10980 3495
rect 10940 3445 10950 3465
rect 10970 3445 10980 3465
rect 10940 3415 10980 3445
rect 10940 3395 10950 3415
rect 10970 3395 10980 3415
rect 10940 3365 10980 3395
rect 10940 3345 10950 3365
rect 10970 3345 10980 3365
rect 10940 3315 10980 3345
rect 10940 3295 10950 3315
rect 10970 3295 10980 3315
rect 10940 3265 10980 3295
rect 10940 3245 10950 3265
rect 10970 3245 10980 3265
rect 10940 3230 10980 3245
rect 11000 3565 11040 3580
rect 11000 3545 11010 3565
rect 11030 3545 11040 3565
rect 11000 3515 11040 3545
rect 11000 3495 11010 3515
rect 11030 3495 11040 3515
rect 11000 3465 11040 3495
rect 11000 3445 11010 3465
rect 11030 3445 11040 3465
rect 11000 3415 11040 3445
rect 11000 3395 11010 3415
rect 11030 3395 11040 3415
rect 11000 3365 11040 3395
rect 11000 3345 11010 3365
rect 11030 3345 11040 3365
rect 11000 3315 11040 3345
rect 11000 3295 11010 3315
rect 11030 3295 11040 3315
rect 11000 3265 11040 3295
rect 11000 3245 11010 3265
rect 11030 3245 11040 3265
rect 11000 3230 11040 3245
rect 11060 3565 11100 3580
rect 11060 3545 11070 3565
rect 11090 3545 11100 3565
rect 11060 3515 11100 3545
rect 11060 3495 11070 3515
rect 11090 3495 11100 3515
rect 11060 3465 11100 3495
rect 11060 3445 11070 3465
rect 11090 3445 11100 3465
rect 11060 3415 11100 3445
rect 11060 3395 11070 3415
rect 11090 3395 11100 3415
rect 11060 3365 11100 3395
rect 11060 3345 11070 3365
rect 11090 3345 11100 3365
rect 11060 3315 11100 3345
rect 11060 3295 11070 3315
rect 11090 3295 11100 3315
rect 11060 3265 11100 3295
rect 11060 3245 11070 3265
rect 11090 3245 11100 3265
rect 11060 3230 11100 3245
rect 11220 3560 11260 3575
rect 11220 3540 11230 3560
rect 11250 3540 11260 3560
rect 11220 3510 11260 3540
rect 11220 3490 11230 3510
rect 11250 3490 11260 3510
rect 11220 3460 11260 3490
rect 11220 3440 11230 3460
rect 11250 3440 11260 3460
rect 11220 3410 11260 3440
rect 11220 3390 11230 3410
rect 11250 3390 11260 3410
rect 11220 3360 11260 3390
rect 11220 3340 11230 3360
rect 11250 3340 11260 3360
rect 11220 3310 11260 3340
rect 11220 3290 11230 3310
rect 11250 3290 11260 3310
rect 11220 3260 11260 3290
rect 11220 3240 11230 3260
rect 11250 3240 11260 3260
rect 11220 3210 11260 3240
rect 11220 3190 11230 3210
rect 11250 3190 11260 3210
rect 11220 3175 11260 3190
rect 11280 3560 11320 3575
rect 11280 3540 11290 3560
rect 11310 3540 11320 3560
rect 11280 3510 11320 3540
rect 11280 3490 11290 3510
rect 11310 3490 11320 3510
rect 11280 3460 11320 3490
rect 11280 3440 11290 3460
rect 11310 3440 11320 3460
rect 11280 3410 11320 3440
rect 11280 3390 11290 3410
rect 11310 3390 11320 3410
rect 11280 3360 11320 3390
rect 11280 3340 11290 3360
rect 11310 3340 11320 3360
rect 11280 3310 11320 3340
rect 11280 3290 11290 3310
rect 11310 3290 11320 3310
rect 11280 3260 11320 3290
rect 11280 3240 11290 3260
rect 11310 3240 11320 3260
rect 11280 3210 11320 3240
rect 11280 3190 11290 3210
rect 11310 3190 11320 3210
rect 11280 3175 11320 3190
rect 11340 3560 11380 3575
rect 11340 3540 11350 3560
rect 11370 3540 11380 3560
rect 11340 3510 11380 3540
rect 11340 3490 11350 3510
rect 11370 3490 11380 3510
rect 11340 3460 11380 3490
rect 11340 3440 11350 3460
rect 11370 3440 11380 3460
rect 11340 3410 11380 3440
rect 11340 3390 11350 3410
rect 11370 3390 11380 3410
rect 11340 3360 11380 3390
rect 11340 3340 11350 3360
rect 11370 3340 11380 3360
rect 11340 3310 11380 3340
rect 11340 3290 11350 3310
rect 11370 3290 11380 3310
rect 11340 3260 11380 3290
rect 11340 3240 11350 3260
rect 11370 3240 11380 3260
rect 11340 3210 11380 3240
rect 11340 3190 11350 3210
rect 11370 3190 11380 3210
rect 11340 3175 11380 3190
rect 11400 3560 11440 3575
rect 11400 3540 11410 3560
rect 11430 3540 11440 3560
rect 11400 3510 11440 3540
rect 11400 3490 11410 3510
rect 11430 3490 11440 3510
rect 11400 3460 11440 3490
rect 11400 3440 11410 3460
rect 11430 3440 11440 3460
rect 11400 3410 11440 3440
rect 11400 3390 11410 3410
rect 11430 3390 11440 3410
rect 11400 3360 11440 3390
rect 11400 3340 11410 3360
rect 11430 3340 11440 3360
rect 11400 3310 11440 3340
rect 11400 3290 11410 3310
rect 11430 3290 11440 3310
rect 11400 3260 11440 3290
rect 11400 3240 11410 3260
rect 11430 3240 11440 3260
rect 11400 3210 11440 3240
rect 11400 3190 11410 3210
rect 11430 3190 11440 3210
rect 11400 3175 11440 3190
rect 11460 3560 11500 3575
rect 11460 3540 11470 3560
rect 11490 3540 11500 3560
rect 11460 3510 11500 3540
rect 11460 3490 11470 3510
rect 11490 3490 11500 3510
rect 11460 3460 11500 3490
rect 11460 3440 11470 3460
rect 11490 3440 11500 3460
rect 11460 3410 11500 3440
rect 11460 3390 11470 3410
rect 11490 3390 11500 3410
rect 11460 3360 11500 3390
rect 11460 3340 11470 3360
rect 11490 3340 11500 3360
rect 11460 3310 11500 3340
rect 11460 3290 11470 3310
rect 11490 3290 11500 3310
rect 11460 3260 11500 3290
rect 11460 3240 11470 3260
rect 11490 3240 11500 3260
rect 11460 3210 11500 3240
rect 11460 3190 11470 3210
rect 11490 3190 11500 3210
rect 11460 3175 11500 3190
rect 11520 3560 11560 3575
rect 11520 3540 11530 3560
rect 11550 3540 11560 3560
rect 11520 3510 11560 3540
rect 11520 3490 11530 3510
rect 11550 3490 11560 3510
rect 11520 3460 11560 3490
rect 11520 3440 11530 3460
rect 11550 3440 11560 3460
rect 11520 3410 11560 3440
rect 11520 3390 11530 3410
rect 11550 3390 11560 3410
rect 11520 3360 11560 3390
rect 11520 3340 11530 3360
rect 11550 3340 11560 3360
rect 11520 3310 11560 3340
rect 11520 3290 11530 3310
rect 11550 3290 11560 3310
rect 11520 3260 11560 3290
rect 11520 3240 11530 3260
rect 11550 3240 11560 3260
rect 11520 3210 11560 3240
rect 11520 3190 11530 3210
rect 11550 3190 11560 3210
rect 11520 3175 11560 3190
rect 11580 3560 11620 3575
rect 11580 3540 11590 3560
rect 11610 3540 11620 3560
rect 11580 3510 11620 3540
rect 11580 3490 11590 3510
rect 11610 3490 11620 3510
rect 11580 3460 11620 3490
rect 11580 3440 11590 3460
rect 11610 3440 11620 3460
rect 11580 3410 11620 3440
rect 11580 3390 11590 3410
rect 11610 3390 11620 3410
rect 11580 3360 11620 3390
rect 11580 3340 11590 3360
rect 11610 3340 11620 3360
rect 11580 3310 11620 3340
rect 11580 3290 11590 3310
rect 11610 3290 11620 3310
rect 11580 3260 11620 3290
rect 11580 3240 11590 3260
rect 11610 3240 11620 3260
rect 11580 3210 11620 3240
rect 11580 3190 11590 3210
rect 11610 3190 11620 3210
rect 11580 3175 11620 3190
rect 11640 3560 11680 3575
rect 11640 3540 11650 3560
rect 11670 3540 11680 3560
rect 11640 3510 11680 3540
rect 11640 3490 11650 3510
rect 11670 3490 11680 3510
rect 11640 3460 11680 3490
rect 11640 3440 11650 3460
rect 11670 3440 11680 3460
rect 11640 3410 11680 3440
rect 11640 3390 11650 3410
rect 11670 3390 11680 3410
rect 11640 3360 11680 3390
rect 11640 3340 11650 3360
rect 11670 3340 11680 3360
rect 11640 3310 11680 3340
rect 11640 3290 11650 3310
rect 11670 3290 11680 3310
rect 11640 3260 11680 3290
rect 11640 3240 11650 3260
rect 11670 3240 11680 3260
rect 11640 3210 11680 3240
rect 11640 3190 11650 3210
rect 11670 3190 11680 3210
rect 11640 3175 11680 3190
rect 11700 3560 11740 3575
rect 11700 3540 11710 3560
rect 11730 3540 11740 3560
rect 11700 3510 11740 3540
rect 11700 3490 11710 3510
rect 11730 3490 11740 3510
rect 11700 3460 11740 3490
rect 11700 3440 11710 3460
rect 11730 3440 11740 3460
rect 11700 3410 11740 3440
rect 11700 3390 11710 3410
rect 11730 3390 11740 3410
rect 11700 3360 11740 3390
rect 11700 3340 11710 3360
rect 11730 3340 11740 3360
rect 11700 3310 11740 3340
rect 11700 3290 11710 3310
rect 11730 3290 11740 3310
rect 11700 3260 11740 3290
rect 11700 3240 11710 3260
rect 11730 3240 11740 3260
rect 11700 3210 11740 3240
rect 11700 3190 11710 3210
rect 11730 3190 11740 3210
rect 11700 3175 11740 3190
rect 11760 3560 11800 3575
rect 11760 3540 11770 3560
rect 11790 3540 11800 3560
rect 11760 3510 11800 3540
rect 11760 3490 11770 3510
rect 11790 3490 11800 3510
rect 11760 3460 11800 3490
rect 11760 3440 11770 3460
rect 11790 3440 11800 3460
rect 11760 3410 11800 3440
rect 11760 3390 11770 3410
rect 11790 3390 11800 3410
rect 11760 3360 11800 3390
rect 11760 3340 11770 3360
rect 11790 3340 11800 3360
rect 11760 3310 11800 3340
rect 11760 3290 11770 3310
rect 11790 3290 11800 3310
rect 11760 3260 11800 3290
rect 11760 3240 11770 3260
rect 11790 3240 11800 3260
rect 11760 3210 11800 3240
rect 11760 3190 11770 3210
rect 11790 3190 11800 3210
rect 11760 3175 11800 3190
rect 11820 3560 11860 3575
rect 11820 3540 11830 3560
rect 11850 3540 11860 3560
rect 11820 3510 11860 3540
rect 11820 3490 11830 3510
rect 11850 3490 11860 3510
rect 11820 3460 11860 3490
rect 11820 3440 11830 3460
rect 11850 3440 11860 3460
rect 11820 3410 11860 3440
rect 11820 3390 11830 3410
rect 11850 3390 11860 3410
rect 11820 3360 11860 3390
rect 11820 3340 11830 3360
rect 11850 3340 11860 3360
rect 11820 3310 11860 3340
rect 11820 3290 11830 3310
rect 11850 3290 11860 3310
rect 11820 3260 11860 3290
rect 11820 3240 11830 3260
rect 11850 3240 11860 3260
rect 11820 3210 11860 3240
rect 11820 3190 11830 3210
rect 11850 3190 11860 3210
rect 11820 3175 11860 3190
rect 11880 3560 11920 3575
rect 11880 3540 11890 3560
rect 11910 3540 11920 3560
rect 11880 3510 11920 3540
rect 11880 3490 11890 3510
rect 11910 3490 11920 3510
rect 11880 3460 11920 3490
rect 11880 3440 11890 3460
rect 11910 3440 11920 3460
rect 11880 3410 11920 3440
rect 11880 3390 11890 3410
rect 11910 3390 11920 3410
rect 11880 3360 11920 3390
rect 11880 3340 11890 3360
rect 11910 3340 11920 3360
rect 11880 3310 11920 3340
rect 11880 3290 11890 3310
rect 11910 3290 11920 3310
rect 11880 3260 11920 3290
rect 11880 3240 11890 3260
rect 11910 3240 11920 3260
rect 11880 3210 11920 3240
rect 11880 3190 11890 3210
rect 11910 3190 11920 3210
rect 11880 3175 11920 3190
rect 11940 3560 11980 3575
rect 11940 3540 11950 3560
rect 11970 3540 11980 3560
rect 11940 3510 11980 3540
rect 11940 3490 11950 3510
rect 11970 3490 11980 3510
rect 11940 3460 11980 3490
rect 11940 3440 11950 3460
rect 11970 3440 11980 3460
rect 11940 3410 11980 3440
rect 11940 3390 11950 3410
rect 11970 3390 11980 3410
rect 11940 3360 11980 3390
rect 11940 3340 11950 3360
rect 11970 3340 11980 3360
rect 11940 3310 11980 3340
rect 11940 3290 11950 3310
rect 11970 3290 11980 3310
rect 11940 3260 11980 3290
rect 11940 3240 11950 3260
rect 11970 3240 11980 3260
rect 11940 3210 11980 3240
rect 11940 3190 11950 3210
rect 11970 3190 11980 3210
rect 11940 3175 11980 3190
rect 12000 3560 12040 3575
rect 12000 3540 12010 3560
rect 12030 3540 12040 3560
rect 12000 3510 12040 3540
rect 12000 3490 12010 3510
rect 12030 3490 12040 3510
rect 12000 3460 12040 3490
rect 12000 3440 12010 3460
rect 12030 3440 12040 3460
rect 12000 3410 12040 3440
rect 12000 3390 12010 3410
rect 12030 3390 12040 3410
rect 12000 3360 12040 3390
rect 12000 3340 12010 3360
rect 12030 3340 12040 3360
rect 12000 3310 12040 3340
rect 12000 3290 12010 3310
rect 12030 3290 12040 3310
rect 12000 3260 12040 3290
rect 12000 3240 12010 3260
rect 12030 3240 12040 3260
rect 12000 3210 12040 3240
rect 12000 3190 12010 3210
rect 12030 3190 12040 3210
rect 12000 3175 12040 3190
rect 12060 3560 12100 3575
rect 12060 3540 12070 3560
rect 12090 3540 12100 3560
rect 12060 3510 12100 3540
rect 12060 3490 12070 3510
rect 12090 3490 12100 3510
rect 12060 3460 12100 3490
rect 12060 3440 12070 3460
rect 12090 3440 12100 3460
rect 12060 3410 12100 3440
rect 12060 3390 12070 3410
rect 12090 3390 12100 3410
rect 12060 3360 12100 3390
rect 12060 3340 12070 3360
rect 12090 3340 12100 3360
rect 12060 3310 12100 3340
rect 12060 3290 12070 3310
rect 12090 3290 12100 3310
rect 12060 3260 12100 3290
rect 12060 3240 12070 3260
rect 12090 3240 12100 3260
rect 12060 3210 12100 3240
rect 12060 3190 12070 3210
rect 12090 3190 12100 3210
rect 12060 3175 12100 3190
rect 12120 3560 12160 3575
rect 12120 3540 12130 3560
rect 12150 3540 12160 3560
rect 12120 3510 12160 3540
rect 12120 3490 12130 3510
rect 12150 3490 12160 3510
rect 12120 3460 12160 3490
rect 12120 3440 12130 3460
rect 12150 3440 12160 3460
rect 12120 3410 12160 3440
rect 12120 3390 12130 3410
rect 12150 3390 12160 3410
rect 12120 3360 12160 3390
rect 12120 3340 12130 3360
rect 12150 3340 12160 3360
rect 12120 3310 12160 3340
rect 12120 3290 12130 3310
rect 12150 3290 12160 3310
rect 12120 3260 12160 3290
rect 12120 3240 12130 3260
rect 12150 3240 12160 3260
rect 12120 3210 12160 3240
rect 12120 3190 12130 3210
rect 12150 3190 12160 3210
rect 12120 3175 12160 3190
rect 12180 3560 12220 3575
rect 12180 3540 12190 3560
rect 12210 3540 12220 3560
rect 12180 3510 12220 3540
rect 12180 3490 12190 3510
rect 12210 3490 12220 3510
rect 12180 3460 12220 3490
rect 12180 3440 12190 3460
rect 12210 3440 12220 3460
rect 12180 3410 12220 3440
rect 12180 3390 12190 3410
rect 12210 3390 12220 3410
rect 12180 3360 12220 3390
rect 12180 3340 12190 3360
rect 12210 3340 12220 3360
rect 12180 3310 12220 3340
rect 12180 3290 12190 3310
rect 12210 3290 12220 3310
rect 12180 3260 12220 3290
rect 12180 3240 12190 3260
rect 12210 3240 12220 3260
rect 12180 3210 12220 3240
rect 12180 3190 12190 3210
rect 12210 3190 12220 3210
rect 12180 3175 12220 3190
rect 12240 3560 12280 3575
rect 12240 3540 12250 3560
rect 12270 3540 12280 3560
rect 12240 3510 12280 3540
rect 12240 3490 12250 3510
rect 12270 3490 12280 3510
rect 12240 3460 12280 3490
rect 12240 3440 12250 3460
rect 12270 3440 12280 3460
rect 12240 3410 12280 3440
rect 12240 3390 12250 3410
rect 12270 3390 12280 3410
rect 12240 3360 12280 3390
rect 12240 3340 12250 3360
rect 12270 3340 12280 3360
rect 12240 3310 12280 3340
rect 12240 3290 12250 3310
rect 12270 3290 12280 3310
rect 12240 3260 12280 3290
rect 12240 3240 12250 3260
rect 12270 3240 12280 3260
rect 12240 3210 12280 3240
rect 12240 3190 12250 3210
rect 12270 3190 12280 3210
rect 12240 3175 12280 3190
rect 12300 3560 12340 3575
rect 12300 3540 12310 3560
rect 12330 3540 12340 3560
rect 12300 3510 12340 3540
rect 12300 3490 12310 3510
rect 12330 3490 12340 3510
rect 12300 3460 12340 3490
rect 12300 3440 12310 3460
rect 12330 3440 12340 3460
rect 12300 3410 12340 3440
rect 12300 3390 12310 3410
rect 12330 3390 12340 3410
rect 12300 3360 12340 3390
rect 12300 3340 12310 3360
rect 12330 3340 12340 3360
rect 12300 3310 12340 3340
rect 12300 3290 12310 3310
rect 12330 3290 12340 3310
rect 12300 3260 12340 3290
rect 12300 3240 12310 3260
rect 12330 3240 12340 3260
rect 12300 3210 12340 3240
rect 12300 3190 12310 3210
rect 12330 3190 12340 3210
rect 12300 3175 12340 3190
rect 12360 3560 12400 3575
rect 12360 3540 12370 3560
rect 12390 3540 12400 3560
rect 12360 3510 12400 3540
rect 12360 3490 12370 3510
rect 12390 3490 12400 3510
rect 12360 3460 12400 3490
rect 12360 3440 12370 3460
rect 12390 3440 12400 3460
rect 12360 3410 12400 3440
rect 12360 3390 12370 3410
rect 12390 3390 12400 3410
rect 12360 3360 12400 3390
rect 12360 3340 12370 3360
rect 12390 3340 12400 3360
rect 12360 3310 12400 3340
rect 12360 3290 12370 3310
rect 12390 3290 12400 3310
rect 12360 3260 12400 3290
rect 12360 3240 12370 3260
rect 12390 3240 12400 3260
rect 12360 3210 12400 3240
rect 12360 3190 12370 3210
rect 12390 3190 12400 3210
rect 12360 3175 12400 3190
rect 12420 3560 12460 3575
rect 12420 3540 12430 3560
rect 12450 3540 12460 3560
rect 12420 3510 12460 3540
rect 12420 3490 12430 3510
rect 12450 3490 12460 3510
rect 12420 3460 12460 3490
rect 12420 3440 12430 3460
rect 12450 3440 12460 3460
rect 12420 3410 12460 3440
rect 12420 3390 12430 3410
rect 12450 3390 12460 3410
rect 12420 3360 12460 3390
rect 12420 3340 12430 3360
rect 12450 3340 12460 3360
rect 12420 3310 12460 3340
rect 12420 3290 12430 3310
rect 12450 3290 12460 3310
rect 12420 3260 12460 3290
rect 12420 3240 12430 3260
rect 12450 3240 12460 3260
rect 12420 3210 12460 3240
rect 12420 3190 12430 3210
rect 12450 3190 12460 3210
rect 12420 3175 12460 3190
rect 12480 3560 12520 3575
rect 12480 3540 12490 3560
rect 12510 3540 12520 3560
rect 12480 3510 12520 3540
rect 12480 3490 12490 3510
rect 12510 3490 12520 3510
rect 12480 3460 12520 3490
rect 12480 3440 12490 3460
rect 12510 3440 12520 3460
rect 12480 3410 12520 3440
rect 12480 3390 12490 3410
rect 12510 3390 12520 3410
rect 12480 3360 12520 3390
rect 12480 3340 12490 3360
rect 12510 3340 12520 3360
rect 12480 3310 12520 3340
rect 12480 3290 12490 3310
rect 12510 3290 12520 3310
rect 12480 3260 12520 3290
rect 12480 3240 12490 3260
rect 12510 3240 12520 3260
rect 12480 3210 12520 3240
rect 12480 3190 12490 3210
rect 12510 3190 12520 3210
rect 12480 3175 12520 3190
rect 12540 3560 12580 3575
rect 12540 3540 12550 3560
rect 12570 3540 12580 3560
rect 18455 3550 18480 3580
rect 12540 3510 12580 3540
rect 12540 3490 12550 3510
rect 12570 3490 12580 3510
rect 12540 3460 12580 3490
rect 12540 3440 12550 3460
rect 12570 3440 12580 3460
rect 12540 3410 12580 3440
rect 12540 3390 12550 3410
rect 12570 3390 12580 3410
rect 12540 3360 12580 3390
rect 12540 3340 12550 3360
rect 12570 3340 12580 3360
rect 18320 3515 18360 3550
rect 18320 3495 18330 3515
rect 18350 3495 18360 3515
rect 18320 3465 18360 3495
rect 18320 3445 18330 3465
rect 18350 3445 18360 3465
rect 18320 3415 18360 3445
rect 18320 3395 18330 3415
rect 18350 3395 18360 3415
rect 18320 3365 18360 3395
rect 12540 3310 12580 3340
rect 12540 3290 12550 3310
rect 12570 3290 12580 3310
rect 18320 3345 18330 3365
rect 18350 3345 18360 3365
rect 18320 3315 18360 3345
rect 18320 3295 18330 3315
rect 18350 3295 18360 3315
rect 12540 3260 12580 3290
rect 12540 3240 12550 3260
rect 12570 3240 12580 3260
rect 17990 3265 18030 3293
rect 17990 3245 18000 3265
rect 18020 3245 18030 3265
rect 12540 3210 12580 3240
rect 12540 3190 12550 3210
rect 12570 3190 12580 3210
rect 12540 3175 12580 3190
rect 12890 3225 12930 3240
rect 12890 3205 12900 3225
rect 12920 3205 12930 3225
rect 12890 3175 12930 3205
rect 12890 3155 12900 3175
rect 12920 3155 12930 3175
rect 12890 3125 12930 3155
rect 12890 3105 12900 3125
rect 12920 3105 12930 3125
rect 12890 3075 12930 3105
rect 12890 3055 12900 3075
rect 12920 3055 12930 3075
rect 12890 3025 12930 3055
rect 12890 3005 12900 3025
rect 12920 3005 12930 3025
rect 12890 2975 12930 3005
rect 12890 2955 12900 2975
rect 12920 2955 12930 2975
rect 12890 2940 12930 2955
rect 12945 3225 12985 3240
rect 12945 3205 12955 3225
rect 12975 3205 12985 3225
rect 12945 3175 12985 3205
rect 12945 3155 12955 3175
rect 12975 3155 12985 3175
rect 12945 3125 12985 3155
rect 12945 3105 12955 3125
rect 12975 3105 12985 3125
rect 12945 3075 12985 3105
rect 12945 3055 12955 3075
rect 12975 3055 12985 3075
rect 12945 3025 12985 3055
rect 12945 3005 12955 3025
rect 12975 3005 12985 3025
rect 12945 2975 12985 3005
rect 12945 2955 12955 2975
rect 12975 2955 12985 2975
rect 12945 2940 12985 2955
rect 13000 3225 13040 3240
rect 13000 3205 13010 3225
rect 13030 3205 13040 3225
rect 13000 3175 13040 3205
rect 13000 3155 13010 3175
rect 13030 3155 13040 3175
rect 13000 3125 13040 3155
rect 13000 3105 13010 3125
rect 13030 3105 13040 3125
rect 13000 3075 13040 3105
rect 13000 3055 13010 3075
rect 13030 3055 13040 3075
rect 13000 3025 13040 3055
rect 13000 3005 13010 3025
rect 13030 3005 13040 3025
rect 13000 2975 13040 3005
rect 13000 2955 13010 2975
rect 13030 2955 13040 2975
rect 13000 2940 13040 2955
rect 13055 3225 13095 3240
rect 13055 3205 13065 3225
rect 13085 3205 13095 3225
rect 13055 3175 13095 3205
rect 13055 3155 13065 3175
rect 13085 3155 13095 3175
rect 13055 3125 13095 3155
rect 13055 3105 13065 3125
rect 13085 3105 13095 3125
rect 13055 3075 13095 3105
rect 13055 3055 13065 3075
rect 13085 3055 13095 3075
rect 13055 3025 13095 3055
rect 13055 3005 13065 3025
rect 13085 3005 13095 3025
rect 13055 2975 13095 3005
rect 13055 2955 13065 2975
rect 13085 2955 13095 2975
rect 13055 2940 13095 2955
rect 13110 3225 13150 3240
rect 13110 3205 13120 3225
rect 13140 3205 13150 3225
rect 13110 3175 13150 3205
rect 13110 3155 13120 3175
rect 13140 3155 13150 3175
rect 13110 3125 13150 3155
rect 13110 3105 13120 3125
rect 13140 3105 13150 3125
rect 13110 3075 13150 3105
rect 13110 3055 13120 3075
rect 13140 3055 13150 3075
rect 13110 3025 13150 3055
rect 13110 3005 13120 3025
rect 13140 3005 13150 3025
rect 13110 2975 13150 3005
rect 13110 2955 13120 2975
rect 13140 2955 13150 2975
rect 13110 2940 13150 2955
rect 13165 3225 13205 3240
rect 13165 3205 13175 3225
rect 13195 3205 13205 3225
rect 13165 3175 13205 3205
rect 13165 3155 13175 3175
rect 13195 3155 13205 3175
rect 13165 3125 13205 3155
rect 13165 3105 13175 3125
rect 13195 3105 13205 3125
rect 13165 3075 13205 3105
rect 13165 3055 13175 3075
rect 13195 3055 13205 3075
rect 13165 3025 13205 3055
rect 13165 3005 13175 3025
rect 13195 3005 13205 3025
rect 13165 2975 13205 3005
rect 13165 2955 13175 2975
rect 13195 2955 13205 2975
rect 13165 2940 13205 2955
rect 13220 3225 13260 3240
rect 13220 3205 13230 3225
rect 13250 3205 13260 3225
rect 13220 3175 13260 3205
rect 13220 3155 13230 3175
rect 13250 3155 13260 3175
rect 13220 3125 13260 3155
rect 13220 3105 13230 3125
rect 13250 3105 13260 3125
rect 13220 3075 13260 3105
rect 13220 3055 13230 3075
rect 13250 3055 13260 3075
rect 13220 3025 13260 3055
rect 13220 3005 13230 3025
rect 13250 3005 13260 3025
rect 13220 2975 13260 3005
rect 13220 2955 13230 2975
rect 13250 2955 13260 2975
rect 13220 2940 13260 2955
rect 13275 3225 13315 3240
rect 13275 3205 13285 3225
rect 13305 3205 13315 3225
rect 13275 3175 13315 3205
rect 13275 3155 13285 3175
rect 13305 3155 13315 3175
rect 13275 3125 13315 3155
rect 13275 3105 13285 3125
rect 13305 3105 13315 3125
rect 13275 3075 13315 3105
rect 13275 3055 13285 3075
rect 13305 3055 13315 3075
rect 13275 3025 13315 3055
rect 13275 3005 13285 3025
rect 13305 3005 13315 3025
rect 13275 2975 13315 3005
rect 13275 2955 13285 2975
rect 13305 2955 13315 2975
rect 13275 2940 13315 2955
rect 13330 3225 13370 3240
rect 13330 3205 13340 3225
rect 13360 3205 13370 3225
rect 13330 3175 13370 3205
rect 13330 3155 13340 3175
rect 13360 3155 13370 3175
rect 13330 3125 13370 3155
rect 13330 3105 13340 3125
rect 13360 3105 13370 3125
rect 13330 3075 13370 3105
rect 13330 3055 13340 3075
rect 13360 3055 13370 3075
rect 13330 3025 13370 3055
rect 13330 3005 13340 3025
rect 13360 3005 13370 3025
rect 13330 2975 13370 3005
rect 13330 2955 13340 2975
rect 13360 2955 13370 2975
rect 13330 2940 13370 2955
rect 13385 3225 13425 3240
rect 13385 3205 13395 3225
rect 13415 3205 13425 3225
rect 13385 3175 13425 3205
rect 13385 3155 13395 3175
rect 13415 3155 13425 3175
rect 13385 3125 13425 3155
rect 13385 3105 13395 3125
rect 13415 3105 13425 3125
rect 13385 3075 13425 3105
rect 13385 3055 13395 3075
rect 13415 3055 13425 3075
rect 13385 3025 13425 3055
rect 13385 3005 13395 3025
rect 13415 3005 13425 3025
rect 13385 2975 13425 3005
rect 13385 2955 13395 2975
rect 13415 2955 13425 2975
rect 13385 2940 13425 2955
rect 13440 3225 13480 3240
rect 13440 3205 13450 3225
rect 13470 3205 13480 3225
rect 13440 3175 13480 3205
rect 13440 3155 13450 3175
rect 13470 3155 13480 3175
rect 13440 3125 13480 3155
rect 13440 3105 13450 3125
rect 13470 3105 13480 3125
rect 13440 3075 13480 3105
rect 13440 3055 13450 3075
rect 13470 3055 13480 3075
rect 13440 3025 13480 3055
rect 13440 3005 13450 3025
rect 13470 3005 13480 3025
rect 13440 2975 13480 3005
rect 13440 2955 13450 2975
rect 13470 2955 13480 2975
rect 13440 2940 13480 2955
rect 13495 3225 13535 3240
rect 13495 3205 13505 3225
rect 13525 3205 13535 3225
rect 13495 3175 13535 3205
rect 13495 3155 13505 3175
rect 13525 3155 13535 3175
rect 13495 3125 13535 3155
rect 13495 3105 13505 3125
rect 13525 3105 13535 3125
rect 13495 3075 13535 3105
rect 13495 3055 13505 3075
rect 13525 3055 13535 3075
rect 13495 3025 13535 3055
rect 13495 3005 13505 3025
rect 13525 3005 13535 3025
rect 13495 2975 13535 3005
rect 13495 2955 13505 2975
rect 13525 2955 13535 2975
rect 13495 2940 13535 2955
rect 13550 3225 13590 3240
rect 13550 3205 13560 3225
rect 13580 3205 13590 3225
rect 13550 3175 13590 3205
rect 13550 3155 13560 3175
rect 13580 3155 13590 3175
rect 13550 3125 13590 3155
rect 13550 3105 13560 3125
rect 13580 3105 13590 3125
rect 13550 3075 13590 3105
rect 13550 3055 13560 3075
rect 13580 3055 13590 3075
rect 13550 3025 13590 3055
rect 13550 3005 13560 3025
rect 13580 3005 13590 3025
rect 13550 2975 13590 3005
rect 13550 2955 13560 2975
rect 13580 2955 13590 2975
rect 13550 2940 13590 2955
rect 13605 3225 13645 3240
rect 13605 3205 13615 3225
rect 13635 3205 13645 3225
rect 13605 3175 13645 3205
rect 13605 3155 13615 3175
rect 13635 3155 13645 3175
rect 13605 3125 13645 3155
rect 13605 3105 13615 3125
rect 13635 3105 13645 3125
rect 13605 3075 13645 3105
rect 13605 3055 13615 3075
rect 13635 3055 13645 3075
rect 13605 3025 13645 3055
rect 13605 3005 13615 3025
rect 13635 3005 13645 3025
rect 13605 2975 13645 3005
rect 13605 2955 13615 2975
rect 13635 2955 13645 2975
rect 13605 2940 13645 2955
rect 13660 3225 13700 3240
rect 13660 3205 13670 3225
rect 13690 3205 13700 3225
rect 13660 3175 13700 3205
rect 13660 3155 13670 3175
rect 13690 3155 13700 3175
rect 13660 3125 13700 3155
rect 13660 3105 13670 3125
rect 13690 3105 13700 3125
rect 13660 3075 13700 3105
rect 13660 3055 13670 3075
rect 13690 3055 13700 3075
rect 13660 3025 13700 3055
rect 13660 3005 13670 3025
rect 13690 3005 13700 3025
rect 13660 2975 13700 3005
rect 13660 2955 13670 2975
rect 13690 2955 13700 2975
rect 13660 2940 13700 2955
rect 13715 3225 13755 3240
rect 13715 3205 13725 3225
rect 13745 3205 13755 3225
rect 13715 3175 13755 3205
rect 13715 3155 13725 3175
rect 13745 3155 13755 3175
rect 13715 3125 13755 3155
rect 13715 3105 13725 3125
rect 13745 3105 13755 3125
rect 13715 3075 13755 3105
rect 13715 3055 13725 3075
rect 13745 3055 13755 3075
rect 13715 3025 13755 3055
rect 13715 3005 13725 3025
rect 13745 3005 13755 3025
rect 13715 2975 13755 3005
rect 13715 2955 13725 2975
rect 13745 2955 13755 2975
rect 13715 2940 13755 2955
rect 13770 3225 13810 3240
rect 13770 3205 13780 3225
rect 13800 3205 13810 3225
rect 13770 3175 13810 3205
rect 13770 3155 13780 3175
rect 13800 3155 13810 3175
rect 13770 3125 13810 3155
rect 13770 3105 13780 3125
rect 13800 3105 13810 3125
rect 13770 3075 13810 3105
rect 13770 3055 13780 3075
rect 13800 3055 13810 3075
rect 13770 3025 13810 3055
rect 13770 3005 13780 3025
rect 13800 3005 13810 3025
rect 13770 2975 13810 3005
rect 13770 2955 13780 2975
rect 13800 2955 13810 2975
rect 13770 2940 13810 2955
rect 13825 3225 13865 3240
rect 13825 3205 13835 3225
rect 13855 3205 13865 3225
rect 13825 3175 13865 3205
rect 13825 3155 13835 3175
rect 13855 3155 13865 3175
rect 13825 3125 13865 3155
rect 13825 3105 13835 3125
rect 13855 3105 13865 3125
rect 13825 3075 13865 3105
rect 13825 3055 13835 3075
rect 13855 3055 13865 3075
rect 13825 3025 13865 3055
rect 13825 3005 13835 3025
rect 13855 3005 13865 3025
rect 13825 2975 13865 3005
rect 13825 2955 13835 2975
rect 13855 2955 13865 2975
rect 13825 2940 13865 2955
rect 13880 3225 13920 3240
rect 13880 3205 13890 3225
rect 13910 3205 13920 3225
rect 13880 3175 13920 3205
rect 13880 3155 13890 3175
rect 13910 3155 13920 3175
rect 13880 3125 13920 3155
rect 13880 3105 13890 3125
rect 13910 3105 13920 3125
rect 13880 3075 13920 3105
rect 13880 3055 13890 3075
rect 13910 3055 13920 3075
rect 13880 3025 13920 3055
rect 13880 3005 13890 3025
rect 13910 3005 13920 3025
rect 13880 2975 13920 3005
rect 13880 2955 13890 2975
rect 13910 2955 13920 2975
rect 13880 2940 13920 2955
rect 13935 3225 13975 3240
rect 13935 3205 13945 3225
rect 13965 3205 13975 3225
rect 13935 3175 13975 3205
rect 13935 3155 13945 3175
rect 13965 3155 13975 3175
rect 13935 3125 13975 3155
rect 13935 3105 13945 3125
rect 13965 3105 13975 3125
rect 13935 3075 13975 3105
rect 13935 3055 13945 3075
rect 13965 3055 13975 3075
rect 13935 3025 13975 3055
rect 13935 3005 13945 3025
rect 13965 3005 13975 3025
rect 13935 2975 13975 3005
rect 13935 2955 13945 2975
rect 13965 2955 13975 2975
rect 13935 2940 13975 2955
rect 13990 3225 14030 3240
rect 13990 3205 14000 3225
rect 14020 3205 14030 3225
rect 13990 3175 14030 3205
rect 13990 3155 14000 3175
rect 14020 3155 14030 3175
rect 13990 3125 14030 3155
rect 13990 3105 14000 3125
rect 14020 3105 14030 3125
rect 13990 3075 14030 3105
rect 13990 3055 14000 3075
rect 14020 3055 14030 3075
rect 13990 3025 14030 3055
rect 13990 3005 14000 3025
rect 14020 3005 14030 3025
rect 13990 2975 14030 3005
rect 13990 2955 14000 2975
rect 14020 2955 14030 2975
rect 13990 2940 14030 2955
rect 14045 3225 14085 3240
rect 14045 3205 14055 3225
rect 14075 3205 14085 3225
rect 14045 3175 14085 3205
rect 14045 3155 14055 3175
rect 14075 3155 14085 3175
rect 14045 3125 14085 3155
rect 14045 3105 14055 3125
rect 14075 3105 14085 3125
rect 14045 3075 14085 3105
rect 14045 3055 14055 3075
rect 14075 3055 14085 3075
rect 14045 3025 14085 3055
rect 14045 3005 14055 3025
rect 14075 3005 14085 3025
rect 14045 2975 14085 3005
rect 14045 2955 14055 2975
rect 14075 2955 14085 2975
rect 14045 2940 14085 2955
rect 14100 3225 14140 3240
rect 17990 3230 18030 3245
rect 18050 3270 18090 3293
rect 18050 3250 18060 3270
rect 18080 3250 18090 3270
rect 18050 3230 18090 3250
rect 18110 3270 18150 3293
rect 18110 3250 18120 3270
rect 18140 3250 18150 3270
rect 18110 3230 18150 3250
rect 18170 3265 18210 3293
rect 18170 3245 18180 3265
rect 18200 3245 18210 3265
rect 18170 3230 18210 3245
rect 18320 3265 18360 3295
rect 18320 3245 18330 3265
rect 18350 3245 18360 3265
rect 18320 3230 18360 3245
rect 18380 3515 18420 3550
rect 18380 3495 18390 3515
rect 18410 3495 18420 3515
rect 18380 3465 18420 3495
rect 18380 3445 18390 3465
rect 18410 3445 18420 3465
rect 18380 3415 18420 3445
rect 18380 3395 18390 3415
rect 18410 3395 18420 3415
rect 18380 3365 18420 3395
rect 18380 3345 18390 3365
rect 18410 3345 18420 3365
rect 18380 3315 18420 3345
rect 18380 3295 18390 3315
rect 18410 3295 18420 3315
rect 18380 3265 18420 3295
rect 18380 3245 18390 3265
rect 18410 3245 18420 3265
rect 18380 3230 18420 3245
rect 18440 3515 18480 3550
rect 18440 3495 18450 3515
rect 18470 3495 18480 3515
rect 18440 3465 18480 3495
rect 18440 3445 18450 3465
rect 18470 3445 18480 3465
rect 18440 3415 18480 3445
rect 18440 3395 18450 3415
rect 18470 3395 18480 3415
rect 18440 3365 18480 3395
rect 18440 3345 18450 3365
rect 18470 3345 18480 3365
rect 18440 3315 18480 3345
rect 18440 3295 18450 3315
rect 18470 3295 18480 3315
rect 18440 3265 18480 3295
rect 18440 3245 18450 3265
rect 18470 3245 18480 3265
rect 18440 3230 18480 3245
rect 18500 3565 18540 3580
rect 18500 3545 18510 3565
rect 18530 3545 18540 3565
rect 18500 3515 18540 3545
rect 18500 3495 18510 3515
rect 18530 3495 18540 3515
rect 18500 3465 18540 3495
rect 18500 3445 18510 3465
rect 18530 3445 18540 3465
rect 18500 3415 18540 3445
rect 18500 3395 18510 3415
rect 18530 3395 18540 3415
rect 18500 3365 18540 3395
rect 18500 3345 18510 3365
rect 18530 3345 18540 3365
rect 18500 3315 18540 3345
rect 18500 3295 18510 3315
rect 18530 3295 18540 3315
rect 18500 3265 18540 3295
rect 18500 3245 18510 3265
rect 18530 3245 18540 3265
rect 18500 3230 18540 3245
rect 18560 3565 18600 3580
rect 18560 3545 18570 3565
rect 18590 3545 18600 3565
rect 18560 3515 18600 3545
rect 18560 3495 18570 3515
rect 18590 3495 18600 3515
rect 18560 3465 18600 3495
rect 18560 3445 18570 3465
rect 18590 3445 18600 3465
rect 18560 3415 18600 3445
rect 18560 3395 18570 3415
rect 18590 3395 18600 3415
rect 18560 3365 18600 3395
rect 18560 3345 18570 3365
rect 18590 3345 18600 3365
rect 18560 3315 18600 3345
rect 18560 3295 18570 3315
rect 18590 3295 18600 3315
rect 18560 3265 18600 3295
rect 18560 3245 18570 3265
rect 18590 3245 18600 3265
rect 18560 3230 18600 3245
rect 18720 3560 18760 3575
rect 18720 3540 18730 3560
rect 18750 3540 18760 3560
rect 18720 3510 18760 3540
rect 18720 3490 18730 3510
rect 18750 3490 18760 3510
rect 18720 3460 18760 3490
rect 18720 3440 18730 3460
rect 18750 3440 18760 3460
rect 18720 3410 18760 3440
rect 18720 3390 18730 3410
rect 18750 3390 18760 3410
rect 18720 3360 18760 3390
rect 18720 3340 18730 3360
rect 18750 3340 18760 3360
rect 18720 3310 18760 3340
rect 18720 3290 18730 3310
rect 18750 3290 18760 3310
rect 18720 3260 18760 3290
rect 18720 3240 18730 3260
rect 18750 3240 18760 3260
rect 14100 3205 14110 3225
rect 14130 3205 14140 3225
rect 14100 3175 14140 3205
rect 18720 3210 18760 3240
rect 18720 3190 18730 3210
rect 18750 3190 18760 3210
rect 18720 3175 18760 3190
rect 18780 3560 18820 3575
rect 18780 3540 18790 3560
rect 18810 3540 18820 3560
rect 18780 3510 18820 3540
rect 18780 3490 18790 3510
rect 18810 3490 18820 3510
rect 18780 3460 18820 3490
rect 18780 3440 18790 3460
rect 18810 3440 18820 3460
rect 18780 3410 18820 3440
rect 18780 3390 18790 3410
rect 18810 3390 18820 3410
rect 18780 3360 18820 3390
rect 18780 3340 18790 3360
rect 18810 3340 18820 3360
rect 18780 3310 18820 3340
rect 18780 3290 18790 3310
rect 18810 3290 18820 3310
rect 18780 3260 18820 3290
rect 18780 3240 18790 3260
rect 18810 3240 18820 3260
rect 18780 3210 18820 3240
rect 18780 3190 18790 3210
rect 18810 3190 18820 3210
rect 18780 3175 18820 3190
rect 18840 3560 18880 3575
rect 18840 3540 18850 3560
rect 18870 3540 18880 3560
rect 18840 3510 18880 3540
rect 18840 3490 18850 3510
rect 18870 3490 18880 3510
rect 18840 3460 18880 3490
rect 18840 3440 18850 3460
rect 18870 3440 18880 3460
rect 18840 3410 18880 3440
rect 18840 3390 18850 3410
rect 18870 3390 18880 3410
rect 18840 3360 18880 3390
rect 18840 3340 18850 3360
rect 18870 3340 18880 3360
rect 18840 3310 18880 3340
rect 18840 3290 18850 3310
rect 18870 3290 18880 3310
rect 18840 3260 18880 3290
rect 18840 3240 18850 3260
rect 18870 3240 18880 3260
rect 18840 3210 18880 3240
rect 18840 3190 18850 3210
rect 18870 3190 18880 3210
rect 18840 3175 18880 3190
rect 18900 3560 18940 3575
rect 18900 3540 18910 3560
rect 18930 3540 18940 3560
rect 18900 3510 18940 3540
rect 18900 3490 18910 3510
rect 18930 3490 18940 3510
rect 18900 3460 18940 3490
rect 18900 3440 18910 3460
rect 18930 3440 18940 3460
rect 18900 3410 18940 3440
rect 18900 3390 18910 3410
rect 18930 3390 18940 3410
rect 18900 3360 18940 3390
rect 18900 3340 18910 3360
rect 18930 3340 18940 3360
rect 18900 3310 18940 3340
rect 18900 3290 18910 3310
rect 18930 3290 18940 3310
rect 18900 3260 18940 3290
rect 18900 3240 18910 3260
rect 18930 3240 18940 3260
rect 18900 3210 18940 3240
rect 18900 3190 18910 3210
rect 18930 3190 18940 3210
rect 18900 3175 18940 3190
rect 18960 3560 19000 3575
rect 18960 3540 18970 3560
rect 18990 3540 19000 3560
rect 18960 3510 19000 3540
rect 18960 3490 18970 3510
rect 18990 3490 19000 3510
rect 18960 3460 19000 3490
rect 18960 3440 18970 3460
rect 18990 3440 19000 3460
rect 18960 3410 19000 3440
rect 18960 3390 18970 3410
rect 18990 3390 19000 3410
rect 18960 3360 19000 3390
rect 18960 3340 18970 3360
rect 18990 3340 19000 3360
rect 18960 3310 19000 3340
rect 18960 3290 18970 3310
rect 18990 3290 19000 3310
rect 18960 3260 19000 3290
rect 18960 3240 18970 3260
rect 18990 3240 19000 3260
rect 18960 3210 19000 3240
rect 18960 3190 18970 3210
rect 18990 3190 19000 3210
rect 18960 3175 19000 3190
rect 19020 3560 19060 3575
rect 19020 3540 19030 3560
rect 19050 3540 19060 3560
rect 19020 3510 19060 3540
rect 19020 3490 19030 3510
rect 19050 3490 19060 3510
rect 19020 3460 19060 3490
rect 19020 3440 19030 3460
rect 19050 3440 19060 3460
rect 19020 3410 19060 3440
rect 19020 3390 19030 3410
rect 19050 3390 19060 3410
rect 19020 3360 19060 3390
rect 19020 3340 19030 3360
rect 19050 3340 19060 3360
rect 19020 3310 19060 3340
rect 19020 3290 19030 3310
rect 19050 3290 19060 3310
rect 19020 3260 19060 3290
rect 19020 3240 19030 3260
rect 19050 3240 19060 3260
rect 19020 3210 19060 3240
rect 19020 3190 19030 3210
rect 19050 3190 19060 3210
rect 19020 3175 19060 3190
rect 19080 3560 19120 3575
rect 19080 3540 19090 3560
rect 19110 3540 19120 3560
rect 19080 3510 19120 3540
rect 19080 3490 19090 3510
rect 19110 3490 19120 3510
rect 19080 3460 19120 3490
rect 19080 3440 19090 3460
rect 19110 3440 19120 3460
rect 19080 3410 19120 3440
rect 19080 3390 19090 3410
rect 19110 3390 19120 3410
rect 19080 3360 19120 3390
rect 19080 3340 19090 3360
rect 19110 3340 19120 3360
rect 19080 3310 19120 3340
rect 19080 3290 19090 3310
rect 19110 3290 19120 3310
rect 19080 3260 19120 3290
rect 19080 3240 19090 3260
rect 19110 3240 19120 3260
rect 19080 3210 19120 3240
rect 19080 3190 19090 3210
rect 19110 3190 19120 3210
rect 19080 3175 19120 3190
rect 19140 3560 19180 3575
rect 19140 3540 19150 3560
rect 19170 3540 19180 3560
rect 19140 3510 19180 3540
rect 19140 3490 19150 3510
rect 19170 3490 19180 3510
rect 19140 3460 19180 3490
rect 19140 3440 19150 3460
rect 19170 3440 19180 3460
rect 19140 3410 19180 3440
rect 19140 3390 19150 3410
rect 19170 3390 19180 3410
rect 19140 3360 19180 3390
rect 19140 3340 19150 3360
rect 19170 3340 19180 3360
rect 19140 3310 19180 3340
rect 19140 3290 19150 3310
rect 19170 3290 19180 3310
rect 19140 3260 19180 3290
rect 19140 3240 19150 3260
rect 19170 3240 19180 3260
rect 19140 3210 19180 3240
rect 19140 3190 19150 3210
rect 19170 3190 19180 3210
rect 19140 3175 19180 3190
rect 19200 3560 19240 3575
rect 19200 3540 19210 3560
rect 19230 3540 19240 3560
rect 19200 3510 19240 3540
rect 19200 3490 19210 3510
rect 19230 3490 19240 3510
rect 19200 3460 19240 3490
rect 19200 3440 19210 3460
rect 19230 3440 19240 3460
rect 19200 3410 19240 3440
rect 19200 3390 19210 3410
rect 19230 3390 19240 3410
rect 19200 3360 19240 3390
rect 19200 3340 19210 3360
rect 19230 3340 19240 3360
rect 19200 3310 19240 3340
rect 19200 3290 19210 3310
rect 19230 3290 19240 3310
rect 19200 3260 19240 3290
rect 19200 3240 19210 3260
rect 19230 3240 19240 3260
rect 19200 3210 19240 3240
rect 19200 3190 19210 3210
rect 19230 3190 19240 3210
rect 19200 3175 19240 3190
rect 19260 3560 19300 3575
rect 19260 3540 19270 3560
rect 19290 3540 19300 3560
rect 19260 3510 19300 3540
rect 19260 3490 19270 3510
rect 19290 3490 19300 3510
rect 19260 3460 19300 3490
rect 19260 3440 19270 3460
rect 19290 3440 19300 3460
rect 19260 3410 19300 3440
rect 19260 3390 19270 3410
rect 19290 3390 19300 3410
rect 19260 3360 19300 3390
rect 19260 3340 19270 3360
rect 19290 3340 19300 3360
rect 19260 3310 19300 3340
rect 19260 3290 19270 3310
rect 19290 3290 19300 3310
rect 19260 3260 19300 3290
rect 19260 3240 19270 3260
rect 19290 3240 19300 3260
rect 19260 3210 19300 3240
rect 19260 3190 19270 3210
rect 19290 3190 19300 3210
rect 19260 3175 19300 3190
rect 19320 3560 19360 3575
rect 19320 3540 19330 3560
rect 19350 3540 19360 3560
rect 19320 3510 19360 3540
rect 19320 3490 19330 3510
rect 19350 3490 19360 3510
rect 19320 3460 19360 3490
rect 19320 3440 19330 3460
rect 19350 3440 19360 3460
rect 19320 3410 19360 3440
rect 19320 3390 19330 3410
rect 19350 3390 19360 3410
rect 19320 3360 19360 3390
rect 19320 3340 19330 3360
rect 19350 3340 19360 3360
rect 19320 3310 19360 3340
rect 19320 3290 19330 3310
rect 19350 3290 19360 3310
rect 19320 3260 19360 3290
rect 19320 3240 19330 3260
rect 19350 3240 19360 3260
rect 19320 3210 19360 3240
rect 19320 3190 19330 3210
rect 19350 3190 19360 3210
rect 19320 3175 19360 3190
rect 19380 3560 19420 3575
rect 19380 3540 19390 3560
rect 19410 3540 19420 3560
rect 19380 3510 19420 3540
rect 19380 3490 19390 3510
rect 19410 3490 19420 3510
rect 19380 3460 19420 3490
rect 19380 3440 19390 3460
rect 19410 3440 19420 3460
rect 19380 3410 19420 3440
rect 19380 3390 19390 3410
rect 19410 3390 19420 3410
rect 19380 3360 19420 3390
rect 19380 3340 19390 3360
rect 19410 3340 19420 3360
rect 19380 3310 19420 3340
rect 19380 3290 19390 3310
rect 19410 3290 19420 3310
rect 19380 3260 19420 3290
rect 19380 3240 19390 3260
rect 19410 3240 19420 3260
rect 19380 3210 19420 3240
rect 19380 3190 19390 3210
rect 19410 3190 19420 3210
rect 19380 3175 19420 3190
rect 19440 3560 19480 3575
rect 19440 3540 19450 3560
rect 19470 3540 19480 3560
rect 19440 3510 19480 3540
rect 19440 3490 19450 3510
rect 19470 3490 19480 3510
rect 19440 3460 19480 3490
rect 19440 3440 19450 3460
rect 19470 3440 19480 3460
rect 19440 3410 19480 3440
rect 19440 3390 19450 3410
rect 19470 3390 19480 3410
rect 19440 3360 19480 3390
rect 19440 3340 19450 3360
rect 19470 3340 19480 3360
rect 19440 3310 19480 3340
rect 19440 3290 19450 3310
rect 19470 3290 19480 3310
rect 19440 3260 19480 3290
rect 19440 3240 19450 3260
rect 19470 3240 19480 3260
rect 19440 3210 19480 3240
rect 19440 3190 19450 3210
rect 19470 3190 19480 3210
rect 19440 3175 19480 3190
rect 19500 3560 19540 3575
rect 19500 3540 19510 3560
rect 19530 3540 19540 3560
rect 19500 3510 19540 3540
rect 19500 3490 19510 3510
rect 19530 3490 19540 3510
rect 19500 3460 19540 3490
rect 19500 3440 19510 3460
rect 19530 3440 19540 3460
rect 19500 3410 19540 3440
rect 19500 3390 19510 3410
rect 19530 3390 19540 3410
rect 19500 3360 19540 3390
rect 19500 3340 19510 3360
rect 19530 3340 19540 3360
rect 19500 3310 19540 3340
rect 19500 3290 19510 3310
rect 19530 3290 19540 3310
rect 19500 3260 19540 3290
rect 19500 3240 19510 3260
rect 19530 3240 19540 3260
rect 19500 3210 19540 3240
rect 19500 3190 19510 3210
rect 19530 3190 19540 3210
rect 19500 3175 19540 3190
rect 19560 3560 19600 3575
rect 19560 3540 19570 3560
rect 19590 3540 19600 3560
rect 19560 3510 19600 3540
rect 19560 3490 19570 3510
rect 19590 3490 19600 3510
rect 19560 3460 19600 3490
rect 19560 3440 19570 3460
rect 19590 3440 19600 3460
rect 19560 3410 19600 3440
rect 19560 3390 19570 3410
rect 19590 3390 19600 3410
rect 19560 3360 19600 3390
rect 19560 3340 19570 3360
rect 19590 3340 19600 3360
rect 19560 3310 19600 3340
rect 19560 3290 19570 3310
rect 19590 3290 19600 3310
rect 19560 3260 19600 3290
rect 19560 3240 19570 3260
rect 19590 3240 19600 3260
rect 19560 3210 19600 3240
rect 19560 3190 19570 3210
rect 19590 3190 19600 3210
rect 19560 3175 19600 3190
rect 19620 3560 19660 3575
rect 19620 3540 19630 3560
rect 19650 3540 19660 3560
rect 19620 3510 19660 3540
rect 19620 3490 19630 3510
rect 19650 3490 19660 3510
rect 19620 3460 19660 3490
rect 19620 3440 19630 3460
rect 19650 3440 19660 3460
rect 19620 3410 19660 3440
rect 19620 3390 19630 3410
rect 19650 3390 19660 3410
rect 19620 3360 19660 3390
rect 19620 3340 19630 3360
rect 19650 3340 19660 3360
rect 19620 3310 19660 3340
rect 19620 3290 19630 3310
rect 19650 3290 19660 3310
rect 19620 3260 19660 3290
rect 19620 3240 19630 3260
rect 19650 3240 19660 3260
rect 19620 3210 19660 3240
rect 19620 3190 19630 3210
rect 19650 3190 19660 3210
rect 19620 3175 19660 3190
rect 19680 3560 19720 3575
rect 19680 3540 19690 3560
rect 19710 3540 19720 3560
rect 19680 3510 19720 3540
rect 19680 3490 19690 3510
rect 19710 3490 19720 3510
rect 19680 3460 19720 3490
rect 19680 3440 19690 3460
rect 19710 3440 19720 3460
rect 19680 3410 19720 3440
rect 19680 3390 19690 3410
rect 19710 3390 19720 3410
rect 19680 3360 19720 3390
rect 19680 3340 19690 3360
rect 19710 3340 19720 3360
rect 19680 3310 19720 3340
rect 19680 3290 19690 3310
rect 19710 3290 19720 3310
rect 19680 3260 19720 3290
rect 19680 3240 19690 3260
rect 19710 3240 19720 3260
rect 19680 3210 19720 3240
rect 19680 3190 19690 3210
rect 19710 3190 19720 3210
rect 19680 3175 19720 3190
rect 19740 3560 19780 3575
rect 19740 3540 19750 3560
rect 19770 3540 19780 3560
rect 19740 3510 19780 3540
rect 19740 3490 19750 3510
rect 19770 3490 19780 3510
rect 19740 3460 19780 3490
rect 19740 3440 19750 3460
rect 19770 3440 19780 3460
rect 19740 3410 19780 3440
rect 19740 3390 19750 3410
rect 19770 3390 19780 3410
rect 19740 3360 19780 3390
rect 19740 3340 19750 3360
rect 19770 3340 19780 3360
rect 19740 3310 19780 3340
rect 19740 3290 19750 3310
rect 19770 3290 19780 3310
rect 19740 3260 19780 3290
rect 19740 3240 19750 3260
rect 19770 3240 19780 3260
rect 19740 3210 19780 3240
rect 19740 3190 19750 3210
rect 19770 3190 19780 3210
rect 19740 3175 19780 3190
rect 19800 3560 19840 3575
rect 19800 3540 19810 3560
rect 19830 3540 19840 3560
rect 19800 3510 19840 3540
rect 19800 3490 19810 3510
rect 19830 3490 19840 3510
rect 19800 3460 19840 3490
rect 19800 3440 19810 3460
rect 19830 3440 19840 3460
rect 19800 3410 19840 3440
rect 19800 3390 19810 3410
rect 19830 3390 19840 3410
rect 19800 3360 19840 3390
rect 19800 3340 19810 3360
rect 19830 3340 19840 3360
rect 19800 3310 19840 3340
rect 19800 3290 19810 3310
rect 19830 3290 19840 3310
rect 19800 3260 19840 3290
rect 19800 3240 19810 3260
rect 19830 3240 19840 3260
rect 19800 3210 19840 3240
rect 19800 3190 19810 3210
rect 19830 3190 19840 3210
rect 19800 3175 19840 3190
rect 19860 3560 19900 3575
rect 19860 3540 19870 3560
rect 19890 3540 19900 3560
rect 19860 3510 19900 3540
rect 19860 3490 19870 3510
rect 19890 3490 19900 3510
rect 19860 3460 19900 3490
rect 19860 3440 19870 3460
rect 19890 3440 19900 3460
rect 19860 3410 19900 3440
rect 19860 3390 19870 3410
rect 19890 3390 19900 3410
rect 19860 3360 19900 3390
rect 19860 3340 19870 3360
rect 19890 3340 19900 3360
rect 19860 3310 19900 3340
rect 19860 3290 19870 3310
rect 19890 3290 19900 3310
rect 19860 3260 19900 3290
rect 19860 3240 19870 3260
rect 19890 3240 19900 3260
rect 19860 3210 19900 3240
rect 19860 3190 19870 3210
rect 19890 3190 19900 3210
rect 19860 3175 19900 3190
rect 19920 3560 19960 3575
rect 19920 3540 19930 3560
rect 19950 3540 19960 3560
rect 19920 3510 19960 3540
rect 19920 3490 19930 3510
rect 19950 3490 19960 3510
rect 19920 3460 19960 3490
rect 19920 3440 19930 3460
rect 19950 3440 19960 3460
rect 19920 3410 19960 3440
rect 19920 3390 19930 3410
rect 19950 3390 19960 3410
rect 19920 3360 19960 3390
rect 19920 3340 19930 3360
rect 19950 3340 19960 3360
rect 19920 3310 19960 3340
rect 19920 3290 19930 3310
rect 19950 3290 19960 3310
rect 19920 3260 19960 3290
rect 19920 3240 19930 3260
rect 19950 3240 19960 3260
rect 19920 3210 19960 3240
rect 19920 3190 19930 3210
rect 19950 3190 19960 3210
rect 19920 3175 19960 3190
rect 19980 3560 20020 3575
rect 19980 3540 19990 3560
rect 20010 3540 20020 3560
rect 19980 3510 20020 3540
rect 19980 3490 19990 3510
rect 20010 3490 20020 3510
rect 19980 3460 20020 3490
rect 19980 3440 19990 3460
rect 20010 3440 20020 3460
rect 19980 3410 20020 3440
rect 19980 3390 19990 3410
rect 20010 3390 20020 3410
rect 19980 3360 20020 3390
rect 19980 3340 19990 3360
rect 20010 3340 20020 3360
rect 19980 3310 20020 3340
rect 19980 3290 19990 3310
rect 20010 3290 20020 3310
rect 19980 3260 20020 3290
rect 19980 3240 19990 3260
rect 20010 3240 20020 3260
rect 19980 3210 20020 3240
rect 19980 3190 19990 3210
rect 20010 3190 20020 3210
rect 19980 3175 20020 3190
rect 20040 3560 20080 3575
rect 20040 3540 20050 3560
rect 20070 3540 20080 3560
rect 20040 3510 20080 3540
rect 20040 3490 20050 3510
rect 20070 3490 20080 3510
rect 20040 3460 20080 3490
rect 20040 3440 20050 3460
rect 20070 3440 20080 3460
rect 20040 3410 20080 3440
rect 20040 3390 20050 3410
rect 20070 3390 20080 3410
rect 20040 3360 20080 3390
rect 20040 3340 20050 3360
rect 20070 3340 20080 3360
rect 20040 3310 20080 3340
rect 20040 3290 20050 3310
rect 20070 3290 20080 3310
rect 20040 3260 20080 3290
rect 20040 3240 20050 3260
rect 20070 3240 20080 3260
rect 20040 3210 20080 3240
rect 20040 3190 20050 3210
rect 20070 3190 20080 3210
rect 20040 3175 20080 3190
rect 20390 3225 20430 3240
rect 20390 3205 20400 3225
rect 20420 3205 20430 3225
rect 20390 3175 20430 3205
rect 14100 3155 14110 3175
rect 14130 3155 14140 3175
rect 14100 3125 14140 3155
rect 20390 3155 20400 3175
rect 20420 3155 20430 3175
rect 14100 3105 14110 3125
rect 14130 3105 14140 3125
rect 20390 3125 20430 3155
rect 14100 3075 14140 3105
rect 14100 3055 14110 3075
rect 14130 3055 14140 3075
rect 14100 3025 14140 3055
rect 14100 3005 14110 3025
rect 14130 3005 14140 3025
rect 14100 2975 14140 3005
rect 14100 2955 14110 2975
rect 14130 2955 14140 2975
rect 14100 2940 14140 2955
rect 20390 3105 20400 3125
rect 20420 3105 20430 3125
rect 20390 3075 20430 3105
rect 20390 3055 20400 3075
rect 20420 3055 20430 3075
rect 20390 3025 20430 3055
rect 20390 3005 20400 3025
rect 20420 3005 20430 3025
rect 20390 2975 20430 3005
rect 20390 2955 20400 2975
rect 20420 2955 20430 2975
rect 11220 2880 11260 2895
rect 11220 2860 11230 2880
rect 11250 2860 11260 2880
rect 11220 2830 11260 2860
rect 11220 2810 11230 2830
rect 11250 2810 11260 2830
rect 11220 2780 11260 2810
rect 11220 2760 11230 2780
rect 11250 2760 11260 2780
rect 11220 2730 11260 2760
rect 11220 2710 11230 2730
rect 11250 2710 11260 2730
rect 11220 2680 11260 2710
rect 11220 2660 11230 2680
rect 11250 2660 11260 2680
rect 11220 2630 11260 2660
rect 9680 2605 9720 2620
rect 9680 2585 9690 2605
rect 9710 2585 9720 2605
rect 9680 2555 9720 2585
rect 9680 2535 9690 2555
rect 9710 2535 9720 2555
rect 9680 2520 9720 2535
rect 9735 2605 9775 2620
rect 9735 2585 9745 2605
rect 9765 2585 9775 2605
rect 9735 2555 9775 2585
rect 9735 2535 9745 2555
rect 9765 2535 9775 2555
rect 9735 2520 9775 2535
rect 9790 2605 9830 2620
rect 9790 2585 9800 2605
rect 9820 2585 9830 2605
rect 9790 2555 9830 2585
rect 9790 2535 9800 2555
rect 9820 2535 9830 2555
rect 9790 2520 9830 2535
rect 9845 2605 9885 2620
rect 9845 2585 9855 2605
rect 9875 2585 9885 2605
rect 9845 2555 9885 2585
rect 9845 2535 9855 2555
rect 9875 2535 9885 2555
rect 9845 2520 9885 2535
rect 9900 2605 9940 2620
rect 9900 2585 9910 2605
rect 9930 2585 9940 2605
rect 9900 2555 9940 2585
rect 9900 2535 9910 2555
rect 9930 2535 9940 2555
rect 9900 2520 9940 2535
rect 9955 2605 9995 2620
rect 9955 2585 9965 2605
rect 9985 2585 9995 2605
rect 9955 2555 9995 2585
rect 9955 2535 9965 2555
rect 9985 2535 9995 2555
rect 9955 2520 9995 2535
rect 10010 2605 10050 2620
rect 10010 2585 10020 2605
rect 10040 2585 10050 2605
rect 10010 2555 10050 2585
rect 10010 2535 10020 2555
rect 10040 2535 10050 2555
rect 10010 2520 10050 2535
rect 10065 2605 10105 2620
rect 10065 2585 10075 2605
rect 10095 2585 10105 2605
rect 10065 2555 10105 2585
rect 10065 2535 10075 2555
rect 10095 2535 10105 2555
rect 10065 2520 10105 2535
rect 10120 2605 10160 2620
rect 10120 2585 10130 2605
rect 10150 2585 10160 2605
rect 10120 2555 10160 2585
rect 10120 2535 10130 2555
rect 10150 2535 10160 2555
rect 10120 2520 10160 2535
rect 10175 2605 10215 2620
rect 10175 2585 10185 2605
rect 10205 2585 10215 2605
rect 10175 2555 10215 2585
rect 10175 2535 10185 2555
rect 10205 2535 10215 2555
rect 10175 2520 10215 2535
rect 10230 2605 10270 2620
rect 10230 2585 10240 2605
rect 10260 2585 10270 2605
rect 10230 2555 10270 2585
rect 10230 2535 10240 2555
rect 10260 2535 10270 2555
rect 10230 2520 10270 2535
rect 10285 2605 10325 2620
rect 10285 2585 10295 2605
rect 10315 2585 10325 2605
rect 10285 2555 10325 2585
rect 10285 2535 10295 2555
rect 10315 2535 10325 2555
rect 10285 2520 10325 2535
rect 10340 2605 10380 2620
rect 10340 2585 10350 2605
rect 10370 2585 10380 2605
rect 10340 2555 10380 2585
rect 10340 2535 10350 2555
rect 10370 2535 10380 2555
rect 10340 2520 10380 2535
rect 10395 2605 10435 2620
rect 10395 2585 10405 2605
rect 10425 2585 10435 2605
rect 10395 2555 10435 2585
rect 10395 2535 10405 2555
rect 10425 2535 10435 2555
rect 10395 2520 10435 2535
rect 10450 2605 10490 2620
rect 10450 2585 10460 2605
rect 10480 2585 10490 2605
rect 10450 2555 10490 2585
rect 10450 2535 10460 2555
rect 10480 2535 10490 2555
rect 10450 2520 10490 2535
rect 10505 2605 10545 2620
rect 10505 2585 10515 2605
rect 10535 2585 10545 2605
rect 10505 2555 10545 2585
rect 10505 2535 10515 2555
rect 10535 2535 10545 2555
rect 10505 2520 10545 2535
rect 10560 2605 10600 2620
rect 10560 2585 10570 2605
rect 10590 2585 10600 2605
rect 10560 2555 10600 2585
rect 10560 2535 10570 2555
rect 10590 2535 10600 2555
rect 10560 2520 10600 2535
rect 10615 2605 10655 2620
rect 10615 2585 10625 2605
rect 10645 2585 10655 2605
rect 10615 2555 10655 2585
rect 10615 2535 10625 2555
rect 10645 2535 10655 2555
rect 10615 2520 10655 2535
rect 10670 2605 10710 2620
rect 10670 2585 10680 2605
rect 10700 2585 10710 2605
rect 10670 2555 10710 2585
rect 10670 2535 10680 2555
rect 10700 2535 10710 2555
rect 10670 2520 10710 2535
rect 10725 2605 10765 2620
rect 10725 2585 10735 2605
rect 10755 2585 10765 2605
rect 10725 2555 10765 2585
rect 10725 2535 10735 2555
rect 10755 2535 10765 2555
rect 10725 2520 10765 2535
rect 10780 2605 10820 2620
rect 10780 2585 10790 2605
rect 10810 2585 10820 2605
rect 10780 2555 10820 2585
rect 10780 2535 10790 2555
rect 10810 2535 10820 2555
rect 10780 2520 10820 2535
rect 10835 2605 10875 2620
rect 10835 2585 10845 2605
rect 10865 2585 10875 2605
rect 10835 2555 10875 2585
rect 10835 2535 10845 2555
rect 10865 2535 10875 2555
rect 10835 2520 10875 2535
rect 10890 2605 10930 2620
rect 10890 2585 10900 2605
rect 10920 2585 10930 2605
rect 10890 2555 10930 2585
rect 10890 2535 10900 2555
rect 10920 2535 10930 2555
rect 10890 2520 10930 2535
rect 11220 2610 11230 2630
rect 11250 2610 11260 2630
rect 11220 2580 11260 2610
rect 11220 2560 11230 2580
rect 11250 2560 11260 2580
rect 11220 2530 11260 2560
rect 11220 2510 11230 2530
rect 11250 2510 11260 2530
rect 11220 2495 11260 2510
rect 11280 2880 11320 2895
rect 11280 2860 11290 2880
rect 11310 2860 11320 2880
rect 11280 2830 11320 2860
rect 11280 2810 11290 2830
rect 11310 2810 11320 2830
rect 11280 2780 11320 2810
rect 11280 2760 11290 2780
rect 11310 2760 11320 2780
rect 11280 2730 11320 2760
rect 11280 2710 11290 2730
rect 11310 2710 11320 2730
rect 11280 2680 11320 2710
rect 11280 2660 11290 2680
rect 11310 2660 11320 2680
rect 11280 2630 11320 2660
rect 11280 2610 11290 2630
rect 11310 2610 11320 2630
rect 11280 2580 11320 2610
rect 11280 2560 11290 2580
rect 11310 2560 11320 2580
rect 11280 2530 11320 2560
rect 11280 2510 11290 2530
rect 11310 2510 11320 2530
rect 11280 2495 11320 2510
rect 11340 2880 11380 2895
rect 11340 2860 11350 2880
rect 11370 2860 11380 2880
rect 11340 2830 11380 2860
rect 11340 2810 11350 2830
rect 11370 2810 11380 2830
rect 11340 2780 11380 2810
rect 11340 2760 11350 2780
rect 11370 2760 11380 2780
rect 11340 2730 11380 2760
rect 11340 2710 11350 2730
rect 11370 2710 11380 2730
rect 11340 2680 11380 2710
rect 11340 2660 11350 2680
rect 11370 2660 11380 2680
rect 11340 2630 11380 2660
rect 11340 2610 11350 2630
rect 11370 2610 11380 2630
rect 11340 2580 11380 2610
rect 11340 2560 11350 2580
rect 11370 2560 11380 2580
rect 11340 2530 11380 2560
rect 11340 2510 11350 2530
rect 11370 2510 11380 2530
rect 11340 2495 11380 2510
rect 11400 2880 11440 2895
rect 11400 2860 11410 2880
rect 11430 2860 11440 2880
rect 11400 2830 11440 2860
rect 11400 2810 11410 2830
rect 11430 2810 11440 2830
rect 11400 2780 11440 2810
rect 11400 2760 11410 2780
rect 11430 2760 11440 2780
rect 11400 2730 11440 2760
rect 11400 2710 11410 2730
rect 11430 2710 11440 2730
rect 11400 2680 11440 2710
rect 11400 2660 11410 2680
rect 11430 2660 11440 2680
rect 11400 2630 11440 2660
rect 11400 2610 11410 2630
rect 11430 2610 11440 2630
rect 11400 2580 11440 2610
rect 11400 2560 11410 2580
rect 11430 2560 11440 2580
rect 11400 2530 11440 2560
rect 11400 2510 11410 2530
rect 11430 2510 11440 2530
rect 11400 2495 11440 2510
rect 11460 2880 11500 2895
rect 11460 2860 11470 2880
rect 11490 2860 11500 2880
rect 11460 2830 11500 2860
rect 11460 2810 11470 2830
rect 11490 2810 11500 2830
rect 11460 2780 11500 2810
rect 11460 2760 11470 2780
rect 11490 2760 11500 2780
rect 11460 2730 11500 2760
rect 11460 2710 11470 2730
rect 11490 2710 11500 2730
rect 11460 2680 11500 2710
rect 11460 2660 11470 2680
rect 11490 2660 11500 2680
rect 11460 2630 11500 2660
rect 11460 2610 11470 2630
rect 11490 2610 11500 2630
rect 11460 2580 11500 2610
rect 11460 2560 11470 2580
rect 11490 2560 11500 2580
rect 11460 2530 11500 2560
rect 11460 2510 11470 2530
rect 11490 2510 11500 2530
rect 11460 2495 11500 2510
rect 11520 2880 11560 2895
rect 11520 2860 11530 2880
rect 11550 2860 11560 2880
rect 11520 2830 11560 2860
rect 11520 2810 11530 2830
rect 11550 2810 11560 2830
rect 11520 2780 11560 2810
rect 11520 2760 11530 2780
rect 11550 2760 11560 2780
rect 11520 2730 11560 2760
rect 11520 2710 11530 2730
rect 11550 2710 11560 2730
rect 11520 2680 11560 2710
rect 11520 2660 11530 2680
rect 11550 2660 11560 2680
rect 11520 2630 11560 2660
rect 11520 2610 11530 2630
rect 11550 2610 11560 2630
rect 11520 2580 11560 2610
rect 11520 2560 11530 2580
rect 11550 2560 11560 2580
rect 11520 2530 11560 2560
rect 11520 2510 11530 2530
rect 11550 2510 11560 2530
rect 11520 2495 11560 2510
rect 11580 2880 11620 2895
rect 11580 2860 11590 2880
rect 11610 2860 11620 2880
rect 11580 2830 11620 2860
rect 11580 2810 11590 2830
rect 11610 2810 11620 2830
rect 11580 2780 11620 2810
rect 11580 2760 11590 2780
rect 11610 2760 11620 2780
rect 11580 2730 11620 2760
rect 11580 2710 11590 2730
rect 11610 2710 11620 2730
rect 11580 2680 11620 2710
rect 11580 2660 11590 2680
rect 11610 2660 11620 2680
rect 11580 2630 11620 2660
rect 11580 2610 11590 2630
rect 11610 2610 11620 2630
rect 11580 2580 11620 2610
rect 11580 2560 11590 2580
rect 11610 2560 11620 2580
rect 11580 2530 11620 2560
rect 11580 2510 11590 2530
rect 11610 2510 11620 2530
rect 11580 2495 11620 2510
rect 11640 2880 11680 2895
rect 11640 2860 11650 2880
rect 11670 2860 11680 2880
rect 11640 2830 11680 2860
rect 11640 2810 11650 2830
rect 11670 2810 11680 2830
rect 11640 2780 11680 2810
rect 11640 2760 11650 2780
rect 11670 2760 11680 2780
rect 11640 2730 11680 2760
rect 11640 2710 11650 2730
rect 11670 2710 11680 2730
rect 11640 2680 11680 2710
rect 11640 2660 11650 2680
rect 11670 2660 11680 2680
rect 11640 2630 11680 2660
rect 11640 2610 11650 2630
rect 11670 2610 11680 2630
rect 11640 2580 11680 2610
rect 11640 2560 11650 2580
rect 11670 2560 11680 2580
rect 11640 2530 11680 2560
rect 11640 2510 11650 2530
rect 11670 2510 11680 2530
rect 11640 2495 11680 2510
rect 11700 2880 11740 2895
rect 11700 2860 11710 2880
rect 11730 2860 11740 2880
rect 11700 2830 11740 2860
rect 11700 2810 11710 2830
rect 11730 2810 11740 2830
rect 11700 2780 11740 2810
rect 11700 2760 11710 2780
rect 11730 2760 11740 2780
rect 11700 2730 11740 2760
rect 11700 2710 11710 2730
rect 11730 2710 11740 2730
rect 11700 2680 11740 2710
rect 11700 2660 11710 2680
rect 11730 2660 11740 2680
rect 11700 2630 11740 2660
rect 11700 2610 11710 2630
rect 11730 2610 11740 2630
rect 11700 2580 11740 2610
rect 11700 2560 11710 2580
rect 11730 2560 11740 2580
rect 11700 2530 11740 2560
rect 11700 2510 11710 2530
rect 11730 2510 11740 2530
rect 11700 2495 11740 2510
rect 11760 2880 11800 2895
rect 11760 2860 11770 2880
rect 11790 2860 11800 2880
rect 11760 2830 11800 2860
rect 11760 2810 11770 2830
rect 11790 2810 11800 2830
rect 11760 2780 11800 2810
rect 11760 2760 11770 2780
rect 11790 2760 11800 2780
rect 11760 2730 11800 2760
rect 11760 2710 11770 2730
rect 11790 2710 11800 2730
rect 11760 2680 11800 2710
rect 11760 2660 11770 2680
rect 11790 2660 11800 2680
rect 11760 2630 11800 2660
rect 11760 2610 11770 2630
rect 11790 2610 11800 2630
rect 11760 2580 11800 2610
rect 11760 2560 11770 2580
rect 11790 2560 11800 2580
rect 11760 2530 11800 2560
rect 11760 2510 11770 2530
rect 11790 2510 11800 2530
rect 11760 2495 11800 2510
rect 11820 2880 11860 2895
rect 11820 2860 11830 2880
rect 11850 2860 11860 2880
rect 11820 2830 11860 2860
rect 11820 2810 11830 2830
rect 11850 2810 11860 2830
rect 11820 2780 11860 2810
rect 11820 2760 11830 2780
rect 11850 2760 11860 2780
rect 11820 2730 11860 2760
rect 11820 2710 11830 2730
rect 11850 2710 11860 2730
rect 11820 2680 11860 2710
rect 11820 2660 11830 2680
rect 11850 2660 11860 2680
rect 11820 2630 11860 2660
rect 11820 2610 11830 2630
rect 11850 2610 11860 2630
rect 11820 2580 11860 2610
rect 11820 2560 11830 2580
rect 11850 2560 11860 2580
rect 11820 2530 11860 2560
rect 11820 2510 11830 2530
rect 11850 2510 11860 2530
rect 11820 2495 11860 2510
rect 11880 2880 11920 2895
rect 11880 2860 11890 2880
rect 11910 2860 11920 2880
rect 11880 2830 11920 2860
rect 11880 2810 11890 2830
rect 11910 2810 11920 2830
rect 11880 2780 11920 2810
rect 11880 2760 11890 2780
rect 11910 2760 11920 2780
rect 11880 2730 11920 2760
rect 11880 2710 11890 2730
rect 11910 2710 11920 2730
rect 11880 2680 11920 2710
rect 11880 2660 11890 2680
rect 11910 2660 11920 2680
rect 11880 2630 11920 2660
rect 11880 2610 11890 2630
rect 11910 2610 11920 2630
rect 11880 2580 11920 2610
rect 11880 2560 11890 2580
rect 11910 2560 11920 2580
rect 11880 2530 11920 2560
rect 11880 2510 11890 2530
rect 11910 2510 11920 2530
rect 11880 2495 11920 2510
rect 11940 2880 11980 2895
rect 11940 2860 11950 2880
rect 11970 2860 11980 2880
rect 11940 2830 11980 2860
rect 11940 2810 11950 2830
rect 11970 2810 11980 2830
rect 11940 2780 11980 2810
rect 11940 2760 11950 2780
rect 11970 2760 11980 2780
rect 11940 2730 11980 2760
rect 11940 2710 11950 2730
rect 11970 2710 11980 2730
rect 11940 2680 11980 2710
rect 11940 2660 11950 2680
rect 11970 2660 11980 2680
rect 11940 2630 11980 2660
rect 11940 2610 11950 2630
rect 11970 2610 11980 2630
rect 11940 2580 11980 2610
rect 11940 2560 11950 2580
rect 11970 2560 11980 2580
rect 11940 2530 11980 2560
rect 11940 2510 11950 2530
rect 11970 2510 11980 2530
rect 11940 2495 11980 2510
rect 12000 2880 12040 2895
rect 12000 2860 12010 2880
rect 12030 2860 12040 2880
rect 12000 2830 12040 2860
rect 12000 2810 12010 2830
rect 12030 2810 12040 2830
rect 12000 2780 12040 2810
rect 12000 2760 12010 2780
rect 12030 2760 12040 2780
rect 12000 2730 12040 2760
rect 12000 2710 12010 2730
rect 12030 2710 12040 2730
rect 12000 2680 12040 2710
rect 12000 2660 12010 2680
rect 12030 2660 12040 2680
rect 12000 2630 12040 2660
rect 12000 2610 12010 2630
rect 12030 2610 12040 2630
rect 12000 2580 12040 2610
rect 12000 2560 12010 2580
rect 12030 2560 12040 2580
rect 12000 2530 12040 2560
rect 12000 2510 12010 2530
rect 12030 2510 12040 2530
rect 12000 2495 12040 2510
rect 12060 2880 12100 2895
rect 12060 2860 12070 2880
rect 12090 2860 12100 2880
rect 12060 2830 12100 2860
rect 12060 2810 12070 2830
rect 12090 2810 12100 2830
rect 12060 2780 12100 2810
rect 12060 2760 12070 2780
rect 12090 2760 12100 2780
rect 12060 2730 12100 2760
rect 12060 2710 12070 2730
rect 12090 2710 12100 2730
rect 12060 2680 12100 2710
rect 12060 2660 12070 2680
rect 12090 2660 12100 2680
rect 12060 2630 12100 2660
rect 12060 2610 12070 2630
rect 12090 2610 12100 2630
rect 12060 2580 12100 2610
rect 12060 2560 12070 2580
rect 12090 2560 12100 2580
rect 12060 2530 12100 2560
rect 12060 2510 12070 2530
rect 12090 2510 12100 2530
rect 12060 2495 12100 2510
rect 12120 2880 12160 2895
rect 12120 2860 12130 2880
rect 12150 2860 12160 2880
rect 12120 2830 12160 2860
rect 12120 2810 12130 2830
rect 12150 2810 12160 2830
rect 12120 2780 12160 2810
rect 12120 2760 12130 2780
rect 12150 2760 12160 2780
rect 12120 2730 12160 2760
rect 12120 2710 12130 2730
rect 12150 2710 12160 2730
rect 12120 2680 12160 2710
rect 12120 2660 12130 2680
rect 12150 2660 12160 2680
rect 12120 2630 12160 2660
rect 12120 2610 12130 2630
rect 12150 2610 12160 2630
rect 12120 2580 12160 2610
rect 12120 2560 12130 2580
rect 12150 2560 12160 2580
rect 12120 2530 12160 2560
rect 12120 2510 12130 2530
rect 12150 2510 12160 2530
rect 12120 2495 12160 2510
rect 12180 2880 12220 2895
rect 12180 2860 12190 2880
rect 12210 2860 12220 2880
rect 12180 2830 12220 2860
rect 12180 2810 12190 2830
rect 12210 2810 12220 2830
rect 12180 2780 12220 2810
rect 12180 2760 12190 2780
rect 12210 2760 12220 2780
rect 12180 2730 12220 2760
rect 12180 2710 12190 2730
rect 12210 2710 12220 2730
rect 12180 2680 12220 2710
rect 12180 2660 12190 2680
rect 12210 2660 12220 2680
rect 12180 2630 12220 2660
rect 12180 2610 12190 2630
rect 12210 2610 12220 2630
rect 12180 2580 12220 2610
rect 12180 2560 12190 2580
rect 12210 2560 12220 2580
rect 12180 2530 12220 2560
rect 12180 2510 12190 2530
rect 12210 2510 12220 2530
rect 12180 2495 12220 2510
rect 12240 2880 12280 2895
rect 12240 2860 12250 2880
rect 12270 2860 12280 2880
rect 12240 2830 12280 2860
rect 12240 2810 12250 2830
rect 12270 2810 12280 2830
rect 12240 2780 12280 2810
rect 12240 2760 12250 2780
rect 12270 2760 12280 2780
rect 12240 2730 12280 2760
rect 12240 2710 12250 2730
rect 12270 2710 12280 2730
rect 12240 2680 12280 2710
rect 12240 2660 12250 2680
rect 12270 2660 12280 2680
rect 12240 2630 12280 2660
rect 12240 2610 12250 2630
rect 12270 2610 12280 2630
rect 12240 2580 12280 2610
rect 12240 2560 12250 2580
rect 12270 2560 12280 2580
rect 12240 2530 12280 2560
rect 12240 2510 12250 2530
rect 12270 2510 12280 2530
rect 12240 2495 12280 2510
rect 12300 2880 12340 2895
rect 12300 2860 12310 2880
rect 12330 2860 12340 2880
rect 12300 2830 12340 2860
rect 12300 2810 12310 2830
rect 12330 2810 12340 2830
rect 12300 2780 12340 2810
rect 12300 2760 12310 2780
rect 12330 2760 12340 2780
rect 12300 2730 12340 2760
rect 12300 2710 12310 2730
rect 12330 2710 12340 2730
rect 12300 2680 12340 2710
rect 12300 2660 12310 2680
rect 12330 2660 12340 2680
rect 12300 2630 12340 2660
rect 12300 2610 12310 2630
rect 12330 2610 12340 2630
rect 12300 2580 12340 2610
rect 12300 2560 12310 2580
rect 12330 2560 12340 2580
rect 12300 2530 12340 2560
rect 12300 2510 12310 2530
rect 12330 2510 12340 2530
rect 12300 2495 12340 2510
rect 12360 2880 12400 2895
rect 12360 2860 12370 2880
rect 12390 2860 12400 2880
rect 12360 2830 12400 2860
rect 12360 2810 12370 2830
rect 12390 2810 12400 2830
rect 12360 2780 12400 2810
rect 12360 2760 12370 2780
rect 12390 2760 12400 2780
rect 12360 2730 12400 2760
rect 12360 2710 12370 2730
rect 12390 2710 12400 2730
rect 12360 2680 12400 2710
rect 12360 2660 12370 2680
rect 12390 2660 12400 2680
rect 12360 2630 12400 2660
rect 12360 2610 12370 2630
rect 12390 2610 12400 2630
rect 12360 2580 12400 2610
rect 12360 2560 12370 2580
rect 12390 2560 12400 2580
rect 12360 2530 12400 2560
rect 12360 2510 12370 2530
rect 12390 2510 12400 2530
rect 12360 2495 12400 2510
rect 12420 2880 12460 2895
rect 12420 2860 12430 2880
rect 12450 2860 12460 2880
rect 12420 2830 12460 2860
rect 12420 2810 12430 2830
rect 12450 2810 12460 2830
rect 12420 2780 12460 2810
rect 12420 2760 12430 2780
rect 12450 2760 12460 2780
rect 12420 2730 12460 2760
rect 12420 2710 12430 2730
rect 12450 2710 12460 2730
rect 12420 2680 12460 2710
rect 12420 2660 12430 2680
rect 12450 2660 12460 2680
rect 12420 2630 12460 2660
rect 12420 2610 12430 2630
rect 12450 2610 12460 2630
rect 12420 2580 12460 2610
rect 12420 2560 12430 2580
rect 12450 2560 12460 2580
rect 12420 2530 12460 2560
rect 12420 2510 12430 2530
rect 12450 2510 12460 2530
rect 12420 2495 12460 2510
rect 12480 2880 12520 2895
rect 12480 2860 12490 2880
rect 12510 2860 12520 2880
rect 12480 2830 12520 2860
rect 12480 2810 12490 2830
rect 12510 2810 12520 2830
rect 12480 2780 12520 2810
rect 12480 2760 12490 2780
rect 12510 2760 12520 2780
rect 12480 2730 12520 2760
rect 12480 2710 12490 2730
rect 12510 2710 12520 2730
rect 12480 2680 12520 2710
rect 12480 2660 12490 2680
rect 12510 2660 12520 2680
rect 12480 2630 12520 2660
rect 12480 2610 12490 2630
rect 12510 2610 12520 2630
rect 12480 2580 12520 2610
rect 12480 2560 12490 2580
rect 12510 2560 12520 2580
rect 12480 2530 12520 2560
rect 12480 2510 12490 2530
rect 12510 2510 12520 2530
rect 12480 2495 12520 2510
rect 12540 2880 12580 2895
rect 20390 2940 20430 2955
rect 20445 3225 20485 3240
rect 20445 3205 20455 3225
rect 20475 3205 20485 3225
rect 20445 3175 20485 3205
rect 20445 3155 20455 3175
rect 20475 3155 20485 3175
rect 20445 3125 20485 3155
rect 20445 3105 20455 3125
rect 20475 3105 20485 3125
rect 20445 3075 20485 3105
rect 20445 3055 20455 3075
rect 20475 3055 20485 3075
rect 20445 3025 20485 3055
rect 20445 3005 20455 3025
rect 20475 3005 20485 3025
rect 20445 2975 20485 3005
rect 20445 2955 20455 2975
rect 20475 2955 20485 2975
rect 20445 2940 20485 2955
rect 20500 3225 20540 3240
rect 20500 3205 20510 3225
rect 20530 3205 20540 3225
rect 20500 3175 20540 3205
rect 20500 3155 20510 3175
rect 20530 3155 20540 3175
rect 20500 3125 20540 3155
rect 20500 3105 20510 3125
rect 20530 3105 20540 3125
rect 20500 3075 20540 3105
rect 20500 3055 20510 3075
rect 20530 3055 20540 3075
rect 20500 3025 20540 3055
rect 20500 3005 20510 3025
rect 20530 3005 20540 3025
rect 20500 2975 20540 3005
rect 20500 2955 20510 2975
rect 20530 2955 20540 2975
rect 20500 2940 20540 2955
rect 20555 3225 20595 3240
rect 20555 3205 20565 3225
rect 20585 3205 20595 3225
rect 20555 3175 20595 3205
rect 20555 3155 20565 3175
rect 20585 3155 20595 3175
rect 20555 3125 20595 3155
rect 20555 3105 20565 3125
rect 20585 3105 20595 3125
rect 20555 3075 20595 3105
rect 20555 3055 20565 3075
rect 20585 3055 20595 3075
rect 20555 3025 20595 3055
rect 20555 3005 20565 3025
rect 20585 3005 20595 3025
rect 20555 2975 20595 3005
rect 20555 2955 20565 2975
rect 20585 2955 20595 2975
rect 20555 2940 20595 2955
rect 20610 3225 20650 3240
rect 20610 3205 20620 3225
rect 20640 3205 20650 3225
rect 20610 3175 20650 3205
rect 20610 3155 20620 3175
rect 20640 3155 20650 3175
rect 20610 3125 20650 3155
rect 20610 3105 20620 3125
rect 20640 3105 20650 3125
rect 20610 3075 20650 3105
rect 20610 3055 20620 3075
rect 20640 3055 20650 3075
rect 20610 3025 20650 3055
rect 20610 3005 20620 3025
rect 20640 3005 20650 3025
rect 20610 2975 20650 3005
rect 20610 2955 20620 2975
rect 20640 2955 20650 2975
rect 20610 2940 20650 2955
rect 20665 3225 20705 3240
rect 20665 3205 20675 3225
rect 20695 3205 20705 3225
rect 20665 3175 20705 3205
rect 20665 3155 20675 3175
rect 20695 3155 20705 3175
rect 20665 3125 20705 3155
rect 20665 3105 20675 3125
rect 20695 3105 20705 3125
rect 20665 3075 20705 3105
rect 20665 3055 20675 3075
rect 20695 3055 20705 3075
rect 20665 3025 20705 3055
rect 20665 3005 20675 3025
rect 20695 3005 20705 3025
rect 20665 2975 20705 3005
rect 20665 2955 20675 2975
rect 20695 2955 20705 2975
rect 20665 2940 20705 2955
rect 20720 3225 20760 3240
rect 20720 3205 20730 3225
rect 20750 3205 20760 3225
rect 20720 3175 20760 3205
rect 20720 3155 20730 3175
rect 20750 3155 20760 3175
rect 20720 3125 20760 3155
rect 20720 3105 20730 3125
rect 20750 3105 20760 3125
rect 20720 3075 20760 3105
rect 20720 3055 20730 3075
rect 20750 3055 20760 3075
rect 20720 3025 20760 3055
rect 20720 3005 20730 3025
rect 20750 3005 20760 3025
rect 20720 2975 20760 3005
rect 20720 2955 20730 2975
rect 20750 2955 20760 2975
rect 20720 2940 20760 2955
rect 20775 3225 20815 3240
rect 20775 3205 20785 3225
rect 20805 3205 20815 3225
rect 20775 3175 20815 3205
rect 20775 3155 20785 3175
rect 20805 3155 20815 3175
rect 20775 3125 20815 3155
rect 20775 3105 20785 3125
rect 20805 3105 20815 3125
rect 20775 3075 20815 3105
rect 20775 3055 20785 3075
rect 20805 3055 20815 3075
rect 20775 3025 20815 3055
rect 20775 3005 20785 3025
rect 20805 3005 20815 3025
rect 20775 2975 20815 3005
rect 20775 2955 20785 2975
rect 20805 2955 20815 2975
rect 20775 2940 20815 2955
rect 20830 3225 20870 3240
rect 20830 3205 20840 3225
rect 20860 3205 20870 3225
rect 20830 3175 20870 3205
rect 20830 3155 20840 3175
rect 20860 3155 20870 3175
rect 20830 3125 20870 3155
rect 20830 3105 20840 3125
rect 20860 3105 20870 3125
rect 20830 3075 20870 3105
rect 20830 3055 20840 3075
rect 20860 3055 20870 3075
rect 20830 3025 20870 3055
rect 20830 3005 20840 3025
rect 20860 3005 20870 3025
rect 20830 2975 20870 3005
rect 20830 2955 20840 2975
rect 20860 2955 20870 2975
rect 20830 2940 20870 2955
rect 20885 3225 20925 3240
rect 20885 3205 20895 3225
rect 20915 3205 20925 3225
rect 20885 3175 20925 3205
rect 20885 3155 20895 3175
rect 20915 3155 20925 3175
rect 20885 3125 20925 3155
rect 20885 3105 20895 3125
rect 20915 3105 20925 3125
rect 20885 3075 20925 3105
rect 20885 3055 20895 3075
rect 20915 3055 20925 3075
rect 20885 3025 20925 3055
rect 20885 3005 20895 3025
rect 20915 3005 20925 3025
rect 20885 2975 20925 3005
rect 20885 2955 20895 2975
rect 20915 2955 20925 2975
rect 20885 2940 20925 2955
rect 20940 3225 20980 3240
rect 20940 3205 20950 3225
rect 20970 3205 20980 3225
rect 20940 3175 20980 3205
rect 20940 3155 20950 3175
rect 20970 3155 20980 3175
rect 20940 3125 20980 3155
rect 20940 3105 20950 3125
rect 20970 3105 20980 3125
rect 20940 3075 20980 3105
rect 20940 3055 20950 3075
rect 20970 3055 20980 3075
rect 20940 3025 20980 3055
rect 20940 3005 20950 3025
rect 20970 3005 20980 3025
rect 20940 2975 20980 3005
rect 20940 2955 20950 2975
rect 20970 2955 20980 2975
rect 20940 2940 20980 2955
rect 20995 3225 21035 3240
rect 20995 3205 21005 3225
rect 21025 3205 21035 3225
rect 20995 3175 21035 3205
rect 20995 3155 21005 3175
rect 21025 3155 21035 3175
rect 20995 3125 21035 3155
rect 20995 3105 21005 3125
rect 21025 3105 21035 3125
rect 20995 3075 21035 3105
rect 20995 3055 21005 3075
rect 21025 3055 21035 3075
rect 20995 3025 21035 3055
rect 20995 3005 21005 3025
rect 21025 3005 21035 3025
rect 20995 2975 21035 3005
rect 20995 2955 21005 2975
rect 21025 2955 21035 2975
rect 20995 2940 21035 2955
rect 21050 3225 21090 3240
rect 21050 3205 21060 3225
rect 21080 3205 21090 3225
rect 21050 3175 21090 3205
rect 21050 3155 21060 3175
rect 21080 3155 21090 3175
rect 21050 3125 21090 3155
rect 21050 3105 21060 3125
rect 21080 3105 21090 3125
rect 21050 3075 21090 3105
rect 21050 3055 21060 3075
rect 21080 3055 21090 3075
rect 21050 3025 21090 3055
rect 21050 3005 21060 3025
rect 21080 3005 21090 3025
rect 21050 2975 21090 3005
rect 21050 2955 21060 2975
rect 21080 2955 21090 2975
rect 21050 2940 21090 2955
rect 21105 3225 21145 3240
rect 21105 3205 21115 3225
rect 21135 3205 21145 3225
rect 21105 3175 21145 3205
rect 21105 3155 21115 3175
rect 21135 3155 21145 3175
rect 21105 3125 21145 3155
rect 21105 3105 21115 3125
rect 21135 3105 21145 3125
rect 21105 3075 21145 3105
rect 21105 3055 21115 3075
rect 21135 3055 21145 3075
rect 21105 3025 21145 3055
rect 21105 3005 21115 3025
rect 21135 3005 21145 3025
rect 21105 2975 21145 3005
rect 21105 2955 21115 2975
rect 21135 2955 21145 2975
rect 21105 2940 21145 2955
rect 21160 3225 21200 3240
rect 21160 3205 21170 3225
rect 21190 3205 21200 3225
rect 21160 3175 21200 3205
rect 21160 3155 21170 3175
rect 21190 3155 21200 3175
rect 21160 3125 21200 3155
rect 21160 3105 21170 3125
rect 21190 3105 21200 3125
rect 21160 3075 21200 3105
rect 21160 3055 21170 3075
rect 21190 3055 21200 3075
rect 21160 3025 21200 3055
rect 21160 3005 21170 3025
rect 21190 3005 21200 3025
rect 21160 2975 21200 3005
rect 21160 2955 21170 2975
rect 21190 2955 21200 2975
rect 21160 2940 21200 2955
rect 21215 3225 21255 3240
rect 21215 3205 21225 3225
rect 21245 3205 21255 3225
rect 21215 3175 21255 3205
rect 21215 3155 21225 3175
rect 21245 3155 21255 3175
rect 21215 3125 21255 3155
rect 21215 3105 21225 3125
rect 21245 3105 21255 3125
rect 21215 3075 21255 3105
rect 21215 3055 21225 3075
rect 21245 3055 21255 3075
rect 21215 3025 21255 3055
rect 21215 3005 21225 3025
rect 21245 3005 21255 3025
rect 21215 2975 21255 3005
rect 21215 2955 21225 2975
rect 21245 2955 21255 2975
rect 21215 2940 21255 2955
rect 21270 3225 21310 3240
rect 21270 3205 21280 3225
rect 21300 3205 21310 3225
rect 21270 3175 21310 3205
rect 21270 3155 21280 3175
rect 21300 3155 21310 3175
rect 21270 3125 21310 3155
rect 21270 3105 21280 3125
rect 21300 3105 21310 3125
rect 21270 3075 21310 3105
rect 21270 3055 21280 3075
rect 21300 3055 21310 3075
rect 21270 3025 21310 3055
rect 21270 3005 21280 3025
rect 21300 3005 21310 3025
rect 21270 2975 21310 3005
rect 21270 2955 21280 2975
rect 21300 2955 21310 2975
rect 21270 2940 21310 2955
rect 21325 3225 21365 3240
rect 21325 3205 21335 3225
rect 21355 3205 21365 3225
rect 21325 3175 21365 3205
rect 21325 3155 21335 3175
rect 21355 3155 21365 3175
rect 21325 3125 21365 3155
rect 21325 3105 21335 3125
rect 21355 3105 21365 3125
rect 21325 3075 21365 3105
rect 21325 3055 21335 3075
rect 21355 3055 21365 3075
rect 21325 3025 21365 3055
rect 21325 3005 21335 3025
rect 21355 3005 21365 3025
rect 21325 2975 21365 3005
rect 21325 2955 21335 2975
rect 21355 2955 21365 2975
rect 21325 2940 21365 2955
rect 21380 3225 21420 3240
rect 21380 3205 21390 3225
rect 21410 3205 21420 3225
rect 21380 3175 21420 3205
rect 21380 3155 21390 3175
rect 21410 3155 21420 3175
rect 21380 3125 21420 3155
rect 21380 3105 21390 3125
rect 21410 3105 21420 3125
rect 21380 3075 21420 3105
rect 21380 3055 21390 3075
rect 21410 3055 21420 3075
rect 21380 3025 21420 3055
rect 21380 3005 21390 3025
rect 21410 3005 21420 3025
rect 21380 2975 21420 3005
rect 21380 2955 21390 2975
rect 21410 2955 21420 2975
rect 21380 2940 21420 2955
rect 21435 3225 21475 3240
rect 21435 3205 21445 3225
rect 21465 3205 21475 3225
rect 21435 3175 21475 3205
rect 21435 3155 21445 3175
rect 21465 3155 21475 3175
rect 21435 3125 21475 3155
rect 21435 3105 21445 3125
rect 21465 3105 21475 3125
rect 21435 3075 21475 3105
rect 21435 3055 21445 3075
rect 21465 3055 21475 3075
rect 21435 3025 21475 3055
rect 21435 3005 21445 3025
rect 21465 3005 21475 3025
rect 21435 2975 21475 3005
rect 21435 2955 21445 2975
rect 21465 2955 21475 2975
rect 21435 2940 21475 2955
rect 21490 3225 21530 3240
rect 21490 3205 21500 3225
rect 21520 3205 21530 3225
rect 21490 3175 21530 3205
rect 21490 3155 21500 3175
rect 21520 3155 21530 3175
rect 21490 3125 21530 3155
rect 21490 3105 21500 3125
rect 21520 3105 21530 3125
rect 21490 3075 21530 3105
rect 21490 3055 21500 3075
rect 21520 3055 21530 3075
rect 21490 3025 21530 3055
rect 21490 3005 21500 3025
rect 21520 3005 21530 3025
rect 21490 2975 21530 3005
rect 21490 2955 21500 2975
rect 21520 2955 21530 2975
rect 21490 2940 21530 2955
rect 21545 3225 21585 3240
rect 21545 3205 21555 3225
rect 21575 3205 21585 3225
rect 21545 3175 21585 3205
rect 21545 3155 21555 3175
rect 21575 3155 21585 3175
rect 21545 3125 21585 3155
rect 21545 3105 21555 3125
rect 21575 3105 21585 3125
rect 21545 3075 21585 3105
rect 21545 3055 21555 3075
rect 21575 3055 21585 3075
rect 21545 3025 21585 3055
rect 21545 3005 21555 3025
rect 21575 3005 21585 3025
rect 21545 2975 21585 3005
rect 21545 2955 21555 2975
rect 21575 2955 21585 2975
rect 21545 2940 21585 2955
rect 21600 3225 21640 3240
rect 21600 3205 21610 3225
rect 21630 3205 21640 3225
rect 21600 3175 21640 3205
rect 21600 3155 21610 3175
rect 21630 3155 21640 3175
rect 21600 3125 21640 3155
rect 21600 3105 21610 3125
rect 21630 3105 21640 3125
rect 21600 3075 21640 3105
rect 21600 3055 21610 3075
rect 21630 3055 21640 3075
rect 21600 3025 21640 3055
rect 21600 3005 21610 3025
rect 21630 3005 21640 3025
rect 21600 2975 21640 3005
rect 21600 2955 21610 2975
rect 21630 2955 21640 2975
rect 21600 2940 21640 2955
rect 12540 2860 12550 2880
rect 12570 2860 12580 2880
rect 12540 2830 12580 2860
rect 18720 2880 18760 2895
rect 18720 2860 18730 2880
rect 18750 2860 18760 2880
rect 12540 2810 12550 2830
rect 12570 2810 12580 2830
rect 12540 2780 12580 2810
rect 12540 2760 12550 2780
rect 12570 2760 12580 2780
rect 12540 2730 12580 2760
rect 12540 2710 12550 2730
rect 12570 2710 12580 2730
rect 12540 2680 12580 2710
rect 18720 2830 18760 2860
rect 18720 2810 18730 2830
rect 18750 2810 18760 2830
rect 18720 2780 18760 2810
rect 18720 2760 18730 2780
rect 18750 2760 18760 2780
rect 18720 2730 18760 2760
rect 18720 2710 18730 2730
rect 18750 2710 18760 2730
rect 12540 2660 12550 2680
rect 12570 2660 12580 2680
rect 12540 2630 12580 2660
rect 18720 2680 18760 2710
rect 18720 2660 18730 2680
rect 18750 2660 18760 2680
rect 12540 2610 12550 2630
rect 12570 2610 12580 2630
rect 18720 2630 18760 2660
rect 12540 2580 12580 2610
rect 12540 2560 12550 2580
rect 12570 2560 12580 2580
rect 12540 2530 12580 2560
rect 12540 2510 12550 2530
rect 12570 2510 12580 2530
rect 12890 2605 12930 2620
rect 12890 2585 12900 2605
rect 12920 2585 12930 2605
rect 12890 2555 12930 2585
rect 12890 2535 12900 2555
rect 12920 2535 12930 2555
rect 12890 2520 12930 2535
rect 12945 2605 12985 2620
rect 12945 2585 12955 2605
rect 12975 2585 12985 2605
rect 12945 2555 12985 2585
rect 12945 2535 12955 2555
rect 12975 2535 12985 2555
rect 12945 2520 12985 2535
rect 13000 2605 13040 2620
rect 13000 2585 13010 2605
rect 13030 2585 13040 2605
rect 13000 2555 13040 2585
rect 13000 2535 13010 2555
rect 13030 2535 13040 2555
rect 13000 2520 13040 2535
rect 13055 2605 13095 2620
rect 13055 2585 13065 2605
rect 13085 2585 13095 2605
rect 13055 2555 13095 2585
rect 13055 2535 13065 2555
rect 13085 2535 13095 2555
rect 13055 2520 13095 2535
rect 13110 2605 13150 2620
rect 13110 2585 13120 2605
rect 13140 2585 13150 2605
rect 13110 2555 13150 2585
rect 13110 2535 13120 2555
rect 13140 2535 13150 2555
rect 13110 2520 13150 2535
rect 13165 2605 13205 2620
rect 13165 2585 13175 2605
rect 13195 2585 13205 2605
rect 13165 2555 13205 2585
rect 13165 2535 13175 2555
rect 13195 2535 13205 2555
rect 13165 2520 13205 2535
rect 13220 2605 13260 2620
rect 13220 2585 13230 2605
rect 13250 2585 13260 2605
rect 13220 2555 13260 2585
rect 13220 2535 13230 2555
rect 13250 2535 13260 2555
rect 13220 2520 13260 2535
rect 13275 2605 13315 2620
rect 13275 2585 13285 2605
rect 13305 2585 13315 2605
rect 13275 2555 13315 2585
rect 13275 2535 13285 2555
rect 13305 2535 13315 2555
rect 13275 2520 13315 2535
rect 13330 2605 13370 2620
rect 13330 2585 13340 2605
rect 13360 2585 13370 2605
rect 13330 2555 13370 2585
rect 13330 2535 13340 2555
rect 13360 2535 13370 2555
rect 13330 2520 13370 2535
rect 13385 2605 13425 2620
rect 13385 2585 13395 2605
rect 13415 2585 13425 2605
rect 13385 2555 13425 2585
rect 13385 2535 13395 2555
rect 13415 2535 13425 2555
rect 13385 2520 13425 2535
rect 13440 2605 13480 2620
rect 13440 2585 13450 2605
rect 13470 2585 13480 2605
rect 13440 2555 13480 2585
rect 13440 2535 13450 2555
rect 13470 2535 13480 2555
rect 13440 2520 13480 2535
rect 13495 2605 13535 2620
rect 13495 2585 13505 2605
rect 13525 2585 13535 2605
rect 13495 2555 13535 2585
rect 13495 2535 13505 2555
rect 13525 2535 13535 2555
rect 13495 2520 13535 2535
rect 13550 2605 13590 2620
rect 13550 2585 13560 2605
rect 13580 2585 13590 2605
rect 13550 2555 13590 2585
rect 13550 2535 13560 2555
rect 13580 2535 13590 2555
rect 13550 2520 13590 2535
rect 13605 2605 13645 2620
rect 13605 2585 13615 2605
rect 13635 2585 13645 2605
rect 13605 2555 13645 2585
rect 13605 2535 13615 2555
rect 13635 2535 13645 2555
rect 13605 2520 13645 2535
rect 13660 2605 13700 2620
rect 13660 2585 13670 2605
rect 13690 2585 13700 2605
rect 13660 2555 13700 2585
rect 13660 2535 13670 2555
rect 13690 2535 13700 2555
rect 13660 2520 13700 2535
rect 13715 2605 13755 2620
rect 13715 2585 13725 2605
rect 13745 2585 13755 2605
rect 13715 2555 13755 2585
rect 13715 2535 13725 2555
rect 13745 2535 13755 2555
rect 13715 2520 13755 2535
rect 13770 2605 13810 2620
rect 13770 2585 13780 2605
rect 13800 2585 13810 2605
rect 13770 2555 13810 2585
rect 13770 2535 13780 2555
rect 13800 2535 13810 2555
rect 13770 2520 13810 2535
rect 13825 2605 13865 2620
rect 13825 2585 13835 2605
rect 13855 2585 13865 2605
rect 13825 2555 13865 2585
rect 13825 2535 13835 2555
rect 13855 2535 13865 2555
rect 13825 2520 13865 2535
rect 13880 2605 13920 2620
rect 13880 2585 13890 2605
rect 13910 2585 13920 2605
rect 13880 2555 13920 2585
rect 13880 2535 13890 2555
rect 13910 2535 13920 2555
rect 13880 2520 13920 2535
rect 13935 2605 13975 2620
rect 13935 2585 13945 2605
rect 13965 2585 13975 2605
rect 13935 2555 13975 2585
rect 13935 2535 13945 2555
rect 13965 2535 13975 2555
rect 13935 2520 13975 2535
rect 13990 2605 14030 2620
rect 13990 2585 14000 2605
rect 14020 2585 14030 2605
rect 13990 2555 14030 2585
rect 13990 2535 14000 2555
rect 14020 2535 14030 2555
rect 13990 2520 14030 2535
rect 14045 2605 14085 2620
rect 14045 2585 14055 2605
rect 14075 2585 14085 2605
rect 14045 2555 14085 2585
rect 14045 2535 14055 2555
rect 14075 2535 14085 2555
rect 14045 2520 14085 2535
rect 14100 2605 14140 2620
rect 14100 2585 14110 2605
rect 14130 2585 14140 2605
rect 14100 2555 14140 2585
rect 14100 2535 14110 2555
rect 14130 2535 14140 2555
rect 14100 2520 14140 2535
rect 17180 2605 17220 2620
rect 17180 2585 17190 2605
rect 17210 2585 17220 2605
rect 17180 2555 17220 2585
rect 17180 2535 17190 2555
rect 17210 2535 17220 2555
rect 17180 2520 17220 2535
rect 17235 2605 17275 2620
rect 17235 2585 17245 2605
rect 17265 2585 17275 2605
rect 17235 2555 17275 2585
rect 17235 2535 17245 2555
rect 17265 2535 17275 2555
rect 17235 2520 17275 2535
rect 17290 2605 17330 2620
rect 17290 2585 17300 2605
rect 17320 2585 17330 2605
rect 17290 2555 17330 2585
rect 17290 2535 17300 2555
rect 17320 2535 17330 2555
rect 17290 2520 17330 2535
rect 17345 2605 17385 2620
rect 17345 2585 17355 2605
rect 17375 2585 17385 2605
rect 17345 2555 17385 2585
rect 17345 2535 17355 2555
rect 17375 2535 17385 2555
rect 17345 2520 17385 2535
rect 17400 2605 17440 2620
rect 17400 2585 17410 2605
rect 17430 2585 17440 2605
rect 17400 2555 17440 2585
rect 17400 2535 17410 2555
rect 17430 2535 17440 2555
rect 17400 2520 17440 2535
rect 17455 2605 17495 2620
rect 17455 2585 17465 2605
rect 17485 2585 17495 2605
rect 17455 2555 17495 2585
rect 17455 2535 17465 2555
rect 17485 2535 17495 2555
rect 17455 2520 17495 2535
rect 17510 2605 17550 2620
rect 17510 2585 17520 2605
rect 17540 2585 17550 2605
rect 17510 2555 17550 2585
rect 17510 2535 17520 2555
rect 17540 2535 17550 2555
rect 17510 2520 17550 2535
rect 17565 2605 17605 2620
rect 17565 2585 17575 2605
rect 17595 2585 17605 2605
rect 17565 2555 17605 2585
rect 17565 2535 17575 2555
rect 17595 2535 17605 2555
rect 17565 2520 17605 2535
rect 17620 2605 17660 2620
rect 17620 2585 17630 2605
rect 17650 2585 17660 2605
rect 17620 2555 17660 2585
rect 17620 2535 17630 2555
rect 17650 2535 17660 2555
rect 17620 2520 17660 2535
rect 17675 2605 17715 2620
rect 17675 2585 17685 2605
rect 17705 2585 17715 2605
rect 17675 2555 17715 2585
rect 17675 2535 17685 2555
rect 17705 2535 17715 2555
rect 17675 2520 17715 2535
rect 17730 2605 17770 2620
rect 17730 2585 17740 2605
rect 17760 2585 17770 2605
rect 17730 2555 17770 2585
rect 17730 2535 17740 2555
rect 17760 2535 17770 2555
rect 17730 2520 17770 2535
rect 17785 2605 17825 2620
rect 17785 2585 17795 2605
rect 17815 2585 17825 2605
rect 17785 2555 17825 2585
rect 17785 2535 17795 2555
rect 17815 2535 17825 2555
rect 17785 2520 17825 2535
rect 17840 2605 17880 2620
rect 17840 2585 17850 2605
rect 17870 2585 17880 2605
rect 17840 2555 17880 2585
rect 17840 2535 17850 2555
rect 17870 2535 17880 2555
rect 17840 2520 17880 2535
rect 17895 2605 17935 2620
rect 17895 2585 17905 2605
rect 17925 2585 17935 2605
rect 17895 2555 17935 2585
rect 17895 2535 17905 2555
rect 17925 2535 17935 2555
rect 17895 2520 17935 2535
rect 17950 2605 17990 2620
rect 17950 2585 17960 2605
rect 17980 2585 17990 2605
rect 17950 2555 17990 2585
rect 17950 2535 17960 2555
rect 17980 2535 17990 2555
rect 17950 2520 17990 2535
rect 18005 2605 18045 2620
rect 18005 2585 18015 2605
rect 18035 2585 18045 2605
rect 18005 2555 18045 2585
rect 18005 2535 18015 2555
rect 18035 2535 18045 2555
rect 18005 2520 18045 2535
rect 18060 2605 18100 2620
rect 18060 2585 18070 2605
rect 18090 2585 18100 2605
rect 18060 2555 18100 2585
rect 18060 2535 18070 2555
rect 18090 2535 18100 2555
rect 18060 2520 18100 2535
rect 18115 2605 18155 2620
rect 18115 2585 18125 2605
rect 18145 2585 18155 2605
rect 18115 2555 18155 2585
rect 18115 2535 18125 2555
rect 18145 2535 18155 2555
rect 18115 2520 18155 2535
rect 18170 2605 18210 2620
rect 18170 2585 18180 2605
rect 18200 2585 18210 2605
rect 18170 2555 18210 2585
rect 18170 2535 18180 2555
rect 18200 2535 18210 2555
rect 18170 2520 18210 2535
rect 18225 2605 18265 2620
rect 18225 2585 18235 2605
rect 18255 2585 18265 2605
rect 18225 2555 18265 2585
rect 18225 2535 18235 2555
rect 18255 2535 18265 2555
rect 18225 2520 18265 2535
rect 18280 2605 18320 2620
rect 18280 2585 18290 2605
rect 18310 2585 18320 2605
rect 18280 2555 18320 2585
rect 18280 2535 18290 2555
rect 18310 2535 18320 2555
rect 18280 2520 18320 2535
rect 18335 2605 18375 2620
rect 18335 2585 18345 2605
rect 18365 2585 18375 2605
rect 18335 2555 18375 2585
rect 18335 2535 18345 2555
rect 18365 2535 18375 2555
rect 18335 2520 18375 2535
rect 18390 2605 18430 2620
rect 18390 2585 18400 2605
rect 18420 2585 18430 2605
rect 18390 2555 18430 2585
rect 18390 2535 18400 2555
rect 18420 2535 18430 2555
rect 18390 2520 18430 2535
rect 18720 2610 18730 2630
rect 18750 2610 18760 2630
rect 18720 2580 18760 2610
rect 18720 2560 18730 2580
rect 18750 2560 18760 2580
rect 18720 2530 18760 2560
rect 12540 2495 12580 2510
rect 18720 2510 18730 2530
rect 18750 2510 18760 2530
rect 18720 2495 18760 2510
rect 18780 2880 18820 2895
rect 18780 2860 18790 2880
rect 18810 2860 18820 2880
rect 18780 2830 18820 2860
rect 18780 2810 18790 2830
rect 18810 2810 18820 2830
rect 18780 2780 18820 2810
rect 18780 2760 18790 2780
rect 18810 2760 18820 2780
rect 18780 2730 18820 2760
rect 18780 2710 18790 2730
rect 18810 2710 18820 2730
rect 18780 2680 18820 2710
rect 18780 2660 18790 2680
rect 18810 2660 18820 2680
rect 18780 2630 18820 2660
rect 18780 2610 18790 2630
rect 18810 2610 18820 2630
rect 18780 2580 18820 2610
rect 18780 2560 18790 2580
rect 18810 2560 18820 2580
rect 18780 2530 18820 2560
rect 18780 2510 18790 2530
rect 18810 2510 18820 2530
rect 18780 2495 18820 2510
rect 18840 2880 18880 2895
rect 18840 2860 18850 2880
rect 18870 2860 18880 2880
rect 18840 2830 18880 2860
rect 18840 2810 18850 2830
rect 18870 2810 18880 2830
rect 18840 2780 18880 2810
rect 18840 2760 18850 2780
rect 18870 2760 18880 2780
rect 18840 2730 18880 2760
rect 18840 2710 18850 2730
rect 18870 2710 18880 2730
rect 18840 2680 18880 2710
rect 18840 2660 18850 2680
rect 18870 2660 18880 2680
rect 18840 2630 18880 2660
rect 18840 2610 18850 2630
rect 18870 2610 18880 2630
rect 18840 2580 18880 2610
rect 18840 2560 18850 2580
rect 18870 2560 18880 2580
rect 18840 2530 18880 2560
rect 18840 2510 18850 2530
rect 18870 2510 18880 2530
rect 18840 2495 18880 2510
rect 18900 2880 18940 2895
rect 18900 2860 18910 2880
rect 18930 2860 18940 2880
rect 18900 2830 18940 2860
rect 18900 2810 18910 2830
rect 18930 2810 18940 2830
rect 18900 2780 18940 2810
rect 18900 2760 18910 2780
rect 18930 2760 18940 2780
rect 18900 2730 18940 2760
rect 18900 2710 18910 2730
rect 18930 2710 18940 2730
rect 18900 2680 18940 2710
rect 18900 2660 18910 2680
rect 18930 2660 18940 2680
rect 18900 2630 18940 2660
rect 18900 2610 18910 2630
rect 18930 2610 18940 2630
rect 18900 2580 18940 2610
rect 18900 2560 18910 2580
rect 18930 2560 18940 2580
rect 18900 2530 18940 2560
rect 18900 2510 18910 2530
rect 18930 2510 18940 2530
rect 18900 2495 18940 2510
rect 18960 2880 19000 2895
rect 18960 2860 18970 2880
rect 18990 2860 19000 2880
rect 18960 2830 19000 2860
rect 18960 2810 18970 2830
rect 18990 2810 19000 2830
rect 18960 2780 19000 2810
rect 18960 2760 18970 2780
rect 18990 2760 19000 2780
rect 18960 2730 19000 2760
rect 18960 2710 18970 2730
rect 18990 2710 19000 2730
rect 18960 2680 19000 2710
rect 18960 2660 18970 2680
rect 18990 2660 19000 2680
rect 18960 2630 19000 2660
rect 18960 2610 18970 2630
rect 18990 2610 19000 2630
rect 18960 2580 19000 2610
rect 18960 2560 18970 2580
rect 18990 2560 19000 2580
rect 18960 2530 19000 2560
rect 18960 2510 18970 2530
rect 18990 2510 19000 2530
rect 18960 2495 19000 2510
rect 19020 2880 19060 2895
rect 19020 2860 19030 2880
rect 19050 2860 19060 2880
rect 19020 2830 19060 2860
rect 19020 2810 19030 2830
rect 19050 2810 19060 2830
rect 19020 2780 19060 2810
rect 19020 2760 19030 2780
rect 19050 2760 19060 2780
rect 19020 2730 19060 2760
rect 19020 2710 19030 2730
rect 19050 2710 19060 2730
rect 19020 2680 19060 2710
rect 19020 2660 19030 2680
rect 19050 2660 19060 2680
rect 19020 2630 19060 2660
rect 19020 2610 19030 2630
rect 19050 2610 19060 2630
rect 19020 2580 19060 2610
rect 19020 2560 19030 2580
rect 19050 2560 19060 2580
rect 19020 2530 19060 2560
rect 19020 2510 19030 2530
rect 19050 2510 19060 2530
rect 19020 2495 19060 2510
rect 19080 2880 19120 2895
rect 19080 2860 19090 2880
rect 19110 2860 19120 2880
rect 19080 2830 19120 2860
rect 19080 2810 19090 2830
rect 19110 2810 19120 2830
rect 19080 2780 19120 2810
rect 19080 2760 19090 2780
rect 19110 2760 19120 2780
rect 19080 2730 19120 2760
rect 19080 2710 19090 2730
rect 19110 2710 19120 2730
rect 19080 2680 19120 2710
rect 19080 2660 19090 2680
rect 19110 2660 19120 2680
rect 19080 2630 19120 2660
rect 19080 2610 19090 2630
rect 19110 2610 19120 2630
rect 19080 2580 19120 2610
rect 19080 2560 19090 2580
rect 19110 2560 19120 2580
rect 19080 2530 19120 2560
rect 19080 2510 19090 2530
rect 19110 2510 19120 2530
rect 19080 2495 19120 2510
rect 19140 2880 19180 2895
rect 19140 2860 19150 2880
rect 19170 2860 19180 2880
rect 19140 2830 19180 2860
rect 19140 2810 19150 2830
rect 19170 2810 19180 2830
rect 19140 2780 19180 2810
rect 19140 2760 19150 2780
rect 19170 2760 19180 2780
rect 19140 2730 19180 2760
rect 19140 2710 19150 2730
rect 19170 2710 19180 2730
rect 19140 2680 19180 2710
rect 19140 2660 19150 2680
rect 19170 2660 19180 2680
rect 19140 2630 19180 2660
rect 19140 2610 19150 2630
rect 19170 2610 19180 2630
rect 19140 2580 19180 2610
rect 19140 2560 19150 2580
rect 19170 2560 19180 2580
rect 19140 2530 19180 2560
rect 19140 2510 19150 2530
rect 19170 2510 19180 2530
rect 19140 2495 19180 2510
rect 19200 2880 19240 2895
rect 19200 2860 19210 2880
rect 19230 2860 19240 2880
rect 19200 2830 19240 2860
rect 19200 2810 19210 2830
rect 19230 2810 19240 2830
rect 19200 2780 19240 2810
rect 19200 2760 19210 2780
rect 19230 2760 19240 2780
rect 19200 2730 19240 2760
rect 19200 2710 19210 2730
rect 19230 2710 19240 2730
rect 19200 2680 19240 2710
rect 19200 2660 19210 2680
rect 19230 2660 19240 2680
rect 19200 2630 19240 2660
rect 19200 2610 19210 2630
rect 19230 2610 19240 2630
rect 19200 2580 19240 2610
rect 19200 2560 19210 2580
rect 19230 2560 19240 2580
rect 19200 2530 19240 2560
rect 19200 2510 19210 2530
rect 19230 2510 19240 2530
rect 19200 2495 19240 2510
rect 19260 2880 19300 2895
rect 19260 2860 19270 2880
rect 19290 2860 19300 2880
rect 19260 2830 19300 2860
rect 19260 2810 19270 2830
rect 19290 2810 19300 2830
rect 19260 2780 19300 2810
rect 19260 2760 19270 2780
rect 19290 2760 19300 2780
rect 19260 2730 19300 2760
rect 19260 2710 19270 2730
rect 19290 2710 19300 2730
rect 19260 2680 19300 2710
rect 19260 2660 19270 2680
rect 19290 2660 19300 2680
rect 19260 2630 19300 2660
rect 19260 2610 19270 2630
rect 19290 2610 19300 2630
rect 19260 2580 19300 2610
rect 19260 2560 19270 2580
rect 19290 2560 19300 2580
rect 19260 2530 19300 2560
rect 19260 2510 19270 2530
rect 19290 2510 19300 2530
rect 19260 2495 19300 2510
rect 19320 2880 19360 2895
rect 19320 2860 19330 2880
rect 19350 2860 19360 2880
rect 19320 2830 19360 2860
rect 19320 2810 19330 2830
rect 19350 2810 19360 2830
rect 19320 2780 19360 2810
rect 19320 2760 19330 2780
rect 19350 2760 19360 2780
rect 19320 2730 19360 2760
rect 19320 2710 19330 2730
rect 19350 2710 19360 2730
rect 19320 2680 19360 2710
rect 19320 2660 19330 2680
rect 19350 2660 19360 2680
rect 19320 2630 19360 2660
rect 19320 2610 19330 2630
rect 19350 2610 19360 2630
rect 19320 2580 19360 2610
rect 19320 2560 19330 2580
rect 19350 2560 19360 2580
rect 19320 2530 19360 2560
rect 19320 2510 19330 2530
rect 19350 2510 19360 2530
rect 19320 2495 19360 2510
rect 19380 2880 19420 2895
rect 19380 2860 19390 2880
rect 19410 2860 19420 2880
rect 19380 2830 19420 2860
rect 19380 2810 19390 2830
rect 19410 2810 19420 2830
rect 19380 2780 19420 2810
rect 19380 2760 19390 2780
rect 19410 2760 19420 2780
rect 19380 2730 19420 2760
rect 19380 2710 19390 2730
rect 19410 2710 19420 2730
rect 19380 2680 19420 2710
rect 19380 2660 19390 2680
rect 19410 2660 19420 2680
rect 19380 2630 19420 2660
rect 19380 2610 19390 2630
rect 19410 2610 19420 2630
rect 19380 2580 19420 2610
rect 19380 2560 19390 2580
rect 19410 2560 19420 2580
rect 19380 2530 19420 2560
rect 19380 2510 19390 2530
rect 19410 2510 19420 2530
rect 19380 2495 19420 2510
rect 19440 2880 19480 2895
rect 19440 2860 19450 2880
rect 19470 2860 19480 2880
rect 19440 2830 19480 2860
rect 19440 2810 19450 2830
rect 19470 2810 19480 2830
rect 19440 2780 19480 2810
rect 19440 2760 19450 2780
rect 19470 2760 19480 2780
rect 19440 2730 19480 2760
rect 19440 2710 19450 2730
rect 19470 2710 19480 2730
rect 19440 2680 19480 2710
rect 19440 2660 19450 2680
rect 19470 2660 19480 2680
rect 19440 2630 19480 2660
rect 19440 2610 19450 2630
rect 19470 2610 19480 2630
rect 19440 2580 19480 2610
rect 19440 2560 19450 2580
rect 19470 2560 19480 2580
rect 19440 2530 19480 2560
rect 19440 2510 19450 2530
rect 19470 2510 19480 2530
rect 19440 2495 19480 2510
rect 19500 2880 19540 2895
rect 19500 2860 19510 2880
rect 19530 2860 19540 2880
rect 19500 2830 19540 2860
rect 19500 2810 19510 2830
rect 19530 2810 19540 2830
rect 19500 2780 19540 2810
rect 19500 2760 19510 2780
rect 19530 2760 19540 2780
rect 19500 2730 19540 2760
rect 19500 2710 19510 2730
rect 19530 2710 19540 2730
rect 19500 2680 19540 2710
rect 19500 2660 19510 2680
rect 19530 2660 19540 2680
rect 19500 2630 19540 2660
rect 19500 2610 19510 2630
rect 19530 2610 19540 2630
rect 19500 2580 19540 2610
rect 19500 2560 19510 2580
rect 19530 2560 19540 2580
rect 19500 2530 19540 2560
rect 19500 2510 19510 2530
rect 19530 2510 19540 2530
rect 19500 2495 19540 2510
rect 19560 2880 19600 2895
rect 19560 2860 19570 2880
rect 19590 2860 19600 2880
rect 19560 2830 19600 2860
rect 19560 2810 19570 2830
rect 19590 2810 19600 2830
rect 19560 2780 19600 2810
rect 19560 2760 19570 2780
rect 19590 2760 19600 2780
rect 19560 2730 19600 2760
rect 19560 2710 19570 2730
rect 19590 2710 19600 2730
rect 19560 2680 19600 2710
rect 19560 2660 19570 2680
rect 19590 2660 19600 2680
rect 19560 2630 19600 2660
rect 19560 2610 19570 2630
rect 19590 2610 19600 2630
rect 19560 2580 19600 2610
rect 19560 2560 19570 2580
rect 19590 2560 19600 2580
rect 19560 2530 19600 2560
rect 19560 2510 19570 2530
rect 19590 2510 19600 2530
rect 19560 2495 19600 2510
rect 19620 2880 19660 2895
rect 19620 2860 19630 2880
rect 19650 2860 19660 2880
rect 19620 2830 19660 2860
rect 19620 2810 19630 2830
rect 19650 2810 19660 2830
rect 19620 2780 19660 2810
rect 19620 2760 19630 2780
rect 19650 2760 19660 2780
rect 19620 2730 19660 2760
rect 19620 2710 19630 2730
rect 19650 2710 19660 2730
rect 19620 2680 19660 2710
rect 19620 2660 19630 2680
rect 19650 2660 19660 2680
rect 19620 2630 19660 2660
rect 19620 2610 19630 2630
rect 19650 2610 19660 2630
rect 19620 2580 19660 2610
rect 19620 2560 19630 2580
rect 19650 2560 19660 2580
rect 19620 2530 19660 2560
rect 19620 2510 19630 2530
rect 19650 2510 19660 2530
rect 19620 2495 19660 2510
rect 19680 2880 19720 2895
rect 19680 2860 19690 2880
rect 19710 2860 19720 2880
rect 19680 2830 19720 2860
rect 19680 2810 19690 2830
rect 19710 2810 19720 2830
rect 19680 2780 19720 2810
rect 19680 2760 19690 2780
rect 19710 2760 19720 2780
rect 19680 2730 19720 2760
rect 19680 2710 19690 2730
rect 19710 2710 19720 2730
rect 19680 2680 19720 2710
rect 19680 2660 19690 2680
rect 19710 2660 19720 2680
rect 19680 2630 19720 2660
rect 19680 2610 19690 2630
rect 19710 2610 19720 2630
rect 19680 2580 19720 2610
rect 19680 2560 19690 2580
rect 19710 2560 19720 2580
rect 19680 2530 19720 2560
rect 19680 2510 19690 2530
rect 19710 2510 19720 2530
rect 19680 2495 19720 2510
rect 19740 2880 19780 2895
rect 19740 2860 19750 2880
rect 19770 2860 19780 2880
rect 19740 2830 19780 2860
rect 19740 2810 19750 2830
rect 19770 2810 19780 2830
rect 19740 2780 19780 2810
rect 19740 2760 19750 2780
rect 19770 2760 19780 2780
rect 19740 2730 19780 2760
rect 19740 2710 19750 2730
rect 19770 2710 19780 2730
rect 19740 2680 19780 2710
rect 19740 2660 19750 2680
rect 19770 2660 19780 2680
rect 19740 2630 19780 2660
rect 19740 2610 19750 2630
rect 19770 2610 19780 2630
rect 19740 2580 19780 2610
rect 19740 2560 19750 2580
rect 19770 2560 19780 2580
rect 19740 2530 19780 2560
rect 19740 2510 19750 2530
rect 19770 2510 19780 2530
rect 19740 2495 19780 2510
rect 19800 2880 19840 2895
rect 19800 2860 19810 2880
rect 19830 2860 19840 2880
rect 19800 2830 19840 2860
rect 19800 2810 19810 2830
rect 19830 2810 19840 2830
rect 19800 2780 19840 2810
rect 19800 2760 19810 2780
rect 19830 2760 19840 2780
rect 19800 2730 19840 2760
rect 19800 2710 19810 2730
rect 19830 2710 19840 2730
rect 19800 2680 19840 2710
rect 19800 2660 19810 2680
rect 19830 2660 19840 2680
rect 19800 2630 19840 2660
rect 19800 2610 19810 2630
rect 19830 2610 19840 2630
rect 19800 2580 19840 2610
rect 19800 2560 19810 2580
rect 19830 2560 19840 2580
rect 19800 2530 19840 2560
rect 19800 2510 19810 2530
rect 19830 2510 19840 2530
rect 19800 2495 19840 2510
rect 19860 2880 19900 2895
rect 19860 2860 19870 2880
rect 19890 2860 19900 2880
rect 19860 2830 19900 2860
rect 19860 2810 19870 2830
rect 19890 2810 19900 2830
rect 19860 2780 19900 2810
rect 19860 2760 19870 2780
rect 19890 2760 19900 2780
rect 19860 2730 19900 2760
rect 19860 2710 19870 2730
rect 19890 2710 19900 2730
rect 19860 2680 19900 2710
rect 19860 2660 19870 2680
rect 19890 2660 19900 2680
rect 19860 2630 19900 2660
rect 19860 2610 19870 2630
rect 19890 2610 19900 2630
rect 19860 2580 19900 2610
rect 19860 2560 19870 2580
rect 19890 2560 19900 2580
rect 19860 2530 19900 2560
rect 19860 2510 19870 2530
rect 19890 2510 19900 2530
rect 19860 2495 19900 2510
rect 19920 2880 19960 2895
rect 19920 2860 19930 2880
rect 19950 2860 19960 2880
rect 19920 2830 19960 2860
rect 19920 2810 19930 2830
rect 19950 2810 19960 2830
rect 19920 2780 19960 2810
rect 19920 2760 19930 2780
rect 19950 2760 19960 2780
rect 19920 2730 19960 2760
rect 19920 2710 19930 2730
rect 19950 2710 19960 2730
rect 19920 2680 19960 2710
rect 19920 2660 19930 2680
rect 19950 2660 19960 2680
rect 19920 2630 19960 2660
rect 19920 2610 19930 2630
rect 19950 2610 19960 2630
rect 19920 2580 19960 2610
rect 19920 2560 19930 2580
rect 19950 2560 19960 2580
rect 19920 2530 19960 2560
rect 19920 2510 19930 2530
rect 19950 2510 19960 2530
rect 19920 2495 19960 2510
rect 19980 2880 20020 2895
rect 19980 2860 19990 2880
rect 20010 2860 20020 2880
rect 19980 2830 20020 2860
rect 19980 2810 19990 2830
rect 20010 2810 20020 2830
rect 19980 2780 20020 2810
rect 19980 2760 19990 2780
rect 20010 2760 20020 2780
rect 19980 2730 20020 2760
rect 19980 2710 19990 2730
rect 20010 2710 20020 2730
rect 19980 2680 20020 2710
rect 19980 2660 19990 2680
rect 20010 2660 20020 2680
rect 19980 2630 20020 2660
rect 19980 2610 19990 2630
rect 20010 2610 20020 2630
rect 19980 2580 20020 2610
rect 19980 2560 19990 2580
rect 20010 2560 20020 2580
rect 19980 2530 20020 2560
rect 19980 2510 19990 2530
rect 20010 2510 20020 2530
rect 19980 2495 20020 2510
rect 20040 2880 20080 2895
rect 20040 2860 20050 2880
rect 20070 2860 20080 2880
rect 20040 2830 20080 2860
rect 20040 2810 20050 2830
rect 20070 2810 20080 2830
rect 20040 2780 20080 2810
rect 20040 2760 20050 2780
rect 20070 2760 20080 2780
rect 20040 2730 20080 2760
rect 20040 2710 20050 2730
rect 20070 2710 20080 2730
rect 20040 2680 20080 2710
rect 20040 2660 20050 2680
rect 20070 2660 20080 2680
rect 20040 2630 20080 2660
rect 20040 2610 20050 2630
rect 20070 2610 20080 2630
rect 20040 2580 20080 2610
rect 20040 2560 20050 2580
rect 20070 2560 20080 2580
rect 20040 2530 20080 2560
rect 20040 2510 20050 2530
rect 20070 2510 20080 2530
rect 20390 2605 20430 2620
rect 20390 2585 20400 2605
rect 20420 2585 20430 2605
rect 20390 2555 20430 2585
rect 20390 2535 20400 2555
rect 20420 2535 20430 2555
rect 20390 2520 20430 2535
rect 20445 2605 20485 2620
rect 20445 2585 20455 2605
rect 20475 2585 20485 2605
rect 20445 2555 20485 2585
rect 20445 2535 20455 2555
rect 20475 2535 20485 2555
rect 20445 2520 20485 2535
rect 20500 2605 20540 2620
rect 20500 2585 20510 2605
rect 20530 2585 20540 2605
rect 20500 2555 20540 2585
rect 20500 2535 20510 2555
rect 20530 2535 20540 2555
rect 20500 2520 20540 2535
rect 20555 2605 20595 2620
rect 20555 2585 20565 2605
rect 20585 2585 20595 2605
rect 20555 2555 20595 2585
rect 20555 2535 20565 2555
rect 20585 2535 20595 2555
rect 20555 2520 20595 2535
rect 20610 2605 20650 2620
rect 20610 2585 20620 2605
rect 20640 2585 20650 2605
rect 20610 2555 20650 2585
rect 20610 2535 20620 2555
rect 20640 2535 20650 2555
rect 20610 2520 20650 2535
rect 20665 2605 20705 2620
rect 20665 2585 20675 2605
rect 20695 2585 20705 2605
rect 20665 2555 20705 2585
rect 20665 2535 20675 2555
rect 20695 2535 20705 2555
rect 20665 2520 20705 2535
rect 20720 2605 20760 2620
rect 20720 2585 20730 2605
rect 20750 2585 20760 2605
rect 20720 2555 20760 2585
rect 20720 2535 20730 2555
rect 20750 2535 20760 2555
rect 20720 2520 20760 2535
rect 20775 2605 20815 2620
rect 20775 2585 20785 2605
rect 20805 2585 20815 2605
rect 20775 2555 20815 2585
rect 20775 2535 20785 2555
rect 20805 2535 20815 2555
rect 20775 2520 20815 2535
rect 20830 2605 20870 2620
rect 20830 2585 20840 2605
rect 20860 2585 20870 2605
rect 20830 2555 20870 2585
rect 20830 2535 20840 2555
rect 20860 2535 20870 2555
rect 20830 2520 20870 2535
rect 20885 2605 20925 2620
rect 20885 2585 20895 2605
rect 20915 2585 20925 2605
rect 20885 2555 20925 2585
rect 20885 2535 20895 2555
rect 20915 2535 20925 2555
rect 20885 2520 20925 2535
rect 20940 2605 20980 2620
rect 20940 2585 20950 2605
rect 20970 2585 20980 2605
rect 20940 2555 20980 2585
rect 20940 2535 20950 2555
rect 20970 2535 20980 2555
rect 20940 2520 20980 2535
rect 20995 2605 21035 2620
rect 20995 2585 21005 2605
rect 21025 2585 21035 2605
rect 20995 2555 21035 2585
rect 20995 2535 21005 2555
rect 21025 2535 21035 2555
rect 20995 2520 21035 2535
rect 21050 2605 21090 2620
rect 21050 2585 21060 2605
rect 21080 2585 21090 2605
rect 21050 2555 21090 2585
rect 21050 2535 21060 2555
rect 21080 2535 21090 2555
rect 21050 2520 21090 2535
rect 21105 2605 21145 2620
rect 21105 2585 21115 2605
rect 21135 2585 21145 2605
rect 21105 2555 21145 2585
rect 21105 2535 21115 2555
rect 21135 2535 21145 2555
rect 21105 2520 21145 2535
rect 21160 2605 21200 2620
rect 21160 2585 21170 2605
rect 21190 2585 21200 2605
rect 21160 2555 21200 2585
rect 21160 2535 21170 2555
rect 21190 2535 21200 2555
rect 21160 2520 21200 2535
rect 21215 2605 21255 2620
rect 21215 2585 21225 2605
rect 21245 2585 21255 2605
rect 21215 2555 21255 2585
rect 21215 2535 21225 2555
rect 21245 2535 21255 2555
rect 21215 2520 21255 2535
rect 21270 2605 21310 2620
rect 21270 2585 21280 2605
rect 21300 2585 21310 2605
rect 21270 2555 21310 2585
rect 21270 2535 21280 2555
rect 21300 2535 21310 2555
rect 21270 2520 21310 2535
rect 21325 2605 21365 2620
rect 21325 2585 21335 2605
rect 21355 2585 21365 2605
rect 21325 2555 21365 2585
rect 21325 2535 21335 2555
rect 21355 2535 21365 2555
rect 21325 2520 21365 2535
rect 21380 2605 21420 2620
rect 21380 2585 21390 2605
rect 21410 2585 21420 2605
rect 21380 2555 21420 2585
rect 21380 2535 21390 2555
rect 21410 2535 21420 2555
rect 21380 2520 21420 2535
rect 21435 2605 21475 2620
rect 21435 2585 21445 2605
rect 21465 2585 21475 2605
rect 21435 2555 21475 2585
rect 21435 2535 21445 2555
rect 21465 2535 21475 2555
rect 21435 2520 21475 2535
rect 21490 2605 21530 2620
rect 21490 2585 21500 2605
rect 21520 2585 21530 2605
rect 21490 2555 21530 2585
rect 21490 2535 21500 2555
rect 21520 2535 21530 2555
rect 21490 2520 21530 2535
rect 21545 2605 21585 2620
rect 21545 2585 21555 2605
rect 21575 2585 21585 2605
rect 21545 2555 21585 2585
rect 21545 2535 21555 2555
rect 21575 2535 21585 2555
rect 21545 2520 21585 2535
rect 21600 2605 21640 2620
rect 21600 2585 21610 2605
rect 21630 2585 21640 2605
rect 21600 2555 21640 2585
rect 21600 2535 21610 2555
rect 21630 2535 21640 2555
rect 21600 2520 21640 2535
rect 20040 2495 20080 2510
rect 9680 2155 9720 2170
rect 9680 2135 9690 2155
rect 9710 2135 9720 2155
rect 9680 2105 9720 2135
rect 9680 2085 9690 2105
rect 9710 2085 9720 2105
rect 9680 2055 9720 2085
rect 9680 2035 9690 2055
rect 9710 2035 9720 2055
rect 9680 2020 9720 2035
rect 9735 2155 9775 2170
rect 9735 2135 9745 2155
rect 9765 2135 9775 2155
rect 9735 2105 9775 2135
rect 9735 2085 9745 2105
rect 9765 2085 9775 2105
rect 9735 2055 9775 2085
rect 9735 2035 9745 2055
rect 9765 2035 9775 2055
rect 9735 2020 9775 2035
rect 9790 2155 9830 2170
rect 9790 2135 9800 2155
rect 9820 2135 9830 2155
rect 9790 2105 9830 2135
rect 9790 2085 9800 2105
rect 9820 2085 9830 2105
rect 9790 2055 9830 2085
rect 9790 2035 9800 2055
rect 9820 2035 9830 2055
rect 9790 2020 9830 2035
rect 9845 2155 9885 2170
rect 9845 2135 9855 2155
rect 9875 2135 9885 2155
rect 9845 2105 9885 2135
rect 9845 2085 9855 2105
rect 9875 2085 9885 2105
rect 9845 2055 9885 2085
rect 9845 2035 9855 2055
rect 9875 2035 9885 2055
rect 9845 2020 9885 2035
rect 9900 2155 9940 2170
rect 9900 2135 9910 2155
rect 9930 2135 9940 2155
rect 9900 2105 9940 2135
rect 9900 2085 9910 2105
rect 9930 2085 9940 2105
rect 9900 2055 9940 2085
rect 9900 2035 9910 2055
rect 9930 2035 9940 2055
rect 9900 2020 9940 2035
rect 9955 2155 9995 2170
rect 9955 2135 9965 2155
rect 9985 2135 9995 2155
rect 9955 2105 9995 2135
rect 9955 2085 9965 2105
rect 9985 2085 9995 2105
rect 9955 2055 9995 2085
rect 9955 2035 9965 2055
rect 9985 2035 9995 2055
rect 9955 2020 9995 2035
rect 10010 2155 10050 2170
rect 10010 2135 10020 2155
rect 10040 2135 10050 2155
rect 10010 2105 10050 2135
rect 10010 2085 10020 2105
rect 10040 2085 10050 2105
rect 10010 2055 10050 2085
rect 10010 2035 10020 2055
rect 10040 2035 10050 2055
rect 10010 2020 10050 2035
rect 10065 2155 10105 2170
rect 10065 2135 10075 2155
rect 10095 2135 10105 2155
rect 10065 2105 10105 2135
rect 10065 2085 10075 2105
rect 10095 2085 10105 2105
rect 10065 2055 10105 2085
rect 10065 2035 10075 2055
rect 10095 2035 10105 2055
rect 10065 2020 10105 2035
rect 10120 2155 10160 2170
rect 10120 2135 10130 2155
rect 10150 2135 10160 2155
rect 10120 2105 10160 2135
rect 10120 2085 10130 2105
rect 10150 2085 10160 2105
rect 10120 2055 10160 2085
rect 10120 2035 10130 2055
rect 10150 2035 10160 2055
rect 10120 2020 10160 2035
rect 10175 2155 10215 2170
rect 10175 2135 10185 2155
rect 10205 2135 10215 2155
rect 10175 2105 10215 2135
rect 10175 2085 10185 2105
rect 10205 2085 10215 2105
rect 10175 2055 10215 2085
rect 10175 2035 10185 2055
rect 10205 2035 10215 2055
rect 10175 2020 10215 2035
rect 10230 2155 10270 2170
rect 10230 2135 10240 2155
rect 10260 2135 10270 2155
rect 10230 2105 10270 2135
rect 10230 2085 10240 2105
rect 10260 2085 10270 2105
rect 10230 2055 10270 2085
rect 10230 2035 10240 2055
rect 10260 2035 10270 2055
rect 10230 2020 10270 2035
rect 10285 2155 10325 2170
rect 10285 2135 10295 2155
rect 10315 2135 10325 2155
rect 10285 2105 10325 2135
rect 10285 2085 10295 2105
rect 10315 2085 10325 2105
rect 10285 2055 10325 2085
rect 10285 2035 10295 2055
rect 10315 2035 10325 2055
rect 10285 2020 10325 2035
rect 10340 2155 10380 2170
rect 10340 2135 10350 2155
rect 10370 2135 10380 2155
rect 10340 2105 10380 2135
rect 10340 2085 10350 2105
rect 10370 2085 10380 2105
rect 10340 2055 10380 2085
rect 10340 2035 10350 2055
rect 10370 2035 10380 2055
rect 10340 2020 10380 2035
rect 10395 2155 10435 2170
rect 10395 2135 10405 2155
rect 10425 2135 10435 2155
rect 10395 2105 10435 2135
rect 10395 2085 10405 2105
rect 10425 2085 10435 2105
rect 10395 2055 10435 2085
rect 10395 2035 10405 2055
rect 10425 2035 10435 2055
rect 10395 2020 10435 2035
rect 10450 2155 10490 2170
rect 10450 2135 10460 2155
rect 10480 2135 10490 2155
rect 10450 2105 10490 2135
rect 10450 2085 10460 2105
rect 10480 2085 10490 2105
rect 10450 2055 10490 2085
rect 10450 2035 10460 2055
rect 10480 2035 10490 2055
rect 10450 2020 10490 2035
rect 10505 2155 10545 2170
rect 10505 2135 10515 2155
rect 10535 2135 10545 2155
rect 10505 2105 10545 2135
rect 10505 2085 10515 2105
rect 10535 2085 10545 2105
rect 10505 2055 10545 2085
rect 10505 2035 10515 2055
rect 10535 2035 10545 2055
rect 10505 2020 10545 2035
rect 10560 2155 10600 2170
rect 10560 2135 10570 2155
rect 10590 2135 10600 2155
rect 10560 2105 10600 2135
rect 10560 2085 10570 2105
rect 10590 2085 10600 2105
rect 10560 2055 10600 2085
rect 10560 2035 10570 2055
rect 10590 2035 10600 2055
rect 10560 2020 10600 2035
rect 10615 2155 10655 2170
rect 10615 2135 10625 2155
rect 10645 2135 10655 2155
rect 10615 2105 10655 2135
rect 10615 2085 10625 2105
rect 10645 2085 10655 2105
rect 10615 2055 10655 2085
rect 10615 2035 10625 2055
rect 10645 2035 10655 2055
rect 10615 2020 10655 2035
rect 10670 2155 10710 2170
rect 10670 2135 10680 2155
rect 10700 2135 10710 2155
rect 10670 2105 10710 2135
rect 10670 2085 10680 2105
rect 10700 2085 10710 2105
rect 10670 2055 10710 2085
rect 10670 2035 10680 2055
rect 10700 2035 10710 2055
rect 10670 2020 10710 2035
rect 10725 2155 10765 2170
rect 10725 2135 10735 2155
rect 10755 2135 10765 2155
rect 10725 2105 10765 2135
rect 10725 2085 10735 2105
rect 10755 2085 10765 2105
rect 10725 2055 10765 2085
rect 10725 2035 10735 2055
rect 10755 2035 10765 2055
rect 10725 2020 10765 2035
rect 10780 2155 10820 2170
rect 10780 2135 10790 2155
rect 10810 2135 10820 2155
rect 10780 2105 10820 2135
rect 10780 2085 10790 2105
rect 10810 2085 10820 2105
rect 10780 2055 10820 2085
rect 10780 2035 10790 2055
rect 10810 2035 10820 2055
rect 10780 2020 10820 2035
rect 10835 2155 10875 2170
rect 10835 2135 10845 2155
rect 10865 2135 10875 2155
rect 10835 2105 10875 2135
rect 10835 2085 10845 2105
rect 10865 2085 10875 2105
rect 10835 2055 10875 2085
rect 10835 2035 10845 2055
rect 10865 2035 10875 2055
rect 10835 2020 10875 2035
rect 10890 2155 10930 2170
rect 12890 2155 12930 2170
rect 10890 2135 10900 2155
rect 10920 2135 10930 2155
rect 10890 2105 10930 2135
rect 12890 2135 12900 2155
rect 12920 2135 12930 2155
rect 10890 2085 10900 2105
rect 10920 2085 10930 2105
rect 10890 2055 10930 2085
rect 10890 2035 10900 2055
rect 10920 2035 10930 2055
rect 10890 2020 10930 2035
rect 11275 2115 11315 2130
rect 11275 2095 11285 2115
rect 11305 2095 11315 2115
rect 11275 2065 11315 2095
rect 11275 2045 11285 2065
rect 11305 2045 11315 2065
rect 11275 2015 11315 2045
rect 11275 1995 11285 2015
rect 11305 1995 11315 2015
rect 11275 1980 11315 1995
rect 11330 2115 11370 2130
rect 11330 2095 11340 2115
rect 11360 2095 11370 2115
rect 11330 2065 11370 2095
rect 11330 2045 11340 2065
rect 11360 2045 11370 2065
rect 11330 2015 11370 2045
rect 11330 1995 11340 2015
rect 11360 1995 11370 2015
rect 11330 1980 11370 1995
rect 11385 2115 11425 2130
rect 11385 2095 11395 2115
rect 11415 2095 11425 2115
rect 11385 2065 11425 2095
rect 11385 2045 11395 2065
rect 11415 2045 11425 2065
rect 11385 2015 11425 2045
rect 11385 1995 11395 2015
rect 11415 1995 11425 2015
rect 11385 1980 11425 1995
rect 11440 2115 11480 2130
rect 11440 2095 11450 2115
rect 11470 2095 11480 2115
rect 11440 2065 11480 2095
rect 11440 2045 11450 2065
rect 11470 2045 11480 2065
rect 11440 2015 11480 2045
rect 11440 1995 11450 2015
rect 11470 1995 11480 2015
rect 11440 1980 11480 1995
rect 11495 2115 11535 2130
rect 11495 2095 11505 2115
rect 11525 2095 11535 2115
rect 11495 2065 11535 2095
rect 11495 2045 11505 2065
rect 11525 2045 11535 2065
rect 11495 2015 11535 2045
rect 11495 1995 11505 2015
rect 11525 1995 11535 2015
rect 11495 1980 11535 1995
rect 11550 2115 11590 2130
rect 11550 2095 11560 2115
rect 11580 2095 11590 2115
rect 11550 2065 11590 2095
rect 11550 2045 11560 2065
rect 11580 2045 11590 2065
rect 11550 2015 11590 2045
rect 11550 1995 11560 2015
rect 11580 1995 11590 2015
rect 11550 1980 11590 1995
rect 11605 2115 11645 2130
rect 11605 2095 11615 2115
rect 11635 2095 11645 2115
rect 11605 2065 11645 2095
rect 11605 2045 11615 2065
rect 11635 2045 11645 2065
rect 11605 2015 11645 2045
rect 11605 1995 11615 2015
rect 11635 1995 11645 2015
rect 11605 1980 11645 1995
rect 11660 2115 11700 2130
rect 11660 2095 11670 2115
rect 11690 2095 11700 2115
rect 11660 2065 11700 2095
rect 11660 2045 11670 2065
rect 11690 2045 11700 2065
rect 11660 2015 11700 2045
rect 11660 1995 11670 2015
rect 11690 1995 11700 2015
rect 11660 1980 11700 1995
rect 11715 2115 11755 2130
rect 11715 2095 11725 2115
rect 11745 2095 11755 2115
rect 11715 2065 11755 2095
rect 11715 2045 11725 2065
rect 11745 2045 11755 2065
rect 11715 2015 11755 2045
rect 11715 1995 11725 2015
rect 11745 1995 11755 2015
rect 11715 1980 11755 1995
rect 11770 2115 11810 2130
rect 11770 2095 11780 2115
rect 11800 2095 11810 2115
rect 11770 2065 11810 2095
rect 11770 2045 11780 2065
rect 11800 2045 11810 2065
rect 11770 2015 11810 2045
rect 11770 1995 11780 2015
rect 11800 1995 11810 2015
rect 11770 1980 11810 1995
rect 11825 2115 11865 2130
rect 11825 2095 11835 2115
rect 11855 2095 11865 2115
rect 11825 2065 11865 2095
rect 11825 2045 11835 2065
rect 11855 2045 11865 2065
rect 11825 2015 11865 2045
rect 11825 1995 11835 2015
rect 11855 1995 11865 2015
rect 11825 1980 11865 1995
rect 11880 2115 11920 2130
rect 11880 2095 11890 2115
rect 11910 2095 11920 2115
rect 11880 2065 11920 2095
rect 11880 2045 11890 2065
rect 11910 2045 11920 2065
rect 11880 2015 11920 2045
rect 11880 1995 11890 2015
rect 11910 1995 11920 2015
rect 11880 1980 11920 1995
rect 11935 2115 11975 2130
rect 11935 2095 11945 2115
rect 11965 2095 11975 2115
rect 11935 2065 11975 2095
rect 11935 2045 11945 2065
rect 11965 2045 11975 2065
rect 11935 2015 11975 2045
rect 11935 1995 11945 2015
rect 11965 1995 11975 2015
rect 11935 1980 11975 1995
rect 11990 2115 12030 2130
rect 11990 2095 12000 2115
rect 12020 2095 12030 2115
rect 11990 2065 12030 2095
rect 11990 2045 12000 2065
rect 12020 2045 12030 2065
rect 11990 2015 12030 2045
rect 11990 1995 12000 2015
rect 12020 1995 12030 2015
rect 11990 1980 12030 1995
rect 12045 2115 12085 2130
rect 12045 2095 12055 2115
rect 12075 2095 12085 2115
rect 12045 2065 12085 2095
rect 12045 2045 12055 2065
rect 12075 2045 12085 2065
rect 12045 2015 12085 2045
rect 12045 1995 12055 2015
rect 12075 1995 12085 2015
rect 12045 1980 12085 1995
rect 12100 2115 12140 2130
rect 12100 2095 12110 2115
rect 12130 2095 12140 2115
rect 12100 2065 12140 2095
rect 12100 2045 12110 2065
rect 12130 2045 12140 2065
rect 12100 2015 12140 2045
rect 12100 1995 12110 2015
rect 12130 1995 12140 2015
rect 12100 1980 12140 1995
rect 12155 2115 12195 2130
rect 12155 2095 12165 2115
rect 12185 2095 12195 2115
rect 12155 2065 12195 2095
rect 12155 2045 12165 2065
rect 12185 2045 12195 2065
rect 12155 2015 12195 2045
rect 12155 1995 12165 2015
rect 12185 1995 12195 2015
rect 12155 1980 12195 1995
rect 12210 2115 12250 2130
rect 12210 2095 12220 2115
rect 12240 2095 12250 2115
rect 12210 2065 12250 2095
rect 12210 2045 12220 2065
rect 12240 2045 12250 2065
rect 12210 2015 12250 2045
rect 12210 1995 12220 2015
rect 12240 1995 12250 2015
rect 12210 1980 12250 1995
rect 12265 2115 12305 2130
rect 12265 2095 12275 2115
rect 12295 2095 12305 2115
rect 12265 2065 12305 2095
rect 12265 2045 12275 2065
rect 12295 2045 12305 2065
rect 12265 2015 12305 2045
rect 12265 1995 12275 2015
rect 12295 1995 12305 2015
rect 12265 1980 12305 1995
rect 12320 2115 12360 2130
rect 12320 2095 12330 2115
rect 12350 2095 12360 2115
rect 12320 2065 12360 2095
rect 12320 2045 12330 2065
rect 12350 2045 12360 2065
rect 12320 2015 12360 2045
rect 12320 1995 12330 2015
rect 12350 1995 12360 2015
rect 12320 1980 12360 1995
rect 12375 2115 12415 2130
rect 12375 2095 12385 2115
rect 12405 2095 12415 2115
rect 12375 2065 12415 2095
rect 12375 2045 12385 2065
rect 12405 2045 12415 2065
rect 12375 2015 12415 2045
rect 12375 1995 12385 2015
rect 12405 1995 12415 2015
rect 12375 1980 12415 1995
rect 12430 2115 12470 2130
rect 12430 2095 12440 2115
rect 12460 2095 12470 2115
rect 12430 2065 12470 2095
rect 12430 2045 12440 2065
rect 12460 2045 12470 2065
rect 12430 2015 12470 2045
rect 12430 1995 12440 2015
rect 12460 1995 12470 2015
rect 12430 1980 12470 1995
rect 12485 2115 12525 2130
rect 12485 2095 12495 2115
rect 12515 2095 12525 2115
rect 12485 2065 12525 2095
rect 12485 2045 12495 2065
rect 12515 2045 12525 2065
rect 12485 2015 12525 2045
rect 12890 2105 12930 2135
rect 12890 2085 12900 2105
rect 12920 2085 12930 2105
rect 12890 2055 12930 2085
rect 12890 2035 12900 2055
rect 12920 2035 12930 2055
rect 12890 2020 12930 2035
rect 12945 2155 12985 2170
rect 12945 2135 12955 2155
rect 12975 2135 12985 2155
rect 12945 2105 12985 2135
rect 12945 2085 12955 2105
rect 12975 2085 12985 2105
rect 12945 2055 12985 2085
rect 12945 2035 12955 2055
rect 12975 2035 12985 2055
rect 12945 2020 12985 2035
rect 13000 2155 13040 2170
rect 13000 2135 13010 2155
rect 13030 2135 13040 2155
rect 13000 2105 13040 2135
rect 13000 2085 13010 2105
rect 13030 2085 13040 2105
rect 13000 2055 13040 2085
rect 13000 2035 13010 2055
rect 13030 2035 13040 2055
rect 13000 2020 13040 2035
rect 13055 2155 13095 2170
rect 13055 2135 13065 2155
rect 13085 2135 13095 2155
rect 13055 2105 13095 2135
rect 13055 2085 13065 2105
rect 13085 2085 13095 2105
rect 13055 2055 13095 2085
rect 13055 2035 13065 2055
rect 13085 2035 13095 2055
rect 13055 2020 13095 2035
rect 13110 2155 13150 2170
rect 13110 2135 13120 2155
rect 13140 2135 13150 2155
rect 13110 2105 13150 2135
rect 13110 2085 13120 2105
rect 13140 2085 13150 2105
rect 13110 2055 13150 2085
rect 13110 2035 13120 2055
rect 13140 2035 13150 2055
rect 13110 2020 13150 2035
rect 13165 2155 13205 2170
rect 13165 2135 13175 2155
rect 13195 2135 13205 2155
rect 13165 2105 13205 2135
rect 13165 2085 13175 2105
rect 13195 2085 13205 2105
rect 13165 2055 13205 2085
rect 13165 2035 13175 2055
rect 13195 2035 13205 2055
rect 13165 2020 13205 2035
rect 13220 2155 13260 2170
rect 13220 2135 13230 2155
rect 13250 2135 13260 2155
rect 13220 2105 13260 2135
rect 13220 2085 13230 2105
rect 13250 2085 13260 2105
rect 13220 2055 13260 2085
rect 13220 2035 13230 2055
rect 13250 2035 13260 2055
rect 13220 2020 13260 2035
rect 13275 2155 13315 2170
rect 13275 2135 13285 2155
rect 13305 2135 13315 2155
rect 13275 2105 13315 2135
rect 13275 2085 13285 2105
rect 13305 2085 13315 2105
rect 13275 2055 13315 2085
rect 13275 2035 13285 2055
rect 13305 2035 13315 2055
rect 13275 2020 13315 2035
rect 13330 2155 13370 2170
rect 13330 2135 13340 2155
rect 13360 2135 13370 2155
rect 13330 2105 13370 2135
rect 13330 2085 13340 2105
rect 13360 2085 13370 2105
rect 13330 2055 13370 2085
rect 13330 2035 13340 2055
rect 13360 2035 13370 2055
rect 13330 2020 13370 2035
rect 13385 2155 13425 2170
rect 13385 2135 13395 2155
rect 13415 2135 13425 2155
rect 13385 2105 13425 2135
rect 13385 2085 13395 2105
rect 13415 2085 13425 2105
rect 13385 2055 13425 2085
rect 13385 2035 13395 2055
rect 13415 2035 13425 2055
rect 13385 2020 13425 2035
rect 13440 2155 13480 2170
rect 13440 2135 13450 2155
rect 13470 2135 13480 2155
rect 13440 2105 13480 2135
rect 13440 2085 13450 2105
rect 13470 2085 13480 2105
rect 13440 2055 13480 2085
rect 13440 2035 13450 2055
rect 13470 2035 13480 2055
rect 13440 2020 13480 2035
rect 13495 2155 13535 2170
rect 13495 2135 13505 2155
rect 13525 2135 13535 2155
rect 13495 2105 13535 2135
rect 13495 2085 13505 2105
rect 13525 2085 13535 2105
rect 13495 2055 13535 2085
rect 13495 2035 13505 2055
rect 13525 2035 13535 2055
rect 13495 2020 13535 2035
rect 13550 2155 13590 2170
rect 13550 2135 13560 2155
rect 13580 2135 13590 2155
rect 13550 2105 13590 2135
rect 13550 2085 13560 2105
rect 13580 2085 13590 2105
rect 13550 2055 13590 2085
rect 13550 2035 13560 2055
rect 13580 2035 13590 2055
rect 13550 2020 13590 2035
rect 13605 2155 13645 2170
rect 13605 2135 13615 2155
rect 13635 2135 13645 2155
rect 13605 2105 13645 2135
rect 13605 2085 13615 2105
rect 13635 2085 13645 2105
rect 13605 2055 13645 2085
rect 13605 2035 13615 2055
rect 13635 2035 13645 2055
rect 13605 2020 13645 2035
rect 13660 2155 13700 2170
rect 13660 2135 13670 2155
rect 13690 2135 13700 2155
rect 13660 2105 13700 2135
rect 13660 2085 13670 2105
rect 13690 2085 13700 2105
rect 13660 2055 13700 2085
rect 13660 2035 13670 2055
rect 13690 2035 13700 2055
rect 13660 2020 13700 2035
rect 13715 2155 13755 2170
rect 13715 2135 13725 2155
rect 13745 2135 13755 2155
rect 13715 2105 13755 2135
rect 13715 2085 13725 2105
rect 13745 2085 13755 2105
rect 13715 2055 13755 2085
rect 13715 2035 13725 2055
rect 13745 2035 13755 2055
rect 13715 2020 13755 2035
rect 13770 2155 13810 2170
rect 13770 2135 13780 2155
rect 13800 2135 13810 2155
rect 13770 2105 13810 2135
rect 13770 2085 13780 2105
rect 13800 2085 13810 2105
rect 13770 2055 13810 2085
rect 13770 2035 13780 2055
rect 13800 2035 13810 2055
rect 13770 2020 13810 2035
rect 13825 2155 13865 2170
rect 13825 2135 13835 2155
rect 13855 2135 13865 2155
rect 13825 2105 13865 2135
rect 13825 2085 13835 2105
rect 13855 2085 13865 2105
rect 13825 2055 13865 2085
rect 13825 2035 13835 2055
rect 13855 2035 13865 2055
rect 13825 2020 13865 2035
rect 13880 2155 13920 2170
rect 13880 2135 13890 2155
rect 13910 2135 13920 2155
rect 13880 2105 13920 2135
rect 13880 2085 13890 2105
rect 13910 2085 13920 2105
rect 13880 2055 13920 2085
rect 13880 2035 13890 2055
rect 13910 2035 13920 2055
rect 13880 2020 13920 2035
rect 13935 2155 13975 2170
rect 13935 2135 13945 2155
rect 13965 2135 13975 2155
rect 13935 2105 13975 2135
rect 13935 2085 13945 2105
rect 13965 2085 13975 2105
rect 13935 2055 13975 2085
rect 13935 2035 13945 2055
rect 13965 2035 13975 2055
rect 13935 2020 13975 2035
rect 13990 2155 14030 2170
rect 13990 2135 14000 2155
rect 14020 2135 14030 2155
rect 13990 2105 14030 2135
rect 13990 2085 14000 2105
rect 14020 2085 14030 2105
rect 13990 2055 14030 2085
rect 13990 2035 14000 2055
rect 14020 2035 14030 2055
rect 13990 2020 14030 2035
rect 14045 2155 14085 2170
rect 14045 2135 14055 2155
rect 14075 2135 14085 2155
rect 14045 2105 14085 2135
rect 14045 2085 14055 2105
rect 14075 2085 14085 2105
rect 14045 2055 14085 2085
rect 14045 2035 14055 2055
rect 14075 2035 14085 2055
rect 14045 2020 14085 2035
rect 14100 2155 14140 2170
rect 14100 2135 14110 2155
rect 14130 2135 14140 2155
rect 14100 2105 14140 2135
rect 14100 2085 14110 2105
rect 14130 2085 14140 2105
rect 14100 2055 14140 2085
rect 14100 2035 14110 2055
rect 14130 2035 14140 2055
rect 14100 2020 14140 2035
rect 17180 2155 17220 2170
rect 17180 2135 17190 2155
rect 17210 2135 17220 2155
rect 17180 2105 17220 2135
rect 17180 2085 17190 2105
rect 17210 2085 17220 2105
rect 17180 2055 17220 2085
rect 17180 2035 17190 2055
rect 17210 2035 17220 2055
rect 17180 2020 17220 2035
rect 17235 2155 17275 2170
rect 17235 2135 17245 2155
rect 17265 2135 17275 2155
rect 17235 2105 17275 2135
rect 17235 2085 17245 2105
rect 17265 2085 17275 2105
rect 17235 2055 17275 2085
rect 17235 2035 17245 2055
rect 17265 2035 17275 2055
rect 17235 2020 17275 2035
rect 17290 2155 17330 2170
rect 17290 2135 17300 2155
rect 17320 2135 17330 2155
rect 17290 2105 17330 2135
rect 17290 2085 17300 2105
rect 17320 2085 17330 2105
rect 17290 2055 17330 2085
rect 17290 2035 17300 2055
rect 17320 2035 17330 2055
rect 17290 2020 17330 2035
rect 17345 2155 17385 2170
rect 17345 2135 17355 2155
rect 17375 2135 17385 2155
rect 17345 2105 17385 2135
rect 17345 2085 17355 2105
rect 17375 2085 17385 2105
rect 17345 2055 17385 2085
rect 17345 2035 17355 2055
rect 17375 2035 17385 2055
rect 17345 2020 17385 2035
rect 17400 2155 17440 2170
rect 17400 2135 17410 2155
rect 17430 2135 17440 2155
rect 17400 2105 17440 2135
rect 17400 2085 17410 2105
rect 17430 2085 17440 2105
rect 17400 2055 17440 2085
rect 17400 2035 17410 2055
rect 17430 2035 17440 2055
rect 17400 2020 17440 2035
rect 17455 2155 17495 2170
rect 17455 2135 17465 2155
rect 17485 2135 17495 2155
rect 17455 2105 17495 2135
rect 17455 2085 17465 2105
rect 17485 2085 17495 2105
rect 17455 2055 17495 2085
rect 17455 2035 17465 2055
rect 17485 2035 17495 2055
rect 17455 2020 17495 2035
rect 17510 2155 17550 2170
rect 17510 2135 17520 2155
rect 17540 2135 17550 2155
rect 17510 2105 17550 2135
rect 17510 2085 17520 2105
rect 17540 2085 17550 2105
rect 17510 2055 17550 2085
rect 17510 2035 17520 2055
rect 17540 2035 17550 2055
rect 17510 2020 17550 2035
rect 17565 2155 17605 2170
rect 17565 2135 17575 2155
rect 17595 2135 17605 2155
rect 17565 2105 17605 2135
rect 17565 2085 17575 2105
rect 17595 2085 17605 2105
rect 17565 2055 17605 2085
rect 17565 2035 17575 2055
rect 17595 2035 17605 2055
rect 17565 2020 17605 2035
rect 17620 2155 17660 2170
rect 17620 2135 17630 2155
rect 17650 2135 17660 2155
rect 17620 2105 17660 2135
rect 17620 2085 17630 2105
rect 17650 2085 17660 2105
rect 17620 2055 17660 2085
rect 17620 2035 17630 2055
rect 17650 2035 17660 2055
rect 17620 2020 17660 2035
rect 17675 2155 17715 2170
rect 17675 2135 17685 2155
rect 17705 2135 17715 2155
rect 17675 2105 17715 2135
rect 17675 2085 17685 2105
rect 17705 2085 17715 2105
rect 17675 2055 17715 2085
rect 17675 2035 17685 2055
rect 17705 2035 17715 2055
rect 17675 2020 17715 2035
rect 17730 2155 17770 2170
rect 17730 2135 17740 2155
rect 17760 2135 17770 2155
rect 17730 2105 17770 2135
rect 17730 2085 17740 2105
rect 17760 2085 17770 2105
rect 17730 2055 17770 2085
rect 17730 2035 17740 2055
rect 17760 2035 17770 2055
rect 17730 2020 17770 2035
rect 17785 2155 17825 2170
rect 17785 2135 17795 2155
rect 17815 2135 17825 2155
rect 17785 2105 17825 2135
rect 17785 2085 17795 2105
rect 17815 2085 17825 2105
rect 17785 2055 17825 2085
rect 17785 2035 17795 2055
rect 17815 2035 17825 2055
rect 17785 2020 17825 2035
rect 17840 2155 17880 2170
rect 17840 2135 17850 2155
rect 17870 2135 17880 2155
rect 17840 2105 17880 2135
rect 17840 2085 17850 2105
rect 17870 2085 17880 2105
rect 17840 2055 17880 2085
rect 17840 2035 17850 2055
rect 17870 2035 17880 2055
rect 17840 2020 17880 2035
rect 17895 2155 17935 2170
rect 17895 2135 17905 2155
rect 17925 2135 17935 2155
rect 17895 2105 17935 2135
rect 17895 2085 17905 2105
rect 17925 2085 17935 2105
rect 17895 2055 17935 2085
rect 17895 2035 17905 2055
rect 17925 2035 17935 2055
rect 17895 2020 17935 2035
rect 17950 2155 17990 2170
rect 17950 2135 17960 2155
rect 17980 2135 17990 2155
rect 17950 2105 17990 2135
rect 17950 2085 17960 2105
rect 17980 2085 17990 2105
rect 17950 2055 17990 2085
rect 17950 2035 17960 2055
rect 17980 2035 17990 2055
rect 17950 2020 17990 2035
rect 18005 2155 18045 2170
rect 18005 2135 18015 2155
rect 18035 2135 18045 2155
rect 18005 2105 18045 2135
rect 18005 2085 18015 2105
rect 18035 2085 18045 2105
rect 18005 2055 18045 2085
rect 18005 2035 18015 2055
rect 18035 2035 18045 2055
rect 18005 2020 18045 2035
rect 18060 2155 18100 2170
rect 18060 2135 18070 2155
rect 18090 2135 18100 2155
rect 18060 2105 18100 2135
rect 18060 2085 18070 2105
rect 18090 2085 18100 2105
rect 18060 2055 18100 2085
rect 18060 2035 18070 2055
rect 18090 2035 18100 2055
rect 18060 2020 18100 2035
rect 18115 2155 18155 2170
rect 18115 2135 18125 2155
rect 18145 2135 18155 2155
rect 18115 2105 18155 2135
rect 18115 2085 18125 2105
rect 18145 2085 18155 2105
rect 18115 2055 18155 2085
rect 18115 2035 18125 2055
rect 18145 2035 18155 2055
rect 18115 2020 18155 2035
rect 18170 2155 18210 2170
rect 18170 2135 18180 2155
rect 18200 2135 18210 2155
rect 18170 2105 18210 2135
rect 18170 2085 18180 2105
rect 18200 2085 18210 2105
rect 18170 2055 18210 2085
rect 18170 2035 18180 2055
rect 18200 2035 18210 2055
rect 18170 2020 18210 2035
rect 18225 2155 18265 2170
rect 18225 2135 18235 2155
rect 18255 2135 18265 2155
rect 18225 2105 18265 2135
rect 18225 2085 18235 2105
rect 18255 2085 18265 2105
rect 18225 2055 18265 2085
rect 18225 2035 18235 2055
rect 18255 2035 18265 2055
rect 18225 2020 18265 2035
rect 18280 2155 18320 2170
rect 18280 2135 18290 2155
rect 18310 2135 18320 2155
rect 18280 2105 18320 2135
rect 18280 2085 18290 2105
rect 18310 2085 18320 2105
rect 18280 2055 18320 2085
rect 18280 2035 18290 2055
rect 18310 2035 18320 2055
rect 18280 2020 18320 2035
rect 18335 2155 18375 2170
rect 18335 2135 18345 2155
rect 18365 2135 18375 2155
rect 18335 2105 18375 2135
rect 18335 2085 18345 2105
rect 18365 2085 18375 2105
rect 18335 2055 18375 2085
rect 18335 2035 18345 2055
rect 18365 2035 18375 2055
rect 18335 2020 18375 2035
rect 18390 2155 18430 2170
rect 20390 2155 20430 2170
rect 18390 2135 18400 2155
rect 18420 2135 18430 2155
rect 18390 2105 18430 2135
rect 20390 2135 20400 2155
rect 20420 2135 20430 2155
rect 18390 2085 18400 2105
rect 18420 2085 18430 2105
rect 18390 2055 18430 2085
rect 18390 2035 18400 2055
rect 18420 2035 18430 2055
rect 18390 2020 18430 2035
rect 18775 2115 18815 2130
rect 18775 2095 18785 2115
rect 18805 2095 18815 2115
rect 18775 2065 18815 2095
rect 18775 2045 18785 2065
rect 18805 2045 18815 2065
rect 12485 1995 12495 2015
rect 12515 1995 12525 2015
rect 18775 2015 18815 2045
rect 12485 1980 12525 1995
rect 18775 1995 18785 2015
rect 18805 1995 18815 2015
rect 18775 1980 18815 1995
rect 18830 2115 18870 2130
rect 18830 2095 18840 2115
rect 18860 2095 18870 2115
rect 18830 2065 18870 2095
rect 18830 2045 18840 2065
rect 18860 2045 18870 2065
rect 18830 2015 18870 2045
rect 18830 1995 18840 2015
rect 18860 1995 18870 2015
rect 18830 1980 18870 1995
rect 18885 2115 18925 2130
rect 18885 2095 18895 2115
rect 18915 2095 18925 2115
rect 18885 2065 18925 2095
rect 18885 2045 18895 2065
rect 18915 2045 18925 2065
rect 18885 2015 18925 2045
rect 18885 1995 18895 2015
rect 18915 1995 18925 2015
rect 18885 1980 18925 1995
rect 18940 2115 18980 2130
rect 18940 2095 18950 2115
rect 18970 2095 18980 2115
rect 18940 2065 18980 2095
rect 18940 2045 18950 2065
rect 18970 2045 18980 2065
rect 18940 2015 18980 2045
rect 18940 1995 18950 2015
rect 18970 1995 18980 2015
rect 18940 1980 18980 1995
rect 18995 2115 19035 2130
rect 18995 2095 19005 2115
rect 19025 2095 19035 2115
rect 18995 2065 19035 2095
rect 18995 2045 19005 2065
rect 19025 2045 19035 2065
rect 18995 2015 19035 2045
rect 18995 1995 19005 2015
rect 19025 1995 19035 2015
rect 18995 1980 19035 1995
rect 19050 2115 19090 2130
rect 19050 2095 19060 2115
rect 19080 2095 19090 2115
rect 19050 2065 19090 2095
rect 19050 2045 19060 2065
rect 19080 2045 19090 2065
rect 19050 2015 19090 2045
rect 19050 1995 19060 2015
rect 19080 1995 19090 2015
rect 19050 1980 19090 1995
rect 19105 2115 19145 2130
rect 19105 2095 19115 2115
rect 19135 2095 19145 2115
rect 19105 2065 19145 2095
rect 19105 2045 19115 2065
rect 19135 2045 19145 2065
rect 19105 2015 19145 2045
rect 19105 1995 19115 2015
rect 19135 1995 19145 2015
rect 19105 1980 19145 1995
rect 19160 2115 19200 2130
rect 19160 2095 19170 2115
rect 19190 2095 19200 2115
rect 19160 2065 19200 2095
rect 19160 2045 19170 2065
rect 19190 2045 19200 2065
rect 19160 2015 19200 2045
rect 19160 1995 19170 2015
rect 19190 1995 19200 2015
rect 19160 1980 19200 1995
rect 19215 2115 19255 2130
rect 19215 2095 19225 2115
rect 19245 2095 19255 2115
rect 19215 2065 19255 2095
rect 19215 2045 19225 2065
rect 19245 2045 19255 2065
rect 19215 2015 19255 2045
rect 19215 1995 19225 2015
rect 19245 1995 19255 2015
rect 19215 1980 19255 1995
rect 19270 2115 19310 2130
rect 19270 2095 19280 2115
rect 19300 2095 19310 2115
rect 19270 2065 19310 2095
rect 19270 2045 19280 2065
rect 19300 2045 19310 2065
rect 19270 2015 19310 2045
rect 19270 1995 19280 2015
rect 19300 1995 19310 2015
rect 19270 1980 19310 1995
rect 19325 2115 19365 2130
rect 19325 2095 19335 2115
rect 19355 2095 19365 2115
rect 19325 2065 19365 2095
rect 19325 2045 19335 2065
rect 19355 2045 19365 2065
rect 19325 2015 19365 2045
rect 19325 1995 19335 2015
rect 19355 1995 19365 2015
rect 19325 1980 19365 1995
rect 19380 2115 19420 2130
rect 19380 2095 19390 2115
rect 19410 2095 19420 2115
rect 19380 2065 19420 2095
rect 19380 2045 19390 2065
rect 19410 2045 19420 2065
rect 19380 2015 19420 2045
rect 19380 1995 19390 2015
rect 19410 1995 19420 2015
rect 19380 1980 19420 1995
rect 19435 2115 19475 2130
rect 19435 2095 19445 2115
rect 19465 2095 19475 2115
rect 19435 2065 19475 2095
rect 19435 2045 19445 2065
rect 19465 2045 19475 2065
rect 19435 2015 19475 2045
rect 19435 1995 19445 2015
rect 19465 1995 19475 2015
rect 19435 1980 19475 1995
rect 19490 2115 19530 2130
rect 19490 2095 19500 2115
rect 19520 2095 19530 2115
rect 19490 2065 19530 2095
rect 19490 2045 19500 2065
rect 19520 2045 19530 2065
rect 19490 2015 19530 2045
rect 19490 1995 19500 2015
rect 19520 1995 19530 2015
rect 19490 1980 19530 1995
rect 19545 2115 19585 2130
rect 19545 2095 19555 2115
rect 19575 2095 19585 2115
rect 19545 2065 19585 2095
rect 19545 2045 19555 2065
rect 19575 2045 19585 2065
rect 19545 2015 19585 2045
rect 19545 1995 19555 2015
rect 19575 1995 19585 2015
rect 19545 1980 19585 1995
rect 19600 2115 19640 2130
rect 19600 2095 19610 2115
rect 19630 2095 19640 2115
rect 19600 2065 19640 2095
rect 19600 2045 19610 2065
rect 19630 2045 19640 2065
rect 19600 2015 19640 2045
rect 19600 1995 19610 2015
rect 19630 1995 19640 2015
rect 19600 1980 19640 1995
rect 19655 2115 19695 2130
rect 19655 2095 19665 2115
rect 19685 2095 19695 2115
rect 19655 2065 19695 2095
rect 19655 2045 19665 2065
rect 19685 2045 19695 2065
rect 19655 2015 19695 2045
rect 19655 1995 19665 2015
rect 19685 1995 19695 2015
rect 19655 1980 19695 1995
rect 19710 2115 19750 2130
rect 19710 2095 19720 2115
rect 19740 2095 19750 2115
rect 19710 2065 19750 2095
rect 19710 2045 19720 2065
rect 19740 2045 19750 2065
rect 19710 2015 19750 2045
rect 19710 1995 19720 2015
rect 19740 1995 19750 2015
rect 19710 1980 19750 1995
rect 19765 2115 19805 2130
rect 19765 2095 19775 2115
rect 19795 2095 19805 2115
rect 19765 2065 19805 2095
rect 19765 2045 19775 2065
rect 19795 2045 19805 2065
rect 19765 2015 19805 2045
rect 19765 1995 19775 2015
rect 19795 1995 19805 2015
rect 19765 1980 19805 1995
rect 19820 2115 19860 2130
rect 19820 2095 19830 2115
rect 19850 2095 19860 2115
rect 19820 2065 19860 2095
rect 19820 2045 19830 2065
rect 19850 2045 19860 2065
rect 19820 2015 19860 2045
rect 19820 1995 19830 2015
rect 19850 1995 19860 2015
rect 19820 1980 19860 1995
rect 19875 2115 19915 2130
rect 19875 2095 19885 2115
rect 19905 2095 19915 2115
rect 19875 2065 19915 2095
rect 19875 2045 19885 2065
rect 19905 2045 19915 2065
rect 19875 2015 19915 2045
rect 19875 1995 19885 2015
rect 19905 1995 19915 2015
rect 19875 1980 19915 1995
rect 19930 2115 19970 2130
rect 19930 2095 19940 2115
rect 19960 2095 19970 2115
rect 19930 2065 19970 2095
rect 19930 2045 19940 2065
rect 19960 2045 19970 2065
rect 19930 2015 19970 2045
rect 19930 1995 19940 2015
rect 19960 1995 19970 2015
rect 19930 1980 19970 1995
rect 19985 2115 20025 2130
rect 19985 2095 19995 2115
rect 20015 2095 20025 2115
rect 19985 2065 20025 2095
rect 19985 2045 19995 2065
rect 20015 2045 20025 2065
rect 19985 2015 20025 2045
rect 20390 2105 20430 2135
rect 20390 2085 20400 2105
rect 20420 2085 20430 2105
rect 20390 2055 20430 2085
rect 20390 2035 20400 2055
rect 20420 2035 20430 2055
rect 20390 2020 20430 2035
rect 20445 2155 20485 2170
rect 20445 2135 20455 2155
rect 20475 2135 20485 2155
rect 20445 2105 20485 2135
rect 20445 2085 20455 2105
rect 20475 2085 20485 2105
rect 20445 2055 20485 2085
rect 20445 2035 20455 2055
rect 20475 2035 20485 2055
rect 20445 2020 20485 2035
rect 20500 2155 20540 2170
rect 20500 2135 20510 2155
rect 20530 2135 20540 2155
rect 20500 2105 20540 2135
rect 20500 2085 20510 2105
rect 20530 2085 20540 2105
rect 20500 2055 20540 2085
rect 20500 2035 20510 2055
rect 20530 2035 20540 2055
rect 20500 2020 20540 2035
rect 20555 2155 20595 2170
rect 20555 2135 20565 2155
rect 20585 2135 20595 2155
rect 20555 2105 20595 2135
rect 20555 2085 20565 2105
rect 20585 2085 20595 2105
rect 20555 2055 20595 2085
rect 20555 2035 20565 2055
rect 20585 2035 20595 2055
rect 20555 2020 20595 2035
rect 20610 2155 20650 2170
rect 20610 2135 20620 2155
rect 20640 2135 20650 2155
rect 20610 2105 20650 2135
rect 20610 2085 20620 2105
rect 20640 2085 20650 2105
rect 20610 2055 20650 2085
rect 20610 2035 20620 2055
rect 20640 2035 20650 2055
rect 20610 2020 20650 2035
rect 20665 2155 20705 2170
rect 20665 2135 20675 2155
rect 20695 2135 20705 2155
rect 20665 2105 20705 2135
rect 20665 2085 20675 2105
rect 20695 2085 20705 2105
rect 20665 2055 20705 2085
rect 20665 2035 20675 2055
rect 20695 2035 20705 2055
rect 20665 2020 20705 2035
rect 20720 2155 20760 2170
rect 20720 2135 20730 2155
rect 20750 2135 20760 2155
rect 20720 2105 20760 2135
rect 20720 2085 20730 2105
rect 20750 2085 20760 2105
rect 20720 2055 20760 2085
rect 20720 2035 20730 2055
rect 20750 2035 20760 2055
rect 20720 2020 20760 2035
rect 20775 2155 20815 2170
rect 20775 2135 20785 2155
rect 20805 2135 20815 2155
rect 20775 2105 20815 2135
rect 20775 2085 20785 2105
rect 20805 2085 20815 2105
rect 20775 2055 20815 2085
rect 20775 2035 20785 2055
rect 20805 2035 20815 2055
rect 20775 2020 20815 2035
rect 20830 2155 20870 2170
rect 20830 2135 20840 2155
rect 20860 2135 20870 2155
rect 20830 2105 20870 2135
rect 20830 2085 20840 2105
rect 20860 2085 20870 2105
rect 20830 2055 20870 2085
rect 20830 2035 20840 2055
rect 20860 2035 20870 2055
rect 20830 2020 20870 2035
rect 20885 2155 20925 2170
rect 20885 2135 20895 2155
rect 20915 2135 20925 2155
rect 20885 2105 20925 2135
rect 20885 2085 20895 2105
rect 20915 2085 20925 2105
rect 20885 2055 20925 2085
rect 20885 2035 20895 2055
rect 20915 2035 20925 2055
rect 20885 2020 20925 2035
rect 20940 2155 20980 2170
rect 20940 2135 20950 2155
rect 20970 2135 20980 2155
rect 20940 2105 20980 2135
rect 20940 2085 20950 2105
rect 20970 2085 20980 2105
rect 20940 2055 20980 2085
rect 20940 2035 20950 2055
rect 20970 2035 20980 2055
rect 20940 2020 20980 2035
rect 20995 2155 21035 2170
rect 20995 2135 21005 2155
rect 21025 2135 21035 2155
rect 20995 2105 21035 2135
rect 20995 2085 21005 2105
rect 21025 2085 21035 2105
rect 20995 2055 21035 2085
rect 20995 2035 21005 2055
rect 21025 2035 21035 2055
rect 20995 2020 21035 2035
rect 21050 2155 21090 2170
rect 21050 2135 21060 2155
rect 21080 2135 21090 2155
rect 21050 2105 21090 2135
rect 21050 2085 21060 2105
rect 21080 2085 21090 2105
rect 21050 2055 21090 2085
rect 21050 2035 21060 2055
rect 21080 2035 21090 2055
rect 21050 2020 21090 2035
rect 21105 2155 21145 2170
rect 21105 2135 21115 2155
rect 21135 2135 21145 2155
rect 21105 2105 21145 2135
rect 21105 2085 21115 2105
rect 21135 2085 21145 2105
rect 21105 2055 21145 2085
rect 21105 2035 21115 2055
rect 21135 2035 21145 2055
rect 21105 2020 21145 2035
rect 21160 2155 21200 2170
rect 21160 2135 21170 2155
rect 21190 2135 21200 2155
rect 21160 2105 21200 2135
rect 21160 2085 21170 2105
rect 21190 2085 21200 2105
rect 21160 2055 21200 2085
rect 21160 2035 21170 2055
rect 21190 2035 21200 2055
rect 21160 2020 21200 2035
rect 21215 2155 21255 2170
rect 21215 2135 21225 2155
rect 21245 2135 21255 2155
rect 21215 2105 21255 2135
rect 21215 2085 21225 2105
rect 21245 2085 21255 2105
rect 21215 2055 21255 2085
rect 21215 2035 21225 2055
rect 21245 2035 21255 2055
rect 21215 2020 21255 2035
rect 21270 2155 21310 2170
rect 21270 2135 21280 2155
rect 21300 2135 21310 2155
rect 21270 2105 21310 2135
rect 21270 2085 21280 2105
rect 21300 2085 21310 2105
rect 21270 2055 21310 2085
rect 21270 2035 21280 2055
rect 21300 2035 21310 2055
rect 21270 2020 21310 2035
rect 21325 2155 21365 2170
rect 21325 2135 21335 2155
rect 21355 2135 21365 2155
rect 21325 2105 21365 2135
rect 21325 2085 21335 2105
rect 21355 2085 21365 2105
rect 21325 2055 21365 2085
rect 21325 2035 21335 2055
rect 21355 2035 21365 2055
rect 21325 2020 21365 2035
rect 21380 2155 21420 2170
rect 21380 2135 21390 2155
rect 21410 2135 21420 2155
rect 21380 2105 21420 2135
rect 21380 2085 21390 2105
rect 21410 2085 21420 2105
rect 21380 2055 21420 2085
rect 21380 2035 21390 2055
rect 21410 2035 21420 2055
rect 21380 2020 21420 2035
rect 21435 2155 21475 2170
rect 21435 2135 21445 2155
rect 21465 2135 21475 2155
rect 21435 2105 21475 2135
rect 21435 2085 21445 2105
rect 21465 2085 21475 2105
rect 21435 2055 21475 2085
rect 21435 2035 21445 2055
rect 21465 2035 21475 2055
rect 21435 2020 21475 2035
rect 21490 2155 21530 2170
rect 21490 2135 21500 2155
rect 21520 2135 21530 2155
rect 21490 2105 21530 2135
rect 21490 2085 21500 2105
rect 21520 2085 21530 2105
rect 21490 2055 21530 2085
rect 21490 2035 21500 2055
rect 21520 2035 21530 2055
rect 21490 2020 21530 2035
rect 21545 2155 21585 2170
rect 21545 2135 21555 2155
rect 21575 2135 21585 2155
rect 21545 2105 21585 2135
rect 21545 2085 21555 2105
rect 21575 2085 21585 2105
rect 21545 2055 21585 2085
rect 21545 2035 21555 2055
rect 21575 2035 21585 2055
rect 21545 2020 21585 2035
rect 21600 2155 21640 2170
rect 21600 2135 21610 2155
rect 21630 2135 21640 2155
rect 21600 2105 21640 2135
rect 21600 2085 21610 2105
rect 21630 2085 21640 2105
rect 21600 2055 21640 2085
rect 21600 2035 21610 2055
rect 21630 2035 21640 2055
rect 21600 2020 21640 2035
rect 19985 1995 19995 2015
rect 20015 1995 20025 2015
rect 19985 1980 20025 1995
rect 20490 1840 20530 1855
rect 20490 1820 20500 1840
rect 20520 1820 20530 1840
rect 20490 1790 20530 1820
rect 20490 1770 20500 1790
rect 20520 1770 20530 1790
rect 20490 1740 20530 1770
rect 20490 1720 20500 1740
rect 20520 1720 20530 1740
rect 20490 1705 20530 1720
rect 20545 1840 20585 1855
rect 20545 1820 20555 1840
rect 20575 1820 20585 1840
rect 20545 1790 20585 1820
rect 20545 1770 20555 1790
rect 20575 1770 20585 1790
rect 20545 1740 20585 1770
rect 20545 1720 20555 1740
rect 20575 1720 20585 1740
rect 20545 1705 20585 1720
rect 20600 1840 20640 1855
rect 20600 1820 20610 1840
rect 20630 1820 20640 1840
rect 20600 1790 20640 1820
rect 20600 1770 20610 1790
rect 20630 1770 20640 1790
rect 20600 1740 20640 1770
rect 20600 1720 20610 1740
rect 20630 1720 20640 1740
rect 20600 1705 20640 1720
rect 20655 1840 20695 1855
rect 20655 1820 20665 1840
rect 20685 1820 20695 1840
rect 20655 1790 20695 1820
rect 20655 1770 20665 1790
rect 20685 1770 20695 1790
rect 20655 1740 20695 1770
rect 20655 1720 20665 1740
rect 20685 1720 20695 1740
rect 20655 1705 20695 1720
rect 20710 1840 20750 1855
rect 20710 1820 20720 1840
rect 20740 1820 20750 1840
rect 20710 1790 20750 1820
rect 20710 1770 20720 1790
rect 20740 1770 20750 1790
rect 20710 1740 20750 1770
rect 20710 1720 20720 1740
rect 20740 1720 20750 1740
rect 20710 1705 20750 1720
rect 20765 1840 20805 1855
rect 20765 1820 20775 1840
rect 20795 1820 20805 1840
rect 20765 1790 20805 1820
rect 20765 1770 20775 1790
rect 20795 1770 20805 1790
rect 20765 1740 20805 1770
rect 20765 1720 20775 1740
rect 20795 1720 20805 1740
rect 20765 1705 20805 1720
rect 20820 1840 20860 1855
rect 20820 1820 20830 1840
rect 20850 1820 20860 1840
rect 20820 1790 20860 1820
rect 20820 1770 20830 1790
rect 20850 1770 20860 1790
rect 20820 1740 20860 1770
rect 20820 1720 20830 1740
rect 20850 1720 20860 1740
rect 20820 1705 20860 1720
rect 3165 1650 3205 1665
rect 3165 1630 3175 1650
rect 3195 1630 3205 1650
rect 3165 1615 3205 1630
rect 3225 1650 3265 1665
rect 3225 1630 3235 1650
rect 3255 1630 3265 1650
rect 3225 1615 3265 1630
rect 3285 1650 3325 1665
rect 3285 1630 3295 1650
rect 3315 1630 3325 1650
rect 3285 1615 3325 1630
rect 3345 1650 3385 1665
rect 3345 1630 3355 1650
rect 3375 1630 3385 1650
rect 3345 1615 3385 1630
rect 3405 1650 3445 1665
rect 3405 1630 3415 1650
rect 3435 1630 3445 1650
rect 3405 1615 3445 1630
rect 3465 1650 3505 1665
rect 3465 1630 3475 1650
rect 3495 1630 3505 1650
rect 3465 1615 3505 1630
rect 3525 1650 3565 1665
rect 3525 1630 3535 1650
rect 3555 1630 3565 1650
rect 3525 1615 3565 1630
rect 3585 1650 3625 1665
rect 3585 1630 3595 1650
rect 3615 1630 3625 1650
rect 3585 1615 3625 1630
rect 3645 1650 3685 1665
rect 3645 1630 3655 1650
rect 3675 1630 3685 1650
rect 3645 1615 3685 1630
rect 3705 1650 3745 1665
rect 3705 1630 3715 1650
rect 3735 1630 3745 1650
rect 3705 1615 3745 1630
rect 3765 1650 3805 1665
rect 3765 1630 3775 1650
rect 3795 1630 3805 1650
rect 3765 1615 3805 1630
rect 4205 1650 4245 1665
rect 4205 1630 4215 1650
rect 4235 1630 4245 1650
rect 4205 1615 4245 1630
rect 4265 1650 4305 1665
rect 4265 1630 4275 1650
rect 4295 1630 4305 1650
rect 4265 1615 4305 1630
rect 4325 1650 4365 1665
rect 4325 1630 4335 1650
rect 4355 1630 4365 1650
rect 4325 1615 4365 1630
rect 4385 1650 4425 1665
rect 4385 1630 4395 1650
rect 4415 1630 4425 1650
rect 4385 1615 4425 1630
rect 4445 1650 4485 1665
rect 4445 1630 4455 1650
rect 4475 1630 4485 1650
rect 4445 1615 4485 1630
rect 4505 1650 4545 1665
rect 4505 1630 4515 1650
rect 4535 1630 4545 1650
rect 4505 1615 4545 1630
rect 4565 1650 4605 1665
rect 4565 1630 4575 1650
rect 4595 1630 4605 1650
rect 4565 1615 4605 1630
rect 4625 1650 4665 1665
rect 4625 1630 4635 1650
rect 4655 1630 4665 1650
rect 4625 1615 4665 1630
rect 4685 1650 4725 1665
rect 4685 1630 4695 1650
rect 4715 1630 4725 1650
rect 4685 1615 4725 1630
rect 4745 1650 4785 1665
rect 4745 1630 4755 1650
rect 4775 1630 4785 1650
rect 4745 1615 4785 1630
rect 4805 1650 4845 1665
rect 4805 1630 4815 1650
rect 4835 1630 4845 1650
rect 4805 1615 4845 1630
rect 11030 1650 11070 1665
rect 11030 1630 11040 1650
rect 11060 1630 11070 1650
rect 11030 1600 11070 1630
rect 11030 1580 11040 1600
rect 11060 1580 11070 1600
rect 11030 1550 11070 1580
rect 11030 1530 11040 1550
rect 11060 1530 11070 1550
rect 11030 1515 11070 1530
rect 11085 1650 11125 1665
rect 11085 1630 11095 1650
rect 11115 1630 11125 1650
rect 11085 1600 11125 1630
rect 11085 1580 11095 1600
rect 11115 1580 11125 1600
rect 11085 1550 11125 1580
rect 11085 1530 11095 1550
rect 11115 1530 11125 1550
rect 11085 1515 11125 1530
rect 11140 1650 11180 1665
rect 11140 1630 11150 1650
rect 11170 1630 11180 1650
rect 11140 1600 11180 1630
rect 11140 1580 11150 1600
rect 11170 1580 11180 1600
rect 11140 1550 11180 1580
rect 11140 1530 11150 1550
rect 11170 1530 11180 1550
rect 11140 1515 11180 1530
rect 11195 1650 11235 1665
rect 11195 1630 11205 1650
rect 11225 1630 11235 1650
rect 11195 1600 11235 1630
rect 11195 1580 11205 1600
rect 11225 1580 11235 1600
rect 11195 1550 11235 1580
rect 11195 1530 11205 1550
rect 11225 1530 11235 1550
rect 11195 1515 11235 1530
rect 11250 1650 11290 1665
rect 11250 1630 11260 1650
rect 11280 1630 11290 1650
rect 11250 1600 11290 1630
rect 11250 1580 11260 1600
rect 11280 1580 11290 1600
rect 11250 1550 11290 1580
rect 11250 1530 11260 1550
rect 11280 1530 11290 1550
rect 11250 1515 11290 1530
rect 11305 1650 11345 1665
rect 11305 1630 11315 1650
rect 11335 1630 11345 1650
rect 11305 1600 11345 1630
rect 11305 1580 11315 1600
rect 11335 1580 11345 1600
rect 11305 1550 11345 1580
rect 11305 1530 11315 1550
rect 11335 1530 11345 1550
rect 11305 1515 11345 1530
rect 11360 1650 11400 1665
rect 11360 1630 11370 1650
rect 11390 1630 11400 1650
rect 11360 1600 11400 1630
rect 11360 1580 11370 1600
rect 11390 1580 11400 1600
rect 11360 1550 11400 1580
rect 11360 1530 11370 1550
rect 11390 1530 11400 1550
rect 11360 1515 11400 1530
rect 11415 1650 11455 1665
rect 11415 1630 11425 1650
rect 11445 1630 11455 1650
rect 11415 1600 11455 1630
rect 11415 1580 11425 1600
rect 11445 1580 11455 1600
rect 11415 1550 11455 1580
rect 11415 1530 11425 1550
rect 11445 1530 11455 1550
rect 11415 1515 11455 1530
rect 11470 1650 11510 1665
rect 11470 1630 11480 1650
rect 11500 1630 11510 1650
rect 11470 1600 11510 1630
rect 11470 1580 11480 1600
rect 11500 1580 11510 1600
rect 11470 1550 11510 1580
rect 11470 1530 11480 1550
rect 11500 1530 11510 1550
rect 11470 1515 11510 1530
rect 11525 1650 11565 1665
rect 11525 1630 11535 1650
rect 11555 1630 11565 1650
rect 11525 1600 11565 1630
rect 11525 1580 11535 1600
rect 11555 1580 11565 1600
rect 11525 1550 11565 1580
rect 11525 1530 11535 1550
rect 11555 1530 11565 1550
rect 11525 1515 11565 1530
rect 11580 1650 11620 1665
rect 11580 1630 11590 1650
rect 11610 1630 11620 1650
rect 11580 1600 11620 1630
rect 11580 1580 11590 1600
rect 11610 1580 11620 1600
rect 11580 1550 11620 1580
rect 11580 1530 11590 1550
rect 11610 1530 11620 1550
rect 11580 1515 11620 1530
rect 11635 1650 11675 1665
rect 11635 1630 11645 1650
rect 11665 1630 11675 1650
rect 11635 1600 11675 1630
rect 11635 1580 11645 1600
rect 11665 1580 11675 1600
rect 11635 1550 11675 1580
rect 11635 1530 11645 1550
rect 11665 1530 11675 1550
rect 11635 1515 11675 1530
rect 11690 1650 11730 1665
rect 11770 1650 11810 1665
rect 11690 1630 11700 1650
rect 11720 1630 11730 1650
rect 11770 1630 11780 1650
rect 11800 1630 11810 1650
rect 11690 1600 11730 1630
rect 11770 1600 11810 1630
rect 11690 1580 11700 1600
rect 11720 1580 11730 1600
rect 11770 1580 11780 1600
rect 11800 1580 11810 1600
rect 11690 1550 11730 1580
rect 11770 1550 11810 1580
rect 11690 1530 11700 1550
rect 11720 1530 11730 1550
rect 11770 1530 11780 1550
rect 11800 1530 11810 1550
rect 11690 1515 11730 1530
rect 11770 1515 11810 1530
rect 11825 1650 11865 1665
rect 11825 1630 11835 1650
rect 11855 1630 11865 1650
rect 11825 1600 11865 1630
rect 11825 1580 11835 1600
rect 11855 1580 11865 1600
rect 11825 1550 11865 1580
rect 11825 1530 11835 1550
rect 11855 1530 11865 1550
rect 11825 1515 11865 1530
rect 11880 1650 11920 1665
rect 11880 1630 11890 1650
rect 11910 1630 11920 1650
rect 11880 1600 11920 1630
rect 11880 1580 11890 1600
rect 11910 1580 11920 1600
rect 11880 1550 11920 1580
rect 11880 1530 11890 1550
rect 11910 1530 11920 1550
rect 11880 1515 11920 1530
rect 11935 1650 11975 1665
rect 11935 1630 11945 1650
rect 11965 1630 11975 1650
rect 11935 1600 11975 1630
rect 11935 1580 11945 1600
rect 11965 1580 11975 1600
rect 11935 1550 11975 1580
rect 11935 1530 11945 1550
rect 11965 1530 11975 1550
rect 11935 1515 11975 1530
rect 11990 1650 12030 1665
rect 12070 1650 12110 1665
rect 11990 1630 12000 1650
rect 12020 1630 12030 1650
rect 12070 1630 12080 1650
rect 12100 1630 12110 1650
rect 11990 1600 12030 1630
rect 12070 1600 12110 1630
rect 11990 1580 12000 1600
rect 12020 1580 12030 1600
rect 12070 1580 12080 1600
rect 12100 1580 12110 1600
rect 11990 1550 12030 1580
rect 12070 1550 12110 1580
rect 11990 1530 12000 1550
rect 12020 1530 12030 1550
rect 12070 1530 12080 1550
rect 12100 1530 12110 1550
rect 11990 1515 12030 1530
rect 12070 1515 12110 1530
rect 12125 1650 12165 1665
rect 12125 1630 12135 1650
rect 12155 1630 12165 1650
rect 12125 1600 12165 1630
rect 12125 1580 12135 1600
rect 12155 1580 12165 1600
rect 12125 1550 12165 1580
rect 12125 1530 12135 1550
rect 12155 1530 12165 1550
rect 12125 1515 12165 1530
rect 12180 1650 12220 1665
rect 12180 1630 12190 1650
rect 12210 1630 12220 1650
rect 12180 1600 12220 1630
rect 12180 1580 12190 1600
rect 12210 1580 12220 1600
rect 12180 1550 12220 1580
rect 12180 1530 12190 1550
rect 12210 1530 12220 1550
rect 12180 1515 12220 1530
rect 12235 1650 12275 1665
rect 12235 1630 12245 1650
rect 12265 1630 12275 1650
rect 12235 1600 12275 1630
rect 12235 1580 12245 1600
rect 12265 1580 12275 1600
rect 12235 1550 12275 1580
rect 12235 1530 12245 1550
rect 12265 1530 12275 1550
rect 12235 1515 12275 1530
rect 12290 1650 12330 1665
rect 12290 1630 12300 1650
rect 12320 1630 12330 1650
rect 12290 1600 12330 1630
rect 12290 1580 12300 1600
rect 12320 1580 12330 1600
rect 12290 1550 12330 1580
rect 12290 1530 12300 1550
rect 12320 1530 12330 1550
rect 12290 1515 12330 1530
rect 12345 1650 12385 1665
rect 12345 1630 12355 1650
rect 12375 1630 12385 1650
rect 12345 1600 12385 1630
rect 12345 1580 12355 1600
rect 12375 1580 12385 1600
rect 12345 1550 12385 1580
rect 12345 1530 12355 1550
rect 12375 1530 12385 1550
rect 12345 1515 12385 1530
rect 12400 1650 12440 1665
rect 12400 1630 12410 1650
rect 12430 1630 12440 1650
rect 12400 1600 12440 1630
rect 12400 1580 12410 1600
rect 12430 1580 12440 1600
rect 12400 1550 12440 1580
rect 12400 1530 12410 1550
rect 12430 1530 12440 1550
rect 12400 1515 12440 1530
rect 12455 1650 12495 1665
rect 12455 1630 12465 1650
rect 12485 1630 12495 1650
rect 12455 1600 12495 1630
rect 12455 1580 12465 1600
rect 12485 1580 12495 1600
rect 12455 1550 12495 1580
rect 12455 1530 12465 1550
rect 12485 1530 12495 1550
rect 12455 1515 12495 1530
rect 12510 1650 12550 1665
rect 12510 1630 12520 1650
rect 12540 1630 12550 1650
rect 12510 1600 12550 1630
rect 12510 1580 12520 1600
rect 12540 1580 12550 1600
rect 12510 1550 12550 1580
rect 12510 1530 12520 1550
rect 12540 1530 12550 1550
rect 12510 1515 12550 1530
rect 12565 1650 12605 1665
rect 12565 1630 12575 1650
rect 12595 1630 12605 1650
rect 12565 1600 12605 1630
rect 12565 1580 12575 1600
rect 12595 1580 12605 1600
rect 12565 1550 12605 1580
rect 12565 1530 12575 1550
rect 12595 1530 12605 1550
rect 12565 1515 12605 1530
rect 12620 1650 12660 1665
rect 12620 1630 12630 1650
rect 12650 1630 12660 1650
rect 12620 1600 12660 1630
rect 12620 1580 12630 1600
rect 12650 1580 12660 1600
rect 12620 1550 12660 1580
rect 12620 1530 12630 1550
rect 12650 1530 12660 1550
rect 12620 1515 12660 1530
rect 12675 1650 12715 1665
rect 12675 1630 12685 1650
rect 12705 1630 12715 1650
rect 12675 1600 12715 1630
rect 12675 1580 12685 1600
rect 12705 1580 12715 1600
rect 12675 1550 12715 1580
rect 12675 1530 12685 1550
rect 12705 1530 12715 1550
rect 12675 1515 12715 1530
rect 12730 1650 12770 1665
rect 12730 1630 12740 1650
rect 12760 1630 12770 1650
rect 12730 1600 12770 1630
rect 12730 1580 12740 1600
rect 12760 1580 12770 1600
rect 12730 1550 12770 1580
rect 12730 1530 12740 1550
rect 12760 1530 12770 1550
rect 12730 1515 12770 1530
rect 18530 1650 18570 1665
rect 18530 1630 18540 1650
rect 18560 1630 18570 1650
rect 18530 1600 18570 1630
rect 18530 1580 18540 1600
rect 18560 1580 18570 1600
rect 18530 1550 18570 1580
rect 18530 1530 18540 1550
rect 18560 1530 18570 1550
rect 18530 1515 18570 1530
rect 18585 1650 18625 1665
rect 18585 1630 18595 1650
rect 18615 1630 18625 1650
rect 18585 1600 18625 1630
rect 18585 1580 18595 1600
rect 18615 1580 18625 1600
rect 18585 1550 18625 1580
rect 18585 1530 18595 1550
rect 18615 1530 18625 1550
rect 18585 1515 18625 1530
rect 18640 1650 18680 1665
rect 18640 1630 18650 1650
rect 18670 1630 18680 1650
rect 18640 1600 18680 1630
rect 18640 1580 18650 1600
rect 18670 1580 18680 1600
rect 18640 1550 18680 1580
rect 18640 1530 18650 1550
rect 18670 1530 18680 1550
rect 18640 1515 18680 1530
rect 18695 1650 18735 1665
rect 18695 1630 18705 1650
rect 18725 1630 18735 1650
rect 18695 1600 18735 1630
rect 18695 1580 18705 1600
rect 18725 1580 18735 1600
rect 18695 1550 18735 1580
rect 18695 1530 18705 1550
rect 18725 1530 18735 1550
rect 18695 1515 18735 1530
rect 18750 1650 18790 1665
rect 18750 1630 18760 1650
rect 18780 1630 18790 1650
rect 18750 1600 18790 1630
rect 18750 1580 18760 1600
rect 18780 1580 18790 1600
rect 18750 1550 18790 1580
rect 18750 1530 18760 1550
rect 18780 1530 18790 1550
rect 18750 1515 18790 1530
rect 18805 1650 18845 1665
rect 18805 1630 18815 1650
rect 18835 1630 18845 1650
rect 18805 1600 18845 1630
rect 18805 1580 18815 1600
rect 18835 1580 18845 1600
rect 18805 1550 18845 1580
rect 18805 1530 18815 1550
rect 18835 1530 18845 1550
rect 18805 1515 18845 1530
rect 18860 1650 18900 1665
rect 18860 1630 18870 1650
rect 18890 1630 18900 1650
rect 18860 1600 18900 1630
rect 18860 1580 18870 1600
rect 18890 1580 18900 1600
rect 18860 1550 18900 1580
rect 18860 1530 18870 1550
rect 18890 1530 18900 1550
rect 18860 1515 18900 1530
rect 18915 1650 18955 1665
rect 18915 1630 18925 1650
rect 18945 1630 18955 1650
rect 18915 1600 18955 1630
rect 18915 1580 18925 1600
rect 18945 1580 18955 1600
rect 18915 1550 18955 1580
rect 18915 1530 18925 1550
rect 18945 1530 18955 1550
rect 18915 1515 18955 1530
rect 18970 1650 19010 1665
rect 18970 1630 18980 1650
rect 19000 1630 19010 1650
rect 18970 1600 19010 1630
rect 18970 1580 18980 1600
rect 19000 1580 19010 1600
rect 18970 1550 19010 1580
rect 18970 1530 18980 1550
rect 19000 1530 19010 1550
rect 18970 1515 19010 1530
rect 19025 1650 19065 1665
rect 19025 1630 19035 1650
rect 19055 1630 19065 1650
rect 19025 1600 19065 1630
rect 19025 1580 19035 1600
rect 19055 1580 19065 1600
rect 19025 1550 19065 1580
rect 19025 1530 19035 1550
rect 19055 1530 19065 1550
rect 19025 1515 19065 1530
rect 19080 1650 19120 1665
rect 19080 1630 19090 1650
rect 19110 1630 19120 1650
rect 19080 1600 19120 1630
rect 19080 1580 19090 1600
rect 19110 1580 19120 1600
rect 19080 1550 19120 1580
rect 19080 1530 19090 1550
rect 19110 1530 19120 1550
rect 19080 1515 19120 1530
rect 19135 1650 19175 1665
rect 19135 1630 19145 1650
rect 19165 1630 19175 1650
rect 19135 1600 19175 1630
rect 19135 1580 19145 1600
rect 19165 1580 19175 1600
rect 19135 1550 19175 1580
rect 19135 1530 19145 1550
rect 19165 1530 19175 1550
rect 19135 1515 19175 1530
rect 19190 1650 19230 1665
rect 19270 1650 19310 1665
rect 19190 1630 19200 1650
rect 19220 1630 19230 1650
rect 19270 1630 19280 1650
rect 19300 1630 19310 1650
rect 19190 1600 19230 1630
rect 19270 1600 19310 1630
rect 19190 1580 19200 1600
rect 19220 1580 19230 1600
rect 19270 1580 19280 1600
rect 19300 1580 19310 1600
rect 19190 1550 19230 1580
rect 19270 1550 19310 1580
rect 19190 1530 19200 1550
rect 19220 1530 19230 1550
rect 19270 1530 19280 1550
rect 19300 1530 19310 1550
rect 19190 1515 19230 1530
rect 19270 1515 19310 1530
rect 19325 1650 19365 1665
rect 19325 1630 19335 1650
rect 19355 1630 19365 1650
rect 19325 1600 19365 1630
rect 19325 1580 19335 1600
rect 19355 1580 19365 1600
rect 19325 1550 19365 1580
rect 19325 1530 19335 1550
rect 19355 1530 19365 1550
rect 19325 1515 19365 1530
rect 19380 1650 19420 1665
rect 19380 1630 19390 1650
rect 19410 1630 19420 1650
rect 19380 1600 19420 1630
rect 19380 1580 19390 1600
rect 19410 1580 19420 1600
rect 19380 1550 19420 1580
rect 19380 1530 19390 1550
rect 19410 1530 19420 1550
rect 19380 1515 19420 1530
rect 19435 1650 19475 1665
rect 19435 1630 19445 1650
rect 19465 1630 19475 1650
rect 19435 1600 19475 1630
rect 19435 1580 19445 1600
rect 19465 1580 19475 1600
rect 19435 1550 19475 1580
rect 19435 1530 19445 1550
rect 19465 1530 19475 1550
rect 19435 1515 19475 1530
rect 19490 1650 19530 1665
rect 19570 1650 19610 1665
rect 19490 1630 19500 1650
rect 19520 1630 19530 1650
rect 19570 1630 19580 1650
rect 19600 1630 19610 1650
rect 19490 1600 19530 1630
rect 19570 1600 19610 1630
rect 19490 1580 19500 1600
rect 19520 1580 19530 1600
rect 19570 1580 19580 1600
rect 19600 1580 19610 1600
rect 19490 1550 19530 1580
rect 19570 1550 19610 1580
rect 19490 1530 19500 1550
rect 19520 1530 19530 1550
rect 19570 1530 19580 1550
rect 19600 1530 19610 1550
rect 19490 1515 19530 1530
rect 19570 1515 19610 1530
rect 19625 1650 19665 1665
rect 19625 1630 19635 1650
rect 19655 1630 19665 1650
rect 19625 1600 19665 1630
rect 19625 1580 19635 1600
rect 19655 1580 19665 1600
rect 19625 1550 19665 1580
rect 19625 1530 19635 1550
rect 19655 1530 19665 1550
rect 19625 1515 19665 1530
rect 19680 1650 19720 1665
rect 19680 1630 19690 1650
rect 19710 1630 19720 1650
rect 19680 1600 19720 1630
rect 19680 1580 19690 1600
rect 19710 1580 19720 1600
rect 19680 1550 19720 1580
rect 19680 1530 19690 1550
rect 19710 1530 19720 1550
rect 19680 1515 19720 1530
rect 19735 1650 19775 1665
rect 19735 1630 19745 1650
rect 19765 1630 19775 1650
rect 19735 1600 19775 1630
rect 19735 1580 19745 1600
rect 19765 1580 19775 1600
rect 19735 1550 19775 1580
rect 19735 1530 19745 1550
rect 19765 1530 19775 1550
rect 19735 1515 19775 1530
rect 19790 1650 19830 1665
rect 19790 1630 19800 1650
rect 19820 1630 19830 1650
rect 19790 1600 19830 1630
rect 19790 1580 19800 1600
rect 19820 1580 19830 1600
rect 19790 1550 19830 1580
rect 19790 1530 19800 1550
rect 19820 1530 19830 1550
rect 19790 1515 19830 1530
rect 19845 1650 19885 1665
rect 19845 1630 19855 1650
rect 19875 1630 19885 1650
rect 19845 1600 19885 1630
rect 19845 1580 19855 1600
rect 19875 1580 19885 1600
rect 19845 1550 19885 1580
rect 19845 1530 19855 1550
rect 19875 1530 19885 1550
rect 19845 1515 19885 1530
rect 19900 1650 19940 1665
rect 19900 1630 19910 1650
rect 19930 1630 19940 1650
rect 19900 1600 19940 1630
rect 19900 1580 19910 1600
rect 19930 1580 19940 1600
rect 19900 1550 19940 1580
rect 19900 1530 19910 1550
rect 19930 1530 19940 1550
rect 19900 1515 19940 1530
rect 19955 1650 19995 1665
rect 19955 1630 19965 1650
rect 19985 1630 19995 1650
rect 19955 1600 19995 1630
rect 19955 1580 19965 1600
rect 19985 1580 19995 1600
rect 19955 1550 19995 1580
rect 19955 1530 19965 1550
rect 19985 1530 19995 1550
rect 19955 1515 19995 1530
rect 20010 1650 20050 1665
rect 20010 1630 20020 1650
rect 20040 1630 20050 1650
rect 20010 1600 20050 1630
rect 20010 1580 20020 1600
rect 20040 1580 20050 1600
rect 20010 1550 20050 1580
rect 20010 1530 20020 1550
rect 20040 1530 20050 1550
rect 20010 1515 20050 1530
rect 20065 1650 20105 1665
rect 20065 1630 20075 1650
rect 20095 1630 20105 1650
rect 20065 1600 20105 1630
rect 20065 1580 20075 1600
rect 20095 1580 20105 1600
rect 20065 1550 20105 1580
rect 20065 1530 20075 1550
rect 20095 1530 20105 1550
rect 20065 1515 20105 1530
rect 20120 1650 20160 1665
rect 20120 1630 20130 1650
rect 20150 1630 20160 1650
rect 20120 1600 20160 1630
rect 20120 1580 20130 1600
rect 20150 1580 20160 1600
rect 20120 1550 20160 1580
rect 20120 1530 20130 1550
rect 20150 1530 20160 1550
rect 20120 1515 20160 1530
rect 20175 1650 20215 1665
rect 20175 1630 20185 1650
rect 20205 1630 20215 1650
rect 20175 1600 20215 1630
rect 20175 1580 20185 1600
rect 20205 1580 20215 1600
rect 20175 1550 20215 1580
rect 20175 1530 20185 1550
rect 20205 1530 20215 1550
rect 20175 1515 20215 1530
rect 20230 1650 20270 1665
rect 20230 1630 20240 1650
rect 20260 1630 20270 1650
rect 20230 1600 20270 1630
rect 20230 1580 20240 1600
rect 20260 1580 20270 1600
rect 20230 1550 20270 1580
rect 20230 1530 20240 1550
rect 20260 1530 20270 1550
rect 20230 1515 20270 1530
rect 20395 1505 20435 1520
rect 20395 1485 20405 1505
rect 20425 1485 20435 1505
rect 20395 1455 20435 1485
rect 2835 1440 2875 1455
rect 2835 1420 2845 1440
rect 2865 1420 2875 1440
rect 2835 1390 2875 1420
rect 2835 1370 2845 1390
rect 2865 1370 2875 1390
rect 2835 1340 2875 1370
rect 2835 1320 2845 1340
rect 2865 1320 2875 1340
rect 2835 1290 2875 1320
rect 2835 1270 2845 1290
rect 2865 1270 2875 1290
rect 2835 1240 2875 1270
rect 2835 1220 2845 1240
rect 2865 1220 2875 1240
rect 2835 1205 2875 1220
rect 3375 1440 3415 1455
rect 3375 1420 3385 1440
rect 3405 1420 3415 1440
rect 3375 1390 3415 1420
rect 3375 1370 3385 1390
rect 3405 1370 3415 1390
rect 3375 1340 3415 1370
rect 3375 1320 3385 1340
rect 3405 1320 3415 1340
rect 3375 1290 3415 1320
rect 3375 1270 3385 1290
rect 3405 1270 3415 1290
rect 3375 1240 3415 1270
rect 3375 1220 3385 1240
rect 3405 1220 3415 1240
rect 3375 1205 3415 1220
rect 3915 1440 3955 1455
rect 3915 1420 3925 1440
rect 3945 1420 3955 1440
rect 3915 1390 3955 1420
rect 3915 1370 3925 1390
rect 3945 1370 3955 1390
rect 3915 1340 3955 1370
rect 3915 1320 3925 1340
rect 3945 1320 3955 1340
rect 3915 1290 3955 1320
rect 3915 1270 3925 1290
rect 3945 1270 3955 1290
rect 3915 1240 3955 1270
rect 3915 1220 3925 1240
rect 3945 1220 3955 1240
rect 3915 1205 3955 1220
rect 4055 1440 4095 1455
rect 4055 1420 4065 1440
rect 4085 1420 4095 1440
rect 4055 1390 4095 1420
rect 4055 1370 4065 1390
rect 4085 1370 4095 1390
rect 4055 1340 4095 1370
rect 4055 1320 4065 1340
rect 4085 1320 4095 1340
rect 4055 1290 4095 1320
rect 4055 1270 4065 1290
rect 4085 1270 4095 1290
rect 4055 1240 4095 1270
rect 4055 1220 4065 1240
rect 4085 1220 4095 1240
rect 4055 1205 4095 1220
rect 4595 1440 4635 1455
rect 4595 1420 4605 1440
rect 4625 1420 4635 1440
rect 4595 1390 4635 1420
rect 4595 1370 4605 1390
rect 4625 1370 4635 1390
rect 4595 1340 4635 1370
rect 4595 1320 4605 1340
rect 4625 1320 4635 1340
rect 4595 1290 4635 1320
rect 4595 1270 4605 1290
rect 4625 1270 4635 1290
rect 4595 1240 4635 1270
rect 4595 1220 4605 1240
rect 4625 1220 4635 1240
rect 4595 1205 4635 1220
rect 5135 1440 5175 1455
rect 5135 1420 5145 1440
rect 5165 1420 5175 1440
rect 20395 1435 20405 1455
rect 20425 1435 20435 1455
rect 5135 1390 5175 1420
rect 20395 1405 20435 1435
rect 5135 1370 5145 1390
rect 5165 1370 5175 1390
rect 20395 1385 20405 1405
rect 20425 1385 20435 1405
rect 20395 1370 20435 1385
rect 20450 1505 20490 1520
rect 20450 1485 20460 1505
rect 20480 1485 20490 1505
rect 20450 1455 20490 1485
rect 20450 1435 20460 1455
rect 20480 1435 20490 1455
rect 20450 1405 20490 1435
rect 20450 1385 20460 1405
rect 20480 1385 20490 1405
rect 20450 1370 20490 1385
rect 20505 1505 20545 1520
rect 20505 1485 20515 1505
rect 20535 1485 20545 1505
rect 20505 1455 20545 1485
rect 20505 1435 20515 1455
rect 20535 1435 20545 1455
rect 20505 1405 20545 1435
rect 20505 1385 20515 1405
rect 20535 1385 20545 1405
rect 20505 1370 20545 1385
rect 20560 1505 20600 1520
rect 20560 1485 20570 1505
rect 20590 1485 20600 1505
rect 20560 1455 20600 1485
rect 20560 1435 20570 1455
rect 20590 1435 20600 1455
rect 20560 1405 20600 1435
rect 20560 1385 20570 1405
rect 20590 1385 20600 1405
rect 20560 1370 20600 1385
rect 20615 1505 20655 1520
rect 20695 1505 20735 1520
rect 20615 1485 20625 1505
rect 20645 1485 20655 1505
rect 20695 1485 20705 1505
rect 20725 1485 20735 1505
rect 20615 1455 20655 1485
rect 20695 1455 20735 1485
rect 20615 1435 20625 1455
rect 20645 1435 20655 1455
rect 20695 1435 20705 1455
rect 20725 1435 20735 1455
rect 20615 1405 20655 1435
rect 20695 1405 20735 1435
rect 20615 1385 20625 1405
rect 20645 1385 20655 1405
rect 20695 1385 20705 1405
rect 20725 1385 20735 1405
rect 20615 1370 20655 1385
rect 20695 1370 20735 1385
rect 20750 1505 20790 1520
rect 20750 1485 20760 1505
rect 20780 1485 20790 1505
rect 20750 1455 20790 1485
rect 20750 1435 20760 1455
rect 20780 1435 20790 1455
rect 20750 1405 20790 1435
rect 20750 1385 20760 1405
rect 20780 1385 20790 1405
rect 20750 1370 20790 1385
rect 20805 1505 20845 1520
rect 20805 1485 20815 1505
rect 20835 1485 20845 1505
rect 20805 1455 20845 1485
rect 20805 1435 20815 1455
rect 20835 1435 20845 1455
rect 20805 1405 20845 1435
rect 20805 1385 20815 1405
rect 20835 1385 20845 1405
rect 20805 1370 20845 1385
rect 20860 1505 20900 1520
rect 20860 1485 20870 1505
rect 20890 1485 20900 1505
rect 20860 1455 20900 1485
rect 20860 1435 20870 1455
rect 20890 1435 20900 1455
rect 20860 1405 20900 1435
rect 20860 1385 20870 1405
rect 20890 1385 20900 1405
rect 20860 1370 20900 1385
rect 20915 1505 20955 1520
rect 20915 1485 20925 1505
rect 20945 1485 20955 1505
rect 20915 1455 20955 1485
rect 20915 1435 20925 1455
rect 20945 1435 20955 1455
rect 20915 1405 20955 1435
rect 20915 1385 20925 1405
rect 20945 1385 20955 1405
rect 20915 1370 20955 1385
rect 5135 1340 5175 1370
rect 5135 1320 5145 1340
rect 5165 1320 5175 1340
rect 5135 1290 5175 1320
rect 5135 1270 5145 1290
rect 5165 1270 5175 1290
rect 5135 1240 5175 1270
rect 12925 1255 12965 1270
rect 5135 1220 5145 1240
rect 5165 1220 5175 1240
rect 5135 1205 5175 1220
rect 12925 1235 12935 1255
rect 12955 1235 12965 1255
rect 12925 1210 12965 1235
rect 12925 1190 12935 1210
rect 12955 1190 12965 1210
rect 11205 1160 11245 1175
rect 11205 1140 11215 1160
rect 11235 1140 11245 1160
rect 11205 1110 11245 1140
rect 11205 1090 11215 1110
rect 11235 1090 11245 1110
rect 2945 1060 2985 1075
rect 2945 1040 2955 1060
rect 2975 1040 2985 1060
rect 2945 1010 2985 1040
rect 2945 990 2955 1010
rect 2975 990 2985 1010
rect 2945 975 2985 990
rect 3985 1060 4025 1075
rect 3985 1040 3995 1060
rect 4015 1040 4025 1060
rect 3985 1010 4025 1040
rect 3985 990 3995 1010
rect 4015 990 4025 1010
rect 3985 975 4025 990
rect 5025 1060 5065 1075
rect 5025 1040 5035 1060
rect 5055 1040 5065 1060
rect 5025 1010 5065 1040
rect 5025 990 5035 1010
rect 5055 990 5065 1010
rect 5025 975 5065 990
rect 11205 1060 11245 1090
rect 11205 1040 11215 1060
rect 11235 1040 11245 1060
rect 11205 1010 11245 1040
rect 11205 990 11215 1010
rect 11235 990 11245 1010
rect 11205 960 11245 990
rect 11205 940 11215 960
rect 11235 940 11245 960
rect 11205 925 11245 940
rect 11260 1160 11300 1175
rect 11260 1140 11270 1160
rect 11290 1140 11300 1160
rect 11260 1110 11300 1140
rect 11260 1090 11270 1110
rect 11290 1090 11300 1110
rect 11260 1060 11300 1090
rect 11260 1040 11270 1060
rect 11290 1040 11300 1060
rect 11260 1010 11300 1040
rect 11260 990 11270 1010
rect 11290 990 11300 1010
rect 11260 960 11300 990
rect 11260 940 11270 960
rect 11290 940 11300 960
rect 11260 925 11300 940
rect 11315 1160 11355 1175
rect 11315 1140 11325 1160
rect 11345 1140 11355 1160
rect 11315 1110 11355 1140
rect 11315 1090 11325 1110
rect 11345 1090 11355 1110
rect 11315 1060 11355 1090
rect 11315 1040 11325 1060
rect 11345 1040 11355 1060
rect 11315 1010 11355 1040
rect 11315 990 11325 1010
rect 11345 990 11355 1010
rect 11315 960 11355 990
rect 11315 940 11325 960
rect 11345 940 11355 960
rect 11315 925 11355 940
rect 11370 1160 11410 1175
rect 11370 1140 11380 1160
rect 11400 1140 11410 1160
rect 11370 1110 11410 1140
rect 11370 1090 11380 1110
rect 11400 1090 11410 1110
rect 11370 1060 11410 1090
rect 11370 1040 11380 1060
rect 11400 1040 11410 1060
rect 11370 1010 11410 1040
rect 11370 990 11380 1010
rect 11400 990 11410 1010
rect 11370 960 11410 990
rect 11370 940 11380 960
rect 11400 940 11410 960
rect 11370 925 11410 940
rect 11425 1160 11465 1175
rect 11425 1140 11435 1160
rect 11455 1140 11465 1160
rect 11425 1110 11465 1140
rect 11425 1090 11435 1110
rect 11455 1090 11465 1110
rect 11425 1060 11465 1090
rect 11425 1040 11435 1060
rect 11455 1040 11465 1060
rect 11425 1010 11465 1040
rect 11425 990 11435 1010
rect 11455 990 11465 1010
rect 11425 960 11465 990
rect 11425 940 11435 960
rect 11455 940 11465 960
rect 11425 925 11465 940
rect 11480 1160 11520 1175
rect 11480 1140 11490 1160
rect 11510 1140 11520 1160
rect 11480 1110 11520 1140
rect 11480 1090 11490 1110
rect 11510 1090 11520 1110
rect 11480 1060 11520 1090
rect 11480 1040 11490 1060
rect 11510 1040 11520 1060
rect 11480 1010 11520 1040
rect 11480 990 11490 1010
rect 11510 990 11520 1010
rect 11480 960 11520 990
rect 11480 940 11490 960
rect 11510 940 11520 960
rect 11480 925 11520 940
rect 11535 1160 11575 1175
rect 11535 1140 11545 1160
rect 11565 1140 11575 1160
rect 11535 1110 11575 1140
rect 11535 1090 11545 1110
rect 11565 1090 11575 1110
rect 11535 1060 11575 1090
rect 11535 1040 11545 1060
rect 11565 1040 11575 1060
rect 11535 1010 11575 1040
rect 11535 990 11545 1010
rect 11565 990 11575 1010
rect 11535 960 11575 990
rect 11535 940 11545 960
rect 11565 940 11575 960
rect 11535 925 11575 940
rect 11590 1160 11630 1175
rect 11590 1140 11600 1160
rect 11620 1140 11630 1160
rect 11590 1110 11630 1140
rect 11590 1090 11600 1110
rect 11620 1090 11630 1110
rect 11590 1060 11630 1090
rect 11590 1040 11600 1060
rect 11620 1040 11630 1060
rect 11590 1010 11630 1040
rect 11590 990 11600 1010
rect 11620 990 11630 1010
rect 11590 960 11630 990
rect 11590 940 11600 960
rect 11620 940 11630 960
rect 11590 925 11630 940
rect 11645 1160 11685 1175
rect 11645 1140 11655 1160
rect 11675 1140 11685 1160
rect 11645 1110 11685 1140
rect 11645 1090 11655 1110
rect 11675 1090 11685 1110
rect 11645 1060 11685 1090
rect 11645 1040 11655 1060
rect 11675 1040 11685 1060
rect 11645 1010 11685 1040
rect 11645 990 11655 1010
rect 11675 990 11685 1010
rect 11645 960 11685 990
rect 11645 940 11655 960
rect 11675 940 11685 960
rect 11645 925 11685 940
rect 11700 1160 11740 1175
rect 11700 1140 11710 1160
rect 11730 1140 11740 1160
rect 11700 1110 11740 1140
rect 11700 1090 11710 1110
rect 11730 1090 11740 1110
rect 11700 1060 11740 1090
rect 11700 1040 11710 1060
rect 11730 1040 11740 1060
rect 11700 1010 11740 1040
rect 11700 990 11710 1010
rect 11730 990 11740 1010
rect 11700 960 11740 990
rect 11700 940 11710 960
rect 11730 940 11740 960
rect 11700 925 11740 940
rect 11755 1160 11795 1175
rect 11755 1140 11765 1160
rect 11785 1140 11795 1160
rect 11755 1110 11795 1140
rect 11755 1090 11765 1110
rect 11785 1090 11795 1110
rect 11755 1060 11795 1090
rect 11755 1040 11765 1060
rect 11785 1040 11795 1060
rect 11755 1010 11795 1040
rect 11755 990 11765 1010
rect 11785 990 11795 1010
rect 11755 960 11795 990
rect 11755 940 11765 960
rect 11785 940 11795 960
rect 11755 925 11795 940
rect 11810 1160 11850 1175
rect 11810 1140 11820 1160
rect 11840 1140 11850 1160
rect 11810 1110 11850 1140
rect 11810 1090 11820 1110
rect 11840 1090 11850 1110
rect 11810 1060 11850 1090
rect 11810 1040 11820 1060
rect 11840 1040 11850 1060
rect 11810 1010 11850 1040
rect 11810 990 11820 1010
rect 11840 990 11850 1010
rect 11810 960 11850 990
rect 11810 940 11820 960
rect 11840 940 11850 960
rect 11810 925 11850 940
rect 11865 1160 11905 1175
rect 11865 1140 11875 1160
rect 11895 1140 11905 1160
rect 11865 1110 11905 1140
rect 11865 1090 11875 1110
rect 11895 1090 11905 1110
rect 11865 1060 11905 1090
rect 11865 1040 11875 1060
rect 11895 1040 11905 1060
rect 11865 1010 11905 1040
rect 11865 990 11875 1010
rect 11895 990 11905 1010
rect 11865 960 11905 990
rect 11865 940 11875 960
rect 11895 940 11905 960
rect 11865 925 11905 940
rect 11920 1160 11960 1175
rect 11920 1140 11930 1160
rect 11950 1140 11960 1160
rect 11920 1110 11960 1140
rect 11920 1090 11930 1110
rect 11950 1090 11960 1110
rect 11920 1060 11960 1090
rect 11920 1040 11930 1060
rect 11950 1040 11960 1060
rect 11920 1010 11960 1040
rect 11920 990 11930 1010
rect 11950 990 11960 1010
rect 11920 960 11960 990
rect 11920 940 11930 960
rect 11950 940 11960 960
rect 11920 925 11960 940
rect 11975 1160 12015 1175
rect 11975 1140 11985 1160
rect 12005 1140 12015 1160
rect 11975 1110 12015 1140
rect 11975 1090 11985 1110
rect 12005 1090 12015 1110
rect 11975 1060 12015 1090
rect 11975 1040 11985 1060
rect 12005 1040 12015 1060
rect 11975 1010 12015 1040
rect 11975 990 11985 1010
rect 12005 990 12015 1010
rect 11975 960 12015 990
rect 11975 940 11985 960
rect 12005 940 12015 960
rect 11975 925 12015 940
rect 12030 1160 12070 1175
rect 12030 1140 12040 1160
rect 12060 1140 12070 1160
rect 12030 1110 12070 1140
rect 12030 1090 12040 1110
rect 12060 1090 12070 1110
rect 12030 1060 12070 1090
rect 12030 1040 12040 1060
rect 12060 1040 12070 1060
rect 12030 1010 12070 1040
rect 12030 990 12040 1010
rect 12060 990 12070 1010
rect 12030 960 12070 990
rect 12030 940 12040 960
rect 12060 940 12070 960
rect 12030 925 12070 940
rect 12085 1160 12125 1175
rect 12085 1140 12095 1160
rect 12115 1140 12125 1160
rect 12085 1110 12125 1140
rect 12085 1090 12095 1110
rect 12115 1090 12125 1110
rect 12085 1060 12125 1090
rect 12085 1040 12095 1060
rect 12115 1040 12125 1060
rect 12085 1010 12125 1040
rect 12085 990 12095 1010
rect 12115 990 12125 1010
rect 12085 960 12125 990
rect 12085 940 12095 960
rect 12115 940 12125 960
rect 12085 925 12125 940
rect 12140 1160 12180 1175
rect 12140 1140 12150 1160
rect 12170 1140 12180 1160
rect 12140 1110 12180 1140
rect 12140 1090 12150 1110
rect 12170 1090 12180 1110
rect 12140 1060 12180 1090
rect 12140 1040 12150 1060
rect 12170 1040 12180 1060
rect 12140 1010 12180 1040
rect 12140 990 12150 1010
rect 12170 990 12180 1010
rect 12140 960 12180 990
rect 12140 940 12150 960
rect 12170 940 12180 960
rect 12140 925 12180 940
rect 12195 1160 12235 1175
rect 12195 1140 12205 1160
rect 12225 1140 12235 1160
rect 12195 1110 12235 1140
rect 12195 1090 12205 1110
rect 12225 1090 12235 1110
rect 12195 1060 12235 1090
rect 12195 1040 12205 1060
rect 12225 1040 12235 1060
rect 12195 1010 12235 1040
rect 12195 990 12205 1010
rect 12225 990 12235 1010
rect 12195 960 12235 990
rect 12195 940 12205 960
rect 12225 940 12235 960
rect 12195 925 12235 940
rect 12250 1160 12290 1175
rect 12250 1140 12260 1160
rect 12280 1140 12290 1160
rect 12250 1110 12290 1140
rect 12250 1090 12260 1110
rect 12280 1090 12290 1110
rect 12250 1060 12290 1090
rect 12250 1040 12260 1060
rect 12280 1040 12290 1060
rect 12250 1010 12290 1040
rect 12250 990 12260 1010
rect 12280 990 12290 1010
rect 12250 960 12290 990
rect 12250 940 12260 960
rect 12280 940 12290 960
rect 12250 925 12290 940
rect 12305 1160 12345 1175
rect 12305 1140 12315 1160
rect 12335 1140 12345 1160
rect 12305 1110 12345 1140
rect 12305 1090 12315 1110
rect 12335 1090 12345 1110
rect 12305 1060 12345 1090
rect 12305 1040 12315 1060
rect 12335 1040 12345 1060
rect 12305 1010 12345 1040
rect 12305 990 12315 1010
rect 12335 990 12345 1010
rect 12305 960 12345 990
rect 12305 940 12315 960
rect 12335 940 12345 960
rect 12305 925 12345 940
rect 12360 1160 12400 1175
rect 12360 1140 12370 1160
rect 12390 1140 12400 1160
rect 12360 1110 12400 1140
rect 12360 1090 12370 1110
rect 12390 1090 12400 1110
rect 12360 1060 12400 1090
rect 12360 1040 12370 1060
rect 12390 1040 12400 1060
rect 12360 1010 12400 1040
rect 12360 990 12370 1010
rect 12390 990 12400 1010
rect 12360 960 12400 990
rect 12360 940 12370 960
rect 12390 940 12400 960
rect 12360 925 12400 940
rect 12415 1160 12455 1175
rect 12415 1140 12425 1160
rect 12445 1140 12455 1160
rect 12415 1110 12455 1140
rect 12415 1090 12425 1110
rect 12445 1090 12455 1110
rect 12415 1060 12455 1090
rect 12415 1040 12425 1060
rect 12445 1040 12455 1060
rect 12415 1010 12455 1040
rect 12415 990 12425 1010
rect 12445 990 12455 1010
rect 12415 960 12455 990
rect 12415 940 12425 960
rect 12445 940 12455 960
rect 12415 925 12455 940
rect 12470 1160 12510 1175
rect 12470 1140 12480 1160
rect 12500 1140 12510 1160
rect 12470 1110 12510 1140
rect 12470 1090 12480 1110
rect 12500 1090 12510 1110
rect 12470 1060 12510 1090
rect 12470 1040 12480 1060
rect 12500 1040 12510 1060
rect 12470 1010 12510 1040
rect 12470 990 12480 1010
rect 12500 990 12510 1010
rect 12470 960 12510 990
rect 12470 940 12480 960
rect 12500 940 12510 960
rect 12470 925 12510 940
rect 12525 1160 12565 1175
rect 12525 1140 12535 1160
rect 12555 1140 12565 1160
rect 12525 1110 12565 1140
rect 12525 1090 12535 1110
rect 12555 1090 12565 1110
rect 12525 1060 12565 1090
rect 12525 1040 12535 1060
rect 12555 1040 12565 1060
rect 12525 1010 12565 1040
rect 12525 990 12535 1010
rect 12555 990 12565 1010
rect 12525 960 12565 990
rect 12525 940 12535 960
rect 12555 940 12565 960
rect 12525 925 12565 940
rect 12580 1160 12620 1175
rect 12580 1140 12590 1160
rect 12610 1140 12620 1160
rect 12580 1110 12620 1140
rect 12580 1090 12590 1110
rect 12610 1090 12620 1110
rect 12580 1060 12620 1090
rect 12580 1040 12590 1060
rect 12610 1040 12620 1060
rect 12580 1010 12620 1040
rect 12580 990 12590 1010
rect 12610 990 12620 1010
rect 12925 1165 12965 1190
rect 12925 1145 12935 1165
rect 12955 1145 12965 1165
rect 12925 1115 12965 1145
rect 12925 1095 12935 1115
rect 12955 1095 12965 1115
rect 12925 1070 12965 1095
rect 12925 1050 12935 1070
rect 12955 1050 12965 1070
rect 12925 1025 12965 1050
rect 12925 1005 12935 1025
rect 12955 1005 12965 1025
rect 12925 990 12965 1005
rect 13025 1255 13065 1270
rect 13025 1235 13035 1255
rect 13055 1235 13065 1255
rect 13025 1210 13065 1235
rect 13025 1190 13035 1210
rect 13055 1190 13065 1210
rect 13025 1165 13065 1190
rect 13025 1145 13035 1165
rect 13055 1145 13065 1165
rect 13025 1115 13065 1145
rect 13025 1095 13035 1115
rect 13055 1095 13065 1115
rect 13025 1070 13065 1095
rect 13025 1050 13035 1070
rect 13055 1050 13065 1070
rect 13025 1025 13065 1050
rect 13025 1005 13035 1025
rect 13055 1005 13065 1025
rect 13025 990 13065 1005
rect 13125 1255 13165 1270
rect 13125 1235 13135 1255
rect 13155 1235 13165 1255
rect 13125 1210 13165 1235
rect 13125 1190 13135 1210
rect 13155 1190 13165 1210
rect 13125 1165 13165 1190
rect 13125 1145 13135 1165
rect 13155 1145 13165 1165
rect 13125 1115 13165 1145
rect 13125 1095 13135 1115
rect 13155 1095 13165 1115
rect 13125 1070 13165 1095
rect 13125 1050 13135 1070
rect 13155 1050 13165 1070
rect 13125 1025 13165 1050
rect 13125 1005 13135 1025
rect 13155 1005 13165 1025
rect 13125 990 13165 1005
rect 13225 1255 13265 1270
rect 13225 1235 13235 1255
rect 13255 1235 13265 1255
rect 13225 1210 13265 1235
rect 13225 1190 13235 1210
rect 13255 1190 13265 1210
rect 13225 1165 13265 1190
rect 13225 1145 13235 1165
rect 13255 1145 13265 1165
rect 13225 1115 13265 1145
rect 13225 1095 13235 1115
rect 13255 1095 13265 1115
rect 13225 1070 13265 1095
rect 13225 1050 13235 1070
rect 13255 1050 13265 1070
rect 13225 1025 13265 1050
rect 13225 1005 13235 1025
rect 13255 1005 13265 1025
rect 13225 990 13265 1005
rect 13325 1255 13365 1270
rect 13325 1235 13335 1255
rect 13355 1235 13365 1255
rect 13325 1210 13365 1235
rect 13325 1190 13335 1210
rect 13355 1190 13365 1210
rect 13325 1165 13365 1190
rect 13325 1145 13335 1165
rect 13355 1145 13365 1165
rect 13325 1115 13365 1145
rect 13325 1095 13335 1115
rect 13355 1095 13365 1115
rect 13325 1070 13365 1095
rect 13325 1050 13335 1070
rect 13355 1050 13365 1070
rect 13325 1025 13365 1050
rect 13325 1005 13335 1025
rect 13355 1005 13365 1025
rect 13325 990 13365 1005
rect 13425 1255 13465 1270
rect 13425 1235 13435 1255
rect 13455 1235 13465 1255
rect 13425 1210 13465 1235
rect 13425 1190 13435 1210
rect 13455 1190 13465 1210
rect 13425 1165 13465 1190
rect 13425 1145 13435 1165
rect 13455 1145 13465 1165
rect 13425 1115 13465 1145
rect 13425 1095 13435 1115
rect 13455 1095 13465 1115
rect 13425 1070 13465 1095
rect 13425 1050 13435 1070
rect 13455 1050 13465 1070
rect 13425 1025 13465 1050
rect 13425 1005 13435 1025
rect 13455 1005 13465 1025
rect 13425 990 13465 1005
rect 13525 1255 13565 1270
rect 13525 1235 13535 1255
rect 13555 1235 13565 1255
rect 13525 1210 13565 1235
rect 13525 1190 13535 1210
rect 13555 1190 13565 1210
rect 13525 1165 13565 1190
rect 13525 1145 13535 1165
rect 13555 1145 13565 1165
rect 13525 1115 13565 1145
rect 13525 1095 13535 1115
rect 13555 1095 13565 1115
rect 13525 1070 13565 1095
rect 13525 1050 13535 1070
rect 13555 1050 13565 1070
rect 13525 1025 13565 1050
rect 13525 1005 13535 1025
rect 13555 1005 13565 1025
rect 13525 990 13565 1005
rect 13625 1255 13665 1270
rect 13625 1235 13635 1255
rect 13655 1235 13665 1255
rect 13625 1210 13665 1235
rect 13625 1190 13635 1210
rect 13655 1190 13665 1210
rect 13625 1165 13665 1190
rect 13625 1145 13635 1165
rect 13655 1145 13665 1165
rect 13625 1115 13665 1145
rect 13625 1095 13635 1115
rect 13655 1095 13665 1115
rect 13625 1070 13665 1095
rect 13625 1050 13635 1070
rect 13655 1050 13665 1070
rect 13625 1025 13665 1050
rect 13625 1005 13635 1025
rect 13655 1005 13665 1025
rect 13625 990 13665 1005
rect 13725 1255 13765 1270
rect 13725 1235 13735 1255
rect 13755 1235 13765 1255
rect 13725 1210 13765 1235
rect 13725 1190 13735 1210
rect 13755 1190 13765 1210
rect 13725 1165 13765 1190
rect 13725 1145 13735 1165
rect 13755 1145 13765 1165
rect 13725 1115 13765 1145
rect 13725 1095 13735 1115
rect 13755 1095 13765 1115
rect 13725 1070 13765 1095
rect 13725 1050 13735 1070
rect 13755 1050 13765 1070
rect 13725 1025 13765 1050
rect 13725 1005 13735 1025
rect 13755 1005 13765 1025
rect 13725 990 13765 1005
rect 13825 1255 13865 1270
rect 13825 1235 13835 1255
rect 13855 1235 13865 1255
rect 13825 1210 13865 1235
rect 13825 1190 13835 1210
rect 13855 1190 13865 1210
rect 13825 1165 13865 1190
rect 13825 1145 13835 1165
rect 13855 1145 13865 1165
rect 13825 1115 13865 1145
rect 13825 1095 13835 1115
rect 13855 1095 13865 1115
rect 13825 1070 13865 1095
rect 13825 1050 13835 1070
rect 13855 1050 13865 1070
rect 13825 1025 13865 1050
rect 13825 1005 13835 1025
rect 13855 1005 13865 1025
rect 13825 990 13865 1005
rect 13925 1255 13965 1270
rect 13925 1235 13935 1255
rect 13955 1235 13965 1255
rect 13925 1210 13965 1235
rect 13925 1190 13935 1210
rect 13955 1190 13965 1210
rect 13925 1165 13965 1190
rect 13925 1145 13935 1165
rect 13955 1145 13965 1165
rect 13925 1115 13965 1145
rect 13925 1095 13935 1115
rect 13955 1095 13965 1115
rect 13925 1070 13965 1095
rect 13925 1050 13935 1070
rect 13955 1050 13965 1070
rect 13925 1025 13965 1050
rect 13925 1005 13935 1025
rect 13955 1005 13965 1025
rect 13925 990 13965 1005
rect 14025 1255 14065 1270
rect 14025 1235 14035 1255
rect 14055 1235 14065 1255
rect 14025 1210 14065 1235
rect 14025 1190 14035 1210
rect 14055 1190 14065 1210
rect 14025 1165 14065 1190
rect 14025 1145 14035 1165
rect 14055 1145 14065 1165
rect 14025 1115 14065 1145
rect 14025 1095 14035 1115
rect 14055 1095 14065 1115
rect 14025 1070 14065 1095
rect 14025 1050 14035 1070
rect 14055 1050 14065 1070
rect 14025 1025 14065 1050
rect 14025 1005 14035 1025
rect 14055 1005 14065 1025
rect 14025 990 14065 1005
rect 14125 1255 14165 1270
rect 14125 1235 14135 1255
rect 14155 1235 14165 1255
rect 14125 1210 14165 1235
rect 14125 1190 14135 1210
rect 14155 1190 14165 1210
rect 14125 1165 14165 1190
rect 14125 1145 14135 1165
rect 14155 1145 14165 1165
rect 14125 1115 14165 1145
rect 14125 1095 14135 1115
rect 14155 1095 14165 1115
rect 14125 1070 14165 1095
rect 14125 1050 14135 1070
rect 14155 1050 14165 1070
rect 14125 1025 14165 1050
rect 14125 1005 14135 1025
rect 14155 1005 14165 1025
rect 14125 990 14165 1005
rect 18705 1210 18745 1225
rect 18705 1190 18715 1210
rect 18735 1190 18745 1210
rect 18705 1160 18745 1190
rect 18705 1140 18715 1160
rect 18735 1140 18745 1160
rect 18705 1110 18745 1140
rect 18705 1090 18715 1110
rect 18735 1090 18745 1110
rect 18705 1060 18745 1090
rect 18705 1040 18715 1060
rect 18735 1040 18745 1060
rect 18705 1010 18745 1040
rect 18705 990 18715 1010
rect 18735 990 18745 1010
rect 12580 960 12620 990
rect 12580 940 12590 960
rect 12610 940 12620 960
rect 12580 925 12620 940
rect 18705 975 18745 990
rect 18760 1210 18800 1225
rect 18760 1190 18770 1210
rect 18790 1190 18800 1210
rect 18760 1160 18800 1190
rect 18760 1140 18770 1160
rect 18790 1140 18800 1160
rect 18760 1110 18800 1140
rect 18760 1090 18770 1110
rect 18790 1090 18800 1110
rect 18760 1060 18800 1090
rect 18760 1040 18770 1060
rect 18790 1040 18800 1060
rect 18760 1010 18800 1040
rect 18760 990 18770 1010
rect 18790 990 18800 1010
rect 18760 975 18800 990
rect 18815 1210 18855 1225
rect 18815 1190 18825 1210
rect 18845 1190 18855 1210
rect 18815 1160 18855 1190
rect 18815 1140 18825 1160
rect 18845 1140 18855 1160
rect 18815 1110 18855 1140
rect 18815 1090 18825 1110
rect 18845 1090 18855 1110
rect 18815 1060 18855 1090
rect 18815 1040 18825 1060
rect 18845 1040 18855 1060
rect 18815 1010 18855 1040
rect 18815 990 18825 1010
rect 18845 990 18855 1010
rect 18815 975 18855 990
rect 18870 1210 18910 1225
rect 18870 1190 18880 1210
rect 18900 1190 18910 1210
rect 18870 1160 18910 1190
rect 18870 1140 18880 1160
rect 18900 1140 18910 1160
rect 18870 1110 18910 1140
rect 18870 1090 18880 1110
rect 18900 1090 18910 1110
rect 18870 1060 18910 1090
rect 18870 1040 18880 1060
rect 18900 1040 18910 1060
rect 18870 1010 18910 1040
rect 18870 990 18880 1010
rect 18900 990 18910 1010
rect 18870 975 18910 990
rect 18925 1210 18965 1225
rect 18925 1190 18935 1210
rect 18955 1190 18965 1210
rect 18925 1160 18965 1190
rect 18925 1140 18935 1160
rect 18955 1140 18965 1160
rect 18925 1110 18965 1140
rect 18925 1090 18935 1110
rect 18955 1090 18965 1110
rect 18925 1060 18965 1090
rect 18925 1040 18935 1060
rect 18955 1040 18965 1060
rect 18925 1010 18965 1040
rect 18925 990 18935 1010
rect 18955 990 18965 1010
rect 18925 975 18965 990
rect 18980 1210 19020 1225
rect 18980 1190 18990 1210
rect 19010 1190 19020 1210
rect 18980 1160 19020 1190
rect 18980 1140 18990 1160
rect 19010 1140 19020 1160
rect 18980 1110 19020 1140
rect 18980 1090 18990 1110
rect 19010 1090 19020 1110
rect 18980 1060 19020 1090
rect 18980 1040 18990 1060
rect 19010 1040 19020 1060
rect 18980 1010 19020 1040
rect 18980 990 18990 1010
rect 19010 990 19020 1010
rect 18980 975 19020 990
rect 19035 1210 19075 1225
rect 19035 1190 19045 1210
rect 19065 1190 19075 1210
rect 19035 1160 19075 1190
rect 19035 1140 19045 1160
rect 19065 1140 19075 1160
rect 19035 1110 19075 1140
rect 19035 1090 19045 1110
rect 19065 1090 19075 1110
rect 19035 1060 19075 1090
rect 19035 1040 19045 1060
rect 19065 1040 19075 1060
rect 19035 1010 19075 1040
rect 19035 990 19045 1010
rect 19065 990 19075 1010
rect 19035 975 19075 990
rect 19090 1210 19130 1225
rect 19090 1190 19100 1210
rect 19120 1190 19130 1210
rect 19090 1160 19130 1190
rect 19090 1140 19100 1160
rect 19120 1140 19130 1160
rect 19090 1110 19130 1140
rect 19090 1090 19100 1110
rect 19120 1090 19130 1110
rect 19090 1060 19130 1090
rect 19090 1040 19100 1060
rect 19120 1040 19130 1060
rect 19090 1010 19130 1040
rect 19090 990 19100 1010
rect 19120 990 19130 1010
rect 19090 975 19130 990
rect 19145 1210 19185 1225
rect 19145 1190 19155 1210
rect 19175 1190 19185 1210
rect 19145 1160 19185 1190
rect 19145 1140 19155 1160
rect 19175 1140 19185 1160
rect 19145 1110 19185 1140
rect 19145 1090 19155 1110
rect 19175 1090 19185 1110
rect 19145 1060 19185 1090
rect 19145 1040 19155 1060
rect 19175 1040 19185 1060
rect 19145 1010 19185 1040
rect 19145 990 19155 1010
rect 19175 990 19185 1010
rect 19145 975 19185 990
rect 19200 1210 19240 1225
rect 19200 1190 19210 1210
rect 19230 1190 19240 1210
rect 19200 1160 19240 1190
rect 19200 1140 19210 1160
rect 19230 1140 19240 1160
rect 19200 1110 19240 1140
rect 19200 1090 19210 1110
rect 19230 1090 19240 1110
rect 19200 1060 19240 1090
rect 19200 1040 19210 1060
rect 19230 1040 19240 1060
rect 19200 1010 19240 1040
rect 19200 990 19210 1010
rect 19230 990 19240 1010
rect 19200 975 19240 990
rect 19255 1210 19295 1225
rect 19255 1190 19265 1210
rect 19285 1190 19295 1210
rect 19255 1160 19295 1190
rect 19255 1140 19265 1160
rect 19285 1140 19295 1160
rect 19255 1110 19295 1140
rect 19255 1090 19265 1110
rect 19285 1090 19295 1110
rect 19255 1060 19295 1090
rect 19255 1040 19265 1060
rect 19285 1040 19295 1060
rect 19255 1010 19295 1040
rect 19255 990 19265 1010
rect 19285 990 19295 1010
rect 19255 975 19295 990
rect 19310 1210 19350 1225
rect 19310 1190 19320 1210
rect 19340 1190 19350 1210
rect 19310 1160 19350 1190
rect 19310 1140 19320 1160
rect 19340 1140 19350 1160
rect 19310 1110 19350 1140
rect 19310 1090 19320 1110
rect 19340 1090 19350 1110
rect 19310 1060 19350 1090
rect 19310 1040 19320 1060
rect 19340 1040 19350 1060
rect 19310 1010 19350 1040
rect 19310 990 19320 1010
rect 19340 990 19350 1010
rect 19310 975 19350 990
rect 19365 1210 19405 1225
rect 19365 1190 19375 1210
rect 19395 1190 19405 1210
rect 19365 1160 19405 1190
rect 19365 1140 19375 1160
rect 19395 1140 19405 1160
rect 19365 1110 19405 1140
rect 19365 1090 19375 1110
rect 19395 1090 19405 1110
rect 19365 1060 19405 1090
rect 19365 1040 19375 1060
rect 19395 1040 19405 1060
rect 19365 1010 19405 1040
rect 19365 990 19375 1010
rect 19395 990 19405 1010
rect 19365 975 19405 990
rect 19420 1210 19460 1225
rect 19420 1190 19430 1210
rect 19450 1190 19460 1210
rect 19420 1160 19460 1190
rect 19420 1140 19430 1160
rect 19450 1140 19460 1160
rect 19420 1110 19460 1140
rect 19420 1090 19430 1110
rect 19450 1090 19460 1110
rect 19420 1060 19460 1090
rect 19420 1040 19430 1060
rect 19450 1040 19460 1060
rect 19420 1010 19460 1040
rect 19420 990 19430 1010
rect 19450 990 19460 1010
rect 19420 975 19460 990
rect 19475 1210 19515 1225
rect 19475 1190 19485 1210
rect 19505 1190 19515 1210
rect 19475 1160 19515 1190
rect 19475 1140 19485 1160
rect 19505 1140 19515 1160
rect 19475 1110 19515 1140
rect 19475 1090 19485 1110
rect 19505 1090 19515 1110
rect 19475 1060 19515 1090
rect 19475 1040 19485 1060
rect 19505 1040 19515 1060
rect 19475 1010 19515 1040
rect 19475 990 19485 1010
rect 19505 990 19515 1010
rect 19475 975 19515 990
rect 19530 1210 19570 1225
rect 19530 1190 19540 1210
rect 19560 1190 19570 1210
rect 19530 1160 19570 1190
rect 19530 1140 19540 1160
rect 19560 1140 19570 1160
rect 19530 1110 19570 1140
rect 19530 1090 19540 1110
rect 19560 1090 19570 1110
rect 19530 1060 19570 1090
rect 19530 1040 19540 1060
rect 19560 1040 19570 1060
rect 19530 1010 19570 1040
rect 19530 990 19540 1010
rect 19560 990 19570 1010
rect 19530 975 19570 990
rect 19585 1210 19625 1225
rect 19585 1190 19595 1210
rect 19615 1190 19625 1210
rect 19585 1160 19625 1190
rect 19585 1140 19595 1160
rect 19615 1140 19625 1160
rect 19585 1110 19625 1140
rect 19585 1090 19595 1110
rect 19615 1090 19625 1110
rect 19585 1060 19625 1090
rect 19585 1040 19595 1060
rect 19615 1040 19625 1060
rect 19585 1010 19625 1040
rect 19585 990 19595 1010
rect 19615 990 19625 1010
rect 19585 975 19625 990
rect 19640 1210 19680 1225
rect 19640 1190 19650 1210
rect 19670 1190 19680 1210
rect 19640 1160 19680 1190
rect 19640 1140 19650 1160
rect 19670 1140 19680 1160
rect 19640 1110 19680 1140
rect 19640 1090 19650 1110
rect 19670 1090 19680 1110
rect 19640 1060 19680 1090
rect 19640 1040 19650 1060
rect 19670 1040 19680 1060
rect 19640 1010 19680 1040
rect 19640 990 19650 1010
rect 19670 990 19680 1010
rect 19640 975 19680 990
rect 19695 1210 19735 1225
rect 19695 1190 19705 1210
rect 19725 1190 19735 1210
rect 19695 1160 19735 1190
rect 19695 1140 19705 1160
rect 19725 1140 19735 1160
rect 19695 1110 19735 1140
rect 19695 1090 19705 1110
rect 19725 1090 19735 1110
rect 19695 1060 19735 1090
rect 19695 1040 19705 1060
rect 19725 1040 19735 1060
rect 19695 1010 19735 1040
rect 19695 990 19705 1010
rect 19725 990 19735 1010
rect 19695 975 19735 990
rect 19750 1210 19790 1225
rect 19750 1190 19760 1210
rect 19780 1190 19790 1210
rect 19750 1160 19790 1190
rect 19750 1140 19760 1160
rect 19780 1140 19790 1160
rect 19750 1110 19790 1140
rect 19750 1090 19760 1110
rect 19780 1090 19790 1110
rect 19750 1060 19790 1090
rect 19750 1040 19760 1060
rect 19780 1040 19790 1060
rect 19750 1010 19790 1040
rect 19750 990 19760 1010
rect 19780 990 19790 1010
rect 19750 975 19790 990
rect 19805 1210 19845 1225
rect 19805 1190 19815 1210
rect 19835 1190 19845 1210
rect 19805 1160 19845 1190
rect 19805 1140 19815 1160
rect 19835 1140 19845 1160
rect 19805 1110 19845 1140
rect 19805 1090 19815 1110
rect 19835 1090 19845 1110
rect 19805 1060 19845 1090
rect 19805 1040 19815 1060
rect 19835 1040 19845 1060
rect 19805 1010 19845 1040
rect 19805 990 19815 1010
rect 19835 990 19845 1010
rect 19805 975 19845 990
rect 19860 1210 19900 1225
rect 19860 1190 19870 1210
rect 19890 1190 19900 1210
rect 19860 1160 19900 1190
rect 19860 1140 19870 1160
rect 19890 1140 19900 1160
rect 19860 1110 19900 1140
rect 19860 1090 19870 1110
rect 19890 1090 19900 1110
rect 19860 1060 19900 1090
rect 19860 1040 19870 1060
rect 19890 1040 19900 1060
rect 19860 1010 19900 1040
rect 19860 990 19870 1010
rect 19890 990 19900 1010
rect 19860 975 19900 990
rect 19915 1210 19955 1225
rect 19915 1190 19925 1210
rect 19945 1190 19955 1210
rect 19915 1160 19955 1190
rect 19915 1140 19925 1160
rect 19945 1140 19955 1160
rect 19915 1110 19955 1140
rect 19915 1090 19925 1110
rect 19945 1090 19955 1110
rect 19915 1060 19955 1090
rect 19915 1040 19925 1060
rect 19945 1040 19955 1060
rect 19915 1010 19955 1040
rect 19915 990 19925 1010
rect 19945 990 19955 1010
rect 19915 975 19955 990
rect 19970 1210 20010 1225
rect 19970 1190 19980 1210
rect 20000 1190 20010 1210
rect 19970 1160 20010 1190
rect 19970 1140 19980 1160
rect 20000 1140 20010 1160
rect 19970 1110 20010 1140
rect 19970 1090 19980 1110
rect 20000 1090 20010 1110
rect 19970 1060 20010 1090
rect 19970 1040 19980 1060
rect 20000 1040 20010 1060
rect 19970 1010 20010 1040
rect 19970 990 19980 1010
rect 20000 990 20010 1010
rect 19970 975 20010 990
rect 20025 1210 20065 1225
rect 20025 1190 20035 1210
rect 20055 1190 20065 1210
rect 20025 1160 20065 1190
rect 20025 1140 20035 1160
rect 20055 1140 20065 1160
rect 20025 1110 20065 1140
rect 20025 1090 20035 1110
rect 20055 1090 20065 1110
rect 20025 1060 20065 1090
rect 20025 1040 20035 1060
rect 20055 1040 20065 1060
rect 20025 1010 20065 1040
rect 20025 990 20035 1010
rect 20055 990 20065 1010
rect 20025 975 20065 990
rect 20080 1210 20120 1225
rect 20080 1190 20090 1210
rect 20110 1190 20120 1210
rect 20080 1160 20120 1190
rect 20080 1140 20090 1160
rect 20110 1140 20120 1160
rect 20080 1110 20120 1140
rect 20080 1090 20090 1110
rect 20110 1090 20120 1110
rect 20080 1060 20120 1090
rect 20080 1040 20090 1060
rect 20110 1040 20120 1060
rect 20080 1010 20120 1040
rect 20545 1165 20585 1180
rect 20545 1145 20555 1165
rect 20575 1145 20585 1165
rect 20545 1115 20585 1145
rect 20545 1095 20555 1115
rect 20575 1095 20585 1115
rect 20545 1065 20585 1095
rect 20545 1045 20555 1065
rect 20575 1045 20585 1065
rect 20545 1030 20585 1045
rect 20600 1165 20640 1180
rect 20600 1145 20610 1165
rect 20630 1145 20640 1165
rect 20600 1115 20640 1145
rect 20600 1095 20610 1115
rect 20630 1095 20640 1115
rect 20600 1065 20640 1095
rect 20600 1045 20610 1065
rect 20630 1045 20640 1065
rect 20600 1030 20640 1045
rect 20655 1165 20695 1180
rect 20655 1145 20665 1165
rect 20685 1145 20695 1165
rect 20655 1115 20695 1145
rect 20655 1095 20665 1115
rect 20685 1095 20695 1115
rect 20655 1065 20695 1095
rect 20655 1045 20665 1065
rect 20685 1045 20695 1065
rect 20655 1030 20695 1045
rect 20710 1165 20750 1180
rect 20710 1145 20720 1165
rect 20740 1145 20750 1165
rect 20710 1115 20750 1145
rect 20710 1095 20720 1115
rect 20740 1095 20750 1115
rect 20710 1065 20750 1095
rect 20710 1045 20720 1065
rect 20740 1045 20750 1065
rect 20710 1030 20750 1045
rect 20765 1165 20805 1180
rect 20765 1145 20775 1165
rect 20795 1145 20805 1165
rect 20765 1115 20805 1145
rect 20765 1095 20775 1115
rect 20795 1095 20805 1115
rect 20765 1065 20805 1095
rect 20765 1045 20775 1065
rect 20795 1045 20805 1065
rect 20765 1030 20805 1045
rect 20080 990 20090 1010
rect 20110 990 20120 1010
rect 20080 975 20120 990
rect 2995 865 3035 880
rect 2995 845 3005 865
rect 3025 845 3035 865
rect 2995 815 3035 845
rect 2995 795 3005 815
rect 3025 795 3035 815
rect 2995 780 3035 795
rect 3085 865 3125 880
rect 3085 845 3095 865
rect 3115 845 3125 865
rect 3085 815 3125 845
rect 3085 795 3095 815
rect 3115 795 3125 815
rect 3085 780 3125 795
rect 3175 865 3215 880
rect 3175 845 3185 865
rect 3205 845 3215 865
rect 3175 815 3215 845
rect 3175 795 3185 815
rect 3205 795 3215 815
rect 3175 780 3215 795
rect 3265 865 3305 880
rect 3265 845 3275 865
rect 3295 845 3305 865
rect 3265 815 3305 845
rect 3265 795 3275 815
rect 3295 795 3305 815
rect 3265 780 3305 795
rect 3355 865 3395 880
rect 3355 845 3365 865
rect 3385 845 3395 865
rect 3355 815 3395 845
rect 3355 795 3365 815
rect 3385 795 3395 815
rect 3355 780 3395 795
rect 3445 865 3485 880
rect 3445 845 3455 865
rect 3475 845 3485 865
rect 3445 815 3485 845
rect 3445 795 3455 815
rect 3475 795 3485 815
rect 3445 780 3485 795
rect 3535 865 3575 880
rect 3535 845 3545 865
rect 3565 845 3575 865
rect 3535 815 3575 845
rect 3535 795 3545 815
rect 3565 795 3575 815
rect 3535 780 3575 795
rect 3625 865 3665 880
rect 3625 845 3635 865
rect 3655 845 3665 865
rect 3625 815 3665 845
rect 3625 795 3635 815
rect 3655 795 3665 815
rect 3625 780 3665 795
rect 3715 865 3755 880
rect 3715 845 3725 865
rect 3745 845 3755 865
rect 3715 815 3755 845
rect 3715 795 3725 815
rect 3745 795 3755 815
rect 3715 780 3755 795
rect 3805 865 3845 880
rect 3805 845 3815 865
rect 3835 845 3845 865
rect 3805 815 3845 845
rect 3805 795 3815 815
rect 3835 795 3845 815
rect 3805 780 3845 795
rect 3895 865 3935 880
rect 3895 845 3905 865
rect 3925 845 3935 865
rect 3895 815 3935 845
rect 3895 795 3905 815
rect 3925 795 3935 815
rect 3895 780 3935 795
rect 3985 865 4025 880
rect 3985 845 3995 865
rect 4015 845 4025 865
rect 3985 815 4025 845
rect 3985 795 3995 815
rect 4015 795 4025 815
rect 3985 780 4025 795
rect 4075 865 4115 880
rect 4075 845 4085 865
rect 4105 845 4115 865
rect 4075 815 4115 845
rect 4075 795 4085 815
rect 4105 795 4115 815
rect 4075 780 4115 795
rect 4165 865 4205 880
rect 4165 845 4175 865
rect 4195 845 4205 865
rect 4165 815 4205 845
rect 4165 795 4175 815
rect 4195 795 4205 815
rect 4165 780 4205 795
rect 4255 865 4295 880
rect 4255 845 4265 865
rect 4285 845 4295 865
rect 4255 815 4295 845
rect 4255 795 4265 815
rect 4285 795 4295 815
rect 4255 780 4295 795
rect 4345 865 4385 880
rect 4345 845 4355 865
rect 4375 845 4385 865
rect 4345 815 4385 845
rect 4345 795 4355 815
rect 4375 795 4385 815
rect 4345 780 4385 795
rect 4435 865 4475 880
rect 4435 845 4445 865
rect 4465 845 4475 865
rect 4435 815 4475 845
rect 4435 795 4445 815
rect 4465 795 4475 815
rect 4435 780 4475 795
rect 4525 865 4565 880
rect 4525 845 4535 865
rect 4555 845 4565 865
rect 4525 815 4565 845
rect 4525 795 4535 815
rect 4555 795 4565 815
rect 4525 780 4565 795
rect 4615 865 4655 880
rect 4615 845 4625 865
rect 4645 845 4655 865
rect 4615 815 4655 845
rect 4615 795 4625 815
rect 4645 795 4655 815
rect 4615 780 4655 795
rect 4705 865 4745 880
rect 4705 845 4715 865
rect 4735 845 4745 865
rect 4705 815 4745 845
rect 4705 795 4715 815
rect 4735 795 4745 815
rect 4705 780 4745 795
rect 4795 865 4835 880
rect 4795 845 4805 865
rect 4825 845 4835 865
rect 4795 815 4835 845
rect 4795 795 4805 815
rect 4825 795 4835 815
rect 4795 780 4835 795
rect 4885 865 4925 880
rect 4885 845 4895 865
rect 4915 845 4925 865
rect 4885 815 4925 845
rect 4885 795 4895 815
rect 4915 795 4925 815
rect 4885 780 4925 795
rect 4975 865 5015 880
rect 4975 845 4985 865
rect 5005 845 5015 865
rect 4975 815 5015 845
rect 4975 795 4985 815
rect 5005 795 5015 815
rect 4975 780 5015 795
rect 9275 -745 9315 -730
rect 9275 -765 9285 -745
rect 9305 -765 9315 -745
rect 9275 -790 9315 -765
rect 9275 -810 9285 -790
rect 9305 -810 9315 -790
rect 9275 -835 9315 -810
rect 9275 -855 9285 -835
rect 9305 -855 9315 -835
rect 9275 -885 9315 -855
rect 9275 -905 9285 -885
rect 9305 -905 9315 -885
rect 9275 -930 9315 -905
rect 9275 -950 9285 -930
rect 9305 -950 9315 -930
rect 9275 -975 9315 -950
rect 9275 -995 9285 -975
rect 9305 -995 9315 -975
rect 9275 -1010 9315 -995
rect 9375 -745 9415 -730
rect 9375 -765 9385 -745
rect 9405 -765 9415 -745
rect 9375 -790 9415 -765
rect 9375 -810 9385 -790
rect 9405 -810 9415 -790
rect 9375 -835 9415 -810
rect 9375 -855 9385 -835
rect 9405 -855 9415 -835
rect 9375 -885 9415 -855
rect 9375 -905 9385 -885
rect 9405 -905 9415 -885
rect 9375 -930 9415 -905
rect 9375 -950 9385 -930
rect 9405 -950 9415 -930
rect 9375 -975 9415 -950
rect 9375 -995 9385 -975
rect 9405 -995 9415 -975
rect 9375 -1010 9415 -995
rect 9475 -745 9515 -730
rect 9475 -765 9485 -745
rect 9505 -765 9515 -745
rect 9475 -790 9515 -765
rect 9475 -810 9485 -790
rect 9505 -810 9515 -790
rect 9475 -835 9515 -810
rect 9475 -855 9485 -835
rect 9505 -855 9515 -835
rect 9475 -885 9515 -855
rect 9475 -905 9485 -885
rect 9505 -905 9515 -885
rect 9475 -930 9515 -905
rect 9475 -950 9485 -930
rect 9505 -950 9515 -930
rect 9475 -975 9515 -950
rect 9475 -995 9485 -975
rect 9505 -995 9515 -975
rect 9475 -1010 9515 -995
rect 9575 -745 9615 -730
rect 9575 -765 9585 -745
rect 9605 -765 9615 -745
rect 9575 -790 9615 -765
rect 9575 -810 9585 -790
rect 9605 -810 9615 -790
rect 9575 -835 9615 -810
rect 9575 -855 9585 -835
rect 9605 -855 9615 -835
rect 9575 -885 9615 -855
rect 9575 -905 9585 -885
rect 9605 -905 9615 -885
rect 9575 -930 9615 -905
rect 9575 -950 9585 -930
rect 9605 -950 9615 -930
rect 9575 -975 9615 -950
rect 9575 -995 9585 -975
rect 9605 -995 9615 -975
rect 9575 -1010 9615 -995
rect 9675 -745 9715 -730
rect 9675 -765 9685 -745
rect 9705 -765 9715 -745
rect 9675 -790 9715 -765
rect 9675 -810 9685 -790
rect 9705 -810 9715 -790
rect 9675 -835 9715 -810
rect 9675 -855 9685 -835
rect 9705 -855 9715 -835
rect 9675 -885 9715 -855
rect 9675 -905 9685 -885
rect 9705 -905 9715 -885
rect 9675 -930 9715 -905
rect 9675 -950 9685 -930
rect 9705 -950 9715 -930
rect 9675 -975 9715 -950
rect 9675 -995 9685 -975
rect 9705 -995 9715 -975
rect 9675 -1010 9715 -995
rect 9775 -745 9815 -730
rect 9775 -765 9785 -745
rect 9805 -765 9815 -745
rect 9775 -790 9815 -765
rect 9775 -810 9785 -790
rect 9805 -810 9815 -790
rect 9775 -835 9815 -810
rect 9775 -855 9785 -835
rect 9805 -855 9815 -835
rect 9775 -885 9815 -855
rect 9775 -905 9785 -885
rect 9805 -905 9815 -885
rect 9775 -930 9815 -905
rect 9775 -950 9785 -930
rect 9805 -950 9815 -930
rect 9775 -975 9815 -950
rect 9775 -995 9785 -975
rect 9805 -995 9815 -975
rect 9775 -1010 9815 -995
rect 9875 -745 9915 -730
rect 9875 -765 9885 -745
rect 9905 -765 9915 -745
rect 9875 -790 9915 -765
rect 9875 -810 9885 -790
rect 9905 -810 9915 -790
rect 9875 -835 9915 -810
rect 9875 -855 9885 -835
rect 9905 -855 9915 -835
rect 9875 -885 9915 -855
rect 9875 -905 9885 -885
rect 9905 -905 9915 -885
rect 9875 -930 9915 -905
rect 9875 -950 9885 -930
rect 9905 -950 9915 -930
rect 9875 -975 9915 -950
rect 9875 -995 9885 -975
rect 9905 -995 9915 -975
rect 9875 -1010 9915 -995
rect 9975 -745 10015 -730
rect 9975 -765 9985 -745
rect 10005 -765 10015 -745
rect 9975 -790 10015 -765
rect 9975 -810 9985 -790
rect 10005 -810 10015 -790
rect 9975 -835 10015 -810
rect 9975 -855 9985 -835
rect 10005 -855 10015 -835
rect 9975 -885 10015 -855
rect 9975 -905 9985 -885
rect 10005 -905 10015 -885
rect 9975 -930 10015 -905
rect 9975 -950 9985 -930
rect 10005 -950 10015 -930
rect 9975 -975 10015 -950
rect 9975 -995 9985 -975
rect 10005 -995 10015 -975
rect 9975 -1010 10015 -995
rect 10075 -745 10115 -730
rect 10075 -765 10085 -745
rect 10105 -765 10115 -745
rect 10075 -790 10115 -765
rect 10075 -810 10085 -790
rect 10105 -810 10115 -790
rect 10075 -835 10115 -810
rect 10075 -855 10085 -835
rect 10105 -855 10115 -835
rect 10075 -885 10115 -855
rect 10075 -905 10085 -885
rect 10105 -905 10115 -885
rect 10075 -930 10115 -905
rect 10075 -950 10085 -930
rect 10105 -950 10115 -930
rect 10075 -975 10115 -950
rect 10075 -995 10085 -975
rect 10105 -995 10115 -975
rect 10075 -1010 10115 -995
rect 10175 -745 10215 -730
rect 10175 -765 10185 -745
rect 10205 -765 10215 -745
rect 10175 -790 10215 -765
rect 10175 -810 10185 -790
rect 10205 -810 10215 -790
rect 10175 -835 10215 -810
rect 10175 -855 10185 -835
rect 10205 -855 10215 -835
rect 10175 -885 10215 -855
rect 10175 -905 10185 -885
rect 10205 -905 10215 -885
rect 10175 -930 10215 -905
rect 10175 -950 10185 -930
rect 10205 -950 10215 -930
rect 10175 -975 10215 -950
rect 10175 -995 10185 -975
rect 10205 -995 10215 -975
rect 10175 -1010 10215 -995
rect 10275 -745 10315 -730
rect 10275 -765 10285 -745
rect 10305 -765 10315 -745
rect 10275 -790 10315 -765
rect 10275 -810 10285 -790
rect 10305 -810 10315 -790
rect 10275 -835 10315 -810
rect 10275 -855 10285 -835
rect 10305 -855 10315 -835
rect 10275 -885 10315 -855
rect 10275 -905 10285 -885
rect 10305 -905 10315 -885
rect 10275 -930 10315 -905
rect 10275 -950 10285 -930
rect 10305 -950 10315 -930
rect 10275 -975 10315 -950
rect 10275 -995 10285 -975
rect 10305 -995 10315 -975
rect 10275 -1010 10315 -995
rect 10375 -745 10415 -730
rect 10375 -765 10385 -745
rect 10405 -765 10415 -745
rect 10375 -790 10415 -765
rect 10375 -810 10385 -790
rect 10405 -810 10415 -790
rect 10375 -835 10415 -810
rect 10375 -855 10385 -835
rect 10405 -855 10415 -835
rect 10375 -885 10415 -855
rect 10375 -905 10385 -885
rect 10405 -905 10415 -885
rect 10375 -930 10415 -905
rect 10375 -950 10385 -930
rect 10405 -950 10415 -930
rect 10375 -975 10415 -950
rect 10375 -995 10385 -975
rect 10405 -995 10415 -975
rect 10375 -1010 10415 -995
rect 10475 -745 10515 -730
rect 10475 -765 10485 -745
rect 10505 -765 10515 -745
rect 10475 -790 10515 -765
rect 10475 -810 10485 -790
rect 10505 -810 10515 -790
rect 10475 -835 10515 -810
rect 10475 -855 10485 -835
rect 10505 -855 10515 -835
rect 10475 -885 10515 -855
rect 10475 -905 10485 -885
rect 10505 -905 10515 -885
rect 10475 -930 10515 -905
rect 10475 -950 10485 -930
rect 10505 -950 10515 -930
rect 10475 -975 10515 -950
rect 10475 -995 10485 -975
rect 10505 -995 10515 -975
rect 10475 -1010 10515 -995
<< pdiff >>
rect 2995 2915 3035 2930
rect 2995 2895 3005 2915
rect 3025 2895 3035 2915
rect 2995 2865 3035 2895
rect 2995 2845 3005 2865
rect 3025 2845 3035 2865
rect 2995 2830 3035 2845
rect 3085 2915 3125 2930
rect 3085 2895 3095 2915
rect 3115 2895 3125 2915
rect 3085 2865 3125 2895
rect 3085 2845 3095 2865
rect 3115 2845 3125 2865
rect 3085 2830 3125 2845
rect 3175 2915 3215 2930
rect 3175 2895 3185 2915
rect 3205 2895 3215 2915
rect 3175 2865 3215 2895
rect 3175 2845 3185 2865
rect 3205 2845 3215 2865
rect 3175 2830 3215 2845
rect 3265 2915 3305 2930
rect 3265 2895 3275 2915
rect 3295 2895 3305 2915
rect 3265 2865 3305 2895
rect 3265 2845 3275 2865
rect 3295 2845 3305 2865
rect 3265 2830 3305 2845
rect 3355 2915 3395 2930
rect 3355 2895 3365 2915
rect 3385 2895 3395 2915
rect 3355 2865 3395 2895
rect 3355 2845 3365 2865
rect 3385 2845 3395 2865
rect 3355 2830 3395 2845
rect 3445 2915 3485 2930
rect 3445 2895 3455 2915
rect 3475 2895 3485 2915
rect 3445 2865 3485 2895
rect 3445 2845 3455 2865
rect 3475 2845 3485 2865
rect 3445 2830 3485 2845
rect 3535 2915 3575 2930
rect 3535 2895 3545 2915
rect 3565 2895 3575 2915
rect 3535 2865 3575 2895
rect 3535 2845 3545 2865
rect 3565 2845 3575 2865
rect 3535 2830 3575 2845
rect 3625 2915 3665 2930
rect 3625 2895 3635 2915
rect 3655 2895 3665 2915
rect 3625 2865 3665 2895
rect 3625 2845 3635 2865
rect 3655 2845 3665 2865
rect 3625 2830 3665 2845
rect 3715 2915 3755 2930
rect 3715 2895 3725 2915
rect 3745 2895 3755 2915
rect 3715 2865 3755 2895
rect 3715 2845 3725 2865
rect 3745 2845 3755 2865
rect 3715 2830 3755 2845
rect 3805 2915 3845 2930
rect 3805 2895 3815 2915
rect 3835 2895 3845 2915
rect 3805 2865 3845 2895
rect 3805 2845 3815 2865
rect 3835 2845 3845 2865
rect 3805 2830 3845 2845
rect 3895 2915 3935 2930
rect 3895 2895 3905 2915
rect 3925 2895 3935 2915
rect 3895 2865 3935 2895
rect 3895 2845 3905 2865
rect 3925 2845 3935 2865
rect 3895 2830 3935 2845
rect 3985 2915 4025 2930
rect 3985 2895 3995 2915
rect 4015 2895 4025 2915
rect 3985 2865 4025 2895
rect 3985 2845 3995 2865
rect 4015 2845 4025 2865
rect 3985 2830 4025 2845
rect 4075 2915 4115 2930
rect 4075 2895 4085 2915
rect 4105 2895 4115 2915
rect 4075 2865 4115 2895
rect 4075 2845 4085 2865
rect 4105 2845 4115 2865
rect 4075 2830 4115 2845
rect 4165 2915 4205 2930
rect 4165 2895 4175 2915
rect 4195 2895 4205 2915
rect 4165 2865 4205 2895
rect 4165 2845 4175 2865
rect 4195 2845 4205 2865
rect 4165 2830 4205 2845
rect 4255 2915 4295 2930
rect 4255 2895 4265 2915
rect 4285 2895 4295 2915
rect 4255 2865 4295 2895
rect 4255 2845 4265 2865
rect 4285 2845 4295 2865
rect 4255 2830 4295 2845
rect 4345 2915 4385 2930
rect 4345 2895 4355 2915
rect 4375 2895 4385 2915
rect 4345 2865 4385 2895
rect 4345 2845 4355 2865
rect 4375 2845 4385 2865
rect 4345 2830 4385 2845
rect 4435 2915 4475 2930
rect 4435 2895 4445 2915
rect 4465 2895 4475 2915
rect 4435 2865 4475 2895
rect 4435 2845 4445 2865
rect 4465 2845 4475 2865
rect 4435 2830 4475 2845
rect 4525 2915 4565 2930
rect 4525 2895 4535 2915
rect 4555 2895 4565 2915
rect 4525 2865 4565 2895
rect 4525 2845 4535 2865
rect 4555 2845 4565 2865
rect 4525 2830 4565 2845
rect 4615 2915 4655 2930
rect 4615 2895 4625 2915
rect 4645 2895 4655 2915
rect 4615 2865 4655 2895
rect 4615 2845 4625 2865
rect 4645 2845 4655 2865
rect 4615 2830 4655 2845
rect 4705 2915 4745 2930
rect 4705 2895 4715 2915
rect 4735 2895 4745 2915
rect 4705 2865 4745 2895
rect 4705 2845 4715 2865
rect 4735 2845 4745 2865
rect 4705 2830 4745 2845
rect 4795 2915 4835 2930
rect 4795 2895 4805 2915
rect 4825 2895 4835 2915
rect 4795 2865 4835 2895
rect 4795 2845 4805 2865
rect 4825 2845 4835 2865
rect 4795 2830 4835 2845
rect 4885 2915 4925 2930
rect 4885 2895 4895 2915
rect 4915 2895 4925 2915
rect 4885 2865 4925 2895
rect 4885 2845 4895 2865
rect 4915 2845 4925 2865
rect 4885 2830 4925 2845
rect 4975 2915 5015 2930
rect 4975 2895 4985 2915
rect 5005 2895 5015 2915
rect 4975 2865 5015 2895
rect 4975 2845 4985 2865
rect 5005 2845 5015 2865
rect 4975 2830 5015 2845
rect 3175 2685 3215 2700
rect 3175 2665 3185 2685
rect 3205 2665 3215 2685
rect 3175 2635 3215 2665
rect 3175 2615 3185 2635
rect 3205 2615 3215 2635
rect 3175 2585 3215 2615
rect 3175 2565 3185 2585
rect 3205 2565 3215 2585
rect 3175 2535 3215 2565
rect 3175 2515 3185 2535
rect 3205 2515 3215 2535
rect 3175 2485 3215 2515
rect 3175 2465 3185 2485
rect 3205 2465 3215 2485
rect 3175 2435 3215 2465
rect 3175 2415 3185 2435
rect 3205 2415 3215 2435
rect 3175 2400 3215 2415
rect 3265 2685 3305 2700
rect 3265 2665 3275 2685
rect 3295 2665 3305 2685
rect 3265 2635 3305 2665
rect 3265 2615 3275 2635
rect 3295 2615 3305 2635
rect 3265 2585 3305 2615
rect 3265 2565 3275 2585
rect 3295 2565 3305 2585
rect 3265 2535 3305 2565
rect 3265 2515 3275 2535
rect 3295 2515 3305 2535
rect 3265 2485 3305 2515
rect 3265 2465 3275 2485
rect 3295 2465 3305 2485
rect 3265 2435 3305 2465
rect 3265 2415 3275 2435
rect 3295 2415 3305 2435
rect 3265 2400 3305 2415
rect 3355 2685 3395 2700
rect 3355 2665 3365 2685
rect 3385 2665 3395 2685
rect 3355 2635 3395 2665
rect 3355 2615 3365 2635
rect 3385 2615 3395 2635
rect 3355 2585 3395 2615
rect 3355 2565 3365 2585
rect 3385 2565 3395 2585
rect 3355 2535 3395 2565
rect 3355 2515 3365 2535
rect 3385 2515 3395 2535
rect 3355 2485 3395 2515
rect 3355 2465 3365 2485
rect 3385 2465 3395 2485
rect 3355 2435 3395 2465
rect 3355 2415 3365 2435
rect 3385 2415 3395 2435
rect 3355 2400 3395 2415
rect 3445 2685 3485 2700
rect 3445 2665 3455 2685
rect 3475 2665 3485 2685
rect 3445 2635 3485 2665
rect 3445 2615 3455 2635
rect 3475 2615 3485 2635
rect 3445 2585 3485 2615
rect 3445 2565 3455 2585
rect 3475 2565 3485 2585
rect 3445 2535 3485 2565
rect 3445 2515 3455 2535
rect 3475 2515 3485 2535
rect 3445 2485 3485 2515
rect 3445 2465 3455 2485
rect 3475 2465 3485 2485
rect 3445 2435 3485 2465
rect 3445 2415 3455 2435
rect 3475 2415 3485 2435
rect 3445 2400 3485 2415
rect 3535 2685 3575 2700
rect 3535 2665 3545 2685
rect 3565 2665 3575 2685
rect 3535 2635 3575 2665
rect 3535 2615 3545 2635
rect 3565 2615 3575 2635
rect 3535 2585 3575 2615
rect 3535 2565 3545 2585
rect 3565 2565 3575 2585
rect 3535 2535 3575 2565
rect 3535 2515 3545 2535
rect 3565 2515 3575 2535
rect 3535 2485 3575 2515
rect 3535 2465 3545 2485
rect 3565 2465 3575 2485
rect 3535 2435 3575 2465
rect 3535 2415 3545 2435
rect 3565 2415 3575 2435
rect 3535 2400 3575 2415
rect 3625 2685 3665 2700
rect 3625 2665 3635 2685
rect 3655 2665 3665 2685
rect 3625 2635 3665 2665
rect 3625 2615 3635 2635
rect 3655 2615 3665 2635
rect 3625 2585 3665 2615
rect 3625 2565 3635 2585
rect 3655 2565 3665 2585
rect 3625 2535 3665 2565
rect 3625 2515 3635 2535
rect 3655 2515 3665 2535
rect 3625 2485 3665 2515
rect 3625 2465 3635 2485
rect 3655 2465 3665 2485
rect 3625 2435 3665 2465
rect 3625 2415 3635 2435
rect 3655 2415 3665 2435
rect 3625 2400 3665 2415
rect 3715 2685 3755 2700
rect 3715 2665 3725 2685
rect 3745 2665 3755 2685
rect 3715 2635 3755 2665
rect 3715 2615 3725 2635
rect 3745 2615 3755 2635
rect 3715 2585 3755 2615
rect 3715 2565 3725 2585
rect 3745 2565 3755 2585
rect 3715 2535 3755 2565
rect 3715 2515 3725 2535
rect 3745 2515 3755 2535
rect 3715 2485 3755 2515
rect 3715 2465 3725 2485
rect 3745 2465 3755 2485
rect 3715 2435 3755 2465
rect 3715 2415 3725 2435
rect 3745 2415 3755 2435
rect 3715 2400 3755 2415
rect 3805 2685 3845 2700
rect 3805 2665 3815 2685
rect 3835 2665 3845 2685
rect 3805 2635 3845 2665
rect 3805 2615 3815 2635
rect 3835 2615 3845 2635
rect 3805 2585 3845 2615
rect 3805 2565 3815 2585
rect 3835 2565 3845 2585
rect 3805 2535 3845 2565
rect 3805 2515 3815 2535
rect 3835 2515 3845 2535
rect 3805 2485 3845 2515
rect 3805 2465 3815 2485
rect 3835 2465 3845 2485
rect 3805 2435 3845 2465
rect 3805 2415 3815 2435
rect 3835 2415 3845 2435
rect 3805 2400 3845 2415
rect 3895 2685 3935 2700
rect 3895 2665 3905 2685
rect 3925 2665 3935 2685
rect 3895 2635 3935 2665
rect 3895 2615 3905 2635
rect 3925 2615 3935 2635
rect 3895 2585 3935 2615
rect 3895 2565 3905 2585
rect 3925 2565 3935 2585
rect 3895 2535 3935 2565
rect 3895 2515 3905 2535
rect 3925 2515 3935 2535
rect 3895 2485 3935 2515
rect 3895 2465 3905 2485
rect 3925 2465 3935 2485
rect 3895 2435 3935 2465
rect 3895 2415 3905 2435
rect 3925 2415 3935 2435
rect 3895 2400 3935 2415
rect 3985 2685 4025 2700
rect 3985 2665 3995 2685
rect 4015 2665 4025 2685
rect 3985 2635 4025 2665
rect 3985 2615 3995 2635
rect 4015 2615 4025 2635
rect 3985 2585 4025 2615
rect 3985 2565 3995 2585
rect 4015 2565 4025 2585
rect 3985 2535 4025 2565
rect 3985 2515 3995 2535
rect 4015 2515 4025 2535
rect 3985 2485 4025 2515
rect 3985 2465 3995 2485
rect 4015 2465 4025 2485
rect 3985 2435 4025 2465
rect 3985 2415 3995 2435
rect 4015 2415 4025 2435
rect 3985 2400 4025 2415
rect 4075 2685 4115 2700
rect 4075 2665 4085 2685
rect 4105 2665 4115 2685
rect 4075 2635 4115 2665
rect 4075 2615 4085 2635
rect 4105 2615 4115 2635
rect 4075 2585 4115 2615
rect 4075 2565 4085 2585
rect 4105 2565 4115 2585
rect 4075 2535 4115 2565
rect 4075 2515 4085 2535
rect 4105 2515 4115 2535
rect 4075 2485 4115 2515
rect 4075 2465 4085 2485
rect 4105 2465 4115 2485
rect 4075 2435 4115 2465
rect 4075 2415 4085 2435
rect 4105 2415 4115 2435
rect 4075 2400 4115 2415
rect 4165 2685 4205 2700
rect 4165 2665 4175 2685
rect 4195 2665 4205 2685
rect 4165 2635 4205 2665
rect 4165 2615 4175 2635
rect 4195 2615 4205 2635
rect 4165 2585 4205 2615
rect 4165 2565 4175 2585
rect 4195 2565 4205 2585
rect 4165 2535 4205 2565
rect 4165 2515 4175 2535
rect 4195 2515 4205 2535
rect 4165 2485 4205 2515
rect 4165 2465 4175 2485
rect 4195 2465 4205 2485
rect 4165 2435 4205 2465
rect 4165 2415 4175 2435
rect 4195 2415 4205 2435
rect 4165 2400 4205 2415
rect 4255 2685 4295 2700
rect 4255 2665 4265 2685
rect 4285 2665 4295 2685
rect 4255 2635 4295 2665
rect 4255 2615 4265 2635
rect 4285 2615 4295 2635
rect 4255 2585 4295 2615
rect 4255 2565 4265 2585
rect 4285 2565 4295 2585
rect 4255 2535 4295 2565
rect 4255 2515 4265 2535
rect 4285 2515 4295 2535
rect 4255 2485 4295 2515
rect 4255 2465 4265 2485
rect 4285 2465 4295 2485
rect 4255 2435 4295 2465
rect 4255 2415 4265 2435
rect 4285 2415 4295 2435
rect 4255 2400 4295 2415
rect 4345 2685 4385 2700
rect 4345 2665 4355 2685
rect 4375 2665 4385 2685
rect 4345 2635 4385 2665
rect 4345 2615 4355 2635
rect 4375 2615 4385 2635
rect 4345 2585 4385 2615
rect 4345 2565 4355 2585
rect 4375 2565 4385 2585
rect 4345 2535 4385 2565
rect 4345 2515 4355 2535
rect 4375 2515 4385 2535
rect 4345 2485 4385 2515
rect 4345 2465 4355 2485
rect 4375 2465 4385 2485
rect 4345 2435 4385 2465
rect 4345 2415 4355 2435
rect 4375 2415 4385 2435
rect 4345 2400 4385 2415
rect 4435 2685 4475 2700
rect 4435 2665 4445 2685
rect 4465 2665 4475 2685
rect 4435 2635 4475 2665
rect 4435 2615 4445 2635
rect 4465 2615 4475 2635
rect 4435 2585 4475 2615
rect 4435 2565 4445 2585
rect 4465 2565 4475 2585
rect 4435 2535 4475 2565
rect 4435 2515 4445 2535
rect 4465 2515 4475 2535
rect 4435 2485 4475 2515
rect 4435 2465 4445 2485
rect 4465 2465 4475 2485
rect 4435 2435 4475 2465
rect 4435 2415 4445 2435
rect 4465 2415 4475 2435
rect 4435 2400 4475 2415
rect 4525 2685 4565 2700
rect 4525 2665 4535 2685
rect 4555 2665 4565 2685
rect 4525 2635 4565 2665
rect 4525 2615 4535 2635
rect 4555 2615 4565 2635
rect 4525 2585 4565 2615
rect 4525 2565 4535 2585
rect 4555 2565 4565 2585
rect 4525 2535 4565 2565
rect 4525 2515 4535 2535
rect 4555 2515 4565 2535
rect 4525 2485 4565 2515
rect 4525 2465 4535 2485
rect 4555 2465 4565 2485
rect 4525 2435 4565 2465
rect 4525 2415 4535 2435
rect 4555 2415 4565 2435
rect 4525 2400 4565 2415
rect 4615 2685 4655 2700
rect 4615 2665 4625 2685
rect 4645 2665 4655 2685
rect 4615 2635 4655 2665
rect 4615 2615 4625 2635
rect 4645 2615 4655 2635
rect 4615 2585 4655 2615
rect 4615 2565 4625 2585
rect 4645 2565 4655 2585
rect 4615 2535 4655 2565
rect 4615 2515 4625 2535
rect 4645 2515 4655 2535
rect 4615 2485 4655 2515
rect 4615 2465 4625 2485
rect 4645 2465 4655 2485
rect 4615 2435 4655 2465
rect 4615 2415 4625 2435
rect 4645 2415 4655 2435
rect 4615 2400 4655 2415
rect 4705 2685 4745 2700
rect 4705 2665 4715 2685
rect 4735 2665 4745 2685
rect 4705 2635 4745 2665
rect 4705 2615 4715 2635
rect 4735 2615 4745 2635
rect 4705 2585 4745 2615
rect 4705 2565 4715 2585
rect 4735 2565 4745 2585
rect 4705 2535 4745 2565
rect 4705 2515 4715 2535
rect 4735 2515 4745 2535
rect 4705 2485 4745 2515
rect 4705 2465 4715 2485
rect 4735 2465 4745 2485
rect 4705 2435 4745 2465
rect 4705 2415 4715 2435
rect 4735 2415 4745 2435
rect 4705 2400 4745 2415
rect 4795 2685 4835 2700
rect 4795 2665 4805 2685
rect 4825 2665 4835 2685
rect 4795 2635 4835 2665
rect 4795 2615 4805 2635
rect 4825 2615 4835 2635
rect 4795 2585 4835 2615
rect 4795 2565 4805 2585
rect 4825 2565 4835 2585
rect 4795 2535 4835 2565
rect 4795 2515 4805 2535
rect 4825 2515 4835 2535
rect 4795 2485 4835 2515
rect 4795 2465 4805 2485
rect 4825 2465 4835 2485
rect 4795 2435 4835 2465
rect 4795 2415 4805 2435
rect 4825 2415 4835 2435
rect 4795 2400 4835 2415
rect 2565 1985 2605 2000
rect 2565 1965 2575 1985
rect 2595 1965 2605 1985
rect 2565 1935 2605 1965
rect 2565 1915 2575 1935
rect 2595 1915 2605 1935
rect 2565 1900 2605 1915
rect 2620 1985 2660 2000
rect 2620 1965 2630 1985
rect 2650 1965 2660 1985
rect 2620 1935 2660 1965
rect 2620 1915 2630 1935
rect 2650 1915 2660 1935
rect 2620 1900 2660 1915
rect 2675 1985 2715 2000
rect 2675 1965 2685 1985
rect 2705 1965 2715 1985
rect 2675 1935 2715 1965
rect 2675 1915 2685 1935
rect 2705 1915 2715 1935
rect 2675 1900 2715 1915
rect 2745 1985 2785 2000
rect 2745 1965 2755 1985
rect 2775 1965 2785 1985
rect 2745 1935 2785 1965
rect 2745 1915 2755 1935
rect 2775 1915 2785 1935
rect 2745 1900 2785 1915
rect 2805 1985 2845 2000
rect 2805 1965 2815 1985
rect 2835 1965 2845 1985
rect 2805 1935 2845 1965
rect 2805 1915 2815 1935
rect 2835 1915 2845 1935
rect 2805 1900 2845 1915
rect 2865 1985 2905 2000
rect 2865 1965 2875 1985
rect 2895 1965 2905 1985
rect 2865 1935 2905 1965
rect 2865 1915 2875 1935
rect 2895 1915 2905 1935
rect 2865 1900 2905 1915
rect 2925 1985 2965 2000
rect 2925 1965 2935 1985
rect 2955 1965 2965 1985
rect 2925 1935 2965 1965
rect 2925 1915 2935 1935
rect 2955 1915 2965 1935
rect 2925 1900 2965 1915
rect 2985 1985 3025 2000
rect 2985 1965 2995 1985
rect 3015 1965 3025 1985
rect 2985 1935 3025 1965
rect 2985 1915 2995 1935
rect 3015 1915 3025 1935
rect 2985 1900 3025 1915
rect 3045 1985 3085 2000
rect 3045 1965 3055 1985
rect 3075 1965 3085 1985
rect 3045 1935 3085 1965
rect 3045 1915 3055 1935
rect 3075 1915 3085 1935
rect 3045 1900 3085 1915
rect 3105 1985 3145 2000
rect 3105 1965 3115 1985
rect 3135 1965 3145 1985
rect 3105 1935 3145 1965
rect 3105 1915 3115 1935
rect 3135 1915 3145 1935
rect 3105 1900 3145 1915
rect 3165 1985 3205 2000
rect 3165 1965 3175 1985
rect 3195 1965 3205 1985
rect 3165 1935 3205 1965
rect 3165 1915 3175 1935
rect 3195 1915 3205 1935
rect 3165 1900 3205 1915
rect 3225 1985 3265 2000
rect 3225 1965 3235 1985
rect 3255 1965 3265 1985
rect 3225 1935 3265 1965
rect 3225 1915 3235 1935
rect 3255 1915 3265 1935
rect 3225 1900 3265 1915
rect 3285 1985 3325 2000
rect 3285 1965 3295 1985
rect 3315 1965 3325 1985
rect 3285 1935 3325 1965
rect 3285 1915 3295 1935
rect 3315 1915 3325 1935
rect 3285 1900 3325 1915
rect 3345 1985 3385 2000
rect 3345 1965 3355 1985
rect 3375 1965 3385 1985
rect 3345 1935 3385 1965
rect 3345 1915 3355 1935
rect 3375 1915 3385 1935
rect 3345 1900 3385 1915
rect 3405 1985 3445 2000
rect 3405 1965 3415 1985
rect 3435 1965 3445 1985
rect 3405 1935 3445 1965
rect 3405 1915 3415 1935
rect 3435 1915 3445 1935
rect 3405 1900 3445 1915
rect 3465 1985 3505 2000
rect 3465 1965 3475 1985
rect 3495 1965 3505 1985
rect 3465 1935 3505 1965
rect 3465 1915 3475 1935
rect 3495 1915 3505 1935
rect 3465 1900 3505 1915
rect 3525 1985 3565 2000
rect 3525 1965 3535 1985
rect 3555 1965 3565 1985
rect 3525 1935 3565 1965
rect 3525 1915 3535 1935
rect 3555 1915 3565 1935
rect 3525 1900 3565 1915
rect 3585 1985 3625 2000
rect 3585 1965 3595 1985
rect 3615 1965 3625 1985
rect 3585 1935 3625 1965
rect 3585 1915 3595 1935
rect 3615 1915 3625 1935
rect 3585 1900 3625 1915
rect 3645 1985 3685 2000
rect 3645 1965 3655 1985
rect 3675 1965 3685 1985
rect 3645 1935 3685 1965
rect 3645 1915 3655 1935
rect 3675 1915 3685 1935
rect 3645 1900 3685 1915
rect 3705 1985 3745 2000
rect 3705 1965 3715 1985
rect 3735 1965 3745 1985
rect 3705 1935 3745 1965
rect 3705 1915 3715 1935
rect 3735 1915 3745 1935
rect 3705 1900 3745 1915
rect 3765 1985 3805 2000
rect 3765 1965 3775 1985
rect 3795 1965 3805 1985
rect 3765 1935 3805 1965
rect 3765 1915 3775 1935
rect 3795 1915 3805 1935
rect 3765 1900 3805 1915
rect 3825 1985 3865 2000
rect 3825 1965 3835 1985
rect 3855 1965 3865 1985
rect 3825 1935 3865 1965
rect 3825 1915 3835 1935
rect 3855 1915 3865 1935
rect 3825 1900 3865 1915
rect 3885 1985 3925 2000
rect 3885 1965 3895 1985
rect 3915 1965 3925 1985
rect 3885 1935 3925 1965
rect 3885 1915 3895 1935
rect 3915 1915 3925 1935
rect 3885 1900 3925 1915
rect 3945 1985 3985 2000
rect 4025 1985 4065 2000
rect 3945 1965 3955 1985
rect 3975 1965 3985 1985
rect 4025 1965 4035 1985
rect 4055 1965 4065 1985
rect 3945 1935 3985 1965
rect 4025 1935 4065 1965
rect 3945 1915 3955 1935
rect 3975 1915 3985 1935
rect 4025 1915 4035 1935
rect 4055 1915 4065 1935
rect 3945 1900 3985 1915
rect 4025 1900 4065 1915
rect 4085 1985 4125 2000
rect 4085 1965 4095 1985
rect 4115 1965 4125 1985
rect 4085 1935 4125 1965
rect 4085 1915 4095 1935
rect 4115 1915 4125 1935
rect 4085 1900 4125 1915
rect 4145 1985 4185 2000
rect 4145 1965 4155 1985
rect 4175 1965 4185 1985
rect 4145 1935 4185 1965
rect 4145 1915 4155 1935
rect 4175 1915 4185 1935
rect 4145 1900 4185 1915
rect 4205 1985 4245 2000
rect 4205 1965 4215 1985
rect 4235 1965 4245 1985
rect 4205 1935 4245 1965
rect 4205 1915 4215 1935
rect 4235 1915 4245 1935
rect 4205 1900 4245 1915
rect 4265 1985 4305 2000
rect 4265 1965 4275 1985
rect 4295 1965 4305 1985
rect 4265 1935 4305 1965
rect 4265 1915 4275 1935
rect 4295 1915 4305 1935
rect 4265 1900 4305 1915
rect 4325 1985 4365 2000
rect 4325 1965 4335 1985
rect 4355 1965 4365 1985
rect 4325 1935 4365 1965
rect 4325 1915 4335 1935
rect 4355 1915 4365 1935
rect 4325 1900 4365 1915
rect 4385 1985 4425 2000
rect 4385 1965 4395 1985
rect 4415 1965 4425 1985
rect 4385 1935 4425 1965
rect 4385 1915 4395 1935
rect 4415 1915 4425 1935
rect 4385 1900 4425 1915
rect 4445 1985 4485 2000
rect 4445 1965 4455 1985
rect 4475 1965 4485 1985
rect 4445 1935 4485 1965
rect 4445 1915 4455 1935
rect 4475 1915 4485 1935
rect 4445 1900 4485 1915
rect 4505 1985 4545 2000
rect 4505 1965 4515 1985
rect 4535 1965 4545 1985
rect 4505 1935 4545 1965
rect 4505 1915 4515 1935
rect 4535 1915 4545 1935
rect 4505 1900 4545 1915
rect 4565 1985 4605 2000
rect 4565 1965 4575 1985
rect 4595 1965 4605 1985
rect 4565 1935 4605 1965
rect 4565 1915 4575 1935
rect 4595 1915 4605 1935
rect 4565 1900 4605 1915
rect 4625 1985 4665 2000
rect 4625 1965 4635 1985
rect 4655 1965 4665 1985
rect 4625 1935 4665 1965
rect 4625 1915 4635 1935
rect 4655 1915 4665 1935
rect 4625 1900 4665 1915
rect 4685 1985 4725 2000
rect 4685 1965 4695 1985
rect 4715 1965 4725 1985
rect 4685 1935 4725 1965
rect 4685 1915 4695 1935
rect 4715 1915 4725 1935
rect 4685 1900 4725 1915
rect 4745 1985 4785 2000
rect 4745 1965 4755 1985
rect 4775 1965 4785 1985
rect 4745 1935 4785 1965
rect 4745 1915 4755 1935
rect 4775 1915 4785 1935
rect 4745 1900 4785 1915
rect 4805 1985 4845 2000
rect 4805 1965 4815 1985
rect 4835 1965 4845 1985
rect 4805 1935 4845 1965
rect 4805 1915 4815 1935
rect 4835 1915 4845 1935
rect 4805 1900 4845 1915
rect 4865 1985 4905 2000
rect 4865 1965 4875 1985
rect 4895 1965 4905 1985
rect 4865 1935 4905 1965
rect 4865 1915 4875 1935
rect 4895 1915 4905 1935
rect 4865 1900 4905 1915
rect 4925 1985 4965 2000
rect 4925 1965 4935 1985
rect 4955 1965 4965 1985
rect 4925 1935 4965 1965
rect 4925 1915 4935 1935
rect 4955 1915 4965 1935
rect 4925 1900 4965 1915
rect 4985 1985 5025 2000
rect 4985 1965 4995 1985
rect 5015 1965 5025 1985
rect 4985 1935 5025 1965
rect 4985 1915 4995 1935
rect 5015 1915 5025 1935
rect 4985 1900 5025 1915
rect 5045 1985 5085 2000
rect 5045 1965 5055 1985
rect 5075 1965 5085 1985
rect 5045 1935 5085 1965
rect 5045 1915 5055 1935
rect 5075 1915 5085 1935
rect 5045 1900 5085 1915
rect 5105 1985 5145 2000
rect 5105 1965 5115 1985
rect 5135 1965 5145 1985
rect 5105 1935 5145 1965
rect 5105 1915 5115 1935
rect 5135 1915 5145 1935
rect 5105 1900 5145 1915
rect 5165 1985 5205 2000
rect 5165 1965 5175 1985
rect 5195 1965 5205 1985
rect 5165 1935 5205 1965
rect 5165 1915 5175 1935
rect 5195 1915 5205 1935
rect 5165 1900 5205 1915
rect 5225 1985 5265 2000
rect 5225 1965 5235 1985
rect 5255 1965 5265 1985
rect 5225 1935 5265 1965
rect 5225 1915 5235 1935
rect 5255 1915 5265 1935
rect 5225 1900 5265 1915
<< ndiffc >>
rect 10830 3495 10850 3515
rect 10830 3445 10850 3465
rect 10830 3395 10850 3415
rect 10830 3345 10850 3365
rect 10830 3295 10850 3315
rect 10500 3245 10520 3265
rect 10560 3250 10580 3270
rect 10620 3250 10640 3270
rect 10680 3245 10700 3265
rect 10830 3245 10850 3265
rect 10890 3495 10910 3515
rect 10890 3445 10910 3465
rect 10890 3395 10910 3415
rect 10890 3345 10910 3365
rect 10890 3295 10910 3315
rect 10890 3245 10910 3265
rect 10950 3495 10970 3515
rect 10950 3445 10970 3465
rect 10950 3395 10970 3415
rect 10950 3345 10970 3365
rect 10950 3295 10970 3315
rect 10950 3245 10970 3265
rect 11010 3545 11030 3565
rect 11010 3495 11030 3515
rect 11010 3445 11030 3465
rect 11010 3395 11030 3415
rect 11010 3345 11030 3365
rect 11010 3295 11030 3315
rect 11010 3245 11030 3265
rect 11070 3545 11090 3565
rect 11070 3495 11090 3515
rect 11070 3445 11090 3465
rect 11070 3395 11090 3415
rect 11070 3345 11090 3365
rect 11070 3295 11090 3315
rect 11070 3245 11090 3265
rect 11230 3540 11250 3560
rect 11230 3490 11250 3510
rect 11230 3440 11250 3460
rect 11230 3390 11250 3410
rect 11230 3340 11250 3360
rect 11230 3290 11250 3310
rect 11230 3240 11250 3260
rect 11230 3190 11250 3210
rect 11290 3540 11310 3560
rect 11290 3490 11310 3510
rect 11290 3440 11310 3460
rect 11290 3390 11310 3410
rect 11290 3340 11310 3360
rect 11290 3290 11310 3310
rect 11290 3240 11310 3260
rect 11290 3190 11310 3210
rect 11350 3540 11370 3560
rect 11350 3490 11370 3510
rect 11350 3440 11370 3460
rect 11350 3390 11370 3410
rect 11350 3340 11370 3360
rect 11350 3290 11370 3310
rect 11350 3240 11370 3260
rect 11350 3190 11370 3210
rect 11410 3540 11430 3560
rect 11410 3490 11430 3510
rect 11410 3440 11430 3460
rect 11410 3390 11430 3410
rect 11410 3340 11430 3360
rect 11410 3290 11430 3310
rect 11410 3240 11430 3260
rect 11410 3190 11430 3210
rect 11470 3540 11490 3560
rect 11470 3490 11490 3510
rect 11470 3440 11490 3460
rect 11470 3390 11490 3410
rect 11470 3340 11490 3360
rect 11470 3290 11490 3310
rect 11470 3240 11490 3260
rect 11470 3190 11490 3210
rect 11530 3540 11550 3560
rect 11530 3490 11550 3510
rect 11530 3440 11550 3460
rect 11530 3390 11550 3410
rect 11530 3340 11550 3360
rect 11530 3290 11550 3310
rect 11530 3240 11550 3260
rect 11530 3190 11550 3210
rect 11590 3540 11610 3560
rect 11590 3490 11610 3510
rect 11590 3440 11610 3460
rect 11590 3390 11610 3410
rect 11590 3340 11610 3360
rect 11590 3290 11610 3310
rect 11590 3240 11610 3260
rect 11590 3190 11610 3210
rect 11650 3540 11670 3560
rect 11650 3490 11670 3510
rect 11650 3440 11670 3460
rect 11650 3390 11670 3410
rect 11650 3340 11670 3360
rect 11650 3290 11670 3310
rect 11650 3240 11670 3260
rect 11650 3190 11670 3210
rect 11710 3540 11730 3560
rect 11710 3490 11730 3510
rect 11710 3440 11730 3460
rect 11710 3390 11730 3410
rect 11710 3340 11730 3360
rect 11710 3290 11730 3310
rect 11710 3240 11730 3260
rect 11710 3190 11730 3210
rect 11770 3540 11790 3560
rect 11770 3490 11790 3510
rect 11770 3440 11790 3460
rect 11770 3390 11790 3410
rect 11770 3340 11790 3360
rect 11770 3290 11790 3310
rect 11770 3240 11790 3260
rect 11770 3190 11790 3210
rect 11830 3540 11850 3560
rect 11830 3490 11850 3510
rect 11830 3440 11850 3460
rect 11830 3390 11850 3410
rect 11830 3340 11850 3360
rect 11830 3290 11850 3310
rect 11830 3240 11850 3260
rect 11830 3190 11850 3210
rect 11890 3540 11910 3560
rect 11890 3490 11910 3510
rect 11890 3440 11910 3460
rect 11890 3390 11910 3410
rect 11890 3340 11910 3360
rect 11890 3290 11910 3310
rect 11890 3240 11910 3260
rect 11890 3190 11910 3210
rect 11950 3540 11970 3560
rect 11950 3490 11970 3510
rect 11950 3440 11970 3460
rect 11950 3390 11970 3410
rect 11950 3340 11970 3360
rect 11950 3290 11970 3310
rect 11950 3240 11970 3260
rect 11950 3190 11970 3210
rect 12010 3540 12030 3560
rect 12010 3490 12030 3510
rect 12010 3440 12030 3460
rect 12010 3390 12030 3410
rect 12010 3340 12030 3360
rect 12010 3290 12030 3310
rect 12010 3240 12030 3260
rect 12010 3190 12030 3210
rect 12070 3540 12090 3560
rect 12070 3490 12090 3510
rect 12070 3440 12090 3460
rect 12070 3390 12090 3410
rect 12070 3340 12090 3360
rect 12070 3290 12090 3310
rect 12070 3240 12090 3260
rect 12070 3190 12090 3210
rect 12130 3540 12150 3560
rect 12130 3490 12150 3510
rect 12130 3440 12150 3460
rect 12130 3390 12150 3410
rect 12130 3340 12150 3360
rect 12130 3290 12150 3310
rect 12130 3240 12150 3260
rect 12130 3190 12150 3210
rect 12190 3540 12210 3560
rect 12190 3490 12210 3510
rect 12190 3440 12210 3460
rect 12190 3390 12210 3410
rect 12190 3340 12210 3360
rect 12190 3290 12210 3310
rect 12190 3240 12210 3260
rect 12190 3190 12210 3210
rect 12250 3540 12270 3560
rect 12250 3490 12270 3510
rect 12250 3440 12270 3460
rect 12250 3390 12270 3410
rect 12250 3340 12270 3360
rect 12250 3290 12270 3310
rect 12250 3240 12270 3260
rect 12250 3190 12270 3210
rect 12310 3540 12330 3560
rect 12310 3490 12330 3510
rect 12310 3440 12330 3460
rect 12310 3390 12330 3410
rect 12310 3340 12330 3360
rect 12310 3290 12330 3310
rect 12310 3240 12330 3260
rect 12310 3190 12330 3210
rect 12370 3540 12390 3560
rect 12370 3490 12390 3510
rect 12370 3440 12390 3460
rect 12370 3390 12390 3410
rect 12370 3340 12390 3360
rect 12370 3290 12390 3310
rect 12370 3240 12390 3260
rect 12370 3190 12390 3210
rect 12430 3540 12450 3560
rect 12430 3490 12450 3510
rect 12430 3440 12450 3460
rect 12430 3390 12450 3410
rect 12430 3340 12450 3360
rect 12430 3290 12450 3310
rect 12430 3240 12450 3260
rect 12430 3190 12450 3210
rect 12490 3540 12510 3560
rect 12490 3490 12510 3510
rect 12490 3440 12510 3460
rect 12490 3390 12510 3410
rect 12490 3340 12510 3360
rect 12490 3290 12510 3310
rect 12490 3240 12510 3260
rect 12490 3190 12510 3210
rect 12550 3540 12570 3560
rect 12550 3490 12570 3510
rect 12550 3440 12570 3460
rect 12550 3390 12570 3410
rect 12550 3340 12570 3360
rect 18330 3495 18350 3515
rect 18330 3445 18350 3465
rect 18330 3395 18350 3415
rect 12550 3290 12570 3310
rect 18330 3345 18350 3365
rect 18330 3295 18350 3315
rect 12550 3240 12570 3260
rect 18000 3245 18020 3265
rect 12550 3190 12570 3210
rect 12900 3205 12920 3225
rect 12900 3155 12920 3175
rect 12900 3105 12920 3125
rect 12900 3055 12920 3075
rect 12900 3005 12920 3025
rect 12900 2955 12920 2975
rect 12955 3205 12975 3225
rect 12955 3155 12975 3175
rect 12955 3105 12975 3125
rect 12955 3055 12975 3075
rect 12955 3005 12975 3025
rect 12955 2955 12975 2975
rect 13010 3205 13030 3225
rect 13010 3155 13030 3175
rect 13010 3105 13030 3125
rect 13010 3055 13030 3075
rect 13010 3005 13030 3025
rect 13010 2955 13030 2975
rect 13065 3205 13085 3225
rect 13065 3155 13085 3175
rect 13065 3105 13085 3125
rect 13065 3055 13085 3075
rect 13065 3005 13085 3025
rect 13065 2955 13085 2975
rect 13120 3205 13140 3225
rect 13120 3155 13140 3175
rect 13120 3105 13140 3125
rect 13120 3055 13140 3075
rect 13120 3005 13140 3025
rect 13120 2955 13140 2975
rect 13175 3205 13195 3225
rect 13175 3155 13195 3175
rect 13175 3105 13195 3125
rect 13175 3055 13195 3075
rect 13175 3005 13195 3025
rect 13175 2955 13195 2975
rect 13230 3205 13250 3225
rect 13230 3155 13250 3175
rect 13230 3105 13250 3125
rect 13230 3055 13250 3075
rect 13230 3005 13250 3025
rect 13230 2955 13250 2975
rect 13285 3205 13305 3225
rect 13285 3155 13305 3175
rect 13285 3105 13305 3125
rect 13285 3055 13305 3075
rect 13285 3005 13305 3025
rect 13285 2955 13305 2975
rect 13340 3205 13360 3225
rect 13340 3155 13360 3175
rect 13340 3105 13360 3125
rect 13340 3055 13360 3075
rect 13340 3005 13360 3025
rect 13340 2955 13360 2975
rect 13395 3205 13415 3225
rect 13395 3155 13415 3175
rect 13395 3105 13415 3125
rect 13395 3055 13415 3075
rect 13395 3005 13415 3025
rect 13395 2955 13415 2975
rect 13450 3205 13470 3225
rect 13450 3155 13470 3175
rect 13450 3105 13470 3125
rect 13450 3055 13470 3075
rect 13450 3005 13470 3025
rect 13450 2955 13470 2975
rect 13505 3205 13525 3225
rect 13505 3155 13525 3175
rect 13505 3105 13525 3125
rect 13505 3055 13525 3075
rect 13505 3005 13525 3025
rect 13505 2955 13525 2975
rect 13560 3205 13580 3225
rect 13560 3155 13580 3175
rect 13560 3105 13580 3125
rect 13560 3055 13580 3075
rect 13560 3005 13580 3025
rect 13560 2955 13580 2975
rect 13615 3205 13635 3225
rect 13615 3155 13635 3175
rect 13615 3105 13635 3125
rect 13615 3055 13635 3075
rect 13615 3005 13635 3025
rect 13615 2955 13635 2975
rect 13670 3205 13690 3225
rect 13670 3155 13690 3175
rect 13670 3105 13690 3125
rect 13670 3055 13690 3075
rect 13670 3005 13690 3025
rect 13670 2955 13690 2975
rect 13725 3205 13745 3225
rect 13725 3155 13745 3175
rect 13725 3105 13745 3125
rect 13725 3055 13745 3075
rect 13725 3005 13745 3025
rect 13725 2955 13745 2975
rect 13780 3205 13800 3225
rect 13780 3155 13800 3175
rect 13780 3105 13800 3125
rect 13780 3055 13800 3075
rect 13780 3005 13800 3025
rect 13780 2955 13800 2975
rect 13835 3205 13855 3225
rect 13835 3155 13855 3175
rect 13835 3105 13855 3125
rect 13835 3055 13855 3075
rect 13835 3005 13855 3025
rect 13835 2955 13855 2975
rect 13890 3205 13910 3225
rect 13890 3155 13910 3175
rect 13890 3105 13910 3125
rect 13890 3055 13910 3075
rect 13890 3005 13910 3025
rect 13890 2955 13910 2975
rect 13945 3205 13965 3225
rect 13945 3155 13965 3175
rect 13945 3105 13965 3125
rect 13945 3055 13965 3075
rect 13945 3005 13965 3025
rect 13945 2955 13965 2975
rect 14000 3205 14020 3225
rect 14000 3155 14020 3175
rect 14000 3105 14020 3125
rect 14000 3055 14020 3075
rect 14000 3005 14020 3025
rect 14000 2955 14020 2975
rect 14055 3205 14075 3225
rect 14055 3155 14075 3175
rect 14055 3105 14075 3125
rect 14055 3055 14075 3075
rect 14055 3005 14075 3025
rect 14055 2955 14075 2975
rect 18060 3250 18080 3270
rect 18120 3250 18140 3270
rect 18180 3245 18200 3265
rect 18330 3245 18350 3265
rect 18390 3495 18410 3515
rect 18390 3445 18410 3465
rect 18390 3395 18410 3415
rect 18390 3345 18410 3365
rect 18390 3295 18410 3315
rect 18390 3245 18410 3265
rect 18450 3495 18470 3515
rect 18450 3445 18470 3465
rect 18450 3395 18470 3415
rect 18450 3345 18470 3365
rect 18450 3295 18470 3315
rect 18450 3245 18470 3265
rect 18510 3545 18530 3565
rect 18510 3495 18530 3515
rect 18510 3445 18530 3465
rect 18510 3395 18530 3415
rect 18510 3345 18530 3365
rect 18510 3295 18530 3315
rect 18510 3245 18530 3265
rect 18570 3545 18590 3565
rect 18570 3495 18590 3515
rect 18570 3445 18590 3465
rect 18570 3395 18590 3415
rect 18570 3345 18590 3365
rect 18570 3295 18590 3315
rect 18570 3245 18590 3265
rect 18730 3540 18750 3560
rect 18730 3490 18750 3510
rect 18730 3440 18750 3460
rect 18730 3390 18750 3410
rect 18730 3340 18750 3360
rect 18730 3290 18750 3310
rect 18730 3240 18750 3260
rect 14110 3205 14130 3225
rect 18730 3190 18750 3210
rect 18790 3540 18810 3560
rect 18790 3490 18810 3510
rect 18790 3440 18810 3460
rect 18790 3390 18810 3410
rect 18790 3340 18810 3360
rect 18790 3290 18810 3310
rect 18790 3240 18810 3260
rect 18790 3190 18810 3210
rect 18850 3540 18870 3560
rect 18850 3490 18870 3510
rect 18850 3440 18870 3460
rect 18850 3390 18870 3410
rect 18850 3340 18870 3360
rect 18850 3290 18870 3310
rect 18850 3240 18870 3260
rect 18850 3190 18870 3210
rect 18910 3540 18930 3560
rect 18910 3490 18930 3510
rect 18910 3440 18930 3460
rect 18910 3390 18930 3410
rect 18910 3340 18930 3360
rect 18910 3290 18930 3310
rect 18910 3240 18930 3260
rect 18910 3190 18930 3210
rect 18970 3540 18990 3560
rect 18970 3490 18990 3510
rect 18970 3440 18990 3460
rect 18970 3390 18990 3410
rect 18970 3340 18990 3360
rect 18970 3290 18990 3310
rect 18970 3240 18990 3260
rect 18970 3190 18990 3210
rect 19030 3540 19050 3560
rect 19030 3490 19050 3510
rect 19030 3440 19050 3460
rect 19030 3390 19050 3410
rect 19030 3340 19050 3360
rect 19030 3290 19050 3310
rect 19030 3240 19050 3260
rect 19030 3190 19050 3210
rect 19090 3540 19110 3560
rect 19090 3490 19110 3510
rect 19090 3440 19110 3460
rect 19090 3390 19110 3410
rect 19090 3340 19110 3360
rect 19090 3290 19110 3310
rect 19090 3240 19110 3260
rect 19090 3190 19110 3210
rect 19150 3540 19170 3560
rect 19150 3490 19170 3510
rect 19150 3440 19170 3460
rect 19150 3390 19170 3410
rect 19150 3340 19170 3360
rect 19150 3290 19170 3310
rect 19150 3240 19170 3260
rect 19150 3190 19170 3210
rect 19210 3540 19230 3560
rect 19210 3490 19230 3510
rect 19210 3440 19230 3460
rect 19210 3390 19230 3410
rect 19210 3340 19230 3360
rect 19210 3290 19230 3310
rect 19210 3240 19230 3260
rect 19210 3190 19230 3210
rect 19270 3540 19290 3560
rect 19270 3490 19290 3510
rect 19270 3440 19290 3460
rect 19270 3390 19290 3410
rect 19270 3340 19290 3360
rect 19270 3290 19290 3310
rect 19270 3240 19290 3260
rect 19270 3190 19290 3210
rect 19330 3540 19350 3560
rect 19330 3490 19350 3510
rect 19330 3440 19350 3460
rect 19330 3390 19350 3410
rect 19330 3340 19350 3360
rect 19330 3290 19350 3310
rect 19330 3240 19350 3260
rect 19330 3190 19350 3210
rect 19390 3540 19410 3560
rect 19390 3490 19410 3510
rect 19390 3440 19410 3460
rect 19390 3390 19410 3410
rect 19390 3340 19410 3360
rect 19390 3290 19410 3310
rect 19390 3240 19410 3260
rect 19390 3190 19410 3210
rect 19450 3540 19470 3560
rect 19450 3490 19470 3510
rect 19450 3440 19470 3460
rect 19450 3390 19470 3410
rect 19450 3340 19470 3360
rect 19450 3290 19470 3310
rect 19450 3240 19470 3260
rect 19450 3190 19470 3210
rect 19510 3540 19530 3560
rect 19510 3490 19530 3510
rect 19510 3440 19530 3460
rect 19510 3390 19530 3410
rect 19510 3340 19530 3360
rect 19510 3290 19530 3310
rect 19510 3240 19530 3260
rect 19510 3190 19530 3210
rect 19570 3540 19590 3560
rect 19570 3490 19590 3510
rect 19570 3440 19590 3460
rect 19570 3390 19590 3410
rect 19570 3340 19590 3360
rect 19570 3290 19590 3310
rect 19570 3240 19590 3260
rect 19570 3190 19590 3210
rect 19630 3540 19650 3560
rect 19630 3490 19650 3510
rect 19630 3440 19650 3460
rect 19630 3390 19650 3410
rect 19630 3340 19650 3360
rect 19630 3290 19650 3310
rect 19630 3240 19650 3260
rect 19630 3190 19650 3210
rect 19690 3540 19710 3560
rect 19690 3490 19710 3510
rect 19690 3440 19710 3460
rect 19690 3390 19710 3410
rect 19690 3340 19710 3360
rect 19690 3290 19710 3310
rect 19690 3240 19710 3260
rect 19690 3190 19710 3210
rect 19750 3540 19770 3560
rect 19750 3490 19770 3510
rect 19750 3440 19770 3460
rect 19750 3390 19770 3410
rect 19750 3340 19770 3360
rect 19750 3290 19770 3310
rect 19750 3240 19770 3260
rect 19750 3190 19770 3210
rect 19810 3540 19830 3560
rect 19810 3490 19830 3510
rect 19810 3440 19830 3460
rect 19810 3390 19830 3410
rect 19810 3340 19830 3360
rect 19810 3290 19830 3310
rect 19810 3240 19830 3260
rect 19810 3190 19830 3210
rect 19870 3540 19890 3560
rect 19870 3490 19890 3510
rect 19870 3440 19890 3460
rect 19870 3390 19890 3410
rect 19870 3340 19890 3360
rect 19870 3290 19890 3310
rect 19870 3240 19890 3260
rect 19870 3190 19890 3210
rect 19930 3540 19950 3560
rect 19930 3490 19950 3510
rect 19930 3440 19950 3460
rect 19930 3390 19950 3410
rect 19930 3340 19950 3360
rect 19930 3290 19950 3310
rect 19930 3240 19950 3260
rect 19930 3190 19950 3210
rect 19990 3540 20010 3560
rect 19990 3490 20010 3510
rect 19990 3440 20010 3460
rect 19990 3390 20010 3410
rect 19990 3340 20010 3360
rect 19990 3290 20010 3310
rect 19990 3240 20010 3260
rect 19990 3190 20010 3210
rect 20050 3540 20070 3560
rect 20050 3490 20070 3510
rect 20050 3440 20070 3460
rect 20050 3390 20070 3410
rect 20050 3340 20070 3360
rect 20050 3290 20070 3310
rect 20050 3240 20070 3260
rect 20050 3190 20070 3210
rect 20400 3205 20420 3225
rect 14110 3155 14130 3175
rect 20400 3155 20420 3175
rect 14110 3105 14130 3125
rect 14110 3055 14130 3075
rect 14110 3005 14130 3025
rect 14110 2955 14130 2975
rect 20400 3105 20420 3125
rect 20400 3055 20420 3075
rect 20400 3005 20420 3025
rect 20400 2955 20420 2975
rect 11230 2860 11250 2880
rect 11230 2810 11250 2830
rect 11230 2760 11250 2780
rect 11230 2710 11250 2730
rect 11230 2660 11250 2680
rect 9690 2585 9710 2605
rect 9690 2535 9710 2555
rect 9745 2585 9765 2605
rect 9745 2535 9765 2555
rect 9800 2585 9820 2605
rect 9800 2535 9820 2555
rect 9855 2585 9875 2605
rect 9855 2535 9875 2555
rect 9910 2585 9930 2605
rect 9910 2535 9930 2555
rect 9965 2585 9985 2605
rect 9965 2535 9985 2555
rect 10020 2585 10040 2605
rect 10020 2535 10040 2555
rect 10075 2585 10095 2605
rect 10075 2535 10095 2555
rect 10130 2585 10150 2605
rect 10130 2535 10150 2555
rect 10185 2585 10205 2605
rect 10185 2535 10205 2555
rect 10240 2585 10260 2605
rect 10240 2535 10260 2555
rect 10295 2585 10315 2605
rect 10295 2535 10315 2555
rect 10350 2585 10370 2605
rect 10350 2535 10370 2555
rect 10405 2585 10425 2605
rect 10405 2535 10425 2555
rect 10460 2585 10480 2605
rect 10460 2535 10480 2555
rect 10515 2585 10535 2605
rect 10515 2535 10535 2555
rect 10570 2585 10590 2605
rect 10570 2535 10590 2555
rect 10625 2585 10645 2605
rect 10625 2535 10645 2555
rect 10680 2585 10700 2605
rect 10680 2535 10700 2555
rect 10735 2585 10755 2605
rect 10735 2535 10755 2555
rect 10790 2585 10810 2605
rect 10790 2535 10810 2555
rect 10845 2585 10865 2605
rect 10845 2535 10865 2555
rect 10900 2585 10920 2605
rect 10900 2535 10920 2555
rect 11230 2610 11250 2630
rect 11230 2560 11250 2580
rect 11230 2510 11250 2530
rect 11290 2860 11310 2880
rect 11290 2810 11310 2830
rect 11290 2760 11310 2780
rect 11290 2710 11310 2730
rect 11290 2660 11310 2680
rect 11290 2610 11310 2630
rect 11290 2560 11310 2580
rect 11290 2510 11310 2530
rect 11350 2860 11370 2880
rect 11350 2810 11370 2830
rect 11350 2760 11370 2780
rect 11350 2710 11370 2730
rect 11350 2660 11370 2680
rect 11350 2610 11370 2630
rect 11350 2560 11370 2580
rect 11350 2510 11370 2530
rect 11410 2860 11430 2880
rect 11410 2810 11430 2830
rect 11410 2760 11430 2780
rect 11410 2710 11430 2730
rect 11410 2660 11430 2680
rect 11410 2610 11430 2630
rect 11410 2560 11430 2580
rect 11410 2510 11430 2530
rect 11470 2860 11490 2880
rect 11470 2810 11490 2830
rect 11470 2760 11490 2780
rect 11470 2710 11490 2730
rect 11470 2660 11490 2680
rect 11470 2610 11490 2630
rect 11470 2560 11490 2580
rect 11470 2510 11490 2530
rect 11530 2860 11550 2880
rect 11530 2810 11550 2830
rect 11530 2760 11550 2780
rect 11530 2710 11550 2730
rect 11530 2660 11550 2680
rect 11530 2610 11550 2630
rect 11530 2560 11550 2580
rect 11530 2510 11550 2530
rect 11590 2860 11610 2880
rect 11590 2810 11610 2830
rect 11590 2760 11610 2780
rect 11590 2710 11610 2730
rect 11590 2660 11610 2680
rect 11590 2610 11610 2630
rect 11590 2560 11610 2580
rect 11590 2510 11610 2530
rect 11650 2860 11670 2880
rect 11650 2810 11670 2830
rect 11650 2760 11670 2780
rect 11650 2710 11670 2730
rect 11650 2660 11670 2680
rect 11650 2610 11670 2630
rect 11650 2560 11670 2580
rect 11650 2510 11670 2530
rect 11710 2860 11730 2880
rect 11710 2810 11730 2830
rect 11710 2760 11730 2780
rect 11710 2710 11730 2730
rect 11710 2660 11730 2680
rect 11710 2610 11730 2630
rect 11710 2560 11730 2580
rect 11710 2510 11730 2530
rect 11770 2860 11790 2880
rect 11770 2810 11790 2830
rect 11770 2760 11790 2780
rect 11770 2710 11790 2730
rect 11770 2660 11790 2680
rect 11770 2610 11790 2630
rect 11770 2560 11790 2580
rect 11770 2510 11790 2530
rect 11830 2860 11850 2880
rect 11830 2810 11850 2830
rect 11830 2760 11850 2780
rect 11830 2710 11850 2730
rect 11830 2660 11850 2680
rect 11830 2610 11850 2630
rect 11830 2560 11850 2580
rect 11830 2510 11850 2530
rect 11890 2860 11910 2880
rect 11890 2810 11910 2830
rect 11890 2760 11910 2780
rect 11890 2710 11910 2730
rect 11890 2660 11910 2680
rect 11890 2610 11910 2630
rect 11890 2560 11910 2580
rect 11890 2510 11910 2530
rect 11950 2860 11970 2880
rect 11950 2810 11970 2830
rect 11950 2760 11970 2780
rect 11950 2710 11970 2730
rect 11950 2660 11970 2680
rect 11950 2610 11970 2630
rect 11950 2560 11970 2580
rect 11950 2510 11970 2530
rect 12010 2860 12030 2880
rect 12010 2810 12030 2830
rect 12010 2760 12030 2780
rect 12010 2710 12030 2730
rect 12010 2660 12030 2680
rect 12010 2610 12030 2630
rect 12010 2560 12030 2580
rect 12010 2510 12030 2530
rect 12070 2860 12090 2880
rect 12070 2810 12090 2830
rect 12070 2760 12090 2780
rect 12070 2710 12090 2730
rect 12070 2660 12090 2680
rect 12070 2610 12090 2630
rect 12070 2560 12090 2580
rect 12070 2510 12090 2530
rect 12130 2860 12150 2880
rect 12130 2810 12150 2830
rect 12130 2760 12150 2780
rect 12130 2710 12150 2730
rect 12130 2660 12150 2680
rect 12130 2610 12150 2630
rect 12130 2560 12150 2580
rect 12130 2510 12150 2530
rect 12190 2860 12210 2880
rect 12190 2810 12210 2830
rect 12190 2760 12210 2780
rect 12190 2710 12210 2730
rect 12190 2660 12210 2680
rect 12190 2610 12210 2630
rect 12190 2560 12210 2580
rect 12190 2510 12210 2530
rect 12250 2860 12270 2880
rect 12250 2810 12270 2830
rect 12250 2760 12270 2780
rect 12250 2710 12270 2730
rect 12250 2660 12270 2680
rect 12250 2610 12270 2630
rect 12250 2560 12270 2580
rect 12250 2510 12270 2530
rect 12310 2860 12330 2880
rect 12310 2810 12330 2830
rect 12310 2760 12330 2780
rect 12310 2710 12330 2730
rect 12310 2660 12330 2680
rect 12310 2610 12330 2630
rect 12310 2560 12330 2580
rect 12310 2510 12330 2530
rect 12370 2860 12390 2880
rect 12370 2810 12390 2830
rect 12370 2760 12390 2780
rect 12370 2710 12390 2730
rect 12370 2660 12390 2680
rect 12370 2610 12390 2630
rect 12370 2560 12390 2580
rect 12370 2510 12390 2530
rect 12430 2860 12450 2880
rect 12430 2810 12450 2830
rect 12430 2760 12450 2780
rect 12430 2710 12450 2730
rect 12430 2660 12450 2680
rect 12430 2610 12450 2630
rect 12430 2560 12450 2580
rect 12430 2510 12450 2530
rect 12490 2860 12510 2880
rect 12490 2810 12510 2830
rect 12490 2760 12510 2780
rect 12490 2710 12510 2730
rect 12490 2660 12510 2680
rect 12490 2610 12510 2630
rect 12490 2560 12510 2580
rect 12490 2510 12510 2530
rect 20455 3205 20475 3225
rect 20455 3155 20475 3175
rect 20455 3105 20475 3125
rect 20455 3055 20475 3075
rect 20455 3005 20475 3025
rect 20455 2955 20475 2975
rect 20510 3205 20530 3225
rect 20510 3155 20530 3175
rect 20510 3105 20530 3125
rect 20510 3055 20530 3075
rect 20510 3005 20530 3025
rect 20510 2955 20530 2975
rect 20565 3205 20585 3225
rect 20565 3155 20585 3175
rect 20565 3105 20585 3125
rect 20565 3055 20585 3075
rect 20565 3005 20585 3025
rect 20565 2955 20585 2975
rect 20620 3205 20640 3225
rect 20620 3155 20640 3175
rect 20620 3105 20640 3125
rect 20620 3055 20640 3075
rect 20620 3005 20640 3025
rect 20620 2955 20640 2975
rect 20675 3205 20695 3225
rect 20675 3155 20695 3175
rect 20675 3105 20695 3125
rect 20675 3055 20695 3075
rect 20675 3005 20695 3025
rect 20675 2955 20695 2975
rect 20730 3205 20750 3225
rect 20730 3155 20750 3175
rect 20730 3105 20750 3125
rect 20730 3055 20750 3075
rect 20730 3005 20750 3025
rect 20730 2955 20750 2975
rect 20785 3205 20805 3225
rect 20785 3155 20805 3175
rect 20785 3105 20805 3125
rect 20785 3055 20805 3075
rect 20785 3005 20805 3025
rect 20785 2955 20805 2975
rect 20840 3205 20860 3225
rect 20840 3155 20860 3175
rect 20840 3105 20860 3125
rect 20840 3055 20860 3075
rect 20840 3005 20860 3025
rect 20840 2955 20860 2975
rect 20895 3205 20915 3225
rect 20895 3155 20915 3175
rect 20895 3105 20915 3125
rect 20895 3055 20915 3075
rect 20895 3005 20915 3025
rect 20895 2955 20915 2975
rect 20950 3205 20970 3225
rect 20950 3155 20970 3175
rect 20950 3105 20970 3125
rect 20950 3055 20970 3075
rect 20950 3005 20970 3025
rect 20950 2955 20970 2975
rect 21005 3205 21025 3225
rect 21005 3155 21025 3175
rect 21005 3105 21025 3125
rect 21005 3055 21025 3075
rect 21005 3005 21025 3025
rect 21005 2955 21025 2975
rect 21060 3205 21080 3225
rect 21060 3155 21080 3175
rect 21060 3105 21080 3125
rect 21060 3055 21080 3075
rect 21060 3005 21080 3025
rect 21060 2955 21080 2975
rect 21115 3205 21135 3225
rect 21115 3155 21135 3175
rect 21115 3105 21135 3125
rect 21115 3055 21135 3075
rect 21115 3005 21135 3025
rect 21115 2955 21135 2975
rect 21170 3205 21190 3225
rect 21170 3155 21190 3175
rect 21170 3105 21190 3125
rect 21170 3055 21190 3075
rect 21170 3005 21190 3025
rect 21170 2955 21190 2975
rect 21225 3205 21245 3225
rect 21225 3155 21245 3175
rect 21225 3105 21245 3125
rect 21225 3055 21245 3075
rect 21225 3005 21245 3025
rect 21225 2955 21245 2975
rect 21280 3205 21300 3225
rect 21280 3155 21300 3175
rect 21280 3105 21300 3125
rect 21280 3055 21300 3075
rect 21280 3005 21300 3025
rect 21280 2955 21300 2975
rect 21335 3205 21355 3225
rect 21335 3155 21355 3175
rect 21335 3105 21355 3125
rect 21335 3055 21355 3075
rect 21335 3005 21355 3025
rect 21335 2955 21355 2975
rect 21390 3205 21410 3225
rect 21390 3155 21410 3175
rect 21390 3105 21410 3125
rect 21390 3055 21410 3075
rect 21390 3005 21410 3025
rect 21390 2955 21410 2975
rect 21445 3205 21465 3225
rect 21445 3155 21465 3175
rect 21445 3105 21465 3125
rect 21445 3055 21465 3075
rect 21445 3005 21465 3025
rect 21445 2955 21465 2975
rect 21500 3205 21520 3225
rect 21500 3155 21520 3175
rect 21500 3105 21520 3125
rect 21500 3055 21520 3075
rect 21500 3005 21520 3025
rect 21500 2955 21520 2975
rect 21555 3205 21575 3225
rect 21555 3155 21575 3175
rect 21555 3105 21575 3125
rect 21555 3055 21575 3075
rect 21555 3005 21575 3025
rect 21555 2955 21575 2975
rect 21610 3205 21630 3225
rect 21610 3155 21630 3175
rect 21610 3105 21630 3125
rect 21610 3055 21630 3075
rect 21610 3005 21630 3025
rect 21610 2955 21630 2975
rect 12550 2860 12570 2880
rect 18730 2860 18750 2880
rect 12550 2810 12570 2830
rect 12550 2760 12570 2780
rect 12550 2710 12570 2730
rect 18730 2810 18750 2830
rect 18730 2760 18750 2780
rect 18730 2710 18750 2730
rect 12550 2660 12570 2680
rect 18730 2660 18750 2680
rect 12550 2610 12570 2630
rect 12550 2560 12570 2580
rect 12550 2510 12570 2530
rect 12900 2585 12920 2605
rect 12900 2535 12920 2555
rect 12955 2585 12975 2605
rect 12955 2535 12975 2555
rect 13010 2585 13030 2605
rect 13010 2535 13030 2555
rect 13065 2585 13085 2605
rect 13065 2535 13085 2555
rect 13120 2585 13140 2605
rect 13120 2535 13140 2555
rect 13175 2585 13195 2605
rect 13175 2535 13195 2555
rect 13230 2585 13250 2605
rect 13230 2535 13250 2555
rect 13285 2585 13305 2605
rect 13285 2535 13305 2555
rect 13340 2585 13360 2605
rect 13340 2535 13360 2555
rect 13395 2585 13415 2605
rect 13395 2535 13415 2555
rect 13450 2585 13470 2605
rect 13450 2535 13470 2555
rect 13505 2585 13525 2605
rect 13505 2535 13525 2555
rect 13560 2585 13580 2605
rect 13560 2535 13580 2555
rect 13615 2585 13635 2605
rect 13615 2535 13635 2555
rect 13670 2585 13690 2605
rect 13670 2535 13690 2555
rect 13725 2585 13745 2605
rect 13725 2535 13745 2555
rect 13780 2585 13800 2605
rect 13780 2535 13800 2555
rect 13835 2585 13855 2605
rect 13835 2535 13855 2555
rect 13890 2585 13910 2605
rect 13890 2535 13910 2555
rect 13945 2585 13965 2605
rect 13945 2535 13965 2555
rect 14000 2585 14020 2605
rect 14000 2535 14020 2555
rect 14055 2585 14075 2605
rect 14055 2535 14075 2555
rect 14110 2585 14130 2605
rect 14110 2535 14130 2555
rect 17190 2585 17210 2605
rect 17190 2535 17210 2555
rect 17245 2585 17265 2605
rect 17245 2535 17265 2555
rect 17300 2585 17320 2605
rect 17300 2535 17320 2555
rect 17355 2585 17375 2605
rect 17355 2535 17375 2555
rect 17410 2585 17430 2605
rect 17410 2535 17430 2555
rect 17465 2585 17485 2605
rect 17465 2535 17485 2555
rect 17520 2585 17540 2605
rect 17520 2535 17540 2555
rect 17575 2585 17595 2605
rect 17575 2535 17595 2555
rect 17630 2585 17650 2605
rect 17630 2535 17650 2555
rect 17685 2585 17705 2605
rect 17685 2535 17705 2555
rect 17740 2585 17760 2605
rect 17740 2535 17760 2555
rect 17795 2585 17815 2605
rect 17795 2535 17815 2555
rect 17850 2585 17870 2605
rect 17850 2535 17870 2555
rect 17905 2585 17925 2605
rect 17905 2535 17925 2555
rect 17960 2585 17980 2605
rect 17960 2535 17980 2555
rect 18015 2585 18035 2605
rect 18015 2535 18035 2555
rect 18070 2585 18090 2605
rect 18070 2535 18090 2555
rect 18125 2585 18145 2605
rect 18125 2535 18145 2555
rect 18180 2585 18200 2605
rect 18180 2535 18200 2555
rect 18235 2585 18255 2605
rect 18235 2535 18255 2555
rect 18290 2585 18310 2605
rect 18290 2535 18310 2555
rect 18345 2585 18365 2605
rect 18345 2535 18365 2555
rect 18400 2585 18420 2605
rect 18400 2535 18420 2555
rect 18730 2610 18750 2630
rect 18730 2560 18750 2580
rect 18730 2510 18750 2530
rect 18790 2860 18810 2880
rect 18790 2810 18810 2830
rect 18790 2760 18810 2780
rect 18790 2710 18810 2730
rect 18790 2660 18810 2680
rect 18790 2610 18810 2630
rect 18790 2560 18810 2580
rect 18790 2510 18810 2530
rect 18850 2860 18870 2880
rect 18850 2810 18870 2830
rect 18850 2760 18870 2780
rect 18850 2710 18870 2730
rect 18850 2660 18870 2680
rect 18850 2610 18870 2630
rect 18850 2560 18870 2580
rect 18850 2510 18870 2530
rect 18910 2860 18930 2880
rect 18910 2810 18930 2830
rect 18910 2760 18930 2780
rect 18910 2710 18930 2730
rect 18910 2660 18930 2680
rect 18910 2610 18930 2630
rect 18910 2560 18930 2580
rect 18910 2510 18930 2530
rect 18970 2860 18990 2880
rect 18970 2810 18990 2830
rect 18970 2760 18990 2780
rect 18970 2710 18990 2730
rect 18970 2660 18990 2680
rect 18970 2610 18990 2630
rect 18970 2560 18990 2580
rect 18970 2510 18990 2530
rect 19030 2860 19050 2880
rect 19030 2810 19050 2830
rect 19030 2760 19050 2780
rect 19030 2710 19050 2730
rect 19030 2660 19050 2680
rect 19030 2610 19050 2630
rect 19030 2560 19050 2580
rect 19030 2510 19050 2530
rect 19090 2860 19110 2880
rect 19090 2810 19110 2830
rect 19090 2760 19110 2780
rect 19090 2710 19110 2730
rect 19090 2660 19110 2680
rect 19090 2610 19110 2630
rect 19090 2560 19110 2580
rect 19090 2510 19110 2530
rect 19150 2860 19170 2880
rect 19150 2810 19170 2830
rect 19150 2760 19170 2780
rect 19150 2710 19170 2730
rect 19150 2660 19170 2680
rect 19150 2610 19170 2630
rect 19150 2560 19170 2580
rect 19150 2510 19170 2530
rect 19210 2860 19230 2880
rect 19210 2810 19230 2830
rect 19210 2760 19230 2780
rect 19210 2710 19230 2730
rect 19210 2660 19230 2680
rect 19210 2610 19230 2630
rect 19210 2560 19230 2580
rect 19210 2510 19230 2530
rect 19270 2860 19290 2880
rect 19270 2810 19290 2830
rect 19270 2760 19290 2780
rect 19270 2710 19290 2730
rect 19270 2660 19290 2680
rect 19270 2610 19290 2630
rect 19270 2560 19290 2580
rect 19270 2510 19290 2530
rect 19330 2860 19350 2880
rect 19330 2810 19350 2830
rect 19330 2760 19350 2780
rect 19330 2710 19350 2730
rect 19330 2660 19350 2680
rect 19330 2610 19350 2630
rect 19330 2560 19350 2580
rect 19330 2510 19350 2530
rect 19390 2860 19410 2880
rect 19390 2810 19410 2830
rect 19390 2760 19410 2780
rect 19390 2710 19410 2730
rect 19390 2660 19410 2680
rect 19390 2610 19410 2630
rect 19390 2560 19410 2580
rect 19390 2510 19410 2530
rect 19450 2860 19470 2880
rect 19450 2810 19470 2830
rect 19450 2760 19470 2780
rect 19450 2710 19470 2730
rect 19450 2660 19470 2680
rect 19450 2610 19470 2630
rect 19450 2560 19470 2580
rect 19450 2510 19470 2530
rect 19510 2860 19530 2880
rect 19510 2810 19530 2830
rect 19510 2760 19530 2780
rect 19510 2710 19530 2730
rect 19510 2660 19530 2680
rect 19510 2610 19530 2630
rect 19510 2560 19530 2580
rect 19510 2510 19530 2530
rect 19570 2860 19590 2880
rect 19570 2810 19590 2830
rect 19570 2760 19590 2780
rect 19570 2710 19590 2730
rect 19570 2660 19590 2680
rect 19570 2610 19590 2630
rect 19570 2560 19590 2580
rect 19570 2510 19590 2530
rect 19630 2860 19650 2880
rect 19630 2810 19650 2830
rect 19630 2760 19650 2780
rect 19630 2710 19650 2730
rect 19630 2660 19650 2680
rect 19630 2610 19650 2630
rect 19630 2560 19650 2580
rect 19630 2510 19650 2530
rect 19690 2860 19710 2880
rect 19690 2810 19710 2830
rect 19690 2760 19710 2780
rect 19690 2710 19710 2730
rect 19690 2660 19710 2680
rect 19690 2610 19710 2630
rect 19690 2560 19710 2580
rect 19690 2510 19710 2530
rect 19750 2860 19770 2880
rect 19750 2810 19770 2830
rect 19750 2760 19770 2780
rect 19750 2710 19770 2730
rect 19750 2660 19770 2680
rect 19750 2610 19770 2630
rect 19750 2560 19770 2580
rect 19750 2510 19770 2530
rect 19810 2860 19830 2880
rect 19810 2810 19830 2830
rect 19810 2760 19830 2780
rect 19810 2710 19830 2730
rect 19810 2660 19830 2680
rect 19810 2610 19830 2630
rect 19810 2560 19830 2580
rect 19810 2510 19830 2530
rect 19870 2860 19890 2880
rect 19870 2810 19890 2830
rect 19870 2760 19890 2780
rect 19870 2710 19890 2730
rect 19870 2660 19890 2680
rect 19870 2610 19890 2630
rect 19870 2560 19890 2580
rect 19870 2510 19890 2530
rect 19930 2860 19950 2880
rect 19930 2810 19950 2830
rect 19930 2760 19950 2780
rect 19930 2710 19950 2730
rect 19930 2660 19950 2680
rect 19930 2610 19950 2630
rect 19930 2560 19950 2580
rect 19930 2510 19950 2530
rect 19990 2860 20010 2880
rect 19990 2810 20010 2830
rect 19990 2760 20010 2780
rect 19990 2710 20010 2730
rect 19990 2660 20010 2680
rect 19990 2610 20010 2630
rect 19990 2560 20010 2580
rect 19990 2510 20010 2530
rect 20050 2860 20070 2880
rect 20050 2810 20070 2830
rect 20050 2760 20070 2780
rect 20050 2710 20070 2730
rect 20050 2660 20070 2680
rect 20050 2610 20070 2630
rect 20050 2560 20070 2580
rect 20050 2510 20070 2530
rect 20400 2585 20420 2605
rect 20400 2535 20420 2555
rect 20455 2585 20475 2605
rect 20455 2535 20475 2555
rect 20510 2585 20530 2605
rect 20510 2535 20530 2555
rect 20565 2585 20585 2605
rect 20565 2535 20585 2555
rect 20620 2585 20640 2605
rect 20620 2535 20640 2555
rect 20675 2585 20695 2605
rect 20675 2535 20695 2555
rect 20730 2585 20750 2605
rect 20730 2535 20750 2555
rect 20785 2585 20805 2605
rect 20785 2535 20805 2555
rect 20840 2585 20860 2605
rect 20840 2535 20860 2555
rect 20895 2585 20915 2605
rect 20895 2535 20915 2555
rect 20950 2585 20970 2605
rect 20950 2535 20970 2555
rect 21005 2585 21025 2605
rect 21005 2535 21025 2555
rect 21060 2585 21080 2605
rect 21060 2535 21080 2555
rect 21115 2585 21135 2605
rect 21115 2535 21135 2555
rect 21170 2585 21190 2605
rect 21170 2535 21190 2555
rect 21225 2585 21245 2605
rect 21225 2535 21245 2555
rect 21280 2585 21300 2605
rect 21280 2535 21300 2555
rect 21335 2585 21355 2605
rect 21335 2535 21355 2555
rect 21390 2585 21410 2605
rect 21390 2535 21410 2555
rect 21445 2585 21465 2605
rect 21445 2535 21465 2555
rect 21500 2585 21520 2605
rect 21500 2535 21520 2555
rect 21555 2585 21575 2605
rect 21555 2535 21575 2555
rect 21610 2585 21630 2605
rect 21610 2535 21630 2555
rect 9690 2135 9710 2155
rect 9690 2085 9710 2105
rect 9690 2035 9710 2055
rect 9745 2135 9765 2155
rect 9745 2085 9765 2105
rect 9745 2035 9765 2055
rect 9800 2135 9820 2155
rect 9800 2085 9820 2105
rect 9800 2035 9820 2055
rect 9855 2135 9875 2155
rect 9855 2085 9875 2105
rect 9855 2035 9875 2055
rect 9910 2135 9930 2155
rect 9910 2085 9930 2105
rect 9910 2035 9930 2055
rect 9965 2135 9985 2155
rect 9965 2085 9985 2105
rect 9965 2035 9985 2055
rect 10020 2135 10040 2155
rect 10020 2085 10040 2105
rect 10020 2035 10040 2055
rect 10075 2135 10095 2155
rect 10075 2085 10095 2105
rect 10075 2035 10095 2055
rect 10130 2135 10150 2155
rect 10130 2085 10150 2105
rect 10130 2035 10150 2055
rect 10185 2135 10205 2155
rect 10185 2085 10205 2105
rect 10185 2035 10205 2055
rect 10240 2135 10260 2155
rect 10240 2085 10260 2105
rect 10240 2035 10260 2055
rect 10295 2135 10315 2155
rect 10295 2085 10315 2105
rect 10295 2035 10315 2055
rect 10350 2135 10370 2155
rect 10350 2085 10370 2105
rect 10350 2035 10370 2055
rect 10405 2135 10425 2155
rect 10405 2085 10425 2105
rect 10405 2035 10425 2055
rect 10460 2135 10480 2155
rect 10460 2085 10480 2105
rect 10460 2035 10480 2055
rect 10515 2135 10535 2155
rect 10515 2085 10535 2105
rect 10515 2035 10535 2055
rect 10570 2135 10590 2155
rect 10570 2085 10590 2105
rect 10570 2035 10590 2055
rect 10625 2135 10645 2155
rect 10625 2085 10645 2105
rect 10625 2035 10645 2055
rect 10680 2135 10700 2155
rect 10680 2085 10700 2105
rect 10680 2035 10700 2055
rect 10735 2135 10755 2155
rect 10735 2085 10755 2105
rect 10735 2035 10755 2055
rect 10790 2135 10810 2155
rect 10790 2085 10810 2105
rect 10790 2035 10810 2055
rect 10845 2135 10865 2155
rect 10845 2085 10865 2105
rect 10845 2035 10865 2055
rect 10900 2135 10920 2155
rect 12900 2135 12920 2155
rect 10900 2085 10920 2105
rect 10900 2035 10920 2055
rect 11285 2095 11305 2115
rect 11285 2045 11305 2065
rect 11285 1995 11305 2015
rect 11340 2095 11360 2115
rect 11340 2045 11360 2065
rect 11340 1995 11360 2015
rect 11395 2095 11415 2115
rect 11395 2045 11415 2065
rect 11395 1995 11415 2015
rect 11450 2095 11470 2115
rect 11450 2045 11470 2065
rect 11450 1995 11470 2015
rect 11505 2095 11525 2115
rect 11505 2045 11525 2065
rect 11505 1995 11525 2015
rect 11560 2095 11580 2115
rect 11560 2045 11580 2065
rect 11560 1995 11580 2015
rect 11615 2095 11635 2115
rect 11615 2045 11635 2065
rect 11615 1995 11635 2015
rect 11670 2095 11690 2115
rect 11670 2045 11690 2065
rect 11670 1995 11690 2015
rect 11725 2095 11745 2115
rect 11725 2045 11745 2065
rect 11725 1995 11745 2015
rect 11780 2095 11800 2115
rect 11780 2045 11800 2065
rect 11780 1995 11800 2015
rect 11835 2095 11855 2115
rect 11835 2045 11855 2065
rect 11835 1995 11855 2015
rect 11890 2095 11910 2115
rect 11890 2045 11910 2065
rect 11890 1995 11910 2015
rect 11945 2095 11965 2115
rect 11945 2045 11965 2065
rect 11945 1995 11965 2015
rect 12000 2095 12020 2115
rect 12000 2045 12020 2065
rect 12000 1995 12020 2015
rect 12055 2095 12075 2115
rect 12055 2045 12075 2065
rect 12055 1995 12075 2015
rect 12110 2095 12130 2115
rect 12110 2045 12130 2065
rect 12110 1995 12130 2015
rect 12165 2095 12185 2115
rect 12165 2045 12185 2065
rect 12165 1995 12185 2015
rect 12220 2095 12240 2115
rect 12220 2045 12240 2065
rect 12220 1995 12240 2015
rect 12275 2095 12295 2115
rect 12275 2045 12295 2065
rect 12275 1995 12295 2015
rect 12330 2095 12350 2115
rect 12330 2045 12350 2065
rect 12330 1995 12350 2015
rect 12385 2095 12405 2115
rect 12385 2045 12405 2065
rect 12385 1995 12405 2015
rect 12440 2095 12460 2115
rect 12440 2045 12460 2065
rect 12440 1995 12460 2015
rect 12495 2095 12515 2115
rect 12495 2045 12515 2065
rect 12900 2085 12920 2105
rect 12900 2035 12920 2055
rect 12955 2135 12975 2155
rect 12955 2085 12975 2105
rect 12955 2035 12975 2055
rect 13010 2135 13030 2155
rect 13010 2085 13030 2105
rect 13010 2035 13030 2055
rect 13065 2135 13085 2155
rect 13065 2085 13085 2105
rect 13065 2035 13085 2055
rect 13120 2135 13140 2155
rect 13120 2085 13140 2105
rect 13120 2035 13140 2055
rect 13175 2135 13195 2155
rect 13175 2085 13195 2105
rect 13175 2035 13195 2055
rect 13230 2135 13250 2155
rect 13230 2085 13250 2105
rect 13230 2035 13250 2055
rect 13285 2135 13305 2155
rect 13285 2085 13305 2105
rect 13285 2035 13305 2055
rect 13340 2135 13360 2155
rect 13340 2085 13360 2105
rect 13340 2035 13360 2055
rect 13395 2135 13415 2155
rect 13395 2085 13415 2105
rect 13395 2035 13415 2055
rect 13450 2135 13470 2155
rect 13450 2085 13470 2105
rect 13450 2035 13470 2055
rect 13505 2135 13525 2155
rect 13505 2085 13525 2105
rect 13505 2035 13525 2055
rect 13560 2135 13580 2155
rect 13560 2085 13580 2105
rect 13560 2035 13580 2055
rect 13615 2135 13635 2155
rect 13615 2085 13635 2105
rect 13615 2035 13635 2055
rect 13670 2135 13690 2155
rect 13670 2085 13690 2105
rect 13670 2035 13690 2055
rect 13725 2135 13745 2155
rect 13725 2085 13745 2105
rect 13725 2035 13745 2055
rect 13780 2135 13800 2155
rect 13780 2085 13800 2105
rect 13780 2035 13800 2055
rect 13835 2135 13855 2155
rect 13835 2085 13855 2105
rect 13835 2035 13855 2055
rect 13890 2135 13910 2155
rect 13890 2085 13910 2105
rect 13890 2035 13910 2055
rect 13945 2135 13965 2155
rect 13945 2085 13965 2105
rect 13945 2035 13965 2055
rect 14000 2135 14020 2155
rect 14000 2085 14020 2105
rect 14000 2035 14020 2055
rect 14055 2135 14075 2155
rect 14055 2085 14075 2105
rect 14055 2035 14075 2055
rect 14110 2135 14130 2155
rect 14110 2085 14130 2105
rect 14110 2035 14130 2055
rect 17190 2135 17210 2155
rect 17190 2085 17210 2105
rect 17190 2035 17210 2055
rect 17245 2135 17265 2155
rect 17245 2085 17265 2105
rect 17245 2035 17265 2055
rect 17300 2135 17320 2155
rect 17300 2085 17320 2105
rect 17300 2035 17320 2055
rect 17355 2135 17375 2155
rect 17355 2085 17375 2105
rect 17355 2035 17375 2055
rect 17410 2135 17430 2155
rect 17410 2085 17430 2105
rect 17410 2035 17430 2055
rect 17465 2135 17485 2155
rect 17465 2085 17485 2105
rect 17465 2035 17485 2055
rect 17520 2135 17540 2155
rect 17520 2085 17540 2105
rect 17520 2035 17540 2055
rect 17575 2135 17595 2155
rect 17575 2085 17595 2105
rect 17575 2035 17595 2055
rect 17630 2135 17650 2155
rect 17630 2085 17650 2105
rect 17630 2035 17650 2055
rect 17685 2135 17705 2155
rect 17685 2085 17705 2105
rect 17685 2035 17705 2055
rect 17740 2135 17760 2155
rect 17740 2085 17760 2105
rect 17740 2035 17760 2055
rect 17795 2135 17815 2155
rect 17795 2085 17815 2105
rect 17795 2035 17815 2055
rect 17850 2135 17870 2155
rect 17850 2085 17870 2105
rect 17850 2035 17870 2055
rect 17905 2135 17925 2155
rect 17905 2085 17925 2105
rect 17905 2035 17925 2055
rect 17960 2135 17980 2155
rect 17960 2085 17980 2105
rect 17960 2035 17980 2055
rect 18015 2135 18035 2155
rect 18015 2085 18035 2105
rect 18015 2035 18035 2055
rect 18070 2135 18090 2155
rect 18070 2085 18090 2105
rect 18070 2035 18090 2055
rect 18125 2135 18145 2155
rect 18125 2085 18145 2105
rect 18125 2035 18145 2055
rect 18180 2135 18200 2155
rect 18180 2085 18200 2105
rect 18180 2035 18200 2055
rect 18235 2135 18255 2155
rect 18235 2085 18255 2105
rect 18235 2035 18255 2055
rect 18290 2135 18310 2155
rect 18290 2085 18310 2105
rect 18290 2035 18310 2055
rect 18345 2135 18365 2155
rect 18345 2085 18365 2105
rect 18345 2035 18365 2055
rect 18400 2135 18420 2155
rect 20400 2135 20420 2155
rect 18400 2085 18420 2105
rect 18400 2035 18420 2055
rect 18785 2095 18805 2115
rect 18785 2045 18805 2065
rect 12495 1995 12515 2015
rect 18785 1995 18805 2015
rect 18840 2095 18860 2115
rect 18840 2045 18860 2065
rect 18840 1995 18860 2015
rect 18895 2095 18915 2115
rect 18895 2045 18915 2065
rect 18895 1995 18915 2015
rect 18950 2095 18970 2115
rect 18950 2045 18970 2065
rect 18950 1995 18970 2015
rect 19005 2095 19025 2115
rect 19005 2045 19025 2065
rect 19005 1995 19025 2015
rect 19060 2095 19080 2115
rect 19060 2045 19080 2065
rect 19060 1995 19080 2015
rect 19115 2095 19135 2115
rect 19115 2045 19135 2065
rect 19115 1995 19135 2015
rect 19170 2095 19190 2115
rect 19170 2045 19190 2065
rect 19170 1995 19190 2015
rect 19225 2095 19245 2115
rect 19225 2045 19245 2065
rect 19225 1995 19245 2015
rect 19280 2095 19300 2115
rect 19280 2045 19300 2065
rect 19280 1995 19300 2015
rect 19335 2095 19355 2115
rect 19335 2045 19355 2065
rect 19335 1995 19355 2015
rect 19390 2095 19410 2115
rect 19390 2045 19410 2065
rect 19390 1995 19410 2015
rect 19445 2095 19465 2115
rect 19445 2045 19465 2065
rect 19445 1995 19465 2015
rect 19500 2095 19520 2115
rect 19500 2045 19520 2065
rect 19500 1995 19520 2015
rect 19555 2095 19575 2115
rect 19555 2045 19575 2065
rect 19555 1995 19575 2015
rect 19610 2095 19630 2115
rect 19610 2045 19630 2065
rect 19610 1995 19630 2015
rect 19665 2095 19685 2115
rect 19665 2045 19685 2065
rect 19665 1995 19685 2015
rect 19720 2095 19740 2115
rect 19720 2045 19740 2065
rect 19720 1995 19740 2015
rect 19775 2095 19795 2115
rect 19775 2045 19795 2065
rect 19775 1995 19795 2015
rect 19830 2095 19850 2115
rect 19830 2045 19850 2065
rect 19830 1995 19850 2015
rect 19885 2095 19905 2115
rect 19885 2045 19905 2065
rect 19885 1995 19905 2015
rect 19940 2095 19960 2115
rect 19940 2045 19960 2065
rect 19940 1995 19960 2015
rect 19995 2095 20015 2115
rect 19995 2045 20015 2065
rect 20400 2085 20420 2105
rect 20400 2035 20420 2055
rect 20455 2135 20475 2155
rect 20455 2085 20475 2105
rect 20455 2035 20475 2055
rect 20510 2135 20530 2155
rect 20510 2085 20530 2105
rect 20510 2035 20530 2055
rect 20565 2135 20585 2155
rect 20565 2085 20585 2105
rect 20565 2035 20585 2055
rect 20620 2135 20640 2155
rect 20620 2085 20640 2105
rect 20620 2035 20640 2055
rect 20675 2135 20695 2155
rect 20675 2085 20695 2105
rect 20675 2035 20695 2055
rect 20730 2135 20750 2155
rect 20730 2085 20750 2105
rect 20730 2035 20750 2055
rect 20785 2135 20805 2155
rect 20785 2085 20805 2105
rect 20785 2035 20805 2055
rect 20840 2135 20860 2155
rect 20840 2085 20860 2105
rect 20840 2035 20860 2055
rect 20895 2135 20915 2155
rect 20895 2085 20915 2105
rect 20895 2035 20915 2055
rect 20950 2135 20970 2155
rect 20950 2085 20970 2105
rect 20950 2035 20970 2055
rect 21005 2135 21025 2155
rect 21005 2085 21025 2105
rect 21005 2035 21025 2055
rect 21060 2135 21080 2155
rect 21060 2085 21080 2105
rect 21060 2035 21080 2055
rect 21115 2135 21135 2155
rect 21115 2085 21135 2105
rect 21115 2035 21135 2055
rect 21170 2135 21190 2155
rect 21170 2085 21190 2105
rect 21170 2035 21190 2055
rect 21225 2135 21245 2155
rect 21225 2085 21245 2105
rect 21225 2035 21245 2055
rect 21280 2135 21300 2155
rect 21280 2085 21300 2105
rect 21280 2035 21300 2055
rect 21335 2135 21355 2155
rect 21335 2085 21355 2105
rect 21335 2035 21355 2055
rect 21390 2135 21410 2155
rect 21390 2085 21410 2105
rect 21390 2035 21410 2055
rect 21445 2135 21465 2155
rect 21445 2085 21465 2105
rect 21445 2035 21465 2055
rect 21500 2135 21520 2155
rect 21500 2085 21520 2105
rect 21500 2035 21520 2055
rect 21555 2135 21575 2155
rect 21555 2085 21575 2105
rect 21555 2035 21575 2055
rect 21610 2135 21630 2155
rect 21610 2085 21630 2105
rect 21610 2035 21630 2055
rect 19995 1995 20015 2015
rect 20500 1820 20520 1840
rect 20500 1770 20520 1790
rect 20500 1720 20520 1740
rect 20555 1820 20575 1840
rect 20555 1770 20575 1790
rect 20555 1720 20575 1740
rect 20610 1820 20630 1840
rect 20610 1770 20630 1790
rect 20610 1720 20630 1740
rect 20665 1820 20685 1840
rect 20665 1770 20685 1790
rect 20665 1720 20685 1740
rect 20720 1820 20740 1840
rect 20720 1770 20740 1790
rect 20720 1720 20740 1740
rect 20775 1820 20795 1840
rect 20775 1770 20795 1790
rect 20775 1720 20795 1740
rect 20830 1820 20850 1840
rect 20830 1770 20850 1790
rect 20830 1720 20850 1740
rect 3175 1630 3195 1650
rect 3235 1630 3255 1650
rect 3295 1630 3315 1650
rect 3355 1630 3375 1650
rect 3415 1630 3435 1650
rect 3475 1630 3495 1650
rect 3535 1630 3555 1650
rect 3595 1630 3615 1650
rect 3655 1630 3675 1650
rect 3715 1630 3735 1650
rect 3775 1630 3795 1650
rect 4215 1630 4235 1650
rect 4275 1630 4295 1650
rect 4335 1630 4355 1650
rect 4395 1630 4415 1650
rect 4455 1630 4475 1650
rect 4515 1630 4535 1650
rect 4575 1630 4595 1650
rect 4635 1630 4655 1650
rect 4695 1630 4715 1650
rect 4755 1630 4775 1650
rect 4815 1630 4835 1650
rect 11040 1630 11060 1650
rect 11040 1580 11060 1600
rect 11040 1530 11060 1550
rect 11095 1630 11115 1650
rect 11095 1580 11115 1600
rect 11095 1530 11115 1550
rect 11150 1630 11170 1650
rect 11150 1580 11170 1600
rect 11150 1530 11170 1550
rect 11205 1630 11225 1650
rect 11205 1580 11225 1600
rect 11205 1530 11225 1550
rect 11260 1630 11280 1650
rect 11260 1580 11280 1600
rect 11260 1530 11280 1550
rect 11315 1630 11335 1650
rect 11315 1580 11335 1600
rect 11315 1530 11335 1550
rect 11370 1630 11390 1650
rect 11370 1580 11390 1600
rect 11370 1530 11390 1550
rect 11425 1630 11445 1650
rect 11425 1580 11445 1600
rect 11425 1530 11445 1550
rect 11480 1630 11500 1650
rect 11480 1580 11500 1600
rect 11480 1530 11500 1550
rect 11535 1630 11555 1650
rect 11535 1580 11555 1600
rect 11535 1530 11555 1550
rect 11590 1630 11610 1650
rect 11590 1580 11610 1600
rect 11590 1530 11610 1550
rect 11645 1630 11665 1650
rect 11645 1580 11665 1600
rect 11645 1530 11665 1550
rect 11700 1630 11720 1650
rect 11780 1630 11800 1650
rect 11700 1580 11720 1600
rect 11780 1580 11800 1600
rect 11700 1530 11720 1550
rect 11780 1530 11800 1550
rect 11835 1630 11855 1650
rect 11835 1580 11855 1600
rect 11835 1530 11855 1550
rect 11890 1630 11910 1650
rect 11890 1580 11910 1600
rect 11890 1530 11910 1550
rect 11945 1630 11965 1650
rect 11945 1580 11965 1600
rect 11945 1530 11965 1550
rect 12000 1630 12020 1650
rect 12080 1630 12100 1650
rect 12000 1580 12020 1600
rect 12080 1580 12100 1600
rect 12000 1530 12020 1550
rect 12080 1530 12100 1550
rect 12135 1630 12155 1650
rect 12135 1580 12155 1600
rect 12135 1530 12155 1550
rect 12190 1630 12210 1650
rect 12190 1580 12210 1600
rect 12190 1530 12210 1550
rect 12245 1630 12265 1650
rect 12245 1580 12265 1600
rect 12245 1530 12265 1550
rect 12300 1630 12320 1650
rect 12300 1580 12320 1600
rect 12300 1530 12320 1550
rect 12355 1630 12375 1650
rect 12355 1580 12375 1600
rect 12355 1530 12375 1550
rect 12410 1630 12430 1650
rect 12410 1580 12430 1600
rect 12410 1530 12430 1550
rect 12465 1630 12485 1650
rect 12465 1580 12485 1600
rect 12465 1530 12485 1550
rect 12520 1630 12540 1650
rect 12520 1580 12540 1600
rect 12520 1530 12540 1550
rect 12575 1630 12595 1650
rect 12575 1580 12595 1600
rect 12575 1530 12595 1550
rect 12630 1630 12650 1650
rect 12630 1580 12650 1600
rect 12630 1530 12650 1550
rect 12685 1630 12705 1650
rect 12685 1580 12705 1600
rect 12685 1530 12705 1550
rect 12740 1630 12760 1650
rect 12740 1580 12760 1600
rect 12740 1530 12760 1550
rect 18540 1630 18560 1650
rect 18540 1580 18560 1600
rect 18540 1530 18560 1550
rect 18595 1630 18615 1650
rect 18595 1580 18615 1600
rect 18595 1530 18615 1550
rect 18650 1630 18670 1650
rect 18650 1580 18670 1600
rect 18650 1530 18670 1550
rect 18705 1630 18725 1650
rect 18705 1580 18725 1600
rect 18705 1530 18725 1550
rect 18760 1630 18780 1650
rect 18760 1580 18780 1600
rect 18760 1530 18780 1550
rect 18815 1630 18835 1650
rect 18815 1580 18835 1600
rect 18815 1530 18835 1550
rect 18870 1630 18890 1650
rect 18870 1580 18890 1600
rect 18870 1530 18890 1550
rect 18925 1630 18945 1650
rect 18925 1580 18945 1600
rect 18925 1530 18945 1550
rect 18980 1630 19000 1650
rect 18980 1580 19000 1600
rect 18980 1530 19000 1550
rect 19035 1630 19055 1650
rect 19035 1580 19055 1600
rect 19035 1530 19055 1550
rect 19090 1630 19110 1650
rect 19090 1580 19110 1600
rect 19090 1530 19110 1550
rect 19145 1630 19165 1650
rect 19145 1580 19165 1600
rect 19145 1530 19165 1550
rect 19200 1630 19220 1650
rect 19280 1630 19300 1650
rect 19200 1580 19220 1600
rect 19280 1580 19300 1600
rect 19200 1530 19220 1550
rect 19280 1530 19300 1550
rect 19335 1630 19355 1650
rect 19335 1580 19355 1600
rect 19335 1530 19355 1550
rect 19390 1630 19410 1650
rect 19390 1580 19410 1600
rect 19390 1530 19410 1550
rect 19445 1630 19465 1650
rect 19445 1580 19465 1600
rect 19445 1530 19465 1550
rect 19500 1630 19520 1650
rect 19580 1630 19600 1650
rect 19500 1580 19520 1600
rect 19580 1580 19600 1600
rect 19500 1530 19520 1550
rect 19580 1530 19600 1550
rect 19635 1630 19655 1650
rect 19635 1580 19655 1600
rect 19635 1530 19655 1550
rect 19690 1630 19710 1650
rect 19690 1580 19710 1600
rect 19690 1530 19710 1550
rect 19745 1630 19765 1650
rect 19745 1580 19765 1600
rect 19745 1530 19765 1550
rect 19800 1630 19820 1650
rect 19800 1580 19820 1600
rect 19800 1530 19820 1550
rect 19855 1630 19875 1650
rect 19855 1580 19875 1600
rect 19855 1530 19875 1550
rect 19910 1630 19930 1650
rect 19910 1580 19930 1600
rect 19910 1530 19930 1550
rect 19965 1630 19985 1650
rect 19965 1580 19985 1600
rect 19965 1530 19985 1550
rect 20020 1630 20040 1650
rect 20020 1580 20040 1600
rect 20020 1530 20040 1550
rect 20075 1630 20095 1650
rect 20075 1580 20095 1600
rect 20075 1530 20095 1550
rect 20130 1630 20150 1650
rect 20130 1580 20150 1600
rect 20130 1530 20150 1550
rect 20185 1630 20205 1650
rect 20185 1580 20205 1600
rect 20185 1530 20205 1550
rect 20240 1630 20260 1650
rect 20240 1580 20260 1600
rect 20240 1530 20260 1550
rect 20405 1485 20425 1505
rect 2845 1420 2865 1440
rect 2845 1370 2865 1390
rect 2845 1320 2865 1340
rect 2845 1270 2865 1290
rect 2845 1220 2865 1240
rect 3385 1420 3405 1440
rect 3385 1370 3405 1390
rect 3385 1320 3405 1340
rect 3385 1270 3405 1290
rect 3385 1220 3405 1240
rect 3925 1420 3945 1440
rect 3925 1370 3945 1390
rect 3925 1320 3945 1340
rect 3925 1270 3945 1290
rect 3925 1220 3945 1240
rect 4065 1420 4085 1440
rect 4065 1370 4085 1390
rect 4065 1320 4085 1340
rect 4065 1270 4085 1290
rect 4065 1220 4085 1240
rect 4605 1420 4625 1440
rect 4605 1370 4625 1390
rect 4605 1320 4625 1340
rect 4605 1270 4625 1290
rect 4605 1220 4625 1240
rect 5145 1420 5165 1440
rect 20405 1435 20425 1455
rect 5145 1370 5165 1390
rect 20405 1385 20425 1405
rect 20460 1485 20480 1505
rect 20460 1435 20480 1455
rect 20460 1385 20480 1405
rect 20515 1485 20535 1505
rect 20515 1435 20535 1455
rect 20515 1385 20535 1405
rect 20570 1485 20590 1505
rect 20570 1435 20590 1455
rect 20570 1385 20590 1405
rect 20625 1485 20645 1505
rect 20705 1485 20725 1505
rect 20625 1435 20645 1455
rect 20705 1435 20725 1455
rect 20625 1385 20645 1405
rect 20705 1385 20725 1405
rect 20760 1485 20780 1505
rect 20760 1435 20780 1455
rect 20760 1385 20780 1405
rect 20815 1485 20835 1505
rect 20815 1435 20835 1455
rect 20815 1385 20835 1405
rect 20870 1485 20890 1505
rect 20870 1435 20890 1455
rect 20870 1385 20890 1405
rect 20925 1485 20945 1505
rect 20925 1435 20945 1455
rect 20925 1385 20945 1405
rect 5145 1320 5165 1340
rect 5145 1270 5165 1290
rect 5145 1220 5165 1240
rect 12935 1235 12955 1255
rect 12935 1190 12955 1210
rect 11215 1140 11235 1160
rect 11215 1090 11235 1110
rect 2955 1040 2975 1060
rect 2955 990 2975 1010
rect 3995 1040 4015 1060
rect 3995 990 4015 1010
rect 5035 1040 5055 1060
rect 5035 990 5055 1010
rect 11215 1040 11235 1060
rect 11215 990 11235 1010
rect 11215 940 11235 960
rect 11270 1140 11290 1160
rect 11270 1090 11290 1110
rect 11270 1040 11290 1060
rect 11270 990 11290 1010
rect 11270 940 11290 960
rect 11325 1140 11345 1160
rect 11325 1090 11345 1110
rect 11325 1040 11345 1060
rect 11325 990 11345 1010
rect 11325 940 11345 960
rect 11380 1140 11400 1160
rect 11380 1090 11400 1110
rect 11380 1040 11400 1060
rect 11380 990 11400 1010
rect 11380 940 11400 960
rect 11435 1140 11455 1160
rect 11435 1090 11455 1110
rect 11435 1040 11455 1060
rect 11435 990 11455 1010
rect 11435 940 11455 960
rect 11490 1140 11510 1160
rect 11490 1090 11510 1110
rect 11490 1040 11510 1060
rect 11490 990 11510 1010
rect 11490 940 11510 960
rect 11545 1140 11565 1160
rect 11545 1090 11565 1110
rect 11545 1040 11565 1060
rect 11545 990 11565 1010
rect 11545 940 11565 960
rect 11600 1140 11620 1160
rect 11600 1090 11620 1110
rect 11600 1040 11620 1060
rect 11600 990 11620 1010
rect 11600 940 11620 960
rect 11655 1140 11675 1160
rect 11655 1090 11675 1110
rect 11655 1040 11675 1060
rect 11655 990 11675 1010
rect 11655 940 11675 960
rect 11710 1140 11730 1160
rect 11710 1090 11730 1110
rect 11710 1040 11730 1060
rect 11710 990 11730 1010
rect 11710 940 11730 960
rect 11765 1140 11785 1160
rect 11765 1090 11785 1110
rect 11765 1040 11785 1060
rect 11765 990 11785 1010
rect 11765 940 11785 960
rect 11820 1140 11840 1160
rect 11820 1090 11840 1110
rect 11820 1040 11840 1060
rect 11820 990 11840 1010
rect 11820 940 11840 960
rect 11875 1140 11895 1160
rect 11875 1090 11895 1110
rect 11875 1040 11895 1060
rect 11875 990 11895 1010
rect 11875 940 11895 960
rect 11930 1140 11950 1160
rect 11930 1090 11950 1110
rect 11930 1040 11950 1060
rect 11930 990 11950 1010
rect 11930 940 11950 960
rect 11985 1140 12005 1160
rect 11985 1090 12005 1110
rect 11985 1040 12005 1060
rect 11985 990 12005 1010
rect 11985 940 12005 960
rect 12040 1140 12060 1160
rect 12040 1090 12060 1110
rect 12040 1040 12060 1060
rect 12040 990 12060 1010
rect 12040 940 12060 960
rect 12095 1140 12115 1160
rect 12095 1090 12115 1110
rect 12095 1040 12115 1060
rect 12095 990 12115 1010
rect 12095 940 12115 960
rect 12150 1140 12170 1160
rect 12150 1090 12170 1110
rect 12150 1040 12170 1060
rect 12150 990 12170 1010
rect 12150 940 12170 960
rect 12205 1140 12225 1160
rect 12205 1090 12225 1110
rect 12205 1040 12225 1060
rect 12205 990 12225 1010
rect 12205 940 12225 960
rect 12260 1140 12280 1160
rect 12260 1090 12280 1110
rect 12260 1040 12280 1060
rect 12260 990 12280 1010
rect 12260 940 12280 960
rect 12315 1140 12335 1160
rect 12315 1090 12335 1110
rect 12315 1040 12335 1060
rect 12315 990 12335 1010
rect 12315 940 12335 960
rect 12370 1140 12390 1160
rect 12370 1090 12390 1110
rect 12370 1040 12390 1060
rect 12370 990 12390 1010
rect 12370 940 12390 960
rect 12425 1140 12445 1160
rect 12425 1090 12445 1110
rect 12425 1040 12445 1060
rect 12425 990 12445 1010
rect 12425 940 12445 960
rect 12480 1140 12500 1160
rect 12480 1090 12500 1110
rect 12480 1040 12500 1060
rect 12480 990 12500 1010
rect 12480 940 12500 960
rect 12535 1140 12555 1160
rect 12535 1090 12555 1110
rect 12535 1040 12555 1060
rect 12535 990 12555 1010
rect 12535 940 12555 960
rect 12590 1140 12610 1160
rect 12590 1090 12610 1110
rect 12590 1040 12610 1060
rect 12590 990 12610 1010
rect 12935 1145 12955 1165
rect 12935 1095 12955 1115
rect 12935 1050 12955 1070
rect 12935 1005 12955 1025
rect 13035 1235 13055 1255
rect 13035 1190 13055 1210
rect 13035 1145 13055 1165
rect 13035 1095 13055 1115
rect 13035 1050 13055 1070
rect 13035 1005 13055 1025
rect 13135 1235 13155 1255
rect 13135 1190 13155 1210
rect 13135 1145 13155 1165
rect 13135 1095 13155 1115
rect 13135 1050 13155 1070
rect 13135 1005 13155 1025
rect 13235 1235 13255 1255
rect 13235 1190 13255 1210
rect 13235 1145 13255 1165
rect 13235 1095 13255 1115
rect 13235 1050 13255 1070
rect 13235 1005 13255 1025
rect 13335 1235 13355 1255
rect 13335 1190 13355 1210
rect 13335 1145 13355 1165
rect 13335 1095 13355 1115
rect 13335 1050 13355 1070
rect 13335 1005 13355 1025
rect 13435 1235 13455 1255
rect 13435 1190 13455 1210
rect 13435 1145 13455 1165
rect 13435 1095 13455 1115
rect 13435 1050 13455 1070
rect 13435 1005 13455 1025
rect 13535 1235 13555 1255
rect 13535 1190 13555 1210
rect 13535 1145 13555 1165
rect 13535 1095 13555 1115
rect 13535 1050 13555 1070
rect 13535 1005 13555 1025
rect 13635 1235 13655 1255
rect 13635 1190 13655 1210
rect 13635 1145 13655 1165
rect 13635 1095 13655 1115
rect 13635 1050 13655 1070
rect 13635 1005 13655 1025
rect 13735 1235 13755 1255
rect 13735 1190 13755 1210
rect 13735 1145 13755 1165
rect 13735 1095 13755 1115
rect 13735 1050 13755 1070
rect 13735 1005 13755 1025
rect 13835 1235 13855 1255
rect 13835 1190 13855 1210
rect 13835 1145 13855 1165
rect 13835 1095 13855 1115
rect 13835 1050 13855 1070
rect 13835 1005 13855 1025
rect 13935 1235 13955 1255
rect 13935 1190 13955 1210
rect 13935 1145 13955 1165
rect 13935 1095 13955 1115
rect 13935 1050 13955 1070
rect 13935 1005 13955 1025
rect 14035 1235 14055 1255
rect 14035 1190 14055 1210
rect 14035 1145 14055 1165
rect 14035 1095 14055 1115
rect 14035 1050 14055 1070
rect 14035 1005 14055 1025
rect 14135 1235 14155 1255
rect 14135 1190 14155 1210
rect 14135 1145 14155 1165
rect 14135 1095 14155 1115
rect 14135 1050 14155 1070
rect 14135 1005 14155 1025
rect 18715 1190 18735 1210
rect 18715 1140 18735 1160
rect 18715 1090 18735 1110
rect 18715 1040 18735 1060
rect 18715 990 18735 1010
rect 12590 940 12610 960
rect 18770 1190 18790 1210
rect 18770 1140 18790 1160
rect 18770 1090 18790 1110
rect 18770 1040 18790 1060
rect 18770 990 18790 1010
rect 18825 1190 18845 1210
rect 18825 1140 18845 1160
rect 18825 1090 18845 1110
rect 18825 1040 18845 1060
rect 18825 990 18845 1010
rect 18880 1190 18900 1210
rect 18880 1140 18900 1160
rect 18880 1090 18900 1110
rect 18880 1040 18900 1060
rect 18880 990 18900 1010
rect 18935 1190 18955 1210
rect 18935 1140 18955 1160
rect 18935 1090 18955 1110
rect 18935 1040 18955 1060
rect 18935 990 18955 1010
rect 18990 1190 19010 1210
rect 18990 1140 19010 1160
rect 18990 1090 19010 1110
rect 18990 1040 19010 1060
rect 18990 990 19010 1010
rect 19045 1190 19065 1210
rect 19045 1140 19065 1160
rect 19045 1090 19065 1110
rect 19045 1040 19065 1060
rect 19045 990 19065 1010
rect 19100 1190 19120 1210
rect 19100 1140 19120 1160
rect 19100 1090 19120 1110
rect 19100 1040 19120 1060
rect 19100 990 19120 1010
rect 19155 1190 19175 1210
rect 19155 1140 19175 1160
rect 19155 1090 19175 1110
rect 19155 1040 19175 1060
rect 19155 990 19175 1010
rect 19210 1190 19230 1210
rect 19210 1140 19230 1160
rect 19210 1090 19230 1110
rect 19210 1040 19230 1060
rect 19210 990 19230 1010
rect 19265 1190 19285 1210
rect 19265 1140 19285 1160
rect 19265 1090 19285 1110
rect 19265 1040 19285 1060
rect 19265 990 19285 1010
rect 19320 1190 19340 1210
rect 19320 1140 19340 1160
rect 19320 1090 19340 1110
rect 19320 1040 19340 1060
rect 19320 990 19340 1010
rect 19375 1190 19395 1210
rect 19375 1140 19395 1160
rect 19375 1090 19395 1110
rect 19375 1040 19395 1060
rect 19375 990 19395 1010
rect 19430 1190 19450 1210
rect 19430 1140 19450 1160
rect 19430 1090 19450 1110
rect 19430 1040 19450 1060
rect 19430 990 19450 1010
rect 19485 1190 19505 1210
rect 19485 1140 19505 1160
rect 19485 1090 19505 1110
rect 19485 1040 19505 1060
rect 19485 990 19505 1010
rect 19540 1190 19560 1210
rect 19540 1140 19560 1160
rect 19540 1090 19560 1110
rect 19540 1040 19560 1060
rect 19540 990 19560 1010
rect 19595 1190 19615 1210
rect 19595 1140 19615 1160
rect 19595 1090 19615 1110
rect 19595 1040 19615 1060
rect 19595 990 19615 1010
rect 19650 1190 19670 1210
rect 19650 1140 19670 1160
rect 19650 1090 19670 1110
rect 19650 1040 19670 1060
rect 19650 990 19670 1010
rect 19705 1190 19725 1210
rect 19705 1140 19725 1160
rect 19705 1090 19725 1110
rect 19705 1040 19725 1060
rect 19705 990 19725 1010
rect 19760 1190 19780 1210
rect 19760 1140 19780 1160
rect 19760 1090 19780 1110
rect 19760 1040 19780 1060
rect 19760 990 19780 1010
rect 19815 1190 19835 1210
rect 19815 1140 19835 1160
rect 19815 1090 19835 1110
rect 19815 1040 19835 1060
rect 19815 990 19835 1010
rect 19870 1190 19890 1210
rect 19870 1140 19890 1160
rect 19870 1090 19890 1110
rect 19870 1040 19890 1060
rect 19870 990 19890 1010
rect 19925 1190 19945 1210
rect 19925 1140 19945 1160
rect 19925 1090 19945 1110
rect 19925 1040 19945 1060
rect 19925 990 19945 1010
rect 19980 1190 20000 1210
rect 19980 1140 20000 1160
rect 19980 1090 20000 1110
rect 19980 1040 20000 1060
rect 19980 990 20000 1010
rect 20035 1190 20055 1210
rect 20035 1140 20055 1160
rect 20035 1090 20055 1110
rect 20035 1040 20055 1060
rect 20035 990 20055 1010
rect 20090 1190 20110 1210
rect 20090 1140 20110 1160
rect 20090 1090 20110 1110
rect 20090 1040 20110 1060
rect 20555 1145 20575 1165
rect 20555 1095 20575 1115
rect 20555 1045 20575 1065
rect 20610 1145 20630 1165
rect 20610 1095 20630 1115
rect 20610 1045 20630 1065
rect 20665 1145 20685 1165
rect 20665 1095 20685 1115
rect 20665 1045 20685 1065
rect 20720 1145 20740 1165
rect 20720 1095 20740 1115
rect 20720 1045 20740 1065
rect 20775 1145 20795 1165
rect 20775 1095 20795 1115
rect 20775 1045 20795 1065
rect 20090 990 20110 1010
rect 3005 845 3025 865
rect 3005 795 3025 815
rect 3095 845 3115 865
rect 3095 795 3115 815
rect 3185 845 3205 865
rect 3185 795 3205 815
rect 3275 845 3295 865
rect 3275 795 3295 815
rect 3365 845 3385 865
rect 3365 795 3385 815
rect 3455 845 3475 865
rect 3455 795 3475 815
rect 3545 845 3565 865
rect 3545 795 3565 815
rect 3635 845 3655 865
rect 3635 795 3655 815
rect 3725 845 3745 865
rect 3725 795 3745 815
rect 3815 845 3835 865
rect 3815 795 3835 815
rect 3905 845 3925 865
rect 3905 795 3925 815
rect 3995 845 4015 865
rect 3995 795 4015 815
rect 4085 845 4105 865
rect 4085 795 4105 815
rect 4175 845 4195 865
rect 4175 795 4195 815
rect 4265 845 4285 865
rect 4265 795 4285 815
rect 4355 845 4375 865
rect 4355 795 4375 815
rect 4445 845 4465 865
rect 4445 795 4465 815
rect 4535 845 4555 865
rect 4535 795 4555 815
rect 4625 845 4645 865
rect 4625 795 4645 815
rect 4715 845 4735 865
rect 4715 795 4735 815
rect 4805 845 4825 865
rect 4805 795 4825 815
rect 4895 845 4915 865
rect 4895 795 4915 815
rect 4985 845 5005 865
rect 4985 795 5005 815
rect -2925 -410 -2905 -390
rect 9285 -765 9305 -745
rect 9285 -810 9305 -790
rect 9285 -855 9305 -835
rect 9285 -905 9305 -885
rect 9285 -950 9305 -930
rect 9285 -995 9305 -975
rect 9385 -765 9405 -745
rect 9385 -810 9405 -790
rect 9385 -855 9405 -835
rect 9385 -905 9405 -885
rect 9385 -950 9405 -930
rect 9385 -995 9405 -975
rect 9485 -765 9505 -745
rect 9485 -810 9505 -790
rect 9485 -855 9505 -835
rect 9485 -905 9505 -885
rect 9485 -950 9505 -930
rect 9485 -995 9505 -975
rect 9585 -765 9605 -745
rect 9585 -810 9605 -790
rect 9585 -855 9605 -835
rect 9585 -905 9605 -885
rect 9585 -950 9605 -930
rect 9585 -995 9605 -975
rect 9685 -765 9705 -745
rect 9685 -810 9705 -790
rect 9685 -855 9705 -835
rect 9685 -905 9705 -885
rect 9685 -950 9705 -930
rect 9685 -995 9705 -975
rect 9785 -765 9805 -745
rect 9785 -810 9805 -790
rect 9785 -855 9805 -835
rect 9785 -905 9805 -885
rect 9785 -950 9805 -930
rect 9785 -995 9805 -975
rect 9885 -765 9905 -745
rect 9885 -810 9905 -790
rect 9885 -855 9905 -835
rect 9885 -905 9905 -885
rect 9885 -950 9905 -930
rect 9885 -995 9905 -975
rect 9985 -765 10005 -745
rect 9985 -810 10005 -790
rect 9985 -855 10005 -835
rect 9985 -905 10005 -885
rect 9985 -950 10005 -930
rect 9985 -995 10005 -975
rect 10085 -765 10105 -745
rect 10085 -810 10105 -790
rect 10085 -855 10105 -835
rect 10085 -905 10105 -885
rect 10085 -950 10105 -930
rect 10085 -995 10105 -975
rect 10185 -765 10205 -745
rect 10185 -810 10205 -790
rect 10185 -855 10205 -835
rect 10185 -905 10205 -885
rect 10185 -950 10205 -930
rect 10185 -995 10205 -975
rect 10285 -765 10305 -745
rect 10285 -810 10305 -790
rect 10285 -855 10305 -835
rect 10285 -905 10305 -885
rect 10285 -950 10305 -930
rect 10285 -995 10305 -975
rect 10385 -765 10405 -745
rect 10385 -810 10405 -790
rect 10385 -855 10405 -835
rect 10385 -905 10405 -885
rect 10385 -950 10405 -930
rect 10385 -995 10405 -975
rect 10485 -765 10505 -745
rect 10485 -810 10505 -790
rect 10485 -855 10505 -835
rect 10485 -905 10505 -885
rect 10485 -950 10505 -930
rect 10485 -995 10505 -975
<< pdiffc >>
rect 3005 2895 3025 2915
rect 3005 2845 3025 2865
rect 3095 2895 3115 2915
rect 3095 2845 3115 2865
rect 3185 2895 3205 2915
rect 3185 2845 3205 2865
rect 3275 2895 3295 2915
rect 3275 2845 3295 2865
rect 3365 2895 3385 2915
rect 3365 2845 3385 2865
rect 3455 2895 3475 2915
rect 3455 2845 3475 2865
rect 3545 2895 3565 2915
rect 3545 2845 3565 2865
rect 3635 2895 3655 2915
rect 3635 2845 3655 2865
rect 3725 2895 3745 2915
rect 3725 2845 3745 2865
rect 3815 2895 3835 2915
rect 3815 2845 3835 2865
rect 3905 2895 3925 2915
rect 3905 2845 3925 2865
rect 3995 2895 4015 2915
rect 3995 2845 4015 2865
rect 4085 2895 4105 2915
rect 4085 2845 4105 2865
rect 4175 2895 4195 2915
rect 4175 2845 4195 2865
rect 4265 2895 4285 2915
rect 4265 2845 4285 2865
rect 4355 2895 4375 2915
rect 4355 2845 4375 2865
rect 4445 2895 4465 2915
rect 4445 2845 4465 2865
rect 4535 2895 4555 2915
rect 4535 2845 4555 2865
rect 4625 2895 4645 2915
rect 4625 2845 4645 2865
rect 4715 2895 4735 2915
rect 4715 2845 4735 2865
rect 4805 2895 4825 2915
rect 4805 2845 4825 2865
rect 4895 2895 4915 2915
rect 4895 2845 4915 2865
rect 4985 2895 5005 2915
rect 4985 2845 5005 2865
rect 3185 2665 3205 2685
rect 3185 2615 3205 2635
rect 3185 2565 3205 2585
rect 3185 2515 3205 2535
rect 3185 2465 3205 2485
rect 3185 2415 3205 2435
rect 3275 2665 3295 2685
rect 3275 2615 3295 2635
rect 3275 2565 3295 2585
rect 3275 2515 3295 2535
rect 3275 2465 3295 2485
rect 3275 2415 3295 2435
rect 3365 2665 3385 2685
rect 3365 2615 3385 2635
rect 3365 2565 3385 2585
rect 3365 2515 3385 2535
rect 3365 2465 3385 2485
rect 3365 2415 3385 2435
rect 3455 2665 3475 2685
rect 3455 2615 3475 2635
rect 3455 2565 3475 2585
rect 3455 2515 3475 2535
rect 3455 2465 3475 2485
rect 3455 2415 3475 2435
rect 3545 2665 3565 2685
rect 3545 2615 3565 2635
rect 3545 2565 3565 2585
rect 3545 2515 3565 2535
rect 3545 2465 3565 2485
rect 3545 2415 3565 2435
rect 3635 2665 3655 2685
rect 3635 2615 3655 2635
rect 3635 2565 3655 2585
rect 3635 2515 3655 2535
rect 3635 2465 3655 2485
rect 3635 2415 3655 2435
rect 3725 2665 3745 2685
rect 3725 2615 3745 2635
rect 3725 2565 3745 2585
rect 3725 2515 3745 2535
rect 3725 2465 3745 2485
rect 3725 2415 3745 2435
rect 3815 2665 3835 2685
rect 3815 2615 3835 2635
rect 3815 2565 3835 2585
rect 3815 2515 3835 2535
rect 3815 2465 3835 2485
rect 3815 2415 3835 2435
rect 3905 2665 3925 2685
rect 3905 2615 3925 2635
rect 3905 2565 3925 2585
rect 3905 2515 3925 2535
rect 3905 2465 3925 2485
rect 3905 2415 3925 2435
rect 3995 2665 4015 2685
rect 3995 2615 4015 2635
rect 3995 2565 4015 2585
rect 3995 2515 4015 2535
rect 3995 2465 4015 2485
rect 3995 2415 4015 2435
rect 4085 2665 4105 2685
rect 4085 2615 4105 2635
rect 4085 2565 4105 2585
rect 4085 2515 4105 2535
rect 4085 2465 4105 2485
rect 4085 2415 4105 2435
rect 4175 2665 4195 2685
rect 4175 2615 4195 2635
rect 4175 2565 4195 2585
rect 4175 2515 4195 2535
rect 4175 2465 4195 2485
rect 4175 2415 4195 2435
rect 4265 2665 4285 2685
rect 4265 2615 4285 2635
rect 4265 2565 4285 2585
rect 4265 2515 4285 2535
rect 4265 2465 4285 2485
rect 4265 2415 4285 2435
rect 4355 2665 4375 2685
rect 4355 2615 4375 2635
rect 4355 2565 4375 2585
rect 4355 2515 4375 2535
rect 4355 2465 4375 2485
rect 4355 2415 4375 2435
rect 4445 2665 4465 2685
rect 4445 2615 4465 2635
rect 4445 2565 4465 2585
rect 4445 2515 4465 2535
rect 4445 2465 4465 2485
rect 4445 2415 4465 2435
rect 4535 2665 4555 2685
rect 4535 2615 4555 2635
rect 4535 2565 4555 2585
rect 4535 2515 4555 2535
rect 4535 2465 4555 2485
rect 4535 2415 4555 2435
rect 4625 2665 4645 2685
rect 4625 2615 4645 2635
rect 4625 2565 4645 2585
rect 4625 2515 4645 2535
rect 4625 2465 4645 2485
rect 4625 2415 4645 2435
rect 4715 2665 4735 2685
rect 4715 2615 4735 2635
rect 4715 2565 4735 2585
rect 4715 2515 4735 2535
rect 4715 2465 4735 2485
rect 4715 2415 4735 2435
rect 4805 2665 4825 2685
rect 4805 2615 4825 2635
rect 4805 2565 4825 2585
rect 4805 2515 4825 2535
rect 4805 2465 4825 2485
rect 4805 2415 4825 2435
rect 2575 1965 2595 1985
rect 2575 1915 2595 1935
rect 2630 1965 2650 1985
rect 2630 1915 2650 1935
rect 2685 1965 2705 1985
rect 2685 1915 2705 1935
rect 2755 1965 2775 1985
rect 2755 1915 2775 1935
rect 2815 1965 2835 1985
rect 2815 1915 2835 1935
rect 2875 1965 2895 1985
rect 2875 1915 2895 1935
rect 2935 1965 2955 1985
rect 2935 1915 2955 1935
rect 2995 1965 3015 1985
rect 2995 1915 3015 1935
rect 3055 1965 3075 1985
rect 3055 1915 3075 1935
rect 3115 1965 3135 1985
rect 3115 1915 3135 1935
rect 3175 1965 3195 1985
rect 3175 1915 3195 1935
rect 3235 1965 3255 1985
rect 3235 1915 3255 1935
rect 3295 1965 3315 1985
rect 3295 1915 3315 1935
rect 3355 1965 3375 1985
rect 3355 1915 3375 1935
rect 3415 1965 3435 1985
rect 3415 1915 3435 1935
rect 3475 1965 3495 1985
rect 3475 1915 3495 1935
rect 3535 1965 3555 1985
rect 3535 1915 3555 1935
rect 3595 1965 3615 1985
rect 3595 1915 3615 1935
rect 3655 1965 3675 1985
rect 3655 1915 3675 1935
rect 3715 1965 3735 1985
rect 3715 1915 3735 1935
rect 3775 1965 3795 1985
rect 3775 1915 3795 1935
rect 3835 1965 3855 1985
rect 3835 1915 3855 1935
rect 3895 1965 3915 1985
rect 3895 1915 3915 1935
rect 3955 1965 3975 1985
rect 4035 1965 4055 1985
rect 3955 1915 3975 1935
rect 4035 1915 4055 1935
rect 4095 1965 4115 1985
rect 4095 1915 4115 1935
rect 4155 1965 4175 1985
rect 4155 1915 4175 1935
rect 4215 1965 4235 1985
rect 4215 1915 4235 1935
rect 4275 1965 4295 1985
rect 4275 1915 4295 1935
rect 4335 1965 4355 1985
rect 4335 1915 4355 1935
rect 4395 1965 4415 1985
rect 4395 1915 4415 1935
rect 4455 1965 4475 1985
rect 4455 1915 4475 1935
rect 4515 1965 4535 1985
rect 4515 1915 4535 1935
rect 4575 1965 4595 1985
rect 4575 1915 4595 1935
rect 4635 1965 4655 1985
rect 4635 1915 4655 1935
rect 4695 1965 4715 1985
rect 4695 1915 4715 1935
rect 4755 1965 4775 1985
rect 4755 1915 4775 1935
rect 4815 1965 4835 1985
rect 4815 1915 4835 1935
rect 4875 1965 4895 1985
rect 4875 1915 4895 1935
rect 4935 1965 4955 1985
rect 4935 1915 4955 1935
rect 4995 1965 5015 1985
rect 4995 1915 5015 1935
rect 5055 1965 5075 1985
rect 5055 1915 5075 1935
rect 5115 1965 5135 1985
rect 5115 1915 5135 1935
rect 5175 1965 5195 1985
rect 5175 1915 5195 1935
rect 5235 1965 5255 1985
rect 5235 1915 5255 1935
<< psubdiff >>
rect 10780 3515 10820 3550
rect 10780 3495 10790 3515
rect 10810 3495 10820 3515
rect 10780 3465 10820 3495
rect 10780 3445 10790 3465
rect 10810 3445 10820 3465
rect 10780 3415 10820 3445
rect 10780 3395 10790 3415
rect 10810 3395 10820 3415
rect 10780 3365 10820 3395
rect 10780 3345 10790 3365
rect 10810 3345 10820 3365
rect 10780 3315 10820 3345
rect 10780 3295 10790 3315
rect 10810 3295 10820 3315
rect 10450 3265 10490 3293
rect 10450 3245 10460 3265
rect 10480 3245 10490 3265
rect 10450 3230 10490 3245
rect 10710 3265 10750 3293
rect 10710 3245 10720 3265
rect 10740 3245 10750 3265
rect 10710 3230 10750 3245
rect 10780 3265 10820 3295
rect 10780 3245 10790 3265
rect 10810 3245 10820 3265
rect 10780 3230 10820 3245
rect 11100 3565 11140 3580
rect 11100 3545 11110 3565
rect 11130 3545 11140 3565
rect 11100 3515 11140 3545
rect 11100 3495 11110 3515
rect 11130 3495 11140 3515
rect 11100 3465 11140 3495
rect 11100 3445 11110 3465
rect 11130 3445 11140 3465
rect 11100 3415 11140 3445
rect 11100 3395 11110 3415
rect 11130 3395 11140 3415
rect 11100 3365 11140 3395
rect 11100 3345 11110 3365
rect 11130 3345 11140 3365
rect 11100 3315 11140 3345
rect 11100 3295 11110 3315
rect 11130 3295 11140 3315
rect 11100 3265 11140 3295
rect 11100 3245 11110 3265
rect 11130 3245 11140 3265
rect 11100 3230 11140 3245
rect 11180 3560 11220 3575
rect 11180 3540 11190 3560
rect 11210 3540 11220 3560
rect 11180 3510 11220 3540
rect 11180 3490 11190 3510
rect 11210 3490 11220 3510
rect 11180 3460 11220 3490
rect 11180 3440 11190 3460
rect 11210 3440 11220 3460
rect 11180 3410 11220 3440
rect 11180 3390 11190 3410
rect 11210 3390 11220 3410
rect 11180 3360 11220 3390
rect 11180 3340 11190 3360
rect 11210 3340 11220 3360
rect 11180 3310 11220 3340
rect 11180 3290 11190 3310
rect 11210 3290 11220 3310
rect 11180 3260 11220 3290
rect 11180 3240 11190 3260
rect 11210 3240 11220 3260
rect 11180 3210 11220 3240
rect 11180 3190 11190 3210
rect 11210 3190 11220 3210
rect 11180 3175 11220 3190
rect 12580 3560 12620 3575
rect 12580 3540 12590 3560
rect 12610 3540 12620 3560
rect 12580 3510 12620 3540
rect 12580 3490 12590 3510
rect 12610 3490 12620 3510
rect 12580 3460 12620 3490
rect 12580 3440 12590 3460
rect 12610 3440 12620 3460
rect 12580 3410 12620 3440
rect 12580 3390 12590 3410
rect 12610 3390 12620 3410
rect 12580 3360 12620 3390
rect 12580 3340 12590 3360
rect 12610 3340 12620 3360
rect 18280 3515 18320 3550
rect 18280 3495 18290 3515
rect 18310 3495 18320 3515
rect 18280 3465 18320 3495
rect 18280 3445 18290 3465
rect 18310 3445 18320 3465
rect 18280 3415 18320 3445
rect 18280 3395 18290 3415
rect 18310 3395 18320 3415
rect 18280 3365 18320 3395
rect 12580 3310 12620 3340
rect 12580 3290 12590 3310
rect 12610 3290 12620 3310
rect 18280 3345 18290 3365
rect 18310 3345 18320 3365
rect 18280 3315 18320 3345
rect 18280 3295 18290 3315
rect 18310 3295 18320 3315
rect 12580 3260 12620 3290
rect 12580 3240 12590 3260
rect 12610 3240 12620 3260
rect 17950 3265 17990 3293
rect 17950 3245 17960 3265
rect 17980 3245 17990 3265
rect 12580 3210 12620 3240
rect 12580 3190 12590 3210
rect 12610 3190 12620 3210
rect 12580 3175 12620 3190
rect 12850 3225 12890 3240
rect 12850 3205 12860 3225
rect 12880 3205 12890 3225
rect 12850 3175 12890 3205
rect 12850 3155 12860 3175
rect 12880 3155 12890 3175
rect 12850 3125 12890 3155
rect 12850 3105 12860 3125
rect 12880 3105 12890 3125
rect 12850 3075 12890 3105
rect 12850 3055 12860 3075
rect 12880 3055 12890 3075
rect 12850 3025 12890 3055
rect 12850 3005 12860 3025
rect 12880 3005 12890 3025
rect 12850 2975 12890 3005
rect 12850 2955 12860 2975
rect 12880 2955 12890 2975
rect 905 2910 1125 2920
rect 905 2880 920 2910
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1125 2910
rect 905 2870 1125 2880
rect 12850 2940 12890 2955
rect 14140 3225 14180 3240
rect 17950 3230 17990 3245
rect 18210 3265 18250 3293
rect 18210 3245 18220 3265
rect 18240 3245 18250 3265
rect 18210 3230 18250 3245
rect 18280 3265 18320 3295
rect 18280 3245 18290 3265
rect 18310 3245 18320 3265
rect 18280 3230 18320 3245
rect 18600 3565 18640 3580
rect 18600 3545 18610 3565
rect 18630 3545 18640 3565
rect 18600 3515 18640 3545
rect 18600 3495 18610 3515
rect 18630 3495 18640 3515
rect 18600 3465 18640 3495
rect 18600 3445 18610 3465
rect 18630 3445 18640 3465
rect 18600 3415 18640 3445
rect 18600 3395 18610 3415
rect 18630 3395 18640 3415
rect 18600 3365 18640 3395
rect 18600 3345 18610 3365
rect 18630 3345 18640 3365
rect 18600 3315 18640 3345
rect 18600 3295 18610 3315
rect 18630 3295 18640 3315
rect 18600 3265 18640 3295
rect 18600 3245 18610 3265
rect 18630 3245 18640 3265
rect 18600 3230 18640 3245
rect 18680 3560 18720 3575
rect 18680 3540 18690 3560
rect 18710 3540 18720 3560
rect 18680 3510 18720 3540
rect 18680 3490 18690 3510
rect 18710 3490 18720 3510
rect 18680 3460 18720 3490
rect 18680 3440 18690 3460
rect 18710 3440 18720 3460
rect 18680 3410 18720 3440
rect 18680 3390 18690 3410
rect 18710 3390 18720 3410
rect 18680 3360 18720 3390
rect 18680 3340 18690 3360
rect 18710 3340 18720 3360
rect 18680 3310 18720 3340
rect 18680 3290 18690 3310
rect 18710 3290 18720 3310
rect 18680 3260 18720 3290
rect 18680 3240 18690 3260
rect 18710 3240 18720 3260
rect 14140 3205 14150 3225
rect 14170 3205 14180 3225
rect 14140 3175 14180 3205
rect 18680 3210 18720 3240
rect 18680 3190 18690 3210
rect 18710 3190 18720 3210
rect 18680 3175 18720 3190
rect 20080 3560 20120 3575
rect 20080 3540 20090 3560
rect 20110 3540 20120 3560
rect 20080 3510 20120 3540
rect 20080 3490 20090 3510
rect 20110 3490 20120 3510
rect 20080 3460 20120 3490
rect 20080 3440 20090 3460
rect 20110 3440 20120 3460
rect 20080 3410 20120 3440
rect 20080 3390 20090 3410
rect 20110 3390 20120 3410
rect 20080 3360 20120 3390
rect 20080 3340 20090 3360
rect 20110 3340 20120 3360
rect 20080 3310 20120 3340
rect 20080 3290 20090 3310
rect 20110 3290 20120 3310
rect 20080 3260 20120 3290
rect 20080 3240 20090 3260
rect 20110 3240 20120 3260
rect 20080 3210 20120 3240
rect 20080 3190 20090 3210
rect 20110 3190 20120 3210
rect 20080 3175 20120 3190
rect 20350 3225 20390 3240
rect 20350 3205 20360 3225
rect 20380 3205 20390 3225
rect 20350 3175 20390 3205
rect 14140 3155 14150 3175
rect 14170 3155 14180 3175
rect 14140 3125 14180 3155
rect 20350 3155 20360 3175
rect 20380 3155 20390 3175
rect 14140 3105 14150 3125
rect 14170 3105 14180 3125
rect 20350 3125 20390 3155
rect 14140 3075 14180 3105
rect 14140 3055 14150 3075
rect 14170 3055 14180 3075
rect 14140 3025 14180 3055
rect 14140 3005 14150 3025
rect 14170 3005 14180 3025
rect 14140 2975 14180 3005
rect 14140 2955 14150 2975
rect 14170 2955 14180 2975
rect 14140 2940 14180 2955
rect 20350 3105 20360 3125
rect 20380 3105 20390 3125
rect 20350 3075 20390 3105
rect 20350 3055 20360 3075
rect 20380 3055 20390 3075
rect 20350 3025 20390 3055
rect 20350 3005 20360 3025
rect 20380 3005 20390 3025
rect 20350 2975 20390 3005
rect 20350 2955 20360 2975
rect 20380 2955 20390 2975
rect 11180 2880 11220 2895
rect 11180 2860 11190 2880
rect 11210 2860 11220 2880
rect 11180 2830 11220 2860
rect 11180 2810 11190 2830
rect 11210 2810 11220 2830
rect 11180 2780 11220 2810
rect 11180 2760 11190 2780
rect 11210 2760 11220 2780
rect 11180 2730 11220 2760
rect 11180 2710 11190 2730
rect 11210 2710 11220 2730
rect 11180 2680 11220 2710
rect 11180 2660 11190 2680
rect 11210 2660 11220 2680
rect 11180 2630 11220 2660
rect 9640 2605 9680 2620
rect 9640 2585 9650 2605
rect 9670 2585 9680 2605
rect 9640 2555 9680 2585
rect 9640 2535 9650 2555
rect 9670 2535 9680 2555
rect 9640 2520 9680 2535
rect 10930 2605 10970 2620
rect 10930 2585 10940 2605
rect 10960 2585 10970 2605
rect 10930 2555 10970 2585
rect 10930 2535 10940 2555
rect 10960 2535 10970 2555
rect 10930 2520 10970 2535
rect 11180 2610 11190 2630
rect 11210 2610 11220 2630
rect 11180 2580 11220 2610
rect 11180 2560 11190 2580
rect 11210 2560 11220 2580
rect 11180 2530 11220 2560
rect 11180 2510 11190 2530
rect 11210 2510 11220 2530
rect 11180 2495 11220 2510
rect 12580 2880 12620 2895
rect 20350 2940 20390 2955
rect 21640 3225 21680 3240
rect 21640 3205 21650 3225
rect 21670 3205 21680 3225
rect 21640 3175 21680 3205
rect 21640 3155 21650 3175
rect 21670 3155 21680 3175
rect 21640 3125 21680 3155
rect 21640 3105 21650 3125
rect 21670 3105 21680 3125
rect 21640 3075 21680 3105
rect 21640 3055 21650 3075
rect 21670 3055 21680 3075
rect 21640 3025 21680 3055
rect 21640 3005 21650 3025
rect 21670 3005 21680 3025
rect 21640 2975 21680 3005
rect 21640 2955 21650 2975
rect 21670 2955 21680 2975
rect 21640 2940 21680 2955
rect 12580 2860 12590 2880
rect 12610 2860 12620 2880
rect 12580 2830 12620 2860
rect 18680 2880 18720 2895
rect 18680 2860 18690 2880
rect 18710 2860 18720 2880
rect 12580 2810 12590 2830
rect 12610 2810 12620 2830
rect 12580 2780 12620 2810
rect 12580 2760 12590 2780
rect 12610 2760 12620 2780
rect 12580 2730 12620 2760
rect 12580 2710 12590 2730
rect 12610 2710 12620 2730
rect 12580 2680 12620 2710
rect 18680 2830 18720 2860
rect 18680 2810 18690 2830
rect 18710 2810 18720 2830
rect 18680 2780 18720 2810
rect 18680 2760 18690 2780
rect 18710 2760 18720 2780
rect 18680 2730 18720 2760
rect 18680 2710 18690 2730
rect 18710 2710 18720 2730
rect 12580 2660 12590 2680
rect 12610 2660 12620 2680
rect 12580 2630 12620 2660
rect 18680 2680 18720 2710
rect 18680 2660 18690 2680
rect 18710 2660 18720 2680
rect 12580 2610 12590 2630
rect 12610 2610 12620 2630
rect 18680 2630 18720 2660
rect 12580 2580 12620 2610
rect 12580 2560 12590 2580
rect 12610 2560 12620 2580
rect 12580 2530 12620 2560
rect 12580 2510 12590 2530
rect 12610 2510 12620 2530
rect 12850 2605 12890 2620
rect 12850 2585 12860 2605
rect 12880 2585 12890 2605
rect 12850 2555 12890 2585
rect 12850 2535 12860 2555
rect 12880 2535 12890 2555
rect 12850 2520 12890 2535
rect 14140 2605 14180 2620
rect 14140 2585 14150 2605
rect 14170 2585 14180 2605
rect 14140 2555 14180 2585
rect 14140 2535 14150 2555
rect 14170 2535 14180 2555
rect 14140 2520 14180 2535
rect 17140 2605 17180 2620
rect 17140 2585 17150 2605
rect 17170 2585 17180 2605
rect 17140 2555 17180 2585
rect 17140 2535 17150 2555
rect 17170 2535 17180 2555
rect 17140 2520 17180 2535
rect 18430 2605 18470 2620
rect 18430 2585 18440 2605
rect 18460 2585 18470 2605
rect 18430 2555 18470 2585
rect 18430 2535 18440 2555
rect 18460 2535 18470 2555
rect 18430 2520 18470 2535
rect 18680 2610 18690 2630
rect 18710 2610 18720 2630
rect 18680 2580 18720 2610
rect 18680 2560 18690 2580
rect 18710 2560 18720 2580
rect 18680 2530 18720 2560
rect 12580 2495 12620 2510
rect 18680 2510 18690 2530
rect 18710 2510 18720 2530
rect 18680 2495 18720 2510
rect 20080 2880 20120 2895
rect 20080 2860 20090 2880
rect 20110 2860 20120 2880
rect 20080 2830 20120 2860
rect 20080 2810 20090 2830
rect 20110 2810 20120 2830
rect 20080 2780 20120 2810
rect 20080 2760 20090 2780
rect 20110 2760 20120 2780
rect 20080 2730 20120 2760
rect 20080 2710 20090 2730
rect 20110 2710 20120 2730
rect 20080 2680 20120 2710
rect 20080 2660 20090 2680
rect 20110 2660 20120 2680
rect 20080 2630 20120 2660
rect 20080 2610 20090 2630
rect 20110 2610 20120 2630
rect 20080 2580 20120 2610
rect 20080 2560 20090 2580
rect 20110 2560 20120 2580
rect 20080 2530 20120 2560
rect 20080 2510 20090 2530
rect 20110 2510 20120 2530
rect 20350 2605 20390 2620
rect 20350 2585 20360 2605
rect 20380 2585 20390 2605
rect 20350 2555 20390 2585
rect 20350 2535 20360 2555
rect 20380 2535 20390 2555
rect 20350 2520 20390 2535
rect 21640 2605 21680 2620
rect 21640 2585 21650 2605
rect 21670 2585 21680 2605
rect 21640 2555 21680 2585
rect 21640 2535 21650 2555
rect 21670 2535 21680 2555
rect 21640 2520 21680 2535
rect 20080 2495 20120 2510
rect 9640 2155 9680 2170
rect 9640 2135 9650 2155
rect 9670 2135 9680 2155
rect 9640 2105 9680 2135
rect 9640 2085 9650 2105
rect 9670 2085 9680 2105
rect 9640 2055 9680 2085
rect 9640 2035 9650 2055
rect 9670 2035 9680 2055
rect 9640 2020 9680 2035
rect 10930 2155 10970 2170
rect 12850 2155 12890 2170
rect 10930 2135 10940 2155
rect 10960 2135 10970 2155
rect 10930 2105 10970 2135
rect 12850 2135 12860 2155
rect 12880 2135 12890 2155
rect 10930 2085 10940 2105
rect 10960 2085 10970 2105
rect 10930 2055 10970 2085
rect 10930 2035 10940 2055
rect 10960 2035 10970 2055
rect 10930 2020 10970 2035
rect 11235 2115 11275 2130
rect 11235 2095 11245 2115
rect 11265 2095 11275 2115
rect 11235 2065 11275 2095
rect 11235 2045 11245 2065
rect 11265 2045 11275 2065
rect 11235 2015 11275 2045
rect 11235 1995 11245 2015
rect 11265 1995 11275 2015
rect 11235 1980 11275 1995
rect 12525 2115 12565 2130
rect 12525 2095 12535 2115
rect 12555 2095 12565 2115
rect 12525 2065 12565 2095
rect 12525 2045 12535 2065
rect 12555 2045 12565 2065
rect 12525 2015 12565 2045
rect 12850 2105 12890 2135
rect 12850 2085 12860 2105
rect 12880 2085 12890 2105
rect 12850 2055 12890 2085
rect 12850 2035 12860 2055
rect 12880 2035 12890 2055
rect 12850 2020 12890 2035
rect 14140 2155 14180 2170
rect 14140 2135 14150 2155
rect 14170 2135 14180 2155
rect 14140 2105 14180 2135
rect 14140 2085 14150 2105
rect 14170 2085 14180 2105
rect 14140 2055 14180 2085
rect 14140 2035 14150 2055
rect 14170 2035 14180 2055
rect 14140 2020 14180 2035
rect 17140 2155 17180 2170
rect 17140 2135 17150 2155
rect 17170 2135 17180 2155
rect 17140 2105 17180 2135
rect 17140 2085 17150 2105
rect 17170 2085 17180 2105
rect 17140 2055 17180 2085
rect 17140 2035 17150 2055
rect 17170 2035 17180 2055
rect 17140 2020 17180 2035
rect 18430 2155 18470 2170
rect 20350 2155 20390 2170
rect 18430 2135 18440 2155
rect 18460 2135 18470 2155
rect 18430 2105 18470 2135
rect 20350 2135 20360 2155
rect 20380 2135 20390 2155
rect 18430 2085 18440 2105
rect 18460 2085 18470 2105
rect 18430 2055 18470 2085
rect 18430 2035 18440 2055
rect 18460 2035 18470 2055
rect 18430 2020 18470 2035
rect 18735 2115 18775 2130
rect 18735 2095 18745 2115
rect 18765 2095 18775 2115
rect 18735 2065 18775 2095
rect 18735 2045 18745 2065
rect 18765 2045 18775 2065
rect 12525 1995 12535 2015
rect 12555 1995 12565 2015
rect 18735 2015 18775 2045
rect 12525 1980 12565 1995
rect 18735 1995 18745 2015
rect 18765 1995 18775 2015
rect 18735 1980 18775 1995
rect 20025 2115 20065 2130
rect 20025 2095 20035 2115
rect 20055 2095 20065 2115
rect 20025 2065 20065 2095
rect 20025 2045 20035 2065
rect 20055 2045 20065 2065
rect 20025 2015 20065 2045
rect 20350 2105 20390 2135
rect 20350 2085 20360 2105
rect 20380 2085 20390 2105
rect 20350 2055 20390 2085
rect 20350 2035 20360 2055
rect 20380 2035 20390 2055
rect 20350 2020 20390 2035
rect 21640 2155 21680 2170
rect 21640 2135 21650 2155
rect 21670 2135 21680 2155
rect 21640 2105 21680 2135
rect 21640 2085 21650 2105
rect 21670 2085 21680 2105
rect 21640 2055 21680 2085
rect 21640 2035 21650 2055
rect 21670 2035 21680 2055
rect 21640 2020 21680 2035
rect 20025 1995 20035 2015
rect 20055 1995 20065 2015
rect 20025 1980 20065 1995
rect 20450 1840 20490 1855
rect 20450 1820 20460 1840
rect 20480 1820 20490 1840
rect 20450 1790 20490 1820
rect 20450 1770 20460 1790
rect 20480 1770 20490 1790
rect -50 1715 100 1730
rect -50 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 100 1715
rect 20450 1740 20490 1770
rect 20450 1720 20460 1740
rect 20480 1720 20490 1740
rect -50 1680 100 1695
rect 20450 1705 20490 1720
rect 20860 1840 20900 1855
rect 20860 1820 20870 1840
rect 20890 1820 20900 1840
rect 20860 1790 20900 1820
rect 20860 1770 20870 1790
rect 20890 1770 20900 1790
rect 20860 1740 20900 1770
rect 20860 1720 20870 1740
rect 20890 1720 20900 1740
rect 20860 1705 20900 1720
rect 3980 1650 4030 1665
rect 3980 1630 3995 1650
rect 4015 1630 4030 1650
rect 3980 1615 4030 1630
rect 10990 1650 11030 1665
rect 10990 1630 11000 1650
rect 11020 1630 11030 1650
rect 10990 1600 11030 1630
rect 10990 1580 11000 1600
rect 11020 1580 11030 1600
rect 10990 1550 11030 1580
rect 10990 1530 11000 1550
rect 11020 1530 11030 1550
rect 10990 1515 11030 1530
rect 11730 1650 11770 1665
rect 11730 1630 11740 1650
rect 11760 1630 11770 1650
rect 11730 1600 11770 1630
rect 11730 1580 11740 1600
rect 11760 1580 11770 1600
rect 11730 1550 11770 1580
rect 11730 1530 11740 1550
rect 11760 1530 11770 1550
rect 11730 1515 11770 1530
rect 12030 1650 12070 1665
rect 12030 1630 12040 1650
rect 12060 1630 12070 1650
rect 12030 1600 12070 1630
rect 12030 1580 12040 1600
rect 12060 1580 12070 1600
rect 12030 1550 12070 1580
rect 12030 1530 12040 1550
rect 12060 1530 12070 1550
rect 12030 1515 12070 1530
rect 12770 1650 12810 1665
rect 12770 1630 12780 1650
rect 12800 1630 12810 1650
rect 12770 1600 12810 1630
rect 12770 1580 12780 1600
rect 12800 1580 12810 1600
rect 12770 1550 12810 1580
rect 12770 1530 12780 1550
rect 12800 1530 12810 1550
rect 12770 1515 12810 1530
rect 18490 1650 18530 1665
rect 18490 1630 18500 1650
rect 18520 1630 18530 1650
rect 18490 1600 18530 1630
rect 18490 1580 18500 1600
rect 18520 1580 18530 1600
rect 18490 1550 18530 1580
rect 18490 1530 18500 1550
rect 18520 1530 18530 1550
rect 18490 1515 18530 1530
rect 19230 1650 19270 1665
rect 19230 1630 19240 1650
rect 19260 1630 19270 1650
rect 19230 1600 19270 1630
rect 19230 1580 19240 1600
rect 19260 1580 19270 1600
rect 19230 1550 19270 1580
rect 19230 1530 19240 1550
rect 19260 1530 19270 1550
rect 19230 1515 19270 1530
rect 19530 1650 19570 1665
rect 19530 1630 19540 1650
rect 19560 1630 19570 1650
rect 19530 1600 19570 1630
rect 19530 1580 19540 1600
rect 19560 1580 19570 1600
rect 19530 1550 19570 1580
rect 19530 1530 19540 1550
rect 19560 1530 19570 1550
rect 19530 1515 19570 1530
rect 20270 1650 20310 1665
rect 20270 1630 20280 1650
rect 20300 1630 20310 1650
rect 20270 1600 20310 1630
rect 20270 1580 20280 1600
rect 20300 1580 20310 1600
rect 20270 1550 20310 1580
rect 20270 1530 20280 1550
rect 20300 1530 20310 1550
rect 20270 1515 20310 1530
rect 20355 1505 20395 1520
rect 20355 1485 20365 1505
rect 20385 1485 20395 1505
rect 20355 1455 20395 1485
rect 20355 1435 20365 1455
rect 20385 1435 20395 1455
rect 20355 1405 20395 1435
rect 20355 1385 20365 1405
rect 20385 1385 20395 1405
rect 20355 1370 20395 1385
rect 20655 1505 20695 1520
rect 20655 1485 20665 1505
rect 20685 1485 20695 1505
rect 20655 1455 20695 1485
rect 20655 1435 20665 1455
rect 20685 1435 20695 1455
rect 20655 1405 20695 1435
rect 20655 1385 20665 1405
rect 20685 1385 20695 1405
rect 20655 1370 20695 1385
rect 20955 1505 20995 1520
rect 20955 1485 20965 1505
rect 20985 1485 20995 1505
rect 20955 1455 20995 1485
rect 20955 1435 20965 1455
rect 20985 1435 20995 1455
rect 20955 1405 20995 1435
rect 20955 1385 20965 1405
rect 20985 1385 20995 1405
rect 20955 1370 20995 1385
rect 12885 1255 12925 1270
rect 12885 1235 12895 1255
rect 12915 1235 12925 1255
rect 12885 1210 12925 1235
rect 12885 1190 12895 1210
rect 12915 1190 12925 1210
rect 11165 1160 11205 1175
rect 11165 1140 11175 1160
rect 11195 1140 11205 1160
rect 11165 1110 11205 1140
rect 11165 1090 11175 1110
rect 11195 1090 11205 1110
rect 5065 1060 5105 1075
rect 5065 1040 5075 1060
rect 5095 1040 5105 1060
rect 5065 1010 5105 1040
rect 5065 990 5075 1010
rect 5095 990 5105 1010
rect 5065 975 5105 990
rect 11165 1060 11205 1090
rect 11165 1040 11175 1060
rect 11195 1040 11205 1060
rect 11165 1010 11205 1040
rect 11165 990 11175 1010
rect 11195 990 11205 1010
rect 11165 960 11205 990
rect 11165 940 11175 960
rect 11195 940 11205 960
rect 11165 925 11205 940
rect 12620 1160 12660 1175
rect 12620 1140 12630 1160
rect 12650 1140 12660 1160
rect 12620 1110 12660 1140
rect 12620 1090 12630 1110
rect 12650 1090 12660 1110
rect 12620 1060 12660 1090
rect 12620 1040 12630 1060
rect 12650 1040 12660 1060
rect 12620 1010 12660 1040
rect 12620 990 12630 1010
rect 12650 990 12660 1010
rect 12885 1165 12925 1190
rect 12885 1145 12895 1165
rect 12915 1145 12925 1165
rect 12885 1115 12925 1145
rect 12885 1095 12895 1115
rect 12915 1095 12925 1115
rect 12885 1070 12925 1095
rect 12885 1050 12895 1070
rect 12915 1050 12925 1070
rect 12885 1025 12925 1050
rect 12885 1005 12895 1025
rect 12915 1005 12925 1025
rect 12885 990 12925 1005
rect 14165 1255 14205 1270
rect 14165 1235 14175 1255
rect 14195 1235 14205 1255
rect 14165 1210 14205 1235
rect 14165 1190 14175 1210
rect 14195 1190 14205 1210
rect 14165 1165 14205 1190
rect 14165 1145 14175 1165
rect 14195 1145 14205 1165
rect 14165 1115 14205 1145
rect 14165 1095 14175 1115
rect 14195 1095 14205 1115
rect 14165 1070 14205 1095
rect 14165 1050 14175 1070
rect 14195 1050 14205 1070
rect 14165 1025 14205 1050
rect 14165 1005 14175 1025
rect 14195 1005 14205 1025
rect 14165 990 14205 1005
rect 18665 1210 18705 1225
rect 18665 1190 18675 1210
rect 18695 1190 18705 1210
rect 18665 1160 18705 1190
rect 18665 1140 18675 1160
rect 18695 1140 18705 1160
rect 18665 1110 18705 1140
rect 18665 1090 18675 1110
rect 18695 1090 18705 1110
rect 18665 1060 18705 1090
rect 18665 1040 18675 1060
rect 18695 1040 18705 1060
rect 18665 1010 18705 1040
rect 18665 990 18675 1010
rect 18695 990 18705 1010
rect 12620 960 12660 990
rect 12620 940 12630 960
rect 12650 940 12660 960
rect 12620 925 12660 940
rect 18665 975 18705 990
rect 20120 1210 20160 1225
rect 20120 1190 20130 1210
rect 20150 1190 20160 1210
rect 20120 1160 20160 1190
rect 20120 1140 20130 1160
rect 20150 1140 20160 1160
rect 20120 1110 20160 1140
rect 20120 1090 20130 1110
rect 20150 1090 20160 1110
rect 20120 1060 20160 1090
rect 20120 1040 20130 1060
rect 20150 1040 20160 1060
rect 20120 1010 20160 1040
rect 20505 1165 20545 1180
rect 20505 1145 20515 1165
rect 20535 1145 20545 1165
rect 20505 1115 20545 1145
rect 20505 1095 20515 1115
rect 20535 1095 20545 1115
rect 20505 1065 20545 1095
rect 20505 1045 20515 1065
rect 20535 1045 20545 1065
rect 20505 1030 20545 1045
rect 20805 1165 20845 1180
rect 20805 1145 20815 1165
rect 20835 1145 20845 1165
rect 20805 1115 20845 1145
rect 20805 1095 20815 1115
rect 20835 1095 20845 1115
rect 20805 1065 20845 1095
rect 20805 1045 20815 1065
rect 20835 1045 20845 1065
rect 20805 1030 20845 1045
rect 20120 990 20130 1010
rect 20150 990 20160 1010
rect 20120 975 20160 990
rect 2955 865 2995 880
rect 2955 845 2965 865
rect 2985 845 2995 865
rect 2955 815 2995 845
rect 2955 795 2965 815
rect 2985 795 2995 815
rect 2955 780 2995 795
rect 5015 865 5055 880
rect 5015 845 5025 865
rect 5045 845 5055 865
rect 5015 815 5055 845
rect 5015 795 5025 815
rect 5045 795 5055 815
rect 5015 780 5055 795
rect 9235 -745 9275 -730
rect 9235 -765 9245 -745
rect 9265 -765 9275 -745
rect 9235 -790 9275 -765
rect 9235 -810 9245 -790
rect 9265 -810 9275 -790
rect 9235 -835 9275 -810
rect 9235 -855 9245 -835
rect 9265 -855 9275 -835
rect 9235 -885 9275 -855
rect 9235 -905 9245 -885
rect 9265 -905 9275 -885
rect 9235 -930 9275 -905
rect 9235 -950 9245 -930
rect 9265 -950 9275 -930
rect 9235 -975 9275 -950
rect 9235 -995 9245 -975
rect 9265 -995 9275 -975
rect 9235 -1010 9275 -995
rect 10515 -745 10555 -730
rect 10515 -765 10525 -745
rect 10545 -765 10555 -745
rect 10515 -790 10555 -765
rect 10515 -810 10525 -790
rect 10545 -810 10555 -790
rect 10515 -835 10555 -810
rect 10515 -855 10525 -835
rect 10545 -855 10555 -835
rect 10515 -885 10555 -855
rect 10515 -905 10525 -885
rect 10545 -905 10555 -885
rect 10515 -930 10555 -905
rect 10515 -950 10525 -930
rect 10545 -950 10555 -930
rect 10515 -975 10555 -950
rect 10515 -995 10525 -975
rect 10545 -995 10555 -975
rect 10515 -1010 10555 -995
<< nsubdiff >>
rect 2955 2915 2995 2930
rect 2955 2895 2965 2915
rect 2985 2895 2995 2915
rect 2955 2865 2995 2895
rect 2955 2845 2965 2865
rect 2985 2845 2995 2865
rect 2955 2830 2995 2845
rect 5015 2915 5055 2930
rect 5015 2895 5025 2915
rect 5045 2895 5055 2915
rect 5015 2865 5055 2895
rect 5015 2845 5025 2865
rect 5045 2845 5055 2865
rect 5015 2830 5055 2845
rect 3135 2685 3175 2700
rect 3135 2665 3145 2685
rect 3165 2665 3175 2685
rect 3135 2635 3175 2665
rect 3135 2615 3145 2635
rect 3165 2615 3175 2635
rect 3135 2585 3175 2615
rect 3135 2565 3145 2585
rect 3165 2565 3175 2585
rect 3135 2535 3175 2565
rect 3135 2515 3145 2535
rect 3165 2515 3175 2535
rect 3135 2485 3175 2515
rect 3135 2465 3145 2485
rect 3165 2465 3175 2485
rect 3135 2435 3175 2465
rect 3135 2415 3145 2435
rect 3165 2415 3175 2435
rect 3135 2400 3175 2415
rect 4835 2685 4875 2700
rect 4835 2665 4845 2685
rect 4865 2665 4875 2685
rect 4835 2635 4875 2665
rect 4835 2615 4845 2635
rect 4865 2615 4875 2635
rect 4835 2585 4875 2615
rect 4835 2565 4845 2585
rect 4865 2565 4875 2585
rect 4835 2535 4875 2565
rect 4835 2515 4845 2535
rect 4865 2515 4875 2535
rect 4835 2485 4875 2515
rect 4835 2465 4845 2485
rect 4865 2465 4875 2485
rect 4835 2435 4875 2465
rect 4835 2415 4845 2435
rect 4865 2415 4875 2435
rect 4835 2400 4875 2415
rect 3985 1985 4025 2000
rect 3985 1965 3995 1985
rect 4015 1965 4025 1985
rect 3985 1935 4025 1965
rect 3985 1915 3995 1935
rect 4015 1915 4025 1935
rect 3985 1900 4025 1915
<< psubdiffcont >>
rect 10790 3495 10810 3515
rect 10790 3445 10810 3465
rect 10790 3395 10810 3415
rect 10790 3345 10810 3365
rect 10790 3295 10810 3315
rect 10460 3245 10480 3265
rect 10720 3245 10740 3265
rect 10790 3245 10810 3265
rect 11110 3545 11130 3565
rect 11110 3495 11130 3515
rect 11110 3445 11130 3465
rect 11110 3395 11130 3415
rect 11110 3345 11130 3365
rect 11110 3295 11130 3315
rect 11110 3245 11130 3265
rect 11190 3540 11210 3560
rect 11190 3490 11210 3510
rect 11190 3440 11210 3460
rect 11190 3390 11210 3410
rect 11190 3340 11210 3360
rect 11190 3290 11210 3310
rect 11190 3240 11210 3260
rect 11190 3190 11210 3210
rect 12590 3540 12610 3560
rect 12590 3490 12610 3510
rect 12590 3440 12610 3460
rect 12590 3390 12610 3410
rect 12590 3340 12610 3360
rect 18290 3495 18310 3515
rect 18290 3445 18310 3465
rect 18290 3395 18310 3415
rect 12590 3290 12610 3310
rect 18290 3345 18310 3365
rect 18290 3295 18310 3315
rect 12590 3240 12610 3260
rect 17960 3245 17980 3265
rect 12590 3190 12610 3210
rect 12860 3205 12880 3225
rect 12860 3155 12880 3175
rect 12860 3105 12880 3125
rect 12860 3055 12880 3075
rect 12860 3005 12880 3025
rect 12860 2955 12880 2975
rect 920 2880 950 2910
rect 1000 2880 1030 2910
rect 1080 2880 1110 2910
rect 18220 3245 18240 3265
rect 18290 3245 18310 3265
rect 18610 3545 18630 3565
rect 18610 3495 18630 3515
rect 18610 3445 18630 3465
rect 18610 3395 18630 3415
rect 18610 3345 18630 3365
rect 18610 3295 18630 3315
rect 18610 3245 18630 3265
rect 18690 3540 18710 3560
rect 18690 3490 18710 3510
rect 18690 3440 18710 3460
rect 18690 3390 18710 3410
rect 18690 3340 18710 3360
rect 18690 3290 18710 3310
rect 18690 3240 18710 3260
rect 14150 3205 14170 3225
rect 18690 3190 18710 3210
rect 20090 3540 20110 3560
rect 20090 3490 20110 3510
rect 20090 3440 20110 3460
rect 20090 3390 20110 3410
rect 20090 3340 20110 3360
rect 20090 3290 20110 3310
rect 20090 3240 20110 3260
rect 20090 3190 20110 3210
rect 20360 3205 20380 3225
rect 14150 3155 14170 3175
rect 20360 3155 20380 3175
rect 14150 3105 14170 3125
rect 14150 3055 14170 3075
rect 14150 3005 14170 3025
rect 14150 2955 14170 2975
rect 20360 3105 20380 3125
rect 20360 3055 20380 3075
rect 20360 3005 20380 3025
rect 20360 2955 20380 2975
rect 11190 2860 11210 2880
rect 11190 2810 11210 2830
rect 11190 2760 11210 2780
rect 11190 2710 11210 2730
rect 11190 2660 11210 2680
rect 9650 2585 9670 2605
rect 9650 2535 9670 2555
rect 10940 2585 10960 2605
rect 10940 2535 10960 2555
rect 11190 2610 11210 2630
rect 11190 2560 11210 2580
rect 11190 2510 11210 2530
rect 21650 3205 21670 3225
rect 21650 3155 21670 3175
rect 21650 3105 21670 3125
rect 21650 3055 21670 3075
rect 21650 3005 21670 3025
rect 21650 2955 21670 2975
rect 12590 2860 12610 2880
rect 18690 2860 18710 2880
rect 12590 2810 12610 2830
rect 12590 2760 12610 2780
rect 12590 2710 12610 2730
rect 18690 2810 18710 2830
rect 18690 2760 18710 2780
rect 18690 2710 18710 2730
rect 12590 2660 12610 2680
rect 18690 2660 18710 2680
rect 12590 2610 12610 2630
rect 12590 2560 12610 2580
rect 12590 2510 12610 2530
rect 12860 2585 12880 2605
rect 12860 2535 12880 2555
rect 14150 2585 14170 2605
rect 14150 2535 14170 2555
rect 17150 2585 17170 2605
rect 17150 2535 17170 2555
rect 18440 2585 18460 2605
rect 18440 2535 18460 2555
rect 18690 2610 18710 2630
rect 18690 2560 18710 2580
rect 18690 2510 18710 2530
rect 20090 2860 20110 2880
rect 20090 2810 20110 2830
rect 20090 2760 20110 2780
rect 20090 2710 20110 2730
rect 20090 2660 20110 2680
rect 20090 2610 20110 2630
rect 20090 2560 20110 2580
rect 20090 2510 20110 2530
rect 20360 2585 20380 2605
rect 20360 2535 20380 2555
rect 21650 2585 21670 2605
rect 21650 2535 21670 2555
rect 9650 2135 9670 2155
rect 9650 2085 9670 2105
rect 9650 2035 9670 2055
rect 10940 2135 10960 2155
rect 12860 2135 12880 2155
rect 10940 2085 10960 2105
rect 10940 2035 10960 2055
rect 11245 2095 11265 2115
rect 11245 2045 11265 2065
rect 11245 1995 11265 2015
rect 12535 2095 12555 2115
rect 12535 2045 12555 2065
rect 12860 2085 12880 2105
rect 12860 2035 12880 2055
rect 14150 2135 14170 2155
rect 14150 2085 14170 2105
rect 14150 2035 14170 2055
rect 17150 2135 17170 2155
rect 17150 2085 17170 2105
rect 17150 2035 17170 2055
rect 18440 2135 18460 2155
rect 20360 2135 20380 2155
rect 18440 2085 18460 2105
rect 18440 2035 18460 2055
rect 18745 2095 18765 2115
rect 18745 2045 18765 2065
rect 12535 1995 12555 2015
rect 18745 1995 18765 2015
rect 20035 2095 20055 2115
rect 20035 2045 20055 2065
rect 20360 2085 20380 2105
rect 20360 2035 20380 2055
rect 21650 2135 21670 2155
rect 21650 2085 21670 2105
rect 21650 2035 21670 2055
rect 20035 1995 20055 2015
rect 20460 1820 20480 1840
rect 20460 1770 20480 1790
rect -35 1695 -15 1715
rect 15 1695 35 1715
rect 65 1695 85 1715
rect 20460 1720 20480 1740
rect 20870 1820 20890 1840
rect 20870 1770 20890 1790
rect 20870 1720 20890 1740
rect 3995 1630 4015 1650
rect 11000 1630 11020 1650
rect 11000 1580 11020 1600
rect 11000 1530 11020 1550
rect 11740 1630 11760 1650
rect 11740 1580 11760 1600
rect 11740 1530 11760 1550
rect 12040 1630 12060 1650
rect 12040 1580 12060 1600
rect 12040 1530 12060 1550
rect 12780 1630 12800 1650
rect 12780 1580 12800 1600
rect 12780 1530 12800 1550
rect 18500 1630 18520 1650
rect 18500 1580 18520 1600
rect 18500 1530 18520 1550
rect 19240 1630 19260 1650
rect 19240 1580 19260 1600
rect 19240 1530 19260 1550
rect 19540 1630 19560 1650
rect 19540 1580 19560 1600
rect 19540 1530 19560 1550
rect 20280 1630 20300 1650
rect 20280 1580 20300 1600
rect 20280 1530 20300 1550
rect 20365 1485 20385 1505
rect 20365 1435 20385 1455
rect 20365 1385 20385 1405
rect 20665 1485 20685 1505
rect 20665 1435 20685 1455
rect 20665 1385 20685 1405
rect 20965 1485 20985 1505
rect 20965 1435 20985 1455
rect 20965 1385 20985 1405
rect 12895 1235 12915 1255
rect 12895 1190 12915 1210
rect 11175 1140 11195 1160
rect 11175 1090 11195 1110
rect 5075 1040 5095 1060
rect 5075 990 5095 1010
rect 11175 1040 11195 1060
rect 11175 990 11195 1010
rect 11175 940 11195 960
rect 12630 1140 12650 1160
rect 12630 1090 12650 1110
rect 12630 1040 12650 1060
rect 12630 990 12650 1010
rect 12895 1145 12915 1165
rect 12895 1095 12915 1115
rect 12895 1050 12915 1070
rect 12895 1005 12915 1025
rect 14175 1235 14195 1255
rect 14175 1190 14195 1210
rect 14175 1145 14195 1165
rect 14175 1095 14195 1115
rect 14175 1050 14195 1070
rect 14175 1005 14195 1025
rect 18675 1190 18695 1210
rect 18675 1140 18695 1160
rect 18675 1090 18695 1110
rect 18675 1040 18695 1060
rect 18675 990 18695 1010
rect 12630 940 12650 960
rect 20130 1190 20150 1210
rect 20130 1140 20150 1160
rect 20130 1090 20150 1110
rect 20130 1040 20150 1060
rect 20515 1145 20535 1165
rect 20515 1095 20535 1115
rect 20515 1045 20535 1065
rect 20815 1145 20835 1165
rect 20815 1095 20835 1115
rect 20815 1045 20835 1065
rect 20130 990 20150 1010
rect 2965 845 2985 865
rect 2965 795 2985 815
rect 5025 845 5045 865
rect 5025 795 5045 815
rect 9245 -765 9265 -745
rect 9245 -810 9265 -790
rect 9245 -855 9265 -835
rect 9245 -905 9265 -885
rect 9245 -950 9265 -930
rect 9245 -995 9265 -975
rect 10525 -765 10545 -745
rect 10525 -810 10545 -790
rect 10525 -855 10545 -835
rect 10525 -905 10545 -885
rect 10525 -950 10545 -930
rect 10525 -995 10545 -975
<< nsubdiffcont >>
rect 2965 2895 2985 2915
rect 2965 2845 2985 2865
rect 5025 2895 5045 2915
rect 5025 2845 5045 2865
rect 3145 2665 3165 2685
rect 3145 2615 3165 2635
rect 3145 2565 3165 2585
rect 3145 2515 3165 2535
rect 3145 2465 3165 2485
rect 3145 2415 3165 2435
rect 4845 2665 4865 2685
rect 4845 2615 4865 2635
rect 4845 2565 4865 2585
rect 4845 2515 4865 2535
rect 4845 2465 4865 2485
rect 4845 2415 4865 2435
rect 3995 1965 4015 1985
rect 3995 1915 4015 1935
<< poly >>
rect 11180 3620 11220 3630
rect 10905 3605 10945 3615
rect 10905 3585 10915 3605
rect 10935 3585 10945 3605
rect 11180 3600 11190 3620
rect 11210 3600 11220 3620
rect 12580 3620 12620 3630
rect 12580 3600 12590 3620
rect 12610 3600 12620 3620
rect 18680 3620 18720 3630
rect 10905 3575 10945 3585
rect 10980 3580 11000 3595
rect 11040 3580 11060 3595
rect 11180 3585 11280 3600
rect 10860 3550 10880 3565
rect 10920 3550 10940 3575
rect 10450 3340 10490 3350
rect 10450 3320 10460 3340
rect 10480 3320 10490 3340
rect 10710 3340 10750 3350
rect 10710 3320 10720 3340
rect 10740 3320 10750 3340
rect 10450 3305 10550 3320
rect 10530 3293 10550 3305
rect 10590 3293 10610 3308
rect 10650 3305 10750 3320
rect 10650 3293 10670 3305
rect 11260 3575 11280 3585
rect 11320 3575 11340 3590
rect 11380 3575 11400 3590
rect 11440 3575 11460 3590
rect 11500 3575 11520 3590
rect 11560 3575 11580 3590
rect 11620 3575 11640 3590
rect 11680 3575 11700 3590
rect 11740 3575 11760 3590
rect 11800 3575 11820 3590
rect 11860 3575 11880 3590
rect 11920 3575 11940 3590
rect 11980 3575 12000 3590
rect 12040 3575 12060 3590
rect 12100 3575 12120 3590
rect 12160 3575 12180 3590
rect 12220 3575 12240 3590
rect 12280 3575 12300 3590
rect 12340 3575 12360 3590
rect 12400 3575 12420 3590
rect 12460 3575 12480 3590
rect 12520 3585 12620 3600
rect 18405 3605 18445 3615
rect 18405 3585 18415 3605
rect 18435 3585 18445 3605
rect 18680 3600 18690 3620
rect 18710 3600 18720 3620
rect 20080 3620 20120 3630
rect 20080 3600 20090 3620
rect 20110 3600 20120 3620
rect 12520 3575 12540 3585
rect 18405 3575 18445 3585
rect 18480 3580 18500 3595
rect 18540 3580 18560 3595
rect 18680 3585 18780 3600
rect 10530 3215 10550 3230
rect 10590 3215 10610 3230
rect 10650 3215 10670 3230
rect 10860 3220 10880 3230
rect 10580 3205 10620 3215
rect 10580 3185 10590 3205
rect 10610 3185 10620 3205
rect 10580 3175 10620 3185
rect 10780 3205 10880 3220
rect 10920 3215 10940 3230
rect 10905 3205 10940 3215
rect 10780 3185 10790 3205
rect 10810 3185 10820 3205
rect 10780 3175 10820 3185
rect 10905 3185 10910 3205
rect 10930 3185 10940 3205
rect 10905 3175 10940 3185
rect 10980 3215 11000 3230
rect 11040 3220 11060 3230
rect 10980 3205 11015 3215
rect 11040 3205 11140 3220
rect 10980 3185 10990 3205
rect 11010 3185 11015 3205
rect 10980 3175 11015 3185
rect 11100 3185 11110 3205
rect 11130 3185 11140 3205
rect 11100 3175 11140 3185
rect 18360 3550 18380 3565
rect 18420 3550 18440 3575
rect 17950 3340 17990 3350
rect 17950 3320 17960 3340
rect 17980 3320 17990 3340
rect 18210 3340 18250 3350
rect 18210 3320 18220 3340
rect 18240 3320 18250 3340
rect 17950 3305 18050 3320
rect 18030 3293 18050 3305
rect 18090 3293 18110 3308
rect 18150 3305 18250 3320
rect 18150 3293 18170 3305
rect 12930 3240 12945 3255
rect 12985 3240 13000 3255
rect 13040 3240 13055 3255
rect 13095 3240 13110 3255
rect 13150 3240 13165 3255
rect 13205 3240 13220 3255
rect 13260 3240 13275 3255
rect 13315 3240 13330 3255
rect 13370 3240 13385 3255
rect 13425 3240 13440 3255
rect 13480 3240 13495 3255
rect 13535 3240 13550 3255
rect 13590 3240 13605 3255
rect 13645 3240 13660 3255
rect 13700 3240 13715 3255
rect 13755 3240 13770 3255
rect 13810 3240 13825 3255
rect 13865 3240 13880 3255
rect 13920 3240 13935 3255
rect 13975 3240 13990 3255
rect 14030 3240 14045 3255
rect 14085 3240 14100 3255
rect 11260 3160 11280 3175
rect 11320 3165 11340 3175
rect 11380 3165 11400 3175
rect 11440 3165 11460 3175
rect 11500 3165 11520 3175
rect 11560 3165 11580 3175
rect 11620 3165 11640 3175
rect 11680 3165 11700 3175
rect 11740 3165 11760 3175
rect 11800 3165 11820 3175
rect 11860 3165 11880 3175
rect 11920 3165 11940 3175
rect 11980 3165 12000 3175
rect 12040 3165 12060 3175
rect 12100 3165 12120 3175
rect 12160 3165 12180 3175
rect 12220 3165 12240 3175
rect 12280 3165 12300 3175
rect 12340 3165 12360 3175
rect 12400 3165 12420 3175
rect 12460 3165 12480 3175
rect 11320 3150 12480 3165
rect 12520 3160 12540 3175
rect 11823 3130 11831 3150
rect 11849 3130 11857 3150
rect 11823 3120 11857 3130
rect 3140 2975 3175 2985
rect 3140 2955 3145 2975
rect 3165 2955 3175 2975
rect 3140 2945 3175 2955
rect 4835 2975 4870 2985
rect 4835 2955 4845 2975
rect 4865 2955 4870 2975
rect 4835 2945 4870 2955
rect 3035 2930 3085 2945
rect 3125 2930 3175 2945
rect 3215 2930 3265 2945
rect 3305 2930 3355 2945
rect 3395 2930 3445 2945
rect 3485 2930 3535 2945
rect 3575 2930 3625 2945
rect 3665 2930 3715 2945
rect 3755 2930 3805 2945
rect 3845 2930 3895 2945
rect 3935 2930 3985 2945
rect 4025 2930 4075 2945
rect 4115 2930 4165 2945
rect 4205 2930 4255 2945
rect 4295 2930 4345 2945
rect 4385 2930 4435 2945
rect 4475 2930 4525 2945
rect 4565 2930 4615 2945
rect 4655 2930 4705 2945
rect 4745 2930 4795 2945
rect 4835 2930 4885 2945
rect 4925 2930 4975 2945
rect 11180 2940 11220 2950
rect 11180 2920 11190 2940
rect 11210 2920 11220 2940
rect 12580 2940 12620 2950
rect 18760 3575 18780 3585
rect 18820 3575 18840 3590
rect 18880 3575 18900 3590
rect 18940 3575 18960 3590
rect 19000 3575 19020 3590
rect 19060 3575 19080 3590
rect 19120 3575 19140 3590
rect 19180 3575 19200 3590
rect 19240 3575 19260 3590
rect 19300 3575 19320 3590
rect 19360 3575 19380 3590
rect 19420 3575 19440 3590
rect 19480 3575 19500 3590
rect 19540 3575 19560 3590
rect 19600 3575 19620 3590
rect 19660 3575 19680 3590
rect 19720 3575 19740 3590
rect 19780 3575 19800 3590
rect 19840 3575 19860 3590
rect 19900 3575 19920 3590
rect 19960 3575 19980 3590
rect 20020 3585 20120 3600
rect 20020 3575 20040 3585
rect 18030 3215 18050 3230
rect 18090 3215 18110 3230
rect 18150 3215 18170 3230
rect 18360 3220 18380 3230
rect 18080 3205 18120 3215
rect 18080 3185 18090 3205
rect 18110 3185 18120 3205
rect 18080 3175 18120 3185
rect 18280 3205 18380 3220
rect 18420 3215 18440 3230
rect 18405 3205 18440 3215
rect 18280 3185 18290 3205
rect 18310 3185 18320 3205
rect 18280 3175 18320 3185
rect 18405 3185 18410 3205
rect 18430 3185 18440 3205
rect 18405 3175 18440 3185
rect 18480 3215 18500 3230
rect 18540 3220 18560 3230
rect 18480 3205 18515 3215
rect 18540 3205 18640 3220
rect 18480 3185 18490 3205
rect 18510 3185 18515 3205
rect 18480 3175 18515 3185
rect 18600 3185 18610 3205
rect 18630 3185 18640 3205
rect 18600 3175 18640 3185
rect 20430 3240 20445 3255
rect 20485 3240 20500 3255
rect 20540 3240 20555 3255
rect 20595 3240 20610 3255
rect 20650 3240 20665 3255
rect 20705 3240 20720 3255
rect 20760 3240 20775 3255
rect 20815 3240 20830 3255
rect 20870 3240 20885 3255
rect 20925 3240 20940 3255
rect 20980 3240 20995 3255
rect 21035 3240 21050 3255
rect 21090 3240 21105 3255
rect 21145 3240 21160 3255
rect 21200 3240 21215 3255
rect 21255 3240 21270 3255
rect 21310 3240 21325 3255
rect 21365 3240 21380 3255
rect 21420 3240 21435 3255
rect 21475 3240 21490 3255
rect 21530 3240 21545 3255
rect 21585 3240 21600 3255
rect 18760 3160 18780 3175
rect 18820 3165 18840 3175
rect 18880 3165 18900 3175
rect 18940 3165 18960 3175
rect 19000 3165 19020 3175
rect 19060 3165 19080 3175
rect 19120 3165 19140 3175
rect 19180 3165 19200 3175
rect 19240 3165 19260 3175
rect 19300 3165 19320 3175
rect 19360 3165 19380 3175
rect 19420 3165 19440 3175
rect 19480 3165 19500 3175
rect 19540 3165 19560 3175
rect 19600 3165 19620 3175
rect 19660 3165 19680 3175
rect 19720 3165 19740 3175
rect 19780 3165 19800 3175
rect 19840 3165 19860 3175
rect 19900 3165 19920 3175
rect 19960 3165 19980 3175
rect 18820 3150 19980 3165
rect 20020 3160 20040 3175
rect 19323 3130 19331 3150
rect 19349 3130 19357 3150
rect 19323 3120 19357 3130
rect 18680 2940 18720 2950
rect 12580 2920 12590 2940
rect 12610 2920 12620 2940
rect 12930 2930 12945 2940
rect 11180 2905 11280 2920
rect 11260 2895 11280 2905
rect 11320 2895 11340 2910
rect 11380 2895 11400 2910
rect 11440 2895 11460 2910
rect 11500 2895 11520 2910
rect 11560 2895 11580 2910
rect 11620 2895 11640 2910
rect 11680 2895 11700 2910
rect 11740 2895 11760 2910
rect 11800 2895 11820 2910
rect 11860 2895 11880 2910
rect 11920 2895 11940 2910
rect 11980 2895 12000 2910
rect 12040 2895 12060 2910
rect 12100 2895 12120 2910
rect 12160 2895 12180 2910
rect 12220 2895 12240 2910
rect 12280 2895 12300 2910
rect 12340 2895 12360 2910
rect 12400 2895 12420 2910
rect 12460 2895 12480 2910
rect 12520 2905 12620 2920
rect 12850 2915 12945 2930
rect 12985 2930 13000 2940
rect 13040 2930 13055 2940
rect 13095 2930 13110 2940
rect 13150 2930 13165 2940
rect 13205 2930 13220 2940
rect 13260 2930 13275 2940
rect 13315 2930 13330 2940
rect 13370 2930 13385 2940
rect 13425 2930 13440 2940
rect 13480 2930 13495 2940
rect 13535 2930 13550 2940
rect 13590 2930 13605 2940
rect 13645 2930 13660 2940
rect 13700 2930 13715 2940
rect 13755 2930 13770 2940
rect 13810 2930 13825 2940
rect 13865 2930 13880 2940
rect 13920 2930 13935 2940
rect 13975 2930 13990 2940
rect 14030 2930 14045 2940
rect 12985 2915 14045 2930
rect 14085 2930 14100 2940
rect 14085 2915 14180 2930
rect 12520 2895 12540 2905
rect 12850 2895 12860 2915
rect 12880 2895 12890 2915
rect 3035 2815 3085 2830
rect 2995 2805 3085 2815
rect 3125 2820 3175 2830
rect 3215 2820 3265 2830
rect 3305 2820 3355 2830
rect 3395 2820 3445 2830
rect 3485 2820 3535 2830
rect 3575 2820 3625 2830
rect 3665 2820 3715 2830
rect 3755 2820 3805 2830
rect 3845 2820 3895 2830
rect 3935 2820 3985 2830
rect 4025 2820 4075 2830
rect 4115 2820 4165 2830
rect 4205 2820 4255 2830
rect 4295 2820 4345 2830
rect 4385 2820 4435 2830
rect 4475 2820 4525 2830
rect 4565 2820 4615 2830
rect 4655 2820 4705 2830
rect 4745 2820 4795 2830
rect 4835 2820 4885 2830
rect 3125 2805 4885 2820
rect 4925 2815 4975 2830
rect 4925 2805 5015 2815
rect 2995 2785 3005 2805
rect 3025 2800 3085 2805
rect 4925 2800 4985 2805
rect 3025 2785 3035 2800
rect 2995 2775 3035 2785
rect 4975 2785 4985 2800
rect 5005 2785 5015 2805
rect 4975 2775 5015 2785
rect 3175 2745 3215 2755
rect 3175 2725 3185 2745
rect 3205 2730 3215 2745
rect 4795 2745 4835 2755
rect 4795 2730 4805 2745
rect 3205 2725 3265 2730
rect 3175 2715 3265 2725
rect 4745 2725 4805 2730
rect 4825 2725 4835 2745
rect 4745 2715 4835 2725
rect 3215 2700 3265 2715
rect 3305 2700 3355 2715
rect 3395 2700 3445 2715
rect 3485 2700 3535 2715
rect 3575 2700 3625 2715
rect 3665 2700 3715 2715
rect 3755 2700 3805 2715
rect 3845 2700 3895 2715
rect 3935 2700 3985 2715
rect 4025 2700 4075 2715
rect 4115 2700 4165 2715
rect 4205 2700 4255 2715
rect 4295 2700 4345 2715
rect 4385 2700 4435 2715
rect 4475 2700 4525 2715
rect 4565 2700 4615 2715
rect 4655 2700 4705 2715
rect 4745 2700 4795 2715
rect 9720 2620 9735 2635
rect 9775 2620 9790 2635
rect 9830 2620 9845 2635
rect 9885 2620 9900 2635
rect 9940 2620 9955 2635
rect 9995 2620 10010 2635
rect 10050 2620 10065 2635
rect 10105 2620 10120 2635
rect 10160 2620 10175 2635
rect 10215 2620 10230 2635
rect 10270 2620 10285 2635
rect 10325 2620 10340 2635
rect 10380 2620 10395 2635
rect 10435 2620 10450 2635
rect 10490 2620 10505 2635
rect 10545 2620 10560 2635
rect 10600 2620 10615 2635
rect 10655 2620 10670 2635
rect 10710 2620 10725 2635
rect 10765 2620 10780 2635
rect 10820 2620 10835 2635
rect 10875 2620 10890 2635
rect 9720 2510 9735 2520
rect 9640 2495 9735 2510
rect 9775 2510 9790 2520
rect 9830 2510 9845 2520
rect 9885 2510 9900 2520
rect 9940 2510 9955 2520
rect 9995 2510 10010 2520
rect 10050 2510 10065 2520
rect 10105 2510 10120 2520
rect 10160 2510 10175 2520
rect 10215 2510 10230 2520
rect 10270 2510 10285 2520
rect 10325 2510 10340 2520
rect 10380 2510 10395 2520
rect 10435 2510 10450 2520
rect 10490 2510 10505 2520
rect 10545 2510 10560 2520
rect 10600 2510 10615 2520
rect 10655 2510 10670 2520
rect 10710 2510 10725 2520
rect 10765 2510 10780 2520
rect 10820 2510 10835 2520
rect 9775 2495 10835 2510
rect 10875 2510 10890 2520
rect 10875 2495 10970 2510
rect 12850 2885 12890 2895
rect 13058 2895 13066 2915
rect 13084 2895 13092 2915
rect 13058 2885 13092 2895
rect 14140 2895 14150 2915
rect 14170 2895 14180 2915
rect 18680 2920 18690 2940
rect 18710 2920 18720 2940
rect 20080 2940 20120 2950
rect 20080 2920 20090 2940
rect 20110 2920 20120 2940
rect 20430 2930 20445 2940
rect 18680 2905 18780 2920
rect 18760 2895 18780 2905
rect 18820 2895 18840 2910
rect 18880 2895 18900 2910
rect 18940 2895 18960 2910
rect 19000 2895 19020 2910
rect 19060 2895 19080 2910
rect 19120 2895 19140 2910
rect 19180 2895 19200 2910
rect 19240 2895 19260 2910
rect 19300 2895 19320 2910
rect 19360 2895 19380 2910
rect 19420 2895 19440 2910
rect 19480 2895 19500 2910
rect 19540 2895 19560 2910
rect 19600 2895 19620 2910
rect 19660 2895 19680 2910
rect 19720 2895 19740 2910
rect 19780 2895 19800 2910
rect 19840 2895 19860 2910
rect 19900 2895 19920 2910
rect 19960 2895 19980 2910
rect 20020 2905 20120 2920
rect 20350 2915 20445 2930
rect 20485 2930 20500 2940
rect 20540 2930 20555 2940
rect 20595 2930 20610 2940
rect 20650 2930 20665 2940
rect 20705 2930 20720 2940
rect 20760 2930 20775 2940
rect 20815 2930 20830 2940
rect 20870 2930 20885 2940
rect 20925 2930 20940 2940
rect 20980 2930 20995 2940
rect 21035 2930 21050 2940
rect 21090 2930 21105 2940
rect 21145 2930 21160 2940
rect 21200 2930 21215 2940
rect 21255 2930 21270 2940
rect 21310 2930 21325 2940
rect 21365 2930 21380 2940
rect 21420 2930 21435 2940
rect 21475 2930 21490 2940
rect 21530 2930 21545 2940
rect 20485 2915 21545 2930
rect 21585 2930 21600 2940
rect 21585 2915 21680 2930
rect 20020 2895 20040 2905
rect 20350 2895 20360 2915
rect 20380 2895 20390 2915
rect 14140 2885 14180 2895
rect 12930 2620 12945 2635
rect 12985 2620 13000 2635
rect 13040 2620 13055 2635
rect 13095 2620 13110 2635
rect 13150 2620 13165 2635
rect 13205 2620 13220 2635
rect 13260 2620 13275 2635
rect 13315 2620 13330 2635
rect 13370 2620 13385 2635
rect 13425 2620 13440 2635
rect 13480 2620 13495 2635
rect 13535 2620 13550 2635
rect 13590 2620 13605 2635
rect 13645 2620 13660 2635
rect 13700 2620 13715 2635
rect 13755 2620 13770 2635
rect 13810 2620 13825 2635
rect 13865 2620 13880 2635
rect 13920 2620 13935 2635
rect 13975 2620 13990 2635
rect 14030 2620 14045 2635
rect 14085 2620 14100 2635
rect 17220 2620 17235 2635
rect 17275 2620 17290 2635
rect 17330 2620 17345 2635
rect 17385 2620 17400 2635
rect 17440 2620 17455 2635
rect 17495 2620 17510 2635
rect 17550 2620 17565 2635
rect 17605 2620 17620 2635
rect 17660 2620 17675 2635
rect 17715 2620 17730 2635
rect 17770 2620 17785 2635
rect 17825 2620 17840 2635
rect 17880 2620 17895 2635
rect 17935 2620 17950 2635
rect 17990 2620 18005 2635
rect 18045 2620 18060 2635
rect 18100 2620 18115 2635
rect 18155 2620 18170 2635
rect 18210 2620 18225 2635
rect 18265 2620 18280 2635
rect 18320 2620 18335 2635
rect 18375 2620 18390 2635
rect 12930 2510 12945 2520
rect 12850 2495 12945 2510
rect 12985 2510 13000 2520
rect 13040 2510 13055 2520
rect 13095 2510 13110 2520
rect 13150 2510 13165 2520
rect 13205 2510 13220 2520
rect 13260 2510 13275 2520
rect 13315 2510 13330 2520
rect 13370 2510 13385 2520
rect 13425 2510 13440 2520
rect 13480 2510 13495 2520
rect 13535 2510 13550 2520
rect 13590 2510 13605 2520
rect 13645 2510 13660 2520
rect 13700 2510 13715 2520
rect 13755 2510 13770 2520
rect 13810 2510 13825 2520
rect 13865 2510 13880 2520
rect 13920 2510 13935 2520
rect 13975 2510 13990 2520
rect 14030 2510 14045 2520
rect 12985 2495 14045 2510
rect 14085 2510 14100 2520
rect 17220 2510 17235 2520
rect 14085 2495 14180 2510
rect 9640 2475 9650 2495
rect 9670 2475 9680 2495
rect 9640 2465 9680 2475
rect 10820 2445 10835 2495
rect 10930 2475 10940 2495
rect 10960 2475 10970 2495
rect 11260 2480 11280 2495
rect 11320 2485 11340 2495
rect 11380 2485 11400 2495
rect 11440 2485 11460 2495
rect 11500 2485 11520 2495
rect 11560 2485 11580 2495
rect 11620 2485 11640 2495
rect 11680 2485 11700 2495
rect 11740 2485 11760 2495
rect 11800 2485 11820 2495
rect 11860 2485 11880 2495
rect 11920 2485 11940 2495
rect 11980 2485 12000 2495
rect 12040 2485 12060 2495
rect 12100 2485 12120 2495
rect 12160 2485 12180 2495
rect 12220 2485 12240 2495
rect 12280 2485 12300 2495
rect 12340 2485 12360 2495
rect 12400 2485 12420 2495
rect 12460 2485 12480 2495
rect 10930 2465 10970 2475
rect 11320 2470 12480 2485
rect 12520 2480 12540 2495
rect 12850 2475 12860 2495
rect 12880 2475 12890 2495
rect 11823 2450 11831 2470
rect 11849 2450 11857 2470
rect 12850 2465 12890 2475
rect 10813 2435 10847 2445
rect 11823 2440 11857 2450
rect 12985 2445 13000 2495
rect 14140 2475 14150 2495
rect 14170 2475 14180 2495
rect 14140 2465 14180 2475
rect 17140 2495 17235 2510
rect 17275 2510 17290 2520
rect 17330 2510 17345 2520
rect 17385 2510 17400 2520
rect 17440 2510 17455 2520
rect 17495 2510 17510 2520
rect 17550 2510 17565 2520
rect 17605 2510 17620 2520
rect 17660 2510 17675 2520
rect 17715 2510 17730 2520
rect 17770 2510 17785 2520
rect 17825 2510 17840 2520
rect 17880 2510 17895 2520
rect 17935 2510 17950 2520
rect 17990 2510 18005 2520
rect 18045 2510 18060 2520
rect 18100 2510 18115 2520
rect 18155 2510 18170 2520
rect 18210 2510 18225 2520
rect 18265 2510 18280 2520
rect 18320 2510 18335 2520
rect 17275 2495 18335 2510
rect 18375 2510 18390 2520
rect 18375 2495 18470 2510
rect 20350 2885 20390 2895
rect 20558 2895 20566 2915
rect 20584 2895 20592 2915
rect 20558 2885 20592 2895
rect 21640 2895 21650 2915
rect 21670 2895 21680 2915
rect 21640 2885 21680 2895
rect 20430 2620 20445 2635
rect 20485 2620 20500 2635
rect 20540 2620 20555 2635
rect 20595 2620 20610 2635
rect 20650 2620 20665 2635
rect 20705 2620 20720 2635
rect 20760 2620 20775 2635
rect 20815 2620 20830 2635
rect 20870 2620 20885 2635
rect 20925 2620 20940 2635
rect 20980 2620 20995 2635
rect 21035 2620 21050 2635
rect 21090 2620 21105 2635
rect 21145 2620 21160 2635
rect 21200 2620 21215 2635
rect 21255 2620 21270 2635
rect 21310 2620 21325 2635
rect 21365 2620 21380 2635
rect 21420 2620 21435 2635
rect 21475 2620 21490 2635
rect 21530 2620 21545 2635
rect 21585 2620 21600 2635
rect 20430 2510 20445 2520
rect 20350 2495 20445 2510
rect 20485 2510 20500 2520
rect 20540 2510 20555 2520
rect 20595 2510 20610 2520
rect 20650 2510 20665 2520
rect 20705 2510 20720 2520
rect 20760 2510 20775 2520
rect 20815 2510 20830 2520
rect 20870 2510 20885 2520
rect 20925 2510 20940 2520
rect 20980 2510 20995 2520
rect 21035 2510 21050 2520
rect 21090 2510 21105 2520
rect 21145 2510 21160 2520
rect 21200 2510 21215 2520
rect 21255 2510 21270 2520
rect 21310 2510 21325 2520
rect 21365 2510 21380 2520
rect 21420 2510 21435 2520
rect 21475 2510 21490 2520
rect 21530 2510 21545 2520
rect 20485 2495 21545 2510
rect 21585 2510 21600 2520
rect 21585 2495 21680 2510
rect 17140 2475 17150 2495
rect 17170 2475 17180 2495
rect 17140 2465 17180 2475
rect 18320 2445 18335 2495
rect 18430 2475 18440 2495
rect 18460 2475 18470 2495
rect 18760 2480 18780 2495
rect 18820 2485 18840 2495
rect 18880 2485 18900 2495
rect 18940 2485 18960 2495
rect 19000 2485 19020 2495
rect 19060 2485 19080 2495
rect 19120 2485 19140 2495
rect 19180 2485 19200 2495
rect 19240 2485 19260 2495
rect 19300 2485 19320 2495
rect 19360 2485 19380 2495
rect 19420 2485 19440 2495
rect 19480 2485 19500 2495
rect 19540 2485 19560 2495
rect 19600 2485 19620 2495
rect 19660 2485 19680 2495
rect 19720 2485 19740 2495
rect 19780 2485 19800 2495
rect 19840 2485 19860 2495
rect 19900 2485 19920 2495
rect 19960 2485 19980 2495
rect 18430 2465 18470 2475
rect 18820 2470 19980 2485
rect 20020 2480 20040 2495
rect 20350 2475 20360 2495
rect 20380 2475 20390 2495
rect 19323 2450 19331 2470
rect 19349 2450 19357 2470
rect 20350 2465 20390 2475
rect 10813 2415 10821 2435
rect 10839 2415 10847 2435
rect 10813 2405 10847 2415
rect 12973 2435 13007 2445
rect 12973 2415 12981 2435
rect 12999 2415 13007 2435
rect 12973 2405 13007 2415
rect 18313 2435 18347 2445
rect 19323 2440 19357 2450
rect 20485 2445 20500 2495
rect 21640 2475 21650 2495
rect 21670 2475 21680 2495
rect 21640 2465 21680 2475
rect 18313 2415 18321 2435
rect 18339 2415 18347 2435
rect 18313 2405 18347 2415
rect 20473 2435 20507 2445
rect 20473 2415 20481 2435
rect 20499 2415 20507 2435
rect 20473 2405 20507 2415
rect 3215 2385 3265 2400
rect 3305 2390 3355 2400
rect 3395 2390 3445 2400
rect 3485 2390 3535 2400
rect 3575 2390 3625 2400
rect 3665 2390 3715 2400
rect 3755 2390 3805 2400
rect 3845 2390 3895 2400
rect 3935 2390 3985 2400
rect 4025 2390 4075 2400
rect 4115 2390 4165 2400
rect 4205 2390 4255 2400
rect 4295 2390 4345 2400
rect 4385 2390 4435 2400
rect 4475 2390 4525 2400
rect 4565 2390 4615 2400
rect 4655 2390 4705 2400
rect 3305 2375 4705 2390
rect 4745 2385 4795 2400
rect 3355 2370 3395 2375
rect 3355 2350 3365 2370
rect 3385 2350 3395 2370
rect 3355 2340 3395 2350
rect 3885 2355 3895 2375
rect 3915 2355 3925 2375
rect 3885 2345 3925 2355
rect 10813 2275 10847 2285
rect 10813 2255 10821 2275
rect 10839 2255 10847 2275
rect 10813 2245 10847 2255
rect 12973 2275 13007 2285
rect 12973 2255 12981 2275
rect 12999 2255 13007 2275
rect 12973 2245 13007 2255
rect 18313 2275 18347 2285
rect 18313 2255 18321 2275
rect 18339 2255 18347 2275
rect 18313 2245 18347 2255
rect 20473 2275 20507 2285
rect 20473 2255 20481 2275
rect 20499 2255 20507 2275
rect 20473 2245 20507 2255
rect 9640 2215 9680 2225
rect 9640 2195 9650 2215
rect 9670 2195 9680 2215
rect 10820 2195 10835 2245
rect 10930 2215 10970 2225
rect 10930 2195 10940 2215
rect 10960 2195 10970 2215
rect 9640 2180 9735 2195
rect 9720 2170 9735 2180
rect 9775 2180 10835 2195
rect 9775 2170 9790 2180
rect 9830 2170 9845 2180
rect 9885 2170 9900 2180
rect 9940 2170 9955 2180
rect 9995 2170 10010 2180
rect 10050 2170 10065 2180
rect 10105 2170 10120 2180
rect 10160 2170 10175 2180
rect 10215 2170 10230 2180
rect 10270 2170 10285 2180
rect 10325 2170 10340 2180
rect 10380 2170 10395 2180
rect 10435 2170 10450 2180
rect 10490 2170 10505 2180
rect 10545 2170 10560 2180
rect 10600 2170 10615 2180
rect 10655 2170 10670 2180
rect 10710 2170 10725 2180
rect 10765 2170 10780 2180
rect 10820 2170 10835 2180
rect 10875 2180 10970 2195
rect 12850 2215 12890 2225
rect 12850 2195 12860 2215
rect 12880 2195 12890 2215
rect 12985 2195 13000 2245
rect 14140 2215 14180 2225
rect 14140 2195 14150 2215
rect 14170 2195 14180 2215
rect 12850 2180 12945 2195
rect 10875 2170 10890 2180
rect 12930 2170 12945 2180
rect 12985 2180 14045 2195
rect 12985 2170 13000 2180
rect 13040 2170 13055 2180
rect 13095 2170 13110 2180
rect 13150 2170 13165 2180
rect 13205 2170 13220 2180
rect 13260 2170 13275 2180
rect 13315 2170 13330 2180
rect 13370 2170 13385 2180
rect 13425 2170 13440 2180
rect 13480 2170 13495 2180
rect 13535 2170 13550 2180
rect 13590 2170 13605 2180
rect 13645 2170 13660 2180
rect 13700 2170 13715 2180
rect 13755 2170 13770 2180
rect 13810 2170 13825 2180
rect 13865 2170 13880 2180
rect 13920 2170 13935 2180
rect 13975 2170 13990 2180
rect 14030 2170 14045 2180
rect 14085 2180 14180 2195
rect 17140 2215 17180 2225
rect 17140 2195 17150 2215
rect 17170 2195 17180 2215
rect 18320 2195 18335 2245
rect 18430 2215 18470 2225
rect 18430 2195 18440 2215
rect 18460 2195 18470 2215
rect 17140 2180 17235 2195
rect 14085 2170 14100 2180
rect 17220 2170 17235 2180
rect 17275 2180 18335 2195
rect 17275 2170 17290 2180
rect 17330 2170 17345 2180
rect 17385 2170 17400 2180
rect 17440 2170 17455 2180
rect 17495 2170 17510 2180
rect 17550 2170 17565 2180
rect 17605 2170 17620 2180
rect 17660 2170 17675 2180
rect 17715 2170 17730 2180
rect 17770 2170 17785 2180
rect 17825 2170 17840 2180
rect 17880 2170 17895 2180
rect 17935 2170 17950 2180
rect 17990 2170 18005 2180
rect 18045 2170 18060 2180
rect 18100 2170 18115 2180
rect 18155 2170 18170 2180
rect 18210 2170 18225 2180
rect 18265 2170 18280 2180
rect 18320 2170 18335 2180
rect 18375 2180 18470 2195
rect 20350 2215 20390 2225
rect 20350 2195 20360 2215
rect 20380 2195 20390 2215
rect 20485 2195 20500 2245
rect 21640 2215 21680 2225
rect 21640 2195 21650 2215
rect 21670 2195 21680 2215
rect 20350 2180 20445 2195
rect 18375 2170 18390 2180
rect 20430 2170 20445 2180
rect 20485 2180 21545 2195
rect 20485 2170 20500 2180
rect 20540 2170 20555 2180
rect 20595 2170 20610 2180
rect 20650 2170 20665 2180
rect 20705 2170 20720 2180
rect 20760 2170 20775 2180
rect 20815 2170 20830 2180
rect 20870 2170 20885 2180
rect 20925 2170 20940 2180
rect 20980 2170 20995 2180
rect 21035 2170 21050 2180
rect 21090 2170 21105 2180
rect 21145 2170 21160 2180
rect 21200 2170 21215 2180
rect 21255 2170 21270 2180
rect 21310 2170 21325 2180
rect 21365 2170 21380 2180
rect 21420 2170 21435 2180
rect 21475 2170 21490 2180
rect 21530 2170 21545 2180
rect 21585 2180 21680 2195
rect 21585 2170 21600 2180
rect 11315 2130 11330 2145
rect 11370 2140 12430 2155
rect 11370 2130 11385 2140
rect 11425 2130 11440 2140
rect 11480 2130 11495 2140
rect 11535 2130 11550 2140
rect 11590 2130 11605 2140
rect 11645 2130 11660 2140
rect 11700 2130 11715 2140
rect 11755 2130 11770 2140
rect 11810 2130 11825 2140
rect 11865 2130 11880 2140
rect 11920 2130 11935 2140
rect 11975 2130 11990 2140
rect 12030 2130 12045 2140
rect 12085 2130 12100 2140
rect 12140 2130 12155 2140
rect 12195 2130 12210 2140
rect 12250 2130 12265 2140
rect 12305 2130 12320 2140
rect 12360 2130 12375 2140
rect 12415 2130 12430 2140
rect 12470 2130 12485 2145
rect 2605 2000 2620 2015
rect 2660 2000 2675 2015
rect 2785 2000 2805 2015
rect 2845 2000 2865 2015
rect 2905 2000 2925 2015
rect 2965 2000 2985 2015
rect 3025 2000 3045 2015
rect 3085 2000 3105 2015
rect 3145 2000 3165 2015
rect 3205 2000 3225 2015
rect 3265 2000 3285 2015
rect 3325 2000 3345 2015
rect 3385 2000 3405 2015
rect 3445 2000 3465 2015
rect 3505 2000 3525 2015
rect 3565 2000 3585 2015
rect 3625 2000 3645 2015
rect 3685 2000 3705 2015
rect 3745 2000 3765 2015
rect 3805 2000 3825 2015
rect 3865 2000 3885 2015
rect 3925 2000 3945 2015
rect 4065 2000 4085 2015
rect 4125 2000 4145 2015
rect 4185 2000 4205 2015
rect 4245 2000 4265 2015
rect 4305 2000 4325 2015
rect 4365 2000 4385 2015
rect 4425 2000 4445 2015
rect 4485 2000 4505 2015
rect 4545 2000 4565 2015
rect 4605 2000 4625 2015
rect 4665 2000 4685 2015
rect 4725 2000 4745 2015
rect 4785 2000 4805 2015
rect 4845 2000 4865 2015
rect 4905 2000 4925 2015
rect 4965 2000 4985 2015
rect 5025 2000 5045 2015
rect 5085 2000 5105 2015
rect 5145 2000 5165 2015
rect 5205 2000 5225 2015
rect 9720 2005 9735 2020
rect 9775 2005 9790 2020
rect 9830 2005 9845 2020
rect 9885 2005 9900 2020
rect 9940 2005 9955 2020
rect 9995 2005 10010 2020
rect 10050 2005 10065 2020
rect 10105 2005 10120 2020
rect 10160 2005 10175 2020
rect 10215 2005 10230 2020
rect 10270 2005 10285 2020
rect 10325 2005 10340 2020
rect 10380 2005 10395 2020
rect 10435 2005 10450 2020
rect 10490 2005 10505 2020
rect 10545 2005 10560 2020
rect 10600 2005 10615 2020
rect 10655 2005 10670 2020
rect 10710 2005 10725 2020
rect 10765 2005 10780 2020
rect 10820 2005 10835 2020
rect 10875 2005 10890 2020
rect 18815 2130 18830 2145
rect 18870 2140 19930 2155
rect 18870 2130 18885 2140
rect 18925 2130 18940 2140
rect 18980 2130 18995 2140
rect 19035 2130 19050 2140
rect 19090 2130 19105 2140
rect 19145 2130 19160 2140
rect 19200 2130 19215 2140
rect 19255 2130 19270 2140
rect 19310 2130 19325 2140
rect 19365 2130 19380 2140
rect 19420 2130 19435 2140
rect 19475 2130 19490 2140
rect 19530 2130 19545 2140
rect 19585 2130 19600 2140
rect 19640 2130 19655 2140
rect 19695 2130 19710 2140
rect 19750 2130 19765 2140
rect 19805 2130 19820 2140
rect 19860 2130 19875 2140
rect 19915 2130 19930 2140
rect 19970 2130 19985 2145
rect 12930 2005 12945 2020
rect 12985 2005 13000 2020
rect 13040 2005 13055 2020
rect 13095 2005 13110 2020
rect 13150 2005 13165 2020
rect 13205 2005 13220 2020
rect 13260 2005 13275 2020
rect 13315 2005 13330 2020
rect 13370 2005 13385 2020
rect 13425 2005 13440 2020
rect 13480 2005 13495 2020
rect 13535 2005 13550 2020
rect 13590 2005 13605 2020
rect 13645 2005 13660 2020
rect 13700 2005 13715 2020
rect 13755 2005 13770 2020
rect 13810 2005 13825 2020
rect 13865 2005 13880 2020
rect 13920 2005 13935 2020
rect 13975 2005 13990 2020
rect 14030 2005 14045 2020
rect 14085 2005 14100 2020
rect 17220 2005 17235 2020
rect 17275 2005 17290 2020
rect 17330 2005 17345 2020
rect 17385 2005 17400 2020
rect 17440 2005 17455 2020
rect 17495 2005 17510 2020
rect 17550 2005 17565 2020
rect 17605 2005 17620 2020
rect 17660 2005 17675 2020
rect 17715 2005 17730 2020
rect 17770 2005 17785 2020
rect 17825 2005 17840 2020
rect 17880 2005 17895 2020
rect 17935 2005 17950 2020
rect 17990 2005 18005 2020
rect 18045 2005 18060 2020
rect 18100 2005 18115 2020
rect 18155 2005 18170 2020
rect 18210 2005 18225 2020
rect 18265 2005 18280 2020
rect 18320 2005 18335 2020
rect 18375 2005 18390 2020
rect 20430 2005 20445 2020
rect 20485 2005 20500 2020
rect 20540 2005 20555 2020
rect 20595 2005 20610 2020
rect 20650 2005 20665 2020
rect 20705 2005 20720 2020
rect 20760 2005 20775 2020
rect 20815 2005 20830 2020
rect 20870 2005 20885 2020
rect 20925 2005 20940 2020
rect 20980 2005 20995 2020
rect 21035 2005 21050 2020
rect 21090 2005 21105 2020
rect 21145 2005 21160 2020
rect 21200 2005 21215 2020
rect 21255 2005 21270 2020
rect 21310 2005 21325 2020
rect 21365 2005 21380 2020
rect 21420 2005 21435 2020
rect 21475 2005 21490 2020
rect 21530 2005 21545 2020
rect 21585 2005 21600 2020
rect 11315 1970 11330 1980
rect 11235 1955 11330 1970
rect 11370 1965 11385 1980
rect 11425 1965 11440 1980
rect 11480 1965 11495 1980
rect 11535 1965 11550 1980
rect 11590 1965 11605 1980
rect 11645 1965 11660 1980
rect 11700 1965 11715 1980
rect 11755 1965 11770 1980
rect 11810 1965 11825 1980
rect 11865 1965 11880 1980
rect 11920 1965 11935 1980
rect 11975 1965 11990 1980
rect 12030 1965 12045 1980
rect 12085 1965 12100 1980
rect 12140 1965 12155 1980
rect 12195 1965 12210 1980
rect 12250 1965 12265 1980
rect 12305 1965 12320 1980
rect 12360 1965 12375 1980
rect 12415 1965 12430 1980
rect 12470 1970 12485 1980
rect 18815 1970 18830 1980
rect 12470 1955 12565 1970
rect 11235 1935 11245 1955
rect 11265 1935 11275 1955
rect 11235 1925 11275 1935
rect 12525 1935 12535 1955
rect 12555 1935 12565 1955
rect 12525 1925 12565 1935
rect 18735 1955 18830 1970
rect 18870 1965 18885 1980
rect 18925 1965 18940 1980
rect 18980 1965 18995 1980
rect 19035 1965 19050 1980
rect 19090 1965 19105 1980
rect 19145 1965 19160 1980
rect 19200 1965 19215 1980
rect 19255 1965 19270 1980
rect 19310 1965 19325 1980
rect 19365 1965 19380 1980
rect 19420 1965 19435 1980
rect 19475 1965 19490 1980
rect 19530 1965 19545 1980
rect 19585 1965 19600 1980
rect 19640 1965 19655 1980
rect 19695 1965 19710 1980
rect 19750 1965 19765 1980
rect 19805 1965 19820 1980
rect 19860 1965 19875 1980
rect 19915 1965 19930 1980
rect 19970 1970 19985 1980
rect 19970 1955 20065 1970
rect 18735 1935 18745 1955
rect 18765 1935 18775 1955
rect 18735 1925 18775 1935
rect 20025 1935 20035 1955
rect 20055 1935 20065 1955
rect 20025 1925 20065 1935
rect 20450 1900 20490 1910
rect 2605 1890 2620 1900
rect 2660 1890 2675 1900
rect 2605 1875 2675 1890
rect 2785 1885 2805 1900
rect 2845 1885 2865 1900
rect 2905 1890 2925 1900
rect 2965 1890 2985 1900
rect 3025 1890 3045 1900
rect 3085 1890 3105 1900
rect 2765 1875 2805 1885
rect 2620 1855 2630 1875
rect 2650 1855 2660 1875
rect 2620 1845 2660 1855
rect 2765 1855 2775 1875
rect 2795 1855 2805 1875
rect 2765 1845 2805 1855
rect 2835 1875 2875 1885
rect 2905 1875 3105 1890
rect 3145 1890 3165 1900
rect 3205 1890 3225 1900
rect 3145 1875 3225 1890
rect 3265 1890 3285 1900
rect 3325 1890 3345 1900
rect 3385 1890 3405 1900
rect 3445 1890 3465 1900
rect 3265 1875 3465 1890
rect 3505 1890 3525 1900
rect 3565 1890 3585 1900
rect 3505 1875 3585 1890
rect 3625 1890 3645 1900
rect 3685 1890 3705 1900
rect 3745 1890 3765 1900
rect 3805 1890 3825 1900
rect 3625 1875 3825 1890
rect 3865 1885 3885 1900
rect 3925 1890 3945 1900
rect 4065 1890 4085 1900
rect 3855 1875 3895 1885
rect 3925 1875 4085 1890
rect 4125 1885 4145 1900
rect 4185 1890 4205 1900
rect 4245 1890 4265 1900
rect 4305 1890 4325 1900
rect 4365 1890 4385 1900
rect 4115 1875 4155 1885
rect 4185 1875 4385 1890
rect 4425 1890 4445 1900
rect 4485 1890 4505 1900
rect 4425 1875 4505 1890
rect 4545 1890 4565 1900
rect 4605 1890 4625 1900
rect 4665 1890 4685 1900
rect 4725 1890 4745 1900
rect 4545 1875 4745 1890
rect 4785 1890 4805 1900
rect 4845 1890 4865 1900
rect 4785 1875 4865 1890
rect 4905 1890 4925 1900
rect 4965 1890 4985 1900
rect 5025 1890 5045 1900
rect 5085 1890 5105 1900
rect 4905 1875 5105 1890
rect 5145 1885 5165 1900
rect 5205 1885 5225 1900
rect 5135 1875 5175 1885
rect 2835 1855 2845 1875
rect 2865 1855 2875 1875
rect 2835 1845 2875 1855
rect 2925 1855 2935 1875
rect 2955 1855 2965 1875
rect 2925 1845 2965 1855
rect 3165 1855 3175 1875
rect 3195 1855 3205 1875
rect 3165 1845 3205 1855
rect 3285 1855 3295 1875
rect 3315 1855 3325 1875
rect 3285 1845 3325 1855
rect 3525 1855 3535 1875
rect 3555 1855 3565 1875
rect 3525 1845 3565 1855
rect 3645 1855 3655 1875
rect 3675 1855 3685 1875
rect 3645 1845 3685 1855
rect 3855 1855 3865 1875
rect 3885 1855 3895 1875
rect 3855 1845 3895 1855
rect 3985 1870 4025 1875
rect 3985 1850 3995 1870
rect 4015 1850 4025 1870
rect 3985 1840 4025 1850
rect 4115 1855 4125 1875
rect 4145 1855 4155 1875
rect 4115 1845 4155 1855
rect 4325 1855 4335 1875
rect 4355 1855 4365 1875
rect 4325 1845 4365 1855
rect 4445 1855 4455 1875
rect 4475 1855 4485 1875
rect 4445 1845 4485 1855
rect 4685 1855 4695 1875
rect 4715 1855 4725 1875
rect 4685 1845 4725 1855
rect 4805 1855 4815 1875
rect 4835 1855 4845 1875
rect 4805 1845 4845 1855
rect 5045 1855 5055 1875
rect 5075 1855 5085 1875
rect 5045 1845 5085 1855
rect 5135 1855 5145 1875
rect 5165 1855 5175 1875
rect 5135 1845 5175 1855
rect 5205 1875 5245 1885
rect 5205 1855 5215 1875
rect 5235 1855 5245 1875
rect 20450 1880 20460 1900
rect 20480 1880 20490 1900
rect 20860 1900 20900 1910
rect 20860 1880 20870 1900
rect 20890 1880 20900 1900
rect 20450 1865 20545 1880
rect 20530 1855 20545 1865
rect 20585 1855 20600 1870
rect 20640 1855 20655 1870
rect 20695 1855 20710 1870
rect 20750 1855 20765 1870
rect 20805 1865 20900 1880
rect 20805 1855 20820 1865
rect 5205 1845 5245 1855
rect 3225 1755 3265 1765
rect 3225 1735 3235 1755
rect 3255 1735 3265 1755
rect 3225 1720 3265 1735
rect 4745 1755 4785 1765
rect 4745 1735 4755 1755
rect 4775 1735 4785 1755
rect 4745 1720 4785 1735
rect 3225 1705 3765 1720
rect 3205 1665 3225 1680
rect 3265 1665 3285 1705
rect 3325 1665 3345 1705
rect 3385 1665 3405 1680
rect 3445 1665 3465 1680
rect 3505 1665 3525 1705
rect 3565 1665 3585 1705
rect 3625 1665 3645 1680
rect 3685 1665 3705 1680
rect 3745 1665 3765 1705
rect 4245 1705 4785 1720
rect 11237 1710 11269 1720
rect 4245 1665 4265 1705
rect 4305 1665 4325 1680
rect 4365 1665 4385 1680
rect 4425 1665 4445 1705
rect 4485 1665 4505 1705
rect 4545 1665 4565 1680
rect 4605 1665 4625 1680
rect 4665 1665 4685 1705
rect 4725 1665 4745 1705
rect 11237 1690 11243 1710
rect 11260 1690 11269 1710
rect 11457 1710 11489 1720
rect 11457 1690 11463 1710
rect 11480 1690 11489 1710
rect 11180 1680 11269 1690
rect 11400 1680 11489 1690
rect 11601 1710 11635 1720
rect 11601 1690 11610 1710
rect 11627 1690 11635 1710
rect 11867 1710 11899 1720
rect 11867 1695 11876 1710
rect 11601 1680 11635 1690
rect 11865 1690 11876 1695
rect 11893 1690 11899 1710
rect 12277 1710 12309 1720
rect 12277 1690 12283 1710
rect 12300 1690 12309 1710
rect 12497 1710 12529 1720
rect 12497 1690 12503 1710
rect 12520 1690 12529 1710
rect 11865 1680 11899 1690
rect 12220 1680 12309 1690
rect 12440 1680 12529 1690
rect 12641 1710 12675 1720
rect 12641 1690 12650 1710
rect 12667 1690 12675 1710
rect 18737 1710 18769 1720
rect 18737 1690 18743 1710
rect 18760 1690 18769 1710
rect 18957 1710 18989 1720
rect 18957 1690 18963 1710
rect 18980 1690 18989 1710
rect 12641 1680 12675 1690
rect 18680 1680 18769 1690
rect 18900 1680 18989 1690
rect 19101 1710 19135 1720
rect 19101 1690 19110 1710
rect 19127 1690 19135 1710
rect 19367 1710 19399 1720
rect 19367 1695 19376 1710
rect 19101 1680 19135 1690
rect 19365 1690 19376 1695
rect 19393 1690 19399 1710
rect 19777 1710 19809 1720
rect 19777 1690 19783 1710
rect 19800 1690 19809 1710
rect 19997 1710 20029 1720
rect 19997 1690 20003 1710
rect 20020 1690 20029 1710
rect 19365 1680 19399 1690
rect 19720 1680 19809 1690
rect 19940 1680 20029 1690
rect 20141 1710 20175 1720
rect 20141 1690 20150 1710
rect 20167 1690 20175 1710
rect 20530 1690 20545 1705
rect 20585 1695 20600 1705
rect 20640 1695 20655 1705
rect 20695 1695 20710 1705
rect 20750 1695 20765 1705
rect 20141 1680 20175 1690
rect 20585 1685 20765 1695
rect 20805 1690 20820 1705
rect 20566 1680 20765 1685
rect 4785 1665 4805 1680
rect 11070 1665 11085 1680
rect 11125 1665 11140 1680
rect 11180 1675 11250 1680
rect 11180 1665 11195 1675
rect 11235 1665 11250 1675
rect 11290 1665 11305 1680
rect 11345 1665 11360 1680
rect 11400 1675 11470 1680
rect 11400 1665 11415 1675
rect 11455 1665 11470 1675
rect 11510 1665 11525 1680
rect 11565 1665 11580 1680
rect 11620 1665 11635 1680
rect 11675 1665 11690 1680
rect 11810 1665 11825 1680
rect 11865 1665 11880 1680
rect 11920 1665 11935 1680
rect 11975 1665 11990 1680
rect 12110 1665 12125 1680
rect 12165 1665 12180 1680
rect 12220 1675 12290 1680
rect 12220 1665 12235 1675
rect 12275 1665 12290 1675
rect 12330 1665 12345 1680
rect 12385 1665 12400 1680
rect 12440 1675 12510 1680
rect 12440 1665 12455 1675
rect 12495 1665 12510 1675
rect 12550 1665 12565 1680
rect 12605 1665 12620 1680
rect 12660 1665 12675 1680
rect 12715 1665 12730 1680
rect 18570 1665 18585 1680
rect 18625 1665 18640 1680
rect 18680 1675 18750 1680
rect 18680 1665 18695 1675
rect 18735 1665 18750 1675
rect 18790 1665 18805 1680
rect 18845 1665 18860 1680
rect 18900 1675 18970 1680
rect 18900 1665 18915 1675
rect 18955 1665 18970 1675
rect 19010 1665 19025 1680
rect 19065 1665 19080 1680
rect 19120 1665 19135 1680
rect 19175 1665 19190 1680
rect 19310 1665 19325 1680
rect 19365 1665 19380 1680
rect 19420 1665 19435 1680
rect 19475 1665 19490 1680
rect 19610 1665 19625 1680
rect 19665 1665 19680 1680
rect 19720 1675 19790 1680
rect 19720 1665 19735 1675
rect 19775 1665 19790 1675
rect 19830 1665 19845 1680
rect 19885 1665 19900 1680
rect 19940 1675 20010 1680
rect 19940 1665 19955 1675
rect 19995 1665 20010 1675
rect 20050 1665 20065 1680
rect 20105 1665 20120 1680
rect 20160 1665 20175 1680
rect 20215 1665 20230 1680
rect 20566 1675 20600 1680
rect 3205 1600 3225 1615
rect 3265 1600 3285 1615
rect 3325 1600 3345 1615
rect 3165 1590 3225 1600
rect 3165 1570 3175 1590
rect 3195 1575 3225 1590
rect 3385 1575 3405 1615
rect 3445 1575 3465 1615
rect 3505 1600 3525 1615
rect 3565 1600 3585 1615
rect 3625 1575 3645 1615
rect 3685 1575 3705 1615
rect 3745 1600 3765 1615
rect 4245 1600 4265 1615
rect 3195 1570 3705 1575
rect 3165 1560 3705 1570
rect 4305 1575 4325 1615
rect 4365 1575 4385 1615
rect 4425 1600 4445 1615
rect 4485 1600 4505 1615
rect 4545 1575 4565 1615
rect 4605 1575 4625 1615
rect 4665 1600 4685 1615
rect 4725 1600 4745 1615
rect 4785 1600 4805 1615
rect 4785 1590 4845 1600
rect 4785 1575 4815 1590
rect 4305 1570 4815 1575
rect 4835 1570 4845 1590
rect 4305 1560 4845 1570
rect 20566 1655 20571 1675
rect 20591 1670 20600 1675
rect 20591 1655 20598 1670
rect 20566 1645 20598 1655
rect 20471 1565 20503 1575
rect 20471 1545 20476 1565
rect 20496 1550 20503 1565
rect 20847 1565 20879 1575
rect 20847 1550 20854 1565
rect 20496 1545 20505 1550
rect 20471 1535 20505 1545
rect 20845 1545 20854 1550
rect 20874 1545 20879 1565
rect 20845 1535 20879 1545
rect 20435 1520 20450 1535
rect 20490 1520 20505 1535
rect 20545 1520 20560 1535
rect 20600 1520 20615 1535
rect 20735 1520 20750 1535
rect 20790 1520 20805 1535
rect 20845 1520 20860 1535
rect 20900 1520 20915 1535
rect 11070 1505 11085 1515
rect 2925 1495 2965 1505
rect 2925 1475 2935 1495
rect 2955 1475 2965 1495
rect 2925 1470 2965 1475
rect 3045 1495 3085 1505
rect 3045 1475 3055 1495
rect 3075 1475 3085 1495
rect 3045 1470 3085 1475
rect 3165 1495 3205 1505
rect 3165 1475 3175 1495
rect 3195 1475 3205 1495
rect 3165 1470 3205 1475
rect 3285 1495 3325 1505
rect 3285 1475 3295 1495
rect 3315 1475 3325 1495
rect 3285 1470 3325 1475
rect 3525 1495 3565 1505
rect 3525 1475 3535 1495
rect 3555 1475 3565 1495
rect 3525 1470 3565 1475
rect 3645 1495 3685 1505
rect 3645 1475 3655 1495
rect 3675 1475 3685 1495
rect 3645 1470 3685 1475
rect 3765 1495 3805 1505
rect 3765 1475 3775 1495
rect 3795 1475 3805 1495
rect 3765 1470 3805 1475
rect 4205 1495 4245 1505
rect 4205 1475 4215 1495
rect 4235 1475 4245 1495
rect 4205 1470 4245 1475
rect 4325 1495 4365 1505
rect 4325 1475 4335 1495
rect 4355 1475 4365 1495
rect 4325 1470 4365 1475
rect 4445 1495 4485 1505
rect 4445 1475 4455 1495
rect 4475 1475 4485 1495
rect 4445 1470 4485 1475
rect 4685 1495 4725 1505
rect 4685 1475 4695 1495
rect 4715 1475 4725 1495
rect 4685 1470 4725 1475
rect 4805 1495 4845 1505
rect 4805 1475 4815 1495
rect 4835 1475 4845 1495
rect 4805 1470 4845 1475
rect 4925 1495 4965 1505
rect 4925 1475 4935 1495
rect 4955 1475 4965 1495
rect 4925 1470 4965 1475
rect 5045 1495 5085 1505
rect 5045 1475 5055 1495
rect 5075 1475 5085 1495
rect 5045 1470 5085 1475
rect 10990 1490 11085 1505
rect 11125 1500 11140 1515
rect 11180 1500 11195 1515
rect 11235 1500 11250 1515
rect 11290 1505 11305 1515
rect 11345 1505 11360 1515
rect 11106 1490 11140 1500
rect 11290 1490 11360 1505
rect 11400 1500 11415 1515
rect 11455 1500 11470 1515
rect 11510 1505 11525 1515
rect 11565 1505 11580 1515
rect 11510 1490 11580 1505
rect 11620 1500 11635 1515
rect 11675 1505 11690 1515
rect 11810 1505 11825 1515
rect 11675 1490 11825 1505
rect 11865 1500 11880 1515
rect 11920 1500 11935 1515
rect 11975 1505 11990 1515
rect 12110 1505 12125 1515
rect 11920 1490 11954 1500
rect 11975 1490 12125 1505
rect 12165 1500 12180 1515
rect 12220 1500 12235 1515
rect 12275 1500 12290 1515
rect 12330 1505 12345 1515
rect 12385 1505 12400 1515
rect 12146 1490 12180 1500
rect 12330 1490 12400 1505
rect 12440 1500 12455 1515
rect 12495 1500 12510 1515
rect 12550 1505 12565 1515
rect 12605 1505 12620 1515
rect 12550 1490 12620 1505
rect 12660 1500 12675 1515
rect 12715 1505 12730 1515
rect 18570 1505 18585 1515
rect 12715 1490 12810 1505
rect 10990 1470 11000 1490
rect 11020 1470 11030 1490
rect 2875 1455 3375 1470
rect 3415 1455 3915 1470
rect 4095 1455 4595 1470
rect 4635 1455 5135 1470
rect 10990 1460 11030 1470
rect 11106 1470 11112 1490
rect 11129 1470 11138 1490
rect 11106 1460 11138 1470
rect 11305 1470 11315 1490
rect 11335 1470 11345 1490
rect 11305 1460 11345 1470
rect 11525 1470 11535 1490
rect 11555 1470 11565 1490
rect 11525 1460 11565 1470
rect 11730 1470 11740 1490
rect 11760 1470 11770 1490
rect 11730 1460 11770 1470
rect 11922 1470 11928 1490
rect 11945 1470 11954 1490
rect 11922 1460 11954 1470
rect 12030 1470 12040 1490
rect 12060 1470 12070 1490
rect 12030 1460 12070 1470
rect 12146 1470 12152 1490
rect 12169 1470 12178 1490
rect 12146 1460 12178 1470
rect 12345 1470 12355 1490
rect 12375 1470 12385 1490
rect 12345 1460 12385 1470
rect 12565 1470 12575 1490
rect 12595 1470 12605 1490
rect 12565 1460 12605 1470
rect 12770 1470 12780 1490
rect 12800 1470 12810 1490
rect 12770 1460 12810 1470
rect 18490 1490 18585 1505
rect 18625 1500 18640 1515
rect 18680 1500 18695 1515
rect 18735 1500 18750 1515
rect 18790 1505 18805 1515
rect 18845 1505 18860 1515
rect 18606 1490 18640 1500
rect 18790 1490 18860 1505
rect 18900 1500 18915 1515
rect 18955 1500 18970 1515
rect 19010 1505 19025 1515
rect 19065 1505 19080 1515
rect 19010 1490 19080 1505
rect 19120 1500 19135 1515
rect 19175 1505 19190 1515
rect 19310 1505 19325 1515
rect 19175 1490 19325 1505
rect 19365 1500 19380 1515
rect 19420 1500 19435 1515
rect 19475 1505 19490 1515
rect 19610 1505 19625 1515
rect 19420 1490 19454 1500
rect 19475 1490 19625 1505
rect 19665 1500 19680 1515
rect 19720 1500 19735 1515
rect 19775 1500 19790 1515
rect 19830 1505 19845 1515
rect 19885 1505 19900 1515
rect 19646 1490 19680 1500
rect 19830 1490 19900 1505
rect 19940 1500 19955 1515
rect 19995 1500 20010 1515
rect 20050 1505 20065 1515
rect 20105 1505 20120 1515
rect 20050 1490 20120 1505
rect 20160 1500 20175 1515
rect 20215 1505 20230 1515
rect 20215 1490 20310 1505
rect 18490 1470 18500 1490
rect 18520 1470 18530 1490
rect 18490 1460 18530 1470
rect 18606 1470 18612 1490
rect 18629 1470 18638 1490
rect 18606 1460 18638 1470
rect 18805 1470 18815 1490
rect 18835 1470 18845 1490
rect 18805 1460 18845 1470
rect 19025 1470 19035 1490
rect 19055 1470 19065 1490
rect 19025 1460 19065 1470
rect 19230 1470 19240 1490
rect 19260 1470 19270 1490
rect 19230 1460 19270 1470
rect 19422 1470 19428 1490
rect 19445 1470 19454 1490
rect 19422 1460 19454 1470
rect 19530 1470 19540 1490
rect 19560 1470 19570 1490
rect 19530 1460 19570 1470
rect 19646 1470 19652 1490
rect 19669 1470 19678 1490
rect 19646 1460 19678 1470
rect 19845 1470 19855 1490
rect 19875 1470 19885 1490
rect 19845 1460 19885 1470
rect 20065 1470 20075 1490
rect 20095 1470 20105 1490
rect 20065 1460 20105 1470
rect 20270 1470 20280 1490
rect 20300 1470 20310 1490
rect 20270 1460 20310 1470
rect 20435 1360 20450 1370
rect 20355 1345 20450 1360
rect 20490 1355 20505 1370
rect 20545 1355 20560 1370
rect 20526 1345 20560 1355
rect 20600 1360 20615 1370
rect 20735 1360 20750 1370
rect 20600 1345 20750 1360
rect 20790 1355 20805 1370
rect 20845 1355 20860 1370
rect 20900 1360 20915 1370
rect 20790 1345 20824 1355
rect 20900 1345 20995 1360
rect 20355 1325 20365 1345
rect 20385 1325 20395 1345
rect 13128 1315 13162 1325
rect 20355 1315 20395 1325
rect 20526 1325 20533 1345
rect 20553 1340 20560 1345
rect 20553 1325 20558 1340
rect 20526 1315 20558 1325
rect 20655 1325 20665 1345
rect 20685 1325 20695 1345
rect 20790 1340 20797 1345
rect 20655 1315 20695 1325
rect 20792 1325 20797 1340
rect 20817 1325 20824 1345
rect 20792 1315 20824 1325
rect 20955 1325 20965 1345
rect 20985 1325 20995 1345
rect 20955 1315 20995 1325
rect 13128 1295 13136 1315
rect 13154 1295 13162 1315
rect 12965 1270 13025 1285
rect 13065 1280 14025 1295
rect 20095 1285 20135 1295
rect 13065 1270 13125 1280
rect 13165 1270 13225 1280
rect 13265 1270 13325 1280
rect 13365 1270 13425 1280
rect 13465 1270 13525 1280
rect 13565 1270 13625 1280
rect 13665 1270 13725 1280
rect 13765 1270 13825 1280
rect 13865 1270 13925 1280
rect 13965 1270 14025 1280
rect 14065 1270 14125 1285
rect 20095 1280 20105 1285
rect 19315 1270 19345 1280
rect 12595 1235 12635 1245
rect 12595 1230 12605 1235
rect 11815 1220 11845 1230
rect 2875 1190 3375 1205
rect 3415 1190 3915 1205
rect 4095 1190 4595 1205
rect 4635 1190 5135 1205
rect 11815 1200 11820 1220
rect 11840 1200 11845 1220
rect 12510 1215 12605 1230
rect 12625 1215 12635 1235
rect 11245 1175 11260 1190
rect 11300 1185 12360 1200
rect 11300 1175 11315 1185
rect 11355 1175 11370 1185
rect 11410 1175 11425 1185
rect 11465 1175 11480 1185
rect 11520 1175 11535 1185
rect 11575 1175 11590 1185
rect 11630 1175 11645 1185
rect 11685 1175 11700 1185
rect 11740 1175 11755 1185
rect 11795 1175 11810 1185
rect 11850 1175 11865 1185
rect 11905 1175 11920 1185
rect 11960 1175 11975 1185
rect 12015 1175 12030 1185
rect 12070 1175 12085 1185
rect 12125 1175 12140 1185
rect 12180 1175 12195 1185
rect 12235 1175 12250 1185
rect 12290 1175 12305 1185
rect 12345 1175 12360 1185
rect 12400 1185 12470 1200
rect 12400 1175 12415 1185
rect 12455 1175 12470 1185
rect 12510 1175 12525 1215
rect 12595 1205 12635 1215
rect 12565 1175 12580 1190
rect 3025 1120 3065 1130
rect 3025 1100 3035 1120
rect 3055 1100 3065 1120
rect 3025 1090 3065 1100
rect 3105 1120 3145 1130
rect 3105 1100 3115 1120
rect 3135 1100 3145 1120
rect 3105 1090 3145 1100
rect 3185 1120 3225 1130
rect 3185 1100 3195 1120
rect 3215 1100 3225 1120
rect 3185 1090 3225 1100
rect 3265 1120 3305 1130
rect 3265 1100 3275 1120
rect 3295 1100 3305 1120
rect 3265 1090 3305 1100
rect 3345 1120 3385 1130
rect 3345 1100 3355 1120
rect 3375 1100 3385 1120
rect 3345 1090 3385 1100
rect 3425 1120 3465 1130
rect 3425 1100 3435 1120
rect 3455 1100 3465 1120
rect 3425 1090 3465 1100
rect 3505 1120 3545 1130
rect 3505 1100 3515 1120
rect 3535 1100 3545 1120
rect 3505 1090 3545 1100
rect 3585 1120 3625 1130
rect 3585 1100 3595 1120
rect 3615 1100 3625 1120
rect 3585 1090 3625 1100
rect 3665 1120 3705 1130
rect 3665 1100 3675 1120
rect 3695 1100 3705 1120
rect 3665 1090 3705 1100
rect 3745 1120 3785 1130
rect 3745 1100 3755 1120
rect 3775 1100 3785 1120
rect 3745 1090 3785 1100
rect 3825 1120 3865 1130
rect 3825 1100 3835 1120
rect 3855 1100 3865 1120
rect 3825 1090 3865 1100
rect 3905 1120 3945 1130
rect 3905 1100 3915 1120
rect 3935 1100 3945 1120
rect 3905 1090 3945 1100
rect 4065 1120 4105 1130
rect 4065 1100 4075 1120
rect 4095 1100 4105 1120
rect 4065 1090 4105 1100
rect 4145 1120 4185 1130
rect 4145 1100 4155 1120
rect 4175 1100 4185 1120
rect 4145 1090 4185 1100
rect 4225 1120 4265 1130
rect 4225 1100 4235 1120
rect 4255 1100 4265 1120
rect 4225 1090 4265 1100
rect 4305 1120 4345 1130
rect 4305 1100 4315 1120
rect 4335 1100 4345 1120
rect 4305 1090 4345 1100
rect 4385 1120 4425 1130
rect 4385 1100 4395 1120
rect 4415 1100 4425 1120
rect 4385 1090 4425 1100
rect 4465 1120 4505 1130
rect 4465 1100 4475 1120
rect 4495 1100 4505 1120
rect 4465 1090 4505 1100
rect 4545 1120 4585 1130
rect 4545 1100 4555 1120
rect 4575 1100 4585 1120
rect 4545 1090 4585 1100
rect 4625 1120 4665 1130
rect 4625 1100 4635 1120
rect 4655 1100 4665 1120
rect 4625 1090 4665 1100
rect 4705 1120 4745 1130
rect 4705 1100 4715 1120
rect 4735 1100 4745 1120
rect 4705 1090 4745 1100
rect 4785 1120 4825 1130
rect 4785 1100 4795 1120
rect 4815 1100 4825 1120
rect 4785 1090 4825 1100
rect 4865 1120 4905 1130
rect 4865 1100 4875 1120
rect 4895 1100 4905 1120
rect 4865 1090 4905 1100
rect 4945 1120 4985 1130
rect 4945 1100 4955 1120
rect 4975 1100 4985 1120
rect 4945 1090 4985 1100
rect 2985 1075 3985 1090
rect 4025 1075 5025 1090
rect 2985 960 3985 975
rect 4025 960 5025 975
rect 2995 925 3035 935
rect 2995 905 3005 925
rect 3025 905 3035 925
rect 4975 925 5015 935
rect 19315 1250 19320 1270
rect 19340 1250 19345 1270
rect 20010 1265 20105 1280
rect 20125 1265 20135 1285
rect 18745 1225 18760 1240
rect 18800 1235 19860 1250
rect 18800 1225 18815 1235
rect 18855 1225 18870 1235
rect 18910 1225 18925 1235
rect 18965 1225 18980 1235
rect 19020 1225 19035 1235
rect 19075 1225 19090 1235
rect 19130 1225 19145 1235
rect 19185 1225 19200 1235
rect 19240 1225 19255 1235
rect 19295 1225 19310 1235
rect 19350 1225 19365 1235
rect 19405 1225 19420 1235
rect 19460 1225 19475 1235
rect 19515 1225 19530 1235
rect 19570 1225 19585 1235
rect 19625 1225 19640 1235
rect 19680 1225 19695 1235
rect 19735 1225 19750 1235
rect 19790 1225 19805 1235
rect 19845 1225 19860 1235
rect 19900 1235 19970 1250
rect 19900 1225 19915 1235
rect 19955 1225 19970 1235
rect 20010 1225 20025 1265
rect 20095 1255 20135 1265
rect 20065 1225 20080 1240
rect 12965 980 13025 990
rect 12885 965 13025 980
rect 13065 975 13125 990
rect 13165 975 13225 990
rect 13265 975 13325 990
rect 13365 975 13425 990
rect 13465 975 13525 990
rect 13565 975 13625 990
rect 13665 975 13725 990
rect 13765 975 13825 990
rect 13865 975 13925 990
rect 13965 975 14025 990
rect 14065 980 14125 990
rect 14065 965 14205 980
rect 20585 1180 20600 1195
rect 20640 1180 20655 1195
rect 20695 1180 20710 1195
rect 20750 1180 20765 1195
rect 20585 1020 20600 1030
rect 20505 1005 20600 1020
rect 20640 1020 20655 1030
rect 20695 1020 20710 1030
rect 20640 1015 20710 1020
rect 20750 1020 20765 1030
rect 20640 1005 20725 1015
rect 20750 1005 20845 1020
rect 20505 985 20515 1005
rect 20535 985 20545 1005
rect 20505 975 20545 985
rect 20685 985 20695 1005
rect 20715 985 20725 1005
rect 20685 975 20725 985
rect 20805 985 20815 1005
rect 20835 985 20845 1005
rect 20805 975 20845 985
rect 12885 945 12895 965
rect 12915 945 12925 965
rect 12885 935 12925 945
rect 14165 945 14175 965
rect 14195 945 14205 965
rect 18745 960 18760 975
rect 18800 960 18815 975
rect 18855 960 18870 975
rect 18910 960 18925 975
rect 18965 960 18980 975
rect 19020 960 19035 975
rect 19075 960 19090 975
rect 19130 960 19145 975
rect 19185 960 19200 975
rect 19240 960 19255 975
rect 19295 960 19310 975
rect 19350 960 19365 975
rect 19405 960 19420 975
rect 19460 960 19475 975
rect 19515 960 19530 975
rect 19570 960 19585 975
rect 19625 960 19640 975
rect 19680 960 19695 975
rect 19735 960 19750 975
rect 19790 960 19805 975
rect 19845 960 19860 975
rect 19900 960 19915 975
rect 19955 960 19970 975
rect 20010 960 20025 975
rect 20065 960 20080 975
rect 14165 935 14205 945
rect 18665 950 18760 960
rect 18665 930 18675 950
rect 18695 945 18760 950
rect 20065 950 20160 960
rect 20065 945 20130 950
rect 18695 930 18705 945
rect 4975 905 4985 925
rect 5005 905 5015 925
rect 11245 910 11260 925
rect 11300 910 11315 925
rect 11355 910 11370 925
rect 11410 910 11425 925
rect 11465 910 11480 925
rect 11520 910 11535 925
rect 11575 910 11590 925
rect 11630 910 11645 925
rect 11685 910 11700 925
rect 11740 910 11755 925
rect 11795 910 11810 925
rect 11850 910 11865 925
rect 11905 910 11920 925
rect 11960 910 11975 925
rect 12015 910 12030 925
rect 12070 910 12085 925
rect 12125 910 12140 925
rect 12180 910 12195 925
rect 12235 910 12250 925
rect 12290 910 12305 925
rect 12345 910 12360 925
rect 12400 910 12415 925
rect 12455 910 12470 925
rect 12510 910 12525 925
rect 12565 910 12580 925
rect 18665 920 18705 930
rect 20120 930 20130 945
rect 20150 930 20160 950
rect 20120 920 20160 930
rect 2995 890 3085 905
rect 3035 880 3085 890
rect 3125 890 4885 905
rect 3125 880 3175 890
rect 3215 880 3265 890
rect 3305 880 3355 890
rect 3395 880 3445 890
rect 3485 880 3535 890
rect 3575 880 3625 890
rect 3665 880 3715 890
rect 3755 880 3805 890
rect 3845 880 3895 890
rect 3935 880 3985 890
rect 4025 880 4075 890
rect 4115 880 4165 890
rect 4205 880 4255 890
rect 4295 880 4345 890
rect 4385 880 4435 890
rect 4475 880 4525 890
rect 4565 880 4615 890
rect 4655 880 4705 890
rect 4745 880 4795 890
rect 4835 880 4885 890
rect 4925 890 5015 905
rect 11165 900 11260 910
rect 4925 880 4975 890
rect 11165 880 11175 900
rect 11195 895 11260 900
rect 12565 900 12660 910
rect 12565 895 12630 900
rect 11195 880 11205 895
rect 11165 870 11205 880
rect 12620 880 12630 895
rect 12650 880 12660 900
rect 12620 870 12660 880
rect 3035 765 3085 780
rect 3125 755 3175 780
rect 3215 765 3265 780
rect 3305 765 3355 780
rect 3395 765 3445 780
rect 3485 765 3535 780
rect 3575 765 3625 780
rect 3665 765 3715 780
rect 3755 765 3805 780
rect 3845 765 3895 780
rect 3935 765 3985 780
rect 4025 765 4075 780
rect 4115 765 4165 780
rect 4205 765 4255 780
rect 4295 765 4345 780
rect 4385 765 4435 780
rect 4475 765 4525 780
rect 4565 765 4615 780
rect 4655 765 4705 780
rect 4745 765 4795 780
rect 4835 765 4885 780
rect 4925 765 4975 780
rect 3125 750 3140 755
rect 3130 735 3140 750
rect 3160 750 3175 755
rect 3160 735 3170 750
rect 3130 725 3170 735
rect 9315 -730 9375 -715
rect 9415 -720 10375 -705
rect 9415 -730 9475 -720
rect 9515 -730 9575 -720
rect 9615 -730 9675 -720
rect 9715 -730 9775 -720
rect 9815 -730 9875 -720
rect 9915 -730 9975 -720
rect 10015 -730 10075 -720
rect 10115 -730 10175 -720
rect 10215 -730 10275 -720
rect 10315 -730 10375 -720
rect 10415 -730 10475 -715
rect 9315 -1020 9375 -1010
rect 9235 -1035 9375 -1020
rect 9415 -1025 9475 -1010
rect 9515 -1025 9575 -1010
rect 9615 -1025 9675 -1010
rect 9715 -1025 9775 -1010
rect 9815 -1025 9875 -1010
rect 9915 -1025 9975 -1010
rect 10015 -1025 10075 -1010
rect 10115 -1025 10175 -1010
rect 10215 -1025 10275 -1010
rect 10315 -1025 10375 -1010
rect 10415 -1020 10475 -1010
rect 10415 -1035 10555 -1020
rect 9235 -1055 9245 -1035
rect 9265 -1055 9275 -1035
rect 9235 -1065 9275 -1055
rect 10515 -1055 10525 -1035
rect 10545 -1055 10555 -1035
rect 10515 -1065 10555 -1055
<< polycont >>
rect 10915 3585 10935 3605
rect 11190 3600 11210 3620
rect 12590 3600 12610 3620
rect 10460 3320 10480 3340
rect 10720 3320 10740 3340
rect 18415 3585 18435 3605
rect 18690 3600 18710 3620
rect 20090 3600 20110 3620
rect 10590 3185 10610 3205
rect 10790 3185 10810 3205
rect 10910 3185 10930 3205
rect 10990 3185 11010 3205
rect 11110 3185 11130 3205
rect 17960 3320 17980 3340
rect 18220 3320 18240 3340
rect 11831 3130 11849 3150
rect 3145 2955 3165 2975
rect 4845 2955 4865 2975
rect 11190 2920 11210 2940
rect 18090 3185 18110 3205
rect 18290 3185 18310 3205
rect 18410 3185 18430 3205
rect 18490 3185 18510 3205
rect 18610 3185 18630 3205
rect 19331 3130 19349 3150
rect 12590 2920 12610 2940
rect 12860 2895 12880 2915
rect 3005 2785 3025 2805
rect 4985 2785 5005 2805
rect 3185 2725 3205 2745
rect 4805 2725 4825 2745
rect 13066 2895 13084 2915
rect 14150 2895 14170 2915
rect 18690 2920 18710 2940
rect 20090 2920 20110 2940
rect 20360 2895 20380 2915
rect 9650 2475 9670 2495
rect 10940 2475 10960 2495
rect 12860 2475 12880 2495
rect 11831 2450 11849 2470
rect 14150 2475 14170 2495
rect 20566 2895 20584 2915
rect 21650 2895 21670 2915
rect 17150 2475 17170 2495
rect 18440 2475 18460 2495
rect 20360 2475 20380 2495
rect 19331 2450 19349 2470
rect 10821 2415 10839 2435
rect 12981 2415 12999 2435
rect 21650 2475 21670 2495
rect 18321 2415 18339 2435
rect 20481 2415 20499 2435
rect 3365 2350 3385 2370
rect 3895 2355 3915 2375
rect 10821 2255 10839 2275
rect 12981 2255 12999 2275
rect 18321 2255 18339 2275
rect 20481 2255 20499 2275
rect 9650 2195 9670 2215
rect 10940 2195 10960 2215
rect 12860 2195 12880 2215
rect 14150 2195 14170 2215
rect 17150 2195 17170 2215
rect 18440 2195 18460 2215
rect 20360 2195 20380 2215
rect 21650 2195 21670 2215
rect 11245 1935 11265 1955
rect 12535 1935 12555 1955
rect 18745 1935 18765 1955
rect 20035 1935 20055 1955
rect 2630 1855 2650 1875
rect 2775 1855 2795 1875
rect 2845 1855 2865 1875
rect 2935 1855 2955 1875
rect 3175 1855 3195 1875
rect 3295 1855 3315 1875
rect 3535 1855 3555 1875
rect 3655 1855 3675 1875
rect 3865 1855 3885 1875
rect 3995 1850 4015 1870
rect 4125 1855 4145 1875
rect 4335 1855 4355 1875
rect 4455 1855 4475 1875
rect 4695 1855 4715 1875
rect 4815 1855 4835 1875
rect 5055 1855 5075 1875
rect 5145 1855 5165 1875
rect 5215 1855 5235 1875
rect 20460 1880 20480 1900
rect 20870 1880 20890 1900
rect 3235 1735 3255 1755
rect 4755 1735 4775 1755
rect 11243 1690 11260 1710
rect 11463 1690 11480 1710
rect 11610 1690 11627 1710
rect 11876 1690 11893 1710
rect 12283 1690 12300 1710
rect 12503 1690 12520 1710
rect 12650 1690 12667 1710
rect 18743 1690 18760 1710
rect 18963 1690 18980 1710
rect 19110 1690 19127 1710
rect 19376 1690 19393 1710
rect 19783 1690 19800 1710
rect 20003 1690 20020 1710
rect 20150 1690 20167 1710
rect 3175 1570 3195 1590
rect 4815 1570 4835 1590
rect 20571 1655 20591 1675
rect 20476 1545 20496 1565
rect 20854 1545 20874 1565
rect 2935 1475 2955 1495
rect 3055 1475 3075 1495
rect 3175 1475 3195 1495
rect 3295 1475 3315 1495
rect 3535 1475 3555 1495
rect 3655 1475 3675 1495
rect 3775 1475 3795 1495
rect 4215 1475 4235 1495
rect 4335 1475 4355 1495
rect 4455 1475 4475 1495
rect 4695 1475 4715 1495
rect 4815 1475 4835 1495
rect 4935 1475 4955 1495
rect 5055 1475 5075 1495
rect 11000 1470 11020 1490
rect 11112 1470 11129 1490
rect 11315 1470 11335 1490
rect 11535 1470 11555 1490
rect 11740 1470 11760 1490
rect 11928 1470 11945 1490
rect 12040 1470 12060 1490
rect 12152 1470 12169 1490
rect 12355 1470 12375 1490
rect 12575 1470 12595 1490
rect 12780 1470 12800 1490
rect 18500 1470 18520 1490
rect 18612 1470 18629 1490
rect 18815 1470 18835 1490
rect 19035 1470 19055 1490
rect 19240 1470 19260 1490
rect 19428 1470 19445 1490
rect 19540 1470 19560 1490
rect 19652 1470 19669 1490
rect 19855 1470 19875 1490
rect 20075 1470 20095 1490
rect 20280 1470 20300 1490
rect 20365 1325 20385 1345
rect 20533 1325 20553 1345
rect 20665 1325 20685 1345
rect 20797 1325 20817 1345
rect 20965 1325 20985 1345
rect 13136 1295 13154 1315
rect 11820 1200 11840 1220
rect 12605 1215 12625 1235
rect 3035 1100 3055 1120
rect 3115 1100 3135 1120
rect 3195 1100 3215 1120
rect 3275 1100 3295 1120
rect 3355 1100 3375 1120
rect 3435 1100 3455 1120
rect 3515 1100 3535 1120
rect 3595 1100 3615 1120
rect 3675 1100 3695 1120
rect 3755 1100 3775 1120
rect 3835 1100 3855 1120
rect 3915 1100 3935 1120
rect 4075 1100 4095 1120
rect 4155 1100 4175 1120
rect 4235 1100 4255 1120
rect 4315 1100 4335 1120
rect 4395 1100 4415 1120
rect 4475 1100 4495 1120
rect 4555 1100 4575 1120
rect 4635 1100 4655 1120
rect 4715 1100 4735 1120
rect 4795 1100 4815 1120
rect 4875 1100 4895 1120
rect 4955 1100 4975 1120
rect 3005 905 3025 925
rect 19320 1250 19340 1270
rect 20105 1265 20125 1285
rect 20515 985 20535 1005
rect 20695 985 20715 1005
rect 20815 985 20835 1005
rect 12895 945 12915 965
rect 14175 945 14195 965
rect 18675 930 18695 950
rect 4985 905 5005 925
rect 20130 930 20150 950
rect 11175 880 11195 900
rect 12630 880 12650 900
rect 3140 735 3160 755
rect 9245 -1055 9265 -1035
rect 10525 -1055 10545 -1035
<< xpolycontact >>
rect 91 3170 311 3205
rect 925 3170 1145 3205
rect 1306 3165 1526 3200
rect 2110 3165 2330 3200
rect 91 3110 311 3145
rect 925 3110 1145 3145
rect 1306 3105 1526 3140
rect 2110 3105 2330 3140
rect 91 3030 311 3065
rect 895 3030 1115 3065
rect 1306 3045 1526 3080
rect 2110 3045 2330 3080
rect 91 2970 311 3005
rect 895 2970 1115 3005
rect 1306 2985 1526 3020
rect 2110 2985 2330 3020
rect 1306 2925 1526 2960
rect 2110 2925 2330 2960
rect 1306 2865 1526 2900
rect 2110 2865 2330 2900
rect 96 2820 315 2855
rect 504 2820 724 2855
rect 1306 2805 1526 2840
rect 1740 2805 1960 2840
rect 96 2760 315 2795
rect 504 2760 724 2795
rect 13095 2695 13315 2836
rect 13455 2695 13675 2836
rect 20595 2695 20815 2836
rect 20955 2695 21175 2836
rect 9845 2345 10065 2380
rect 10415 2345 10635 2380
rect 13185 2345 13405 2380
rect 13755 2345 13975 2380
rect 17345 2345 17565 2380
rect 17915 2345 18135 2380
rect 20685 2345 20905 2380
rect 21255 2345 21475 2380
rect 9845 2285 10065 2320
rect 10415 2285 10635 2320
rect 13185 2285 13405 2320
rect 13755 2285 13975 2320
rect 17345 2285 17565 2320
rect 17915 2285 18135 2320
rect 20685 2285 20905 2320
rect 21255 2285 21475 2320
rect 13060 1395 13280 1430
rect 13805 1395 14025 1430
<< ppolyres >>
rect 315 2820 504 2855
rect 315 2760 504 2795
rect 13315 2695 13455 2836
rect 20815 2695 20955 2836
<< xpolyres >>
rect 311 3170 925 3205
rect 1526 3165 2110 3200
rect 311 3110 925 3145
rect 1526 3105 2110 3140
rect 311 3030 895 3065
rect 1526 3045 2110 3080
rect 311 2970 895 3005
rect 1526 2985 2110 3020
rect 1526 2925 2110 2960
rect 1526 2865 2110 2900
rect 1526 2805 1740 2840
rect 10065 2345 10415 2380
rect 13405 2345 13755 2380
rect 17565 2345 17915 2380
rect 20905 2345 21255 2380
rect 10065 2285 10415 2320
rect 13405 2285 13755 2320
rect 17565 2285 17915 2320
rect 20905 2285 21255 2320
rect 13280 1395 13805 1430
<< locali >>
rect 11180 3620 11220 3630
rect 10905 3605 11030 3615
rect 10905 3585 10915 3605
rect 10935 3595 11030 3605
rect 10935 3585 10945 3595
rect 10905 3575 10945 3585
rect 11010 3575 11030 3595
rect 11180 3600 11190 3620
rect 11210 3600 11220 3620
rect 11180 3590 11220 3600
rect 11340 3620 11380 3630
rect 11340 3600 11350 3620
rect 11370 3600 11380 3620
rect 11340 3590 11380 3600
rect 11460 3620 11500 3630
rect 11460 3600 11470 3620
rect 11490 3600 11500 3620
rect 11460 3590 11500 3600
rect 11580 3620 11620 3630
rect 11580 3600 11590 3620
rect 11610 3600 11620 3620
rect 11580 3590 11620 3600
rect 11700 3620 11740 3630
rect 11700 3600 11710 3620
rect 11730 3600 11740 3620
rect 11700 3590 11740 3600
rect 11820 3620 11860 3630
rect 11820 3600 11830 3620
rect 11850 3600 11860 3620
rect 11820 3590 11860 3600
rect 11940 3620 11980 3630
rect 11940 3600 11950 3620
rect 11970 3600 11980 3620
rect 11940 3590 11980 3600
rect 12060 3620 12100 3630
rect 12060 3600 12070 3620
rect 12090 3600 12100 3620
rect 12060 3590 12100 3600
rect 12180 3620 12220 3630
rect 12180 3600 12190 3620
rect 12210 3600 12220 3620
rect 12180 3590 12220 3600
rect 12300 3620 12340 3630
rect 12300 3600 12310 3620
rect 12330 3600 12340 3620
rect 12300 3590 12340 3600
rect 12420 3620 12460 3630
rect 12420 3600 12430 3620
rect 12450 3600 12460 3620
rect 12420 3590 12460 3600
rect 12580 3620 12620 3630
rect 12580 3600 12590 3620
rect 12610 3600 12620 3620
rect 18680 3620 18720 3630
rect 12580 3590 12620 3600
rect 18405 3605 18530 3615
rect 11005 3565 11035 3575
rect 11005 3545 11010 3565
rect 11030 3545 11035 3565
rect 1266 3495 1296 3525
rect 10785 3515 10855 3545
rect 10785 3495 10790 3515
rect 10810 3495 10830 3515
rect 10850 3495 10855 3515
rect 4445 3465 4475 3495
rect 10785 3465 10855 3495
rect -10 3415 20 3445
rect 945 3415 975 3445
rect 1645 3415 1675 3445
rect 2475 3420 2505 3450
rect 10785 3445 10790 3465
rect 10810 3445 10830 3465
rect 10850 3445 10855 3465
rect 5145 3415 5175 3445
rect 10785 3415 10855 3445
rect 10785 3395 10790 3415
rect 10810 3395 10830 3415
rect 10850 3395 10855 3415
rect -55 3360 -25 3390
rect 2695 3360 2725 3390
rect 10785 3365 10855 3395
rect 10450 3340 10490 3350
rect 1210 3310 1240 3340
rect 3140 3310 3170 3340
rect 3395 3305 3425 3335
rect 5365 3305 5395 3335
rect 10450 3320 10460 3340
rect 10480 3320 10490 3340
rect 10450 3310 10490 3320
rect 10710 3340 10750 3350
rect 10710 3320 10720 3340
rect 10740 3320 10750 3340
rect 10710 3310 10750 3320
rect 10785 3345 10790 3365
rect 10810 3345 10830 3365
rect 10850 3345 10855 3365
rect 10785 3315 10855 3345
rect 10460 3288 10480 3310
rect 10720 3288 10740 3310
rect 10785 3295 10790 3315
rect 10810 3295 10830 3315
rect 10850 3295 10855 3315
rect 1165 3255 1195 3285
rect 4890 3255 4920 3285
rect 5415 3255 5445 3285
rect 10455 3265 10525 3288
rect 10455 3245 10460 3265
rect 10480 3245 10500 3265
rect 10520 3245 10525 3265
rect 2740 3210 2770 3240
rect 10455 3235 10525 3245
rect 10555 3270 10585 3288
rect 10555 3250 10560 3270
rect 10580 3250 10585 3270
rect 10555 3235 10585 3250
rect 10615 3270 10645 3288
rect 10615 3250 10620 3270
rect 10640 3250 10645 3270
rect 10615 3235 10645 3250
rect 10675 3265 10745 3288
rect 10675 3245 10680 3265
rect 10700 3245 10720 3265
rect 10740 3245 10745 3265
rect 10675 3235 10745 3245
rect 10785 3265 10855 3295
rect 10785 3245 10790 3265
rect 10810 3245 10830 3265
rect 10850 3245 10855 3265
rect 10785 3235 10855 3245
rect 10885 3515 10915 3545
rect 10885 3495 10890 3515
rect 10910 3495 10915 3515
rect 10885 3465 10915 3495
rect 10885 3445 10890 3465
rect 10910 3445 10915 3465
rect 10885 3415 10915 3445
rect 10885 3395 10890 3415
rect 10910 3395 10915 3415
rect 10885 3365 10915 3395
rect 10885 3345 10890 3365
rect 10910 3345 10915 3365
rect 10885 3315 10915 3345
rect 10885 3295 10890 3315
rect 10910 3295 10915 3315
rect 10885 3265 10915 3295
rect 10885 3245 10890 3265
rect 10910 3245 10915 3265
rect 10885 3235 10915 3245
rect 10945 3515 10975 3545
rect 10945 3495 10950 3515
rect 10970 3495 10975 3515
rect 10945 3465 10975 3495
rect 10945 3445 10950 3465
rect 10970 3445 10975 3465
rect 10945 3415 10975 3445
rect 10945 3395 10950 3415
rect 10970 3395 10975 3415
rect 10945 3365 10975 3395
rect 10945 3345 10950 3365
rect 10970 3345 10975 3365
rect 10945 3315 10975 3345
rect 10945 3295 10950 3315
rect 10970 3295 10975 3315
rect 10945 3265 10975 3295
rect 10945 3245 10950 3265
rect 10970 3245 10975 3265
rect 10945 3235 10975 3245
rect 11005 3515 11035 3545
rect 11005 3495 11010 3515
rect 11030 3495 11035 3515
rect 11005 3465 11035 3495
rect 11005 3445 11010 3465
rect 11030 3445 11035 3465
rect 11005 3415 11035 3445
rect 11005 3395 11010 3415
rect 11030 3395 11035 3415
rect 11005 3365 11035 3395
rect 11005 3345 11010 3365
rect 11030 3345 11035 3365
rect 11005 3315 11035 3345
rect 11005 3295 11010 3315
rect 11030 3295 11035 3315
rect 11005 3265 11035 3295
rect 11005 3245 11010 3265
rect 11030 3245 11035 3265
rect 11005 3235 11035 3245
rect 11065 3565 11135 3575
rect 11190 3570 11210 3590
rect 11350 3570 11370 3590
rect 11470 3570 11490 3590
rect 11590 3570 11610 3590
rect 11710 3570 11730 3590
rect 11830 3570 11850 3590
rect 11950 3570 11970 3590
rect 12070 3570 12090 3590
rect 12190 3570 12210 3590
rect 12310 3570 12330 3590
rect 12430 3570 12450 3590
rect 12590 3570 12610 3590
rect 18405 3585 18415 3605
rect 18435 3595 18530 3605
rect 18435 3585 18445 3595
rect 18405 3575 18445 3585
rect 18510 3575 18530 3595
rect 18680 3600 18690 3620
rect 18710 3600 18720 3620
rect 18680 3590 18720 3600
rect 18840 3620 18880 3630
rect 18840 3600 18850 3620
rect 18870 3600 18880 3620
rect 18840 3590 18880 3600
rect 18960 3620 19000 3630
rect 18960 3600 18970 3620
rect 18990 3600 19000 3620
rect 18960 3590 19000 3600
rect 19080 3620 19120 3630
rect 19080 3600 19090 3620
rect 19110 3600 19120 3620
rect 19080 3590 19120 3600
rect 19200 3620 19240 3630
rect 19200 3600 19210 3620
rect 19230 3600 19240 3620
rect 19200 3590 19240 3600
rect 19320 3620 19360 3630
rect 19320 3600 19330 3620
rect 19350 3600 19360 3620
rect 19320 3590 19360 3600
rect 19440 3620 19480 3630
rect 19440 3600 19450 3620
rect 19470 3600 19480 3620
rect 19440 3590 19480 3600
rect 19560 3620 19600 3630
rect 19560 3600 19570 3620
rect 19590 3600 19600 3620
rect 19560 3590 19600 3600
rect 19680 3620 19720 3630
rect 19680 3600 19690 3620
rect 19710 3600 19720 3620
rect 19680 3590 19720 3600
rect 19800 3620 19840 3630
rect 19800 3600 19810 3620
rect 19830 3600 19840 3620
rect 19800 3590 19840 3600
rect 19920 3620 19960 3630
rect 19920 3600 19930 3620
rect 19950 3600 19960 3620
rect 19920 3590 19960 3600
rect 20080 3620 20120 3630
rect 20080 3600 20090 3620
rect 20110 3600 20120 3620
rect 20080 3590 20120 3600
rect 11065 3545 11070 3565
rect 11090 3545 11110 3565
rect 11130 3545 11135 3565
rect 11065 3515 11135 3545
rect 11065 3495 11070 3515
rect 11090 3495 11110 3515
rect 11130 3495 11135 3515
rect 11065 3465 11135 3495
rect 11065 3445 11070 3465
rect 11090 3445 11110 3465
rect 11130 3445 11135 3465
rect 11065 3415 11135 3445
rect 11065 3395 11070 3415
rect 11090 3395 11110 3415
rect 11130 3395 11135 3415
rect 11065 3365 11135 3395
rect 11065 3345 11070 3365
rect 11090 3345 11110 3365
rect 11130 3345 11135 3365
rect 11065 3315 11135 3345
rect 11065 3295 11070 3315
rect 11090 3295 11110 3315
rect 11130 3295 11135 3315
rect 11065 3265 11135 3295
rect 11065 3245 11070 3265
rect 11090 3245 11110 3265
rect 11130 3245 11135 3265
rect 11065 3235 11135 3245
rect 11185 3560 11255 3570
rect 11185 3540 11190 3560
rect 11210 3540 11230 3560
rect 11250 3540 11255 3560
rect 11185 3510 11255 3540
rect 11185 3490 11190 3510
rect 11210 3490 11230 3510
rect 11250 3490 11255 3510
rect 11185 3460 11255 3490
rect 11185 3440 11190 3460
rect 11210 3440 11230 3460
rect 11250 3440 11255 3460
rect 11185 3410 11255 3440
rect 11185 3390 11190 3410
rect 11210 3390 11230 3410
rect 11250 3390 11255 3410
rect 11185 3360 11255 3390
rect 11185 3340 11190 3360
rect 11210 3340 11230 3360
rect 11250 3340 11255 3360
rect 11185 3310 11255 3340
rect 11185 3290 11190 3310
rect 11210 3290 11230 3310
rect 11250 3290 11255 3310
rect 11185 3260 11255 3290
rect 11185 3240 11190 3260
rect 11210 3240 11230 3260
rect 11250 3240 11255 3260
rect 10620 3215 10640 3235
rect 10790 3215 10810 3235
rect 11110 3215 11130 3235
rect 10580 3205 10640 3215
rect 46 3200 91 3205
rect 46 3175 56 3200
rect 81 3175 91 3200
rect 46 3170 91 3175
rect 1110 3145 1145 3170
rect 1261 3195 1306 3200
rect 1261 3170 1271 3195
rect 1296 3170 1306 3195
rect 1261 3165 1306 3170
rect 2330 3165 2370 3200
rect 10580 3185 10590 3205
rect 10610 3195 10640 3205
rect 10780 3205 10820 3215
rect 10610 3185 10620 3195
rect 46 3140 91 3145
rect 46 3115 56 3140
rect 81 3115 91 3140
rect 46 3110 91 3115
rect 1261 3135 1306 3140
rect 1261 3110 1271 3135
rect 1296 3110 1306 3135
rect 1261 3105 1306 3110
rect 1165 3070 1195 3100
rect 2295 3080 2330 3105
rect 46 3060 91 3065
rect 46 3035 56 3060
rect 81 3035 91 3060
rect 46 3030 91 3035
rect 1080 3005 1115 3030
rect 46 3000 91 3005
rect 46 2975 56 3000
rect 81 2975 91 3000
rect 46 2970 91 2975
rect 1266 3045 1306 3080
rect 910 2910 1120 2915
rect 910 2880 920 2910
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1120 2910
rect 910 2875 1120 2880
rect 1266 2900 1286 3045
rect 2350 3020 2370 3165
rect 2625 3155 2655 3185
rect 4445 3155 4475 3185
rect 10580 3175 10620 3185
rect 10780 3185 10790 3205
rect 10810 3185 10820 3205
rect 10780 3175 10820 3185
rect 10905 3205 10940 3215
rect 10905 3185 10910 3205
rect 10930 3185 10940 3205
rect 10905 3175 10940 3185
rect 10980 3205 11015 3215
rect 10980 3185 10990 3205
rect 11010 3185 11015 3205
rect 10980 3175 11015 3185
rect 11100 3205 11140 3215
rect 11100 3185 11110 3205
rect 11130 3185 11140 3205
rect 11100 3175 11140 3185
rect 11185 3210 11255 3240
rect 11185 3190 11190 3210
rect 11210 3190 11230 3210
rect 11250 3190 11255 3210
rect 11185 3180 11255 3190
rect 11285 3560 11315 3570
rect 11285 3540 11290 3560
rect 11310 3540 11315 3560
rect 11285 3510 11315 3540
rect 11285 3490 11290 3510
rect 11310 3490 11315 3510
rect 11285 3460 11315 3490
rect 11285 3440 11290 3460
rect 11310 3440 11315 3460
rect 11285 3410 11315 3440
rect 11285 3390 11290 3410
rect 11310 3390 11315 3410
rect 11285 3360 11315 3390
rect 11285 3340 11290 3360
rect 11310 3340 11315 3360
rect 11285 3310 11315 3340
rect 11285 3290 11290 3310
rect 11310 3290 11315 3310
rect 11285 3260 11315 3290
rect 11285 3240 11290 3260
rect 11310 3240 11315 3260
rect 11285 3210 11315 3240
rect 11285 3190 11290 3210
rect 11310 3190 11315 3210
rect 11285 3180 11315 3190
rect 11345 3560 11375 3570
rect 11345 3540 11350 3560
rect 11370 3540 11375 3560
rect 11345 3510 11375 3540
rect 11345 3490 11350 3510
rect 11370 3490 11375 3510
rect 11345 3460 11375 3490
rect 11345 3440 11350 3460
rect 11370 3440 11375 3460
rect 11345 3410 11375 3440
rect 11345 3390 11350 3410
rect 11370 3390 11375 3410
rect 11345 3360 11375 3390
rect 11345 3340 11350 3360
rect 11370 3340 11375 3360
rect 11345 3310 11375 3340
rect 11345 3290 11350 3310
rect 11370 3290 11375 3310
rect 11345 3260 11375 3290
rect 11345 3240 11350 3260
rect 11370 3240 11375 3260
rect 11345 3210 11375 3240
rect 11345 3190 11350 3210
rect 11370 3190 11375 3210
rect 11345 3180 11375 3190
rect 11405 3560 11435 3570
rect 11405 3540 11410 3560
rect 11430 3540 11435 3560
rect 11405 3510 11435 3540
rect 11405 3490 11410 3510
rect 11430 3490 11435 3510
rect 11405 3460 11435 3490
rect 11405 3440 11410 3460
rect 11430 3440 11435 3460
rect 11405 3410 11435 3440
rect 11405 3390 11410 3410
rect 11430 3390 11435 3410
rect 11405 3360 11435 3390
rect 11405 3340 11410 3360
rect 11430 3340 11435 3360
rect 11405 3310 11435 3340
rect 11405 3290 11410 3310
rect 11430 3290 11435 3310
rect 11405 3260 11435 3290
rect 11405 3240 11410 3260
rect 11430 3240 11435 3260
rect 11405 3210 11435 3240
rect 11405 3190 11410 3210
rect 11430 3190 11435 3210
rect 11405 3180 11435 3190
rect 11465 3560 11495 3570
rect 11465 3540 11470 3560
rect 11490 3540 11495 3560
rect 11465 3510 11495 3540
rect 11465 3490 11470 3510
rect 11490 3490 11495 3510
rect 11465 3460 11495 3490
rect 11465 3440 11470 3460
rect 11490 3440 11495 3460
rect 11465 3410 11495 3440
rect 11465 3390 11470 3410
rect 11490 3390 11495 3410
rect 11465 3360 11495 3390
rect 11465 3340 11470 3360
rect 11490 3340 11495 3360
rect 11465 3310 11495 3340
rect 11465 3290 11470 3310
rect 11490 3290 11495 3310
rect 11465 3260 11495 3290
rect 11465 3240 11470 3260
rect 11490 3240 11495 3260
rect 11465 3210 11495 3240
rect 11465 3190 11470 3210
rect 11490 3190 11495 3210
rect 11465 3180 11495 3190
rect 11525 3560 11555 3570
rect 11525 3540 11530 3560
rect 11550 3540 11555 3560
rect 11525 3510 11555 3540
rect 11525 3490 11530 3510
rect 11550 3490 11555 3510
rect 11525 3460 11555 3490
rect 11525 3440 11530 3460
rect 11550 3440 11555 3460
rect 11525 3410 11555 3440
rect 11525 3390 11530 3410
rect 11550 3390 11555 3410
rect 11525 3360 11555 3390
rect 11525 3340 11530 3360
rect 11550 3340 11555 3360
rect 11525 3310 11555 3340
rect 11525 3290 11530 3310
rect 11550 3290 11555 3310
rect 11525 3260 11555 3290
rect 11525 3240 11530 3260
rect 11550 3240 11555 3260
rect 11525 3210 11555 3240
rect 11525 3190 11530 3210
rect 11550 3190 11555 3210
rect 11525 3180 11555 3190
rect 11585 3560 11615 3570
rect 11585 3540 11590 3560
rect 11610 3540 11615 3560
rect 11585 3510 11615 3540
rect 11585 3490 11590 3510
rect 11610 3490 11615 3510
rect 11585 3460 11615 3490
rect 11585 3440 11590 3460
rect 11610 3440 11615 3460
rect 11585 3410 11615 3440
rect 11585 3390 11590 3410
rect 11610 3390 11615 3410
rect 11585 3360 11615 3390
rect 11585 3340 11590 3360
rect 11610 3340 11615 3360
rect 11585 3310 11615 3340
rect 11585 3290 11590 3310
rect 11610 3290 11615 3310
rect 11585 3260 11615 3290
rect 11585 3240 11590 3260
rect 11610 3240 11615 3260
rect 11585 3210 11615 3240
rect 11585 3190 11590 3210
rect 11610 3190 11615 3210
rect 11585 3180 11615 3190
rect 11645 3560 11675 3570
rect 11645 3540 11650 3560
rect 11670 3540 11675 3560
rect 11645 3510 11675 3540
rect 11645 3490 11650 3510
rect 11670 3490 11675 3510
rect 11645 3460 11675 3490
rect 11645 3440 11650 3460
rect 11670 3440 11675 3460
rect 11645 3410 11675 3440
rect 11645 3390 11650 3410
rect 11670 3390 11675 3410
rect 11645 3360 11675 3390
rect 11645 3340 11650 3360
rect 11670 3340 11675 3360
rect 11645 3310 11675 3340
rect 11645 3290 11650 3310
rect 11670 3290 11675 3310
rect 11645 3260 11675 3290
rect 11645 3240 11650 3260
rect 11670 3240 11675 3260
rect 11645 3210 11675 3240
rect 11645 3190 11650 3210
rect 11670 3190 11675 3210
rect 11645 3180 11675 3190
rect 11705 3560 11735 3570
rect 11705 3540 11710 3560
rect 11730 3540 11735 3560
rect 11705 3510 11735 3540
rect 11705 3490 11710 3510
rect 11730 3490 11735 3510
rect 11705 3460 11735 3490
rect 11705 3440 11710 3460
rect 11730 3440 11735 3460
rect 11705 3410 11735 3440
rect 11705 3390 11710 3410
rect 11730 3390 11735 3410
rect 11705 3360 11735 3390
rect 11705 3340 11710 3360
rect 11730 3340 11735 3360
rect 11705 3310 11735 3340
rect 11705 3290 11710 3310
rect 11730 3290 11735 3310
rect 11705 3260 11735 3290
rect 11705 3240 11710 3260
rect 11730 3240 11735 3260
rect 11705 3210 11735 3240
rect 11705 3190 11710 3210
rect 11730 3190 11735 3210
rect 11705 3180 11735 3190
rect 11765 3560 11795 3570
rect 11765 3540 11770 3560
rect 11790 3540 11795 3560
rect 11765 3510 11795 3540
rect 11765 3490 11770 3510
rect 11790 3490 11795 3510
rect 11765 3460 11795 3490
rect 11765 3440 11770 3460
rect 11790 3440 11795 3460
rect 11765 3410 11795 3440
rect 11765 3390 11770 3410
rect 11790 3390 11795 3410
rect 11765 3360 11795 3390
rect 11765 3340 11770 3360
rect 11790 3340 11795 3360
rect 11765 3310 11795 3340
rect 11765 3290 11770 3310
rect 11790 3290 11795 3310
rect 11765 3260 11795 3290
rect 11765 3240 11770 3260
rect 11790 3240 11795 3260
rect 11765 3210 11795 3240
rect 11765 3190 11770 3210
rect 11790 3190 11795 3210
rect 11765 3180 11795 3190
rect 11825 3560 11855 3570
rect 11825 3540 11830 3560
rect 11850 3540 11855 3560
rect 11825 3510 11855 3540
rect 11825 3490 11830 3510
rect 11850 3490 11855 3510
rect 11825 3460 11855 3490
rect 11825 3440 11830 3460
rect 11850 3440 11855 3460
rect 11825 3410 11855 3440
rect 11825 3390 11830 3410
rect 11850 3390 11855 3410
rect 11825 3360 11855 3390
rect 11825 3340 11830 3360
rect 11850 3340 11855 3360
rect 11825 3310 11855 3340
rect 11825 3290 11830 3310
rect 11850 3290 11855 3310
rect 11825 3260 11855 3290
rect 11825 3240 11830 3260
rect 11850 3240 11855 3260
rect 11825 3210 11855 3240
rect 11825 3190 11830 3210
rect 11850 3190 11855 3210
rect 11825 3180 11855 3190
rect 11885 3560 11915 3570
rect 11885 3540 11890 3560
rect 11910 3540 11915 3560
rect 11885 3510 11915 3540
rect 11885 3490 11890 3510
rect 11910 3490 11915 3510
rect 11885 3460 11915 3490
rect 11885 3440 11890 3460
rect 11910 3440 11915 3460
rect 11885 3410 11915 3440
rect 11885 3390 11890 3410
rect 11910 3390 11915 3410
rect 11885 3360 11915 3390
rect 11885 3340 11890 3360
rect 11910 3340 11915 3360
rect 11885 3310 11915 3340
rect 11885 3290 11890 3310
rect 11910 3290 11915 3310
rect 11885 3260 11915 3290
rect 11885 3240 11890 3260
rect 11910 3240 11915 3260
rect 11885 3210 11915 3240
rect 11885 3190 11890 3210
rect 11910 3190 11915 3210
rect 11885 3180 11915 3190
rect 11945 3560 11975 3570
rect 11945 3540 11950 3560
rect 11970 3540 11975 3560
rect 11945 3510 11975 3540
rect 11945 3490 11950 3510
rect 11970 3490 11975 3510
rect 11945 3460 11975 3490
rect 11945 3440 11950 3460
rect 11970 3440 11975 3460
rect 11945 3410 11975 3440
rect 11945 3390 11950 3410
rect 11970 3390 11975 3410
rect 11945 3360 11975 3390
rect 11945 3340 11950 3360
rect 11970 3340 11975 3360
rect 11945 3310 11975 3340
rect 11945 3290 11950 3310
rect 11970 3290 11975 3310
rect 11945 3260 11975 3290
rect 11945 3240 11950 3260
rect 11970 3240 11975 3260
rect 11945 3210 11975 3240
rect 11945 3190 11950 3210
rect 11970 3190 11975 3210
rect 11945 3180 11975 3190
rect 12005 3560 12035 3570
rect 12005 3540 12010 3560
rect 12030 3540 12035 3560
rect 12005 3510 12035 3540
rect 12005 3490 12010 3510
rect 12030 3490 12035 3510
rect 12005 3460 12035 3490
rect 12005 3440 12010 3460
rect 12030 3440 12035 3460
rect 12005 3410 12035 3440
rect 12005 3390 12010 3410
rect 12030 3390 12035 3410
rect 12005 3360 12035 3390
rect 12005 3340 12010 3360
rect 12030 3340 12035 3360
rect 12005 3310 12035 3340
rect 12005 3290 12010 3310
rect 12030 3290 12035 3310
rect 12005 3260 12035 3290
rect 12005 3240 12010 3260
rect 12030 3240 12035 3260
rect 12005 3210 12035 3240
rect 12005 3190 12010 3210
rect 12030 3190 12035 3210
rect 12005 3180 12035 3190
rect 12065 3560 12095 3570
rect 12065 3540 12070 3560
rect 12090 3540 12095 3560
rect 12065 3510 12095 3540
rect 12065 3490 12070 3510
rect 12090 3490 12095 3510
rect 12065 3460 12095 3490
rect 12065 3440 12070 3460
rect 12090 3440 12095 3460
rect 12065 3410 12095 3440
rect 12065 3390 12070 3410
rect 12090 3390 12095 3410
rect 12065 3360 12095 3390
rect 12065 3340 12070 3360
rect 12090 3340 12095 3360
rect 12065 3310 12095 3340
rect 12065 3290 12070 3310
rect 12090 3290 12095 3310
rect 12065 3260 12095 3290
rect 12065 3240 12070 3260
rect 12090 3240 12095 3260
rect 12065 3210 12095 3240
rect 12065 3190 12070 3210
rect 12090 3190 12095 3210
rect 12065 3180 12095 3190
rect 12125 3560 12155 3570
rect 12125 3540 12130 3560
rect 12150 3540 12155 3560
rect 12125 3510 12155 3540
rect 12125 3490 12130 3510
rect 12150 3490 12155 3510
rect 12125 3460 12155 3490
rect 12125 3440 12130 3460
rect 12150 3440 12155 3460
rect 12125 3410 12155 3440
rect 12125 3390 12130 3410
rect 12150 3390 12155 3410
rect 12125 3360 12155 3390
rect 12125 3340 12130 3360
rect 12150 3340 12155 3360
rect 12125 3310 12155 3340
rect 12125 3290 12130 3310
rect 12150 3290 12155 3310
rect 12125 3260 12155 3290
rect 12125 3240 12130 3260
rect 12150 3240 12155 3260
rect 12125 3210 12155 3240
rect 12125 3190 12130 3210
rect 12150 3190 12155 3210
rect 12125 3180 12155 3190
rect 12185 3560 12215 3570
rect 12185 3540 12190 3560
rect 12210 3540 12215 3560
rect 12185 3510 12215 3540
rect 12185 3490 12190 3510
rect 12210 3490 12215 3510
rect 12185 3460 12215 3490
rect 12185 3440 12190 3460
rect 12210 3440 12215 3460
rect 12185 3410 12215 3440
rect 12185 3390 12190 3410
rect 12210 3390 12215 3410
rect 12185 3360 12215 3390
rect 12185 3340 12190 3360
rect 12210 3340 12215 3360
rect 12185 3310 12215 3340
rect 12185 3290 12190 3310
rect 12210 3290 12215 3310
rect 12185 3260 12215 3290
rect 12185 3240 12190 3260
rect 12210 3240 12215 3260
rect 12185 3210 12215 3240
rect 12185 3190 12190 3210
rect 12210 3190 12215 3210
rect 12185 3180 12215 3190
rect 12245 3560 12275 3570
rect 12245 3540 12250 3560
rect 12270 3540 12275 3560
rect 12245 3510 12275 3540
rect 12245 3490 12250 3510
rect 12270 3490 12275 3510
rect 12245 3460 12275 3490
rect 12245 3440 12250 3460
rect 12270 3440 12275 3460
rect 12245 3410 12275 3440
rect 12245 3390 12250 3410
rect 12270 3390 12275 3410
rect 12245 3360 12275 3390
rect 12245 3340 12250 3360
rect 12270 3340 12275 3360
rect 12245 3310 12275 3340
rect 12245 3290 12250 3310
rect 12270 3290 12275 3310
rect 12245 3260 12275 3290
rect 12245 3240 12250 3260
rect 12270 3240 12275 3260
rect 12245 3210 12275 3240
rect 12245 3190 12250 3210
rect 12270 3190 12275 3210
rect 12245 3180 12275 3190
rect 12305 3560 12335 3570
rect 12305 3540 12310 3560
rect 12330 3540 12335 3560
rect 12305 3510 12335 3540
rect 12305 3490 12310 3510
rect 12330 3490 12335 3510
rect 12305 3460 12335 3490
rect 12305 3440 12310 3460
rect 12330 3440 12335 3460
rect 12305 3410 12335 3440
rect 12305 3390 12310 3410
rect 12330 3390 12335 3410
rect 12305 3360 12335 3390
rect 12305 3340 12310 3360
rect 12330 3340 12335 3360
rect 12305 3310 12335 3340
rect 12305 3290 12310 3310
rect 12330 3290 12335 3310
rect 12305 3260 12335 3290
rect 12305 3240 12310 3260
rect 12330 3240 12335 3260
rect 12305 3210 12335 3240
rect 12305 3190 12310 3210
rect 12330 3190 12335 3210
rect 12305 3180 12335 3190
rect 12365 3560 12395 3570
rect 12365 3540 12370 3560
rect 12390 3540 12395 3560
rect 12365 3510 12395 3540
rect 12365 3490 12370 3510
rect 12390 3490 12395 3510
rect 12365 3460 12395 3490
rect 12365 3440 12370 3460
rect 12390 3440 12395 3460
rect 12365 3410 12395 3440
rect 12365 3390 12370 3410
rect 12390 3390 12395 3410
rect 12365 3360 12395 3390
rect 12365 3340 12370 3360
rect 12390 3340 12395 3360
rect 12365 3310 12395 3340
rect 12365 3290 12370 3310
rect 12390 3290 12395 3310
rect 12365 3260 12395 3290
rect 12365 3240 12370 3260
rect 12390 3240 12395 3260
rect 12365 3210 12395 3240
rect 12365 3190 12370 3210
rect 12390 3190 12395 3210
rect 12365 3180 12395 3190
rect 12425 3560 12455 3570
rect 12425 3540 12430 3560
rect 12450 3540 12455 3560
rect 12425 3510 12455 3540
rect 12425 3490 12430 3510
rect 12450 3490 12455 3510
rect 12425 3460 12455 3490
rect 12425 3440 12430 3460
rect 12450 3440 12455 3460
rect 12425 3410 12455 3440
rect 12425 3390 12430 3410
rect 12450 3390 12455 3410
rect 12425 3360 12455 3390
rect 12425 3340 12430 3360
rect 12450 3340 12455 3360
rect 12425 3310 12455 3340
rect 12425 3290 12430 3310
rect 12450 3290 12455 3310
rect 12425 3260 12455 3290
rect 12425 3240 12430 3260
rect 12450 3240 12455 3260
rect 12425 3210 12455 3240
rect 12425 3190 12430 3210
rect 12450 3190 12455 3210
rect 12425 3180 12455 3190
rect 12485 3560 12515 3570
rect 12485 3540 12490 3560
rect 12510 3540 12515 3560
rect 12485 3510 12515 3540
rect 12485 3490 12490 3510
rect 12510 3490 12515 3510
rect 12485 3460 12515 3490
rect 12485 3440 12490 3460
rect 12510 3440 12515 3460
rect 12485 3410 12515 3440
rect 12485 3390 12490 3410
rect 12510 3390 12515 3410
rect 12485 3360 12515 3390
rect 12485 3340 12490 3360
rect 12510 3340 12515 3360
rect 12485 3310 12515 3340
rect 12485 3290 12490 3310
rect 12510 3290 12515 3310
rect 12485 3260 12515 3290
rect 12485 3240 12490 3260
rect 12510 3240 12515 3260
rect 12485 3210 12515 3240
rect 12485 3190 12490 3210
rect 12510 3190 12515 3210
rect 12485 3180 12515 3190
rect 12545 3560 12615 3570
rect 12545 3540 12550 3560
rect 12570 3540 12590 3560
rect 12610 3540 12615 3560
rect 18505 3565 18535 3575
rect 18505 3545 18510 3565
rect 18530 3545 18535 3565
rect 12545 3510 12615 3540
rect 12545 3490 12550 3510
rect 12570 3490 12590 3510
rect 12610 3490 12615 3510
rect 12545 3460 12615 3490
rect 12545 3440 12550 3460
rect 12570 3440 12590 3460
rect 12610 3440 12615 3460
rect 12545 3410 12615 3440
rect 12545 3390 12550 3410
rect 12570 3390 12590 3410
rect 12610 3390 12615 3410
rect 12545 3360 12615 3390
rect 12545 3340 12550 3360
rect 12570 3340 12590 3360
rect 12610 3340 12615 3360
rect 18285 3515 18355 3545
rect 18285 3495 18290 3515
rect 18310 3495 18330 3515
rect 18350 3495 18355 3515
rect 18285 3465 18355 3495
rect 18285 3445 18290 3465
rect 18310 3445 18330 3465
rect 18350 3445 18355 3465
rect 18285 3415 18355 3445
rect 18285 3395 18290 3415
rect 18310 3395 18330 3415
rect 18350 3395 18355 3415
rect 18285 3365 18355 3395
rect 12545 3310 12615 3340
rect 17950 3340 17990 3350
rect 17950 3320 17960 3340
rect 17980 3320 17990 3340
rect 17950 3310 17990 3320
rect 18210 3340 18250 3350
rect 18210 3320 18220 3340
rect 18240 3320 18250 3340
rect 18210 3310 18250 3320
rect 18285 3345 18290 3365
rect 18310 3345 18330 3365
rect 18350 3345 18355 3365
rect 18285 3315 18355 3345
rect 12545 3290 12550 3310
rect 12570 3290 12590 3310
rect 12610 3290 12615 3310
rect 12545 3260 12615 3290
rect 12545 3240 12550 3260
rect 12570 3240 12590 3260
rect 12610 3240 12615 3260
rect 12945 3285 12985 3295
rect 12945 3265 12955 3285
rect 12975 3265 12985 3285
rect 12945 3255 12985 3265
rect 13055 3285 13095 3295
rect 13055 3265 13065 3285
rect 13085 3265 13095 3285
rect 13055 3255 13095 3265
rect 13165 3285 13205 3295
rect 13165 3265 13175 3285
rect 13195 3265 13205 3285
rect 13165 3255 13205 3265
rect 13275 3285 13315 3295
rect 13275 3265 13285 3285
rect 13305 3265 13315 3285
rect 13275 3255 13315 3265
rect 13385 3285 13425 3295
rect 13385 3265 13395 3285
rect 13415 3265 13425 3285
rect 13385 3255 13425 3265
rect 13495 3285 13535 3295
rect 13495 3265 13505 3285
rect 13525 3265 13535 3285
rect 13495 3255 13535 3265
rect 13605 3285 13645 3295
rect 13605 3265 13615 3285
rect 13635 3265 13645 3285
rect 13605 3255 13645 3265
rect 13715 3285 13755 3295
rect 13715 3265 13725 3285
rect 13745 3265 13755 3285
rect 13715 3255 13755 3265
rect 13825 3285 13865 3295
rect 13825 3265 13835 3285
rect 13855 3265 13865 3285
rect 13825 3255 13865 3265
rect 13935 3285 13975 3295
rect 13935 3265 13945 3285
rect 13965 3265 13975 3285
rect 13935 3255 13975 3265
rect 14045 3285 14085 3295
rect 17960 3288 17980 3310
rect 18220 3288 18240 3310
rect 18285 3295 18290 3315
rect 18310 3295 18330 3315
rect 18350 3295 18355 3315
rect 14045 3265 14055 3285
rect 14075 3265 14085 3285
rect 14045 3255 14085 3265
rect 17955 3265 18025 3288
rect 12545 3210 12615 3240
rect 12955 3235 12975 3255
rect 13065 3235 13085 3255
rect 13175 3235 13195 3255
rect 13285 3235 13305 3255
rect 13395 3235 13415 3255
rect 13505 3235 13525 3255
rect 13615 3235 13635 3255
rect 13725 3235 13745 3255
rect 13835 3235 13855 3255
rect 13945 3235 13965 3255
rect 14055 3235 14075 3255
rect 17955 3245 17960 3265
rect 17980 3245 18000 3265
rect 18020 3245 18025 3265
rect 17955 3235 18025 3245
rect 18055 3270 18085 3288
rect 18055 3250 18060 3270
rect 18080 3250 18085 3270
rect 18055 3235 18085 3250
rect 18115 3270 18145 3288
rect 18115 3250 18120 3270
rect 18140 3250 18145 3270
rect 18115 3235 18145 3250
rect 18175 3265 18245 3288
rect 18175 3245 18180 3265
rect 18200 3245 18220 3265
rect 18240 3245 18245 3265
rect 18175 3235 18245 3245
rect 18285 3265 18355 3295
rect 18285 3245 18290 3265
rect 18310 3245 18330 3265
rect 18350 3245 18355 3265
rect 18285 3235 18355 3245
rect 18385 3515 18415 3545
rect 18385 3495 18390 3515
rect 18410 3495 18415 3515
rect 18385 3465 18415 3495
rect 18385 3445 18390 3465
rect 18410 3445 18415 3465
rect 18385 3415 18415 3445
rect 18385 3395 18390 3415
rect 18410 3395 18415 3415
rect 18385 3365 18415 3395
rect 18385 3345 18390 3365
rect 18410 3345 18415 3365
rect 18385 3315 18415 3345
rect 18385 3295 18390 3315
rect 18410 3295 18415 3315
rect 18385 3265 18415 3295
rect 18385 3245 18390 3265
rect 18410 3245 18415 3265
rect 18385 3235 18415 3245
rect 18445 3515 18475 3545
rect 18445 3495 18450 3515
rect 18470 3495 18475 3515
rect 18445 3465 18475 3495
rect 18445 3445 18450 3465
rect 18470 3445 18475 3465
rect 18445 3415 18475 3445
rect 18445 3395 18450 3415
rect 18470 3395 18475 3415
rect 18445 3365 18475 3395
rect 18445 3345 18450 3365
rect 18470 3345 18475 3365
rect 18445 3315 18475 3345
rect 18445 3295 18450 3315
rect 18470 3295 18475 3315
rect 18445 3265 18475 3295
rect 18445 3245 18450 3265
rect 18470 3245 18475 3265
rect 18445 3235 18475 3245
rect 18505 3515 18535 3545
rect 18505 3495 18510 3515
rect 18530 3495 18535 3515
rect 18505 3465 18535 3495
rect 18505 3445 18510 3465
rect 18530 3445 18535 3465
rect 18505 3415 18535 3445
rect 18505 3395 18510 3415
rect 18530 3395 18535 3415
rect 18505 3365 18535 3395
rect 18505 3345 18510 3365
rect 18530 3345 18535 3365
rect 18505 3315 18535 3345
rect 18505 3295 18510 3315
rect 18530 3295 18535 3315
rect 18505 3265 18535 3295
rect 18505 3245 18510 3265
rect 18530 3245 18535 3265
rect 18505 3235 18535 3245
rect 18565 3565 18635 3575
rect 18690 3570 18710 3590
rect 18850 3570 18870 3590
rect 18970 3570 18990 3590
rect 19090 3570 19110 3590
rect 19210 3570 19230 3590
rect 19330 3570 19350 3590
rect 19450 3570 19470 3590
rect 19570 3570 19590 3590
rect 19690 3570 19710 3590
rect 19810 3570 19830 3590
rect 19930 3570 19950 3590
rect 20090 3570 20110 3590
rect 18565 3545 18570 3565
rect 18590 3545 18610 3565
rect 18630 3545 18635 3565
rect 18565 3515 18635 3545
rect 18565 3495 18570 3515
rect 18590 3495 18610 3515
rect 18630 3495 18635 3515
rect 18565 3465 18635 3495
rect 18565 3445 18570 3465
rect 18590 3445 18610 3465
rect 18630 3445 18635 3465
rect 18565 3415 18635 3445
rect 18565 3395 18570 3415
rect 18590 3395 18610 3415
rect 18630 3395 18635 3415
rect 18565 3365 18635 3395
rect 18565 3345 18570 3365
rect 18590 3345 18610 3365
rect 18630 3345 18635 3365
rect 18565 3315 18635 3345
rect 18565 3295 18570 3315
rect 18590 3295 18610 3315
rect 18630 3295 18635 3315
rect 18565 3265 18635 3295
rect 18565 3245 18570 3265
rect 18590 3245 18610 3265
rect 18630 3245 18635 3265
rect 18565 3235 18635 3245
rect 18685 3560 18755 3570
rect 18685 3540 18690 3560
rect 18710 3540 18730 3560
rect 18750 3540 18755 3560
rect 18685 3510 18755 3540
rect 18685 3490 18690 3510
rect 18710 3490 18730 3510
rect 18750 3490 18755 3510
rect 18685 3460 18755 3490
rect 18685 3440 18690 3460
rect 18710 3440 18730 3460
rect 18750 3440 18755 3460
rect 18685 3410 18755 3440
rect 18685 3390 18690 3410
rect 18710 3390 18730 3410
rect 18750 3390 18755 3410
rect 18685 3360 18755 3390
rect 18685 3340 18690 3360
rect 18710 3340 18730 3360
rect 18750 3340 18755 3360
rect 18685 3310 18755 3340
rect 18685 3290 18690 3310
rect 18710 3290 18730 3310
rect 18750 3290 18755 3310
rect 18685 3260 18755 3290
rect 18685 3240 18690 3260
rect 18710 3240 18730 3260
rect 18750 3240 18755 3260
rect 12545 3190 12550 3210
rect 12570 3190 12590 3210
rect 12610 3190 12615 3210
rect 12545 3180 12615 3190
rect 12855 3225 12925 3235
rect 12855 3205 12860 3225
rect 12880 3205 12900 3225
rect 12920 3205 12925 3225
rect 11290 3160 11310 3180
rect 11410 3160 11430 3180
rect 11530 3160 11550 3180
rect 11650 3160 11670 3180
rect 11770 3160 11790 3180
rect 11890 3160 11910 3180
rect 12010 3160 12030 3180
rect 12130 3160 12150 3180
rect 12250 3160 12270 3180
rect 12370 3160 12390 3180
rect 12490 3160 12510 3180
rect 12855 3175 12925 3205
rect 11280 3150 11320 3160
rect 3140 3110 3170 3140
rect 4840 3110 4870 3140
rect 5320 3110 5350 3140
rect 11280 3130 11290 3150
rect 11310 3130 11320 3150
rect 11280 3120 11320 3130
rect 11400 3150 11440 3160
rect 11400 3130 11410 3150
rect 11430 3130 11440 3150
rect 11400 3120 11440 3130
rect 11520 3150 11560 3160
rect 11520 3130 11530 3150
rect 11550 3130 11560 3150
rect 11520 3120 11560 3130
rect 11640 3150 11680 3160
rect 11640 3130 11650 3150
rect 11670 3130 11680 3150
rect 11640 3120 11680 3130
rect 11760 3150 11800 3160
rect 11760 3130 11770 3150
rect 11790 3130 11800 3150
rect 11760 3120 11800 3130
rect 11823 3150 11857 3160
rect 11823 3130 11831 3150
rect 11849 3130 11857 3150
rect 11823 3120 11857 3130
rect 11880 3150 11920 3160
rect 11880 3130 11890 3150
rect 11910 3130 11920 3150
rect 11880 3120 11920 3130
rect 12000 3150 12040 3160
rect 12000 3130 12010 3150
rect 12030 3130 12040 3150
rect 12000 3120 12040 3130
rect 12120 3150 12160 3160
rect 12120 3130 12130 3150
rect 12150 3130 12160 3150
rect 12120 3120 12160 3130
rect 12240 3150 12280 3160
rect 12240 3130 12250 3150
rect 12270 3130 12280 3150
rect 12240 3120 12280 3130
rect 12360 3150 12400 3160
rect 12360 3130 12370 3150
rect 12390 3130 12400 3150
rect 12360 3120 12400 3130
rect 12480 3150 12520 3160
rect 12480 3130 12490 3150
rect 12510 3130 12520 3150
rect 12480 3120 12520 3130
rect 12855 3155 12860 3175
rect 12880 3155 12900 3175
rect 12920 3155 12925 3175
rect 12855 3125 12925 3155
rect 12855 3105 12860 3125
rect 12880 3105 12900 3125
rect 12920 3105 12925 3125
rect 3990 3050 4020 3080
rect 12855 3075 12925 3105
rect 12855 3055 12860 3075
rect 12880 3055 12900 3075
rect 12920 3055 12925 3075
rect 2330 2985 2370 3020
rect 3450 3005 3480 3035
rect 3810 3005 3840 3035
rect 4350 3005 4380 3035
rect 4710 3005 4740 3035
rect 12855 3025 12925 3055
rect 12855 3005 12860 3025
rect 12880 3005 12900 3025
rect 12920 3005 12925 3025
rect 1306 2960 1341 2985
rect 2330 2955 2375 2960
rect 2330 2930 2340 2955
rect 2365 2930 2375 2955
rect 2330 2925 2375 2930
rect 2430 2925 2460 2955
rect 2520 2945 2560 2985
rect 3080 2975 3120 2985
rect 3080 2955 3090 2975
rect 3110 2955 3120 2975
rect 3080 2945 3120 2955
rect 3140 2975 3175 2985
rect 3140 2955 3145 2975
rect 3165 2955 3175 2975
rect 3140 2945 3175 2955
rect 3265 2975 3305 2985
rect 3265 2955 3275 2975
rect 3295 2955 3305 2975
rect 3265 2945 3305 2955
rect 3445 2975 3485 2985
rect 3445 2955 3455 2975
rect 3475 2955 3485 2975
rect 3445 2945 3485 2955
rect 3625 2975 3665 2985
rect 3625 2955 3635 2975
rect 3655 2955 3665 2975
rect 3625 2945 3665 2955
rect 3805 2975 3845 2985
rect 3805 2955 3815 2975
rect 3835 2955 3845 2975
rect 3805 2945 3845 2955
rect 3985 2975 4025 2985
rect 3985 2955 3995 2975
rect 4015 2955 4025 2975
rect 3985 2945 4025 2955
rect 4165 2975 4205 2985
rect 4165 2955 4175 2975
rect 4195 2955 4205 2975
rect 4165 2945 4205 2955
rect 4345 2975 4385 2985
rect 4345 2955 4355 2975
rect 4375 2955 4385 2975
rect 4345 2945 4385 2955
rect 4525 2975 4565 2985
rect 4525 2955 4535 2975
rect 4555 2955 4565 2975
rect 4525 2945 4565 2955
rect 4705 2975 4745 2985
rect 4705 2955 4715 2975
rect 4735 2955 4745 2975
rect 4705 2945 4745 2955
rect 4835 2975 4870 2985
rect 4835 2955 4845 2975
rect 4865 2955 4870 2975
rect 4835 2945 4870 2955
rect 4890 2975 4925 2985
rect 4890 2955 4895 2975
rect 4915 2955 4925 2975
rect 4890 2945 4925 2955
rect 12855 2975 12925 3005
rect 12855 2955 12860 2975
rect 12880 2955 12900 2975
rect 12920 2955 12925 2975
rect 3095 2925 3115 2945
rect 3275 2925 3295 2945
rect 3455 2925 3475 2945
rect 3635 2925 3655 2945
rect 3815 2925 3835 2945
rect 3995 2925 4015 2945
rect 4175 2925 4195 2945
rect 4355 2925 4375 2945
rect 4535 2925 4555 2945
rect 4715 2925 4735 2945
rect 4895 2925 4915 2945
rect 11180 2940 11220 2950
rect 2960 2915 3030 2925
rect 1266 2865 1306 2900
rect 2330 2895 2375 2905
rect 2330 2870 2340 2895
rect 2365 2870 2375 2895
rect 2330 2860 2375 2870
rect 2960 2895 2965 2915
rect 2985 2895 3005 2915
rect 3025 2895 3030 2915
rect 2960 2865 3030 2895
rect -55 2825 -25 2855
rect 51 2850 96 2855
rect 51 2825 61 2850
rect 86 2825 96 2850
rect 51 2820 96 2825
rect 724 2850 769 2855
rect 724 2825 734 2850
rect 759 2825 769 2850
rect 724 2820 769 2825
rect 1210 2820 1240 2850
rect 2960 2845 2965 2865
rect 2985 2845 3005 2865
rect 3025 2845 3030 2865
rect 1261 2835 1306 2840
rect 1261 2810 1271 2835
rect 1296 2810 1306 2835
rect 1261 2805 1306 2810
rect 1960 2835 2005 2840
rect 1960 2810 1970 2835
rect 1995 2810 2005 2835
rect 1960 2805 2005 2810
rect 2330 2800 2370 2840
rect 2960 2835 3030 2845
rect 3090 2915 3120 2925
rect 3090 2895 3095 2915
rect 3115 2895 3120 2915
rect 3090 2865 3120 2895
rect 3090 2845 3095 2865
rect 3115 2845 3120 2865
rect 3090 2835 3120 2845
rect 3180 2915 3210 2925
rect 3180 2895 3185 2915
rect 3205 2895 3210 2915
rect 3180 2865 3210 2895
rect 3180 2845 3185 2865
rect 3205 2845 3210 2865
rect 3180 2835 3210 2845
rect 3270 2915 3300 2925
rect 3270 2895 3275 2915
rect 3295 2895 3300 2915
rect 3270 2865 3300 2895
rect 3270 2845 3275 2865
rect 3295 2845 3300 2865
rect 3270 2835 3300 2845
rect 3360 2915 3390 2925
rect 3360 2895 3365 2915
rect 3385 2895 3390 2915
rect 3360 2865 3390 2895
rect 3360 2845 3365 2865
rect 3385 2845 3390 2865
rect 3360 2835 3390 2845
rect 3450 2915 3480 2925
rect 3450 2895 3455 2915
rect 3475 2895 3480 2915
rect 3450 2865 3480 2895
rect 3450 2845 3455 2865
rect 3475 2845 3480 2865
rect 3450 2835 3480 2845
rect 3540 2915 3570 2925
rect 3540 2895 3545 2915
rect 3565 2895 3570 2915
rect 3540 2865 3570 2895
rect 3540 2845 3545 2865
rect 3565 2845 3570 2865
rect 3540 2835 3570 2845
rect 3630 2915 3660 2925
rect 3630 2895 3635 2915
rect 3655 2895 3660 2915
rect 3630 2865 3660 2895
rect 3630 2845 3635 2865
rect 3655 2845 3660 2865
rect 3630 2835 3660 2845
rect 3720 2915 3750 2925
rect 3720 2895 3725 2915
rect 3745 2895 3750 2915
rect 3720 2865 3750 2895
rect 3720 2845 3725 2865
rect 3745 2845 3750 2865
rect 3720 2835 3750 2845
rect 3810 2915 3840 2925
rect 3810 2895 3815 2915
rect 3835 2895 3840 2915
rect 3810 2865 3840 2895
rect 3810 2845 3815 2865
rect 3835 2845 3840 2865
rect 3810 2835 3840 2845
rect 3900 2915 3930 2925
rect 3900 2895 3905 2915
rect 3925 2895 3930 2915
rect 3900 2865 3930 2895
rect 3900 2845 3905 2865
rect 3925 2845 3930 2865
rect 3900 2835 3930 2845
rect 3990 2915 4020 2925
rect 3990 2895 3995 2915
rect 4015 2895 4020 2915
rect 3990 2865 4020 2895
rect 3990 2845 3995 2865
rect 4015 2845 4020 2865
rect 3990 2835 4020 2845
rect 4080 2915 4110 2925
rect 4080 2895 4085 2915
rect 4105 2895 4110 2915
rect 4080 2865 4110 2895
rect 4080 2845 4085 2865
rect 4105 2845 4110 2865
rect 4080 2835 4110 2845
rect 4170 2915 4200 2925
rect 4170 2895 4175 2915
rect 4195 2895 4200 2915
rect 4170 2865 4200 2895
rect 4170 2845 4175 2865
rect 4195 2845 4200 2865
rect 4170 2835 4200 2845
rect 4260 2915 4290 2925
rect 4260 2895 4265 2915
rect 4285 2895 4290 2915
rect 4260 2865 4290 2895
rect 4260 2845 4265 2865
rect 4285 2845 4290 2865
rect 4260 2835 4290 2845
rect 4350 2915 4380 2925
rect 4350 2895 4355 2915
rect 4375 2895 4380 2915
rect 4350 2865 4380 2895
rect 4350 2845 4355 2865
rect 4375 2845 4380 2865
rect 4350 2835 4380 2845
rect 4440 2915 4470 2925
rect 4440 2895 4445 2915
rect 4465 2895 4470 2915
rect 4440 2865 4470 2895
rect 4440 2845 4445 2865
rect 4465 2845 4470 2865
rect 4440 2835 4470 2845
rect 4530 2915 4560 2925
rect 4530 2895 4535 2915
rect 4555 2895 4560 2915
rect 4530 2865 4560 2895
rect 4530 2845 4535 2865
rect 4555 2845 4560 2865
rect 4530 2835 4560 2845
rect 4620 2915 4650 2925
rect 4620 2895 4625 2915
rect 4645 2895 4650 2915
rect 4620 2865 4650 2895
rect 4620 2845 4625 2865
rect 4645 2845 4650 2865
rect 4620 2835 4650 2845
rect 4710 2915 4740 2925
rect 4710 2895 4715 2915
rect 4735 2895 4740 2915
rect 4710 2865 4740 2895
rect 4710 2845 4715 2865
rect 4735 2845 4740 2865
rect 4710 2835 4740 2845
rect 4800 2915 4830 2925
rect 4800 2895 4805 2915
rect 4825 2895 4830 2915
rect 4800 2865 4830 2895
rect 4800 2845 4805 2865
rect 4825 2845 4830 2865
rect 4800 2835 4830 2845
rect 4890 2915 4920 2925
rect 4890 2895 4895 2915
rect 4915 2895 4920 2915
rect 4890 2865 4920 2895
rect 4890 2845 4895 2865
rect 4915 2845 4920 2865
rect 4890 2835 4920 2845
rect 4980 2915 5050 2925
rect 4980 2895 4985 2915
rect 5005 2895 5025 2915
rect 5045 2895 5050 2915
rect 11180 2920 11190 2940
rect 11210 2920 11220 2940
rect 11180 2910 11220 2920
rect 11340 2940 11380 2950
rect 11340 2920 11350 2940
rect 11370 2920 11380 2940
rect 11340 2910 11380 2920
rect 11460 2940 11500 2950
rect 11460 2920 11470 2940
rect 11490 2920 11500 2940
rect 11460 2910 11500 2920
rect 11580 2940 11620 2950
rect 11580 2920 11590 2940
rect 11610 2920 11620 2940
rect 11580 2910 11620 2920
rect 11700 2940 11740 2950
rect 11700 2920 11710 2940
rect 11730 2920 11740 2940
rect 11700 2910 11740 2920
rect 11820 2940 11860 2950
rect 11820 2920 11830 2940
rect 11850 2920 11860 2940
rect 11820 2910 11860 2920
rect 11940 2940 11980 2950
rect 11940 2920 11950 2940
rect 11970 2920 11980 2940
rect 11940 2910 11980 2920
rect 12060 2940 12100 2950
rect 12060 2920 12070 2940
rect 12090 2920 12100 2940
rect 12060 2910 12100 2920
rect 12180 2940 12220 2950
rect 12180 2920 12190 2940
rect 12210 2920 12220 2940
rect 12180 2910 12220 2920
rect 12300 2940 12340 2950
rect 12300 2920 12310 2940
rect 12330 2920 12340 2940
rect 12300 2910 12340 2920
rect 12420 2940 12460 2950
rect 12420 2920 12430 2940
rect 12450 2920 12460 2940
rect 12420 2910 12460 2920
rect 12480 2910 12520 2950
rect 12580 2940 12620 2950
rect 12855 2945 12925 2955
rect 12950 3225 12980 3235
rect 12950 3205 12955 3225
rect 12975 3205 12980 3225
rect 12950 3175 12980 3205
rect 12950 3155 12955 3175
rect 12975 3155 12980 3175
rect 12950 3125 12980 3155
rect 12950 3105 12955 3125
rect 12975 3105 12980 3125
rect 12950 3075 12980 3105
rect 12950 3055 12955 3075
rect 12975 3055 12980 3075
rect 12950 3025 12980 3055
rect 12950 3005 12955 3025
rect 12975 3005 12980 3025
rect 12950 2975 12980 3005
rect 12950 2955 12955 2975
rect 12975 2955 12980 2975
rect 12950 2945 12980 2955
rect 13005 3225 13035 3235
rect 13005 3205 13010 3225
rect 13030 3205 13035 3225
rect 13005 3175 13035 3205
rect 13005 3155 13010 3175
rect 13030 3155 13035 3175
rect 13005 3125 13035 3155
rect 13005 3105 13010 3125
rect 13030 3105 13035 3125
rect 13005 3075 13035 3105
rect 13005 3055 13010 3075
rect 13030 3055 13035 3075
rect 13005 3025 13035 3055
rect 13005 3005 13010 3025
rect 13030 3005 13035 3025
rect 13005 2975 13035 3005
rect 13005 2955 13010 2975
rect 13030 2955 13035 2975
rect 13005 2945 13035 2955
rect 13060 3225 13090 3235
rect 13060 3205 13065 3225
rect 13085 3205 13090 3225
rect 13060 3175 13090 3205
rect 13060 3155 13065 3175
rect 13085 3155 13090 3175
rect 13060 3125 13090 3155
rect 13060 3105 13065 3125
rect 13085 3105 13090 3125
rect 13060 3075 13090 3105
rect 13060 3055 13065 3075
rect 13085 3055 13090 3075
rect 13060 3025 13090 3055
rect 13060 3005 13065 3025
rect 13085 3005 13090 3025
rect 13060 2975 13090 3005
rect 13060 2955 13065 2975
rect 13085 2955 13090 2975
rect 13060 2945 13090 2955
rect 13115 3225 13145 3235
rect 13115 3205 13120 3225
rect 13140 3205 13145 3225
rect 13115 3175 13145 3205
rect 13115 3155 13120 3175
rect 13140 3155 13145 3175
rect 13115 3125 13145 3155
rect 13115 3105 13120 3125
rect 13140 3105 13145 3125
rect 13115 3075 13145 3105
rect 13115 3055 13120 3075
rect 13140 3055 13145 3075
rect 13115 3025 13145 3055
rect 13115 3005 13120 3025
rect 13140 3005 13145 3025
rect 13115 2975 13145 3005
rect 13115 2955 13120 2975
rect 13140 2955 13145 2975
rect 13115 2945 13145 2955
rect 13170 3225 13200 3235
rect 13170 3205 13175 3225
rect 13195 3205 13200 3225
rect 13170 3175 13200 3205
rect 13170 3155 13175 3175
rect 13195 3155 13200 3175
rect 13170 3125 13200 3155
rect 13170 3105 13175 3125
rect 13195 3105 13200 3125
rect 13170 3075 13200 3105
rect 13170 3055 13175 3075
rect 13195 3055 13200 3075
rect 13170 3025 13200 3055
rect 13170 3005 13175 3025
rect 13195 3005 13200 3025
rect 13170 2975 13200 3005
rect 13170 2955 13175 2975
rect 13195 2955 13200 2975
rect 13170 2945 13200 2955
rect 13225 3225 13255 3235
rect 13225 3205 13230 3225
rect 13250 3205 13255 3225
rect 13225 3175 13255 3205
rect 13225 3155 13230 3175
rect 13250 3155 13255 3175
rect 13225 3125 13255 3155
rect 13225 3105 13230 3125
rect 13250 3105 13255 3125
rect 13225 3075 13255 3105
rect 13225 3055 13230 3075
rect 13250 3055 13255 3075
rect 13225 3025 13255 3055
rect 13225 3005 13230 3025
rect 13250 3005 13255 3025
rect 13225 2975 13255 3005
rect 13225 2955 13230 2975
rect 13250 2955 13255 2975
rect 13225 2945 13255 2955
rect 13280 3225 13310 3235
rect 13280 3205 13285 3225
rect 13305 3205 13310 3225
rect 13280 3175 13310 3205
rect 13280 3155 13285 3175
rect 13305 3155 13310 3175
rect 13280 3125 13310 3155
rect 13280 3105 13285 3125
rect 13305 3105 13310 3125
rect 13280 3075 13310 3105
rect 13280 3055 13285 3075
rect 13305 3055 13310 3075
rect 13280 3025 13310 3055
rect 13280 3005 13285 3025
rect 13305 3005 13310 3025
rect 13280 2975 13310 3005
rect 13280 2955 13285 2975
rect 13305 2955 13310 2975
rect 13280 2945 13310 2955
rect 13335 3225 13365 3235
rect 13335 3205 13340 3225
rect 13360 3205 13365 3225
rect 13335 3175 13365 3205
rect 13335 3155 13340 3175
rect 13360 3155 13365 3175
rect 13335 3125 13365 3155
rect 13335 3105 13340 3125
rect 13360 3105 13365 3125
rect 13335 3075 13365 3105
rect 13335 3055 13340 3075
rect 13360 3055 13365 3075
rect 13335 3025 13365 3055
rect 13335 3005 13340 3025
rect 13360 3005 13365 3025
rect 13335 2975 13365 3005
rect 13335 2955 13340 2975
rect 13360 2955 13365 2975
rect 13335 2945 13365 2955
rect 13390 3225 13420 3235
rect 13390 3205 13395 3225
rect 13415 3205 13420 3225
rect 13390 3175 13420 3205
rect 13390 3155 13395 3175
rect 13415 3155 13420 3175
rect 13390 3125 13420 3155
rect 13390 3105 13395 3125
rect 13415 3105 13420 3125
rect 13390 3075 13420 3105
rect 13390 3055 13395 3075
rect 13415 3055 13420 3075
rect 13390 3025 13420 3055
rect 13390 3005 13395 3025
rect 13415 3005 13420 3025
rect 13390 2975 13420 3005
rect 13390 2955 13395 2975
rect 13415 2955 13420 2975
rect 13390 2945 13420 2955
rect 13445 3225 13475 3235
rect 13445 3205 13450 3225
rect 13470 3205 13475 3225
rect 13445 3175 13475 3205
rect 13445 3155 13450 3175
rect 13470 3155 13475 3175
rect 13445 3125 13475 3155
rect 13445 3105 13450 3125
rect 13470 3105 13475 3125
rect 13445 3075 13475 3105
rect 13445 3055 13450 3075
rect 13470 3055 13475 3075
rect 13445 3025 13475 3055
rect 13445 3005 13450 3025
rect 13470 3005 13475 3025
rect 13445 2975 13475 3005
rect 13445 2955 13450 2975
rect 13470 2955 13475 2975
rect 13445 2945 13475 2955
rect 13500 3225 13530 3235
rect 13500 3205 13505 3225
rect 13525 3205 13530 3225
rect 13500 3175 13530 3205
rect 13500 3155 13505 3175
rect 13525 3155 13530 3175
rect 13500 3125 13530 3155
rect 13500 3105 13505 3125
rect 13525 3105 13530 3125
rect 13500 3075 13530 3105
rect 13500 3055 13505 3075
rect 13525 3055 13530 3075
rect 13500 3025 13530 3055
rect 13500 3005 13505 3025
rect 13525 3005 13530 3025
rect 13500 2975 13530 3005
rect 13500 2955 13505 2975
rect 13525 2955 13530 2975
rect 13500 2945 13530 2955
rect 13555 3225 13585 3235
rect 13555 3205 13560 3225
rect 13580 3205 13585 3225
rect 13555 3175 13585 3205
rect 13555 3155 13560 3175
rect 13580 3155 13585 3175
rect 13555 3125 13585 3155
rect 13555 3105 13560 3125
rect 13580 3105 13585 3125
rect 13555 3075 13585 3105
rect 13555 3055 13560 3075
rect 13580 3055 13585 3075
rect 13555 3025 13585 3055
rect 13555 3005 13560 3025
rect 13580 3005 13585 3025
rect 13555 2975 13585 3005
rect 13555 2955 13560 2975
rect 13580 2955 13585 2975
rect 13555 2945 13585 2955
rect 13610 3225 13640 3235
rect 13610 3205 13615 3225
rect 13635 3205 13640 3225
rect 13610 3175 13640 3205
rect 13610 3155 13615 3175
rect 13635 3155 13640 3175
rect 13610 3125 13640 3155
rect 13610 3105 13615 3125
rect 13635 3105 13640 3125
rect 13610 3075 13640 3105
rect 13610 3055 13615 3075
rect 13635 3055 13640 3075
rect 13610 3025 13640 3055
rect 13610 3005 13615 3025
rect 13635 3005 13640 3025
rect 13610 2975 13640 3005
rect 13610 2955 13615 2975
rect 13635 2955 13640 2975
rect 13610 2945 13640 2955
rect 13665 3225 13695 3235
rect 13665 3205 13670 3225
rect 13690 3205 13695 3225
rect 13665 3175 13695 3205
rect 13665 3155 13670 3175
rect 13690 3155 13695 3175
rect 13665 3125 13695 3155
rect 13665 3105 13670 3125
rect 13690 3105 13695 3125
rect 13665 3075 13695 3105
rect 13665 3055 13670 3075
rect 13690 3055 13695 3075
rect 13665 3025 13695 3055
rect 13665 3005 13670 3025
rect 13690 3005 13695 3025
rect 13665 2975 13695 3005
rect 13665 2955 13670 2975
rect 13690 2955 13695 2975
rect 13665 2945 13695 2955
rect 13720 3225 13750 3235
rect 13720 3205 13725 3225
rect 13745 3205 13750 3225
rect 13720 3175 13750 3205
rect 13720 3155 13725 3175
rect 13745 3155 13750 3175
rect 13720 3125 13750 3155
rect 13720 3105 13725 3125
rect 13745 3105 13750 3125
rect 13720 3075 13750 3105
rect 13720 3055 13725 3075
rect 13745 3055 13750 3075
rect 13720 3025 13750 3055
rect 13720 3005 13725 3025
rect 13745 3005 13750 3025
rect 13720 2975 13750 3005
rect 13720 2955 13725 2975
rect 13745 2955 13750 2975
rect 13720 2945 13750 2955
rect 13775 3225 13805 3235
rect 13775 3205 13780 3225
rect 13800 3205 13805 3225
rect 13775 3175 13805 3205
rect 13775 3155 13780 3175
rect 13800 3155 13805 3175
rect 13775 3125 13805 3155
rect 13775 3105 13780 3125
rect 13800 3105 13805 3125
rect 13775 3075 13805 3105
rect 13775 3055 13780 3075
rect 13800 3055 13805 3075
rect 13775 3025 13805 3055
rect 13775 3005 13780 3025
rect 13800 3005 13805 3025
rect 13775 2975 13805 3005
rect 13775 2955 13780 2975
rect 13800 2955 13805 2975
rect 13775 2945 13805 2955
rect 13830 3225 13860 3235
rect 13830 3205 13835 3225
rect 13855 3205 13860 3225
rect 13830 3175 13860 3205
rect 13830 3155 13835 3175
rect 13855 3155 13860 3175
rect 13830 3125 13860 3155
rect 13830 3105 13835 3125
rect 13855 3105 13860 3125
rect 13830 3075 13860 3105
rect 13830 3055 13835 3075
rect 13855 3055 13860 3075
rect 13830 3025 13860 3055
rect 13830 3005 13835 3025
rect 13855 3005 13860 3025
rect 13830 2975 13860 3005
rect 13830 2955 13835 2975
rect 13855 2955 13860 2975
rect 13830 2945 13860 2955
rect 13885 3225 13915 3235
rect 13885 3205 13890 3225
rect 13910 3205 13915 3225
rect 13885 3175 13915 3205
rect 13885 3155 13890 3175
rect 13910 3155 13915 3175
rect 13885 3125 13915 3155
rect 13885 3105 13890 3125
rect 13910 3105 13915 3125
rect 13885 3075 13915 3105
rect 13885 3055 13890 3075
rect 13910 3055 13915 3075
rect 13885 3025 13915 3055
rect 13885 3005 13890 3025
rect 13910 3005 13915 3025
rect 13885 2975 13915 3005
rect 13885 2955 13890 2975
rect 13910 2955 13915 2975
rect 13885 2945 13915 2955
rect 13940 3225 13970 3235
rect 13940 3205 13945 3225
rect 13965 3205 13970 3225
rect 13940 3175 13970 3205
rect 13940 3155 13945 3175
rect 13965 3155 13970 3175
rect 13940 3125 13970 3155
rect 13940 3105 13945 3125
rect 13965 3105 13970 3125
rect 13940 3075 13970 3105
rect 13940 3055 13945 3075
rect 13965 3055 13970 3075
rect 13940 3025 13970 3055
rect 13940 3005 13945 3025
rect 13965 3005 13970 3025
rect 13940 2975 13970 3005
rect 13940 2955 13945 2975
rect 13965 2955 13970 2975
rect 13940 2945 13970 2955
rect 13995 3225 14025 3235
rect 13995 3205 14000 3225
rect 14020 3205 14025 3225
rect 13995 3175 14025 3205
rect 13995 3155 14000 3175
rect 14020 3155 14025 3175
rect 13995 3125 14025 3155
rect 13995 3105 14000 3125
rect 14020 3105 14025 3125
rect 13995 3075 14025 3105
rect 13995 3055 14000 3075
rect 14020 3055 14025 3075
rect 13995 3025 14025 3055
rect 13995 3005 14000 3025
rect 14020 3005 14025 3025
rect 13995 2975 14025 3005
rect 13995 2955 14000 2975
rect 14020 2955 14025 2975
rect 13995 2945 14025 2955
rect 14050 3225 14080 3235
rect 14050 3205 14055 3225
rect 14075 3205 14080 3225
rect 14050 3175 14080 3205
rect 14050 3155 14055 3175
rect 14075 3155 14080 3175
rect 14050 3125 14080 3155
rect 14050 3105 14055 3125
rect 14075 3105 14080 3125
rect 14050 3075 14080 3105
rect 14050 3055 14055 3075
rect 14075 3055 14080 3075
rect 14050 3025 14080 3055
rect 14050 3005 14055 3025
rect 14075 3005 14080 3025
rect 14050 2975 14080 3005
rect 14050 2955 14055 2975
rect 14075 2955 14080 2975
rect 14050 2945 14080 2955
rect 14105 3225 14175 3235
rect 14105 3205 14110 3225
rect 14130 3205 14150 3225
rect 14170 3205 14175 3225
rect 18120 3215 18140 3235
rect 18290 3215 18310 3235
rect 18610 3215 18630 3235
rect 14105 3175 14175 3205
rect 18080 3205 18140 3215
rect 18080 3185 18090 3205
rect 18110 3195 18140 3205
rect 18280 3205 18320 3215
rect 18110 3185 18120 3195
rect 18080 3175 18120 3185
rect 18280 3185 18290 3205
rect 18310 3185 18320 3205
rect 18280 3175 18320 3185
rect 18405 3205 18440 3215
rect 18405 3185 18410 3205
rect 18430 3185 18440 3205
rect 18405 3175 18440 3185
rect 18480 3205 18515 3215
rect 18480 3185 18490 3205
rect 18510 3185 18515 3205
rect 18480 3175 18515 3185
rect 18600 3205 18640 3215
rect 18600 3185 18610 3205
rect 18630 3185 18640 3205
rect 18600 3175 18640 3185
rect 18685 3210 18755 3240
rect 18685 3190 18690 3210
rect 18710 3190 18730 3210
rect 18750 3190 18755 3210
rect 18685 3180 18755 3190
rect 18785 3560 18815 3570
rect 18785 3540 18790 3560
rect 18810 3540 18815 3560
rect 18785 3510 18815 3540
rect 18785 3490 18790 3510
rect 18810 3490 18815 3510
rect 18785 3460 18815 3490
rect 18785 3440 18790 3460
rect 18810 3440 18815 3460
rect 18785 3410 18815 3440
rect 18785 3390 18790 3410
rect 18810 3390 18815 3410
rect 18785 3360 18815 3390
rect 18785 3340 18790 3360
rect 18810 3340 18815 3360
rect 18785 3310 18815 3340
rect 18785 3290 18790 3310
rect 18810 3290 18815 3310
rect 18785 3260 18815 3290
rect 18785 3240 18790 3260
rect 18810 3240 18815 3260
rect 18785 3210 18815 3240
rect 18785 3190 18790 3210
rect 18810 3190 18815 3210
rect 18785 3180 18815 3190
rect 18845 3560 18875 3570
rect 18845 3540 18850 3560
rect 18870 3540 18875 3560
rect 18845 3510 18875 3540
rect 18845 3490 18850 3510
rect 18870 3490 18875 3510
rect 18845 3460 18875 3490
rect 18845 3440 18850 3460
rect 18870 3440 18875 3460
rect 18845 3410 18875 3440
rect 18845 3390 18850 3410
rect 18870 3390 18875 3410
rect 18845 3360 18875 3390
rect 18845 3340 18850 3360
rect 18870 3340 18875 3360
rect 18845 3310 18875 3340
rect 18845 3290 18850 3310
rect 18870 3290 18875 3310
rect 18845 3260 18875 3290
rect 18845 3240 18850 3260
rect 18870 3240 18875 3260
rect 18845 3210 18875 3240
rect 18845 3190 18850 3210
rect 18870 3190 18875 3210
rect 18845 3180 18875 3190
rect 18905 3560 18935 3570
rect 18905 3540 18910 3560
rect 18930 3540 18935 3560
rect 18905 3510 18935 3540
rect 18905 3490 18910 3510
rect 18930 3490 18935 3510
rect 18905 3460 18935 3490
rect 18905 3440 18910 3460
rect 18930 3440 18935 3460
rect 18905 3410 18935 3440
rect 18905 3390 18910 3410
rect 18930 3390 18935 3410
rect 18905 3360 18935 3390
rect 18905 3340 18910 3360
rect 18930 3340 18935 3360
rect 18905 3310 18935 3340
rect 18905 3290 18910 3310
rect 18930 3290 18935 3310
rect 18905 3260 18935 3290
rect 18905 3240 18910 3260
rect 18930 3240 18935 3260
rect 18905 3210 18935 3240
rect 18905 3190 18910 3210
rect 18930 3190 18935 3210
rect 18905 3180 18935 3190
rect 18965 3560 18995 3570
rect 18965 3540 18970 3560
rect 18990 3540 18995 3560
rect 18965 3510 18995 3540
rect 18965 3490 18970 3510
rect 18990 3490 18995 3510
rect 18965 3460 18995 3490
rect 18965 3440 18970 3460
rect 18990 3440 18995 3460
rect 18965 3410 18995 3440
rect 18965 3390 18970 3410
rect 18990 3390 18995 3410
rect 18965 3360 18995 3390
rect 18965 3340 18970 3360
rect 18990 3340 18995 3360
rect 18965 3310 18995 3340
rect 18965 3290 18970 3310
rect 18990 3290 18995 3310
rect 18965 3260 18995 3290
rect 18965 3240 18970 3260
rect 18990 3240 18995 3260
rect 18965 3210 18995 3240
rect 18965 3190 18970 3210
rect 18990 3190 18995 3210
rect 18965 3180 18995 3190
rect 19025 3560 19055 3570
rect 19025 3540 19030 3560
rect 19050 3540 19055 3560
rect 19025 3510 19055 3540
rect 19025 3490 19030 3510
rect 19050 3490 19055 3510
rect 19025 3460 19055 3490
rect 19025 3440 19030 3460
rect 19050 3440 19055 3460
rect 19025 3410 19055 3440
rect 19025 3390 19030 3410
rect 19050 3390 19055 3410
rect 19025 3360 19055 3390
rect 19025 3340 19030 3360
rect 19050 3340 19055 3360
rect 19025 3310 19055 3340
rect 19025 3290 19030 3310
rect 19050 3290 19055 3310
rect 19025 3260 19055 3290
rect 19025 3240 19030 3260
rect 19050 3240 19055 3260
rect 19025 3210 19055 3240
rect 19025 3190 19030 3210
rect 19050 3190 19055 3210
rect 19025 3180 19055 3190
rect 19085 3560 19115 3570
rect 19085 3540 19090 3560
rect 19110 3540 19115 3560
rect 19085 3510 19115 3540
rect 19085 3490 19090 3510
rect 19110 3490 19115 3510
rect 19085 3460 19115 3490
rect 19085 3440 19090 3460
rect 19110 3440 19115 3460
rect 19085 3410 19115 3440
rect 19085 3390 19090 3410
rect 19110 3390 19115 3410
rect 19085 3360 19115 3390
rect 19085 3340 19090 3360
rect 19110 3340 19115 3360
rect 19085 3310 19115 3340
rect 19085 3290 19090 3310
rect 19110 3290 19115 3310
rect 19085 3260 19115 3290
rect 19085 3240 19090 3260
rect 19110 3240 19115 3260
rect 19085 3210 19115 3240
rect 19085 3190 19090 3210
rect 19110 3190 19115 3210
rect 19085 3180 19115 3190
rect 19145 3560 19175 3570
rect 19145 3540 19150 3560
rect 19170 3540 19175 3560
rect 19145 3510 19175 3540
rect 19145 3490 19150 3510
rect 19170 3490 19175 3510
rect 19145 3460 19175 3490
rect 19145 3440 19150 3460
rect 19170 3440 19175 3460
rect 19145 3410 19175 3440
rect 19145 3390 19150 3410
rect 19170 3390 19175 3410
rect 19145 3360 19175 3390
rect 19145 3340 19150 3360
rect 19170 3340 19175 3360
rect 19145 3310 19175 3340
rect 19145 3290 19150 3310
rect 19170 3290 19175 3310
rect 19145 3260 19175 3290
rect 19145 3240 19150 3260
rect 19170 3240 19175 3260
rect 19145 3210 19175 3240
rect 19145 3190 19150 3210
rect 19170 3190 19175 3210
rect 19145 3180 19175 3190
rect 19205 3560 19235 3570
rect 19205 3540 19210 3560
rect 19230 3540 19235 3560
rect 19205 3510 19235 3540
rect 19205 3490 19210 3510
rect 19230 3490 19235 3510
rect 19205 3460 19235 3490
rect 19205 3440 19210 3460
rect 19230 3440 19235 3460
rect 19205 3410 19235 3440
rect 19205 3390 19210 3410
rect 19230 3390 19235 3410
rect 19205 3360 19235 3390
rect 19205 3340 19210 3360
rect 19230 3340 19235 3360
rect 19205 3310 19235 3340
rect 19205 3290 19210 3310
rect 19230 3290 19235 3310
rect 19205 3260 19235 3290
rect 19205 3240 19210 3260
rect 19230 3240 19235 3260
rect 19205 3210 19235 3240
rect 19205 3190 19210 3210
rect 19230 3190 19235 3210
rect 19205 3180 19235 3190
rect 19265 3560 19295 3570
rect 19265 3540 19270 3560
rect 19290 3540 19295 3560
rect 19265 3510 19295 3540
rect 19265 3490 19270 3510
rect 19290 3490 19295 3510
rect 19265 3460 19295 3490
rect 19265 3440 19270 3460
rect 19290 3440 19295 3460
rect 19265 3410 19295 3440
rect 19265 3390 19270 3410
rect 19290 3390 19295 3410
rect 19265 3360 19295 3390
rect 19265 3340 19270 3360
rect 19290 3340 19295 3360
rect 19265 3310 19295 3340
rect 19265 3290 19270 3310
rect 19290 3290 19295 3310
rect 19265 3260 19295 3290
rect 19265 3240 19270 3260
rect 19290 3240 19295 3260
rect 19265 3210 19295 3240
rect 19265 3190 19270 3210
rect 19290 3190 19295 3210
rect 19265 3180 19295 3190
rect 19325 3560 19355 3570
rect 19325 3540 19330 3560
rect 19350 3540 19355 3560
rect 19325 3510 19355 3540
rect 19325 3490 19330 3510
rect 19350 3490 19355 3510
rect 19325 3460 19355 3490
rect 19325 3440 19330 3460
rect 19350 3440 19355 3460
rect 19325 3410 19355 3440
rect 19325 3390 19330 3410
rect 19350 3390 19355 3410
rect 19325 3360 19355 3390
rect 19325 3340 19330 3360
rect 19350 3340 19355 3360
rect 19325 3310 19355 3340
rect 19325 3290 19330 3310
rect 19350 3290 19355 3310
rect 19325 3260 19355 3290
rect 19325 3240 19330 3260
rect 19350 3240 19355 3260
rect 19325 3210 19355 3240
rect 19325 3190 19330 3210
rect 19350 3190 19355 3210
rect 19325 3180 19355 3190
rect 19385 3560 19415 3570
rect 19385 3540 19390 3560
rect 19410 3540 19415 3560
rect 19385 3510 19415 3540
rect 19385 3490 19390 3510
rect 19410 3490 19415 3510
rect 19385 3460 19415 3490
rect 19385 3440 19390 3460
rect 19410 3440 19415 3460
rect 19385 3410 19415 3440
rect 19385 3390 19390 3410
rect 19410 3390 19415 3410
rect 19385 3360 19415 3390
rect 19385 3340 19390 3360
rect 19410 3340 19415 3360
rect 19385 3310 19415 3340
rect 19385 3290 19390 3310
rect 19410 3290 19415 3310
rect 19385 3260 19415 3290
rect 19385 3240 19390 3260
rect 19410 3240 19415 3260
rect 19385 3210 19415 3240
rect 19385 3190 19390 3210
rect 19410 3190 19415 3210
rect 19385 3180 19415 3190
rect 19445 3560 19475 3570
rect 19445 3540 19450 3560
rect 19470 3540 19475 3560
rect 19445 3510 19475 3540
rect 19445 3490 19450 3510
rect 19470 3490 19475 3510
rect 19445 3460 19475 3490
rect 19445 3440 19450 3460
rect 19470 3440 19475 3460
rect 19445 3410 19475 3440
rect 19445 3390 19450 3410
rect 19470 3390 19475 3410
rect 19445 3360 19475 3390
rect 19445 3340 19450 3360
rect 19470 3340 19475 3360
rect 19445 3310 19475 3340
rect 19445 3290 19450 3310
rect 19470 3290 19475 3310
rect 19445 3260 19475 3290
rect 19445 3240 19450 3260
rect 19470 3240 19475 3260
rect 19445 3210 19475 3240
rect 19445 3190 19450 3210
rect 19470 3190 19475 3210
rect 19445 3180 19475 3190
rect 19505 3560 19535 3570
rect 19505 3540 19510 3560
rect 19530 3540 19535 3560
rect 19505 3510 19535 3540
rect 19505 3490 19510 3510
rect 19530 3490 19535 3510
rect 19505 3460 19535 3490
rect 19505 3440 19510 3460
rect 19530 3440 19535 3460
rect 19505 3410 19535 3440
rect 19505 3390 19510 3410
rect 19530 3390 19535 3410
rect 19505 3360 19535 3390
rect 19505 3340 19510 3360
rect 19530 3340 19535 3360
rect 19505 3310 19535 3340
rect 19505 3290 19510 3310
rect 19530 3290 19535 3310
rect 19505 3260 19535 3290
rect 19505 3240 19510 3260
rect 19530 3240 19535 3260
rect 19505 3210 19535 3240
rect 19505 3190 19510 3210
rect 19530 3190 19535 3210
rect 19505 3180 19535 3190
rect 19565 3560 19595 3570
rect 19565 3540 19570 3560
rect 19590 3540 19595 3560
rect 19565 3510 19595 3540
rect 19565 3490 19570 3510
rect 19590 3490 19595 3510
rect 19565 3460 19595 3490
rect 19565 3440 19570 3460
rect 19590 3440 19595 3460
rect 19565 3410 19595 3440
rect 19565 3390 19570 3410
rect 19590 3390 19595 3410
rect 19565 3360 19595 3390
rect 19565 3340 19570 3360
rect 19590 3340 19595 3360
rect 19565 3310 19595 3340
rect 19565 3290 19570 3310
rect 19590 3290 19595 3310
rect 19565 3260 19595 3290
rect 19565 3240 19570 3260
rect 19590 3240 19595 3260
rect 19565 3210 19595 3240
rect 19565 3190 19570 3210
rect 19590 3190 19595 3210
rect 19565 3180 19595 3190
rect 19625 3560 19655 3570
rect 19625 3540 19630 3560
rect 19650 3540 19655 3560
rect 19625 3510 19655 3540
rect 19625 3490 19630 3510
rect 19650 3490 19655 3510
rect 19625 3460 19655 3490
rect 19625 3440 19630 3460
rect 19650 3440 19655 3460
rect 19625 3410 19655 3440
rect 19625 3390 19630 3410
rect 19650 3390 19655 3410
rect 19625 3360 19655 3390
rect 19625 3340 19630 3360
rect 19650 3340 19655 3360
rect 19625 3310 19655 3340
rect 19625 3290 19630 3310
rect 19650 3290 19655 3310
rect 19625 3260 19655 3290
rect 19625 3240 19630 3260
rect 19650 3240 19655 3260
rect 19625 3210 19655 3240
rect 19625 3190 19630 3210
rect 19650 3190 19655 3210
rect 19625 3180 19655 3190
rect 19685 3560 19715 3570
rect 19685 3540 19690 3560
rect 19710 3540 19715 3560
rect 19685 3510 19715 3540
rect 19685 3490 19690 3510
rect 19710 3490 19715 3510
rect 19685 3460 19715 3490
rect 19685 3440 19690 3460
rect 19710 3440 19715 3460
rect 19685 3410 19715 3440
rect 19685 3390 19690 3410
rect 19710 3390 19715 3410
rect 19685 3360 19715 3390
rect 19685 3340 19690 3360
rect 19710 3340 19715 3360
rect 19685 3310 19715 3340
rect 19685 3290 19690 3310
rect 19710 3290 19715 3310
rect 19685 3260 19715 3290
rect 19685 3240 19690 3260
rect 19710 3240 19715 3260
rect 19685 3210 19715 3240
rect 19685 3190 19690 3210
rect 19710 3190 19715 3210
rect 19685 3180 19715 3190
rect 19745 3560 19775 3570
rect 19745 3540 19750 3560
rect 19770 3540 19775 3560
rect 19745 3510 19775 3540
rect 19745 3490 19750 3510
rect 19770 3490 19775 3510
rect 19745 3460 19775 3490
rect 19745 3440 19750 3460
rect 19770 3440 19775 3460
rect 19745 3410 19775 3440
rect 19745 3390 19750 3410
rect 19770 3390 19775 3410
rect 19745 3360 19775 3390
rect 19745 3340 19750 3360
rect 19770 3340 19775 3360
rect 19745 3310 19775 3340
rect 19745 3290 19750 3310
rect 19770 3290 19775 3310
rect 19745 3260 19775 3290
rect 19745 3240 19750 3260
rect 19770 3240 19775 3260
rect 19745 3210 19775 3240
rect 19745 3190 19750 3210
rect 19770 3190 19775 3210
rect 19745 3180 19775 3190
rect 19805 3560 19835 3570
rect 19805 3540 19810 3560
rect 19830 3540 19835 3560
rect 19805 3510 19835 3540
rect 19805 3490 19810 3510
rect 19830 3490 19835 3510
rect 19805 3460 19835 3490
rect 19805 3440 19810 3460
rect 19830 3440 19835 3460
rect 19805 3410 19835 3440
rect 19805 3390 19810 3410
rect 19830 3390 19835 3410
rect 19805 3360 19835 3390
rect 19805 3340 19810 3360
rect 19830 3340 19835 3360
rect 19805 3310 19835 3340
rect 19805 3290 19810 3310
rect 19830 3290 19835 3310
rect 19805 3260 19835 3290
rect 19805 3240 19810 3260
rect 19830 3240 19835 3260
rect 19805 3210 19835 3240
rect 19805 3190 19810 3210
rect 19830 3190 19835 3210
rect 19805 3180 19835 3190
rect 19865 3560 19895 3570
rect 19865 3540 19870 3560
rect 19890 3540 19895 3560
rect 19865 3510 19895 3540
rect 19865 3490 19870 3510
rect 19890 3490 19895 3510
rect 19865 3460 19895 3490
rect 19865 3440 19870 3460
rect 19890 3440 19895 3460
rect 19865 3410 19895 3440
rect 19865 3390 19870 3410
rect 19890 3390 19895 3410
rect 19865 3360 19895 3390
rect 19865 3340 19870 3360
rect 19890 3340 19895 3360
rect 19865 3310 19895 3340
rect 19865 3290 19870 3310
rect 19890 3290 19895 3310
rect 19865 3260 19895 3290
rect 19865 3240 19870 3260
rect 19890 3240 19895 3260
rect 19865 3210 19895 3240
rect 19865 3190 19870 3210
rect 19890 3190 19895 3210
rect 19865 3180 19895 3190
rect 19925 3560 19955 3570
rect 19925 3540 19930 3560
rect 19950 3540 19955 3560
rect 19925 3510 19955 3540
rect 19925 3490 19930 3510
rect 19950 3490 19955 3510
rect 19925 3460 19955 3490
rect 19925 3440 19930 3460
rect 19950 3440 19955 3460
rect 19925 3410 19955 3440
rect 19925 3390 19930 3410
rect 19950 3390 19955 3410
rect 19925 3360 19955 3390
rect 19925 3340 19930 3360
rect 19950 3340 19955 3360
rect 19925 3310 19955 3340
rect 19925 3290 19930 3310
rect 19950 3290 19955 3310
rect 19925 3260 19955 3290
rect 19925 3240 19930 3260
rect 19950 3240 19955 3260
rect 19925 3210 19955 3240
rect 19925 3190 19930 3210
rect 19950 3190 19955 3210
rect 19925 3180 19955 3190
rect 19985 3560 20015 3570
rect 19985 3540 19990 3560
rect 20010 3540 20015 3560
rect 19985 3510 20015 3540
rect 19985 3490 19990 3510
rect 20010 3490 20015 3510
rect 19985 3460 20015 3490
rect 19985 3440 19990 3460
rect 20010 3440 20015 3460
rect 19985 3410 20015 3440
rect 19985 3390 19990 3410
rect 20010 3390 20015 3410
rect 19985 3360 20015 3390
rect 19985 3340 19990 3360
rect 20010 3340 20015 3360
rect 19985 3310 20015 3340
rect 19985 3290 19990 3310
rect 20010 3290 20015 3310
rect 19985 3260 20015 3290
rect 19985 3240 19990 3260
rect 20010 3240 20015 3260
rect 19985 3210 20015 3240
rect 19985 3190 19990 3210
rect 20010 3190 20015 3210
rect 19985 3180 20015 3190
rect 20045 3560 20115 3570
rect 20045 3540 20050 3560
rect 20070 3540 20090 3560
rect 20110 3540 20115 3560
rect 20045 3510 20115 3540
rect 20045 3490 20050 3510
rect 20070 3490 20090 3510
rect 20110 3490 20115 3510
rect 20045 3460 20115 3490
rect 20045 3440 20050 3460
rect 20070 3440 20090 3460
rect 20110 3440 20115 3460
rect 20045 3410 20115 3440
rect 20045 3390 20050 3410
rect 20070 3390 20090 3410
rect 20110 3390 20115 3410
rect 20045 3360 20115 3390
rect 20045 3340 20050 3360
rect 20070 3340 20090 3360
rect 20110 3340 20115 3360
rect 20045 3310 20115 3340
rect 20045 3290 20050 3310
rect 20070 3290 20090 3310
rect 20110 3290 20115 3310
rect 20045 3260 20115 3290
rect 20045 3240 20050 3260
rect 20070 3240 20090 3260
rect 20110 3240 20115 3260
rect 20445 3285 20485 3295
rect 20445 3265 20455 3285
rect 20475 3265 20485 3285
rect 20445 3255 20485 3265
rect 20555 3285 20595 3295
rect 20555 3265 20565 3285
rect 20585 3265 20595 3285
rect 20555 3255 20595 3265
rect 20665 3285 20705 3295
rect 20665 3265 20675 3285
rect 20695 3265 20705 3285
rect 20665 3255 20705 3265
rect 20775 3285 20815 3295
rect 20775 3265 20785 3285
rect 20805 3265 20815 3285
rect 20775 3255 20815 3265
rect 20885 3285 20925 3295
rect 20885 3265 20895 3285
rect 20915 3265 20925 3285
rect 20885 3255 20925 3265
rect 20995 3285 21035 3295
rect 20995 3265 21005 3285
rect 21025 3265 21035 3285
rect 20995 3255 21035 3265
rect 21105 3285 21145 3295
rect 21105 3265 21115 3285
rect 21135 3265 21145 3285
rect 21105 3255 21145 3265
rect 21215 3285 21255 3295
rect 21215 3265 21225 3285
rect 21245 3265 21255 3285
rect 21215 3255 21255 3265
rect 21325 3285 21365 3295
rect 21325 3265 21335 3285
rect 21355 3265 21365 3285
rect 21325 3255 21365 3265
rect 21435 3285 21475 3295
rect 21435 3265 21445 3285
rect 21465 3265 21475 3285
rect 21435 3255 21475 3265
rect 21545 3285 21585 3295
rect 21545 3265 21555 3285
rect 21575 3265 21585 3285
rect 21545 3255 21585 3265
rect 20045 3210 20115 3240
rect 20455 3235 20475 3255
rect 20565 3235 20585 3255
rect 20675 3235 20695 3255
rect 20785 3235 20805 3255
rect 20895 3235 20915 3255
rect 21005 3235 21025 3255
rect 21115 3235 21135 3255
rect 21225 3235 21245 3255
rect 21335 3235 21355 3255
rect 21445 3235 21465 3255
rect 21555 3235 21575 3255
rect 20045 3190 20050 3210
rect 20070 3190 20090 3210
rect 20110 3190 20115 3210
rect 20045 3180 20115 3190
rect 20355 3225 20425 3235
rect 20355 3205 20360 3225
rect 20380 3205 20400 3225
rect 20420 3205 20425 3225
rect 14105 3155 14110 3175
rect 14130 3155 14150 3175
rect 14170 3155 14175 3175
rect 18790 3160 18810 3180
rect 18910 3160 18930 3180
rect 19030 3160 19050 3180
rect 19150 3160 19170 3180
rect 19270 3160 19290 3180
rect 19390 3160 19410 3180
rect 19510 3160 19530 3180
rect 19630 3160 19650 3180
rect 19750 3160 19770 3180
rect 19870 3160 19890 3180
rect 19990 3160 20010 3180
rect 20355 3175 20425 3205
rect 14105 3125 14175 3155
rect 14105 3105 14110 3125
rect 14130 3105 14150 3125
rect 14170 3105 14175 3125
rect 18780 3150 18820 3160
rect 18780 3130 18790 3150
rect 18810 3130 18820 3150
rect 18780 3120 18820 3130
rect 18900 3150 18940 3160
rect 18900 3130 18910 3150
rect 18930 3130 18940 3150
rect 18900 3120 18940 3130
rect 19020 3150 19060 3160
rect 19020 3130 19030 3150
rect 19050 3130 19060 3150
rect 19020 3120 19060 3130
rect 19140 3150 19180 3160
rect 19140 3130 19150 3150
rect 19170 3130 19180 3150
rect 19140 3120 19180 3130
rect 19260 3150 19300 3160
rect 19260 3130 19270 3150
rect 19290 3130 19300 3150
rect 19260 3120 19300 3130
rect 19323 3150 19357 3160
rect 19323 3130 19331 3150
rect 19349 3130 19357 3150
rect 19323 3120 19357 3130
rect 19380 3150 19420 3160
rect 19380 3130 19390 3150
rect 19410 3130 19420 3150
rect 19380 3120 19420 3130
rect 19500 3150 19540 3160
rect 19500 3130 19510 3150
rect 19530 3130 19540 3150
rect 19500 3120 19540 3130
rect 19620 3150 19660 3160
rect 19620 3130 19630 3150
rect 19650 3130 19660 3150
rect 19620 3120 19660 3130
rect 19740 3150 19780 3160
rect 19740 3130 19750 3150
rect 19770 3130 19780 3150
rect 19740 3120 19780 3130
rect 19860 3150 19900 3160
rect 19860 3130 19870 3150
rect 19890 3130 19900 3150
rect 19860 3120 19900 3130
rect 19980 3150 20020 3160
rect 19980 3130 19990 3150
rect 20010 3130 20020 3150
rect 19980 3120 20020 3130
rect 20355 3155 20360 3175
rect 20380 3155 20400 3175
rect 20420 3155 20425 3175
rect 20355 3125 20425 3155
rect 14105 3075 14175 3105
rect 14105 3055 14110 3075
rect 14130 3055 14150 3075
rect 14170 3055 14175 3075
rect 14105 3025 14175 3055
rect 14105 3005 14110 3025
rect 14130 3005 14150 3025
rect 14170 3005 14175 3025
rect 14105 2975 14175 3005
rect 14105 2955 14110 2975
rect 14130 2955 14150 2975
rect 14170 2955 14175 2975
rect 14105 2945 14175 2955
rect 20355 3105 20360 3125
rect 20380 3105 20400 3125
rect 20420 3105 20425 3125
rect 20355 3075 20425 3105
rect 20355 3055 20360 3075
rect 20380 3055 20400 3075
rect 20420 3055 20425 3075
rect 20355 3025 20425 3055
rect 20355 3005 20360 3025
rect 20380 3005 20400 3025
rect 20420 3005 20425 3025
rect 20355 2975 20425 3005
rect 20355 2955 20360 2975
rect 20380 2955 20400 2975
rect 20420 2955 20425 2975
rect 12580 2920 12590 2940
rect 12610 2920 12620 2940
rect 12860 2925 12880 2945
rect 13010 2925 13030 2945
rect 13120 2925 13140 2945
rect 13230 2925 13250 2945
rect 13340 2925 13360 2945
rect 13450 2925 13470 2945
rect 13560 2925 13580 2945
rect 13670 2925 13690 2945
rect 13780 2925 13800 2945
rect 13890 2925 13910 2945
rect 14000 2925 14020 2945
rect 14150 2925 14170 2945
rect 18680 2940 18720 2950
rect 12580 2910 12620 2920
rect 12850 2915 12890 2925
rect 4980 2865 5050 2895
rect 11190 2890 11210 2910
rect 11350 2890 11370 2910
rect 11470 2890 11490 2910
rect 11590 2890 11610 2910
rect 11710 2890 11730 2910
rect 11830 2890 11850 2910
rect 11950 2890 11970 2910
rect 12070 2890 12090 2910
rect 12190 2890 12210 2910
rect 12310 2890 12330 2910
rect 12430 2890 12450 2910
rect 12590 2890 12610 2910
rect 12850 2895 12860 2915
rect 12880 2895 12890 2915
rect 4980 2845 4985 2865
rect 5005 2845 5025 2865
rect 5045 2845 5050 2865
rect 4980 2835 5050 2845
rect 11185 2880 11255 2890
rect 11185 2860 11190 2880
rect 11210 2860 11230 2880
rect 11250 2860 11255 2880
rect 3005 2815 3025 2835
rect 3185 2815 3205 2835
rect 3365 2815 3385 2835
rect 3545 2815 3565 2835
rect 3725 2815 3745 2835
rect 3905 2815 3925 2835
rect 4085 2815 4105 2835
rect 4265 2815 4285 2835
rect 4445 2815 4465 2835
rect 4625 2815 4645 2835
rect 4805 2815 4825 2835
rect 4985 2815 5005 2835
rect 11185 2830 11255 2860
rect 2995 2805 3035 2815
rect -10 2765 20 2795
rect 51 2790 96 2795
rect 51 2765 61 2790
rect 86 2765 96 2790
rect 51 2760 96 2765
rect 724 2790 769 2795
rect 724 2765 734 2790
rect 759 2765 769 2790
rect 724 2760 769 2765
rect 2620 2755 2660 2795
rect 2995 2785 3005 2805
rect 3025 2785 3035 2805
rect 2995 2775 3035 2785
rect 3175 2805 3215 2815
rect 3175 2785 3185 2805
rect 3205 2785 3215 2805
rect 3175 2775 3215 2785
rect 3355 2805 3395 2815
rect 3355 2785 3365 2805
rect 3385 2785 3395 2805
rect 3355 2775 3395 2785
rect 3535 2805 3575 2815
rect 3535 2785 3545 2805
rect 3565 2785 3575 2805
rect 3535 2775 3575 2785
rect 3715 2805 3755 2815
rect 3715 2785 3725 2805
rect 3745 2785 3755 2805
rect 3715 2775 3755 2785
rect 3895 2805 3935 2815
rect 3895 2785 3905 2805
rect 3925 2785 3935 2805
rect 3895 2775 3935 2785
rect 4075 2805 4115 2815
rect 4075 2785 4085 2805
rect 4105 2785 4115 2805
rect 4075 2775 4115 2785
rect 4255 2805 4295 2815
rect 4255 2785 4265 2805
rect 4285 2785 4295 2805
rect 4255 2775 4295 2785
rect 4435 2805 4475 2815
rect 4435 2785 4445 2805
rect 4465 2785 4475 2805
rect 4435 2775 4475 2785
rect 4615 2805 4655 2815
rect 4615 2785 4625 2805
rect 4645 2785 4655 2805
rect 4615 2775 4655 2785
rect 4795 2805 4835 2815
rect 4795 2785 4805 2805
rect 4825 2785 4835 2805
rect 4795 2775 4835 2785
rect 4975 2805 5015 2815
rect 4975 2785 4985 2805
rect 5005 2785 5015 2805
rect 4975 2775 5015 2785
rect 11185 2810 11190 2830
rect 11210 2810 11230 2830
rect 11250 2810 11255 2830
rect 11185 2780 11255 2810
rect 11185 2760 11190 2780
rect 11210 2760 11230 2780
rect 11250 2760 11255 2780
rect 1266 2715 1296 2745
rect 2150 2710 2190 2750
rect 3175 2745 3215 2755
rect 3175 2725 3185 2745
rect 3205 2725 3215 2745
rect 3175 2715 3215 2725
rect 3355 2745 3395 2755
rect 3355 2725 3365 2745
rect 3385 2725 3395 2745
rect 3355 2715 3395 2725
rect 3535 2745 3575 2755
rect 3535 2725 3545 2745
rect 3565 2725 3575 2745
rect 3535 2715 3575 2725
rect 3715 2745 3755 2755
rect 3715 2725 3725 2745
rect 3745 2725 3755 2745
rect 3715 2715 3755 2725
rect 3895 2745 3935 2755
rect 3895 2725 3905 2745
rect 3925 2725 3935 2745
rect 3895 2715 3935 2725
rect 4075 2745 4115 2755
rect 4075 2725 4085 2745
rect 4105 2725 4115 2745
rect 4075 2715 4115 2725
rect 4255 2745 4295 2755
rect 4255 2725 4265 2745
rect 4285 2725 4295 2745
rect 4255 2715 4295 2725
rect 4435 2745 4475 2755
rect 4435 2725 4445 2745
rect 4465 2725 4475 2745
rect 4435 2715 4475 2725
rect 4615 2745 4655 2755
rect 4615 2725 4625 2745
rect 4645 2725 4655 2745
rect 4615 2715 4655 2725
rect 4795 2745 4835 2755
rect 4795 2725 4805 2745
rect 4825 2725 4835 2745
rect 4795 2715 4835 2725
rect 11185 2730 11255 2760
rect 650 2055 775 2700
rect 1330 2055 1455 2700
rect 2010 2055 2135 2700
rect 3185 2695 3205 2715
rect 3365 2695 3385 2715
rect 3545 2695 3565 2715
rect 3725 2695 3745 2715
rect 3905 2695 3925 2715
rect 4085 2695 4105 2715
rect 4265 2695 4285 2715
rect 4445 2695 4465 2715
rect 4625 2695 4645 2715
rect 4805 2695 4825 2715
rect 11185 2710 11190 2730
rect 11210 2710 11230 2730
rect 11250 2710 11255 2730
rect 3140 2685 3210 2695
rect 3140 2665 3145 2685
rect 3165 2665 3185 2685
rect 3205 2665 3210 2685
rect 3140 2635 3210 2665
rect 3140 2615 3145 2635
rect 3165 2615 3185 2635
rect 3205 2615 3210 2635
rect 3140 2585 3210 2615
rect 3140 2565 3145 2585
rect 3165 2565 3185 2585
rect 3205 2565 3210 2585
rect 3140 2535 3210 2565
rect 3140 2515 3145 2535
rect 3165 2515 3185 2535
rect 3205 2515 3210 2535
rect 3140 2485 3210 2515
rect 3140 2465 3145 2485
rect 3165 2465 3185 2485
rect 3205 2465 3210 2485
rect 3140 2435 3210 2465
rect 3140 2415 3145 2435
rect 3165 2415 3185 2435
rect 3205 2415 3210 2435
rect 3140 2405 3210 2415
rect 3270 2685 3300 2695
rect 3270 2665 3275 2685
rect 3295 2665 3300 2685
rect 3270 2635 3300 2665
rect 3270 2615 3275 2635
rect 3295 2615 3300 2635
rect 3270 2585 3300 2615
rect 3270 2565 3275 2585
rect 3295 2565 3300 2585
rect 3270 2535 3300 2565
rect 3270 2515 3275 2535
rect 3295 2515 3300 2535
rect 3270 2485 3300 2515
rect 3270 2465 3275 2485
rect 3295 2465 3300 2485
rect 3270 2435 3300 2465
rect 3270 2415 3275 2435
rect 3295 2415 3300 2435
rect 3270 2405 3300 2415
rect 3360 2685 3390 2695
rect 3360 2665 3365 2685
rect 3385 2665 3390 2685
rect 3360 2635 3390 2665
rect 3360 2615 3365 2635
rect 3385 2615 3390 2635
rect 3360 2585 3390 2615
rect 3360 2565 3365 2585
rect 3385 2565 3390 2585
rect 3360 2535 3390 2565
rect 3360 2515 3365 2535
rect 3385 2515 3390 2535
rect 3360 2485 3390 2515
rect 3360 2465 3365 2485
rect 3385 2465 3390 2485
rect 3360 2435 3390 2465
rect 3360 2415 3365 2435
rect 3385 2415 3390 2435
rect 3360 2405 3390 2415
rect 3450 2685 3480 2695
rect 3450 2665 3455 2685
rect 3475 2665 3480 2685
rect 3450 2635 3480 2665
rect 3450 2615 3455 2635
rect 3475 2615 3480 2635
rect 3450 2585 3480 2615
rect 3450 2565 3455 2585
rect 3475 2565 3480 2585
rect 3450 2535 3480 2565
rect 3450 2515 3455 2535
rect 3475 2515 3480 2535
rect 3450 2485 3480 2515
rect 3450 2465 3455 2485
rect 3475 2465 3480 2485
rect 3450 2435 3480 2465
rect 3450 2415 3455 2435
rect 3475 2415 3480 2435
rect 3450 2405 3480 2415
rect 3540 2685 3570 2695
rect 3540 2665 3545 2685
rect 3565 2665 3570 2685
rect 3540 2635 3570 2665
rect 3540 2615 3545 2635
rect 3565 2615 3570 2635
rect 3540 2585 3570 2615
rect 3540 2565 3545 2585
rect 3565 2565 3570 2585
rect 3540 2535 3570 2565
rect 3540 2515 3545 2535
rect 3565 2515 3570 2535
rect 3540 2485 3570 2515
rect 3540 2465 3545 2485
rect 3565 2465 3570 2485
rect 3540 2435 3570 2465
rect 3540 2415 3545 2435
rect 3565 2415 3570 2435
rect 3540 2405 3570 2415
rect 3630 2685 3660 2695
rect 3630 2665 3635 2685
rect 3655 2665 3660 2685
rect 3630 2635 3660 2665
rect 3630 2615 3635 2635
rect 3655 2615 3660 2635
rect 3630 2585 3660 2615
rect 3630 2565 3635 2585
rect 3655 2565 3660 2585
rect 3630 2535 3660 2565
rect 3630 2515 3635 2535
rect 3655 2515 3660 2535
rect 3630 2485 3660 2515
rect 3630 2465 3635 2485
rect 3655 2465 3660 2485
rect 3630 2435 3660 2465
rect 3630 2415 3635 2435
rect 3655 2415 3660 2435
rect 3630 2405 3660 2415
rect 3720 2685 3750 2695
rect 3720 2665 3725 2685
rect 3745 2665 3750 2685
rect 3720 2635 3750 2665
rect 3720 2615 3725 2635
rect 3745 2615 3750 2635
rect 3720 2585 3750 2615
rect 3720 2565 3725 2585
rect 3745 2565 3750 2585
rect 3720 2535 3750 2565
rect 3720 2515 3725 2535
rect 3745 2515 3750 2535
rect 3720 2485 3750 2515
rect 3720 2465 3725 2485
rect 3745 2465 3750 2485
rect 3720 2435 3750 2465
rect 3720 2415 3725 2435
rect 3745 2415 3750 2435
rect 3720 2405 3750 2415
rect 3810 2685 3840 2695
rect 3810 2665 3815 2685
rect 3835 2665 3840 2685
rect 3810 2635 3840 2665
rect 3810 2615 3815 2635
rect 3835 2615 3840 2635
rect 3810 2585 3840 2615
rect 3810 2565 3815 2585
rect 3835 2565 3840 2585
rect 3810 2535 3840 2565
rect 3810 2515 3815 2535
rect 3835 2515 3840 2535
rect 3810 2485 3840 2515
rect 3810 2465 3815 2485
rect 3835 2465 3840 2485
rect 3810 2435 3840 2465
rect 3810 2415 3815 2435
rect 3835 2415 3840 2435
rect 3810 2405 3840 2415
rect 3900 2685 3930 2695
rect 3900 2665 3905 2685
rect 3925 2665 3930 2685
rect 3900 2635 3930 2665
rect 3900 2615 3905 2635
rect 3925 2615 3930 2635
rect 3900 2585 3930 2615
rect 3900 2565 3905 2585
rect 3925 2565 3930 2585
rect 3900 2535 3930 2565
rect 3900 2515 3905 2535
rect 3925 2515 3930 2535
rect 3900 2485 3930 2515
rect 3900 2465 3905 2485
rect 3925 2465 3930 2485
rect 3900 2435 3930 2465
rect 3900 2415 3905 2435
rect 3925 2415 3930 2435
rect 3900 2405 3930 2415
rect 3990 2685 4020 2695
rect 3990 2665 3995 2685
rect 4015 2665 4020 2685
rect 3990 2635 4020 2665
rect 3990 2615 3995 2635
rect 4015 2615 4020 2635
rect 3990 2585 4020 2615
rect 3990 2565 3995 2585
rect 4015 2565 4020 2585
rect 3990 2535 4020 2565
rect 3990 2515 3995 2535
rect 4015 2515 4020 2535
rect 3990 2485 4020 2515
rect 3990 2465 3995 2485
rect 4015 2465 4020 2485
rect 3990 2435 4020 2465
rect 3990 2415 3995 2435
rect 4015 2415 4020 2435
rect 3990 2405 4020 2415
rect 4080 2685 4110 2695
rect 4080 2665 4085 2685
rect 4105 2665 4110 2685
rect 4080 2635 4110 2665
rect 4080 2615 4085 2635
rect 4105 2615 4110 2635
rect 4080 2585 4110 2615
rect 4080 2565 4085 2585
rect 4105 2565 4110 2585
rect 4080 2535 4110 2565
rect 4080 2515 4085 2535
rect 4105 2515 4110 2535
rect 4080 2485 4110 2515
rect 4080 2465 4085 2485
rect 4105 2465 4110 2485
rect 4080 2435 4110 2465
rect 4080 2415 4085 2435
rect 4105 2415 4110 2435
rect 4080 2405 4110 2415
rect 4170 2685 4200 2695
rect 4170 2665 4175 2685
rect 4195 2665 4200 2685
rect 4170 2635 4200 2665
rect 4170 2615 4175 2635
rect 4195 2615 4200 2635
rect 4170 2585 4200 2615
rect 4170 2565 4175 2585
rect 4195 2565 4200 2585
rect 4170 2535 4200 2565
rect 4170 2515 4175 2535
rect 4195 2515 4200 2535
rect 4170 2485 4200 2515
rect 4170 2465 4175 2485
rect 4195 2465 4200 2485
rect 4170 2435 4200 2465
rect 4170 2415 4175 2435
rect 4195 2415 4200 2435
rect 4170 2405 4200 2415
rect 4260 2685 4290 2695
rect 4260 2665 4265 2685
rect 4285 2665 4290 2685
rect 4260 2635 4290 2665
rect 4260 2615 4265 2635
rect 4285 2615 4290 2635
rect 4260 2585 4290 2615
rect 4260 2565 4265 2585
rect 4285 2565 4290 2585
rect 4260 2535 4290 2565
rect 4260 2515 4265 2535
rect 4285 2515 4290 2535
rect 4260 2485 4290 2515
rect 4260 2465 4265 2485
rect 4285 2465 4290 2485
rect 4260 2435 4290 2465
rect 4260 2415 4265 2435
rect 4285 2415 4290 2435
rect 4260 2405 4290 2415
rect 4350 2685 4380 2695
rect 4350 2665 4355 2685
rect 4375 2665 4380 2685
rect 4350 2635 4380 2665
rect 4350 2615 4355 2635
rect 4375 2615 4380 2635
rect 4350 2585 4380 2615
rect 4350 2565 4355 2585
rect 4375 2565 4380 2585
rect 4350 2535 4380 2565
rect 4350 2515 4355 2535
rect 4375 2515 4380 2535
rect 4350 2485 4380 2515
rect 4350 2465 4355 2485
rect 4375 2465 4380 2485
rect 4350 2435 4380 2465
rect 4350 2415 4355 2435
rect 4375 2415 4380 2435
rect 4350 2405 4380 2415
rect 4440 2685 4470 2695
rect 4440 2665 4445 2685
rect 4465 2665 4470 2685
rect 4440 2635 4470 2665
rect 4440 2615 4445 2635
rect 4465 2615 4470 2635
rect 4440 2585 4470 2615
rect 4440 2565 4445 2585
rect 4465 2565 4470 2585
rect 4440 2535 4470 2565
rect 4440 2515 4445 2535
rect 4465 2515 4470 2535
rect 4440 2485 4470 2515
rect 4440 2465 4445 2485
rect 4465 2465 4470 2485
rect 4440 2435 4470 2465
rect 4440 2415 4445 2435
rect 4465 2415 4470 2435
rect 4440 2405 4470 2415
rect 4530 2685 4560 2695
rect 4530 2665 4535 2685
rect 4555 2665 4560 2685
rect 4530 2635 4560 2665
rect 4530 2615 4535 2635
rect 4555 2615 4560 2635
rect 4530 2585 4560 2615
rect 4530 2565 4535 2585
rect 4555 2565 4560 2585
rect 4530 2535 4560 2565
rect 4530 2515 4535 2535
rect 4555 2515 4560 2535
rect 4530 2485 4560 2515
rect 4530 2465 4535 2485
rect 4555 2465 4560 2485
rect 4530 2435 4560 2465
rect 4530 2415 4535 2435
rect 4555 2415 4560 2435
rect 4530 2405 4560 2415
rect 4620 2685 4650 2695
rect 4620 2665 4625 2685
rect 4645 2665 4650 2685
rect 4620 2635 4650 2665
rect 4620 2615 4625 2635
rect 4645 2615 4650 2635
rect 4620 2585 4650 2615
rect 4620 2565 4625 2585
rect 4645 2565 4650 2585
rect 4620 2535 4650 2565
rect 4620 2515 4625 2535
rect 4645 2515 4650 2535
rect 4620 2485 4650 2515
rect 4620 2465 4625 2485
rect 4645 2465 4650 2485
rect 4620 2435 4650 2465
rect 4620 2415 4625 2435
rect 4645 2415 4650 2435
rect 4620 2405 4650 2415
rect 4710 2685 4740 2695
rect 4710 2665 4715 2685
rect 4735 2665 4740 2685
rect 4710 2635 4740 2665
rect 4710 2615 4715 2635
rect 4735 2615 4740 2635
rect 4710 2585 4740 2615
rect 4710 2565 4715 2585
rect 4735 2565 4740 2585
rect 4710 2535 4740 2565
rect 4710 2515 4715 2535
rect 4735 2515 4740 2535
rect 4710 2485 4740 2515
rect 4710 2465 4715 2485
rect 4735 2465 4740 2485
rect 4710 2435 4740 2465
rect 4710 2415 4715 2435
rect 4735 2415 4740 2435
rect 4710 2405 4740 2415
rect 4800 2685 4870 2695
rect 4800 2665 4805 2685
rect 4825 2665 4845 2685
rect 4865 2665 4870 2685
rect 11185 2680 11255 2710
rect 4800 2635 4870 2665
rect 9735 2665 9775 2675
rect 9735 2645 9745 2665
rect 9765 2645 9775 2665
rect 9735 2635 9775 2645
rect 9845 2665 9885 2675
rect 9845 2645 9855 2665
rect 9875 2645 9885 2665
rect 9845 2635 9885 2645
rect 9955 2665 9995 2675
rect 9955 2645 9965 2665
rect 9985 2645 9995 2665
rect 9955 2635 9995 2645
rect 10065 2665 10105 2675
rect 10065 2645 10075 2665
rect 10095 2645 10105 2665
rect 10065 2635 10105 2645
rect 10175 2665 10215 2675
rect 10175 2645 10185 2665
rect 10205 2645 10215 2665
rect 10175 2635 10215 2645
rect 10285 2665 10325 2675
rect 10285 2645 10295 2665
rect 10315 2645 10325 2665
rect 10285 2635 10325 2645
rect 10395 2665 10435 2675
rect 10395 2645 10405 2665
rect 10425 2645 10435 2665
rect 10395 2635 10435 2645
rect 10505 2665 10545 2675
rect 10505 2645 10515 2665
rect 10535 2645 10545 2665
rect 10505 2635 10545 2645
rect 10615 2665 10655 2675
rect 10615 2645 10625 2665
rect 10645 2645 10655 2665
rect 10615 2635 10655 2645
rect 10725 2665 10765 2675
rect 10725 2645 10735 2665
rect 10755 2645 10765 2665
rect 10725 2635 10765 2645
rect 10835 2665 10875 2675
rect 10835 2645 10845 2665
rect 10865 2645 10875 2665
rect 10835 2635 10875 2645
rect 11185 2660 11190 2680
rect 11210 2660 11230 2680
rect 11250 2660 11255 2680
rect 4800 2615 4805 2635
rect 4825 2615 4845 2635
rect 4865 2615 4870 2635
rect 9745 2615 9765 2635
rect 9855 2615 9875 2635
rect 9965 2615 9985 2635
rect 10075 2615 10095 2635
rect 10185 2615 10205 2635
rect 10295 2615 10315 2635
rect 10405 2615 10425 2635
rect 10515 2615 10535 2635
rect 10625 2615 10645 2635
rect 10735 2615 10755 2635
rect 10845 2615 10865 2635
rect 11185 2630 11255 2660
rect 4800 2585 4870 2615
rect 4800 2565 4805 2585
rect 4825 2565 4845 2585
rect 4865 2565 4870 2585
rect 4800 2535 4870 2565
rect 4800 2515 4805 2535
rect 4825 2515 4845 2535
rect 4865 2515 4870 2535
rect 9645 2605 9715 2615
rect 9645 2585 9650 2605
rect 9670 2585 9690 2605
rect 9710 2585 9715 2605
rect 9645 2555 9715 2585
rect 9645 2535 9650 2555
rect 9670 2535 9690 2555
rect 9710 2535 9715 2555
rect 9645 2525 9715 2535
rect 9740 2605 9770 2615
rect 9740 2585 9745 2605
rect 9765 2585 9770 2605
rect 9740 2555 9770 2585
rect 9740 2535 9745 2555
rect 9765 2535 9770 2555
rect 9740 2525 9770 2535
rect 9795 2605 9825 2615
rect 9795 2585 9800 2605
rect 9820 2585 9825 2605
rect 9795 2555 9825 2585
rect 9795 2535 9800 2555
rect 9820 2535 9825 2555
rect 9795 2525 9825 2535
rect 9850 2605 9880 2615
rect 9850 2585 9855 2605
rect 9875 2585 9880 2605
rect 9850 2555 9880 2585
rect 9850 2535 9855 2555
rect 9875 2535 9880 2555
rect 9850 2525 9880 2535
rect 9905 2605 9935 2615
rect 9905 2585 9910 2605
rect 9930 2585 9935 2605
rect 9905 2555 9935 2585
rect 9905 2535 9910 2555
rect 9930 2535 9935 2555
rect 9905 2525 9935 2535
rect 9960 2605 9990 2615
rect 9960 2585 9965 2605
rect 9985 2585 9990 2605
rect 9960 2555 9990 2585
rect 9960 2535 9965 2555
rect 9985 2535 9990 2555
rect 9960 2525 9990 2535
rect 10015 2605 10045 2615
rect 10015 2585 10020 2605
rect 10040 2585 10045 2605
rect 10015 2555 10045 2585
rect 10015 2535 10020 2555
rect 10040 2535 10045 2555
rect 10015 2525 10045 2535
rect 10070 2605 10100 2615
rect 10070 2585 10075 2605
rect 10095 2585 10100 2605
rect 10070 2555 10100 2585
rect 10070 2535 10075 2555
rect 10095 2535 10100 2555
rect 10070 2525 10100 2535
rect 10125 2605 10155 2615
rect 10125 2585 10130 2605
rect 10150 2585 10155 2605
rect 10125 2555 10155 2585
rect 10125 2535 10130 2555
rect 10150 2535 10155 2555
rect 10125 2525 10155 2535
rect 10180 2605 10210 2615
rect 10180 2585 10185 2605
rect 10205 2585 10210 2605
rect 10180 2555 10210 2585
rect 10180 2535 10185 2555
rect 10205 2535 10210 2555
rect 10180 2525 10210 2535
rect 10235 2605 10265 2615
rect 10235 2585 10240 2605
rect 10260 2585 10265 2605
rect 10235 2555 10265 2585
rect 10235 2535 10240 2555
rect 10260 2535 10265 2555
rect 10235 2525 10265 2535
rect 10290 2605 10320 2615
rect 10290 2585 10295 2605
rect 10315 2585 10320 2605
rect 10290 2555 10320 2585
rect 10290 2535 10295 2555
rect 10315 2535 10320 2555
rect 10290 2525 10320 2535
rect 10345 2605 10375 2615
rect 10345 2585 10350 2605
rect 10370 2585 10375 2605
rect 10345 2555 10375 2585
rect 10345 2535 10350 2555
rect 10370 2535 10375 2555
rect 10345 2525 10375 2535
rect 10400 2605 10430 2615
rect 10400 2585 10405 2605
rect 10425 2585 10430 2605
rect 10400 2555 10430 2585
rect 10400 2535 10405 2555
rect 10425 2535 10430 2555
rect 10400 2525 10430 2535
rect 10455 2605 10485 2615
rect 10455 2585 10460 2605
rect 10480 2585 10485 2605
rect 10455 2555 10485 2585
rect 10455 2535 10460 2555
rect 10480 2535 10485 2555
rect 10455 2525 10485 2535
rect 10510 2605 10540 2615
rect 10510 2585 10515 2605
rect 10535 2585 10540 2605
rect 10510 2555 10540 2585
rect 10510 2535 10515 2555
rect 10535 2535 10540 2555
rect 10510 2525 10540 2535
rect 10565 2605 10595 2615
rect 10565 2585 10570 2605
rect 10590 2585 10595 2605
rect 10565 2555 10595 2585
rect 10565 2535 10570 2555
rect 10590 2535 10595 2555
rect 10565 2525 10595 2535
rect 10620 2605 10650 2615
rect 10620 2585 10625 2605
rect 10645 2585 10650 2605
rect 10620 2555 10650 2585
rect 10620 2535 10625 2555
rect 10645 2535 10650 2555
rect 10620 2525 10650 2535
rect 10675 2605 10705 2615
rect 10675 2585 10680 2605
rect 10700 2585 10705 2605
rect 10675 2555 10705 2585
rect 10675 2535 10680 2555
rect 10700 2535 10705 2555
rect 10675 2525 10705 2535
rect 10730 2605 10760 2615
rect 10730 2585 10735 2605
rect 10755 2585 10760 2605
rect 10730 2555 10760 2585
rect 10730 2535 10735 2555
rect 10755 2535 10760 2555
rect 10730 2525 10760 2535
rect 10785 2605 10815 2615
rect 10785 2585 10790 2605
rect 10810 2585 10815 2605
rect 10785 2555 10815 2585
rect 10785 2535 10790 2555
rect 10810 2535 10815 2555
rect 10785 2525 10815 2535
rect 10840 2605 10870 2615
rect 10840 2585 10845 2605
rect 10865 2585 10870 2605
rect 10840 2555 10870 2585
rect 10840 2535 10845 2555
rect 10865 2535 10870 2555
rect 10840 2525 10870 2535
rect 10895 2605 10965 2615
rect 10895 2585 10900 2605
rect 10920 2585 10940 2605
rect 10960 2585 10965 2605
rect 10895 2555 10965 2585
rect 10895 2535 10900 2555
rect 10920 2535 10940 2555
rect 10960 2535 10965 2555
rect 10895 2525 10965 2535
rect 11185 2610 11190 2630
rect 11210 2610 11230 2630
rect 11250 2610 11255 2630
rect 11185 2580 11255 2610
rect 11185 2560 11190 2580
rect 11210 2560 11230 2580
rect 11250 2560 11255 2580
rect 11185 2530 11255 2560
rect 4800 2485 4870 2515
rect 9650 2505 9670 2525
rect 9800 2505 9820 2525
rect 9910 2505 9930 2525
rect 10020 2505 10040 2525
rect 10130 2505 10150 2525
rect 10240 2505 10260 2525
rect 10350 2505 10370 2525
rect 10460 2505 10480 2525
rect 10570 2505 10590 2525
rect 10680 2505 10700 2525
rect 10790 2505 10810 2525
rect 10940 2505 10960 2525
rect 11185 2510 11190 2530
rect 11210 2510 11230 2530
rect 11250 2510 11255 2530
rect 4800 2465 4805 2485
rect 4825 2465 4845 2485
rect 4865 2465 4870 2485
rect 9640 2495 9680 2505
rect 9640 2475 9650 2495
rect 9670 2475 9680 2495
rect 9640 2465 9680 2475
rect 9790 2495 9830 2505
rect 9790 2475 9800 2495
rect 9820 2475 9830 2495
rect 9790 2465 9830 2475
rect 9900 2495 9940 2505
rect 9900 2475 9910 2495
rect 9930 2475 9940 2495
rect 9900 2465 9940 2475
rect 10010 2495 10050 2505
rect 10010 2475 10020 2495
rect 10040 2475 10050 2495
rect 10010 2465 10050 2475
rect 10120 2495 10160 2505
rect 10120 2475 10130 2495
rect 10150 2475 10160 2495
rect 10120 2465 10160 2475
rect 10230 2495 10270 2505
rect 10230 2475 10240 2495
rect 10260 2475 10270 2495
rect 10230 2465 10270 2475
rect 10340 2495 10380 2505
rect 10340 2475 10350 2495
rect 10370 2475 10380 2495
rect 10340 2465 10380 2475
rect 10450 2495 10490 2505
rect 10450 2475 10460 2495
rect 10480 2475 10490 2495
rect 10450 2465 10490 2475
rect 10560 2495 10600 2505
rect 10560 2475 10570 2495
rect 10590 2475 10600 2495
rect 10560 2465 10600 2475
rect 10670 2495 10710 2505
rect 10670 2475 10680 2495
rect 10700 2475 10710 2495
rect 10670 2465 10710 2475
rect 10780 2495 10820 2505
rect 10780 2475 10790 2495
rect 10810 2475 10820 2495
rect 10780 2465 10820 2475
rect 10930 2495 10970 2505
rect 11185 2500 11255 2510
rect 11285 2880 11315 2890
rect 11285 2860 11290 2880
rect 11310 2860 11315 2880
rect 11285 2830 11315 2860
rect 11285 2810 11290 2830
rect 11310 2810 11315 2830
rect 11285 2780 11315 2810
rect 11285 2760 11290 2780
rect 11310 2760 11315 2780
rect 11285 2730 11315 2760
rect 11285 2710 11290 2730
rect 11310 2710 11315 2730
rect 11285 2680 11315 2710
rect 11285 2660 11290 2680
rect 11310 2660 11315 2680
rect 11285 2630 11315 2660
rect 11285 2610 11290 2630
rect 11310 2610 11315 2630
rect 11285 2580 11315 2610
rect 11285 2560 11290 2580
rect 11310 2560 11315 2580
rect 11285 2530 11315 2560
rect 11285 2510 11290 2530
rect 11310 2510 11315 2530
rect 11285 2500 11315 2510
rect 11345 2880 11375 2890
rect 11345 2860 11350 2880
rect 11370 2860 11375 2880
rect 11345 2830 11375 2860
rect 11345 2810 11350 2830
rect 11370 2810 11375 2830
rect 11345 2780 11375 2810
rect 11345 2760 11350 2780
rect 11370 2760 11375 2780
rect 11345 2730 11375 2760
rect 11345 2710 11350 2730
rect 11370 2710 11375 2730
rect 11345 2680 11375 2710
rect 11345 2660 11350 2680
rect 11370 2660 11375 2680
rect 11345 2630 11375 2660
rect 11345 2610 11350 2630
rect 11370 2610 11375 2630
rect 11345 2580 11375 2610
rect 11345 2560 11350 2580
rect 11370 2560 11375 2580
rect 11345 2530 11375 2560
rect 11345 2510 11350 2530
rect 11370 2510 11375 2530
rect 11345 2500 11375 2510
rect 11405 2880 11435 2890
rect 11405 2860 11410 2880
rect 11430 2860 11435 2880
rect 11405 2830 11435 2860
rect 11405 2810 11410 2830
rect 11430 2810 11435 2830
rect 11405 2780 11435 2810
rect 11405 2760 11410 2780
rect 11430 2760 11435 2780
rect 11405 2730 11435 2760
rect 11405 2710 11410 2730
rect 11430 2710 11435 2730
rect 11405 2680 11435 2710
rect 11405 2660 11410 2680
rect 11430 2660 11435 2680
rect 11405 2630 11435 2660
rect 11405 2610 11410 2630
rect 11430 2610 11435 2630
rect 11405 2580 11435 2610
rect 11405 2560 11410 2580
rect 11430 2560 11435 2580
rect 11405 2530 11435 2560
rect 11405 2510 11410 2530
rect 11430 2510 11435 2530
rect 11405 2500 11435 2510
rect 11465 2880 11495 2890
rect 11465 2860 11470 2880
rect 11490 2860 11495 2880
rect 11465 2830 11495 2860
rect 11465 2810 11470 2830
rect 11490 2810 11495 2830
rect 11465 2780 11495 2810
rect 11465 2760 11470 2780
rect 11490 2760 11495 2780
rect 11465 2730 11495 2760
rect 11465 2710 11470 2730
rect 11490 2710 11495 2730
rect 11465 2680 11495 2710
rect 11465 2660 11470 2680
rect 11490 2660 11495 2680
rect 11465 2630 11495 2660
rect 11465 2610 11470 2630
rect 11490 2610 11495 2630
rect 11465 2580 11495 2610
rect 11465 2560 11470 2580
rect 11490 2560 11495 2580
rect 11465 2530 11495 2560
rect 11465 2510 11470 2530
rect 11490 2510 11495 2530
rect 11465 2500 11495 2510
rect 11525 2880 11555 2890
rect 11525 2860 11530 2880
rect 11550 2860 11555 2880
rect 11525 2830 11555 2860
rect 11525 2810 11530 2830
rect 11550 2810 11555 2830
rect 11525 2780 11555 2810
rect 11525 2760 11530 2780
rect 11550 2760 11555 2780
rect 11525 2730 11555 2760
rect 11525 2710 11530 2730
rect 11550 2710 11555 2730
rect 11525 2680 11555 2710
rect 11525 2660 11530 2680
rect 11550 2660 11555 2680
rect 11525 2630 11555 2660
rect 11525 2610 11530 2630
rect 11550 2610 11555 2630
rect 11525 2580 11555 2610
rect 11525 2560 11530 2580
rect 11550 2560 11555 2580
rect 11525 2530 11555 2560
rect 11525 2510 11530 2530
rect 11550 2510 11555 2530
rect 11525 2500 11555 2510
rect 11585 2880 11615 2890
rect 11585 2860 11590 2880
rect 11610 2860 11615 2880
rect 11585 2830 11615 2860
rect 11585 2810 11590 2830
rect 11610 2810 11615 2830
rect 11585 2780 11615 2810
rect 11585 2760 11590 2780
rect 11610 2760 11615 2780
rect 11585 2730 11615 2760
rect 11585 2710 11590 2730
rect 11610 2710 11615 2730
rect 11585 2680 11615 2710
rect 11585 2660 11590 2680
rect 11610 2660 11615 2680
rect 11585 2630 11615 2660
rect 11585 2610 11590 2630
rect 11610 2610 11615 2630
rect 11585 2580 11615 2610
rect 11585 2560 11590 2580
rect 11610 2560 11615 2580
rect 11585 2530 11615 2560
rect 11585 2510 11590 2530
rect 11610 2510 11615 2530
rect 11585 2500 11615 2510
rect 11645 2880 11675 2890
rect 11645 2860 11650 2880
rect 11670 2860 11675 2880
rect 11645 2830 11675 2860
rect 11645 2810 11650 2830
rect 11670 2810 11675 2830
rect 11645 2780 11675 2810
rect 11645 2760 11650 2780
rect 11670 2760 11675 2780
rect 11645 2730 11675 2760
rect 11645 2710 11650 2730
rect 11670 2710 11675 2730
rect 11645 2680 11675 2710
rect 11645 2660 11650 2680
rect 11670 2660 11675 2680
rect 11645 2630 11675 2660
rect 11645 2610 11650 2630
rect 11670 2610 11675 2630
rect 11645 2580 11675 2610
rect 11645 2560 11650 2580
rect 11670 2560 11675 2580
rect 11645 2530 11675 2560
rect 11645 2510 11650 2530
rect 11670 2510 11675 2530
rect 11645 2500 11675 2510
rect 11705 2880 11735 2890
rect 11705 2860 11710 2880
rect 11730 2860 11735 2880
rect 11705 2830 11735 2860
rect 11705 2810 11710 2830
rect 11730 2810 11735 2830
rect 11705 2780 11735 2810
rect 11705 2760 11710 2780
rect 11730 2760 11735 2780
rect 11705 2730 11735 2760
rect 11705 2710 11710 2730
rect 11730 2710 11735 2730
rect 11705 2680 11735 2710
rect 11705 2660 11710 2680
rect 11730 2660 11735 2680
rect 11705 2630 11735 2660
rect 11705 2610 11710 2630
rect 11730 2610 11735 2630
rect 11705 2580 11735 2610
rect 11705 2560 11710 2580
rect 11730 2560 11735 2580
rect 11705 2530 11735 2560
rect 11705 2510 11710 2530
rect 11730 2510 11735 2530
rect 11705 2500 11735 2510
rect 11765 2880 11795 2890
rect 11765 2860 11770 2880
rect 11790 2860 11795 2880
rect 11765 2830 11795 2860
rect 11765 2810 11770 2830
rect 11790 2810 11795 2830
rect 11765 2780 11795 2810
rect 11765 2760 11770 2780
rect 11790 2760 11795 2780
rect 11765 2730 11795 2760
rect 11765 2710 11770 2730
rect 11790 2710 11795 2730
rect 11765 2680 11795 2710
rect 11765 2660 11770 2680
rect 11790 2660 11795 2680
rect 11765 2630 11795 2660
rect 11765 2610 11770 2630
rect 11790 2610 11795 2630
rect 11765 2580 11795 2610
rect 11765 2560 11770 2580
rect 11790 2560 11795 2580
rect 11765 2530 11795 2560
rect 11765 2510 11770 2530
rect 11790 2510 11795 2530
rect 11765 2500 11795 2510
rect 11825 2880 11855 2890
rect 11825 2860 11830 2880
rect 11850 2860 11855 2880
rect 11825 2830 11855 2860
rect 11825 2810 11830 2830
rect 11850 2810 11855 2830
rect 11825 2780 11855 2810
rect 11825 2760 11830 2780
rect 11850 2760 11855 2780
rect 11825 2730 11855 2760
rect 11825 2710 11830 2730
rect 11850 2710 11855 2730
rect 11825 2680 11855 2710
rect 11825 2660 11830 2680
rect 11850 2660 11855 2680
rect 11825 2630 11855 2660
rect 11825 2610 11830 2630
rect 11850 2610 11855 2630
rect 11825 2580 11855 2610
rect 11825 2560 11830 2580
rect 11850 2560 11855 2580
rect 11825 2530 11855 2560
rect 11825 2510 11830 2530
rect 11850 2510 11855 2530
rect 11825 2500 11855 2510
rect 11885 2880 11915 2890
rect 11885 2860 11890 2880
rect 11910 2860 11915 2880
rect 11885 2830 11915 2860
rect 11885 2810 11890 2830
rect 11910 2810 11915 2830
rect 11885 2780 11915 2810
rect 11885 2760 11890 2780
rect 11910 2760 11915 2780
rect 11885 2730 11915 2760
rect 11885 2710 11890 2730
rect 11910 2710 11915 2730
rect 11885 2680 11915 2710
rect 11885 2660 11890 2680
rect 11910 2660 11915 2680
rect 11885 2630 11915 2660
rect 11885 2610 11890 2630
rect 11910 2610 11915 2630
rect 11885 2580 11915 2610
rect 11885 2560 11890 2580
rect 11910 2560 11915 2580
rect 11885 2530 11915 2560
rect 11885 2510 11890 2530
rect 11910 2510 11915 2530
rect 11885 2500 11915 2510
rect 11945 2880 11975 2890
rect 11945 2860 11950 2880
rect 11970 2860 11975 2880
rect 11945 2830 11975 2860
rect 11945 2810 11950 2830
rect 11970 2810 11975 2830
rect 11945 2780 11975 2810
rect 11945 2760 11950 2780
rect 11970 2760 11975 2780
rect 11945 2730 11975 2760
rect 11945 2710 11950 2730
rect 11970 2710 11975 2730
rect 11945 2680 11975 2710
rect 11945 2660 11950 2680
rect 11970 2660 11975 2680
rect 11945 2630 11975 2660
rect 11945 2610 11950 2630
rect 11970 2610 11975 2630
rect 11945 2580 11975 2610
rect 11945 2560 11950 2580
rect 11970 2560 11975 2580
rect 11945 2530 11975 2560
rect 11945 2510 11950 2530
rect 11970 2510 11975 2530
rect 11945 2500 11975 2510
rect 12005 2880 12035 2890
rect 12005 2860 12010 2880
rect 12030 2860 12035 2880
rect 12005 2830 12035 2860
rect 12005 2810 12010 2830
rect 12030 2810 12035 2830
rect 12005 2780 12035 2810
rect 12005 2760 12010 2780
rect 12030 2760 12035 2780
rect 12005 2730 12035 2760
rect 12005 2710 12010 2730
rect 12030 2710 12035 2730
rect 12005 2680 12035 2710
rect 12005 2660 12010 2680
rect 12030 2660 12035 2680
rect 12005 2630 12035 2660
rect 12005 2610 12010 2630
rect 12030 2610 12035 2630
rect 12005 2580 12035 2610
rect 12005 2560 12010 2580
rect 12030 2560 12035 2580
rect 12005 2530 12035 2560
rect 12005 2510 12010 2530
rect 12030 2510 12035 2530
rect 12005 2500 12035 2510
rect 12065 2880 12095 2890
rect 12065 2860 12070 2880
rect 12090 2860 12095 2880
rect 12065 2830 12095 2860
rect 12065 2810 12070 2830
rect 12090 2810 12095 2830
rect 12065 2780 12095 2810
rect 12065 2760 12070 2780
rect 12090 2760 12095 2780
rect 12065 2730 12095 2760
rect 12065 2710 12070 2730
rect 12090 2710 12095 2730
rect 12065 2680 12095 2710
rect 12065 2660 12070 2680
rect 12090 2660 12095 2680
rect 12065 2630 12095 2660
rect 12065 2610 12070 2630
rect 12090 2610 12095 2630
rect 12065 2580 12095 2610
rect 12065 2560 12070 2580
rect 12090 2560 12095 2580
rect 12065 2530 12095 2560
rect 12065 2510 12070 2530
rect 12090 2510 12095 2530
rect 12065 2500 12095 2510
rect 12125 2880 12155 2890
rect 12125 2860 12130 2880
rect 12150 2860 12155 2880
rect 12125 2830 12155 2860
rect 12125 2810 12130 2830
rect 12150 2810 12155 2830
rect 12125 2780 12155 2810
rect 12125 2760 12130 2780
rect 12150 2760 12155 2780
rect 12125 2730 12155 2760
rect 12125 2710 12130 2730
rect 12150 2710 12155 2730
rect 12125 2680 12155 2710
rect 12125 2660 12130 2680
rect 12150 2660 12155 2680
rect 12125 2630 12155 2660
rect 12125 2610 12130 2630
rect 12150 2610 12155 2630
rect 12125 2580 12155 2610
rect 12125 2560 12130 2580
rect 12150 2560 12155 2580
rect 12125 2530 12155 2560
rect 12125 2510 12130 2530
rect 12150 2510 12155 2530
rect 12125 2500 12155 2510
rect 12185 2880 12215 2890
rect 12185 2860 12190 2880
rect 12210 2860 12215 2880
rect 12185 2830 12215 2860
rect 12185 2810 12190 2830
rect 12210 2810 12215 2830
rect 12185 2780 12215 2810
rect 12185 2760 12190 2780
rect 12210 2760 12215 2780
rect 12185 2730 12215 2760
rect 12185 2710 12190 2730
rect 12210 2710 12215 2730
rect 12185 2680 12215 2710
rect 12185 2660 12190 2680
rect 12210 2660 12215 2680
rect 12185 2630 12215 2660
rect 12185 2610 12190 2630
rect 12210 2610 12215 2630
rect 12185 2580 12215 2610
rect 12185 2560 12190 2580
rect 12210 2560 12215 2580
rect 12185 2530 12215 2560
rect 12185 2510 12190 2530
rect 12210 2510 12215 2530
rect 12185 2500 12215 2510
rect 12245 2880 12275 2890
rect 12245 2860 12250 2880
rect 12270 2860 12275 2880
rect 12245 2830 12275 2860
rect 12245 2810 12250 2830
rect 12270 2810 12275 2830
rect 12245 2780 12275 2810
rect 12245 2760 12250 2780
rect 12270 2760 12275 2780
rect 12245 2730 12275 2760
rect 12245 2710 12250 2730
rect 12270 2710 12275 2730
rect 12245 2680 12275 2710
rect 12245 2660 12250 2680
rect 12270 2660 12275 2680
rect 12245 2630 12275 2660
rect 12245 2610 12250 2630
rect 12270 2610 12275 2630
rect 12245 2580 12275 2610
rect 12245 2560 12250 2580
rect 12270 2560 12275 2580
rect 12245 2530 12275 2560
rect 12245 2510 12250 2530
rect 12270 2510 12275 2530
rect 12245 2500 12275 2510
rect 12305 2880 12335 2890
rect 12305 2860 12310 2880
rect 12330 2860 12335 2880
rect 12305 2830 12335 2860
rect 12305 2810 12310 2830
rect 12330 2810 12335 2830
rect 12305 2780 12335 2810
rect 12305 2760 12310 2780
rect 12330 2760 12335 2780
rect 12305 2730 12335 2760
rect 12305 2710 12310 2730
rect 12330 2710 12335 2730
rect 12305 2680 12335 2710
rect 12305 2660 12310 2680
rect 12330 2660 12335 2680
rect 12305 2630 12335 2660
rect 12305 2610 12310 2630
rect 12330 2610 12335 2630
rect 12305 2580 12335 2610
rect 12305 2560 12310 2580
rect 12330 2560 12335 2580
rect 12305 2530 12335 2560
rect 12305 2510 12310 2530
rect 12330 2510 12335 2530
rect 12305 2500 12335 2510
rect 12365 2880 12395 2890
rect 12365 2860 12370 2880
rect 12390 2860 12395 2880
rect 12365 2830 12395 2860
rect 12365 2810 12370 2830
rect 12390 2810 12395 2830
rect 12365 2780 12395 2810
rect 12365 2760 12370 2780
rect 12390 2760 12395 2780
rect 12365 2730 12395 2760
rect 12365 2710 12370 2730
rect 12390 2710 12395 2730
rect 12365 2680 12395 2710
rect 12365 2660 12370 2680
rect 12390 2660 12395 2680
rect 12365 2630 12395 2660
rect 12365 2610 12370 2630
rect 12390 2610 12395 2630
rect 12365 2580 12395 2610
rect 12365 2560 12370 2580
rect 12390 2560 12395 2580
rect 12365 2530 12395 2560
rect 12365 2510 12370 2530
rect 12390 2510 12395 2530
rect 12365 2500 12395 2510
rect 12425 2880 12455 2890
rect 12425 2860 12430 2880
rect 12450 2860 12455 2880
rect 12425 2830 12455 2860
rect 12425 2810 12430 2830
rect 12450 2810 12455 2830
rect 12425 2780 12455 2810
rect 12425 2760 12430 2780
rect 12450 2760 12455 2780
rect 12425 2730 12455 2760
rect 12425 2710 12430 2730
rect 12450 2710 12455 2730
rect 12425 2680 12455 2710
rect 12425 2660 12430 2680
rect 12450 2660 12455 2680
rect 12425 2630 12455 2660
rect 12425 2610 12430 2630
rect 12450 2610 12455 2630
rect 12425 2580 12455 2610
rect 12425 2560 12430 2580
rect 12450 2560 12455 2580
rect 12425 2530 12455 2560
rect 12425 2510 12430 2530
rect 12450 2510 12455 2530
rect 12425 2500 12455 2510
rect 12485 2880 12515 2890
rect 12485 2860 12490 2880
rect 12510 2860 12515 2880
rect 12485 2830 12515 2860
rect 12485 2810 12490 2830
rect 12510 2810 12515 2830
rect 12485 2780 12515 2810
rect 12485 2760 12490 2780
rect 12510 2760 12515 2780
rect 12485 2730 12515 2760
rect 12485 2710 12490 2730
rect 12510 2710 12515 2730
rect 12485 2680 12515 2710
rect 12485 2660 12490 2680
rect 12510 2660 12515 2680
rect 12485 2630 12515 2660
rect 12485 2610 12490 2630
rect 12510 2610 12515 2630
rect 12485 2580 12515 2610
rect 12485 2560 12490 2580
rect 12510 2560 12515 2580
rect 12485 2530 12515 2560
rect 12485 2510 12490 2530
rect 12510 2510 12515 2530
rect 12485 2500 12515 2510
rect 12545 2880 12615 2890
rect 12850 2885 12890 2895
rect 13000 2915 13040 2925
rect 13000 2895 13010 2915
rect 13030 2895 13040 2915
rect 13000 2885 13040 2895
rect 13058 2915 13092 2925
rect 13058 2895 13066 2915
rect 13084 2895 13092 2915
rect 13058 2885 13092 2895
rect 13110 2915 13150 2925
rect 13110 2895 13120 2915
rect 13140 2895 13150 2915
rect 13110 2885 13150 2895
rect 13220 2915 13260 2925
rect 13220 2895 13230 2915
rect 13250 2895 13260 2915
rect 13220 2885 13260 2895
rect 13330 2915 13370 2925
rect 13330 2895 13340 2915
rect 13360 2895 13370 2915
rect 13330 2885 13370 2895
rect 13440 2915 13480 2925
rect 13440 2895 13450 2915
rect 13470 2895 13480 2915
rect 13440 2885 13480 2895
rect 13550 2915 13590 2925
rect 13550 2895 13560 2915
rect 13580 2895 13590 2915
rect 13550 2885 13590 2895
rect 13660 2915 13700 2925
rect 13660 2895 13670 2915
rect 13690 2895 13700 2915
rect 13660 2885 13700 2895
rect 13770 2915 13810 2925
rect 13770 2895 13780 2915
rect 13800 2895 13810 2915
rect 13770 2885 13810 2895
rect 13880 2915 13920 2925
rect 13880 2895 13890 2915
rect 13910 2895 13920 2915
rect 13880 2885 13920 2895
rect 13990 2915 14030 2925
rect 13990 2895 14000 2915
rect 14020 2895 14030 2915
rect 13990 2885 14030 2895
rect 14140 2915 14180 2925
rect 14140 2895 14150 2915
rect 14170 2895 14180 2915
rect 18680 2920 18690 2940
rect 18710 2920 18720 2940
rect 18680 2910 18720 2920
rect 18840 2940 18880 2950
rect 18840 2920 18850 2940
rect 18870 2920 18880 2940
rect 18840 2910 18880 2920
rect 18960 2940 19000 2950
rect 18960 2920 18970 2940
rect 18990 2920 19000 2940
rect 18960 2910 19000 2920
rect 19080 2940 19120 2950
rect 19080 2920 19090 2940
rect 19110 2920 19120 2940
rect 19080 2910 19120 2920
rect 19200 2940 19240 2950
rect 19200 2920 19210 2940
rect 19230 2920 19240 2940
rect 19200 2910 19240 2920
rect 19320 2940 19360 2950
rect 19320 2920 19330 2940
rect 19350 2920 19360 2940
rect 19320 2910 19360 2920
rect 19440 2940 19480 2950
rect 19440 2920 19450 2940
rect 19470 2920 19480 2940
rect 19440 2910 19480 2920
rect 19560 2940 19600 2950
rect 19560 2920 19570 2940
rect 19590 2920 19600 2940
rect 19560 2910 19600 2920
rect 19680 2940 19720 2950
rect 19680 2920 19690 2940
rect 19710 2920 19720 2940
rect 19680 2910 19720 2920
rect 19800 2940 19840 2950
rect 19800 2920 19810 2940
rect 19830 2920 19840 2940
rect 19800 2910 19840 2920
rect 19920 2940 19960 2950
rect 19920 2920 19930 2940
rect 19950 2920 19960 2940
rect 19920 2910 19960 2920
rect 19980 2910 20020 2950
rect 20080 2940 20120 2950
rect 20355 2945 20425 2955
rect 20450 3225 20480 3235
rect 20450 3205 20455 3225
rect 20475 3205 20480 3225
rect 20450 3175 20480 3205
rect 20450 3155 20455 3175
rect 20475 3155 20480 3175
rect 20450 3125 20480 3155
rect 20450 3105 20455 3125
rect 20475 3105 20480 3125
rect 20450 3075 20480 3105
rect 20450 3055 20455 3075
rect 20475 3055 20480 3075
rect 20450 3025 20480 3055
rect 20450 3005 20455 3025
rect 20475 3005 20480 3025
rect 20450 2975 20480 3005
rect 20450 2955 20455 2975
rect 20475 2955 20480 2975
rect 20450 2945 20480 2955
rect 20505 3225 20535 3235
rect 20505 3205 20510 3225
rect 20530 3205 20535 3225
rect 20505 3175 20535 3205
rect 20505 3155 20510 3175
rect 20530 3155 20535 3175
rect 20505 3125 20535 3155
rect 20505 3105 20510 3125
rect 20530 3105 20535 3125
rect 20505 3075 20535 3105
rect 20505 3055 20510 3075
rect 20530 3055 20535 3075
rect 20505 3025 20535 3055
rect 20505 3005 20510 3025
rect 20530 3005 20535 3025
rect 20505 2975 20535 3005
rect 20505 2955 20510 2975
rect 20530 2955 20535 2975
rect 20505 2945 20535 2955
rect 20560 3225 20590 3235
rect 20560 3205 20565 3225
rect 20585 3205 20590 3225
rect 20560 3175 20590 3205
rect 20560 3155 20565 3175
rect 20585 3155 20590 3175
rect 20560 3125 20590 3155
rect 20560 3105 20565 3125
rect 20585 3105 20590 3125
rect 20560 3075 20590 3105
rect 20560 3055 20565 3075
rect 20585 3055 20590 3075
rect 20560 3025 20590 3055
rect 20560 3005 20565 3025
rect 20585 3005 20590 3025
rect 20560 2975 20590 3005
rect 20560 2955 20565 2975
rect 20585 2955 20590 2975
rect 20560 2945 20590 2955
rect 20615 3225 20645 3235
rect 20615 3205 20620 3225
rect 20640 3205 20645 3225
rect 20615 3175 20645 3205
rect 20615 3155 20620 3175
rect 20640 3155 20645 3175
rect 20615 3125 20645 3155
rect 20615 3105 20620 3125
rect 20640 3105 20645 3125
rect 20615 3075 20645 3105
rect 20615 3055 20620 3075
rect 20640 3055 20645 3075
rect 20615 3025 20645 3055
rect 20615 3005 20620 3025
rect 20640 3005 20645 3025
rect 20615 2975 20645 3005
rect 20615 2955 20620 2975
rect 20640 2955 20645 2975
rect 20615 2945 20645 2955
rect 20670 3225 20700 3235
rect 20670 3205 20675 3225
rect 20695 3205 20700 3225
rect 20670 3175 20700 3205
rect 20670 3155 20675 3175
rect 20695 3155 20700 3175
rect 20670 3125 20700 3155
rect 20670 3105 20675 3125
rect 20695 3105 20700 3125
rect 20670 3075 20700 3105
rect 20670 3055 20675 3075
rect 20695 3055 20700 3075
rect 20670 3025 20700 3055
rect 20670 3005 20675 3025
rect 20695 3005 20700 3025
rect 20670 2975 20700 3005
rect 20670 2955 20675 2975
rect 20695 2955 20700 2975
rect 20670 2945 20700 2955
rect 20725 3225 20755 3235
rect 20725 3205 20730 3225
rect 20750 3205 20755 3225
rect 20725 3175 20755 3205
rect 20725 3155 20730 3175
rect 20750 3155 20755 3175
rect 20725 3125 20755 3155
rect 20725 3105 20730 3125
rect 20750 3105 20755 3125
rect 20725 3075 20755 3105
rect 20725 3055 20730 3075
rect 20750 3055 20755 3075
rect 20725 3025 20755 3055
rect 20725 3005 20730 3025
rect 20750 3005 20755 3025
rect 20725 2975 20755 3005
rect 20725 2955 20730 2975
rect 20750 2955 20755 2975
rect 20725 2945 20755 2955
rect 20780 3225 20810 3235
rect 20780 3205 20785 3225
rect 20805 3205 20810 3225
rect 20780 3175 20810 3205
rect 20780 3155 20785 3175
rect 20805 3155 20810 3175
rect 20780 3125 20810 3155
rect 20780 3105 20785 3125
rect 20805 3105 20810 3125
rect 20780 3075 20810 3105
rect 20780 3055 20785 3075
rect 20805 3055 20810 3075
rect 20780 3025 20810 3055
rect 20780 3005 20785 3025
rect 20805 3005 20810 3025
rect 20780 2975 20810 3005
rect 20780 2955 20785 2975
rect 20805 2955 20810 2975
rect 20780 2945 20810 2955
rect 20835 3225 20865 3235
rect 20835 3205 20840 3225
rect 20860 3205 20865 3225
rect 20835 3175 20865 3205
rect 20835 3155 20840 3175
rect 20860 3155 20865 3175
rect 20835 3125 20865 3155
rect 20835 3105 20840 3125
rect 20860 3105 20865 3125
rect 20835 3075 20865 3105
rect 20835 3055 20840 3075
rect 20860 3055 20865 3075
rect 20835 3025 20865 3055
rect 20835 3005 20840 3025
rect 20860 3005 20865 3025
rect 20835 2975 20865 3005
rect 20835 2955 20840 2975
rect 20860 2955 20865 2975
rect 20835 2945 20865 2955
rect 20890 3225 20920 3235
rect 20890 3205 20895 3225
rect 20915 3205 20920 3225
rect 20890 3175 20920 3205
rect 20890 3155 20895 3175
rect 20915 3155 20920 3175
rect 20890 3125 20920 3155
rect 20890 3105 20895 3125
rect 20915 3105 20920 3125
rect 20890 3075 20920 3105
rect 20890 3055 20895 3075
rect 20915 3055 20920 3075
rect 20890 3025 20920 3055
rect 20890 3005 20895 3025
rect 20915 3005 20920 3025
rect 20890 2975 20920 3005
rect 20890 2955 20895 2975
rect 20915 2955 20920 2975
rect 20890 2945 20920 2955
rect 20945 3225 20975 3235
rect 20945 3205 20950 3225
rect 20970 3205 20975 3225
rect 20945 3175 20975 3205
rect 20945 3155 20950 3175
rect 20970 3155 20975 3175
rect 20945 3125 20975 3155
rect 20945 3105 20950 3125
rect 20970 3105 20975 3125
rect 20945 3075 20975 3105
rect 20945 3055 20950 3075
rect 20970 3055 20975 3075
rect 20945 3025 20975 3055
rect 20945 3005 20950 3025
rect 20970 3005 20975 3025
rect 20945 2975 20975 3005
rect 20945 2955 20950 2975
rect 20970 2955 20975 2975
rect 20945 2945 20975 2955
rect 21000 3225 21030 3235
rect 21000 3205 21005 3225
rect 21025 3205 21030 3225
rect 21000 3175 21030 3205
rect 21000 3155 21005 3175
rect 21025 3155 21030 3175
rect 21000 3125 21030 3155
rect 21000 3105 21005 3125
rect 21025 3105 21030 3125
rect 21000 3075 21030 3105
rect 21000 3055 21005 3075
rect 21025 3055 21030 3075
rect 21000 3025 21030 3055
rect 21000 3005 21005 3025
rect 21025 3005 21030 3025
rect 21000 2975 21030 3005
rect 21000 2955 21005 2975
rect 21025 2955 21030 2975
rect 21000 2945 21030 2955
rect 21055 3225 21085 3235
rect 21055 3205 21060 3225
rect 21080 3205 21085 3225
rect 21055 3175 21085 3205
rect 21055 3155 21060 3175
rect 21080 3155 21085 3175
rect 21055 3125 21085 3155
rect 21055 3105 21060 3125
rect 21080 3105 21085 3125
rect 21055 3075 21085 3105
rect 21055 3055 21060 3075
rect 21080 3055 21085 3075
rect 21055 3025 21085 3055
rect 21055 3005 21060 3025
rect 21080 3005 21085 3025
rect 21055 2975 21085 3005
rect 21055 2955 21060 2975
rect 21080 2955 21085 2975
rect 21055 2945 21085 2955
rect 21110 3225 21140 3235
rect 21110 3205 21115 3225
rect 21135 3205 21140 3225
rect 21110 3175 21140 3205
rect 21110 3155 21115 3175
rect 21135 3155 21140 3175
rect 21110 3125 21140 3155
rect 21110 3105 21115 3125
rect 21135 3105 21140 3125
rect 21110 3075 21140 3105
rect 21110 3055 21115 3075
rect 21135 3055 21140 3075
rect 21110 3025 21140 3055
rect 21110 3005 21115 3025
rect 21135 3005 21140 3025
rect 21110 2975 21140 3005
rect 21110 2955 21115 2975
rect 21135 2955 21140 2975
rect 21110 2945 21140 2955
rect 21165 3225 21195 3235
rect 21165 3205 21170 3225
rect 21190 3205 21195 3225
rect 21165 3175 21195 3205
rect 21165 3155 21170 3175
rect 21190 3155 21195 3175
rect 21165 3125 21195 3155
rect 21165 3105 21170 3125
rect 21190 3105 21195 3125
rect 21165 3075 21195 3105
rect 21165 3055 21170 3075
rect 21190 3055 21195 3075
rect 21165 3025 21195 3055
rect 21165 3005 21170 3025
rect 21190 3005 21195 3025
rect 21165 2975 21195 3005
rect 21165 2955 21170 2975
rect 21190 2955 21195 2975
rect 21165 2945 21195 2955
rect 21220 3225 21250 3235
rect 21220 3205 21225 3225
rect 21245 3205 21250 3225
rect 21220 3175 21250 3205
rect 21220 3155 21225 3175
rect 21245 3155 21250 3175
rect 21220 3125 21250 3155
rect 21220 3105 21225 3125
rect 21245 3105 21250 3125
rect 21220 3075 21250 3105
rect 21220 3055 21225 3075
rect 21245 3055 21250 3075
rect 21220 3025 21250 3055
rect 21220 3005 21225 3025
rect 21245 3005 21250 3025
rect 21220 2975 21250 3005
rect 21220 2955 21225 2975
rect 21245 2955 21250 2975
rect 21220 2945 21250 2955
rect 21275 3225 21305 3235
rect 21275 3205 21280 3225
rect 21300 3205 21305 3225
rect 21275 3175 21305 3205
rect 21275 3155 21280 3175
rect 21300 3155 21305 3175
rect 21275 3125 21305 3155
rect 21275 3105 21280 3125
rect 21300 3105 21305 3125
rect 21275 3075 21305 3105
rect 21275 3055 21280 3075
rect 21300 3055 21305 3075
rect 21275 3025 21305 3055
rect 21275 3005 21280 3025
rect 21300 3005 21305 3025
rect 21275 2975 21305 3005
rect 21275 2955 21280 2975
rect 21300 2955 21305 2975
rect 21275 2945 21305 2955
rect 21330 3225 21360 3235
rect 21330 3205 21335 3225
rect 21355 3205 21360 3225
rect 21330 3175 21360 3205
rect 21330 3155 21335 3175
rect 21355 3155 21360 3175
rect 21330 3125 21360 3155
rect 21330 3105 21335 3125
rect 21355 3105 21360 3125
rect 21330 3075 21360 3105
rect 21330 3055 21335 3075
rect 21355 3055 21360 3075
rect 21330 3025 21360 3055
rect 21330 3005 21335 3025
rect 21355 3005 21360 3025
rect 21330 2975 21360 3005
rect 21330 2955 21335 2975
rect 21355 2955 21360 2975
rect 21330 2945 21360 2955
rect 21385 3225 21415 3235
rect 21385 3205 21390 3225
rect 21410 3205 21415 3225
rect 21385 3175 21415 3205
rect 21385 3155 21390 3175
rect 21410 3155 21415 3175
rect 21385 3125 21415 3155
rect 21385 3105 21390 3125
rect 21410 3105 21415 3125
rect 21385 3075 21415 3105
rect 21385 3055 21390 3075
rect 21410 3055 21415 3075
rect 21385 3025 21415 3055
rect 21385 3005 21390 3025
rect 21410 3005 21415 3025
rect 21385 2975 21415 3005
rect 21385 2955 21390 2975
rect 21410 2955 21415 2975
rect 21385 2945 21415 2955
rect 21440 3225 21470 3235
rect 21440 3205 21445 3225
rect 21465 3205 21470 3225
rect 21440 3175 21470 3205
rect 21440 3155 21445 3175
rect 21465 3155 21470 3175
rect 21440 3125 21470 3155
rect 21440 3105 21445 3125
rect 21465 3105 21470 3125
rect 21440 3075 21470 3105
rect 21440 3055 21445 3075
rect 21465 3055 21470 3075
rect 21440 3025 21470 3055
rect 21440 3005 21445 3025
rect 21465 3005 21470 3025
rect 21440 2975 21470 3005
rect 21440 2955 21445 2975
rect 21465 2955 21470 2975
rect 21440 2945 21470 2955
rect 21495 3225 21525 3235
rect 21495 3205 21500 3225
rect 21520 3205 21525 3225
rect 21495 3175 21525 3205
rect 21495 3155 21500 3175
rect 21520 3155 21525 3175
rect 21495 3125 21525 3155
rect 21495 3105 21500 3125
rect 21520 3105 21525 3125
rect 21495 3075 21525 3105
rect 21495 3055 21500 3075
rect 21520 3055 21525 3075
rect 21495 3025 21525 3055
rect 21495 3005 21500 3025
rect 21520 3005 21525 3025
rect 21495 2975 21525 3005
rect 21495 2955 21500 2975
rect 21520 2955 21525 2975
rect 21495 2945 21525 2955
rect 21550 3225 21580 3235
rect 21550 3205 21555 3225
rect 21575 3205 21580 3225
rect 21550 3175 21580 3205
rect 21550 3155 21555 3175
rect 21575 3155 21580 3175
rect 21550 3125 21580 3155
rect 21550 3105 21555 3125
rect 21575 3105 21580 3125
rect 21550 3075 21580 3105
rect 21550 3055 21555 3075
rect 21575 3055 21580 3075
rect 21550 3025 21580 3055
rect 21550 3005 21555 3025
rect 21575 3005 21580 3025
rect 21550 2975 21580 3005
rect 21550 2955 21555 2975
rect 21575 2955 21580 2975
rect 21550 2945 21580 2955
rect 21605 3225 21675 3235
rect 21605 3205 21610 3225
rect 21630 3205 21650 3225
rect 21670 3205 21675 3225
rect 21605 3175 21675 3205
rect 21605 3155 21610 3175
rect 21630 3155 21650 3175
rect 21670 3155 21675 3175
rect 21605 3125 21675 3155
rect 21605 3105 21610 3125
rect 21630 3105 21650 3125
rect 21670 3105 21675 3125
rect 21605 3075 21675 3105
rect 21605 3055 21610 3075
rect 21630 3055 21650 3075
rect 21670 3055 21675 3075
rect 21605 3025 21675 3055
rect 21605 3005 21610 3025
rect 21630 3005 21650 3025
rect 21670 3005 21675 3025
rect 21605 2975 21675 3005
rect 21605 2955 21610 2975
rect 21630 2955 21650 2975
rect 21670 2955 21675 2975
rect 21605 2945 21675 2955
rect 20080 2920 20090 2940
rect 20110 2920 20120 2940
rect 20360 2925 20380 2945
rect 20510 2925 20530 2945
rect 20620 2925 20640 2945
rect 20730 2925 20750 2945
rect 20840 2925 20860 2945
rect 20950 2925 20970 2945
rect 21060 2925 21080 2945
rect 21170 2925 21190 2945
rect 21280 2925 21300 2945
rect 21390 2925 21410 2945
rect 21500 2925 21520 2945
rect 21650 2925 21670 2945
rect 20080 2910 20120 2920
rect 20350 2915 20390 2925
rect 14140 2885 14180 2895
rect 18690 2890 18710 2910
rect 18850 2890 18870 2910
rect 18970 2890 18990 2910
rect 19090 2890 19110 2910
rect 19210 2890 19230 2910
rect 19330 2890 19350 2910
rect 19450 2890 19470 2910
rect 19570 2890 19590 2910
rect 19690 2890 19710 2910
rect 19810 2890 19830 2910
rect 19930 2890 19950 2910
rect 20090 2890 20110 2910
rect 20350 2895 20360 2915
rect 20380 2895 20390 2915
rect 12545 2860 12550 2880
rect 12570 2860 12590 2880
rect 12610 2860 12615 2880
rect 12545 2830 12615 2860
rect 18685 2880 18755 2890
rect 18685 2860 18690 2880
rect 18710 2860 18730 2880
rect 18750 2860 18755 2880
rect 12545 2810 12550 2830
rect 12570 2810 12590 2830
rect 12610 2810 12615 2830
rect 12545 2780 12615 2810
rect 12545 2760 12550 2780
rect 12570 2760 12590 2780
rect 12610 2760 12615 2780
rect 12545 2730 12615 2760
rect 12545 2710 12550 2730
rect 12570 2710 12590 2730
rect 12610 2710 12615 2730
rect 12545 2680 12615 2710
rect 13055 2695 13095 2836
rect 18685 2830 18755 2860
rect 18685 2810 18690 2830
rect 18710 2810 18730 2830
rect 18750 2810 18755 2830
rect 18685 2780 18755 2810
rect 18685 2760 18690 2780
rect 18710 2760 18730 2780
rect 18750 2760 18755 2780
rect 18685 2730 18755 2760
rect 18685 2710 18690 2730
rect 18710 2710 18730 2730
rect 18750 2710 18755 2730
rect 12545 2660 12550 2680
rect 12570 2660 12590 2680
rect 12610 2660 12615 2680
rect 18685 2680 18755 2710
rect 12545 2630 12615 2660
rect 12945 2665 12985 2675
rect 12945 2645 12955 2665
rect 12975 2645 12985 2665
rect 12945 2635 12985 2645
rect 13055 2665 13095 2675
rect 13055 2645 13065 2665
rect 13085 2645 13095 2665
rect 13055 2635 13095 2645
rect 13165 2665 13205 2675
rect 13165 2645 13175 2665
rect 13195 2645 13205 2665
rect 13165 2635 13205 2645
rect 13275 2665 13315 2675
rect 13275 2645 13285 2665
rect 13305 2645 13315 2665
rect 13275 2635 13315 2645
rect 13385 2665 13425 2675
rect 13385 2645 13395 2665
rect 13415 2645 13425 2665
rect 13385 2635 13425 2645
rect 13495 2665 13535 2675
rect 13495 2645 13505 2665
rect 13525 2645 13535 2665
rect 13495 2635 13535 2645
rect 13605 2665 13645 2675
rect 13605 2645 13615 2665
rect 13635 2645 13645 2665
rect 13605 2635 13645 2645
rect 13715 2665 13755 2675
rect 13715 2645 13725 2665
rect 13745 2645 13755 2665
rect 13715 2635 13755 2645
rect 13825 2665 13865 2675
rect 13825 2645 13835 2665
rect 13855 2645 13865 2665
rect 13825 2635 13865 2645
rect 13935 2665 13975 2675
rect 13935 2645 13945 2665
rect 13965 2645 13975 2665
rect 13935 2635 13975 2645
rect 14045 2665 14085 2675
rect 14045 2645 14055 2665
rect 14075 2645 14085 2665
rect 14045 2635 14085 2645
rect 17235 2665 17275 2675
rect 17235 2645 17245 2665
rect 17265 2645 17275 2665
rect 17235 2635 17275 2645
rect 17345 2665 17385 2675
rect 17345 2645 17355 2665
rect 17375 2645 17385 2665
rect 17345 2635 17385 2645
rect 17455 2665 17495 2675
rect 17455 2645 17465 2665
rect 17485 2645 17495 2665
rect 17455 2635 17495 2645
rect 17565 2665 17605 2675
rect 17565 2645 17575 2665
rect 17595 2645 17605 2665
rect 17565 2635 17605 2645
rect 17675 2665 17715 2675
rect 17675 2645 17685 2665
rect 17705 2645 17715 2665
rect 17675 2635 17715 2645
rect 17785 2665 17825 2675
rect 17785 2645 17795 2665
rect 17815 2645 17825 2665
rect 17785 2635 17825 2645
rect 17895 2665 17935 2675
rect 17895 2645 17905 2665
rect 17925 2645 17935 2665
rect 17895 2635 17935 2645
rect 18005 2665 18045 2675
rect 18005 2645 18015 2665
rect 18035 2645 18045 2665
rect 18005 2635 18045 2645
rect 18115 2665 18155 2675
rect 18115 2645 18125 2665
rect 18145 2645 18155 2665
rect 18115 2635 18155 2645
rect 18225 2665 18265 2675
rect 18225 2645 18235 2665
rect 18255 2645 18265 2665
rect 18225 2635 18265 2645
rect 18335 2665 18375 2675
rect 18335 2645 18345 2665
rect 18365 2645 18375 2665
rect 18335 2635 18375 2645
rect 18685 2660 18690 2680
rect 18710 2660 18730 2680
rect 18750 2660 18755 2680
rect 12545 2610 12550 2630
rect 12570 2610 12590 2630
rect 12610 2610 12615 2630
rect 12955 2615 12975 2635
rect 13065 2615 13085 2635
rect 13175 2615 13195 2635
rect 13285 2615 13305 2635
rect 13395 2615 13415 2635
rect 13505 2615 13525 2635
rect 13615 2615 13635 2635
rect 13725 2615 13745 2635
rect 13835 2615 13855 2635
rect 13945 2615 13965 2635
rect 14055 2615 14075 2635
rect 17245 2615 17265 2635
rect 17355 2615 17375 2635
rect 17465 2615 17485 2635
rect 17575 2615 17595 2635
rect 17685 2615 17705 2635
rect 17795 2615 17815 2635
rect 17905 2615 17925 2635
rect 18015 2615 18035 2635
rect 18125 2615 18145 2635
rect 18235 2615 18255 2635
rect 18345 2615 18365 2635
rect 18685 2630 18755 2660
rect 12545 2580 12615 2610
rect 12545 2560 12550 2580
rect 12570 2560 12590 2580
rect 12610 2560 12615 2580
rect 12545 2530 12615 2560
rect 12545 2510 12550 2530
rect 12570 2510 12590 2530
rect 12610 2510 12615 2530
rect 12855 2605 12925 2615
rect 12855 2585 12860 2605
rect 12880 2585 12900 2605
rect 12920 2585 12925 2605
rect 12855 2555 12925 2585
rect 12855 2535 12860 2555
rect 12880 2535 12900 2555
rect 12920 2535 12925 2555
rect 12855 2525 12925 2535
rect 12950 2605 12980 2615
rect 12950 2585 12955 2605
rect 12975 2585 12980 2605
rect 12950 2555 12980 2585
rect 12950 2535 12955 2555
rect 12975 2535 12980 2555
rect 12950 2525 12980 2535
rect 13005 2605 13035 2615
rect 13005 2585 13010 2605
rect 13030 2585 13035 2605
rect 13005 2555 13035 2585
rect 13005 2535 13010 2555
rect 13030 2535 13035 2555
rect 13005 2525 13035 2535
rect 13060 2605 13090 2615
rect 13060 2585 13065 2605
rect 13085 2585 13090 2605
rect 13060 2555 13090 2585
rect 13060 2535 13065 2555
rect 13085 2535 13090 2555
rect 13060 2525 13090 2535
rect 13115 2605 13145 2615
rect 13115 2585 13120 2605
rect 13140 2585 13145 2605
rect 13115 2555 13145 2585
rect 13115 2535 13120 2555
rect 13140 2535 13145 2555
rect 13115 2525 13145 2535
rect 13170 2605 13200 2615
rect 13170 2585 13175 2605
rect 13195 2585 13200 2605
rect 13170 2555 13200 2585
rect 13170 2535 13175 2555
rect 13195 2535 13200 2555
rect 13170 2525 13200 2535
rect 13225 2605 13255 2615
rect 13225 2585 13230 2605
rect 13250 2585 13255 2605
rect 13225 2555 13255 2585
rect 13225 2535 13230 2555
rect 13250 2535 13255 2555
rect 13225 2525 13255 2535
rect 13280 2605 13310 2615
rect 13280 2585 13285 2605
rect 13305 2585 13310 2605
rect 13280 2555 13310 2585
rect 13280 2535 13285 2555
rect 13305 2535 13310 2555
rect 13280 2525 13310 2535
rect 13335 2605 13365 2615
rect 13335 2585 13340 2605
rect 13360 2585 13365 2605
rect 13335 2555 13365 2585
rect 13335 2535 13340 2555
rect 13360 2535 13365 2555
rect 13335 2525 13365 2535
rect 13390 2605 13420 2615
rect 13390 2585 13395 2605
rect 13415 2585 13420 2605
rect 13390 2555 13420 2585
rect 13390 2535 13395 2555
rect 13415 2535 13420 2555
rect 13390 2525 13420 2535
rect 13445 2605 13475 2615
rect 13445 2585 13450 2605
rect 13470 2585 13475 2605
rect 13445 2555 13475 2585
rect 13445 2535 13450 2555
rect 13470 2535 13475 2555
rect 13445 2525 13475 2535
rect 13500 2605 13530 2615
rect 13500 2585 13505 2605
rect 13525 2585 13530 2605
rect 13500 2555 13530 2585
rect 13500 2535 13505 2555
rect 13525 2535 13530 2555
rect 13500 2525 13530 2535
rect 13555 2605 13585 2615
rect 13555 2585 13560 2605
rect 13580 2585 13585 2605
rect 13555 2555 13585 2585
rect 13555 2535 13560 2555
rect 13580 2535 13585 2555
rect 13555 2525 13585 2535
rect 13610 2605 13640 2615
rect 13610 2585 13615 2605
rect 13635 2585 13640 2605
rect 13610 2555 13640 2585
rect 13610 2535 13615 2555
rect 13635 2535 13640 2555
rect 13610 2525 13640 2535
rect 13665 2605 13695 2615
rect 13665 2585 13670 2605
rect 13690 2585 13695 2605
rect 13665 2555 13695 2585
rect 13665 2535 13670 2555
rect 13690 2535 13695 2555
rect 13665 2525 13695 2535
rect 13720 2605 13750 2615
rect 13720 2585 13725 2605
rect 13745 2585 13750 2605
rect 13720 2555 13750 2585
rect 13720 2535 13725 2555
rect 13745 2535 13750 2555
rect 13720 2525 13750 2535
rect 13775 2605 13805 2615
rect 13775 2585 13780 2605
rect 13800 2585 13805 2605
rect 13775 2555 13805 2585
rect 13775 2535 13780 2555
rect 13800 2535 13805 2555
rect 13775 2525 13805 2535
rect 13830 2605 13860 2615
rect 13830 2585 13835 2605
rect 13855 2585 13860 2605
rect 13830 2555 13860 2585
rect 13830 2535 13835 2555
rect 13855 2535 13860 2555
rect 13830 2525 13860 2535
rect 13885 2605 13915 2615
rect 13885 2585 13890 2605
rect 13910 2585 13915 2605
rect 13885 2555 13915 2585
rect 13885 2535 13890 2555
rect 13910 2535 13915 2555
rect 13885 2525 13915 2535
rect 13940 2605 13970 2615
rect 13940 2585 13945 2605
rect 13965 2585 13970 2605
rect 13940 2555 13970 2585
rect 13940 2535 13945 2555
rect 13965 2535 13970 2555
rect 13940 2525 13970 2535
rect 13995 2605 14025 2615
rect 13995 2585 14000 2605
rect 14020 2585 14025 2605
rect 13995 2555 14025 2585
rect 13995 2535 14000 2555
rect 14020 2535 14025 2555
rect 13995 2525 14025 2535
rect 14050 2605 14080 2615
rect 14050 2585 14055 2605
rect 14075 2585 14080 2605
rect 14050 2555 14080 2585
rect 14050 2535 14055 2555
rect 14075 2535 14080 2555
rect 14050 2525 14080 2535
rect 14105 2605 14175 2615
rect 14105 2585 14110 2605
rect 14130 2585 14150 2605
rect 14170 2585 14175 2605
rect 14105 2555 14175 2585
rect 14105 2535 14110 2555
rect 14130 2535 14150 2555
rect 14170 2535 14175 2555
rect 14105 2525 14175 2535
rect 17145 2605 17215 2615
rect 17145 2585 17150 2605
rect 17170 2585 17190 2605
rect 17210 2585 17215 2605
rect 17145 2555 17215 2585
rect 17145 2535 17150 2555
rect 17170 2535 17190 2555
rect 17210 2535 17215 2555
rect 17145 2525 17215 2535
rect 17240 2605 17270 2615
rect 17240 2585 17245 2605
rect 17265 2585 17270 2605
rect 17240 2555 17270 2585
rect 17240 2535 17245 2555
rect 17265 2535 17270 2555
rect 17240 2525 17270 2535
rect 17295 2605 17325 2615
rect 17295 2585 17300 2605
rect 17320 2585 17325 2605
rect 17295 2555 17325 2585
rect 17295 2535 17300 2555
rect 17320 2535 17325 2555
rect 17295 2525 17325 2535
rect 17350 2605 17380 2615
rect 17350 2585 17355 2605
rect 17375 2585 17380 2605
rect 17350 2555 17380 2585
rect 17350 2535 17355 2555
rect 17375 2535 17380 2555
rect 17350 2525 17380 2535
rect 17405 2605 17435 2615
rect 17405 2585 17410 2605
rect 17430 2585 17435 2605
rect 17405 2555 17435 2585
rect 17405 2535 17410 2555
rect 17430 2535 17435 2555
rect 17405 2525 17435 2535
rect 17460 2605 17490 2615
rect 17460 2585 17465 2605
rect 17485 2585 17490 2605
rect 17460 2555 17490 2585
rect 17460 2535 17465 2555
rect 17485 2535 17490 2555
rect 17460 2525 17490 2535
rect 17515 2605 17545 2615
rect 17515 2585 17520 2605
rect 17540 2585 17545 2605
rect 17515 2555 17545 2585
rect 17515 2535 17520 2555
rect 17540 2535 17545 2555
rect 17515 2525 17545 2535
rect 17570 2605 17600 2615
rect 17570 2585 17575 2605
rect 17595 2585 17600 2605
rect 17570 2555 17600 2585
rect 17570 2535 17575 2555
rect 17595 2535 17600 2555
rect 17570 2525 17600 2535
rect 17625 2605 17655 2615
rect 17625 2585 17630 2605
rect 17650 2585 17655 2605
rect 17625 2555 17655 2585
rect 17625 2535 17630 2555
rect 17650 2535 17655 2555
rect 17625 2525 17655 2535
rect 17680 2605 17710 2615
rect 17680 2585 17685 2605
rect 17705 2585 17710 2605
rect 17680 2555 17710 2585
rect 17680 2535 17685 2555
rect 17705 2535 17710 2555
rect 17680 2525 17710 2535
rect 17735 2605 17765 2615
rect 17735 2585 17740 2605
rect 17760 2585 17765 2605
rect 17735 2555 17765 2585
rect 17735 2535 17740 2555
rect 17760 2535 17765 2555
rect 17735 2525 17765 2535
rect 17790 2605 17820 2615
rect 17790 2585 17795 2605
rect 17815 2585 17820 2605
rect 17790 2555 17820 2585
rect 17790 2535 17795 2555
rect 17815 2535 17820 2555
rect 17790 2525 17820 2535
rect 17845 2605 17875 2615
rect 17845 2585 17850 2605
rect 17870 2585 17875 2605
rect 17845 2555 17875 2585
rect 17845 2535 17850 2555
rect 17870 2535 17875 2555
rect 17845 2525 17875 2535
rect 17900 2605 17930 2615
rect 17900 2585 17905 2605
rect 17925 2585 17930 2605
rect 17900 2555 17930 2585
rect 17900 2535 17905 2555
rect 17925 2535 17930 2555
rect 17900 2525 17930 2535
rect 17955 2605 17985 2615
rect 17955 2585 17960 2605
rect 17980 2585 17985 2605
rect 17955 2555 17985 2585
rect 17955 2535 17960 2555
rect 17980 2535 17985 2555
rect 17955 2525 17985 2535
rect 18010 2605 18040 2615
rect 18010 2585 18015 2605
rect 18035 2585 18040 2605
rect 18010 2555 18040 2585
rect 18010 2535 18015 2555
rect 18035 2535 18040 2555
rect 18010 2525 18040 2535
rect 18065 2605 18095 2615
rect 18065 2585 18070 2605
rect 18090 2585 18095 2605
rect 18065 2555 18095 2585
rect 18065 2535 18070 2555
rect 18090 2535 18095 2555
rect 18065 2525 18095 2535
rect 18120 2605 18150 2615
rect 18120 2585 18125 2605
rect 18145 2585 18150 2605
rect 18120 2555 18150 2585
rect 18120 2535 18125 2555
rect 18145 2535 18150 2555
rect 18120 2525 18150 2535
rect 18175 2605 18205 2615
rect 18175 2585 18180 2605
rect 18200 2585 18205 2605
rect 18175 2555 18205 2585
rect 18175 2535 18180 2555
rect 18200 2535 18205 2555
rect 18175 2525 18205 2535
rect 18230 2605 18260 2615
rect 18230 2585 18235 2605
rect 18255 2585 18260 2605
rect 18230 2555 18260 2585
rect 18230 2535 18235 2555
rect 18255 2535 18260 2555
rect 18230 2525 18260 2535
rect 18285 2605 18315 2615
rect 18285 2585 18290 2605
rect 18310 2585 18315 2605
rect 18285 2555 18315 2585
rect 18285 2535 18290 2555
rect 18310 2535 18315 2555
rect 18285 2525 18315 2535
rect 18340 2605 18370 2615
rect 18340 2585 18345 2605
rect 18365 2585 18370 2605
rect 18340 2555 18370 2585
rect 18340 2535 18345 2555
rect 18365 2535 18370 2555
rect 18340 2525 18370 2535
rect 18395 2605 18465 2615
rect 18395 2585 18400 2605
rect 18420 2585 18440 2605
rect 18460 2585 18465 2605
rect 18395 2555 18465 2585
rect 18395 2535 18400 2555
rect 18420 2535 18440 2555
rect 18460 2535 18465 2555
rect 18395 2525 18465 2535
rect 18685 2610 18690 2630
rect 18710 2610 18730 2630
rect 18750 2610 18755 2630
rect 18685 2580 18755 2610
rect 18685 2560 18690 2580
rect 18710 2560 18730 2580
rect 18750 2560 18755 2580
rect 18685 2530 18755 2560
rect 12545 2500 12615 2510
rect 12860 2505 12880 2525
rect 13010 2505 13030 2525
rect 13120 2505 13140 2525
rect 13230 2505 13250 2525
rect 13340 2505 13360 2525
rect 13450 2505 13470 2525
rect 13560 2505 13580 2525
rect 13670 2505 13690 2525
rect 13780 2505 13800 2525
rect 13890 2505 13910 2525
rect 14000 2505 14020 2525
rect 14150 2505 14170 2525
rect 17150 2505 17170 2525
rect 17300 2505 17320 2525
rect 17410 2505 17430 2525
rect 17520 2505 17540 2525
rect 17630 2505 17650 2525
rect 17740 2505 17760 2525
rect 17850 2505 17870 2525
rect 17960 2505 17980 2525
rect 18070 2505 18090 2525
rect 18180 2505 18200 2525
rect 18290 2505 18310 2525
rect 18440 2505 18460 2525
rect 18685 2510 18690 2530
rect 18710 2510 18730 2530
rect 18750 2510 18755 2530
rect 10930 2475 10940 2495
rect 10960 2475 10970 2495
rect 11290 2480 11310 2500
rect 11410 2480 11430 2500
rect 11530 2480 11550 2500
rect 11650 2480 11670 2500
rect 11770 2480 11790 2500
rect 11890 2480 11910 2500
rect 12010 2480 12030 2500
rect 12130 2480 12150 2500
rect 12250 2480 12270 2500
rect 12370 2480 12390 2500
rect 12490 2480 12510 2500
rect 12850 2495 12890 2505
rect 10930 2465 10970 2475
rect 11280 2470 11320 2480
rect 4800 2435 4870 2465
rect 11280 2450 11290 2470
rect 11310 2450 11320 2470
rect 4800 2415 4805 2435
rect 4825 2415 4845 2435
rect 4865 2415 4870 2435
rect 4800 2405 4870 2415
rect 10813 2435 10847 2445
rect 11280 2440 11320 2450
rect 11400 2470 11440 2480
rect 11400 2450 11410 2470
rect 11430 2450 11440 2470
rect 11400 2440 11440 2450
rect 11520 2470 11560 2480
rect 11520 2450 11530 2470
rect 11550 2450 11560 2470
rect 11520 2440 11560 2450
rect 11640 2470 11680 2480
rect 11640 2450 11650 2470
rect 11670 2450 11680 2470
rect 11640 2440 11680 2450
rect 11760 2470 11800 2480
rect 11760 2450 11770 2470
rect 11790 2450 11800 2470
rect 11760 2440 11800 2450
rect 11823 2470 11857 2480
rect 11823 2450 11831 2470
rect 11849 2450 11857 2470
rect 11823 2440 11857 2450
rect 11880 2470 11920 2480
rect 11880 2450 11890 2470
rect 11910 2450 11920 2470
rect 11880 2440 11920 2450
rect 12000 2470 12040 2480
rect 12000 2450 12010 2470
rect 12030 2450 12040 2470
rect 12000 2440 12040 2450
rect 12120 2470 12160 2480
rect 12120 2450 12130 2470
rect 12150 2450 12160 2470
rect 12120 2440 12160 2450
rect 12240 2470 12280 2480
rect 12240 2450 12250 2470
rect 12270 2450 12280 2470
rect 12240 2440 12280 2450
rect 12360 2470 12400 2480
rect 12360 2450 12370 2470
rect 12390 2450 12400 2470
rect 12360 2440 12400 2450
rect 12480 2470 12520 2480
rect 12480 2450 12490 2470
rect 12510 2450 12520 2470
rect 12850 2475 12860 2495
rect 12880 2475 12890 2495
rect 12850 2465 12890 2475
rect 13000 2495 13040 2505
rect 13000 2475 13010 2495
rect 13030 2475 13040 2495
rect 13000 2465 13040 2475
rect 13110 2495 13150 2505
rect 13110 2475 13120 2495
rect 13140 2475 13150 2495
rect 13110 2465 13150 2475
rect 13220 2495 13260 2505
rect 13220 2475 13230 2495
rect 13250 2475 13260 2495
rect 13220 2465 13260 2475
rect 13330 2495 13370 2505
rect 13330 2475 13340 2495
rect 13360 2475 13370 2495
rect 13330 2465 13370 2475
rect 13440 2495 13480 2505
rect 13440 2475 13450 2495
rect 13470 2475 13480 2495
rect 13440 2465 13480 2475
rect 13550 2495 13590 2505
rect 13550 2475 13560 2495
rect 13580 2475 13590 2495
rect 13550 2465 13590 2475
rect 13660 2495 13700 2505
rect 13660 2475 13670 2495
rect 13690 2475 13700 2495
rect 13660 2465 13700 2475
rect 13770 2495 13810 2505
rect 13770 2475 13780 2495
rect 13800 2475 13810 2495
rect 13770 2465 13810 2475
rect 13880 2495 13920 2505
rect 13880 2475 13890 2495
rect 13910 2475 13920 2495
rect 13880 2465 13920 2475
rect 13990 2495 14030 2505
rect 13990 2475 14000 2495
rect 14020 2475 14030 2495
rect 13990 2465 14030 2475
rect 14140 2495 14180 2505
rect 14140 2475 14150 2495
rect 14170 2475 14180 2495
rect 14140 2465 14180 2475
rect 17140 2495 17180 2505
rect 17140 2475 17150 2495
rect 17170 2475 17180 2495
rect 17140 2465 17180 2475
rect 17290 2495 17330 2505
rect 17290 2475 17300 2495
rect 17320 2475 17330 2495
rect 17290 2465 17330 2475
rect 17400 2495 17440 2505
rect 17400 2475 17410 2495
rect 17430 2475 17440 2495
rect 17400 2465 17440 2475
rect 17510 2495 17550 2505
rect 17510 2475 17520 2495
rect 17540 2475 17550 2495
rect 17510 2465 17550 2475
rect 17620 2495 17660 2505
rect 17620 2475 17630 2495
rect 17650 2475 17660 2495
rect 17620 2465 17660 2475
rect 17730 2495 17770 2505
rect 17730 2475 17740 2495
rect 17760 2475 17770 2495
rect 17730 2465 17770 2475
rect 17840 2495 17880 2505
rect 17840 2475 17850 2495
rect 17870 2475 17880 2495
rect 17840 2465 17880 2475
rect 17950 2495 17990 2505
rect 17950 2475 17960 2495
rect 17980 2475 17990 2495
rect 17950 2465 17990 2475
rect 18060 2495 18100 2505
rect 18060 2475 18070 2495
rect 18090 2475 18100 2495
rect 18060 2465 18100 2475
rect 18170 2495 18210 2505
rect 18170 2475 18180 2495
rect 18200 2475 18210 2495
rect 18170 2465 18210 2475
rect 18280 2495 18320 2505
rect 18280 2475 18290 2495
rect 18310 2475 18320 2495
rect 18280 2465 18320 2475
rect 18430 2495 18470 2505
rect 18685 2500 18755 2510
rect 18785 2880 18815 2890
rect 18785 2860 18790 2880
rect 18810 2860 18815 2880
rect 18785 2830 18815 2860
rect 18785 2810 18790 2830
rect 18810 2810 18815 2830
rect 18785 2780 18815 2810
rect 18785 2760 18790 2780
rect 18810 2760 18815 2780
rect 18785 2730 18815 2760
rect 18785 2710 18790 2730
rect 18810 2710 18815 2730
rect 18785 2680 18815 2710
rect 18785 2660 18790 2680
rect 18810 2660 18815 2680
rect 18785 2630 18815 2660
rect 18785 2610 18790 2630
rect 18810 2610 18815 2630
rect 18785 2580 18815 2610
rect 18785 2560 18790 2580
rect 18810 2560 18815 2580
rect 18785 2530 18815 2560
rect 18785 2510 18790 2530
rect 18810 2510 18815 2530
rect 18785 2500 18815 2510
rect 18845 2880 18875 2890
rect 18845 2860 18850 2880
rect 18870 2860 18875 2880
rect 18845 2830 18875 2860
rect 18845 2810 18850 2830
rect 18870 2810 18875 2830
rect 18845 2780 18875 2810
rect 18845 2760 18850 2780
rect 18870 2760 18875 2780
rect 18845 2730 18875 2760
rect 18845 2710 18850 2730
rect 18870 2710 18875 2730
rect 18845 2680 18875 2710
rect 18845 2660 18850 2680
rect 18870 2660 18875 2680
rect 18845 2630 18875 2660
rect 18845 2610 18850 2630
rect 18870 2610 18875 2630
rect 18845 2580 18875 2610
rect 18845 2560 18850 2580
rect 18870 2560 18875 2580
rect 18845 2530 18875 2560
rect 18845 2510 18850 2530
rect 18870 2510 18875 2530
rect 18845 2500 18875 2510
rect 18905 2880 18935 2890
rect 18905 2860 18910 2880
rect 18930 2860 18935 2880
rect 18905 2830 18935 2860
rect 18905 2810 18910 2830
rect 18930 2810 18935 2830
rect 18905 2780 18935 2810
rect 18905 2760 18910 2780
rect 18930 2760 18935 2780
rect 18905 2730 18935 2760
rect 18905 2710 18910 2730
rect 18930 2710 18935 2730
rect 18905 2680 18935 2710
rect 18905 2660 18910 2680
rect 18930 2660 18935 2680
rect 18905 2630 18935 2660
rect 18905 2610 18910 2630
rect 18930 2610 18935 2630
rect 18905 2580 18935 2610
rect 18905 2560 18910 2580
rect 18930 2560 18935 2580
rect 18905 2530 18935 2560
rect 18905 2510 18910 2530
rect 18930 2510 18935 2530
rect 18905 2500 18935 2510
rect 18965 2880 18995 2890
rect 18965 2860 18970 2880
rect 18990 2860 18995 2880
rect 18965 2830 18995 2860
rect 18965 2810 18970 2830
rect 18990 2810 18995 2830
rect 18965 2780 18995 2810
rect 18965 2760 18970 2780
rect 18990 2760 18995 2780
rect 18965 2730 18995 2760
rect 18965 2710 18970 2730
rect 18990 2710 18995 2730
rect 18965 2680 18995 2710
rect 18965 2660 18970 2680
rect 18990 2660 18995 2680
rect 18965 2630 18995 2660
rect 18965 2610 18970 2630
rect 18990 2610 18995 2630
rect 18965 2580 18995 2610
rect 18965 2560 18970 2580
rect 18990 2560 18995 2580
rect 18965 2530 18995 2560
rect 18965 2510 18970 2530
rect 18990 2510 18995 2530
rect 18965 2500 18995 2510
rect 19025 2880 19055 2890
rect 19025 2860 19030 2880
rect 19050 2860 19055 2880
rect 19025 2830 19055 2860
rect 19025 2810 19030 2830
rect 19050 2810 19055 2830
rect 19025 2780 19055 2810
rect 19025 2760 19030 2780
rect 19050 2760 19055 2780
rect 19025 2730 19055 2760
rect 19025 2710 19030 2730
rect 19050 2710 19055 2730
rect 19025 2680 19055 2710
rect 19025 2660 19030 2680
rect 19050 2660 19055 2680
rect 19025 2630 19055 2660
rect 19025 2610 19030 2630
rect 19050 2610 19055 2630
rect 19025 2580 19055 2610
rect 19025 2560 19030 2580
rect 19050 2560 19055 2580
rect 19025 2530 19055 2560
rect 19025 2510 19030 2530
rect 19050 2510 19055 2530
rect 19025 2500 19055 2510
rect 19085 2880 19115 2890
rect 19085 2860 19090 2880
rect 19110 2860 19115 2880
rect 19085 2830 19115 2860
rect 19085 2810 19090 2830
rect 19110 2810 19115 2830
rect 19085 2780 19115 2810
rect 19085 2760 19090 2780
rect 19110 2760 19115 2780
rect 19085 2730 19115 2760
rect 19085 2710 19090 2730
rect 19110 2710 19115 2730
rect 19085 2680 19115 2710
rect 19085 2660 19090 2680
rect 19110 2660 19115 2680
rect 19085 2630 19115 2660
rect 19085 2610 19090 2630
rect 19110 2610 19115 2630
rect 19085 2580 19115 2610
rect 19085 2560 19090 2580
rect 19110 2560 19115 2580
rect 19085 2530 19115 2560
rect 19085 2510 19090 2530
rect 19110 2510 19115 2530
rect 19085 2500 19115 2510
rect 19145 2880 19175 2890
rect 19145 2860 19150 2880
rect 19170 2860 19175 2880
rect 19145 2830 19175 2860
rect 19145 2810 19150 2830
rect 19170 2810 19175 2830
rect 19145 2780 19175 2810
rect 19145 2760 19150 2780
rect 19170 2760 19175 2780
rect 19145 2730 19175 2760
rect 19145 2710 19150 2730
rect 19170 2710 19175 2730
rect 19145 2680 19175 2710
rect 19145 2660 19150 2680
rect 19170 2660 19175 2680
rect 19145 2630 19175 2660
rect 19145 2610 19150 2630
rect 19170 2610 19175 2630
rect 19145 2580 19175 2610
rect 19145 2560 19150 2580
rect 19170 2560 19175 2580
rect 19145 2530 19175 2560
rect 19145 2510 19150 2530
rect 19170 2510 19175 2530
rect 19145 2500 19175 2510
rect 19205 2880 19235 2890
rect 19205 2860 19210 2880
rect 19230 2860 19235 2880
rect 19205 2830 19235 2860
rect 19205 2810 19210 2830
rect 19230 2810 19235 2830
rect 19205 2780 19235 2810
rect 19205 2760 19210 2780
rect 19230 2760 19235 2780
rect 19205 2730 19235 2760
rect 19205 2710 19210 2730
rect 19230 2710 19235 2730
rect 19205 2680 19235 2710
rect 19205 2660 19210 2680
rect 19230 2660 19235 2680
rect 19205 2630 19235 2660
rect 19205 2610 19210 2630
rect 19230 2610 19235 2630
rect 19205 2580 19235 2610
rect 19205 2560 19210 2580
rect 19230 2560 19235 2580
rect 19205 2530 19235 2560
rect 19205 2510 19210 2530
rect 19230 2510 19235 2530
rect 19205 2500 19235 2510
rect 19265 2880 19295 2890
rect 19265 2860 19270 2880
rect 19290 2860 19295 2880
rect 19265 2830 19295 2860
rect 19265 2810 19270 2830
rect 19290 2810 19295 2830
rect 19265 2780 19295 2810
rect 19265 2760 19270 2780
rect 19290 2760 19295 2780
rect 19265 2730 19295 2760
rect 19265 2710 19270 2730
rect 19290 2710 19295 2730
rect 19265 2680 19295 2710
rect 19265 2660 19270 2680
rect 19290 2660 19295 2680
rect 19265 2630 19295 2660
rect 19265 2610 19270 2630
rect 19290 2610 19295 2630
rect 19265 2580 19295 2610
rect 19265 2560 19270 2580
rect 19290 2560 19295 2580
rect 19265 2530 19295 2560
rect 19265 2510 19270 2530
rect 19290 2510 19295 2530
rect 19265 2500 19295 2510
rect 19325 2880 19355 2890
rect 19325 2860 19330 2880
rect 19350 2860 19355 2880
rect 19325 2830 19355 2860
rect 19325 2810 19330 2830
rect 19350 2810 19355 2830
rect 19325 2780 19355 2810
rect 19325 2760 19330 2780
rect 19350 2760 19355 2780
rect 19325 2730 19355 2760
rect 19325 2710 19330 2730
rect 19350 2710 19355 2730
rect 19325 2680 19355 2710
rect 19325 2660 19330 2680
rect 19350 2660 19355 2680
rect 19325 2630 19355 2660
rect 19325 2610 19330 2630
rect 19350 2610 19355 2630
rect 19325 2580 19355 2610
rect 19325 2560 19330 2580
rect 19350 2560 19355 2580
rect 19325 2530 19355 2560
rect 19325 2510 19330 2530
rect 19350 2510 19355 2530
rect 19325 2500 19355 2510
rect 19385 2880 19415 2890
rect 19385 2860 19390 2880
rect 19410 2860 19415 2880
rect 19385 2830 19415 2860
rect 19385 2810 19390 2830
rect 19410 2810 19415 2830
rect 19385 2780 19415 2810
rect 19385 2760 19390 2780
rect 19410 2760 19415 2780
rect 19385 2730 19415 2760
rect 19385 2710 19390 2730
rect 19410 2710 19415 2730
rect 19385 2680 19415 2710
rect 19385 2660 19390 2680
rect 19410 2660 19415 2680
rect 19385 2630 19415 2660
rect 19385 2610 19390 2630
rect 19410 2610 19415 2630
rect 19385 2580 19415 2610
rect 19385 2560 19390 2580
rect 19410 2560 19415 2580
rect 19385 2530 19415 2560
rect 19385 2510 19390 2530
rect 19410 2510 19415 2530
rect 19385 2500 19415 2510
rect 19445 2880 19475 2890
rect 19445 2860 19450 2880
rect 19470 2860 19475 2880
rect 19445 2830 19475 2860
rect 19445 2810 19450 2830
rect 19470 2810 19475 2830
rect 19445 2780 19475 2810
rect 19445 2760 19450 2780
rect 19470 2760 19475 2780
rect 19445 2730 19475 2760
rect 19445 2710 19450 2730
rect 19470 2710 19475 2730
rect 19445 2680 19475 2710
rect 19445 2660 19450 2680
rect 19470 2660 19475 2680
rect 19445 2630 19475 2660
rect 19445 2610 19450 2630
rect 19470 2610 19475 2630
rect 19445 2580 19475 2610
rect 19445 2560 19450 2580
rect 19470 2560 19475 2580
rect 19445 2530 19475 2560
rect 19445 2510 19450 2530
rect 19470 2510 19475 2530
rect 19445 2500 19475 2510
rect 19505 2880 19535 2890
rect 19505 2860 19510 2880
rect 19530 2860 19535 2880
rect 19505 2830 19535 2860
rect 19505 2810 19510 2830
rect 19530 2810 19535 2830
rect 19505 2780 19535 2810
rect 19505 2760 19510 2780
rect 19530 2760 19535 2780
rect 19505 2730 19535 2760
rect 19505 2710 19510 2730
rect 19530 2710 19535 2730
rect 19505 2680 19535 2710
rect 19505 2660 19510 2680
rect 19530 2660 19535 2680
rect 19505 2630 19535 2660
rect 19505 2610 19510 2630
rect 19530 2610 19535 2630
rect 19505 2580 19535 2610
rect 19505 2560 19510 2580
rect 19530 2560 19535 2580
rect 19505 2530 19535 2560
rect 19505 2510 19510 2530
rect 19530 2510 19535 2530
rect 19505 2500 19535 2510
rect 19565 2880 19595 2890
rect 19565 2860 19570 2880
rect 19590 2860 19595 2880
rect 19565 2830 19595 2860
rect 19565 2810 19570 2830
rect 19590 2810 19595 2830
rect 19565 2780 19595 2810
rect 19565 2760 19570 2780
rect 19590 2760 19595 2780
rect 19565 2730 19595 2760
rect 19565 2710 19570 2730
rect 19590 2710 19595 2730
rect 19565 2680 19595 2710
rect 19565 2660 19570 2680
rect 19590 2660 19595 2680
rect 19565 2630 19595 2660
rect 19565 2610 19570 2630
rect 19590 2610 19595 2630
rect 19565 2580 19595 2610
rect 19565 2560 19570 2580
rect 19590 2560 19595 2580
rect 19565 2530 19595 2560
rect 19565 2510 19570 2530
rect 19590 2510 19595 2530
rect 19565 2500 19595 2510
rect 19625 2880 19655 2890
rect 19625 2860 19630 2880
rect 19650 2860 19655 2880
rect 19625 2830 19655 2860
rect 19625 2810 19630 2830
rect 19650 2810 19655 2830
rect 19625 2780 19655 2810
rect 19625 2760 19630 2780
rect 19650 2760 19655 2780
rect 19625 2730 19655 2760
rect 19625 2710 19630 2730
rect 19650 2710 19655 2730
rect 19625 2680 19655 2710
rect 19625 2660 19630 2680
rect 19650 2660 19655 2680
rect 19625 2630 19655 2660
rect 19625 2610 19630 2630
rect 19650 2610 19655 2630
rect 19625 2580 19655 2610
rect 19625 2560 19630 2580
rect 19650 2560 19655 2580
rect 19625 2530 19655 2560
rect 19625 2510 19630 2530
rect 19650 2510 19655 2530
rect 19625 2500 19655 2510
rect 19685 2880 19715 2890
rect 19685 2860 19690 2880
rect 19710 2860 19715 2880
rect 19685 2830 19715 2860
rect 19685 2810 19690 2830
rect 19710 2810 19715 2830
rect 19685 2780 19715 2810
rect 19685 2760 19690 2780
rect 19710 2760 19715 2780
rect 19685 2730 19715 2760
rect 19685 2710 19690 2730
rect 19710 2710 19715 2730
rect 19685 2680 19715 2710
rect 19685 2660 19690 2680
rect 19710 2660 19715 2680
rect 19685 2630 19715 2660
rect 19685 2610 19690 2630
rect 19710 2610 19715 2630
rect 19685 2580 19715 2610
rect 19685 2560 19690 2580
rect 19710 2560 19715 2580
rect 19685 2530 19715 2560
rect 19685 2510 19690 2530
rect 19710 2510 19715 2530
rect 19685 2500 19715 2510
rect 19745 2880 19775 2890
rect 19745 2860 19750 2880
rect 19770 2860 19775 2880
rect 19745 2830 19775 2860
rect 19745 2810 19750 2830
rect 19770 2810 19775 2830
rect 19745 2780 19775 2810
rect 19745 2760 19750 2780
rect 19770 2760 19775 2780
rect 19745 2730 19775 2760
rect 19745 2710 19750 2730
rect 19770 2710 19775 2730
rect 19745 2680 19775 2710
rect 19745 2660 19750 2680
rect 19770 2660 19775 2680
rect 19745 2630 19775 2660
rect 19745 2610 19750 2630
rect 19770 2610 19775 2630
rect 19745 2580 19775 2610
rect 19745 2560 19750 2580
rect 19770 2560 19775 2580
rect 19745 2530 19775 2560
rect 19745 2510 19750 2530
rect 19770 2510 19775 2530
rect 19745 2500 19775 2510
rect 19805 2880 19835 2890
rect 19805 2860 19810 2880
rect 19830 2860 19835 2880
rect 19805 2830 19835 2860
rect 19805 2810 19810 2830
rect 19830 2810 19835 2830
rect 19805 2780 19835 2810
rect 19805 2760 19810 2780
rect 19830 2760 19835 2780
rect 19805 2730 19835 2760
rect 19805 2710 19810 2730
rect 19830 2710 19835 2730
rect 19805 2680 19835 2710
rect 19805 2660 19810 2680
rect 19830 2660 19835 2680
rect 19805 2630 19835 2660
rect 19805 2610 19810 2630
rect 19830 2610 19835 2630
rect 19805 2580 19835 2610
rect 19805 2560 19810 2580
rect 19830 2560 19835 2580
rect 19805 2530 19835 2560
rect 19805 2510 19810 2530
rect 19830 2510 19835 2530
rect 19805 2500 19835 2510
rect 19865 2880 19895 2890
rect 19865 2860 19870 2880
rect 19890 2860 19895 2880
rect 19865 2830 19895 2860
rect 19865 2810 19870 2830
rect 19890 2810 19895 2830
rect 19865 2780 19895 2810
rect 19865 2760 19870 2780
rect 19890 2760 19895 2780
rect 19865 2730 19895 2760
rect 19865 2710 19870 2730
rect 19890 2710 19895 2730
rect 19865 2680 19895 2710
rect 19865 2660 19870 2680
rect 19890 2660 19895 2680
rect 19865 2630 19895 2660
rect 19865 2610 19870 2630
rect 19890 2610 19895 2630
rect 19865 2580 19895 2610
rect 19865 2560 19870 2580
rect 19890 2560 19895 2580
rect 19865 2530 19895 2560
rect 19865 2510 19870 2530
rect 19890 2510 19895 2530
rect 19865 2500 19895 2510
rect 19925 2880 19955 2890
rect 19925 2860 19930 2880
rect 19950 2860 19955 2880
rect 19925 2830 19955 2860
rect 19925 2810 19930 2830
rect 19950 2810 19955 2830
rect 19925 2780 19955 2810
rect 19925 2760 19930 2780
rect 19950 2760 19955 2780
rect 19925 2730 19955 2760
rect 19925 2710 19930 2730
rect 19950 2710 19955 2730
rect 19925 2680 19955 2710
rect 19925 2660 19930 2680
rect 19950 2660 19955 2680
rect 19925 2630 19955 2660
rect 19925 2610 19930 2630
rect 19950 2610 19955 2630
rect 19925 2580 19955 2610
rect 19925 2560 19930 2580
rect 19950 2560 19955 2580
rect 19925 2530 19955 2560
rect 19925 2510 19930 2530
rect 19950 2510 19955 2530
rect 19925 2500 19955 2510
rect 19985 2880 20015 2890
rect 19985 2860 19990 2880
rect 20010 2860 20015 2880
rect 19985 2830 20015 2860
rect 19985 2810 19990 2830
rect 20010 2810 20015 2830
rect 19985 2780 20015 2810
rect 19985 2760 19990 2780
rect 20010 2760 20015 2780
rect 19985 2730 20015 2760
rect 19985 2710 19990 2730
rect 20010 2710 20015 2730
rect 19985 2680 20015 2710
rect 19985 2660 19990 2680
rect 20010 2660 20015 2680
rect 19985 2630 20015 2660
rect 19985 2610 19990 2630
rect 20010 2610 20015 2630
rect 19985 2580 20015 2610
rect 19985 2560 19990 2580
rect 20010 2560 20015 2580
rect 19985 2530 20015 2560
rect 19985 2510 19990 2530
rect 20010 2510 20015 2530
rect 19985 2500 20015 2510
rect 20045 2880 20115 2890
rect 20350 2885 20390 2895
rect 20500 2915 20540 2925
rect 20500 2895 20510 2915
rect 20530 2895 20540 2915
rect 20500 2885 20540 2895
rect 20558 2915 20592 2925
rect 20558 2895 20566 2915
rect 20584 2895 20592 2915
rect 20558 2885 20592 2895
rect 20610 2915 20650 2925
rect 20610 2895 20620 2915
rect 20640 2895 20650 2915
rect 20610 2885 20650 2895
rect 20720 2915 20760 2925
rect 20720 2895 20730 2915
rect 20750 2895 20760 2915
rect 20720 2885 20760 2895
rect 20830 2915 20870 2925
rect 20830 2895 20840 2915
rect 20860 2895 20870 2915
rect 20830 2885 20870 2895
rect 20940 2915 20980 2925
rect 20940 2895 20950 2915
rect 20970 2895 20980 2915
rect 20940 2885 20980 2895
rect 21050 2915 21090 2925
rect 21050 2895 21060 2915
rect 21080 2895 21090 2915
rect 21050 2885 21090 2895
rect 21160 2915 21200 2925
rect 21160 2895 21170 2915
rect 21190 2895 21200 2915
rect 21160 2885 21200 2895
rect 21270 2915 21310 2925
rect 21270 2895 21280 2915
rect 21300 2895 21310 2915
rect 21270 2885 21310 2895
rect 21380 2915 21420 2925
rect 21380 2895 21390 2915
rect 21410 2895 21420 2915
rect 21380 2885 21420 2895
rect 21490 2915 21530 2925
rect 21490 2895 21500 2915
rect 21520 2895 21530 2915
rect 21490 2885 21530 2895
rect 21640 2915 21680 2925
rect 21640 2895 21650 2915
rect 21670 2895 21680 2915
rect 21640 2885 21680 2895
rect 20045 2860 20050 2880
rect 20070 2860 20090 2880
rect 20110 2860 20115 2880
rect 20045 2830 20115 2860
rect 20045 2810 20050 2830
rect 20070 2810 20090 2830
rect 20110 2810 20115 2830
rect 20045 2780 20115 2810
rect 20045 2760 20050 2780
rect 20070 2760 20090 2780
rect 20110 2760 20115 2780
rect 20045 2730 20115 2760
rect 20045 2710 20050 2730
rect 20070 2710 20090 2730
rect 20110 2710 20115 2730
rect 20045 2680 20115 2710
rect 20555 2695 20595 2836
rect 20045 2660 20050 2680
rect 20070 2660 20090 2680
rect 20110 2660 20115 2680
rect 20045 2630 20115 2660
rect 20445 2665 20485 2675
rect 20445 2645 20455 2665
rect 20475 2645 20485 2665
rect 20445 2635 20485 2645
rect 20555 2665 20595 2675
rect 20555 2645 20565 2665
rect 20585 2645 20595 2665
rect 20555 2635 20595 2645
rect 20665 2665 20705 2675
rect 20665 2645 20675 2665
rect 20695 2645 20705 2665
rect 20665 2635 20705 2645
rect 20775 2665 20815 2675
rect 20775 2645 20785 2665
rect 20805 2645 20815 2665
rect 20775 2635 20815 2645
rect 20885 2665 20925 2675
rect 20885 2645 20895 2665
rect 20915 2645 20925 2665
rect 20885 2635 20925 2645
rect 20995 2665 21035 2675
rect 20995 2645 21005 2665
rect 21025 2645 21035 2665
rect 20995 2635 21035 2645
rect 21105 2665 21145 2675
rect 21105 2645 21115 2665
rect 21135 2645 21145 2665
rect 21105 2635 21145 2645
rect 21215 2665 21255 2675
rect 21215 2645 21225 2665
rect 21245 2645 21255 2665
rect 21215 2635 21255 2645
rect 21325 2665 21365 2675
rect 21325 2645 21335 2665
rect 21355 2645 21365 2665
rect 21325 2635 21365 2645
rect 21435 2665 21475 2675
rect 21435 2645 21445 2665
rect 21465 2645 21475 2665
rect 21435 2635 21475 2645
rect 21545 2665 21585 2675
rect 21545 2645 21555 2665
rect 21575 2645 21585 2665
rect 21545 2635 21585 2645
rect 20045 2610 20050 2630
rect 20070 2610 20090 2630
rect 20110 2610 20115 2630
rect 20455 2615 20475 2635
rect 20565 2615 20585 2635
rect 20675 2615 20695 2635
rect 20785 2615 20805 2635
rect 20895 2615 20915 2635
rect 21005 2615 21025 2635
rect 21115 2615 21135 2635
rect 21225 2615 21245 2635
rect 21335 2615 21355 2635
rect 21445 2615 21465 2635
rect 21555 2615 21575 2635
rect 20045 2580 20115 2610
rect 20045 2560 20050 2580
rect 20070 2560 20090 2580
rect 20110 2560 20115 2580
rect 20045 2530 20115 2560
rect 20045 2510 20050 2530
rect 20070 2510 20090 2530
rect 20110 2510 20115 2530
rect 20355 2605 20425 2615
rect 20355 2585 20360 2605
rect 20380 2585 20400 2605
rect 20420 2585 20425 2605
rect 20355 2555 20425 2585
rect 20355 2535 20360 2555
rect 20380 2535 20400 2555
rect 20420 2535 20425 2555
rect 20355 2525 20425 2535
rect 20450 2605 20480 2615
rect 20450 2585 20455 2605
rect 20475 2585 20480 2605
rect 20450 2555 20480 2585
rect 20450 2535 20455 2555
rect 20475 2535 20480 2555
rect 20450 2525 20480 2535
rect 20505 2605 20535 2615
rect 20505 2585 20510 2605
rect 20530 2585 20535 2605
rect 20505 2555 20535 2585
rect 20505 2535 20510 2555
rect 20530 2535 20535 2555
rect 20505 2525 20535 2535
rect 20560 2605 20590 2615
rect 20560 2585 20565 2605
rect 20585 2585 20590 2605
rect 20560 2555 20590 2585
rect 20560 2535 20565 2555
rect 20585 2535 20590 2555
rect 20560 2525 20590 2535
rect 20615 2605 20645 2615
rect 20615 2585 20620 2605
rect 20640 2585 20645 2605
rect 20615 2555 20645 2585
rect 20615 2535 20620 2555
rect 20640 2535 20645 2555
rect 20615 2525 20645 2535
rect 20670 2605 20700 2615
rect 20670 2585 20675 2605
rect 20695 2585 20700 2605
rect 20670 2555 20700 2585
rect 20670 2535 20675 2555
rect 20695 2535 20700 2555
rect 20670 2525 20700 2535
rect 20725 2605 20755 2615
rect 20725 2585 20730 2605
rect 20750 2585 20755 2605
rect 20725 2555 20755 2585
rect 20725 2535 20730 2555
rect 20750 2535 20755 2555
rect 20725 2525 20755 2535
rect 20780 2605 20810 2615
rect 20780 2585 20785 2605
rect 20805 2585 20810 2605
rect 20780 2555 20810 2585
rect 20780 2535 20785 2555
rect 20805 2535 20810 2555
rect 20780 2525 20810 2535
rect 20835 2605 20865 2615
rect 20835 2585 20840 2605
rect 20860 2585 20865 2605
rect 20835 2555 20865 2585
rect 20835 2535 20840 2555
rect 20860 2535 20865 2555
rect 20835 2525 20865 2535
rect 20890 2605 20920 2615
rect 20890 2585 20895 2605
rect 20915 2585 20920 2605
rect 20890 2555 20920 2585
rect 20890 2535 20895 2555
rect 20915 2535 20920 2555
rect 20890 2525 20920 2535
rect 20945 2605 20975 2615
rect 20945 2585 20950 2605
rect 20970 2585 20975 2605
rect 20945 2555 20975 2585
rect 20945 2535 20950 2555
rect 20970 2535 20975 2555
rect 20945 2525 20975 2535
rect 21000 2605 21030 2615
rect 21000 2585 21005 2605
rect 21025 2585 21030 2605
rect 21000 2555 21030 2585
rect 21000 2535 21005 2555
rect 21025 2535 21030 2555
rect 21000 2525 21030 2535
rect 21055 2605 21085 2615
rect 21055 2585 21060 2605
rect 21080 2585 21085 2605
rect 21055 2555 21085 2585
rect 21055 2535 21060 2555
rect 21080 2535 21085 2555
rect 21055 2525 21085 2535
rect 21110 2605 21140 2615
rect 21110 2585 21115 2605
rect 21135 2585 21140 2605
rect 21110 2555 21140 2585
rect 21110 2535 21115 2555
rect 21135 2535 21140 2555
rect 21110 2525 21140 2535
rect 21165 2605 21195 2615
rect 21165 2585 21170 2605
rect 21190 2585 21195 2605
rect 21165 2555 21195 2585
rect 21165 2535 21170 2555
rect 21190 2535 21195 2555
rect 21165 2525 21195 2535
rect 21220 2605 21250 2615
rect 21220 2585 21225 2605
rect 21245 2585 21250 2605
rect 21220 2555 21250 2585
rect 21220 2535 21225 2555
rect 21245 2535 21250 2555
rect 21220 2525 21250 2535
rect 21275 2605 21305 2615
rect 21275 2585 21280 2605
rect 21300 2585 21305 2605
rect 21275 2555 21305 2585
rect 21275 2535 21280 2555
rect 21300 2535 21305 2555
rect 21275 2525 21305 2535
rect 21330 2605 21360 2615
rect 21330 2585 21335 2605
rect 21355 2585 21360 2605
rect 21330 2555 21360 2585
rect 21330 2535 21335 2555
rect 21355 2535 21360 2555
rect 21330 2525 21360 2535
rect 21385 2605 21415 2615
rect 21385 2585 21390 2605
rect 21410 2585 21415 2605
rect 21385 2555 21415 2585
rect 21385 2535 21390 2555
rect 21410 2535 21415 2555
rect 21385 2525 21415 2535
rect 21440 2605 21470 2615
rect 21440 2585 21445 2605
rect 21465 2585 21470 2605
rect 21440 2555 21470 2585
rect 21440 2535 21445 2555
rect 21465 2535 21470 2555
rect 21440 2525 21470 2535
rect 21495 2605 21525 2615
rect 21495 2585 21500 2605
rect 21520 2585 21525 2605
rect 21495 2555 21525 2585
rect 21495 2535 21500 2555
rect 21520 2535 21525 2555
rect 21495 2525 21525 2535
rect 21550 2605 21580 2615
rect 21550 2585 21555 2605
rect 21575 2585 21580 2605
rect 21550 2555 21580 2585
rect 21550 2535 21555 2555
rect 21575 2535 21580 2555
rect 21550 2525 21580 2535
rect 21605 2605 21675 2615
rect 21605 2585 21610 2605
rect 21630 2585 21650 2605
rect 21670 2585 21675 2605
rect 21605 2555 21675 2585
rect 21605 2535 21610 2555
rect 21630 2535 21650 2555
rect 21670 2535 21675 2555
rect 21605 2525 21675 2535
rect 20045 2500 20115 2510
rect 20360 2505 20380 2525
rect 20510 2505 20530 2525
rect 20620 2505 20640 2525
rect 20730 2505 20750 2525
rect 20840 2505 20860 2525
rect 20950 2505 20970 2525
rect 21060 2505 21080 2525
rect 21170 2505 21190 2525
rect 21280 2505 21300 2525
rect 21390 2505 21410 2525
rect 21500 2505 21520 2525
rect 21650 2505 21670 2525
rect 18430 2475 18440 2495
rect 18460 2475 18470 2495
rect 18790 2480 18810 2500
rect 18910 2480 18930 2500
rect 19030 2480 19050 2500
rect 19150 2480 19170 2500
rect 19270 2480 19290 2500
rect 19390 2480 19410 2500
rect 19510 2480 19530 2500
rect 19630 2480 19650 2500
rect 19750 2480 19770 2500
rect 19870 2480 19890 2500
rect 19990 2480 20010 2500
rect 20350 2495 20390 2505
rect 18430 2465 18470 2475
rect 18780 2470 18820 2480
rect 12480 2440 12520 2450
rect 18780 2450 18790 2470
rect 18810 2450 18820 2470
rect 10813 2415 10821 2435
rect 10839 2415 10847 2435
rect 10813 2405 10847 2415
rect 12973 2435 13007 2445
rect 12973 2415 12981 2435
rect 12999 2415 13007 2435
rect 12973 2405 13007 2415
rect 18313 2435 18347 2445
rect 18780 2440 18820 2450
rect 18900 2470 18940 2480
rect 18900 2450 18910 2470
rect 18930 2450 18940 2470
rect 18900 2440 18940 2450
rect 19020 2470 19060 2480
rect 19020 2450 19030 2470
rect 19050 2450 19060 2470
rect 19020 2440 19060 2450
rect 19140 2470 19180 2480
rect 19140 2450 19150 2470
rect 19170 2450 19180 2470
rect 19140 2440 19180 2450
rect 19260 2470 19300 2480
rect 19260 2450 19270 2470
rect 19290 2450 19300 2470
rect 19260 2440 19300 2450
rect 19323 2470 19357 2480
rect 19323 2450 19331 2470
rect 19349 2450 19357 2470
rect 19323 2440 19357 2450
rect 19380 2470 19420 2480
rect 19380 2450 19390 2470
rect 19410 2450 19420 2470
rect 19380 2440 19420 2450
rect 19500 2470 19540 2480
rect 19500 2450 19510 2470
rect 19530 2450 19540 2470
rect 19500 2440 19540 2450
rect 19620 2470 19660 2480
rect 19620 2450 19630 2470
rect 19650 2450 19660 2470
rect 19620 2440 19660 2450
rect 19740 2470 19780 2480
rect 19740 2450 19750 2470
rect 19770 2450 19780 2470
rect 19740 2440 19780 2450
rect 19860 2470 19900 2480
rect 19860 2450 19870 2470
rect 19890 2450 19900 2470
rect 19860 2440 19900 2450
rect 19980 2470 20020 2480
rect 19980 2450 19990 2470
rect 20010 2450 20020 2470
rect 20350 2475 20360 2495
rect 20380 2475 20390 2495
rect 20350 2465 20390 2475
rect 20500 2495 20540 2505
rect 20500 2475 20510 2495
rect 20530 2475 20540 2495
rect 20500 2465 20540 2475
rect 20610 2495 20650 2505
rect 20610 2475 20620 2495
rect 20640 2475 20650 2495
rect 20610 2465 20650 2475
rect 20720 2495 20760 2505
rect 20720 2475 20730 2495
rect 20750 2475 20760 2495
rect 20720 2465 20760 2475
rect 20830 2495 20870 2505
rect 20830 2475 20840 2495
rect 20860 2475 20870 2495
rect 20830 2465 20870 2475
rect 20940 2495 20980 2505
rect 20940 2475 20950 2495
rect 20970 2475 20980 2495
rect 20940 2465 20980 2475
rect 21050 2495 21090 2505
rect 21050 2475 21060 2495
rect 21080 2475 21090 2495
rect 21050 2465 21090 2475
rect 21160 2495 21200 2505
rect 21160 2475 21170 2495
rect 21190 2475 21200 2495
rect 21160 2465 21200 2475
rect 21270 2495 21310 2505
rect 21270 2475 21280 2495
rect 21300 2475 21310 2495
rect 21270 2465 21310 2475
rect 21380 2495 21420 2505
rect 21380 2475 21390 2495
rect 21410 2475 21420 2495
rect 21380 2465 21420 2475
rect 21490 2495 21530 2505
rect 21490 2475 21500 2495
rect 21520 2475 21530 2495
rect 21490 2465 21530 2475
rect 21640 2495 21680 2505
rect 21640 2475 21650 2495
rect 21670 2475 21680 2495
rect 21640 2465 21680 2475
rect 19980 2440 20020 2450
rect 18313 2415 18321 2435
rect 18339 2415 18347 2435
rect 18313 2405 18347 2415
rect 20473 2435 20507 2445
rect 20473 2415 20481 2435
rect 20499 2415 20507 2435
rect 20473 2405 20507 2415
rect 3275 2385 3295 2405
rect 3455 2385 3475 2405
rect 3265 2375 3305 2385
rect 3265 2355 3275 2375
rect 3295 2355 3305 2375
rect 3265 2345 3305 2355
rect 3355 2370 3395 2380
rect 3355 2350 3365 2370
rect 3385 2350 3395 2370
rect 2625 2315 2655 2345
rect 3355 2340 3395 2350
rect 3445 2375 3485 2385
rect 3445 2355 3455 2375
rect 3475 2355 3485 2375
rect 3445 2345 3485 2355
rect 3635 2340 3655 2405
rect 3815 2385 3835 2405
rect 3995 2385 4015 2405
rect 4175 2385 4195 2405
rect 3805 2375 3845 2385
rect 3805 2355 3815 2375
rect 3835 2355 3845 2375
rect 3805 2345 3845 2355
rect 3885 2375 3925 2385
rect 3885 2355 3895 2375
rect 3915 2355 3925 2375
rect 3885 2345 3925 2355
rect 3985 2375 4025 2385
rect 3985 2355 3995 2375
rect 4015 2355 4025 2375
rect 3985 2345 4025 2355
rect 4165 2375 4205 2385
rect 4165 2355 4175 2375
rect 4195 2355 4205 2375
rect 4165 2345 4205 2355
rect 4355 2340 4375 2405
rect 4535 2385 4555 2405
rect 4715 2385 4735 2405
rect 4525 2375 4565 2385
rect 4525 2355 4535 2375
rect 4555 2355 4565 2375
rect 4525 2345 4565 2355
rect 4705 2375 4745 2385
rect 4705 2355 4715 2375
rect 4735 2355 4745 2375
rect 4705 2345 4745 2355
rect 9800 2375 9845 2380
rect 9800 2350 9810 2375
rect 9835 2350 9845 2375
rect 9800 2345 9845 2350
rect 10635 2375 10680 2380
rect 10635 2350 10645 2375
rect 10670 2350 10680 2375
rect 10635 2345 10680 2350
rect 13140 2375 13185 2380
rect 13140 2350 13150 2375
rect 13175 2350 13185 2375
rect 13140 2345 13185 2350
rect 13975 2375 14020 2380
rect 13975 2350 13985 2375
rect 14010 2350 14020 2375
rect 13975 2345 14020 2350
rect 17300 2375 17345 2380
rect 17300 2350 17310 2375
rect 17335 2350 17345 2375
rect 17300 2345 17345 2350
rect 18135 2375 18180 2380
rect 18135 2350 18145 2375
rect 18170 2350 18180 2375
rect 18135 2345 18180 2350
rect 20640 2375 20685 2380
rect 20640 2350 20650 2375
rect 20675 2350 20685 2375
rect 20640 2345 20685 2350
rect 21475 2375 21520 2380
rect 21475 2350 21485 2375
rect 21510 2350 21520 2375
rect 21475 2345 21520 2350
rect 3625 2330 3665 2340
rect 3625 2310 3635 2330
rect 3655 2310 3665 2330
rect 3625 2300 3665 2310
rect 4345 2330 4385 2340
rect 4345 2310 4355 2330
rect 4375 2310 4385 2330
rect 4345 2300 4385 2310
rect 9800 2315 9845 2320
rect 2740 2260 2770 2290
rect 3445 2285 3485 2295
rect 3445 2265 3455 2285
rect 3475 2265 3485 2285
rect 3445 2255 3485 2265
rect 4525 2285 4565 2295
rect 9800 2290 9810 2315
rect 9835 2290 9845 2315
rect 4525 2265 4535 2285
rect 4555 2265 4565 2285
rect 4525 2255 4565 2265
rect 5275 2260 5305 2290
rect 9800 2285 9845 2290
rect 10635 2315 10680 2320
rect 10635 2290 10645 2315
rect 10670 2290 10680 2315
rect 10635 2285 10680 2290
rect 13140 2315 13185 2320
rect 13140 2290 13150 2315
rect 13175 2290 13185 2315
rect 13140 2285 13185 2290
rect 13975 2315 14020 2320
rect 13975 2290 13985 2315
rect 14010 2290 14020 2315
rect 13975 2285 14020 2290
rect 17300 2315 17345 2320
rect 17300 2290 17310 2315
rect 17335 2290 17345 2315
rect 17300 2285 17345 2290
rect 18135 2315 18180 2320
rect 18135 2290 18145 2315
rect 18170 2290 18180 2315
rect 18135 2285 18180 2290
rect 20640 2315 20685 2320
rect 20640 2290 20650 2315
rect 20675 2290 20685 2315
rect 20640 2285 20685 2290
rect 21475 2315 21520 2320
rect 21475 2290 21485 2315
rect 21510 2290 21520 2315
rect 21475 2285 21520 2290
rect 10813 2275 10847 2285
rect 10813 2255 10821 2275
rect 10839 2255 10847 2275
rect 10813 2245 10847 2255
rect 12973 2275 13007 2285
rect 12973 2255 12981 2275
rect 12999 2255 13007 2275
rect 12973 2245 13007 2255
rect 18313 2275 18347 2285
rect 18313 2255 18321 2275
rect 18339 2255 18347 2275
rect 18313 2245 18347 2255
rect 20473 2275 20507 2285
rect 20473 2255 20481 2275
rect 20499 2255 20507 2275
rect 20473 2245 20507 2255
rect 2430 2215 2460 2245
rect 3810 2215 3840 2245
rect 9640 2215 9680 2225
rect 2335 2170 2365 2200
rect 9640 2195 9650 2215
rect 9670 2195 9680 2215
rect 9640 2185 9680 2195
rect 9790 2215 9830 2225
rect 9790 2195 9800 2215
rect 9820 2195 9830 2215
rect 9790 2185 9830 2195
rect 9900 2215 9940 2225
rect 9900 2195 9910 2215
rect 9930 2195 9940 2215
rect 9900 2185 9940 2195
rect 10010 2215 10050 2225
rect 10010 2195 10020 2215
rect 10040 2195 10050 2215
rect 10010 2185 10050 2195
rect 10120 2215 10160 2225
rect 10120 2195 10130 2215
rect 10150 2195 10160 2215
rect 10120 2185 10160 2195
rect 10230 2215 10270 2225
rect 10230 2195 10240 2215
rect 10260 2195 10270 2215
rect 10230 2185 10270 2195
rect 10340 2215 10380 2225
rect 10340 2195 10350 2215
rect 10370 2195 10380 2215
rect 10340 2185 10380 2195
rect 10450 2215 10490 2225
rect 10450 2195 10460 2215
rect 10480 2195 10490 2215
rect 10450 2185 10490 2195
rect 10560 2215 10600 2225
rect 10560 2195 10570 2215
rect 10590 2195 10600 2215
rect 10560 2185 10600 2195
rect 10670 2215 10710 2225
rect 10670 2195 10680 2215
rect 10700 2195 10710 2215
rect 10670 2185 10710 2195
rect 10780 2215 10820 2225
rect 10780 2195 10790 2215
rect 10810 2195 10820 2215
rect 10780 2185 10820 2195
rect 10930 2215 10970 2225
rect 10930 2195 10940 2215
rect 10960 2195 10970 2215
rect 10930 2185 10970 2195
rect 12850 2215 12890 2225
rect 12850 2195 12860 2215
rect 12880 2195 12890 2215
rect 12850 2185 12890 2195
rect 13000 2215 13040 2225
rect 13000 2195 13010 2215
rect 13030 2195 13040 2215
rect 13000 2185 13040 2195
rect 13110 2215 13150 2225
rect 13110 2195 13120 2215
rect 13140 2195 13150 2215
rect 13110 2185 13150 2195
rect 13220 2215 13260 2225
rect 13220 2195 13230 2215
rect 13250 2195 13260 2215
rect 13220 2185 13260 2195
rect 13330 2215 13370 2225
rect 13330 2195 13340 2215
rect 13360 2195 13370 2215
rect 13330 2185 13370 2195
rect 13440 2215 13480 2225
rect 13440 2195 13450 2215
rect 13470 2195 13480 2215
rect 13440 2185 13480 2195
rect 13550 2215 13590 2225
rect 13550 2195 13560 2215
rect 13580 2195 13590 2215
rect 13550 2185 13590 2195
rect 13660 2215 13700 2225
rect 13660 2195 13670 2215
rect 13690 2195 13700 2215
rect 13660 2185 13700 2195
rect 13770 2215 13810 2225
rect 13770 2195 13780 2215
rect 13800 2195 13810 2215
rect 13770 2185 13810 2195
rect 13880 2215 13920 2225
rect 13880 2195 13890 2215
rect 13910 2195 13920 2215
rect 13880 2185 13920 2195
rect 13990 2215 14030 2225
rect 13990 2195 14000 2215
rect 14020 2195 14030 2215
rect 13990 2185 14030 2195
rect 14140 2215 14180 2225
rect 14140 2195 14150 2215
rect 14170 2195 14180 2215
rect 14140 2185 14180 2195
rect 17140 2215 17180 2225
rect 17140 2195 17150 2215
rect 17170 2195 17180 2215
rect 17140 2185 17180 2195
rect 17290 2215 17330 2225
rect 17290 2195 17300 2215
rect 17320 2195 17330 2215
rect 17290 2185 17330 2195
rect 17400 2215 17440 2225
rect 17400 2195 17410 2215
rect 17430 2195 17440 2215
rect 17400 2185 17440 2195
rect 17510 2215 17550 2225
rect 17510 2195 17520 2215
rect 17540 2195 17550 2215
rect 17510 2185 17550 2195
rect 17620 2215 17660 2225
rect 17620 2195 17630 2215
rect 17650 2195 17660 2215
rect 17620 2185 17660 2195
rect 17730 2215 17770 2225
rect 17730 2195 17740 2215
rect 17760 2195 17770 2215
rect 17730 2185 17770 2195
rect 17840 2215 17880 2225
rect 17840 2195 17850 2215
rect 17870 2195 17880 2215
rect 17840 2185 17880 2195
rect 17950 2215 17990 2225
rect 17950 2195 17960 2215
rect 17980 2195 17990 2215
rect 17950 2185 17990 2195
rect 18060 2215 18100 2225
rect 18060 2195 18070 2215
rect 18090 2195 18100 2215
rect 18060 2185 18100 2195
rect 18170 2215 18210 2225
rect 18170 2195 18180 2215
rect 18200 2195 18210 2215
rect 18170 2185 18210 2195
rect 18280 2215 18320 2225
rect 18280 2195 18290 2215
rect 18310 2195 18320 2215
rect 18280 2185 18320 2195
rect 18430 2215 18470 2225
rect 18430 2195 18440 2215
rect 18460 2195 18470 2215
rect 18430 2185 18470 2195
rect 20350 2215 20390 2225
rect 20350 2195 20360 2215
rect 20380 2195 20390 2215
rect 20350 2185 20390 2195
rect 20500 2215 20540 2225
rect 20500 2195 20510 2215
rect 20530 2195 20540 2215
rect 20500 2185 20540 2195
rect 20610 2215 20650 2225
rect 20610 2195 20620 2215
rect 20640 2195 20650 2215
rect 20610 2185 20650 2195
rect 20720 2215 20760 2225
rect 20720 2195 20730 2215
rect 20750 2195 20760 2215
rect 20720 2185 20760 2195
rect 20830 2215 20870 2225
rect 20830 2195 20840 2215
rect 20860 2195 20870 2215
rect 20830 2185 20870 2195
rect 20940 2215 20980 2225
rect 20940 2195 20950 2215
rect 20970 2195 20980 2215
rect 20940 2185 20980 2195
rect 21050 2215 21090 2225
rect 21050 2195 21060 2215
rect 21080 2195 21090 2215
rect 21050 2185 21090 2195
rect 21160 2215 21200 2225
rect 21160 2195 21170 2215
rect 21190 2195 21200 2215
rect 21160 2185 21200 2195
rect 21270 2215 21310 2225
rect 21270 2195 21280 2215
rect 21300 2195 21310 2215
rect 21270 2185 21310 2195
rect 21380 2215 21420 2225
rect 21380 2195 21390 2215
rect 21410 2195 21420 2215
rect 21380 2185 21420 2195
rect 21490 2215 21530 2225
rect 21490 2195 21500 2215
rect 21520 2195 21530 2215
rect 21490 2185 21530 2195
rect 21640 2215 21680 2225
rect 21640 2195 21650 2215
rect 21670 2195 21680 2215
rect 21640 2185 21680 2195
rect 9650 2165 9670 2185
rect 9800 2165 9820 2185
rect 9910 2165 9930 2185
rect 10020 2165 10040 2185
rect 10130 2165 10150 2185
rect 10240 2165 10260 2185
rect 10350 2165 10370 2185
rect 10460 2165 10480 2185
rect 10570 2165 10590 2185
rect 10680 2165 10700 2185
rect 10790 2165 10810 2185
rect 10940 2165 10960 2185
rect 11330 2175 11370 2185
rect 9645 2155 9715 2165
rect 2385 2120 2415 2150
rect 3630 2120 3660 2150
rect 4090 2115 4120 2145
rect 5320 2115 5350 2145
rect 9645 2135 9650 2155
rect 9670 2135 9690 2155
rect 9710 2135 9715 2155
rect 9645 2105 9715 2135
rect 2745 2090 2785 2100
rect 2745 2070 2755 2090
rect 2775 2070 2785 2090
rect 2745 2060 2785 2070
rect 2865 2090 2905 2100
rect 2865 2070 2875 2090
rect 2895 2070 2905 2090
rect 2865 2060 2905 2070
rect 2985 2090 3025 2100
rect 2985 2070 2995 2090
rect 3015 2070 3025 2090
rect 2985 2060 3025 2070
rect 3105 2090 3145 2100
rect 3105 2070 3115 2090
rect 3135 2070 3145 2090
rect 3105 2060 3145 2070
rect 3225 2090 3265 2100
rect 3225 2070 3235 2090
rect 3255 2070 3265 2090
rect 3225 2060 3265 2070
rect 3345 2090 3385 2100
rect 3345 2070 3355 2090
rect 3375 2070 3385 2090
rect 3345 2060 3385 2070
rect 3465 2090 3505 2100
rect 3465 2070 3475 2090
rect 3495 2070 3505 2090
rect 3465 2060 3505 2070
rect 3585 2090 3625 2100
rect 3585 2070 3595 2090
rect 3615 2070 3625 2090
rect 3585 2060 3625 2070
rect 3705 2090 3745 2100
rect 3705 2070 3715 2090
rect 3735 2070 3745 2090
rect 3705 2060 3745 2070
rect 3825 2090 3865 2100
rect 3825 2070 3835 2090
rect 3855 2070 3865 2090
rect 3825 2060 3865 2070
rect 3985 2090 4025 2100
rect 3985 2070 3995 2090
rect 4015 2070 4025 2090
rect 3985 2060 4025 2070
rect 4145 2090 4185 2100
rect 4145 2070 4155 2090
rect 4175 2070 4185 2090
rect 4145 2060 4185 2070
rect 4265 2090 4305 2100
rect 4265 2070 4275 2090
rect 4295 2070 4305 2090
rect 4265 2060 4305 2070
rect 4385 2090 4425 2100
rect 4385 2070 4395 2090
rect 4415 2070 4425 2090
rect 4385 2060 4425 2070
rect 4505 2090 4545 2100
rect 4505 2070 4515 2090
rect 4535 2070 4545 2090
rect 4505 2060 4545 2070
rect 4625 2090 4665 2100
rect 4625 2070 4635 2090
rect 4655 2070 4665 2090
rect 4625 2060 4665 2070
rect 4745 2090 4785 2100
rect 4745 2070 4755 2090
rect 4775 2070 4785 2090
rect 4745 2060 4785 2070
rect 4865 2090 4905 2100
rect 4865 2070 4875 2090
rect 4895 2070 4905 2090
rect 4865 2060 4905 2070
rect 4985 2090 5025 2100
rect 4985 2070 4995 2090
rect 5015 2070 5025 2090
rect 4985 2060 5025 2070
rect 5105 2090 5145 2100
rect 5105 2070 5115 2090
rect 5135 2070 5145 2090
rect 5105 2060 5145 2070
rect 5225 2090 5265 2100
rect 5225 2070 5235 2090
rect 5255 2070 5265 2090
rect 5225 2060 5265 2070
rect 9645 2085 9650 2105
rect 9670 2085 9690 2105
rect 9710 2085 9715 2105
rect 125 2015 2135 2055
rect 2620 2045 2660 2055
rect 2620 2025 2630 2045
rect 2650 2025 2660 2045
rect 2620 2015 2660 2025
rect -45 1715 130 1725
rect -45 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 130 1715
rect -45 1685 130 1695
rect 650 1375 775 2015
rect 1330 1375 1455 2015
rect 2010 1375 2135 2015
rect 2630 1995 2650 2015
rect 2755 1995 2775 2060
rect 2805 2045 2845 2055
rect 2805 2025 2815 2045
rect 2835 2025 2845 2045
rect 2805 2015 2845 2025
rect 2815 1995 2835 2015
rect 2875 1995 2895 2060
rect 2995 1995 3015 2060
rect 3115 1995 3135 2060
rect 3165 2045 3205 2055
rect 3165 2025 3175 2045
rect 3195 2025 3205 2045
rect 3165 2015 3205 2025
rect 3175 1995 3195 2015
rect 3235 1995 3255 2060
rect 3355 1995 3375 2060
rect 3475 1995 3495 2060
rect 3525 2045 3565 2055
rect 3525 2025 3535 2045
rect 3555 2025 3565 2045
rect 3525 2015 3565 2025
rect 3535 1995 3555 2015
rect 3595 1995 3615 2060
rect 3715 1995 3735 2060
rect 3835 1995 3855 2060
rect 3885 2045 3925 2055
rect 3885 2025 3895 2045
rect 3915 2025 3925 2045
rect 3885 2015 3925 2025
rect 3895 1995 3915 2015
rect 3995 1995 4015 2060
rect 4085 2045 4125 2055
rect 4085 2025 4095 2045
rect 4115 2025 4125 2045
rect 4085 2015 4125 2025
rect 4095 1995 4115 2015
rect 4155 1995 4175 2060
rect 4275 1995 4295 2060
rect 4395 1995 4415 2060
rect 4445 2045 4485 2055
rect 4445 2025 4455 2045
rect 4475 2025 4485 2045
rect 4445 2015 4485 2025
rect 4455 1995 4475 2015
rect 4515 1995 4535 2060
rect 4635 1995 4655 2060
rect 4755 1995 4775 2060
rect 4805 2045 4845 2055
rect 4805 2025 4815 2045
rect 4835 2025 4845 2045
rect 4805 2015 4845 2025
rect 4815 1995 4835 2015
rect 4875 1995 4895 2060
rect 4995 1995 5015 2060
rect 5115 1995 5135 2060
rect 5165 2045 5205 2055
rect 5165 2025 5175 2045
rect 5195 2025 5205 2045
rect 5165 2015 5205 2025
rect 5175 1995 5195 2015
rect 5235 1995 5255 2060
rect 9645 2055 9715 2085
rect 9645 2035 9650 2055
rect 9670 2035 9690 2055
rect 9710 2035 9715 2055
rect 9645 2025 9715 2035
rect 9740 2155 9770 2165
rect 9740 2135 9745 2155
rect 9765 2135 9770 2155
rect 9740 2105 9770 2135
rect 9740 2085 9745 2105
rect 9765 2085 9770 2105
rect 9740 2055 9770 2085
rect 9740 2035 9745 2055
rect 9765 2035 9770 2055
rect 9740 2025 9770 2035
rect 9795 2155 9825 2165
rect 9795 2135 9800 2155
rect 9820 2135 9825 2155
rect 9795 2105 9825 2135
rect 9795 2085 9800 2105
rect 9820 2085 9825 2105
rect 9795 2055 9825 2085
rect 9795 2035 9800 2055
rect 9820 2035 9825 2055
rect 9795 2025 9825 2035
rect 9850 2155 9880 2165
rect 9850 2135 9855 2155
rect 9875 2135 9880 2155
rect 9850 2105 9880 2135
rect 9850 2085 9855 2105
rect 9875 2085 9880 2105
rect 9850 2055 9880 2085
rect 9850 2035 9855 2055
rect 9875 2035 9880 2055
rect 9850 2025 9880 2035
rect 9905 2155 9935 2165
rect 9905 2135 9910 2155
rect 9930 2135 9935 2155
rect 9905 2105 9935 2135
rect 9905 2085 9910 2105
rect 9930 2085 9935 2105
rect 9905 2055 9935 2085
rect 9905 2035 9910 2055
rect 9930 2035 9935 2055
rect 9905 2025 9935 2035
rect 9960 2155 9990 2165
rect 9960 2135 9965 2155
rect 9985 2135 9990 2155
rect 9960 2105 9990 2135
rect 9960 2085 9965 2105
rect 9985 2085 9990 2105
rect 9960 2055 9990 2085
rect 9960 2035 9965 2055
rect 9985 2035 9990 2055
rect 9960 2025 9990 2035
rect 10015 2155 10045 2165
rect 10015 2135 10020 2155
rect 10040 2135 10045 2155
rect 10015 2105 10045 2135
rect 10015 2085 10020 2105
rect 10040 2085 10045 2105
rect 10015 2055 10045 2085
rect 10015 2035 10020 2055
rect 10040 2035 10045 2055
rect 10015 2025 10045 2035
rect 10070 2155 10100 2165
rect 10070 2135 10075 2155
rect 10095 2135 10100 2155
rect 10070 2105 10100 2135
rect 10070 2085 10075 2105
rect 10095 2085 10100 2105
rect 10070 2055 10100 2085
rect 10070 2035 10075 2055
rect 10095 2035 10100 2055
rect 10070 2025 10100 2035
rect 10125 2155 10155 2165
rect 10125 2135 10130 2155
rect 10150 2135 10155 2155
rect 10125 2105 10155 2135
rect 10125 2085 10130 2105
rect 10150 2085 10155 2105
rect 10125 2055 10155 2085
rect 10125 2035 10130 2055
rect 10150 2035 10155 2055
rect 10125 2025 10155 2035
rect 10180 2155 10210 2165
rect 10180 2135 10185 2155
rect 10205 2135 10210 2155
rect 10180 2105 10210 2135
rect 10180 2085 10185 2105
rect 10205 2085 10210 2105
rect 10180 2055 10210 2085
rect 10180 2035 10185 2055
rect 10205 2035 10210 2055
rect 10180 2025 10210 2035
rect 10235 2155 10265 2165
rect 10235 2135 10240 2155
rect 10260 2135 10265 2155
rect 10235 2105 10265 2135
rect 10235 2085 10240 2105
rect 10260 2085 10265 2105
rect 10235 2055 10265 2085
rect 10235 2035 10240 2055
rect 10260 2035 10265 2055
rect 10235 2025 10265 2035
rect 10290 2155 10320 2165
rect 10290 2135 10295 2155
rect 10315 2135 10320 2155
rect 10290 2105 10320 2135
rect 10290 2085 10295 2105
rect 10315 2085 10320 2105
rect 10290 2055 10320 2085
rect 10290 2035 10295 2055
rect 10315 2035 10320 2055
rect 10290 2025 10320 2035
rect 10345 2155 10375 2165
rect 10345 2135 10350 2155
rect 10370 2135 10375 2155
rect 10345 2105 10375 2135
rect 10345 2085 10350 2105
rect 10370 2085 10375 2105
rect 10345 2055 10375 2085
rect 10345 2035 10350 2055
rect 10370 2035 10375 2055
rect 10345 2025 10375 2035
rect 10400 2155 10430 2165
rect 10400 2135 10405 2155
rect 10425 2135 10430 2155
rect 10400 2105 10430 2135
rect 10400 2085 10405 2105
rect 10425 2085 10430 2105
rect 10400 2055 10430 2085
rect 10400 2035 10405 2055
rect 10425 2035 10430 2055
rect 10400 2025 10430 2035
rect 10455 2155 10485 2165
rect 10455 2135 10460 2155
rect 10480 2135 10485 2155
rect 10455 2105 10485 2135
rect 10455 2085 10460 2105
rect 10480 2085 10485 2105
rect 10455 2055 10485 2085
rect 10455 2035 10460 2055
rect 10480 2035 10485 2055
rect 10455 2025 10485 2035
rect 10510 2155 10540 2165
rect 10510 2135 10515 2155
rect 10535 2135 10540 2155
rect 10510 2105 10540 2135
rect 10510 2085 10515 2105
rect 10535 2085 10540 2105
rect 10510 2055 10540 2085
rect 10510 2035 10515 2055
rect 10535 2035 10540 2055
rect 10510 2025 10540 2035
rect 10565 2155 10595 2165
rect 10565 2135 10570 2155
rect 10590 2135 10595 2155
rect 10565 2105 10595 2135
rect 10565 2085 10570 2105
rect 10590 2085 10595 2105
rect 10565 2055 10595 2085
rect 10565 2035 10570 2055
rect 10590 2035 10595 2055
rect 10565 2025 10595 2035
rect 10620 2155 10650 2165
rect 10620 2135 10625 2155
rect 10645 2135 10650 2155
rect 10620 2105 10650 2135
rect 10620 2085 10625 2105
rect 10645 2085 10650 2105
rect 10620 2055 10650 2085
rect 10620 2035 10625 2055
rect 10645 2035 10650 2055
rect 10620 2025 10650 2035
rect 10675 2155 10705 2165
rect 10675 2135 10680 2155
rect 10700 2135 10705 2155
rect 10675 2105 10705 2135
rect 10675 2085 10680 2105
rect 10700 2085 10705 2105
rect 10675 2055 10705 2085
rect 10675 2035 10680 2055
rect 10700 2035 10705 2055
rect 10675 2025 10705 2035
rect 10730 2155 10760 2165
rect 10730 2135 10735 2155
rect 10755 2135 10760 2155
rect 10730 2105 10760 2135
rect 10730 2085 10735 2105
rect 10755 2085 10760 2105
rect 10730 2055 10760 2085
rect 10730 2035 10735 2055
rect 10755 2035 10760 2055
rect 10730 2025 10760 2035
rect 10785 2155 10815 2165
rect 10785 2135 10790 2155
rect 10810 2135 10815 2155
rect 10785 2105 10815 2135
rect 10785 2085 10790 2105
rect 10810 2085 10815 2105
rect 10785 2055 10815 2085
rect 10785 2035 10790 2055
rect 10810 2035 10815 2055
rect 10785 2025 10815 2035
rect 10840 2155 10870 2165
rect 10840 2135 10845 2155
rect 10865 2135 10870 2155
rect 10840 2105 10870 2135
rect 10840 2085 10845 2105
rect 10865 2085 10870 2105
rect 10840 2055 10870 2085
rect 10840 2035 10845 2055
rect 10865 2035 10870 2055
rect 10840 2025 10870 2035
rect 10895 2155 10965 2165
rect 10895 2135 10900 2155
rect 10920 2135 10940 2155
rect 10960 2135 10965 2155
rect 11330 2155 11340 2175
rect 11360 2155 11370 2175
rect 11330 2145 11370 2155
rect 11440 2175 11480 2185
rect 11440 2155 11450 2175
rect 11470 2155 11480 2175
rect 11440 2145 11480 2155
rect 11550 2175 11590 2185
rect 11550 2155 11560 2175
rect 11580 2155 11590 2175
rect 11550 2145 11590 2155
rect 11660 2175 11700 2185
rect 11660 2155 11670 2175
rect 11690 2155 11700 2175
rect 11660 2145 11700 2155
rect 11770 2175 11810 2185
rect 11770 2155 11780 2175
rect 11800 2155 11810 2175
rect 11770 2145 11810 2155
rect 11880 2175 11920 2185
rect 11880 2155 11890 2175
rect 11910 2155 11920 2175
rect 11880 2145 11920 2155
rect 11990 2175 12030 2185
rect 11990 2155 12000 2175
rect 12020 2155 12030 2175
rect 11990 2145 12030 2155
rect 12100 2175 12140 2185
rect 12100 2155 12110 2175
rect 12130 2155 12140 2175
rect 12100 2145 12140 2155
rect 12210 2175 12250 2185
rect 12210 2155 12220 2175
rect 12240 2155 12250 2175
rect 12210 2145 12250 2155
rect 12320 2175 12360 2185
rect 12320 2155 12330 2175
rect 12350 2155 12360 2175
rect 12320 2145 12360 2155
rect 12430 2175 12470 2185
rect 12430 2155 12440 2175
rect 12460 2155 12470 2175
rect 12860 2165 12880 2185
rect 13010 2165 13030 2185
rect 13120 2165 13140 2185
rect 13230 2165 13250 2185
rect 13340 2165 13360 2185
rect 13450 2165 13470 2185
rect 13560 2165 13580 2185
rect 13670 2165 13690 2185
rect 13780 2165 13800 2185
rect 13890 2165 13910 2185
rect 14000 2165 14020 2185
rect 14150 2165 14170 2185
rect 17150 2165 17170 2185
rect 17300 2165 17320 2185
rect 17410 2165 17430 2185
rect 17520 2165 17540 2185
rect 17630 2165 17650 2185
rect 17740 2165 17760 2185
rect 17850 2165 17870 2185
rect 17960 2165 17980 2185
rect 18070 2165 18090 2185
rect 18180 2165 18200 2185
rect 18290 2165 18310 2185
rect 18440 2165 18460 2185
rect 18830 2175 18870 2185
rect 12430 2145 12470 2155
rect 12855 2155 12925 2165
rect 10895 2105 10965 2135
rect 11340 2125 11360 2145
rect 11450 2125 11470 2145
rect 11560 2125 11580 2145
rect 11670 2125 11690 2145
rect 11780 2125 11800 2145
rect 11890 2125 11910 2145
rect 12000 2125 12020 2145
rect 12110 2125 12130 2145
rect 12220 2125 12240 2145
rect 12330 2125 12350 2145
rect 12440 2125 12460 2145
rect 12855 2135 12860 2155
rect 12880 2135 12900 2155
rect 12920 2135 12925 2155
rect 10895 2085 10900 2105
rect 10920 2085 10940 2105
rect 10960 2085 10965 2105
rect 10895 2055 10965 2085
rect 10895 2035 10900 2055
rect 10920 2035 10940 2055
rect 10960 2035 10965 2055
rect 10895 2025 10965 2035
rect 11240 2115 11310 2125
rect 11240 2095 11245 2115
rect 11265 2095 11285 2115
rect 11305 2095 11310 2115
rect 11240 2065 11310 2095
rect 11240 2045 11245 2065
rect 11265 2045 11285 2065
rect 11305 2045 11310 2065
rect 9745 2005 9765 2025
rect 9855 2005 9875 2025
rect 9965 2005 9985 2025
rect 10075 2005 10095 2025
rect 10185 2005 10205 2025
rect 10295 2005 10315 2025
rect 10405 2005 10425 2025
rect 10515 2005 10535 2025
rect 10625 2005 10645 2025
rect 10735 2005 10755 2025
rect 10845 2005 10865 2025
rect 11240 2015 11310 2045
rect 9735 1995 9775 2005
rect 2570 1985 2600 1995
rect 2570 1965 2575 1985
rect 2595 1965 2600 1985
rect 2570 1935 2600 1965
rect 2570 1915 2575 1935
rect 2595 1915 2600 1935
rect 2570 1905 2600 1915
rect 2625 1985 2655 1995
rect 2625 1965 2630 1985
rect 2650 1965 2655 1985
rect 2625 1935 2655 1965
rect 2625 1915 2630 1935
rect 2650 1915 2655 1935
rect 2625 1905 2655 1915
rect 2680 1985 2710 1995
rect 2680 1965 2685 1985
rect 2705 1965 2710 1985
rect 2680 1935 2710 1965
rect 2680 1915 2685 1935
rect 2705 1915 2710 1935
rect 2680 1905 2710 1915
rect 2750 1985 2780 1995
rect 2750 1965 2755 1985
rect 2775 1965 2780 1985
rect 2750 1935 2780 1965
rect 2750 1915 2755 1935
rect 2775 1915 2780 1935
rect 2750 1905 2780 1915
rect 2810 1985 2840 1995
rect 2810 1965 2815 1985
rect 2835 1965 2840 1985
rect 2810 1935 2840 1965
rect 2810 1915 2815 1935
rect 2835 1915 2840 1935
rect 2810 1905 2840 1915
rect 2870 1985 2900 1995
rect 2870 1965 2875 1985
rect 2895 1965 2900 1985
rect 2870 1935 2900 1965
rect 2870 1915 2875 1935
rect 2895 1915 2900 1935
rect 2870 1905 2900 1915
rect 2930 1985 2960 1995
rect 2930 1965 2935 1985
rect 2955 1965 2960 1985
rect 2930 1935 2960 1965
rect 2930 1915 2935 1935
rect 2955 1915 2960 1935
rect 2930 1905 2960 1915
rect 2990 1985 3020 1995
rect 2990 1965 2995 1985
rect 3015 1965 3020 1985
rect 2990 1935 3020 1965
rect 2990 1915 2995 1935
rect 3015 1915 3020 1935
rect 2990 1905 3020 1915
rect 3050 1985 3080 1995
rect 3050 1965 3055 1985
rect 3075 1965 3080 1985
rect 3050 1935 3080 1965
rect 3050 1915 3055 1935
rect 3075 1915 3080 1935
rect 3050 1905 3080 1915
rect 3110 1985 3140 1995
rect 3110 1965 3115 1985
rect 3135 1965 3140 1985
rect 3110 1935 3140 1965
rect 3110 1915 3115 1935
rect 3135 1915 3140 1935
rect 3110 1905 3140 1915
rect 3170 1985 3200 1995
rect 3170 1965 3175 1985
rect 3195 1965 3200 1985
rect 3170 1935 3200 1965
rect 3170 1915 3175 1935
rect 3195 1915 3200 1935
rect 3170 1905 3200 1915
rect 3230 1985 3260 1995
rect 3230 1965 3235 1985
rect 3255 1965 3260 1985
rect 3230 1935 3260 1965
rect 3230 1915 3235 1935
rect 3255 1915 3260 1935
rect 3230 1905 3260 1915
rect 3290 1985 3320 1995
rect 3290 1965 3295 1985
rect 3315 1965 3320 1985
rect 3290 1935 3320 1965
rect 3290 1915 3295 1935
rect 3315 1915 3320 1935
rect 3290 1905 3320 1915
rect 3350 1985 3380 1995
rect 3350 1965 3355 1985
rect 3375 1965 3380 1985
rect 3350 1935 3380 1965
rect 3350 1915 3355 1935
rect 3375 1915 3380 1935
rect 3350 1905 3380 1915
rect 3410 1985 3440 1995
rect 3410 1965 3415 1985
rect 3435 1965 3440 1985
rect 3410 1935 3440 1965
rect 3410 1915 3415 1935
rect 3435 1915 3440 1935
rect 3410 1905 3440 1915
rect 3470 1985 3500 1995
rect 3470 1965 3475 1985
rect 3495 1965 3500 1985
rect 3470 1935 3500 1965
rect 3470 1915 3475 1935
rect 3495 1915 3500 1935
rect 3470 1905 3500 1915
rect 3530 1985 3560 1995
rect 3530 1965 3535 1985
rect 3555 1965 3560 1985
rect 3530 1935 3560 1965
rect 3530 1915 3535 1935
rect 3555 1915 3560 1935
rect 3530 1905 3560 1915
rect 3590 1985 3620 1995
rect 3590 1965 3595 1985
rect 3615 1965 3620 1985
rect 3590 1935 3620 1965
rect 3590 1915 3595 1935
rect 3615 1915 3620 1935
rect 3590 1905 3620 1915
rect 3650 1985 3680 1995
rect 3650 1965 3655 1985
rect 3675 1965 3680 1985
rect 3650 1935 3680 1965
rect 3650 1915 3655 1935
rect 3675 1915 3680 1935
rect 3650 1905 3680 1915
rect 3710 1985 3740 1995
rect 3710 1965 3715 1985
rect 3735 1965 3740 1985
rect 3710 1935 3740 1965
rect 3710 1915 3715 1935
rect 3735 1915 3740 1935
rect 3710 1905 3740 1915
rect 3770 1985 3800 1995
rect 3770 1965 3775 1985
rect 3795 1965 3800 1985
rect 3770 1935 3800 1965
rect 3770 1915 3775 1935
rect 3795 1915 3800 1935
rect 3770 1905 3800 1915
rect 3830 1985 3860 1995
rect 3830 1965 3835 1985
rect 3855 1965 3860 1985
rect 3830 1935 3860 1965
rect 3830 1915 3835 1935
rect 3855 1915 3860 1935
rect 3830 1905 3860 1915
rect 3890 1985 3920 1995
rect 3890 1965 3895 1985
rect 3915 1965 3920 1985
rect 3890 1935 3920 1965
rect 3890 1915 3895 1935
rect 3915 1915 3920 1935
rect 3890 1905 3920 1915
rect 3950 1985 4060 1995
rect 3950 1965 3955 1985
rect 3975 1965 3995 1985
rect 4015 1965 4035 1985
rect 4055 1965 4060 1985
rect 3950 1935 4060 1965
rect 3950 1915 3955 1935
rect 3975 1915 3995 1935
rect 4015 1915 4035 1935
rect 4055 1915 4060 1935
rect 3950 1905 4060 1915
rect 4090 1985 4120 1995
rect 4090 1965 4095 1985
rect 4115 1965 4120 1985
rect 4090 1935 4120 1965
rect 4090 1915 4095 1935
rect 4115 1915 4120 1935
rect 4090 1905 4120 1915
rect 4150 1985 4180 1995
rect 4150 1965 4155 1985
rect 4175 1965 4180 1985
rect 4150 1935 4180 1965
rect 4150 1915 4155 1935
rect 4175 1915 4180 1935
rect 4150 1905 4180 1915
rect 4210 1985 4240 1995
rect 4210 1965 4215 1985
rect 4235 1965 4240 1985
rect 4210 1935 4240 1965
rect 4210 1915 4215 1935
rect 4235 1915 4240 1935
rect 4210 1905 4240 1915
rect 4270 1985 4300 1995
rect 4270 1965 4275 1985
rect 4295 1965 4300 1985
rect 4270 1935 4300 1965
rect 4270 1915 4275 1935
rect 4295 1915 4300 1935
rect 4270 1905 4300 1915
rect 4330 1985 4360 1995
rect 4330 1965 4335 1985
rect 4355 1965 4360 1985
rect 4330 1935 4360 1965
rect 4330 1915 4335 1935
rect 4355 1915 4360 1935
rect 4330 1905 4360 1915
rect 4390 1985 4420 1995
rect 4390 1965 4395 1985
rect 4415 1965 4420 1985
rect 4390 1935 4420 1965
rect 4390 1915 4395 1935
rect 4415 1915 4420 1935
rect 4390 1905 4420 1915
rect 4450 1985 4480 1995
rect 4450 1965 4455 1985
rect 4475 1965 4480 1985
rect 4450 1935 4480 1965
rect 4450 1915 4455 1935
rect 4475 1915 4480 1935
rect 4450 1905 4480 1915
rect 4510 1985 4540 1995
rect 4510 1965 4515 1985
rect 4535 1965 4540 1985
rect 4510 1935 4540 1965
rect 4510 1915 4515 1935
rect 4535 1915 4540 1935
rect 4510 1905 4540 1915
rect 4570 1985 4600 1995
rect 4570 1965 4575 1985
rect 4595 1965 4600 1985
rect 4570 1935 4600 1965
rect 4570 1915 4575 1935
rect 4595 1915 4600 1935
rect 4570 1905 4600 1915
rect 4630 1985 4660 1995
rect 4630 1965 4635 1985
rect 4655 1965 4660 1985
rect 4630 1935 4660 1965
rect 4630 1915 4635 1935
rect 4655 1915 4660 1935
rect 4630 1905 4660 1915
rect 4690 1985 4720 1995
rect 4690 1965 4695 1985
rect 4715 1965 4720 1985
rect 4690 1935 4720 1965
rect 4690 1915 4695 1935
rect 4715 1915 4720 1935
rect 4690 1905 4720 1915
rect 4750 1985 4780 1995
rect 4750 1965 4755 1985
rect 4775 1965 4780 1985
rect 4750 1935 4780 1965
rect 4750 1915 4755 1935
rect 4775 1915 4780 1935
rect 4750 1905 4780 1915
rect 4810 1985 4840 1995
rect 4810 1965 4815 1985
rect 4835 1965 4840 1985
rect 4810 1935 4840 1965
rect 4810 1915 4815 1935
rect 4835 1915 4840 1935
rect 4810 1905 4840 1915
rect 4870 1985 4900 1995
rect 4870 1965 4875 1985
rect 4895 1965 4900 1985
rect 4870 1935 4900 1965
rect 4870 1915 4875 1935
rect 4895 1915 4900 1935
rect 4870 1905 4900 1915
rect 4930 1985 4960 1995
rect 4930 1965 4935 1985
rect 4955 1965 4960 1985
rect 4930 1935 4960 1965
rect 4930 1915 4935 1935
rect 4955 1915 4960 1935
rect 4930 1905 4960 1915
rect 4990 1985 5020 1995
rect 4990 1965 4995 1985
rect 5015 1965 5020 1985
rect 4990 1935 5020 1965
rect 4990 1915 4995 1935
rect 5015 1915 5020 1935
rect 4990 1905 5020 1915
rect 5050 1985 5080 1995
rect 5050 1965 5055 1985
rect 5075 1965 5080 1985
rect 5050 1935 5080 1965
rect 5050 1915 5055 1935
rect 5075 1915 5080 1935
rect 5050 1905 5080 1915
rect 5110 1985 5140 1995
rect 5110 1965 5115 1985
rect 5135 1965 5140 1985
rect 5110 1935 5140 1965
rect 5110 1915 5115 1935
rect 5135 1915 5140 1935
rect 5110 1905 5140 1915
rect 5170 1985 5200 1995
rect 5170 1965 5175 1985
rect 5195 1965 5200 1985
rect 5170 1935 5200 1965
rect 5170 1915 5175 1935
rect 5195 1915 5200 1935
rect 5170 1905 5200 1915
rect 5230 1985 5260 1995
rect 5230 1965 5235 1985
rect 5255 1965 5260 1985
rect 9735 1975 9745 1995
rect 9763 1975 9775 1995
rect 9735 1965 9775 1975
rect 9845 1995 9885 2005
rect 9845 1975 9855 1995
rect 9873 1975 9885 1995
rect 9845 1965 9885 1975
rect 9955 1995 9995 2005
rect 9955 1975 9965 1995
rect 9983 1975 9995 1995
rect 9955 1965 9995 1975
rect 10065 1995 10105 2005
rect 10065 1975 10075 1995
rect 10093 1975 10105 1995
rect 10065 1965 10105 1975
rect 10175 1995 10215 2005
rect 10175 1975 10185 1995
rect 10203 1975 10215 1995
rect 10175 1965 10215 1975
rect 10285 1995 10325 2005
rect 10285 1975 10295 1995
rect 10313 1975 10325 1995
rect 10285 1965 10325 1975
rect 10395 1995 10435 2005
rect 10395 1975 10405 1995
rect 10423 1975 10435 1995
rect 10395 1965 10435 1975
rect 10505 1995 10545 2005
rect 10505 1975 10515 1995
rect 10533 1975 10545 1995
rect 10505 1965 10545 1975
rect 10615 1995 10655 2005
rect 10615 1975 10625 1995
rect 10643 1975 10655 1995
rect 10615 1965 10655 1975
rect 10725 1995 10765 2005
rect 10725 1975 10735 1995
rect 10753 1975 10765 1995
rect 10725 1965 10765 1975
rect 10835 1995 10875 2005
rect 10835 1975 10845 1995
rect 10863 1975 10875 1995
rect 11240 1995 11245 2015
rect 11265 1995 11285 2015
rect 11305 1995 11310 2015
rect 11240 1985 11310 1995
rect 11335 2115 11365 2125
rect 11335 2095 11340 2115
rect 11360 2095 11365 2115
rect 11335 2065 11365 2095
rect 11335 2045 11340 2065
rect 11360 2045 11365 2065
rect 11335 2015 11365 2045
rect 11335 1995 11340 2015
rect 11360 1995 11365 2015
rect 11335 1985 11365 1995
rect 11390 2115 11420 2125
rect 11390 2095 11395 2115
rect 11415 2095 11420 2115
rect 11390 2065 11420 2095
rect 11390 2045 11395 2065
rect 11415 2045 11420 2065
rect 11390 2015 11420 2045
rect 11390 1995 11395 2015
rect 11415 1995 11420 2015
rect 11390 1985 11420 1995
rect 11445 2115 11475 2125
rect 11445 2095 11450 2115
rect 11470 2095 11475 2115
rect 11445 2065 11475 2095
rect 11445 2045 11450 2065
rect 11470 2045 11475 2065
rect 11445 2015 11475 2045
rect 11445 1995 11450 2015
rect 11470 1995 11475 2015
rect 11445 1985 11475 1995
rect 11500 2115 11530 2125
rect 11500 2095 11505 2115
rect 11525 2095 11530 2115
rect 11500 2065 11530 2095
rect 11500 2045 11505 2065
rect 11525 2045 11530 2065
rect 11500 2015 11530 2045
rect 11500 1995 11505 2015
rect 11525 1995 11530 2015
rect 11500 1985 11530 1995
rect 11555 2115 11585 2125
rect 11555 2095 11560 2115
rect 11580 2095 11585 2115
rect 11555 2065 11585 2095
rect 11555 2045 11560 2065
rect 11580 2045 11585 2065
rect 11555 2015 11585 2045
rect 11555 1995 11560 2015
rect 11580 1995 11585 2015
rect 11555 1985 11585 1995
rect 11610 2115 11640 2125
rect 11610 2095 11615 2115
rect 11635 2095 11640 2115
rect 11610 2065 11640 2095
rect 11610 2045 11615 2065
rect 11635 2045 11640 2065
rect 11610 2015 11640 2045
rect 11610 1995 11615 2015
rect 11635 1995 11640 2015
rect 11610 1985 11640 1995
rect 11665 2115 11695 2125
rect 11665 2095 11670 2115
rect 11690 2095 11695 2115
rect 11665 2065 11695 2095
rect 11665 2045 11670 2065
rect 11690 2045 11695 2065
rect 11665 2015 11695 2045
rect 11665 1995 11670 2015
rect 11690 1995 11695 2015
rect 11665 1985 11695 1995
rect 11720 2115 11750 2125
rect 11720 2095 11725 2115
rect 11745 2095 11750 2115
rect 11720 2065 11750 2095
rect 11720 2045 11725 2065
rect 11745 2045 11750 2065
rect 11720 2015 11750 2045
rect 11720 1995 11725 2015
rect 11745 1995 11750 2015
rect 11720 1985 11750 1995
rect 11775 2115 11805 2125
rect 11775 2095 11780 2115
rect 11800 2095 11805 2115
rect 11775 2065 11805 2095
rect 11775 2045 11780 2065
rect 11800 2045 11805 2065
rect 11775 2015 11805 2045
rect 11775 1995 11780 2015
rect 11800 1995 11805 2015
rect 11775 1985 11805 1995
rect 11830 2115 11860 2125
rect 11830 2095 11835 2115
rect 11855 2095 11860 2115
rect 11830 2065 11860 2095
rect 11830 2045 11835 2065
rect 11855 2045 11860 2065
rect 11830 2015 11860 2045
rect 11830 1995 11835 2015
rect 11855 1995 11860 2015
rect 11830 1985 11860 1995
rect 11885 2115 11915 2125
rect 11885 2095 11890 2115
rect 11910 2095 11915 2115
rect 11885 2065 11915 2095
rect 11885 2045 11890 2065
rect 11910 2045 11915 2065
rect 11885 2015 11915 2045
rect 11885 1995 11890 2015
rect 11910 1995 11915 2015
rect 11885 1985 11915 1995
rect 11940 2115 11970 2125
rect 11940 2095 11945 2115
rect 11965 2095 11970 2115
rect 11940 2065 11970 2095
rect 11940 2045 11945 2065
rect 11965 2045 11970 2065
rect 11940 2015 11970 2045
rect 11940 1995 11945 2015
rect 11965 1995 11970 2015
rect 11940 1985 11970 1995
rect 11995 2115 12025 2125
rect 11995 2095 12000 2115
rect 12020 2095 12025 2115
rect 11995 2065 12025 2095
rect 11995 2045 12000 2065
rect 12020 2045 12025 2065
rect 11995 2015 12025 2045
rect 11995 1995 12000 2015
rect 12020 1995 12025 2015
rect 11995 1985 12025 1995
rect 12050 2115 12080 2125
rect 12050 2095 12055 2115
rect 12075 2095 12080 2115
rect 12050 2065 12080 2095
rect 12050 2045 12055 2065
rect 12075 2045 12080 2065
rect 12050 2015 12080 2045
rect 12050 1995 12055 2015
rect 12075 1995 12080 2015
rect 12050 1985 12080 1995
rect 12105 2115 12135 2125
rect 12105 2095 12110 2115
rect 12130 2095 12135 2115
rect 12105 2065 12135 2095
rect 12105 2045 12110 2065
rect 12130 2045 12135 2065
rect 12105 2015 12135 2045
rect 12105 1995 12110 2015
rect 12130 1995 12135 2015
rect 12105 1985 12135 1995
rect 12160 2115 12190 2125
rect 12160 2095 12165 2115
rect 12185 2095 12190 2115
rect 12160 2065 12190 2095
rect 12160 2045 12165 2065
rect 12185 2045 12190 2065
rect 12160 2015 12190 2045
rect 12160 1995 12165 2015
rect 12185 1995 12190 2015
rect 12160 1985 12190 1995
rect 12215 2115 12245 2125
rect 12215 2095 12220 2115
rect 12240 2095 12245 2115
rect 12215 2065 12245 2095
rect 12215 2045 12220 2065
rect 12240 2045 12245 2065
rect 12215 2015 12245 2045
rect 12215 1995 12220 2015
rect 12240 1995 12245 2015
rect 12215 1985 12245 1995
rect 12270 2115 12300 2125
rect 12270 2095 12275 2115
rect 12295 2095 12300 2115
rect 12270 2065 12300 2095
rect 12270 2045 12275 2065
rect 12295 2045 12300 2065
rect 12270 2015 12300 2045
rect 12270 1995 12275 2015
rect 12295 1995 12300 2015
rect 12270 1985 12300 1995
rect 12325 2115 12355 2125
rect 12325 2095 12330 2115
rect 12350 2095 12355 2115
rect 12325 2065 12355 2095
rect 12325 2045 12330 2065
rect 12350 2045 12355 2065
rect 12325 2015 12355 2045
rect 12325 1995 12330 2015
rect 12350 1995 12355 2015
rect 12325 1985 12355 1995
rect 12380 2115 12410 2125
rect 12380 2095 12385 2115
rect 12405 2095 12410 2115
rect 12380 2065 12410 2095
rect 12380 2045 12385 2065
rect 12405 2045 12410 2065
rect 12380 2015 12410 2045
rect 12380 1995 12385 2015
rect 12405 1995 12410 2015
rect 12380 1985 12410 1995
rect 12435 2115 12465 2125
rect 12435 2095 12440 2115
rect 12460 2095 12465 2115
rect 12435 2065 12465 2095
rect 12435 2045 12440 2065
rect 12460 2045 12465 2065
rect 12435 2015 12465 2045
rect 12435 1995 12440 2015
rect 12460 1995 12465 2015
rect 12435 1985 12465 1995
rect 12490 2115 12560 2125
rect 12490 2095 12495 2115
rect 12515 2095 12535 2115
rect 12555 2095 12560 2115
rect 12490 2065 12560 2095
rect 12490 2045 12495 2065
rect 12515 2045 12535 2065
rect 12555 2045 12560 2065
rect 12490 2015 12560 2045
rect 12855 2105 12925 2135
rect 12855 2085 12860 2105
rect 12880 2085 12900 2105
rect 12920 2085 12925 2105
rect 12855 2055 12925 2085
rect 12855 2035 12860 2055
rect 12880 2035 12900 2055
rect 12920 2035 12925 2055
rect 12855 2025 12925 2035
rect 12950 2155 12980 2165
rect 12950 2135 12955 2155
rect 12975 2135 12980 2155
rect 12950 2105 12980 2135
rect 12950 2085 12955 2105
rect 12975 2085 12980 2105
rect 12950 2055 12980 2085
rect 12950 2035 12955 2055
rect 12975 2035 12980 2055
rect 12950 2025 12980 2035
rect 13005 2155 13035 2165
rect 13005 2135 13010 2155
rect 13030 2135 13035 2155
rect 13005 2105 13035 2135
rect 13005 2085 13010 2105
rect 13030 2085 13035 2105
rect 13005 2055 13035 2085
rect 13005 2035 13010 2055
rect 13030 2035 13035 2055
rect 13005 2025 13035 2035
rect 13060 2155 13090 2165
rect 13060 2135 13065 2155
rect 13085 2135 13090 2155
rect 13060 2105 13090 2135
rect 13060 2085 13065 2105
rect 13085 2085 13090 2105
rect 13060 2055 13090 2085
rect 13060 2035 13065 2055
rect 13085 2035 13090 2055
rect 13060 2025 13090 2035
rect 13115 2155 13145 2165
rect 13115 2135 13120 2155
rect 13140 2135 13145 2155
rect 13115 2105 13145 2135
rect 13115 2085 13120 2105
rect 13140 2085 13145 2105
rect 13115 2055 13145 2085
rect 13115 2035 13120 2055
rect 13140 2035 13145 2055
rect 13115 2025 13145 2035
rect 13170 2155 13200 2165
rect 13170 2135 13175 2155
rect 13195 2135 13200 2155
rect 13170 2105 13200 2135
rect 13170 2085 13175 2105
rect 13195 2085 13200 2105
rect 13170 2055 13200 2085
rect 13170 2035 13175 2055
rect 13195 2035 13200 2055
rect 13170 2025 13200 2035
rect 13225 2155 13255 2165
rect 13225 2135 13230 2155
rect 13250 2135 13255 2155
rect 13225 2105 13255 2135
rect 13225 2085 13230 2105
rect 13250 2085 13255 2105
rect 13225 2055 13255 2085
rect 13225 2035 13230 2055
rect 13250 2035 13255 2055
rect 13225 2025 13255 2035
rect 13280 2155 13310 2165
rect 13280 2135 13285 2155
rect 13305 2135 13310 2155
rect 13280 2105 13310 2135
rect 13280 2085 13285 2105
rect 13305 2085 13310 2105
rect 13280 2055 13310 2085
rect 13280 2035 13285 2055
rect 13305 2035 13310 2055
rect 13280 2025 13310 2035
rect 13335 2155 13365 2165
rect 13335 2135 13340 2155
rect 13360 2135 13365 2155
rect 13335 2105 13365 2135
rect 13335 2085 13340 2105
rect 13360 2085 13365 2105
rect 13335 2055 13365 2085
rect 13335 2035 13340 2055
rect 13360 2035 13365 2055
rect 13335 2025 13365 2035
rect 13390 2155 13420 2165
rect 13390 2135 13395 2155
rect 13415 2135 13420 2155
rect 13390 2105 13420 2135
rect 13390 2085 13395 2105
rect 13415 2085 13420 2105
rect 13390 2055 13420 2085
rect 13390 2035 13395 2055
rect 13415 2035 13420 2055
rect 13390 2025 13420 2035
rect 13445 2155 13475 2165
rect 13445 2135 13450 2155
rect 13470 2135 13475 2155
rect 13445 2105 13475 2135
rect 13445 2085 13450 2105
rect 13470 2085 13475 2105
rect 13445 2055 13475 2085
rect 13445 2035 13450 2055
rect 13470 2035 13475 2055
rect 13445 2025 13475 2035
rect 13500 2155 13530 2165
rect 13500 2135 13505 2155
rect 13525 2135 13530 2155
rect 13500 2105 13530 2135
rect 13500 2085 13505 2105
rect 13525 2085 13530 2105
rect 13500 2055 13530 2085
rect 13500 2035 13505 2055
rect 13525 2035 13530 2055
rect 13500 2025 13530 2035
rect 13555 2155 13585 2165
rect 13555 2135 13560 2155
rect 13580 2135 13585 2155
rect 13555 2105 13585 2135
rect 13555 2085 13560 2105
rect 13580 2085 13585 2105
rect 13555 2055 13585 2085
rect 13555 2035 13560 2055
rect 13580 2035 13585 2055
rect 13555 2025 13585 2035
rect 13610 2155 13640 2165
rect 13610 2135 13615 2155
rect 13635 2135 13640 2155
rect 13610 2105 13640 2135
rect 13610 2085 13615 2105
rect 13635 2085 13640 2105
rect 13610 2055 13640 2085
rect 13610 2035 13615 2055
rect 13635 2035 13640 2055
rect 13610 2025 13640 2035
rect 13665 2155 13695 2165
rect 13665 2135 13670 2155
rect 13690 2135 13695 2155
rect 13665 2105 13695 2135
rect 13665 2085 13670 2105
rect 13690 2085 13695 2105
rect 13665 2055 13695 2085
rect 13665 2035 13670 2055
rect 13690 2035 13695 2055
rect 13665 2025 13695 2035
rect 13720 2155 13750 2165
rect 13720 2135 13725 2155
rect 13745 2135 13750 2155
rect 13720 2105 13750 2135
rect 13720 2085 13725 2105
rect 13745 2085 13750 2105
rect 13720 2055 13750 2085
rect 13720 2035 13725 2055
rect 13745 2035 13750 2055
rect 13720 2025 13750 2035
rect 13775 2155 13805 2165
rect 13775 2135 13780 2155
rect 13800 2135 13805 2155
rect 13775 2105 13805 2135
rect 13775 2085 13780 2105
rect 13800 2085 13805 2105
rect 13775 2055 13805 2085
rect 13775 2035 13780 2055
rect 13800 2035 13805 2055
rect 13775 2025 13805 2035
rect 13830 2155 13860 2165
rect 13830 2135 13835 2155
rect 13855 2135 13860 2155
rect 13830 2105 13860 2135
rect 13830 2085 13835 2105
rect 13855 2085 13860 2105
rect 13830 2055 13860 2085
rect 13830 2035 13835 2055
rect 13855 2035 13860 2055
rect 13830 2025 13860 2035
rect 13885 2155 13915 2165
rect 13885 2135 13890 2155
rect 13910 2135 13915 2155
rect 13885 2105 13915 2135
rect 13885 2085 13890 2105
rect 13910 2085 13915 2105
rect 13885 2055 13915 2085
rect 13885 2035 13890 2055
rect 13910 2035 13915 2055
rect 13885 2025 13915 2035
rect 13940 2155 13970 2165
rect 13940 2135 13945 2155
rect 13965 2135 13970 2155
rect 13940 2105 13970 2135
rect 13940 2085 13945 2105
rect 13965 2085 13970 2105
rect 13940 2055 13970 2085
rect 13940 2035 13945 2055
rect 13965 2035 13970 2055
rect 13940 2025 13970 2035
rect 13995 2155 14025 2165
rect 13995 2135 14000 2155
rect 14020 2135 14025 2155
rect 13995 2105 14025 2135
rect 13995 2085 14000 2105
rect 14020 2085 14025 2105
rect 13995 2055 14025 2085
rect 13995 2035 14000 2055
rect 14020 2035 14025 2055
rect 13995 2025 14025 2035
rect 14050 2155 14080 2165
rect 14050 2135 14055 2155
rect 14075 2135 14080 2155
rect 14050 2105 14080 2135
rect 14050 2085 14055 2105
rect 14075 2085 14080 2105
rect 14050 2055 14080 2085
rect 14050 2035 14055 2055
rect 14075 2035 14080 2055
rect 14050 2025 14080 2035
rect 14105 2155 14175 2165
rect 14105 2135 14110 2155
rect 14130 2135 14150 2155
rect 14170 2135 14175 2155
rect 14105 2105 14175 2135
rect 14105 2085 14110 2105
rect 14130 2085 14150 2105
rect 14170 2085 14175 2105
rect 14105 2055 14175 2085
rect 14105 2035 14110 2055
rect 14130 2035 14150 2055
rect 14170 2035 14175 2055
rect 14105 2025 14175 2035
rect 17145 2155 17215 2165
rect 17145 2135 17150 2155
rect 17170 2135 17190 2155
rect 17210 2135 17215 2155
rect 17145 2105 17215 2135
rect 17145 2085 17150 2105
rect 17170 2085 17190 2105
rect 17210 2085 17215 2105
rect 17145 2055 17215 2085
rect 17145 2035 17150 2055
rect 17170 2035 17190 2055
rect 17210 2035 17215 2055
rect 17145 2025 17215 2035
rect 17240 2155 17270 2165
rect 17240 2135 17245 2155
rect 17265 2135 17270 2155
rect 17240 2105 17270 2135
rect 17240 2085 17245 2105
rect 17265 2085 17270 2105
rect 17240 2055 17270 2085
rect 17240 2035 17245 2055
rect 17265 2035 17270 2055
rect 17240 2025 17270 2035
rect 17295 2155 17325 2165
rect 17295 2135 17300 2155
rect 17320 2135 17325 2155
rect 17295 2105 17325 2135
rect 17295 2085 17300 2105
rect 17320 2085 17325 2105
rect 17295 2055 17325 2085
rect 17295 2035 17300 2055
rect 17320 2035 17325 2055
rect 17295 2025 17325 2035
rect 17350 2155 17380 2165
rect 17350 2135 17355 2155
rect 17375 2135 17380 2155
rect 17350 2105 17380 2135
rect 17350 2085 17355 2105
rect 17375 2085 17380 2105
rect 17350 2055 17380 2085
rect 17350 2035 17355 2055
rect 17375 2035 17380 2055
rect 17350 2025 17380 2035
rect 17405 2155 17435 2165
rect 17405 2135 17410 2155
rect 17430 2135 17435 2155
rect 17405 2105 17435 2135
rect 17405 2085 17410 2105
rect 17430 2085 17435 2105
rect 17405 2055 17435 2085
rect 17405 2035 17410 2055
rect 17430 2035 17435 2055
rect 17405 2025 17435 2035
rect 17460 2155 17490 2165
rect 17460 2135 17465 2155
rect 17485 2135 17490 2155
rect 17460 2105 17490 2135
rect 17460 2085 17465 2105
rect 17485 2085 17490 2105
rect 17460 2055 17490 2085
rect 17460 2035 17465 2055
rect 17485 2035 17490 2055
rect 17460 2025 17490 2035
rect 17515 2155 17545 2165
rect 17515 2135 17520 2155
rect 17540 2135 17545 2155
rect 17515 2105 17545 2135
rect 17515 2085 17520 2105
rect 17540 2085 17545 2105
rect 17515 2055 17545 2085
rect 17515 2035 17520 2055
rect 17540 2035 17545 2055
rect 17515 2025 17545 2035
rect 17570 2155 17600 2165
rect 17570 2135 17575 2155
rect 17595 2135 17600 2155
rect 17570 2105 17600 2135
rect 17570 2085 17575 2105
rect 17595 2085 17600 2105
rect 17570 2055 17600 2085
rect 17570 2035 17575 2055
rect 17595 2035 17600 2055
rect 17570 2025 17600 2035
rect 17625 2155 17655 2165
rect 17625 2135 17630 2155
rect 17650 2135 17655 2155
rect 17625 2105 17655 2135
rect 17625 2085 17630 2105
rect 17650 2085 17655 2105
rect 17625 2055 17655 2085
rect 17625 2035 17630 2055
rect 17650 2035 17655 2055
rect 17625 2025 17655 2035
rect 17680 2155 17710 2165
rect 17680 2135 17685 2155
rect 17705 2135 17710 2155
rect 17680 2105 17710 2135
rect 17680 2085 17685 2105
rect 17705 2085 17710 2105
rect 17680 2055 17710 2085
rect 17680 2035 17685 2055
rect 17705 2035 17710 2055
rect 17680 2025 17710 2035
rect 17735 2155 17765 2165
rect 17735 2135 17740 2155
rect 17760 2135 17765 2155
rect 17735 2105 17765 2135
rect 17735 2085 17740 2105
rect 17760 2085 17765 2105
rect 17735 2055 17765 2085
rect 17735 2035 17740 2055
rect 17760 2035 17765 2055
rect 17735 2025 17765 2035
rect 17790 2155 17820 2165
rect 17790 2135 17795 2155
rect 17815 2135 17820 2155
rect 17790 2105 17820 2135
rect 17790 2085 17795 2105
rect 17815 2085 17820 2105
rect 17790 2055 17820 2085
rect 17790 2035 17795 2055
rect 17815 2035 17820 2055
rect 17790 2025 17820 2035
rect 17845 2155 17875 2165
rect 17845 2135 17850 2155
rect 17870 2135 17875 2155
rect 17845 2105 17875 2135
rect 17845 2085 17850 2105
rect 17870 2085 17875 2105
rect 17845 2055 17875 2085
rect 17845 2035 17850 2055
rect 17870 2035 17875 2055
rect 17845 2025 17875 2035
rect 17900 2155 17930 2165
rect 17900 2135 17905 2155
rect 17925 2135 17930 2155
rect 17900 2105 17930 2135
rect 17900 2085 17905 2105
rect 17925 2085 17930 2105
rect 17900 2055 17930 2085
rect 17900 2035 17905 2055
rect 17925 2035 17930 2055
rect 17900 2025 17930 2035
rect 17955 2155 17985 2165
rect 17955 2135 17960 2155
rect 17980 2135 17985 2155
rect 17955 2105 17985 2135
rect 17955 2085 17960 2105
rect 17980 2085 17985 2105
rect 17955 2055 17985 2085
rect 17955 2035 17960 2055
rect 17980 2035 17985 2055
rect 17955 2025 17985 2035
rect 18010 2155 18040 2165
rect 18010 2135 18015 2155
rect 18035 2135 18040 2155
rect 18010 2105 18040 2135
rect 18010 2085 18015 2105
rect 18035 2085 18040 2105
rect 18010 2055 18040 2085
rect 18010 2035 18015 2055
rect 18035 2035 18040 2055
rect 18010 2025 18040 2035
rect 18065 2155 18095 2165
rect 18065 2135 18070 2155
rect 18090 2135 18095 2155
rect 18065 2105 18095 2135
rect 18065 2085 18070 2105
rect 18090 2085 18095 2105
rect 18065 2055 18095 2085
rect 18065 2035 18070 2055
rect 18090 2035 18095 2055
rect 18065 2025 18095 2035
rect 18120 2155 18150 2165
rect 18120 2135 18125 2155
rect 18145 2135 18150 2155
rect 18120 2105 18150 2135
rect 18120 2085 18125 2105
rect 18145 2085 18150 2105
rect 18120 2055 18150 2085
rect 18120 2035 18125 2055
rect 18145 2035 18150 2055
rect 18120 2025 18150 2035
rect 18175 2155 18205 2165
rect 18175 2135 18180 2155
rect 18200 2135 18205 2155
rect 18175 2105 18205 2135
rect 18175 2085 18180 2105
rect 18200 2085 18205 2105
rect 18175 2055 18205 2085
rect 18175 2035 18180 2055
rect 18200 2035 18205 2055
rect 18175 2025 18205 2035
rect 18230 2155 18260 2165
rect 18230 2135 18235 2155
rect 18255 2135 18260 2155
rect 18230 2105 18260 2135
rect 18230 2085 18235 2105
rect 18255 2085 18260 2105
rect 18230 2055 18260 2085
rect 18230 2035 18235 2055
rect 18255 2035 18260 2055
rect 18230 2025 18260 2035
rect 18285 2155 18315 2165
rect 18285 2135 18290 2155
rect 18310 2135 18315 2155
rect 18285 2105 18315 2135
rect 18285 2085 18290 2105
rect 18310 2085 18315 2105
rect 18285 2055 18315 2085
rect 18285 2035 18290 2055
rect 18310 2035 18315 2055
rect 18285 2025 18315 2035
rect 18340 2155 18370 2165
rect 18340 2135 18345 2155
rect 18365 2135 18370 2155
rect 18340 2105 18370 2135
rect 18340 2085 18345 2105
rect 18365 2085 18370 2105
rect 18340 2055 18370 2085
rect 18340 2035 18345 2055
rect 18365 2035 18370 2055
rect 18340 2025 18370 2035
rect 18395 2155 18465 2165
rect 18395 2135 18400 2155
rect 18420 2135 18440 2155
rect 18460 2135 18465 2155
rect 18830 2155 18840 2175
rect 18860 2155 18870 2175
rect 18830 2145 18870 2155
rect 18940 2175 18980 2185
rect 18940 2155 18950 2175
rect 18970 2155 18980 2175
rect 18940 2145 18980 2155
rect 19050 2175 19090 2185
rect 19050 2155 19060 2175
rect 19080 2155 19090 2175
rect 19050 2145 19090 2155
rect 19160 2175 19200 2185
rect 19160 2155 19170 2175
rect 19190 2155 19200 2175
rect 19160 2145 19200 2155
rect 19270 2175 19310 2185
rect 19270 2155 19280 2175
rect 19300 2155 19310 2175
rect 19270 2145 19310 2155
rect 19380 2175 19420 2185
rect 19380 2155 19390 2175
rect 19410 2155 19420 2175
rect 19380 2145 19420 2155
rect 19490 2175 19530 2185
rect 19490 2155 19500 2175
rect 19520 2155 19530 2175
rect 19490 2145 19530 2155
rect 19600 2175 19640 2185
rect 19600 2155 19610 2175
rect 19630 2155 19640 2175
rect 19600 2145 19640 2155
rect 19710 2175 19750 2185
rect 19710 2155 19720 2175
rect 19740 2155 19750 2175
rect 19710 2145 19750 2155
rect 19820 2175 19860 2185
rect 19820 2155 19830 2175
rect 19850 2155 19860 2175
rect 19820 2145 19860 2155
rect 19930 2175 19970 2185
rect 19930 2155 19940 2175
rect 19960 2155 19970 2175
rect 20360 2165 20380 2185
rect 20510 2165 20530 2185
rect 20620 2165 20640 2185
rect 20730 2165 20750 2185
rect 20840 2165 20860 2185
rect 20950 2165 20970 2185
rect 21060 2165 21080 2185
rect 21170 2165 21190 2185
rect 21280 2165 21300 2185
rect 21390 2165 21410 2185
rect 21500 2165 21520 2185
rect 21650 2165 21670 2185
rect 19930 2145 19970 2155
rect 20355 2155 20425 2165
rect 18395 2105 18465 2135
rect 18840 2125 18860 2145
rect 18950 2125 18970 2145
rect 19060 2125 19080 2145
rect 19170 2125 19190 2145
rect 19280 2125 19300 2145
rect 19390 2125 19410 2145
rect 19500 2125 19520 2145
rect 19610 2125 19630 2145
rect 19720 2125 19740 2145
rect 19830 2125 19850 2145
rect 19940 2125 19960 2145
rect 20355 2135 20360 2155
rect 20380 2135 20400 2155
rect 20420 2135 20425 2155
rect 18395 2085 18400 2105
rect 18420 2085 18440 2105
rect 18460 2085 18465 2105
rect 18395 2055 18465 2085
rect 18395 2035 18400 2055
rect 18420 2035 18440 2055
rect 18460 2035 18465 2055
rect 18395 2025 18465 2035
rect 18740 2115 18810 2125
rect 18740 2095 18745 2115
rect 18765 2095 18785 2115
rect 18805 2095 18810 2115
rect 18740 2065 18810 2095
rect 18740 2045 18745 2065
rect 18765 2045 18785 2065
rect 18805 2045 18810 2065
rect 12490 1995 12495 2015
rect 12515 1995 12535 2015
rect 12555 1995 12560 2015
rect 12955 2005 12975 2025
rect 13065 2005 13085 2025
rect 13175 2005 13195 2025
rect 13285 2005 13305 2025
rect 13395 2005 13415 2025
rect 13505 2005 13525 2025
rect 13615 2005 13635 2025
rect 13725 2005 13745 2025
rect 13835 2005 13855 2025
rect 13945 2005 13965 2025
rect 14055 2005 14075 2025
rect 17245 2005 17265 2025
rect 17355 2005 17375 2025
rect 17465 2005 17485 2025
rect 17575 2005 17595 2025
rect 17685 2005 17705 2025
rect 17795 2005 17815 2025
rect 17905 2005 17925 2025
rect 18015 2005 18035 2025
rect 18125 2005 18145 2025
rect 18235 2005 18255 2025
rect 18345 2005 18365 2025
rect 18740 2015 18810 2045
rect 12490 1985 12560 1995
rect 12945 1995 12985 2005
rect 10835 1965 10875 1975
rect 11245 1965 11265 1985
rect 11395 1965 11415 1985
rect 11505 1965 11525 1985
rect 11615 1965 11635 1985
rect 11725 1965 11745 1985
rect 11835 1965 11855 1985
rect 11945 1965 11965 1985
rect 12055 1965 12075 1985
rect 12165 1965 12185 1985
rect 12275 1965 12295 1985
rect 12385 1965 12405 1985
rect 12535 1965 12555 1985
rect 12945 1975 12957 1995
rect 12975 1975 12985 1995
rect 12945 1965 12985 1975
rect 13055 1995 13095 2005
rect 13055 1975 13067 1995
rect 13085 1975 13095 1995
rect 13055 1965 13095 1975
rect 13165 1995 13205 2005
rect 13165 1975 13177 1995
rect 13195 1975 13205 1995
rect 13165 1965 13205 1975
rect 13275 1995 13315 2005
rect 13275 1975 13287 1995
rect 13305 1975 13315 1995
rect 13275 1965 13315 1975
rect 13385 1995 13425 2005
rect 13385 1975 13397 1995
rect 13415 1975 13425 1995
rect 13385 1965 13425 1975
rect 13495 1995 13535 2005
rect 13495 1975 13507 1995
rect 13525 1975 13535 1995
rect 13495 1965 13535 1975
rect 13605 1995 13645 2005
rect 13605 1975 13617 1995
rect 13635 1975 13645 1995
rect 13605 1965 13645 1975
rect 13715 1995 13755 2005
rect 13715 1975 13727 1995
rect 13745 1975 13755 1995
rect 13715 1965 13755 1975
rect 13825 1995 13865 2005
rect 13825 1975 13837 1995
rect 13855 1975 13865 1995
rect 13825 1965 13865 1975
rect 13935 1995 13975 2005
rect 13935 1975 13947 1995
rect 13965 1975 13975 1995
rect 13935 1965 13975 1975
rect 14045 1995 14085 2005
rect 14045 1975 14057 1995
rect 14075 1975 14085 1995
rect 14045 1965 14085 1975
rect 17235 1995 17275 2005
rect 17235 1975 17245 1995
rect 17263 1975 17275 1995
rect 17235 1965 17275 1975
rect 17345 1995 17385 2005
rect 17345 1975 17355 1995
rect 17373 1975 17385 1995
rect 17345 1965 17385 1975
rect 17455 1995 17495 2005
rect 17455 1975 17465 1995
rect 17483 1975 17495 1995
rect 17455 1965 17495 1975
rect 17565 1995 17605 2005
rect 17565 1975 17575 1995
rect 17593 1975 17605 1995
rect 17565 1965 17605 1975
rect 17675 1995 17715 2005
rect 17675 1975 17685 1995
rect 17703 1975 17715 1995
rect 17675 1965 17715 1975
rect 17785 1995 17825 2005
rect 17785 1975 17795 1995
rect 17813 1975 17825 1995
rect 17785 1965 17825 1975
rect 17895 1995 17935 2005
rect 17895 1975 17905 1995
rect 17923 1975 17935 1995
rect 17895 1965 17935 1975
rect 18005 1995 18045 2005
rect 18005 1975 18015 1995
rect 18033 1975 18045 1995
rect 18005 1965 18045 1975
rect 18115 1995 18155 2005
rect 18115 1975 18125 1995
rect 18143 1975 18155 1995
rect 18115 1965 18155 1975
rect 18225 1995 18265 2005
rect 18225 1975 18235 1995
rect 18253 1975 18265 1995
rect 18225 1965 18265 1975
rect 18335 1995 18375 2005
rect 18335 1975 18345 1995
rect 18363 1975 18375 1995
rect 18740 1995 18745 2015
rect 18765 1995 18785 2015
rect 18805 1995 18810 2015
rect 18740 1985 18810 1995
rect 18835 2115 18865 2125
rect 18835 2095 18840 2115
rect 18860 2095 18865 2115
rect 18835 2065 18865 2095
rect 18835 2045 18840 2065
rect 18860 2045 18865 2065
rect 18835 2015 18865 2045
rect 18835 1995 18840 2015
rect 18860 1995 18865 2015
rect 18835 1985 18865 1995
rect 18890 2115 18920 2125
rect 18890 2095 18895 2115
rect 18915 2095 18920 2115
rect 18890 2065 18920 2095
rect 18890 2045 18895 2065
rect 18915 2045 18920 2065
rect 18890 2015 18920 2045
rect 18890 1995 18895 2015
rect 18915 1995 18920 2015
rect 18890 1985 18920 1995
rect 18945 2115 18975 2125
rect 18945 2095 18950 2115
rect 18970 2095 18975 2115
rect 18945 2065 18975 2095
rect 18945 2045 18950 2065
rect 18970 2045 18975 2065
rect 18945 2015 18975 2045
rect 18945 1995 18950 2015
rect 18970 1995 18975 2015
rect 18945 1985 18975 1995
rect 19000 2115 19030 2125
rect 19000 2095 19005 2115
rect 19025 2095 19030 2115
rect 19000 2065 19030 2095
rect 19000 2045 19005 2065
rect 19025 2045 19030 2065
rect 19000 2015 19030 2045
rect 19000 1995 19005 2015
rect 19025 1995 19030 2015
rect 19000 1985 19030 1995
rect 19055 2115 19085 2125
rect 19055 2095 19060 2115
rect 19080 2095 19085 2115
rect 19055 2065 19085 2095
rect 19055 2045 19060 2065
rect 19080 2045 19085 2065
rect 19055 2015 19085 2045
rect 19055 1995 19060 2015
rect 19080 1995 19085 2015
rect 19055 1985 19085 1995
rect 19110 2115 19140 2125
rect 19110 2095 19115 2115
rect 19135 2095 19140 2115
rect 19110 2065 19140 2095
rect 19110 2045 19115 2065
rect 19135 2045 19140 2065
rect 19110 2015 19140 2045
rect 19110 1995 19115 2015
rect 19135 1995 19140 2015
rect 19110 1985 19140 1995
rect 19165 2115 19195 2125
rect 19165 2095 19170 2115
rect 19190 2095 19195 2115
rect 19165 2065 19195 2095
rect 19165 2045 19170 2065
rect 19190 2045 19195 2065
rect 19165 2015 19195 2045
rect 19165 1995 19170 2015
rect 19190 1995 19195 2015
rect 19165 1985 19195 1995
rect 19220 2115 19250 2125
rect 19220 2095 19225 2115
rect 19245 2095 19250 2115
rect 19220 2065 19250 2095
rect 19220 2045 19225 2065
rect 19245 2045 19250 2065
rect 19220 2015 19250 2045
rect 19220 1995 19225 2015
rect 19245 1995 19250 2015
rect 19220 1985 19250 1995
rect 19275 2115 19305 2125
rect 19275 2095 19280 2115
rect 19300 2095 19305 2115
rect 19275 2065 19305 2095
rect 19275 2045 19280 2065
rect 19300 2045 19305 2065
rect 19275 2015 19305 2045
rect 19275 1995 19280 2015
rect 19300 1995 19305 2015
rect 19275 1985 19305 1995
rect 19330 2115 19360 2125
rect 19330 2095 19335 2115
rect 19355 2095 19360 2115
rect 19330 2065 19360 2095
rect 19330 2045 19335 2065
rect 19355 2045 19360 2065
rect 19330 2015 19360 2045
rect 19330 1995 19335 2015
rect 19355 1995 19360 2015
rect 19330 1985 19360 1995
rect 19385 2115 19415 2125
rect 19385 2095 19390 2115
rect 19410 2095 19415 2115
rect 19385 2065 19415 2095
rect 19385 2045 19390 2065
rect 19410 2045 19415 2065
rect 19385 2015 19415 2045
rect 19385 1995 19390 2015
rect 19410 1995 19415 2015
rect 19385 1985 19415 1995
rect 19440 2115 19470 2125
rect 19440 2095 19445 2115
rect 19465 2095 19470 2115
rect 19440 2065 19470 2095
rect 19440 2045 19445 2065
rect 19465 2045 19470 2065
rect 19440 2015 19470 2045
rect 19440 1995 19445 2015
rect 19465 1995 19470 2015
rect 19440 1985 19470 1995
rect 19495 2115 19525 2125
rect 19495 2095 19500 2115
rect 19520 2095 19525 2115
rect 19495 2065 19525 2095
rect 19495 2045 19500 2065
rect 19520 2045 19525 2065
rect 19495 2015 19525 2045
rect 19495 1995 19500 2015
rect 19520 1995 19525 2015
rect 19495 1985 19525 1995
rect 19550 2115 19580 2125
rect 19550 2095 19555 2115
rect 19575 2095 19580 2115
rect 19550 2065 19580 2095
rect 19550 2045 19555 2065
rect 19575 2045 19580 2065
rect 19550 2015 19580 2045
rect 19550 1995 19555 2015
rect 19575 1995 19580 2015
rect 19550 1985 19580 1995
rect 19605 2115 19635 2125
rect 19605 2095 19610 2115
rect 19630 2095 19635 2115
rect 19605 2065 19635 2095
rect 19605 2045 19610 2065
rect 19630 2045 19635 2065
rect 19605 2015 19635 2045
rect 19605 1995 19610 2015
rect 19630 1995 19635 2015
rect 19605 1985 19635 1995
rect 19660 2115 19690 2125
rect 19660 2095 19665 2115
rect 19685 2095 19690 2115
rect 19660 2065 19690 2095
rect 19660 2045 19665 2065
rect 19685 2045 19690 2065
rect 19660 2015 19690 2045
rect 19660 1995 19665 2015
rect 19685 1995 19690 2015
rect 19660 1985 19690 1995
rect 19715 2115 19745 2125
rect 19715 2095 19720 2115
rect 19740 2095 19745 2115
rect 19715 2065 19745 2095
rect 19715 2045 19720 2065
rect 19740 2045 19745 2065
rect 19715 2015 19745 2045
rect 19715 1995 19720 2015
rect 19740 1995 19745 2015
rect 19715 1985 19745 1995
rect 19770 2115 19800 2125
rect 19770 2095 19775 2115
rect 19795 2095 19800 2115
rect 19770 2065 19800 2095
rect 19770 2045 19775 2065
rect 19795 2045 19800 2065
rect 19770 2015 19800 2045
rect 19770 1995 19775 2015
rect 19795 1995 19800 2015
rect 19770 1985 19800 1995
rect 19825 2115 19855 2125
rect 19825 2095 19830 2115
rect 19850 2095 19855 2115
rect 19825 2065 19855 2095
rect 19825 2045 19830 2065
rect 19850 2045 19855 2065
rect 19825 2015 19855 2045
rect 19825 1995 19830 2015
rect 19850 1995 19855 2015
rect 19825 1985 19855 1995
rect 19880 2115 19910 2125
rect 19880 2095 19885 2115
rect 19905 2095 19910 2115
rect 19880 2065 19910 2095
rect 19880 2045 19885 2065
rect 19905 2045 19910 2065
rect 19880 2015 19910 2045
rect 19880 1995 19885 2015
rect 19905 1995 19910 2015
rect 19880 1985 19910 1995
rect 19935 2115 19965 2125
rect 19935 2095 19940 2115
rect 19960 2095 19965 2115
rect 19935 2065 19965 2095
rect 19935 2045 19940 2065
rect 19960 2045 19965 2065
rect 19935 2015 19965 2045
rect 19935 1995 19940 2015
rect 19960 1995 19965 2015
rect 19935 1985 19965 1995
rect 19990 2115 20060 2125
rect 19990 2095 19995 2115
rect 20015 2095 20035 2115
rect 20055 2095 20060 2115
rect 19990 2065 20060 2095
rect 19990 2045 19995 2065
rect 20015 2045 20035 2065
rect 20055 2045 20060 2065
rect 19990 2015 20060 2045
rect 20355 2105 20425 2135
rect 20355 2085 20360 2105
rect 20380 2085 20400 2105
rect 20420 2085 20425 2105
rect 20355 2055 20425 2085
rect 20355 2035 20360 2055
rect 20380 2035 20400 2055
rect 20420 2035 20425 2055
rect 20355 2025 20425 2035
rect 20450 2155 20480 2165
rect 20450 2135 20455 2155
rect 20475 2135 20480 2155
rect 20450 2105 20480 2135
rect 20450 2085 20455 2105
rect 20475 2085 20480 2105
rect 20450 2055 20480 2085
rect 20450 2035 20455 2055
rect 20475 2035 20480 2055
rect 20450 2025 20480 2035
rect 20505 2155 20535 2165
rect 20505 2135 20510 2155
rect 20530 2135 20535 2155
rect 20505 2105 20535 2135
rect 20505 2085 20510 2105
rect 20530 2085 20535 2105
rect 20505 2055 20535 2085
rect 20505 2035 20510 2055
rect 20530 2035 20535 2055
rect 20505 2025 20535 2035
rect 20560 2155 20590 2165
rect 20560 2135 20565 2155
rect 20585 2135 20590 2155
rect 20560 2105 20590 2135
rect 20560 2085 20565 2105
rect 20585 2085 20590 2105
rect 20560 2055 20590 2085
rect 20560 2035 20565 2055
rect 20585 2035 20590 2055
rect 20560 2025 20590 2035
rect 20615 2155 20645 2165
rect 20615 2135 20620 2155
rect 20640 2135 20645 2155
rect 20615 2105 20645 2135
rect 20615 2085 20620 2105
rect 20640 2085 20645 2105
rect 20615 2055 20645 2085
rect 20615 2035 20620 2055
rect 20640 2035 20645 2055
rect 20615 2025 20645 2035
rect 20670 2155 20700 2165
rect 20670 2135 20675 2155
rect 20695 2135 20700 2155
rect 20670 2105 20700 2135
rect 20670 2085 20675 2105
rect 20695 2085 20700 2105
rect 20670 2055 20700 2085
rect 20670 2035 20675 2055
rect 20695 2035 20700 2055
rect 20670 2025 20700 2035
rect 20725 2155 20755 2165
rect 20725 2135 20730 2155
rect 20750 2135 20755 2155
rect 20725 2105 20755 2135
rect 20725 2085 20730 2105
rect 20750 2085 20755 2105
rect 20725 2055 20755 2085
rect 20725 2035 20730 2055
rect 20750 2035 20755 2055
rect 20725 2025 20755 2035
rect 20780 2155 20810 2165
rect 20780 2135 20785 2155
rect 20805 2135 20810 2155
rect 20780 2105 20810 2135
rect 20780 2085 20785 2105
rect 20805 2085 20810 2105
rect 20780 2055 20810 2085
rect 20780 2035 20785 2055
rect 20805 2035 20810 2055
rect 20780 2025 20810 2035
rect 20835 2155 20865 2165
rect 20835 2135 20840 2155
rect 20860 2135 20865 2155
rect 20835 2105 20865 2135
rect 20835 2085 20840 2105
rect 20860 2085 20865 2105
rect 20835 2055 20865 2085
rect 20835 2035 20840 2055
rect 20860 2035 20865 2055
rect 20835 2025 20865 2035
rect 20890 2155 20920 2165
rect 20890 2135 20895 2155
rect 20915 2135 20920 2155
rect 20890 2105 20920 2135
rect 20890 2085 20895 2105
rect 20915 2085 20920 2105
rect 20890 2055 20920 2085
rect 20890 2035 20895 2055
rect 20915 2035 20920 2055
rect 20890 2025 20920 2035
rect 20945 2155 20975 2165
rect 20945 2135 20950 2155
rect 20970 2135 20975 2155
rect 20945 2105 20975 2135
rect 20945 2085 20950 2105
rect 20970 2085 20975 2105
rect 20945 2055 20975 2085
rect 20945 2035 20950 2055
rect 20970 2035 20975 2055
rect 20945 2025 20975 2035
rect 21000 2155 21030 2165
rect 21000 2135 21005 2155
rect 21025 2135 21030 2155
rect 21000 2105 21030 2135
rect 21000 2085 21005 2105
rect 21025 2085 21030 2105
rect 21000 2055 21030 2085
rect 21000 2035 21005 2055
rect 21025 2035 21030 2055
rect 21000 2025 21030 2035
rect 21055 2155 21085 2165
rect 21055 2135 21060 2155
rect 21080 2135 21085 2155
rect 21055 2105 21085 2135
rect 21055 2085 21060 2105
rect 21080 2085 21085 2105
rect 21055 2055 21085 2085
rect 21055 2035 21060 2055
rect 21080 2035 21085 2055
rect 21055 2025 21085 2035
rect 21110 2155 21140 2165
rect 21110 2135 21115 2155
rect 21135 2135 21140 2155
rect 21110 2105 21140 2135
rect 21110 2085 21115 2105
rect 21135 2085 21140 2105
rect 21110 2055 21140 2085
rect 21110 2035 21115 2055
rect 21135 2035 21140 2055
rect 21110 2025 21140 2035
rect 21165 2155 21195 2165
rect 21165 2135 21170 2155
rect 21190 2135 21195 2155
rect 21165 2105 21195 2135
rect 21165 2085 21170 2105
rect 21190 2085 21195 2105
rect 21165 2055 21195 2085
rect 21165 2035 21170 2055
rect 21190 2035 21195 2055
rect 21165 2025 21195 2035
rect 21220 2155 21250 2165
rect 21220 2135 21225 2155
rect 21245 2135 21250 2155
rect 21220 2105 21250 2135
rect 21220 2085 21225 2105
rect 21245 2085 21250 2105
rect 21220 2055 21250 2085
rect 21220 2035 21225 2055
rect 21245 2035 21250 2055
rect 21220 2025 21250 2035
rect 21275 2155 21305 2165
rect 21275 2135 21280 2155
rect 21300 2135 21305 2155
rect 21275 2105 21305 2135
rect 21275 2085 21280 2105
rect 21300 2085 21305 2105
rect 21275 2055 21305 2085
rect 21275 2035 21280 2055
rect 21300 2035 21305 2055
rect 21275 2025 21305 2035
rect 21330 2155 21360 2165
rect 21330 2135 21335 2155
rect 21355 2135 21360 2155
rect 21330 2105 21360 2135
rect 21330 2085 21335 2105
rect 21355 2085 21360 2105
rect 21330 2055 21360 2085
rect 21330 2035 21335 2055
rect 21355 2035 21360 2055
rect 21330 2025 21360 2035
rect 21385 2155 21415 2165
rect 21385 2135 21390 2155
rect 21410 2135 21415 2155
rect 21385 2105 21415 2135
rect 21385 2085 21390 2105
rect 21410 2085 21415 2105
rect 21385 2055 21415 2085
rect 21385 2035 21390 2055
rect 21410 2035 21415 2055
rect 21385 2025 21415 2035
rect 21440 2155 21470 2165
rect 21440 2135 21445 2155
rect 21465 2135 21470 2155
rect 21440 2105 21470 2135
rect 21440 2085 21445 2105
rect 21465 2085 21470 2105
rect 21440 2055 21470 2085
rect 21440 2035 21445 2055
rect 21465 2035 21470 2055
rect 21440 2025 21470 2035
rect 21495 2155 21525 2165
rect 21495 2135 21500 2155
rect 21520 2135 21525 2155
rect 21495 2105 21525 2135
rect 21495 2085 21500 2105
rect 21520 2085 21525 2105
rect 21495 2055 21525 2085
rect 21495 2035 21500 2055
rect 21520 2035 21525 2055
rect 21495 2025 21525 2035
rect 21550 2155 21580 2165
rect 21550 2135 21555 2155
rect 21575 2135 21580 2155
rect 21550 2105 21580 2135
rect 21550 2085 21555 2105
rect 21575 2085 21580 2105
rect 21550 2055 21580 2085
rect 21550 2035 21555 2055
rect 21575 2035 21580 2055
rect 21550 2025 21580 2035
rect 21605 2155 21675 2165
rect 21605 2135 21610 2155
rect 21630 2135 21650 2155
rect 21670 2135 21675 2155
rect 21605 2105 21675 2135
rect 21605 2085 21610 2105
rect 21630 2085 21650 2105
rect 21670 2085 21675 2105
rect 21605 2055 21675 2085
rect 21605 2035 21610 2055
rect 21630 2035 21650 2055
rect 21670 2035 21675 2055
rect 21605 2025 21675 2035
rect 19990 1995 19995 2015
rect 20015 1995 20035 2015
rect 20055 1995 20060 2015
rect 20455 2005 20475 2025
rect 20565 2005 20585 2025
rect 20675 2005 20695 2025
rect 20785 2005 20805 2025
rect 20895 2005 20915 2025
rect 21005 2005 21025 2025
rect 21115 2005 21135 2025
rect 21225 2005 21245 2025
rect 21335 2005 21355 2025
rect 21445 2005 21465 2025
rect 21555 2005 21575 2025
rect 19990 1985 20060 1995
rect 20445 1995 20485 2005
rect 18335 1965 18375 1975
rect 18745 1965 18765 1985
rect 18895 1965 18915 1985
rect 19005 1965 19025 1985
rect 19115 1965 19135 1985
rect 19225 1965 19245 1985
rect 19335 1965 19355 1985
rect 19445 1965 19465 1985
rect 19555 1965 19575 1985
rect 19665 1965 19685 1985
rect 19775 1965 19795 1985
rect 19885 1965 19905 1985
rect 20035 1965 20055 1985
rect 20445 1975 20457 1995
rect 20475 1975 20485 1995
rect 20445 1965 20485 1975
rect 20555 1995 20595 2005
rect 20555 1975 20567 1995
rect 20585 1975 20595 1995
rect 20555 1965 20595 1975
rect 20665 1995 20705 2005
rect 20665 1975 20677 1995
rect 20695 1975 20705 1995
rect 20665 1965 20705 1975
rect 20775 1995 20815 2005
rect 20775 1975 20787 1995
rect 20805 1975 20815 1995
rect 20775 1965 20815 1975
rect 20885 1995 20925 2005
rect 20885 1975 20897 1995
rect 20915 1975 20925 1995
rect 20885 1965 20925 1975
rect 20995 1995 21035 2005
rect 20995 1975 21007 1995
rect 21025 1975 21035 1995
rect 20995 1965 21035 1975
rect 21105 1995 21145 2005
rect 21105 1975 21117 1995
rect 21135 1975 21145 1995
rect 21105 1965 21145 1975
rect 21215 1995 21255 2005
rect 21215 1975 21227 1995
rect 21245 1975 21255 1995
rect 21215 1965 21255 1975
rect 21325 1995 21365 2005
rect 21325 1975 21337 1995
rect 21355 1975 21365 1995
rect 21325 1965 21365 1975
rect 21435 1995 21475 2005
rect 21435 1975 21447 1995
rect 21465 1975 21475 1995
rect 21435 1965 21475 1975
rect 21545 1995 21585 2005
rect 21545 1975 21557 1995
rect 21575 1975 21585 1995
rect 21545 1965 21585 1975
rect 5230 1935 5260 1965
rect 5230 1915 5235 1935
rect 5255 1915 5260 1935
rect 11235 1955 11275 1965
rect 11235 1935 11245 1955
rect 11265 1935 11275 1955
rect 11235 1925 11275 1935
rect 11385 1955 11425 1965
rect 11385 1935 11395 1955
rect 11415 1935 11425 1955
rect 11385 1925 11425 1935
rect 11495 1955 11535 1965
rect 11495 1935 11505 1955
rect 11525 1935 11535 1955
rect 11495 1925 11535 1935
rect 11605 1955 11645 1965
rect 11605 1935 11615 1955
rect 11635 1935 11645 1955
rect 11605 1925 11645 1935
rect 11715 1955 11755 1965
rect 11715 1935 11725 1955
rect 11745 1935 11755 1955
rect 11715 1925 11755 1935
rect 11825 1955 11865 1965
rect 11825 1935 11835 1955
rect 11855 1935 11865 1955
rect 11825 1925 11865 1935
rect 11935 1955 11975 1965
rect 11935 1935 11945 1955
rect 11965 1935 11975 1955
rect 11935 1925 11975 1935
rect 12045 1955 12085 1965
rect 12045 1935 12055 1955
rect 12075 1935 12085 1955
rect 12045 1925 12085 1935
rect 12155 1955 12195 1965
rect 12155 1935 12165 1955
rect 12185 1935 12195 1955
rect 12155 1925 12195 1935
rect 12265 1955 12305 1965
rect 12265 1935 12275 1955
rect 12295 1935 12305 1955
rect 12265 1925 12305 1935
rect 12375 1955 12415 1965
rect 12375 1935 12385 1955
rect 12405 1935 12415 1955
rect 12375 1925 12415 1935
rect 12525 1955 12565 1965
rect 12525 1935 12535 1955
rect 12555 1935 12565 1955
rect 12525 1925 12565 1935
rect 18735 1955 18775 1965
rect 18735 1935 18745 1955
rect 18765 1935 18775 1955
rect 18735 1925 18775 1935
rect 18885 1955 18925 1965
rect 18885 1935 18895 1955
rect 18915 1935 18925 1955
rect 18885 1925 18925 1935
rect 18995 1955 19035 1965
rect 18995 1935 19005 1955
rect 19025 1935 19035 1955
rect 18995 1925 19035 1935
rect 19105 1955 19145 1965
rect 19105 1935 19115 1955
rect 19135 1935 19145 1955
rect 19105 1925 19145 1935
rect 19215 1955 19255 1965
rect 19215 1935 19225 1955
rect 19245 1935 19255 1955
rect 19215 1925 19255 1935
rect 19325 1955 19365 1965
rect 19325 1935 19335 1955
rect 19355 1935 19365 1955
rect 19325 1925 19365 1935
rect 19435 1955 19475 1965
rect 19435 1935 19445 1955
rect 19465 1935 19475 1955
rect 19435 1925 19475 1935
rect 19545 1955 19585 1965
rect 19545 1935 19555 1955
rect 19575 1935 19585 1955
rect 19545 1925 19585 1935
rect 19655 1955 19695 1965
rect 19655 1935 19665 1955
rect 19685 1935 19695 1955
rect 19655 1925 19695 1935
rect 19765 1955 19805 1965
rect 19765 1935 19775 1955
rect 19795 1935 19805 1955
rect 19765 1925 19805 1935
rect 19875 1955 19915 1965
rect 19875 1935 19885 1955
rect 19905 1935 19915 1955
rect 19875 1925 19915 1935
rect 20025 1955 20065 1965
rect 20025 1935 20035 1955
rect 20055 1935 20065 1955
rect 20025 1925 20065 1935
rect 5230 1905 5260 1915
rect 2575 1885 2595 1905
rect 2685 1885 2705 1905
rect 2755 1885 2775 1905
rect 2935 1885 2955 1905
rect 3055 1885 3075 1905
rect 3295 1885 3315 1905
rect 3415 1885 3435 1905
rect 3655 1885 3675 1905
rect 3775 1885 3795 1905
rect 2565 1875 2600 1885
rect 2565 1855 2575 1875
rect 2595 1855 2600 1875
rect 2565 1845 2600 1855
rect 2620 1875 2660 1885
rect 2620 1855 2630 1875
rect 2650 1855 2660 1875
rect 2620 1845 2660 1855
rect 2680 1875 2715 1885
rect 2680 1855 2685 1875
rect 2705 1855 2715 1875
rect 2680 1845 2715 1855
rect 2755 1875 2805 1885
rect 2755 1855 2775 1875
rect 2795 1855 2805 1875
rect 2755 1845 2805 1855
rect 2835 1875 2875 1885
rect 2835 1855 2845 1875
rect 2865 1855 2875 1875
rect 2835 1845 2875 1855
rect 2925 1875 2965 1885
rect 2925 1855 2935 1875
rect 2955 1855 2965 1875
rect 2925 1845 2965 1855
rect 3045 1875 3085 1885
rect 3045 1855 3055 1875
rect 3075 1855 3085 1875
rect 3045 1845 3085 1855
rect 3165 1875 3205 1885
rect 3165 1855 3175 1875
rect 3195 1855 3205 1875
rect 3165 1845 3205 1855
rect 3285 1875 3325 1885
rect 3285 1855 3295 1875
rect 3315 1855 3325 1875
rect 3285 1845 3325 1855
rect 3405 1875 3445 1885
rect 3405 1855 3415 1875
rect 3435 1855 3445 1875
rect 3405 1845 3445 1855
rect 3525 1875 3565 1885
rect 3525 1855 3535 1875
rect 3555 1855 3565 1875
rect 3525 1845 3565 1855
rect 3645 1875 3685 1885
rect 3645 1855 3655 1875
rect 3675 1855 3685 1875
rect 3645 1845 3685 1855
rect 3765 1875 3805 1885
rect 3765 1855 3775 1875
rect 3795 1855 3805 1875
rect 3765 1845 3805 1855
rect 3855 1875 3895 1885
rect 3995 1880 4015 1905
rect 4215 1885 4235 1905
rect 4335 1885 4355 1905
rect 4575 1885 4595 1905
rect 4695 1885 4715 1905
rect 4935 1885 4955 1905
rect 5055 1885 5075 1905
rect 5235 1885 5255 1905
rect 3855 1855 3865 1875
rect 3885 1855 3895 1875
rect 3855 1845 3895 1855
rect 3985 1870 4025 1880
rect 3985 1850 3995 1870
rect 4015 1850 4025 1870
rect 3985 1840 4025 1850
rect 4115 1875 4155 1885
rect 4115 1855 4125 1875
rect 4145 1855 4155 1875
rect 4115 1845 4155 1855
rect 4205 1875 4245 1885
rect 4205 1855 4215 1875
rect 4235 1855 4245 1875
rect 4205 1845 4245 1855
rect 4325 1875 4365 1885
rect 4325 1855 4335 1875
rect 4355 1855 4365 1875
rect 4325 1845 4365 1855
rect 4445 1875 4485 1885
rect 4445 1855 4455 1875
rect 4475 1855 4485 1875
rect 4445 1845 4485 1855
rect 4565 1875 4605 1885
rect 4565 1855 4575 1875
rect 4595 1855 4605 1875
rect 4565 1845 4605 1855
rect 4685 1875 4725 1885
rect 4685 1855 4695 1875
rect 4715 1855 4725 1875
rect 4685 1845 4725 1855
rect 4805 1875 4845 1885
rect 4805 1855 4815 1875
rect 4835 1855 4845 1875
rect 4805 1845 4845 1855
rect 4925 1875 4965 1885
rect 4925 1855 4935 1875
rect 4955 1855 4965 1875
rect 4925 1845 4965 1855
rect 5045 1875 5085 1885
rect 5045 1855 5055 1875
rect 5075 1855 5085 1875
rect 5045 1845 5085 1855
rect 5135 1875 5175 1885
rect 5135 1855 5145 1875
rect 5165 1855 5175 1875
rect 5135 1845 5175 1855
rect 5205 1875 5255 1885
rect 5205 1855 5215 1875
rect 5235 1855 5255 1875
rect 20450 1900 20490 1910
rect 20450 1880 20460 1900
rect 20480 1880 20490 1900
rect 20450 1870 20490 1880
rect 20545 1900 20585 1910
rect 20545 1880 20555 1900
rect 20575 1880 20585 1900
rect 20545 1870 20585 1880
rect 20655 1900 20695 1910
rect 20655 1880 20665 1900
rect 20685 1880 20695 1900
rect 20655 1870 20695 1880
rect 20765 1900 20805 1910
rect 20765 1880 20775 1900
rect 20795 1880 20805 1900
rect 20765 1870 20805 1880
rect 20860 1900 20900 1910
rect 20860 1880 20870 1900
rect 20890 1880 20900 1900
rect 20860 1870 20900 1880
rect 5205 1845 5255 1855
rect 20460 1850 20480 1870
rect 20555 1850 20575 1870
rect 20665 1850 20685 1870
rect 20775 1850 20795 1870
rect 20870 1850 20890 1870
rect 20455 1840 20525 1850
rect 2475 1790 2505 1820
rect 2835 1785 2875 1825
rect 3045 1815 3085 1825
rect 3045 1795 3055 1815
rect 3075 1795 3085 1815
rect 3045 1785 3085 1795
rect 3165 1785 3205 1825
rect 3405 1815 3445 1825
rect 3405 1795 3415 1815
rect 3435 1795 3445 1815
rect 3405 1785 3445 1795
rect 3525 1785 3565 1825
rect 3765 1815 3805 1825
rect 3765 1795 3775 1815
rect 3795 1795 3805 1815
rect 3765 1785 3805 1795
rect 3855 1785 3895 1825
rect 4115 1785 4155 1825
rect 4205 1815 4245 1825
rect 4205 1795 4215 1815
rect 4235 1795 4245 1815
rect 4205 1785 4245 1795
rect 4445 1785 4485 1825
rect 4565 1815 4605 1825
rect 4565 1795 4575 1815
rect 4595 1795 4605 1815
rect 4565 1785 4605 1795
rect 4805 1785 4845 1825
rect 4925 1815 4965 1825
rect 4925 1795 4935 1815
rect 4955 1795 4965 1815
rect 4925 1785 4965 1795
rect 5135 1785 5175 1825
rect 20455 1820 20460 1840
rect 20480 1820 20500 1840
rect 20520 1820 20525 1840
rect 5365 1790 5395 1820
rect 20455 1790 20525 1820
rect 11190 1770 11230 1780
rect 2430 1730 2460 1760
rect 2570 1730 2600 1760
rect 2680 1730 2710 1760
rect 2805 1735 2835 1765
rect 3225 1755 3265 1765
rect 3225 1735 3235 1755
rect 3255 1735 3265 1755
rect 3225 1725 3265 1735
rect 3285 1755 3325 1765
rect 3285 1735 3295 1755
rect 3315 1735 3325 1755
rect 3285 1725 3325 1735
rect 3525 1755 3565 1765
rect 3525 1735 3535 1755
rect 3555 1735 3565 1755
rect 3525 1725 3565 1735
rect 3765 1755 3805 1765
rect 3765 1735 3775 1755
rect 3795 1735 3805 1755
rect 3765 1725 3805 1735
rect 4205 1755 4245 1765
rect 4205 1735 4215 1755
rect 4235 1735 4245 1755
rect 4205 1725 4245 1735
rect 4445 1755 4485 1765
rect 4445 1735 4455 1755
rect 4475 1735 4485 1755
rect 4445 1725 4485 1735
rect 4685 1755 4725 1765
rect 4685 1735 4695 1755
rect 4715 1735 4725 1755
rect 4685 1725 4725 1735
rect 4745 1755 4785 1765
rect 4745 1735 4755 1755
rect 4775 1735 4785 1755
rect 4745 1725 4785 1735
rect 5275 1730 5305 1760
rect 11085 1755 11125 1765
rect 11085 1735 11095 1755
rect 11115 1735 11125 1755
rect 11190 1750 11200 1770
rect 11220 1750 11230 1770
rect 11410 1770 11450 1780
rect 11190 1740 11230 1750
rect 11305 1755 11345 1765
rect 11085 1725 11125 1735
rect 3165 1710 3205 1720
rect 2805 1680 2835 1710
rect 3165 1690 3175 1710
rect 3195 1690 3205 1710
rect 3165 1680 3205 1690
rect 2385 1635 2415 1665
rect 2625 1635 2655 1665
rect 3175 1660 3195 1680
rect 3295 1660 3315 1725
rect 3405 1710 3445 1720
rect 3405 1690 3415 1710
rect 3435 1690 3445 1710
rect 3405 1680 3445 1690
rect 3415 1660 3435 1680
rect 3535 1660 3555 1725
rect 3645 1710 3685 1720
rect 3645 1690 3655 1710
rect 3675 1690 3685 1710
rect 3645 1680 3685 1690
rect 3655 1660 3675 1680
rect 3775 1660 3795 1725
rect 4215 1660 4235 1725
rect 4325 1710 4365 1720
rect 4325 1690 4335 1710
rect 4355 1690 4365 1710
rect 4325 1680 4365 1690
rect 4335 1660 4355 1680
rect 4455 1660 4475 1725
rect 4565 1710 4605 1720
rect 4565 1690 4575 1710
rect 4595 1690 4605 1710
rect 4565 1680 4605 1690
rect 4575 1660 4595 1680
rect 4695 1660 4715 1725
rect 4805 1710 4845 1720
rect 4805 1690 4815 1710
rect 4835 1690 4845 1710
rect 4805 1680 4845 1690
rect 4815 1660 4835 1680
rect 11095 1660 11115 1725
rect 11200 1660 11220 1740
rect 11305 1735 11315 1755
rect 11335 1735 11345 1755
rect 11410 1750 11420 1770
rect 11440 1750 11450 1770
rect 11640 1770 11680 1780
rect 11410 1740 11450 1750
rect 11525 1755 11565 1765
rect 11305 1725 11345 1735
rect 11237 1710 11269 1720
rect 11237 1690 11243 1710
rect 11260 1690 11269 1710
rect 11237 1680 11269 1690
rect 11315 1660 11335 1725
rect 11420 1660 11440 1740
rect 11525 1735 11535 1755
rect 11555 1735 11565 1755
rect 11640 1750 11650 1770
rect 11670 1750 11680 1770
rect 12230 1770 12270 1780
rect 11640 1740 11680 1750
rect 12125 1755 12165 1765
rect 11525 1725 11565 1735
rect 11457 1710 11489 1720
rect 11457 1690 11463 1710
rect 11480 1690 11489 1710
rect 11457 1680 11489 1690
rect 11535 1660 11555 1725
rect 11601 1710 11633 1720
rect 11601 1690 11610 1710
rect 11627 1690 11633 1710
rect 11601 1680 11633 1690
rect 11650 1660 11670 1740
rect 12125 1735 12135 1755
rect 12155 1735 12165 1755
rect 12230 1750 12240 1770
rect 12260 1750 12270 1770
rect 12450 1770 12490 1780
rect 12230 1740 12270 1750
rect 12345 1755 12385 1765
rect 12125 1725 12165 1735
rect 11820 1710 11850 1720
rect 11820 1690 11825 1710
rect 11845 1690 11850 1710
rect 11820 1680 11850 1690
rect 11867 1710 11899 1720
rect 11867 1690 11876 1710
rect 11893 1690 11899 1710
rect 11867 1680 11899 1690
rect 11950 1710 11980 1720
rect 11950 1690 11955 1710
rect 11975 1690 11980 1710
rect 11950 1680 11980 1690
rect 11830 1660 11850 1680
rect 11950 1660 11970 1680
rect 12135 1660 12155 1725
rect 12240 1660 12260 1740
rect 12345 1735 12355 1755
rect 12375 1735 12385 1755
rect 12450 1750 12460 1770
rect 12480 1750 12490 1770
rect 12680 1770 12720 1780
rect 12450 1740 12490 1750
rect 12565 1755 12605 1765
rect 12345 1725 12385 1735
rect 12277 1710 12309 1720
rect 12277 1690 12283 1710
rect 12300 1690 12309 1710
rect 12277 1680 12309 1690
rect 12355 1660 12375 1725
rect 12460 1660 12480 1740
rect 12565 1735 12575 1755
rect 12595 1735 12605 1755
rect 12680 1750 12690 1770
rect 12710 1750 12720 1770
rect 18690 1770 18730 1780
rect 12680 1740 12720 1750
rect 18585 1755 18625 1765
rect 12565 1725 12605 1735
rect 12497 1710 12529 1720
rect 12497 1690 12503 1710
rect 12520 1690 12529 1710
rect 12497 1680 12529 1690
rect 12575 1660 12595 1725
rect 12641 1710 12673 1720
rect 12641 1690 12650 1710
rect 12667 1690 12673 1710
rect 12641 1680 12673 1690
rect 12690 1660 12710 1740
rect 18585 1735 18595 1755
rect 18615 1735 18625 1755
rect 18690 1750 18700 1770
rect 18720 1750 18730 1770
rect 18910 1770 18950 1780
rect 18690 1740 18730 1750
rect 18805 1755 18845 1765
rect 18585 1725 18625 1735
rect 18595 1660 18615 1725
rect 18700 1660 18720 1740
rect 18805 1735 18815 1755
rect 18835 1735 18845 1755
rect 18910 1750 18920 1770
rect 18940 1750 18950 1770
rect 19140 1770 19180 1780
rect 18910 1740 18950 1750
rect 19025 1755 19065 1765
rect 18805 1725 18845 1735
rect 18737 1710 18769 1720
rect 18737 1690 18743 1710
rect 18760 1690 18769 1710
rect 18737 1680 18769 1690
rect 18815 1660 18835 1725
rect 18920 1660 18940 1740
rect 19025 1735 19035 1755
rect 19055 1735 19065 1755
rect 19140 1750 19150 1770
rect 19170 1750 19180 1770
rect 19730 1770 19770 1780
rect 19140 1740 19180 1750
rect 19625 1755 19665 1765
rect 19025 1725 19065 1735
rect 18957 1710 18989 1720
rect 18957 1690 18963 1710
rect 18980 1690 18989 1710
rect 18957 1680 18989 1690
rect 19035 1660 19055 1725
rect 19101 1710 19133 1720
rect 19101 1690 19110 1710
rect 19127 1690 19133 1710
rect 19101 1680 19133 1690
rect 19150 1660 19170 1740
rect 19625 1735 19635 1755
rect 19655 1735 19665 1755
rect 19730 1750 19740 1770
rect 19760 1750 19770 1770
rect 19950 1770 19990 1780
rect 19730 1740 19770 1750
rect 19845 1755 19885 1765
rect 19625 1725 19665 1735
rect 19320 1710 19350 1720
rect 19320 1690 19325 1710
rect 19345 1690 19350 1710
rect 19320 1680 19350 1690
rect 19367 1710 19399 1720
rect 19367 1690 19376 1710
rect 19393 1690 19399 1710
rect 19367 1680 19399 1690
rect 19450 1710 19480 1720
rect 19450 1690 19455 1710
rect 19475 1690 19480 1710
rect 19450 1680 19480 1690
rect 19330 1660 19350 1680
rect 19450 1660 19470 1680
rect 19635 1660 19655 1725
rect 19740 1660 19760 1740
rect 19845 1735 19855 1755
rect 19875 1735 19885 1755
rect 19950 1750 19960 1770
rect 19980 1750 19990 1770
rect 20180 1770 20220 1780
rect 19950 1740 19990 1750
rect 20065 1755 20105 1765
rect 19845 1725 19885 1735
rect 19777 1710 19809 1720
rect 19777 1690 19783 1710
rect 19800 1690 19809 1710
rect 19777 1680 19809 1690
rect 19855 1660 19875 1725
rect 19960 1660 19980 1740
rect 20065 1735 20075 1755
rect 20095 1735 20105 1755
rect 20180 1750 20190 1770
rect 20210 1750 20220 1770
rect 20180 1740 20220 1750
rect 20455 1770 20460 1790
rect 20480 1770 20500 1790
rect 20520 1770 20525 1790
rect 20455 1740 20525 1770
rect 20065 1725 20105 1735
rect 19997 1710 20029 1720
rect 19997 1690 20003 1710
rect 20020 1690 20029 1710
rect 19997 1680 20029 1690
rect 20075 1660 20095 1725
rect 20141 1710 20173 1720
rect 20141 1690 20150 1710
rect 20167 1690 20173 1710
rect 20141 1680 20173 1690
rect 20190 1660 20210 1740
rect 20455 1720 20460 1740
rect 20480 1720 20500 1740
rect 20520 1720 20525 1740
rect 20455 1710 20525 1720
rect 20550 1840 20580 1850
rect 20550 1820 20555 1840
rect 20575 1820 20580 1840
rect 20550 1790 20580 1820
rect 20550 1770 20555 1790
rect 20575 1770 20580 1790
rect 20550 1740 20580 1770
rect 20550 1720 20555 1740
rect 20575 1720 20580 1740
rect 20550 1710 20580 1720
rect 20605 1840 20635 1850
rect 20605 1820 20610 1840
rect 20630 1820 20635 1840
rect 20605 1790 20635 1820
rect 20605 1770 20610 1790
rect 20630 1770 20635 1790
rect 20605 1740 20635 1770
rect 20605 1720 20610 1740
rect 20630 1720 20635 1740
rect 20605 1710 20635 1720
rect 20660 1840 20690 1850
rect 20660 1820 20665 1840
rect 20685 1820 20690 1840
rect 20660 1790 20690 1820
rect 20660 1770 20665 1790
rect 20685 1770 20690 1790
rect 20660 1740 20690 1770
rect 20660 1720 20665 1740
rect 20685 1720 20690 1740
rect 20660 1710 20690 1720
rect 20715 1840 20745 1850
rect 20715 1820 20720 1840
rect 20740 1820 20745 1840
rect 20715 1790 20745 1820
rect 20715 1770 20720 1790
rect 20740 1770 20745 1790
rect 20715 1740 20745 1770
rect 20715 1720 20720 1740
rect 20740 1720 20745 1740
rect 20715 1710 20745 1720
rect 20770 1840 20800 1850
rect 20770 1820 20775 1840
rect 20795 1820 20800 1840
rect 20770 1790 20800 1820
rect 20770 1770 20775 1790
rect 20795 1770 20800 1790
rect 20770 1740 20800 1770
rect 20770 1720 20775 1740
rect 20795 1720 20800 1740
rect 20770 1710 20800 1720
rect 20825 1840 20895 1850
rect 20825 1820 20830 1840
rect 20850 1820 20870 1840
rect 20890 1820 20895 1840
rect 20825 1790 20895 1820
rect 20825 1770 20830 1790
rect 20850 1770 20870 1790
rect 20890 1770 20895 1790
rect 20825 1740 20895 1770
rect 20825 1720 20830 1740
rect 20850 1720 20870 1740
rect 20890 1720 20895 1740
rect 20825 1710 20895 1720
rect 20615 1690 20635 1710
rect 20720 1690 20740 1710
rect 20566 1675 20598 1685
rect 3170 1650 3200 1660
rect 3170 1630 3175 1650
rect 3195 1630 3200 1650
rect 3170 1620 3200 1630
rect 3230 1650 3260 1660
rect 3230 1630 3235 1650
rect 3255 1630 3260 1650
rect 3230 1620 3260 1630
rect 3290 1650 3320 1660
rect 3290 1630 3295 1650
rect 3315 1630 3320 1650
rect 3290 1620 3320 1630
rect 3350 1650 3380 1660
rect 3350 1630 3355 1650
rect 3375 1630 3380 1650
rect 3350 1620 3380 1630
rect 3410 1650 3440 1660
rect 3410 1630 3415 1650
rect 3435 1630 3440 1650
rect 3410 1620 3440 1630
rect 3470 1650 3500 1660
rect 3470 1630 3475 1650
rect 3495 1630 3500 1650
rect 3470 1620 3500 1630
rect 3530 1650 3560 1660
rect 3530 1630 3535 1650
rect 3555 1630 3560 1650
rect 3530 1620 3560 1630
rect 3590 1650 3620 1660
rect 3590 1630 3595 1650
rect 3615 1630 3620 1650
rect 3590 1620 3620 1630
rect 3650 1650 3680 1660
rect 3650 1630 3655 1650
rect 3675 1630 3680 1650
rect 3650 1620 3680 1630
rect 3710 1650 3740 1660
rect 3710 1630 3715 1650
rect 3735 1630 3740 1650
rect 3710 1620 3740 1630
rect 3770 1650 3800 1660
rect 3770 1630 3775 1650
rect 3795 1630 3800 1650
rect 3770 1620 3800 1630
rect 3985 1650 4025 1660
rect 3985 1630 3995 1650
rect 4015 1630 4025 1650
rect 3985 1620 4025 1630
rect 4210 1650 4240 1660
rect 4210 1630 4215 1650
rect 4235 1630 4240 1650
rect 4210 1620 4240 1630
rect 4270 1650 4300 1660
rect 4270 1630 4275 1650
rect 4295 1630 4300 1650
rect 4270 1620 4300 1630
rect 4330 1650 4360 1660
rect 4330 1630 4335 1650
rect 4355 1630 4360 1650
rect 4330 1620 4360 1630
rect 4390 1650 4420 1660
rect 4390 1630 4395 1650
rect 4415 1630 4420 1650
rect 4390 1620 4420 1630
rect 4450 1650 4480 1660
rect 4450 1630 4455 1650
rect 4475 1630 4480 1650
rect 4450 1620 4480 1630
rect 4510 1650 4540 1660
rect 4510 1630 4515 1650
rect 4535 1630 4540 1650
rect 4510 1620 4540 1630
rect 4570 1650 4600 1660
rect 4570 1630 4575 1650
rect 4595 1630 4600 1650
rect 4570 1620 4600 1630
rect 4630 1650 4660 1660
rect 4630 1630 4635 1650
rect 4655 1630 4660 1650
rect 4630 1620 4660 1630
rect 4690 1650 4720 1660
rect 4690 1630 4695 1650
rect 4715 1630 4720 1650
rect 4690 1620 4720 1630
rect 4750 1650 4780 1660
rect 4750 1630 4755 1650
rect 4775 1630 4780 1650
rect 4750 1620 4780 1630
rect 4810 1650 4840 1660
rect 4810 1630 4815 1650
rect 4835 1630 4840 1650
rect 4810 1620 4840 1630
rect 10990 1650 11065 1660
rect 10990 1630 11000 1650
rect 11020 1630 11040 1650
rect 11060 1630 11065 1650
rect 2335 1565 2365 1595
rect 3165 1590 3205 1600
rect 3165 1570 3175 1590
rect 3195 1570 3205 1590
rect 3165 1560 3205 1570
rect 3235 1550 3255 1620
rect 3355 1550 3375 1620
rect 3475 1550 3495 1620
rect 3595 1550 3615 1620
rect 3715 1550 3735 1620
rect 4275 1550 4295 1620
rect 4395 1550 4415 1620
rect 4515 1550 4535 1620
rect 4635 1550 4655 1620
rect 4755 1550 4775 1620
rect 10990 1600 11065 1630
rect 4805 1590 4845 1600
rect 4805 1570 4815 1590
rect 4835 1570 4845 1590
rect 4805 1560 4845 1570
rect 5415 1565 5445 1595
rect 10990 1580 11000 1600
rect 11020 1580 11040 1600
rect 11060 1580 11065 1600
rect 10990 1550 11065 1580
rect 3225 1540 3265 1550
rect 3225 1520 3235 1540
rect 3255 1520 3265 1540
rect 3225 1510 3265 1520
rect 3345 1540 3385 1550
rect 3345 1520 3355 1540
rect 3375 1520 3385 1540
rect 3345 1510 3385 1520
rect 3465 1540 3505 1550
rect 3465 1520 3475 1540
rect 3495 1520 3505 1540
rect 3465 1510 3505 1520
rect 3585 1540 3625 1550
rect 3585 1520 3595 1540
rect 3615 1520 3625 1540
rect 3585 1510 3625 1520
rect 3705 1540 3745 1550
rect 3705 1520 3715 1540
rect 3735 1520 3745 1540
rect 3705 1510 3745 1520
rect 4265 1540 4305 1550
rect 4265 1520 4275 1540
rect 4295 1520 4305 1540
rect 4265 1510 4305 1520
rect 4385 1540 4425 1550
rect 4385 1520 4395 1540
rect 4415 1520 4425 1540
rect 4385 1510 4425 1520
rect 4505 1540 4545 1550
rect 4505 1520 4515 1540
rect 4535 1520 4545 1540
rect 4505 1510 4545 1520
rect 4625 1540 4665 1550
rect 4625 1520 4635 1540
rect 4655 1520 4665 1540
rect 4625 1510 4665 1520
rect 4745 1540 4785 1550
rect 4745 1520 4755 1540
rect 4775 1520 4785 1540
rect 10990 1530 11000 1550
rect 11020 1530 11040 1550
rect 11060 1530 11065 1550
rect 10990 1520 11065 1530
rect 11090 1650 11120 1660
rect 11090 1630 11095 1650
rect 11115 1630 11120 1650
rect 11090 1600 11120 1630
rect 11090 1580 11095 1600
rect 11115 1580 11120 1600
rect 11090 1550 11120 1580
rect 11090 1530 11095 1550
rect 11115 1530 11120 1550
rect 11090 1520 11120 1530
rect 11145 1650 11175 1660
rect 11145 1630 11150 1650
rect 11170 1630 11175 1650
rect 11145 1600 11175 1630
rect 11145 1580 11150 1600
rect 11170 1580 11175 1600
rect 11145 1550 11175 1580
rect 11145 1530 11150 1550
rect 11170 1530 11175 1550
rect 11145 1520 11175 1530
rect 11200 1650 11230 1660
rect 11200 1630 11205 1650
rect 11225 1630 11230 1650
rect 11200 1600 11230 1630
rect 11200 1580 11205 1600
rect 11225 1580 11230 1600
rect 11200 1550 11230 1580
rect 11200 1530 11205 1550
rect 11225 1530 11230 1550
rect 11200 1520 11230 1530
rect 11255 1650 11285 1660
rect 11255 1630 11260 1650
rect 11280 1630 11285 1650
rect 11255 1600 11285 1630
rect 11255 1580 11260 1600
rect 11280 1580 11285 1600
rect 11255 1550 11285 1580
rect 11255 1530 11260 1550
rect 11280 1530 11285 1550
rect 11255 1520 11285 1530
rect 11310 1650 11340 1660
rect 11310 1630 11315 1650
rect 11335 1630 11340 1650
rect 11310 1600 11340 1630
rect 11310 1580 11315 1600
rect 11335 1580 11340 1600
rect 11310 1550 11340 1580
rect 11310 1530 11315 1550
rect 11335 1530 11340 1550
rect 11310 1520 11340 1530
rect 11365 1650 11395 1660
rect 11365 1630 11370 1650
rect 11390 1630 11395 1650
rect 11365 1600 11395 1630
rect 11365 1580 11370 1600
rect 11390 1580 11395 1600
rect 11365 1550 11395 1580
rect 11365 1530 11370 1550
rect 11390 1530 11395 1550
rect 11365 1520 11395 1530
rect 11420 1650 11450 1660
rect 11420 1630 11425 1650
rect 11445 1630 11450 1650
rect 11420 1600 11450 1630
rect 11420 1580 11425 1600
rect 11445 1580 11450 1600
rect 11420 1550 11450 1580
rect 11420 1530 11425 1550
rect 11445 1530 11450 1550
rect 11420 1520 11450 1530
rect 11475 1650 11505 1660
rect 11475 1630 11480 1650
rect 11500 1630 11505 1650
rect 11475 1600 11505 1630
rect 11475 1580 11480 1600
rect 11500 1580 11505 1600
rect 11475 1550 11505 1580
rect 11475 1530 11480 1550
rect 11500 1530 11505 1550
rect 11475 1520 11505 1530
rect 11530 1650 11560 1660
rect 11530 1630 11535 1650
rect 11555 1630 11560 1650
rect 11530 1600 11560 1630
rect 11530 1580 11535 1600
rect 11555 1580 11560 1600
rect 11530 1550 11560 1580
rect 11530 1530 11535 1550
rect 11555 1530 11560 1550
rect 11530 1520 11560 1530
rect 11585 1650 11615 1660
rect 11585 1630 11590 1650
rect 11610 1630 11615 1650
rect 11585 1600 11615 1630
rect 11585 1580 11590 1600
rect 11610 1580 11615 1600
rect 11585 1550 11615 1580
rect 11585 1530 11590 1550
rect 11610 1530 11615 1550
rect 11585 1520 11615 1530
rect 11640 1650 11670 1660
rect 11640 1630 11645 1650
rect 11665 1630 11670 1650
rect 11640 1600 11670 1630
rect 11640 1580 11645 1600
rect 11665 1580 11670 1600
rect 11640 1550 11670 1580
rect 11640 1530 11645 1550
rect 11665 1530 11670 1550
rect 11640 1520 11670 1530
rect 11695 1650 11805 1660
rect 11695 1630 11700 1650
rect 11720 1630 11740 1650
rect 11760 1630 11780 1650
rect 11800 1630 11805 1650
rect 11695 1600 11805 1630
rect 11695 1580 11700 1600
rect 11720 1580 11740 1600
rect 11760 1580 11780 1600
rect 11800 1580 11805 1600
rect 11695 1550 11805 1580
rect 11695 1530 11700 1550
rect 11720 1530 11740 1550
rect 11760 1530 11780 1550
rect 11800 1530 11805 1550
rect 11695 1520 11805 1530
rect 11830 1650 11860 1660
rect 11830 1630 11835 1650
rect 11855 1630 11860 1650
rect 11830 1600 11860 1630
rect 11830 1580 11835 1600
rect 11855 1580 11860 1600
rect 11830 1550 11860 1580
rect 11830 1530 11835 1550
rect 11855 1530 11860 1550
rect 11830 1520 11860 1530
rect 11885 1650 11915 1660
rect 11885 1630 11890 1650
rect 11910 1630 11915 1650
rect 11885 1600 11915 1630
rect 11885 1580 11890 1600
rect 11910 1580 11915 1600
rect 11885 1550 11915 1580
rect 11885 1530 11890 1550
rect 11910 1530 11915 1550
rect 11885 1520 11915 1530
rect 11940 1650 11970 1660
rect 11940 1630 11945 1650
rect 11965 1630 11970 1650
rect 11940 1600 11970 1630
rect 11940 1580 11945 1600
rect 11965 1580 11970 1600
rect 11940 1550 11970 1580
rect 11940 1530 11945 1550
rect 11965 1530 11970 1550
rect 11940 1520 11970 1530
rect 11995 1650 12105 1660
rect 11995 1630 12000 1650
rect 12020 1630 12040 1650
rect 12060 1630 12080 1650
rect 12100 1630 12105 1650
rect 11995 1600 12105 1630
rect 11995 1580 12000 1600
rect 12020 1580 12040 1600
rect 12060 1580 12080 1600
rect 12100 1580 12105 1600
rect 11995 1550 12105 1580
rect 11995 1530 12000 1550
rect 12020 1530 12040 1550
rect 12060 1530 12080 1550
rect 12100 1530 12105 1550
rect 11995 1520 12105 1530
rect 12130 1650 12160 1660
rect 12130 1630 12135 1650
rect 12155 1630 12160 1650
rect 12130 1600 12160 1630
rect 12130 1580 12135 1600
rect 12155 1580 12160 1600
rect 12130 1550 12160 1580
rect 12130 1530 12135 1550
rect 12155 1530 12160 1550
rect 12130 1520 12160 1530
rect 12185 1650 12215 1660
rect 12185 1630 12190 1650
rect 12210 1630 12215 1650
rect 12185 1600 12215 1630
rect 12185 1580 12190 1600
rect 12210 1580 12215 1600
rect 12185 1550 12215 1580
rect 12185 1530 12190 1550
rect 12210 1530 12215 1550
rect 12185 1520 12215 1530
rect 12240 1650 12270 1660
rect 12240 1630 12245 1650
rect 12265 1630 12270 1650
rect 12240 1600 12270 1630
rect 12240 1580 12245 1600
rect 12265 1580 12270 1600
rect 12240 1550 12270 1580
rect 12240 1530 12245 1550
rect 12265 1530 12270 1550
rect 12240 1520 12270 1530
rect 12295 1650 12325 1660
rect 12295 1630 12300 1650
rect 12320 1630 12325 1650
rect 12295 1600 12325 1630
rect 12295 1580 12300 1600
rect 12320 1580 12325 1600
rect 12295 1550 12325 1580
rect 12295 1530 12300 1550
rect 12320 1530 12325 1550
rect 12295 1520 12325 1530
rect 12350 1650 12380 1660
rect 12350 1630 12355 1650
rect 12375 1630 12380 1650
rect 12350 1600 12380 1630
rect 12350 1580 12355 1600
rect 12375 1580 12380 1600
rect 12350 1550 12380 1580
rect 12350 1530 12355 1550
rect 12375 1530 12380 1550
rect 12350 1520 12380 1530
rect 12405 1650 12435 1660
rect 12405 1630 12410 1650
rect 12430 1630 12435 1650
rect 12405 1600 12435 1630
rect 12405 1580 12410 1600
rect 12430 1580 12435 1600
rect 12405 1550 12435 1580
rect 12405 1530 12410 1550
rect 12430 1530 12435 1550
rect 12405 1520 12435 1530
rect 12460 1650 12490 1660
rect 12460 1630 12465 1650
rect 12485 1630 12490 1650
rect 12460 1600 12490 1630
rect 12460 1580 12465 1600
rect 12485 1580 12490 1600
rect 12460 1550 12490 1580
rect 12460 1530 12465 1550
rect 12485 1530 12490 1550
rect 12460 1520 12490 1530
rect 12515 1650 12545 1660
rect 12515 1630 12520 1650
rect 12540 1630 12545 1650
rect 12515 1600 12545 1630
rect 12515 1580 12520 1600
rect 12540 1580 12545 1600
rect 12515 1550 12545 1580
rect 12515 1530 12520 1550
rect 12540 1530 12545 1550
rect 12515 1520 12545 1530
rect 12570 1650 12600 1660
rect 12570 1630 12575 1650
rect 12595 1630 12600 1650
rect 12570 1600 12600 1630
rect 12570 1580 12575 1600
rect 12595 1580 12600 1600
rect 12570 1550 12600 1580
rect 12570 1530 12575 1550
rect 12595 1530 12600 1550
rect 12570 1520 12600 1530
rect 12625 1650 12655 1660
rect 12625 1630 12630 1650
rect 12650 1630 12655 1650
rect 12625 1600 12655 1630
rect 12625 1580 12630 1600
rect 12650 1580 12655 1600
rect 12625 1550 12655 1580
rect 12625 1530 12630 1550
rect 12650 1530 12655 1550
rect 12625 1520 12655 1530
rect 12680 1650 12710 1660
rect 12680 1630 12685 1650
rect 12705 1630 12710 1650
rect 12680 1600 12710 1630
rect 12680 1580 12685 1600
rect 12705 1580 12710 1600
rect 12680 1550 12710 1580
rect 12680 1530 12685 1550
rect 12705 1530 12710 1550
rect 12680 1520 12710 1530
rect 12735 1650 12810 1660
rect 12735 1630 12740 1650
rect 12760 1630 12780 1650
rect 12800 1630 12810 1650
rect 12735 1600 12810 1630
rect 12735 1580 12740 1600
rect 12760 1580 12780 1600
rect 12800 1580 12810 1600
rect 12735 1550 12810 1580
rect 12735 1530 12740 1550
rect 12760 1530 12780 1550
rect 12800 1530 12810 1550
rect 12735 1520 12810 1530
rect 18490 1650 18565 1660
rect 18490 1630 18500 1650
rect 18520 1630 18540 1650
rect 18560 1630 18565 1650
rect 18490 1600 18565 1630
rect 18490 1580 18500 1600
rect 18520 1580 18540 1600
rect 18560 1580 18565 1600
rect 18490 1550 18565 1580
rect 18490 1530 18500 1550
rect 18520 1530 18540 1550
rect 18560 1530 18565 1550
rect 18490 1520 18565 1530
rect 18590 1650 18620 1660
rect 18590 1630 18595 1650
rect 18615 1630 18620 1650
rect 18590 1600 18620 1630
rect 18590 1580 18595 1600
rect 18615 1580 18620 1600
rect 18590 1550 18620 1580
rect 18590 1530 18595 1550
rect 18615 1530 18620 1550
rect 18590 1520 18620 1530
rect 18645 1650 18675 1660
rect 18645 1630 18650 1650
rect 18670 1630 18675 1650
rect 18645 1600 18675 1630
rect 18645 1580 18650 1600
rect 18670 1580 18675 1600
rect 18645 1550 18675 1580
rect 18645 1530 18650 1550
rect 18670 1530 18675 1550
rect 18645 1520 18675 1530
rect 18700 1650 18730 1660
rect 18700 1630 18705 1650
rect 18725 1630 18730 1650
rect 18700 1600 18730 1630
rect 18700 1580 18705 1600
rect 18725 1580 18730 1600
rect 18700 1550 18730 1580
rect 18700 1530 18705 1550
rect 18725 1530 18730 1550
rect 18700 1520 18730 1530
rect 18755 1650 18785 1660
rect 18755 1630 18760 1650
rect 18780 1630 18785 1650
rect 18755 1600 18785 1630
rect 18755 1580 18760 1600
rect 18780 1580 18785 1600
rect 18755 1550 18785 1580
rect 18755 1530 18760 1550
rect 18780 1530 18785 1550
rect 18755 1520 18785 1530
rect 18810 1650 18840 1660
rect 18810 1630 18815 1650
rect 18835 1630 18840 1650
rect 18810 1600 18840 1630
rect 18810 1580 18815 1600
rect 18835 1580 18840 1600
rect 18810 1550 18840 1580
rect 18810 1530 18815 1550
rect 18835 1530 18840 1550
rect 18810 1520 18840 1530
rect 18865 1650 18895 1660
rect 18865 1630 18870 1650
rect 18890 1630 18895 1650
rect 18865 1600 18895 1630
rect 18865 1580 18870 1600
rect 18890 1580 18895 1600
rect 18865 1550 18895 1580
rect 18865 1530 18870 1550
rect 18890 1530 18895 1550
rect 18865 1520 18895 1530
rect 18920 1650 18950 1660
rect 18920 1630 18925 1650
rect 18945 1630 18950 1650
rect 18920 1600 18950 1630
rect 18920 1580 18925 1600
rect 18945 1580 18950 1600
rect 18920 1550 18950 1580
rect 18920 1530 18925 1550
rect 18945 1530 18950 1550
rect 18920 1520 18950 1530
rect 18975 1650 19005 1660
rect 18975 1630 18980 1650
rect 19000 1630 19005 1650
rect 18975 1600 19005 1630
rect 18975 1580 18980 1600
rect 19000 1580 19005 1600
rect 18975 1550 19005 1580
rect 18975 1530 18980 1550
rect 19000 1530 19005 1550
rect 18975 1520 19005 1530
rect 19030 1650 19060 1660
rect 19030 1630 19035 1650
rect 19055 1630 19060 1650
rect 19030 1600 19060 1630
rect 19030 1580 19035 1600
rect 19055 1580 19060 1600
rect 19030 1550 19060 1580
rect 19030 1530 19035 1550
rect 19055 1530 19060 1550
rect 19030 1520 19060 1530
rect 19085 1650 19115 1660
rect 19085 1630 19090 1650
rect 19110 1630 19115 1650
rect 19085 1600 19115 1630
rect 19085 1580 19090 1600
rect 19110 1580 19115 1600
rect 19085 1550 19115 1580
rect 19085 1530 19090 1550
rect 19110 1530 19115 1550
rect 19085 1520 19115 1530
rect 19140 1650 19170 1660
rect 19140 1630 19145 1650
rect 19165 1630 19170 1650
rect 19140 1600 19170 1630
rect 19140 1580 19145 1600
rect 19165 1580 19170 1600
rect 19140 1550 19170 1580
rect 19140 1530 19145 1550
rect 19165 1530 19170 1550
rect 19140 1520 19170 1530
rect 19195 1650 19305 1660
rect 19195 1630 19200 1650
rect 19220 1630 19240 1650
rect 19260 1630 19280 1650
rect 19300 1630 19305 1650
rect 19195 1600 19305 1630
rect 19195 1580 19200 1600
rect 19220 1580 19240 1600
rect 19260 1580 19280 1600
rect 19300 1580 19305 1600
rect 19195 1550 19305 1580
rect 19195 1530 19200 1550
rect 19220 1530 19240 1550
rect 19260 1530 19280 1550
rect 19300 1530 19305 1550
rect 19195 1520 19305 1530
rect 19330 1650 19360 1660
rect 19330 1630 19335 1650
rect 19355 1630 19360 1650
rect 19330 1600 19360 1630
rect 19330 1580 19335 1600
rect 19355 1580 19360 1600
rect 19330 1550 19360 1580
rect 19330 1530 19335 1550
rect 19355 1530 19360 1550
rect 19330 1520 19360 1530
rect 19385 1650 19415 1660
rect 19385 1630 19390 1650
rect 19410 1630 19415 1650
rect 19385 1600 19415 1630
rect 19385 1580 19390 1600
rect 19410 1580 19415 1600
rect 19385 1550 19415 1580
rect 19385 1530 19390 1550
rect 19410 1530 19415 1550
rect 19385 1520 19415 1530
rect 19440 1650 19470 1660
rect 19440 1630 19445 1650
rect 19465 1630 19470 1650
rect 19440 1600 19470 1630
rect 19440 1580 19445 1600
rect 19465 1580 19470 1600
rect 19440 1550 19470 1580
rect 19440 1530 19445 1550
rect 19465 1530 19470 1550
rect 19440 1520 19470 1530
rect 19495 1650 19605 1660
rect 19495 1630 19500 1650
rect 19520 1630 19540 1650
rect 19560 1630 19580 1650
rect 19600 1630 19605 1650
rect 19495 1600 19605 1630
rect 19495 1580 19500 1600
rect 19520 1580 19540 1600
rect 19560 1580 19580 1600
rect 19600 1580 19605 1600
rect 19495 1550 19605 1580
rect 19495 1530 19500 1550
rect 19520 1530 19540 1550
rect 19560 1530 19580 1550
rect 19600 1530 19605 1550
rect 19495 1520 19605 1530
rect 19630 1650 19660 1660
rect 19630 1630 19635 1650
rect 19655 1630 19660 1650
rect 19630 1600 19660 1630
rect 19630 1580 19635 1600
rect 19655 1580 19660 1600
rect 19630 1550 19660 1580
rect 19630 1530 19635 1550
rect 19655 1530 19660 1550
rect 19630 1520 19660 1530
rect 19685 1650 19715 1660
rect 19685 1630 19690 1650
rect 19710 1630 19715 1650
rect 19685 1600 19715 1630
rect 19685 1580 19690 1600
rect 19710 1580 19715 1600
rect 19685 1550 19715 1580
rect 19685 1530 19690 1550
rect 19710 1530 19715 1550
rect 19685 1520 19715 1530
rect 19740 1650 19770 1660
rect 19740 1630 19745 1650
rect 19765 1630 19770 1650
rect 19740 1600 19770 1630
rect 19740 1580 19745 1600
rect 19765 1580 19770 1600
rect 19740 1550 19770 1580
rect 19740 1530 19745 1550
rect 19765 1530 19770 1550
rect 19740 1520 19770 1530
rect 19795 1650 19825 1660
rect 19795 1630 19800 1650
rect 19820 1630 19825 1650
rect 19795 1600 19825 1630
rect 19795 1580 19800 1600
rect 19820 1580 19825 1600
rect 19795 1550 19825 1580
rect 19795 1530 19800 1550
rect 19820 1530 19825 1550
rect 19795 1520 19825 1530
rect 19850 1650 19880 1660
rect 19850 1630 19855 1650
rect 19875 1630 19880 1650
rect 19850 1600 19880 1630
rect 19850 1580 19855 1600
rect 19875 1580 19880 1600
rect 19850 1550 19880 1580
rect 19850 1530 19855 1550
rect 19875 1530 19880 1550
rect 19850 1520 19880 1530
rect 19905 1650 19935 1660
rect 19905 1630 19910 1650
rect 19930 1630 19935 1650
rect 19905 1600 19935 1630
rect 19905 1580 19910 1600
rect 19930 1580 19935 1600
rect 19905 1550 19935 1580
rect 19905 1530 19910 1550
rect 19930 1530 19935 1550
rect 19905 1520 19935 1530
rect 19960 1650 19990 1660
rect 19960 1630 19965 1650
rect 19985 1630 19990 1650
rect 19960 1600 19990 1630
rect 19960 1580 19965 1600
rect 19985 1580 19990 1600
rect 19960 1550 19990 1580
rect 19960 1530 19965 1550
rect 19985 1530 19990 1550
rect 19960 1520 19990 1530
rect 20015 1650 20045 1660
rect 20015 1630 20020 1650
rect 20040 1630 20045 1650
rect 20015 1600 20045 1630
rect 20015 1580 20020 1600
rect 20040 1580 20045 1600
rect 20015 1550 20045 1580
rect 20015 1530 20020 1550
rect 20040 1530 20045 1550
rect 20015 1520 20045 1530
rect 20070 1650 20100 1660
rect 20070 1630 20075 1650
rect 20095 1630 20100 1650
rect 20070 1600 20100 1630
rect 20070 1580 20075 1600
rect 20095 1580 20100 1600
rect 20070 1550 20100 1580
rect 20070 1530 20075 1550
rect 20095 1530 20100 1550
rect 20070 1520 20100 1530
rect 20125 1650 20155 1660
rect 20125 1630 20130 1650
rect 20150 1630 20155 1650
rect 20125 1600 20155 1630
rect 20125 1580 20130 1600
rect 20150 1580 20155 1600
rect 20125 1550 20155 1580
rect 20125 1530 20130 1550
rect 20150 1530 20155 1550
rect 20125 1520 20155 1530
rect 20180 1650 20210 1660
rect 20180 1630 20185 1650
rect 20205 1630 20210 1650
rect 20180 1600 20210 1630
rect 20180 1580 20185 1600
rect 20205 1580 20210 1600
rect 20180 1550 20210 1580
rect 20180 1530 20185 1550
rect 20205 1530 20210 1550
rect 20180 1520 20210 1530
rect 20235 1650 20310 1660
rect 20235 1630 20240 1650
rect 20260 1630 20280 1650
rect 20300 1630 20310 1650
rect 20566 1655 20571 1675
rect 20591 1655 20598 1675
rect 20566 1645 20598 1655
rect 20615 1680 20655 1690
rect 20615 1660 20625 1680
rect 20645 1660 20655 1680
rect 20615 1650 20655 1660
rect 20710 1680 20750 1690
rect 20710 1660 20720 1680
rect 20740 1660 20750 1680
rect 20710 1650 20750 1660
rect 20235 1600 20310 1630
rect 20235 1580 20240 1600
rect 20260 1580 20280 1600
rect 20300 1580 20310 1600
rect 20510 1625 20550 1635
rect 20510 1605 20520 1625
rect 20540 1605 20550 1625
rect 20510 1595 20550 1605
rect 20800 1625 20840 1635
rect 20800 1605 20810 1625
rect 20830 1605 20840 1625
rect 20800 1595 20840 1605
rect 20235 1550 20310 1580
rect 20235 1530 20240 1550
rect 20260 1530 20280 1550
rect 20300 1530 20310 1550
rect 20471 1565 20503 1575
rect 20471 1545 20476 1565
rect 20496 1545 20503 1565
rect 20471 1535 20503 1545
rect 20235 1520 20310 1530
rect 4745 1510 4785 1520
rect 2925 1495 2965 1505
rect 2835 1480 2875 1490
rect 2835 1460 2845 1480
rect 2865 1460 2875 1480
rect 2925 1475 2935 1495
rect 2955 1475 2965 1495
rect 2925 1465 2965 1475
rect 3045 1495 3085 1505
rect 3045 1475 3055 1495
rect 3075 1475 3085 1495
rect 3045 1465 3085 1475
rect 3165 1495 3205 1505
rect 3165 1475 3175 1495
rect 3195 1475 3205 1495
rect 3165 1465 3205 1475
rect 3285 1495 3325 1505
rect 3285 1475 3295 1495
rect 3315 1475 3325 1495
rect 3285 1465 3325 1475
rect 3525 1495 3565 1505
rect 3525 1475 3535 1495
rect 3555 1475 3565 1495
rect 3525 1465 3565 1475
rect 3645 1495 3685 1505
rect 3645 1475 3655 1495
rect 3675 1475 3685 1495
rect 3645 1465 3685 1475
rect 3765 1495 3805 1505
rect 3765 1475 3775 1495
rect 3795 1475 3805 1495
rect 4205 1495 4245 1505
rect 3765 1465 3805 1475
rect 3915 1480 3955 1490
rect 2835 1450 2875 1460
rect 3915 1460 3925 1480
rect 3945 1460 3955 1480
rect 3915 1450 3955 1460
rect 4055 1480 4095 1490
rect 4055 1460 4065 1480
rect 4085 1460 4095 1480
rect 4205 1475 4215 1495
rect 4235 1475 4245 1495
rect 4205 1465 4245 1475
rect 4325 1495 4365 1505
rect 4325 1475 4335 1495
rect 4355 1475 4365 1495
rect 4325 1465 4365 1475
rect 4445 1495 4485 1505
rect 4445 1475 4455 1495
rect 4475 1475 4485 1495
rect 4445 1465 4485 1475
rect 4685 1495 4725 1505
rect 4685 1475 4695 1495
rect 4715 1475 4725 1495
rect 4685 1465 4725 1475
rect 4805 1495 4845 1505
rect 4805 1475 4815 1495
rect 4835 1475 4845 1495
rect 4805 1465 4845 1475
rect 4925 1495 4965 1505
rect 4925 1475 4935 1495
rect 4955 1475 4965 1495
rect 4925 1465 4965 1475
rect 5045 1495 5085 1505
rect 11000 1500 11020 1520
rect 5045 1475 5055 1495
rect 5075 1475 5085 1495
rect 10990 1490 11030 1500
rect 5045 1465 5085 1475
rect 5135 1480 5175 1490
rect 4055 1450 4095 1460
rect 5135 1460 5145 1480
rect 5165 1460 5175 1480
rect 10990 1470 11000 1490
rect 11020 1470 11030 1490
rect 10990 1460 11030 1470
rect 11106 1490 11138 1500
rect 11106 1470 11112 1490
rect 11129 1470 11138 1490
rect 11106 1460 11138 1470
rect 5135 1450 5175 1460
rect 125 1335 2135 1375
rect 650 690 775 1335
rect 1330 690 1455 1335
rect 2010 695 2135 1335
rect 2840 1440 2870 1450
rect 2840 1420 2845 1440
rect 2865 1420 2870 1440
rect 2840 1390 2870 1420
rect 2840 1370 2845 1390
rect 2865 1370 2870 1390
rect 2840 1340 2870 1370
rect 2840 1320 2845 1340
rect 2865 1320 2870 1340
rect 2840 1290 2870 1320
rect 2840 1270 2845 1290
rect 2865 1270 2870 1290
rect 2840 1240 2870 1270
rect 2840 1220 2845 1240
rect 2865 1220 2870 1240
rect 2840 1210 2870 1220
rect 3380 1440 3410 1450
rect 3380 1420 3385 1440
rect 3405 1420 3410 1440
rect 3380 1390 3410 1420
rect 3380 1370 3385 1390
rect 3405 1370 3410 1390
rect 3380 1340 3410 1370
rect 3380 1320 3385 1340
rect 3405 1320 3410 1340
rect 3380 1290 3410 1320
rect 3380 1270 3385 1290
rect 3405 1270 3410 1290
rect 3380 1240 3410 1270
rect 3380 1220 3385 1240
rect 3405 1220 3410 1240
rect 3380 1210 3410 1220
rect 3920 1440 3950 1450
rect 3920 1420 3925 1440
rect 3945 1420 3950 1440
rect 3920 1390 3950 1420
rect 3920 1370 3925 1390
rect 3945 1370 3950 1390
rect 3920 1340 3950 1370
rect 3920 1320 3925 1340
rect 3945 1320 3950 1340
rect 3920 1290 3950 1320
rect 3920 1270 3925 1290
rect 3945 1270 3950 1290
rect 3920 1240 3950 1270
rect 3920 1220 3925 1240
rect 3945 1220 3950 1240
rect 3920 1210 3950 1220
rect 4060 1440 4090 1450
rect 4060 1420 4065 1440
rect 4085 1420 4090 1440
rect 4060 1390 4090 1420
rect 4060 1370 4065 1390
rect 4085 1370 4090 1390
rect 4060 1340 4090 1370
rect 4060 1320 4065 1340
rect 4085 1320 4090 1340
rect 4060 1290 4090 1320
rect 4060 1270 4065 1290
rect 4085 1270 4090 1290
rect 4060 1240 4090 1270
rect 4060 1220 4065 1240
rect 4085 1220 4090 1240
rect 4060 1210 4090 1220
rect 4600 1440 4630 1450
rect 4600 1420 4605 1440
rect 4625 1420 4630 1440
rect 4600 1390 4630 1420
rect 4600 1370 4605 1390
rect 4625 1370 4630 1390
rect 4600 1340 4630 1370
rect 4600 1320 4605 1340
rect 4625 1320 4630 1340
rect 4600 1290 4630 1320
rect 4600 1270 4605 1290
rect 4625 1270 4630 1290
rect 4600 1240 4630 1270
rect 4600 1220 4605 1240
rect 4625 1220 4630 1240
rect 4600 1210 4630 1220
rect 5140 1440 5170 1450
rect 11155 1440 11175 1520
rect 11260 1440 11280 1520
rect 11305 1490 11345 1500
rect 11305 1470 11315 1490
rect 11335 1470 11345 1490
rect 11305 1460 11345 1470
rect 11370 1440 11390 1520
rect 11480 1440 11500 1520
rect 11525 1490 11565 1500
rect 11525 1470 11535 1490
rect 11555 1470 11565 1490
rect 11525 1460 11565 1470
rect 11590 1440 11610 1520
rect 11740 1500 11760 1520
rect 11830 1500 11850 1520
rect 11885 1500 11905 1520
rect 12040 1500 12060 1520
rect 11730 1490 11770 1500
rect 11730 1470 11740 1490
rect 11760 1470 11770 1490
rect 11730 1460 11770 1470
rect 11825 1490 11855 1500
rect 11825 1470 11830 1490
rect 11850 1470 11855 1490
rect 11825 1460 11855 1470
rect 11875 1490 11905 1500
rect 11875 1470 11880 1490
rect 11900 1470 11905 1490
rect 11875 1460 11905 1470
rect 11922 1490 11954 1500
rect 11922 1470 11928 1490
rect 11945 1470 11954 1490
rect 11922 1460 11954 1470
rect 12030 1490 12070 1500
rect 12030 1470 12040 1490
rect 12060 1470 12070 1490
rect 12030 1460 12070 1470
rect 12146 1490 12178 1500
rect 12146 1470 12152 1490
rect 12169 1470 12178 1490
rect 12146 1460 12178 1470
rect 12195 1440 12215 1520
rect 12300 1440 12320 1520
rect 12345 1490 12385 1500
rect 12345 1470 12355 1490
rect 12375 1470 12385 1490
rect 12345 1460 12385 1470
rect 12410 1440 12430 1520
rect 12520 1440 12540 1520
rect 12565 1490 12605 1500
rect 12565 1470 12575 1490
rect 12595 1470 12605 1490
rect 12565 1460 12605 1470
rect 12630 1440 12650 1520
rect 12780 1500 12800 1520
rect 18500 1500 18520 1520
rect 12770 1490 12810 1500
rect 12770 1470 12780 1490
rect 12800 1470 12810 1490
rect 12770 1460 12810 1470
rect 18490 1490 18530 1500
rect 18490 1470 18500 1490
rect 18520 1470 18530 1490
rect 18490 1460 18530 1470
rect 18606 1490 18638 1500
rect 18606 1470 18612 1490
rect 18629 1470 18638 1490
rect 18606 1460 18638 1470
rect 18655 1440 18675 1520
rect 18760 1440 18780 1520
rect 18805 1490 18845 1500
rect 18805 1470 18815 1490
rect 18835 1470 18845 1490
rect 18805 1460 18845 1470
rect 18870 1440 18890 1520
rect 18980 1440 19000 1520
rect 19025 1490 19065 1500
rect 19025 1470 19035 1490
rect 19055 1470 19065 1490
rect 19025 1460 19065 1470
rect 19090 1440 19110 1520
rect 19240 1500 19260 1520
rect 19330 1500 19350 1520
rect 19385 1500 19405 1520
rect 19540 1500 19560 1520
rect 19230 1490 19270 1500
rect 19230 1470 19240 1490
rect 19260 1470 19270 1490
rect 19230 1460 19270 1470
rect 19325 1490 19355 1500
rect 19325 1470 19330 1490
rect 19350 1470 19355 1490
rect 19325 1460 19355 1470
rect 19375 1490 19405 1500
rect 19375 1470 19380 1490
rect 19400 1470 19405 1490
rect 19375 1460 19405 1470
rect 19422 1490 19454 1500
rect 19422 1470 19428 1490
rect 19445 1470 19454 1490
rect 19422 1460 19454 1470
rect 19530 1490 19570 1500
rect 19530 1470 19540 1490
rect 19560 1470 19570 1490
rect 19530 1460 19570 1470
rect 19646 1490 19678 1500
rect 19646 1470 19652 1490
rect 19669 1470 19678 1490
rect 19646 1460 19678 1470
rect 19695 1440 19715 1520
rect 19800 1440 19820 1520
rect 19845 1490 19885 1500
rect 19845 1470 19855 1490
rect 19875 1470 19885 1490
rect 19845 1460 19885 1470
rect 19910 1440 19930 1520
rect 20020 1440 20040 1520
rect 20065 1490 20105 1500
rect 20065 1470 20075 1490
rect 20095 1470 20105 1490
rect 20065 1460 20105 1470
rect 20130 1440 20150 1520
rect 20280 1500 20300 1520
rect 20520 1515 20540 1595
rect 20560 1565 20600 1575
rect 20560 1545 20570 1565
rect 20590 1545 20600 1565
rect 20560 1535 20600 1545
rect 20570 1515 20590 1535
rect 20810 1515 20830 1595
rect 20847 1565 20879 1575
rect 20847 1545 20854 1565
rect 20874 1545 20879 1565
rect 20847 1535 20879 1545
rect 20355 1505 20430 1515
rect 20270 1490 20310 1500
rect 20270 1470 20280 1490
rect 20300 1470 20310 1490
rect 20270 1460 20310 1470
rect 20355 1485 20365 1505
rect 20385 1485 20405 1505
rect 20425 1485 20430 1505
rect 20355 1455 20430 1485
rect 5140 1420 5145 1440
rect 5165 1420 5170 1440
rect 5140 1390 5170 1420
rect 11145 1430 11185 1440
rect 11145 1410 11155 1430
rect 11175 1410 11185 1430
rect 11145 1400 11185 1410
rect 11250 1430 11290 1440
rect 11250 1410 11260 1430
rect 11280 1410 11290 1430
rect 11250 1400 11290 1410
rect 11360 1430 11400 1440
rect 11360 1410 11370 1430
rect 11390 1410 11400 1430
rect 11360 1400 11400 1410
rect 11470 1430 11510 1440
rect 11470 1410 11480 1430
rect 11500 1410 11510 1430
rect 11470 1400 11510 1410
rect 11580 1430 11620 1440
rect 11580 1410 11590 1430
rect 11610 1410 11620 1430
rect 11580 1400 11620 1410
rect 12185 1430 12225 1440
rect 12185 1410 12195 1430
rect 12215 1410 12225 1430
rect 12185 1400 12225 1410
rect 12290 1430 12330 1440
rect 12290 1410 12300 1430
rect 12320 1410 12330 1430
rect 12290 1400 12330 1410
rect 12400 1430 12440 1440
rect 12400 1410 12410 1430
rect 12430 1410 12440 1430
rect 12400 1400 12440 1410
rect 12510 1430 12550 1440
rect 12510 1410 12520 1430
rect 12540 1410 12550 1430
rect 12510 1400 12550 1410
rect 12620 1430 12660 1440
rect 18645 1430 18685 1440
rect 12620 1410 12630 1430
rect 12650 1410 12660 1430
rect 12620 1400 12660 1410
rect 13015 1425 13060 1430
rect 13015 1400 13025 1425
rect 13050 1400 13060 1425
rect 13015 1395 13060 1400
rect 14025 1425 14070 1430
rect 14025 1400 14035 1425
rect 14060 1400 14070 1425
rect 18645 1410 18655 1430
rect 18675 1410 18685 1430
rect 18645 1400 18685 1410
rect 18750 1430 18790 1440
rect 18750 1410 18760 1430
rect 18780 1410 18790 1430
rect 18750 1400 18790 1410
rect 18860 1430 18900 1440
rect 18860 1410 18870 1430
rect 18890 1410 18900 1430
rect 18860 1400 18900 1410
rect 18970 1430 19010 1440
rect 18970 1410 18980 1430
rect 19000 1410 19010 1430
rect 18970 1400 19010 1410
rect 19080 1430 19120 1440
rect 19080 1410 19090 1430
rect 19110 1410 19120 1430
rect 19080 1400 19120 1410
rect 19685 1430 19725 1440
rect 19685 1410 19695 1430
rect 19715 1410 19725 1430
rect 19685 1400 19725 1410
rect 19790 1430 19830 1440
rect 19790 1410 19800 1430
rect 19820 1410 19830 1430
rect 19790 1400 19830 1410
rect 19900 1430 19940 1440
rect 19900 1410 19910 1430
rect 19930 1410 19940 1430
rect 19900 1400 19940 1410
rect 20010 1430 20050 1440
rect 20010 1410 20020 1430
rect 20040 1410 20050 1430
rect 20010 1400 20050 1410
rect 20120 1430 20160 1440
rect 20120 1410 20130 1430
rect 20150 1410 20160 1430
rect 20120 1400 20160 1410
rect 20355 1435 20365 1455
rect 20385 1435 20405 1455
rect 20425 1435 20430 1455
rect 20355 1405 20430 1435
rect 14025 1395 14070 1400
rect 5140 1370 5145 1390
rect 5165 1370 5170 1390
rect 5140 1340 5170 1370
rect 19310 1350 19350 1390
rect 20355 1385 20365 1405
rect 20385 1385 20405 1405
rect 20425 1385 20430 1405
rect 20355 1375 20430 1385
rect 20455 1505 20485 1515
rect 20455 1485 20460 1505
rect 20480 1485 20485 1505
rect 20455 1455 20485 1485
rect 20455 1435 20460 1455
rect 20480 1435 20485 1455
rect 20455 1405 20485 1435
rect 20455 1385 20460 1405
rect 20480 1385 20485 1405
rect 20455 1375 20485 1385
rect 20510 1505 20540 1515
rect 20510 1485 20515 1505
rect 20535 1485 20540 1505
rect 20510 1455 20540 1485
rect 20510 1435 20515 1455
rect 20535 1435 20540 1455
rect 20510 1405 20540 1435
rect 20510 1385 20515 1405
rect 20535 1385 20540 1405
rect 20510 1375 20540 1385
rect 20565 1505 20595 1515
rect 20565 1485 20570 1505
rect 20590 1485 20595 1505
rect 20565 1455 20595 1485
rect 20565 1435 20570 1455
rect 20590 1435 20595 1455
rect 20565 1405 20595 1435
rect 20565 1385 20570 1405
rect 20590 1385 20595 1405
rect 20565 1375 20595 1385
rect 20620 1505 20730 1515
rect 20620 1485 20625 1505
rect 20645 1485 20665 1505
rect 20685 1485 20705 1505
rect 20725 1485 20730 1505
rect 20620 1455 20730 1485
rect 20620 1435 20625 1455
rect 20645 1435 20665 1455
rect 20685 1435 20705 1455
rect 20725 1435 20730 1455
rect 20620 1405 20730 1435
rect 20620 1385 20625 1405
rect 20645 1385 20665 1405
rect 20685 1385 20705 1405
rect 20725 1385 20730 1405
rect 20620 1375 20730 1385
rect 20755 1505 20785 1515
rect 20755 1485 20760 1505
rect 20780 1485 20785 1505
rect 20755 1455 20785 1485
rect 20755 1435 20760 1455
rect 20780 1435 20785 1455
rect 20755 1405 20785 1435
rect 20755 1385 20760 1405
rect 20780 1385 20785 1405
rect 20755 1375 20785 1385
rect 20810 1505 20840 1515
rect 20810 1485 20815 1505
rect 20835 1485 20840 1505
rect 20810 1455 20840 1485
rect 20810 1435 20815 1455
rect 20835 1435 20840 1455
rect 20810 1405 20840 1435
rect 20810 1385 20815 1405
rect 20835 1385 20840 1405
rect 20810 1375 20840 1385
rect 20865 1505 20895 1515
rect 20865 1485 20870 1505
rect 20890 1485 20895 1505
rect 20865 1455 20895 1485
rect 20865 1435 20870 1455
rect 20890 1435 20895 1455
rect 20865 1405 20895 1435
rect 20865 1385 20870 1405
rect 20890 1385 20895 1405
rect 20865 1375 20895 1385
rect 20920 1505 20995 1515
rect 20920 1485 20925 1505
rect 20945 1485 20965 1505
rect 20985 1485 20995 1505
rect 20920 1455 20995 1485
rect 20920 1435 20925 1455
rect 20945 1435 20965 1455
rect 20985 1435 20995 1455
rect 20920 1405 20995 1435
rect 20920 1385 20925 1405
rect 20945 1385 20965 1405
rect 20985 1385 20995 1405
rect 20920 1375 20995 1385
rect 20365 1355 20385 1375
rect 20355 1345 20395 1355
rect 5140 1320 5145 1340
rect 5165 1320 5170 1340
rect 5140 1290 5170 1320
rect 11810 1300 11850 1340
rect 13025 1315 13065 1325
rect 13025 1295 13035 1315
rect 13055 1295 13065 1315
rect 5140 1270 5145 1290
rect 5165 1270 5170 1290
rect 5140 1240 5170 1270
rect 11315 1250 11355 1290
rect 11880 1250 11920 1290
rect 13025 1285 13065 1295
rect 13128 1315 13162 1325
rect 13128 1295 13136 1315
rect 13154 1295 13162 1315
rect 13128 1285 13162 1295
rect 13225 1315 13265 1325
rect 13225 1295 13235 1315
rect 13255 1295 13265 1315
rect 13225 1285 13265 1295
rect 13425 1315 13465 1325
rect 13425 1295 13435 1315
rect 13455 1295 13465 1315
rect 13425 1285 13465 1295
rect 13625 1315 13665 1325
rect 13625 1295 13635 1315
rect 13655 1295 13665 1315
rect 13625 1285 13665 1295
rect 13825 1315 13865 1325
rect 13825 1295 13835 1315
rect 13855 1295 13865 1315
rect 13825 1285 13865 1295
rect 14025 1315 14065 1325
rect 14025 1295 14035 1315
rect 14055 1295 14065 1315
rect 18815 1300 18855 1340
rect 19380 1300 19420 1340
rect 20355 1325 20365 1345
rect 20385 1325 20395 1345
rect 20355 1315 20395 1325
rect 20455 1295 20475 1375
rect 20526 1345 20558 1355
rect 20526 1325 20533 1345
rect 20553 1325 20558 1345
rect 20526 1315 20558 1325
rect 20575 1295 20595 1375
rect 20665 1355 20685 1375
rect 20655 1345 20695 1355
rect 20655 1325 20665 1345
rect 20685 1325 20695 1345
rect 20655 1315 20695 1325
rect 20755 1295 20775 1375
rect 20792 1345 20824 1355
rect 20792 1325 20797 1345
rect 20817 1325 20824 1345
rect 20792 1315 20824 1325
rect 20875 1295 20895 1375
rect 20965 1355 20985 1375
rect 20955 1345 20995 1355
rect 20955 1325 20965 1345
rect 20985 1325 20995 1345
rect 20955 1315 20995 1325
rect 14025 1285 14065 1295
rect 20095 1285 20135 1295
rect 13035 1265 13055 1285
rect 13235 1265 13255 1285
rect 13435 1265 13455 1285
rect 13635 1265 13655 1285
rect 13835 1265 13855 1285
rect 14035 1265 14055 1285
rect 18815 1270 18855 1280
rect 12890 1255 12960 1265
rect 5140 1220 5145 1240
rect 5165 1220 5170 1240
rect 12595 1235 12635 1245
rect 5140 1210 5170 1220
rect 11315 1220 11355 1230
rect 3385 1190 3405 1210
rect 4605 1190 4625 1210
rect 11315 1200 11325 1220
rect 11345 1200 11355 1220
rect 11315 1190 11355 1200
rect 11425 1220 11465 1230
rect 11425 1200 11435 1220
rect 11455 1200 11465 1220
rect 11425 1190 11465 1200
rect 11535 1220 11575 1230
rect 11535 1200 11545 1220
rect 11565 1200 11575 1220
rect 11535 1190 11575 1200
rect 11645 1220 11685 1230
rect 11645 1200 11655 1220
rect 11675 1200 11685 1220
rect 11645 1190 11685 1200
rect 11755 1220 11795 1230
rect 11755 1200 11765 1220
rect 11785 1200 11795 1220
rect 11755 1190 11795 1200
rect 11815 1220 11845 1230
rect 11815 1200 11820 1220
rect 11840 1200 11845 1220
rect 11815 1190 11845 1200
rect 11865 1220 11905 1230
rect 11865 1200 11875 1220
rect 11895 1200 11905 1220
rect 11865 1190 11905 1200
rect 11975 1220 12015 1230
rect 11975 1200 11985 1220
rect 12005 1200 12015 1220
rect 11975 1190 12015 1200
rect 12085 1220 12125 1230
rect 12085 1200 12095 1220
rect 12115 1200 12125 1220
rect 12085 1190 12125 1200
rect 12195 1220 12235 1230
rect 12195 1200 12205 1220
rect 12225 1200 12235 1220
rect 12195 1190 12235 1200
rect 12305 1220 12345 1230
rect 12305 1200 12315 1220
rect 12335 1200 12345 1220
rect 12305 1190 12345 1200
rect 12415 1220 12455 1230
rect 12415 1200 12425 1220
rect 12445 1200 12455 1220
rect 12415 1190 12455 1200
rect 12525 1220 12565 1230
rect 12525 1200 12535 1220
rect 12555 1200 12565 1220
rect 12595 1215 12605 1235
rect 12625 1215 12635 1235
rect 12595 1205 12635 1215
rect 12890 1235 12895 1255
rect 12915 1235 12935 1255
rect 12955 1235 12960 1255
rect 12890 1210 12960 1235
rect 12525 1190 12565 1200
rect 12890 1190 12895 1210
rect 12915 1190 12935 1210
rect 12955 1190 12960 1210
rect 3375 1180 3415 1190
rect 3375 1160 3385 1180
rect 3405 1160 3415 1180
rect 3375 1150 3415 1160
rect 3990 1155 4020 1185
rect 4595 1180 4635 1190
rect 4595 1160 4605 1180
rect 4625 1160 4635 1180
rect 11325 1170 11345 1190
rect 11435 1170 11455 1190
rect 11545 1170 11565 1190
rect 11655 1170 11675 1190
rect 11765 1170 11785 1190
rect 11875 1170 11895 1190
rect 11985 1170 12005 1190
rect 12095 1170 12115 1190
rect 12205 1170 12225 1190
rect 12315 1170 12335 1190
rect 12425 1170 12445 1190
rect 12535 1170 12555 1190
rect 4595 1150 4635 1160
rect 11170 1160 11240 1170
rect 11170 1140 11175 1160
rect 11195 1140 11215 1160
rect 11235 1140 11240 1160
rect 2945 1120 2985 1130
rect 2945 1100 2955 1120
rect 2975 1100 2985 1120
rect 2945 1090 2985 1100
rect 3025 1120 3065 1130
rect 3025 1100 3035 1120
rect 3055 1100 3065 1120
rect 3025 1090 3065 1100
rect 3105 1120 3145 1130
rect 3105 1100 3115 1120
rect 3135 1100 3145 1120
rect 3105 1090 3145 1100
rect 3185 1120 3225 1130
rect 3185 1100 3195 1120
rect 3215 1100 3225 1120
rect 3185 1090 3225 1100
rect 3265 1120 3305 1130
rect 3265 1100 3275 1120
rect 3295 1100 3305 1120
rect 3265 1090 3305 1100
rect 3345 1120 3385 1130
rect 3345 1100 3355 1120
rect 3375 1100 3385 1120
rect 3345 1090 3385 1100
rect 3425 1120 3465 1130
rect 3425 1100 3435 1120
rect 3455 1100 3465 1120
rect 3425 1090 3465 1100
rect 3505 1120 3545 1130
rect 3505 1100 3515 1120
rect 3535 1100 3545 1120
rect 3505 1090 3545 1100
rect 3585 1120 3625 1130
rect 3585 1100 3595 1120
rect 3615 1100 3625 1120
rect 3585 1090 3625 1100
rect 3665 1120 3705 1130
rect 3665 1100 3675 1120
rect 3695 1100 3705 1120
rect 3665 1090 3705 1100
rect 3745 1120 3785 1130
rect 3745 1100 3755 1120
rect 3775 1100 3785 1120
rect 3745 1090 3785 1100
rect 3825 1120 3865 1130
rect 3825 1100 3835 1120
rect 3855 1100 3865 1120
rect 3825 1090 3865 1100
rect 3905 1120 3945 1130
rect 3905 1100 3915 1120
rect 3935 1100 3945 1120
rect 3905 1090 3945 1100
rect 3985 1120 4025 1130
rect 3985 1100 3995 1120
rect 4015 1100 4025 1120
rect 3985 1090 4025 1100
rect 4065 1120 4105 1130
rect 4065 1100 4075 1120
rect 4095 1100 4105 1120
rect 4065 1090 4105 1100
rect 4145 1120 4185 1130
rect 4145 1100 4155 1120
rect 4175 1100 4185 1120
rect 4145 1090 4185 1100
rect 4225 1120 4265 1130
rect 4225 1100 4235 1120
rect 4255 1100 4265 1120
rect 4225 1090 4265 1100
rect 4305 1120 4345 1130
rect 4305 1100 4315 1120
rect 4335 1100 4345 1120
rect 4305 1090 4345 1100
rect 4385 1120 4425 1130
rect 4385 1100 4395 1120
rect 4415 1100 4425 1120
rect 4385 1090 4425 1100
rect 4465 1120 4505 1130
rect 4465 1100 4475 1120
rect 4495 1100 4505 1120
rect 4465 1090 4505 1100
rect 4545 1120 4585 1130
rect 4545 1100 4555 1120
rect 4575 1100 4585 1120
rect 4545 1090 4585 1100
rect 4625 1120 4665 1130
rect 4625 1100 4635 1120
rect 4655 1100 4665 1120
rect 4625 1090 4665 1100
rect 4705 1120 4745 1130
rect 4705 1100 4715 1120
rect 4735 1100 4745 1120
rect 4705 1090 4745 1100
rect 4785 1120 4825 1130
rect 4785 1100 4795 1120
rect 4815 1100 4825 1120
rect 4785 1090 4825 1100
rect 4865 1120 4905 1130
rect 4865 1100 4875 1120
rect 4895 1100 4905 1120
rect 4865 1090 4905 1100
rect 4945 1120 4985 1130
rect 4945 1100 4955 1120
rect 4975 1100 4985 1120
rect 4945 1090 4985 1100
rect 11170 1110 11240 1140
rect 11170 1090 11175 1110
rect 11195 1090 11215 1110
rect 11235 1090 11240 1110
rect 2955 1070 2975 1090
rect 3995 1070 4015 1090
rect 2950 1060 2980 1070
rect 2950 1045 2955 1060
rect 2935 1040 2955 1045
rect 2975 1040 2980 1060
rect 2625 1010 2655 1040
rect 2910 1035 2980 1040
rect 2910 1015 2915 1035
rect 2935 1015 2980 1035
rect 2910 1010 2980 1015
rect 2935 1005 2955 1010
rect 2950 990 2955 1005
rect 2975 990 2980 1010
rect 2950 980 2980 990
rect 3990 1060 4020 1070
rect 3990 1040 3995 1060
rect 4015 1040 4020 1060
rect 3990 1010 4020 1040
rect 3990 990 3995 1010
rect 4015 990 4020 1010
rect 3990 980 4020 990
rect 5030 1060 5100 1070
rect 5030 1040 5035 1060
rect 5055 1040 5075 1060
rect 5095 1045 5100 1060
rect 11170 1060 11240 1090
rect 5095 1040 5150 1045
rect 5030 1035 5150 1040
rect 5030 1015 5120 1035
rect 5140 1015 5150 1035
rect 5030 1010 5150 1015
rect 5030 990 5035 1010
rect 5055 990 5075 1010
rect 5095 1005 5150 1010
rect 11170 1040 11175 1060
rect 11195 1040 11215 1060
rect 11235 1040 11240 1060
rect 11170 1010 11240 1040
rect 5095 990 5100 1005
rect 5030 980 5100 990
rect 11170 990 11175 1010
rect 11195 990 11215 1010
rect 11235 990 11240 1010
rect 11170 960 11240 990
rect 11170 940 11175 960
rect 11195 940 11215 960
rect 11235 940 11240 960
rect 2995 925 3035 935
rect 2995 905 3005 925
rect 3025 905 3035 925
rect 2995 895 3035 905
rect 3175 925 3215 935
rect 3175 905 3185 925
rect 3205 905 3215 925
rect 3175 895 3215 905
rect 3355 925 3395 935
rect 3355 905 3365 925
rect 3385 905 3395 925
rect 3355 895 3395 905
rect 3535 925 3575 935
rect 3535 905 3545 925
rect 3565 905 3575 925
rect 3535 895 3575 905
rect 3715 925 3755 935
rect 3715 905 3725 925
rect 3745 905 3755 925
rect 3715 895 3755 905
rect 3895 925 3935 935
rect 3895 905 3905 925
rect 3925 905 3935 925
rect 3895 895 3935 905
rect 4075 925 4115 935
rect 4075 905 4085 925
rect 4105 905 4115 925
rect 4075 895 4115 905
rect 4255 925 4295 935
rect 4255 905 4265 925
rect 4285 905 4295 925
rect 4255 895 4295 905
rect 4435 925 4475 935
rect 4435 905 4445 925
rect 4465 905 4475 925
rect 4435 895 4475 905
rect 4615 925 4655 935
rect 4615 905 4625 925
rect 4645 905 4655 925
rect 4615 895 4655 905
rect 4795 925 4835 935
rect 4795 905 4805 925
rect 4825 905 4835 925
rect 4795 895 4835 905
rect 4975 925 5015 935
rect 11170 930 11240 940
rect 11265 1160 11295 1170
rect 11265 1140 11270 1160
rect 11290 1140 11295 1160
rect 11265 1110 11295 1140
rect 11265 1090 11270 1110
rect 11290 1090 11295 1110
rect 11265 1060 11295 1090
rect 11265 1040 11270 1060
rect 11290 1040 11295 1060
rect 11265 1010 11295 1040
rect 11265 990 11270 1010
rect 11290 990 11295 1010
rect 11265 960 11295 990
rect 11265 940 11270 960
rect 11290 940 11295 960
rect 11265 930 11295 940
rect 11320 1160 11350 1170
rect 11320 1140 11325 1160
rect 11345 1140 11350 1160
rect 11320 1110 11350 1140
rect 11320 1090 11325 1110
rect 11345 1090 11350 1110
rect 11320 1060 11350 1090
rect 11320 1040 11325 1060
rect 11345 1040 11350 1060
rect 11320 1010 11350 1040
rect 11320 990 11325 1010
rect 11345 990 11350 1010
rect 11320 960 11350 990
rect 11320 940 11325 960
rect 11345 940 11350 960
rect 11320 930 11350 940
rect 11375 1160 11405 1170
rect 11375 1140 11380 1160
rect 11400 1140 11405 1160
rect 11375 1110 11405 1140
rect 11375 1090 11380 1110
rect 11400 1090 11405 1110
rect 11375 1060 11405 1090
rect 11375 1040 11380 1060
rect 11400 1040 11405 1060
rect 11375 1010 11405 1040
rect 11375 990 11380 1010
rect 11400 990 11405 1010
rect 11375 960 11405 990
rect 11375 940 11380 960
rect 11400 940 11405 960
rect 11375 930 11405 940
rect 11430 1160 11460 1170
rect 11430 1140 11435 1160
rect 11455 1140 11460 1160
rect 11430 1110 11460 1140
rect 11430 1090 11435 1110
rect 11455 1090 11460 1110
rect 11430 1060 11460 1090
rect 11430 1040 11435 1060
rect 11455 1040 11460 1060
rect 11430 1010 11460 1040
rect 11430 990 11435 1010
rect 11455 990 11460 1010
rect 11430 960 11460 990
rect 11430 940 11435 960
rect 11455 940 11460 960
rect 11430 930 11460 940
rect 11485 1160 11515 1170
rect 11485 1140 11490 1160
rect 11510 1140 11515 1160
rect 11485 1110 11515 1140
rect 11485 1090 11490 1110
rect 11510 1090 11515 1110
rect 11485 1060 11515 1090
rect 11485 1040 11490 1060
rect 11510 1040 11515 1060
rect 11485 1010 11515 1040
rect 11485 990 11490 1010
rect 11510 990 11515 1010
rect 11485 960 11515 990
rect 11485 940 11490 960
rect 11510 940 11515 960
rect 11485 930 11515 940
rect 11540 1160 11570 1170
rect 11540 1140 11545 1160
rect 11565 1140 11570 1160
rect 11540 1110 11570 1140
rect 11540 1090 11545 1110
rect 11565 1090 11570 1110
rect 11540 1060 11570 1090
rect 11540 1040 11545 1060
rect 11565 1040 11570 1060
rect 11540 1010 11570 1040
rect 11540 990 11545 1010
rect 11565 990 11570 1010
rect 11540 960 11570 990
rect 11540 940 11545 960
rect 11565 940 11570 960
rect 11540 930 11570 940
rect 11595 1160 11625 1170
rect 11595 1140 11600 1160
rect 11620 1140 11625 1160
rect 11595 1110 11625 1140
rect 11595 1090 11600 1110
rect 11620 1090 11625 1110
rect 11595 1060 11625 1090
rect 11595 1040 11600 1060
rect 11620 1040 11625 1060
rect 11595 1010 11625 1040
rect 11595 990 11600 1010
rect 11620 990 11625 1010
rect 11595 960 11625 990
rect 11595 940 11600 960
rect 11620 940 11625 960
rect 11595 930 11625 940
rect 11650 1160 11680 1170
rect 11650 1140 11655 1160
rect 11675 1140 11680 1160
rect 11650 1110 11680 1140
rect 11650 1090 11655 1110
rect 11675 1090 11680 1110
rect 11650 1060 11680 1090
rect 11650 1040 11655 1060
rect 11675 1040 11680 1060
rect 11650 1010 11680 1040
rect 11650 990 11655 1010
rect 11675 990 11680 1010
rect 11650 960 11680 990
rect 11650 940 11655 960
rect 11675 940 11680 960
rect 11650 930 11680 940
rect 11705 1160 11735 1170
rect 11705 1140 11710 1160
rect 11730 1140 11735 1160
rect 11705 1110 11735 1140
rect 11705 1090 11710 1110
rect 11730 1090 11735 1110
rect 11705 1060 11735 1090
rect 11705 1040 11710 1060
rect 11730 1040 11735 1060
rect 11705 1010 11735 1040
rect 11705 990 11710 1010
rect 11730 990 11735 1010
rect 11705 960 11735 990
rect 11705 940 11710 960
rect 11730 940 11735 960
rect 11705 930 11735 940
rect 11760 1160 11790 1170
rect 11760 1140 11765 1160
rect 11785 1140 11790 1160
rect 11760 1110 11790 1140
rect 11760 1090 11765 1110
rect 11785 1090 11790 1110
rect 11760 1060 11790 1090
rect 11760 1040 11765 1060
rect 11785 1040 11790 1060
rect 11760 1010 11790 1040
rect 11760 990 11765 1010
rect 11785 990 11790 1010
rect 11760 960 11790 990
rect 11760 940 11765 960
rect 11785 940 11790 960
rect 11760 930 11790 940
rect 11815 1160 11845 1170
rect 11815 1140 11820 1160
rect 11840 1140 11845 1160
rect 11815 1110 11845 1140
rect 11815 1090 11820 1110
rect 11840 1090 11845 1110
rect 11815 1060 11845 1090
rect 11815 1040 11820 1060
rect 11840 1040 11845 1060
rect 11815 1010 11845 1040
rect 11815 990 11820 1010
rect 11840 990 11845 1010
rect 11815 960 11845 990
rect 11815 940 11820 960
rect 11840 940 11845 960
rect 11815 930 11845 940
rect 11870 1160 11900 1170
rect 11870 1140 11875 1160
rect 11895 1140 11900 1160
rect 11870 1110 11900 1140
rect 11870 1090 11875 1110
rect 11895 1090 11900 1110
rect 11870 1060 11900 1090
rect 11870 1040 11875 1060
rect 11895 1040 11900 1060
rect 11870 1010 11900 1040
rect 11870 990 11875 1010
rect 11895 990 11900 1010
rect 11870 960 11900 990
rect 11870 940 11875 960
rect 11895 940 11900 960
rect 11870 930 11900 940
rect 11925 1160 11955 1170
rect 11925 1140 11930 1160
rect 11950 1140 11955 1160
rect 11925 1110 11955 1140
rect 11925 1090 11930 1110
rect 11950 1090 11955 1110
rect 11925 1060 11955 1090
rect 11925 1040 11930 1060
rect 11950 1040 11955 1060
rect 11925 1010 11955 1040
rect 11925 990 11930 1010
rect 11950 990 11955 1010
rect 11925 960 11955 990
rect 11925 940 11930 960
rect 11950 940 11955 960
rect 11925 930 11955 940
rect 11980 1160 12010 1170
rect 11980 1140 11985 1160
rect 12005 1140 12010 1160
rect 11980 1110 12010 1140
rect 11980 1090 11985 1110
rect 12005 1090 12010 1110
rect 11980 1060 12010 1090
rect 11980 1040 11985 1060
rect 12005 1040 12010 1060
rect 11980 1010 12010 1040
rect 11980 990 11985 1010
rect 12005 990 12010 1010
rect 11980 960 12010 990
rect 11980 940 11985 960
rect 12005 940 12010 960
rect 11980 930 12010 940
rect 12035 1160 12065 1170
rect 12035 1140 12040 1160
rect 12060 1140 12065 1160
rect 12035 1110 12065 1140
rect 12035 1090 12040 1110
rect 12060 1090 12065 1110
rect 12035 1060 12065 1090
rect 12035 1040 12040 1060
rect 12060 1040 12065 1060
rect 12035 1010 12065 1040
rect 12035 990 12040 1010
rect 12060 990 12065 1010
rect 12035 960 12065 990
rect 12035 940 12040 960
rect 12060 940 12065 960
rect 12035 930 12065 940
rect 12090 1160 12120 1170
rect 12090 1140 12095 1160
rect 12115 1140 12120 1160
rect 12090 1110 12120 1140
rect 12090 1090 12095 1110
rect 12115 1090 12120 1110
rect 12090 1060 12120 1090
rect 12090 1040 12095 1060
rect 12115 1040 12120 1060
rect 12090 1010 12120 1040
rect 12090 990 12095 1010
rect 12115 990 12120 1010
rect 12090 960 12120 990
rect 12090 940 12095 960
rect 12115 940 12120 960
rect 12090 930 12120 940
rect 12145 1160 12175 1170
rect 12145 1140 12150 1160
rect 12170 1140 12175 1160
rect 12145 1110 12175 1140
rect 12145 1090 12150 1110
rect 12170 1090 12175 1110
rect 12145 1060 12175 1090
rect 12145 1040 12150 1060
rect 12170 1040 12175 1060
rect 12145 1010 12175 1040
rect 12145 990 12150 1010
rect 12170 990 12175 1010
rect 12145 960 12175 990
rect 12145 940 12150 960
rect 12170 940 12175 960
rect 12145 930 12175 940
rect 12200 1160 12230 1170
rect 12200 1140 12205 1160
rect 12225 1140 12230 1160
rect 12200 1110 12230 1140
rect 12200 1090 12205 1110
rect 12225 1090 12230 1110
rect 12200 1060 12230 1090
rect 12200 1040 12205 1060
rect 12225 1040 12230 1060
rect 12200 1010 12230 1040
rect 12200 990 12205 1010
rect 12225 990 12230 1010
rect 12200 960 12230 990
rect 12200 940 12205 960
rect 12225 940 12230 960
rect 12200 930 12230 940
rect 12255 1160 12285 1170
rect 12255 1140 12260 1160
rect 12280 1140 12285 1160
rect 12255 1110 12285 1140
rect 12255 1090 12260 1110
rect 12280 1090 12285 1110
rect 12255 1060 12285 1090
rect 12255 1040 12260 1060
rect 12280 1040 12285 1060
rect 12255 1010 12285 1040
rect 12255 990 12260 1010
rect 12280 990 12285 1010
rect 12255 960 12285 990
rect 12255 940 12260 960
rect 12280 940 12285 960
rect 12255 930 12285 940
rect 12310 1160 12340 1170
rect 12310 1140 12315 1160
rect 12335 1140 12340 1160
rect 12310 1110 12340 1140
rect 12310 1090 12315 1110
rect 12335 1090 12340 1110
rect 12310 1060 12340 1090
rect 12310 1040 12315 1060
rect 12335 1040 12340 1060
rect 12310 1010 12340 1040
rect 12310 990 12315 1010
rect 12335 990 12340 1010
rect 12310 960 12340 990
rect 12310 940 12315 960
rect 12335 940 12340 960
rect 12310 930 12340 940
rect 12365 1160 12395 1170
rect 12365 1140 12370 1160
rect 12390 1140 12395 1160
rect 12365 1110 12395 1140
rect 12365 1090 12370 1110
rect 12390 1090 12395 1110
rect 12365 1060 12395 1090
rect 12365 1040 12370 1060
rect 12390 1040 12395 1060
rect 12365 1010 12395 1040
rect 12365 990 12370 1010
rect 12390 990 12395 1010
rect 12365 960 12395 990
rect 12365 940 12370 960
rect 12390 940 12395 960
rect 12365 930 12395 940
rect 12420 1160 12450 1170
rect 12420 1140 12425 1160
rect 12445 1140 12450 1160
rect 12420 1110 12450 1140
rect 12420 1090 12425 1110
rect 12445 1090 12450 1110
rect 12420 1060 12450 1090
rect 12420 1040 12425 1060
rect 12445 1040 12450 1060
rect 12420 1010 12450 1040
rect 12420 990 12425 1010
rect 12445 990 12450 1010
rect 12420 960 12450 990
rect 12420 940 12425 960
rect 12445 940 12450 960
rect 12420 930 12450 940
rect 12475 1160 12505 1170
rect 12475 1140 12480 1160
rect 12500 1140 12505 1160
rect 12475 1110 12505 1140
rect 12475 1090 12480 1110
rect 12500 1090 12505 1110
rect 12475 1060 12505 1090
rect 12475 1040 12480 1060
rect 12500 1040 12505 1060
rect 12475 1010 12505 1040
rect 12475 990 12480 1010
rect 12500 990 12505 1010
rect 12475 960 12505 990
rect 12475 940 12480 960
rect 12500 940 12505 960
rect 12475 930 12505 940
rect 12530 1160 12560 1170
rect 12530 1140 12535 1160
rect 12555 1140 12560 1160
rect 12530 1110 12560 1140
rect 12530 1090 12535 1110
rect 12555 1090 12560 1110
rect 12530 1060 12560 1090
rect 12530 1040 12535 1060
rect 12555 1040 12560 1060
rect 12530 1010 12560 1040
rect 12530 990 12535 1010
rect 12555 990 12560 1010
rect 12530 960 12560 990
rect 12530 940 12535 960
rect 12555 940 12560 960
rect 12530 930 12560 940
rect 12585 1160 12655 1170
rect 12585 1140 12590 1160
rect 12610 1140 12630 1160
rect 12650 1140 12655 1160
rect 12585 1110 12655 1140
rect 12585 1090 12590 1110
rect 12610 1090 12630 1110
rect 12650 1090 12655 1110
rect 12585 1060 12655 1090
rect 12585 1040 12590 1060
rect 12610 1040 12630 1060
rect 12650 1040 12655 1060
rect 12585 1010 12655 1040
rect 12585 990 12590 1010
rect 12610 990 12630 1010
rect 12650 990 12655 1010
rect 12890 1165 12960 1190
rect 12890 1145 12895 1165
rect 12915 1145 12935 1165
rect 12955 1145 12960 1165
rect 12890 1115 12960 1145
rect 12890 1095 12895 1115
rect 12915 1095 12935 1115
rect 12955 1095 12960 1115
rect 12890 1070 12960 1095
rect 12890 1050 12895 1070
rect 12915 1050 12935 1070
rect 12955 1050 12960 1070
rect 12890 1025 12960 1050
rect 12890 1005 12895 1025
rect 12915 1005 12935 1025
rect 12955 1005 12960 1025
rect 12890 995 12960 1005
rect 13030 1255 13060 1265
rect 13030 1235 13035 1255
rect 13055 1235 13060 1255
rect 13030 1210 13060 1235
rect 13030 1190 13035 1210
rect 13055 1190 13060 1210
rect 13030 1165 13060 1190
rect 13030 1145 13035 1165
rect 13055 1145 13060 1165
rect 13030 1115 13060 1145
rect 13030 1095 13035 1115
rect 13055 1095 13060 1115
rect 13030 1070 13060 1095
rect 13030 1050 13035 1070
rect 13055 1050 13060 1070
rect 13030 1025 13060 1050
rect 13030 1005 13035 1025
rect 13055 1005 13060 1025
rect 13030 995 13060 1005
rect 13130 1255 13160 1265
rect 13130 1235 13135 1255
rect 13155 1235 13160 1255
rect 13130 1210 13160 1235
rect 13130 1190 13135 1210
rect 13155 1190 13160 1210
rect 13130 1165 13160 1190
rect 13130 1145 13135 1165
rect 13155 1145 13160 1165
rect 13130 1115 13160 1145
rect 13130 1095 13135 1115
rect 13155 1095 13160 1115
rect 13130 1070 13160 1095
rect 13130 1050 13135 1070
rect 13155 1050 13160 1070
rect 13130 1025 13160 1050
rect 13130 1005 13135 1025
rect 13155 1005 13160 1025
rect 13130 995 13160 1005
rect 13230 1255 13260 1265
rect 13230 1235 13235 1255
rect 13255 1235 13260 1255
rect 13230 1210 13260 1235
rect 13230 1190 13235 1210
rect 13255 1190 13260 1210
rect 13230 1165 13260 1190
rect 13230 1145 13235 1165
rect 13255 1145 13260 1165
rect 13230 1115 13260 1145
rect 13230 1095 13235 1115
rect 13255 1095 13260 1115
rect 13230 1070 13260 1095
rect 13230 1050 13235 1070
rect 13255 1050 13260 1070
rect 13230 1025 13260 1050
rect 13230 1005 13235 1025
rect 13255 1005 13260 1025
rect 13230 995 13260 1005
rect 13330 1255 13360 1265
rect 13330 1235 13335 1255
rect 13355 1235 13360 1255
rect 13330 1210 13360 1235
rect 13330 1190 13335 1210
rect 13355 1190 13360 1210
rect 13330 1165 13360 1190
rect 13330 1145 13335 1165
rect 13355 1145 13360 1165
rect 13330 1115 13360 1145
rect 13330 1095 13335 1115
rect 13355 1095 13360 1115
rect 13330 1070 13360 1095
rect 13330 1050 13335 1070
rect 13355 1050 13360 1070
rect 13330 1025 13360 1050
rect 13330 1005 13335 1025
rect 13355 1005 13360 1025
rect 13330 995 13360 1005
rect 13430 1255 13460 1265
rect 13430 1235 13435 1255
rect 13455 1235 13460 1255
rect 13430 1210 13460 1235
rect 13430 1190 13435 1210
rect 13455 1190 13460 1210
rect 13430 1165 13460 1190
rect 13430 1145 13435 1165
rect 13455 1145 13460 1165
rect 13430 1115 13460 1145
rect 13430 1095 13435 1115
rect 13455 1095 13460 1115
rect 13430 1070 13460 1095
rect 13430 1050 13435 1070
rect 13455 1050 13460 1070
rect 13430 1025 13460 1050
rect 13430 1005 13435 1025
rect 13455 1005 13460 1025
rect 13430 995 13460 1005
rect 13530 1255 13560 1265
rect 13530 1235 13535 1255
rect 13555 1235 13560 1255
rect 13530 1210 13560 1235
rect 13530 1190 13535 1210
rect 13555 1190 13560 1210
rect 13530 1165 13560 1190
rect 13530 1145 13535 1165
rect 13555 1145 13560 1165
rect 13530 1115 13560 1145
rect 13530 1095 13535 1115
rect 13555 1095 13560 1115
rect 13530 1070 13560 1095
rect 13530 1050 13535 1070
rect 13555 1050 13560 1070
rect 13530 1025 13560 1050
rect 13530 1005 13535 1025
rect 13555 1005 13560 1025
rect 13530 995 13560 1005
rect 13630 1255 13660 1265
rect 13630 1235 13635 1255
rect 13655 1235 13660 1255
rect 13630 1210 13660 1235
rect 13630 1190 13635 1210
rect 13655 1190 13660 1210
rect 13630 1165 13660 1190
rect 13630 1145 13635 1165
rect 13655 1145 13660 1165
rect 13630 1115 13660 1145
rect 13630 1095 13635 1115
rect 13655 1095 13660 1115
rect 13630 1070 13660 1095
rect 13630 1050 13635 1070
rect 13655 1050 13660 1070
rect 13630 1025 13660 1050
rect 13630 1005 13635 1025
rect 13655 1005 13660 1025
rect 13630 995 13660 1005
rect 13730 1255 13760 1265
rect 13730 1235 13735 1255
rect 13755 1235 13760 1255
rect 13730 1210 13760 1235
rect 13730 1190 13735 1210
rect 13755 1190 13760 1210
rect 13730 1165 13760 1190
rect 13730 1145 13735 1165
rect 13755 1145 13760 1165
rect 13730 1115 13760 1145
rect 13730 1095 13735 1115
rect 13755 1095 13760 1115
rect 13730 1070 13760 1095
rect 13730 1050 13735 1070
rect 13755 1050 13760 1070
rect 13730 1025 13760 1050
rect 13730 1005 13735 1025
rect 13755 1005 13760 1025
rect 13730 995 13760 1005
rect 13830 1255 13860 1265
rect 13830 1235 13835 1255
rect 13855 1235 13860 1255
rect 13830 1210 13860 1235
rect 13830 1190 13835 1210
rect 13855 1190 13860 1210
rect 13830 1165 13860 1190
rect 13830 1145 13835 1165
rect 13855 1145 13860 1165
rect 13830 1115 13860 1145
rect 13830 1095 13835 1115
rect 13855 1095 13860 1115
rect 13830 1070 13860 1095
rect 13830 1050 13835 1070
rect 13855 1050 13860 1070
rect 13830 1025 13860 1050
rect 13830 1005 13835 1025
rect 13855 1005 13860 1025
rect 13830 995 13860 1005
rect 13930 1255 13960 1265
rect 13930 1235 13935 1255
rect 13955 1235 13960 1255
rect 13930 1210 13960 1235
rect 13930 1190 13935 1210
rect 13955 1190 13960 1210
rect 13930 1165 13960 1190
rect 13930 1145 13935 1165
rect 13955 1145 13960 1165
rect 13930 1115 13960 1145
rect 13930 1095 13935 1115
rect 13955 1095 13960 1115
rect 13930 1070 13960 1095
rect 13930 1050 13935 1070
rect 13955 1050 13960 1070
rect 13930 1025 13960 1050
rect 13930 1005 13935 1025
rect 13955 1005 13960 1025
rect 13930 995 13960 1005
rect 14030 1255 14060 1265
rect 14030 1235 14035 1255
rect 14055 1235 14060 1255
rect 14030 1210 14060 1235
rect 14030 1190 14035 1210
rect 14055 1190 14060 1210
rect 14030 1165 14060 1190
rect 14030 1145 14035 1165
rect 14055 1145 14060 1165
rect 14030 1115 14060 1145
rect 14030 1095 14035 1115
rect 14055 1095 14060 1115
rect 14030 1070 14060 1095
rect 14030 1050 14035 1070
rect 14055 1050 14060 1070
rect 14030 1025 14060 1050
rect 14030 1005 14035 1025
rect 14055 1005 14060 1025
rect 14030 995 14060 1005
rect 14130 1255 14200 1265
rect 14130 1235 14135 1255
rect 14155 1235 14175 1255
rect 14195 1235 14200 1255
rect 18815 1250 18825 1270
rect 18845 1250 18855 1270
rect 18815 1240 18855 1250
rect 18925 1270 18965 1280
rect 18925 1250 18935 1270
rect 18955 1250 18965 1270
rect 18925 1240 18965 1250
rect 19035 1270 19075 1280
rect 19035 1250 19045 1270
rect 19065 1250 19075 1270
rect 19035 1240 19075 1250
rect 19145 1270 19185 1280
rect 19145 1250 19155 1270
rect 19175 1250 19185 1270
rect 19145 1240 19185 1250
rect 19255 1270 19295 1280
rect 19255 1250 19265 1270
rect 19285 1250 19295 1270
rect 19255 1240 19295 1250
rect 19315 1270 19345 1280
rect 19315 1250 19320 1270
rect 19340 1250 19345 1270
rect 19315 1240 19345 1250
rect 19365 1270 19405 1280
rect 19365 1250 19375 1270
rect 19395 1250 19405 1270
rect 19365 1240 19405 1250
rect 19475 1270 19515 1280
rect 19475 1250 19485 1270
rect 19505 1250 19515 1270
rect 19475 1240 19515 1250
rect 19585 1270 19625 1280
rect 19585 1250 19595 1270
rect 19615 1250 19625 1270
rect 19585 1240 19625 1250
rect 19695 1270 19735 1280
rect 19695 1250 19705 1270
rect 19725 1250 19735 1270
rect 19695 1240 19735 1250
rect 19805 1270 19845 1280
rect 19805 1250 19815 1270
rect 19835 1250 19845 1270
rect 19805 1240 19845 1250
rect 19915 1270 19955 1280
rect 19915 1250 19925 1270
rect 19945 1250 19955 1270
rect 19915 1240 19955 1250
rect 20025 1270 20065 1280
rect 20025 1250 20035 1270
rect 20055 1250 20065 1270
rect 20095 1265 20105 1285
rect 20125 1265 20135 1285
rect 20095 1255 20135 1265
rect 20445 1285 20485 1295
rect 20445 1265 20455 1285
rect 20475 1265 20485 1285
rect 20445 1255 20485 1265
rect 20560 1285 20600 1295
rect 20560 1265 20570 1285
rect 20590 1265 20600 1285
rect 20560 1255 20600 1265
rect 20750 1285 20790 1295
rect 20750 1265 20760 1285
rect 20780 1265 20790 1285
rect 20750 1255 20790 1265
rect 20865 1285 20905 1295
rect 20865 1265 20875 1285
rect 20895 1265 20905 1285
rect 20865 1255 20905 1265
rect 20025 1240 20065 1250
rect 14130 1210 14200 1235
rect 18825 1220 18845 1240
rect 18935 1220 18955 1240
rect 19045 1220 19065 1240
rect 19155 1220 19175 1240
rect 19265 1220 19285 1240
rect 19375 1220 19395 1240
rect 19485 1220 19505 1240
rect 19595 1220 19615 1240
rect 19705 1220 19725 1240
rect 19815 1220 19835 1240
rect 19925 1220 19945 1240
rect 20035 1220 20055 1240
rect 20600 1225 20640 1235
rect 14130 1190 14135 1210
rect 14155 1190 14175 1210
rect 14195 1190 14200 1210
rect 14130 1165 14200 1190
rect 14130 1145 14135 1165
rect 14155 1145 14175 1165
rect 14195 1145 14200 1165
rect 14130 1115 14200 1145
rect 14130 1095 14135 1115
rect 14155 1095 14175 1115
rect 14195 1095 14200 1115
rect 14130 1070 14200 1095
rect 14130 1050 14135 1070
rect 14155 1050 14175 1070
rect 14195 1050 14200 1070
rect 14130 1025 14200 1050
rect 14130 1005 14135 1025
rect 14155 1005 14175 1025
rect 14195 1005 14200 1025
rect 14130 995 14200 1005
rect 18670 1210 18740 1220
rect 18670 1190 18675 1210
rect 18695 1190 18715 1210
rect 18735 1190 18740 1210
rect 18670 1160 18740 1190
rect 18670 1140 18675 1160
rect 18695 1140 18715 1160
rect 18735 1140 18740 1160
rect 18670 1110 18740 1140
rect 18670 1090 18675 1110
rect 18695 1090 18715 1110
rect 18735 1090 18740 1110
rect 18670 1060 18740 1090
rect 18670 1040 18675 1060
rect 18695 1040 18715 1060
rect 18735 1040 18740 1060
rect 18670 1010 18740 1040
rect 12585 960 12655 990
rect 12895 975 12915 995
rect 13135 975 13155 995
rect 13335 975 13355 995
rect 13535 975 13555 995
rect 13735 975 13755 995
rect 13935 975 13955 995
rect 14175 975 14195 995
rect 18670 990 18675 1010
rect 18695 990 18715 1010
rect 18735 990 18740 1010
rect 18670 980 18740 990
rect 18765 1210 18795 1220
rect 18765 1190 18770 1210
rect 18790 1190 18795 1210
rect 18765 1160 18795 1190
rect 18765 1140 18770 1160
rect 18790 1140 18795 1160
rect 18765 1110 18795 1140
rect 18765 1090 18770 1110
rect 18790 1090 18795 1110
rect 18765 1060 18795 1090
rect 18765 1040 18770 1060
rect 18790 1040 18795 1060
rect 18765 1010 18795 1040
rect 18765 990 18770 1010
rect 18790 990 18795 1010
rect 18765 980 18795 990
rect 18820 1210 18850 1220
rect 18820 1190 18825 1210
rect 18845 1190 18850 1210
rect 18820 1160 18850 1190
rect 18820 1140 18825 1160
rect 18845 1140 18850 1160
rect 18820 1110 18850 1140
rect 18820 1090 18825 1110
rect 18845 1090 18850 1110
rect 18820 1060 18850 1090
rect 18820 1040 18825 1060
rect 18845 1040 18850 1060
rect 18820 1010 18850 1040
rect 18820 990 18825 1010
rect 18845 990 18850 1010
rect 18820 980 18850 990
rect 18875 1210 18905 1220
rect 18875 1190 18880 1210
rect 18900 1190 18905 1210
rect 18875 1160 18905 1190
rect 18875 1140 18880 1160
rect 18900 1140 18905 1160
rect 18875 1110 18905 1140
rect 18875 1090 18880 1110
rect 18900 1090 18905 1110
rect 18875 1060 18905 1090
rect 18875 1040 18880 1060
rect 18900 1040 18905 1060
rect 18875 1010 18905 1040
rect 18875 990 18880 1010
rect 18900 990 18905 1010
rect 18875 980 18905 990
rect 18930 1210 18960 1220
rect 18930 1190 18935 1210
rect 18955 1190 18960 1210
rect 18930 1160 18960 1190
rect 18930 1140 18935 1160
rect 18955 1140 18960 1160
rect 18930 1110 18960 1140
rect 18930 1090 18935 1110
rect 18955 1090 18960 1110
rect 18930 1060 18960 1090
rect 18930 1040 18935 1060
rect 18955 1040 18960 1060
rect 18930 1010 18960 1040
rect 18930 990 18935 1010
rect 18955 990 18960 1010
rect 18930 980 18960 990
rect 18985 1210 19015 1220
rect 18985 1190 18990 1210
rect 19010 1190 19015 1210
rect 18985 1160 19015 1190
rect 18985 1140 18990 1160
rect 19010 1140 19015 1160
rect 18985 1110 19015 1140
rect 18985 1090 18990 1110
rect 19010 1090 19015 1110
rect 18985 1060 19015 1090
rect 18985 1040 18990 1060
rect 19010 1040 19015 1060
rect 18985 1010 19015 1040
rect 18985 990 18990 1010
rect 19010 990 19015 1010
rect 18985 980 19015 990
rect 19040 1210 19070 1220
rect 19040 1190 19045 1210
rect 19065 1190 19070 1210
rect 19040 1160 19070 1190
rect 19040 1140 19045 1160
rect 19065 1140 19070 1160
rect 19040 1110 19070 1140
rect 19040 1090 19045 1110
rect 19065 1090 19070 1110
rect 19040 1060 19070 1090
rect 19040 1040 19045 1060
rect 19065 1040 19070 1060
rect 19040 1010 19070 1040
rect 19040 990 19045 1010
rect 19065 990 19070 1010
rect 19040 980 19070 990
rect 19095 1210 19125 1220
rect 19095 1190 19100 1210
rect 19120 1190 19125 1210
rect 19095 1160 19125 1190
rect 19095 1140 19100 1160
rect 19120 1140 19125 1160
rect 19095 1110 19125 1140
rect 19095 1090 19100 1110
rect 19120 1090 19125 1110
rect 19095 1060 19125 1090
rect 19095 1040 19100 1060
rect 19120 1040 19125 1060
rect 19095 1010 19125 1040
rect 19095 990 19100 1010
rect 19120 990 19125 1010
rect 19095 980 19125 990
rect 19150 1210 19180 1220
rect 19150 1190 19155 1210
rect 19175 1190 19180 1210
rect 19150 1160 19180 1190
rect 19150 1140 19155 1160
rect 19175 1140 19180 1160
rect 19150 1110 19180 1140
rect 19150 1090 19155 1110
rect 19175 1090 19180 1110
rect 19150 1060 19180 1090
rect 19150 1040 19155 1060
rect 19175 1040 19180 1060
rect 19150 1010 19180 1040
rect 19150 990 19155 1010
rect 19175 990 19180 1010
rect 19150 980 19180 990
rect 19205 1210 19235 1220
rect 19205 1190 19210 1210
rect 19230 1190 19235 1210
rect 19205 1160 19235 1190
rect 19205 1140 19210 1160
rect 19230 1140 19235 1160
rect 19205 1110 19235 1140
rect 19205 1090 19210 1110
rect 19230 1090 19235 1110
rect 19205 1060 19235 1090
rect 19205 1040 19210 1060
rect 19230 1040 19235 1060
rect 19205 1010 19235 1040
rect 19205 990 19210 1010
rect 19230 990 19235 1010
rect 19205 980 19235 990
rect 19260 1210 19290 1220
rect 19260 1190 19265 1210
rect 19285 1190 19290 1210
rect 19260 1160 19290 1190
rect 19260 1140 19265 1160
rect 19285 1140 19290 1160
rect 19260 1110 19290 1140
rect 19260 1090 19265 1110
rect 19285 1090 19290 1110
rect 19260 1060 19290 1090
rect 19260 1040 19265 1060
rect 19285 1040 19290 1060
rect 19260 1010 19290 1040
rect 19260 990 19265 1010
rect 19285 990 19290 1010
rect 19260 980 19290 990
rect 19315 1210 19345 1220
rect 19315 1190 19320 1210
rect 19340 1190 19345 1210
rect 19315 1160 19345 1190
rect 19315 1140 19320 1160
rect 19340 1140 19345 1160
rect 19315 1110 19345 1140
rect 19315 1090 19320 1110
rect 19340 1090 19345 1110
rect 19315 1060 19345 1090
rect 19315 1040 19320 1060
rect 19340 1040 19345 1060
rect 19315 1010 19345 1040
rect 19315 990 19320 1010
rect 19340 990 19345 1010
rect 19315 980 19345 990
rect 19370 1210 19400 1220
rect 19370 1190 19375 1210
rect 19395 1190 19400 1210
rect 19370 1160 19400 1190
rect 19370 1140 19375 1160
rect 19395 1140 19400 1160
rect 19370 1110 19400 1140
rect 19370 1090 19375 1110
rect 19395 1090 19400 1110
rect 19370 1060 19400 1090
rect 19370 1040 19375 1060
rect 19395 1040 19400 1060
rect 19370 1010 19400 1040
rect 19370 990 19375 1010
rect 19395 990 19400 1010
rect 19370 980 19400 990
rect 19425 1210 19455 1220
rect 19425 1190 19430 1210
rect 19450 1190 19455 1210
rect 19425 1160 19455 1190
rect 19425 1140 19430 1160
rect 19450 1140 19455 1160
rect 19425 1110 19455 1140
rect 19425 1090 19430 1110
rect 19450 1090 19455 1110
rect 19425 1060 19455 1090
rect 19425 1040 19430 1060
rect 19450 1040 19455 1060
rect 19425 1010 19455 1040
rect 19425 990 19430 1010
rect 19450 990 19455 1010
rect 19425 980 19455 990
rect 19480 1210 19510 1220
rect 19480 1190 19485 1210
rect 19505 1190 19510 1210
rect 19480 1160 19510 1190
rect 19480 1140 19485 1160
rect 19505 1140 19510 1160
rect 19480 1110 19510 1140
rect 19480 1090 19485 1110
rect 19505 1090 19510 1110
rect 19480 1060 19510 1090
rect 19480 1040 19485 1060
rect 19505 1040 19510 1060
rect 19480 1010 19510 1040
rect 19480 990 19485 1010
rect 19505 990 19510 1010
rect 19480 980 19510 990
rect 19535 1210 19565 1220
rect 19535 1190 19540 1210
rect 19560 1190 19565 1210
rect 19535 1160 19565 1190
rect 19535 1140 19540 1160
rect 19560 1140 19565 1160
rect 19535 1110 19565 1140
rect 19535 1090 19540 1110
rect 19560 1090 19565 1110
rect 19535 1060 19565 1090
rect 19535 1040 19540 1060
rect 19560 1040 19565 1060
rect 19535 1010 19565 1040
rect 19535 990 19540 1010
rect 19560 990 19565 1010
rect 19535 980 19565 990
rect 19590 1210 19620 1220
rect 19590 1190 19595 1210
rect 19615 1190 19620 1210
rect 19590 1160 19620 1190
rect 19590 1140 19595 1160
rect 19615 1140 19620 1160
rect 19590 1110 19620 1140
rect 19590 1090 19595 1110
rect 19615 1090 19620 1110
rect 19590 1060 19620 1090
rect 19590 1040 19595 1060
rect 19615 1040 19620 1060
rect 19590 1010 19620 1040
rect 19590 990 19595 1010
rect 19615 990 19620 1010
rect 19590 980 19620 990
rect 19645 1210 19675 1220
rect 19645 1190 19650 1210
rect 19670 1190 19675 1210
rect 19645 1160 19675 1190
rect 19645 1140 19650 1160
rect 19670 1140 19675 1160
rect 19645 1110 19675 1140
rect 19645 1090 19650 1110
rect 19670 1090 19675 1110
rect 19645 1060 19675 1090
rect 19645 1040 19650 1060
rect 19670 1040 19675 1060
rect 19645 1010 19675 1040
rect 19645 990 19650 1010
rect 19670 990 19675 1010
rect 19645 980 19675 990
rect 19700 1210 19730 1220
rect 19700 1190 19705 1210
rect 19725 1190 19730 1210
rect 19700 1160 19730 1190
rect 19700 1140 19705 1160
rect 19725 1140 19730 1160
rect 19700 1110 19730 1140
rect 19700 1090 19705 1110
rect 19725 1090 19730 1110
rect 19700 1060 19730 1090
rect 19700 1040 19705 1060
rect 19725 1040 19730 1060
rect 19700 1010 19730 1040
rect 19700 990 19705 1010
rect 19725 990 19730 1010
rect 19700 980 19730 990
rect 19755 1210 19785 1220
rect 19755 1190 19760 1210
rect 19780 1190 19785 1210
rect 19755 1160 19785 1190
rect 19755 1140 19760 1160
rect 19780 1140 19785 1160
rect 19755 1110 19785 1140
rect 19755 1090 19760 1110
rect 19780 1090 19785 1110
rect 19755 1060 19785 1090
rect 19755 1040 19760 1060
rect 19780 1040 19785 1060
rect 19755 1010 19785 1040
rect 19755 990 19760 1010
rect 19780 990 19785 1010
rect 19755 980 19785 990
rect 19810 1210 19840 1220
rect 19810 1190 19815 1210
rect 19835 1190 19840 1210
rect 19810 1160 19840 1190
rect 19810 1140 19815 1160
rect 19835 1140 19840 1160
rect 19810 1110 19840 1140
rect 19810 1090 19815 1110
rect 19835 1090 19840 1110
rect 19810 1060 19840 1090
rect 19810 1040 19815 1060
rect 19835 1040 19840 1060
rect 19810 1010 19840 1040
rect 19810 990 19815 1010
rect 19835 990 19840 1010
rect 19810 980 19840 990
rect 19865 1210 19895 1220
rect 19865 1190 19870 1210
rect 19890 1190 19895 1210
rect 19865 1160 19895 1190
rect 19865 1140 19870 1160
rect 19890 1140 19895 1160
rect 19865 1110 19895 1140
rect 19865 1090 19870 1110
rect 19890 1090 19895 1110
rect 19865 1060 19895 1090
rect 19865 1040 19870 1060
rect 19890 1040 19895 1060
rect 19865 1010 19895 1040
rect 19865 990 19870 1010
rect 19890 990 19895 1010
rect 19865 980 19895 990
rect 19920 1210 19950 1220
rect 19920 1190 19925 1210
rect 19945 1190 19950 1210
rect 19920 1160 19950 1190
rect 19920 1140 19925 1160
rect 19945 1140 19950 1160
rect 19920 1110 19950 1140
rect 19920 1090 19925 1110
rect 19945 1090 19950 1110
rect 19920 1060 19950 1090
rect 19920 1040 19925 1060
rect 19945 1040 19950 1060
rect 19920 1010 19950 1040
rect 19920 990 19925 1010
rect 19945 990 19950 1010
rect 19920 980 19950 990
rect 19975 1210 20005 1220
rect 19975 1190 19980 1210
rect 20000 1190 20005 1210
rect 19975 1160 20005 1190
rect 19975 1140 19980 1160
rect 20000 1140 20005 1160
rect 19975 1110 20005 1140
rect 19975 1090 19980 1110
rect 20000 1090 20005 1110
rect 19975 1060 20005 1090
rect 19975 1040 19980 1060
rect 20000 1040 20005 1060
rect 19975 1010 20005 1040
rect 19975 990 19980 1010
rect 20000 990 20005 1010
rect 19975 980 20005 990
rect 20030 1210 20060 1220
rect 20030 1190 20035 1210
rect 20055 1190 20060 1210
rect 20030 1160 20060 1190
rect 20030 1140 20035 1160
rect 20055 1140 20060 1160
rect 20030 1110 20060 1140
rect 20030 1090 20035 1110
rect 20055 1090 20060 1110
rect 20030 1060 20060 1090
rect 20030 1040 20035 1060
rect 20055 1040 20060 1060
rect 20030 1010 20060 1040
rect 20030 990 20035 1010
rect 20055 990 20060 1010
rect 20030 980 20060 990
rect 20085 1210 20155 1220
rect 20085 1190 20090 1210
rect 20110 1190 20130 1210
rect 20150 1190 20155 1210
rect 20600 1205 20610 1225
rect 20630 1205 20640 1225
rect 20600 1195 20640 1205
rect 20660 1225 20690 1235
rect 20660 1205 20665 1225
rect 20685 1205 20690 1225
rect 20660 1195 20690 1205
rect 20710 1225 20750 1235
rect 20710 1205 20720 1225
rect 20740 1205 20750 1225
rect 20710 1195 20750 1205
rect 20085 1160 20155 1190
rect 20610 1175 20630 1195
rect 20720 1175 20740 1195
rect 20085 1140 20090 1160
rect 20110 1140 20130 1160
rect 20150 1140 20155 1160
rect 20085 1110 20155 1140
rect 20085 1090 20090 1110
rect 20110 1090 20130 1110
rect 20150 1090 20155 1110
rect 20085 1060 20155 1090
rect 20085 1040 20090 1060
rect 20110 1040 20130 1060
rect 20150 1040 20155 1060
rect 20085 1010 20155 1040
rect 20510 1165 20580 1175
rect 20510 1145 20515 1165
rect 20535 1145 20555 1165
rect 20575 1145 20580 1165
rect 20510 1115 20580 1145
rect 20510 1095 20515 1115
rect 20535 1095 20555 1115
rect 20575 1095 20580 1115
rect 20510 1065 20580 1095
rect 20510 1045 20515 1065
rect 20535 1045 20555 1065
rect 20575 1045 20580 1065
rect 20510 1035 20580 1045
rect 20605 1165 20635 1175
rect 20605 1145 20610 1165
rect 20630 1145 20635 1165
rect 20605 1115 20635 1145
rect 20605 1095 20610 1115
rect 20630 1095 20635 1115
rect 20605 1065 20635 1095
rect 20605 1045 20610 1065
rect 20630 1045 20635 1065
rect 20605 1035 20635 1045
rect 20660 1165 20690 1175
rect 20660 1145 20665 1165
rect 20685 1145 20690 1165
rect 20660 1115 20690 1145
rect 20660 1095 20665 1115
rect 20685 1095 20690 1115
rect 20660 1065 20690 1095
rect 20660 1045 20665 1065
rect 20685 1045 20690 1065
rect 20660 1035 20690 1045
rect 20715 1165 20745 1175
rect 20715 1145 20720 1165
rect 20740 1145 20745 1165
rect 20715 1115 20745 1145
rect 20715 1095 20720 1115
rect 20740 1095 20745 1115
rect 20715 1065 20745 1095
rect 20715 1045 20720 1065
rect 20740 1045 20745 1065
rect 20715 1035 20745 1045
rect 20770 1165 20840 1175
rect 20770 1145 20775 1165
rect 20795 1145 20815 1165
rect 20835 1145 20840 1165
rect 20770 1115 20840 1145
rect 20770 1095 20775 1115
rect 20795 1095 20815 1115
rect 20835 1095 20840 1115
rect 20770 1065 20840 1095
rect 20770 1045 20775 1065
rect 20795 1045 20815 1065
rect 20835 1045 20840 1065
rect 20770 1035 20840 1045
rect 20515 1015 20535 1035
rect 20720 1015 20740 1035
rect 20815 1015 20835 1035
rect 20085 990 20090 1010
rect 20110 990 20130 1010
rect 20150 990 20155 1010
rect 20085 980 20155 990
rect 20505 1005 20545 1015
rect 20505 985 20515 1005
rect 20535 985 20545 1005
rect 12585 940 12590 960
rect 12610 940 12630 960
rect 12650 940 12655 960
rect 12585 930 12655 940
rect 12885 965 12925 975
rect 12885 945 12895 965
rect 12915 945 12925 965
rect 12885 935 12925 945
rect 13125 965 13165 975
rect 13125 945 13135 965
rect 13155 945 13165 965
rect 13125 935 13165 945
rect 13325 965 13365 975
rect 13325 945 13335 965
rect 13355 945 13365 965
rect 13325 935 13365 945
rect 13525 965 13565 975
rect 13525 945 13535 965
rect 13555 945 13565 965
rect 13525 935 13565 945
rect 13725 965 13765 975
rect 13725 945 13735 965
rect 13755 945 13765 965
rect 13725 935 13765 945
rect 13925 965 13965 975
rect 13925 945 13935 965
rect 13955 945 13965 965
rect 13925 935 13965 945
rect 14165 965 14205 975
rect 14165 945 14175 965
rect 14195 945 14205 965
rect 18675 960 18695 980
rect 18770 960 18790 980
rect 18880 960 18900 980
rect 18990 960 19010 980
rect 19100 960 19120 980
rect 19210 960 19230 980
rect 19320 960 19340 980
rect 19430 960 19450 980
rect 19540 960 19560 980
rect 19650 960 19670 980
rect 19760 960 19780 980
rect 19870 960 19890 980
rect 19980 960 20000 980
rect 20130 960 20150 980
rect 20505 975 20545 985
rect 20685 1005 20740 1015
rect 20685 985 20695 1005
rect 20715 995 20740 1005
rect 20805 1005 20845 1015
rect 20715 985 20725 995
rect 20685 975 20725 985
rect 20805 985 20815 1005
rect 20835 985 20845 1005
rect 20805 975 20845 985
rect 14165 935 14205 945
rect 18665 950 18705 960
rect 18665 930 18675 950
rect 18695 930 18705 950
rect 4975 905 4985 925
rect 5005 905 5015 925
rect 11175 910 11195 930
rect 11270 910 11290 930
rect 11380 910 11400 930
rect 11490 910 11510 930
rect 11600 910 11620 930
rect 11710 910 11730 930
rect 11820 910 11840 930
rect 11930 910 11950 930
rect 12040 910 12060 930
rect 12150 910 12170 930
rect 12260 910 12280 930
rect 12370 910 12390 930
rect 12480 910 12500 930
rect 12630 910 12650 930
rect 18665 920 18705 930
rect 18760 950 18800 960
rect 18760 930 18770 950
rect 18790 930 18800 950
rect 18760 920 18800 930
rect 18870 950 18910 960
rect 18870 930 18880 950
rect 18900 930 18910 950
rect 18870 920 18910 930
rect 18980 950 19020 960
rect 18980 930 18990 950
rect 19010 930 19020 950
rect 18980 920 19020 930
rect 19090 950 19130 960
rect 19090 930 19100 950
rect 19120 930 19130 950
rect 19090 920 19130 930
rect 19200 950 19240 960
rect 19200 930 19210 950
rect 19230 930 19240 950
rect 19200 920 19240 930
rect 19310 950 19350 960
rect 19310 930 19320 950
rect 19340 930 19350 950
rect 19310 920 19350 930
rect 19420 950 19460 960
rect 19420 930 19430 950
rect 19450 930 19460 950
rect 19420 920 19460 930
rect 19530 950 19570 960
rect 19530 930 19540 950
rect 19560 930 19570 950
rect 19530 920 19570 930
rect 19640 950 19680 960
rect 19640 930 19650 950
rect 19670 930 19680 950
rect 19640 920 19680 930
rect 19750 950 19790 960
rect 19750 930 19760 950
rect 19780 930 19790 950
rect 19750 920 19790 930
rect 19860 950 19900 960
rect 19860 930 19870 950
rect 19890 930 19900 950
rect 19860 920 19900 930
rect 19970 950 20010 960
rect 19970 930 19980 950
rect 20000 930 20010 950
rect 19970 920 20010 930
rect 20120 950 20160 960
rect 20120 930 20130 950
rect 20150 930 20160 950
rect 20120 920 20160 930
rect 4975 895 5015 905
rect 11165 900 11205 910
rect 3005 875 3025 895
rect 3185 875 3205 895
rect 3365 875 3385 895
rect 3545 875 3565 895
rect 3725 875 3745 895
rect 3905 875 3925 895
rect 4085 875 4105 895
rect 4265 875 4285 895
rect 4445 875 4465 895
rect 4625 875 4645 895
rect 4805 875 4825 895
rect 4985 875 5005 895
rect 11165 880 11175 900
rect 11195 880 11205 900
rect 2960 865 3030 875
rect 2960 845 2965 865
rect 2985 845 3005 865
rect 3025 845 3030 865
rect 2960 815 3030 845
rect 2960 795 2965 815
rect 2985 795 3005 815
rect 3025 795 3030 815
rect 2960 785 3030 795
rect 3090 865 3120 875
rect 3090 845 3095 865
rect 3115 845 3120 865
rect 3090 815 3120 845
rect 3090 795 3095 815
rect 3115 795 3120 815
rect 3090 785 3120 795
rect 3180 865 3210 875
rect 3180 845 3185 865
rect 3205 845 3210 865
rect 3180 815 3210 845
rect 3180 795 3185 815
rect 3205 795 3210 815
rect 3180 785 3210 795
rect 3270 865 3300 875
rect 3270 845 3275 865
rect 3295 845 3300 865
rect 3270 815 3300 845
rect 3270 795 3275 815
rect 3295 795 3300 815
rect 3270 785 3300 795
rect 3360 865 3390 875
rect 3360 845 3365 865
rect 3385 845 3390 865
rect 3360 815 3390 845
rect 3360 795 3365 815
rect 3385 795 3390 815
rect 3360 785 3390 795
rect 3450 865 3480 875
rect 3450 845 3455 865
rect 3475 845 3480 865
rect 3450 815 3480 845
rect 3450 795 3455 815
rect 3475 795 3480 815
rect 3450 785 3480 795
rect 3540 865 3570 875
rect 3540 845 3545 865
rect 3565 845 3570 865
rect 3540 815 3570 845
rect 3540 795 3545 815
rect 3565 795 3570 815
rect 3540 785 3570 795
rect 3630 865 3660 875
rect 3630 845 3635 865
rect 3655 845 3660 865
rect 3630 815 3660 845
rect 3630 795 3635 815
rect 3655 795 3660 815
rect 3630 785 3660 795
rect 3720 865 3750 875
rect 3720 845 3725 865
rect 3745 845 3750 865
rect 3720 815 3750 845
rect 3720 795 3725 815
rect 3745 795 3750 815
rect 3720 785 3750 795
rect 3810 865 3840 875
rect 3810 845 3815 865
rect 3835 845 3840 865
rect 3810 815 3840 845
rect 3810 795 3815 815
rect 3835 795 3840 815
rect 3810 785 3840 795
rect 3900 865 3930 875
rect 3900 845 3905 865
rect 3925 845 3930 865
rect 3900 815 3930 845
rect 3900 795 3905 815
rect 3925 795 3930 815
rect 3900 785 3930 795
rect 3990 865 4020 875
rect 3990 845 3995 865
rect 4015 845 4020 865
rect 3990 815 4020 845
rect 3990 795 3995 815
rect 4015 795 4020 815
rect 3990 785 4020 795
rect 4080 865 4110 875
rect 4080 845 4085 865
rect 4105 845 4110 865
rect 4080 815 4110 845
rect 4080 795 4085 815
rect 4105 795 4110 815
rect 4080 785 4110 795
rect 4170 865 4200 875
rect 4170 845 4175 865
rect 4195 845 4200 865
rect 4170 815 4200 845
rect 4170 795 4175 815
rect 4195 795 4200 815
rect 4170 785 4200 795
rect 4260 865 4290 875
rect 4260 845 4265 865
rect 4285 845 4290 865
rect 4260 815 4290 845
rect 4260 795 4265 815
rect 4285 795 4290 815
rect 4260 785 4290 795
rect 4350 865 4380 875
rect 4350 845 4355 865
rect 4375 845 4380 865
rect 4350 815 4380 845
rect 4350 795 4355 815
rect 4375 795 4380 815
rect 4350 785 4380 795
rect 4440 865 4470 875
rect 4440 845 4445 865
rect 4465 845 4470 865
rect 4440 815 4470 845
rect 4440 795 4445 815
rect 4465 795 4470 815
rect 4440 785 4470 795
rect 4530 865 4560 875
rect 4530 845 4535 865
rect 4555 845 4560 865
rect 4530 815 4560 845
rect 4530 795 4535 815
rect 4555 795 4560 815
rect 4530 785 4560 795
rect 4620 865 4650 875
rect 4620 845 4625 865
rect 4645 845 4650 865
rect 4620 815 4650 845
rect 4620 795 4625 815
rect 4645 795 4650 815
rect 4620 785 4650 795
rect 4710 865 4740 875
rect 4710 845 4715 865
rect 4735 845 4740 865
rect 4710 815 4740 845
rect 4710 795 4715 815
rect 4735 795 4740 815
rect 4710 785 4740 795
rect 4800 865 4830 875
rect 4800 845 4805 865
rect 4825 845 4830 865
rect 4800 815 4830 845
rect 4800 795 4805 815
rect 4825 795 4830 815
rect 4800 785 4830 795
rect 4890 865 4920 875
rect 4890 845 4895 865
rect 4915 845 4920 865
rect 4890 815 4920 845
rect 4890 795 4895 815
rect 4915 795 4920 815
rect 4890 785 4920 795
rect 4980 865 5050 875
rect 11165 870 11205 880
rect 11260 900 11300 910
rect 11260 880 11270 900
rect 11290 880 11300 900
rect 11260 870 11300 880
rect 11370 900 11410 910
rect 11370 880 11380 900
rect 11400 880 11410 900
rect 11370 870 11410 880
rect 11480 900 11520 910
rect 11480 880 11490 900
rect 11510 880 11520 900
rect 11480 870 11520 880
rect 11590 900 11630 910
rect 11590 880 11600 900
rect 11620 880 11630 900
rect 11590 870 11630 880
rect 11700 900 11740 910
rect 11700 880 11710 900
rect 11730 880 11740 900
rect 11700 870 11740 880
rect 11810 900 11850 910
rect 11810 880 11820 900
rect 11840 880 11850 900
rect 11810 870 11850 880
rect 11920 900 11960 910
rect 11920 880 11930 900
rect 11950 880 11960 900
rect 11920 870 11960 880
rect 12030 900 12070 910
rect 12030 880 12040 900
rect 12060 880 12070 900
rect 12030 870 12070 880
rect 12140 900 12180 910
rect 12140 880 12150 900
rect 12170 880 12180 900
rect 12140 870 12180 880
rect 12250 900 12290 910
rect 12250 880 12260 900
rect 12280 880 12290 900
rect 12250 870 12290 880
rect 12360 900 12400 910
rect 12360 880 12370 900
rect 12390 880 12400 900
rect 12360 870 12400 880
rect 12470 900 12510 910
rect 12470 880 12480 900
rect 12500 880 12510 900
rect 12470 870 12510 880
rect 12620 900 12660 910
rect 12620 880 12630 900
rect 12650 880 12660 900
rect 12620 870 12660 880
rect 4980 845 4985 865
rect 5005 845 5025 865
rect 5045 845 5050 865
rect 4980 815 5050 845
rect 4980 795 4985 815
rect 5005 795 5025 815
rect 5045 795 5050 815
rect 4980 785 5050 795
rect 3095 765 3115 785
rect 3275 765 3295 785
rect 3455 765 3475 785
rect 3635 765 3655 785
rect 3815 765 3835 785
rect 3995 765 4015 785
rect 4175 765 4195 785
rect 4355 765 4375 785
rect 4535 765 4555 785
rect 4715 765 4735 785
rect 4895 765 4915 785
rect 2525 730 2555 760
rect 3095 755 3170 765
rect 3095 745 3140 755
rect 3130 735 3140 745
rect 3160 735 3170 755
rect 3130 725 3170 735
rect 3265 755 3305 765
rect 3265 735 3275 755
rect 3295 735 3305 755
rect 3265 725 3305 735
rect 3445 755 3485 765
rect 3445 735 3455 755
rect 3475 735 3485 755
rect 3445 725 3485 735
rect 3625 755 3665 765
rect 3625 735 3635 755
rect 3655 735 3665 755
rect 3625 725 3665 735
rect 3805 755 3845 765
rect 3805 735 3815 755
rect 3835 735 3845 755
rect 3805 725 3845 735
rect 3985 755 4025 765
rect 3985 735 3995 755
rect 4015 735 4025 755
rect 3985 725 4025 735
rect 4165 755 4205 765
rect 4165 735 4175 755
rect 4195 735 4205 755
rect 4165 725 4205 735
rect 4345 755 4385 765
rect 4345 735 4355 755
rect 4375 735 4385 755
rect 4345 725 4385 735
rect 4525 755 4565 765
rect 4525 735 4535 755
rect 4555 735 4565 755
rect 4525 725 4565 735
rect 4705 755 4745 765
rect 4705 735 4715 755
rect 4735 735 4745 755
rect 4705 725 4745 735
rect 4885 755 4925 765
rect 4885 735 4895 755
rect 4915 735 4925 755
rect 4885 725 4925 735
rect 3450 675 3480 705
rect 3810 675 3840 705
rect 4170 675 4200 705
rect 9375 -685 9415 -675
rect 9375 -705 9385 -685
rect 9405 -705 9415 -685
rect 9375 -715 9415 -705
rect 9575 -685 9615 -675
rect 9575 -705 9585 -685
rect 9605 -705 9615 -685
rect 9575 -715 9615 -705
rect 9775 -685 9815 -675
rect 9775 -705 9785 -685
rect 9805 -705 9815 -685
rect 9775 -715 9815 -705
rect 9975 -685 10015 -675
rect 9975 -705 9985 -685
rect 10005 -705 10015 -685
rect 9975 -715 10015 -705
rect 10175 -685 10215 -675
rect 10175 -705 10185 -685
rect 10205 -705 10215 -685
rect 10175 -715 10215 -705
rect 10375 -685 10415 -675
rect 10375 -705 10385 -685
rect 10405 -705 10415 -685
rect 10375 -715 10415 -705
rect 9385 -735 9405 -715
rect 9585 -735 9605 -715
rect 9785 -735 9805 -715
rect 9985 -735 10005 -715
rect 10185 -735 10205 -715
rect 10385 -735 10405 -715
rect 9240 -745 9310 -735
rect 9240 -765 9245 -745
rect 9265 -765 9285 -745
rect 9305 -765 9310 -745
rect 9240 -790 9310 -765
rect 9240 -810 9245 -790
rect 9265 -810 9285 -790
rect 9305 -810 9310 -790
rect 9240 -835 9310 -810
rect 9240 -855 9245 -835
rect 9265 -855 9285 -835
rect 9305 -855 9310 -835
rect 9240 -885 9310 -855
rect 9240 -905 9245 -885
rect 9265 -905 9285 -885
rect 9305 -905 9310 -885
rect 9240 -930 9310 -905
rect 9240 -950 9245 -930
rect 9265 -950 9285 -930
rect 9305 -950 9310 -930
rect 9240 -975 9310 -950
rect 9240 -995 9245 -975
rect 9265 -995 9285 -975
rect 9305 -995 9310 -975
rect 9240 -1005 9310 -995
rect 9380 -745 9410 -735
rect 9380 -765 9385 -745
rect 9405 -765 9410 -745
rect 9380 -790 9410 -765
rect 9380 -810 9385 -790
rect 9405 -810 9410 -790
rect 9380 -835 9410 -810
rect 9380 -855 9385 -835
rect 9405 -855 9410 -835
rect 9380 -885 9410 -855
rect 9380 -905 9385 -885
rect 9405 -905 9410 -885
rect 9380 -930 9410 -905
rect 9380 -950 9385 -930
rect 9405 -950 9410 -930
rect 9380 -975 9410 -950
rect 9380 -995 9385 -975
rect 9405 -995 9410 -975
rect 9380 -1005 9410 -995
rect 9480 -745 9510 -735
rect 9480 -765 9485 -745
rect 9505 -765 9510 -745
rect 9480 -790 9510 -765
rect 9480 -810 9485 -790
rect 9505 -810 9510 -790
rect 9480 -835 9510 -810
rect 9480 -855 9485 -835
rect 9505 -855 9510 -835
rect 9480 -885 9510 -855
rect 9480 -905 9485 -885
rect 9505 -905 9510 -885
rect 9480 -930 9510 -905
rect 9480 -950 9485 -930
rect 9505 -950 9510 -930
rect 9480 -975 9510 -950
rect 9480 -995 9485 -975
rect 9505 -995 9510 -975
rect 9480 -1005 9510 -995
rect 9580 -745 9610 -735
rect 9580 -765 9585 -745
rect 9605 -765 9610 -745
rect 9580 -790 9610 -765
rect 9580 -810 9585 -790
rect 9605 -810 9610 -790
rect 9580 -835 9610 -810
rect 9580 -855 9585 -835
rect 9605 -855 9610 -835
rect 9580 -885 9610 -855
rect 9580 -905 9585 -885
rect 9605 -905 9610 -885
rect 9580 -930 9610 -905
rect 9580 -950 9585 -930
rect 9605 -950 9610 -930
rect 9580 -975 9610 -950
rect 9580 -995 9585 -975
rect 9605 -995 9610 -975
rect 9580 -1005 9610 -995
rect 9680 -745 9710 -735
rect 9680 -765 9685 -745
rect 9705 -765 9710 -745
rect 9680 -790 9710 -765
rect 9680 -810 9685 -790
rect 9705 -810 9710 -790
rect 9680 -835 9710 -810
rect 9680 -855 9685 -835
rect 9705 -855 9710 -835
rect 9680 -885 9710 -855
rect 9680 -905 9685 -885
rect 9705 -905 9710 -885
rect 9680 -930 9710 -905
rect 9680 -950 9685 -930
rect 9705 -950 9710 -930
rect 9680 -975 9710 -950
rect 9680 -995 9685 -975
rect 9705 -995 9710 -975
rect 9680 -1005 9710 -995
rect 9780 -745 9810 -735
rect 9780 -765 9785 -745
rect 9805 -765 9810 -745
rect 9780 -790 9810 -765
rect 9780 -810 9785 -790
rect 9805 -810 9810 -790
rect 9780 -835 9810 -810
rect 9780 -855 9785 -835
rect 9805 -855 9810 -835
rect 9780 -885 9810 -855
rect 9780 -905 9785 -885
rect 9805 -905 9810 -885
rect 9780 -930 9810 -905
rect 9780 -950 9785 -930
rect 9805 -950 9810 -930
rect 9780 -975 9810 -950
rect 9780 -995 9785 -975
rect 9805 -995 9810 -975
rect 9780 -1005 9810 -995
rect 9880 -745 9910 -735
rect 9880 -765 9885 -745
rect 9905 -765 9910 -745
rect 9880 -790 9910 -765
rect 9880 -810 9885 -790
rect 9905 -810 9910 -790
rect 9880 -835 9910 -810
rect 9880 -855 9885 -835
rect 9905 -855 9910 -835
rect 9880 -885 9910 -855
rect 9880 -905 9885 -885
rect 9905 -905 9910 -885
rect 9880 -930 9910 -905
rect 9880 -950 9885 -930
rect 9905 -950 9910 -930
rect 9880 -975 9910 -950
rect 9880 -995 9885 -975
rect 9905 -995 9910 -975
rect 9880 -1005 9910 -995
rect 9980 -745 10010 -735
rect 9980 -765 9985 -745
rect 10005 -765 10010 -745
rect 9980 -790 10010 -765
rect 9980 -810 9985 -790
rect 10005 -810 10010 -790
rect 9980 -835 10010 -810
rect 9980 -855 9985 -835
rect 10005 -855 10010 -835
rect 9980 -885 10010 -855
rect 9980 -905 9985 -885
rect 10005 -905 10010 -885
rect 9980 -930 10010 -905
rect 9980 -950 9985 -930
rect 10005 -950 10010 -930
rect 9980 -975 10010 -950
rect 9980 -995 9985 -975
rect 10005 -995 10010 -975
rect 9980 -1005 10010 -995
rect 10080 -745 10110 -735
rect 10080 -765 10085 -745
rect 10105 -765 10110 -745
rect 10080 -790 10110 -765
rect 10080 -810 10085 -790
rect 10105 -810 10110 -790
rect 10080 -835 10110 -810
rect 10080 -855 10085 -835
rect 10105 -855 10110 -835
rect 10080 -885 10110 -855
rect 10080 -905 10085 -885
rect 10105 -905 10110 -885
rect 10080 -930 10110 -905
rect 10080 -950 10085 -930
rect 10105 -950 10110 -930
rect 10080 -975 10110 -950
rect 10080 -995 10085 -975
rect 10105 -995 10110 -975
rect 10080 -1005 10110 -995
rect 10180 -745 10210 -735
rect 10180 -765 10185 -745
rect 10205 -765 10210 -745
rect 10180 -790 10210 -765
rect 10180 -810 10185 -790
rect 10205 -810 10210 -790
rect 10180 -835 10210 -810
rect 10180 -855 10185 -835
rect 10205 -855 10210 -835
rect 10180 -885 10210 -855
rect 10180 -905 10185 -885
rect 10205 -905 10210 -885
rect 10180 -930 10210 -905
rect 10180 -950 10185 -930
rect 10205 -950 10210 -930
rect 10180 -975 10210 -950
rect 10180 -995 10185 -975
rect 10205 -995 10210 -975
rect 10180 -1005 10210 -995
rect 10280 -745 10310 -735
rect 10280 -765 10285 -745
rect 10305 -765 10310 -745
rect 10280 -790 10310 -765
rect 10280 -810 10285 -790
rect 10305 -810 10310 -790
rect 10280 -835 10310 -810
rect 10280 -855 10285 -835
rect 10305 -855 10310 -835
rect 10280 -885 10310 -855
rect 10280 -905 10285 -885
rect 10305 -905 10310 -885
rect 10280 -930 10310 -905
rect 10280 -950 10285 -930
rect 10305 -950 10310 -930
rect 10280 -975 10310 -950
rect 10280 -995 10285 -975
rect 10305 -995 10310 -975
rect 10280 -1005 10310 -995
rect 10380 -745 10410 -735
rect 10380 -765 10385 -745
rect 10405 -765 10410 -745
rect 10380 -790 10410 -765
rect 10380 -810 10385 -790
rect 10405 -810 10410 -790
rect 10380 -835 10410 -810
rect 10380 -855 10385 -835
rect 10405 -855 10410 -835
rect 10380 -885 10410 -855
rect 10380 -905 10385 -885
rect 10405 -905 10410 -885
rect 10380 -930 10410 -905
rect 10380 -950 10385 -930
rect 10405 -950 10410 -930
rect 10380 -975 10410 -950
rect 10380 -995 10385 -975
rect 10405 -995 10410 -975
rect 10380 -1005 10410 -995
rect 10480 -745 10550 -735
rect 10480 -765 10485 -745
rect 10505 -765 10525 -745
rect 10545 -765 10550 -745
rect 10480 -790 10550 -765
rect 10480 -810 10485 -790
rect 10505 -810 10525 -790
rect 10545 -810 10550 -790
rect 10480 -835 10550 -810
rect 10480 -855 10485 -835
rect 10505 -855 10525 -835
rect 10545 -855 10550 -835
rect 10480 -885 10550 -855
rect 10480 -905 10485 -885
rect 10505 -905 10525 -885
rect 10545 -905 10550 -885
rect 10480 -930 10550 -905
rect 10480 -950 10485 -930
rect 10505 -950 10525 -930
rect 10545 -950 10550 -930
rect 10480 -975 10550 -950
rect 10480 -995 10485 -975
rect 10505 -995 10525 -975
rect 10545 -995 10550 -975
rect 10480 -1005 10550 -995
rect 9245 -1025 9265 -1005
rect 9485 -1025 9505 -1005
rect 9685 -1025 9705 -1005
rect 9885 -1025 9905 -1005
rect 10085 -1025 10105 -1005
rect 10285 -1025 10305 -1005
rect 10525 -1025 10545 -1005
rect 9235 -1035 9275 -1025
rect 9235 -1055 9245 -1035
rect 9265 -1055 9275 -1035
rect 9235 -1065 9275 -1055
rect 9475 -1035 9515 -1025
rect 9475 -1055 9485 -1035
rect 9505 -1055 9515 -1035
rect 9475 -1065 9515 -1055
rect 9675 -1035 9715 -1025
rect 9675 -1055 9685 -1035
rect 9705 -1055 9715 -1035
rect 9675 -1065 9715 -1055
rect 9875 -1035 9915 -1025
rect 9875 -1055 9885 -1035
rect 9905 -1055 9915 -1035
rect 9875 -1065 9915 -1055
rect 10075 -1035 10115 -1025
rect 10075 -1055 10085 -1035
rect 10105 -1055 10115 -1035
rect 10075 -1065 10115 -1055
rect 10275 -1035 10315 -1025
rect 10275 -1055 10285 -1035
rect 10305 -1055 10315 -1035
rect 10275 -1065 10315 -1055
rect 10515 -1035 10555 -1025
rect 10515 -1055 10525 -1035
rect 10545 -1055 10555 -1035
rect 10515 -1065 10555 -1055
<< viali >>
rect 11350 3600 11370 3620
rect 11470 3600 11490 3620
rect 11590 3600 11610 3620
rect 11710 3600 11730 3620
rect 11830 3600 11850 3620
rect 11950 3600 11970 3620
rect 12070 3600 12090 3620
rect 12190 3600 12210 3620
rect 12310 3600 12330 3620
rect 12430 3600 12450 3620
rect 18850 3600 18870 3620
rect 18970 3600 18990 3620
rect 19090 3600 19110 3620
rect 19210 3600 19230 3620
rect 19330 3600 19350 3620
rect 19450 3600 19470 3620
rect 19570 3600 19590 3620
rect 19690 3600 19710 3620
rect 19810 3600 19830 3620
rect 19930 3600 19950 3620
rect 56 3175 81 3200
rect 1271 3170 1296 3195
rect 10590 3185 10610 3205
rect 56 3115 81 3140
rect 1271 3110 1296 3135
rect 56 3035 81 3060
rect 56 2975 81 3000
rect 920 2880 950 2910
rect 1000 2880 1030 2910
rect 1080 2880 1110 2910
rect 10910 3185 10930 3205
rect 10990 3185 11010 3205
rect 12955 3265 12975 3285
rect 13065 3265 13085 3285
rect 13175 3265 13195 3285
rect 13285 3265 13305 3285
rect 13395 3265 13415 3285
rect 13505 3265 13525 3285
rect 13615 3265 13635 3285
rect 13725 3265 13745 3285
rect 13835 3265 13855 3285
rect 13945 3265 13965 3285
rect 14055 3265 14075 3285
rect 11290 3130 11310 3150
rect 11410 3130 11430 3150
rect 11530 3130 11550 3150
rect 11650 3130 11670 3150
rect 11770 3130 11790 3150
rect 11831 3130 11849 3150
rect 11890 3130 11910 3150
rect 12010 3130 12030 3150
rect 12130 3130 12150 3150
rect 12250 3130 12270 3150
rect 12370 3130 12390 3150
rect 12490 3130 12510 3150
rect 2340 2930 2365 2955
rect 3090 2955 3110 2975
rect 3145 2955 3165 2975
rect 3275 2955 3295 2975
rect 3455 2955 3475 2975
rect 3635 2955 3655 2975
rect 3815 2955 3835 2975
rect 3995 2955 4015 2975
rect 4175 2955 4195 2975
rect 4355 2955 4375 2975
rect 4535 2955 4555 2975
rect 4715 2955 4735 2975
rect 4845 2955 4865 2975
rect 4895 2955 4915 2975
rect 2340 2870 2365 2895
rect 61 2825 86 2850
rect 734 2825 759 2850
rect 1271 2810 1296 2835
rect 1970 2810 1995 2835
rect 11350 2920 11370 2940
rect 11470 2920 11490 2940
rect 11590 2920 11610 2940
rect 11710 2920 11730 2940
rect 11830 2920 11850 2940
rect 11950 2920 11970 2940
rect 12070 2920 12090 2940
rect 12190 2920 12210 2940
rect 12310 2920 12330 2940
rect 12430 2920 12450 2940
rect 18090 3185 18110 3205
rect 18410 3185 18430 3205
rect 18490 3185 18510 3205
rect 20455 3265 20475 3285
rect 20565 3265 20585 3285
rect 20675 3265 20695 3285
rect 20785 3265 20805 3285
rect 20895 3265 20915 3285
rect 21005 3265 21025 3285
rect 21115 3265 21135 3285
rect 21225 3265 21245 3285
rect 21335 3265 21355 3285
rect 21445 3265 21465 3285
rect 21555 3265 21575 3285
rect 18790 3130 18810 3150
rect 18910 3130 18930 3150
rect 19030 3130 19050 3150
rect 19150 3130 19170 3150
rect 19270 3130 19290 3150
rect 19331 3130 19349 3150
rect 19390 3130 19410 3150
rect 19510 3130 19530 3150
rect 19630 3130 19650 3150
rect 19750 3130 19770 3150
rect 19870 3130 19890 3150
rect 19990 3130 20010 3150
rect 61 2765 86 2790
rect 734 2765 759 2790
rect 3005 2785 3025 2805
rect 3185 2785 3205 2805
rect 3365 2785 3385 2805
rect 3545 2785 3565 2805
rect 3725 2785 3745 2805
rect 3905 2785 3925 2805
rect 4085 2785 4105 2805
rect 4265 2785 4285 2805
rect 4445 2785 4465 2805
rect 4625 2785 4645 2805
rect 4805 2785 4825 2805
rect 4985 2785 5005 2805
rect 3185 2725 3205 2745
rect 3365 2725 3385 2745
rect 3545 2725 3565 2745
rect 3725 2725 3745 2745
rect 3905 2725 3925 2745
rect 4085 2725 4105 2745
rect 4265 2725 4285 2745
rect 4445 2725 4465 2745
rect 4625 2725 4645 2745
rect 4805 2725 4825 2745
rect 9745 2645 9765 2665
rect 9855 2645 9875 2665
rect 9965 2645 9985 2665
rect 10075 2645 10095 2665
rect 10185 2645 10205 2665
rect 10295 2645 10315 2665
rect 10405 2645 10425 2665
rect 10515 2645 10535 2665
rect 10625 2645 10645 2665
rect 10735 2645 10755 2665
rect 10845 2645 10865 2665
rect 9800 2475 9820 2495
rect 9910 2475 9930 2495
rect 10020 2475 10040 2495
rect 10130 2475 10150 2495
rect 10240 2475 10260 2495
rect 10350 2475 10370 2495
rect 10460 2475 10480 2495
rect 10570 2475 10590 2495
rect 10680 2475 10700 2495
rect 10790 2475 10810 2495
rect 13010 2895 13030 2915
rect 13066 2895 13084 2915
rect 13120 2895 13140 2915
rect 13230 2895 13250 2915
rect 13340 2895 13360 2915
rect 13450 2895 13470 2915
rect 13560 2895 13580 2915
rect 13670 2895 13690 2915
rect 13780 2895 13800 2915
rect 13890 2895 13910 2915
rect 14000 2895 14020 2915
rect 18850 2920 18870 2940
rect 18970 2920 18990 2940
rect 19090 2920 19110 2940
rect 19210 2920 19230 2940
rect 19330 2920 19350 2940
rect 19450 2920 19470 2940
rect 19570 2920 19590 2940
rect 19690 2920 19710 2940
rect 19810 2920 19830 2940
rect 19930 2920 19950 2940
rect 12955 2645 12975 2665
rect 13065 2645 13085 2665
rect 13175 2645 13195 2665
rect 13285 2645 13305 2665
rect 13395 2645 13415 2665
rect 13505 2645 13525 2665
rect 13615 2645 13635 2665
rect 13725 2645 13745 2665
rect 13835 2645 13855 2665
rect 13945 2645 13965 2665
rect 14055 2645 14075 2665
rect 17245 2645 17265 2665
rect 17355 2645 17375 2665
rect 17465 2645 17485 2665
rect 17575 2645 17595 2665
rect 17685 2645 17705 2665
rect 17795 2645 17815 2665
rect 17905 2645 17925 2665
rect 18015 2645 18035 2665
rect 18125 2645 18145 2665
rect 18235 2645 18255 2665
rect 18345 2645 18365 2665
rect 11290 2450 11310 2470
rect 11410 2450 11430 2470
rect 11530 2450 11550 2470
rect 11650 2450 11670 2470
rect 11770 2450 11790 2470
rect 11831 2450 11849 2470
rect 11890 2450 11910 2470
rect 12010 2450 12030 2470
rect 12130 2450 12150 2470
rect 12250 2450 12270 2470
rect 12370 2450 12390 2470
rect 12490 2450 12510 2470
rect 13010 2475 13030 2495
rect 13120 2475 13140 2495
rect 13230 2475 13250 2495
rect 13340 2475 13360 2495
rect 13450 2475 13470 2495
rect 13560 2475 13580 2495
rect 13670 2475 13690 2495
rect 13780 2475 13800 2495
rect 13890 2475 13910 2495
rect 14000 2475 14020 2495
rect 17300 2475 17320 2495
rect 17410 2475 17430 2495
rect 17520 2475 17540 2495
rect 17630 2475 17650 2495
rect 17740 2475 17760 2495
rect 17850 2475 17870 2495
rect 17960 2475 17980 2495
rect 18070 2475 18090 2495
rect 18180 2475 18200 2495
rect 18290 2475 18310 2495
rect 20510 2895 20530 2915
rect 20566 2895 20584 2915
rect 20620 2895 20640 2915
rect 20730 2895 20750 2915
rect 20840 2895 20860 2915
rect 20950 2895 20970 2915
rect 21060 2895 21080 2915
rect 21170 2895 21190 2915
rect 21280 2895 21300 2915
rect 21390 2895 21410 2915
rect 21500 2895 21520 2915
rect 20455 2645 20475 2665
rect 20565 2645 20585 2665
rect 20675 2645 20695 2665
rect 20785 2645 20805 2665
rect 20895 2645 20915 2665
rect 21005 2645 21025 2665
rect 21115 2645 21135 2665
rect 21225 2645 21245 2665
rect 21335 2645 21355 2665
rect 21445 2645 21465 2665
rect 21555 2645 21575 2665
rect 18790 2450 18810 2470
rect 10821 2415 10839 2435
rect 12981 2415 12999 2435
rect 18910 2450 18930 2470
rect 19030 2450 19050 2470
rect 19150 2450 19170 2470
rect 19270 2450 19290 2470
rect 19331 2450 19349 2470
rect 19390 2450 19410 2470
rect 19510 2450 19530 2470
rect 19630 2450 19650 2470
rect 19750 2450 19770 2470
rect 19870 2450 19890 2470
rect 19990 2450 20010 2470
rect 20510 2475 20530 2495
rect 20620 2475 20640 2495
rect 20730 2475 20750 2495
rect 20840 2475 20860 2495
rect 20950 2475 20970 2495
rect 21060 2475 21080 2495
rect 21170 2475 21190 2495
rect 21280 2475 21300 2495
rect 21390 2475 21410 2495
rect 21500 2475 21520 2495
rect 18321 2415 18339 2435
rect 20481 2415 20499 2435
rect 3275 2355 3295 2375
rect 3365 2350 3385 2370
rect 3455 2355 3475 2375
rect 3815 2355 3835 2375
rect 3895 2355 3915 2375
rect 3995 2355 4015 2375
rect 4175 2355 4195 2375
rect 4535 2355 4555 2375
rect 4715 2355 4735 2375
rect 9810 2350 9835 2375
rect 10645 2350 10670 2375
rect 13150 2350 13175 2375
rect 13985 2350 14010 2375
rect 17310 2350 17335 2375
rect 18145 2350 18170 2375
rect 20650 2350 20675 2375
rect 21485 2350 21510 2375
rect 3635 2310 3655 2330
rect 4355 2310 4375 2330
rect 3455 2265 3475 2285
rect 9810 2290 9835 2315
rect 4535 2265 4555 2285
rect 10645 2290 10670 2315
rect 13150 2290 13175 2315
rect 13985 2290 14010 2315
rect 17310 2290 17335 2315
rect 18145 2290 18170 2315
rect 20650 2290 20675 2315
rect 21485 2290 21510 2315
rect 10821 2255 10839 2275
rect 12981 2255 12999 2275
rect 18321 2255 18339 2275
rect 20481 2255 20499 2275
rect 9800 2195 9820 2215
rect 9910 2195 9930 2215
rect 10020 2195 10040 2215
rect 10130 2195 10150 2215
rect 10240 2195 10260 2215
rect 10350 2195 10370 2215
rect 10460 2195 10480 2215
rect 10570 2195 10590 2215
rect 10680 2195 10700 2215
rect 10790 2195 10810 2215
rect 13010 2195 13030 2215
rect 13120 2195 13140 2215
rect 13230 2195 13250 2215
rect 13340 2195 13360 2215
rect 13450 2195 13470 2215
rect 13560 2195 13580 2215
rect 13670 2195 13690 2215
rect 13780 2195 13800 2215
rect 13890 2195 13910 2215
rect 14000 2195 14020 2215
rect 17300 2195 17320 2215
rect 17410 2195 17430 2215
rect 17520 2195 17540 2215
rect 17630 2195 17650 2215
rect 17740 2195 17760 2215
rect 17850 2195 17870 2215
rect 17960 2195 17980 2215
rect 18070 2195 18090 2215
rect 18180 2195 18200 2215
rect 18290 2195 18310 2215
rect 20510 2195 20530 2215
rect 20620 2195 20640 2215
rect 20730 2195 20750 2215
rect 20840 2195 20860 2215
rect 20950 2195 20970 2215
rect 21060 2195 21080 2215
rect 21170 2195 21190 2215
rect 21280 2195 21300 2215
rect 21390 2195 21410 2215
rect 21500 2195 21520 2215
rect 2755 2070 2775 2090
rect 2875 2070 2895 2090
rect 2995 2070 3015 2090
rect 3115 2070 3135 2090
rect 3235 2070 3255 2090
rect 3355 2070 3375 2090
rect 3475 2070 3495 2090
rect 3595 2070 3615 2090
rect 3715 2070 3735 2090
rect 3835 2070 3855 2090
rect 3995 2070 4015 2090
rect 4155 2070 4175 2090
rect 4275 2070 4295 2090
rect 4395 2070 4415 2090
rect 4515 2070 4535 2090
rect 4635 2070 4655 2090
rect 4755 2070 4775 2090
rect 4875 2070 4895 2090
rect 4995 2070 5015 2090
rect 5115 2070 5135 2090
rect 5235 2070 5255 2090
rect 2630 2025 2650 2045
rect -35 1695 -15 1715
rect 2815 2025 2835 2045
rect 3175 2025 3195 2045
rect 3535 2025 3555 2045
rect 3895 2025 3915 2045
rect 4095 2025 4115 2045
rect 4455 2025 4475 2045
rect 4815 2025 4835 2045
rect 5175 2025 5195 2045
rect 11340 2155 11360 2175
rect 11450 2155 11470 2175
rect 11560 2155 11580 2175
rect 11670 2155 11690 2175
rect 11780 2155 11800 2175
rect 11890 2155 11910 2175
rect 12000 2155 12020 2175
rect 12110 2155 12130 2175
rect 12220 2155 12240 2175
rect 12330 2155 12350 2175
rect 12440 2155 12460 2175
rect 9745 1975 9763 1995
rect 9855 1975 9873 1995
rect 9965 1975 9983 1995
rect 10075 1975 10093 1995
rect 10185 1975 10203 1995
rect 10295 1975 10313 1995
rect 10405 1975 10423 1995
rect 10515 1975 10533 1995
rect 10625 1975 10643 1995
rect 10735 1975 10753 1995
rect 10845 1975 10863 1995
rect 18840 2155 18860 2175
rect 18950 2155 18970 2175
rect 19060 2155 19080 2175
rect 19170 2155 19190 2175
rect 19280 2155 19300 2175
rect 19390 2155 19410 2175
rect 19500 2155 19520 2175
rect 19610 2155 19630 2175
rect 19720 2155 19740 2175
rect 19830 2155 19850 2175
rect 19940 2155 19960 2175
rect 12957 1975 12975 1995
rect 13067 1975 13085 1995
rect 13177 1975 13195 1995
rect 13287 1975 13305 1995
rect 13397 1975 13415 1995
rect 13507 1975 13525 1995
rect 13617 1975 13635 1995
rect 13727 1975 13745 1995
rect 13837 1975 13855 1995
rect 13947 1975 13965 1995
rect 14057 1975 14075 1995
rect 17245 1975 17263 1995
rect 17355 1975 17373 1995
rect 17465 1975 17483 1995
rect 17575 1975 17593 1995
rect 17685 1975 17703 1995
rect 17795 1975 17813 1995
rect 17905 1975 17923 1995
rect 18015 1975 18033 1995
rect 18125 1975 18143 1995
rect 18235 1975 18253 1995
rect 18345 1975 18363 1995
rect 20457 1975 20475 1995
rect 20567 1975 20585 1995
rect 20677 1975 20695 1995
rect 20787 1975 20805 1995
rect 20897 1975 20915 1995
rect 21007 1975 21025 1995
rect 21117 1975 21135 1995
rect 21227 1975 21245 1995
rect 21337 1975 21355 1995
rect 21447 1975 21465 1995
rect 21557 1975 21575 1995
rect 11395 1935 11415 1955
rect 11505 1935 11525 1955
rect 11615 1935 11635 1955
rect 11725 1935 11745 1955
rect 11835 1935 11855 1955
rect 11945 1935 11965 1955
rect 12055 1935 12075 1955
rect 12165 1935 12185 1955
rect 12275 1935 12295 1955
rect 12385 1935 12405 1955
rect 18895 1935 18915 1955
rect 19005 1935 19025 1955
rect 19115 1935 19135 1955
rect 19225 1935 19245 1955
rect 19335 1935 19355 1955
rect 19445 1935 19465 1955
rect 19555 1935 19575 1955
rect 19665 1935 19685 1955
rect 19775 1935 19795 1955
rect 19885 1935 19905 1955
rect 2575 1855 2595 1875
rect 2630 1855 2650 1875
rect 2685 1855 2705 1875
rect 2845 1855 2865 1875
rect 2935 1855 2955 1875
rect 3055 1855 3075 1875
rect 3175 1855 3195 1875
rect 3295 1855 3315 1875
rect 3415 1855 3435 1875
rect 3535 1855 3555 1875
rect 3655 1855 3675 1875
rect 3775 1855 3795 1875
rect 3865 1855 3885 1875
rect 4125 1855 4145 1875
rect 4215 1855 4235 1875
rect 4335 1855 4355 1875
rect 4455 1855 4475 1875
rect 4575 1855 4595 1875
rect 4695 1855 4715 1875
rect 4815 1855 4835 1875
rect 4935 1855 4955 1875
rect 5055 1855 5075 1875
rect 5145 1855 5165 1875
rect 20555 1880 20575 1900
rect 20665 1880 20685 1900
rect 20775 1880 20795 1900
rect 3055 1795 3075 1815
rect 3415 1795 3435 1815
rect 3775 1795 3795 1815
rect 4215 1795 4235 1815
rect 4575 1795 4595 1815
rect 4935 1795 4955 1815
rect 3235 1735 3255 1755
rect 3295 1735 3315 1755
rect 3535 1735 3555 1755
rect 3775 1735 3795 1755
rect 4215 1735 4235 1755
rect 4455 1735 4475 1755
rect 4695 1735 4715 1755
rect 4755 1735 4775 1755
rect 11095 1735 11115 1755
rect 11200 1750 11220 1770
rect 3175 1690 3195 1710
rect 3415 1690 3435 1710
rect 3655 1690 3675 1710
rect 4335 1690 4355 1710
rect 4575 1690 4595 1710
rect 4815 1690 4835 1710
rect 11315 1735 11335 1755
rect 11420 1750 11440 1770
rect 11243 1690 11260 1710
rect 11535 1735 11555 1755
rect 11650 1750 11670 1770
rect 11463 1690 11480 1710
rect 11610 1690 11627 1710
rect 12135 1735 12155 1755
rect 12240 1750 12260 1770
rect 11825 1690 11845 1710
rect 11876 1690 11893 1710
rect 11955 1690 11975 1710
rect 12355 1735 12375 1755
rect 12460 1750 12480 1770
rect 12283 1690 12300 1710
rect 12575 1735 12595 1755
rect 12690 1750 12710 1770
rect 12503 1690 12520 1710
rect 12650 1690 12667 1710
rect 18595 1735 18615 1755
rect 18700 1750 18720 1770
rect 18815 1735 18835 1755
rect 18920 1750 18940 1770
rect 18743 1690 18760 1710
rect 19035 1735 19055 1755
rect 19150 1750 19170 1770
rect 18963 1690 18980 1710
rect 19110 1690 19127 1710
rect 19635 1735 19655 1755
rect 19740 1750 19760 1770
rect 19325 1690 19345 1710
rect 19376 1690 19393 1710
rect 19455 1690 19475 1710
rect 19855 1735 19875 1755
rect 19960 1750 19980 1770
rect 19783 1690 19800 1710
rect 20075 1735 20095 1755
rect 20190 1750 20210 1770
rect 20003 1690 20020 1710
rect 20150 1690 20167 1710
rect 3995 1630 4015 1650
rect 3175 1570 3195 1590
rect 4815 1570 4835 1590
rect 3235 1520 3255 1540
rect 3355 1520 3375 1540
rect 3475 1520 3495 1540
rect 3595 1520 3615 1540
rect 3715 1520 3735 1540
rect 4275 1520 4295 1540
rect 4395 1520 4415 1540
rect 4515 1520 4535 1540
rect 4635 1520 4655 1540
rect 4755 1520 4775 1540
rect 20571 1655 20591 1675
rect 20625 1660 20645 1680
rect 20720 1660 20740 1680
rect 20520 1605 20540 1625
rect 20810 1605 20830 1625
rect 20476 1545 20496 1565
rect 2845 1460 2865 1480
rect 2935 1475 2955 1495
rect 3055 1475 3075 1495
rect 3175 1475 3195 1495
rect 3295 1475 3315 1495
rect 3535 1475 3555 1495
rect 3655 1475 3675 1495
rect 3775 1475 3795 1495
rect 3925 1460 3945 1480
rect 4065 1460 4085 1480
rect 4215 1475 4235 1495
rect 4335 1475 4355 1495
rect 4455 1475 4475 1495
rect 4695 1475 4715 1495
rect 4815 1475 4835 1495
rect 4935 1475 4955 1495
rect 5055 1475 5075 1495
rect 5145 1460 5165 1480
rect 11112 1470 11129 1490
rect 11315 1470 11335 1490
rect 11535 1470 11555 1490
rect 11830 1470 11850 1490
rect 11880 1470 11900 1490
rect 11928 1470 11945 1490
rect 12152 1470 12169 1490
rect 12355 1470 12375 1490
rect 12575 1470 12595 1490
rect 18612 1470 18629 1490
rect 18815 1470 18835 1490
rect 19035 1470 19055 1490
rect 19330 1470 19350 1490
rect 19380 1470 19400 1490
rect 19428 1470 19445 1490
rect 19652 1470 19669 1490
rect 19855 1470 19875 1490
rect 20075 1470 20095 1490
rect 20570 1545 20590 1565
rect 20854 1545 20874 1565
rect 11155 1410 11175 1430
rect 11260 1410 11280 1430
rect 11370 1410 11390 1430
rect 11480 1410 11500 1430
rect 11590 1410 11610 1430
rect 12195 1410 12215 1430
rect 12300 1410 12320 1430
rect 12410 1410 12430 1430
rect 12520 1410 12540 1430
rect 12630 1410 12650 1430
rect 13025 1400 13050 1425
rect 14035 1400 14060 1425
rect 18655 1410 18675 1430
rect 18760 1410 18780 1430
rect 18870 1410 18890 1430
rect 18980 1410 19000 1430
rect 19090 1410 19110 1430
rect 19695 1410 19715 1430
rect 19800 1410 19820 1430
rect 19910 1410 19930 1430
rect 20020 1410 20040 1430
rect 20130 1410 20150 1430
rect 13035 1295 13055 1315
rect 13136 1295 13154 1315
rect 13235 1295 13255 1315
rect 13435 1295 13455 1315
rect 13635 1295 13655 1315
rect 13835 1295 13855 1315
rect 14035 1295 14055 1315
rect 20533 1325 20553 1345
rect 20797 1325 20817 1345
rect 11325 1200 11345 1220
rect 11435 1200 11455 1220
rect 11545 1200 11565 1220
rect 11655 1200 11675 1220
rect 11765 1200 11785 1220
rect 11820 1200 11840 1220
rect 11875 1200 11895 1220
rect 11985 1200 12005 1220
rect 12095 1200 12115 1220
rect 12205 1200 12225 1220
rect 12315 1200 12335 1220
rect 12425 1200 12445 1220
rect 12535 1200 12555 1220
rect 12605 1215 12625 1235
rect 3385 1160 3405 1180
rect 4605 1160 4625 1180
rect 2955 1100 2975 1120
rect 3035 1100 3055 1120
rect 3115 1100 3135 1120
rect 3195 1100 3215 1120
rect 3275 1100 3295 1120
rect 3355 1100 3375 1120
rect 3435 1100 3455 1120
rect 3515 1100 3535 1120
rect 3595 1100 3615 1120
rect 3675 1100 3695 1120
rect 3755 1100 3775 1120
rect 3835 1100 3855 1120
rect 3915 1100 3935 1120
rect 3995 1100 4015 1120
rect 4075 1100 4095 1120
rect 4155 1100 4175 1120
rect 4235 1100 4255 1120
rect 4315 1100 4335 1120
rect 4395 1100 4415 1120
rect 4475 1100 4495 1120
rect 4555 1100 4575 1120
rect 4635 1100 4655 1120
rect 4715 1100 4735 1120
rect 4795 1100 4815 1120
rect 4875 1100 4895 1120
rect 4955 1100 4975 1120
rect 2915 1015 2935 1035
rect 5120 1015 5140 1035
rect 3005 905 3025 925
rect 3185 905 3205 925
rect 3365 905 3385 925
rect 3545 905 3565 925
rect 3725 905 3745 925
rect 3905 905 3925 925
rect 4085 905 4105 925
rect 4265 905 4285 925
rect 4445 905 4465 925
rect 4625 905 4645 925
rect 4805 905 4825 925
rect 18825 1250 18845 1270
rect 18935 1250 18955 1270
rect 19045 1250 19065 1270
rect 19155 1250 19175 1270
rect 19265 1250 19285 1270
rect 19320 1250 19340 1270
rect 19375 1250 19395 1270
rect 19485 1250 19505 1270
rect 19595 1250 19615 1270
rect 19705 1250 19725 1270
rect 19815 1250 19835 1270
rect 19925 1250 19945 1270
rect 20035 1250 20055 1270
rect 20105 1265 20125 1285
rect 20455 1265 20475 1285
rect 20570 1265 20590 1285
rect 20760 1265 20780 1285
rect 20875 1265 20895 1285
rect 20610 1205 20630 1225
rect 20665 1205 20685 1225
rect 20720 1205 20740 1225
rect 13135 945 13155 965
rect 13335 945 13355 965
rect 13535 945 13555 965
rect 13735 945 13755 965
rect 13935 945 13955 965
rect 18675 930 18695 950
rect 4985 905 5005 925
rect 18770 930 18790 950
rect 18880 930 18900 950
rect 18990 930 19010 950
rect 19100 930 19120 950
rect 19210 930 19230 950
rect 19320 930 19340 950
rect 19430 930 19450 950
rect 19540 930 19560 950
rect 19650 930 19670 950
rect 19760 930 19780 950
rect 19870 930 19890 950
rect 19980 930 20000 950
rect 20130 930 20150 950
rect 11175 880 11195 900
rect 11270 880 11290 900
rect 11380 880 11400 900
rect 11490 880 11510 900
rect 11600 880 11620 900
rect 11710 880 11730 900
rect 11820 880 11840 900
rect 11930 880 11950 900
rect 12040 880 12060 900
rect 12150 880 12170 900
rect 12260 880 12280 900
rect 12370 880 12390 900
rect 12480 880 12500 900
rect 12630 880 12650 900
rect 3140 735 3160 755
rect 3275 735 3295 755
rect 3455 735 3475 755
rect 3635 735 3655 755
rect 3815 735 3835 755
rect 3995 735 4015 755
rect 4175 735 4195 755
rect 4355 735 4375 755
rect 4535 735 4555 755
rect 4715 735 4735 755
rect 4895 735 4915 755
rect 9385 -705 9405 -685
rect 9585 -705 9605 -685
rect 9785 -705 9805 -685
rect 9985 -705 10005 -685
rect 10185 -705 10205 -685
rect 10385 -705 10405 -685
rect 9485 -1055 9505 -1035
rect 9685 -1055 9705 -1035
rect 9885 -1055 9905 -1035
rect 10085 -1055 10105 -1035
rect 10285 -1055 10305 -1035
<< metal1 >>
rect 11340 3625 11380 3630
rect 11340 3595 11345 3625
rect 11375 3595 11380 3625
rect 11340 3590 11380 3595
rect 11460 3625 11500 3630
rect 11460 3595 11465 3625
rect 11495 3595 11500 3625
rect 11460 3590 11500 3595
rect 11580 3625 11620 3630
rect 11580 3595 11585 3625
rect 11615 3595 11620 3625
rect 11580 3590 11620 3595
rect 11700 3625 11740 3630
rect 11700 3595 11705 3625
rect 11735 3595 11740 3625
rect 11700 3590 11740 3595
rect 11820 3625 11860 3630
rect 11820 3595 11825 3625
rect 11855 3595 11860 3625
rect 11820 3590 11860 3595
rect 11940 3625 11980 3630
rect 11940 3595 11945 3625
rect 11975 3595 11980 3625
rect 11940 3590 11980 3595
rect 12060 3625 12100 3630
rect 12060 3595 12065 3625
rect 12095 3595 12100 3625
rect 12060 3590 12100 3595
rect 12180 3625 12220 3630
rect 12180 3595 12185 3625
rect 12215 3595 12220 3625
rect 12180 3590 12220 3595
rect 12300 3625 12340 3630
rect 12300 3595 12305 3625
rect 12335 3595 12340 3625
rect 12300 3590 12340 3595
rect 12420 3625 12460 3630
rect 12420 3595 12425 3625
rect 12455 3595 12460 3625
rect 12420 3590 12460 3595
rect 18840 3625 18880 3630
rect 18840 3595 18845 3625
rect 18875 3595 18880 3625
rect 18840 3590 18880 3595
rect 18960 3625 19000 3630
rect 18960 3595 18965 3625
rect 18995 3595 19000 3625
rect 18960 3590 19000 3595
rect 19080 3625 19120 3630
rect 19080 3595 19085 3625
rect 19115 3595 19120 3625
rect 19080 3590 19120 3595
rect 19200 3625 19240 3630
rect 19200 3595 19205 3625
rect 19235 3595 19240 3625
rect 19200 3590 19240 3595
rect 19320 3625 19360 3630
rect 19320 3595 19325 3625
rect 19355 3595 19360 3625
rect 19320 3590 19360 3595
rect 19440 3625 19480 3630
rect 19440 3595 19445 3625
rect 19475 3595 19480 3625
rect 19440 3590 19480 3595
rect 19560 3625 19600 3630
rect 19560 3595 19565 3625
rect 19595 3595 19600 3625
rect 19560 3590 19600 3595
rect 19680 3625 19720 3630
rect 19680 3595 19685 3625
rect 19715 3595 19720 3625
rect 19680 3590 19720 3595
rect 19800 3625 19840 3630
rect 19800 3595 19805 3625
rect 19835 3595 19840 3625
rect 19800 3590 19840 3595
rect 19920 3625 19960 3630
rect 19920 3595 19925 3625
rect 19955 3595 19960 3625
rect 19920 3590 19960 3595
rect 1261 3525 1301 3530
rect 1261 3495 1266 3525
rect 1296 3495 1301 3525
rect 1261 3490 1301 3495
rect 4440 3495 4480 3500
rect -15 3445 25 3450
rect -15 3415 -10 3445
rect 20 3415 25 3445
rect -15 3410 25 3415
rect 940 3445 980 3450
rect 940 3415 945 3445
rect 975 3415 980 3445
rect 940 3410 980 3415
rect -60 3390 -20 3395
rect -60 3360 -55 3390
rect -25 3360 -20 3390
rect -60 3355 -20 3360
rect -50 2860 -30 3355
rect -60 2855 -20 2860
rect -60 2825 -55 2855
rect -25 2825 -20 2855
rect -60 2820 -20 2825
rect -5 2800 15 3410
rect 1205 3340 1245 3345
rect 1205 3310 1210 3340
rect 1240 3310 1245 3340
rect 1205 3305 1245 3310
rect 1160 3285 1200 3290
rect 1160 3255 1165 3285
rect 1195 3255 1200 3285
rect 1160 3250 1200 3255
rect 46 3170 51 3205
rect 86 3170 91 3205
rect 46 3110 51 3145
rect 86 3110 91 3145
rect 1170 3105 1190 3250
rect 1160 3100 1200 3105
rect 1160 3070 1165 3100
rect 1195 3070 1200 3100
rect 1160 3065 1200 3070
rect 46 3030 51 3065
rect 86 3030 91 3065
rect 46 2970 51 3005
rect 86 2970 91 3005
rect 905 2910 1125 2920
rect 905 2880 920 2910
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1125 2910
rect 905 2870 1125 2880
rect 1215 2855 1235 3305
rect 1271 3200 1291 3490
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect 1635 3445 1685 3455
rect 1635 3415 1645 3445
rect 1675 3415 1685 3445
rect 2470 3450 2510 3455
rect 2470 3420 2475 3450
rect 2505 3420 2510 3450
rect 2470 3415 2510 3420
rect 1635 3405 1685 3415
rect 1261 3165 1266 3200
rect 1301 3165 1306 3200
rect 1271 3140 1291 3165
rect 1261 3105 1266 3140
rect 1301 3105 1306 3140
rect 2330 2925 2335 2960
rect 2370 2925 2375 2960
rect 2425 2955 2465 2960
rect 2425 2925 2430 2955
rect 2460 2925 2465 2955
rect 2425 2920 2465 2925
rect 2330 2900 2375 2905
rect 2330 2865 2335 2900
rect 2370 2865 2375 2900
rect 2330 2860 2375 2865
rect 51 2820 56 2855
rect 91 2820 96 2855
rect 724 2820 729 2855
rect 764 2820 769 2855
rect 1205 2850 1245 2855
rect 1205 2820 1210 2850
rect 1240 2820 1245 2850
rect 2340 2840 2360 2860
rect 1205 2815 1245 2820
rect 1261 2805 1266 2840
rect 1301 2805 1306 2840
rect 1960 2805 1965 2840
rect 2000 2805 2005 2840
rect 2330 2835 2370 2840
rect 2330 2805 2335 2835
rect 2365 2805 2370 2835
rect -15 2795 25 2800
rect -15 2765 -10 2795
rect 20 2765 25 2795
rect -15 2760 25 2765
rect 51 2760 56 2795
rect 91 2760 96 2795
rect 724 2760 729 2795
rect 764 2760 769 2795
rect 1271 2750 1291 2805
rect 2330 2800 2370 2805
rect 1261 2745 1301 2750
rect 1261 2715 1266 2745
rect 1296 2715 1301 2745
rect 1261 2710 1301 2715
rect 2150 2745 2190 2750
rect 2150 2715 2155 2745
rect 2185 2715 2190 2745
rect 2150 2710 2190 2715
rect 275 2200 1985 2550
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1715 -70 1720
rect -45 1720 -5 1725
rect -45 1715 -40 1720
rect -75 1695 -40 1715
rect -75 1690 -70 1695
rect -110 1685 -70 1690
rect -45 1690 -40 1695
rect -10 1690 -5 1720
rect -45 1685 -5 1690
rect 275 1190 625 2200
rect 952 1710 1302 1870
rect 952 1680 1270 1710
rect 1297 1680 1302 1710
rect 952 1520 1302 1680
rect 1330 1190 1455 1345
rect 1635 1190 1985 2200
rect 2160 1190 2180 2710
rect 2340 2205 2360 2800
rect 2435 2250 2455 2920
rect 2425 2245 2465 2250
rect 2425 2215 2430 2245
rect 2460 2215 2465 2245
rect 2425 2210 2465 2215
rect 2330 2200 2370 2205
rect 2330 2170 2335 2200
rect 2365 2170 2370 2200
rect 2330 2165 2370 2170
rect 2340 1600 2360 2165
rect 2380 2150 2420 2155
rect 2380 2120 2385 2150
rect 2415 2120 2420 2150
rect 2380 2115 2420 2120
rect 2390 1670 2410 2115
rect 2435 1765 2455 2210
rect 2480 1825 2500 3415
rect 2690 3390 2730 3395
rect 2690 3360 2695 3390
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 3135 3340 3175 3345
rect 3135 3310 3140 3340
rect 3170 3310 3175 3340
rect 3135 3305 3175 3310
rect 3385 3335 3435 3345
rect 3385 3305 3395 3335
rect 3425 3305 3435 3335
rect 2735 3240 2775 3245
rect 2735 3210 2740 3240
rect 2770 3210 2775 3240
rect 2735 3205 2775 3210
rect 2620 3185 2660 3190
rect 2620 3155 2625 3185
rect 2655 3155 2660 3185
rect 2620 3150 2660 3155
rect 2520 2980 2560 2985
rect 2520 2950 2525 2980
rect 2555 2950 2560 2980
rect 2520 2945 2560 2950
rect 2470 1820 2510 1825
rect 2470 1790 2475 1820
rect 2505 1790 2510 1820
rect 2470 1785 2510 1790
rect 2425 1760 2465 1765
rect 2425 1730 2430 1760
rect 2460 1730 2465 1760
rect 2425 1725 2465 1730
rect 2380 1665 2420 1670
rect 2380 1635 2385 1665
rect 2415 1635 2420 1665
rect 2380 1630 2420 1635
rect 2330 1595 2370 1600
rect 2330 1565 2335 1595
rect 2365 1565 2370 1595
rect 2330 1560 2370 1565
rect 275 840 2180 1190
rect 2530 765 2550 2945
rect 2630 2795 2650 3150
rect 2620 2790 2660 2795
rect 2620 2760 2625 2790
rect 2655 2760 2660 2790
rect 2620 2755 2660 2760
rect 2630 2350 2650 2755
rect 2620 2345 2660 2350
rect 2620 2315 2625 2345
rect 2655 2315 2660 2345
rect 2620 2310 2660 2315
rect 2630 2055 2650 2310
rect 2745 2295 2765 3205
rect 3145 3145 3165 3305
rect 3385 3295 3435 3305
rect 4450 3190 4470 3460
rect 5135 3445 5185 3455
rect 5135 3415 5145 3445
rect 5175 3415 5185 3445
rect 5135 3405 5185 3415
rect 5360 3335 5400 3340
rect 5360 3305 5365 3335
rect 5395 3305 5400 3335
rect 5360 3300 5400 3305
rect 4885 3285 4925 3290
rect 4885 3255 4890 3285
rect 4920 3255 4925 3285
rect 4885 3250 4925 3255
rect 4440 3185 4480 3190
rect 4440 3155 4445 3185
rect 4475 3155 4480 3185
rect 4440 3150 4480 3155
rect 3135 3140 3175 3145
rect 3135 3110 3140 3140
rect 3170 3110 3175 3140
rect 3135 3105 3175 3110
rect 4835 3140 4875 3145
rect 4835 3110 4840 3140
rect 4870 3110 4875 3140
rect 4835 3105 4875 3110
rect 3145 2985 3165 3105
rect 3985 3080 4025 3085
rect 3985 3050 3990 3080
rect 4020 3050 4025 3080
rect 3985 3045 4025 3050
rect 3445 3035 3485 3040
rect 3445 3005 3450 3035
rect 3480 3005 3485 3035
rect 3445 3000 3485 3005
rect 3805 3035 3845 3040
rect 3805 3005 3810 3035
rect 3840 3005 3845 3035
rect 3805 3000 3845 3005
rect 3455 2985 3475 3000
rect 3815 2985 3835 3000
rect 3995 2985 4015 3045
rect 4345 3035 4385 3040
rect 4345 3005 4350 3035
rect 4380 3005 4385 3035
rect 4345 3000 4385 3005
rect 4705 3035 4745 3040
rect 4705 3005 4710 3035
rect 4740 3005 4745 3035
rect 4705 3000 4745 3005
rect 4355 2985 4375 3000
rect 4715 2985 4735 3000
rect 4845 2985 4865 3105
rect 4895 2985 4915 3250
rect 5315 3140 5355 3145
rect 5315 3110 5320 3140
rect 5350 3110 5355 3140
rect 5315 3105 5355 3110
rect 3080 2980 3120 2985
rect 3080 2950 3085 2980
rect 3115 2950 3120 2980
rect 3080 2945 3120 2950
rect 3140 2975 3175 2985
rect 3140 2955 3145 2975
rect 3165 2955 3175 2975
rect 3140 2945 3175 2955
rect 3265 2980 3305 2985
rect 3265 2950 3270 2980
rect 3300 2950 3305 2980
rect 3265 2945 3305 2950
rect 3445 2975 3485 2985
rect 3445 2955 3455 2975
rect 3475 2955 3485 2975
rect 3445 2945 3485 2955
rect 3625 2980 3665 2985
rect 3625 2950 3630 2980
rect 3660 2950 3665 2980
rect 3625 2945 3665 2950
rect 3805 2975 3845 2985
rect 3805 2955 3815 2975
rect 3835 2955 3845 2975
rect 3805 2945 3845 2955
rect 3985 2975 4025 2985
rect 3985 2955 3995 2975
rect 4015 2955 4025 2975
rect 3985 2945 4025 2955
rect 4165 2980 4205 2985
rect 4165 2950 4170 2980
rect 4200 2950 4205 2980
rect 4165 2945 4205 2950
rect 4345 2975 4385 2985
rect 4345 2955 4355 2975
rect 4375 2955 4385 2975
rect 4345 2945 4385 2955
rect 4525 2980 4565 2985
rect 4525 2950 4530 2980
rect 4560 2950 4565 2980
rect 4525 2945 4565 2950
rect 4705 2975 4745 2985
rect 4705 2955 4715 2975
rect 4735 2955 4745 2975
rect 4705 2945 4745 2955
rect 4835 2975 4870 2985
rect 4835 2955 4845 2975
rect 4865 2955 4870 2975
rect 4835 2945 4870 2955
rect 4890 2975 4925 2985
rect 4890 2955 4895 2975
rect 4915 2955 4925 2975
rect 4890 2945 4925 2955
rect 2995 2810 3035 2815
rect 2995 2780 3000 2810
rect 3030 2780 3035 2810
rect 2995 2775 3035 2780
rect 3175 2810 3215 2815
rect 3175 2780 3180 2810
rect 3210 2780 3215 2810
rect 3175 2775 3215 2780
rect 3355 2810 3395 2815
rect 3355 2780 3360 2810
rect 3390 2780 3395 2810
rect 3355 2775 3395 2780
rect 3535 2810 3575 2815
rect 3535 2780 3540 2810
rect 3570 2780 3575 2810
rect 3535 2775 3575 2780
rect 3715 2810 3755 2815
rect 3715 2780 3720 2810
rect 3750 2780 3755 2810
rect 3715 2775 3755 2780
rect 3895 2810 3935 2815
rect 3895 2780 3900 2810
rect 3930 2780 3935 2810
rect 3895 2775 3935 2780
rect 4075 2810 4115 2815
rect 4075 2780 4080 2810
rect 4110 2780 4115 2810
rect 4075 2775 4115 2780
rect 4255 2810 4295 2815
rect 4255 2780 4260 2810
rect 4290 2780 4295 2810
rect 4255 2775 4295 2780
rect 4435 2810 4475 2815
rect 4435 2780 4440 2810
rect 4470 2780 4475 2810
rect 4435 2775 4475 2780
rect 4615 2810 4655 2815
rect 4615 2780 4620 2810
rect 4650 2780 4655 2810
rect 4615 2775 4655 2780
rect 4795 2810 4835 2815
rect 4795 2780 4800 2810
rect 4830 2780 4835 2810
rect 4795 2775 4835 2780
rect 4975 2810 5015 2815
rect 4975 2780 4980 2810
rect 5010 2780 5015 2810
rect 4975 2775 5015 2780
rect 4805 2755 4825 2775
rect 3175 2750 3215 2755
rect 3175 2720 3180 2750
rect 3210 2720 3215 2750
rect 3175 2715 3215 2720
rect 3355 2750 3395 2755
rect 3355 2720 3360 2750
rect 3390 2720 3395 2750
rect 3355 2715 3395 2720
rect 3535 2750 3575 2755
rect 3535 2720 3540 2750
rect 3570 2720 3575 2750
rect 3535 2715 3575 2720
rect 3715 2750 3755 2755
rect 3715 2720 3720 2750
rect 3750 2720 3755 2750
rect 3715 2715 3755 2720
rect 3895 2750 3935 2755
rect 3895 2720 3900 2750
rect 3930 2720 3935 2750
rect 3895 2715 3935 2720
rect 4075 2750 4115 2755
rect 4075 2720 4080 2750
rect 4110 2720 4115 2750
rect 4075 2715 4115 2720
rect 4255 2750 4295 2755
rect 4255 2720 4260 2750
rect 4290 2720 4295 2750
rect 4255 2715 4295 2720
rect 4435 2750 4475 2755
rect 4435 2720 4440 2750
rect 4470 2720 4475 2750
rect 4435 2715 4475 2720
rect 4615 2750 4655 2755
rect 4615 2720 4620 2750
rect 4650 2720 4655 2750
rect 4615 2715 4655 2720
rect 4795 2750 4835 2755
rect 4795 2720 4800 2750
rect 4830 2720 4835 2750
rect 4795 2715 4835 2720
rect 3265 2375 3305 2385
rect 3265 2355 3275 2375
rect 3295 2355 3305 2375
rect 3265 2345 3305 2355
rect 3355 2375 3395 2380
rect 3355 2345 3360 2375
rect 3390 2345 3395 2375
rect 3445 2375 3485 2385
rect 3445 2355 3455 2375
rect 3475 2355 3485 2375
rect 3445 2345 3485 2355
rect 3805 2380 3845 2385
rect 3805 2350 3810 2380
rect 3840 2350 3845 2380
rect 3805 2345 3845 2350
rect 3885 2375 3925 2385
rect 3885 2355 3895 2375
rect 3915 2355 3925 2375
rect 3885 2345 3925 2355
rect 3985 2375 4025 2385
rect 3985 2355 3995 2375
rect 4015 2355 4025 2375
rect 3985 2345 4025 2355
rect 4165 2380 4205 2385
rect 4165 2350 4170 2380
rect 4200 2350 4205 2380
rect 4165 2345 4205 2350
rect 4525 2375 4565 2385
rect 4525 2355 4535 2375
rect 4555 2355 4565 2375
rect 4525 2345 4565 2355
rect 4705 2375 4745 2385
rect 4705 2355 4715 2375
rect 4735 2355 4745 2375
rect 4705 2345 4745 2355
rect 2735 2290 2775 2295
rect 2735 2260 2740 2290
rect 2770 2260 2775 2290
rect 2735 2255 2775 2260
rect 3275 2205 3295 2345
rect 3355 2340 3395 2345
rect 3455 2295 3475 2345
rect 3625 2335 3665 2340
rect 3625 2305 3630 2335
rect 3660 2305 3665 2335
rect 3625 2300 3665 2305
rect 3445 2290 3485 2295
rect 3445 2260 3450 2290
rect 3480 2260 3485 2290
rect 3445 2255 3485 2260
rect 3265 2200 3305 2205
rect 3265 2170 3270 2200
rect 3300 2170 3305 2200
rect 3265 2165 3305 2170
rect 3635 2155 3655 2300
rect 3815 2250 3835 2345
rect 3805 2245 3845 2250
rect 3805 2215 3810 2245
rect 3840 2215 3845 2245
rect 3805 2210 3845 2215
rect 3625 2150 3665 2155
rect 3625 2120 3630 2150
rect 3660 2120 3665 2150
rect 3625 2115 3665 2120
rect 2745 2095 2785 2100
rect 2745 2065 2750 2095
rect 2780 2065 2785 2095
rect 2745 2060 2785 2065
rect 2865 2095 2905 2100
rect 2865 2065 2870 2095
rect 2900 2065 2905 2095
rect 2865 2060 2905 2065
rect 2985 2095 3025 2100
rect 2985 2065 2990 2095
rect 3020 2065 3025 2095
rect 2985 2060 3025 2065
rect 3105 2095 3145 2100
rect 3105 2065 3110 2095
rect 3140 2065 3145 2095
rect 3105 2060 3145 2065
rect 3225 2095 3265 2100
rect 3225 2065 3230 2095
rect 3260 2065 3265 2095
rect 3225 2060 3265 2065
rect 3345 2095 3385 2100
rect 3345 2065 3350 2095
rect 3380 2065 3385 2095
rect 3345 2060 3385 2065
rect 3465 2095 3505 2100
rect 3465 2065 3470 2095
rect 3500 2065 3505 2095
rect 3465 2060 3505 2065
rect 3585 2095 3625 2100
rect 3585 2065 3590 2095
rect 3620 2065 3625 2095
rect 3585 2060 3625 2065
rect 3705 2095 3745 2100
rect 3705 2065 3710 2095
rect 3740 2065 3745 2095
rect 3705 2060 3745 2065
rect 3825 2095 3865 2100
rect 3825 2065 3830 2095
rect 3860 2065 3865 2095
rect 3825 2060 3865 2065
rect 3895 2055 3915 2345
rect 3995 2205 4015 2345
rect 4345 2335 4385 2340
rect 4345 2305 4350 2335
rect 4380 2305 4385 2335
rect 4345 2300 4385 2305
rect 4535 2295 4555 2345
rect 4525 2290 4565 2295
rect 4525 2260 4530 2290
rect 4560 2260 4565 2290
rect 4525 2255 4565 2260
rect 4715 2205 4735 2345
rect 5270 2290 5310 2295
rect 5270 2260 5275 2290
rect 5305 2260 5310 2290
rect 5270 2255 5310 2260
rect 3985 2200 4025 2205
rect 3985 2170 3990 2200
rect 4020 2170 4025 2200
rect 3985 2165 4025 2170
rect 4705 2200 4745 2205
rect 4705 2170 4710 2200
rect 4740 2170 4745 2200
rect 4705 2165 4745 2170
rect 4085 2145 4125 2150
rect 4085 2115 4090 2145
rect 4120 2115 4125 2145
rect 4085 2110 4125 2115
rect 3985 2095 4025 2100
rect 3985 2065 3990 2095
rect 4020 2065 4025 2095
rect 3985 2060 4025 2065
rect 4095 2055 4115 2110
rect 4145 2095 4185 2100
rect 4145 2065 4150 2095
rect 4180 2065 4185 2095
rect 4145 2060 4185 2065
rect 4265 2095 4305 2100
rect 4265 2065 4270 2095
rect 4300 2065 4305 2095
rect 4265 2060 4305 2065
rect 4385 2095 4425 2100
rect 4385 2065 4390 2095
rect 4420 2065 4425 2095
rect 4385 2060 4425 2065
rect 4505 2095 4545 2100
rect 4505 2065 4510 2095
rect 4540 2065 4545 2095
rect 4505 2060 4545 2065
rect 4625 2095 4665 2100
rect 4625 2065 4630 2095
rect 4660 2065 4665 2095
rect 4625 2060 4665 2065
rect 4745 2095 4785 2100
rect 4745 2065 4750 2095
rect 4780 2065 4785 2095
rect 4745 2060 4785 2065
rect 4865 2095 4905 2100
rect 4865 2065 4870 2095
rect 4900 2065 4905 2095
rect 4865 2060 4905 2065
rect 4985 2095 5025 2100
rect 4985 2065 4990 2095
rect 5020 2065 5025 2095
rect 4985 2060 5025 2065
rect 5105 2095 5145 2100
rect 5105 2065 5110 2095
rect 5140 2065 5145 2095
rect 5105 2060 5145 2065
rect 5225 2095 5265 2100
rect 5225 2065 5230 2095
rect 5260 2065 5265 2095
rect 5225 2060 5265 2065
rect 2620 2050 2660 2055
rect 2620 2020 2625 2050
rect 2655 2020 2660 2050
rect 2620 2015 2660 2020
rect 2805 2050 2845 2055
rect 2805 2020 2810 2050
rect 2840 2020 2845 2050
rect 2805 2015 2845 2020
rect 3165 2050 3205 2055
rect 3165 2020 3170 2050
rect 3200 2020 3205 2050
rect 3165 2015 3205 2020
rect 3525 2050 3565 2055
rect 3525 2020 3530 2050
rect 3560 2020 3565 2050
rect 3525 2015 3565 2020
rect 3885 2050 3925 2055
rect 3885 2020 3890 2050
rect 3920 2045 3925 2050
rect 4085 2050 4125 2055
rect 4085 2045 4090 2050
rect 3920 2020 3945 2045
rect 3885 2015 3945 2020
rect 2565 1875 2600 1885
rect 2565 1855 2575 1875
rect 2595 1855 2600 1875
rect 2565 1845 2600 1855
rect 2620 1875 2660 1885
rect 2620 1855 2630 1875
rect 2650 1855 2660 1875
rect 2620 1845 2660 1855
rect 2680 1875 2715 1885
rect 2680 1855 2685 1875
rect 2705 1855 2715 1875
rect 2680 1845 2715 1855
rect 2835 1875 2875 1885
rect 2835 1855 2845 1875
rect 2865 1855 2875 1875
rect 2835 1845 2875 1855
rect 2925 1880 2965 1885
rect 2925 1850 2930 1880
rect 2960 1850 2965 1880
rect 2925 1845 2965 1850
rect 3045 1875 3085 1885
rect 3045 1855 3055 1875
rect 3075 1855 3085 1875
rect 3045 1845 3085 1855
rect 3165 1875 3205 1885
rect 3165 1855 3175 1875
rect 3195 1855 3205 1875
rect 3165 1845 3205 1855
rect 3285 1880 3325 1885
rect 3285 1850 3290 1880
rect 3320 1850 3325 1880
rect 3285 1845 3325 1850
rect 3405 1875 3445 1885
rect 3405 1855 3415 1875
rect 3435 1855 3445 1875
rect 3405 1845 3445 1855
rect 3525 1875 3565 1885
rect 3525 1855 3535 1875
rect 3555 1855 3565 1875
rect 3525 1845 3565 1855
rect 3645 1880 3685 1885
rect 3645 1850 3650 1880
rect 3680 1850 3685 1880
rect 3645 1845 3685 1850
rect 3765 1875 3805 1885
rect 3765 1855 3775 1875
rect 3795 1855 3805 1875
rect 3765 1845 3805 1855
rect 3855 1875 3895 1885
rect 3855 1855 3865 1875
rect 3885 1855 3895 1875
rect 3855 1845 3895 1855
rect 2575 1765 2595 1845
rect 2565 1760 2605 1765
rect 2565 1730 2570 1760
rect 2600 1730 2605 1760
rect 2565 1725 2605 1730
rect 2630 1670 2650 1845
rect 2685 1765 2705 1845
rect 2845 1825 2865 1845
rect 3055 1825 3075 1845
rect 3175 1825 3195 1845
rect 2835 1820 2875 1825
rect 2835 1790 2840 1820
rect 2870 1790 2875 1820
rect 2835 1785 2875 1790
rect 3045 1820 3085 1825
rect 3045 1790 3050 1820
rect 3080 1790 3085 1820
rect 3045 1785 3085 1790
rect 3165 1820 3205 1825
rect 3165 1790 3170 1820
rect 3200 1790 3205 1820
rect 3165 1785 3205 1790
rect 2800 1765 2840 1770
rect 3295 1765 3315 1845
rect 3415 1825 3435 1845
rect 3535 1825 3555 1845
rect 3775 1825 3795 1845
rect 3865 1825 3885 1845
rect 3405 1820 3445 1825
rect 3405 1790 3410 1820
rect 3440 1790 3445 1820
rect 3405 1785 3445 1790
rect 3525 1820 3565 1825
rect 3525 1790 3530 1820
rect 3560 1790 3565 1820
rect 3525 1785 3565 1790
rect 3765 1820 3805 1825
rect 3765 1790 3770 1820
rect 3800 1790 3805 1820
rect 3765 1785 3805 1790
rect 3855 1820 3895 1825
rect 3855 1790 3860 1820
rect 3890 1790 3895 1820
rect 3855 1785 3895 1790
rect 2675 1760 2715 1765
rect 2675 1730 2680 1760
rect 2710 1730 2715 1760
rect 2800 1735 2805 1765
rect 2835 1735 2840 1765
rect 2800 1730 2840 1735
rect 3225 1760 3265 1765
rect 3225 1730 3230 1760
rect 3260 1730 3265 1760
rect 2675 1725 2715 1730
rect 2810 1715 2830 1730
rect 3225 1725 3265 1730
rect 3285 1760 3325 1765
rect 3285 1730 3290 1760
rect 3320 1730 3325 1760
rect 3285 1725 3325 1730
rect 3415 1720 3435 1785
rect 3525 1760 3565 1765
rect 3525 1730 3530 1760
rect 3560 1730 3565 1760
rect 3525 1725 3565 1730
rect 3765 1760 3805 1765
rect 3765 1730 3770 1760
rect 3800 1730 3805 1760
rect 3765 1725 3805 1730
rect 3165 1715 3205 1720
rect 2800 1710 2840 1715
rect 2800 1680 2805 1710
rect 2835 1680 2840 1710
rect 3165 1685 3170 1715
rect 3200 1685 3205 1715
rect 3165 1680 3205 1685
rect 3405 1715 3445 1720
rect 3405 1685 3410 1715
rect 3440 1685 3445 1715
rect 3405 1680 3445 1685
rect 3645 1715 3685 1720
rect 3645 1685 3650 1715
rect 3680 1685 3685 1715
rect 3645 1680 3685 1685
rect 2800 1675 2840 1680
rect 2620 1665 2660 1670
rect 2620 1635 2625 1665
rect 2655 1635 2660 1665
rect 2620 1630 2660 1635
rect 2630 1045 2650 1630
rect 3165 1595 3205 1600
rect 3165 1565 3170 1595
rect 3200 1565 3205 1595
rect 3165 1560 3205 1565
rect 2835 1545 2875 1550
rect 2835 1515 2840 1545
rect 2870 1515 2875 1545
rect 2835 1510 2875 1515
rect 3225 1545 3265 1550
rect 3225 1515 3230 1545
rect 3260 1515 3265 1545
rect 3225 1510 3265 1515
rect 3345 1545 3385 1550
rect 3345 1515 3350 1545
rect 3380 1515 3385 1545
rect 3345 1510 3385 1515
rect 3465 1545 3505 1550
rect 3465 1515 3470 1545
rect 3500 1515 3505 1545
rect 3465 1510 3505 1515
rect 3585 1545 3625 1550
rect 3585 1515 3590 1545
rect 3620 1515 3625 1545
rect 3585 1510 3625 1515
rect 3705 1545 3745 1550
rect 3705 1515 3710 1545
rect 3740 1515 3745 1545
rect 3705 1510 3745 1515
rect 2845 1490 2865 1510
rect 2925 1500 2965 1505
rect 2835 1480 2875 1490
rect 2835 1460 2845 1480
rect 2865 1460 2875 1480
rect 2925 1470 2930 1500
rect 2960 1470 2965 1500
rect 2925 1465 2965 1470
rect 3045 1500 3085 1505
rect 3045 1470 3050 1500
rect 3080 1470 3085 1500
rect 3045 1465 3085 1470
rect 3165 1500 3205 1505
rect 3165 1470 3170 1500
rect 3200 1470 3205 1500
rect 3165 1465 3205 1470
rect 3285 1500 3325 1505
rect 3285 1470 3290 1500
rect 3320 1470 3325 1500
rect 3285 1465 3325 1470
rect 3525 1500 3565 1505
rect 3525 1470 3530 1500
rect 3560 1470 3565 1500
rect 3525 1465 3565 1470
rect 3645 1500 3685 1505
rect 3645 1470 3650 1500
rect 3680 1470 3685 1500
rect 3645 1465 3685 1470
rect 3765 1500 3805 1505
rect 3765 1470 3770 1500
rect 3800 1470 3805 1500
rect 3925 1490 3945 2015
rect 4065 2020 4090 2045
rect 4120 2020 4125 2050
rect 4065 2015 4125 2020
rect 4445 2050 4485 2055
rect 4445 2020 4450 2050
rect 4480 2020 4485 2050
rect 4445 2015 4485 2020
rect 4805 2050 4845 2055
rect 4805 2020 4810 2050
rect 4840 2020 4845 2050
rect 4805 2015 4845 2020
rect 5165 2050 5205 2055
rect 5165 2020 5170 2050
rect 5200 2020 5205 2050
rect 5165 2015 5205 2020
rect 3985 1650 4025 1660
rect 3985 1630 3995 1650
rect 4015 1630 4025 1650
rect 3985 1620 4025 1630
rect 3765 1465 3805 1470
rect 3915 1480 3955 1490
rect 2835 1450 2875 1460
rect 3915 1460 3925 1480
rect 3945 1460 3955 1480
rect 3915 1450 3955 1460
rect 3995 1190 4015 1620
rect 4065 1490 4085 2015
rect 4115 1875 4155 1885
rect 4115 1855 4125 1875
rect 4145 1855 4155 1875
rect 4115 1845 4155 1855
rect 4205 1875 4245 1885
rect 4205 1855 4215 1875
rect 4235 1855 4245 1875
rect 4205 1845 4245 1855
rect 4325 1880 4365 1885
rect 4325 1850 4330 1880
rect 4360 1850 4365 1880
rect 4325 1845 4365 1850
rect 4445 1875 4485 1885
rect 4445 1855 4455 1875
rect 4475 1855 4485 1875
rect 4445 1845 4485 1855
rect 4565 1875 4605 1885
rect 4565 1855 4575 1875
rect 4595 1855 4605 1875
rect 4565 1845 4605 1855
rect 4685 1880 4725 1885
rect 4685 1850 4690 1880
rect 4720 1850 4725 1880
rect 4685 1845 4725 1850
rect 4805 1875 4845 1885
rect 4805 1855 4815 1875
rect 4835 1855 4845 1875
rect 4805 1845 4845 1855
rect 4925 1875 4965 1885
rect 4925 1855 4935 1875
rect 4955 1855 4965 1875
rect 4925 1845 4965 1855
rect 5045 1880 5085 1885
rect 5045 1850 5050 1880
rect 5080 1850 5085 1880
rect 5045 1845 5085 1850
rect 5135 1875 5175 1885
rect 5135 1855 5145 1875
rect 5165 1855 5175 1875
rect 5135 1845 5175 1855
rect 4125 1825 4145 1845
rect 4215 1825 4235 1845
rect 4455 1825 4475 1845
rect 4575 1825 4595 1845
rect 4115 1820 4155 1825
rect 4115 1790 4120 1820
rect 4150 1790 4155 1820
rect 4115 1785 4155 1790
rect 4205 1820 4245 1825
rect 4205 1790 4210 1820
rect 4240 1790 4245 1820
rect 4205 1785 4245 1790
rect 4445 1820 4485 1825
rect 4445 1790 4450 1820
rect 4480 1790 4485 1820
rect 4445 1785 4485 1790
rect 4565 1820 4605 1825
rect 4565 1790 4570 1820
rect 4600 1790 4605 1820
rect 4565 1785 4605 1790
rect 4205 1760 4245 1765
rect 4205 1730 4210 1760
rect 4240 1730 4245 1760
rect 4205 1725 4245 1730
rect 4445 1760 4485 1765
rect 4445 1730 4450 1760
rect 4480 1730 4485 1760
rect 4445 1725 4485 1730
rect 4575 1720 4595 1785
rect 4695 1765 4715 1845
rect 4815 1825 4835 1845
rect 4935 1825 4955 1845
rect 5145 1825 5165 1845
rect 4805 1820 4845 1825
rect 4805 1790 4810 1820
rect 4840 1790 4845 1820
rect 4805 1785 4845 1790
rect 4925 1820 4965 1825
rect 4925 1790 4930 1820
rect 4960 1790 4965 1820
rect 4925 1785 4965 1790
rect 5135 1820 5175 1825
rect 5135 1790 5140 1820
rect 5170 1790 5175 1820
rect 5135 1785 5175 1790
rect 5280 1765 5300 2255
rect 5325 2150 5345 3105
rect 5315 2145 5355 2150
rect 5315 2115 5320 2145
rect 5350 2115 5355 2145
rect 5315 2110 5355 2115
rect 5370 1825 5390 3300
rect 12945 3290 12985 3295
rect 5410 3285 5450 3290
rect 5410 3255 5415 3285
rect 5445 3255 5450 3285
rect 12945 3260 12950 3290
rect 12980 3260 12985 3290
rect 12945 3255 12985 3260
rect 13055 3290 13095 3295
rect 13055 3260 13060 3290
rect 13090 3260 13095 3290
rect 13055 3255 13095 3260
rect 13165 3290 13205 3295
rect 13165 3260 13170 3290
rect 13200 3260 13205 3290
rect 13165 3255 13205 3260
rect 13275 3290 13315 3295
rect 13275 3260 13280 3290
rect 13310 3260 13315 3290
rect 13275 3255 13315 3260
rect 13385 3290 13425 3295
rect 13385 3260 13390 3290
rect 13420 3260 13425 3290
rect 13385 3255 13425 3260
rect 13495 3290 13535 3295
rect 13495 3260 13500 3290
rect 13530 3260 13535 3290
rect 13495 3255 13535 3260
rect 13605 3290 13645 3295
rect 13605 3260 13610 3290
rect 13640 3260 13645 3290
rect 13605 3255 13645 3260
rect 13715 3290 13755 3295
rect 13715 3260 13720 3290
rect 13750 3260 13755 3290
rect 13715 3255 13755 3260
rect 13825 3290 13865 3295
rect 13825 3260 13830 3290
rect 13860 3260 13865 3290
rect 13825 3255 13865 3260
rect 13935 3290 13975 3295
rect 13935 3260 13940 3290
rect 13970 3260 13975 3290
rect 13935 3255 13975 3260
rect 14045 3290 14085 3295
rect 14045 3260 14050 3290
rect 14080 3260 14085 3290
rect 14045 3255 14085 3260
rect 20445 3290 20485 3295
rect 20445 3260 20450 3290
rect 20480 3260 20485 3290
rect 20445 3255 20485 3260
rect 20555 3290 20595 3295
rect 20555 3260 20560 3290
rect 20590 3260 20595 3290
rect 20555 3255 20595 3260
rect 20665 3290 20705 3295
rect 20665 3260 20670 3290
rect 20700 3260 20705 3290
rect 20665 3255 20705 3260
rect 20775 3290 20815 3295
rect 20775 3260 20780 3290
rect 20810 3260 20815 3290
rect 20775 3255 20815 3260
rect 20885 3290 20925 3295
rect 20885 3260 20890 3290
rect 20920 3260 20925 3290
rect 20885 3255 20925 3260
rect 20995 3290 21035 3295
rect 20995 3260 21000 3290
rect 21030 3260 21035 3290
rect 20995 3255 21035 3260
rect 21105 3290 21145 3295
rect 21105 3260 21110 3290
rect 21140 3260 21145 3290
rect 21105 3255 21145 3260
rect 21215 3290 21255 3295
rect 21215 3260 21220 3290
rect 21250 3260 21255 3290
rect 21215 3255 21255 3260
rect 21325 3290 21365 3295
rect 21325 3260 21330 3290
rect 21360 3260 21365 3290
rect 21325 3255 21365 3260
rect 21435 3290 21475 3295
rect 21435 3260 21440 3290
rect 21470 3260 21475 3290
rect 21435 3255 21475 3260
rect 21545 3290 21585 3295
rect 21545 3260 21550 3290
rect 21580 3260 21585 3290
rect 21545 3255 21585 3260
rect 5410 3250 5450 3255
rect 5360 1820 5400 1825
rect 5360 1790 5365 1820
rect 5395 1790 5400 1820
rect 5360 1785 5400 1790
rect 4685 1760 4725 1765
rect 4685 1730 4690 1760
rect 4720 1730 4725 1760
rect 4685 1725 4725 1730
rect 4745 1760 4785 1765
rect 4745 1730 4750 1760
rect 4780 1730 4785 1760
rect 4745 1725 4785 1730
rect 5270 1760 5310 1765
rect 5270 1730 5275 1760
rect 5305 1730 5310 1760
rect 5270 1725 5310 1730
rect 4325 1715 4365 1720
rect 4325 1685 4330 1715
rect 4360 1685 4365 1715
rect 4325 1680 4365 1685
rect 4565 1715 4605 1720
rect 4565 1685 4570 1715
rect 4600 1685 4605 1715
rect 4565 1680 4605 1685
rect 4805 1715 4845 1720
rect 4805 1685 4810 1715
rect 4840 1685 4845 1715
rect 4805 1680 4845 1685
rect 5420 1600 5440 3250
rect 10580 3210 10620 3215
rect 10580 3180 10585 3210
rect 10615 3180 10620 3210
rect 10580 3175 10620 3180
rect 10905 3205 10940 3215
rect 10905 3185 10910 3205
rect 10930 3185 10940 3205
rect 10905 3175 10940 3185
rect 10980 3210 11015 3215
rect 10980 3180 10985 3210
rect 10980 3175 11015 3180
rect 18080 3210 18120 3215
rect 18080 3180 18085 3210
rect 18115 3180 18120 3210
rect 18080 3175 18120 3180
rect 18405 3205 18440 3215
rect 18405 3185 18410 3205
rect 18430 3185 18440 3205
rect 18405 3175 18440 3185
rect 18480 3210 18515 3215
rect 18480 3180 18485 3210
rect 18480 3175 18515 3180
rect 10910 3160 10930 3175
rect 10900 3155 10940 3160
rect 10900 3125 10905 3155
rect 10935 3125 10940 3155
rect 10900 3120 10940 3125
rect 9735 2670 9775 2675
rect 9735 2640 9740 2670
rect 9770 2640 9775 2670
rect 9735 2635 9775 2640
rect 9845 2670 9885 2675
rect 9845 2640 9850 2670
rect 9880 2640 9885 2670
rect 9845 2635 9885 2640
rect 9955 2670 9995 2675
rect 9955 2640 9960 2670
rect 9990 2640 9995 2670
rect 9955 2635 9995 2640
rect 10065 2670 10105 2675
rect 10065 2640 10070 2670
rect 10100 2640 10105 2670
rect 10065 2635 10105 2640
rect 10175 2670 10215 2675
rect 10175 2640 10180 2670
rect 10210 2640 10215 2670
rect 10175 2635 10215 2640
rect 10285 2670 10325 2675
rect 10285 2640 10290 2670
rect 10320 2640 10325 2670
rect 10285 2635 10325 2640
rect 10395 2670 10435 2675
rect 10395 2640 10400 2670
rect 10430 2640 10435 2670
rect 10395 2635 10435 2640
rect 10505 2670 10545 2675
rect 10505 2640 10510 2670
rect 10540 2640 10545 2670
rect 10505 2635 10545 2640
rect 10615 2670 10655 2675
rect 10615 2640 10620 2670
rect 10650 2640 10655 2670
rect 10615 2635 10655 2640
rect 10725 2670 10765 2675
rect 10725 2640 10730 2670
rect 10760 2640 10765 2670
rect 10725 2635 10765 2640
rect 10835 2670 10875 2675
rect 10835 2640 10840 2670
rect 10870 2640 10875 2670
rect 10835 2635 10875 2640
rect 9790 2500 9830 2505
rect 9790 2470 9795 2500
rect 9825 2470 9830 2500
rect 9790 2465 9830 2470
rect 9900 2500 9940 2505
rect 9900 2470 9905 2500
rect 9935 2470 9940 2500
rect 9900 2465 9940 2470
rect 10010 2500 10050 2505
rect 10010 2470 10015 2500
rect 10045 2470 10050 2500
rect 10010 2465 10050 2470
rect 10120 2500 10160 2505
rect 10120 2470 10125 2500
rect 10155 2470 10160 2500
rect 10120 2465 10160 2470
rect 10230 2500 10270 2505
rect 10230 2470 10235 2500
rect 10265 2470 10270 2500
rect 10230 2465 10270 2470
rect 10340 2500 10380 2505
rect 10340 2470 10345 2500
rect 10375 2470 10380 2500
rect 10340 2465 10380 2470
rect 10450 2500 10490 2505
rect 10450 2470 10455 2500
rect 10485 2470 10490 2500
rect 10450 2465 10490 2470
rect 10560 2500 10600 2505
rect 10560 2470 10565 2500
rect 10595 2470 10600 2500
rect 10560 2465 10600 2470
rect 10670 2500 10710 2505
rect 10670 2470 10675 2500
rect 10705 2470 10710 2500
rect 10670 2465 10710 2470
rect 10780 2500 10820 2505
rect 10780 2470 10785 2500
rect 10815 2470 10820 2500
rect 10990 2480 11010 3175
rect 18410 3160 18430 3175
rect 11280 3150 11320 3160
rect 11280 3130 11290 3150
rect 11310 3130 11320 3150
rect 11280 3120 11320 3130
rect 11400 3150 11440 3160
rect 11400 3130 11410 3150
rect 11430 3130 11440 3150
rect 11400 3120 11440 3130
rect 11520 3150 11560 3160
rect 11520 3130 11530 3150
rect 11550 3130 11560 3150
rect 11520 3120 11560 3130
rect 11640 3150 11680 3160
rect 11640 3130 11650 3150
rect 11670 3130 11680 3150
rect 11640 3120 11680 3130
rect 11760 3150 11800 3160
rect 11760 3130 11770 3150
rect 11790 3130 11800 3150
rect 11760 3120 11800 3130
rect 11823 3155 11857 3160
rect 11823 3125 11826 3155
rect 11854 3125 11857 3155
rect 11823 3120 11857 3125
rect 11880 3150 11920 3160
rect 11880 3130 11890 3150
rect 11910 3130 11920 3150
rect 11880 3120 11920 3130
rect 12000 3150 12040 3160
rect 12000 3130 12010 3150
rect 12030 3130 12040 3150
rect 12000 3120 12040 3130
rect 12120 3150 12160 3160
rect 12120 3130 12130 3150
rect 12150 3130 12160 3150
rect 12120 3120 12160 3130
rect 12240 3150 12280 3160
rect 12240 3130 12250 3150
rect 12270 3130 12280 3150
rect 12240 3120 12280 3130
rect 12360 3150 12400 3160
rect 12360 3130 12370 3150
rect 12390 3130 12400 3150
rect 12360 3120 12400 3130
rect 12480 3150 12520 3160
rect 12480 3130 12490 3150
rect 12510 3130 12520 3150
rect 12480 3120 12520 3130
rect 18400 3155 18440 3160
rect 18400 3125 18405 3155
rect 18435 3125 18440 3155
rect 18400 3120 18440 3125
rect 11290 3105 11310 3120
rect 11280 3100 11320 3105
rect 11280 3070 11285 3100
rect 11315 3070 11320 3100
rect 11280 3065 11320 3070
rect 11410 3060 11430 3120
rect 11530 3105 11550 3120
rect 11520 3100 11560 3105
rect 11520 3070 11525 3100
rect 11555 3070 11560 3100
rect 11520 3065 11560 3070
rect 11650 3060 11670 3120
rect 11770 3105 11790 3120
rect 11760 3100 11800 3105
rect 11760 3070 11765 3100
rect 11795 3070 11800 3100
rect 11760 3065 11800 3070
rect 11890 3060 11910 3120
rect 12010 3105 12030 3120
rect 12000 3100 12040 3105
rect 12000 3070 12005 3100
rect 12035 3070 12040 3100
rect 12000 3065 12040 3070
rect 12130 3060 12150 3120
rect 12250 3105 12270 3120
rect 12240 3100 12280 3105
rect 12240 3070 12245 3100
rect 12275 3070 12280 3100
rect 12240 3065 12280 3070
rect 12370 3060 12390 3120
rect 12490 3105 12510 3120
rect 12480 3100 12520 3105
rect 12480 3070 12485 3100
rect 12515 3070 12520 3100
rect 12480 3065 12520 3070
rect 11400 3055 11440 3060
rect 11400 3025 11405 3055
rect 11435 3025 11440 3055
rect 11400 3020 11440 3025
rect 11640 3055 11680 3060
rect 11640 3025 11645 3055
rect 11675 3025 11680 3055
rect 11640 3020 11680 3025
rect 11880 3055 11920 3060
rect 11880 3025 11885 3055
rect 11915 3025 11920 3055
rect 11880 3020 11920 3025
rect 12120 3055 12160 3060
rect 12120 3025 12125 3055
rect 12155 3025 12160 3055
rect 12120 3020 12160 3025
rect 12360 3055 12400 3060
rect 12360 3025 12365 3055
rect 12395 3025 12400 3055
rect 12360 3020 12400 3025
rect 11410 3005 11430 3020
rect 11340 3000 11380 3005
rect 11340 2970 11345 3000
rect 11375 2970 11380 3000
rect 11340 2965 11380 2970
rect 11400 3000 11440 3005
rect 11400 2970 11405 3000
rect 11435 2970 11440 3000
rect 11400 2965 11440 2970
rect 11580 3000 11620 3005
rect 11580 2970 11585 3000
rect 11615 2970 11620 3000
rect 11580 2965 11620 2970
rect 11820 3000 11860 3005
rect 11820 2970 11825 3000
rect 11855 2970 11860 3000
rect 11820 2965 11860 2970
rect 12060 3000 12100 3005
rect 12060 2970 12065 3000
rect 12095 2970 12100 3000
rect 12060 2965 12100 2970
rect 12300 3000 12340 3005
rect 12300 2970 12305 3000
rect 12335 2970 12340 3000
rect 12300 2965 12340 2970
rect 11350 2950 11370 2965
rect 11590 2950 11610 2965
rect 11830 2950 11850 2965
rect 12070 2950 12090 2965
rect 12310 2950 12330 2965
rect 12490 2950 12510 3065
rect 11340 2940 11380 2950
rect 11340 2920 11350 2940
rect 11370 2920 11380 2940
rect 11340 2910 11380 2920
rect 11460 2945 11500 2950
rect 11460 2915 11465 2945
rect 11495 2915 11500 2945
rect 11460 2910 11500 2915
rect 11580 2940 11620 2950
rect 11580 2920 11590 2940
rect 11610 2920 11620 2940
rect 11580 2910 11620 2920
rect 11700 2945 11740 2950
rect 11700 2915 11705 2945
rect 11735 2915 11740 2945
rect 11700 2910 11740 2915
rect 11820 2940 11860 2950
rect 11820 2920 11830 2940
rect 11850 2920 11860 2940
rect 11820 2910 11860 2920
rect 11940 2945 11980 2950
rect 11940 2915 11945 2945
rect 11975 2915 11980 2945
rect 11940 2910 11980 2915
rect 12060 2940 12100 2950
rect 12060 2920 12070 2940
rect 12090 2920 12100 2940
rect 12060 2910 12100 2920
rect 12180 2945 12220 2950
rect 12180 2915 12185 2945
rect 12215 2915 12220 2945
rect 12180 2910 12220 2915
rect 12300 2940 12340 2950
rect 12300 2920 12310 2940
rect 12330 2920 12340 2940
rect 12300 2910 12340 2920
rect 12420 2945 12460 2950
rect 12420 2915 12425 2945
rect 12455 2915 12460 2945
rect 12420 2910 12460 2915
rect 12480 2945 12520 2950
rect 12480 2915 12485 2945
rect 12515 2915 12520 2945
rect 12480 2910 12520 2915
rect 13000 2920 13040 2925
rect 13000 2890 13005 2920
rect 13035 2890 13040 2920
rect 13000 2885 13040 2890
rect 13058 2915 13092 2925
rect 13058 2895 13066 2915
rect 13084 2895 13092 2915
rect 13058 2885 13092 2895
rect 13110 2920 13150 2925
rect 13110 2890 13115 2920
rect 13145 2890 13150 2920
rect 13110 2885 13150 2890
rect 13220 2920 13260 2925
rect 13220 2890 13225 2920
rect 13255 2890 13260 2920
rect 13220 2885 13260 2890
rect 13330 2920 13370 2925
rect 13330 2890 13335 2920
rect 13365 2890 13370 2920
rect 13330 2885 13370 2890
rect 13440 2920 13480 2925
rect 13440 2890 13445 2920
rect 13475 2890 13480 2920
rect 13440 2885 13480 2890
rect 13550 2920 13590 2925
rect 13550 2890 13555 2920
rect 13585 2890 13590 2920
rect 13550 2885 13590 2890
rect 13660 2920 13700 2925
rect 13660 2890 13665 2920
rect 13695 2890 13700 2920
rect 13660 2885 13700 2890
rect 13770 2920 13810 2925
rect 13770 2890 13775 2920
rect 13805 2890 13810 2920
rect 13770 2885 13810 2890
rect 13880 2920 13920 2925
rect 13880 2890 13885 2920
rect 13915 2890 13920 2920
rect 13880 2885 13920 2890
rect 13990 2920 14030 2925
rect 13990 2890 13995 2920
rect 14025 2890 14030 2920
rect 13990 2885 14030 2890
rect 13065 2836 13085 2885
rect 13055 2830 13095 2836
rect 13055 2800 13060 2830
rect 13090 2800 13095 2830
rect 13055 2780 13095 2800
rect 13055 2750 13060 2780
rect 13090 2750 13095 2780
rect 12690 2730 12730 2735
rect 12690 2700 12695 2730
rect 12725 2700 12730 2730
rect 12690 2695 12730 2700
rect 13055 2730 13095 2750
rect 13055 2700 13060 2730
rect 13090 2700 13095 2730
rect 13055 2695 13095 2700
rect 10780 2465 10820 2470
rect 10980 2475 11020 2480
rect 9800 2380 9820 2465
rect 10980 2445 10985 2475
rect 11015 2445 11020 2475
rect 10813 2440 10847 2445
rect 10980 2440 11020 2445
rect 11280 2470 11320 2480
rect 11280 2450 11290 2470
rect 11310 2450 11320 2470
rect 11280 2440 11320 2450
rect 11400 2470 11440 2480
rect 11400 2450 11410 2470
rect 11430 2450 11440 2470
rect 11400 2440 11440 2450
rect 11520 2470 11560 2480
rect 11520 2450 11530 2470
rect 11550 2450 11560 2470
rect 11520 2440 11560 2450
rect 11640 2470 11680 2480
rect 11640 2450 11650 2470
rect 11670 2450 11680 2470
rect 11640 2440 11680 2450
rect 11760 2470 11800 2480
rect 11760 2450 11770 2470
rect 11790 2450 11800 2470
rect 11760 2440 11800 2450
rect 11823 2475 11857 2480
rect 11823 2445 11826 2475
rect 11854 2445 11857 2475
rect 11823 2440 11857 2445
rect 11880 2470 11920 2480
rect 11880 2450 11890 2470
rect 11910 2450 11920 2470
rect 11880 2440 11920 2450
rect 12000 2470 12040 2480
rect 12000 2450 12010 2470
rect 12030 2450 12040 2470
rect 12000 2440 12040 2450
rect 12120 2470 12160 2480
rect 12120 2450 12130 2470
rect 12150 2450 12160 2470
rect 12120 2440 12160 2450
rect 12240 2470 12280 2480
rect 12240 2450 12250 2470
rect 12270 2450 12280 2470
rect 12240 2440 12280 2450
rect 12360 2470 12400 2480
rect 12360 2450 12370 2470
rect 12390 2450 12400 2470
rect 12360 2440 12400 2450
rect 12480 2470 12520 2480
rect 12480 2450 12490 2470
rect 12510 2450 12520 2470
rect 12480 2440 12520 2450
rect 10813 2410 10816 2440
rect 10844 2410 10847 2440
rect 11290 2425 11310 2440
rect 10813 2405 10847 2410
rect 11280 2420 11320 2425
rect 9800 2345 9805 2380
rect 9840 2345 9845 2380
rect 10635 2345 10640 2380
rect 10675 2345 10680 2380
rect 10635 2320 10680 2345
rect 9800 2285 9805 2320
rect 9840 2285 9845 2320
rect 10635 2285 10640 2320
rect 10675 2285 10680 2320
rect 10820 2285 10840 2405
rect 11280 2390 11285 2420
rect 11315 2390 11320 2420
rect 11280 2385 11320 2390
rect 11410 2380 11430 2440
rect 11530 2425 11550 2440
rect 11520 2420 11560 2425
rect 11520 2390 11525 2420
rect 11555 2390 11560 2420
rect 11520 2385 11560 2390
rect 11650 2380 11670 2440
rect 11770 2425 11790 2440
rect 11760 2420 11800 2425
rect 11760 2390 11765 2420
rect 11795 2390 11800 2420
rect 11760 2385 11800 2390
rect 11400 2375 11440 2380
rect 11400 2345 11405 2375
rect 11435 2345 11440 2375
rect 11400 2340 11440 2345
rect 11640 2375 11680 2380
rect 11640 2345 11645 2375
rect 11675 2345 11680 2375
rect 11640 2340 11680 2345
rect 9800 2225 9820 2285
rect 10813 2280 10847 2285
rect 10813 2250 10816 2280
rect 10844 2250 10847 2280
rect 10813 2245 10847 2250
rect 11440 2280 11480 2285
rect 11440 2250 11445 2280
rect 11475 2250 11480 2280
rect 11440 2245 11480 2250
rect 11660 2280 11700 2285
rect 11660 2250 11665 2280
rect 11695 2250 11700 2280
rect 11660 2245 11700 2250
rect 11330 2235 11370 2240
rect 9790 2220 9830 2225
rect 9790 2190 9795 2220
rect 9825 2190 9830 2220
rect 9790 2185 9830 2190
rect 9900 2220 9940 2225
rect 9900 2190 9905 2220
rect 9935 2190 9940 2220
rect 9900 2185 9940 2190
rect 10010 2220 10050 2225
rect 10010 2190 10015 2220
rect 10045 2190 10050 2220
rect 10010 2185 10050 2190
rect 10120 2220 10160 2225
rect 10120 2190 10125 2220
rect 10155 2190 10160 2220
rect 10120 2185 10160 2190
rect 10230 2220 10270 2225
rect 10230 2190 10235 2220
rect 10265 2190 10270 2220
rect 10230 2185 10270 2190
rect 10340 2220 10380 2225
rect 10340 2190 10345 2220
rect 10375 2190 10380 2220
rect 10340 2185 10380 2190
rect 10450 2220 10490 2225
rect 10450 2190 10455 2220
rect 10485 2190 10490 2220
rect 10450 2185 10490 2190
rect 10560 2220 10600 2225
rect 10560 2190 10565 2220
rect 10595 2190 10600 2220
rect 10560 2185 10600 2190
rect 10670 2220 10710 2225
rect 10670 2190 10675 2220
rect 10705 2190 10710 2220
rect 10670 2185 10710 2190
rect 10780 2220 10820 2225
rect 10780 2190 10785 2220
rect 10815 2190 10820 2220
rect 11330 2205 11335 2235
rect 11365 2205 11370 2235
rect 11330 2200 11370 2205
rect 10780 2185 10820 2190
rect 11340 2185 11360 2200
rect 11450 2185 11470 2245
rect 11550 2235 11590 2240
rect 11550 2205 11555 2235
rect 11585 2205 11590 2235
rect 11550 2200 11590 2205
rect 11560 2185 11580 2200
rect 11670 2185 11690 2245
rect 11770 2240 11790 2385
rect 11890 2380 11910 2440
rect 12010 2425 12030 2440
rect 12000 2420 12040 2425
rect 12000 2390 12005 2420
rect 12035 2390 12040 2420
rect 12000 2385 12040 2390
rect 12130 2380 12150 2440
rect 12250 2425 12270 2440
rect 12240 2420 12280 2425
rect 12240 2390 12245 2420
rect 12275 2390 12280 2420
rect 12240 2385 12280 2390
rect 12370 2380 12390 2440
rect 12490 2425 12510 2440
rect 12480 2420 12520 2425
rect 12480 2390 12485 2420
rect 12515 2390 12520 2420
rect 12480 2385 12520 2390
rect 12700 2380 12720 2695
rect 12945 2670 12985 2675
rect 12945 2640 12950 2670
rect 12980 2640 12985 2670
rect 12945 2635 12985 2640
rect 13055 2670 13095 2675
rect 13055 2640 13060 2670
rect 13090 2640 13095 2670
rect 13055 2635 13095 2640
rect 13165 2670 13205 2675
rect 13165 2640 13170 2670
rect 13200 2640 13205 2670
rect 13165 2635 13205 2640
rect 13275 2670 13315 2675
rect 13275 2640 13280 2670
rect 13310 2640 13315 2670
rect 13275 2635 13315 2640
rect 13385 2670 13425 2675
rect 13385 2640 13390 2670
rect 13420 2640 13425 2670
rect 13385 2635 13425 2640
rect 13495 2670 13535 2675
rect 13495 2640 13500 2670
rect 13530 2640 13535 2670
rect 13495 2635 13535 2640
rect 13605 2670 13645 2675
rect 13605 2640 13610 2670
rect 13640 2640 13645 2670
rect 13605 2635 13645 2640
rect 13715 2670 13755 2675
rect 13715 2640 13720 2670
rect 13750 2640 13755 2670
rect 13715 2635 13755 2640
rect 13825 2670 13865 2675
rect 13825 2640 13830 2670
rect 13860 2640 13865 2670
rect 13825 2635 13865 2640
rect 13935 2670 13975 2675
rect 13935 2640 13940 2670
rect 13970 2640 13975 2670
rect 13935 2635 13975 2640
rect 14045 2670 14085 2675
rect 14045 2640 14050 2670
rect 14080 2640 14085 2670
rect 14045 2635 14085 2640
rect 17235 2670 17275 2675
rect 17235 2640 17240 2670
rect 17270 2640 17275 2670
rect 17235 2635 17275 2640
rect 17345 2670 17385 2675
rect 17345 2640 17350 2670
rect 17380 2640 17385 2670
rect 17345 2635 17385 2640
rect 17455 2670 17495 2675
rect 17455 2640 17460 2670
rect 17490 2640 17495 2670
rect 17455 2635 17495 2640
rect 17565 2670 17605 2675
rect 17565 2640 17570 2670
rect 17600 2640 17605 2670
rect 17565 2635 17605 2640
rect 17675 2670 17715 2675
rect 17675 2640 17680 2670
rect 17710 2640 17715 2670
rect 17675 2635 17715 2640
rect 17785 2670 17825 2675
rect 17785 2640 17790 2670
rect 17820 2640 17825 2670
rect 17785 2635 17825 2640
rect 17895 2670 17935 2675
rect 17895 2640 17900 2670
rect 17930 2640 17935 2670
rect 17895 2635 17935 2640
rect 18005 2670 18045 2675
rect 18005 2640 18010 2670
rect 18040 2640 18045 2670
rect 18005 2635 18045 2640
rect 18115 2670 18155 2675
rect 18115 2640 18120 2670
rect 18150 2640 18155 2670
rect 18115 2635 18155 2640
rect 18225 2670 18265 2675
rect 18225 2640 18230 2670
rect 18260 2640 18265 2670
rect 18225 2635 18265 2640
rect 18335 2670 18375 2675
rect 18335 2640 18340 2670
rect 18370 2640 18375 2670
rect 18335 2635 18375 2640
rect 13000 2500 13040 2505
rect 13000 2470 13005 2500
rect 13035 2470 13040 2500
rect 13000 2465 13040 2470
rect 13110 2500 13150 2505
rect 13110 2470 13115 2500
rect 13145 2470 13150 2500
rect 13110 2465 13150 2470
rect 13220 2500 13260 2505
rect 13220 2470 13225 2500
rect 13255 2470 13260 2500
rect 13220 2465 13260 2470
rect 13330 2500 13370 2505
rect 13330 2470 13335 2500
rect 13365 2470 13370 2500
rect 13330 2465 13370 2470
rect 13440 2500 13480 2505
rect 13440 2470 13445 2500
rect 13475 2470 13480 2500
rect 13440 2465 13480 2470
rect 13550 2500 13590 2505
rect 13550 2470 13555 2500
rect 13585 2470 13590 2500
rect 13550 2465 13590 2470
rect 13660 2500 13700 2505
rect 13660 2470 13665 2500
rect 13695 2470 13700 2500
rect 13660 2465 13700 2470
rect 13770 2500 13810 2505
rect 13770 2470 13775 2500
rect 13805 2470 13810 2500
rect 13770 2465 13810 2470
rect 13880 2500 13920 2505
rect 13880 2470 13885 2500
rect 13915 2470 13920 2500
rect 13880 2465 13920 2470
rect 13990 2500 14030 2505
rect 13990 2470 13995 2500
rect 14025 2470 14030 2500
rect 13990 2465 14030 2470
rect 17290 2500 17330 2505
rect 17290 2470 17295 2500
rect 17325 2470 17330 2500
rect 17290 2465 17330 2470
rect 17400 2500 17440 2505
rect 17400 2470 17405 2500
rect 17435 2470 17440 2500
rect 17400 2465 17440 2470
rect 17510 2500 17550 2505
rect 17510 2470 17515 2500
rect 17545 2470 17550 2500
rect 17510 2465 17550 2470
rect 17620 2500 17660 2505
rect 17620 2470 17625 2500
rect 17655 2470 17660 2500
rect 17620 2465 17660 2470
rect 17730 2500 17770 2505
rect 17730 2470 17735 2500
rect 17765 2470 17770 2500
rect 17730 2465 17770 2470
rect 17840 2500 17880 2505
rect 17840 2470 17845 2500
rect 17875 2470 17880 2500
rect 17840 2465 17880 2470
rect 17950 2500 17990 2505
rect 17950 2470 17955 2500
rect 17985 2470 17990 2500
rect 17950 2465 17990 2470
rect 18060 2500 18100 2505
rect 18060 2470 18065 2500
rect 18095 2470 18100 2500
rect 18060 2465 18100 2470
rect 18170 2500 18210 2505
rect 18170 2470 18175 2500
rect 18205 2470 18210 2500
rect 18170 2465 18210 2470
rect 18280 2500 18320 2505
rect 18280 2470 18285 2500
rect 18315 2470 18320 2500
rect 18490 2480 18510 3175
rect 18780 3150 18820 3160
rect 18780 3130 18790 3150
rect 18810 3130 18820 3150
rect 18780 3120 18820 3130
rect 18900 3150 18940 3160
rect 18900 3130 18910 3150
rect 18930 3130 18940 3150
rect 18900 3120 18940 3130
rect 19020 3150 19060 3160
rect 19020 3130 19030 3150
rect 19050 3130 19060 3150
rect 19020 3120 19060 3130
rect 19140 3150 19180 3160
rect 19140 3130 19150 3150
rect 19170 3130 19180 3150
rect 19140 3120 19180 3130
rect 19260 3150 19300 3160
rect 19260 3130 19270 3150
rect 19290 3130 19300 3150
rect 19260 3120 19300 3130
rect 19323 3155 19357 3160
rect 19323 3125 19326 3155
rect 19354 3125 19357 3155
rect 19323 3120 19357 3125
rect 19380 3150 19420 3160
rect 19380 3130 19390 3150
rect 19410 3130 19420 3150
rect 19380 3120 19420 3130
rect 19500 3150 19540 3160
rect 19500 3130 19510 3150
rect 19530 3130 19540 3150
rect 19500 3120 19540 3130
rect 19620 3150 19660 3160
rect 19620 3130 19630 3150
rect 19650 3130 19660 3150
rect 19620 3120 19660 3130
rect 19740 3150 19780 3160
rect 19740 3130 19750 3150
rect 19770 3130 19780 3150
rect 19740 3120 19780 3130
rect 19860 3150 19900 3160
rect 19860 3130 19870 3150
rect 19890 3130 19900 3150
rect 19860 3120 19900 3130
rect 19980 3150 20020 3160
rect 19980 3130 19990 3150
rect 20010 3130 20020 3150
rect 19980 3120 20020 3130
rect 18790 3105 18810 3120
rect 18780 3100 18820 3105
rect 18780 3070 18785 3100
rect 18815 3070 18820 3100
rect 18780 3065 18820 3070
rect 18910 3060 18930 3120
rect 19030 3105 19050 3120
rect 19020 3100 19060 3105
rect 19020 3070 19025 3100
rect 19055 3070 19060 3100
rect 19020 3065 19060 3070
rect 19150 3060 19170 3120
rect 19270 3105 19290 3120
rect 19260 3100 19300 3105
rect 19260 3070 19265 3100
rect 19295 3070 19300 3100
rect 19260 3065 19300 3070
rect 19390 3060 19410 3120
rect 19510 3105 19530 3120
rect 19500 3100 19540 3105
rect 19500 3070 19505 3100
rect 19535 3070 19540 3100
rect 19500 3065 19540 3070
rect 19630 3060 19650 3120
rect 19750 3105 19770 3120
rect 19740 3100 19780 3105
rect 19740 3070 19745 3100
rect 19775 3070 19780 3100
rect 19740 3065 19780 3070
rect 19870 3060 19890 3120
rect 19990 3105 20010 3120
rect 19980 3100 20020 3105
rect 19980 3070 19985 3100
rect 20015 3070 20020 3100
rect 19980 3065 20020 3070
rect 18900 3055 18940 3060
rect 18900 3025 18905 3055
rect 18935 3025 18940 3055
rect 18900 3020 18940 3025
rect 19140 3055 19180 3060
rect 19140 3025 19145 3055
rect 19175 3025 19180 3055
rect 19140 3020 19180 3025
rect 19380 3055 19420 3060
rect 19380 3025 19385 3055
rect 19415 3025 19420 3055
rect 19380 3020 19420 3025
rect 19620 3055 19660 3060
rect 19620 3025 19625 3055
rect 19655 3025 19660 3055
rect 19620 3020 19660 3025
rect 19860 3055 19900 3060
rect 19860 3025 19865 3055
rect 19895 3025 19900 3055
rect 19860 3020 19900 3025
rect 18910 3005 18930 3020
rect 18840 3000 18880 3005
rect 18840 2970 18845 3000
rect 18875 2970 18880 3000
rect 18840 2965 18880 2970
rect 18900 3000 18940 3005
rect 18900 2970 18905 3000
rect 18935 2970 18940 3000
rect 18900 2965 18940 2970
rect 19080 3000 19120 3005
rect 19080 2970 19085 3000
rect 19115 2970 19120 3000
rect 19080 2965 19120 2970
rect 19320 3000 19360 3005
rect 19320 2970 19325 3000
rect 19355 2970 19360 3000
rect 19320 2965 19360 2970
rect 19560 3000 19600 3005
rect 19560 2970 19565 3000
rect 19595 2970 19600 3000
rect 19560 2965 19600 2970
rect 19800 3000 19840 3005
rect 19800 2970 19805 3000
rect 19835 2970 19840 3000
rect 19800 2965 19840 2970
rect 18850 2950 18870 2965
rect 19090 2950 19110 2965
rect 19330 2950 19350 2965
rect 19570 2950 19590 2965
rect 19810 2950 19830 2965
rect 19990 2950 20010 3065
rect 18840 2940 18880 2950
rect 18840 2920 18850 2940
rect 18870 2920 18880 2940
rect 18840 2910 18880 2920
rect 18960 2945 19000 2950
rect 18960 2915 18965 2945
rect 18995 2915 19000 2945
rect 18960 2910 19000 2915
rect 19080 2940 19120 2950
rect 19080 2920 19090 2940
rect 19110 2920 19120 2940
rect 19080 2910 19120 2920
rect 19200 2945 19240 2950
rect 19200 2915 19205 2945
rect 19235 2915 19240 2945
rect 19200 2910 19240 2915
rect 19320 2940 19360 2950
rect 19320 2920 19330 2940
rect 19350 2920 19360 2940
rect 19320 2910 19360 2920
rect 19440 2945 19480 2950
rect 19440 2915 19445 2945
rect 19475 2915 19480 2945
rect 19440 2910 19480 2915
rect 19560 2940 19600 2950
rect 19560 2920 19570 2940
rect 19590 2920 19600 2940
rect 19560 2910 19600 2920
rect 19680 2945 19720 2950
rect 19680 2915 19685 2945
rect 19715 2915 19720 2945
rect 19680 2910 19720 2915
rect 19800 2940 19840 2950
rect 19800 2920 19810 2940
rect 19830 2920 19840 2940
rect 19800 2910 19840 2920
rect 19920 2945 19960 2950
rect 19920 2915 19925 2945
rect 19955 2915 19960 2945
rect 19920 2910 19960 2915
rect 19980 2945 20020 2950
rect 19980 2915 19985 2945
rect 20015 2915 20020 2945
rect 19980 2910 20020 2915
rect 20500 2920 20540 2925
rect 20500 2890 20505 2920
rect 20535 2890 20540 2920
rect 20500 2885 20540 2890
rect 20558 2915 20592 2925
rect 20558 2895 20566 2915
rect 20584 2895 20592 2915
rect 20558 2885 20592 2895
rect 20610 2920 20650 2925
rect 20610 2890 20615 2920
rect 20645 2890 20650 2920
rect 20610 2885 20650 2890
rect 20720 2920 20760 2925
rect 20720 2890 20725 2920
rect 20755 2890 20760 2920
rect 20720 2885 20760 2890
rect 20830 2920 20870 2925
rect 20830 2890 20835 2920
rect 20865 2890 20870 2920
rect 20830 2885 20870 2890
rect 20940 2920 20980 2925
rect 20940 2890 20945 2920
rect 20975 2890 20980 2920
rect 20940 2885 20980 2890
rect 21050 2920 21090 2925
rect 21050 2890 21055 2920
rect 21085 2890 21090 2920
rect 21050 2885 21090 2890
rect 21160 2920 21200 2925
rect 21160 2890 21165 2920
rect 21195 2890 21200 2920
rect 21160 2885 21200 2890
rect 21270 2920 21310 2925
rect 21270 2890 21275 2920
rect 21305 2890 21310 2920
rect 21270 2885 21310 2890
rect 21380 2920 21420 2925
rect 21380 2890 21385 2920
rect 21415 2890 21420 2920
rect 21380 2885 21420 2890
rect 21490 2920 21530 2925
rect 21490 2890 21495 2920
rect 21525 2890 21530 2920
rect 21490 2885 21530 2890
rect 20565 2836 20585 2885
rect 20555 2830 20595 2836
rect 20555 2800 20560 2830
rect 20590 2800 20595 2830
rect 20555 2780 20595 2800
rect 20555 2750 20560 2780
rect 20590 2750 20595 2780
rect 20190 2730 20230 2735
rect 20190 2700 20195 2730
rect 20225 2700 20230 2730
rect 20190 2695 20230 2700
rect 20555 2730 20595 2750
rect 20555 2700 20560 2730
rect 20590 2700 20595 2730
rect 20555 2695 20595 2700
rect 18280 2465 18320 2470
rect 18480 2475 18520 2480
rect 12973 2440 13007 2445
rect 12973 2410 12976 2440
rect 13004 2410 13007 2440
rect 12973 2405 13007 2410
rect 12980 2380 13000 2405
rect 14000 2380 14020 2465
rect 11880 2375 11920 2380
rect 11880 2345 11885 2375
rect 11915 2345 11920 2375
rect 11880 2340 11920 2345
rect 12120 2375 12160 2380
rect 12120 2345 12125 2375
rect 12155 2345 12160 2375
rect 12120 2340 12160 2345
rect 12360 2375 12400 2380
rect 12360 2345 12365 2375
rect 12395 2345 12400 2375
rect 12360 2340 12400 2345
rect 12690 2375 12730 2380
rect 12690 2345 12695 2375
rect 12725 2345 12730 2375
rect 12690 2340 12730 2345
rect 12970 2375 13010 2380
rect 12970 2345 12975 2375
rect 13005 2345 13010 2375
rect 12970 2340 13010 2345
rect 13140 2345 13145 2380
rect 13180 2345 13185 2380
rect 13974 2345 13980 2380
rect 14015 2345 14020 2380
rect 17300 2380 17320 2465
rect 18480 2445 18485 2475
rect 18515 2445 18520 2475
rect 18313 2440 18347 2445
rect 18480 2440 18520 2445
rect 18780 2470 18820 2480
rect 18780 2450 18790 2470
rect 18810 2450 18820 2470
rect 18780 2440 18820 2450
rect 18900 2470 18940 2480
rect 18900 2450 18910 2470
rect 18930 2450 18940 2470
rect 18900 2440 18940 2450
rect 19020 2470 19060 2480
rect 19020 2450 19030 2470
rect 19050 2450 19060 2470
rect 19020 2440 19060 2450
rect 19140 2470 19180 2480
rect 19140 2450 19150 2470
rect 19170 2450 19180 2470
rect 19140 2440 19180 2450
rect 19260 2470 19300 2480
rect 19260 2450 19270 2470
rect 19290 2450 19300 2470
rect 19260 2440 19300 2450
rect 19323 2475 19357 2480
rect 19323 2445 19326 2475
rect 19354 2445 19357 2475
rect 19323 2440 19357 2445
rect 19380 2470 19420 2480
rect 19380 2450 19390 2470
rect 19410 2450 19420 2470
rect 19380 2440 19420 2450
rect 19500 2470 19540 2480
rect 19500 2450 19510 2470
rect 19530 2450 19540 2470
rect 19500 2440 19540 2450
rect 19620 2470 19660 2480
rect 19620 2450 19630 2470
rect 19650 2450 19660 2470
rect 19620 2440 19660 2450
rect 19740 2470 19780 2480
rect 19740 2450 19750 2470
rect 19770 2450 19780 2470
rect 19740 2440 19780 2450
rect 19860 2470 19900 2480
rect 19860 2450 19870 2470
rect 19890 2450 19900 2470
rect 19860 2440 19900 2450
rect 19980 2470 20020 2480
rect 19980 2450 19990 2470
rect 20010 2450 20020 2470
rect 19980 2440 20020 2450
rect 18313 2410 18316 2440
rect 18344 2410 18347 2440
rect 18790 2425 18810 2440
rect 18313 2405 18347 2410
rect 18780 2420 18820 2425
rect 17300 2345 17305 2380
rect 17340 2345 17345 2380
rect 18135 2345 18140 2380
rect 18175 2345 18180 2380
rect 12120 2285 12140 2340
rect 12815 2325 12855 2330
rect 12815 2295 12820 2325
rect 12850 2295 12855 2325
rect 12815 2290 12855 2295
rect 11880 2280 11920 2285
rect 11880 2250 11885 2280
rect 11915 2250 11920 2280
rect 11880 2245 11920 2250
rect 12100 2280 12140 2285
rect 12100 2250 12105 2280
rect 12135 2250 12140 2280
rect 12100 2245 12140 2250
rect 12320 2280 12360 2285
rect 12320 2250 12325 2280
rect 12355 2250 12360 2280
rect 12320 2245 12360 2250
rect 11770 2235 11810 2240
rect 11770 2205 11775 2235
rect 11805 2205 11810 2235
rect 11770 2200 11810 2205
rect 11780 2185 11800 2200
rect 11890 2185 11910 2245
rect 11990 2235 12030 2240
rect 11990 2205 11995 2235
rect 12025 2205 12030 2235
rect 11990 2200 12030 2205
rect 12000 2185 12020 2200
rect 12110 2185 12130 2245
rect 12210 2235 12250 2240
rect 12210 2205 12215 2235
rect 12245 2205 12250 2235
rect 12210 2200 12250 2205
rect 12220 2185 12240 2200
rect 12330 2185 12350 2245
rect 12430 2235 12470 2240
rect 12430 2205 12435 2235
rect 12465 2205 12470 2235
rect 12430 2200 12470 2205
rect 12440 2185 12460 2200
rect 11330 2175 11370 2185
rect 11330 2155 11340 2175
rect 11360 2155 11370 2175
rect 11330 2145 11370 2155
rect 11440 2175 11480 2185
rect 11440 2155 11450 2175
rect 11470 2155 11480 2175
rect 11440 2145 11480 2155
rect 11550 2175 11590 2185
rect 11550 2155 11560 2175
rect 11580 2155 11590 2175
rect 11550 2145 11590 2155
rect 11660 2175 11700 2185
rect 11660 2155 11670 2175
rect 11690 2155 11700 2175
rect 11660 2145 11700 2155
rect 11770 2175 11810 2185
rect 11770 2155 11780 2175
rect 11800 2155 11810 2175
rect 11770 2145 11810 2155
rect 11880 2175 11920 2185
rect 11880 2155 11890 2175
rect 11910 2155 11920 2175
rect 11880 2145 11920 2155
rect 11990 2175 12030 2185
rect 11990 2155 12000 2175
rect 12020 2155 12030 2175
rect 11990 2145 12030 2155
rect 12100 2175 12140 2185
rect 12100 2155 12110 2175
rect 12130 2155 12140 2175
rect 12100 2145 12140 2155
rect 12210 2175 12250 2185
rect 12210 2155 12220 2175
rect 12240 2155 12250 2175
rect 12210 2145 12250 2155
rect 12320 2175 12360 2185
rect 12320 2155 12330 2175
rect 12350 2155 12360 2175
rect 12320 2145 12360 2155
rect 12430 2175 12470 2185
rect 12430 2155 12440 2175
rect 12460 2155 12470 2175
rect 12430 2145 12470 2155
rect 9735 2000 9775 2005
rect 9735 1970 9740 2000
rect 9770 1970 9775 2000
rect 9735 1965 9775 1970
rect 9845 2000 9885 2005
rect 9845 1970 9850 2000
rect 9880 1970 9885 2000
rect 9845 1965 9885 1970
rect 9955 2000 9995 2005
rect 9955 1970 9960 2000
rect 9990 1970 9995 2000
rect 9955 1965 9995 1970
rect 10065 2000 10105 2005
rect 10065 1970 10070 2000
rect 10100 1970 10105 2000
rect 10065 1965 10105 1970
rect 10175 2000 10215 2005
rect 10175 1970 10180 2000
rect 10210 1970 10215 2000
rect 10175 1965 10215 1970
rect 10285 2000 10325 2005
rect 10285 1970 10290 2000
rect 10320 1970 10325 2000
rect 10285 1965 10325 1970
rect 10395 2000 10435 2005
rect 10395 1970 10400 2000
rect 10430 1970 10435 2000
rect 10395 1965 10435 1970
rect 10505 2000 10545 2005
rect 10505 1970 10510 2000
rect 10540 1970 10545 2000
rect 10505 1965 10545 1970
rect 10615 2000 10655 2005
rect 10615 1970 10620 2000
rect 10650 1970 10655 2000
rect 10615 1965 10655 1970
rect 10725 2000 10765 2005
rect 10725 1970 10730 2000
rect 10760 1970 10765 2000
rect 10725 1965 10765 1970
rect 10835 2000 10875 2005
rect 10835 1970 10840 2000
rect 10870 1970 10875 2000
rect 10835 1965 10875 1970
rect 11385 1960 11425 1965
rect 11385 1930 11390 1960
rect 11420 1930 11425 1960
rect 11385 1925 11425 1930
rect 11495 1955 11535 1965
rect 11495 1935 11505 1955
rect 11525 1935 11535 1955
rect 11495 1925 11535 1935
rect 11605 1960 11645 1965
rect 11605 1930 11610 1960
rect 11640 1930 11645 1960
rect 11605 1925 11645 1930
rect 11715 1955 11755 1965
rect 11715 1935 11725 1955
rect 11745 1935 11755 1955
rect 11715 1925 11755 1935
rect 11825 1960 11865 1965
rect 11825 1930 11830 1960
rect 11860 1930 11865 1960
rect 11825 1925 11865 1930
rect 11935 1955 11975 1965
rect 11935 1935 11945 1955
rect 11965 1935 11975 1955
rect 11935 1925 11975 1935
rect 12045 1960 12085 1965
rect 12045 1930 12050 1960
rect 12080 1930 12085 1960
rect 12045 1925 12085 1930
rect 12155 1955 12195 1965
rect 12155 1935 12165 1955
rect 12185 1935 12195 1955
rect 12155 1925 12195 1935
rect 12245 1960 12305 1965
rect 12245 1930 12270 1960
rect 12300 1930 12305 1960
rect 12245 1925 12305 1930
rect 12375 1955 12415 1965
rect 12375 1935 12385 1955
rect 12405 1935 12415 1955
rect 12375 1925 12415 1935
rect 11505 1910 11525 1925
rect 11725 1910 11745 1925
rect 11945 1910 11965 1925
rect 12165 1910 12185 1925
rect 11495 1905 11555 1910
rect 11495 1875 11500 1905
rect 11530 1875 11555 1905
rect 11495 1870 11555 1875
rect 11715 1905 11755 1910
rect 11715 1875 11720 1905
rect 11750 1875 11755 1905
rect 11715 1870 11755 1875
rect 11935 1905 11975 1910
rect 11935 1875 11940 1905
rect 11970 1875 11975 1905
rect 11935 1870 11975 1875
rect 12155 1905 12195 1910
rect 12155 1875 12160 1905
rect 12190 1875 12195 1905
rect 12155 1870 12195 1875
rect 11190 1850 11230 1855
rect 11190 1820 11195 1850
rect 11225 1820 11230 1850
rect 11190 1815 11230 1820
rect 11410 1850 11450 1855
rect 11410 1820 11415 1850
rect 11445 1820 11450 1850
rect 11410 1815 11450 1820
rect 11200 1780 11220 1815
rect 11420 1780 11440 1815
rect 11190 1770 11230 1780
rect 11085 1760 11125 1765
rect 11085 1730 11090 1760
rect 11120 1730 11125 1760
rect 11190 1750 11200 1770
rect 11220 1750 11230 1770
rect 11410 1770 11450 1780
rect 11190 1740 11230 1750
rect 11305 1760 11345 1765
rect 11085 1725 11125 1730
rect 11305 1730 11310 1760
rect 11340 1730 11345 1760
rect 11410 1750 11420 1770
rect 11440 1750 11450 1770
rect 11535 1765 11555 1870
rect 12245 1855 12265 1925
rect 12385 1910 12405 1925
rect 12375 1905 12415 1910
rect 12375 1875 12380 1905
rect 12410 1875 12415 1905
rect 12375 1870 12415 1875
rect 11640 1850 11680 1855
rect 11640 1820 11645 1850
rect 11675 1820 11680 1850
rect 11640 1815 11680 1820
rect 12230 1850 12270 1855
rect 12230 1820 12235 1850
rect 12265 1820 12270 1850
rect 12230 1815 12270 1820
rect 12450 1850 12490 1855
rect 12450 1820 12455 1850
rect 12485 1820 12490 1850
rect 12450 1815 12490 1820
rect 12680 1850 12720 1855
rect 12680 1820 12685 1850
rect 12715 1820 12720 1850
rect 12680 1815 12720 1820
rect 11650 1780 11670 1815
rect 11820 1805 11860 1810
rect 11640 1770 11680 1780
rect 11820 1775 11825 1805
rect 11855 1775 11860 1805
rect 11820 1770 11860 1775
rect 11940 1805 11980 1810
rect 11940 1775 11945 1805
rect 11975 1775 11980 1805
rect 12240 1780 12260 1815
rect 12460 1780 12480 1815
rect 12690 1780 12710 1815
rect 11940 1770 11980 1775
rect 12230 1770 12270 1780
rect 11410 1740 11450 1750
rect 11525 1760 11565 1765
rect 11305 1725 11345 1730
rect 11525 1730 11530 1760
rect 11560 1730 11565 1760
rect 11640 1750 11650 1770
rect 11670 1750 11680 1770
rect 11640 1740 11680 1750
rect 11525 1725 11565 1730
rect 11830 1720 11850 1770
rect 11950 1720 11970 1770
rect 12125 1760 12165 1765
rect 12125 1730 12130 1760
rect 12160 1730 12165 1760
rect 12230 1750 12240 1770
rect 12260 1750 12270 1770
rect 12450 1770 12490 1780
rect 12230 1740 12270 1750
rect 12345 1760 12385 1765
rect 12125 1725 12165 1730
rect 12345 1730 12350 1760
rect 12380 1730 12385 1760
rect 12450 1750 12460 1770
rect 12480 1750 12490 1770
rect 12680 1770 12720 1780
rect 12450 1740 12490 1750
rect 12565 1760 12605 1765
rect 12345 1725 12385 1730
rect 12565 1730 12570 1760
rect 12600 1730 12605 1760
rect 12680 1750 12690 1770
rect 12710 1750 12720 1770
rect 12680 1740 12720 1750
rect 12565 1725 12605 1730
rect 11237 1715 11269 1720
rect 11237 1685 11240 1715
rect 11266 1685 11269 1715
rect 11237 1680 11269 1685
rect 11457 1715 11489 1720
rect 11457 1685 11460 1715
rect 11486 1685 11489 1715
rect 11457 1680 11489 1685
rect 11601 1715 11633 1720
rect 11601 1685 11604 1715
rect 11630 1685 11633 1715
rect 11601 1680 11633 1685
rect 11820 1710 11850 1720
rect 11820 1690 11825 1710
rect 11845 1690 11850 1710
rect 11820 1680 11850 1690
rect 11867 1715 11899 1720
rect 11867 1685 11870 1715
rect 11896 1685 11899 1715
rect 11867 1680 11899 1685
rect 11950 1710 11980 1720
rect 11950 1690 11955 1710
rect 11975 1690 11980 1710
rect 11950 1680 11980 1690
rect 12277 1715 12309 1720
rect 12277 1685 12280 1715
rect 12306 1685 12309 1715
rect 12277 1680 12309 1685
rect 12497 1715 12529 1720
rect 12497 1685 12500 1715
rect 12526 1685 12529 1715
rect 12497 1680 12529 1685
rect 12641 1715 12673 1720
rect 12641 1685 12644 1715
rect 12670 1685 12673 1715
rect 12641 1680 12673 1685
rect 4805 1595 4845 1600
rect 4805 1565 4810 1595
rect 4840 1565 4845 1595
rect 4805 1560 4845 1565
rect 5410 1595 5450 1600
rect 5410 1565 5415 1595
rect 5445 1565 5450 1595
rect 12825 1575 12845 2290
rect 12980 2285 13000 2340
rect 13140 2320 13185 2345
rect 18135 2320 18180 2345
rect 13140 2285 13145 2320
rect 13180 2285 13185 2320
rect 13975 2285 13980 2320
rect 14015 2285 14020 2320
rect 12973 2280 13007 2285
rect 12973 2250 12976 2280
rect 13004 2250 13007 2280
rect 12973 2245 13007 2250
rect 14000 2225 14020 2285
rect 17300 2285 17305 2320
rect 17340 2285 17345 2320
rect 18135 2285 18140 2320
rect 18175 2285 18180 2320
rect 18320 2285 18340 2405
rect 18780 2390 18785 2420
rect 18815 2390 18820 2420
rect 18780 2385 18820 2390
rect 18910 2380 18930 2440
rect 19030 2425 19050 2440
rect 19020 2420 19060 2425
rect 19020 2390 19025 2420
rect 19055 2390 19060 2420
rect 19020 2385 19060 2390
rect 19150 2380 19170 2440
rect 19270 2425 19290 2440
rect 19260 2420 19300 2425
rect 19260 2390 19265 2420
rect 19295 2390 19300 2420
rect 19260 2385 19300 2390
rect 18900 2375 18940 2380
rect 18900 2345 18905 2375
rect 18935 2345 18940 2375
rect 18900 2340 18940 2345
rect 19140 2375 19180 2380
rect 19140 2345 19145 2375
rect 19175 2345 19180 2375
rect 19140 2340 19180 2345
rect 17300 2225 17320 2285
rect 18313 2280 18347 2285
rect 18313 2250 18316 2280
rect 18344 2250 18347 2280
rect 18313 2245 18347 2250
rect 18940 2280 18980 2285
rect 18940 2250 18945 2280
rect 18975 2250 18980 2280
rect 18940 2245 18980 2250
rect 19160 2280 19200 2285
rect 19160 2250 19165 2280
rect 19195 2250 19200 2280
rect 19160 2245 19200 2250
rect 18830 2235 18870 2240
rect 13000 2220 13040 2225
rect 13000 2190 13005 2220
rect 13035 2190 13040 2220
rect 13000 2185 13040 2190
rect 13110 2220 13150 2225
rect 13110 2190 13115 2220
rect 13145 2190 13150 2220
rect 13110 2185 13150 2190
rect 13220 2220 13260 2225
rect 13220 2190 13225 2220
rect 13255 2190 13260 2220
rect 13220 2185 13260 2190
rect 13330 2220 13370 2225
rect 13330 2190 13335 2220
rect 13365 2190 13370 2220
rect 13330 2185 13370 2190
rect 13440 2220 13480 2225
rect 13440 2190 13445 2220
rect 13475 2190 13480 2220
rect 13440 2185 13480 2190
rect 13550 2220 13590 2225
rect 13550 2190 13555 2220
rect 13585 2190 13590 2220
rect 13550 2185 13590 2190
rect 13660 2220 13700 2225
rect 13660 2190 13665 2220
rect 13695 2190 13700 2220
rect 13660 2185 13700 2190
rect 13770 2220 13810 2225
rect 13770 2190 13775 2220
rect 13805 2190 13810 2220
rect 13770 2185 13810 2190
rect 13880 2220 13920 2225
rect 13880 2190 13885 2220
rect 13915 2190 13920 2220
rect 13880 2185 13920 2190
rect 13990 2220 14030 2225
rect 13990 2190 13995 2220
rect 14025 2190 14030 2220
rect 13990 2185 14030 2190
rect 17290 2220 17330 2225
rect 17290 2190 17295 2220
rect 17325 2190 17330 2220
rect 17290 2185 17330 2190
rect 17400 2220 17440 2225
rect 17400 2190 17405 2220
rect 17435 2190 17440 2220
rect 17400 2185 17440 2190
rect 17510 2220 17550 2225
rect 17510 2190 17515 2220
rect 17545 2190 17550 2220
rect 17510 2185 17550 2190
rect 17620 2220 17660 2225
rect 17620 2190 17625 2220
rect 17655 2190 17660 2220
rect 17620 2185 17660 2190
rect 17730 2220 17770 2225
rect 17730 2190 17735 2220
rect 17765 2190 17770 2220
rect 17730 2185 17770 2190
rect 17840 2220 17880 2225
rect 17840 2190 17845 2220
rect 17875 2190 17880 2220
rect 17840 2185 17880 2190
rect 17950 2220 17990 2225
rect 17950 2190 17955 2220
rect 17985 2190 17990 2220
rect 17950 2185 17990 2190
rect 18060 2220 18100 2225
rect 18060 2190 18065 2220
rect 18095 2190 18100 2220
rect 18060 2185 18100 2190
rect 18170 2220 18210 2225
rect 18170 2190 18175 2220
rect 18205 2190 18210 2220
rect 18170 2185 18210 2190
rect 18280 2220 18320 2225
rect 18280 2190 18285 2220
rect 18315 2190 18320 2220
rect 18830 2205 18835 2235
rect 18865 2205 18870 2235
rect 18830 2200 18870 2205
rect 18280 2185 18320 2190
rect 18840 2185 18860 2200
rect 18950 2185 18970 2245
rect 19050 2235 19090 2240
rect 19050 2205 19055 2235
rect 19085 2205 19090 2235
rect 19050 2200 19090 2205
rect 19060 2185 19080 2200
rect 19170 2185 19190 2245
rect 19270 2240 19290 2385
rect 19390 2380 19410 2440
rect 19510 2425 19530 2440
rect 19500 2420 19540 2425
rect 19500 2390 19505 2420
rect 19535 2390 19540 2420
rect 19500 2385 19540 2390
rect 19630 2380 19650 2440
rect 19750 2425 19770 2440
rect 19740 2420 19780 2425
rect 19740 2390 19745 2420
rect 19775 2390 19780 2420
rect 19740 2385 19780 2390
rect 19870 2380 19890 2440
rect 19990 2425 20010 2440
rect 19980 2420 20020 2425
rect 19980 2390 19985 2420
rect 20015 2390 20020 2420
rect 19980 2385 20020 2390
rect 20200 2380 20220 2695
rect 20445 2670 20485 2675
rect 20445 2640 20450 2670
rect 20480 2640 20485 2670
rect 20445 2635 20485 2640
rect 20555 2670 20595 2675
rect 20555 2640 20560 2670
rect 20590 2640 20595 2670
rect 20555 2635 20595 2640
rect 20665 2670 20705 2675
rect 20665 2640 20670 2670
rect 20700 2640 20705 2670
rect 20665 2635 20705 2640
rect 20775 2670 20815 2675
rect 20775 2640 20780 2670
rect 20810 2640 20815 2670
rect 20775 2635 20815 2640
rect 20885 2670 20925 2675
rect 20885 2640 20890 2670
rect 20920 2640 20925 2670
rect 20885 2635 20925 2640
rect 20995 2670 21035 2675
rect 20995 2640 21000 2670
rect 21030 2640 21035 2670
rect 20995 2635 21035 2640
rect 21105 2670 21145 2675
rect 21105 2640 21110 2670
rect 21140 2640 21145 2670
rect 21105 2635 21145 2640
rect 21215 2670 21255 2675
rect 21215 2640 21220 2670
rect 21250 2640 21255 2670
rect 21215 2635 21255 2640
rect 21325 2670 21365 2675
rect 21325 2640 21330 2670
rect 21360 2640 21365 2670
rect 21325 2635 21365 2640
rect 21435 2670 21475 2675
rect 21435 2640 21440 2670
rect 21470 2640 21475 2670
rect 21435 2635 21475 2640
rect 21545 2670 21585 2675
rect 21545 2640 21550 2670
rect 21580 2640 21585 2670
rect 21545 2635 21585 2640
rect 20500 2500 20540 2505
rect 20500 2470 20505 2500
rect 20535 2470 20540 2500
rect 20500 2465 20540 2470
rect 20610 2500 20650 2505
rect 20610 2470 20615 2500
rect 20645 2470 20650 2500
rect 20610 2465 20650 2470
rect 20720 2500 20760 2505
rect 20720 2470 20725 2500
rect 20755 2470 20760 2500
rect 20720 2465 20760 2470
rect 20830 2500 20870 2505
rect 20830 2470 20835 2500
rect 20865 2470 20870 2500
rect 20830 2465 20870 2470
rect 20940 2500 20980 2505
rect 20940 2470 20945 2500
rect 20975 2470 20980 2500
rect 20940 2465 20980 2470
rect 21050 2500 21090 2505
rect 21050 2470 21055 2500
rect 21085 2470 21090 2500
rect 21050 2465 21090 2470
rect 21160 2500 21200 2505
rect 21160 2470 21165 2500
rect 21195 2470 21200 2500
rect 21160 2465 21200 2470
rect 21270 2500 21310 2505
rect 21270 2470 21275 2500
rect 21305 2470 21310 2500
rect 21270 2465 21310 2470
rect 21380 2500 21420 2505
rect 21380 2470 21385 2500
rect 21415 2470 21420 2500
rect 21380 2465 21420 2470
rect 21490 2500 21530 2505
rect 21490 2470 21495 2500
rect 21525 2470 21530 2500
rect 21490 2465 21530 2470
rect 20473 2440 20507 2445
rect 20473 2410 20476 2440
rect 20504 2410 20507 2440
rect 20473 2405 20507 2410
rect 20480 2380 20500 2405
rect 21500 2380 21520 2465
rect 19380 2375 19420 2380
rect 19380 2345 19385 2375
rect 19415 2345 19420 2375
rect 19380 2340 19420 2345
rect 19620 2375 19660 2380
rect 19620 2345 19625 2375
rect 19655 2345 19660 2375
rect 19620 2340 19660 2345
rect 19860 2375 19900 2380
rect 19860 2345 19865 2375
rect 19895 2345 19900 2375
rect 19860 2340 19900 2345
rect 20190 2375 20230 2380
rect 20190 2345 20195 2375
rect 20225 2345 20230 2375
rect 20190 2340 20230 2345
rect 20470 2375 20510 2380
rect 20470 2345 20475 2375
rect 20505 2345 20510 2375
rect 20470 2340 20510 2345
rect 20640 2345 20645 2380
rect 20680 2345 20685 2380
rect 21474 2345 21480 2380
rect 21515 2345 21520 2380
rect 19620 2285 19640 2340
rect 20315 2325 20355 2330
rect 20315 2295 20320 2325
rect 20350 2295 20355 2325
rect 20315 2290 20355 2295
rect 19380 2280 19420 2285
rect 19380 2250 19385 2280
rect 19415 2250 19420 2280
rect 19380 2245 19420 2250
rect 19600 2280 19640 2285
rect 19600 2250 19605 2280
rect 19635 2250 19640 2280
rect 19600 2245 19640 2250
rect 19820 2280 19860 2285
rect 19820 2250 19825 2280
rect 19855 2250 19860 2280
rect 19820 2245 19860 2250
rect 19270 2235 19310 2240
rect 19270 2205 19275 2235
rect 19305 2205 19310 2235
rect 19270 2200 19310 2205
rect 19280 2185 19300 2200
rect 19390 2185 19410 2245
rect 19490 2235 19530 2240
rect 19490 2205 19495 2235
rect 19525 2205 19530 2235
rect 19490 2200 19530 2205
rect 19500 2185 19520 2200
rect 19610 2185 19630 2245
rect 19710 2235 19750 2240
rect 19710 2205 19715 2235
rect 19745 2205 19750 2235
rect 19710 2200 19750 2205
rect 19720 2185 19740 2200
rect 19830 2185 19850 2245
rect 19930 2235 19970 2240
rect 19930 2205 19935 2235
rect 19965 2205 19970 2235
rect 19930 2200 19970 2205
rect 19940 2185 19960 2200
rect 18830 2175 18870 2185
rect 18830 2155 18840 2175
rect 18860 2155 18870 2175
rect 18830 2145 18870 2155
rect 18940 2175 18980 2185
rect 18940 2155 18950 2175
rect 18970 2155 18980 2175
rect 18940 2145 18980 2155
rect 19050 2175 19090 2185
rect 19050 2155 19060 2175
rect 19080 2155 19090 2175
rect 19050 2145 19090 2155
rect 19160 2175 19200 2185
rect 19160 2155 19170 2175
rect 19190 2155 19200 2175
rect 19160 2145 19200 2155
rect 19270 2175 19310 2185
rect 19270 2155 19280 2175
rect 19300 2155 19310 2175
rect 19270 2145 19310 2155
rect 19380 2175 19420 2185
rect 19380 2155 19390 2175
rect 19410 2155 19420 2175
rect 19380 2145 19420 2155
rect 19490 2175 19530 2185
rect 19490 2155 19500 2175
rect 19520 2155 19530 2175
rect 19490 2145 19530 2155
rect 19600 2175 19640 2185
rect 19600 2155 19610 2175
rect 19630 2155 19640 2175
rect 19600 2145 19640 2155
rect 19710 2175 19750 2185
rect 19710 2155 19720 2175
rect 19740 2155 19750 2175
rect 19710 2145 19750 2155
rect 19820 2175 19860 2185
rect 19820 2155 19830 2175
rect 19850 2155 19860 2175
rect 19820 2145 19860 2155
rect 19930 2175 19970 2185
rect 19930 2155 19940 2175
rect 19960 2155 19970 2175
rect 19930 2145 19970 2155
rect 12945 2000 12985 2005
rect 12945 1970 12950 2000
rect 12980 1970 12985 2000
rect 12945 1965 12985 1970
rect 13055 2000 13095 2005
rect 13055 1970 13060 2000
rect 13090 1970 13095 2000
rect 13055 1965 13095 1970
rect 13165 2000 13205 2005
rect 13165 1970 13170 2000
rect 13200 1970 13205 2000
rect 13165 1965 13205 1970
rect 13275 2000 13315 2005
rect 13275 1970 13280 2000
rect 13310 1970 13315 2000
rect 13275 1965 13315 1970
rect 13385 2000 13425 2005
rect 13385 1970 13390 2000
rect 13420 1970 13425 2000
rect 13385 1965 13425 1970
rect 13495 2000 13535 2005
rect 13495 1970 13500 2000
rect 13530 1970 13535 2000
rect 13495 1965 13535 1970
rect 13605 2000 13645 2005
rect 13605 1970 13610 2000
rect 13640 1970 13645 2000
rect 13605 1965 13645 1970
rect 13715 2000 13755 2005
rect 13715 1970 13720 2000
rect 13750 1970 13755 2000
rect 13715 1965 13755 1970
rect 13825 2000 13865 2005
rect 13825 1970 13830 2000
rect 13860 1970 13865 2000
rect 13825 1965 13865 1970
rect 13935 2000 13975 2005
rect 13935 1970 13940 2000
rect 13970 1970 13975 2000
rect 13935 1965 13975 1970
rect 14045 2000 14085 2005
rect 14045 1970 14050 2000
rect 14080 1970 14085 2000
rect 14045 1965 14085 1970
rect 17235 2000 17275 2005
rect 17235 1970 17240 2000
rect 17270 1970 17275 2000
rect 17235 1965 17275 1970
rect 17345 2000 17385 2005
rect 17345 1970 17350 2000
rect 17380 1970 17385 2000
rect 17345 1965 17385 1970
rect 17455 2000 17495 2005
rect 17455 1970 17460 2000
rect 17490 1970 17495 2000
rect 17455 1965 17495 1970
rect 17565 2000 17605 2005
rect 17565 1970 17570 2000
rect 17600 1970 17605 2000
rect 17565 1965 17605 1970
rect 17675 2000 17715 2005
rect 17675 1970 17680 2000
rect 17710 1970 17715 2000
rect 17675 1965 17715 1970
rect 17785 2000 17825 2005
rect 17785 1970 17790 2000
rect 17820 1970 17825 2000
rect 17785 1965 17825 1970
rect 17895 2000 17935 2005
rect 17895 1970 17900 2000
rect 17930 1970 17935 2000
rect 17895 1965 17935 1970
rect 18005 2000 18045 2005
rect 18005 1970 18010 2000
rect 18040 1970 18045 2000
rect 18005 1965 18045 1970
rect 18115 2000 18155 2005
rect 18115 1970 18120 2000
rect 18150 1970 18155 2000
rect 18115 1965 18155 1970
rect 18225 2000 18265 2005
rect 18225 1970 18230 2000
rect 18260 1970 18265 2000
rect 18225 1965 18265 1970
rect 18335 2000 18375 2005
rect 18335 1970 18340 2000
rect 18370 1970 18375 2000
rect 18335 1965 18375 1970
rect 18885 1960 18925 1965
rect 18885 1930 18890 1960
rect 18920 1930 18925 1960
rect 18885 1925 18925 1930
rect 18995 1955 19035 1965
rect 18995 1935 19005 1955
rect 19025 1935 19035 1955
rect 18995 1925 19035 1935
rect 19105 1960 19145 1965
rect 19105 1930 19110 1960
rect 19140 1930 19145 1960
rect 19105 1925 19145 1930
rect 19215 1955 19255 1965
rect 19215 1935 19225 1955
rect 19245 1935 19255 1955
rect 19215 1925 19255 1935
rect 19325 1960 19365 1965
rect 19325 1930 19330 1960
rect 19360 1930 19365 1960
rect 19325 1925 19365 1930
rect 19435 1955 19475 1965
rect 19435 1935 19445 1955
rect 19465 1935 19475 1955
rect 19435 1925 19475 1935
rect 19545 1960 19585 1965
rect 19545 1930 19550 1960
rect 19580 1930 19585 1960
rect 19545 1925 19585 1930
rect 19655 1955 19695 1965
rect 19655 1935 19665 1955
rect 19685 1935 19695 1955
rect 19655 1925 19695 1935
rect 19745 1960 19805 1965
rect 19745 1930 19770 1960
rect 19800 1930 19805 1960
rect 19745 1925 19805 1930
rect 19875 1955 19915 1965
rect 19875 1935 19885 1955
rect 19905 1935 19915 1955
rect 19875 1925 19915 1935
rect 19005 1910 19025 1925
rect 19225 1910 19245 1925
rect 19445 1910 19465 1925
rect 19665 1910 19685 1925
rect 18995 1905 19055 1910
rect 18995 1875 19000 1905
rect 19030 1875 19055 1905
rect 18995 1870 19055 1875
rect 19215 1905 19255 1910
rect 19215 1875 19220 1905
rect 19250 1875 19255 1905
rect 19215 1870 19255 1875
rect 19435 1905 19475 1910
rect 19435 1875 19440 1905
rect 19470 1875 19475 1905
rect 19435 1870 19475 1875
rect 19655 1905 19695 1910
rect 19655 1875 19660 1905
rect 19690 1875 19695 1905
rect 19655 1870 19695 1875
rect 18690 1850 18730 1855
rect 18690 1820 18695 1850
rect 18725 1820 18730 1850
rect 18690 1815 18730 1820
rect 18910 1850 18950 1855
rect 18910 1820 18915 1850
rect 18945 1820 18950 1850
rect 18910 1815 18950 1820
rect 18700 1780 18720 1815
rect 18920 1780 18940 1815
rect 18690 1770 18730 1780
rect 18585 1760 18625 1765
rect 18585 1730 18590 1760
rect 18620 1730 18625 1760
rect 18690 1750 18700 1770
rect 18720 1750 18730 1770
rect 18910 1770 18950 1780
rect 18690 1740 18730 1750
rect 18805 1760 18845 1765
rect 18585 1725 18625 1730
rect 18805 1730 18810 1760
rect 18840 1730 18845 1760
rect 18910 1750 18920 1770
rect 18940 1750 18950 1770
rect 19035 1765 19055 1870
rect 19745 1855 19765 1925
rect 19885 1910 19905 1925
rect 19875 1905 19915 1910
rect 19875 1875 19880 1905
rect 19910 1875 19915 1905
rect 19875 1870 19915 1875
rect 19140 1850 19180 1855
rect 19140 1820 19145 1850
rect 19175 1820 19180 1850
rect 19140 1815 19180 1820
rect 19730 1850 19770 1855
rect 19730 1820 19735 1850
rect 19765 1820 19770 1850
rect 19730 1815 19770 1820
rect 19950 1850 19990 1855
rect 19950 1820 19955 1850
rect 19985 1820 19990 1850
rect 19950 1815 19990 1820
rect 20180 1850 20220 1855
rect 20180 1820 20185 1850
rect 20215 1820 20220 1850
rect 20180 1815 20220 1820
rect 19150 1780 19170 1815
rect 19320 1805 19360 1810
rect 19140 1770 19180 1780
rect 19320 1775 19325 1805
rect 19355 1775 19360 1805
rect 19320 1770 19360 1775
rect 19440 1805 19480 1810
rect 19440 1775 19445 1805
rect 19475 1775 19480 1805
rect 19740 1780 19760 1815
rect 19960 1780 19980 1815
rect 20190 1780 20210 1815
rect 19440 1770 19480 1775
rect 19730 1770 19770 1780
rect 18910 1740 18950 1750
rect 19025 1760 19065 1765
rect 18805 1725 18845 1730
rect 19025 1730 19030 1760
rect 19060 1730 19065 1760
rect 19140 1750 19150 1770
rect 19170 1750 19180 1770
rect 19140 1740 19180 1750
rect 19025 1725 19065 1730
rect 19330 1720 19350 1770
rect 19450 1720 19470 1770
rect 19625 1760 19665 1765
rect 19625 1730 19630 1760
rect 19660 1730 19665 1760
rect 19730 1750 19740 1770
rect 19760 1750 19770 1770
rect 19950 1770 19990 1780
rect 19730 1740 19770 1750
rect 19845 1760 19885 1765
rect 19625 1725 19665 1730
rect 19845 1730 19850 1760
rect 19880 1730 19885 1760
rect 19950 1750 19960 1770
rect 19980 1750 19990 1770
rect 20180 1770 20220 1780
rect 19950 1740 19990 1750
rect 20065 1760 20105 1765
rect 19845 1725 19885 1730
rect 20065 1730 20070 1760
rect 20100 1730 20105 1760
rect 20180 1750 20190 1770
rect 20210 1750 20220 1770
rect 20180 1740 20220 1750
rect 20065 1725 20105 1730
rect 18737 1715 18769 1720
rect 18737 1685 18740 1715
rect 18766 1685 18769 1715
rect 18737 1680 18769 1685
rect 18957 1715 18989 1720
rect 18957 1685 18960 1715
rect 18986 1685 18989 1715
rect 18957 1680 18989 1685
rect 19101 1715 19133 1720
rect 19101 1685 19104 1715
rect 19130 1685 19133 1715
rect 19101 1680 19133 1685
rect 19320 1710 19350 1720
rect 19320 1690 19325 1710
rect 19345 1690 19350 1710
rect 19320 1680 19350 1690
rect 19367 1715 19399 1720
rect 19367 1685 19370 1715
rect 19396 1685 19399 1715
rect 19367 1680 19399 1685
rect 19450 1710 19480 1720
rect 19450 1690 19455 1710
rect 19475 1690 19480 1710
rect 19450 1680 19480 1690
rect 19777 1715 19809 1720
rect 19777 1685 19780 1715
rect 19806 1685 19809 1715
rect 19777 1680 19809 1685
rect 19997 1715 20029 1720
rect 19997 1685 20000 1715
rect 20026 1685 20029 1715
rect 19997 1680 20029 1685
rect 20141 1715 20173 1720
rect 20141 1685 20144 1715
rect 20170 1685 20173 1715
rect 20141 1680 20173 1685
rect 20325 1575 20345 2290
rect 20480 2285 20500 2340
rect 20640 2320 20685 2345
rect 20640 2285 20645 2320
rect 20680 2285 20685 2320
rect 21475 2285 21480 2320
rect 21515 2285 21520 2320
rect 20473 2280 20507 2285
rect 20473 2250 20476 2280
rect 20504 2250 20507 2280
rect 20473 2245 20507 2250
rect 21500 2225 21520 2285
rect 20500 2220 20540 2225
rect 20500 2190 20505 2220
rect 20535 2190 20540 2220
rect 20500 2185 20540 2190
rect 20610 2220 20650 2225
rect 20610 2190 20615 2220
rect 20645 2190 20650 2220
rect 20610 2185 20650 2190
rect 20720 2220 20760 2225
rect 20720 2190 20725 2220
rect 20755 2190 20760 2220
rect 20720 2185 20760 2190
rect 20830 2220 20870 2225
rect 20830 2190 20835 2220
rect 20865 2190 20870 2220
rect 20830 2185 20870 2190
rect 20940 2220 20980 2225
rect 20940 2190 20945 2220
rect 20975 2190 20980 2220
rect 20940 2185 20980 2190
rect 21050 2220 21090 2225
rect 21050 2190 21055 2220
rect 21085 2190 21090 2220
rect 21050 2185 21090 2190
rect 21160 2220 21200 2225
rect 21160 2190 21165 2220
rect 21195 2190 21200 2220
rect 21160 2185 21200 2190
rect 21270 2220 21310 2225
rect 21270 2190 21275 2220
rect 21305 2190 21310 2220
rect 21270 2185 21310 2190
rect 21380 2220 21420 2225
rect 21380 2190 21385 2220
rect 21415 2190 21420 2220
rect 21380 2185 21420 2190
rect 21490 2220 21530 2225
rect 21490 2190 21495 2220
rect 21525 2190 21530 2220
rect 21490 2185 21530 2190
rect 20445 2000 20485 2005
rect 20445 1970 20450 2000
rect 20480 1970 20485 2000
rect 20445 1965 20485 1970
rect 20555 2000 20595 2005
rect 20555 1970 20560 2000
rect 20590 1970 20595 2000
rect 20555 1965 20595 1970
rect 20665 2000 20705 2005
rect 20665 1970 20670 2000
rect 20700 1970 20705 2000
rect 20665 1965 20705 1970
rect 20775 2000 20815 2005
rect 20775 1970 20780 2000
rect 20810 1970 20815 2000
rect 20775 1965 20815 1970
rect 20885 2000 20925 2005
rect 20885 1970 20890 2000
rect 20920 1970 20925 2000
rect 20885 1965 20925 1970
rect 20995 2000 21035 2005
rect 20995 1970 21000 2000
rect 21030 1970 21035 2000
rect 20995 1965 21035 1970
rect 21105 2000 21145 2005
rect 21105 1970 21110 2000
rect 21140 1970 21145 2000
rect 21105 1965 21145 1970
rect 21215 2000 21255 2005
rect 21215 1970 21220 2000
rect 21250 1970 21255 2000
rect 21215 1965 21255 1970
rect 21325 2000 21365 2005
rect 21325 1970 21330 2000
rect 21360 1970 21365 2000
rect 21325 1965 21365 1970
rect 21435 2000 21475 2005
rect 21435 1970 21440 2000
rect 21470 1970 21475 2000
rect 21435 1965 21475 1970
rect 21545 2000 21585 2005
rect 21545 1970 21550 2000
rect 21580 1970 21585 2000
rect 21545 1965 21585 1970
rect 20545 1905 20585 1910
rect 20545 1875 20550 1905
rect 20580 1875 20585 1905
rect 20545 1870 20585 1875
rect 20655 1905 20695 1910
rect 20655 1875 20660 1905
rect 20690 1875 20695 1905
rect 20655 1870 20695 1875
rect 20765 1905 20805 1910
rect 20765 1875 20770 1905
rect 20800 1875 20805 1905
rect 20765 1870 20805 1875
rect 20566 1680 20598 1685
rect 20566 1650 20570 1680
rect 20596 1650 20598 1680
rect 20615 1680 20655 1690
rect 20615 1660 20625 1680
rect 20645 1660 20655 1680
rect 20615 1650 20655 1660
rect 20710 1680 20750 1690
rect 20710 1660 20720 1680
rect 20740 1660 20750 1680
rect 20710 1650 20750 1660
rect 20566 1645 20598 1650
rect 20510 1630 20550 1635
rect 20510 1600 20515 1630
rect 20545 1600 20550 1630
rect 20510 1595 20550 1600
rect 20570 1575 20590 1645
rect 20625 1635 20645 1650
rect 20720 1635 20740 1650
rect 20616 1630 20656 1635
rect 20616 1600 20621 1630
rect 20651 1600 20656 1630
rect 20616 1595 20656 1600
rect 20710 1630 20750 1635
rect 20710 1600 20715 1630
rect 20745 1600 20750 1630
rect 20710 1595 20750 1600
rect 20800 1630 20840 1635
rect 20800 1600 20805 1630
rect 20835 1600 20840 1630
rect 20800 1595 20840 1600
rect 5410 1560 5450 1565
rect 12815 1570 12855 1575
rect 4265 1545 4305 1550
rect 4265 1515 4270 1545
rect 4300 1515 4305 1545
rect 4265 1510 4305 1515
rect 4385 1545 4425 1550
rect 4385 1515 4390 1545
rect 4420 1515 4425 1545
rect 4385 1510 4425 1515
rect 4505 1545 4545 1550
rect 4505 1515 4510 1545
rect 4540 1515 4545 1545
rect 4505 1510 4545 1515
rect 4625 1545 4665 1550
rect 4625 1515 4630 1545
rect 4660 1515 4665 1545
rect 4625 1510 4665 1515
rect 4745 1545 4785 1550
rect 4745 1515 4750 1545
rect 4780 1515 4785 1545
rect 4745 1510 4785 1515
rect 5135 1545 5175 1550
rect 5135 1515 5140 1545
rect 5170 1515 5175 1545
rect 12815 1540 12820 1570
rect 12850 1540 12855 1570
rect 12815 1535 12855 1540
rect 20315 1570 20355 1575
rect 20315 1540 20320 1570
rect 20350 1540 20355 1570
rect 20315 1535 20355 1540
rect 20471 1570 20503 1575
rect 20471 1540 20475 1570
rect 20501 1540 20503 1570
rect 20471 1535 20503 1540
rect 20560 1565 20600 1575
rect 20560 1545 20570 1565
rect 20590 1545 20600 1565
rect 20560 1535 20600 1545
rect 20847 1570 20879 1575
rect 20847 1540 20849 1570
rect 20875 1540 20879 1570
rect 20847 1535 20879 1540
rect 5135 1510 5175 1515
rect 4205 1500 4245 1505
rect 4055 1480 4095 1490
rect 4055 1460 4065 1480
rect 4085 1460 4095 1480
rect 4205 1470 4210 1500
rect 4240 1470 4245 1500
rect 4205 1465 4245 1470
rect 4325 1500 4365 1505
rect 4325 1470 4330 1500
rect 4360 1470 4365 1500
rect 4325 1465 4365 1470
rect 4445 1500 4485 1505
rect 4445 1470 4450 1500
rect 4480 1470 4485 1500
rect 4445 1465 4485 1470
rect 4685 1500 4725 1505
rect 4685 1470 4690 1500
rect 4720 1470 4725 1500
rect 4685 1465 4725 1470
rect 4805 1500 4845 1505
rect 4805 1470 4810 1500
rect 4840 1470 4845 1500
rect 4805 1465 4845 1470
rect 4925 1500 4965 1505
rect 4925 1470 4930 1500
rect 4960 1470 4965 1500
rect 4925 1465 4965 1470
rect 5045 1500 5085 1505
rect 5045 1470 5050 1500
rect 5080 1470 5085 1500
rect 5145 1490 5165 1510
rect 11106 1495 11138 1500
rect 5045 1465 5085 1470
rect 5135 1480 5175 1490
rect 4055 1450 4095 1460
rect 5135 1460 5145 1480
rect 5165 1460 5175 1480
rect 11106 1465 11109 1495
rect 11135 1465 11138 1495
rect 11106 1460 11138 1465
rect 11305 1495 11345 1500
rect 11305 1465 11310 1495
rect 11340 1465 11345 1495
rect 11305 1460 11345 1465
rect 11525 1495 11565 1500
rect 11525 1465 11530 1495
rect 11560 1465 11565 1495
rect 11525 1460 11565 1465
rect 11825 1490 11855 1500
rect 11825 1470 11830 1490
rect 11850 1470 11855 1490
rect 11825 1460 11855 1470
rect 11875 1490 11905 1500
rect 11875 1470 11880 1490
rect 11900 1470 11905 1490
rect 11875 1460 11905 1470
rect 11922 1495 11954 1500
rect 11922 1465 11925 1495
rect 11951 1465 11954 1495
rect 11922 1460 11954 1465
rect 12146 1495 12178 1500
rect 12146 1465 12149 1495
rect 12175 1465 12178 1495
rect 12146 1460 12178 1465
rect 12345 1495 12385 1500
rect 12345 1465 12350 1495
rect 12380 1465 12385 1495
rect 12345 1460 12385 1465
rect 12565 1495 12605 1500
rect 12565 1465 12570 1495
rect 12600 1465 12605 1495
rect 12565 1460 12605 1465
rect 18606 1495 18638 1500
rect 18606 1465 18609 1495
rect 18635 1465 18638 1495
rect 18606 1460 18638 1465
rect 18805 1495 18845 1500
rect 18805 1465 18810 1495
rect 18840 1465 18845 1495
rect 18805 1460 18845 1465
rect 19025 1495 19065 1500
rect 19025 1465 19030 1495
rect 19060 1465 19065 1495
rect 19025 1460 19065 1465
rect 19325 1490 19355 1500
rect 19325 1470 19330 1490
rect 19350 1470 19355 1490
rect 19325 1460 19355 1470
rect 19375 1490 19405 1500
rect 19375 1470 19380 1490
rect 19400 1470 19405 1490
rect 19375 1460 19405 1470
rect 19422 1495 19454 1500
rect 19422 1465 19425 1495
rect 19451 1465 19454 1495
rect 19422 1460 19454 1465
rect 19646 1495 19678 1500
rect 19646 1465 19649 1495
rect 19675 1465 19678 1495
rect 19646 1460 19678 1465
rect 19845 1495 19885 1500
rect 19845 1465 19850 1495
rect 19880 1465 19885 1495
rect 19845 1460 19885 1465
rect 20065 1495 20105 1500
rect 20065 1465 20070 1495
rect 20100 1465 20105 1495
rect 20065 1460 20105 1465
rect 5135 1450 5175 1460
rect 11145 1435 11185 1440
rect 11145 1405 11150 1435
rect 11180 1405 11185 1435
rect 11145 1400 11185 1405
rect 11250 1435 11290 1440
rect 11250 1405 11255 1435
rect 11285 1405 11290 1435
rect 11250 1400 11290 1405
rect 11360 1435 11400 1440
rect 11360 1405 11365 1435
rect 11395 1405 11400 1435
rect 11360 1400 11400 1405
rect 11470 1435 11510 1440
rect 11470 1405 11475 1435
rect 11505 1405 11510 1435
rect 11470 1400 11510 1405
rect 11580 1435 11620 1440
rect 11580 1405 11585 1435
rect 11615 1405 11620 1435
rect 11580 1400 11620 1405
rect 11830 1340 11850 1460
rect 11810 1335 11850 1340
rect 11810 1305 11815 1335
rect 11845 1305 11850 1335
rect 11810 1300 11850 1305
rect 11315 1285 11355 1290
rect 11315 1255 11320 1285
rect 11350 1255 11355 1285
rect 11315 1250 11355 1255
rect 11325 1230 11345 1250
rect 11820 1230 11840 1300
rect 11880 1290 11900 1460
rect 12185 1435 12225 1440
rect 12185 1405 12190 1435
rect 12220 1405 12225 1435
rect 12185 1400 12225 1405
rect 12290 1435 12330 1440
rect 12290 1405 12295 1435
rect 12325 1405 12330 1435
rect 12290 1400 12330 1405
rect 12400 1435 12440 1440
rect 12400 1405 12405 1435
rect 12435 1405 12440 1435
rect 12400 1400 12440 1405
rect 12510 1435 12550 1440
rect 12510 1405 12515 1435
rect 12545 1405 12550 1435
rect 12510 1400 12550 1405
rect 12620 1435 12660 1440
rect 12620 1405 12625 1435
rect 12655 1405 12660 1435
rect 18645 1435 18685 1440
rect 12620 1400 12660 1405
rect 13015 1395 13020 1430
rect 13055 1395 13060 1430
rect 14025 1395 14030 1430
rect 14065 1395 14070 1430
rect 18645 1405 18650 1435
rect 18680 1405 18685 1435
rect 18645 1400 18685 1405
rect 18750 1435 18790 1440
rect 18750 1405 18755 1435
rect 18785 1405 18790 1435
rect 18750 1400 18790 1405
rect 18860 1435 18900 1440
rect 18860 1405 18865 1435
rect 18895 1405 18900 1435
rect 18860 1400 18900 1405
rect 18970 1435 19010 1440
rect 18970 1405 18975 1435
rect 19005 1405 19010 1435
rect 18970 1400 19010 1405
rect 19080 1435 19120 1440
rect 19080 1405 19085 1435
rect 19115 1405 19120 1435
rect 19080 1400 19120 1405
rect 13030 1380 13050 1395
rect 13020 1375 13060 1380
rect 13020 1345 13025 1375
rect 13055 1345 13060 1375
rect 13020 1340 13060 1345
rect 13125 1375 13165 1380
rect 13125 1345 13130 1375
rect 13160 1345 13165 1375
rect 13125 1340 13165 1345
rect 13135 1325 13155 1340
rect 14035 1325 14055 1395
rect 19330 1390 19350 1460
rect 19310 1385 19350 1390
rect 19310 1355 19315 1385
rect 19345 1355 19350 1385
rect 19310 1350 19350 1355
rect 18815 1335 18855 1340
rect 13025 1320 13065 1325
rect 13025 1290 13030 1320
rect 13060 1290 13065 1320
rect 11880 1285 11920 1290
rect 13025 1285 13065 1290
rect 13128 1315 13162 1325
rect 13128 1295 13136 1315
rect 13154 1295 13162 1315
rect 13128 1285 13162 1295
rect 13225 1320 13265 1325
rect 13225 1290 13230 1320
rect 13260 1290 13265 1320
rect 13225 1285 13265 1290
rect 13425 1320 13465 1325
rect 13425 1290 13430 1320
rect 13460 1290 13465 1320
rect 13425 1285 13465 1290
rect 13625 1320 13665 1325
rect 13625 1290 13630 1320
rect 13660 1290 13665 1320
rect 13625 1285 13665 1290
rect 13825 1320 13865 1325
rect 13825 1290 13830 1320
rect 13860 1290 13865 1320
rect 13825 1285 13865 1290
rect 14025 1320 14065 1325
rect 14025 1290 14030 1320
rect 14060 1290 14065 1320
rect 18815 1305 18820 1335
rect 18850 1305 18855 1335
rect 18815 1300 18855 1305
rect 14025 1285 14065 1290
rect 11880 1255 11885 1285
rect 11915 1255 11920 1285
rect 18825 1280 18845 1300
rect 19320 1280 19340 1350
rect 19380 1340 19400 1460
rect 19685 1435 19725 1440
rect 19685 1405 19690 1435
rect 19720 1405 19725 1435
rect 19685 1400 19725 1405
rect 19790 1435 19830 1440
rect 19790 1405 19795 1435
rect 19825 1405 19830 1435
rect 19790 1400 19830 1405
rect 19900 1435 19940 1440
rect 19900 1405 19905 1435
rect 19935 1405 19940 1435
rect 19900 1400 19940 1405
rect 20010 1435 20050 1440
rect 20010 1405 20015 1435
rect 20045 1405 20050 1435
rect 20010 1400 20050 1405
rect 20120 1435 20160 1440
rect 20120 1405 20125 1435
rect 20155 1405 20160 1435
rect 20120 1400 20160 1405
rect 20526 1350 20558 1355
rect 19380 1335 19420 1340
rect 19380 1305 19385 1335
rect 19415 1305 19420 1335
rect 20526 1320 20528 1350
rect 20554 1320 20558 1350
rect 20526 1315 20558 1320
rect 20792 1350 20824 1355
rect 20792 1320 20796 1350
rect 20822 1320 20824 1350
rect 20792 1315 20824 1320
rect 19380 1300 19420 1305
rect 20095 1290 20135 1295
rect 11880 1250 11920 1255
rect 18815 1270 18855 1280
rect 18815 1250 18825 1270
rect 18845 1250 18855 1270
rect 12595 1240 12635 1245
rect 18815 1240 18855 1250
rect 18925 1275 18965 1280
rect 18925 1245 18930 1275
rect 18960 1245 18965 1275
rect 18925 1240 18965 1245
rect 19035 1275 19075 1280
rect 19035 1245 19040 1275
rect 19070 1245 19075 1275
rect 19035 1240 19075 1245
rect 19145 1275 19185 1280
rect 19145 1245 19150 1275
rect 19180 1245 19185 1275
rect 19145 1240 19185 1245
rect 19255 1275 19295 1280
rect 19255 1245 19260 1275
rect 19290 1245 19295 1275
rect 19255 1240 19295 1245
rect 19315 1270 19345 1280
rect 19315 1250 19320 1270
rect 19340 1250 19345 1270
rect 19315 1240 19345 1250
rect 19365 1275 19405 1280
rect 19365 1245 19370 1275
rect 19400 1245 19405 1275
rect 19365 1240 19405 1245
rect 19475 1275 19515 1280
rect 19475 1245 19480 1275
rect 19510 1245 19515 1275
rect 19475 1240 19515 1245
rect 19585 1275 19625 1280
rect 19585 1245 19590 1275
rect 19620 1245 19625 1275
rect 19585 1240 19625 1245
rect 19695 1275 19735 1280
rect 19695 1245 19700 1275
rect 19730 1245 19735 1275
rect 19695 1240 19735 1245
rect 19805 1275 19845 1280
rect 19805 1245 19810 1275
rect 19840 1245 19845 1275
rect 19805 1240 19845 1245
rect 19915 1275 19955 1280
rect 19915 1245 19920 1275
rect 19950 1245 19955 1275
rect 19915 1240 19955 1245
rect 20025 1275 20065 1280
rect 20025 1245 20030 1275
rect 20060 1245 20065 1275
rect 20095 1260 20100 1290
rect 20130 1260 20135 1290
rect 20095 1255 20135 1260
rect 20445 1290 20485 1295
rect 20445 1260 20450 1290
rect 20480 1260 20485 1290
rect 20445 1255 20485 1260
rect 20560 1290 20600 1295
rect 20560 1260 20565 1290
rect 20595 1260 20600 1290
rect 20560 1255 20600 1260
rect 20655 1290 20695 1295
rect 20655 1260 20660 1290
rect 20690 1260 20695 1290
rect 20655 1255 20695 1260
rect 20750 1290 20790 1295
rect 20750 1260 20755 1290
rect 20785 1260 20790 1290
rect 20750 1255 20790 1260
rect 20865 1290 20905 1295
rect 20865 1260 20870 1290
rect 20900 1260 20905 1290
rect 20865 1255 20905 1260
rect 20025 1240 20065 1245
rect 11315 1220 11355 1230
rect 11315 1200 11325 1220
rect 11345 1200 11355 1220
rect 11315 1190 11355 1200
rect 11425 1225 11465 1230
rect 11425 1195 11430 1225
rect 11460 1195 11465 1225
rect 11425 1190 11465 1195
rect 11535 1225 11575 1230
rect 11535 1195 11540 1225
rect 11570 1195 11575 1225
rect 11535 1190 11575 1195
rect 11645 1225 11685 1230
rect 11645 1195 11650 1225
rect 11680 1195 11685 1225
rect 11645 1190 11685 1195
rect 11755 1225 11795 1230
rect 11755 1195 11760 1225
rect 11790 1195 11795 1225
rect 11755 1190 11795 1195
rect 11815 1220 11845 1230
rect 11815 1200 11820 1220
rect 11840 1200 11845 1220
rect 11815 1190 11845 1200
rect 11865 1225 11905 1230
rect 11865 1195 11870 1225
rect 11900 1195 11905 1225
rect 11865 1190 11905 1195
rect 11975 1225 12015 1230
rect 11975 1195 11980 1225
rect 12010 1195 12015 1225
rect 11975 1190 12015 1195
rect 12085 1225 12125 1230
rect 12085 1195 12090 1225
rect 12120 1195 12125 1225
rect 12085 1190 12125 1195
rect 12195 1225 12235 1230
rect 12195 1195 12200 1225
rect 12230 1195 12235 1225
rect 12195 1190 12235 1195
rect 12305 1225 12345 1230
rect 12305 1195 12310 1225
rect 12340 1195 12345 1225
rect 12305 1190 12345 1195
rect 12415 1225 12455 1230
rect 12415 1195 12420 1225
rect 12450 1195 12455 1225
rect 12415 1190 12455 1195
rect 12525 1225 12565 1230
rect 12525 1195 12530 1225
rect 12560 1195 12565 1225
rect 12595 1210 12600 1240
rect 12630 1210 12635 1240
rect 20665 1235 20685 1255
rect 20875 1235 20895 1255
rect 12595 1205 12635 1210
rect 20600 1230 20640 1235
rect 20600 1200 20605 1230
rect 20635 1200 20640 1230
rect 20600 1195 20640 1200
rect 20660 1230 20690 1235
rect 20660 1195 20690 1200
rect 20710 1230 20750 1235
rect 20710 1200 20715 1230
rect 20745 1200 20750 1230
rect 20710 1195 20750 1200
rect 20865 1230 20905 1235
rect 20865 1200 20870 1230
rect 20900 1200 20905 1230
rect 20865 1195 20905 1200
rect 12525 1190 12565 1195
rect 3375 1185 3415 1190
rect 3375 1155 3380 1185
rect 3410 1155 3415 1185
rect 3375 1150 3415 1155
rect 3985 1185 4025 1190
rect 3985 1155 3990 1185
rect 4020 1155 4025 1185
rect 3985 1150 4025 1155
rect 4595 1185 4635 1190
rect 4595 1155 4600 1185
rect 4630 1155 4635 1185
rect 4595 1150 4635 1155
rect 2945 1125 2985 1130
rect 2945 1095 2950 1125
rect 2980 1095 2985 1125
rect 2945 1090 2985 1095
rect 3025 1125 3065 1130
rect 3025 1095 3030 1125
rect 3060 1095 3065 1125
rect 3025 1090 3065 1095
rect 3105 1125 3145 1130
rect 3105 1095 3110 1125
rect 3140 1095 3145 1125
rect 3105 1090 3145 1095
rect 3185 1125 3225 1130
rect 3185 1095 3190 1125
rect 3220 1095 3225 1125
rect 3185 1090 3225 1095
rect 3265 1125 3305 1130
rect 3265 1095 3270 1125
rect 3300 1095 3305 1125
rect 3265 1090 3305 1095
rect 3345 1125 3385 1130
rect 3345 1095 3350 1125
rect 3380 1095 3385 1125
rect 3345 1090 3385 1095
rect 3425 1125 3465 1130
rect 3425 1095 3430 1125
rect 3460 1095 3465 1125
rect 3425 1090 3465 1095
rect 3505 1125 3545 1130
rect 3505 1095 3510 1125
rect 3540 1095 3545 1125
rect 3505 1090 3545 1095
rect 3585 1125 3625 1130
rect 3585 1095 3590 1125
rect 3620 1095 3625 1125
rect 3585 1090 3625 1095
rect 3665 1125 3705 1130
rect 3665 1095 3670 1125
rect 3700 1095 3705 1125
rect 3665 1090 3705 1095
rect 3745 1125 3785 1130
rect 3745 1095 3750 1125
rect 3780 1095 3785 1125
rect 3745 1090 3785 1095
rect 3825 1125 3865 1130
rect 3825 1095 3830 1125
rect 3860 1095 3865 1125
rect 3825 1090 3865 1095
rect 3905 1125 3945 1130
rect 3905 1095 3910 1125
rect 3940 1095 3945 1125
rect 3905 1090 3945 1095
rect 3985 1125 4025 1130
rect 3985 1095 3990 1125
rect 4020 1095 4025 1125
rect 3985 1090 4025 1095
rect 4065 1125 4105 1130
rect 4065 1095 4070 1125
rect 4100 1095 4105 1125
rect 4065 1090 4105 1095
rect 4145 1125 4185 1130
rect 4145 1095 4150 1125
rect 4180 1095 4185 1125
rect 4145 1090 4185 1095
rect 4225 1125 4265 1130
rect 4225 1095 4230 1125
rect 4260 1095 4265 1125
rect 4225 1090 4265 1095
rect 4305 1125 4345 1130
rect 4305 1095 4310 1125
rect 4340 1095 4345 1125
rect 4305 1090 4345 1095
rect 4385 1125 4425 1130
rect 4385 1095 4390 1125
rect 4420 1095 4425 1125
rect 4385 1090 4425 1095
rect 4465 1125 4505 1130
rect 4465 1095 4470 1125
rect 4500 1095 4505 1125
rect 4465 1090 4505 1095
rect 4545 1125 4585 1130
rect 4545 1095 4550 1125
rect 4580 1095 4585 1125
rect 4545 1090 4585 1095
rect 4625 1125 4665 1130
rect 4625 1095 4630 1125
rect 4660 1095 4665 1125
rect 4625 1090 4665 1095
rect 4705 1125 4745 1130
rect 4705 1095 4710 1125
rect 4740 1095 4745 1125
rect 4705 1090 4745 1095
rect 4785 1125 4825 1130
rect 4785 1095 4790 1125
rect 4820 1095 4825 1125
rect 4785 1090 4825 1095
rect 4865 1125 4905 1130
rect 4865 1095 4870 1125
rect 4900 1095 4905 1125
rect 4865 1090 4905 1095
rect 4945 1125 4985 1130
rect 4945 1095 4950 1125
rect 4980 1095 4985 1125
rect 4945 1090 4985 1095
rect 2620 1040 2660 1045
rect 2620 1010 2625 1040
rect 2655 1010 2660 1040
rect 2620 1005 2660 1010
rect 2905 1040 2945 1045
rect 2905 1010 2910 1040
rect 2940 1010 2945 1040
rect 2905 1005 2945 1010
rect 5110 1040 5150 1045
rect 5110 1010 5115 1040
rect 5145 1010 5150 1040
rect 5110 1005 5150 1010
rect 13125 970 13165 975
rect 13125 940 13130 970
rect 13160 940 13165 970
rect 13125 935 13165 940
rect 13325 970 13365 975
rect 13325 940 13330 970
rect 13360 940 13365 970
rect 13325 935 13365 940
rect 13525 970 13565 975
rect 13525 940 13530 970
rect 13560 940 13565 970
rect 13525 935 13565 940
rect 13725 970 13765 975
rect 13725 940 13730 970
rect 13760 940 13765 970
rect 13725 935 13765 940
rect 13925 970 13965 975
rect 13925 940 13930 970
rect 13960 940 13965 970
rect 13925 935 13965 940
rect 18665 955 18705 960
rect 2995 930 3035 935
rect 2995 900 3000 930
rect 3030 900 3035 930
rect 2995 895 3035 900
rect 3175 930 3215 935
rect 3175 900 3180 930
rect 3210 900 3215 930
rect 3175 895 3215 900
rect 3355 930 3395 935
rect 3355 900 3360 930
rect 3390 900 3395 930
rect 3355 895 3395 900
rect 3535 930 3575 935
rect 3535 900 3540 930
rect 3570 900 3575 930
rect 3535 895 3575 900
rect 3715 930 3755 935
rect 3715 900 3720 930
rect 3750 900 3755 930
rect 3715 895 3755 900
rect 3895 930 3935 935
rect 3895 900 3900 930
rect 3930 900 3935 930
rect 3895 895 3935 900
rect 4075 930 4115 935
rect 4075 900 4080 930
rect 4110 900 4115 930
rect 4075 895 4115 900
rect 4255 930 4295 935
rect 4255 900 4260 930
rect 4290 900 4295 930
rect 4255 895 4295 900
rect 4435 930 4475 935
rect 4435 900 4440 930
rect 4470 900 4475 930
rect 4435 895 4475 900
rect 4615 930 4655 935
rect 4615 900 4620 930
rect 4650 900 4655 930
rect 4615 895 4655 900
rect 4795 930 4835 935
rect 4795 900 4800 930
rect 4830 900 4835 930
rect 4795 895 4835 900
rect 4975 930 5015 935
rect 4975 900 4980 930
rect 5010 900 5015 930
rect 18665 925 18670 955
rect 18700 925 18705 955
rect 18665 920 18705 925
rect 18760 955 18800 960
rect 18760 925 18765 955
rect 18795 925 18800 955
rect 18760 920 18800 925
rect 18870 955 18910 960
rect 18870 925 18875 955
rect 18905 925 18910 955
rect 18870 920 18910 925
rect 18980 955 19020 960
rect 18980 925 18985 955
rect 19015 925 19020 955
rect 18980 920 19020 925
rect 19090 955 19130 960
rect 19090 925 19095 955
rect 19125 925 19130 955
rect 19090 920 19130 925
rect 19200 955 19240 960
rect 19200 925 19205 955
rect 19235 925 19240 955
rect 19200 920 19240 925
rect 19310 955 19350 960
rect 19310 925 19315 955
rect 19345 925 19350 955
rect 19310 920 19350 925
rect 19420 955 19460 960
rect 19420 925 19425 955
rect 19455 925 19460 955
rect 19420 920 19460 925
rect 19530 955 19570 960
rect 19530 925 19535 955
rect 19565 925 19570 955
rect 19530 920 19570 925
rect 19640 955 19680 960
rect 19640 925 19645 955
rect 19675 925 19680 955
rect 19640 920 19680 925
rect 19750 955 19790 960
rect 19750 925 19755 955
rect 19785 925 19790 955
rect 19750 920 19790 925
rect 19860 955 19900 960
rect 19860 925 19865 955
rect 19895 925 19900 955
rect 19860 920 19900 925
rect 19970 955 20010 960
rect 19970 925 19975 955
rect 20005 925 20010 955
rect 19970 920 20010 925
rect 20120 955 20160 960
rect 20120 925 20125 955
rect 20155 925 20160 955
rect 20120 920 20160 925
rect 4975 895 5015 900
rect 11165 905 11205 910
rect 11165 875 11170 905
rect 11200 875 11205 905
rect 11165 870 11205 875
rect 11260 905 11300 910
rect 11260 875 11265 905
rect 11295 875 11300 905
rect 11260 870 11300 875
rect 11370 905 11410 910
rect 11370 875 11375 905
rect 11405 875 11410 905
rect 11370 870 11410 875
rect 11480 905 11520 910
rect 11480 875 11485 905
rect 11515 875 11520 905
rect 11480 870 11520 875
rect 11590 905 11630 910
rect 11590 875 11595 905
rect 11625 875 11630 905
rect 11590 870 11630 875
rect 11700 905 11740 910
rect 11700 875 11705 905
rect 11735 875 11740 905
rect 11700 870 11740 875
rect 11810 905 11850 910
rect 11810 875 11815 905
rect 11845 875 11850 905
rect 11810 870 11850 875
rect 11920 905 11960 910
rect 11920 875 11925 905
rect 11955 875 11960 905
rect 11920 870 11960 875
rect 12030 905 12070 910
rect 12030 875 12035 905
rect 12065 875 12070 905
rect 12030 870 12070 875
rect 12140 905 12180 910
rect 12140 875 12145 905
rect 12175 875 12180 905
rect 12140 870 12180 875
rect 12250 905 12290 910
rect 12250 875 12255 905
rect 12285 875 12290 905
rect 12250 870 12290 875
rect 12360 905 12400 910
rect 12360 875 12365 905
rect 12395 875 12400 905
rect 12360 870 12400 875
rect 12470 905 12510 910
rect 12470 875 12475 905
rect 12505 875 12510 905
rect 12470 870 12510 875
rect 12620 905 12660 910
rect 12620 875 12625 905
rect 12655 875 12660 905
rect 12620 870 12660 875
rect 2520 760 2560 765
rect 2520 730 2525 760
rect 2555 730 2560 760
rect 2520 725 2560 730
rect 3130 760 3170 765
rect 3130 730 3135 760
rect 3165 730 3170 760
rect 3130 725 3170 730
rect 3265 755 3305 765
rect 3265 735 3275 755
rect 3295 735 3305 755
rect 3265 725 3305 735
rect 3445 755 3485 765
rect 3445 735 3455 755
rect 3475 735 3485 755
rect 3445 725 3485 735
rect 3625 760 3665 765
rect 3625 730 3630 760
rect 3660 730 3665 760
rect 3625 725 3665 730
rect 3805 755 3845 765
rect 3805 735 3815 755
rect 3835 735 3845 755
rect 3805 725 3845 735
rect 3985 760 4025 765
rect 3985 730 3990 760
rect 4020 730 4025 760
rect 3985 725 4025 730
rect 4165 755 4205 765
rect 4165 735 4175 755
rect 4195 735 4205 755
rect 4165 725 4205 735
rect 4345 760 4385 765
rect 4345 730 4350 760
rect 4380 730 4385 760
rect 4345 725 4385 730
rect 4525 760 4565 765
rect 4525 730 4530 760
rect 4560 730 4565 760
rect 4525 725 4565 730
rect 4705 760 4745 765
rect 4705 730 4710 760
rect 4740 730 4745 760
rect 4705 725 4745 730
rect 4885 760 4925 765
rect 4885 730 4890 760
rect 4920 730 4925 760
rect 4885 725 4925 730
rect 3275 295 3295 725
rect 3455 710 3475 725
rect 3815 710 3835 725
rect 3445 705 3485 710
rect 3445 675 3450 705
rect 3480 675 3485 705
rect 3445 670 3485 675
rect 3805 705 3845 710
rect 3805 675 3810 705
rect 3840 675 3845 705
rect 3805 670 3845 675
rect 3815 295 3835 670
rect 3995 295 4015 725
rect 4175 710 4195 725
rect 4165 705 4205 710
rect 4165 675 4170 705
rect 4200 675 4205 705
rect 4165 670 4205 675
rect 4715 295 4735 725
rect 9375 -680 9415 -675
rect 9375 -710 9380 -680
rect 9410 -710 9415 -680
rect 9375 -715 9415 -710
rect 9575 -680 9615 -675
rect 9575 -710 9580 -680
rect 9610 -710 9615 -680
rect 9575 -715 9615 -710
rect 9775 -680 9815 -675
rect 9775 -710 9780 -680
rect 9810 -710 9815 -680
rect 9775 -715 9815 -710
rect 9975 -680 10015 -675
rect 9975 -710 9980 -680
rect 10010 -710 10015 -680
rect 9975 -715 10015 -710
rect 10175 -680 10215 -675
rect 10175 -710 10180 -680
rect 10210 -710 10215 -680
rect 10175 -715 10215 -710
rect 10375 -680 10415 -675
rect 10375 -710 10380 -680
rect 10410 -710 10415 -680
rect 10375 -715 10415 -710
rect 9475 -1030 9515 -1025
rect 9475 -1060 9480 -1030
rect 9510 -1060 9515 -1030
rect 9475 -1065 9515 -1060
rect 9675 -1030 9715 -1025
rect 9675 -1060 9680 -1030
rect 9710 -1060 9715 -1030
rect 9675 -1065 9715 -1060
rect 9875 -1030 9915 -1025
rect 9875 -1060 9880 -1030
rect 9910 -1060 9915 -1030
rect 9875 -1065 9915 -1060
rect 10075 -1030 10115 -1025
rect 10075 -1060 10080 -1030
rect 10110 -1060 10115 -1030
rect 10075 -1065 10115 -1060
rect 10275 -1030 10315 -1025
rect 10275 -1060 10280 -1030
rect 10310 -1060 10315 -1030
rect 10275 -1065 10315 -1060
<< via1 >>
rect 11345 3620 11375 3625
rect 11345 3600 11350 3620
rect 11350 3600 11370 3620
rect 11370 3600 11375 3620
rect 11345 3595 11375 3600
rect 11465 3620 11495 3625
rect 11465 3600 11470 3620
rect 11470 3600 11490 3620
rect 11490 3600 11495 3620
rect 11465 3595 11495 3600
rect 11585 3620 11615 3625
rect 11585 3600 11590 3620
rect 11590 3600 11610 3620
rect 11610 3600 11615 3620
rect 11585 3595 11615 3600
rect 11705 3620 11735 3625
rect 11705 3600 11710 3620
rect 11710 3600 11730 3620
rect 11730 3600 11735 3620
rect 11705 3595 11735 3600
rect 11825 3620 11855 3625
rect 11825 3600 11830 3620
rect 11830 3600 11850 3620
rect 11850 3600 11855 3620
rect 11825 3595 11855 3600
rect 11945 3620 11975 3625
rect 11945 3600 11950 3620
rect 11950 3600 11970 3620
rect 11970 3600 11975 3620
rect 11945 3595 11975 3600
rect 12065 3620 12095 3625
rect 12065 3600 12070 3620
rect 12070 3600 12090 3620
rect 12090 3600 12095 3620
rect 12065 3595 12095 3600
rect 12185 3620 12215 3625
rect 12185 3600 12190 3620
rect 12190 3600 12210 3620
rect 12210 3600 12215 3620
rect 12185 3595 12215 3600
rect 12305 3620 12335 3625
rect 12305 3600 12310 3620
rect 12310 3600 12330 3620
rect 12330 3600 12335 3620
rect 12305 3595 12335 3600
rect 12425 3620 12455 3625
rect 12425 3600 12430 3620
rect 12430 3600 12450 3620
rect 12450 3600 12455 3620
rect 12425 3595 12455 3600
rect 18845 3620 18875 3625
rect 18845 3600 18850 3620
rect 18850 3600 18870 3620
rect 18870 3600 18875 3620
rect 18845 3595 18875 3600
rect 18965 3620 18995 3625
rect 18965 3600 18970 3620
rect 18970 3600 18990 3620
rect 18990 3600 18995 3620
rect 18965 3595 18995 3600
rect 19085 3620 19115 3625
rect 19085 3600 19090 3620
rect 19090 3600 19110 3620
rect 19110 3600 19115 3620
rect 19085 3595 19115 3600
rect 19205 3620 19235 3625
rect 19205 3600 19210 3620
rect 19210 3600 19230 3620
rect 19230 3600 19235 3620
rect 19205 3595 19235 3600
rect 19325 3620 19355 3625
rect 19325 3600 19330 3620
rect 19330 3600 19350 3620
rect 19350 3600 19355 3620
rect 19325 3595 19355 3600
rect 19445 3620 19475 3625
rect 19445 3600 19450 3620
rect 19450 3600 19470 3620
rect 19470 3600 19475 3620
rect 19445 3595 19475 3600
rect 19565 3620 19595 3625
rect 19565 3600 19570 3620
rect 19570 3600 19590 3620
rect 19590 3600 19595 3620
rect 19565 3595 19595 3600
rect 19685 3620 19715 3625
rect 19685 3600 19690 3620
rect 19690 3600 19710 3620
rect 19710 3600 19715 3620
rect 19685 3595 19715 3600
rect 19805 3620 19835 3625
rect 19805 3600 19810 3620
rect 19810 3600 19830 3620
rect 19830 3600 19835 3620
rect 19805 3595 19835 3600
rect 19925 3620 19955 3625
rect 19925 3600 19930 3620
rect 19930 3600 19950 3620
rect 19950 3600 19955 3620
rect 19925 3595 19955 3600
rect 1266 3495 1296 3525
rect -10 3415 20 3445
rect 945 3415 975 3445
rect -55 3360 -25 3390
rect -55 2825 -25 2855
rect 1210 3310 1240 3340
rect 1165 3255 1195 3285
rect 51 3200 86 3205
rect 51 3175 56 3200
rect 56 3175 81 3200
rect 81 3175 86 3200
rect 51 3170 86 3175
rect 51 3140 86 3145
rect 51 3115 56 3140
rect 56 3115 81 3140
rect 81 3115 86 3140
rect 51 3110 86 3115
rect 1165 3070 1195 3100
rect 51 3060 86 3065
rect 51 3035 56 3060
rect 56 3035 81 3060
rect 81 3035 86 3060
rect 51 3030 86 3035
rect 51 3000 86 3005
rect 51 2975 56 3000
rect 56 2975 81 3000
rect 81 2975 86 3000
rect 51 2970 86 2975
rect 920 2880 950 2910
rect 1000 2880 1030 2910
rect 1080 2880 1110 2910
rect 4445 3465 4475 3495
rect 1645 3415 1675 3445
rect 2475 3420 2505 3450
rect 1266 3195 1301 3200
rect 1266 3170 1271 3195
rect 1271 3170 1296 3195
rect 1296 3170 1301 3195
rect 1266 3165 1301 3170
rect 1266 3135 1301 3140
rect 1266 3110 1271 3135
rect 1271 3110 1296 3135
rect 1296 3110 1301 3135
rect 1266 3105 1301 3110
rect 2335 2955 2370 2960
rect 2335 2930 2340 2955
rect 2340 2930 2365 2955
rect 2365 2930 2370 2955
rect 2335 2925 2370 2930
rect 2430 2925 2460 2955
rect 2335 2895 2370 2900
rect 2335 2870 2340 2895
rect 2340 2870 2365 2895
rect 2365 2870 2370 2895
rect 2335 2865 2370 2870
rect 56 2850 91 2855
rect 56 2825 61 2850
rect 61 2825 86 2850
rect 86 2825 91 2850
rect 56 2820 91 2825
rect 729 2850 764 2855
rect 729 2825 734 2850
rect 734 2825 759 2850
rect 759 2825 764 2850
rect 729 2820 764 2825
rect 1210 2820 1240 2850
rect 1266 2835 1301 2840
rect 1266 2810 1271 2835
rect 1271 2810 1296 2835
rect 1296 2810 1301 2835
rect 1266 2805 1301 2810
rect 1965 2835 2000 2840
rect 1965 2810 1970 2835
rect 1970 2810 1995 2835
rect 1995 2810 2000 2835
rect 1965 2805 2000 2810
rect 2335 2805 2365 2835
rect -10 2765 20 2795
rect 56 2790 91 2795
rect 56 2765 61 2790
rect 61 2765 86 2790
rect 86 2765 91 2790
rect 56 2760 91 2765
rect 729 2790 764 2795
rect 729 2765 734 2790
rect 734 2765 759 2790
rect 759 2765 764 2790
rect 729 2760 764 2765
rect 1266 2715 1296 2745
rect 2155 2715 2185 2745
rect -105 1690 -75 1720
rect -40 1715 -10 1720
rect -40 1695 -35 1715
rect -35 1695 -15 1715
rect -15 1695 -10 1715
rect -40 1690 -10 1695
rect 1270 1680 1297 1710
rect 2430 2215 2460 2245
rect 2335 2170 2365 2200
rect 2385 2120 2415 2150
rect 2695 3360 2725 3390
rect 3140 3310 3170 3340
rect 3395 3305 3425 3335
rect 2740 3210 2770 3240
rect 2625 3155 2655 3185
rect 2525 2950 2555 2980
rect 2475 1790 2505 1820
rect 2430 1730 2460 1760
rect 2385 1635 2415 1665
rect 2335 1565 2365 1595
rect 2625 2760 2655 2790
rect 2625 2315 2655 2345
rect 5145 3415 5175 3445
rect 5365 3305 5395 3335
rect 4890 3255 4920 3285
rect 4445 3155 4475 3185
rect 3140 3110 3170 3140
rect 4840 3110 4870 3140
rect 3990 3050 4020 3080
rect 3450 3005 3480 3035
rect 3810 3005 3840 3035
rect 4350 3005 4380 3035
rect 4710 3005 4740 3035
rect 5320 3110 5350 3140
rect 3085 2975 3115 2980
rect 3085 2955 3090 2975
rect 3090 2955 3110 2975
rect 3110 2955 3115 2975
rect 3085 2950 3115 2955
rect 3270 2975 3300 2980
rect 3270 2955 3275 2975
rect 3275 2955 3295 2975
rect 3295 2955 3300 2975
rect 3270 2950 3300 2955
rect 3630 2975 3660 2980
rect 3630 2955 3635 2975
rect 3635 2955 3655 2975
rect 3655 2955 3660 2975
rect 3630 2950 3660 2955
rect 4170 2975 4200 2980
rect 4170 2955 4175 2975
rect 4175 2955 4195 2975
rect 4195 2955 4200 2975
rect 4170 2950 4200 2955
rect 4530 2975 4560 2980
rect 4530 2955 4535 2975
rect 4535 2955 4555 2975
rect 4555 2955 4560 2975
rect 4530 2950 4560 2955
rect 3000 2805 3030 2810
rect 3000 2785 3005 2805
rect 3005 2785 3025 2805
rect 3025 2785 3030 2805
rect 3000 2780 3030 2785
rect 3180 2805 3210 2810
rect 3180 2785 3185 2805
rect 3185 2785 3205 2805
rect 3205 2785 3210 2805
rect 3180 2780 3210 2785
rect 3360 2805 3390 2810
rect 3360 2785 3365 2805
rect 3365 2785 3385 2805
rect 3385 2785 3390 2805
rect 3360 2780 3390 2785
rect 3540 2805 3570 2810
rect 3540 2785 3545 2805
rect 3545 2785 3565 2805
rect 3565 2785 3570 2805
rect 3540 2780 3570 2785
rect 3720 2805 3750 2810
rect 3720 2785 3725 2805
rect 3725 2785 3745 2805
rect 3745 2785 3750 2805
rect 3720 2780 3750 2785
rect 3900 2805 3930 2810
rect 3900 2785 3905 2805
rect 3905 2785 3925 2805
rect 3925 2785 3930 2805
rect 3900 2780 3930 2785
rect 4080 2805 4110 2810
rect 4080 2785 4085 2805
rect 4085 2785 4105 2805
rect 4105 2785 4110 2805
rect 4080 2780 4110 2785
rect 4260 2805 4290 2810
rect 4260 2785 4265 2805
rect 4265 2785 4285 2805
rect 4285 2785 4290 2805
rect 4260 2780 4290 2785
rect 4440 2805 4470 2810
rect 4440 2785 4445 2805
rect 4445 2785 4465 2805
rect 4465 2785 4470 2805
rect 4440 2780 4470 2785
rect 4620 2805 4650 2810
rect 4620 2785 4625 2805
rect 4625 2785 4645 2805
rect 4645 2785 4650 2805
rect 4620 2780 4650 2785
rect 4800 2805 4830 2810
rect 4800 2785 4805 2805
rect 4805 2785 4825 2805
rect 4825 2785 4830 2805
rect 4800 2780 4830 2785
rect 4980 2805 5010 2810
rect 4980 2785 4985 2805
rect 4985 2785 5005 2805
rect 5005 2785 5010 2805
rect 4980 2780 5010 2785
rect 3180 2745 3210 2750
rect 3180 2725 3185 2745
rect 3185 2725 3205 2745
rect 3205 2725 3210 2745
rect 3180 2720 3210 2725
rect 3360 2745 3390 2750
rect 3360 2725 3365 2745
rect 3365 2725 3385 2745
rect 3385 2725 3390 2745
rect 3360 2720 3390 2725
rect 3540 2745 3570 2750
rect 3540 2725 3545 2745
rect 3545 2725 3565 2745
rect 3565 2725 3570 2745
rect 3540 2720 3570 2725
rect 3720 2745 3750 2750
rect 3720 2725 3725 2745
rect 3725 2725 3745 2745
rect 3745 2725 3750 2745
rect 3720 2720 3750 2725
rect 3900 2745 3930 2750
rect 3900 2725 3905 2745
rect 3905 2725 3925 2745
rect 3925 2725 3930 2745
rect 3900 2720 3930 2725
rect 4080 2745 4110 2750
rect 4080 2725 4085 2745
rect 4085 2725 4105 2745
rect 4105 2725 4110 2745
rect 4080 2720 4110 2725
rect 4260 2745 4290 2750
rect 4260 2725 4265 2745
rect 4265 2725 4285 2745
rect 4285 2725 4290 2745
rect 4260 2720 4290 2725
rect 4440 2745 4470 2750
rect 4440 2725 4445 2745
rect 4445 2725 4465 2745
rect 4465 2725 4470 2745
rect 4440 2720 4470 2725
rect 4620 2745 4650 2750
rect 4620 2725 4625 2745
rect 4625 2725 4645 2745
rect 4645 2725 4650 2745
rect 4620 2720 4650 2725
rect 4800 2745 4830 2750
rect 4800 2725 4805 2745
rect 4805 2725 4825 2745
rect 4825 2725 4830 2745
rect 4800 2720 4830 2725
rect 3360 2370 3390 2375
rect 3360 2350 3365 2370
rect 3365 2350 3385 2370
rect 3385 2350 3390 2370
rect 3360 2345 3390 2350
rect 3810 2375 3840 2380
rect 3810 2355 3815 2375
rect 3815 2355 3835 2375
rect 3835 2355 3840 2375
rect 3810 2350 3840 2355
rect 4170 2375 4200 2380
rect 4170 2355 4175 2375
rect 4175 2355 4195 2375
rect 4195 2355 4200 2375
rect 4170 2350 4200 2355
rect 2740 2260 2770 2290
rect 3630 2330 3660 2335
rect 3630 2310 3635 2330
rect 3635 2310 3655 2330
rect 3655 2310 3660 2330
rect 3630 2305 3660 2310
rect 3450 2285 3480 2290
rect 3450 2265 3455 2285
rect 3455 2265 3475 2285
rect 3475 2265 3480 2285
rect 3450 2260 3480 2265
rect 3270 2170 3300 2200
rect 3810 2215 3840 2245
rect 3630 2120 3660 2150
rect 2750 2090 2780 2095
rect 2750 2070 2755 2090
rect 2755 2070 2775 2090
rect 2775 2070 2780 2090
rect 2750 2065 2780 2070
rect 2870 2090 2900 2095
rect 2870 2070 2875 2090
rect 2875 2070 2895 2090
rect 2895 2070 2900 2090
rect 2870 2065 2900 2070
rect 2990 2090 3020 2095
rect 2990 2070 2995 2090
rect 2995 2070 3015 2090
rect 3015 2070 3020 2090
rect 2990 2065 3020 2070
rect 3110 2090 3140 2095
rect 3110 2070 3115 2090
rect 3115 2070 3135 2090
rect 3135 2070 3140 2090
rect 3110 2065 3140 2070
rect 3230 2090 3260 2095
rect 3230 2070 3235 2090
rect 3235 2070 3255 2090
rect 3255 2070 3260 2090
rect 3230 2065 3260 2070
rect 3350 2090 3380 2095
rect 3350 2070 3355 2090
rect 3355 2070 3375 2090
rect 3375 2070 3380 2090
rect 3350 2065 3380 2070
rect 3470 2090 3500 2095
rect 3470 2070 3475 2090
rect 3475 2070 3495 2090
rect 3495 2070 3500 2090
rect 3470 2065 3500 2070
rect 3590 2090 3620 2095
rect 3590 2070 3595 2090
rect 3595 2070 3615 2090
rect 3615 2070 3620 2090
rect 3590 2065 3620 2070
rect 3710 2090 3740 2095
rect 3710 2070 3715 2090
rect 3715 2070 3735 2090
rect 3735 2070 3740 2090
rect 3710 2065 3740 2070
rect 3830 2090 3860 2095
rect 3830 2070 3835 2090
rect 3835 2070 3855 2090
rect 3855 2070 3860 2090
rect 3830 2065 3860 2070
rect 4350 2330 4380 2335
rect 4350 2310 4355 2330
rect 4355 2310 4375 2330
rect 4375 2310 4380 2330
rect 4350 2305 4380 2310
rect 4530 2285 4560 2290
rect 4530 2265 4535 2285
rect 4535 2265 4555 2285
rect 4555 2265 4560 2285
rect 4530 2260 4560 2265
rect 5275 2260 5305 2290
rect 3990 2170 4020 2200
rect 4710 2170 4740 2200
rect 4090 2115 4120 2145
rect 3990 2090 4020 2095
rect 3990 2070 3995 2090
rect 3995 2070 4015 2090
rect 4015 2070 4020 2090
rect 3990 2065 4020 2070
rect 4150 2090 4180 2095
rect 4150 2070 4155 2090
rect 4155 2070 4175 2090
rect 4175 2070 4180 2090
rect 4150 2065 4180 2070
rect 4270 2090 4300 2095
rect 4270 2070 4275 2090
rect 4275 2070 4295 2090
rect 4295 2070 4300 2090
rect 4270 2065 4300 2070
rect 4390 2090 4420 2095
rect 4390 2070 4395 2090
rect 4395 2070 4415 2090
rect 4415 2070 4420 2090
rect 4390 2065 4420 2070
rect 4510 2090 4540 2095
rect 4510 2070 4515 2090
rect 4515 2070 4535 2090
rect 4535 2070 4540 2090
rect 4510 2065 4540 2070
rect 4630 2090 4660 2095
rect 4630 2070 4635 2090
rect 4635 2070 4655 2090
rect 4655 2070 4660 2090
rect 4630 2065 4660 2070
rect 4750 2090 4780 2095
rect 4750 2070 4755 2090
rect 4755 2070 4775 2090
rect 4775 2070 4780 2090
rect 4750 2065 4780 2070
rect 4870 2090 4900 2095
rect 4870 2070 4875 2090
rect 4875 2070 4895 2090
rect 4895 2070 4900 2090
rect 4870 2065 4900 2070
rect 4990 2090 5020 2095
rect 4990 2070 4995 2090
rect 4995 2070 5015 2090
rect 5015 2070 5020 2090
rect 4990 2065 5020 2070
rect 5110 2090 5140 2095
rect 5110 2070 5115 2090
rect 5115 2070 5135 2090
rect 5135 2070 5140 2090
rect 5110 2065 5140 2070
rect 5230 2090 5260 2095
rect 5230 2070 5235 2090
rect 5235 2070 5255 2090
rect 5255 2070 5260 2090
rect 5230 2065 5260 2070
rect 2625 2045 2655 2050
rect 2625 2025 2630 2045
rect 2630 2025 2650 2045
rect 2650 2025 2655 2045
rect 2625 2020 2655 2025
rect 2810 2045 2840 2050
rect 2810 2025 2815 2045
rect 2815 2025 2835 2045
rect 2835 2025 2840 2045
rect 2810 2020 2840 2025
rect 3170 2045 3200 2050
rect 3170 2025 3175 2045
rect 3175 2025 3195 2045
rect 3195 2025 3200 2045
rect 3170 2020 3200 2025
rect 3530 2045 3560 2050
rect 3530 2025 3535 2045
rect 3535 2025 3555 2045
rect 3555 2025 3560 2045
rect 3530 2020 3560 2025
rect 3890 2045 3920 2050
rect 4090 2045 4120 2050
rect 3890 2025 3895 2045
rect 3895 2025 3915 2045
rect 3915 2025 3920 2045
rect 3890 2020 3920 2025
rect 2930 1875 2960 1880
rect 2930 1855 2935 1875
rect 2935 1855 2955 1875
rect 2955 1855 2960 1875
rect 2930 1850 2960 1855
rect 3290 1875 3320 1880
rect 3290 1855 3295 1875
rect 3295 1855 3315 1875
rect 3315 1855 3320 1875
rect 3290 1850 3320 1855
rect 3650 1875 3680 1880
rect 3650 1855 3655 1875
rect 3655 1855 3675 1875
rect 3675 1855 3680 1875
rect 3650 1850 3680 1855
rect 2570 1730 2600 1760
rect 2840 1790 2870 1820
rect 3050 1815 3080 1820
rect 3050 1795 3055 1815
rect 3055 1795 3075 1815
rect 3075 1795 3080 1815
rect 3050 1790 3080 1795
rect 3170 1790 3200 1820
rect 3410 1815 3440 1820
rect 3410 1795 3415 1815
rect 3415 1795 3435 1815
rect 3435 1795 3440 1815
rect 3410 1790 3440 1795
rect 3530 1790 3560 1820
rect 3770 1815 3800 1820
rect 3770 1795 3775 1815
rect 3775 1795 3795 1815
rect 3795 1795 3800 1815
rect 3770 1790 3800 1795
rect 3860 1790 3890 1820
rect 2680 1730 2710 1760
rect 2805 1735 2835 1765
rect 3230 1755 3260 1760
rect 3230 1735 3235 1755
rect 3235 1735 3255 1755
rect 3255 1735 3260 1755
rect 3230 1730 3260 1735
rect 3290 1755 3320 1760
rect 3290 1735 3295 1755
rect 3295 1735 3315 1755
rect 3315 1735 3320 1755
rect 3290 1730 3320 1735
rect 3530 1755 3560 1760
rect 3530 1735 3535 1755
rect 3535 1735 3555 1755
rect 3555 1735 3560 1755
rect 3530 1730 3560 1735
rect 3770 1755 3800 1760
rect 3770 1735 3775 1755
rect 3775 1735 3795 1755
rect 3795 1735 3800 1755
rect 3770 1730 3800 1735
rect 2805 1680 2835 1710
rect 3170 1710 3200 1715
rect 3170 1690 3175 1710
rect 3175 1690 3195 1710
rect 3195 1690 3200 1710
rect 3170 1685 3200 1690
rect 3410 1710 3440 1715
rect 3410 1690 3415 1710
rect 3415 1690 3435 1710
rect 3435 1690 3440 1710
rect 3410 1685 3440 1690
rect 3650 1710 3680 1715
rect 3650 1690 3655 1710
rect 3655 1690 3675 1710
rect 3675 1690 3680 1710
rect 3650 1685 3680 1690
rect 2625 1635 2655 1665
rect 3170 1590 3200 1595
rect 3170 1570 3175 1590
rect 3175 1570 3195 1590
rect 3195 1570 3200 1590
rect 3170 1565 3200 1570
rect 2840 1515 2870 1545
rect 3230 1540 3260 1545
rect 3230 1520 3235 1540
rect 3235 1520 3255 1540
rect 3255 1520 3260 1540
rect 3230 1515 3260 1520
rect 3350 1540 3380 1545
rect 3350 1520 3355 1540
rect 3355 1520 3375 1540
rect 3375 1520 3380 1540
rect 3350 1515 3380 1520
rect 3470 1540 3500 1545
rect 3470 1520 3475 1540
rect 3475 1520 3495 1540
rect 3495 1520 3500 1540
rect 3470 1515 3500 1520
rect 3590 1540 3620 1545
rect 3590 1520 3595 1540
rect 3595 1520 3615 1540
rect 3615 1520 3620 1540
rect 3590 1515 3620 1520
rect 3710 1540 3740 1545
rect 3710 1520 3715 1540
rect 3715 1520 3735 1540
rect 3735 1520 3740 1540
rect 3710 1515 3740 1520
rect 2930 1495 2960 1500
rect 2930 1475 2935 1495
rect 2935 1475 2955 1495
rect 2955 1475 2960 1495
rect 2930 1470 2960 1475
rect 3050 1495 3080 1500
rect 3050 1475 3055 1495
rect 3055 1475 3075 1495
rect 3075 1475 3080 1495
rect 3050 1470 3080 1475
rect 3170 1495 3200 1500
rect 3170 1475 3175 1495
rect 3175 1475 3195 1495
rect 3195 1475 3200 1495
rect 3170 1470 3200 1475
rect 3290 1495 3320 1500
rect 3290 1475 3295 1495
rect 3295 1475 3315 1495
rect 3315 1475 3320 1495
rect 3290 1470 3320 1475
rect 3530 1495 3560 1500
rect 3530 1475 3535 1495
rect 3535 1475 3555 1495
rect 3555 1475 3560 1495
rect 3530 1470 3560 1475
rect 3650 1495 3680 1500
rect 3650 1475 3655 1495
rect 3655 1475 3675 1495
rect 3675 1475 3680 1495
rect 3650 1470 3680 1475
rect 3770 1495 3800 1500
rect 3770 1475 3775 1495
rect 3775 1475 3795 1495
rect 3795 1475 3800 1495
rect 3770 1470 3800 1475
rect 4090 2025 4095 2045
rect 4095 2025 4115 2045
rect 4115 2025 4120 2045
rect 4090 2020 4120 2025
rect 4450 2045 4480 2050
rect 4450 2025 4455 2045
rect 4455 2025 4475 2045
rect 4475 2025 4480 2045
rect 4450 2020 4480 2025
rect 4810 2045 4840 2050
rect 4810 2025 4815 2045
rect 4815 2025 4835 2045
rect 4835 2025 4840 2045
rect 4810 2020 4840 2025
rect 5170 2045 5200 2050
rect 5170 2025 5175 2045
rect 5175 2025 5195 2045
rect 5195 2025 5200 2045
rect 5170 2020 5200 2025
rect 4330 1875 4360 1880
rect 4330 1855 4335 1875
rect 4335 1855 4355 1875
rect 4355 1855 4360 1875
rect 4330 1850 4360 1855
rect 4690 1875 4720 1880
rect 4690 1855 4695 1875
rect 4695 1855 4715 1875
rect 4715 1855 4720 1875
rect 4690 1850 4720 1855
rect 5050 1875 5080 1880
rect 5050 1855 5055 1875
rect 5055 1855 5075 1875
rect 5075 1855 5080 1875
rect 5050 1850 5080 1855
rect 4120 1790 4150 1820
rect 4210 1815 4240 1820
rect 4210 1795 4215 1815
rect 4215 1795 4235 1815
rect 4235 1795 4240 1815
rect 4210 1790 4240 1795
rect 4450 1790 4480 1820
rect 4570 1815 4600 1820
rect 4570 1795 4575 1815
rect 4575 1795 4595 1815
rect 4595 1795 4600 1815
rect 4570 1790 4600 1795
rect 4210 1755 4240 1760
rect 4210 1735 4215 1755
rect 4215 1735 4235 1755
rect 4235 1735 4240 1755
rect 4210 1730 4240 1735
rect 4450 1755 4480 1760
rect 4450 1735 4455 1755
rect 4455 1735 4475 1755
rect 4475 1735 4480 1755
rect 4450 1730 4480 1735
rect 4810 1790 4840 1820
rect 4930 1815 4960 1820
rect 4930 1795 4935 1815
rect 4935 1795 4955 1815
rect 4955 1795 4960 1815
rect 4930 1790 4960 1795
rect 5140 1790 5170 1820
rect 5320 2115 5350 2145
rect 5415 3255 5445 3285
rect 12950 3285 12980 3290
rect 12950 3265 12955 3285
rect 12955 3265 12975 3285
rect 12975 3265 12980 3285
rect 12950 3260 12980 3265
rect 13060 3285 13090 3290
rect 13060 3265 13065 3285
rect 13065 3265 13085 3285
rect 13085 3265 13090 3285
rect 13060 3260 13090 3265
rect 13170 3285 13200 3290
rect 13170 3265 13175 3285
rect 13175 3265 13195 3285
rect 13195 3265 13200 3285
rect 13170 3260 13200 3265
rect 13280 3285 13310 3290
rect 13280 3265 13285 3285
rect 13285 3265 13305 3285
rect 13305 3265 13310 3285
rect 13280 3260 13310 3265
rect 13390 3285 13420 3290
rect 13390 3265 13395 3285
rect 13395 3265 13415 3285
rect 13415 3265 13420 3285
rect 13390 3260 13420 3265
rect 13500 3285 13530 3290
rect 13500 3265 13505 3285
rect 13505 3265 13525 3285
rect 13525 3265 13530 3285
rect 13500 3260 13530 3265
rect 13610 3285 13640 3290
rect 13610 3265 13615 3285
rect 13615 3265 13635 3285
rect 13635 3265 13640 3285
rect 13610 3260 13640 3265
rect 13720 3285 13750 3290
rect 13720 3265 13725 3285
rect 13725 3265 13745 3285
rect 13745 3265 13750 3285
rect 13720 3260 13750 3265
rect 13830 3285 13860 3290
rect 13830 3265 13835 3285
rect 13835 3265 13855 3285
rect 13855 3265 13860 3285
rect 13830 3260 13860 3265
rect 13940 3285 13970 3290
rect 13940 3265 13945 3285
rect 13945 3265 13965 3285
rect 13965 3265 13970 3285
rect 13940 3260 13970 3265
rect 14050 3285 14080 3290
rect 14050 3265 14055 3285
rect 14055 3265 14075 3285
rect 14075 3265 14080 3285
rect 14050 3260 14080 3265
rect 20450 3285 20480 3290
rect 20450 3265 20455 3285
rect 20455 3265 20475 3285
rect 20475 3265 20480 3285
rect 20450 3260 20480 3265
rect 20560 3285 20590 3290
rect 20560 3265 20565 3285
rect 20565 3265 20585 3285
rect 20585 3265 20590 3285
rect 20560 3260 20590 3265
rect 20670 3285 20700 3290
rect 20670 3265 20675 3285
rect 20675 3265 20695 3285
rect 20695 3265 20700 3285
rect 20670 3260 20700 3265
rect 20780 3285 20810 3290
rect 20780 3265 20785 3285
rect 20785 3265 20805 3285
rect 20805 3265 20810 3285
rect 20780 3260 20810 3265
rect 20890 3285 20920 3290
rect 20890 3265 20895 3285
rect 20895 3265 20915 3285
rect 20915 3265 20920 3285
rect 20890 3260 20920 3265
rect 21000 3285 21030 3290
rect 21000 3265 21005 3285
rect 21005 3265 21025 3285
rect 21025 3265 21030 3285
rect 21000 3260 21030 3265
rect 21110 3285 21140 3290
rect 21110 3265 21115 3285
rect 21115 3265 21135 3285
rect 21135 3265 21140 3285
rect 21110 3260 21140 3265
rect 21220 3285 21250 3290
rect 21220 3265 21225 3285
rect 21225 3265 21245 3285
rect 21245 3265 21250 3285
rect 21220 3260 21250 3265
rect 21330 3285 21360 3290
rect 21330 3265 21335 3285
rect 21335 3265 21355 3285
rect 21355 3265 21360 3285
rect 21330 3260 21360 3265
rect 21440 3285 21470 3290
rect 21440 3265 21445 3285
rect 21445 3265 21465 3285
rect 21465 3265 21470 3285
rect 21440 3260 21470 3265
rect 21550 3285 21580 3290
rect 21550 3265 21555 3285
rect 21555 3265 21575 3285
rect 21575 3265 21580 3285
rect 21550 3260 21580 3265
rect 5365 1790 5395 1820
rect 4690 1755 4720 1760
rect 4690 1735 4695 1755
rect 4695 1735 4715 1755
rect 4715 1735 4720 1755
rect 4690 1730 4720 1735
rect 4750 1755 4780 1760
rect 4750 1735 4755 1755
rect 4755 1735 4775 1755
rect 4775 1735 4780 1755
rect 4750 1730 4780 1735
rect 5275 1730 5305 1760
rect 4330 1710 4360 1715
rect 4330 1690 4335 1710
rect 4335 1690 4355 1710
rect 4355 1690 4360 1710
rect 4330 1685 4360 1690
rect 4570 1710 4600 1715
rect 4570 1690 4575 1710
rect 4575 1690 4595 1710
rect 4595 1690 4600 1710
rect 4570 1685 4600 1690
rect 4810 1710 4840 1715
rect 4810 1690 4815 1710
rect 4815 1690 4835 1710
rect 4835 1690 4840 1710
rect 4810 1685 4840 1690
rect 10585 3205 10615 3210
rect 10585 3185 10590 3205
rect 10590 3185 10610 3205
rect 10610 3185 10615 3205
rect 10585 3180 10615 3185
rect 10985 3205 11015 3210
rect 10985 3185 10990 3205
rect 10990 3185 11010 3205
rect 11010 3185 11015 3205
rect 10985 3180 11015 3185
rect 18085 3205 18115 3210
rect 18085 3185 18090 3205
rect 18090 3185 18110 3205
rect 18110 3185 18115 3205
rect 18085 3180 18115 3185
rect 18485 3205 18515 3210
rect 18485 3185 18490 3205
rect 18490 3185 18510 3205
rect 18510 3185 18515 3205
rect 18485 3180 18515 3185
rect 10905 3125 10935 3155
rect 9740 2665 9770 2670
rect 9740 2645 9745 2665
rect 9745 2645 9765 2665
rect 9765 2645 9770 2665
rect 9740 2640 9770 2645
rect 9850 2665 9880 2670
rect 9850 2645 9855 2665
rect 9855 2645 9875 2665
rect 9875 2645 9880 2665
rect 9850 2640 9880 2645
rect 9960 2665 9990 2670
rect 9960 2645 9965 2665
rect 9965 2645 9985 2665
rect 9985 2645 9990 2665
rect 9960 2640 9990 2645
rect 10070 2665 10100 2670
rect 10070 2645 10075 2665
rect 10075 2645 10095 2665
rect 10095 2645 10100 2665
rect 10070 2640 10100 2645
rect 10180 2665 10210 2670
rect 10180 2645 10185 2665
rect 10185 2645 10205 2665
rect 10205 2645 10210 2665
rect 10180 2640 10210 2645
rect 10290 2665 10320 2670
rect 10290 2645 10295 2665
rect 10295 2645 10315 2665
rect 10315 2645 10320 2665
rect 10290 2640 10320 2645
rect 10400 2665 10430 2670
rect 10400 2645 10405 2665
rect 10405 2645 10425 2665
rect 10425 2645 10430 2665
rect 10400 2640 10430 2645
rect 10510 2665 10540 2670
rect 10510 2645 10515 2665
rect 10515 2645 10535 2665
rect 10535 2645 10540 2665
rect 10510 2640 10540 2645
rect 10620 2665 10650 2670
rect 10620 2645 10625 2665
rect 10625 2645 10645 2665
rect 10645 2645 10650 2665
rect 10620 2640 10650 2645
rect 10730 2665 10760 2670
rect 10730 2645 10735 2665
rect 10735 2645 10755 2665
rect 10755 2645 10760 2665
rect 10730 2640 10760 2645
rect 10840 2665 10870 2670
rect 10840 2645 10845 2665
rect 10845 2645 10865 2665
rect 10865 2645 10870 2665
rect 10840 2640 10870 2645
rect 9795 2495 9825 2500
rect 9795 2475 9800 2495
rect 9800 2475 9820 2495
rect 9820 2475 9825 2495
rect 9795 2470 9825 2475
rect 9905 2495 9935 2500
rect 9905 2475 9910 2495
rect 9910 2475 9930 2495
rect 9930 2475 9935 2495
rect 9905 2470 9935 2475
rect 10015 2495 10045 2500
rect 10015 2475 10020 2495
rect 10020 2475 10040 2495
rect 10040 2475 10045 2495
rect 10015 2470 10045 2475
rect 10125 2495 10155 2500
rect 10125 2475 10130 2495
rect 10130 2475 10150 2495
rect 10150 2475 10155 2495
rect 10125 2470 10155 2475
rect 10235 2495 10265 2500
rect 10235 2475 10240 2495
rect 10240 2475 10260 2495
rect 10260 2475 10265 2495
rect 10235 2470 10265 2475
rect 10345 2495 10375 2500
rect 10345 2475 10350 2495
rect 10350 2475 10370 2495
rect 10370 2475 10375 2495
rect 10345 2470 10375 2475
rect 10455 2495 10485 2500
rect 10455 2475 10460 2495
rect 10460 2475 10480 2495
rect 10480 2475 10485 2495
rect 10455 2470 10485 2475
rect 10565 2495 10595 2500
rect 10565 2475 10570 2495
rect 10570 2475 10590 2495
rect 10590 2475 10595 2495
rect 10565 2470 10595 2475
rect 10675 2495 10705 2500
rect 10675 2475 10680 2495
rect 10680 2475 10700 2495
rect 10700 2475 10705 2495
rect 10675 2470 10705 2475
rect 10785 2495 10815 2500
rect 10785 2475 10790 2495
rect 10790 2475 10810 2495
rect 10810 2475 10815 2495
rect 10785 2470 10815 2475
rect 11826 3150 11854 3155
rect 11826 3130 11831 3150
rect 11831 3130 11849 3150
rect 11849 3130 11854 3150
rect 11826 3125 11854 3130
rect 18405 3125 18435 3155
rect 11285 3070 11315 3100
rect 11525 3070 11555 3100
rect 11765 3070 11795 3100
rect 12005 3070 12035 3100
rect 12245 3070 12275 3100
rect 12485 3070 12515 3100
rect 11405 3025 11435 3055
rect 11645 3025 11675 3055
rect 11885 3025 11915 3055
rect 12125 3025 12155 3055
rect 12365 3025 12395 3055
rect 11345 2970 11375 3000
rect 11405 2970 11435 3000
rect 11585 2970 11615 3000
rect 11825 2970 11855 3000
rect 12065 2970 12095 3000
rect 12305 2970 12335 3000
rect 11465 2940 11495 2945
rect 11465 2920 11470 2940
rect 11470 2920 11490 2940
rect 11490 2920 11495 2940
rect 11465 2915 11495 2920
rect 11705 2940 11735 2945
rect 11705 2920 11710 2940
rect 11710 2920 11730 2940
rect 11730 2920 11735 2940
rect 11705 2915 11735 2920
rect 11945 2940 11975 2945
rect 11945 2920 11950 2940
rect 11950 2920 11970 2940
rect 11970 2920 11975 2940
rect 11945 2915 11975 2920
rect 12185 2940 12215 2945
rect 12185 2920 12190 2940
rect 12190 2920 12210 2940
rect 12210 2920 12215 2940
rect 12185 2915 12215 2920
rect 12425 2940 12455 2945
rect 12425 2920 12430 2940
rect 12430 2920 12450 2940
rect 12450 2920 12455 2940
rect 12425 2915 12455 2920
rect 12485 2915 12515 2945
rect 13005 2915 13035 2920
rect 13005 2895 13010 2915
rect 13010 2895 13030 2915
rect 13030 2895 13035 2915
rect 13005 2890 13035 2895
rect 13115 2915 13145 2920
rect 13115 2895 13120 2915
rect 13120 2895 13140 2915
rect 13140 2895 13145 2915
rect 13115 2890 13145 2895
rect 13225 2915 13255 2920
rect 13225 2895 13230 2915
rect 13230 2895 13250 2915
rect 13250 2895 13255 2915
rect 13225 2890 13255 2895
rect 13335 2915 13365 2920
rect 13335 2895 13340 2915
rect 13340 2895 13360 2915
rect 13360 2895 13365 2915
rect 13335 2890 13365 2895
rect 13445 2915 13475 2920
rect 13445 2895 13450 2915
rect 13450 2895 13470 2915
rect 13470 2895 13475 2915
rect 13445 2890 13475 2895
rect 13555 2915 13585 2920
rect 13555 2895 13560 2915
rect 13560 2895 13580 2915
rect 13580 2895 13585 2915
rect 13555 2890 13585 2895
rect 13665 2915 13695 2920
rect 13665 2895 13670 2915
rect 13670 2895 13690 2915
rect 13690 2895 13695 2915
rect 13665 2890 13695 2895
rect 13775 2915 13805 2920
rect 13775 2895 13780 2915
rect 13780 2895 13800 2915
rect 13800 2895 13805 2915
rect 13775 2890 13805 2895
rect 13885 2915 13915 2920
rect 13885 2895 13890 2915
rect 13890 2895 13910 2915
rect 13910 2895 13915 2915
rect 13885 2890 13915 2895
rect 13995 2915 14025 2920
rect 13995 2895 14000 2915
rect 14000 2895 14020 2915
rect 14020 2895 14025 2915
rect 13995 2890 14025 2895
rect 13060 2800 13090 2830
rect 13060 2750 13090 2780
rect 12695 2700 12725 2730
rect 13060 2700 13090 2730
rect 10985 2445 11015 2475
rect 11826 2470 11854 2475
rect 11826 2450 11831 2470
rect 11831 2450 11849 2470
rect 11849 2450 11854 2470
rect 11826 2445 11854 2450
rect 10816 2435 10844 2440
rect 10816 2415 10821 2435
rect 10821 2415 10839 2435
rect 10839 2415 10844 2435
rect 10816 2410 10844 2415
rect 9805 2375 9840 2380
rect 9805 2350 9810 2375
rect 9810 2350 9835 2375
rect 9835 2350 9840 2375
rect 9805 2345 9840 2350
rect 10640 2375 10675 2380
rect 10640 2350 10645 2375
rect 10645 2350 10670 2375
rect 10670 2350 10675 2375
rect 10640 2345 10675 2350
rect 9805 2315 9840 2320
rect 9805 2290 9810 2315
rect 9810 2290 9835 2315
rect 9835 2290 9840 2315
rect 9805 2285 9840 2290
rect 10640 2315 10675 2320
rect 10640 2290 10645 2315
rect 10645 2290 10670 2315
rect 10670 2290 10675 2315
rect 10640 2285 10675 2290
rect 11285 2390 11315 2420
rect 11525 2390 11555 2420
rect 11765 2390 11795 2420
rect 11405 2345 11435 2375
rect 11645 2345 11675 2375
rect 10816 2275 10844 2280
rect 10816 2255 10821 2275
rect 10821 2255 10839 2275
rect 10839 2255 10844 2275
rect 10816 2250 10844 2255
rect 11445 2250 11475 2280
rect 11665 2250 11695 2280
rect 9795 2215 9825 2220
rect 9795 2195 9800 2215
rect 9800 2195 9820 2215
rect 9820 2195 9825 2215
rect 9795 2190 9825 2195
rect 9905 2215 9935 2220
rect 9905 2195 9910 2215
rect 9910 2195 9930 2215
rect 9930 2195 9935 2215
rect 9905 2190 9935 2195
rect 10015 2215 10045 2220
rect 10015 2195 10020 2215
rect 10020 2195 10040 2215
rect 10040 2195 10045 2215
rect 10015 2190 10045 2195
rect 10125 2215 10155 2220
rect 10125 2195 10130 2215
rect 10130 2195 10150 2215
rect 10150 2195 10155 2215
rect 10125 2190 10155 2195
rect 10235 2215 10265 2220
rect 10235 2195 10240 2215
rect 10240 2195 10260 2215
rect 10260 2195 10265 2215
rect 10235 2190 10265 2195
rect 10345 2215 10375 2220
rect 10345 2195 10350 2215
rect 10350 2195 10370 2215
rect 10370 2195 10375 2215
rect 10345 2190 10375 2195
rect 10455 2215 10485 2220
rect 10455 2195 10460 2215
rect 10460 2195 10480 2215
rect 10480 2195 10485 2215
rect 10455 2190 10485 2195
rect 10565 2215 10595 2220
rect 10565 2195 10570 2215
rect 10570 2195 10590 2215
rect 10590 2195 10595 2215
rect 10565 2190 10595 2195
rect 10675 2215 10705 2220
rect 10675 2195 10680 2215
rect 10680 2195 10700 2215
rect 10700 2195 10705 2215
rect 10675 2190 10705 2195
rect 10785 2215 10815 2220
rect 10785 2195 10790 2215
rect 10790 2195 10810 2215
rect 10810 2195 10815 2215
rect 10785 2190 10815 2195
rect 11335 2205 11365 2235
rect 11555 2205 11585 2235
rect 12005 2390 12035 2420
rect 12245 2390 12275 2420
rect 12485 2390 12515 2420
rect 12950 2665 12980 2670
rect 12950 2645 12955 2665
rect 12955 2645 12975 2665
rect 12975 2645 12980 2665
rect 12950 2640 12980 2645
rect 13060 2665 13090 2670
rect 13060 2645 13065 2665
rect 13065 2645 13085 2665
rect 13085 2645 13090 2665
rect 13060 2640 13090 2645
rect 13170 2665 13200 2670
rect 13170 2645 13175 2665
rect 13175 2645 13195 2665
rect 13195 2645 13200 2665
rect 13170 2640 13200 2645
rect 13280 2665 13310 2670
rect 13280 2645 13285 2665
rect 13285 2645 13305 2665
rect 13305 2645 13310 2665
rect 13280 2640 13310 2645
rect 13390 2665 13420 2670
rect 13390 2645 13395 2665
rect 13395 2645 13415 2665
rect 13415 2645 13420 2665
rect 13390 2640 13420 2645
rect 13500 2665 13530 2670
rect 13500 2645 13505 2665
rect 13505 2645 13525 2665
rect 13525 2645 13530 2665
rect 13500 2640 13530 2645
rect 13610 2665 13640 2670
rect 13610 2645 13615 2665
rect 13615 2645 13635 2665
rect 13635 2645 13640 2665
rect 13610 2640 13640 2645
rect 13720 2665 13750 2670
rect 13720 2645 13725 2665
rect 13725 2645 13745 2665
rect 13745 2645 13750 2665
rect 13720 2640 13750 2645
rect 13830 2665 13860 2670
rect 13830 2645 13835 2665
rect 13835 2645 13855 2665
rect 13855 2645 13860 2665
rect 13830 2640 13860 2645
rect 13940 2665 13970 2670
rect 13940 2645 13945 2665
rect 13945 2645 13965 2665
rect 13965 2645 13970 2665
rect 13940 2640 13970 2645
rect 14050 2665 14080 2670
rect 14050 2645 14055 2665
rect 14055 2645 14075 2665
rect 14075 2645 14080 2665
rect 14050 2640 14080 2645
rect 17240 2665 17270 2670
rect 17240 2645 17245 2665
rect 17245 2645 17265 2665
rect 17265 2645 17270 2665
rect 17240 2640 17270 2645
rect 17350 2665 17380 2670
rect 17350 2645 17355 2665
rect 17355 2645 17375 2665
rect 17375 2645 17380 2665
rect 17350 2640 17380 2645
rect 17460 2665 17490 2670
rect 17460 2645 17465 2665
rect 17465 2645 17485 2665
rect 17485 2645 17490 2665
rect 17460 2640 17490 2645
rect 17570 2665 17600 2670
rect 17570 2645 17575 2665
rect 17575 2645 17595 2665
rect 17595 2645 17600 2665
rect 17570 2640 17600 2645
rect 17680 2665 17710 2670
rect 17680 2645 17685 2665
rect 17685 2645 17705 2665
rect 17705 2645 17710 2665
rect 17680 2640 17710 2645
rect 17790 2665 17820 2670
rect 17790 2645 17795 2665
rect 17795 2645 17815 2665
rect 17815 2645 17820 2665
rect 17790 2640 17820 2645
rect 17900 2665 17930 2670
rect 17900 2645 17905 2665
rect 17905 2645 17925 2665
rect 17925 2645 17930 2665
rect 17900 2640 17930 2645
rect 18010 2665 18040 2670
rect 18010 2645 18015 2665
rect 18015 2645 18035 2665
rect 18035 2645 18040 2665
rect 18010 2640 18040 2645
rect 18120 2665 18150 2670
rect 18120 2645 18125 2665
rect 18125 2645 18145 2665
rect 18145 2645 18150 2665
rect 18120 2640 18150 2645
rect 18230 2665 18260 2670
rect 18230 2645 18235 2665
rect 18235 2645 18255 2665
rect 18255 2645 18260 2665
rect 18230 2640 18260 2645
rect 18340 2665 18370 2670
rect 18340 2645 18345 2665
rect 18345 2645 18365 2665
rect 18365 2645 18370 2665
rect 18340 2640 18370 2645
rect 13005 2495 13035 2500
rect 13005 2475 13010 2495
rect 13010 2475 13030 2495
rect 13030 2475 13035 2495
rect 13005 2470 13035 2475
rect 13115 2495 13145 2500
rect 13115 2475 13120 2495
rect 13120 2475 13140 2495
rect 13140 2475 13145 2495
rect 13115 2470 13145 2475
rect 13225 2495 13255 2500
rect 13225 2475 13230 2495
rect 13230 2475 13250 2495
rect 13250 2475 13255 2495
rect 13225 2470 13255 2475
rect 13335 2495 13365 2500
rect 13335 2475 13340 2495
rect 13340 2475 13360 2495
rect 13360 2475 13365 2495
rect 13335 2470 13365 2475
rect 13445 2495 13475 2500
rect 13445 2475 13450 2495
rect 13450 2475 13470 2495
rect 13470 2475 13475 2495
rect 13445 2470 13475 2475
rect 13555 2495 13585 2500
rect 13555 2475 13560 2495
rect 13560 2475 13580 2495
rect 13580 2475 13585 2495
rect 13555 2470 13585 2475
rect 13665 2495 13695 2500
rect 13665 2475 13670 2495
rect 13670 2475 13690 2495
rect 13690 2475 13695 2495
rect 13665 2470 13695 2475
rect 13775 2495 13805 2500
rect 13775 2475 13780 2495
rect 13780 2475 13800 2495
rect 13800 2475 13805 2495
rect 13775 2470 13805 2475
rect 13885 2495 13915 2500
rect 13885 2475 13890 2495
rect 13890 2475 13910 2495
rect 13910 2475 13915 2495
rect 13885 2470 13915 2475
rect 13995 2495 14025 2500
rect 13995 2475 14000 2495
rect 14000 2475 14020 2495
rect 14020 2475 14025 2495
rect 13995 2470 14025 2475
rect 17295 2495 17325 2500
rect 17295 2475 17300 2495
rect 17300 2475 17320 2495
rect 17320 2475 17325 2495
rect 17295 2470 17325 2475
rect 17405 2495 17435 2500
rect 17405 2475 17410 2495
rect 17410 2475 17430 2495
rect 17430 2475 17435 2495
rect 17405 2470 17435 2475
rect 17515 2495 17545 2500
rect 17515 2475 17520 2495
rect 17520 2475 17540 2495
rect 17540 2475 17545 2495
rect 17515 2470 17545 2475
rect 17625 2495 17655 2500
rect 17625 2475 17630 2495
rect 17630 2475 17650 2495
rect 17650 2475 17655 2495
rect 17625 2470 17655 2475
rect 17735 2495 17765 2500
rect 17735 2475 17740 2495
rect 17740 2475 17760 2495
rect 17760 2475 17765 2495
rect 17735 2470 17765 2475
rect 17845 2495 17875 2500
rect 17845 2475 17850 2495
rect 17850 2475 17870 2495
rect 17870 2475 17875 2495
rect 17845 2470 17875 2475
rect 17955 2495 17985 2500
rect 17955 2475 17960 2495
rect 17960 2475 17980 2495
rect 17980 2475 17985 2495
rect 17955 2470 17985 2475
rect 18065 2495 18095 2500
rect 18065 2475 18070 2495
rect 18070 2475 18090 2495
rect 18090 2475 18095 2495
rect 18065 2470 18095 2475
rect 18175 2495 18205 2500
rect 18175 2475 18180 2495
rect 18180 2475 18200 2495
rect 18200 2475 18205 2495
rect 18175 2470 18205 2475
rect 18285 2495 18315 2500
rect 18285 2475 18290 2495
rect 18290 2475 18310 2495
rect 18310 2475 18315 2495
rect 18285 2470 18315 2475
rect 19326 3150 19354 3155
rect 19326 3130 19331 3150
rect 19331 3130 19349 3150
rect 19349 3130 19354 3150
rect 19326 3125 19354 3130
rect 18785 3070 18815 3100
rect 19025 3070 19055 3100
rect 19265 3070 19295 3100
rect 19505 3070 19535 3100
rect 19745 3070 19775 3100
rect 19985 3070 20015 3100
rect 18905 3025 18935 3055
rect 19145 3025 19175 3055
rect 19385 3025 19415 3055
rect 19625 3025 19655 3055
rect 19865 3025 19895 3055
rect 18845 2970 18875 3000
rect 18905 2970 18935 3000
rect 19085 2970 19115 3000
rect 19325 2970 19355 3000
rect 19565 2970 19595 3000
rect 19805 2970 19835 3000
rect 18965 2940 18995 2945
rect 18965 2920 18970 2940
rect 18970 2920 18990 2940
rect 18990 2920 18995 2940
rect 18965 2915 18995 2920
rect 19205 2940 19235 2945
rect 19205 2920 19210 2940
rect 19210 2920 19230 2940
rect 19230 2920 19235 2940
rect 19205 2915 19235 2920
rect 19445 2940 19475 2945
rect 19445 2920 19450 2940
rect 19450 2920 19470 2940
rect 19470 2920 19475 2940
rect 19445 2915 19475 2920
rect 19685 2940 19715 2945
rect 19685 2920 19690 2940
rect 19690 2920 19710 2940
rect 19710 2920 19715 2940
rect 19685 2915 19715 2920
rect 19925 2940 19955 2945
rect 19925 2920 19930 2940
rect 19930 2920 19950 2940
rect 19950 2920 19955 2940
rect 19925 2915 19955 2920
rect 19985 2915 20015 2945
rect 20505 2915 20535 2920
rect 20505 2895 20510 2915
rect 20510 2895 20530 2915
rect 20530 2895 20535 2915
rect 20505 2890 20535 2895
rect 20615 2915 20645 2920
rect 20615 2895 20620 2915
rect 20620 2895 20640 2915
rect 20640 2895 20645 2915
rect 20615 2890 20645 2895
rect 20725 2915 20755 2920
rect 20725 2895 20730 2915
rect 20730 2895 20750 2915
rect 20750 2895 20755 2915
rect 20725 2890 20755 2895
rect 20835 2915 20865 2920
rect 20835 2895 20840 2915
rect 20840 2895 20860 2915
rect 20860 2895 20865 2915
rect 20835 2890 20865 2895
rect 20945 2915 20975 2920
rect 20945 2895 20950 2915
rect 20950 2895 20970 2915
rect 20970 2895 20975 2915
rect 20945 2890 20975 2895
rect 21055 2915 21085 2920
rect 21055 2895 21060 2915
rect 21060 2895 21080 2915
rect 21080 2895 21085 2915
rect 21055 2890 21085 2895
rect 21165 2915 21195 2920
rect 21165 2895 21170 2915
rect 21170 2895 21190 2915
rect 21190 2895 21195 2915
rect 21165 2890 21195 2895
rect 21275 2915 21305 2920
rect 21275 2895 21280 2915
rect 21280 2895 21300 2915
rect 21300 2895 21305 2915
rect 21275 2890 21305 2895
rect 21385 2915 21415 2920
rect 21385 2895 21390 2915
rect 21390 2895 21410 2915
rect 21410 2895 21415 2915
rect 21385 2890 21415 2895
rect 21495 2915 21525 2920
rect 21495 2895 21500 2915
rect 21500 2895 21520 2915
rect 21520 2895 21525 2915
rect 21495 2890 21525 2895
rect 20560 2800 20590 2830
rect 20560 2750 20590 2780
rect 20195 2700 20225 2730
rect 20560 2700 20590 2730
rect 12976 2435 13004 2440
rect 12976 2415 12981 2435
rect 12981 2415 12999 2435
rect 12999 2415 13004 2435
rect 12976 2410 13004 2415
rect 11885 2345 11915 2375
rect 12125 2345 12155 2375
rect 12365 2345 12395 2375
rect 12695 2345 12725 2375
rect 12975 2345 13005 2375
rect 13145 2375 13180 2380
rect 13145 2350 13150 2375
rect 13150 2350 13175 2375
rect 13175 2350 13180 2375
rect 13145 2345 13180 2350
rect 13980 2375 14015 2380
rect 13980 2350 13985 2375
rect 13985 2350 14010 2375
rect 14010 2350 14015 2375
rect 13980 2345 14015 2350
rect 18485 2445 18515 2475
rect 19326 2470 19354 2475
rect 19326 2450 19331 2470
rect 19331 2450 19349 2470
rect 19349 2450 19354 2470
rect 19326 2445 19354 2450
rect 18316 2435 18344 2440
rect 18316 2415 18321 2435
rect 18321 2415 18339 2435
rect 18339 2415 18344 2435
rect 18316 2410 18344 2415
rect 17305 2375 17340 2380
rect 17305 2350 17310 2375
rect 17310 2350 17335 2375
rect 17335 2350 17340 2375
rect 17305 2345 17340 2350
rect 18140 2375 18175 2380
rect 18140 2350 18145 2375
rect 18145 2350 18170 2375
rect 18170 2350 18175 2375
rect 18140 2345 18175 2350
rect 12820 2295 12850 2325
rect 11885 2250 11915 2280
rect 12105 2250 12135 2280
rect 12325 2250 12355 2280
rect 11775 2205 11805 2235
rect 11995 2205 12025 2235
rect 12215 2205 12245 2235
rect 12435 2205 12465 2235
rect 9740 1995 9770 2000
rect 9740 1975 9745 1995
rect 9745 1975 9763 1995
rect 9763 1975 9770 1995
rect 9740 1970 9770 1975
rect 9850 1995 9880 2000
rect 9850 1975 9855 1995
rect 9855 1975 9873 1995
rect 9873 1975 9880 1995
rect 9850 1970 9880 1975
rect 9960 1995 9990 2000
rect 9960 1975 9965 1995
rect 9965 1975 9983 1995
rect 9983 1975 9990 1995
rect 9960 1970 9990 1975
rect 10070 1995 10100 2000
rect 10070 1975 10075 1995
rect 10075 1975 10093 1995
rect 10093 1975 10100 1995
rect 10070 1970 10100 1975
rect 10180 1995 10210 2000
rect 10180 1975 10185 1995
rect 10185 1975 10203 1995
rect 10203 1975 10210 1995
rect 10180 1970 10210 1975
rect 10290 1995 10320 2000
rect 10290 1975 10295 1995
rect 10295 1975 10313 1995
rect 10313 1975 10320 1995
rect 10290 1970 10320 1975
rect 10400 1995 10430 2000
rect 10400 1975 10405 1995
rect 10405 1975 10423 1995
rect 10423 1975 10430 1995
rect 10400 1970 10430 1975
rect 10510 1995 10540 2000
rect 10510 1975 10515 1995
rect 10515 1975 10533 1995
rect 10533 1975 10540 1995
rect 10510 1970 10540 1975
rect 10620 1995 10650 2000
rect 10620 1975 10625 1995
rect 10625 1975 10643 1995
rect 10643 1975 10650 1995
rect 10620 1970 10650 1975
rect 10730 1995 10760 2000
rect 10730 1975 10735 1995
rect 10735 1975 10753 1995
rect 10753 1975 10760 1995
rect 10730 1970 10760 1975
rect 10840 1995 10870 2000
rect 10840 1975 10845 1995
rect 10845 1975 10863 1995
rect 10863 1975 10870 1995
rect 10840 1970 10870 1975
rect 11390 1955 11420 1960
rect 11390 1935 11395 1955
rect 11395 1935 11415 1955
rect 11415 1935 11420 1955
rect 11390 1930 11420 1935
rect 11610 1955 11640 1960
rect 11610 1935 11615 1955
rect 11615 1935 11635 1955
rect 11635 1935 11640 1955
rect 11610 1930 11640 1935
rect 11830 1955 11860 1960
rect 11830 1935 11835 1955
rect 11835 1935 11855 1955
rect 11855 1935 11860 1955
rect 11830 1930 11860 1935
rect 12050 1955 12080 1960
rect 12050 1935 12055 1955
rect 12055 1935 12075 1955
rect 12075 1935 12080 1955
rect 12050 1930 12080 1935
rect 12270 1955 12300 1960
rect 12270 1935 12275 1955
rect 12275 1935 12295 1955
rect 12295 1935 12300 1955
rect 12270 1930 12300 1935
rect 11500 1875 11530 1905
rect 11720 1875 11750 1905
rect 11940 1875 11970 1905
rect 12160 1875 12190 1905
rect 11195 1820 11225 1850
rect 11415 1820 11445 1850
rect 11090 1755 11120 1760
rect 11090 1735 11095 1755
rect 11095 1735 11115 1755
rect 11115 1735 11120 1755
rect 11090 1730 11120 1735
rect 11310 1755 11340 1760
rect 11310 1735 11315 1755
rect 11315 1735 11335 1755
rect 11335 1735 11340 1755
rect 11310 1730 11340 1735
rect 12380 1875 12410 1905
rect 11645 1820 11675 1850
rect 12235 1820 12265 1850
rect 12455 1820 12485 1850
rect 12685 1820 12715 1850
rect 11825 1775 11855 1805
rect 11945 1775 11975 1805
rect 11530 1755 11560 1760
rect 11530 1735 11535 1755
rect 11535 1735 11555 1755
rect 11555 1735 11560 1755
rect 11530 1730 11560 1735
rect 12130 1755 12160 1760
rect 12130 1735 12135 1755
rect 12135 1735 12155 1755
rect 12155 1735 12160 1755
rect 12130 1730 12160 1735
rect 12350 1755 12380 1760
rect 12350 1735 12355 1755
rect 12355 1735 12375 1755
rect 12375 1735 12380 1755
rect 12350 1730 12380 1735
rect 12570 1755 12600 1760
rect 12570 1735 12575 1755
rect 12575 1735 12595 1755
rect 12595 1735 12600 1755
rect 12570 1730 12600 1735
rect 11240 1710 11266 1715
rect 11240 1690 11243 1710
rect 11243 1690 11260 1710
rect 11260 1690 11266 1710
rect 11240 1685 11266 1690
rect 11460 1710 11486 1715
rect 11460 1690 11463 1710
rect 11463 1690 11480 1710
rect 11480 1690 11486 1710
rect 11460 1685 11486 1690
rect 11604 1710 11630 1715
rect 11604 1690 11610 1710
rect 11610 1690 11627 1710
rect 11627 1690 11630 1710
rect 11604 1685 11630 1690
rect 11870 1710 11896 1715
rect 11870 1690 11876 1710
rect 11876 1690 11893 1710
rect 11893 1690 11896 1710
rect 11870 1685 11896 1690
rect 12280 1710 12306 1715
rect 12280 1690 12283 1710
rect 12283 1690 12300 1710
rect 12300 1690 12306 1710
rect 12280 1685 12306 1690
rect 12500 1710 12526 1715
rect 12500 1690 12503 1710
rect 12503 1690 12520 1710
rect 12520 1690 12526 1710
rect 12500 1685 12526 1690
rect 12644 1710 12670 1715
rect 12644 1690 12650 1710
rect 12650 1690 12667 1710
rect 12667 1690 12670 1710
rect 12644 1685 12670 1690
rect 4810 1590 4840 1595
rect 4810 1570 4815 1590
rect 4815 1570 4835 1590
rect 4835 1570 4840 1590
rect 4810 1565 4840 1570
rect 5415 1565 5445 1595
rect 13145 2315 13180 2320
rect 13145 2290 13150 2315
rect 13150 2290 13175 2315
rect 13175 2290 13180 2315
rect 13145 2285 13180 2290
rect 13980 2315 14015 2320
rect 13980 2290 13985 2315
rect 13985 2290 14010 2315
rect 14010 2290 14015 2315
rect 13980 2285 14015 2290
rect 12976 2275 13004 2280
rect 12976 2255 12981 2275
rect 12981 2255 12999 2275
rect 12999 2255 13004 2275
rect 12976 2250 13004 2255
rect 17305 2315 17340 2320
rect 17305 2290 17310 2315
rect 17310 2290 17335 2315
rect 17335 2290 17340 2315
rect 17305 2285 17340 2290
rect 18140 2315 18175 2320
rect 18140 2290 18145 2315
rect 18145 2290 18170 2315
rect 18170 2290 18175 2315
rect 18140 2285 18175 2290
rect 18785 2390 18815 2420
rect 19025 2390 19055 2420
rect 19265 2390 19295 2420
rect 18905 2345 18935 2375
rect 19145 2345 19175 2375
rect 18316 2275 18344 2280
rect 18316 2255 18321 2275
rect 18321 2255 18339 2275
rect 18339 2255 18344 2275
rect 18316 2250 18344 2255
rect 18945 2250 18975 2280
rect 19165 2250 19195 2280
rect 13005 2215 13035 2220
rect 13005 2195 13010 2215
rect 13010 2195 13030 2215
rect 13030 2195 13035 2215
rect 13005 2190 13035 2195
rect 13115 2215 13145 2220
rect 13115 2195 13120 2215
rect 13120 2195 13140 2215
rect 13140 2195 13145 2215
rect 13115 2190 13145 2195
rect 13225 2215 13255 2220
rect 13225 2195 13230 2215
rect 13230 2195 13250 2215
rect 13250 2195 13255 2215
rect 13225 2190 13255 2195
rect 13335 2215 13365 2220
rect 13335 2195 13340 2215
rect 13340 2195 13360 2215
rect 13360 2195 13365 2215
rect 13335 2190 13365 2195
rect 13445 2215 13475 2220
rect 13445 2195 13450 2215
rect 13450 2195 13470 2215
rect 13470 2195 13475 2215
rect 13445 2190 13475 2195
rect 13555 2215 13585 2220
rect 13555 2195 13560 2215
rect 13560 2195 13580 2215
rect 13580 2195 13585 2215
rect 13555 2190 13585 2195
rect 13665 2215 13695 2220
rect 13665 2195 13670 2215
rect 13670 2195 13690 2215
rect 13690 2195 13695 2215
rect 13665 2190 13695 2195
rect 13775 2215 13805 2220
rect 13775 2195 13780 2215
rect 13780 2195 13800 2215
rect 13800 2195 13805 2215
rect 13775 2190 13805 2195
rect 13885 2215 13915 2220
rect 13885 2195 13890 2215
rect 13890 2195 13910 2215
rect 13910 2195 13915 2215
rect 13885 2190 13915 2195
rect 13995 2215 14025 2220
rect 13995 2195 14000 2215
rect 14000 2195 14020 2215
rect 14020 2195 14025 2215
rect 13995 2190 14025 2195
rect 17295 2215 17325 2220
rect 17295 2195 17300 2215
rect 17300 2195 17320 2215
rect 17320 2195 17325 2215
rect 17295 2190 17325 2195
rect 17405 2215 17435 2220
rect 17405 2195 17410 2215
rect 17410 2195 17430 2215
rect 17430 2195 17435 2215
rect 17405 2190 17435 2195
rect 17515 2215 17545 2220
rect 17515 2195 17520 2215
rect 17520 2195 17540 2215
rect 17540 2195 17545 2215
rect 17515 2190 17545 2195
rect 17625 2215 17655 2220
rect 17625 2195 17630 2215
rect 17630 2195 17650 2215
rect 17650 2195 17655 2215
rect 17625 2190 17655 2195
rect 17735 2215 17765 2220
rect 17735 2195 17740 2215
rect 17740 2195 17760 2215
rect 17760 2195 17765 2215
rect 17735 2190 17765 2195
rect 17845 2215 17875 2220
rect 17845 2195 17850 2215
rect 17850 2195 17870 2215
rect 17870 2195 17875 2215
rect 17845 2190 17875 2195
rect 17955 2215 17985 2220
rect 17955 2195 17960 2215
rect 17960 2195 17980 2215
rect 17980 2195 17985 2215
rect 17955 2190 17985 2195
rect 18065 2215 18095 2220
rect 18065 2195 18070 2215
rect 18070 2195 18090 2215
rect 18090 2195 18095 2215
rect 18065 2190 18095 2195
rect 18175 2215 18205 2220
rect 18175 2195 18180 2215
rect 18180 2195 18200 2215
rect 18200 2195 18205 2215
rect 18175 2190 18205 2195
rect 18285 2215 18315 2220
rect 18285 2195 18290 2215
rect 18290 2195 18310 2215
rect 18310 2195 18315 2215
rect 18285 2190 18315 2195
rect 18835 2205 18865 2235
rect 19055 2205 19085 2235
rect 19505 2390 19535 2420
rect 19745 2390 19775 2420
rect 19985 2390 20015 2420
rect 20450 2665 20480 2670
rect 20450 2645 20455 2665
rect 20455 2645 20475 2665
rect 20475 2645 20480 2665
rect 20450 2640 20480 2645
rect 20560 2665 20590 2670
rect 20560 2645 20565 2665
rect 20565 2645 20585 2665
rect 20585 2645 20590 2665
rect 20560 2640 20590 2645
rect 20670 2665 20700 2670
rect 20670 2645 20675 2665
rect 20675 2645 20695 2665
rect 20695 2645 20700 2665
rect 20670 2640 20700 2645
rect 20780 2665 20810 2670
rect 20780 2645 20785 2665
rect 20785 2645 20805 2665
rect 20805 2645 20810 2665
rect 20780 2640 20810 2645
rect 20890 2665 20920 2670
rect 20890 2645 20895 2665
rect 20895 2645 20915 2665
rect 20915 2645 20920 2665
rect 20890 2640 20920 2645
rect 21000 2665 21030 2670
rect 21000 2645 21005 2665
rect 21005 2645 21025 2665
rect 21025 2645 21030 2665
rect 21000 2640 21030 2645
rect 21110 2665 21140 2670
rect 21110 2645 21115 2665
rect 21115 2645 21135 2665
rect 21135 2645 21140 2665
rect 21110 2640 21140 2645
rect 21220 2665 21250 2670
rect 21220 2645 21225 2665
rect 21225 2645 21245 2665
rect 21245 2645 21250 2665
rect 21220 2640 21250 2645
rect 21330 2665 21360 2670
rect 21330 2645 21335 2665
rect 21335 2645 21355 2665
rect 21355 2645 21360 2665
rect 21330 2640 21360 2645
rect 21440 2665 21470 2670
rect 21440 2645 21445 2665
rect 21445 2645 21465 2665
rect 21465 2645 21470 2665
rect 21440 2640 21470 2645
rect 21550 2665 21580 2670
rect 21550 2645 21555 2665
rect 21555 2645 21575 2665
rect 21575 2645 21580 2665
rect 21550 2640 21580 2645
rect 20505 2495 20535 2500
rect 20505 2475 20510 2495
rect 20510 2475 20530 2495
rect 20530 2475 20535 2495
rect 20505 2470 20535 2475
rect 20615 2495 20645 2500
rect 20615 2475 20620 2495
rect 20620 2475 20640 2495
rect 20640 2475 20645 2495
rect 20615 2470 20645 2475
rect 20725 2495 20755 2500
rect 20725 2475 20730 2495
rect 20730 2475 20750 2495
rect 20750 2475 20755 2495
rect 20725 2470 20755 2475
rect 20835 2495 20865 2500
rect 20835 2475 20840 2495
rect 20840 2475 20860 2495
rect 20860 2475 20865 2495
rect 20835 2470 20865 2475
rect 20945 2495 20975 2500
rect 20945 2475 20950 2495
rect 20950 2475 20970 2495
rect 20970 2475 20975 2495
rect 20945 2470 20975 2475
rect 21055 2495 21085 2500
rect 21055 2475 21060 2495
rect 21060 2475 21080 2495
rect 21080 2475 21085 2495
rect 21055 2470 21085 2475
rect 21165 2495 21195 2500
rect 21165 2475 21170 2495
rect 21170 2475 21190 2495
rect 21190 2475 21195 2495
rect 21165 2470 21195 2475
rect 21275 2495 21305 2500
rect 21275 2475 21280 2495
rect 21280 2475 21300 2495
rect 21300 2475 21305 2495
rect 21275 2470 21305 2475
rect 21385 2495 21415 2500
rect 21385 2475 21390 2495
rect 21390 2475 21410 2495
rect 21410 2475 21415 2495
rect 21385 2470 21415 2475
rect 21495 2495 21525 2500
rect 21495 2475 21500 2495
rect 21500 2475 21520 2495
rect 21520 2475 21525 2495
rect 21495 2470 21525 2475
rect 20476 2435 20504 2440
rect 20476 2415 20481 2435
rect 20481 2415 20499 2435
rect 20499 2415 20504 2435
rect 20476 2410 20504 2415
rect 19385 2345 19415 2375
rect 19625 2345 19655 2375
rect 19865 2345 19895 2375
rect 20195 2345 20225 2375
rect 20475 2345 20505 2375
rect 20645 2375 20680 2380
rect 20645 2350 20650 2375
rect 20650 2350 20675 2375
rect 20675 2350 20680 2375
rect 20645 2345 20680 2350
rect 21480 2375 21515 2380
rect 21480 2350 21485 2375
rect 21485 2350 21510 2375
rect 21510 2350 21515 2375
rect 21480 2345 21515 2350
rect 20320 2295 20350 2325
rect 19385 2250 19415 2280
rect 19605 2250 19635 2280
rect 19825 2250 19855 2280
rect 19275 2205 19305 2235
rect 19495 2205 19525 2235
rect 19715 2205 19745 2235
rect 19935 2205 19965 2235
rect 12950 1995 12980 2000
rect 12950 1975 12957 1995
rect 12957 1975 12975 1995
rect 12975 1975 12980 1995
rect 12950 1970 12980 1975
rect 13060 1995 13090 2000
rect 13060 1975 13067 1995
rect 13067 1975 13085 1995
rect 13085 1975 13090 1995
rect 13060 1970 13090 1975
rect 13170 1995 13200 2000
rect 13170 1975 13177 1995
rect 13177 1975 13195 1995
rect 13195 1975 13200 1995
rect 13170 1970 13200 1975
rect 13280 1995 13310 2000
rect 13280 1975 13287 1995
rect 13287 1975 13305 1995
rect 13305 1975 13310 1995
rect 13280 1970 13310 1975
rect 13390 1995 13420 2000
rect 13390 1975 13397 1995
rect 13397 1975 13415 1995
rect 13415 1975 13420 1995
rect 13390 1970 13420 1975
rect 13500 1995 13530 2000
rect 13500 1975 13507 1995
rect 13507 1975 13525 1995
rect 13525 1975 13530 1995
rect 13500 1970 13530 1975
rect 13610 1995 13640 2000
rect 13610 1975 13617 1995
rect 13617 1975 13635 1995
rect 13635 1975 13640 1995
rect 13610 1970 13640 1975
rect 13720 1995 13750 2000
rect 13720 1975 13727 1995
rect 13727 1975 13745 1995
rect 13745 1975 13750 1995
rect 13720 1970 13750 1975
rect 13830 1995 13860 2000
rect 13830 1975 13837 1995
rect 13837 1975 13855 1995
rect 13855 1975 13860 1995
rect 13830 1970 13860 1975
rect 13940 1995 13970 2000
rect 13940 1975 13947 1995
rect 13947 1975 13965 1995
rect 13965 1975 13970 1995
rect 13940 1970 13970 1975
rect 14050 1995 14080 2000
rect 14050 1975 14057 1995
rect 14057 1975 14075 1995
rect 14075 1975 14080 1995
rect 14050 1970 14080 1975
rect 17240 1995 17270 2000
rect 17240 1975 17245 1995
rect 17245 1975 17263 1995
rect 17263 1975 17270 1995
rect 17240 1970 17270 1975
rect 17350 1995 17380 2000
rect 17350 1975 17355 1995
rect 17355 1975 17373 1995
rect 17373 1975 17380 1995
rect 17350 1970 17380 1975
rect 17460 1995 17490 2000
rect 17460 1975 17465 1995
rect 17465 1975 17483 1995
rect 17483 1975 17490 1995
rect 17460 1970 17490 1975
rect 17570 1995 17600 2000
rect 17570 1975 17575 1995
rect 17575 1975 17593 1995
rect 17593 1975 17600 1995
rect 17570 1970 17600 1975
rect 17680 1995 17710 2000
rect 17680 1975 17685 1995
rect 17685 1975 17703 1995
rect 17703 1975 17710 1995
rect 17680 1970 17710 1975
rect 17790 1995 17820 2000
rect 17790 1975 17795 1995
rect 17795 1975 17813 1995
rect 17813 1975 17820 1995
rect 17790 1970 17820 1975
rect 17900 1995 17930 2000
rect 17900 1975 17905 1995
rect 17905 1975 17923 1995
rect 17923 1975 17930 1995
rect 17900 1970 17930 1975
rect 18010 1995 18040 2000
rect 18010 1975 18015 1995
rect 18015 1975 18033 1995
rect 18033 1975 18040 1995
rect 18010 1970 18040 1975
rect 18120 1995 18150 2000
rect 18120 1975 18125 1995
rect 18125 1975 18143 1995
rect 18143 1975 18150 1995
rect 18120 1970 18150 1975
rect 18230 1995 18260 2000
rect 18230 1975 18235 1995
rect 18235 1975 18253 1995
rect 18253 1975 18260 1995
rect 18230 1970 18260 1975
rect 18340 1995 18370 2000
rect 18340 1975 18345 1995
rect 18345 1975 18363 1995
rect 18363 1975 18370 1995
rect 18340 1970 18370 1975
rect 18890 1955 18920 1960
rect 18890 1935 18895 1955
rect 18895 1935 18915 1955
rect 18915 1935 18920 1955
rect 18890 1930 18920 1935
rect 19110 1955 19140 1960
rect 19110 1935 19115 1955
rect 19115 1935 19135 1955
rect 19135 1935 19140 1955
rect 19110 1930 19140 1935
rect 19330 1955 19360 1960
rect 19330 1935 19335 1955
rect 19335 1935 19355 1955
rect 19355 1935 19360 1955
rect 19330 1930 19360 1935
rect 19550 1955 19580 1960
rect 19550 1935 19555 1955
rect 19555 1935 19575 1955
rect 19575 1935 19580 1955
rect 19550 1930 19580 1935
rect 19770 1955 19800 1960
rect 19770 1935 19775 1955
rect 19775 1935 19795 1955
rect 19795 1935 19800 1955
rect 19770 1930 19800 1935
rect 19000 1875 19030 1905
rect 19220 1875 19250 1905
rect 19440 1875 19470 1905
rect 19660 1875 19690 1905
rect 18695 1820 18725 1850
rect 18915 1820 18945 1850
rect 18590 1755 18620 1760
rect 18590 1735 18595 1755
rect 18595 1735 18615 1755
rect 18615 1735 18620 1755
rect 18590 1730 18620 1735
rect 18810 1755 18840 1760
rect 18810 1735 18815 1755
rect 18815 1735 18835 1755
rect 18835 1735 18840 1755
rect 18810 1730 18840 1735
rect 19880 1875 19910 1905
rect 19145 1820 19175 1850
rect 19735 1820 19765 1850
rect 19955 1820 19985 1850
rect 20185 1820 20215 1850
rect 19325 1775 19355 1805
rect 19445 1775 19475 1805
rect 19030 1755 19060 1760
rect 19030 1735 19035 1755
rect 19035 1735 19055 1755
rect 19055 1735 19060 1755
rect 19030 1730 19060 1735
rect 19630 1755 19660 1760
rect 19630 1735 19635 1755
rect 19635 1735 19655 1755
rect 19655 1735 19660 1755
rect 19630 1730 19660 1735
rect 19850 1755 19880 1760
rect 19850 1735 19855 1755
rect 19855 1735 19875 1755
rect 19875 1735 19880 1755
rect 19850 1730 19880 1735
rect 20070 1755 20100 1760
rect 20070 1735 20075 1755
rect 20075 1735 20095 1755
rect 20095 1735 20100 1755
rect 20070 1730 20100 1735
rect 18740 1710 18766 1715
rect 18740 1690 18743 1710
rect 18743 1690 18760 1710
rect 18760 1690 18766 1710
rect 18740 1685 18766 1690
rect 18960 1710 18986 1715
rect 18960 1690 18963 1710
rect 18963 1690 18980 1710
rect 18980 1690 18986 1710
rect 18960 1685 18986 1690
rect 19104 1710 19130 1715
rect 19104 1690 19110 1710
rect 19110 1690 19127 1710
rect 19127 1690 19130 1710
rect 19104 1685 19130 1690
rect 19370 1710 19396 1715
rect 19370 1690 19376 1710
rect 19376 1690 19393 1710
rect 19393 1690 19396 1710
rect 19370 1685 19396 1690
rect 19780 1710 19806 1715
rect 19780 1690 19783 1710
rect 19783 1690 19800 1710
rect 19800 1690 19806 1710
rect 19780 1685 19806 1690
rect 20000 1710 20026 1715
rect 20000 1690 20003 1710
rect 20003 1690 20020 1710
rect 20020 1690 20026 1710
rect 20000 1685 20026 1690
rect 20144 1710 20170 1715
rect 20144 1690 20150 1710
rect 20150 1690 20167 1710
rect 20167 1690 20170 1710
rect 20144 1685 20170 1690
rect 20645 2315 20680 2320
rect 20645 2290 20650 2315
rect 20650 2290 20675 2315
rect 20675 2290 20680 2315
rect 20645 2285 20680 2290
rect 21480 2315 21515 2320
rect 21480 2290 21485 2315
rect 21485 2290 21510 2315
rect 21510 2290 21515 2315
rect 21480 2285 21515 2290
rect 20476 2275 20504 2280
rect 20476 2255 20481 2275
rect 20481 2255 20499 2275
rect 20499 2255 20504 2275
rect 20476 2250 20504 2255
rect 20505 2215 20535 2220
rect 20505 2195 20510 2215
rect 20510 2195 20530 2215
rect 20530 2195 20535 2215
rect 20505 2190 20535 2195
rect 20615 2215 20645 2220
rect 20615 2195 20620 2215
rect 20620 2195 20640 2215
rect 20640 2195 20645 2215
rect 20615 2190 20645 2195
rect 20725 2215 20755 2220
rect 20725 2195 20730 2215
rect 20730 2195 20750 2215
rect 20750 2195 20755 2215
rect 20725 2190 20755 2195
rect 20835 2215 20865 2220
rect 20835 2195 20840 2215
rect 20840 2195 20860 2215
rect 20860 2195 20865 2215
rect 20835 2190 20865 2195
rect 20945 2215 20975 2220
rect 20945 2195 20950 2215
rect 20950 2195 20970 2215
rect 20970 2195 20975 2215
rect 20945 2190 20975 2195
rect 21055 2215 21085 2220
rect 21055 2195 21060 2215
rect 21060 2195 21080 2215
rect 21080 2195 21085 2215
rect 21055 2190 21085 2195
rect 21165 2215 21195 2220
rect 21165 2195 21170 2215
rect 21170 2195 21190 2215
rect 21190 2195 21195 2215
rect 21165 2190 21195 2195
rect 21275 2215 21305 2220
rect 21275 2195 21280 2215
rect 21280 2195 21300 2215
rect 21300 2195 21305 2215
rect 21275 2190 21305 2195
rect 21385 2215 21415 2220
rect 21385 2195 21390 2215
rect 21390 2195 21410 2215
rect 21410 2195 21415 2215
rect 21385 2190 21415 2195
rect 21495 2215 21525 2220
rect 21495 2195 21500 2215
rect 21500 2195 21520 2215
rect 21520 2195 21525 2215
rect 21495 2190 21525 2195
rect 20450 1995 20480 2000
rect 20450 1975 20457 1995
rect 20457 1975 20475 1995
rect 20475 1975 20480 1995
rect 20450 1970 20480 1975
rect 20560 1995 20590 2000
rect 20560 1975 20567 1995
rect 20567 1975 20585 1995
rect 20585 1975 20590 1995
rect 20560 1970 20590 1975
rect 20670 1995 20700 2000
rect 20670 1975 20677 1995
rect 20677 1975 20695 1995
rect 20695 1975 20700 1995
rect 20670 1970 20700 1975
rect 20780 1995 20810 2000
rect 20780 1975 20787 1995
rect 20787 1975 20805 1995
rect 20805 1975 20810 1995
rect 20780 1970 20810 1975
rect 20890 1995 20920 2000
rect 20890 1975 20897 1995
rect 20897 1975 20915 1995
rect 20915 1975 20920 1995
rect 20890 1970 20920 1975
rect 21000 1995 21030 2000
rect 21000 1975 21007 1995
rect 21007 1975 21025 1995
rect 21025 1975 21030 1995
rect 21000 1970 21030 1975
rect 21110 1995 21140 2000
rect 21110 1975 21117 1995
rect 21117 1975 21135 1995
rect 21135 1975 21140 1995
rect 21110 1970 21140 1975
rect 21220 1995 21250 2000
rect 21220 1975 21227 1995
rect 21227 1975 21245 1995
rect 21245 1975 21250 1995
rect 21220 1970 21250 1975
rect 21330 1995 21360 2000
rect 21330 1975 21337 1995
rect 21337 1975 21355 1995
rect 21355 1975 21360 1995
rect 21330 1970 21360 1975
rect 21440 1995 21470 2000
rect 21440 1975 21447 1995
rect 21447 1975 21465 1995
rect 21465 1975 21470 1995
rect 21440 1970 21470 1975
rect 21550 1995 21580 2000
rect 21550 1975 21557 1995
rect 21557 1975 21575 1995
rect 21575 1975 21580 1995
rect 21550 1970 21580 1975
rect 20550 1900 20580 1905
rect 20550 1880 20555 1900
rect 20555 1880 20575 1900
rect 20575 1880 20580 1900
rect 20550 1875 20580 1880
rect 20660 1900 20690 1905
rect 20660 1880 20665 1900
rect 20665 1880 20685 1900
rect 20685 1880 20690 1900
rect 20660 1875 20690 1880
rect 20770 1900 20800 1905
rect 20770 1880 20775 1900
rect 20775 1880 20795 1900
rect 20795 1880 20800 1900
rect 20770 1875 20800 1880
rect 20570 1675 20596 1680
rect 20570 1655 20571 1675
rect 20571 1655 20591 1675
rect 20591 1655 20596 1675
rect 20570 1650 20596 1655
rect 20515 1625 20545 1630
rect 20515 1605 20520 1625
rect 20520 1605 20540 1625
rect 20540 1605 20545 1625
rect 20515 1600 20545 1605
rect 20621 1600 20651 1630
rect 20715 1600 20745 1630
rect 20805 1625 20835 1630
rect 20805 1605 20810 1625
rect 20810 1605 20830 1625
rect 20830 1605 20835 1625
rect 20805 1600 20835 1605
rect 4270 1540 4300 1545
rect 4270 1520 4275 1540
rect 4275 1520 4295 1540
rect 4295 1520 4300 1540
rect 4270 1515 4300 1520
rect 4390 1540 4420 1545
rect 4390 1520 4395 1540
rect 4395 1520 4415 1540
rect 4415 1520 4420 1540
rect 4390 1515 4420 1520
rect 4510 1540 4540 1545
rect 4510 1520 4515 1540
rect 4515 1520 4535 1540
rect 4535 1520 4540 1540
rect 4510 1515 4540 1520
rect 4630 1540 4660 1545
rect 4630 1520 4635 1540
rect 4635 1520 4655 1540
rect 4655 1520 4660 1540
rect 4630 1515 4660 1520
rect 4750 1540 4780 1545
rect 4750 1520 4755 1540
rect 4755 1520 4775 1540
rect 4775 1520 4780 1540
rect 4750 1515 4780 1520
rect 5140 1515 5170 1545
rect 12820 1540 12850 1570
rect 20320 1540 20350 1570
rect 20475 1565 20501 1570
rect 20475 1545 20476 1565
rect 20476 1545 20496 1565
rect 20496 1545 20501 1565
rect 20475 1540 20501 1545
rect 20849 1565 20875 1570
rect 20849 1545 20854 1565
rect 20854 1545 20874 1565
rect 20874 1545 20875 1565
rect 20849 1540 20875 1545
rect 4210 1495 4240 1500
rect 4210 1475 4215 1495
rect 4215 1475 4235 1495
rect 4235 1475 4240 1495
rect 4210 1470 4240 1475
rect 4330 1495 4360 1500
rect 4330 1475 4335 1495
rect 4335 1475 4355 1495
rect 4355 1475 4360 1495
rect 4330 1470 4360 1475
rect 4450 1495 4480 1500
rect 4450 1475 4455 1495
rect 4455 1475 4475 1495
rect 4475 1475 4480 1495
rect 4450 1470 4480 1475
rect 4690 1495 4720 1500
rect 4690 1475 4695 1495
rect 4695 1475 4715 1495
rect 4715 1475 4720 1495
rect 4690 1470 4720 1475
rect 4810 1495 4840 1500
rect 4810 1475 4815 1495
rect 4815 1475 4835 1495
rect 4835 1475 4840 1495
rect 4810 1470 4840 1475
rect 4930 1495 4960 1500
rect 4930 1475 4935 1495
rect 4935 1475 4955 1495
rect 4955 1475 4960 1495
rect 4930 1470 4960 1475
rect 5050 1495 5080 1500
rect 5050 1475 5055 1495
rect 5055 1475 5075 1495
rect 5075 1475 5080 1495
rect 5050 1470 5080 1475
rect 11109 1490 11135 1495
rect 11109 1470 11112 1490
rect 11112 1470 11129 1490
rect 11129 1470 11135 1490
rect 11109 1465 11135 1470
rect 11310 1490 11340 1495
rect 11310 1470 11315 1490
rect 11315 1470 11335 1490
rect 11335 1470 11340 1490
rect 11310 1465 11340 1470
rect 11530 1490 11560 1495
rect 11530 1470 11535 1490
rect 11535 1470 11555 1490
rect 11555 1470 11560 1490
rect 11530 1465 11560 1470
rect 11925 1490 11951 1495
rect 11925 1470 11928 1490
rect 11928 1470 11945 1490
rect 11945 1470 11951 1490
rect 11925 1465 11951 1470
rect 12149 1490 12175 1495
rect 12149 1470 12152 1490
rect 12152 1470 12169 1490
rect 12169 1470 12175 1490
rect 12149 1465 12175 1470
rect 12350 1490 12380 1495
rect 12350 1470 12355 1490
rect 12355 1470 12375 1490
rect 12375 1470 12380 1490
rect 12350 1465 12380 1470
rect 12570 1490 12600 1495
rect 12570 1470 12575 1490
rect 12575 1470 12595 1490
rect 12595 1470 12600 1490
rect 12570 1465 12600 1470
rect 18609 1490 18635 1495
rect 18609 1470 18612 1490
rect 18612 1470 18629 1490
rect 18629 1470 18635 1490
rect 18609 1465 18635 1470
rect 18810 1490 18840 1495
rect 18810 1470 18815 1490
rect 18815 1470 18835 1490
rect 18835 1470 18840 1490
rect 18810 1465 18840 1470
rect 19030 1490 19060 1495
rect 19030 1470 19035 1490
rect 19035 1470 19055 1490
rect 19055 1470 19060 1490
rect 19030 1465 19060 1470
rect 19425 1490 19451 1495
rect 19425 1470 19428 1490
rect 19428 1470 19445 1490
rect 19445 1470 19451 1490
rect 19425 1465 19451 1470
rect 19649 1490 19675 1495
rect 19649 1470 19652 1490
rect 19652 1470 19669 1490
rect 19669 1470 19675 1490
rect 19649 1465 19675 1470
rect 19850 1490 19880 1495
rect 19850 1470 19855 1490
rect 19855 1470 19875 1490
rect 19875 1470 19880 1490
rect 19850 1465 19880 1470
rect 20070 1490 20100 1495
rect 20070 1470 20075 1490
rect 20075 1470 20095 1490
rect 20095 1470 20100 1490
rect 20070 1465 20100 1470
rect 11150 1430 11180 1435
rect 11150 1410 11155 1430
rect 11155 1410 11175 1430
rect 11175 1410 11180 1430
rect 11150 1405 11180 1410
rect 11255 1430 11285 1435
rect 11255 1410 11260 1430
rect 11260 1410 11280 1430
rect 11280 1410 11285 1430
rect 11255 1405 11285 1410
rect 11365 1430 11395 1435
rect 11365 1410 11370 1430
rect 11370 1410 11390 1430
rect 11390 1410 11395 1430
rect 11365 1405 11395 1410
rect 11475 1430 11505 1435
rect 11475 1410 11480 1430
rect 11480 1410 11500 1430
rect 11500 1410 11505 1430
rect 11475 1405 11505 1410
rect 11585 1430 11615 1435
rect 11585 1410 11590 1430
rect 11590 1410 11610 1430
rect 11610 1410 11615 1430
rect 11585 1405 11615 1410
rect 11815 1305 11845 1335
rect 11320 1255 11350 1285
rect 12190 1430 12220 1435
rect 12190 1410 12195 1430
rect 12195 1410 12215 1430
rect 12215 1410 12220 1430
rect 12190 1405 12220 1410
rect 12295 1430 12325 1435
rect 12295 1410 12300 1430
rect 12300 1410 12320 1430
rect 12320 1410 12325 1430
rect 12295 1405 12325 1410
rect 12405 1430 12435 1435
rect 12405 1410 12410 1430
rect 12410 1410 12430 1430
rect 12430 1410 12435 1430
rect 12405 1405 12435 1410
rect 12515 1430 12545 1435
rect 12515 1410 12520 1430
rect 12520 1410 12540 1430
rect 12540 1410 12545 1430
rect 12515 1405 12545 1410
rect 12625 1430 12655 1435
rect 12625 1410 12630 1430
rect 12630 1410 12650 1430
rect 12650 1410 12655 1430
rect 12625 1405 12655 1410
rect 13020 1425 13055 1430
rect 13020 1400 13025 1425
rect 13025 1400 13050 1425
rect 13050 1400 13055 1425
rect 13020 1395 13055 1400
rect 14030 1425 14065 1430
rect 14030 1400 14035 1425
rect 14035 1400 14060 1425
rect 14060 1400 14065 1425
rect 14030 1395 14065 1400
rect 18650 1430 18680 1435
rect 18650 1410 18655 1430
rect 18655 1410 18675 1430
rect 18675 1410 18680 1430
rect 18650 1405 18680 1410
rect 18755 1430 18785 1435
rect 18755 1410 18760 1430
rect 18760 1410 18780 1430
rect 18780 1410 18785 1430
rect 18755 1405 18785 1410
rect 18865 1430 18895 1435
rect 18865 1410 18870 1430
rect 18870 1410 18890 1430
rect 18890 1410 18895 1430
rect 18865 1405 18895 1410
rect 18975 1430 19005 1435
rect 18975 1410 18980 1430
rect 18980 1410 19000 1430
rect 19000 1410 19005 1430
rect 18975 1405 19005 1410
rect 19085 1430 19115 1435
rect 19085 1410 19090 1430
rect 19090 1410 19110 1430
rect 19110 1410 19115 1430
rect 19085 1405 19115 1410
rect 13025 1345 13055 1375
rect 13130 1345 13160 1375
rect 19315 1355 19345 1385
rect 13030 1315 13060 1320
rect 13030 1295 13035 1315
rect 13035 1295 13055 1315
rect 13055 1295 13060 1315
rect 13030 1290 13060 1295
rect 13230 1315 13260 1320
rect 13230 1295 13235 1315
rect 13235 1295 13255 1315
rect 13255 1295 13260 1315
rect 13230 1290 13260 1295
rect 13430 1315 13460 1320
rect 13430 1295 13435 1315
rect 13435 1295 13455 1315
rect 13455 1295 13460 1315
rect 13430 1290 13460 1295
rect 13630 1315 13660 1320
rect 13630 1295 13635 1315
rect 13635 1295 13655 1315
rect 13655 1295 13660 1315
rect 13630 1290 13660 1295
rect 13830 1315 13860 1320
rect 13830 1295 13835 1315
rect 13835 1295 13855 1315
rect 13855 1295 13860 1315
rect 13830 1290 13860 1295
rect 14030 1315 14060 1320
rect 14030 1295 14035 1315
rect 14035 1295 14055 1315
rect 14055 1295 14060 1315
rect 14030 1290 14060 1295
rect 18820 1305 18850 1335
rect 11885 1255 11915 1285
rect 19690 1430 19720 1435
rect 19690 1410 19695 1430
rect 19695 1410 19715 1430
rect 19715 1410 19720 1430
rect 19690 1405 19720 1410
rect 19795 1430 19825 1435
rect 19795 1410 19800 1430
rect 19800 1410 19820 1430
rect 19820 1410 19825 1430
rect 19795 1405 19825 1410
rect 19905 1430 19935 1435
rect 19905 1410 19910 1430
rect 19910 1410 19930 1430
rect 19930 1410 19935 1430
rect 19905 1405 19935 1410
rect 20015 1430 20045 1435
rect 20015 1410 20020 1430
rect 20020 1410 20040 1430
rect 20040 1410 20045 1430
rect 20015 1405 20045 1410
rect 20125 1430 20155 1435
rect 20125 1410 20130 1430
rect 20130 1410 20150 1430
rect 20150 1410 20155 1430
rect 20125 1405 20155 1410
rect 19385 1305 19415 1335
rect 20528 1345 20554 1350
rect 20528 1325 20533 1345
rect 20533 1325 20553 1345
rect 20553 1325 20554 1345
rect 20528 1320 20554 1325
rect 20796 1345 20822 1350
rect 20796 1325 20797 1345
rect 20797 1325 20817 1345
rect 20817 1325 20822 1345
rect 20796 1320 20822 1325
rect 18930 1270 18960 1275
rect 18930 1250 18935 1270
rect 18935 1250 18955 1270
rect 18955 1250 18960 1270
rect 18930 1245 18960 1250
rect 19040 1270 19070 1275
rect 19040 1250 19045 1270
rect 19045 1250 19065 1270
rect 19065 1250 19070 1270
rect 19040 1245 19070 1250
rect 19150 1270 19180 1275
rect 19150 1250 19155 1270
rect 19155 1250 19175 1270
rect 19175 1250 19180 1270
rect 19150 1245 19180 1250
rect 19260 1270 19290 1275
rect 19260 1250 19265 1270
rect 19265 1250 19285 1270
rect 19285 1250 19290 1270
rect 19260 1245 19290 1250
rect 19370 1270 19400 1275
rect 19370 1250 19375 1270
rect 19375 1250 19395 1270
rect 19395 1250 19400 1270
rect 19370 1245 19400 1250
rect 19480 1270 19510 1275
rect 19480 1250 19485 1270
rect 19485 1250 19505 1270
rect 19505 1250 19510 1270
rect 19480 1245 19510 1250
rect 19590 1270 19620 1275
rect 19590 1250 19595 1270
rect 19595 1250 19615 1270
rect 19615 1250 19620 1270
rect 19590 1245 19620 1250
rect 19700 1270 19730 1275
rect 19700 1250 19705 1270
rect 19705 1250 19725 1270
rect 19725 1250 19730 1270
rect 19700 1245 19730 1250
rect 19810 1270 19840 1275
rect 19810 1250 19815 1270
rect 19815 1250 19835 1270
rect 19835 1250 19840 1270
rect 19810 1245 19840 1250
rect 19920 1270 19950 1275
rect 19920 1250 19925 1270
rect 19925 1250 19945 1270
rect 19945 1250 19950 1270
rect 19920 1245 19950 1250
rect 20030 1270 20060 1275
rect 20030 1250 20035 1270
rect 20035 1250 20055 1270
rect 20055 1250 20060 1270
rect 20030 1245 20060 1250
rect 20100 1285 20130 1290
rect 20100 1265 20105 1285
rect 20105 1265 20125 1285
rect 20125 1265 20130 1285
rect 20100 1260 20130 1265
rect 20450 1285 20480 1290
rect 20450 1265 20455 1285
rect 20455 1265 20475 1285
rect 20475 1265 20480 1285
rect 20450 1260 20480 1265
rect 20565 1285 20595 1290
rect 20565 1265 20570 1285
rect 20570 1265 20590 1285
rect 20590 1265 20595 1285
rect 20565 1260 20595 1265
rect 20660 1260 20690 1290
rect 20755 1285 20785 1290
rect 20755 1265 20760 1285
rect 20760 1265 20780 1285
rect 20780 1265 20785 1285
rect 20755 1260 20785 1265
rect 20870 1285 20900 1290
rect 20870 1265 20875 1285
rect 20875 1265 20895 1285
rect 20895 1265 20900 1285
rect 20870 1260 20900 1265
rect 11430 1220 11460 1225
rect 11430 1200 11435 1220
rect 11435 1200 11455 1220
rect 11455 1200 11460 1220
rect 11430 1195 11460 1200
rect 11540 1220 11570 1225
rect 11540 1200 11545 1220
rect 11545 1200 11565 1220
rect 11565 1200 11570 1220
rect 11540 1195 11570 1200
rect 11650 1220 11680 1225
rect 11650 1200 11655 1220
rect 11655 1200 11675 1220
rect 11675 1200 11680 1220
rect 11650 1195 11680 1200
rect 11760 1220 11790 1225
rect 11760 1200 11765 1220
rect 11765 1200 11785 1220
rect 11785 1200 11790 1220
rect 11760 1195 11790 1200
rect 11870 1220 11900 1225
rect 11870 1200 11875 1220
rect 11875 1200 11895 1220
rect 11895 1200 11900 1220
rect 11870 1195 11900 1200
rect 11980 1220 12010 1225
rect 11980 1200 11985 1220
rect 11985 1200 12005 1220
rect 12005 1200 12010 1220
rect 11980 1195 12010 1200
rect 12090 1220 12120 1225
rect 12090 1200 12095 1220
rect 12095 1200 12115 1220
rect 12115 1200 12120 1220
rect 12090 1195 12120 1200
rect 12200 1220 12230 1225
rect 12200 1200 12205 1220
rect 12205 1200 12225 1220
rect 12225 1200 12230 1220
rect 12200 1195 12230 1200
rect 12310 1220 12340 1225
rect 12310 1200 12315 1220
rect 12315 1200 12335 1220
rect 12335 1200 12340 1220
rect 12310 1195 12340 1200
rect 12420 1220 12450 1225
rect 12420 1200 12425 1220
rect 12425 1200 12445 1220
rect 12445 1200 12450 1220
rect 12420 1195 12450 1200
rect 12530 1220 12560 1225
rect 12530 1200 12535 1220
rect 12535 1200 12555 1220
rect 12555 1200 12560 1220
rect 12530 1195 12560 1200
rect 12600 1235 12630 1240
rect 12600 1215 12605 1235
rect 12605 1215 12625 1235
rect 12625 1215 12630 1235
rect 12600 1210 12630 1215
rect 20605 1225 20635 1230
rect 20605 1205 20610 1225
rect 20610 1205 20630 1225
rect 20630 1205 20635 1225
rect 20605 1200 20635 1205
rect 20660 1225 20690 1230
rect 20660 1205 20665 1225
rect 20665 1205 20685 1225
rect 20685 1205 20690 1225
rect 20660 1200 20690 1205
rect 20715 1225 20745 1230
rect 20715 1205 20720 1225
rect 20720 1205 20740 1225
rect 20740 1205 20745 1225
rect 20715 1200 20745 1205
rect 20870 1200 20900 1230
rect 3380 1180 3410 1185
rect 3380 1160 3385 1180
rect 3385 1160 3405 1180
rect 3405 1160 3410 1180
rect 3380 1155 3410 1160
rect 3990 1155 4020 1185
rect 4600 1180 4630 1185
rect 4600 1160 4605 1180
rect 4605 1160 4625 1180
rect 4625 1160 4630 1180
rect 4600 1155 4630 1160
rect 2950 1120 2980 1125
rect 2950 1100 2955 1120
rect 2955 1100 2975 1120
rect 2975 1100 2980 1120
rect 2950 1095 2980 1100
rect 3030 1120 3060 1125
rect 3030 1100 3035 1120
rect 3035 1100 3055 1120
rect 3055 1100 3060 1120
rect 3030 1095 3060 1100
rect 3110 1120 3140 1125
rect 3110 1100 3115 1120
rect 3115 1100 3135 1120
rect 3135 1100 3140 1120
rect 3110 1095 3140 1100
rect 3190 1120 3220 1125
rect 3190 1100 3195 1120
rect 3195 1100 3215 1120
rect 3215 1100 3220 1120
rect 3190 1095 3220 1100
rect 3270 1120 3300 1125
rect 3270 1100 3275 1120
rect 3275 1100 3295 1120
rect 3295 1100 3300 1120
rect 3270 1095 3300 1100
rect 3350 1120 3380 1125
rect 3350 1100 3355 1120
rect 3355 1100 3375 1120
rect 3375 1100 3380 1120
rect 3350 1095 3380 1100
rect 3430 1120 3460 1125
rect 3430 1100 3435 1120
rect 3435 1100 3455 1120
rect 3455 1100 3460 1120
rect 3430 1095 3460 1100
rect 3510 1120 3540 1125
rect 3510 1100 3515 1120
rect 3515 1100 3535 1120
rect 3535 1100 3540 1120
rect 3510 1095 3540 1100
rect 3590 1120 3620 1125
rect 3590 1100 3595 1120
rect 3595 1100 3615 1120
rect 3615 1100 3620 1120
rect 3590 1095 3620 1100
rect 3670 1120 3700 1125
rect 3670 1100 3675 1120
rect 3675 1100 3695 1120
rect 3695 1100 3700 1120
rect 3670 1095 3700 1100
rect 3750 1120 3780 1125
rect 3750 1100 3755 1120
rect 3755 1100 3775 1120
rect 3775 1100 3780 1120
rect 3750 1095 3780 1100
rect 3830 1120 3860 1125
rect 3830 1100 3835 1120
rect 3835 1100 3855 1120
rect 3855 1100 3860 1120
rect 3830 1095 3860 1100
rect 3910 1120 3940 1125
rect 3910 1100 3915 1120
rect 3915 1100 3935 1120
rect 3935 1100 3940 1120
rect 3910 1095 3940 1100
rect 3990 1120 4020 1125
rect 3990 1100 3995 1120
rect 3995 1100 4015 1120
rect 4015 1100 4020 1120
rect 3990 1095 4020 1100
rect 4070 1120 4100 1125
rect 4070 1100 4075 1120
rect 4075 1100 4095 1120
rect 4095 1100 4100 1120
rect 4070 1095 4100 1100
rect 4150 1120 4180 1125
rect 4150 1100 4155 1120
rect 4155 1100 4175 1120
rect 4175 1100 4180 1120
rect 4150 1095 4180 1100
rect 4230 1120 4260 1125
rect 4230 1100 4235 1120
rect 4235 1100 4255 1120
rect 4255 1100 4260 1120
rect 4230 1095 4260 1100
rect 4310 1120 4340 1125
rect 4310 1100 4315 1120
rect 4315 1100 4335 1120
rect 4335 1100 4340 1120
rect 4310 1095 4340 1100
rect 4390 1120 4420 1125
rect 4390 1100 4395 1120
rect 4395 1100 4415 1120
rect 4415 1100 4420 1120
rect 4390 1095 4420 1100
rect 4470 1120 4500 1125
rect 4470 1100 4475 1120
rect 4475 1100 4495 1120
rect 4495 1100 4500 1120
rect 4470 1095 4500 1100
rect 4550 1120 4580 1125
rect 4550 1100 4555 1120
rect 4555 1100 4575 1120
rect 4575 1100 4580 1120
rect 4550 1095 4580 1100
rect 4630 1120 4660 1125
rect 4630 1100 4635 1120
rect 4635 1100 4655 1120
rect 4655 1100 4660 1120
rect 4630 1095 4660 1100
rect 4710 1120 4740 1125
rect 4710 1100 4715 1120
rect 4715 1100 4735 1120
rect 4735 1100 4740 1120
rect 4710 1095 4740 1100
rect 4790 1120 4820 1125
rect 4790 1100 4795 1120
rect 4795 1100 4815 1120
rect 4815 1100 4820 1120
rect 4790 1095 4820 1100
rect 4870 1120 4900 1125
rect 4870 1100 4875 1120
rect 4875 1100 4895 1120
rect 4895 1100 4900 1120
rect 4870 1095 4900 1100
rect 4950 1120 4980 1125
rect 4950 1100 4955 1120
rect 4955 1100 4975 1120
rect 4975 1100 4980 1120
rect 4950 1095 4980 1100
rect 2625 1010 2655 1040
rect 2910 1035 2940 1040
rect 2910 1015 2915 1035
rect 2915 1015 2935 1035
rect 2935 1015 2940 1035
rect 2910 1010 2940 1015
rect 5115 1035 5145 1040
rect 5115 1015 5120 1035
rect 5120 1015 5140 1035
rect 5140 1015 5145 1035
rect 5115 1010 5145 1015
rect 13130 965 13160 970
rect 13130 945 13135 965
rect 13135 945 13155 965
rect 13155 945 13160 965
rect 13130 940 13160 945
rect 13330 965 13360 970
rect 13330 945 13335 965
rect 13335 945 13355 965
rect 13355 945 13360 965
rect 13330 940 13360 945
rect 13530 965 13560 970
rect 13530 945 13535 965
rect 13535 945 13555 965
rect 13555 945 13560 965
rect 13530 940 13560 945
rect 13730 965 13760 970
rect 13730 945 13735 965
rect 13735 945 13755 965
rect 13755 945 13760 965
rect 13730 940 13760 945
rect 13930 965 13960 970
rect 13930 945 13935 965
rect 13935 945 13955 965
rect 13955 945 13960 965
rect 13930 940 13960 945
rect 3000 925 3030 930
rect 3000 905 3005 925
rect 3005 905 3025 925
rect 3025 905 3030 925
rect 3000 900 3030 905
rect 3180 925 3210 930
rect 3180 905 3185 925
rect 3185 905 3205 925
rect 3205 905 3210 925
rect 3180 900 3210 905
rect 3360 925 3390 930
rect 3360 905 3365 925
rect 3365 905 3385 925
rect 3385 905 3390 925
rect 3360 900 3390 905
rect 3540 925 3570 930
rect 3540 905 3545 925
rect 3545 905 3565 925
rect 3565 905 3570 925
rect 3540 900 3570 905
rect 3720 925 3750 930
rect 3720 905 3725 925
rect 3725 905 3745 925
rect 3745 905 3750 925
rect 3720 900 3750 905
rect 3900 925 3930 930
rect 3900 905 3905 925
rect 3905 905 3925 925
rect 3925 905 3930 925
rect 3900 900 3930 905
rect 4080 925 4110 930
rect 4080 905 4085 925
rect 4085 905 4105 925
rect 4105 905 4110 925
rect 4080 900 4110 905
rect 4260 925 4290 930
rect 4260 905 4265 925
rect 4265 905 4285 925
rect 4285 905 4290 925
rect 4260 900 4290 905
rect 4440 925 4470 930
rect 4440 905 4445 925
rect 4445 905 4465 925
rect 4465 905 4470 925
rect 4440 900 4470 905
rect 4620 925 4650 930
rect 4620 905 4625 925
rect 4625 905 4645 925
rect 4645 905 4650 925
rect 4620 900 4650 905
rect 4800 925 4830 930
rect 4800 905 4805 925
rect 4805 905 4825 925
rect 4825 905 4830 925
rect 4800 900 4830 905
rect 4980 925 5010 930
rect 4980 905 4985 925
rect 4985 905 5005 925
rect 5005 905 5010 925
rect 4980 900 5010 905
rect 18670 950 18700 955
rect 18670 930 18675 950
rect 18675 930 18695 950
rect 18695 930 18700 950
rect 18670 925 18700 930
rect 18765 950 18795 955
rect 18765 930 18770 950
rect 18770 930 18790 950
rect 18790 930 18795 950
rect 18765 925 18795 930
rect 18875 950 18905 955
rect 18875 930 18880 950
rect 18880 930 18900 950
rect 18900 930 18905 950
rect 18875 925 18905 930
rect 18985 950 19015 955
rect 18985 930 18990 950
rect 18990 930 19010 950
rect 19010 930 19015 950
rect 18985 925 19015 930
rect 19095 950 19125 955
rect 19095 930 19100 950
rect 19100 930 19120 950
rect 19120 930 19125 950
rect 19095 925 19125 930
rect 19205 950 19235 955
rect 19205 930 19210 950
rect 19210 930 19230 950
rect 19230 930 19235 950
rect 19205 925 19235 930
rect 19315 950 19345 955
rect 19315 930 19320 950
rect 19320 930 19340 950
rect 19340 930 19345 950
rect 19315 925 19345 930
rect 19425 950 19455 955
rect 19425 930 19430 950
rect 19430 930 19450 950
rect 19450 930 19455 950
rect 19425 925 19455 930
rect 19535 950 19565 955
rect 19535 930 19540 950
rect 19540 930 19560 950
rect 19560 930 19565 950
rect 19535 925 19565 930
rect 19645 950 19675 955
rect 19645 930 19650 950
rect 19650 930 19670 950
rect 19670 930 19675 950
rect 19645 925 19675 930
rect 19755 950 19785 955
rect 19755 930 19760 950
rect 19760 930 19780 950
rect 19780 930 19785 950
rect 19755 925 19785 930
rect 19865 950 19895 955
rect 19865 930 19870 950
rect 19870 930 19890 950
rect 19890 930 19895 950
rect 19865 925 19895 930
rect 19975 950 20005 955
rect 19975 930 19980 950
rect 19980 930 20000 950
rect 20000 930 20005 950
rect 19975 925 20005 930
rect 20125 950 20155 955
rect 20125 930 20130 950
rect 20130 930 20150 950
rect 20150 930 20155 950
rect 20125 925 20155 930
rect 11170 900 11200 905
rect 11170 880 11175 900
rect 11175 880 11195 900
rect 11195 880 11200 900
rect 11170 875 11200 880
rect 11265 900 11295 905
rect 11265 880 11270 900
rect 11270 880 11290 900
rect 11290 880 11295 900
rect 11265 875 11295 880
rect 11375 900 11405 905
rect 11375 880 11380 900
rect 11380 880 11400 900
rect 11400 880 11405 900
rect 11375 875 11405 880
rect 11485 900 11515 905
rect 11485 880 11490 900
rect 11490 880 11510 900
rect 11510 880 11515 900
rect 11485 875 11515 880
rect 11595 900 11625 905
rect 11595 880 11600 900
rect 11600 880 11620 900
rect 11620 880 11625 900
rect 11595 875 11625 880
rect 11705 900 11735 905
rect 11705 880 11710 900
rect 11710 880 11730 900
rect 11730 880 11735 900
rect 11705 875 11735 880
rect 11815 900 11845 905
rect 11815 880 11820 900
rect 11820 880 11840 900
rect 11840 880 11845 900
rect 11815 875 11845 880
rect 11925 900 11955 905
rect 11925 880 11930 900
rect 11930 880 11950 900
rect 11950 880 11955 900
rect 11925 875 11955 880
rect 12035 900 12065 905
rect 12035 880 12040 900
rect 12040 880 12060 900
rect 12060 880 12065 900
rect 12035 875 12065 880
rect 12145 900 12175 905
rect 12145 880 12150 900
rect 12150 880 12170 900
rect 12170 880 12175 900
rect 12145 875 12175 880
rect 12255 900 12285 905
rect 12255 880 12260 900
rect 12260 880 12280 900
rect 12280 880 12285 900
rect 12255 875 12285 880
rect 12365 900 12395 905
rect 12365 880 12370 900
rect 12370 880 12390 900
rect 12390 880 12395 900
rect 12365 875 12395 880
rect 12475 900 12505 905
rect 12475 880 12480 900
rect 12480 880 12500 900
rect 12500 880 12505 900
rect 12475 875 12505 880
rect 12625 900 12655 905
rect 12625 880 12630 900
rect 12630 880 12650 900
rect 12650 880 12655 900
rect 12625 875 12655 880
rect 2525 730 2555 760
rect 3135 755 3165 760
rect 3135 735 3140 755
rect 3140 735 3160 755
rect 3160 735 3165 755
rect 3135 730 3165 735
rect 3630 755 3660 760
rect 3630 735 3635 755
rect 3635 735 3655 755
rect 3655 735 3660 755
rect 3630 730 3660 735
rect 3990 755 4020 760
rect 3990 735 3995 755
rect 3995 735 4015 755
rect 4015 735 4020 755
rect 3990 730 4020 735
rect 4350 755 4380 760
rect 4350 735 4355 755
rect 4355 735 4375 755
rect 4375 735 4380 755
rect 4350 730 4380 735
rect 4530 755 4560 760
rect 4530 735 4535 755
rect 4535 735 4555 755
rect 4555 735 4560 755
rect 4530 730 4560 735
rect 4710 755 4740 760
rect 4710 735 4715 755
rect 4715 735 4735 755
rect 4735 735 4740 755
rect 4710 730 4740 735
rect 4890 755 4920 760
rect 4890 735 4895 755
rect 4895 735 4915 755
rect 4915 735 4920 755
rect 4890 730 4920 735
rect 3450 675 3480 705
rect 3810 675 3840 705
rect 4170 675 4200 705
rect 9380 -685 9410 -680
rect 9380 -705 9385 -685
rect 9385 -705 9405 -685
rect 9405 -705 9410 -685
rect 9380 -710 9410 -705
rect 9580 -685 9610 -680
rect 9580 -705 9585 -685
rect 9585 -705 9605 -685
rect 9605 -705 9610 -685
rect 9580 -710 9610 -705
rect 9780 -685 9810 -680
rect 9780 -705 9785 -685
rect 9785 -705 9805 -685
rect 9805 -705 9810 -685
rect 9780 -710 9810 -705
rect 9980 -685 10010 -680
rect 9980 -705 9985 -685
rect 9985 -705 10005 -685
rect 10005 -705 10010 -685
rect 9980 -710 10010 -705
rect 10180 -685 10210 -680
rect 10180 -705 10185 -685
rect 10185 -705 10205 -685
rect 10205 -705 10210 -685
rect 10180 -710 10210 -705
rect 10380 -685 10410 -680
rect 10380 -705 10385 -685
rect 10385 -705 10405 -685
rect 10405 -705 10410 -685
rect 10380 -710 10410 -705
rect 9480 -1035 9510 -1030
rect 9480 -1055 9485 -1035
rect 9485 -1055 9505 -1035
rect 9505 -1055 9510 -1035
rect 9480 -1060 9510 -1055
rect 9680 -1035 9710 -1030
rect 9680 -1055 9685 -1035
rect 9685 -1055 9705 -1035
rect 9705 -1055 9710 -1035
rect 9680 -1060 9710 -1055
rect 9880 -1035 9910 -1030
rect 9880 -1055 9885 -1035
rect 9885 -1055 9905 -1035
rect 9905 -1055 9910 -1035
rect 9880 -1060 9910 -1055
rect 10080 -1035 10110 -1030
rect 10080 -1055 10085 -1035
rect 10085 -1055 10105 -1035
rect 10105 -1055 10110 -1035
rect 10080 -1060 10110 -1055
rect 10280 -1035 10310 -1030
rect 10280 -1055 10285 -1035
rect 10285 -1055 10305 -1035
rect 10305 -1055 10310 -1035
rect 10280 -1060 10310 -1055
<< metal2 >>
rect -195 4990 -155 4995
rect -195 4960 -190 4990
rect -160 4960 -155 4990
rect -195 4955 -155 4960
rect 5550 4990 5590 4995
rect 5550 4960 5555 4990
rect 5585 4960 5590 4990
rect 5550 4955 5590 4960
rect 11340 3625 11380 3630
rect 11340 3595 11345 3625
rect 11375 3620 11380 3625
rect 11460 3625 11500 3630
rect 11460 3620 11465 3625
rect 11375 3600 11465 3620
rect 11375 3595 11380 3600
rect 11340 3590 11380 3595
rect 11460 3595 11465 3600
rect 11495 3620 11500 3625
rect 11580 3625 11620 3630
rect 11580 3620 11585 3625
rect 11495 3600 11585 3620
rect 11495 3595 11500 3600
rect 11460 3590 11500 3595
rect 11580 3595 11585 3600
rect 11615 3620 11620 3625
rect 11700 3625 11740 3630
rect 11700 3620 11705 3625
rect 11615 3600 11705 3620
rect 11615 3595 11620 3600
rect 11580 3590 11620 3595
rect 11700 3595 11705 3600
rect 11735 3620 11740 3625
rect 11820 3625 11860 3630
rect 11820 3620 11825 3625
rect 11735 3600 11825 3620
rect 11735 3595 11740 3600
rect 11700 3590 11740 3595
rect 11820 3595 11825 3600
rect 11855 3620 11860 3625
rect 11940 3625 11980 3630
rect 11940 3620 11945 3625
rect 11855 3600 11945 3620
rect 11855 3595 11860 3600
rect 11820 3590 11860 3595
rect 11940 3595 11945 3600
rect 11975 3620 11980 3625
rect 12060 3625 12100 3630
rect 12060 3620 12065 3625
rect 11975 3600 12065 3620
rect 11975 3595 11980 3600
rect 11940 3590 11980 3595
rect 12060 3595 12065 3600
rect 12095 3620 12100 3625
rect 12180 3625 12220 3630
rect 12180 3620 12185 3625
rect 12095 3600 12185 3620
rect 12095 3595 12100 3600
rect 12060 3590 12100 3595
rect 12180 3595 12185 3600
rect 12215 3620 12220 3625
rect 12300 3625 12340 3630
rect 12300 3620 12305 3625
rect 12215 3600 12305 3620
rect 12215 3595 12220 3600
rect 12180 3590 12220 3595
rect 12300 3595 12305 3600
rect 12335 3620 12340 3625
rect 12420 3625 12460 3630
rect 12420 3620 12425 3625
rect 12335 3600 12425 3620
rect 12335 3595 12340 3600
rect 12300 3590 12340 3595
rect 12420 3595 12425 3600
rect 12455 3595 12460 3625
rect 12420 3590 12460 3595
rect 18840 3625 18880 3630
rect 18840 3595 18845 3625
rect 18875 3620 18880 3625
rect 18960 3625 19000 3630
rect 18960 3620 18965 3625
rect 18875 3600 18965 3620
rect 18875 3595 18880 3600
rect 18840 3590 18880 3595
rect 18960 3595 18965 3600
rect 18995 3620 19000 3625
rect 19080 3625 19120 3630
rect 19080 3620 19085 3625
rect 18995 3600 19085 3620
rect 18995 3595 19000 3600
rect 18960 3590 19000 3595
rect 19080 3595 19085 3600
rect 19115 3620 19120 3625
rect 19200 3625 19240 3630
rect 19200 3620 19205 3625
rect 19115 3600 19205 3620
rect 19115 3595 19120 3600
rect 19080 3590 19120 3595
rect 19200 3595 19205 3600
rect 19235 3620 19240 3625
rect 19320 3625 19360 3630
rect 19320 3620 19325 3625
rect 19235 3600 19325 3620
rect 19235 3595 19240 3600
rect 19200 3590 19240 3595
rect 19320 3595 19325 3600
rect 19355 3620 19360 3625
rect 19440 3625 19480 3630
rect 19440 3620 19445 3625
rect 19355 3600 19445 3620
rect 19355 3595 19360 3600
rect 19320 3590 19360 3595
rect 19440 3595 19445 3600
rect 19475 3620 19480 3625
rect 19560 3625 19600 3630
rect 19560 3620 19565 3625
rect 19475 3600 19565 3620
rect 19475 3595 19480 3600
rect 19440 3590 19480 3595
rect 19560 3595 19565 3600
rect 19595 3620 19600 3625
rect 19680 3625 19720 3630
rect 19680 3620 19685 3625
rect 19595 3600 19685 3620
rect 19595 3595 19600 3600
rect 19560 3590 19600 3595
rect 19680 3595 19685 3600
rect 19715 3620 19720 3625
rect 19800 3625 19840 3630
rect 19800 3620 19805 3625
rect 19715 3600 19805 3620
rect 19715 3595 19720 3600
rect 19680 3590 19720 3595
rect 19800 3595 19805 3600
rect 19835 3620 19840 3625
rect 19920 3625 19960 3630
rect 19920 3620 19925 3625
rect 19835 3600 19925 3620
rect 19835 3595 19840 3600
rect 19800 3590 19840 3595
rect 19920 3595 19925 3600
rect 19955 3595 19960 3625
rect 19920 3590 19960 3595
rect -110 3525 -70 3530
rect -110 3495 -105 3525
rect -75 3520 -70 3525
rect 1261 3525 1301 3530
rect 1261 3520 1266 3525
rect -75 3500 1266 3520
rect -75 3495 -70 3500
rect -110 3490 -70 3495
rect 1261 3495 1266 3500
rect 1296 3495 1301 3525
rect 1261 3490 1301 3495
rect 4440 3495 4480 3500
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect -15 3445 25 3450
rect -15 3415 -10 3445
rect 20 3440 25 3445
rect 940 3445 980 3450
rect 940 3440 945 3445
rect 20 3420 945 3440
rect 20 3415 25 3420
rect -15 3410 25 3415
rect 940 3415 945 3420
rect 975 3415 980 3445
rect 940 3410 980 3415
rect 1635 3445 1685 3455
rect 2470 3450 2510 3455
rect 2470 3445 2475 3450
rect 1635 3415 1645 3445
rect 1675 3425 2475 3445
rect 1675 3415 1685 3425
rect 2470 3420 2475 3425
rect 2505 3420 2510 3450
rect 2470 3415 2510 3420
rect 5135 3445 5185 3455
rect 5135 3415 5145 3445
rect 5175 3440 5185 3445
rect 5550 3445 5590 3450
rect 5550 3440 5555 3445
rect 5175 3420 5555 3440
rect 5175 3415 5185 3420
rect 1635 3405 1685 3415
rect 5135 3405 5185 3415
rect 5550 3415 5555 3420
rect 5585 3415 5590 3445
rect 5550 3410 5590 3415
rect -60 3390 -20 3395
rect -60 3360 -55 3390
rect -25 3385 -20 3390
rect 2690 3390 2730 3395
rect 2690 3385 2695 3390
rect -25 3365 2695 3385
rect -25 3360 -20 3365
rect -60 3355 -20 3360
rect 2690 3360 2695 3365
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 1205 3340 1245 3345
rect 1205 3310 1210 3340
rect 1240 3335 1245 3340
rect 3135 3340 3175 3345
rect 3135 3335 3140 3340
rect 1240 3315 3140 3335
rect 1240 3310 1245 3315
rect 1205 3305 1245 3310
rect 3135 3310 3140 3315
rect 3170 3310 3175 3340
rect 3135 3305 3175 3310
rect 3385 3335 3435 3345
rect 3385 3305 3395 3335
rect 3425 3330 3435 3335
rect 5360 3335 5400 3340
rect 5360 3330 5365 3335
rect 3425 3310 5365 3330
rect 3425 3305 3435 3310
rect 3385 3295 3435 3305
rect 5360 3305 5365 3310
rect 5395 3305 5400 3335
rect 5360 3300 5400 3305
rect 12945 3290 12985 3295
rect 1160 3285 1200 3290
rect 1160 3255 1165 3285
rect 1195 3280 1200 3285
rect 4885 3285 4925 3290
rect 4885 3280 4890 3285
rect 1195 3260 4890 3280
rect 1195 3255 1200 3260
rect 1160 3250 1200 3255
rect 4885 3255 4890 3260
rect 4920 3280 4925 3285
rect 5410 3285 5450 3290
rect 5410 3280 5415 3285
rect 4920 3260 5415 3280
rect 4920 3255 4925 3260
rect 4885 3250 4925 3255
rect 5410 3255 5415 3260
rect 5445 3255 5450 3285
rect 12945 3260 12950 3290
rect 12980 3285 12985 3290
rect 13055 3290 13095 3295
rect 13055 3285 13060 3290
rect 12980 3265 13060 3285
rect 12980 3260 12985 3265
rect 12945 3255 12985 3260
rect 13055 3260 13060 3265
rect 13090 3285 13095 3290
rect 13165 3290 13205 3295
rect 13165 3285 13170 3290
rect 13090 3265 13170 3285
rect 13090 3260 13095 3265
rect 13055 3255 13095 3260
rect 13165 3260 13170 3265
rect 13200 3285 13205 3290
rect 13275 3290 13315 3295
rect 13275 3285 13280 3290
rect 13200 3265 13280 3285
rect 13200 3260 13205 3265
rect 13165 3255 13205 3260
rect 13275 3260 13280 3265
rect 13310 3285 13315 3290
rect 13385 3290 13425 3295
rect 13385 3285 13390 3290
rect 13310 3265 13390 3285
rect 13310 3260 13315 3265
rect 13275 3255 13315 3260
rect 13385 3260 13390 3265
rect 13420 3285 13425 3290
rect 13495 3290 13535 3295
rect 13495 3285 13500 3290
rect 13420 3265 13500 3285
rect 13420 3260 13425 3265
rect 13385 3255 13425 3260
rect 13495 3260 13500 3265
rect 13530 3285 13535 3290
rect 13605 3290 13645 3295
rect 13605 3285 13610 3290
rect 13530 3265 13610 3285
rect 13530 3260 13535 3265
rect 13495 3255 13535 3260
rect 13605 3260 13610 3265
rect 13640 3285 13645 3290
rect 13715 3290 13755 3295
rect 13715 3285 13720 3290
rect 13640 3265 13720 3285
rect 13640 3260 13645 3265
rect 13605 3255 13645 3260
rect 13715 3260 13720 3265
rect 13750 3285 13755 3290
rect 13825 3290 13865 3295
rect 13825 3285 13830 3290
rect 13750 3265 13830 3285
rect 13750 3260 13755 3265
rect 13715 3255 13755 3260
rect 13825 3260 13830 3265
rect 13860 3285 13865 3290
rect 13935 3290 13975 3295
rect 13935 3285 13940 3290
rect 13860 3265 13940 3285
rect 13860 3260 13865 3265
rect 13825 3255 13865 3260
rect 13935 3260 13940 3265
rect 13970 3285 13975 3290
rect 14045 3290 14085 3295
rect 14045 3285 14050 3290
rect 13970 3265 14050 3285
rect 13970 3260 13975 3265
rect 13935 3255 13975 3260
rect 14045 3260 14050 3265
rect 14080 3260 14085 3290
rect 14045 3255 14085 3260
rect 20445 3290 20485 3295
rect 20445 3260 20450 3290
rect 20480 3285 20485 3290
rect 20555 3290 20595 3295
rect 20555 3285 20560 3290
rect 20480 3265 20560 3285
rect 20480 3260 20485 3265
rect 20445 3255 20485 3260
rect 20555 3260 20560 3265
rect 20590 3285 20595 3290
rect 20665 3290 20705 3295
rect 20665 3285 20670 3290
rect 20590 3265 20670 3285
rect 20590 3260 20595 3265
rect 20555 3255 20595 3260
rect 20665 3260 20670 3265
rect 20700 3285 20705 3290
rect 20775 3290 20815 3295
rect 20775 3285 20780 3290
rect 20700 3265 20780 3285
rect 20700 3260 20705 3265
rect 20665 3255 20705 3260
rect 20775 3260 20780 3265
rect 20810 3285 20815 3290
rect 20885 3290 20925 3295
rect 20885 3285 20890 3290
rect 20810 3265 20890 3285
rect 20810 3260 20815 3265
rect 20775 3255 20815 3260
rect 20885 3260 20890 3265
rect 20920 3285 20925 3290
rect 20995 3290 21035 3295
rect 20995 3285 21000 3290
rect 20920 3265 21000 3285
rect 20920 3260 20925 3265
rect 20885 3255 20925 3260
rect 20995 3260 21000 3265
rect 21030 3285 21035 3290
rect 21105 3290 21145 3295
rect 21105 3285 21110 3290
rect 21030 3265 21110 3285
rect 21030 3260 21035 3265
rect 20995 3255 21035 3260
rect 21105 3260 21110 3265
rect 21140 3285 21145 3290
rect 21215 3290 21255 3295
rect 21215 3285 21220 3290
rect 21140 3265 21220 3285
rect 21140 3260 21145 3265
rect 21105 3255 21145 3260
rect 21215 3260 21220 3265
rect 21250 3285 21255 3290
rect 21325 3290 21365 3295
rect 21325 3285 21330 3290
rect 21250 3265 21330 3285
rect 21250 3260 21255 3265
rect 21215 3255 21255 3260
rect 21325 3260 21330 3265
rect 21360 3285 21365 3290
rect 21435 3290 21475 3295
rect 21435 3285 21440 3290
rect 21360 3265 21440 3285
rect 21360 3260 21365 3265
rect 21325 3255 21365 3260
rect 21435 3260 21440 3265
rect 21470 3285 21475 3290
rect 21545 3290 21585 3295
rect 21545 3285 21550 3290
rect 21470 3265 21550 3285
rect 21470 3260 21475 3265
rect 21435 3255 21475 3260
rect 21545 3260 21550 3265
rect 21580 3260 21585 3290
rect 21545 3255 21585 3260
rect 5410 3250 5450 3255
rect 2735 3240 2775 3245
rect 2735 3235 2740 3240
rect 46 3215 2740 3235
rect 46 3205 91 3215
rect 2735 3210 2740 3215
rect 2770 3210 2775 3240
rect 2735 3205 2775 3210
rect 10580 3210 10620 3215
rect 46 3170 51 3205
rect 86 3170 91 3205
rect 1261 3165 1266 3200
rect 1301 3165 1306 3200
rect 2620 3185 2660 3190
rect 2620 3155 2625 3185
rect 2655 3180 2660 3185
rect 4440 3185 4480 3190
rect 4440 3180 4445 3185
rect 2655 3160 4445 3180
rect 2655 3155 2660 3160
rect 2620 3150 2660 3155
rect 4440 3155 4445 3160
rect 4475 3155 4480 3185
rect 10580 3180 10585 3210
rect 10615 3205 10620 3210
rect 10980 3210 11015 3215
rect 10980 3205 10985 3210
rect 10615 3185 10985 3205
rect 10615 3180 10620 3185
rect 10580 3175 10620 3180
rect 10980 3180 10985 3185
rect 10980 3175 11015 3180
rect 18080 3210 18120 3215
rect 18080 3180 18085 3210
rect 18115 3205 18120 3210
rect 18480 3210 18515 3215
rect 18480 3205 18485 3210
rect 18115 3185 18485 3205
rect 18115 3180 18120 3185
rect 18080 3175 18120 3180
rect 18480 3180 18485 3185
rect 18480 3175 18515 3180
rect 4440 3150 4480 3155
rect 10900 3155 10940 3160
rect -110 3140 -70 3145
rect -110 3110 -105 3140
rect -75 3135 -70 3140
rect 46 3135 51 3145
rect -75 3115 51 3135
rect -75 3110 -70 3115
rect 46 3110 51 3115
rect 86 3110 91 3145
rect 3135 3140 3175 3145
rect -110 3105 -70 3110
rect 1261 3105 1266 3140
rect 1301 3105 1306 3140
rect 3135 3110 3140 3140
rect 3170 3135 3175 3140
rect 4835 3140 4875 3145
rect 4835 3135 4840 3140
rect 3170 3115 4840 3135
rect 3170 3110 3175 3115
rect 3135 3105 3175 3110
rect 4835 3110 4840 3115
rect 4870 3135 4875 3140
rect 5315 3140 5355 3145
rect 5315 3135 5320 3140
rect 4870 3115 5320 3135
rect 4870 3110 4875 3115
rect 4835 3105 4875 3110
rect 5315 3110 5320 3115
rect 5350 3110 5355 3140
rect 10900 3125 10905 3155
rect 10935 3150 10940 3155
rect 11823 3155 11857 3160
rect 11823 3150 11826 3155
rect 10935 3130 11826 3150
rect 10935 3125 10940 3130
rect 10900 3120 10940 3125
rect 11823 3125 11826 3130
rect 11854 3125 11857 3155
rect 11823 3120 11857 3125
rect 18400 3155 18440 3160
rect 18400 3125 18405 3155
rect 18435 3150 18440 3155
rect 19323 3155 19357 3160
rect 19323 3150 19326 3155
rect 18435 3130 19326 3150
rect 18435 3125 18440 3130
rect 18400 3120 18440 3125
rect 19323 3125 19326 3130
rect 19354 3125 19357 3155
rect 19323 3120 19357 3125
rect 5315 3105 5355 3110
rect 1160 3100 1200 3105
rect 1160 3095 1165 3100
rect 46 3075 1165 3095
rect 46 3065 91 3075
rect 1160 3070 1165 3075
rect 1195 3070 1200 3100
rect 11280 3100 11320 3105
rect 1160 3065 1200 3070
rect 3985 3080 4025 3085
rect 46 3030 51 3065
rect 86 3030 91 3065
rect 3985 3050 3990 3080
rect 4020 3075 4025 3080
rect 4020 3055 6100 3075
rect 11280 3070 11285 3100
rect 11315 3095 11320 3100
rect 11520 3100 11560 3105
rect 11520 3095 11525 3100
rect 11315 3075 11525 3095
rect 11315 3070 11320 3075
rect 11280 3065 11320 3070
rect 11520 3070 11525 3075
rect 11555 3095 11560 3100
rect 11760 3100 11800 3105
rect 11760 3095 11765 3100
rect 11555 3075 11765 3095
rect 11555 3070 11560 3075
rect 11520 3065 11560 3070
rect 11760 3070 11765 3075
rect 11795 3095 11800 3100
rect 12000 3100 12040 3105
rect 12000 3095 12005 3100
rect 11795 3075 12005 3095
rect 11795 3070 11800 3075
rect 11760 3065 11800 3070
rect 12000 3070 12005 3075
rect 12035 3095 12040 3100
rect 12240 3100 12280 3105
rect 12240 3095 12245 3100
rect 12035 3075 12245 3095
rect 12035 3070 12040 3075
rect 12000 3065 12040 3070
rect 12240 3070 12245 3075
rect 12275 3095 12280 3100
rect 12480 3100 12520 3105
rect 12480 3095 12485 3100
rect 12275 3075 12485 3095
rect 12275 3070 12280 3075
rect 12240 3065 12280 3070
rect 12480 3070 12485 3075
rect 12515 3070 12520 3100
rect 12480 3065 12520 3070
rect 18780 3100 18820 3105
rect 18780 3070 18785 3100
rect 18815 3095 18820 3100
rect 19020 3100 19060 3105
rect 19020 3095 19025 3100
rect 18815 3075 19025 3095
rect 18815 3070 18820 3075
rect 18780 3065 18820 3070
rect 19020 3070 19025 3075
rect 19055 3095 19060 3100
rect 19260 3100 19300 3105
rect 19260 3095 19265 3100
rect 19055 3075 19265 3095
rect 19055 3070 19060 3075
rect 19020 3065 19060 3070
rect 19260 3070 19265 3075
rect 19295 3095 19300 3100
rect 19500 3100 19540 3105
rect 19500 3095 19505 3100
rect 19295 3075 19505 3095
rect 19295 3070 19300 3075
rect 19260 3065 19300 3070
rect 19500 3070 19505 3075
rect 19535 3095 19540 3100
rect 19740 3100 19780 3105
rect 19740 3095 19745 3100
rect 19535 3075 19745 3095
rect 19535 3070 19540 3075
rect 19500 3065 19540 3070
rect 19740 3070 19745 3075
rect 19775 3095 19780 3100
rect 19980 3100 20020 3105
rect 19980 3095 19985 3100
rect 19775 3075 19985 3095
rect 19775 3070 19780 3075
rect 19740 3065 19780 3070
rect 19980 3070 19985 3075
rect 20015 3070 20020 3100
rect 19980 3065 20020 3070
rect 11400 3055 11440 3060
rect 4020 3050 4025 3055
rect 3985 3045 4025 3050
rect 3445 3035 3485 3040
rect 3445 3005 3450 3035
rect 3480 3030 3485 3035
rect 3805 3035 3845 3040
rect 3805 3030 3810 3035
rect 3480 3010 3810 3030
rect 3480 3005 3485 3010
rect -110 3000 -70 3005
rect -110 2970 -105 3000
rect -75 2995 -70 3000
rect 46 2995 51 3005
rect -75 2975 51 2995
rect -75 2970 -70 2975
rect 46 2970 51 2975
rect 86 2970 91 3005
rect 3445 3000 3485 3005
rect 3805 3005 3810 3010
rect 3840 3030 3845 3035
rect 4345 3035 4385 3040
rect 4345 3030 4350 3035
rect 3840 3010 4350 3030
rect 3840 3005 3845 3010
rect 3805 3000 3845 3005
rect 4345 3005 4350 3010
rect 4380 3030 4385 3035
rect 4705 3035 4745 3040
rect 4705 3030 4710 3035
rect 4380 3010 4710 3030
rect 4380 3005 4385 3010
rect 4345 3000 4385 3005
rect 4705 3005 4710 3010
rect 4740 3030 4745 3035
rect 4740 3010 6100 3030
rect 11400 3025 11405 3055
rect 11435 3050 11440 3055
rect 11640 3055 11680 3060
rect 11640 3050 11645 3055
rect 11435 3030 11645 3050
rect 11435 3025 11440 3030
rect 11400 3020 11440 3025
rect 11640 3025 11645 3030
rect 11675 3050 11680 3055
rect 11880 3055 11920 3060
rect 11880 3050 11885 3055
rect 11675 3030 11885 3050
rect 11675 3025 11680 3030
rect 11640 3020 11680 3025
rect 11880 3025 11885 3030
rect 11915 3050 11920 3055
rect 12120 3055 12160 3060
rect 12120 3050 12125 3055
rect 11915 3030 12125 3050
rect 11915 3025 11920 3030
rect 11880 3020 11920 3025
rect 12120 3025 12125 3030
rect 12155 3050 12160 3055
rect 12360 3055 12400 3060
rect 12360 3050 12365 3055
rect 12155 3030 12365 3050
rect 12155 3025 12160 3030
rect 12120 3020 12160 3025
rect 12360 3025 12365 3030
rect 12395 3025 12400 3055
rect 12360 3020 12400 3025
rect 18900 3055 18940 3060
rect 18900 3025 18905 3055
rect 18935 3050 18940 3055
rect 19140 3055 19180 3060
rect 19140 3050 19145 3055
rect 18935 3030 19145 3050
rect 18935 3025 18940 3030
rect 18900 3020 18940 3025
rect 19140 3025 19145 3030
rect 19175 3050 19180 3055
rect 19380 3055 19420 3060
rect 19380 3050 19385 3055
rect 19175 3030 19385 3050
rect 19175 3025 19180 3030
rect 19140 3020 19180 3025
rect 19380 3025 19385 3030
rect 19415 3050 19420 3055
rect 19620 3055 19660 3060
rect 19620 3050 19625 3055
rect 19415 3030 19625 3050
rect 19415 3025 19420 3030
rect 19380 3020 19420 3025
rect 19620 3025 19625 3030
rect 19655 3050 19660 3055
rect 19860 3055 19900 3060
rect 19860 3050 19865 3055
rect 19655 3030 19865 3050
rect 19655 3025 19660 3030
rect 19620 3020 19660 3025
rect 19860 3025 19865 3030
rect 19895 3025 19900 3055
rect 19860 3020 19900 3025
rect 4740 3005 4745 3010
rect 4705 3000 4745 3005
rect 11340 3000 11380 3005
rect 2520 2980 2560 2985
rect -110 2965 -70 2970
rect 2330 2925 2335 2960
rect 2370 2950 2375 2960
rect 2425 2955 2465 2960
rect 2425 2950 2430 2955
rect 2370 2930 2430 2950
rect 2370 2925 2375 2930
rect 2425 2925 2430 2930
rect 2460 2925 2465 2955
rect 2520 2950 2525 2980
rect 2555 2975 2560 2980
rect 3080 2980 3120 2985
rect 3080 2975 3085 2980
rect 2555 2955 3085 2975
rect 2555 2950 2560 2955
rect 2520 2945 2560 2950
rect 3080 2950 3085 2955
rect 3115 2950 3120 2980
rect 3080 2945 3120 2950
rect 3265 2980 3305 2985
rect 3265 2950 3270 2980
rect 3300 2975 3305 2980
rect 3625 2980 3665 2985
rect 3625 2975 3630 2980
rect 3300 2955 3630 2975
rect 3300 2950 3305 2955
rect 3265 2945 3305 2950
rect 3625 2950 3630 2955
rect 3660 2975 3665 2980
rect 4165 2980 4205 2985
rect 4165 2975 4170 2980
rect 3660 2955 4170 2975
rect 3660 2950 3665 2955
rect 3625 2945 3665 2950
rect 4165 2950 4170 2955
rect 4200 2975 4205 2980
rect 4525 2980 4565 2985
rect 4525 2975 4530 2980
rect 4200 2955 4530 2975
rect 4200 2950 4205 2955
rect 4165 2945 4205 2950
rect 4525 2950 4530 2955
rect 4560 2975 4565 2980
rect 4560 2955 6100 2975
rect 11340 2970 11345 3000
rect 11375 2995 11380 3000
rect 11400 3000 11440 3005
rect 11400 2995 11405 3000
rect 11375 2975 11405 2995
rect 11375 2970 11380 2975
rect 11340 2965 11380 2970
rect 11400 2970 11405 2975
rect 11435 2995 11440 3000
rect 11580 3000 11620 3005
rect 11580 2995 11585 3000
rect 11435 2975 11585 2995
rect 11435 2970 11440 2975
rect 11400 2965 11440 2970
rect 11580 2970 11585 2975
rect 11615 2995 11620 3000
rect 11820 3000 11860 3005
rect 11820 2995 11825 3000
rect 11615 2975 11825 2995
rect 11615 2970 11620 2975
rect 11580 2965 11620 2970
rect 11820 2970 11825 2975
rect 11855 2995 11860 3000
rect 12060 3000 12100 3005
rect 12060 2995 12065 3000
rect 11855 2975 12065 2995
rect 11855 2970 11860 2975
rect 11820 2965 11860 2970
rect 12060 2970 12065 2975
rect 12095 2995 12100 3000
rect 12300 3000 12340 3005
rect 12300 2995 12305 3000
rect 12095 2975 12305 2995
rect 12095 2970 12100 2975
rect 12060 2965 12100 2970
rect 12300 2970 12305 2975
rect 12335 2970 12340 3000
rect 12300 2965 12340 2970
rect 18840 3000 18880 3005
rect 18840 2970 18845 3000
rect 18875 2995 18880 3000
rect 18900 3000 18940 3005
rect 18900 2995 18905 3000
rect 18875 2975 18905 2995
rect 18875 2970 18880 2975
rect 18840 2965 18880 2970
rect 18900 2970 18905 2975
rect 18935 2995 18940 3000
rect 19080 3000 19120 3005
rect 19080 2995 19085 3000
rect 18935 2975 19085 2995
rect 18935 2970 18940 2975
rect 18900 2965 18940 2970
rect 19080 2970 19085 2975
rect 19115 2995 19120 3000
rect 19320 3000 19360 3005
rect 19320 2995 19325 3000
rect 19115 2975 19325 2995
rect 19115 2970 19120 2975
rect 19080 2965 19120 2970
rect 19320 2970 19325 2975
rect 19355 2995 19360 3000
rect 19560 3000 19600 3005
rect 19560 2995 19565 3000
rect 19355 2975 19565 2995
rect 19355 2970 19360 2975
rect 19320 2965 19360 2970
rect 19560 2970 19565 2975
rect 19595 2995 19600 3000
rect 19800 3000 19840 3005
rect 19800 2995 19805 3000
rect 19595 2975 19805 2995
rect 19595 2970 19600 2975
rect 19560 2965 19600 2970
rect 19800 2970 19805 2975
rect 19835 2970 19840 3000
rect 19800 2965 19840 2970
rect 4560 2950 4565 2955
rect 4525 2945 4565 2950
rect 11460 2945 11500 2950
rect 2425 2920 2465 2925
rect -110 2910 -70 2915
rect -110 2880 -105 2910
rect -75 2905 -70 2910
rect 905 2910 1125 2920
rect 11460 2915 11465 2945
rect 11495 2940 11500 2945
rect 11700 2945 11740 2950
rect 11700 2940 11705 2945
rect 11495 2920 11705 2940
rect 11495 2915 11500 2920
rect 11460 2910 11500 2915
rect 11700 2915 11705 2920
rect 11735 2940 11740 2945
rect 11940 2945 11980 2950
rect 11940 2940 11945 2945
rect 11735 2920 11945 2940
rect 11735 2915 11740 2920
rect 11700 2910 11740 2915
rect 11940 2915 11945 2920
rect 11975 2940 11980 2945
rect 12180 2945 12220 2950
rect 12180 2940 12185 2945
rect 11975 2920 12185 2940
rect 11975 2915 11980 2920
rect 11940 2910 11980 2915
rect 12180 2915 12185 2920
rect 12215 2940 12220 2945
rect 12420 2945 12460 2950
rect 12420 2940 12425 2945
rect 12215 2920 12425 2940
rect 12215 2915 12220 2920
rect 12180 2910 12220 2915
rect 12420 2915 12425 2920
rect 12455 2940 12460 2945
rect 12480 2945 12520 2950
rect 12480 2940 12485 2945
rect 12455 2920 12485 2940
rect 12455 2915 12460 2920
rect 12420 2910 12460 2915
rect 12480 2915 12485 2920
rect 12515 2915 12520 2945
rect 18960 2945 19000 2950
rect 12480 2910 12520 2915
rect 13000 2920 13040 2925
rect 905 2905 920 2910
rect -75 2885 920 2905
rect -75 2880 -70 2885
rect -110 2875 -70 2880
rect 905 2880 920 2885
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1125 2910
rect 905 2870 1125 2880
rect 2330 2900 2375 2905
rect 2330 2865 2335 2900
rect 2370 2865 2375 2900
rect 13000 2890 13005 2920
rect 13035 2915 13040 2920
rect 13110 2920 13150 2925
rect 13110 2915 13115 2920
rect 13035 2895 13115 2915
rect 13035 2890 13040 2895
rect 13000 2885 13040 2890
rect 13110 2890 13115 2895
rect 13145 2915 13150 2920
rect 13220 2920 13260 2925
rect 13220 2915 13225 2920
rect 13145 2895 13225 2915
rect 13145 2890 13150 2895
rect 13110 2885 13150 2890
rect 13220 2890 13225 2895
rect 13255 2915 13260 2920
rect 13330 2920 13370 2925
rect 13330 2915 13335 2920
rect 13255 2895 13335 2915
rect 13255 2890 13260 2895
rect 13220 2885 13260 2890
rect 13330 2890 13335 2895
rect 13365 2915 13370 2920
rect 13440 2920 13480 2925
rect 13440 2915 13445 2920
rect 13365 2895 13445 2915
rect 13365 2890 13370 2895
rect 13330 2885 13370 2890
rect 13440 2890 13445 2895
rect 13475 2915 13480 2920
rect 13550 2920 13590 2925
rect 13550 2915 13555 2920
rect 13475 2895 13555 2915
rect 13475 2890 13480 2895
rect 13440 2885 13480 2890
rect 13550 2890 13555 2895
rect 13585 2915 13590 2920
rect 13660 2920 13700 2925
rect 13660 2915 13665 2920
rect 13585 2895 13665 2915
rect 13585 2890 13590 2895
rect 13550 2885 13590 2890
rect 13660 2890 13665 2895
rect 13695 2915 13700 2920
rect 13770 2920 13810 2925
rect 13770 2915 13775 2920
rect 13695 2895 13775 2915
rect 13695 2890 13700 2895
rect 13660 2885 13700 2890
rect 13770 2890 13775 2895
rect 13805 2915 13810 2920
rect 13880 2920 13920 2925
rect 13880 2915 13885 2920
rect 13805 2895 13885 2915
rect 13805 2890 13810 2895
rect 13770 2885 13810 2890
rect 13880 2890 13885 2895
rect 13915 2915 13920 2920
rect 13990 2920 14030 2925
rect 13990 2915 13995 2920
rect 13915 2895 13995 2915
rect 13915 2890 13920 2895
rect 13880 2885 13920 2890
rect 13990 2890 13995 2895
rect 14025 2890 14030 2920
rect 18960 2915 18965 2945
rect 18995 2940 19000 2945
rect 19200 2945 19240 2950
rect 19200 2940 19205 2945
rect 18995 2920 19205 2940
rect 18995 2915 19000 2920
rect 18960 2910 19000 2915
rect 19200 2915 19205 2920
rect 19235 2940 19240 2945
rect 19440 2945 19480 2950
rect 19440 2940 19445 2945
rect 19235 2920 19445 2940
rect 19235 2915 19240 2920
rect 19200 2910 19240 2915
rect 19440 2915 19445 2920
rect 19475 2940 19480 2945
rect 19680 2945 19720 2950
rect 19680 2940 19685 2945
rect 19475 2920 19685 2940
rect 19475 2915 19480 2920
rect 19440 2910 19480 2915
rect 19680 2915 19685 2920
rect 19715 2940 19720 2945
rect 19920 2945 19960 2950
rect 19920 2940 19925 2945
rect 19715 2920 19925 2940
rect 19715 2915 19720 2920
rect 19680 2910 19720 2915
rect 19920 2915 19925 2920
rect 19955 2940 19960 2945
rect 19980 2945 20020 2950
rect 19980 2940 19985 2945
rect 19955 2920 19985 2940
rect 19955 2915 19960 2920
rect 19920 2910 19960 2915
rect 19980 2915 19985 2920
rect 20015 2915 20020 2945
rect 19980 2910 20020 2915
rect 20500 2920 20540 2925
rect 13990 2885 14030 2890
rect 20500 2890 20505 2920
rect 20535 2915 20540 2920
rect 20610 2920 20650 2925
rect 20610 2915 20615 2920
rect 20535 2895 20615 2915
rect 20535 2890 20540 2895
rect 20500 2885 20540 2890
rect 20610 2890 20615 2895
rect 20645 2915 20650 2920
rect 20720 2920 20760 2925
rect 20720 2915 20725 2920
rect 20645 2895 20725 2915
rect 20645 2890 20650 2895
rect 20610 2885 20650 2890
rect 20720 2890 20725 2895
rect 20755 2915 20760 2920
rect 20830 2920 20870 2925
rect 20830 2915 20835 2920
rect 20755 2895 20835 2915
rect 20755 2890 20760 2895
rect 20720 2885 20760 2890
rect 20830 2890 20835 2895
rect 20865 2915 20870 2920
rect 20940 2920 20980 2925
rect 20940 2915 20945 2920
rect 20865 2895 20945 2915
rect 20865 2890 20870 2895
rect 20830 2885 20870 2890
rect 20940 2890 20945 2895
rect 20975 2915 20980 2920
rect 21050 2920 21090 2925
rect 21050 2915 21055 2920
rect 20975 2895 21055 2915
rect 20975 2890 20980 2895
rect 20940 2885 20980 2890
rect 21050 2890 21055 2895
rect 21085 2915 21090 2920
rect 21160 2920 21200 2925
rect 21160 2915 21165 2920
rect 21085 2895 21165 2915
rect 21085 2890 21090 2895
rect 21050 2885 21090 2890
rect 21160 2890 21165 2895
rect 21195 2915 21200 2920
rect 21270 2920 21310 2925
rect 21270 2915 21275 2920
rect 21195 2895 21275 2915
rect 21195 2890 21200 2895
rect 21160 2885 21200 2890
rect 21270 2890 21275 2895
rect 21305 2915 21310 2920
rect 21380 2920 21420 2925
rect 21380 2915 21385 2920
rect 21305 2895 21385 2915
rect 21305 2890 21310 2895
rect 21270 2885 21310 2890
rect 21380 2890 21385 2895
rect 21415 2915 21420 2920
rect 21490 2920 21530 2925
rect 21490 2915 21495 2920
rect 21415 2895 21495 2915
rect 21415 2890 21420 2895
rect 21380 2885 21420 2890
rect 21490 2890 21495 2895
rect 21525 2890 21530 2920
rect 21490 2885 21530 2890
rect 2330 2860 2375 2865
rect -60 2855 -20 2860
rect -60 2825 -55 2855
rect -25 2850 -20 2855
rect 51 2850 56 2855
rect -25 2830 56 2850
rect -25 2825 -20 2830
rect -60 2820 -20 2825
rect 51 2820 56 2830
rect 91 2820 96 2855
rect 724 2820 729 2855
rect 764 2845 769 2855
rect 1205 2850 1245 2855
rect 1205 2845 1210 2850
rect 764 2825 1210 2845
rect 764 2820 769 2825
rect 1205 2820 1210 2825
rect 1240 2820 1245 2850
rect 1205 2815 1245 2820
rect 1261 2805 1266 2840
rect 1301 2805 1306 2840
rect 1960 2805 1965 2840
rect 2000 2830 2005 2840
rect 2330 2835 2370 2840
rect 2330 2830 2335 2835
rect 2000 2810 2335 2830
rect 2000 2805 2005 2810
rect 2330 2805 2335 2810
rect 2365 2805 2370 2835
rect 13055 2830 13095 2836
rect 2330 2800 2370 2805
rect 2995 2810 3035 2815
rect -15 2795 25 2800
rect -15 2765 -10 2795
rect 20 2785 25 2795
rect 51 2785 56 2795
rect 20 2765 56 2785
rect -15 2760 25 2765
rect 51 2760 56 2765
rect 91 2760 96 2795
rect 724 2760 729 2795
rect 764 2785 769 2795
rect 2620 2790 2660 2795
rect 2620 2785 2625 2790
rect 764 2765 2625 2785
rect 764 2760 769 2765
rect 2620 2760 2625 2765
rect 2655 2760 2660 2790
rect 2995 2780 3000 2810
rect 3030 2805 3035 2810
rect 3175 2810 3215 2815
rect 3175 2805 3180 2810
rect 3030 2785 3180 2805
rect 3030 2780 3035 2785
rect 2995 2775 3035 2780
rect 3175 2780 3180 2785
rect 3210 2805 3215 2810
rect 3355 2810 3395 2815
rect 3355 2805 3360 2810
rect 3210 2785 3360 2805
rect 3210 2780 3215 2785
rect 3175 2775 3215 2780
rect 3355 2780 3360 2785
rect 3390 2805 3395 2810
rect 3535 2810 3575 2815
rect 3535 2805 3540 2810
rect 3390 2785 3540 2805
rect 3390 2780 3395 2785
rect 3355 2775 3395 2780
rect 3535 2780 3540 2785
rect 3570 2805 3575 2810
rect 3715 2810 3755 2815
rect 3715 2805 3720 2810
rect 3570 2785 3720 2805
rect 3570 2780 3575 2785
rect 3535 2775 3575 2780
rect 3715 2780 3720 2785
rect 3750 2805 3755 2810
rect 3895 2810 3935 2815
rect 3895 2805 3900 2810
rect 3750 2785 3900 2805
rect 3750 2780 3755 2785
rect 3715 2775 3755 2780
rect 3895 2780 3900 2785
rect 3930 2805 3935 2810
rect 4075 2810 4115 2815
rect 4075 2805 4080 2810
rect 3930 2785 4080 2805
rect 3930 2780 3935 2785
rect 3895 2775 3935 2780
rect 4075 2780 4080 2785
rect 4110 2805 4115 2810
rect 4255 2810 4295 2815
rect 4255 2805 4260 2810
rect 4110 2785 4260 2805
rect 4110 2780 4115 2785
rect 4075 2775 4115 2780
rect 4255 2780 4260 2785
rect 4290 2805 4295 2810
rect 4435 2810 4475 2815
rect 4435 2805 4440 2810
rect 4290 2785 4440 2805
rect 4290 2780 4295 2785
rect 4255 2775 4295 2780
rect 4435 2780 4440 2785
rect 4470 2805 4475 2810
rect 4615 2810 4655 2815
rect 4615 2805 4620 2810
rect 4470 2785 4620 2805
rect 4470 2780 4475 2785
rect 4435 2775 4475 2780
rect 4615 2780 4620 2785
rect 4650 2805 4655 2810
rect 4795 2810 4835 2815
rect 4795 2805 4800 2810
rect 4650 2785 4800 2805
rect 4650 2780 4655 2785
rect 4615 2775 4655 2780
rect 4795 2780 4800 2785
rect 4830 2805 4835 2810
rect 4975 2810 5015 2815
rect 4975 2805 4980 2810
rect 4830 2785 4980 2805
rect 4830 2780 4835 2785
rect 4795 2775 4835 2780
rect 4975 2780 4980 2785
rect 5010 2805 5015 2810
rect 5550 2810 5590 2815
rect 5550 2805 5555 2810
rect 5010 2785 5555 2805
rect 5010 2780 5015 2785
rect 4975 2775 5015 2780
rect 5550 2780 5555 2785
rect 5585 2780 5590 2810
rect 5550 2775 5590 2780
rect 13055 2800 13060 2830
rect 13090 2800 13095 2830
rect 13055 2780 13095 2800
rect 2620 2755 2660 2760
rect 3175 2750 3215 2755
rect 1261 2745 1301 2750
rect 1261 2715 1266 2745
rect 1296 2740 1301 2745
rect 2150 2745 2190 2750
rect 2150 2740 2155 2745
rect 1296 2720 2155 2740
rect 1296 2715 1301 2720
rect 1261 2710 1301 2715
rect 2150 2715 2155 2720
rect 2185 2715 2190 2745
rect 3175 2720 3180 2750
rect 3210 2745 3215 2750
rect 3355 2750 3395 2755
rect 3355 2745 3360 2750
rect 3210 2725 3360 2745
rect 3210 2720 3215 2725
rect 3175 2715 3215 2720
rect 3355 2720 3360 2725
rect 3390 2745 3395 2750
rect 3535 2750 3575 2755
rect 3535 2745 3540 2750
rect 3390 2725 3540 2745
rect 3390 2720 3395 2725
rect 3355 2715 3395 2720
rect 3535 2720 3540 2725
rect 3570 2745 3575 2750
rect 3715 2750 3755 2755
rect 3715 2745 3720 2750
rect 3570 2725 3720 2745
rect 3570 2720 3575 2725
rect 3535 2715 3575 2720
rect 3715 2720 3720 2725
rect 3750 2745 3755 2750
rect 3895 2750 3935 2755
rect 3895 2745 3900 2750
rect 3750 2725 3900 2745
rect 3750 2720 3755 2725
rect 3715 2715 3755 2720
rect 3895 2720 3900 2725
rect 3930 2745 3935 2750
rect 4075 2750 4115 2755
rect 4075 2745 4080 2750
rect 3930 2725 4080 2745
rect 3930 2720 3935 2725
rect 3895 2715 3935 2720
rect 4075 2720 4080 2725
rect 4110 2745 4115 2750
rect 4255 2750 4295 2755
rect 4255 2745 4260 2750
rect 4110 2725 4260 2745
rect 4110 2720 4115 2725
rect 4075 2715 4115 2720
rect 4255 2720 4260 2725
rect 4290 2745 4295 2750
rect 4435 2750 4475 2755
rect 4435 2745 4440 2750
rect 4290 2725 4440 2745
rect 4290 2720 4295 2725
rect 4255 2715 4295 2720
rect 4435 2720 4440 2725
rect 4470 2745 4475 2750
rect 4615 2750 4655 2755
rect 4615 2745 4620 2750
rect 4470 2725 4620 2745
rect 4470 2720 4475 2725
rect 4435 2715 4475 2720
rect 4615 2720 4620 2725
rect 4650 2745 4655 2750
rect 4795 2750 4835 2755
rect 4795 2745 4800 2750
rect 4650 2725 4800 2745
rect 4650 2720 4655 2725
rect 4615 2715 4655 2720
rect 4795 2720 4800 2725
rect 4830 2720 4835 2750
rect 13055 2750 13060 2780
rect 13090 2750 13095 2780
rect 4795 2715 4835 2720
rect 12690 2730 12730 2735
rect 2150 2710 2190 2715
rect 12690 2700 12695 2730
rect 12725 2725 12730 2730
rect 13055 2730 13095 2750
rect 20555 2830 20595 2836
rect 20555 2800 20560 2830
rect 20590 2800 20595 2830
rect 20555 2780 20595 2800
rect 20555 2750 20560 2780
rect 20590 2750 20595 2780
rect 13055 2725 13060 2730
rect 12725 2705 13060 2725
rect 12725 2700 12730 2705
rect 12690 2695 12730 2700
rect 13055 2700 13060 2705
rect 13090 2700 13095 2730
rect 13055 2695 13095 2700
rect 20190 2730 20230 2735
rect 20190 2700 20195 2730
rect 20225 2725 20230 2730
rect 20555 2730 20595 2750
rect 20555 2725 20560 2730
rect 20225 2705 20560 2725
rect 20225 2700 20230 2705
rect 20190 2695 20230 2700
rect 20555 2700 20560 2705
rect 20590 2700 20595 2730
rect 20555 2695 20595 2700
rect 9735 2670 9775 2675
rect 9735 2640 9740 2670
rect 9770 2665 9775 2670
rect 9845 2670 9885 2675
rect 9845 2665 9850 2670
rect 9770 2645 9850 2665
rect 9770 2640 9775 2645
rect 9735 2635 9775 2640
rect 9845 2640 9850 2645
rect 9880 2665 9885 2670
rect 9955 2670 9995 2675
rect 9955 2665 9960 2670
rect 9880 2645 9960 2665
rect 9880 2640 9885 2645
rect 9845 2635 9885 2640
rect 9955 2640 9960 2645
rect 9990 2665 9995 2670
rect 10065 2670 10105 2675
rect 10065 2665 10070 2670
rect 9990 2645 10070 2665
rect 9990 2640 9995 2645
rect 9955 2635 9995 2640
rect 10065 2640 10070 2645
rect 10100 2665 10105 2670
rect 10175 2670 10215 2675
rect 10175 2665 10180 2670
rect 10100 2645 10180 2665
rect 10100 2640 10105 2645
rect 10065 2635 10105 2640
rect 10175 2640 10180 2645
rect 10210 2665 10215 2670
rect 10285 2670 10325 2675
rect 10285 2665 10290 2670
rect 10210 2645 10290 2665
rect 10210 2640 10215 2645
rect 10175 2635 10215 2640
rect 10285 2640 10290 2645
rect 10320 2665 10325 2670
rect 10395 2670 10435 2675
rect 10395 2665 10400 2670
rect 10320 2645 10400 2665
rect 10320 2640 10325 2645
rect 10285 2635 10325 2640
rect 10395 2640 10400 2645
rect 10430 2665 10435 2670
rect 10505 2670 10545 2675
rect 10505 2665 10510 2670
rect 10430 2645 10510 2665
rect 10430 2640 10435 2645
rect 10395 2635 10435 2640
rect 10505 2640 10510 2645
rect 10540 2665 10545 2670
rect 10615 2670 10655 2675
rect 10615 2665 10620 2670
rect 10540 2645 10620 2665
rect 10540 2640 10545 2645
rect 10505 2635 10545 2640
rect 10615 2640 10620 2645
rect 10650 2665 10655 2670
rect 10725 2670 10765 2675
rect 10725 2665 10730 2670
rect 10650 2645 10730 2665
rect 10650 2640 10655 2645
rect 10615 2635 10655 2640
rect 10725 2640 10730 2645
rect 10760 2665 10765 2670
rect 10835 2670 10875 2675
rect 10835 2665 10840 2670
rect 10760 2645 10840 2665
rect 10760 2640 10765 2645
rect 10725 2635 10765 2640
rect 10835 2640 10840 2645
rect 10870 2640 10875 2670
rect 10835 2635 10875 2640
rect 12945 2670 12985 2675
rect 12945 2640 12950 2670
rect 12980 2665 12985 2670
rect 13055 2670 13095 2675
rect 13055 2665 13060 2670
rect 12980 2645 13060 2665
rect 12980 2640 12985 2645
rect 12945 2635 12985 2640
rect 13055 2640 13060 2645
rect 13090 2665 13095 2670
rect 13165 2670 13205 2675
rect 13165 2665 13170 2670
rect 13090 2645 13170 2665
rect 13090 2640 13095 2645
rect 13055 2635 13095 2640
rect 13165 2640 13170 2645
rect 13200 2665 13205 2670
rect 13275 2670 13315 2675
rect 13275 2665 13280 2670
rect 13200 2645 13280 2665
rect 13200 2640 13205 2645
rect 13165 2635 13205 2640
rect 13275 2640 13280 2645
rect 13310 2665 13315 2670
rect 13385 2670 13425 2675
rect 13385 2665 13390 2670
rect 13310 2645 13390 2665
rect 13310 2640 13315 2645
rect 13275 2635 13315 2640
rect 13385 2640 13390 2645
rect 13420 2665 13425 2670
rect 13495 2670 13535 2675
rect 13495 2665 13500 2670
rect 13420 2645 13500 2665
rect 13420 2640 13425 2645
rect 13385 2635 13425 2640
rect 13495 2640 13500 2645
rect 13530 2665 13535 2670
rect 13605 2670 13645 2675
rect 13605 2665 13610 2670
rect 13530 2645 13610 2665
rect 13530 2640 13535 2645
rect 13495 2635 13535 2640
rect 13605 2640 13610 2645
rect 13640 2665 13645 2670
rect 13715 2670 13755 2675
rect 13715 2665 13720 2670
rect 13640 2645 13720 2665
rect 13640 2640 13645 2645
rect 13605 2635 13645 2640
rect 13715 2640 13720 2645
rect 13750 2665 13755 2670
rect 13825 2670 13865 2675
rect 13825 2665 13830 2670
rect 13750 2645 13830 2665
rect 13750 2640 13755 2645
rect 13715 2635 13755 2640
rect 13825 2640 13830 2645
rect 13860 2665 13865 2670
rect 13935 2670 13975 2675
rect 13935 2665 13940 2670
rect 13860 2645 13940 2665
rect 13860 2640 13865 2645
rect 13825 2635 13865 2640
rect 13935 2640 13940 2645
rect 13970 2665 13975 2670
rect 14045 2670 14085 2675
rect 14045 2665 14050 2670
rect 13970 2645 14050 2665
rect 13970 2640 13975 2645
rect 13935 2635 13975 2640
rect 14045 2640 14050 2645
rect 14080 2640 14085 2670
rect 14045 2635 14085 2640
rect 17235 2670 17275 2675
rect 17235 2640 17240 2670
rect 17270 2665 17275 2670
rect 17345 2670 17385 2675
rect 17345 2665 17350 2670
rect 17270 2645 17350 2665
rect 17270 2640 17275 2645
rect 17235 2635 17275 2640
rect 17345 2640 17350 2645
rect 17380 2665 17385 2670
rect 17455 2670 17495 2675
rect 17455 2665 17460 2670
rect 17380 2645 17460 2665
rect 17380 2640 17385 2645
rect 17345 2635 17385 2640
rect 17455 2640 17460 2645
rect 17490 2665 17495 2670
rect 17565 2670 17605 2675
rect 17565 2665 17570 2670
rect 17490 2645 17570 2665
rect 17490 2640 17495 2645
rect 17455 2635 17495 2640
rect 17565 2640 17570 2645
rect 17600 2665 17605 2670
rect 17675 2670 17715 2675
rect 17675 2665 17680 2670
rect 17600 2645 17680 2665
rect 17600 2640 17605 2645
rect 17565 2635 17605 2640
rect 17675 2640 17680 2645
rect 17710 2665 17715 2670
rect 17785 2670 17825 2675
rect 17785 2665 17790 2670
rect 17710 2645 17790 2665
rect 17710 2640 17715 2645
rect 17675 2635 17715 2640
rect 17785 2640 17790 2645
rect 17820 2665 17825 2670
rect 17895 2670 17935 2675
rect 17895 2665 17900 2670
rect 17820 2645 17900 2665
rect 17820 2640 17825 2645
rect 17785 2635 17825 2640
rect 17895 2640 17900 2645
rect 17930 2665 17935 2670
rect 18005 2670 18045 2675
rect 18005 2665 18010 2670
rect 17930 2645 18010 2665
rect 17930 2640 17935 2645
rect 17895 2635 17935 2640
rect 18005 2640 18010 2645
rect 18040 2665 18045 2670
rect 18115 2670 18155 2675
rect 18115 2665 18120 2670
rect 18040 2645 18120 2665
rect 18040 2640 18045 2645
rect 18005 2635 18045 2640
rect 18115 2640 18120 2645
rect 18150 2665 18155 2670
rect 18225 2670 18265 2675
rect 18225 2665 18230 2670
rect 18150 2645 18230 2665
rect 18150 2640 18155 2645
rect 18115 2635 18155 2640
rect 18225 2640 18230 2645
rect 18260 2665 18265 2670
rect 18335 2670 18375 2675
rect 18335 2665 18340 2670
rect 18260 2645 18340 2665
rect 18260 2640 18265 2645
rect 18225 2635 18265 2640
rect 18335 2640 18340 2645
rect 18370 2640 18375 2670
rect 18335 2635 18375 2640
rect 20445 2670 20485 2675
rect 20445 2640 20450 2670
rect 20480 2665 20485 2670
rect 20555 2670 20595 2675
rect 20555 2665 20560 2670
rect 20480 2645 20560 2665
rect 20480 2640 20485 2645
rect 20445 2635 20485 2640
rect 20555 2640 20560 2645
rect 20590 2665 20595 2670
rect 20665 2670 20705 2675
rect 20665 2665 20670 2670
rect 20590 2645 20670 2665
rect 20590 2640 20595 2645
rect 20555 2635 20595 2640
rect 20665 2640 20670 2645
rect 20700 2665 20705 2670
rect 20775 2670 20815 2675
rect 20775 2665 20780 2670
rect 20700 2645 20780 2665
rect 20700 2640 20705 2645
rect 20665 2635 20705 2640
rect 20775 2640 20780 2645
rect 20810 2665 20815 2670
rect 20885 2670 20925 2675
rect 20885 2665 20890 2670
rect 20810 2645 20890 2665
rect 20810 2640 20815 2645
rect 20775 2635 20815 2640
rect 20885 2640 20890 2645
rect 20920 2665 20925 2670
rect 20995 2670 21035 2675
rect 20995 2665 21000 2670
rect 20920 2645 21000 2665
rect 20920 2640 20925 2645
rect 20885 2635 20925 2640
rect 20995 2640 21000 2645
rect 21030 2665 21035 2670
rect 21105 2670 21145 2675
rect 21105 2665 21110 2670
rect 21030 2645 21110 2665
rect 21030 2640 21035 2645
rect 20995 2635 21035 2640
rect 21105 2640 21110 2645
rect 21140 2665 21145 2670
rect 21215 2670 21255 2675
rect 21215 2665 21220 2670
rect 21140 2645 21220 2665
rect 21140 2640 21145 2645
rect 21105 2635 21145 2640
rect 21215 2640 21220 2645
rect 21250 2665 21255 2670
rect 21325 2670 21365 2675
rect 21325 2665 21330 2670
rect 21250 2645 21330 2665
rect 21250 2640 21255 2645
rect 21215 2635 21255 2640
rect 21325 2640 21330 2645
rect 21360 2665 21365 2670
rect 21435 2670 21475 2675
rect 21435 2665 21440 2670
rect 21360 2645 21440 2665
rect 21360 2640 21365 2645
rect 21325 2635 21365 2640
rect 21435 2640 21440 2645
rect 21470 2665 21475 2670
rect 21545 2670 21585 2675
rect 21545 2665 21550 2670
rect 21470 2645 21550 2665
rect 21470 2640 21475 2645
rect 21435 2635 21475 2640
rect 21545 2640 21550 2645
rect 21580 2640 21585 2670
rect 21545 2635 21585 2640
rect 9790 2500 9830 2505
rect 9790 2470 9795 2500
rect 9825 2495 9830 2500
rect 9900 2500 9940 2505
rect 9900 2495 9905 2500
rect 9825 2475 9905 2495
rect 9825 2470 9830 2475
rect 9790 2465 9830 2470
rect 9900 2470 9905 2475
rect 9935 2495 9940 2500
rect 10010 2500 10050 2505
rect 10010 2495 10015 2500
rect 9935 2475 10015 2495
rect 9935 2470 9940 2475
rect 9900 2465 9940 2470
rect 10010 2470 10015 2475
rect 10045 2495 10050 2500
rect 10120 2500 10160 2505
rect 10120 2495 10125 2500
rect 10045 2475 10125 2495
rect 10045 2470 10050 2475
rect 10010 2465 10050 2470
rect 10120 2470 10125 2475
rect 10155 2495 10160 2500
rect 10230 2500 10270 2505
rect 10230 2495 10235 2500
rect 10155 2475 10235 2495
rect 10155 2470 10160 2475
rect 10120 2465 10160 2470
rect 10230 2470 10235 2475
rect 10265 2495 10270 2500
rect 10340 2500 10380 2505
rect 10340 2495 10345 2500
rect 10265 2475 10345 2495
rect 10265 2470 10270 2475
rect 10230 2465 10270 2470
rect 10340 2470 10345 2475
rect 10375 2495 10380 2500
rect 10450 2500 10490 2505
rect 10450 2495 10455 2500
rect 10375 2475 10455 2495
rect 10375 2470 10380 2475
rect 10340 2465 10380 2470
rect 10450 2470 10455 2475
rect 10485 2495 10490 2500
rect 10560 2500 10600 2505
rect 10560 2495 10565 2500
rect 10485 2475 10565 2495
rect 10485 2470 10490 2475
rect 10450 2465 10490 2470
rect 10560 2470 10565 2475
rect 10595 2495 10600 2500
rect 10670 2500 10710 2505
rect 10670 2495 10675 2500
rect 10595 2475 10675 2495
rect 10595 2470 10600 2475
rect 10560 2465 10600 2470
rect 10670 2470 10675 2475
rect 10705 2495 10710 2500
rect 10780 2500 10820 2505
rect 10780 2495 10785 2500
rect 10705 2475 10785 2495
rect 10705 2470 10710 2475
rect 10670 2465 10710 2470
rect 10780 2470 10785 2475
rect 10815 2470 10820 2500
rect 13000 2500 13040 2505
rect 10780 2465 10820 2470
rect 10980 2475 11020 2480
rect 10980 2445 10985 2475
rect 11015 2470 11020 2475
rect 11823 2475 11857 2480
rect 11823 2470 11826 2475
rect 11015 2450 11826 2470
rect 11015 2445 11020 2450
rect 10813 2440 10847 2445
rect 10980 2440 11020 2445
rect 11823 2445 11826 2450
rect 11854 2445 11857 2475
rect 13000 2470 13005 2500
rect 13035 2495 13040 2500
rect 13110 2500 13150 2505
rect 13110 2495 13115 2500
rect 13035 2475 13115 2495
rect 13035 2470 13040 2475
rect 13000 2465 13040 2470
rect 13110 2470 13115 2475
rect 13145 2495 13150 2500
rect 13220 2500 13260 2505
rect 13220 2495 13225 2500
rect 13145 2475 13225 2495
rect 13145 2470 13150 2475
rect 13110 2465 13150 2470
rect 13220 2470 13225 2475
rect 13255 2495 13260 2500
rect 13330 2500 13370 2505
rect 13330 2495 13335 2500
rect 13255 2475 13335 2495
rect 13255 2470 13260 2475
rect 13220 2465 13260 2470
rect 13330 2470 13335 2475
rect 13365 2495 13370 2500
rect 13440 2500 13480 2505
rect 13440 2495 13445 2500
rect 13365 2475 13445 2495
rect 13365 2470 13370 2475
rect 13330 2465 13370 2470
rect 13440 2470 13445 2475
rect 13475 2495 13480 2500
rect 13550 2500 13590 2505
rect 13550 2495 13555 2500
rect 13475 2475 13555 2495
rect 13475 2470 13480 2475
rect 13440 2465 13480 2470
rect 13550 2470 13555 2475
rect 13585 2495 13590 2500
rect 13660 2500 13700 2505
rect 13660 2495 13665 2500
rect 13585 2475 13665 2495
rect 13585 2470 13590 2475
rect 13550 2465 13590 2470
rect 13660 2470 13665 2475
rect 13695 2495 13700 2500
rect 13770 2500 13810 2505
rect 13770 2495 13775 2500
rect 13695 2475 13775 2495
rect 13695 2470 13700 2475
rect 13660 2465 13700 2470
rect 13770 2470 13775 2475
rect 13805 2495 13810 2500
rect 13880 2500 13920 2505
rect 13880 2495 13885 2500
rect 13805 2475 13885 2495
rect 13805 2470 13810 2475
rect 13770 2465 13810 2470
rect 13880 2470 13885 2475
rect 13915 2495 13920 2500
rect 13990 2500 14030 2505
rect 13990 2495 13995 2500
rect 13915 2475 13995 2495
rect 13915 2470 13920 2475
rect 13880 2465 13920 2470
rect 13990 2470 13995 2475
rect 14025 2470 14030 2500
rect 13990 2465 14030 2470
rect 17290 2500 17330 2505
rect 17290 2470 17295 2500
rect 17325 2495 17330 2500
rect 17400 2500 17440 2505
rect 17400 2495 17405 2500
rect 17325 2475 17405 2495
rect 17325 2470 17330 2475
rect 17290 2465 17330 2470
rect 17400 2470 17405 2475
rect 17435 2495 17440 2500
rect 17510 2500 17550 2505
rect 17510 2495 17515 2500
rect 17435 2475 17515 2495
rect 17435 2470 17440 2475
rect 17400 2465 17440 2470
rect 17510 2470 17515 2475
rect 17545 2495 17550 2500
rect 17620 2500 17660 2505
rect 17620 2495 17625 2500
rect 17545 2475 17625 2495
rect 17545 2470 17550 2475
rect 17510 2465 17550 2470
rect 17620 2470 17625 2475
rect 17655 2495 17660 2500
rect 17730 2500 17770 2505
rect 17730 2495 17735 2500
rect 17655 2475 17735 2495
rect 17655 2470 17660 2475
rect 17620 2465 17660 2470
rect 17730 2470 17735 2475
rect 17765 2495 17770 2500
rect 17840 2500 17880 2505
rect 17840 2495 17845 2500
rect 17765 2475 17845 2495
rect 17765 2470 17770 2475
rect 17730 2465 17770 2470
rect 17840 2470 17845 2475
rect 17875 2495 17880 2500
rect 17950 2500 17990 2505
rect 17950 2495 17955 2500
rect 17875 2475 17955 2495
rect 17875 2470 17880 2475
rect 17840 2465 17880 2470
rect 17950 2470 17955 2475
rect 17985 2495 17990 2500
rect 18060 2500 18100 2505
rect 18060 2495 18065 2500
rect 17985 2475 18065 2495
rect 17985 2470 17990 2475
rect 17950 2465 17990 2470
rect 18060 2470 18065 2475
rect 18095 2495 18100 2500
rect 18170 2500 18210 2505
rect 18170 2495 18175 2500
rect 18095 2475 18175 2495
rect 18095 2470 18100 2475
rect 18060 2465 18100 2470
rect 18170 2470 18175 2475
rect 18205 2495 18210 2500
rect 18280 2500 18320 2505
rect 18280 2495 18285 2500
rect 18205 2475 18285 2495
rect 18205 2470 18210 2475
rect 18170 2465 18210 2470
rect 18280 2470 18285 2475
rect 18315 2470 18320 2500
rect 20500 2500 20540 2505
rect 18280 2465 18320 2470
rect 18480 2475 18520 2480
rect 18480 2445 18485 2475
rect 18515 2470 18520 2475
rect 19323 2475 19357 2480
rect 19323 2470 19326 2475
rect 18515 2450 19326 2470
rect 18515 2445 18520 2450
rect 11823 2440 11857 2445
rect 12973 2440 13007 2445
rect 10813 2410 10816 2440
rect 10844 2425 10847 2440
rect 10844 2420 11320 2425
rect 10844 2410 11285 2420
rect 10813 2405 11285 2410
rect 11280 2390 11285 2405
rect 11315 2415 11320 2420
rect 11520 2420 11560 2425
rect 11520 2415 11525 2420
rect 11315 2395 11525 2415
rect 11315 2390 11320 2395
rect 11280 2385 11320 2390
rect 11520 2390 11525 2395
rect 11555 2415 11560 2420
rect 11760 2420 11800 2425
rect 11760 2415 11765 2420
rect 11555 2395 11765 2415
rect 11555 2390 11560 2395
rect 11520 2385 11560 2390
rect 11760 2390 11765 2395
rect 11795 2415 11800 2420
rect 12000 2420 12040 2425
rect 12000 2415 12005 2420
rect 11795 2395 12005 2415
rect 11795 2390 11800 2395
rect 11760 2385 11800 2390
rect 12000 2390 12005 2395
rect 12035 2415 12040 2420
rect 12240 2420 12280 2425
rect 12240 2415 12245 2420
rect 12035 2395 12245 2415
rect 12035 2390 12040 2395
rect 12000 2385 12040 2390
rect 12240 2390 12245 2395
rect 12275 2415 12280 2420
rect 12480 2420 12520 2425
rect 12480 2415 12485 2420
rect 12275 2395 12485 2415
rect 12275 2390 12280 2395
rect 12240 2385 12280 2390
rect 12480 2390 12485 2395
rect 12515 2390 12520 2420
rect 12973 2410 12976 2440
rect 13004 2410 13007 2440
rect 12973 2405 13007 2410
rect 18313 2440 18347 2445
rect 18480 2440 18520 2445
rect 19323 2445 19326 2450
rect 19354 2445 19357 2475
rect 20500 2470 20505 2500
rect 20535 2495 20540 2500
rect 20610 2500 20650 2505
rect 20610 2495 20615 2500
rect 20535 2475 20615 2495
rect 20535 2470 20540 2475
rect 20500 2465 20540 2470
rect 20610 2470 20615 2475
rect 20645 2495 20650 2500
rect 20720 2500 20760 2505
rect 20720 2495 20725 2500
rect 20645 2475 20725 2495
rect 20645 2470 20650 2475
rect 20610 2465 20650 2470
rect 20720 2470 20725 2475
rect 20755 2495 20760 2500
rect 20830 2500 20870 2505
rect 20830 2495 20835 2500
rect 20755 2475 20835 2495
rect 20755 2470 20760 2475
rect 20720 2465 20760 2470
rect 20830 2470 20835 2475
rect 20865 2495 20870 2500
rect 20940 2500 20980 2505
rect 20940 2495 20945 2500
rect 20865 2475 20945 2495
rect 20865 2470 20870 2475
rect 20830 2465 20870 2470
rect 20940 2470 20945 2475
rect 20975 2495 20980 2500
rect 21050 2500 21090 2505
rect 21050 2495 21055 2500
rect 20975 2475 21055 2495
rect 20975 2470 20980 2475
rect 20940 2465 20980 2470
rect 21050 2470 21055 2475
rect 21085 2495 21090 2500
rect 21160 2500 21200 2505
rect 21160 2495 21165 2500
rect 21085 2475 21165 2495
rect 21085 2470 21090 2475
rect 21050 2465 21090 2470
rect 21160 2470 21165 2475
rect 21195 2495 21200 2500
rect 21270 2500 21310 2505
rect 21270 2495 21275 2500
rect 21195 2475 21275 2495
rect 21195 2470 21200 2475
rect 21160 2465 21200 2470
rect 21270 2470 21275 2475
rect 21305 2495 21310 2500
rect 21380 2500 21420 2505
rect 21380 2495 21385 2500
rect 21305 2475 21385 2495
rect 21305 2470 21310 2475
rect 21270 2465 21310 2470
rect 21380 2470 21385 2475
rect 21415 2495 21420 2500
rect 21490 2500 21530 2505
rect 21490 2495 21495 2500
rect 21415 2475 21495 2495
rect 21415 2470 21420 2475
rect 21380 2465 21420 2470
rect 21490 2470 21495 2475
rect 21525 2470 21530 2500
rect 21490 2465 21530 2470
rect 19323 2440 19357 2445
rect 20473 2440 20507 2445
rect 18313 2410 18316 2440
rect 18344 2425 18347 2440
rect 18344 2420 18820 2425
rect 18344 2410 18785 2420
rect 18313 2405 18785 2410
rect 12480 2385 12520 2390
rect 18780 2390 18785 2405
rect 18815 2415 18820 2420
rect 19020 2420 19060 2425
rect 19020 2415 19025 2420
rect 18815 2395 19025 2415
rect 18815 2390 18820 2395
rect 18780 2385 18820 2390
rect 19020 2390 19025 2395
rect 19055 2415 19060 2420
rect 19260 2420 19300 2425
rect 19260 2415 19265 2420
rect 19055 2395 19265 2415
rect 19055 2390 19060 2395
rect 19020 2385 19060 2390
rect 19260 2390 19265 2395
rect 19295 2415 19300 2420
rect 19500 2420 19540 2425
rect 19500 2415 19505 2420
rect 19295 2395 19505 2415
rect 19295 2390 19300 2395
rect 19260 2385 19300 2390
rect 19500 2390 19505 2395
rect 19535 2415 19540 2420
rect 19740 2420 19780 2425
rect 19740 2415 19745 2420
rect 19535 2395 19745 2415
rect 19535 2390 19540 2395
rect 19500 2385 19540 2390
rect 19740 2390 19745 2395
rect 19775 2415 19780 2420
rect 19980 2420 20020 2425
rect 19980 2415 19985 2420
rect 19775 2395 19985 2415
rect 19775 2390 19780 2395
rect 19740 2385 19780 2390
rect 19980 2390 19985 2395
rect 20015 2390 20020 2420
rect 20473 2410 20476 2440
rect 20504 2410 20507 2440
rect 20473 2405 20507 2410
rect 19980 2385 20020 2390
rect 3805 2380 3845 2385
rect 3355 2375 3395 2380
rect 2620 2345 2660 2350
rect 2620 2315 2625 2345
rect 2655 2340 2660 2345
rect 3355 2345 3360 2375
rect 3390 2345 3395 2375
rect 3805 2350 3810 2380
rect 3840 2375 3845 2380
rect 4165 2380 4205 2385
rect 4165 2375 4170 2380
rect 3840 2355 4170 2375
rect 3840 2350 3845 2355
rect 3805 2345 3845 2350
rect 4165 2350 4170 2355
rect 4200 2350 4205 2380
rect 4165 2345 4205 2350
rect 9800 2345 9805 2380
rect 9840 2345 9845 2380
rect 10635 2345 10640 2380
rect 10675 2345 10680 2380
rect 11400 2375 11440 2380
rect 11400 2345 11405 2375
rect 11435 2370 11440 2375
rect 11640 2375 11680 2380
rect 11640 2370 11645 2375
rect 11435 2350 11645 2370
rect 11435 2345 11440 2350
rect 3355 2340 3395 2345
rect 11400 2340 11440 2345
rect 11640 2345 11645 2350
rect 11675 2370 11680 2375
rect 11880 2375 11920 2380
rect 11880 2370 11885 2375
rect 11675 2350 11885 2370
rect 11675 2345 11680 2350
rect 11640 2340 11680 2345
rect 11880 2345 11885 2350
rect 11915 2370 11920 2375
rect 12120 2375 12160 2380
rect 12120 2370 12125 2375
rect 11915 2350 12125 2370
rect 11915 2345 11920 2350
rect 11880 2340 11920 2345
rect 12120 2345 12125 2350
rect 12155 2370 12160 2375
rect 12360 2375 12400 2380
rect 12360 2370 12365 2375
rect 12155 2350 12365 2370
rect 12155 2345 12160 2350
rect 12120 2340 12160 2345
rect 12360 2345 12365 2350
rect 12395 2370 12400 2375
rect 12690 2375 12730 2380
rect 12690 2370 12695 2375
rect 12395 2350 12695 2370
rect 12395 2345 12400 2350
rect 12360 2340 12400 2345
rect 12690 2345 12695 2350
rect 12725 2370 12730 2375
rect 12970 2375 13010 2380
rect 12970 2370 12975 2375
rect 12725 2350 12975 2370
rect 12725 2345 12730 2350
rect 12690 2340 12730 2345
rect 12970 2345 12975 2350
rect 13005 2345 13010 2375
rect 13140 2345 13145 2380
rect 13180 2345 13185 2380
rect 13974 2345 13980 2380
rect 14015 2345 14020 2380
rect 17300 2345 17305 2380
rect 17340 2345 17345 2380
rect 18135 2345 18140 2380
rect 18175 2345 18180 2380
rect 18900 2375 18940 2380
rect 18900 2345 18905 2375
rect 18935 2370 18940 2375
rect 19140 2375 19180 2380
rect 19140 2370 19145 2375
rect 18935 2350 19145 2370
rect 18935 2345 18940 2350
rect 12970 2340 13010 2345
rect 18900 2340 18940 2345
rect 19140 2345 19145 2350
rect 19175 2370 19180 2375
rect 19380 2375 19420 2380
rect 19380 2370 19385 2375
rect 19175 2350 19385 2370
rect 19175 2345 19180 2350
rect 19140 2340 19180 2345
rect 19380 2345 19385 2350
rect 19415 2370 19420 2375
rect 19620 2375 19660 2380
rect 19620 2370 19625 2375
rect 19415 2350 19625 2370
rect 19415 2345 19420 2350
rect 19380 2340 19420 2345
rect 19620 2345 19625 2350
rect 19655 2370 19660 2375
rect 19860 2375 19900 2380
rect 19860 2370 19865 2375
rect 19655 2350 19865 2370
rect 19655 2345 19660 2350
rect 19620 2340 19660 2345
rect 19860 2345 19865 2350
rect 19895 2370 19900 2375
rect 20190 2375 20230 2380
rect 20190 2370 20195 2375
rect 19895 2350 20195 2370
rect 19895 2345 19900 2350
rect 19860 2340 19900 2345
rect 20190 2345 20195 2350
rect 20225 2370 20230 2375
rect 20470 2375 20510 2380
rect 20470 2370 20475 2375
rect 20225 2350 20475 2370
rect 20225 2345 20230 2350
rect 20190 2340 20230 2345
rect 20470 2345 20475 2350
rect 20505 2345 20510 2375
rect 20640 2345 20645 2380
rect 20680 2345 20685 2380
rect 21474 2345 21480 2380
rect 21515 2345 21520 2380
rect 20470 2340 20510 2345
rect 2655 2320 3395 2340
rect 3625 2335 3665 2340
rect 2655 2315 2660 2320
rect 2620 2310 2660 2315
rect 3625 2305 3630 2335
rect 3660 2330 3665 2335
rect 4345 2335 4385 2340
rect 4345 2330 4350 2335
rect 3660 2310 4350 2330
rect 3660 2305 3665 2310
rect 3625 2300 3665 2305
rect 4345 2305 4350 2310
rect 4380 2305 4385 2335
rect 12815 2325 12855 2330
rect 12815 2320 12820 2325
rect 4345 2300 4385 2305
rect 2735 2290 2775 2295
rect 2735 2260 2740 2290
rect 2770 2285 2775 2290
rect 3445 2290 3485 2295
rect 3445 2285 3450 2290
rect 2770 2265 3450 2285
rect 2770 2260 2775 2265
rect 2735 2255 2775 2260
rect 3445 2260 3450 2265
rect 3480 2285 3485 2290
rect 4525 2290 4565 2295
rect 4525 2285 4530 2290
rect 3480 2265 4530 2285
rect 3480 2260 3485 2265
rect 3445 2255 3485 2260
rect 4525 2260 4530 2265
rect 4560 2285 4565 2290
rect 5270 2290 5310 2295
rect 5270 2285 5275 2290
rect 4560 2265 5275 2285
rect 4560 2260 4565 2265
rect 4525 2255 4565 2260
rect 5270 2260 5275 2265
rect 5305 2260 5310 2290
rect 9800 2285 9805 2320
rect 9840 2285 9845 2320
rect 10635 2285 10640 2320
rect 10675 2300 12820 2320
rect 10675 2285 10680 2300
rect 12815 2295 12820 2300
rect 12850 2320 12855 2325
rect 20315 2325 20355 2330
rect 20315 2320 20320 2325
rect 12850 2300 13145 2320
rect 12850 2295 12855 2300
rect 12815 2290 12855 2295
rect 13140 2285 13145 2300
rect 13180 2285 13185 2320
rect 13975 2285 13980 2320
rect 14015 2285 14020 2320
rect 17300 2285 17305 2320
rect 17340 2285 17345 2320
rect 18135 2285 18140 2320
rect 18175 2300 20320 2320
rect 18175 2285 18180 2300
rect 20315 2295 20320 2300
rect 20350 2320 20355 2325
rect 20350 2300 20645 2320
rect 20350 2295 20355 2300
rect 20315 2290 20355 2295
rect 20640 2285 20645 2300
rect 20680 2285 20685 2320
rect 21475 2285 21480 2320
rect 21515 2285 21520 2320
rect 5270 2255 5310 2260
rect 10813 2280 10847 2285
rect 10813 2250 10816 2280
rect 10844 2250 10847 2280
rect 2425 2245 2465 2250
rect 2425 2215 2430 2245
rect 2460 2240 2465 2245
rect 3805 2245 3845 2250
rect 10813 2245 10847 2250
rect 11440 2280 11480 2285
rect 11440 2250 11445 2280
rect 11475 2275 11480 2280
rect 11660 2280 11700 2285
rect 11660 2275 11665 2280
rect 11475 2255 11665 2275
rect 11475 2250 11480 2255
rect 11440 2245 11480 2250
rect 11660 2250 11665 2255
rect 11695 2275 11700 2280
rect 11880 2280 11920 2285
rect 11880 2275 11885 2280
rect 11695 2255 11885 2275
rect 11695 2250 11700 2255
rect 11660 2245 11700 2250
rect 11880 2250 11885 2255
rect 11915 2275 11920 2280
rect 12100 2280 12140 2285
rect 12100 2275 12105 2280
rect 11915 2255 12105 2275
rect 11915 2250 11920 2255
rect 11880 2245 11920 2250
rect 12100 2250 12105 2255
rect 12135 2275 12140 2280
rect 12320 2280 12360 2285
rect 12320 2275 12325 2280
rect 12135 2255 12325 2275
rect 12135 2250 12140 2255
rect 12100 2245 12140 2250
rect 12320 2250 12325 2255
rect 12355 2250 12360 2280
rect 12320 2245 12360 2250
rect 12973 2280 13007 2285
rect 12973 2250 12976 2280
rect 13004 2250 13007 2280
rect 12973 2245 13007 2250
rect 18313 2280 18347 2285
rect 18313 2250 18316 2280
rect 18344 2250 18347 2280
rect 18313 2245 18347 2250
rect 18940 2280 18980 2285
rect 18940 2250 18945 2280
rect 18975 2275 18980 2280
rect 19160 2280 19200 2285
rect 19160 2275 19165 2280
rect 18975 2255 19165 2275
rect 18975 2250 18980 2255
rect 18940 2245 18980 2250
rect 19160 2250 19165 2255
rect 19195 2275 19200 2280
rect 19380 2280 19420 2285
rect 19380 2275 19385 2280
rect 19195 2255 19385 2275
rect 19195 2250 19200 2255
rect 19160 2245 19200 2250
rect 19380 2250 19385 2255
rect 19415 2275 19420 2280
rect 19600 2280 19640 2285
rect 19600 2275 19605 2280
rect 19415 2255 19605 2275
rect 19415 2250 19420 2255
rect 19380 2245 19420 2250
rect 19600 2250 19605 2255
rect 19635 2275 19640 2280
rect 19820 2280 19860 2285
rect 19820 2275 19825 2280
rect 19635 2255 19825 2275
rect 19635 2250 19640 2255
rect 19600 2245 19640 2250
rect 19820 2250 19825 2255
rect 19855 2250 19860 2280
rect 19820 2245 19860 2250
rect 20473 2280 20507 2285
rect 20473 2250 20476 2280
rect 20504 2250 20507 2280
rect 20473 2245 20507 2250
rect 3805 2240 3810 2245
rect 2460 2220 3810 2240
rect 2460 2215 2465 2220
rect 2425 2210 2465 2215
rect 3805 2215 3810 2220
rect 3840 2215 3845 2245
rect 11330 2235 11370 2240
rect 3805 2210 3845 2215
rect 9790 2220 9830 2225
rect 2330 2200 2370 2205
rect 2330 2170 2335 2200
rect 2365 2195 2370 2200
rect 3265 2200 3305 2205
rect 3265 2195 3270 2200
rect 2365 2175 3270 2195
rect 2365 2170 2370 2175
rect 2330 2165 2370 2170
rect 3265 2170 3270 2175
rect 3300 2195 3305 2200
rect 3985 2200 4025 2205
rect 3985 2195 3990 2200
rect 3300 2175 3990 2195
rect 3300 2170 3305 2175
rect 3265 2165 3305 2170
rect 3985 2170 3990 2175
rect 4020 2195 4025 2200
rect 4705 2200 4745 2205
rect 4705 2195 4710 2200
rect 4020 2175 4710 2195
rect 4020 2170 4025 2175
rect 3985 2165 4025 2170
rect 4705 2170 4710 2175
rect 4740 2170 4745 2200
rect 9790 2190 9795 2220
rect 9825 2215 9830 2220
rect 9900 2220 9940 2225
rect 9900 2215 9905 2220
rect 9825 2195 9905 2215
rect 9825 2190 9830 2195
rect 9790 2185 9830 2190
rect 9900 2190 9905 2195
rect 9935 2215 9940 2220
rect 10010 2220 10050 2225
rect 10010 2215 10015 2220
rect 9935 2195 10015 2215
rect 9935 2190 9940 2195
rect 9900 2185 9940 2190
rect 10010 2190 10015 2195
rect 10045 2215 10050 2220
rect 10120 2220 10160 2225
rect 10120 2215 10125 2220
rect 10045 2195 10125 2215
rect 10045 2190 10050 2195
rect 10010 2185 10050 2190
rect 10120 2190 10125 2195
rect 10155 2215 10160 2220
rect 10230 2220 10270 2225
rect 10230 2215 10235 2220
rect 10155 2195 10235 2215
rect 10155 2190 10160 2195
rect 10120 2185 10160 2190
rect 10230 2190 10235 2195
rect 10265 2215 10270 2220
rect 10340 2220 10380 2225
rect 10340 2215 10345 2220
rect 10265 2195 10345 2215
rect 10265 2190 10270 2195
rect 10230 2185 10270 2190
rect 10340 2190 10345 2195
rect 10375 2215 10380 2220
rect 10450 2220 10490 2225
rect 10450 2215 10455 2220
rect 10375 2195 10455 2215
rect 10375 2190 10380 2195
rect 10340 2185 10380 2190
rect 10450 2190 10455 2195
rect 10485 2215 10490 2220
rect 10560 2220 10600 2225
rect 10560 2215 10565 2220
rect 10485 2195 10565 2215
rect 10485 2190 10490 2195
rect 10450 2185 10490 2190
rect 10560 2190 10565 2195
rect 10595 2215 10600 2220
rect 10670 2220 10710 2225
rect 10670 2215 10675 2220
rect 10595 2195 10675 2215
rect 10595 2190 10600 2195
rect 10560 2185 10600 2190
rect 10670 2190 10675 2195
rect 10705 2215 10710 2220
rect 10780 2220 10820 2225
rect 10780 2215 10785 2220
rect 10705 2195 10785 2215
rect 10705 2190 10710 2195
rect 10670 2185 10710 2190
rect 10780 2190 10785 2195
rect 10815 2190 10820 2220
rect 11330 2205 11335 2235
rect 11365 2230 11370 2235
rect 11550 2235 11590 2240
rect 11550 2230 11555 2235
rect 11365 2210 11555 2230
rect 11365 2205 11370 2210
rect 11330 2200 11370 2205
rect 11550 2205 11555 2210
rect 11585 2230 11590 2235
rect 11770 2235 11810 2240
rect 11770 2230 11775 2235
rect 11585 2210 11775 2230
rect 11585 2205 11590 2210
rect 11550 2200 11590 2205
rect 11770 2205 11775 2210
rect 11805 2230 11810 2235
rect 11990 2235 12030 2240
rect 11990 2230 11995 2235
rect 11805 2210 11995 2230
rect 11805 2205 11810 2210
rect 11770 2200 11810 2205
rect 11990 2205 11995 2210
rect 12025 2230 12030 2235
rect 12210 2235 12250 2240
rect 12210 2230 12215 2235
rect 12025 2210 12215 2230
rect 12025 2205 12030 2210
rect 11990 2200 12030 2205
rect 12210 2205 12215 2210
rect 12245 2230 12250 2235
rect 12430 2235 12470 2240
rect 12430 2230 12435 2235
rect 12245 2210 12435 2230
rect 12245 2205 12250 2210
rect 12210 2200 12250 2205
rect 12430 2205 12435 2210
rect 12465 2205 12470 2235
rect 18830 2235 18870 2240
rect 12430 2200 12470 2205
rect 13000 2220 13040 2225
rect 10780 2185 10820 2190
rect 13000 2190 13005 2220
rect 13035 2215 13040 2220
rect 13110 2220 13150 2225
rect 13110 2215 13115 2220
rect 13035 2195 13115 2215
rect 13035 2190 13040 2195
rect 13000 2185 13040 2190
rect 13110 2190 13115 2195
rect 13145 2215 13150 2220
rect 13220 2220 13260 2225
rect 13220 2215 13225 2220
rect 13145 2195 13225 2215
rect 13145 2190 13150 2195
rect 13110 2185 13150 2190
rect 13220 2190 13225 2195
rect 13255 2215 13260 2220
rect 13330 2220 13370 2225
rect 13330 2215 13335 2220
rect 13255 2195 13335 2215
rect 13255 2190 13260 2195
rect 13220 2185 13260 2190
rect 13330 2190 13335 2195
rect 13365 2215 13370 2220
rect 13440 2220 13480 2225
rect 13440 2215 13445 2220
rect 13365 2195 13445 2215
rect 13365 2190 13370 2195
rect 13330 2185 13370 2190
rect 13440 2190 13445 2195
rect 13475 2215 13480 2220
rect 13550 2220 13590 2225
rect 13550 2215 13555 2220
rect 13475 2195 13555 2215
rect 13475 2190 13480 2195
rect 13440 2185 13480 2190
rect 13550 2190 13555 2195
rect 13585 2215 13590 2220
rect 13660 2220 13700 2225
rect 13660 2215 13665 2220
rect 13585 2195 13665 2215
rect 13585 2190 13590 2195
rect 13550 2185 13590 2190
rect 13660 2190 13665 2195
rect 13695 2215 13700 2220
rect 13770 2220 13810 2225
rect 13770 2215 13775 2220
rect 13695 2195 13775 2215
rect 13695 2190 13700 2195
rect 13660 2185 13700 2190
rect 13770 2190 13775 2195
rect 13805 2215 13810 2220
rect 13880 2220 13920 2225
rect 13880 2215 13885 2220
rect 13805 2195 13885 2215
rect 13805 2190 13810 2195
rect 13770 2185 13810 2190
rect 13880 2190 13885 2195
rect 13915 2215 13920 2220
rect 13990 2220 14030 2225
rect 13990 2215 13995 2220
rect 13915 2195 13995 2215
rect 13915 2190 13920 2195
rect 13880 2185 13920 2190
rect 13990 2190 13995 2195
rect 14025 2190 14030 2220
rect 13990 2185 14030 2190
rect 17290 2220 17330 2225
rect 17290 2190 17295 2220
rect 17325 2215 17330 2220
rect 17400 2220 17440 2225
rect 17400 2215 17405 2220
rect 17325 2195 17405 2215
rect 17325 2190 17330 2195
rect 17290 2185 17330 2190
rect 17400 2190 17405 2195
rect 17435 2215 17440 2220
rect 17510 2220 17550 2225
rect 17510 2215 17515 2220
rect 17435 2195 17515 2215
rect 17435 2190 17440 2195
rect 17400 2185 17440 2190
rect 17510 2190 17515 2195
rect 17545 2215 17550 2220
rect 17620 2220 17660 2225
rect 17620 2215 17625 2220
rect 17545 2195 17625 2215
rect 17545 2190 17550 2195
rect 17510 2185 17550 2190
rect 17620 2190 17625 2195
rect 17655 2215 17660 2220
rect 17730 2220 17770 2225
rect 17730 2215 17735 2220
rect 17655 2195 17735 2215
rect 17655 2190 17660 2195
rect 17620 2185 17660 2190
rect 17730 2190 17735 2195
rect 17765 2215 17770 2220
rect 17840 2220 17880 2225
rect 17840 2215 17845 2220
rect 17765 2195 17845 2215
rect 17765 2190 17770 2195
rect 17730 2185 17770 2190
rect 17840 2190 17845 2195
rect 17875 2215 17880 2220
rect 17950 2220 17990 2225
rect 17950 2215 17955 2220
rect 17875 2195 17955 2215
rect 17875 2190 17880 2195
rect 17840 2185 17880 2190
rect 17950 2190 17955 2195
rect 17985 2215 17990 2220
rect 18060 2220 18100 2225
rect 18060 2215 18065 2220
rect 17985 2195 18065 2215
rect 17985 2190 17990 2195
rect 17950 2185 17990 2190
rect 18060 2190 18065 2195
rect 18095 2215 18100 2220
rect 18170 2220 18210 2225
rect 18170 2215 18175 2220
rect 18095 2195 18175 2215
rect 18095 2190 18100 2195
rect 18060 2185 18100 2190
rect 18170 2190 18175 2195
rect 18205 2215 18210 2220
rect 18280 2220 18320 2225
rect 18280 2215 18285 2220
rect 18205 2195 18285 2215
rect 18205 2190 18210 2195
rect 18170 2185 18210 2190
rect 18280 2190 18285 2195
rect 18315 2190 18320 2220
rect 18830 2205 18835 2235
rect 18865 2230 18870 2235
rect 19050 2235 19090 2240
rect 19050 2230 19055 2235
rect 18865 2210 19055 2230
rect 18865 2205 18870 2210
rect 18830 2200 18870 2205
rect 19050 2205 19055 2210
rect 19085 2230 19090 2235
rect 19270 2235 19310 2240
rect 19270 2230 19275 2235
rect 19085 2210 19275 2230
rect 19085 2205 19090 2210
rect 19050 2200 19090 2205
rect 19270 2205 19275 2210
rect 19305 2230 19310 2235
rect 19490 2235 19530 2240
rect 19490 2230 19495 2235
rect 19305 2210 19495 2230
rect 19305 2205 19310 2210
rect 19270 2200 19310 2205
rect 19490 2205 19495 2210
rect 19525 2230 19530 2235
rect 19710 2235 19750 2240
rect 19710 2230 19715 2235
rect 19525 2210 19715 2230
rect 19525 2205 19530 2210
rect 19490 2200 19530 2205
rect 19710 2205 19715 2210
rect 19745 2230 19750 2235
rect 19930 2235 19970 2240
rect 19930 2230 19935 2235
rect 19745 2210 19935 2230
rect 19745 2205 19750 2210
rect 19710 2200 19750 2205
rect 19930 2205 19935 2210
rect 19965 2205 19970 2235
rect 19930 2200 19970 2205
rect 20500 2220 20540 2225
rect 18280 2185 18320 2190
rect 20500 2190 20505 2220
rect 20535 2215 20540 2220
rect 20610 2220 20650 2225
rect 20610 2215 20615 2220
rect 20535 2195 20615 2215
rect 20535 2190 20540 2195
rect 20500 2185 20540 2190
rect 20610 2190 20615 2195
rect 20645 2215 20650 2220
rect 20720 2220 20760 2225
rect 20720 2215 20725 2220
rect 20645 2195 20725 2215
rect 20645 2190 20650 2195
rect 20610 2185 20650 2190
rect 20720 2190 20725 2195
rect 20755 2215 20760 2220
rect 20830 2220 20870 2225
rect 20830 2215 20835 2220
rect 20755 2195 20835 2215
rect 20755 2190 20760 2195
rect 20720 2185 20760 2190
rect 20830 2190 20835 2195
rect 20865 2215 20870 2220
rect 20940 2220 20980 2225
rect 20940 2215 20945 2220
rect 20865 2195 20945 2215
rect 20865 2190 20870 2195
rect 20830 2185 20870 2190
rect 20940 2190 20945 2195
rect 20975 2215 20980 2220
rect 21050 2220 21090 2225
rect 21050 2215 21055 2220
rect 20975 2195 21055 2215
rect 20975 2190 20980 2195
rect 20940 2185 20980 2190
rect 21050 2190 21055 2195
rect 21085 2215 21090 2220
rect 21160 2220 21200 2225
rect 21160 2215 21165 2220
rect 21085 2195 21165 2215
rect 21085 2190 21090 2195
rect 21050 2185 21090 2190
rect 21160 2190 21165 2195
rect 21195 2215 21200 2220
rect 21270 2220 21310 2225
rect 21270 2215 21275 2220
rect 21195 2195 21275 2215
rect 21195 2190 21200 2195
rect 21160 2185 21200 2190
rect 21270 2190 21275 2195
rect 21305 2215 21310 2220
rect 21380 2220 21420 2225
rect 21380 2215 21385 2220
rect 21305 2195 21385 2215
rect 21305 2190 21310 2195
rect 21270 2185 21310 2190
rect 21380 2190 21385 2195
rect 21415 2215 21420 2220
rect 21490 2220 21530 2225
rect 21490 2215 21495 2220
rect 21415 2195 21495 2215
rect 21415 2190 21420 2195
rect 21380 2185 21420 2190
rect 21490 2190 21495 2195
rect 21525 2190 21530 2220
rect 21490 2185 21530 2190
rect 4705 2165 4745 2170
rect 2380 2150 2420 2155
rect 2380 2120 2385 2150
rect 2415 2145 2420 2150
rect 3625 2150 3665 2155
rect 3625 2145 3630 2150
rect 2415 2125 3630 2145
rect 2415 2120 2420 2125
rect 2380 2115 2420 2120
rect 3625 2120 3630 2125
rect 3660 2120 3665 2150
rect 3625 2115 3665 2120
rect 4085 2145 4125 2150
rect 4085 2115 4090 2145
rect 4120 2140 4125 2145
rect 5315 2145 5355 2150
rect 5315 2140 5320 2145
rect 4120 2120 5320 2140
rect 4120 2115 4125 2120
rect 4085 2110 4125 2115
rect 5315 2115 5320 2120
rect 5350 2115 5355 2145
rect 5315 2110 5355 2115
rect 2745 2095 2785 2100
rect 2745 2065 2750 2095
rect 2780 2090 2785 2095
rect 2865 2095 2905 2100
rect 2865 2090 2870 2095
rect 2780 2070 2870 2090
rect 2780 2065 2785 2070
rect 2745 2060 2785 2065
rect 2865 2065 2870 2070
rect 2900 2090 2905 2095
rect 2985 2095 3025 2100
rect 2985 2090 2990 2095
rect 2900 2070 2990 2090
rect 2900 2065 2905 2070
rect 2865 2060 2905 2065
rect 2985 2065 2990 2070
rect 3020 2090 3025 2095
rect 3105 2095 3145 2100
rect 3105 2090 3110 2095
rect 3020 2070 3110 2090
rect 3020 2065 3025 2070
rect 2985 2060 3025 2065
rect 3105 2065 3110 2070
rect 3140 2090 3145 2095
rect 3225 2095 3265 2100
rect 3225 2090 3230 2095
rect 3140 2070 3230 2090
rect 3140 2065 3145 2070
rect 3105 2060 3145 2065
rect 3225 2065 3230 2070
rect 3260 2090 3265 2095
rect 3345 2095 3385 2100
rect 3345 2090 3350 2095
rect 3260 2070 3350 2090
rect 3260 2065 3265 2070
rect 3225 2060 3265 2065
rect 3345 2065 3350 2070
rect 3380 2090 3385 2095
rect 3465 2095 3505 2100
rect 3465 2090 3470 2095
rect 3380 2070 3470 2090
rect 3380 2065 3385 2070
rect 3345 2060 3385 2065
rect 3465 2065 3470 2070
rect 3500 2090 3505 2095
rect 3585 2095 3625 2100
rect 3585 2090 3590 2095
rect 3500 2070 3590 2090
rect 3500 2065 3505 2070
rect 3465 2060 3505 2065
rect 3585 2065 3590 2070
rect 3620 2090 3625 2095
rect 3705 2095 3745 2100
rect 3705 2090 3710 2095
rect 3620 2070 3710 2090
rect 3620 2065 3625 2070
rect 3585 2060 3625 2065
rect 3705 2065 3710 2070
rect 3740 2090 3745 2095
rect 3825 2095 3865 2100
rect 3825 2090 3830 2095
rect 3740 2070 3830 2090
rect 3740 2065 3745 2070
rect 3705 2060 3745 2065
rect 3825 2065 3830 2070
rect 3860 2090 3865 2095
rect 3985 2095 4025 2100
rect 3985 2090 3990 2095
rect 3860 2070 3990 2090
rect 3860 2065 3865 2070
rect 3825 2060 3865 2065
rect 3985 2065 3990 2070
rect 4020 2090 4025 2095
rect 4145 2095 4185 2100
rect 4145 2090 4150 2095
rect 4020 2070 4150 2090
rect 4020 2065 4025 2070
rect 3985 2060 4025 2065
rect 4145 2065 4150 2070
rect 4180 2090 4185 2095
rect 4265 2095 4305 2100
rect 4265 2090 4270 2095
rect 4180 2070 4270 2090
rect 4180 2065 4185 2070
rect 4145 2060 4185 2065
rect 4265 2065 4270 2070
rect 4300 2090 4305 2095
rect 4385 2095 4425 2100
rect 4385 2090 4390 2095
rect 4300 2070 4390 2090
rect 4300 2065 4305 2070
rect 4265 2060 4305 2065
rect 4385 2065 4390 2070
rect 4420 2090 4425 2095
rect 4505 2095 4545 2100
rect 4505 2090 4510 2095
rect 4420 2070 4510 2090
rect 4420 2065 4425 2070
rect 4385 2060 4425 2065
rect 4505 2065 4510 2070
rect 4540 2090 4545 2095
rect 4625 2095 4665 2100
rect 4625 2090 4630 2095
rect 4540 2070 4630 2090
rect 4540 2065 4545 2070
rect 4505 2060 4545 2065
rect 4625 2065 4630 2070
rect 4660 2090 4665 2095
rect 4745 2095 4785 2100
rect 4745 2090 4750 2095
rect 4660 2070 4750 2090
rect 4660 2065 4665 2070
rect 4625 2060 4665 2065
rect 4745 2065 4750 2070
rect 4780 2090 4785 2095
rect 4865 2095 4905 2100
rect 4865 2090 4870 2095
rect 4780 2070 4870 2090
rect 4780 2065 4785 2070
rect 4745 2060 4785 2065
rect 4865 2065 4870 2070
rect 4900 2090 4905 2095
rect 4985 2095 5025 2100
rect 4985 2090 4990 2095
rect 4900 2070 4990 2090
rect 4900 2065 4905 2070
rect 4865 2060 4905 2065
rect 4985 2065 4990 2070
rect 5020 2090 5025 2095
rect 5105 2095 5145 2100
rect 5105 2090 5110 2095
rect 5020 2070 5110 2090
rect 5020 2065 5025 2070
rect 4985 2060 5025 2065
rect 5105 2065 5110 2070
rect 5140 2090 5145 2095
rect 5225 2095 5265 2100
rect 5225 2090 5230 2095
rect 5140 2070 5230 2090
rect 5140 2065 5145 2070
rect 5105 2060 5145 2065
rect 5225 2065 5230 2070
rect 5260 2090 5265 2095
rect 5550 2095 5590 2100
rect 5550 2090 5555 2095
rect 5260 2070 5555 2090
rect 5260 2065 5265 2070
rect 5225 2060 5265 2065
rect 5550 2065 5555 2070
rect 5585 2065 5590 2095
rect 5550 2060 5590 2065
rect 2620 2050 2660 2055
rect 2620 2020 2625 2050
rect 2655 2020 2660 2050
rect 2620 2015 2660 2020
rect 2805 2050 2845 2055
rect 2805 2020 2810 2050
rect 2840 2045 2845 2050
rect 3165 2050 3205 2055
rect 3165 2045 3170 2050
rect 2840 2025 3170 2045
rect 2840 2020 2845 2025
rect 2805 2015 2845 2020
rect 3165 2020 3170 2025
rect 3200 2045 3205 2050
rect 3525 2050 3565 2055
rect 3525 2045 3530 2050
rect 3200 2025 3530 2045
rect 3200 2020 3205 2025
rect 3165 2015 3205 2020
rect 3525 2020 3530 2025
rect 3560 2045 3565 2050
rect 3885 2050 3925 2055
rect 3885 2045 3890 2050
rect 3560 2025 3890 2045
rect 3560 2020 3565 2025
rect 3525 2015 3565 2020
rect 3885 2020 3890 2025
rect 3920 2020 3925 2050
rect 3885 2015 3925 2020
rect 4085 2050 4125 2055
rect 4085 2020 4090 2050
rect 4120 2045 4125 2050
rect 4445 2050 4485 2055
rect 4445 2045 4450 2050
rect 4120 2025 4450 2045
rect 4120 2020 4125 2025
rect 4085 2015 4125 2020
rect 4445 2020 4450 2025
rect 4480 2045 4485 2050
rect 4805 2050 4845 2055
rect 4805 2045 4810 2050
rect 4480 2025 4810 2045
rect 4480 2020 4485 2025
rect 4445 2015 4485 2020
rect 4805 2020 4810 2025
rect 4840 2045 4845 2050
rect 5165 2050 5205 2055
rect 5165 2045 5170 2050
rect 4840 2025 5170 2045
rect 4840 2020 4845 2025
rect 4805 2015 4845 2020
rect 5165 2020 5170 2025
rect 5200 2020 5205 2050
rect 5165 2015 5205 2020
rect 9735 2000 9775 2005
rect 9735 1970 9740 2000
rect 9770 1995 9775 2000
rect 9845 2000 9885 2005
rect 9845 1995 9850 2000
rect 9770 1975 9850 1995
rect 9770 1970 9775 1975
rect 9735 1965 9775 1970
rect 9845 1970 9850 1975
rect 9880 1995 9885 2000
rect 9955 2000 9995 2005
rect 9955 1995 9960 2000
rect 9880 1975 9960 1995
rect 9880 1970 9885 1975
rect 9845 1965 9885 1970
rect 9955 1970 9960 1975
rect 9990 1995 9995 2000
rect 10065 2000 10105 2005
rect 10065 1995 10070 2000
rect 9990 1975 10070 1995
rect 9990 1970 9995 1975
rect 9955 1965 9995 1970
rect 10065 1970 10070 1975
rect 10100 1995 10105 2000
rect 10175 2000 10215 2005
rect 10175 1995 10180 2000
rect 10100 1975 10180 1995
rect 10100 1970 10105 1975
rect 10065 1965 10105 1970
rect 10175 1970 10180 1975
rect 10210 1995 10215 2000
rect 10285 2000 10325 2005
rect 10285 1995 10290 2000
rect 10210 1975 10290 1995
rect 10210 1970 10215 1975
rect 10175 1965 10215 1970
rect 10285 1970 10290 1975
rect 10320 1995 10325 2000
rect 10395 2000 10435 2005
rect 10395 1995 10400 2000
rect 10320 1975 10400 1995
rect 10320 1970 10325 1975
rect 10285 1965 10325 1970
rect 10395 1970 10400 1975
rect 10430 1995 10435 2000
rect 10505 2000 10545 2005
rect 10505 1995 10510 2000
rect 10430 1975 10510 1995
rect 10430 1970 10435 1975
rect 10395 1965 10435 1970
rect 10505 1970 10510 1975
rect 10540 1995 10545 2000
rect 10615 2000 10655 2005
rect 10615 1995 10620 2000
rect 10540 1975 10620 1995
rect 10540 1970 10545 1975
rect 10505 1965 10545 1970
rect 10615 1970 10620 1975
rect 10650 1995 10655 2000
rect 10725 2000 10765 2005
rect 10725 1995 10730 2000
rect 10650 1975 10730 1995
rect 10650 1970 10655 1975
rect 10615 1965 10655 1970
rect 10725 1970 10730 1975
rect 10760 1995 10765 2000
rect 10835 2000 10875 2005
rect 10835 1995 10840 2000
rect 10760 1975 10840 1995
rect 10760 1970 10765 1975
rect 10725 1965 10765 1970
rect 10835 1970 10840 1975
rect 10870 1970 10875 2000
rect 10835 1965 10875 1970
rect 12945 2000 12985 2005
rect 12945 1970 12950 2000
rect 12980 1995 12985 2000
rect 13055 2000 13095 2005
rect 13055 1995 13060 2000
rect 12980 1975 13060 1995
rect 12980 1970 12985 1975
rect 12945 1965 12985 1970
rect 13055 1970 13060 1975
rect 13090 1995 13095 2000
rect 13165 2000 13205 2005
rect 13165 1995 13170 2000
rect 13090 1975 13170 1995
rect 13090 1970 13095 1975
rect 13055 1965 13095 1970
rect 13165 1970 13170 1975
rect 13200 1995 13205 2000
rect 13275 2000 13315 2005
rect 13275 1995 13280 2000
rect 13200 1975 13280 1995
rect 13200 1970 13205 1975
rect 13165 1965 13205 1970
rect 13275 1970 13280 1975
rect 13310 1995 13315 2000
rect 13385 2000 13425 2005
rect 13385 1995 13390 2000
rect 13310 1975 13390 1995
rect 13310 1970 13315 1975
rect 13275 1965 13315 1970
rect 13385 1970 13390 1975
rect 13420 1995 13425 2000
rect 13495 2000 13535 2005
rect 13495 1995 13500 2000
rect 13420 1975 13500 1995
rect 13420 1970 13425 1975
rect 13385 1965 13425 1970
rect 13495 1970 13500 1975
rect 13530 1995 13535 2000
rect 13605 2000 13645 2005
rect 13605 1995 13610 2000
rect 13530 1975 13610 1995
rect 13530 1970 13535 1975
rect 13495 1965 13535 1970
rect 13605 1970 13610 1975
rect 13640 1995 13645 2000
rect 13715 2000 13755 2005
rect 13715 1995 13720 2000
rect 13640 1975 13720 1995
rect 13640 1970 13645 1975
rect 13605 1965 13645 1970
rect 13715 1970 13720 1975
rect 13750 1995 13755 2000
rect 13825 2000 13865 2005
rect 13825 1995 13830 2000
rect 13750 1975 13830 1995
rect 13750 1970 13755 1975
rect 13715 1965 13755 1970
rect 13825 1970 13830 1975
rect 13860 1995 13865 2000
rect 13935 2000 13975 2005
rect 13935 1995 13940 2000
rect 13860 1975 13940 1995
rect 13860 1970 13865 1975
rect 13825 1965 13865 1970
rect 13935 1970 13940 1975
rect 13970 1995 13975 2000
rect 14045 2000 14085 2005
rect 14045 1995 14050 2000
rect 13970 1975 14050 1995
rect 13970 1970 13975 1975
rect 13935 1965 13975 1970
rect 14045 1970 14050 1975
rect 14080 1970 14085 2000
rect 14045 1965 14085 1970
rect 17235 2000 17275 2005
rect 17235 1970 17240 2000
rect 17270 1995 17275 2000
rect 17345 2000 17385 2005
rect 17345 1995 17350 2000
rect 17270 1975 17350 1995
rect 17270 1970 17275 1975
rect 17235 1965 17275 1970
rect 17345 1970 17350 1975
rect 17380 1995 17385 2000
rect 17455 2000 17495 2005
rect 17455 1995 17460 2000
rect 17380 1975 17460 1995
rect 17380 1970 17385 1975
rect 17345 1965 17385 1970
rect 17455 1970 17460 1975
rect 17490 1995 17495 2000
rect 17565 2000 17605 2005
rect 17565 1995 17570 2000
rect 17490 1975 17570 1995
rect 17490 1970 17495 1975
rect 17455 1965 17495 1970
rect 17565 1970 17570 1975
rect 17600 1995 17605 2000
rect 17675 2000 17715 2005
rect 17675 1995 17680 2000
rect 17600 1975 17680 1995
rect 17600 1970 17605 1975
rect 17565 1965 17605 1970
rect 17675 1970 17680 1975
rect 17710 1995 17715 2000
rect 17785 2000 17825 2005
rect 17785 1995 17790 2000
rect 17710 1975 17790 1995
rect 17710 1970 17715 1975
rect 17675 1965 17715 1970
rect 17785 1970 17790 1975
rect 17820 1995 17825 2000
rect 17895 2000 17935 2005
rect 17895 1995 17900 2000
rect 17820 1975 17900 1995
rect 17820 1970 17825 1975
rect 17785 1965 17825 1970
rect 17895 1970 17900 1975
rect 17930 1995 17935 2000
rect 18005 2000 18045 2005
rect 18005 1995 18010 2000
rect 17930 1975 18010 1995
rect 17930 1970 17935 1975
rect 17895 1965 17935 1970
rect 18005 1970 18010 1975
rect 18040 1995 18045 2000
rect 18115 2000 18155 2005
rect 18115 1995 18120 2000
rect 18040 1975 18120 1995
rect 18040 1970 18045 1975
rect 18005 1965 18045 1970
rect 18115 1970 18120 1975
rect 18150 1995 18155 2000
rect 18225 2000 18265 2005
rect 18225 1995 18230 2000
rect 18150 1975 18230 1995
rect 18150 1970 18155 1975
rect 18115 1965 18155 1970
rect 18225 1970 18230 1975
rect 18260 1995 18265 2000
rect 18335 2000 18375 2005
rect 18335 1995 18340 2000
rect 18260 1975 18340 1995
rect 18260 1970 18265 1975
rect 18225 1965 18265 1970
rect 18335 1970 18340 1975
rect 18370 1970 18375 2000
rect 18335 1965 18375 1970
rect 20445 2000 20485 2005
rect 20445 1970 20450 2000
rect 20480 1995 20485 2000
rect 20555 2000 20595 2005
rect 20555 1995 20560 2000
rect 20480 1975 20560 1995
rect 20480 1970 20485 1975
rect 20445 1965 20485 1970
rect 20555 1970 20560 1975
rect 20590 1995 20595 2000
rect 20665 2000 20705 2005
rect 20665 1995 20670 2000
rect 20590 1975 20670 1995
rect 20590 1970 20595 1975
rect 20555 1965 20595 1970
rect 20665 1970 20670 1975
rect 20700 1995 20705 2000
rect 20775 2000 20815 2005
rect 20775 1995 20780 2000
rect 20700 1975 20780 1995
rect 20700 1970 20705 1975
rect 20665 1965 20705 1970
rect 20775 1970 20780 1975
rect 20810 1995 20815 2000
rect 20885 2000 20925 2005
rect 20885 1995 20890 2000
rect 20810 1975 20890 1995
rect 20810 1970 20815 1975
rect 20775 1965 20815 1970
rect 20885 1970 20890 1975
rect 20920 1995 20925 2000
rect 20995 2000 21035 2005
rect 20995 1995 21000 2000
rect 20920 1975 21000 1995
rect 20920 1970 20925 1975
rect 20885 1965 20925 1970
rect 20995 1970 21000 1975
rect 21030 1995 21035 2000
rect 21105 2000 21145 2005
rect 21105 1995 21110 2000
rect 21030 1975 21110 1995
rect 21030 1970 21035 1975
rect 20995 1965 21035 1970
rect 21105 1970 21110 1975
rect 21140 1995 21145 2000
rect 21215 2000 21255 2005
rect 21215 1995 21220 2000
rect 21140 1975 21220 1995
rect 21140 1970 21145 1975
rect 21105 1965 21145 1970
rect 21215 1970 21220 1975
rect 21250 1995 21255 2000
rect 21325 2000 21365 2005
rect 21325 1995 21330 2000
rect 21250 1975 21330 1995
rect 21250 1970 21255 1975
rect 21215 1965 21255 1970
rect 21325 1970 21330 1975
rect 21360 1995 21365 2000
rect 21435 2000 21475 2005
rect 21435 1995 21440 2000
rect 21360 1975 21440 1995
rect 21360 1970 21365 1975
rect 21325 1965 21365 1970
rect 21435 1970 21440 1975
rect 21470 1995 21475 2000
rect 21545 2000 21585 2005
rect 21545 1995 21550 2000
rect 21470 1975 21550 1995
rect 21470 1970 21475 1975
rect 21435 1965 21475 1970
rect 21545 1970 21550 1975
rect 21580 1970 21585 2000
rect 21545 1965 21585 1970
rect 11385 1960 11425 1965
rect 11385 1930 11390 1960
rect 11420 1955 11425 1960
rect 11605 1960 11645 1965
rect 11605 1955 11610 1960
rect 11420 1935 11610 1955
rect 11420 1930 11425 1935
rect 11385 1925 11425 1930
rect 11605 1930 11610 1935
rect 11640 1955 11645 1960
rect 11825 1960 11865 1965
rect 11825 1955 11830 1960
rect 11640 1935 11830 1955
rect 11640 1930 11645 1935
rect 11605 1925 11645 1930
rect 11825 1930 11830 1935
rect 11860 1955 11865 1960
rect 12045 1960 12085 1965
rect 12045 1955 12050 1960
rect 11860 1935 12050 1955
rect 11860 1930 11865 1935
rect 11825 1925 11865 1930
rect 12045 1930 12050 1935
rect 12080 1955 12085 1960
rect 12265 1960 12305 1965
rect 12265 1955 12270 1960
rect 12080 1935 12270 1955
rect 12080 1930 12085 1935
rect 12045 1925 12085 1930
rect 12265 1930 12270 1935
rect 12300 1930 12305 1960
rect 12265 1925 12305 1930
rect 18885 1960 18925 1965
rect 18885 1930 18890 1960
rect 18920 1955 18925 1960
rect 19105 1960 19145 1965
rect 19105 1955 19110 1960
rect 18920 1935 19110 1955
rect 18920 1930 18925 1935
rect 18885 1925 18925 1930
rect 19105 1930 19110 1935
rect 19140 1955 19145 1960
rect 19325 1960 19365 1965
rect 19325 1955 19330 1960
rect 19140 1935 19330 1955
rect 19140 1930 19145 1935
rect 19105 1925 19145 1930
rect 19325 1930 19330 1935
rect 19360 1955 19365 1960
rect 19545 1960 19585 1965
rect 19545 1955 19550 1960
rect 19360 1935 19550 1955
rect 19360 1930 19365 1935
rect 19325 1925 19365 1930
rect 19545 1930 19550 1935
rect 19580 1955 19585 1960
rect 19765 1960 19805 1965
rect 19765 1955 19770 1960
rect 19580 1935 19770 1955
rect 19580 1930 19585 1935
rect 19545 1925 19585 1930
rect 19765 1930 19770 1935
rect 19800 1930 19805 1960
rect 19765 1925 19805 1930
rect 11495 1905 11535 1910
rect 2925 1880 2965 1885
rect 2925 1850 2930 1880
rect 2960 1875 2965 1880
rect 3045 1875 3085 1885
rect 3285 1880 3325 1885
rect 3285 1875 3290 1880
rect 2960 1855 3290 1875
rect 2960 1850 2965 1855
rect 2925 1845 2965 1850
rect 3045 1845 3085 1855
rect 3285 1850 3290 1855
rect 3320 1875 3325 1880
rect 3405 1875 3445 1885
rect 3645 1880 3685 1885
rect 3645 1875 3650 1880
rect 3320 1855 3650 1875
rect 3320 1850 3325 1855
rect 3285 1845 3325 1850
rect 3405 1845 3445 1855
rect 3645 1850 3650 1855
rect 3680 1850 3685 1880
rect 3645 1845 3685 1850
rect 3765 1845 3805 1885
rect 4205 1845 4245 1885
rect 4325 1880 4365 1885
rect 4325 1850 4330 1880
rect 4360 1875 4365 1880
rect 4565 1875 4605 1885
rect 4685 1880 4725 1885
rect 4685 1875 4690 1880
rect 4360 1855 4690 1875
rect 4360 1850 4365 1855
rect 4325 1845 4365 1850
rect 4565 1845 4605 1855
rect 4685 1850 4690 1855
rect 4720 1875 4725 1880
rect 4925 1875 4965 1885
rect 5045 1880 5085 1885
rect 5045 1875 5050 1880
rect 4720 1855 5050 1875
rect 4720 1850 4725 1855
rect 4685 1845 4725 1850
rect 4925 1845 4965 1855
rect 5045 1850 5050 1855
rect 5080 1875 5085 1880
rect 11495 1875 11500 1905
rect 11530 1900 11535 1905
rect 11715 1905 11755 1910
rect 11715 1900 11720 1905
rect 11530 1880 11720 1900
rect 11530 1875 11535 1880
rect 5080 1855 5175 1875
rect 11495 1870 11535 1875
rect 11715 1875 11720 1880
rect 11750 1900 11755 1905
rect 11935 1905 11975 1910
rect 11935 1900 11940 1905
rect 11750 1880 11940 1900
rect 11750 1875 11755 1880
rect 11715 1870 11755 1875
rect 11935 1875 11940 1880
rect 11970 1900 11975 1905
rect 12155 1905 12195 1910
rect 12155 1900 12160 1905
rect 11970 1880 12160 1900
rect 11970 1875 11975 1880
rect 11935 1870 11975 1875
rect 12155 1875 12160 1880
rect 12190 1900 12195 1905
rect 12375 1905 12415 1910
rect 12375 1900 12380 1905
rect 12190 1880 12380 1900
rect 12190 1875 12195 1880
rect 12155 1870 12195 1875
rect 12375 1875 12380 1880
rect 12410 1875 12415 1905
rect 12375 1870 12415 1875
rect 18995 1905 19035 1910
rect 18995 1875 19000 1905
rect 19030 1900 19035 1905
rect 19215 1905 19255 1910
rect 19215 1900 19220 1905
rect 19030 1880 19220 1900
rect 19030 1875 19035 1880
rect 18995 1870 19035 1875
rect 19215 1875 19220 1880
rect 19250 1900 19255 1905
rect 19435 1905 19475 1910
rect 19435 1900 19440 1905
rect 19250 1880 19440 1900
rect 19250 1875 19255 1880
rect 19215 1870 19255 1875
rect 19435 1875 19440 1880
rect 19470 1900 19475 1905
rect 19655 1905 19695 1910
rect 19655 1900 19660 1905
rect 19470 1880 19660 1900
rect 19470 1875 19475 1880
rect 19435 1870 19475 1875
rect 19655 1875 19660 1880
rect 19690 1900 19695 1905
rect 19875 1905 19915 1910
rect 19875 1900 19880 1905
rect 19690 1880 19880 1900
rect 19690 1875 19695 1880
rect 19655 1870 19695 1875
rect 19875 1875 19880 1880
rect 19910 1875 19915 1905
rect 19875 1870 19915 1875
rect 20545 1905 20585 1910
rect 20545 1875 20550 1905
rect 20580 1900 20585 1905
rect 20655 1905 20695 1910
rect 20655 1900 20660 1905
rect 20580 1880 20660 1900
rect 20580 1875 20585 1880
rect 20545 1870 20585 1875
rect 20655 1875 20660 1880
rect 20690 1900 20695 1905
rect 20765 1905 20805 1910
rect 20765 1900 20770 1905
rect 20690 1880 20770 1900
rect 20690 1875 20695 1880
rect 20655 1870 20695 1875
rect 20765 1875 20770 1880
rect 20800 1875 20805 1905
rect 20765 1870 20805 1875
rect 5080 1850 5085 1855
rect 5045 1845 5085 1850
rect 11190 1850 11230 1855
rect 2470 1820 2510 1825
rect 2470 1790 2475 1820
rect 2505 1815 2510 1820
rect 2835 1820 2875 1825
rect 2835 1815 2840 1820
rect 2505 1795 2840 1815
rect 2505 1790 2510 1795
rect 2470 1785 2510 1790
rect 2835 1790 2840 1795
rect 2870 1815 2875 1820
rect 3045 1820 3085 1825
rect 3045 1815 3050 1820
rect 2870 1795 3050 1815
rect 2870 1790 2875 1795
rect 2835 1785 2875 1790
rect 3045 1790 3050 1795
rect 3080 1815 3085 1820
rect 3165 1820 3205 1825
rect 3165 1815 3170 1820
rect 3080 1795 3170 1815
rect 3080 1790 3085 1795
rect 3045 1785 3085 1790
rect 3165 1790 3170 1795
rect 3200 1815 3205 1820
rect 3405 1820 3445 1825
rect 3405 1815 3410 1820
rect 3200 1795 3410 1815
rect 3200 1790 3205 1795
rect 3165 1785 3205 1790
rect 3405 1790 3410 1795
rect 3440 1815 3445 1820
rect 3525 1820 3565 1825
rect 3525 1815 3530 1820
rect 3440 1795 3530 1815
rect 3440 1790 3445 1795
rect 3405 1785 3445 1790
rect 3525 1790 3530 1795
rect 3560 1815 3565 1820
rect 3765 1820 3805 1825
rect 3765 1815 3770 1820
rect 3560 1795 3770 1815
rect 3560 1790 3565 1795
rect 3525 1785 3565 1790
rect 3765 1790 3770 1795
rect 3800 1815 3805 1820
rect 3855 1820 3895 1825
rect 3855 1815 3860 1820
rect 3800 1795 3860 1815
rect 3800 1790 3805 1795
rect 3765 1785 3805 1790
rect 3855 1790 3860 1795
rect 3890 1790 3895 1820
rect 3855 1785 3895 1790
rect 4115 1820 4155 1825
rect 4115 1790 4120 1820
rect 4150 1815 4155 1820
rect 4205 1820 4245 1825
rect 4205 1815 4210 1820
rect 4150 1795 4210 1815
rect 4150 1790 4155 1795
rect 4115 1785 4155 1790
rect 4205 1790 4210 1795
rect 4240 1815 4245 1820
rect 4445 1820 4485 1825
rect 4445 1815 4450 1820
rect 4240 1795 4450 1815
rect 4240 1790 4245 1795
rect 4205 1785 4245 1790
rect 4445 1790 4450 1795
rect 4480 1815 4485 1820
rect 4565 1820 4605 1825
rect 4565 1815 4570 1820
rect 4480 1795 4570 1815
rect 4480 1790 4485 1795
rect 4445 1785 4485 1790
rect 4565 1790 4570 1795
rect 4600 1815 4605 1820
rect 4805 1820 4845 1825
rect 4805 1815 4810 1820
rect 4600 1795 4810 1815
rect 4600 1790 4605 1795
rect 4565 1785 4605 1790
rect 4805 1790 4810 1795
rect 4840 1815 4845 1820
rect 4925 1820 4965 1825
rect 4925 1815 4930 1820
rect 4840 1795 4930 1815
rect 4840 1790 4845 1795
rect 4805 1785 4845 1790
rect 4925 1790 4930 1795
rect 4960 1815 4965 1820
rect 5135 1820 5175 1825
rect 5135 1815 5140 1820
rect 4960 1795 5140 1815
rect 4960 1790 4965 1795
rect 4925 1785 4965 1790
rect 5135 1790 5140 1795
rect 5170 1815 5175 1820
rect 5360 1820 5400 1825
rect 5360 1815 5365 1820
rect 5170 1795 5365 1815
rect 5170 1790 5175 1795
rect 5135 1785 5175 1790
rect 5360 1790 5365 1795
rect 5395 1790 5400 1820
rect 11190 1820 11195 1850
rect 11225 1845 11230 1850
rect 11410 1850 11450 1855
rect 11410 1845 11415 1850
rect 11225 1825 11415 1845
rect 11225 1820 11230 1825
rect 11190 1815 11230 1820
rect 11410 1820 11415 1825
rect 11445 1845 11450 1850
rect 11640 1850 11680 1855
rect 11640 1845 11645 1850
rect 11445 1825 11645 1845
rect 11445 1820 11450 1825
rect 11410 1815 11450 1820
rect 11640 1820 11645 1825
rect 11675 1845 11680 1850
rect 12230 1850 12270 1855
rect 12230 1845 12235 1850
rect 11675 1825 12235 1845
rect 11675 1820 11680 1825
rect 11640 1815 11680 1820
rect 12230 1820 12235 1825
rect 12265 1845 12270 1850
rect 12450 1850 12490 1855
rect 12450 1845 12455 1850
rect 12265 1825 12455 1845
rect 12265 1820 12270 1825
rect 12230 1815 12270 1820
rect 12450 1820 12455 1825
rect 12485 1845 12490 1850
rect 12680 1850 12720 1855
rect 12680 1845 12685 1850
rect 12485 1825 12685 1845
rect 12485 1820 12490 1825
rect 12450 1815 12490 1820
rect 12680 1820 12685 1825
rect 12715 1820 12720 1850
rect 12680 1815 12720 1820
rect 18690 1850 18730 1855
rect 18690 1820 18695 1850
rect 18725 1845 18730 1850
rect 18910 1850 18950 1855
rect 18910 1845 18915 1850
rect 18725 1825 18915 1845
rect 18725 1820 18730 1825
rect 18690 1815 18730 1820
rect 18910 1820 18915 1825
rect 18945 1845 18950 1850
rect 19140 1850 19180 1855
rect 19140 1845 19145 1850
rect 18945 1825 19145 1845
rect 18945 1820 18950 1825
rect 18910 1815 18950 1820
rect 19140 1820 19145 1825
rect 19175 1845 19180 1850
rect 19730 1850 19770 1855
rect 19730 1845 19735 1850
rect 19175 1825 19735 1845
rect 19175 1820 19180 1825
rect 19140 1815 19180 1820
rect 19730 1820 19735 1825
rect 19765 1845 19770 1850
rect 19950 1850 19990 1855
rect 19950 1845 19955 1850
rect 19765 1825 19955 1845
rect 19765 1820 19770 1825
rect 19730 1815 19770 1820
rect 19950 1820 19955 1825
rect 19985 1845 19990 1850
rect 20180 1850 20220 1855
rect 20180 1845 20185 1850
rect 19985 1825 20185 1845
rect 19985 1820 19990 1825
rect 19950 1815 19990 1820
rect 20180 1820 20185 1825
rect 20215 1820 20220 1850
rect 20180 1815 20220 1820
rect 5360 1785 5400 1790
rect 11820 1805 11860 1810
rect 11820 1775 11825 1805
rect 11855 1800 11860 1805
rect 11940 1805 11980 1810
rect 11940 1800 11945 1805
rect 11855 1780 11945 1800
rect 11855 1775 11860 1780
rect 11820 1770 11860 1775
rect 11940 1775 11945 1780
rect 11975 1775 11980 1805
rect 11940 1770 11980 1775
rect 19320 1805 19360 1810
rect 19320 1775 19325 1805
rect 19355 1800 19360 1805
rect 19440 1805 19480 1810
rect 19440 1800 19445 1805
rect 19355 1780 19445 1800
rect 19355 1775 19360 1780
rect 19320 1770 19360 1775
rect 19440 1775 19445 1780
rect 19475 1775 19480 1805
rect 19440 1770 19480 1775
rect 2800 1765 2840 1770
rect 2425 1760 2465 1765
rect 2425 1730 2430 1760
rect 2460 1755 2465 1760
rect 2565 1760 2605 1765
rect 2565 1755 2570 1760
rect 2460 1735 2570 1755
rect 2460 1730 2465 1735
rect 2425 1725 2465 1730
rect 2565 1730 2570 1735
rect 2600 1755 2605 1760
rect 2675 1760 2715 1765
rect 2675 1755 2680 1760
rect 2600 1735 2680 1755
rect 2600 1730 2605 1735
rect 2565 1725 2605 1730
rect 2675 1730 2680 1735
rect 2710 1755 2715 1760
rect 2800 1755 2805 1765
rect 2710 1735 2805 1755
rect 2835 1755 2840 1765
rect 3225 1760 3265 1765
rect 3225 1755 3230 1760
rect 2835 1735 3230 1755
rect 2710 1730 2715 1735
rect 2800 1730 2840 1735
rect 3225 1730 3230 1735
rect 3260 1730 3265 1760
rect 2675 1725 2715 1730
rect 3225 1725 3265 1730
rect 3285 1760 3325 1765
rect 3285 1730 3290 1760
rect 3320 1755 3325 1760
rect 3525 1760 3565 1765
rect 3525 1755 3530 1760
rect 3320 1735 3530 1755
rect 3320 1730 3325 1735
rect 3285 1725 3325 1730
rect 3525 1730 3530 1735
rect 3560 1755 3565 1760
rect 3765 1760 3805 1765
rect 3765 1755 3770 1760
rect 3560 1735 3770 1755
rect 3560 1730 3565 1735
rect 3525 1725 3565 1730
rect 3765 1730 3770 1735
rect 3800 1730 3805 1760
rect 3765 1725 3805 1730
rect 4205 1760 4245 1765
rect 4205 1730 4210 1760
rect 4240 1755 4245 1760
rect 4445 1760 4485 1765
rect 4445 1755 4450 1760
rect 4240 1735 4450 1755
rect 4240 1730 4245 1735
rect 4205 1725 4245 1730
rect 4445 1730 4450 1735
rect 4480 1755 4485 1760
rect 4685 1760 4725 1765
rect 4685 1755 4690 1760
rect 4480 1735 4690 1755
rect 4480 1730 4485 1735
rect 4445 1725 4485 1730
rect 4685 1730 4690 1735
rect 4720 1730 4725 1760
rect 4685 1725 4725 1730
rect 4745 1760 4785 1765
rect 4745 1730 4750 1760
rect 4780 1755 4785 1760
rect 5270 1760 5310 1765
rect 5270 1755 5275 1760
rect 4780 1735 5275 1755
rect 4780 1730 4785 1735
rect 4745 1725 4785 1730
rect 5270 1730 5275 1735
rect 5305 1755 5310 1760
rect 11085 1760 11125 1765
rect 5305 1735 6100 1755
rect 5305 1730 5310 1735
rect 5270 1725 5310 1730
rect 11085 1730 11090 1760
rect 11120 1755 11125 1760
rect 11305 1760 11345 1765
rect 11305 1755 11310 1760
rect 11120 1735 11310 1755
rect 11120 1730 11125 1735
rect 11085 1725 11125 1730
rect 11305 1730 11310 1735
rect 11340 1755 11345 1760
rect 11525 1760 11565 1765
rect 11525 1755 11530 1760
rect 11340 1735 11530 1755
rect 11340 1730 11345 1735
rect 11305 1725 11345 1730
rect 11525 1730 11530 1735
rect 11560 1755 11565 1760
rect 12125 1760 12165 1765
rect 12125 1755 12130 1760
rect 11560 1735 12130 1755
rect 11560 1730 11565 1735
rect 11525 1725 11565 1730
rect 12125 1730 12130 1735
rect 12160 1755 12165 1760
rect 12345 1760 12385 1765
rect 12345 1755 12350 1760
rect 12160 1735 12350 1755
rect 12160 1730 12165 1735
rect 12125 1725 12165 1730
rect 12345 1730 12350 1735
rect 12380 1755 12385 1760
rect 12565 1760 12605 1765
rect 12565 1755 12570 1760
rect 12380 1735 12570 1755
rect 12380 1730 12385 1735
rect 12345 1725 12385 1730
rect 12565 1730 12570 1735
rect 12600 1730 12605 1760
rect 12565 1725 12605 1730
rect 18585 1760 18625 1765
rect 18585 1730 18590 1760
rect 18620 1755 18625 1760
rect 18805 1760 18845 1765
rect 18805 1755 18810 1760
rect 18620 1735 18810 1755
rect 18620 1730 18625 1735
rect 18585 1725 18625 1730
rect 18805 1730 18810 1735
rect 18840 1755 18845 1760
rect 19025 1760 19065 1765
rect 19025 1755 19030 1760
rect 18840 1735 19030 1755
rect 18840 1730 18845 1735
rect 18805 1725 18845 1730
rect 19025 1730 19030 1735
rect 19060 1755 19065 1760
rect 19625 1760 19665 1765
rect 19625 1755 19630 1760
rect 19060 1735 19630 1755
rect 19060 1730 19065 1735
rect 19025 1725 19065 1730
rect 19625 1730 19630 1735
rect 19660 1755 19665 1760
rect 19845 1760 19885 1765
rect 19845 1755 19850 1760
rect 19660 1735 19850 1755
rect 19660 1730 19665 1735
rect 19625 1725 19665 1730
rect 19845 1730 19850 1735
rect 19880 1755 19885 1760
rect 20065 1760 20105 1765
rect 20065 1755 20070 1760
rect 19880 1735 20070 1755
rect 19880 1730 19885 1735
rect 19845 1725 19885 1730
rect 20065 1730 20070 1735
rect 20100 1730 20105 1760
rect 20065 1725 20105 1730
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 1685 -70 1690
rect -45 1720 -5 1725
rect -45 1690 -40 1720
rect -10 1690 -5 1720
rect 3165 1715 3205 1720
rect -45 1685 -5 1690
rect 1262 1710 1302 1715
rect 1262 1680 1270 1710
rect 1297 1705 1302 1710
rect 2800 1710 2840 1715
rect 2800 1705 2805 1710
rect 1297 1685 2805 1705
rect 1297 1680 1302 1685
rect 1262 1675 1302 1680
rect 2800 1680 2805 1685
rect 2835 1680 2840 1710
rect 3165 1685 3170 1715
rect 3200 1710 3205 1715
rect 3405 1715 3445 1720
rect 3405 1710 3410 1715
rect 3200 1690 3410 1710
rect 3200 1685 3205 1690
rect 3165 1680 3205 1685
rect 3405 1685 3410 1690
rect 3440 1710 3445 1715
rect 3645 1715 3685 1720
rect 3645 1710 3650 1715
rect 3440 1690 3650 1710
rect 3440 1685 3445 1690
rect 3405 1680 3445 1685
rect 3645 1685 3650 1690
rect 3680 1685 3685 1715
rect 3645 1680 3685 1685
rect 4325 1715 4365 1720
rect 4325 1685 4330 1715
rect 4360 1710 4365 1715
rect 4565 1715 4605 1720
rect 4565 1710 4570 1715
rect 4360 1690 4570 1710
rect 4360 1685 4365 1690
rect 4325 1680 4365 1685
rect 4565 1685 4570 1690
rect 4600 1710 4605 1715
rect 4805 1715 4845 1720
rect 4805 1710 4810 1715
rect 4600 1690 4810 1710
rect 4600 1685 4605 1690
rect 4565 1680 4605 1685
rect 4805 1685 4810 1690
rect 4840 1685 4845 1715
rect 11237 1715 11269 1720
rect 11237 1710 11240 1715
rect 10910 1690 11240 1710
rect 4805 1680 4845 1685
rect 11237 1685 11240 1690
rect 11266 1710 11269 1715
rect 11457 1715 11489 1720
rect 11457 1710 11460 1715
rect 11266 1690 11460 1710
rect 11266 1685 11269 1690
rect 11237 1680 11269 1685
rect 11457 1685 11460 1690
rect 11486 1710 11489 1715
rect 11601 1715 11633 1720
rect 11601 1710 11604 1715
rect 11486 1690 11604 1710
rect 11486 1685 11489 1690
rect 11457 1680 11489 1685
rect 11601 1685 11604 1690
rect 11630 1710 11633 1715
rect 11867 1715 11899 1720
rect 11867 1710 11870 1715
rect 11630 1690 11870 1710
rect 11630 1685 11633 1690
rect 11601 1680 11633 1685
rect 11867 1685 11870 1690
rect 11896 1710 11899 1715
rect 12277 1715 12309 1720
rect 12277 1710 12280 1715
rect 11896 1690 12280 1710
rect 11896 1685 11899 1690
rect 11867 1680 11899 1685
rect 12277 1685 12280 1690
rect 12306 1710 12309 1715
rect 12497 1715 12529 1720
rect 12497 1710 12500 1715
rect 12306 1690 12500 1710
rect 12306 1685 12309 1690
rect 12277 1680 12309 1685
rect 12497 1685 12500 1690
rect 12526 1710 12529 1715
rect 12641 1715 12673 1720
rect 12641 1710 12644 1715
rect 12526 1690 12644 1710
rect 12526 1685 12529 1690
rect 12497 1680 12529 1685
rect 12641 1685 12644 1690
rect 12670 1685 12673 1715
rect 18737 1715 18769 1720
rect 18737 1710 18740 1715
rect 18410 1690 18740 1710
rect 12641 1680 12673 1685
rect 18737 1685 18740 1690
rect 18766 1710 18769 1715
rect 18957 1715 18989 1720
rect 18957 1710 18960 1715
rect 18766 1690 18960 1710
rect 18766 1685 18769 1690
rect 18737 1680 18769 1685
rect 18957 1685 18960 1690
rect 18986 1710 18989 1715
rect 19101 1715 19133 1720
rect 19101 1710 19104 1715
rect 18986 1690 19104 1710
rect 18986 1685 18989 1690
rect 18957 1680 18989 1685
rect 19101 1685 19104 1690
rect 19130 1710 19133 1715
rect 19367 1715 19399 1720
rect 19367 1710 19370 1715
rect 19130 1690 19370 1710
rect 19130 1685 19133 1690
rect 19101 1680 19133 1685
rect 19367 1685 19370 1690
rect 19396 1710 19399 1715
rect 19777 1715 19809 1720
rect 19777 1710 19780 1715
rect 19396 1690 19780 1710
rect 19396 1685 19399 1690
rect 19367 1680 19399 1685
rect 19777 1685 19780 1690
rect 19806 1710 19809 1715
rect 19997 1715 20029 1720
rect 19997 1710 20000 1715
rect 19806 1690 20000 1710
rect 19806 1685 19809 1690
rect 19777 1680 19809 1685
rect 19997 1685 20000 1690
rect 20026 1710 20029 1715
rect 20141 1715 20173 1720
rect 20141 1710 20144 1715
rect 20026 1690 20144 1710
rect 20026 1685 20029 1690
rect 19997 1680 20029 1685
rect 20141 1685 20144 1690
rect 20170 1685 20173 1715
rect 20141 1680 20173 1685
rect 20566 1680 20598 1685
rect 2800 1675 2840 1680
rect 2380 1665 2420 1670
rect 2380 1635 2385 1665
rect 2415 1660 2420 1665
rect 2620 1665 2660 1670
rect 2620 1660 2625 1665
rect 2415 1640 2625 1660
rect 2415 1635 2420 1640
rect 2380 1630 2420 1635
rect 2620 1635 2625 1640
rect 2655 1635 2660 1665
rect 20566 1650 20570 1680
rect 20596 1650 20598 1680
rect 20566 1645 20598 1650
rect 2620 1630 2660 1635
rect 20510 1630 20550 1635
rect 20510 1600 20515 1630
rect 20545 1625 20550 1630
rect 20616 1630 20656 1635
rect 20616 1625 20621 1630
rect 20545 1605 20621 1625
rect 20545 1600 20550 1605
rect 2330 1595 2370 1600
rect 2330 1565 2335 1595
rect 2365 1590 2370 1595
rect 3165 1595 3205 1600
rect 3165 1590 3170 1595
rect 2365 1570 3170 1590
rect 2365 1565 2370 1570
rect 2330 1560 2370 1565
rect 3165 1565 3170 1570
rect 3200 1565 3205 1595
rect 3165 1560 3205 1565
rect 4805 1595 4845 1600
rect 4805 1565 4810 1595
rect 4840 1590 4845 1595
rect 5410 1595 5450 1600
rect 20510 1595 20550 1600
rect 20616 1600 20621 1605
rect 20651 1600 20656 1630
rect 20616 1595 20656 1600
rect 20710 1630 20750 1635
rect 20710 1600 20715 1630
rect 20745 1625 20750 1630
rect 20800 1630 20840 1635
rect 20800 1625 20805 1630
rect 20745 1605 20805 1625
rect 20745 1600 20750 1605
rect 20710 1595 20750 1600
rect 20800 1600 20805 1605
rect 20835 1600 20840 1630
rect 20800 1595 20840 1600
rect 5410 1590 5415 1595
rect 4840 1570 5415 1590
rect 4840 1565 4845 1570
rect 4805 1560 4845 1565
rect 5410 1565 5415 1570
rect 5445 1565 5450 1595
rect 5410 1560 5450 1565
rect 12815 1570 12855 1575
rect 2835 1545 2875 1550
rect 2835 1515 2840 1545
rect 2870 1540 2875 1545
rect 3225 1545 3265 1550
rect 3225 1540 3230 1545
rect 2870 1520 3230 1540
rect 2870 1515 2875 1520
rect 2835 1510 2875 1515
rect 3225 1515 3230 1520
rect 3260 1540 3265 1545
rect 3345 1545 3385 1550
rect 3345 1540 3350 1545
rect 3260 1520 3350 1540
rect 3260 1515 3265 1520
rect 3225 1510 3265 1515
rect 3345 1515 3350 1520
rect 3380 1540 3385 1545
rect 3465 1545 3505 1550
rect 3465 1540 3470 1545
rect 3380 1520 3470 1540
rect 3380 1515 3385 1520
rect 3345 1510 3385 1515
rect 3465 1515 3470 1520
rect 3500 1540 3505 1545
rect 3585 1545 3625 1550
rect 3585 1540 3590 1545
rect 3500 1520 3590 1540
rect 3500 1515 3505 1520
rect 3465 1510 3505 1515
rect 3585 1515 3590 1520
rect 3620 1540 3625 1545
rect 3705 1545 3745 1550
rect 3705 1540 3710 1545
rect 3620 1520 3710 1540
rect 3620 1515 3625 1520
rect 3585 1510 3625 1515
rect 3705 1515 3710 1520
rect 3740 1515 3745 1545
rect 3705 1510 3745 1515
rect 4265 1545 4305 1550
rect 4265 1515 4270 1545
rect 4300 1540 4305 1545
rect 4385 1545 4425 1550
rect 4385 1540 4390 1545
rect 4300 1520 4390 1540
rect 4300 1515 4305 1520
rect 4265 1510 4305 1515
rect 4385 1515 4390 1520
rect 4420 1540 4425 1545
rect 4505 1545 4545 1550
rect 4505 1540 4510 1545
rect 4420 1520 4510 1540
rect 4420 1515 4425 1520
rect 4385 1510 4425 1515
rect 4505 1515 4510 1520
rect 4540 1540 4545 1545
rect 4625 1545 4665 1550
rect 4625 1540 4630 1545
rect 4540 1520 4630 1540
rect 4540 1515 4545 1520
rect 4505 1510 4545 1515
rect 4625 1515 4630 1520
rect 4660 1540 4665 1545
rect 4745 1545 4785 1550
rect 4745 1540 4750 1545
rect 4660 1520 4750 1540
rect 4660 1515 4665 1520
rect 4625 1510 4665 1515
rect 4745 1515 4750 1520
rect 4780 1540 4785 1545
rect 5135 1545 5175 1550
rect 5135 1540 5140 1545
rect 4780 1520 5140 1540
rect 4780 1515 4785 1520
rect 4745 1510 4785 1515
rect 5135 1515 5140 1520
rect 5170 1515 5175 1545
rect 12815 1540 12820 1570
rect 12850 1540 12855 1570
rect 12815 1535 12855 1540
rect 20315 1570 20355 1575
rect 20315 1540 20320 1570
rect 20350 1565 20355 1570
rect 20471 1570 20503 1575
rect 20471 1565 20475 1570
rect 20350 1545 20475 1565
rect 20350 1540 20355 1545
rect 20315 1535 20355 1540
rect 20471 1540 20475 1545
rect 20501 1565 20503 1570
rect 20847 1570 20879 1575
rect 20847 1565 20849 1570
rect 20501 1545 20849 1565
rect 20501 1540 20503 1545
rect 20471 1535 20503 1540
rect 20847 1540 20849 1545
rect 20875 1540 20879 1570
rect 20847 1535 20879 1540
rect 5135 1510 5175 1515
rect 2925 1500 2965 1505
rect 2925 1470 2930 1500
rect 2960 1495 2965 1500
rect 3045 1500 3085 1505
rect 3045 1495 3050 1500
rect 2960 1475 3050 1495
rect 2960 1470 2965 1475
rect 2925 1465 2965 1470
rect 3045 1470 3050 1475
rect 3080 1495 3085 1500
rect 3165 1500 3205 1505
rect 3165 1495 3170 1500
rect 3080 1475 3170 1495
rect 3080 1470 3085 1475
rect 3045 1465 3085 1470
rect 3165 1470 3170 1475
rect 3200 1495 3205 1500
rect 3285 1500 3325 1505
rect 3285 1495 3290 1500
rect 3200 1475 3290 1495
rect 3200 1470 3205 1475
rect 3165 1465 3205 1470
rect 3285 1470 3290 1475
rect 3320 1495 3325 1500
rect 3525 1500 3565 1505
rect 3525 1495 3530 1500
rect 3320 1475 3530 1495
rect 3320 1470 3325 1475
rect 3285 1465 3325 1470
rect 3525 1470 3530 1475
rect 3560 1495 3565 1500
rect 3645 1500 3685 1505
rect 3645 1495 3650 1500
rect 3560 1475 3650 1495
rect 3560 1470 3565 1475
rect 3525 1465 3565 1470
rect 3645 1470 3650 1475
rect 3680 1495 3685 1500
rect 3765 1500 3805 1505
rect 3765 1495 3770 1500
rect 3680 1475 3770 1495
rect 3680 1470 3685 1475
rect 3645 1465 3685 1470
rect 3765 1470 3770 1475
rect 3800 1495 3805 1500
rect 4205 1500 4245 1505
rect 4205 1495 4210 1500
rect 3800 1475 4210 1495
rect 3800 1470 3805 1475
rect 3765 1465 3805 1470
rect 4205 1470 4210 1475
rect 4240 1495 4245 1500
rect 4325 1500 4365 1505
rect 4325 1495 4330 1500
rect 4240 1475 4330 1495
rect 4240 1470 4245 1475
rect 4205 1465 4245 1470
rect 4325 1470 4330 1475
rect 4360 1495 4365 1500
rect 4445 1500 4485 1505
rect 4445 1495 4450 1500
rect 4360 1475 4450 1495
rect 4360 1470 4365 1475
rect 4325 1465 4365 1470
rect 4445 1470 4450 1475
rect 4480 1495 4485 1500
rect 4685 1500 4725 1505
rect 4685 1495 4690 1500
rect 4480 1475 4690 1495
rect 4480 1470 4485 1475
rect 4445 1465 4485 1470
rect 4685 1470 4690 1475
rect 4720 1495 4725 1500
rect 4805 1500 4845 1505
rect 4805 1495 4810 1500
rect 4720 1475 4810 1495
rect 4720 1470 4725 1475
rect 4685 1465 4725 1470
rect 4805 1470 4810 1475
rect 4840 1495 4845 1500
rect 4925 1500 4965 1505
rect 4925 1495 4930 1500
rect 4840 1475 4930 1495
rect 4840 1470 4845 1475
rect 4805 1465 4845 1470
rect 4925 1470 4930 1475
rect 4960 1495 4965 1500
rect 5045 1500 5085 1505
rect 5045 1495 5050 1500
rect 4960 1475 5050 1495
rect 4960 1470 4965 1475
rect 4925 1465 4965 1470
rect 5045 1470 5050 1475
rect 5080 1495 5085 1500
rect 5550 1500 5590 1505
rect 5550 1495 5555 1500
rect 5080 1475 5555 1495
rect 5080 1470 5085 1475
rect 5045 1465 5085 1470
rect 5550 1470 5555 1475
rect 5585 1470 5590 1500
rect 11106 1495 11138 1500
rect 11106 1490 11109 1495
rect 10910 1470 11109 1490
rect 5550 1465 5590 1470
rect 11106 1465 11109 1470
rect 11135 1490 11138 1495
rect 11305 1495 11345 1500
rect 11305 1490 11310 1495
rect 11135 1470 11310 1490
rect 11135 1465 11138 1470
rect 11106 1460 11138 1465
rect 11305 1465 11310 1470
rect 11340 1490 11345 1495
rect 11525 1495 11565 1500
rect 11525 1490 11530 1495
rect 11340 1470 11530 1490
rect 11340 1465 11345 1470
rect 11305 1460 11345 1465
rect 11525 1465 11530 1470
rect 11560 1490 11565 1495
rect 11922 1495 11954 1500
rect 11922 1490 11925 1495
rect 11560 1470 11925 1490
rect 11560 1465 11565 1470
rect 11525 1460 11565 1465
rect 11922 1465 11925 1470
rect 11951 1490 11954 1495
rect 12146 1495 12178 1500
rect 12146 1490 12149 1495
rect 11951 1470 12149 1490
rect 11951 1465 11954 1470
rect 11922 1460 11954 1465
rect 12146 1465 12149 1470
rect 12175 1490 12178 1495
rect 12345 1495 12385 1500
rect 12345 1490 12350 1495
rect 12175 1470 12350 1490
rect 12175 1465 12178 1470
rect 12146 1460 12178 1465
rect 12345 1465 12350 1470
rect 12380 1490 12385 1495
rect 12565 1495 12605 1500
rect 12565 1490 12570 1495
rect 12380 1470 12570 1490
rect 12380 1465 12385 1470
rect 12345 1460 12385 1465
rect 12565 1465 12570 1470
rect 12600 1465 12605 1495
rect 18606 1495 18638 1500
rect 18606 1490 18609 1495
rect 18410 1470 18609 1490
rect 12565 1460 12605 1465
rect 18606 1465 18609 1470
rect 18635 1490 18638 1495
rect 18805 1495 18845 1500
rect 18805 1490 18810 1495
rect 18635 1470 18810 1490
rect 18635 1465 18638 1470
rect 18606 1460 18638 1465
rect 18805 1465 18810 1470
rect 18840 1490 18845 1495
rect 19025 1495 19065 1500
rect 19025 1490 19030 1495
rect 18840 1470 19030 1490
rect 18840 1465 18845 1470
rect 18805 1460 18845 1465
rect 19025 1465 19030 1470
rect 19060 1490 19065 1495
rect 19422 1495 19454 1500
rect 19422 1490 19425 1495
rect 19060 1470 19425 1490
rect 19060 1465 19065 1470
rect 19025 1460 19065 1465
rect 19422 1465 19425 1470
rect 19451 1490 19454 1495
rect 19646 1495 19678 1500
rect 19646 1490 19649 1495
rect 19451 1470 19649 1490
rect 19451 1465 19454 1470
rect 19422 1460 19454 1465
rect 19646 1465 19649 1470
rect 19675 1490 19678 1495
rect 19845 1495 19885 1500
rect 19845 1490 19850 1495
rect 19675 1470 19850 1490
rect 19675 1465 19678 1470
rect 19646 1460 19678 1465
rect 19845 1465 19850 1470
rect 19880 1490 19885 1495
rect 20065 1495 20105 1500
rect 20065 1490 20070 1495
rect 19880 1470 20070 1490
rect 19880 1465 19885 1470
rect 19845 1460 19885 1465
rect 20065 1465 20070 1470
rect 20100 1465 20105 1495
rect 20065 1460 20105 1465
rect 11145 1435 11185 1440
rect 11145 1405 11150 1435
rect 11180 1430 11185 1435
rect 11250 1435 11290 1440
rect 11250 1430 11255 1435
rect 11180 1410 11255 1430
rect 11180 1405 11185 1410
rect 11145 1400 11185 1405
rect 11250 1405 11255 1410
rect 11285 1430 11290 1435
rect 11360 1435 11400 1440
rect 11360 1430 11365 1435
rect 11285 1410 11365 1430
rect 11285 1405 11290 1410
rect 11250 1400 11290 1405
rect 11360 1405 11365 1410
rect 11395 1430 11400 1435
rect 11470 1435 11510 1440
rect 11470 1430 11475 1435
rect 11395 1410 11475 1430
rect 11395 1405 11400 1410
rect 11360 1400 11400 1405
rect 11470 1405 11475 1410
rect 11505 1430 11510 1435
rect 11580 1435 11620 1440
rect 11580 1430 11585 1435
rect 11505 1410 11585 1430
rect 11505 1405 11510 1410
rect 11470 1400 11510 1405
rect 11580 1405 11585 1410
rect 11615 1430 11620 1435
rect 12185 1435 12225 1440
rect 12185 1430 12190 1435
rect 11615 1410 12190 1430
rect 11615 1405 11620 1410
rect 11580 1400 11620 1405
rect 12185 1405 12190 1410
rect 12220 1430 12225 1435
rect 12290 1435 12330 1440
rect 12290 1430 12295 1435
rect 12220 1410 12295 1430
rect 12220 1405 12225 1410
rect 12185 1400 12225 1405
rect 12290 1405 12295 1410
rect 12325 1430 12330 1435
rect 12400 1435 12440 1440
rect 12400 1430 12405 1435
rect 12325 1410 12405 1430
rect 12325 1405 12330 1410
rect 12290 1400 12330 1405
rect 12400 1405 12405 1410
rect 12435 1430 12440 1435
rect 12510 1435 12550 1440
rect 12510 1430 12515 1435
rect 12435 1410 12515 1430
rect 12435 1405 12440 1410
rect 12400 1400 12440 1405
rect 12510 1405 12515 1410
rect 12545 1430 12550 1435
rect 12620 1435 12660 1440
rect 12620 1430 12625 1435
rect 12545 1410 12625 1430
rect 12545 1405 12550 1410
rect 12510 1400 12550 1405
rect 12620 1405 12625 1410
rect 12655 1405 12660 1435
rect 18645 1435 18685 1440
rect 12620 1400 12660 1405
rect 13015 1395 13020 1430
rect 13055 1395 13060 1430
rect 14025 1395 14030 1430
rect 14065 1395 14070 1430
rect 18645 1405 18650 1435
rect 18680 1430 18685 1435
rect 18750 1435 18790 1440
rect 18750 1430 18755 1435
rect 18680 1410 18755 1430
rect 18680 1405 18685 1410
rect 18645 1400 18685 1405
rect 18750 1405 18755 1410
rect 18785 1430 18790 1435
rect 18860 1435 18900 1440
rect 18860 1430 18865 1435
rect 18785 1410 18865 1430
rect 18785 1405 18790 1410
rect 18750 1400 18790 1405
rect 18860 1405 18865 1410
rect 18895 1430 18900 1435
rect 18970 1435 19010 1440
rect 18970 1430 18975 1435
rect 18895 1410 18975 1430
rect 18895 1405 18900 1410
rect 18860 1400 18900 1405
rect 18970 1405 18975 1410
rect 19005 1430 19010 1435
rect 19080 1435 19120 1440
rect 19080 1430 19085 1435
rect 19005 1410 19085 1430
rect 19005 1405 19010 1410
rect 18970 1400 19010 1405
rect 19080 1405 19085 1410
rect 19115 1430 19120 1435
rect 19685 1435 19725 1440
rect 19685 1430 19690 1435
rect 19115 1410 19690 1430
rect 19115 1405 19120 1410
rect 19080 1400 19120 1405
rect 19685 1405 19690 1410
rect 19720 1430 19725 1435
rect 19790 1435 19830 1440
rect 19790 1430 19795 1435
rect 19720 1410 19795 1430
rect 19720 1405 19725 1410
rect 19685 1400 19725 1405
rect 19790 1405 19795 1410
rect 19825 1430 19830 1435
rect 19900 1435 19940 1440
rect 19900 1430 19905 1435
rect 19825 1410 19905 1430
rect 19825 1405 19830 1410
rect 19790 1400 19830 1405
rect 19900 1405 19905 1410
rect 19935 1430 19940 1435
rect 20010 1435 20050 1440
rect 20010 1430 20015 1435
rect 19935 1410 20015 1430
rect 19935 1405 19940 1410
rect 19900 1400 19940 1405
rect 20010 1405 20015 1410
rect 20045 1430 20050 1435
rect 20120 1435 20160 1440
rect 20120 1430 20125 1435
rect 20045 1410 20125 1430
rect 20045 1405 20050 1410
rect 20010 1400 20050 1405
rect 20120 1405 20125 1410
rect 20155 1405 20160 1435
rect 20120 1400 20160 1405
rect 19310 1385 19350 1390
rect 13020 1375 13060 1380
rect 13020 1345 13025 1375
rect 13055 1370 13060 1375
rect 13125 1375 13165 1380
rect 13125 1370 13130 1375
rect 13055 1350 13130 1370
rect 13055 1345 13060 1350
rect 13020 1340 13060 1345
rect 13125 1345 13130 1350
rect 13160 1345 13165 1375
rect 19310 1355 19315 1385
rect 19345 1355 19350 1385
rect 19310 1350 19350 1355
rect 20526 1350 20558 1355
rect 20526 1345 20528 1350
rect 13125 1340 13165 1345
rect 11810 1335 11850 1340
rect 11810 1305 11815 1335
rect 11845 1305 11850 1335
rect 18815 1335 18855 1340
rect 11810 1300 11850 1305
rect 13025 1320 13065 1325
rect 13025 1290 13030 1320
rect 13060 1315 13065 1320
rect 13225 1320 13265 1325
rect 13225 1315 13230 1320
rect 13060 1295 13230 1315
rect 13060 1290 13065 1295
rect 11315 1285 11355 1290
rect 11315 1255 11320 1285
rect 11350 1280 11355 1285
rect 11880 1285 11920 1290
rect 13025 1285 13065 1290
rect 13225 1290 13230 1295
rect 13260 1315 13265 1320
rect 13425 1320 13465 1325
rect 13425 1315 13430 1320
rect 13260 1295 13430 1315
rect 13260 1290 13265 1295
rect 13225 1285 13265 1290
rect 13425 1290 13430 1295
rect 13460 1315 13465 1320
rect 13625 1320 13665 1325
rect 13625 1315 13630 1320
rect 13460 1295 13630 1315
rect 13460 1290 13465 1295
rect 13425 1285 13465 1290
rect 13625 1290 13630 1295
rect 13660 1315 13665 1320
rect 13825 1320 13865 1325
rect 13825 1315 13830 1320
rect 13660 1295 13830 1315
rect 13660 1290 13665 1295
rect 13625 1285 13665 1290
rect 13825 1290 13830 1295
rect 13860 1315 13865 1320
rect 14025 1320 14065 1325
rect 14025 1315 14030 1320
rect 13860 1295 14030 1315
rect 13860 1290 13865 1295
rect 13825 1285 13865 1290
rect 14025 1290 14030 1295
rect 14060 1290 14065 1320
rect 18815 1305 18820 1335
rect 18850 1330 18855 1335
rect 19380 1335 19420 1340
rect 19380 1330 19385 1335
rect 18850 1310 19385 1330
rect 18850 1305 18855 1310
rect 18815 1300 18855 1305
rect 19380 1305 19385 1310
rect 19415 1305 19420 1335
rect 20525 1325 20528 1345
rect 20526 1320 20528 1325
rect 20554 1345 20558 1350
rect 20792 1350 20824 1355
rect 20792 1345 20796 1350
rect 20554 1325 20796 1345
rect 20554 1320 20558 1325
rect 20526 1315 20558 1320
rect 20792 1320 20796 1325
rect 20822 1345 20824 1350
rect 20822 1325 20825 1345
rect 20822 1320 20824 1325
rect 20792 1315 20824 1320
rect 19380 1300 19420 1305
rect 14025 1285 14065 1290
rect 20095 1290 20135 1295
rect 11880 1280 11885 1285
rect 11350 1260 11885 1280
rect 11350 1255 11355 1260
rect 11315 1250 11355 1255
rect 11880 1255 11885 1260
rect 11915 1255 11920 1285
rect 11880 1250 11920 1255
rect 18925 1275 18965 1280
rect 18925 1245 18930 1275
rect 18960 1270 18965 1275
rect 19035 1275 19075 1280
rect 19035 1270 19040 1275
rect 18960 1250 19040 1270
rect 18960 1245 18965 1250
rect 12595 1240 12635 1245
rect 18925 1240 18965 1245
rect 19035 1245 19040 1250
rect 19070 1270 19075 1275
rect 19145 1275 19185 1280
rect 19145 1270 19150 1275
rect 19070 1250 19150 1270
rect 19070 1245 19075 1250
rect 19035 1240 19075 1245
rect 19145 1245 19150 1250
rect 19180 1270 19185 1275
rect 19255 1275 19295 1280
rect 19255 1270 19260 1275
rect 19180 1250 19260 1270
rect 19180 1245 19185 1250
rect 19145 1240 19185 1245
rect 19255 1245 19260 1250
rect 19290 1270 19295 1275
rect 19365 1275 19405 1280
rect 19365 1270 19370 1275
rect 19290 1250 19370 1270
rect 19290 1245 19295 1250
rect 19255 1240 19295 1245
rect 19365 1245 19370 1250
rect 19400 1270 19405 1275
rect 19475 1275 19515 1280
rect 19475 1270 19480 1275
rect 19400 1250 19480 1270
rect 19400 1245 19405 1250
rect 19365 1240 19405 1245
rect 19475 1245 19480 1250
rect 19510 1270 19515 1275
rect 19585 1275 19625 1280
rect 19585 1270 19590 1275
rect 19510 1250 19590 1270
rect 19510 1245 19515 1250
rect 19475 1240 19515 1245
rect 19585 1245 19590 1250
rect 19620 1270 19625 1275
rect 19695 1275 19735 1280
rect 19695 1270 19700 1275
rect 19620 1250 19700 1270
rect 19620 1245 19625 1250
rect 19585 1240 19625 1245
rect 19695 1245 19700 1250
rect 19730 1270 19735 1275
rect 19805 1275 19845 1280
rect 19805 1270 19810 1275
rect 19730 1250 19810 1270
rect 19730 1245 19735 1250
rect 19695 1240 19735 1245
rect 19805 1245 19810 1250
rect 19840 1270 19845 1275
rect 19915 1275 19955 1280
rect 19915 1270 19920 1275
rect 19840 1250 19920 1270
rect 19840 1245 19845 1250
rect 19805 1240 19845 1245
rect 19915 1245 19920 1250
rect 19950 1270 19955 1275
rect 20025 1275 20065 1280
rect 20025 1270 20030 1275
rect 19950 1250 20030 1270
rect 19950 1245 19955 1250
rect 19915 1240 19955 1245
rect 20025 1245 20030 1250
rect 20060 1245 20065 1275
rect 20095 1260 20100 1290
rect 20130 1285 20135 1290
rect 20445 1290 20485 1295
rect 20445 1285 20450 1290
rect 20130 1265 20450 1285
rect 20130 1260 20135 1265
rect 20095 1255 20135 1260
rect 20445 1260 20450 1265
rect 20480 1285 20485 1290
rect 20560 1290 20600 1295
rect 20560 1285 20565 1290
rect 20480 1265 20565 1285
rect 20480 1260 20485 1265
rect 20445 1255 20485 1260
rect 20560 1260 20565 1265
rect 20595 1260 20600 1290
rect 20560 1255 20600 1260
rect 20655 1290 20695 1295
rect 20655 1260 20660 1290
rect 20690 1285 20695 1290
rect 20750 1290 20790 1295
rect 20750 1285 20755 1290
rect 20690 1265 20755 1285
rect 20690 1260 20695 1265
rect 20655 1255 20695 1260
rect 20750 1260 20755 1265
rect 20785 1260 20790 1290
rect 20750 1255 20790 1260
rect 20865 1290 20905 1295
rect 20865 1260 20870 1290
rect 20900 1260 20905 1290
rect 20865 1255 20905 1260
rect 20025 1240 20065 1245
rect 11425 1225 11465 1230
rect 11425 1195 11430 1225
rect 11460 1220 11465 1225
rect 11535 1225 11575 1230
rect 11535 1220 11540 1225
rect 11460 1200 11540 1220
rect 11460 1195 11465 1200
rect 11425 1190 11465 1195
rect 11535 1195 11540 1200
rect 11570 1220 11575 1225
rect 11645 1225 11685 1230
rect 11645 1220 11650 1225
rect 11570 1200 11650 1220
rect 11570 1195 11575 1200
rect 11535 1190 11575 1195
rect 11645 1195 11650 1200
rect 11680 1220 11685 1225
rect 11755 1225 11795 1230
rect 11755 1220 11760 1225
rect 11680 1200 11760 1220
rect 11680 1195 11685 1200
rect 11645 1190 11685 1195
rect 11755 1195 11760 1200
rect 11790 1220 11795 1225
rect 11865 1225 11905 1230
rect 11865 1220 11870 1225
rect 11790 1200 11870 1220
rect 11790 1195 11795 1200
rect 11755 1190 11795 1195
rect 11865 1195 11870 1200
rect 11900 1220 11905 1225
rect 11975 1225 12015 1230
rect 11975 1220 11980 1225
rect 11900 1200 11980 1220
rect 11900 1195 11905 1200
rect 11865 1190 11905 1195
rect 11975 1195 11980 1200
rect 12010 1220 12015 1225
rect 12085 1225 12125 1230
rect 12085 1220 12090 1225
rect 12010 1200 12090 1220
rect 12010 1195 12015 1200
rect 11975 1190 12015 1195
rect 12085 1195 12090 1200
rect 12120 1220 12125 1225
rect 12195 1225 12235 1230
rect 12195 1220 12200 1225
rect 12120 1200 12200 1220
rect 12120 1195 12125 1200
rect 12085 1190 12125 1195
rect 12195 1195 12200 1200
rect 12230 1220 12235 1225
rect 12305 1225 12345 1230
rect 12305 1220 12310 1225
rect 12230 1200 12310 1220
rect 12230 1195 12235 1200
rect 12195 1190 12235 1195
rect 12305 1195 12310 1200
rect 12340 1220 12345 1225
rect 12415 1225 12455 1230
rect 12415 1220 12420 1225
rect 12340 1200 12420 1220
rect 12340 1195 12345 1200
rect 12305 1190 12345 1195
rect 12415 1195 12420 1200
rect 12450 1220 12455 1225
rect 12525 1225 12565 1230
rect 12525 1220 12530 1225
rect 12450 1200 12530 1220
rect 12450 1195 12455 1200
rect 12415 1190 12455 1195
rect 12525 1195 12530 1200
rect 12560 1195 12565 1225
rect 12595 1210 12600 1240
rect 12630 1235 12635 1240
rect 12630 1215 12695 1235
rect 20600 1230 20640 1235
rect 12630 1210 12635 1215
rect 12595 1205 12635 1210
rect 20600 1200 20605 1230
rect 20635 1225 20640 1230
rect 20660 1230 20690 1235
rect 20635 1205 20660 1225
rect 20635 1200 20640 1205
rect 20600 1195 20640 1200
rect 20660 1195 20690 1200
rect 20710 1230 20750 1235
rect 20710 1200 20715 1230
rect 20745 1225 20750 1230
rect 20865 1230 20905 1235
rect 20865 1225 20870 1230
rect 20745 1205 20870 1225
rect 20745 1200 20750 1205
rect 20710 1195 20750 1200
rect 20865 1200 20870 1205
rect 20900 1200 20905 1230
rect 20865 1195 20905 1200
rect 12525 1190 12565 1195
rect 3375 1185 3415 1190
rect 3375 1155 3380 1185
rect 3410 1180 3415 1185
rect 3985 1185 4025 1190
rect 3985 1180 3990 1185
rect 3410 1160 3990 1180
rect 3410 1155 3415 1160
rect 3375 1150 3415 1155
rect 3985 1155 3990 1160
rect 4020 1180 4025 1185
rect 4595 1185 4635 1190
rect 4595 1180 4600 1185
rect 4020 1160 4600 1180
rect 4020 1155 4025 1160
rect 3985 1150 4025 1155
rect 4595 1155 4600 1160
rect 4630 1180 4635 1185
rect 5465 1185 5505 1190
rect 5465 1180 5470 1185
rect 4630 1160 5470 1180
rect 4630 1155 4635 1160
rect 4595 1150 4635 1155
rect 5465 1155 5470 1160
rect 5500 1155 5505 1185
rect 5465 1150 5505 1155
rect 2945 1125 2985 1130
rect 2945 1095 2950 1125
rect 2980 1120 2985 1125
rect 3025 1125 3065 1130
rect 3025 1120 3030 1125
rect 2980 1100 3030 1120
rect 2980 1095 2985 1100
rect 2945 1090 2985 1095
rect 3025 1095 3030 1100
rect 3060 1120 3065 1125
rect 3105 1125 3145 1130
rect 3105 1120 3110 1125
rect 3060 1100 3110 1120
rect 3060 1095 3065 1100
rect 3025 1090 3065 1095
rect 3105 1095 3110 1100
rect 3140 1120 3145 1125
rect 3185 1125 3225 1130
rect 3185 1120 3190 1125
rect 3140 1100 3190 1120
rect 3140 1095 3145 1100
rect 3105 1090 3145 1095
rect 3185 1095 3190 1100
rect 3220 1120 3225 1125
rect 3265 1125 3305 1130
rect 3265 1120 3270 1125
rect 3220 1100 3270 1120
rect 3220 1095 3225 1100
rect 3185 1090 3225 1095
rect 3265 1095 3270 1100
rect 3300 1120 3305 1125
rect 3345 1125 3385 1130
rect 3345 1120 3350 1125
rect 3300 1100 3350 1120
rect 3300 1095 3305 1100
rect 3265 1090 3305 1095
rect 3345 1095 3350 1100
rect 3380 1120 3385 1125
rect 3425 1125 3465 1130
rect 3425 1120 3430 1125
rect 3380 1100 3430 1120
rect 3380 1095 3385 1100
rect 3345 1090 3385 1095
rect 3425 1095 3430 1100
rect 3460 1120 3465 1125
rect 3505 1125 3545 1130
rect 3505 1120 3510 1125
rect 3460 1100 3510 1120
rect 3460 1095 3465 1100
rect 3425 1090 3465 1095
rect 3505 1095 3510 1100
rect 3540 1120 3545 1125
rect 3585 1125 3625 1130
rect 3585 1120 3590 1125
rect 3540 1100 3590 1120
rect 3540 1095 3545 1100
rect 3505 1090 3545 1095
rect 3585 1095 3590 1100
rect 3620 1120 3625 1125
rect 3665 1125 3705 1130
rect 3665 1120 3670 1125
rect 3620 1100 3670 1120
rect 3620 1095 3625 1100
rect 3585 1090 3625 1095
rect 3665 1095 3670 1100
rect 3700 1120 3705 1125
rect 3745 1125 3785 1130
rect 3745 1120 3750 1125
rect 3700 1100 3750 1120
rect 3700 1095 3705 1100
rect 3665 1090 3705 1095
rect 3745 1095 3750 1100
rect 3780 1120 3785 1125
rect 3825 1125 3865 1130
rect 3825 1120 3830 1125
rect 3780 1100 3830 1120
rect 3780 1095 3785 1100
rect 3745 1090 3785 1095
rect 3825 1095 3830 1100
rect 3860 1120 3865 1125
rect 3905 1125 3945 1130
rect 3905 1120 3910 1125
rect 3860 1100 3910 1120
rect 3860 1095 3865 1100
rect 3825 1090 3865 1095
rect 3905 1095 3910 1100
rect 3940 1095 3945 1125
rect 3905 1090 3945 1095
rect 3985 1125 4025 1130
rect 3985 1095 3990 1125
rect 4020 1120 4025 1125
rect 4065 1125 4105 1130
rect 4065 1120 4070 1125
rect 4020 1100 4070 1120
rect 4020 1095 4025 1100
rect 3985 1090 4025 1095
rect 4065 1095 4070 1100
rect 4100 1120 4105 1125
rect 4145 1125 4185 1130
rect 4145 1120 4150 1125
rect 4100 1100 4150 1120
rect 4100 1095 4105 1100
rect 4065 1090 4105 1095
rect 4145 1095 4150 1100
rect 4180 1120 4185 1125
rect 4225 1125 4265 1130
rect 4225 1120 4230 1125
rect 4180 1100 4230 1120
rect 4180 1095 4185 1100
rect 4145 1090 4185 1095
rect 4225 1095 4230 1100
rect 4260 1120 4265 1125
rect 4305 1125 4345 1130
rect 4305 1120 4310 1125
rect 4260 1100 4310 1120
rect 4260 1095 4265 1100
rect 4225 1090 4265 1095
rect 4305 1095 4310 1100
rect 4340 1120 4345 1125
rect 4385 1125 4425 1130
rect 4385 1120 4390 1125
rect 4340 1100 4390 1120
rect 4340 1095 4345 1100
rect 4305 1090 4345 1095
rect 4385 1095 4390 1100
rect 4420 1120 4425 1125
rect 4465 1125 4505 1130
rect 4465 1120 4470 1125
rect 4420 1100 4470 1120
rect 4420 1095 4425 1100
rect 4385 1090 4425 1095
rect 4465 1095 4470 1100
rect 4500 1120 4505 1125
rect 4545 1125 4585 1130
rect 4545 1120 4550 1125
rect 4500 1100 4550 1120
rect 4500 1095 4505 1100
rect 4465 1090 4505 1095
rect 4545 1095 4550 1100
rect 4580 1120 4585 1125
rect 4625 1125 4665 1130
rect 4625 1120 4630 1125
rect 4580 1100 4630 1120
rect 4580 1095 4585 1100
rect 4545 1090 4585 1095
rect 4625 1095 4630 1100
rect 4660 1120 4665 1125
rect 4705 1125 4745 1130
rect 4705 1120 4710 1125
rect 4660 1100 4710 1120
rect 4660 1095 4665 1100
rect 4625 1090 4665 1095
rect 4705 1095 4710 1100
rect 4740 1120 4745 1125
rect 4785 1125 4825 1130
rect 4785 1120 4790 1125
rect 4740 1100 4790 1120
rect 4740 1095 4745 1100
rect 4705 1090 4745 1095
rect 4785 1095 4790 1100
rect 4820 1120 4825 1125
rect 4865 1125 4905 1130
rect 4865 1120 4870 1125
rect 4820 1100 4870 1120
rect 4820 1095 4825 1100
rect 4785 1090 4825 1095
rect 4865 1095 4870 1100
rect 4900 1120 4905 1125
rect 4945 1125 4985 1130
rect 4945 1120 4950 1125
rect 4900 1100 4950 1120
rect 4900 1095 4905 1100
rect 4865 1090 4905 1095
rect 4945 1095 4950 1100
rect 4980 1095 4985 1125
rect 4945 1090 4985 1095
rect 2620 1040 2660 1045
rect 2620 1010 2625 1040
rect 2655 1035 2660 1040
rect 2905 1040 2945 1045
rect 2905 1035 2910 1040
rect 2655 1015 2910 1035
rect 2655 1010 2660 1015
rect 2620 1005 2660 1010
rect 2905 1010 2910 1015
rect 2940 1010 2945 1040
rect 2905 1005 2945 1010
rect 5110 1040 5150 1045
rect 5110 1010 5115 1040
rect 5145 1035 5150 1040
rect 5465 1040 5505 1045
rect 5465 1035 5470 1040
rect 5145 1015 5470 1035
rect 5145 1010 5150 1015
rect 5110 1005 5150 1010
rect 5465 1010 5470 1015
rect 5500 1010 5505 1040
rect 5465 1005 5505 1010
rect 13125 970 13165 975
rect 13125 940 13130 970
rect 13160 965 13165 970
rect 13325 970 13365 975
rect 13325 965 13330 970
rect 13160 945 13330 965
rect 13160 940 13165 945
rect 13125 935 13165 940
rect 13325 940 13330 945
rect 13360 965 13365 970
rect 13525 970 13565 975
rect 13525 965 13530 970
rect 13360 945 13530 965
rect 13360 940 13365 945
rect 13325 935 13365 940
rect 13525 940 13530 945
rect 13560 965 13565 970
rect 13725 970 13765 975
rect 13725 965 13730 970
rect 13560 945 13730 965
rect 13560 940 13565 945
rect 13525 935 13565 940
rect 13725 940 13730 945
rect 13760 965 13765 970
rect 13925 970 13965 975
rect 13925 965 13930 970
rect 13760 945 13930 965
rect 13760 940 13765 945
rect 13725 935 13765 940
rect 13925 940 13930 945
rect 13960 940 13965 970
rect 13925 935 13965 940
rect 18665 955 18705 960
rect 2995 930 3035 935
rect 2995 900 3000 930
rect 3030 925 3035 930
rect 3175 930 3215 935
rect 3175 925 3180 930
rect 3030 905 3180 925
rect 3030 900 3035 905
rect 2995 895 3035 900
rect 3175 900 3180 905
rect 3210 925 3215 930
rect 3355 930 3395 935
rect 3355 925 3360 930
rect 3210 905 3360 925
rect 3210 900 3215 905
rect 3175 895 3215 900
rect 3355 900 3360 905
rect 3390 925 3395 930
rect 3535 930 3575 935
rect 3535 925 3540 930
rect 3390 905 3540 925
rect 3390 900 3395 905
rect 3355 895 3395 900
rect 3535 900 3540 905
rect 3570 925 3575 930
rect 3715 930 3755 935
rect 3715 925 3720 930
rect 3570 905 3720 925
rect 3570 900 3575 905
rect 3535 895 3575 900
rect 3715 900 3720 905
rect 3750 925 3755 930
rect 3895 930 3935 935
rect 3895 925 3900 930
rect 3750 905 3900 925
rect 3750 900 3755 905
rect 3715 895 3755 900
rect 3895 900 3900 905
rect 3930 925 3935 930
rect 4075 930 4115 935
rect 4075 925 4080 930
rect 3930 905 4080 925
rect 3930 900 3935 905
rect 3895 895 3935 900
rect 4075 900 4080 905
rect 4110 925 4115 930
rect 4255 930 4295 935
rect 4255 925 4260 930
rect 4110 905 4260 925
rect 4110 900 4115 905
rect 4075 895 4115 900
rect 4255 900 4260 905
rect 4290 925 4295 930
rect 4435 930 4475 935
rect 4435 925 4440 930
rect 4290 905 4440 925
rect 4290 900 4295 905
rect 4255 895 4295 900
rect 4435 900 4440 905
rect 4470 925 4475 930
rect 4615 930 4655 935
rect 4615 925 4620 930
rect 4470 905 4620 925
rect 4470 900 4475 905
rect 4435 895 4475 900
rect 4615 900 4620 905
rect 4650 925 4655 930
rect 4795 930 4835 935
rect 4795 925 4800 930
rect 4650 905 4800 925
rect 4650 900 4655 905
rect 4615 895 4655 900
rect 4795 900 4800 905
rect 4830 925 4835 930
rect 4975 930 5015 935
rect 4975 925 4980 930
rect 4830 905 4980 925
rect 4830 900 4835 905
rect 4795 895 4835 900
rect 4975 900 4980 905
rect 5010 925 5015 930
rect 5465 930 5505 935
rect 5465 925 5470 930
rect 5010 905 5470 925
rect 5010 900 5015 905
rect 4975 895 5015 900
rect 5465 900 5470 905
rect 5500 900 5505 930
rect 18665 925 18670 955
rect 18700 950 18705 955
rect 18760 955 18800 960
rect 18760 950 18765 955
rect 18700 930 18765 950
rect 18700 925 18705 930
rect 18665 920 18705 925
rect 18760 925 18765 930
rect 18795 950 18800 955
rect 18870 955 18910 960
rect 18870 950 18875 955
rect 18795 930 18875 950
rect 18795 925 18800 930
rect 18760 920 18800 925
rect 18870 925 18875 930
rect 18905 950 18910 955
rect 18980 955 19020 960
rect 18980 950 18985 955
rect 18905 930 18985 950
rect 18905 925 18910 930
rect 18870 920 18910 925
rect 18980 925 18985 930
rect 19015 950 19020 955
rect 19090 955 19130 960
rect 19090 950 19095 955
rect 19015 930 19095 950
rect 19015 925 19020 930
rect 18980 920 19020 925
rect 19090 925 19095 930
rect 19125 950 19130 955
rect 19200 955 19240 960
rect 19200 950 19205 955
rect 19125 930 19205 950
rect 19125 925 19130 930
rect 19090 920 19130 925
rect 19200 925 19205 930
rect 19235 950 19240 955
rect 19310 955 19350 960
rect 19310 950 19315 955
rect 19235 930 19315 950
rect 19235 925 19240 930
rect 19200 920 19240 925
rect 19310 925 19315 930
rect 19345 950 19350 955
rect 19420 955 19460 960
rect 19420 950 19425 955
rect 19345 930 19425 950
rect 19345 925 19350 930
rect 19310 920 19350 925
rect 19420 925 19425 930
rect 19455 950 19460 955
rect 19530 955 19570 960
rect 19530 950 19535 955
rect 19455 930 19535 950
rect 19455 925 19460 930
rect 19420 920 19460 925
rect 19530 925 19535 930
rect 19565 950 19570 955
rect 19640 955 19680 960
rect 19640 950 19645 955
rect 19565 930 19645 950
rect 19565 925 19570 930
rect 19530 920 19570 925
rect 19640 925 19645 930
rect 19675 950 19680 955
rect 19750 955 19790 960
rect 19750 950 19755 955
rect 19675 930 19755 950
rect 19675 925 19680 930
rect 19640 920 19680 925
rect 19750 925 19755 930
rect 19785 950 19790 955
rect 19860 955 19900 960
rect 19860 950 19865 955
rect 19785 930 19865 950
rect 19785 925 19790 930
rect 19750 920 19790 925
rect 19860 925 19865 930
rect 19895 950 19900 955
rect 19970 955 20010 960
rect 19970 950 19975 955
rect 19895 930 19975 950
rect 19895 925 19900 930
rect 19860 920 19900 925
rect 19970 925 19975 930
rect 20005 950 20010 955
rect 20120 955 20160 960
rect 20120 950 20125 955
rect 20005 930 20125 950
rect 20005 925 20010 930
rect 19970 920 20010 925
rect 20120 925 20125 930
rect 20155 925 20160 955
rect 20120 920 20160 925
rect 5465 895 5505 900
rect 11165 905 11205 910
rect 11165 875 11170 905
rect 11200 900 11205 905
rect 11260 905 11300 910
rect 11260 900 11265 905
rect 11200 880 11265 900
rect 11200 875 11205 880
rect 11165 870 11205 875
rect 11260 875 11265 880
rect 11295 900 11300 905
rect 11370 905 11410 910
rect 11370 900 11375 905
rect 11295 880 11375 900
rect 11295 875 11300 880
rect 11260 870 11300 875
rect 11370 875 11375 880
rect 11405 900 11410 905
rect 11480 905 11520 910
rect 11480 900 11485 905
rect 11405 880 11485 900
rect 11405 875 11410 880
rect 11370 870 11410 875
rect 11480 875 11485 880
rect 11515 900 11520 905
rect 11590 905 11630 910
rect 11590 900 11595 905
rect 11515 880 11595 900
rect 11515 875 11520 880
rect 11480 870 11520 875
rect 11590 875 11595 880
rect 11625 900 11630 905
rect 11700 905 11740 910
rect 11700 900 11705 905
rect 11625 880 11705 900
rect 11625 875 11630 880
rect 11590 870 11630 875
rect 11700 875 11705 880
rect 11735 900 11740 905
rect 11810 905 11850 910
rect 11810 900 11815 905
rect 11735 880 11815 900
rect 11735 875 11740 880
rect 11700 870 11740 875
rect 11810 875 11815 880
rect 11845 900 11850 905
rect 11920 905 11960 910
rect 11920 900 11925 905
rect 11845 880 11925 900
rect 11845 875 11850 880
rect 11810 870 11850 875
rect 11920 875 11925 880
rect 11955 900 11960 905
rect 12030 905 12070 910
rect 12030 900 12035 905
rect 11955 880 12035 900
rect 11955 875 11960 880
rect 11920 870 11960 875
rect 12030 875 12035 880
rect 12065 900 12070 905
rect 12140 905 12180 910
rect 12140 900 12145 905
rect 12065 880 12145 900
rect 12065 875 12070 880
rect 12030 870 12070 875
rect 12140 875 12145 880
rect 12175 900 12180 905
rect 12250 905 12290 910
rect 12250 900 12255 905
rect 12175 880 12255 900
rect 12175 875 12180 880
rect 12140 870 12180 875
rect 12250 875 12255 880
rect 12285 900 12290 905
rect 12360 905 12400 910
rect 12360 900 12365 905
rect 12285 880 12365 900
rect 12285 875 12290 880
rect 12250 870 12290 875
rect 12360 875 12365 880
rect 12395 900 12400 905
rect 12470 905 12510 910
rect 12470 900 12475 905
rect 12395 880 12475 900
rect 12395 875 12400 880
rect 12360 870 12400 875
rect 12470 875 12475 880
rect 12505 900 12510 905
rect 12620 905 12660 910
rect 12620 900 12625 905
rect 12505 880 12625 900
rect 12505 875 12510 880
rect 12470 870 12510 875
rect 12620 875 12625 880
rect 12655 875 12660 905
rect 12620 870 12660 875
rect 2520 760 2560 765
rect 2520 730 2525 760
rect 2555 755 2560 760
rect 3130 760 3170 765
rect 3130 755 3135 760
rect 2555 735 3135 755
rect 2555 730 2560 735
rect 2520 725 2560 730
rect 3130 730 3135 735
rect 3165 730 3170 760
rect 3130 725 3170 730
rect 3625 760 3665 765
rect 3625 730 3630 760
rect 3660 755 3665 760
rect 3985 760 4025 765
rect 3985 755 3990 760
rect 3660 735 3990 755
rect 3660 730 3665 735
rect 3625 725 3665 730
rect 3985 730 3990 735
rect 4020 755 4025 760
rect 4345 760 4385 765
rect 4345 755 4350 760
rect 4020 735 4350 755
rect 4020 730 4025 735
rect 3985 725 4025 730
rect 4345 730 4350 735
rect 4380 730 4385 760
rect 4345 725 4385 730
rect 4525 760 4565 765
rect 4525 730 4530 760
rect 4560 755 4565 760
rect 4705 760 4745 765
rect 4705 755 4710 760
rect 4560 735 4710 755
rect 4560 730 4565 735
rect 4525 725 4565 730
rect 4705 730 4710 735
rect 4740 755 4745 760
rect 4885 760 4925 765
rect 4885 755 4890 760
rect 4740 735 4890 755
rect 4740 730 4745 735
rect 4705 725 4745 730
rect 4885 730 4890 735
rect 4920 730 4925 760
rect 4885 725 4925 730
rect 3445 705 3485 710
rect 3445 675 3450 705
rect 3480 700 3485 705
rect 3805 705 3845 710
rect 3805 700 3810 705
rect 3480 680 3810 700
rect 3480 675 3485 680
rect 3445 670 3485 675
rect 3805 675 3810 680
rect 3840 700 3845 705
rect 4165 705 4205 710
rect 4165 700 4170 705
rect 3840 680 4170 700
rect 3840 675 3845 680
rect 3805 670 3845 675
rect 4165 675 4170 680
rect 4200 675 4205 705
rect 4165 670 4205 675
rect -195 575 -155 580
rect -195 545 -190 575
rect -160 545 -155 575
rect -195 540 -155 545
rect 9375 -680 9415 -675
rect 9375 -710 9380 -680
rect 9410 -685 9415 -680
rect 9575 -680 9615 -675
rect 9575 -685 9580 -680
rect 9410 -705 9580 -685
rect 9410 -710 9415 -705
rect 9375 -715 9415 -710
rect 9575 -710 9580 -705
rect 9610 -685 9615 -680
rect 9775 -680 9815 -675
rect 9775 -685 9780 -680
rect 9610 -705 9780 -685
rect 9610 -710 9615 -705
rect 9575 -715 9615 -710
rect 9775 -710 9780 -705
rect 9810 -685 9815 -680
rect 9975 -680 10015 -675
rect 9975 -685 9980 -680
rect 9810 -705 9980 -685
rect 9810 -710 9815 -705
rect 9775 -715 9815 -710
rect 9975 -710 9980 -705
rect 10010 -685 10015 -680
rect 10175 -680 10215 -675
rect 10175 -685 10180 -680
rect 10010 -705 10180 -685
rect 10010 -710 10015 -705
rect 9975 -715 10015 -710
rect 10175 -710 10180 -705
rect 10210 -685 10215 -680
rect 10375 -680 10415 -675
rect 10375 -685 10380 -680
rect 10210 -705 10380 -685
rect 10210 -710 10215 -705
rect 10175 -715 10215 -710
rect 10375 -710 10380 -705
rect 10410 -710 10415 -680
rect 10375 -715 10415 -710
rect 9475 -1030 9515 -1025
rect 9475 -1060 9480 -1030
rect 9510 -1035 9515 -1030
rect 9675 -1030 9715 -1025
rect 9675 -1035 9680 -1030
rect 9510 -1055 9680 -1035
rect 9510 -1060 9515 -1055
rect 9475 -1065 9515 -1060
rect 9675 -1060 9680 -1055
rect 9710 -1035 9715 -1030
rect 9875 -1030 9915 -1025
rect 9875 -1035 9880 -1030
rect 9710 -1055 9880 -1035
rect 9710 -1060 9715 -1055
rect 9675 -1065 9715 -1060
rect 9875 -1060 9880 -1055
rect 9910 -1035 9915 -1030
rect 10075 -1030 10115 -1025
rect 10075 -1035 10080 -1030
rect 9910 -1055 10080 -1035
rect 9910 -1060 9915 -1055
rect 9875 -1065 9915 -1060
rect 10075 -1060 10080 -1055
rect 10110 -1035 10115 -1030
rect 10275 -1030 10315 -1025
rect 10275 -1035 10280 -1030
rect 10110 -1055 10280 -1035
rect 10110 -1060 10115 -1055
rect 10075 -1065 10115 -1060
rect 10275 -1060 10280 -1055
rect 10310 -1060 10315 -1030
rect 10275 -1065 10315 -1060
<< via2 >>
rect -190 4960 -160 4990
rect 5555 4960 5585 4990
rect -105 3495 -75 3525
rect 4445 3465 4475 3495
rect 945 3415 975 3445
rect 1645 3415 1675 3445
rect 5145 3415 5175 3445
rect 5555 3415 5585 3445
rect 2695 3360 2725 3390
rect 3395 3305 3425 3335
rect -105 3110 -75 3140
rect -105 2970 -75 3000
rect -105 2880 -75 2910
rect 5555 2780 5585 2810
rect 5555 2065 5585 2095
rect -105 1690 -75 1720
rect 5555 1470 5585 1500
rect 5470 1155 5500 1185
rect 5470 1010 5500 1040
rect 5470 900 5500 930
rect -190 545 -160 575
<< metal3 >>
rect -200 4995 -150 5000
rect -200 4955 -195 4995
rect -155 4955 -150 4995
rect -200 4950 -150 4955
rect 5545 4995 5595 5000
rect 5545 4955 5550 4995
rect 5590 4955 5595 4995
rect 5545 4950 5595 4955
rect -195 585 -155 4950
rect -115 4910 -65 4915
rect -115 4870 -110 4910
rect -70 4870 -65 4910
rect -115 4865 -65 4870
rect 5460 4910 5510 4915
rect 5460 4870 5465 4910
rect 5505 4870 5510 4910
rect 5460 4865 5510 4870
rect -110 3525 -70 4865
rect 145 4770 375 4855
rect 495 4770 725 4855
rect 845 4770 1075 4855
rect 1195 4770 1425 4855
rect 1545 4770 1775 4855
rect 145 4720 1775 4770
rect 145 4625 375 4720
rect 495 4625 725 4720
rect 845 4625 1075 4720
rect 1195 4625 1425 4720
rect 1545 4625 1775 4720
rect 1895 4770 2125 4855
rect 2245 4770 2475 4855
rect 2595 4770 2825 4855
rect 2945 4770 3175 4855
rect 3295 4770 3525 4855
rect 1895 4720 3525 4770
rect 1895 4625 2125 4720
rect 2245 4625 2475 4720
rect 2595 4625 2825 4720
rect 2945 4625 3175 4720
rect 3295 4625 3525 4720
rect 3645 4770 3875 4855
rect 3995 4770 4225 4855
rect 4345 4770 4575 4855
rect 4695 4770 4925 4855
rect 5045 4770 5275 4855
rect 3645 4720 5275 4770
rect 3645 4625 3875 4720
rect 3995 4625 4225 4720
rect 4345 4625 4575 4720
rect 4695 4625 4925 4720
rect 5045 4625 5275 4720
rect 935 4505 985 4625
rect 2685 4505 2735 4625
rect 4435 4505 4485 4625
rect 145 4420 375 4505
rect 495 4420 725 4505
rect 845 4420 1075 4505
rect 1195 4420 1425 4505
rect 1545 4420 1775 4505
rect 145 4370 1775 4420
rect 145 4275 375 4370
rect 495 4275 725 4370
rect 845 4275 1075 4370
rect 1195 4275 1425 4370
rect 1545 4275 1775 4370
rect 1895 4420 2125 4505
rect 2245 4420 2475 4505
rect 2595 4420 2825 4505
rect 2945 4420 3175 4505
rect 3295 4420 3525 4505
rect 1895 4370 3525 4420
rect 1895 4275 2125 4370
rect 2245 4275 2475 4370
rect 2595 4275 2825 4370
rect 2945 4275 3175 4370
rect 3295 4275 3525 4370
rect 3645 4420 3875 4505
rect 3995 4420 4225 4505
rect 4345 4420 4575 4505
rect 4695 4420 4925 4505
rect 5045 4420 5275 4505
rect 3645 4370 5275 4420
rect 3645 4275 3875 4370
rect 3995 4275 4225 4370
rect 4345 4275 4575 4370
rect 4695 4275 4925 4370
rect 5045 4275 5275 4370
rect 935 4155 985 4275
rect 2685 4155 2735 4275
rect 4435 4155 4485 4275
rect 145 4070 375 4155
rect 495 4070 725 4155
rect 845 4070 1075 4155
rect 1195 4070 1425 4155
rect 1545 4070 1775 4155
rect 145 4020 1775 4070
rect 145 3925 375 4020
rect 495 3925 725 4020
rect 845 3925 1075 4020
rect 1195 3925 1425 4020
rect 1545 3925 1775 4020
rect 1895 4070 2125 4155
rect 2245 4070 2475 4155
rect 2595 4070 2825 4155
rect 2945 4070 3175 4155
rect 3295 4070 3525 4155
rect 1895 4020 3525 4070
rect 1895 3925 2125 4020
rect 2245 3925 2475 4020
rect 2595 3925 2825 4020
rect 2945 3925 3175 4020
rect 3295 3925 3525 4020
rect 3645 4070 3875 4155
rect 3995 4070 4225 4155
rect 4345 4070 4575 4155
rect 4695 4070 4925 4155
rect 5045 4070 5275 4155
rect 3645 4020 5275 4070
rect 3645 3925 3875 4020
rect 3995 3925 4225 4020
rect 4345 3925 4575 4020
rect 4695 3925 4925 4020
rect 5045 3925 5275 4020
rect 935 3805 985 3925
rect 2685 3805 2735 3925
rect 4435 3805 4485 3925
rect 145 3720 375 3805
rect 495 3720 725 3805
rect 845 3720 1075 3805
rect 1195 3720 1425 3805
rect 1545 3720 1775 3805
rect 145 3670 1775 3720
rect 145 3575 375 3670
rect 495 3575 725 3670
rect 845 3575 1075 3670
rect 1195 3575 1425 3670
rect 1545 3575 1775 3670
rect 1895 3720 2125 3805
rect 2245 3720 2475 3805
rect 2595 3720 2825 3805
rect 2945 3720 3175 3805
rect 3295 3720 3525 3805
rect 1895 3670 3525 3720
rect 1895 3575 2125 3670
rect 2245 3575 2475 3670
rect 2595 3575 2825 3670
rect 2945 3575 3175 3670
rect 3295 3575 3525 3670
rect 3645 3720 3875 3805
rect 3995 3720 4225 3805
rect 4345 3720 4575 3805
rect 4695 3720 4925 3805
rect 5045 3720 5275 3805
rect 3645 3670 5275 3720
rect 3645 3575 3875 3670
rect 3995 3575 4225 3670
rect 4345 3575 4575 3670
rect 4695 3575 4925 3670
rect 5045 3575 5275 3670
rect -110 3495 -105 3525
rect -75 3495 -70 3525
rect -110 3140 -70 3495
rect 940 3445 980 3575
rect 940 3415 945 3445
rect 975 3415 980 3445
rect 940 3410 980 3415
rect 1635 3450 1685 3455
rect 1635 3410 1640 3450
rect 1680 3410 1685 3450
rect 1635 3405 1685 3410
rect 2690 3390 2730 3575
rect 4440 3495 4480 3575
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect 5135 3450 5185 3455
rect 5135 3410 5140 3450
rect 5180 3410 5185 3450
rect 5135 3405 5185 3410
rect 2690 3360 2695 3390
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 3385 3340 3435 3345
rect 3385 3300 3390 3340
rect 3430 3300 3435 3340
rect 3385 3295 3435 3300
rect -110 3110 -105 3140
rect -75 3110 -70 3140
rect -110 3000 -70 3110
rect -110 2970 -105 3000
rect -75 2970 -70 3000
rect -110 2910 -70 2970
rect -110 2880 -105 2910
rect -75 2880 -70 2910
rect -110 1720 -70 2880
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 665 -70 1690
rect 5465 1185 5505 4865
rect 5465 1155 5470 1185
rect 5500 1155 5505 1185
rect 5465 1040 5505 1155
rect 5465 1010 5470 1040
rect 5500 1010 5505 1040
rect 5465 930 5505 1010
rect 5465 900 5470 930
rect 5500 900 5505 930
rect 5465 665 5505 900
rect 5550 3445 5590 4950
rect 5550 3415 5555 3445
rect 5585 3415 5590 3445
rect 5550 2810 5590 3415
rect 5550 2780 5555 2810
rect 5585 2780 5590 2810
rect 5550 2095 5590 2780
rect 5550 2065 5555 2095
rect 5585 2065 5590 2095
rect 5550 1500 5590 2065
rect 5550 1470 5555 1500
rect 5585 1470 5590 1500
rect -115 660 -65 665
rect -115 620 -110 660
rect -70 620 -65 660
rect -115 615 -65 620
rect 5460 660 5510 665
rect 5460 620 5465 660
rect 5505 620 5510 660
rect 5460 615 5510 620
rect 5550 585 5590 1470
rect -200 580 -150 585
rect -200 540 -195 580
rect -155 540 -150 580
rect -200 535 -150 540
rect 5545 580 5595 585
rect 5545 540 5550 580
rect 5590 540 5595 580
rect 5545 535 5595 540
<< via3 >>
rect -195 4990 -155 4995
rect -195 4960 -190 4990
rect -190 4960 -160 4990
rect -160 4960 -155 4990
rect -195 4955 -155 4960
rect 5550 4990 5590 4995
rect 5550 4960 5555 4990
rect 5555 4960 5585 4990
rect 5585 4960 5590 4990
rect 5550 4955 5590 4960
rect -110 4870 -70 4910
rect 5465 4870 5505 4910
rect 1640 3445 1680 3450
rect 1640 3415 1645 3445
rect 1645 3415 1675 3445
rect 1675 3415 1680 3445
rect 1640 3410 1680 3415
rect 5140 3445 5180 3450
rect 5140 3415 5145 3445
rect 5145 3415 5175 3445
rect 5175 3415 5180 3445
rect 5140 3410 5180 3415
rect 3390 3335 3430 3340
rect 3390 3305 3395 3335
rect 3395 3305 3425 3335
rect 3425 3305 3430 3335
rect 3390 3300 3430 3305
rect -110 620 -70 660
rect 5465 620 5505 660
rect -195 575 -155 580
rect -195 545 -190 575
rect -190 545 -160 575
rect -160 545 -155 575
rect -195 540 -155 545
rect 5550 540 5590 580
<< mimcap >>
rect 160 4765 360 4840
rect 160 4725 240 4765
rect 280 4725 360 4765
rect 160 4640 360 4725
rect 510 4765 710 4840
rect 510 4725 590 4765
rect 630 4725 710 4765
rect 510 4640 710 4725
rect 860 4765 1060 4840
rect 860 4725 940 4765
rect 980 4725 1060 4765
rect 860 4640 1060 4725
rect 1210 4765 1410 4840
rect 1210 4725 1290 4765
rect 1330 4725 1410 4765
rect 1210 4640 1410 4725
rect 1560 4765 1760 4840
rect 1560 4725 1640 4765
rect 1680 4725 1760 4765
rect 1560 4640 1760 4725
rect 1910 4765 2110 4840
rect 1910 4725 1990 4765
rect 2030 4725 2110 4765
rect 1910 4640 2110 4725
rect 2260 4765 2460 4840
rect 2260 4725 2340 4765
rect 2380 4725 2460 4765
rect 2260 4640 2460 4725
rect 2610 4765 2810 4840
rect 2610 4725 2690 4765
rect 2730 4725 2810 4765
rect 2610 4640 2810 4725
rect 2960 4765 3160 4840
rect 2960 4725 3040 4765
rect 3080 4725 3160 4765
rect 2960 4640 3160 4725
rect 3310 4765 3510 4840
rect 3310 4725 3390 4765
rect 3430 4725 3510 4765
rect 3310 4640 3510 4725
rect 3660 4765 3860 4840
rect 3660 4725 3740 4765
rect 3780 4725 3860 4765
rect 3660 4640 3860 4725
rect 4010 4765 4210 4840
rect 4010 4725 4090 4765
rect 4130 4725 4210 4765
rect 4010 4640 4210 4725
rect 4360 4765 4560 4840
rect 4360 4725 4440 4765
rect 4480 4725 4560 4765
rect 4360 4640 4560 4725
rect 4710 4765 4910 4840
rect 4710 4725 4790 4765
rect 4830 4725 4910 4765
rect 4710 4640 4910 4725
rect 5060 4765 5260 4840
rect 5060 4725 5140 4765
rect 5180 4725 5260 4765
rect 5060 4640 5260 4725
rect 160 4415 360 4490
rect 160 4375 240 4415
rect 280 4375 360 4415
rect 160 4290 360 4375
rect 510 4415 710 4490
rect 510 4375 590 4415
rect 630 4375 710 4415
rect 510 4290 710 4375
rect 860 4415 1060 4490
rect 860 4375 940 4415
rect 980 4375 1060 4415
rect 860 4290 1060 4375
rect 1210 4415 1410 4490
rect 1210 4375 1290 4415
rect 1330 4375 1410 4415
rect 1210 4290 1410 4375
rect 1560 4415 1760 4490
rect 1560 4375 1640 4415
rect 1680 4375 1760 4415
rect 1560 4290 1760 4375
rect 1910 4415 2110 4490
rect 1910 4375 1990 4415
rect 2030 4375 2110 4415
rect 1910 4290 2110 4375
rect 2260 4415 2460 4490
rect 2260 4375 2340 4415
rect 2380 4375 2460 4415
rect 2260 4290 2460 4375
rect 2610 4415 2810 4490
rect 2610 4375 2690 4415
rect 2730 4375 2810 4415
rect 2610 4290 2810 4375
rect 2960 4415 3160 4490
rect 2960 4375 3040 4415
rect 3080 4375 3160 4415
rect 2960 4290 3160 4375
rect 3310 4415 3510 4490
rect 3310 4375 3390 4415
rect 3430 4375 3510 4415
rect 3310 4290 3510 4375
rect 3660 4415 3860 4490
rect 3660 4375 3740 4415
rect 3780 4375 3860 4415
rect 3660 4290 3860 4375
rect 4010 4415 4210 4490
rect 4010 4375 4090 4415
rect 4130 4375 4210 4415
rect 4010 4290 4210 4375
rect 4360 4415 4560 4490
rect 4360 4375 4440 4415
rect 4480 4375 4560 4415
rect 4360 4290 4560 4375
rect 4710 4415 4910 4490
rect 4710 4375 4790 4415
rect 4830 4375 4910 4415
rect 4710 4290 4910 4375
rect 5060 4415 5260 4490
rect 5060 4375 5140 4415
rect 5180 4375 5260 4415
rect 5060 4290 5260 4375
rect 160 4065 360 4140
rect 160 4025 240 4065
rect 280 4025 360 4065
rect 160 3940 360 4025
rect 510 4065 710 4140
rect 510 4025 590 4065
rect 630 4025 710 4065
rect 510 3940 710 4025
rect 860 4065 1060 4140
rect 860 4025 940 4065
rect 980 4025 1060 4065
rect 860 3940 1060 4025
rect 1210 4065 1410 4140
rect 1210 4025 1290 4065
rect 1330 4025 1410 4065
rect 1210 3940 1410 4025
rect 1560 4065 1760 4140
rect 1560 4025 1640 4065
rect 1680 4025 1760 4065
rect 1560 3940 1760 4025
rect 1910 4065 2110 4140
rect 1910 4025 1990 4065
rect 2030 4025 2110 4065
rect 1910 3940 2110 4025
rect 2260 4065 2460 4140
rect 2260 4025 2340 4065
rect 2380 4025 2460 4065
rect 2260 3940 2460 4025
rect 2610 4065 2810 4140
rect 2610 4025 2690 4065
rect 2730 4025 2810 4065
rect 2610 3940 2810 4025
rect 2960 4065 3160 4140
rect 2960 4025 3040 4065
rect 3080 4025 3160 4065
rect 2960 3940 3160 4025
rect 3310 4065 3510 4140
rect 3310 4025 3390 4065
rect 3430 4025 3510 4065
rect 3310 3940 3510 4025
rect 3660 4065 3860 4140
rect 3660 4025 3740 4065
rect 3780 4025 3860 4065
rect 3660 3940 3860 4025
rect 4010 4065 4210 4140
rect 4010 4025 4090 4065
rect 4130 4025 4210 4065
rect 4010 3940 4210 4025
rect 4360 4065 4560 4140
rect 4360 4025 4440 4065
rect 4480 4025 4560 4065
rect 4360 3940 4560 4025
rect 4710 4065 4910 4140
rect 4710 4025 4790 4065
rect 4830 4025 4910 4065
rect 4710 3940 4910 4025
rect 5060 4065 5260 4140
rect 5060 4025 5140 4065
rect 5180 4025 5260 4065
rect 5060 3940 5260 4025
rect 160 3715 360 3790
rect 160 3675 240 3715
rect 280 3675 360 3715
rect 160 3590 360 3675
rect 510 3715 710 3790
rect 510 3675 590 3715
rect 630 3675 710 3715
rect 510 3590 710 3675
rect 860 3715 1060 3790
rect 860 3675 940 3715
rect 980 3675 1060 3715
rect 860 3590 1060 3675
rect 1210 3715 1410 3790
rect 1210 3675 1290 3715
rect 1330 3675 1410 3715
rect 1210 3590 1410 3675
rect 1560 3715 1760 3790
rect 1560 3675 1640 3715
rect 1680 3675 1760 3715
rect 1560 3590 1760 3675
rect 1910 3715 2110 3790
rect 1910 3675 1990 3715
rect 2030 3675 2110 3715
rect 1910 3590 2110 3675
rect 2260 3715 2460 3790
rect 2260 3675 2340 3715
rect 2380 3675 2460 3715
rect 2260 3590 2460 3675
rect 2610 3715 2810 3790
rect 2610 3675 2690 3715
rect 2730 3675 2810 3715
rect 2610 3590 2810 3675
rect 2960 3715 3160 3790
rect 2960 3675 3040 3715
rect 3080 3675 3160 3715
rect 2960 3590 3160 3675
rect 3310 3715 3510 3790
rect 3310 3675 3390 3715
rect 3430 3675 3510 3715
rect 3310 3590 3510 3675
rect 3660 3715 3860 3790
rect 3660 3675 3740 3715
rect 3780 3675 3860 3715
rect 3660 3590 3860 3675
rect 4010 3715 4210 3790
rect 4010 3675 4090 3715
rect 4130 3675 4210 3715
rect 4010 3590 4210 3675
rect 4360 3715 4560 3790
rect 4360 3675 4440 3715
rect 4480 3675 4560 3715
rect 4360 3590 4560 3675
rect 4710 3715 4910 3790
rect 4710 3675 4790 3715
rect 4830 3675 4910 3715
rect 4710 3590 4910 3675
rect 5060 3715 5260 3790
rect 5060 3675 5140 3715
rect 5180 3675 5260 3715
rect 5060 3590 5260 3675
<< mimcapcontact >>
rect 240 4725 280 4765
rect 590 4725 630 4765
rect 940 4725 980 4765
rect 1290 4725 1330 4765
rect 1640 4725 1680 4765
rect 1990 4725 2030 4765
rect 2340 4725 2380 4765
rect 2690 4725 2730 4765
rect 3040 4725 3080 4765
rect 3390 4725 3430 4765
rect 3740 4725 3780 4765
rect 4090 4725 4130 4765
rect 4440 4725 4480 4765
rect 4790 4725 4830 4765
rect 5140 4725 5180 4765
rect 240 4375 280 4415
rect 590 4375 630 4415
rect 940 4375 980 4415
rect 1290 4375 1330 4415
rect 1640 4375 1680 4415
rect 1990 4375 2030 4415
rect 2340 4375 2380 4415
rect 2690 4375 2730 4415
rect 3040 4375 3080 4415
rect 3390 4375 3430 4415
rect 3740 4375 3780 4415
rect 4090 4375 4130 4415
rect 4440 4375 4480 4415
rect 4790 4375 4830 4415
rect 5140 4375 5180 4415
rect 240 4025 280 4065
rect 590 4025 630 4065
rect 940 4025 980 4065
rect 1290 4025 1330 4065
rect 1640 4025 1680 4065
rect 1990 4025 2030 4065
rect 2340 4025 2380 4065
rect 2690 4025 2730 4065
rect 3040 4025 3080 4065
rect 3390 4025 3430 4065
rect 3740 4025 3780 4065
rect 4090 4025 4130 4065
rect 4440 4025 4480 4065
rect 4790 4025 4830 4065
rect 5140 4025 5180 4065
rect 240 3675 280 3715
rect 590 3675 630 3715
rect 940 3675 980 3715
rect 1290 3675 1330 3715
rect 1640 3675 1680 3715
rect 1990 3675 2030 3715
rect 2340 3675 2380 3715
rect 2690 3675 2730 3715
rect 3040 3675 3080 3715
rect 3390 3675 3430 3715
rect 3740 3675 3780 3715
rect 4090 3675 4130 3715
rect 4440 3675 4480 3715
rect 4790 3675 4830 3715
rect 5140 3675 5180 3715
<< metal4 >>
rect -200 4995 5595 5000
rect -200 4955 -195 4995
rect -155 4955 5550 4995
rect 5590 4955 5595 4995
rect -200 4950 5595 4955
rect -115 4910 5510 4915
rect -115 4870 -110 4910
rect -70 4870 5465 4910
rect 5505 4870 5510 4910
rect -115 4865 5510 4870
rect 235 4765 1685 4770
rect 235 4725 240 4765
rect 280 4725 590 4765
rect 630 4725 940 4765
rect 980 4725 1290 4765
rect 1330 4725 1640 4765
rect 1680 4725 1685 4765
rect 235 4720 1685 4725
rect 1985 4765 3435 4770
rect 1985 4725 1990 4765
rect 2030 4725 2340 4765
rect 2380 4725 2690 4765
rect 2730 4725 3040 4765
rect 3080 4725 3390 4765
rect 3430 4725 3435 4765
rect 1985 4720 3435 4725
rect 3735 4765 5185 4770
rect 3735 4725 3740 4765
rect 3780 4725 4090 4765
rect 4130 4725 4440 4765
rect 4480 4725 4790 4765
rect 4830 4725 5140 4765
rect 5180 4725 5185 4765
rect 3735 4720 5185 4725
rect 935 4420 985 4720
rect 2685 4420 2735 4720
rect 4435 4420 4485 4720
rect 235 4415 1685 4420
rect 235 4375 240 4415
rect 280 4375 590 4415
rect 630 4375 940 4415
rect 980 4375 1290 4415
rect 1330 4375 1640 4415
rect 1680 4375 1685 4415
rect 235 4370 1685 4375
rect 1985 4415 3435 4420
rect 1985 4375 1990 4415
rect 2030 4375 2340 4415
rect 2380 4375 2690 4415
rect 2730 4375 3040 4415
rect 3080 4375 3390 4415
rect 3430 4375 3435 4415
rect 1985 4370 3435 4375
rect 3735 4415 5185 4420
rect 3735 4375 3740 4415
rect 3780 4375 4090 4415
rect 4130 4375 4440 4415
rect 4480 4375 4790 4415
rect 4830 4375 5140 4415
rect 5180 4375 5185 4415
rect 3735 4370 5185 4375
rect 935 4070 985 4370
rect 2685 4070 2735 4370
rect 4435 4070 4485 4370
rect 235 4065 1685 4070
rect 235 4025 240 4065
rect 280 4025 590 4065
rect 630 4025 940 4065
rect 980 4025 1290 4065
rect 1330 4025 1640 4065
rect 1680 4025 1685 4065
rect 235 4020 1685 4025
rect 1985 4065 3435 4070
rect 1985 4025 1990 4065
rect 2030 4025 2340 4065
rect 2380 4025 2690 4065
rect 2730 4025 3040 4065
rect 3080 4025 3390 4065
rect 3430 4025 3435 4065
rect 1985 4020 3435 4025
rect 3735 4065 5185 4070
rect 3735 4025 3740 4065
rect 3780 4025 4090 4065
rect 4130 4025 4440 4065
rect 4480 4025 4790 4065
rect 4830 4025 5140 4065
rect 5180 4025 5185 4065
rect 3735 4020 5185 4025
rect 935 3720 985 4020
rect 2685 3720 2735 4020
rect 4435 3720 4485 4020
rect 235 3715 1685 3720
rect 235 3675 240 3715
rect 280 3675 590 3715
rect 630 3675 940 3715
rect 980 3675 1290 3715
rect 1330 3675 1640 3715
rect 1680 3675 1685 3715
rect 235 3670 1685 3675
rect 1985 3715 3435 3720
rect 1985 3675 1990 3715
rect 2030 3675 2340 3715
rect 2380 3675 2690 3715
rect 2730 3675 3040 3715
rect 3080 3675 3390 3715
rect 3430 3675 3435 3715
rect 1985 3670 3435 3675
rect 3735 3715 5185 3720
rect 3735 3675 3740 3715
rect 3780 3675 4090 3715
rect 4130 3675 4440 3715
rect 4480 3675 4790 3715
rect 4830 3675 5140 3715
rect 5180 3675 5185 3715
rect 3735 3670 5185 3675
rect 1635 3450 1685 3670
rect 1635 3410 1640 3450
rect 1680 3410 1685 3450
rect 1635 3405 1685 3410
rect 3385 3340 3435 3670
rect 5135 3450 5185 3670
rect 5135 3410 5140 3450
rect 5180 3410 5185 3450
rect 5135 3405 5185 3410
rect 3385 3300 3390 3340
rect 3430 3300 3435 3340
rect 3385 3295 3435 3300
rect -115 660 5510 665
rect -115 620 -110 660
rect -70 620 5465 660
rect 5505 620 5510 660
rect -115 615 5510 620
rect -200 580 5595 585
rect -200 540 -195 580
rect -155 540 5550 580
rect 5590 540 5595 580
rect -200 535 5595 540
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 795 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1723858470
transform 1 0 795 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1723858470
transform 1 0 795 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1723858470
transform 1 0 115 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1723858470
transform 1 0 115 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1723858470
transform 1 0 115 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1723858470
transform 1 0 1475 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1723858470
transform 1 0 1475 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1723858470
transform 1 0 1475 0 1 1360
box 0 0 670 670
<< labels >>
flabel metal2 2950 1735 2950 1735 5 FreeSans 400 0 0 -80 Vin-
flabel metal2 2955 1590 2955 1590 1 FreeSans 400 0 0 80 Vin+
flabel metal2 2945 1845 2945 1845 5 FreeSans 400 0 0 -40 V_mir1
flabel metal2 3745 1530 3745 1530 3 FreeSans 400 0 40 0 V_p1
flabel metal1 2650 1155 2650 1155 3 FreeSans 400 0 200 0 START_UP
flabel metal2 3785 1785 3785 1785 5 FreeSans 400 0 0 -40 1st_Vout1
flabel metal2 455 3440 455 3440 1 FreeSans 400 0 0 40 cap_res1
flabel metal3 2730 3375 2730 3375 3 FreeSans 400 0 40 0 cap_res2
flabel metal1 2550 845 2550 845 3 FreeSans 400 0 40 0 NFET_GATE_10uA
flabel metal2 5120 1590 5120 1590 1 FreeSans 400 0 0 80 V_CUR_REF_REG
flabel metal2 4225 1785 4225 1785 5 FreeSans 400 0 0 -40 1st_Vout2
flabel metal2 5065 1845 5065 1845 5 FreeSans 400 0 0 -40 V_mir2
flabel metal2 4265 1530 4265 1530 7 FreeSans 400 0 -40 0 V_p2
flabel metal1 3275 350 3275 350 7 FreeSans 400 0 -400 0 CMFB_NFET_CUR_BIAS
port 8 w
flabel metal1 3825 295 3825 295 5 FreeSans 400 0 0 -200 VB2_CUR_BIAS
port 5 s
flabel metal1 4015 350 4015 350 3 FreeSans 400 0 200 0 ERR_AMP_CUR_BIAS
port 7 e
flabel metal1 4725 295 4725 295 5 FreeSans 400 0 0 -200 VB3_CUR_BIAS
port 6 s
flabel metal1 4985 1110 4985 1110 3 FreeSans 400 0 200 0 START_UP_NFET1
flabel metal2 4115 3135 4115 3135 1 FreeSans 400 0 0 40 PFET_GATE_10uA
flabel metal2 6080 3075 6080 3075 1 FreeSans 400 0 0 200 VB1_CUR_BIAS
port 1 n
flabel metal2 6100 3020 6100 3020 3 FreeSans 400 0 200 0 TAIL_CUR_MIR_BIAS
port 9 e
flabel metal2 6080 2955 6080 2955 5 FreeSans 400 0 0 -200 CMFB_PFET_CUR_BIAS
port 10 s
flabel metal2 6100 1745 6100 1745 3 FreeSans 400 0 200 0 ERR_AMP_REF
port 3 e
flabel metal3 5590 4400 5590 4400 3 FreeSans 800 0 80 0 VDDA
port 4 e
flabel metal3 5505 4175 5505 4175 3 FreeSans 800 0 80 0 GNDA
port 2 e
flabel metal1 2180 1010 2180 1010 3 FreeSans 400 0 40 0 Vbe2
flabel poly 4635 2375 4635 2375 5 FreeSans 400 0 0 -40 V_TOP
<< end >>
