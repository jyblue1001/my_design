magic
tech sky130A
timestamp 1737656614
<< nwell >>
rect -314 88 726 612
<< nmos >>
rect 19 -1 41 42
rect 296 -1 318 42
rect 573 -1 595 42
rect 26 -95 41 -52
rect 303 -95 318 -52
rect 580 -95 595 -52
rect -39 -246 -24 -146
rect 26 -246 41 -146
rect 303 -246 318 -146
rect 580 -246 595 -146
<< pmos >>
rect -246 382 -96 582
rect -46 382 104 582
rect 231 382 381 582
rect 508 382 658 582
rect 26 245 41 331
rect 303 245 318 331
rect 580 245 595 331
rect 19 108 41 194
rect 296 108 318 194
rect 573 108 595 194
<< ndiff >>
rect -31 34 19 42
rect -31 9 -16 34
rect 4 9 19 34
rect -31 -1 19 9
rect 41 34 91 42
rect 41 9 56 34
rect 76 9 91 34
rect 41 -1 91 9
rect 246 34 296 42
rect 246 9 261 34
rect 281 9 296 34
rect 246 -1 296 9
rect 318 34 368 42
rect 318 9 333 34
rect 353 9 368 34
rect 318 -1 368 9
rect 523 34 573 42
rect 523 9 538 34
rect 558 9 573 34
rect 523 -1 573 9
rect 595 34 645 42
rect 595 9 610 34
rect 630 9 645 34
rect 595 -1 645 9
rect -24 -62 26 -52
rect -24 -85 -9 -62
rect 11 -85 26 -62
rect -24 -95 26 -85
rect 41 -62 91 -52
rect 41 -85 56 -62
rect 76 -85 91 -62
rect 41 -95 91 -85
rect 253 -62 303 -52
rect 253 -85 268 -62
rect 288 -85 303 -62
rect 253 -95 303 -85
rect 318 -62 368 -52
rect 318 -85 333 -62
rect 353 -85 368 -62
rect 318 -95 368 -85
rect 530 -62 580 -52
rect 530 -85 545 -62
rect 565 -85 580 -62
rect 530 -95 580 -85
rect 595 -62 645 -52
rect 595 -85 610 -62
rect 630 -85 645 -62
rect 595 -95 645 -85
rect -89 -156 -39 -146
rect -89 -236 -74 -156
rect -54 -236 -39 -156
rect -89 -246 -39 -236
rect -24 -156 26 -146
rect -24 -236 -9 -156
rect 11 -236 26 -156
rect -24 -246 26 -236
rect 41 -156 91 -146
rect 41 -236 56 -156
rect 76 -236 91 -156
rect 41 -246 91 -236
rect 253 -156 303 -146
rect 253 -236 268 -156
rect 288 -236 303 -156
rect 253 -246 303 -236
rect 318 -156 368 -146
rect 318 -236 333 -156
rect 353 -236 368 -156
rect 318 -246 368 -236
rect 530 -156 580 -146
rect 530 -236 545 -156
rect 565 -236 580 -156
rect 530 -246 580 -236
rect 595 -156 645 -146
rect 595 -236 610 -156
rect 630 -236 645 -156
rect 595 -246 645 -236
<< pdiff >>
rect -296 572 -246 582
rect -296 392 -281 572
rect -261 392 -246 572
rect -296 382 -246 392
rect -96 572 -46 582
rect -96 392 -81 572
rect -61 392 -46 572
rect -96 382 -46 392
rect 104 572 154 582
rect 104 392 119 572
rect 139 392 154 572
rect 104 382 154 392
rect 181 572 231 582
rect 181 392 196 572
rect 216 392 231 572
rect 181 382 231 392
rect 381 572 431 582
rect 381 392 396 572
rect 416 392 431 572
rect 381 382 431 392
rect 458 572 508 582
rect 458 392 473 572
rect 493 392 508 572
rect 458 382 508 392
rect 658 572 708 582
rect 658 392 673 572
rect 693 392 708 572
rect 658 382 708 392
rect -24 321 26 331
rect -24 255 -9 321
rect 11 255 26 321
rect -24 245 26 255
rect 41 321 91 331
rect 41 255 56 321
rect 76 255 91 321
rect 41 245 91 255
rect 253 321 303 331
rect 253 255 268 321
rect 288 255 303 321
rect 253 245 303 255
rect 318 321 368 331
rect 318 255 333 321
rect 353 255 368 321
rect 318 245 368 255
rect 530 321 580 331
rect 530 255 545 321
rect 565 255 580 321
rect 530 245 580 255
rect 595 321 645 331
rect 595 255 610 321
rect 630 255 645 321
rect 595 245 645 255
rect -31 186 19 194
rect -31 118 -16 186
rect 4 118 19 186
rect -31 108 19 118
rect 41 186 91 194
rect 41 118 56 186
rect 76 118 91 186
rect 41 108 91 118
rect 246 186 296 194
rect 246 118 261 186
rect 281 118 296 186
rect 246 108 296 118
rect 318 186 368 194
rect 318 118 333 186
rect 353 118 368 186
rect 318 108 368 118
rect 523 186 573 194
rect 523 118 538 186
rect 558 118 573 186
rect 523 108 573 118
rect 595 186 645 194
rect 595 118 610 186
rect 630 118 645 186
rect 595 108 645 118
<< ndiffc >>
rect -16 9 4 34
rect 56 9 76 34
rect 261 9 281 34
rect 333 9 353 34
rect 538 9 558 34
rect 610 9 630 34
rect -9 -85 11 -62
rect 56 -85 76 -62
rect 268 -85 288 -62
rect 333 -85 353 -62
rect 545 -85 565 -62
rect 610 -85 630 -62
rect -74 -236 -54 -156
rect -9 -236 11 -156
rect 56 -236 76 -156
rect 268 -236 288 -156
rect 333 -236 353 -156
rect 545 -236 565 -156
rect 610 -236 630 -156
<< pdiffc >>
rect -281 392 -261 572
rect -81 392 -61 572
rect 119 392 139 572
rect 196 392 216 572
rect 396 392 416 572
rect 473 392 493 572
rect 673 392 693 572
rect -9 255 11 321
rect 56 255 76 321
rect 268 255 288 321
rect 333 255 353 321
rect 545 255 565 321
rect 610 255 630 321
rect -16 118 4 186
rect 56 118 76 186
rect 261 118 281 186
rect 333 118 353 186
rect 538 118 558 186
rect 610 118 630 186
<< psubdiff >>
rect 203 -156 253 -146
rect 203 -236 217 -156
rect 237 -236 253 -156
rect 203 -246 253 -236
<< nsubdiff >>
rect 196 186 246 194
rect 196 118 211 186
rect 231 118 246 186
rect 196 108 246 118
<< psubdiffcont >>
rect 217 -236 237 -156
<< nsubdiffcont >>
rect 211 118 231 186
<< poly >>
rect -246 597 658 612
rect -246 582 -96 597
rect -46 582 104 597
rect 231 582 381 597
rect 508 582 658 597
rect -246 367 -96 382
rect -46 367 104 382
rect 231 367 381 382
rect 508 367 658 382
rect 26 331 41 346
rect 303 331 318 346
rect 580 331 595 346
rect 26 230 41 245
rect 303 230 318 245
rect 580 230 595 245
rect 19 194 41 209
rect 296 194 318 209
rect 573 194 595 209
rect 19 89 41 108
rect 296 89 318 108
rect 573 89 595 108
rect 19 84 81 89
rect -121 74 -81 84
rect -121 54 -111 74
rect -91 54 -81 74
rect -121 44 -81 54
rect 19 64 51 84
rect 71 64 81 84
rect 19 59 81 64
rect 296 84 358 89
rect 296 64 328 84
rect 348 64 358 84
rect 296 59 358 64
rect 573 84 635 89
rect 573 64 605 84
rect 625 64 635 84
rect 573 59 635 64
rect -121 -255 -101 44
rect 19 42 41 59
rect 296 42 318 59
rect 573 42 595 59
rect 19 -16 41 -1
rect 296 -16 318 -1
rect 573 -16 595 -1
rect 26 -52 41 -37
rect 303 -52 318 -37
rect 580 -52 595 -37
rect 26 -110 41 -95
rect 303 -110 318 -95
rect 580 -110 595 -95
rect -39 -146 -24 -131
rect 26 -146 41 -131
rect 303 -146 318 -131
rect 580 -146 595 -131
rect -121 -265 -81 -255
rect -121 -285 -111 -265
rect -91 -285 -81 -265
rect -121 -295 -81 -285
rect -39 -261 -24 -246
rect 26 -261 41 -246
rect 303 -261 318 -246
rect 580 -261 595 -246
rect -39 -276 595 -261
rect -39 -316 -24 -276
rect -295 -331 -24 -316
<< polycont >>
rect -111 54 -91 74
rect 51 64 71 84
rect 328 64 348 84
rect 605 64 625 84
rect -111 -285 -91 -265
<< locali >>
rect -291 572 -251 582
rect -291 392 -281 572
rect -261 392 -251 572
rect -291 -156 -251 392
rect -91 572 -51 582
rect -91 392 -81 572
rect -61 392 -51 572
rect -91 382 -51 392
rect 109 572 149 582
rect 109 392 119 572
rect 139 392 149 572
rect 109 331 149 392
rect 186 572 226 582
rect 186 392 196 572
rect 216 392 226 572
rect 186 382 226 392
rect 386 572 426 582
rect 386 392 396 572
rect 416 392 426 572
rect 386 331 426 392
rect 463 572 503 582
rect 463 392 473 572
rect 493 392 503 572
rect 463 382 503 392
rect 663 572 703 582
rect 663 392 673 572
rect 693 392 703 572
rect 663 331 703 392
rect -19 321 21 331
rect -19 255 -9 321
rect 11 255 21 321
rect -19 245 21 255
rect 46 321 149 331
rect 46 255 56 321
rect 76 297 149 321
rect 258 321 298 331
rect 76 255 86 297
rect -26 186 14 194
rect -26 118 -16 186
rect 4 118 14 186
rect -26 84 14 118
rect 46 186 86 255
rect 258 255 268 321
rect 288 255 298 321
rect 258 245 298 255
rect 323 321 426 331
rect 323 255 333 321
rect 353 297 426 321
rect 535 321 575 331
rect 353 255 363 297
rect 323 186 363 255
rect 535 255 545 321
rect 565 255 575 321
rect 535 245 575 255
rect 600 321 703 331
rect 600 255 610 321
rect 630 297 703 321
rect 630 255 640 297
rect 46 118 56 186
rect 76 118 86 186
rect 201 118 211 186
rect 231 118 261 186
rect 281 118 291 186
rect 46 108 86 118
rect -121 74 14 84
rect -121 54 -111 74
rect -91 64 14 74
rect -91 54 -81 64
rect -121 44 -81 54
rect -26 34 14 64
rect 41 84 81 89
rect 251 84 291 118
rect 323 118 333 186
rect 353 118 363 186
rect 323 108 363 118
rect 528 186 568 194
rect 528 118 538 186
rect 558 118 568 186
rect 41 64 51 84
rect 71 64 291 84
rect 41 59 81 64
rect -26 9 -16 34
rect 4 9 14 34
rect -26 -1 14 9
rect 46 34 86 42
rect 46 9 56 34
rect 76 9 86 34
rect -19 -62 21 -52
rect -19 -85 -9 -62
rect 11 -85 21 -62
rect -19 -95 21 -85
rect 46 -62 86 9
rect 251 34 291 64
rect 318 84 358 89
rect 528 84 568 118
rect 600 186 640 255
rect 600 118 610 186
rect 630 118 640 186
rect 600 108 640 118
rect 318 64 328 84
rect 348 64 568 84
rect 318 59 358 64
rect 251 9 261 34
rect 281 9 291 34
rect 251 -1 291 9
rect 323 34 363 42
rect 323 9 333 34
rect 353 9 363 34
rect 46 -85 56 -62
rect 76 -85 86 -62
rect 46 -156 86 -85
rect 258 -62 298 -52
rect 258 -85 268 -62
rect 288 -85 298 -62
rect 258 -95 298 -85
rect 323 -62 363 9
rect 528 34 568 64
rect 595 84 635 89
rect 595 64 605 84
rect 625 64 737 84
rect 595 59 635 64
rect 528 9 538 34
rect 558 9 568 34
rect 528 -1 568 9
rect 600 34 640 42
rect 600 9 610 34
rect 630 9 640 34
rect 323 -85 333 -62
rect 353 -85 363 -62
rect 323 -156 363 -85
rect 535 -62 575 -52
rect 535 -85 545 -62
rect 565 -85 575 -62
rect 535 -95 575 -85
rect 600 -62 640 9
rect 600 -85 610 -62
rect 630 -85 640 -62
rect -291 -236 -74 -156
rect -54 -236 -44 -156
rect -19 -236 -9 -156
rect 11 -236 21 -156
rect 46 -236 56 -156
rect 76 -236 86 -156
rect 208 -236 217 -156
rect 237 -236 268 -156
rect 288 -236 298 -156
rect 323 -236 333 -156
rect 353 -236 363 -156
rect 535 -156 575 -146
rect 535 -236 545 -156
rect 565 -236 575 -156
rect 600 -156 640 -85
rect 600 -236 610 -156
rect 630 -236 640 -156
rect 657 -255 677 64
rect -121 -265 677 -255
rect -121 -285 -111 -265
rect -91 -275 677 -265
rect -91 -285 -81 -275
rect -121 -295 -81 -285
<< end >>
