* PEX produced on Fri Feb 21 05:46:04 PM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from pfd_cp_lf_magic_3.ext - technology: sky130A

.subckt pfd_cp_lf_magic V_OUT VDDA GNDA F_REF F_VCO I_IN
X0 GNDA.t95 a_6200_5250.t2 a_6200_5250.t3 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X1 a_5970_4630.t6 V_OUT.t8 a_6200_5250.t0 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X2 GNDA.t137 GNDA.t135 GNDA.t137 GNDA.t136 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X3 pfd_8_0.DOWN_b.t1 VDDA.t130 pfd_8_0.DOWN_PFD_b.t3 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X4 a_870_1400.t1 pfd_8_0.QA_b.t3 VDDA.t126 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X5 pfd_8_0.UP_input.t3 pfd_8_0.UP_b.t1 sky130_fd_pr__cap_mim_m3_1 l=6.3 w=5.2
X6 pfd_8_0.DOWN.t2 pfd_8_0.DOWN_b.t2 VDDA.t55 VDDA.t30 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X7 VDDA.t27 pfd_8_0.opamp_out.t10 opamp_cell_4_0.VIN+.t4 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X8 opamp_cell_4_0.n_right.t1 opamp_cell_4_0.VIN+.t6 a_6320_5840.t8 GNDA.t148 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X9 opamp_cell_4_0.n_right.t3 opamp_cell_4_0.n_left.t6 VDDA.t71 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X10 pfd_8_0.opamp_out.t5 opamp_cell_4_0.n_right.t5 VDDA.t65 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X11 pfd_8_0.opamp_out.t9 a_6490_4630.t5 GNDA.t70 GNDA.t69 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X12 a_2350_1400.t0 pfd_8_0.before_Reset.t3 GNDA.t72 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X13 pfd_8_0.DOWN.t1 pfd_8_0.DOWN_b.t3 GNDA.t74 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X14 VDDA.t46 opamp_cell_4_0.p_bias.t7 opamp_cell_4_0.p_bias.t8 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X15 GNDA.t26 I_IN.t3 I_IN.t4 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X16 a_n30_1400.t0 F_REF.t0 VDDA.t129 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X17 GNDA.t153 pfd_8_0.QA.t3 pfd_8_0.QA_b.t2 GNDA.t152 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X18 a_6200_5250.t5 a_6200_5250.t4 GNDA.t93 GNDA.t92 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X19 a_6200_5250.t1 V_OUT.t9 a_5970_4630.t5 VDDA.t84 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X20 VDDA.t17 opamp_cell_4_0.p_bias.t9 a_5970_4630.t2 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X21 VDDA.t122 VDDA.t119 VDDA.t121 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X22 pfd_8_0.DOWN_input.t1 pfd_8_0.DOWN_b.t4 I_IN.t5 VDDA.t40 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X23 VDDA.t118 VDDA.t116 VDDA.t118 VDDA.t117 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X24 VDDA.t57 pfd_8_0.UP_input.t4 V_OUT.t3 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X25 a_1910_2020.t1 pfd_8_0.QB.t3 GNDA.t57 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X26 a_6220_5810.t8 a_6220_5810.t7 GNDA.t51 GNDA.t50 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X27 pfd_8_0.UP.t1 pfd_8_0.UP_PFD_b.t2 VDDA.t128 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X28 a_6320_5840.t12 a_6220_5810.t9 GNDA.t139 GNDA.t138 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X29 pfd_8_0.UP_input.t0 pfd_8_0.UP.t2 pfd_8_0.opamp_out.t0 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X30 pfd_8_0.QA.t2 pfd_8_0.QA_b.t4 GNDA.t76 GNDA.t75 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X31 a_5970_4630.t4 opamp_cell_4_0.p_bias.t10 VDDA.t44 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X32 pfd_8_0.DOWN_input.t0 pfd_8_0.DOWN.t3 I_IN.t0 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X33 a_1390_1400.t1 pfd_8_0.E.t3 pfd_8_0.E_b.t0 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X34 I_IN.t2 I_IN.t1 GNDA.t8 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X35 a_870_640.t0 pfd_8_0.QB_b.t3 VDDA.t21 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X36 VDDA.t115 VDDA.t112 VDDA.t114 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X37 pfd_8_0.opamp_out.t11 a_9360_3514.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X38 V_OUT.t4 loop_filter_2_0.R1_C1.t0 GNDA.t60 sky130_fd_pr__res_xhigh_po_0p35 l=7.52
X39 VDDA.t77 a_2530_190.t2 a_2200_190.t1 VDDA.t76 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X40 GNDA.t134 GNDA.t132 GNDA.t134 GNDA.t133 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0 ps=0 w=1.25 l=0.5
X41 GNDA.t131 GNDA.t128 GNDA.t130 GNDA.t129 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X42 opamp_cell_4_0.p_bias.t6 opamp_cell_4_0.p_bias.t5 VDDA.t19 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X43 VDDA.t111 VDDA.t109 VDDA.t111 VDDA.t110 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X44 V_OUT.t2 pfd_8_0.UP_input.t5 VDDA.t52 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X45 pfd_8_0.DOWN_input.t2 pfd_8_0.DOWN_b.t5 GNDA.t151 GNDA.t150 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X46 GNDA.t12 a_2530_190.t3 a_2200_190.t0 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X47 pfd_8_0.F.t0 pfd_8_0.QB_b.t4 GNDA.t47 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X48 GNDA.t127 GNDA.t124 GNDA.t126 GNDA.t125 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X49 GNDA.t123 GNDA.t120 GNDA.t122 GNDA.t121 sky130_fd_pr__nfet_01v8 ad=0.625 pd=3.5 as=0 ps=0 w=1.25 l=0.5
X50 pfd_8_0.opamp_out.t12 a_9360_6440.t1 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X51 pfd_8_0.UP_b.t2 pfd_8_0.UP.t3 GNDA.t143 GNDA.t142 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X52 GNDA.t145 pfd_8_0.E_b.t3 pfd_8_0.E.t2 GNDA.t144 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X53 GNDA.t39 a_6220_5810.t10 a_6320_5840.t7 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X54 GNDA.t119 GNDA.t116 GNDA.t118 GNDA.t117 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X55 a_1390_640.t0 pfd_8_0.F.t3 pfd_8_0.F_b.t0 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X56 a_2350_1400.t1 pfd_8_0.before_Reset.t4 VDDA.t75 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X57 GNDA.t83 a_6220_5810.t5 a_6220_5810.t6 GNDA.t82 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X58 GNDA.t115 GNDA.t112 GNDA.t114 GNDA.t113 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X59 GNDA.t111 GNDA.t109 GNDA.t111 GNDA.t110 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X60 a_5970_4630.t11 a_5970_4630.t10 a_5970_4630.t11 VDDA.t87 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X61 pfd_8_0.F_b.t1 pfd_8_0.F.t4 GNDA.t14 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X62 VDDA.t73 pfd_8_0.UP_input.t6 V_OUT.t6 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X63 GNDA.t156 loop_filter_2_0.R1_C1.t1 sky130_fd_pr__cap_mim_m3_1 l=60 w=69.8
X64 VDDA.t7 pfd_8_0.F.t5 a_490_640.t1 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X65 VDDA.t108 VDDA.t106 VDDA.t108 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X66 pfd_8_0.QA_b.t1 pfd_8_0.QA.t4 a_n30_1400.t1 VDDA.t80 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X67 GNDA.t108 GNDA.t106 GNDA.t108 GNDA.t107 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X68 GNDA.t78 pfd_8_0.F.t6 pfd_8_0.QB.t1 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X69 pfd_8_0.before_Reset.t2 pfd_8_0.QB.t4 VDDA.t54 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.805 ps=5 w=2 l=0.15
X70 GNDA.t68 a_6490_4630.t6 pfd_8_0.opamp_out.t8 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X71 VDDA.t63 opamp_cell_4_0.n_right.t6 pfd_8_0.opamp_out.t4 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X72 opamp_cell_4_0.VIN+.t3 pfd_8_0.opamp_out.t13 VDDA.t5 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X73 pfd_8_0.UP_input.t1 pfd_8_0.UP_b.t3 pfd_8_0.opamp_out.t1 VDDA.t40 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X74 a_490_1400.t1 pfd_8_0.QA_b.t5 pfd_8_0.QA.t1 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X75 V_OUT.t5 pfd_8_0.UP_input.t7 VDDA.t69 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X76 GNDA.t147 pfd_8_0.Reset.t2 pfd_8_0.E_b.t2 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X77 a_2530_190.t0 a_2350_1400.t2 GNDA.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X78 VDDA.t82 opamp_cell_4_0.n_left.t2 opamp_cell_4_0.n_left.t3 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X79 a_6320_5840.t10 V_OUT.t10 opamp_cell_4_0.n_left.t5 GNDA.t149 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X80 pfd_8_0.E.t0 pfd_8_0.E_b.t4 a_870_1400.t0 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X81 pfd_8_0.UP_b.t0 pfd_8_0.UP.t4 VDDA.t31 VDDA.t30 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X82 pfd_8_0.DOWN_input.t3 pfd_8_0.DOWN.t0 sky130_fd_pr__cap_mim_m3_1 l=3.8 w=2.7
X83 a_5970_4630.t9 a_5970_4630.t7 a_5970_4630.t8 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X84 GNDA.t105 GNDA.t102 GNDA.t104 GNDA.t103 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X85 VDDA.t48 a_1870_190.t2 pfd_8_0.Reset.t1 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X86 pfd_8_0.opamp_out.t7 a_6490_4630.t7 GNDA.t66 GNDA.t65 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X87 pfd_8_0.opamp_out.t3 opamp_cell_4_0.n_right.t7 VDDA.t61 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X88 GNDA.t16 a_1870_190.t3 pfd_8_0.Reset.t0 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X89 VDDA.t105 VDDA.t102 VDDA.t104 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X90 opamp_cell_4_0.p_bias.t4 opamp_cell_4_0.p_bias.t3 VDDA.t37 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X91 opamp_cell_4_0.p_bias.t0 a_6220_5810.t0 GNDA.t20 sky130_fd_pr__res_xhigh_po_5p73 l=1
X92 opamp_cell_4_0.n_left.t1 opamp_cell_4_0.n_left.t0 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X93 GNDA.t157 V_OUT.t7 sky130_fd_pr__cap_mim_m3_1 l=60 w=13.8
X94 opamp_cell_4_0.n_left.t4 V_OUT.t11 a_6320_5840.t11 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X95 a_5970_4630.t1 opamp_cell_4_0.p_bias.t11 VDDA.t15 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X96 pfd_8_0.before_Reset.t1 pfd_8_0.QA.t5 a_1910_2020.t0 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X97 pfd_8_0.UP_PFD_b.t0 pfd_8_0.QA.t6 GNDA.t30 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X98 GNDA.t45 pfd_8_0.E.t4 pfd_8_0.QA.t0 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X99 a_9360_6440.t0 a_6490_4630.t0 GNDA.t19 sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X100 VDDA.t101 VDDA.t99 VDDA.t101 VDDA.t100 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0 ps=0 w=2.5 l=0.5
X101 pfd_8_0.F.t1 pfd_8_0.F_b.t3 a_870_640.t1 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X102 VDDA.t33 pfd_8_0.Reset.t3 a_1390_1400.t0 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X103 GNDA.t101 GNDA.t99 GNDA.t101 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X104 a_2530_190.t1 a_2350_1400.t3 VDDA.t39 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X105 GNDA.t85 a_6220_5810.t3 a_6220_5810.t4 GNDA.t84 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X106 GNDA.t64 a_6490_4630.t8 pfd_8_0.opamp_out.t6 GNDA.t63 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X107 VDDA.t59 opamp_cell_4_0.n_right.t8 pfd_8_0.opamp_out.t2 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X108 VDDA.t98 VDDA.t95 VDDA.t97 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0 ps=0 w=2.5 l=0.5
X109 GNDA.t80 pfd_8_0.F_b.t4 pfd_8_0.F.t2 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X110 GNDA.t3 a_6220_5810.t11 a_6320_5840.t5 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X111 pfd_8_0.QB_b.t1 pfd_8_0.QB.t5 a_n30_640.t0 VDDA.t80 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X112 GNDA.t91 a_6200_5250.t6 a_6490_4630.t4 GNDA.t90 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X113 a_5970_4630.t12 opamp_cell_4_0.VIN+.t7 a_6490_4630.t2 VDDA.t127 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X114 VDDA.t13 opamp_cell_4_0.p_bias.t12 a_5970_4630.t0 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X115 VDDA.t78 pfd_8_0.Reset.t4 a_1390_640.t1 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X116 VDDA.t23 opamp_cell_4_0.p_bias.t1 opamp_cell_4_0.p_bias.t2 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X117 pfd_8_0.UP_input.t2 pfd_8_0.UP.t5 VDDA.t124 VDDA.t123 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X118 opamp_cell_4_0.n_right.t4 a_9360_3514.t1 GNDA.t81 sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X119 VDDA.t94 VDDA.t91 VDDA.t93 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X120 a_6320_5840.t4 a_6320_5840.t2 a_6320_5840.t3 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X121 GNDA.t1 pfd_8_0.QB.t6 pfd_8_0.QB_b.t2 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X122 a_6320_5840.t6 a_6220_5810.t12 GNDA.t37 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X123 GNDA.t62 pfd_8_0.Reset.t5 pfd_8_0.F_b.t2 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X124 GNDA.t28 pfd_8_0.DOWN_input.t4 V_OUT.t1 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X125 a_6320_5840.t1 a_6320_5840.t0 a_6320_5840.t1 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X126 VDDA.t90 VDDA.t88 VDDA.t90 VDDA.t89 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X127 a_6220_5810.t2 a_6220_5810.t1 GNDA.t87 GNDA.t86 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X128 GNDA.t141 I_IN.t6 opamp_cell_4_0.VIN+.t5 GNDA.t140 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X129 pfd_8_0.E.t1 pfd_8_0.QA_b.t6 GNDA.t22 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X130 VDDA.t25 pfd_8_0.QA.t7 pfd_8_0.before_Reset.t0 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X131 a_n30_640.t1 F_VCO.t0 VDDA.t67 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X132 pfd_8_0.UP_PFD_b.t1 pfd_8_0.QA.t8 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X133 a_6490_4630.t3 a_6200_5250.t7 GNDA.t89 GNDA.t88 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X134 a_6490_4630.t1 opamp_cell_4_0.VIN+.t8 a_5970_4630.t3 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X135 VDDA.t125 pfd_8_0.E.t5 a_490_1400.t0 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X136 VDDA.t42 a_2200_190.t2 a_1870_190.t1 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X137 pfd_8_0.QA_b.t0 F_REF.t1 GNDA.t59 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X138 pfd_8_0.QB_b.t0 F_VCO.t1 GNDA.t18 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X139 V_OUT.t0 pfd_8_0.DOWN_input.t5 GNDA.t10 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X140 a_490_640.t0 pfd_8_0.QB_b.t5 pfd_8_0.QB.t2 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X141 VDDA.t11 pfd_8_0.opamp_out.t14 opamp_cell_4_0.VIN+.t2 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X142 GNDA.t49 a_2200_190.t3 a_1870_190.t0 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X143 opamp_cell_4_0.VIN+.t0 I_IN.t7 GNDA.t24 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X144 a_6320_5840.t9 opamp_cell_4_0.VIN+.t9 opamp_cell_4_0.n_right.t0 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X145 VDDA.t50 opamp_cell_4_0.n_left.t7 opamp_cell_4_0.n_right.t2 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X146 pfd_8_0.QB.t0 pfd_8_0.QB_b.t6 GNDA.t43 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X147 pfd_8_0.DOWN_PFD_b.t1 pfd_8_0.QB.t7 VDDA.t79 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X148 pfd_8_0.UP.t0 pfd_8_0.UP_PFD_b.t3 GNDA.t155 GNDA.t154 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X149 GNDA.t98 GNDA.t96 GNDA.t98 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X150 pfd_8_0.DOWN_PFD_b.t0 pfd_8_0.QB.t8 GNDA.t32 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X151 pfd_8_0.E_b.t1 pfd_8_0.E.t6 GNDA.t41 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X152 opamp_cell_4_0.VIN+.t1 pfd_8_0.opamp_out.t15 VDDA.t35 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X153 pfd_8_0.DOWN_b.t0 GNDA.t158 pfd_8_0.DOWN_PFD_b.t2 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
R0 a_6200_5250.n5 a_6200_5250.n4 427.647
R1 a_6200_5250.n1 a_6200_5250.t6 321.334
R2 a_6200_5250.n4 a_6200_5250.n0 210.601
R3 a_6200_5250.n2 a_6200_5250.n1 208.868
R4 a_6200_5250.n3 a_6200_5250.t4 174.056
R5 a_6200_5250.n4 a_6200_5250.n3 152
R6 a_6200_5250.n1 a_6200_5250.t7 112.468
R7 a_6200_5250.n2 a_6200_5250.t2 112.468
R8 a_6200_5250.n3 a_6200_5250.n2 61.5894
R9 a_6200_5250.n0 a_6200_5250.t3 60.0005
R10 a_6200_5250.n0 a_6200_5250.t5 60.0005
R11 a_6200_5250.t0 a_6200_5250.n5 49.2505
R12 a_6200_5250.n5 a_6200_5250.t1 49.2505
R13 GNDA.n397 GNDA.n396 348175
R14 GNDA.n396 GNDA.n395 292776
R15 GNDA.n348 GNDA.t35 25257.7
R16 GNDA.n348 GNDA.n148 15376.3
R17 GNDA.n395 GNDA.t150 2083.03
R18 GNDA.t13 GNDA.t79 1939.79
R19 GNDA.t42 GNDA.t0 1939.79
R20 GNDA.n186 GNDA.n24 1860.65
R21 GNDA.t34 GNDA.t31 1845.16
R22 GNDA.t73 GNDA.t55 1372.04
R23 GNDA.t15 GNDA.n400 1253.76
R24 GNDA.n403 GNDA.n23 1230.11
R25 GNDA.n340 GNDA.n339 1186
R26 GNDA.n185 GNDA.n184 1186
R27 GNDA.n178 GNDA.n177 1186
R28 GNDA.n347 GNDA.n346 1186
R29 GNDA.n350 GNDA.n349 1170
R30 GNDA.n394 GNDA.t55 1064.52
R31 GNDA.n357 GNDA.t34 1064.52
R32 GNDA.n395 GNDA.n26 1052.76
R33 GNDA.t11 GNDA.n402 922.582
R34 GNDA.t48 GNDA.n401 922.582
R35 GNDA.n232 GNDA.t58 783.001
R36 GNDA.t150 GNDA.n394 780.645
R37 GNDA.n357 GNDA.t73 780.645
R38 GNDA.t31 GNDA.n23 780.645
R39 GNDA.n99 GNDA.n98 669.307
R40 GNDA.n102 GNDA.n101 669.307
R41 GNDA.n120 GNDA.n119 669.307
R42 GNDA.n123 GNDA.n122 669.307
R43 GNDA.n147 GNDA.n146 669.307
R44 GNDA.n141 GNDA.n28 669.307
R45 GNDA.n403 GNDA.t11 638.711
R46 GNDA.n402 GNDA.t48 638.711
R47 GNDA.n401 GNDA.t15 638.711
R48 GNDA.n400 GNDA.t61 638.711
R49 GNDA.t46 GNDA.n399 638.711
R50 GNDA.n399 GNDA.t77 638.711
R51 GNDA.t17 GNDA.n397 638.711
R52 GNDA.t144 GNDA.t40 601.333
R53 GNDA.t152 GNDA.t75 601.333
R54 GNDA.t27 GNDA.t100 593.865
R55 GNDA.t9 GNDA.t27 593.865
R56 GNDA.t125 GNDA.t9 593.865
R57 GNDA.t140 GNDA.t97 593.865
R58 GNDA.t23 GNDA.t140 593.865
R59 GNDA.t117 GNDA.t23 593.865
R60 GNDA.t136 GNDA.t25 593.865
R61 GNDA.t25 GNDA.t7 593.865
R62 GNDA.t7 GNDA.t113 593.865
R63 GNDA.n231 GNDA.n230 585.003
R64 GNDA.n399 GNDA.n398 585.003
R65 GNDA.n228 GNDA.n227 585.001
R66 GNDA.n226 GNDA.n225 585.001
R67 GNDA.n224 GNDA.n223 585.001
R68 GNDA.n205 GNDA.n25 585.001
R69 GNDA.n338 GNDA.n337 585.001
R70 GNDA.n187 GNDA.n186 585.001
R71 GNDA.n197 GNDA.n196 585.001
R72 GNDA.n199 GNDA.n198 585.001
R73 GNDA.n201 GNDA.n200 585.001
R74 GNDA.n394 GNDA.n393 585.001
R75 GNDA.n358 GNDA.n357 585.001
R76 GNDA.n363 GNDA.n23 585.001
R77 GNDA.n404 GNDA.n403 585.001
R78 GNDA.n402 GNDA.n19 585.001
R79 GNDA.n401 GNDA.n16 585.001
R80 GNDA.n400 GNDA.n13 585.001
R81 GNDA.n397 GNDA.n2 585.001
R82 GNDA.n145 GNDA.n29 585
R83 GNDA.n143 GNDA.n142 585
R84 GNDA.n44 GNDA.n40 585
R85 GNDA.n42 GNDA.n39 585
R86 GNDA.n61 GNDA.n57 585
R87 GNDA.n59 GNDA.n56 585
R88 GNDA.n72 GNDA.n71 585
R89 GNDA.n71 GNDA.n26 585
R90 GNDA.n75 GNDA.n74 585
R91 GNDA.n77 GNDA.n69 585
R92 GNDA.n79 GNDA.n78 585
R93 GNDA.n78 GNDA.n26 585
R94 GNDA.n376 GNDA.t158 566.966
R95 GNDA.n148 GNDA.t100 566.871
R96 GNDA.n121 GNDA.t125 566.871
R97 GNDA.n121 GNDA.t97 566.871
R98 GNDA.n100 GNDA.t117 566.871
R99 GNDA.n100 GNDA.t136 566.871
R100 GNDA.t113 GNDA.n26 566.871
R101 GNDA.t19 GNDA.n347 564.696
R102 GNDA.n348 GNDA.t81 534.24
R103 GNDA.t61 GNDA.t13 520.431
R104 GNDA.t79 GNDA.t46 520.431
R105 GNDA.t77 GNDA.t42 520.431
R106 GNDA.t0 GNDA.t17 520.431
R107 GNDA.t81 GNDA.t19 509.197
R108 GNDA.t142 GNDA.t35 425.334
R109 GNDA.n200 GNDA.t4 418
R110 GNDA.t154 GNDA.n197 344.668
R111 GNDA.t29 GNDA.n199 344.668
R112 GNDA.n58 GNDA.t135 336.329
R113 GNDA.n58 GNDA.t116 336.329
R114 GNDA.n41 GNDA.t96 336.329
R115 GNDA.n41 GNDA.t124 336.329
R116 GNDA.n349 GNDA.n348 331.702
R117 GNDA.n80 GNDA.t112 320.7
R118 GNDA.n140 GNDA.t99 320.7
R119 GNDA.n149 GNDA.t106 304.634
R120 GNDA.n341 GNDA.t128 304.634
R121 GNDA.n183 GNDA.t102 304.634
R122 GNDA.n179 GNDA.t109 304.634
R123 GNDA.n336 GNDA.t132 292.584
R124 GNDA.n188 GNDA.t120 292.584
R125 GNDA.t71 GNDA.n25 286
R126 GNDA.t33 GNDA.n224 286
R127 GNDA.n148 GNDA.n147 250.349
R128 GNDA.n148 GNDA.n28 250.349
R129 GNDA.n121 GNDA.n120 250.349
R130 GNDA.n122 GNDA.n121 250.349
R131 GNDA.n100 GNDA.n99 250.349
R132 GNDA.n101 GNDA.n100 250.349
R133 GNDA.n76 GNDA.n26 250.349
R134 GNDA.n346 GNDA.t108 245
R135 GNDA.n340 GNDA.t131 245
R136 GNDA.n184 GNDA.t105 245
R137 GNDA.n178 GNDA.t111 245
R138 GNDA.n197 GNDA.t142 227.333
R139 GNDA.n199 GNDA.t154 227.333
R140 GNDA.n200 GNDA.t29 227.333
R141 GNDA.n228 GNDA.n226 205.333
R142 GNDA.n343 GNDA.n151 204.201
R143 GNDA.n181 GNDA.n175 204.201
R144 GNDA.n182 GNDA.n174 204.201
R145 GNDA.n180 GNDA.n176 204.201
R146 GNDA.n342 GNDA.n152 204.201
R147 GNDA.n345 GNDA.n344 204.201
R148 GNDA.n3 GNDA.t1 198.058
R149 GNDA.n445 GNDA.t43 198.058
R150 GNDA.n433 GNDA.t80 198.058
R151 GNDA.n11 GNDA.t14 198.058
R152 GNDA.n257 GNDA.t41 198.058
R153 GNDA.n252 GNDA.t145 198.058
R154 GNDA.n220 GNDA.t76 198.058
R155 GNDA.n238 GNDA.t153 198.058
R156 GNDA.n224 GNDA.t71 198
R157 GNDA.n226 GNDA.t56 198
R158 GNDA.t146 GNDA.n228 198
R159 GNDA.n231 GNDA.t21 198
R160 GNDA.t44 GNDA.n231 198
R161 GNDA.n57 GNDA.n56 197
R162 GNDA.n40 GNDA.n39 197
R163 GNDA.n142 GNDA.n29 197
R164 GNDA.n75 GNDA.n71 197
R165 GNDA.n78 GNDA.n77 197
R166 GNDA.n98 GNDA.n55 185
R167 GNDA.n102 GNDA.n55 185
R168 GNDA.n119 GNDA.n38 185
R169 GNDA.n123 GNDA.n38 185
R170 GNDA.n146 GNDA.n30 185
R171 GNDA.n141 GNDA.n30 185
R172 GNDA.n72 GNDA.n70 185
R173 GNDA.n79 GNDA.n70 185
R174 GNDA.n98 GNDA.n58 166.63
R175 GNDA.n119 GNDA.n41 166.63
R176 GNDA.n351 GNDA.n350 166.119
R177 GNDA.t56 GNDA.t33 161.333
R178 GNDA.t40 GNDA.t146 161.333
R179 GNDA.t21 GNDA.t144 161.333
R180 GNDA.t75 GNDA.t44 161.333
R181 GNDA.t58 GNDA.t152 161.333
R182 GNDA.n337 GNDA.t134 134.501
R183 GNDA.n187 GNDA.t123 134.501
R184 GNDA.n7 GNDA.t78 130.713
R185 GNDA.n232 GNDA.t59 130.001
R186 GNDA.n227 GNDA.t147 130.001
R187 GNDA.n225 GNDA.t57 130.001
R188 GNDA.n223 GNDA.t72 130.001
R189 GNDA.n205 GNDA.t5 130.001
R190 GNDA.n2 GNDA.t18 130.001
R191 GNDA.n13 GNDA.t62 130.001
R192 GNDA.n16 GNDA.t16 130.001
R193 GNDA.n19 GNDA.t49 130.001
R194 GNDA.n404 GNDA.t12 130.001
R195 GNDA.n229 GNDA.t22 130.001
R196 GNDA.n219 GNDA.t45 130.001
R197 GNDA.n8 GNDA.t47 130.001
R198 GNDA.n201 GNDA.t30 122.501
R199 GNDA.n198 GNDA.t155 122.501
R200 GNDA.n196 GNDA.t143 122.501
R201 GNDA.n363 GNDA.t32 122.501
R202 GNDA.n358 GNDA.t74 122.501
R203 GNDA.n393 GNDA.t151 122.501
R204 GNDA.n338 GNDA.t54 112.451
R205 GNDA.n156 GNDA.n155 97.8707
R206 GNDA.n160 GNDA.n159 97.8707
R207 GNDA.n164 GNDA.n163 97.8707
R208 GNDA.n168 GNDA.n167 97.8707
R209 GNDA.n173 GNDA.n172 97.8707
R210 GNDA.n177 GNDA.t50 97.7783
R211 GNDA.n339 GNDA.t129 95.1512
R212 GNDA.n347 GNDA.t107 94.9025
R213 GNDA.n130 GNDA.n129 92.2612
R214 GNDA.n138 GNDA.n137 92.2612
R215 GNDA.n116 GNDA.n115 92.2612
R216 GNDA.n109 GNDA.n50 92.2612
R217 GNDA.n95 GNDA.n94 92.2612
R218 GNDA.n88 GNDA.n68 92.2612
R219 GNDA.n60 GNDA.n55 91.3721
R220 GNDA.n97 GNDA.n96 91.3721
R221 GNDA.n96 GNDA.n54 91.3721
R222 GNDA.n43 GNDA.n38 91.3721
R223 GNDA.n118 GNDA.n117 91.3721
R224 GNDA.n117 GNDA.n37 91.3721
R225 GNDA.n144 GNDA.n30 90.7567
R226 GNDA.n73 GNDA.n70 90.7567
R227 GNDA.t50 GNDA.t53 89.1508
R228 GNDA.n185 GNDA.t121 86.275
R229 GNDA.n350 GNDA.t157 86.0829
R230 GNDA.n147 GNDA.n29 84.306
R231 GNDA.n142 GNDA.n28 84.306
R232 GNDA.n120 GNDA.n40 84.306
R233 GNDA.n122 GNDA.n39 84.306
R234 GNDA.n99 GNDA.n57 84.306
R235 GNDA.n101 GNDA.n56 84.306
R236 GNDA.n76 GNDA.n75 84.306
R237 GNDA.n77 GNDA.n76 84.306
R238 GNDA.n181 GNDA.n180 83.2005
R239 GNDA.n182 GNDA.n181 83.2005
R240 GNDA.n350 GNDA.t156 82.8829
R241 GNDA.n396 GNDA.n24 80.6672
R242 GNDA.t82 GNDA.t110 77.6476
R243 GNDA.n339 GNDA.n338 74.9677
R244 GNDA.t129 GNDA.t69 74.8697
R245 GNDA.t67 GNDA.t107 74.7717
R246 GNDA.t65 GNDA.t67 74.7717
R247 GNDA.t63 GNDA.t65 74.7717
R248 GNDA.t69 GNDA.t63 74.7717
R249 GNDA.t149 GNDA.t148 74.7717
R250 GNDA.t90 GNDA.t88 74.7717
R251 GNDA.t92 GNDA.t103 74.7717
R252 GNDA.n396 GNDA.n25 73.3338
R253 GNDA.t6 GNDA.t133 72.0844
R254 GNDA.t38 GNDA.t94 71.8959
R255 GNDA.n344 GNDA.n343 66.5605
R256 GNDA.n343 GNDA.n342 66.5605
R257 GNDA.t52 GNDA.t138 66.1443
R258 GNDA.n343 GNDA.n150 65.9634
R259 GNDA.n233 GNDA.n232 60.29
R260 GNDA.n227 GNDA.n212 60.29
R261 GNDA.n225 GNDA.n211 60.29
R262 GNDA.n223 GNDA.n208 60.29
R263 GNDA.n276 GNDA.n205 60.29
R264 GNDA.n405 GNDA.n404 60.29
R265 GNDA.n412 GNDA.n19 60.29
R266 GNDA.n418 GNDA.n16 60.29
R267 GNDA.n425 GNDA.n13 60.29
R268 GNDA.n453 GNDA.n2 60.29
R269 GNDA.n151 GNDA.t66 60.0005
R270 GNDA.n151 GNDA.t64 60.0005
R271 GNDA.n175 GNDA.t89 60.0005
R272 GNDA.n175 GNDA.t95 60.0005
R273 GNDA.n174 GNDA.t93 60.0005
R274 GNDA.n174 GNDA.t104 60.0005
R275 GNDA.t111 GNDA.n176 60.0005
R276 GNDA.n176 GNDA.t91 60.0005
R277 GNDA.n152 GNDA.t70 60.0005
R278 GNDA.n152 GNDA.t130 60.0005
R279 GNDA.t108 GNDA.n345 60.0005
R280 GNDA.n345 GNDA.t68 60.0005
R281 GNDA.n202 GNDA.n201 59.5478
R282 GNDA.n198 GNDA.n192 59.5478
R283 GNDA.n196 GNDA.n190 59.5478
R284 GNDA.n381 GNDA.n358 58.9809
R285 GNDA.n364 GNDA.n363 58.9809
R286 GNDA.n393 GNDA.n392 58.9809
R287 GNDA.n246 GNDA.n219 54.4005
R288 GNDA.n229 GNDA.n218 54.4005
R289 GNDA.n438 GNDA.n8 54.4005
R290 GNDA.n440 GNDA.n7 54.4005
R291 GNDA.t84 GNDA.t52 48.8894
R292 GNDA.t4 GNDA.n24 44.0005
R293 GNDA.t94 GNDA.t36 43.1378
R294 GNDA.n181 GNDA.n170 41.6005
R295 GNDA.n83 GNDA.n82 41.3005
R296 GNDA.t2 GNDA.t6 40.3637
R297 GNDA.n333 GNDA.n150 39.4985
R298 GNDA.t110 GNDA.t86 37.3861
R299 GNDA.t86 GNDA.t90 37.3861
R300 GNDA.n349 GNDA.t60 34.0494
R301 GNDA.n233 GNDA.n0 33.0991
R302 GNDA.n454 GNDA.n453 33.0991
R303 GNDA.n130 GNDA.n128 32.0005
R304 GNDA.n128 GNDA.n34 32.0005
R305 GNDA.n136 GNDA.n135 32.0005
R306 GNDA.n135 GNDA.n32 32.0005
R307 GNDA.n131 GNDA.n32 32.0005
R308 GNDA.n45 GNDA.n36 32.0005
R309 GNDA.n114 GNDA.n48 32.0005
R310 GNDA.n110 GNDA.n48 32.0005
R311 GNDA.n110 GNDA.n109 32.0005
R312 GNDA.n108 GNDA.n51 32.0005
R313 GNDA.n104 GNDA.n51 32.0005
R314 GNDA.n103 GNDA.n53 32.0005
R315 GNDA.n62 GNDA.n53 32.0005
R316 GNDA.n93 GNDA.n66 32.0005
R317 GNDA.n89 GNDA.n66 32.0005
R318 GNDA.n87 GNDA.n81 32.0005
R319 GNDA.n294 GNDA.n190 32.0005
R320 GNDA.n294 GNDA.n293 32.0005
R321 GNDA.n293 GNDA.n292 32.0005
R322 GNDA.n289 GNDA.n288 32.0005
R323 GNDA.n288 GNDA.n287 32.0005
R324 GNDA.n287 GNDA.n194 32.0005
R325 GNDA.n283 GNDA.n282 32.0005
R326 GNDA.n282 GNDA.n281 32.0005
R327 GNDA.n281 GNDA.n203 32.0005
R328 GNDA.n277 GNDA.n203 32.0005
R329 GNDA.n275 GNDA.n274 32.0005
R330 GNDA.n274 GNDA.n206 32.0005
R331 GNDA.n270 GNDA.n269 32.0005
R332 GNDA.n269 GNDA.n268 32.0005
R333 GNDA.n268 GNDA.n209 32.0005
R334 GNDA.n264 GNDA.n263 32.0005
R335 GNDA.n263 GNDA.n262 32.0005
R336 GNDA.n259 GNDA.n258 32.0005
R337 GNDA.n258 GNDA.n257 32.0005
R338 GNDA.n257 GNDA.n214 32.0005
R339 GNDA.n253 GNDA.n214 32.0005
R340 GNDA.n253 GNDA.n252 32.0005
R341 GNDA.n252 GNDA.n251 32.0005
R342 GNDA.n251 GNDA.n216 32.0005
R343 GNDA.n245 GNDA.n244 32.0005
R344 GNDA.n244 GNDA.n220 32.0005
R345 GNDA.n240 GNDA.n220 32.0005
R346 GNDA.n240 GNDA.n239 32.0005
R347 GNDA.n239 GNDA.n238 32.0005
R348 GNDA.n238 GNDA.n222 32.0005
R349 GNDA.n234 GNDA.n222 32.0005
R350 GNDA.n333 GNDA.n332 32.0005
R351 GNDA.n332 GNDA.n331 32.0005
R352 GNDA.n331 GNDA.n154 32.0005
R353 GNDA.n327 GNDA.n154 32.0005
R354 GNDA.n327 GNDA.n326 32.0005
R355 GNDA.n326 GNDA.n325 32.0005
R356 GNDA.n325 GNDA.n158 32.0005
R357 GNDA.n321 GNDA.n158 32.0005
R358 GNDA.n321 GNDA.n320 32.0005
R359 GNDA.n320 GNDA.n319 32.0005
R360 GNDA.n319 GNDA.n162 32.0005
R361 GNDA.n315 GNDA.n162 32.0005
R362 GNDA.n315 GNDA.n314 32.0005
R363 GNDA.n314 GNDA.n313 32.0005
R364 GNDA.n313 GNDA.n166 32.0005
R365 GNDA.n309 GNDA.n308 32.0005
R366 GNDA.n308 GNDA.n307 32.0005
R367 GNDA.n307 GNDA.n171 32.0005
R368 GNDA.n302 GNDA.n171 32.0005
R369 GNDA.n302 GNDA.n301 32.0005
R370 GNDA.n301 GNDA.n300 32.0005
R371 GNDA.n391 GNDA.n353 32.0005
R372 GNDA.n387 GNDA.n353 32.0005
R373 GNDA.n387 GNDA.n386 32.0005
R374 GNDA.n386 GNDA.n385 32.0005
R375 GNDA.n385 GNDA.n355 32.0005
R376 GNDA.n381 GNDA.n355 32.0005
R377 GNDA.n381 GNDA.n380 32.0005
R378 GNDA.n380 GNDA.n379 32.0005
R379 GNDA.n379 GNDA.n359 32.0005
R380 GNDA.n374 GNDA.n359 32.0005
R381 GNDA.n374 GNDA.n373 32.0005
R382 GNDA.n373 GNDA.n372 32.0005
R383 GNDA.n372 GNDA.n361 32.0005
R384 GNDA.n368 GNDA.n367 32.0005
R385 GNDA.n367 GNDA.n366 32.0005
R386 GNDA.n366 GNDA.n22 32.0005
R387 GNDA.n406 GNDA.n22 32.0005
R388 GNDA.n410 GNDA.n20 32.0005
R389 GNDA.n411 GNDA.n410 32.0005
R390 GNDA.n413 GNDA.n17 32.0005
R391 GNDA.n417 GNDA.n17 32.0005
R392 GNDA.n420 GNDA.n419 32.0005
R393 GNDA.n420 GNDA.n14 32.0005
R394 GNDA.n424 GNDA.n14 32.0005
R395 GNDA.n427 GNDA.n426 32.0005
R396 GNDA.n427 GNDA.n11 32.0005
R397 GNDA.n431 GNDA.n11 32.0005
R398 GNDA.n432 GNDA.n431 32.0005
R399 GNDA.n433 GNDA.n432 32.0005
R400 GNDA.n433 GNDA.n9 32.0005
R401 GNDA.n437 GNDA.n9 32.0005
R402 GNDA.n441 GNDA.n5 32.0005
R403 GNDA.n445 GNDA.n5 32.0005
R404 GNDA.n446 GNDA.n445 32.0005
R405 GNDA.n447 GNDA.n446 32.0005
R406 GNDA.n447 GNDA.n3 32.0005
R407 GNDA.n451 GNDA.n3 32.0005
R408 GNDA.n452 GNDA.n451 32.0005
R409 GNDA.t148 GNDA.t2 31.6345
R410 GNDA.n103 GNDA.n102 29.0291
R411 GNDA.n124 GNDA.n123 29.0291
R412 GNDA.n292 GNDA.n192 28.8005
R413 GNDA.n276 GNDA.n275 28.8005
R414 GNDA.n186 GNDA.n185 28.7587
R415 GNDA.n341 GNDA.n340 27.2005
R416 GNDA.n346 GNDA.n149 27.2005
R417 GNDA.t53 GNDA.t84 25.8829
R418 GNDA.n124 GNDA.n36 25.6005
R419 GNDA.n94 GNDA.n93 25.6005
R420 GNDA.n89 GNDA.n88 25.6005
R421 GNDA.n202 GNDA.n194 25.6005
R422 GNDA.n211 GNDA.n209 25.6005
R423 GNDA.n262 GNDA.n212 25.6005
R424 GNDA.n247 GNDA.n218 25.6005
R425 GNDA.n247 GNDA.n246 25.6005
R426 GNDA.n184 GNDA.n183 25.6005
R427 GNDA.n179 GNDA.n178 25.6005
R428 GNDA.n309 GNDA.n170 25.6005
R429 GNDA.n300 GNDA 25.6005
R430 GNDA.n392 GNDA.n391 25.6005
R431 GNDA.n364 GNDA.n361 25.6005
R432 GNDA.n405 GNDA.n20 25.6005
R433 GNDA.n418 GNDA.n417 25.6005
R434 GNDA.n425 GNDA.n424 25.6005
R435 GNDA.n439 GNDA.n438 25.6005
R436 GNDA.n337 GNDA.n336 24.8279
R437 GNDA.n188 GNDA.n187 24.8279
R438 GNDA.n155 GNDA.t134 24.0005
R439 GNDA.n155 GNDA.t3 24.0005
R440 GNDA.n159 GNDA.t139 24.0005
R441 GNDA.n159 GNDA.t85 24.0005
R442 GNDA.n163 GNDA.t51 24.0005
R443 GNDA.n163 GNDA.t83 24.0005
R444 GNDA.n167 GNDA.t87 24.0005
R445 GNDA.n167 GNDA.t39 24.0005
R446 GNDA.n172 GNDA.t37 24.0005
R447 GNDA.n172 GNDA.t122 24.0005
R448 GNDA.n440 GNDA.n439 22.4005
R449 GNDA.n140 GNDA.n139 20.9665
R450 GNDA.n115 GNDA.n45 19.2005
R451 GNDA.n115 GNDA.n114 19.2005
R452 GNDA.n270 GNDA.n208 19.2005
R453 GNDA.t20 GNDA.t92 17.8306
R454 GNDA.n177 GNDA.t82 17.2554
R455 GNDA.n412 GNDA.n411 16.0005
R456 GNDA.n413 GNDA.n412 16.0005
R457 GNDA.n298 GNDA 15.7005
R458 GNDA.n141 GNDA.n140 15.6449
R459 GNDA.n80 GNDA.n79 15.6449
R460 GNDA.n129 GNDA.t10 15.0005
R461 GNDA.n129 GNDA.t126 15.0005
R462 GNDA.n137 GNDA.t101 15.0005
R463 GNDA.n137 GNDA.t28 15.0005
R464 GNDA.t98 GNDA.n116 15.0005
R465 GNDA.n116 GNDA.t141 15.0005
R466 GNDA.n50 GNDA.t24 15.0005
R467 GNDA.n50 GNDA.t118 15.0005
R468 GNDA.t137 GNDA.n95 15.0005
R469 GNDA.n95 GNDA.t26 15.0005
R470 GNDA.n68 GNDA.t8 15.0005
R471 GNDA.n68 GNDA.t114 15.0005
R472 GNDA.n96 GNDA.t137 15.0005
R473 GNDA.n55 GNDA.t119 15.0005
R474 GNDA.n117 GNDA.t98 15.0005
R475 GNDA.n38 GNDA.t127 15.0005
R476 GNDA.t101 GNDA.n30 15.0005
R477 GNDA.n70 GNDA.t115 15.0005
R478 GNDA.n81 GNDA.n80 14.4005
R479 GNDA.n342 GNDA.n341 14.0805
R480 GNDA.n344 GNDA.n149 14.0805
R481 GNDA.n392 GNDA.n352 13.9181
R482 GNDA.t36 GNDA.t20 13.8044
R483 GNDA.n298 GNDA.n297 13.1958
R484 GNDA.n297 GNDA.n296 12.8163
R485 GNDA.n124 GNDA.n34 12.8005
R486 GNDA.n138 GNDA.n136 12.8005
R487 GNDA.n94 GNDA.n62 12.8005
R488 GNDA.n88 GNDA.n87 12.8005
R489 GNDA.n208 GNDA.n206 12.8005
R490 GNDA.n183 GNDA.n182 12.8005
R491 GNDA.n180 GNDA.n179 12.8005
R492 GNDA GNDA.n0 12.7806
R493 GNDA GNDA.n454 11.8829
R494 GNDA.n352 GNDA.n351 11.7212
R495 GNDA.n82 GNDA.n27 11.6542
R496 GNDA.n441 GNDA.n440 9.6005
R497 GNDA.n336 GNDA.n335 9.58175
R498 GNDA.n304 GNDA.n188 9.58175
R499 GNDA.n248 GNDA.n247 9.3005
R500 GNDA.n235 GNDA.n234 9.3005
R501 GNDA.n236 GNDA.n222 9.3005
R502 GNDA.n238 GNDA.n237 9.3005
R503 GNDA.n239 GNDA.n221 9.3005
R504 GNDA.n241 GNDA.n240 9.3005
R505 GNDA.n242 GNDA.n220 9.3005
R506 GNDA.n244 GNDA.n243 9.3005
R507 GNDA.n245 GNDA.n217 9.3005
R508 GNDA.n249 GNDA.n216 9.3005
R509 GNDA.n251 GNDA.n250 9.3005
R510 GNDA.n252 GNDA.n215 9.3005
R511 GNDA.n254 GNDA.n253 9.3005
R512 GNDA.n255 GNDA.n214 9.3005
R513 GNDA.n257 GNDA.n256 9.3005
R514 GNDA.n258 GNDA.n213 9.3005
R515 GNDA.n260 GNDA.n259 9.3005
R516 GNDA.n262 GNDA.n261 9.3005
R517 GNDA.n263 GNDA.n210 9.3005
R518 GNDA.n265 GNDA.n264 9.3005
R519 GNDA.n266 GNDA.n209 9.3005
R520 GNDA.n268 GNDA.n267 9.3005
R521 GNDA.n269 GNDA.n207 9.3005
R522 GNDA.n271 GNDA.n270 9.3005
R523 GNDA.n272 GNDA.n206 9.3005
R524 GNDA.n274 GNDA.n273 9.3005
R525 GNDA.n275 GNDA.n204 9.3005
R526 GNDA.n278 GNDA.n277 9.3005
R527 GNDA.n279 GNDA.n203 9.3005
R528 GNDA.n281 GNDA.n280 9.3005
R529 GNDA.n282 GNDA.n195 9.3005
R530 GNDA.n284 GNDA.n283 9.3005
R531 GNDA.n285 GNDA.n194 9.3005
R532 GNDA.n287 GNDA.n286 9.3005
R533 GNDA.n288 GNDA.n193 9.3005
R534 GNDA.n290 GNDA.n289 9.3005
R535 GNDA.n292 GNDA.n291 9.3005
R536 GNDA.n293 GNDA.n191 9.3005
R537 GNDA.n295 GNDA.n294 9.3005
R538 GNDA.n334 GNDA.n333 9.3005
R539 GNDA.n332 GNDA.n153 9.3005
R540 GNDA.n331 GNDA.n330 9.3005
R541 GNDA.n329 GNDA.n154 9.3005
R542 GNDA.n328 GNDA.n327 9.3005
R543 GNDA.n326 GNDA.n157 9.3005
R544 GNDA.n325 GNDA.n324 9.3005
R545 GNDA.n323 GNDA.n158 9.3005
R546 GNDA.n322 GNDA.n321 9.3005
R547 GNDA.n320 GNDA.n161 9.3005
R548 GNDA.n319 GNDA.n318 9.3005
R549 GNDA.n317 GNDA.n162 9.3005
R550 GNDA.n316 GNDA.n315 9.3005
R551 GNDA.n314 GNDA.n165 9.3005
R552 GNDA.n313 GNDA.n312 9.3005
R553 GNDA.n311 GNDA.n166 9.3005
R554 GNDA.n310 GNDA.n309 9.3005
R555 GNDA.n308 GNDA.n169 9.3005
R556 GNDA.n307 GNDA.n306 9.3005
R557 GNDA.n305 GNDA.n171 9.3005
R558 GNDA.n303 GNDA.n302 9.3005
R559 GNDA.n301 GNDA.n189 9.3005
R560 GNDA.n300 GNDA.n299 9.3005
R561 GNDA.n84 GNDA.n83 9.3005
R562 GNDA.n85 GNDA.n81 9.3005
R563 GNDA.n87 GNDA.n86 9.3005
R564 GNDA.n88 GNDA.n67 9.3005
R565 GNDA.n90 GNDA.n89 9.3005
R566 GNDA.n91 GNDA.n66 9.3005
R567 GNDA.n93 GNDA.n92 9.3005
R568 GNDA.n94 GNDA.n65 9.3005
R569 GNDA.n64 GNDA.n62 9.3005
R570 GNDA.n63 GNDA.n53 9.3005
R571 GNDA.n103 GNDA.n52 9.3005
R572 GNDA.n136 GNDA.n31 9.3005
R573 GNDA.n135 GNDA.n134 9.3005
R574 GNDA.n133 GNDA.n32 9.3005
R575 GNDA.n132 GNDA.n131 9.3005
R576 GNDA.n130 GNDA.n33 9.3005
R577 GNDA.n128 GNDA.n127 9.3005
R578 GNDA.n126 GNDA.n34 9.3005
R579 GNDA.n125 GNDA.n124 9.3005
R580 GNDA.n36 GNDA.n35 9.3005
R581 GNDA.n46 GNDA.n45 9.3005
R582 GNDA.n115 GNDA.n47 9.3005
R583 GNDA.n114 GNDA.n113 9.3005
R584 GNDA.n112 GNDA.n48 9.3005
R585 GNDA.n111 GNDA.n110 9.3005
R586 GNDA.n109 GNDA.n49 9.3005
R587 GNDA.n108 GNDA.n107 9.3005
R588 GNDA.n106 GNDA.n51 9.3005
R589 GNDA.n105 GNDA.n104 9.3005
R590 GNDA.n391 GNDA.n390 9.3005
R591 GNDA.n389 GNDA.n353 9.3005
R592 GNDA.n388 GNDA.n387 9.3005
R593 GNDA.n386 GNDA.n354 9.3005
R594 GNDA.n385 GNDA.n384 9.3005
R595 GNDA.n383 GNDA.n355 9.3005
R596 GNDA.n382 GNDA.n381 9.3005
R597 GNDA.n380 GNDA.n356 9.3005
R598 GNDA.n379 GNDA.n378 9.3005
R599 GNDA.n377 GNDA.n359 9.3005
R600 GNDA.n375 GNDA.n374 9.3005
R601 GNDA.n373 GNDA.n360 9.3005
R602 GNDA.n372 GNDA.n371 9.3005
R603 GNDA.n370 GNDA.n361 9.3005
R604 GNDA.n369 GNDA.n368 9.3005
R605 GNDA.n367 GNDA.n362 9.3005
R606 GNDA.n366 GNDA.n365 9.3005
R607 GNDA.n22 GNDA.n21 9.3005
R608 GNDA.n407 GNDA.n406 9.3005
R609 GNDA.n408 GNDA.n20 9.3005
R610 GNDA.n410 GNDA.n409 9.3005
R611 GNDA.n411 GNDA.n18 9.3005
R612 GNDA.n414 GNDA.n413 9.3005
R613 GNDA.n415 GNDA.n17 9.3005
R614 GNDA.n417 GNDA.n416 9.3005
R615 GNDA.n419 GNDA.n15 9.3005
R616 GNDA.n421 GNDA.n420 9.3005
R617 GNDA.n422 GNDA.n14 9.3005
R618 GNDA.n424 GNDA.n423 9.3005
R619 GNDA.n426 GNDA.n12 9.3005
R620 GNDA.n428 GNDA.n427 9.3005
R621 GNDA.n429 GNDA.n11 9.3005
R622 GNDA.n431 GNDA.n430 9.3005
R623 GNDA.n432 GNDA.n10 9.3005
R624 GNDA.n434 GNDA.n433 9.3005
R625 GNDA.n435 GNDA.n9 9.3005
R626 GNDA.n437 GNDA.n436 9.3005
R627 GNDA.n439 GNDA.n6 9.3005
R628 GNDA.n442 GNDA.n441 9.3005
R629 GNDA.n443 GNDA.n5 9.3005
R630 GNDA.n445 GNDA.n444 9.3005
R631 GNDA.n446 GNDA.n4 9.3005
R632 GNDA.n448 GNDA.n447 9.3005
R633 GNDA.n449 GNDA.n3 9.3005
R634 GNDA.n451 GNDA.n450 9.3005
R635 GNDA.n452 GNDA.n1 9.3005
R636 GNDA.t138 GNDA.t149 8.62795
R637 GNDA.t103 GNDA.t121 8.62795
R638 GNDA.n296 GNDA.n190 7.49888
R639 GNDA.n146 GNDA.n145 7.11161
R640 GNDA.n143 GNDA.n141 7.11161
R641 GNDA.n74 GNDA.n72 7.11161
R642 GNDA.n79 GNDA.n69 7.11161
R643 GNDA.n139 GNDA.n138 6.69883
R644 GNDA.n131 GNDA.n130 6.4005
R645 GNDA.n109 GNDA.n108 6.4005
R646 GNDA.n104 GNDA.n103 6.4005
R647 GNDA.n283 GNDA.n202 6.4005
R648 GNDA.n264 GNDA.n211 6.4005
R649 GNDA.n259 GNDA.n212 6.4005
R650 GNDA.n218 GNDA.n216 6.4005
R651 GNDA.n246 GNDA.n245 6.4005
R652 GNDA.n234 GNDA.n233 6.4005
R653 GNDA.n170 GNDA.n166 6.4005
R654 GNDA.n368 GNDA.n364 6.4005
R655 GNDA.n406 GNDA.n405 6.4005
R656 GNDA.n419 GNDA.n418 6.4005
R657 GNDA.n426 GNDA.n425 6.4005
R658 GNDA.n438 GNDA.n437 6.4005
R659 GNDA.n453 GNDA.n452 6.4005
R660 GNDA.n83 GNDA.n81 6.4005
R661 GNDA.n230 GNDA.n229 5.68939
R662 GNDA.n230 GNDA.n219 5.68939
R663 GNDA.n398 GNDA.n8 5.68939
R664 GNDA.n398 GNDA.n7 4.97828
R665 GNDA.n145 GNDA.n144 3.48951
R666 GNDA.n144 GNDA.n143 3.48951
R667 GNDA.n74 GNDA.n73 3.48951
R668 GNDA.n73 GNDA.n69 3.48951
R669 GNDA.n289 GNDA.n192 3.2005
R670 GNDA.n277 GNDA.n276 3.2005
R671 GNDA.t133 GNDA.t54 2.88386
R672 GNDA.t88 GNDA.t38 2.87632
R673 GNDA.n97 GNDA.n61 2.25882
R674 GNDA.n61 GNDA.n60 2.25882
R675 GNDA.n102 GNDA.n54 2.25882
R676 GNDA.n60 GNDA.n59 2.25882
R677 GNDA.n98 GNDA.n97 2.25882
R678 GNDA.n59 GNDA.n54 2.25882
R679 GNDA.n118 GNDA.n44 2.25882
R680 GNDA.n44 GNDA.n43 2.25882
R681 GNDA.n123 GNDA.n37 2.25882
R682 GNDA.n43 GNDA.n42 2.25882
R683 GNDA.n119 GNDA.n118 2.25882
R684 GNDA.n42 GNDA.n37 2.25882
R685 GNDA.n297 GNDA.n27 0.9875
R686 GNDA.n139 GNDA.n31 0.703977
R687 GNDA.n296 GNDA.n295 0.193977
R688 GNDA.n235 GNDA.n0 0.193881
R689 GNDA.n454 GNDA.n1 0.193881
R690 GNDA.n390 GNDA.n352 0.193695
R691 GNDA.n299 GNDA.n298 0.188
R692 GNDA.n295 GNDA.n191 0.15675
R693 GNDA.n291 GNDA.n191 0.15675
R694 GNDA.n291 GNDA.n290 0.15675
R695 GNDA.n290 GNDA.n193 0.15675
R696 GNDA.n286 GNDA.n193 0.15675
R697 GNDA.n286 GNDA.n285 0.15675
R698 GNDA.n285 GNDA.n284 0.15675
R699 GNDA.n284 GNDA.n195 0.15675
R700 GNDA.n280 GNDA.n195 0.15675
R701 GNDA.n280 GNDA.n279 0.15675
R702 GNDA.n279 GNDA.n278 0.15675
R703 GNDA.n278 GNDA.n204 0.15675
R704 GNDA.n273 GNDA.n204 0.15675
R705 GNDA.n273 GNDA.n272 0.15675
R706 GNDA.n272 GNDA.n271 0.15675
R707 GNDA.n271 GNDA.n207 0.15675
R708 GNDA.n267 GNDA.n207 0.15675
R709 GNDA.n267 GNDA.n266 0.15675
R710 GNDA.n266 GNDA.n265 0.15675
R711 GNDA.n265 GNDA.n210 0.15675
R712 GNDA.n261 GNDA.n210 0.15675
R713 GNDA.n261 GNDA.n260 0.15675
R714 GNDA.n260 GNDA.n213 0.15675
R715 GNDA.n256 GNDA.n213 0.15675
R716 GNDA.n256 GNDA.n255 0.15675
R717 GNDA.n255 GNDA.n254 0.15675
R718 GNDA.n254 GNDA.n215 0.15675
R719 GNDA.n250 GNDA.n215 0.15675
R720 GNDA.n250 GNDA.n249 0.15675
R721 GNDA.n249 GNDA.n248 0.15675
R722 GNDA.n248 GNDA.n217 0.15675
R723 GNDA.n243 GNDA.n217 0.15675
R724 GNDA.n243 GNDA.n242 0.15675
R725 GNDA.n242 GNDA.n241 0.15675
R726 GNDA.n241 GNDA.n221 0.15675
R727 GNDA.n237 GNDA.n221 0.15675
R728 GNDA.n237 GNDA.n236 0.15675
R729 GNDA.n236 GNDA.n235 0.15675
R730 GNDA.n334 GNDA.n153 0.15675
R731 GNDA.n330 GNDA.n329 0.15675
R732 GNDA.n329 GNDA.n328 0.15675
R733 GNDA.n328 GNDA.n157 0.15675
R734 GNDA.n324 GNDA.n323 0.15675
R735 GNDA.n323 GNDA.n322 0.15675
R736 GNDA.n322 GNDA.n161 0.15675
R737 GNDA.n318 GNDA.n317 0.15675
R738 GNDA.n317 GNDA.n316 0.15675
R739 GNDA.n316 GNDA.n165 0.15675
R740 GNDA.n312 GNDA.n311 0.15675
R741 GNDA.n311 GNDA.n310 0.15675
R742 GNDA.n310 GNDA.n169 0.15675
R743 GNDA.n306 GNDA.n305 0.15675
R744 GNDA.n303 GNDA.n189 0.15675
R745 GNDA.n299 GNDA.n189 0.15675
R746 GNDA.n134 GNDA.n31 0.15675
R747 GNDA.n134 GNDA.n133 0.15675
R748 GNDA.n133 GNDA.n132 0.15675
R749 GNDA.n132 GNDA.n33 0.15675
R750 GNDA.n127 GNDA.n33 0.15675
R751 GNDA.n127 GNDA.n126 0.15675
R752 GNDA.n126 GNDA.n125 0.15675
R753 GNDA.n125 GNDA.n35 0.15675
R754 GNDA.n46 GNDA.n35 0.15675
R755 GNDA.n47 GNDA.n46 0.15675
R756 GNDA.n113 GNDA.n47 0.15675
R757 GNDA.n113 GNDA.n112 0.15675
R758 GNDA.n112 GNDA.n111 0.15675
R759 GNDA.n111 GNDA.n49 0.15675
R760 GNDA.n107 GNDA.n49 0.15675
R761 GNDA.n107 GNDA.n106 0.15675
R762 GNDA.n106 GNDA.n105 0.15675
R763 GNDA.n105 GNDA.n52 0.15675
R764 GNDA.n63 GNDA.n52 0.15675
R765 GNDA.n64 GNDA.n63 0.15675
R766 GNDA.n65 GNDA.n64 0.15675
R767 GNDA.n92 GNDA.n65 0.15675
R768 GNDA.n92 GNDA.n91 0.15675
R769 GNDA.n91 GNDA.n90 0.15675
R770 GNDA.n90 GNDA.n67 0.15675
R771 GNDA.n86 GNDA.n67 0.15675
R772 GNDA.n86 GNDA.n85 0.15675
R773 GNDA.n85 GNDA.n84 0.15675
R774 GNDA.n390 GNDA.n389 0.15675
R775 GNDA.n389 GNDA.n388 0.15675
R776 GNDA.n388 GNDA.n354 0.15675
R777 GNDA.n384 GNDA.n354 0.15675
R778 GNDA.n384 GNDA.n383 0.15675
R779 GNDA.n383 GNDA.n382 0.15675
R780 GNDA.n382 GNDA.n356 0.15675
R781 GNDA.n378 GNDA.n356 0.15675
R782 GNDA.n378 GNDA.n377 0.15675
R783 GNDA.n375 GNDA.n360 0.15675
R784 GNDA.n371 GNDA.n360 0.15675
R785 GNDA.n371 GNDA.n370 0.15675
R786 GNDA.n370 GNDA.n369 0.15675
R787 GNDA.n369 GNDA.n362 0.15675
R788 GNDA.n365 GNDA.n362 0.15675
R789 GNDA.n365 GNDA.n21 0.15675
R790 GNDA.n407 GNDA.n21 0.15675
R791 GNDA.n408 GNDA.n407 0.15675
R792 GNDA.n409 GNDA.n408 0.15675
R793 GNDA.n409 GNDA.n18 0.15675
R794 GNDA.n414 GNDA.n18 0.15675
R795 GNDA.n415 GNDA.n414 0.15675
R796 GNDA.n416 GNDA.n415 0.15675
R797 GNDA.n416 GNDA.n15 0.15675
R798 GNDA.n421 GNDA.n15 0.15675
R799 GNDA.n422 GNDA.n421 0.15675
R800 GNDA.n423 GNDA.n422 0.15675
R801 GNDA.n423 GNDA.n12 0.15675
R802 GNDA.n428 GNDA.n12 0.15675
R803 GNDA.n429 GNDA.n428 0.15675
R804 GNDA.n430 GNDA.n429 0.15675
R805 GNDA.n430 GNDA.n10 0.15675
R806 GNDA.n434 GNDA.n10 0.15675
R807 GNDA.n435 GNDA.n434 0.15675
R808 GNDA.n436 GNDA.n435 0.15675
R809 GNDA.n436 GNDA.n6 0.15675
R810 GNDA.n442 GNDA.n6 0.15675
R811 GNDA.n443 GNDA.n442 0.15675
R812 GNDA.n444 GNDA.n443 0.15675
R813 GNDA.n444 GNDA.n4 0.15675
R814 GNDA.n448 GNDA.n4 0.15675
R815 GNDA.n449 GNDA.n448 0.15675
R816 GNDA.n450 GNDA.n449 0.15675
R817 GNDA.n450 GNDA.n1 0.15675
R818 GNDA.n351 GNDA.n27 0.1321
R819 GNDA.n335 GNDA.n150 0.131895
R820 GNDA.n84 GNDA 0.1255
R821 GNDA.n377 GNDA.n376 0.109875
R822 GNDA.n156 GNDA.n153 0.09425
R823 GNDA.n160 GNDA.n157 0.09425
R824 GNDA.n164 GNDA.n161 0.09425
R825 GNDA.n168 GNDA.n165 0.09425
R826 GNDA.n173 GNDA.n169 0.09425
R827 GNDA.n305 GNDA.n304 0.09425
R828 GNDA.n335 GNDA.n334 0.063
R829 GNDA.n330 GNDA.n156 0.063
R830 GNDA.n324 GNDA.n160 0.063
R831 GNDA.n318 GNDA.n164 0.063
R832 GNDA.n312 GNDA.n168 0.063
R833 GNDA.n306 GNDA.n173 0.063
R834 GNDA.n304 GNDA.n303 0.063
R835 GNDA.n82 GNDA 0.063
R836 GNDA.n376 GNDA.n375 0.047375
R837 V_OUT.n1 V_OUT.t8 377.567
R838 V_OUT.n0 V_OUT.t10 297.233
R839 V_OUT.n5 V_OUT.n4 242.903
R840 V_OUT.n2 V_OUT.n0 237.851
R841 V_OUT.n2 V_OUT.n1 232.809
R842 V_OUT.n1 V_OUT.t9 216.9
R843 V_OUT.n5 V_OUT.n3 172.502
R844 V_OUT.n9 V_OUT.t4 164.118
R845 V_OUT.n0 V_OUT.t11 136.567
R846 V_OUT.n10 V_OUT.n7 118.35
R847 V_OUT.n7 V_OUT.n6 106.662
R848 V_OUT.n10 V_OUT 50.938
R849 V_OUT.n3 V_OUT.t6 24.6255
R850 V_OUT.n3 V_OUT.t5 24.6255
R851 V_OUT.n4 V_OUT.t3 24.6255
R852 V_OUT.n4 V_OUT.t2 24.6255
R853 V_OUT.n7 V_OUT.n5 22.4005
R854 V_OUT.n6 V_OUT.t1 15.0005
R855 V_OUT.n6 V_OUT.t0 15.0005
R856 V_OUT.n10 V_OUT.n9 9.91717
R857 V_OUT.n9 V_OUT.t7 8.246
R858 V_OUT V_OUT.n2 1.39633
R859 V_OUT.n10 V_OUT.n8 0.0838333
R860 V_OUT V_OUT.n10 0.063
R861 a_5970_4630.n8 a_5970_4630.n6 522.322
R862 a_5970_4630.n3 a_5970_4630.t7 384.967
R863 a_5970_4630.n0 a_5970_4630.t10 384.967
R864 a_5970_4630.n3 a_5970_4630.t9 379.166
R865 a_5970_4630.t11 a_5970_4630.n0 376.56
R866 a_5970_4630.n5 a_5970_4630.n1 315.647
R867 a_5970_4630.n4 a_5970_4630.n2 315.647
R868 a_5970_4630.n11 a_5970_4630.n10 314.502
R869 a_5970_4630.n8 a_5970_4630.n7 160.721
R870 a_5970_4630.n5 a_5970_4630.n4 83.2005
R871 a_5970_4630.n1 a_5970_4630.t3 49.2505
R872 a_5970_4630.n1 a_5970_4630.t6 49.2505
R873 a_5970_4630.n2 a_5970_4630.t5 49.2505
R874 a_5970_4630.n2 a_5970_4630.t8 49.2505
R875 a_5970_4630.t11 a_5970_4630.n11 49.2505
R876 a_5970_4630.n11 a_5970_4630.t12 49.2505
R877 a_5970_4630.n10 a_5970_4630.n9 42.6672
R878 a_5970_4630.n9 a_5970_4630.n8 37.763
R879 a_5970_4630.n9 a_5970_4630.n5 23.4672
R880 a_5970_4630.n6 a_5970_4630.t2 19.7005
R881 a_5970_4630.n6 a_5970_4630.t1 19.7005
R882 a_5970_4630.n7 a_5970_4630.t0 19.7005
R883 a_5970_4630.n7 a_5970_4630.t4 19.7005
R884 a_5970_4630.n4 a_5970_4630.n3 16.0005
R885 a_5970_4630.n10 a_5970_4630.n0 16.0005
R886 VDDA.n468 VDDA.n460 831.25
R887 VDDA.n463 VDDA.n462 831.25
R888 VDDA.n457 VDDA.n449 831.25
R889 VDDA.n452 VDDA.n451 831.25
R890 VDDA.n461 VDDA.n460 585
R891 VDDA.n465 VDDA.n463 585
R892 VDDA.n361 VDDA.n355 585
R893 VDDA.n356 VDDA.n355 585
R894 VDDA.n367 VDDA.n44 585
R895 VDDA.n371 VDDA.n44 585
R896 VDDA.n312 VDDA.n50 585
R897 VDDA.n307 VDDA.n50 585
R898 VDDA.n288 VDDA.n283 585
R899 VDDA.n292 VDDA.n283 585
R900 VDDA.n450 VDDA.n449 585
R901 VDDA.n454 VDDA.n452 585
R902 VDDA.n352 VDDA.n346 585
R903 VDDA.n347 VDDA.n346 585
R904 VDDA.n58 VDDA.n51 585
R905 VDDA.n53 VDDA.n51 585
R906 VDDA.n123 VDDA.n116 585
R907 VDDA.n105 VDDA.n97 585
R908 VDDA.n271 VDDA.n175 585
R909 VDDA.n264 VDDA.n175 585
R910 VDDA.n261 VDDA.n260 585
R911 VDDA.n260 VDDA.n259 585
R912 VDDA.n230 VDDA.n229 585
R913 VDDA.n230 VDDA.n219 585
R914 VDDA.n467 VDDA.t126 465.079
R915 VDDA.t126 VDDA.n466 465.079
R916 VDDA.n456 VDDA.t21 465.079
R917 VDDA.t21 VDDA.n455 465.079
R918 VDDA.t77 VDDA.n336 464.281
R919 VDDA.n338 VDDA.t77 464.281
R920 VDDA.n444 VDDA.t129 464.281
R921 VDDA.t129 VDDA.n443 464.281
R922 VDDA.n481 VDDA.t33 464.281
R923 VDDA.t33 VDDA.n480 464.281
R924 VDDA.n425 VDDA.t54 464.281
R925 VDDA.t54 VDDA.n424 464.281
R926 VDDA.n403 VDDA.t75 464.281
R927 VDDA.t75 VDDA.n402 464.281
R928 VDDA.n333 VDDA.t39 464.281
R929 VDDA.t39 VDDA.n332 464.281
R930 VDDA.t67 VDDA.n433 464.281
R931 VDDA.n434 VDDA.t67 464.281
R932 VDDA.t78 VDDA.n17 464.281
R933 VDDA.n471 VDDA.t78 464.281
R934 VDDA.t48 VDDA.n25 464.281
R935 VDDA.n406 VDDA.t48 464.281
R936 VDDA.t42 VDDA.n321 464.281
R937 VDDA.n322 VDDA.t42 464.281
R938 VDDA.n41 VDDA.t130 415.336
R939 VDDA.n86 VDDA.t106 384.967
R940 VDDA.n128 VDDA.t112 384.967
R941 VDDA.n91 VDDA.t91 384.967
R942 VDDA.n111 VDDA.t88 384.967
R943 VDDA.n123 VDDA.t99 374.878
R944 VDDA.t110 VDDA.t72 360.346
R945 VDDA.t72 VDDA.t68 360.346
R946 VDDA.t68 VDDA.t56 360.346
R947 VDDA.t56 VDDA.t51 360.346
R948 VDDA.t51 VDDA.t103 360.346
R949 VDDA.t10 VDDA.t117 360.346
R950 VDDA.t34 VDDA.t10 360.346
R951 VDDA.t26 VDDA.t34 360.346
R952 VDDA.t4 VDDA.t26 360.346
R953 VDDA.t120 VDDA.t4 360.346
R954 VDDA.n96 VDDA.t95 352.834
R955 VDDA.n225 VDDA.t110 343.966
R956 VDDA.n263 VDDA.t103 343.966
R957 VDDA.t117 VDDA.n263 343.966
R958 VDDA.n269 VDDA.t120 343.966
R959 VDDA.n112 VDDA.t90 341.752
R960 VDDA.n127 VDDA.t115 341.752
R961 VDDA.n87 VDDA.t108 341.752
R962 VDDA.n92 VDDA.t94 341.752
R963 VDDA.n258 VDDA.t116 336.329
R964 VDDA.n258 VDDA.t102 336.329
R965 VDDA.n220 VDDA.t109 320.7
R966 VDDA.n272 VDDA.t119 320.7
R967 VDDA.n85 VDDA.n83 315.647
R968 VDDA.n79 VDDA.n78 315.647
R969 VDDA.n110 VDDA.n109 315.647
R970 VDDA.n90 VDDA.n89 315.647
R971 VDDA.n130 VDDA.n82 315.647
R972 VDDA.n129 VDDA.n84 315.647
R973 VDDA.n24 VDDA.t25 315.25
R974 VDDA.t8 VDDA.t9 314.113
R975 VDDA.t28 VDDA.t80 314.113
R976 VDDA.t107 VDDA.n87 304.659
R977 VDDA.n260 VDDA.n183 291.363
R978 VDDA.n256 VDDA.n181 291.363
R979 VDDA.n257 VDDA.n256 291.363
R980 VDDA.n359 VDDA.n355 290.733
R981 VDDA.n365 VDDA.n44 290.733
R982 VDDA.n310 VDDA.n50 290.733
R983 VDDA.n286 VDDA.n283 290.733
R984 VDDA.n350 VDDA.n346 290.733
R985 VDDA.n52 VDDA.n51 290.733
R986 VDDA.n121 VDDA.n116 290.733
R987 VDDA.n117 VDDA.n116 290.733
R988 VDDA.n103 VDDA.n97 290.733
R989 VDDA.n98 VDDA.n97 290.733
R990 VDDA.n265 VDDA.n175 290.733
R991 VDDA.n230 VDDA.n218 290.733
R992 VDDA.n445 VDDA.n444 243.698
R993 VDDA.n482 VDDA.n481 243.698
R994 VDDA.n426 VDDA.n425 243.698
R995 VDDA.n404 VDDA.n403 243.698
R996 VDDA.n334 VDDA.n333 243.698
R997 VDDA.n434 VDDA.n431 243.698
R998 VDDA.n475 VDDA.n471 243.698
R999 VDDA.n410 VDDA.n406 243.698
R1000 VDDA.n322 VDDA.n319 243.698
R1001 VDDA.n430 VDDA.n1 238.367
R1002 VDDA.n469 VDDA.n468 238.367
R1003 VDDA.n462 VDDA.n429 238.367
R1004 VDDA.n428 VDDA.n16 238.367
R1005 VDDA.n421 VDDA.n19 238.367
R1006 VDDA.n399 VDDA.n27 238.367
R1007 VDDA.n318 VDDA.n35 238.367
R1008 VDDA.n438 VDDA.n2 238.367
R1009 VDDA.n458 VDDA.n457 238.367
R1010 VDDA.n485 VDDA.n484 238.367
R1011 VDDA.n413 VDDA.n412 238.367
R1012 VDDA.n326 VDDA.n31 238.367
R1013 VDDA.n451 VDDA.n447 238.367
R1014 VDDA.n117 VDDA.n88 233.841
R1015 VDDA.n98 VDDA.n94 233.841
R1016 VDDA.n362 VDDA.n361 230.308
R1017 VDDA.n356 VDDA.n315 230.308
R1018 VDDA.n368 VDDA.n367 230.308
R1019 VDDA.n371 VDDA.n370 230.308
R1020 VDDA.n313 VDDA.n312 230.308
R1021 VDDA.n307 VDDA.n46 230.308
R1022 VDDA.n289 VDDA.n288 230.308
R1023 VDDA.n292 VDDA.n291 230.308
R1024 VDDA.n353 VDDA.n352 230.308
R1025 VDDA.n58 VDDA.n48 230.308
R1026 VDDA.n53 VDDA.n47 230.308
R1027 VDDA.n347 VDDA.n344 230.308
R1028 VDDA.n124 VDDA.n123 230.308
R1029 VDDA.n271 VDDA.n270 230.308
R1030 VDDA.n268 VDDA.n264 230.308
R1031 VDDA.n262 VDDA.n261 230.308
R1032 VDDA.n259 VDDA.n178 230.308
R1033 VDDA.t40 VDDA.t30 222.178
R1034 VDDA.n363 VDDA.n343 199.195
R1035 VDDA.n192 VDDA.n191 196.502
R1036 VDDA.n189 VDDA.n188 196.502
R1037 VDDA.n255 VDDA.n254 196.502
R1038 VDDA.n246 VDDA.n211 196.502
R1039 VDDA.n239 VDDA.n214 196.502
R1040 VDDA.n232 VDDA.n231 196.502
R1041 VDDA.n338 VDDA.n317 190.333
R1042 VDDA.n127 VDDA.n126 185.001
R1043 VDDA.n113 VDDA.n112 185.001
R1044 VDDA.n108 VDDA.n92 185.001
R1045 VDDA.n57 VDDA.n56 185
R1046 VDDA.n55 VDDA.n54 185
R1047 VDDA.n351 VDDA.n345 185
R1048 VDDA.n349 VDDA.n348 185
R1049 VDDA.n325 VDDA.n324 185
R1050 VDDA.n323 VDDA.n320 185
R1051 VDDA.n407 VDDA.n26 185
R1052 VDDA.n409 VDDA.n408 185
R1053 VDDA.n472 VDDA.n18 185
R1054 VDDA.n474 VDDA.n473 185
R1055 VDDA.n450 VDDA.n448 185
R1056 VDDA.n454 VDDA.n453 185
R1057 VDDA.n437 VDDA.n436 185
R1058 VDDA.n435 VDDA.n432 185
R1059 VDDA.n287 VDDA.n285 185
R1060 VDDA.n284 VDDA.n282 185
R1061 VDDA.n311 VDDA.n49 185
R1062 VDDA.n309 VDDA.n308 185
R1063 VDDA.n366 VDDA.n364 185
R1064 VDDA.n45 VDDA.n43 185
R1065 VDDA.n360 VDDA.n354 185
R1066 VDDA.n358 VDDA.n357 185
R1067 VDDA.n329 VDDA.n328 185
R1068 VDDA.n331 VDDA.n330 185
R1069 VDDA.n29 VDDA.n28 185
R1070 VDDA.n401 VDDA.n400 185
R1071 VDDA.n21 VDDA.n20 185
R1072 VDDA.n423 VDDA.n422 185
R1073 VDDA.n477 VDDA.n476 185
R1074 VDDA.n479 VDDA.n478 185
R1075 VDDA.n461 VDDA.n459 185
R1076 VDDA.n465 VDDA.n464 185
R1077 VDDA.n440 VDDA.n439 185
R1078 VDDA.n442 VDDA.n441 185
R1079 VDDA.n342 VDDA.n34 185
R1080 VDDA.n343 VDDA.n342 185
R1081 VDDA.n341 VDDA.n340 185
R1082 VDDA.n339 VDDA.n337 185
R1083 VDDA.n343 VDDA.n317 185
R1084 VDDA.n122 VDDA.n115 185
R1085 VDDA.n120 VDDA.n114 185
R1086 VDDA.n125 VDDA.n114 185
R1087 VDDA.n119 VDDA.n118 185
R1088 VDDA.n106 VDDA.n105 185
R1089 VDDA.n107 VDDA.n106 185
R1090 VDDA.n104 VDDA.n95 185
R1091 VDDA.n102 VDDA.n101 185
R1092 VDDA.n100 VDDA.n99 185
R1093 VDDA.n182 VDDA.n179 185
R1094 VDDA.n185 VDDA.n184 185
R1095 VDDA.n177 VDDA.n176 185
R1096 VDDA.n267 VDDA.n266 185
R1097 VDDA.n229 VDDA.n221 185
R1098 VDDA.n225 VDDA.n221 185
R1099 VDDA.n228 VDDA.n227 185
R1100 VDDA.n223 VDDA.n222 185
R1101 VDDA.n224 VDDA.n219 185
R1102 VDDA.n225 VDDA.n224 185
R1103 VDDA.n290 VDDA.t40 172.38
R1104 VDDA.t83 VDDA.n314 172.38
R1105 VDDA.n369 VDDA.t2 172.38
R1106 VDDA.n259 VDDA.n258 166.63
R1107 VDDA.n441 VDDA.n439 150
R1108 VDDA.n464 VDDA.n459 150
R1109 VDDA.n478 VDDA.n476 150
R1110 VDDA.n422 VDDA.n20 150
R1111 VDDA.n400 VDDA.n28 150
R1112 VDDA.n330 VDDA.n328 150
R1113 VDDA.n437 VDDA.n432 150
R1114 VDDA.n453 VDDA.n448 150
R1115 VDDA.n474 VDDA.n18 150
R1116 VDDA.n409 VDDA.n26 150
R1117 VDDA.n325 VDDA.n320 150
R1118 VDDA.n342 VDDA.n341 150
R1119 VDDA.n337 VDDA.n317 150
R1120 VDDA.t22 VDDA.t18 145.038
R1121 VDDA.n335 VDDA.n327 137.904
R1122 VDDA.n411 VDDA.n405 137.904
R1123 VDDA.n290 VDDA.t123 126.412
R1124 VDDA.n314 VDDA.t30 126.412
R1125 VDDA.n369 VDDA.t83 126.412
R1126 VDDA.t2 VDDA.n363 126.412
R1127 VDDA.t125 VDDA.n460 123.126
R1128 VDDA.n463 VDDA.t125 123.126
R1129 VDDA.t7 VDDA.n449 123.126
R1130 VDDA.n452 VDDA.t7 123.126
R1131 VDDA.n357 VDDA.n354 120.001
R1132 VDDA.n364 VDDA.n45 120.001
R1133 VDDA.n308 VDDA.n49 120.001
R1134 VDDA.n285 VDDA.n284 120.001
R1135 VDDA.n348 VDDA.n345 120.001
R1136 VDDA.n56 VDDA.n55 120.001
R1137 VDDA.n115 VDDA.n114 120.001
R1138 VDDA.n118 VDDA.n114 120.001
R1139 VDDA.n106 VDDA.n95 120.001
R1140 VDDA.n101 VDDA.n100 120.001
R1141 VDDA.n267 VDDA.n177 120.001
R1142 VDDA.n184 VDDA.n179 120.001
R1143 VDDA.n227 VDDA.n221 120.001
R1144 VDDA.n224 VDDA.n223 120.001
R1145 VDDA.n161 VDDA.n67 119.737
R1146 VDDA.n154 VDDA.n70 119.737
R1147 VDDA.n147 VDDA.n73 119.737
R1148 VDDA.n140 VDDA.n76 119.737
R1149 VDDA.n132 VDDA.n81 119.737
R1150 VDDA.n126 VDDA.t113 119.656
R1151 VDDA.n125 VDDA.n113 108.779
R1152 VDDA.n483 VDDA.n427 107.258
R1153 VDDA.n483 VDDA.t32 103.427
R1154 VDDA.t20 VDDA.n470 103.427
R1155 VDDA.n470 VDDA.t6 103.427
R1156 VDDA.t66 VDDA.n446 103.427
R1157 VDDA.n427 VDDA.t47 95.7666
R1158 VDDA.t62 VDDA.t107 94.2753
R1159 VDDA.t60 VDDA.t62 94.2753
R1160 VDDA.t58 VDDA.t60 94.2753
R1161 VDDA.t64 VDDA.t58 94.2753
R1162 VDDA.t113 VDDA.t64 94.2753
R1163 VDDA.t49 VDDA.t70 94.2753
R1164 VDDA.t0 VDDA.t92 94.2753
R1165 VDDA.t36 VDDA.n108 94.2753
R1166 VDDA.t87 VDDA.t127 94.2753
R1167 VDDA.t85 VDDA.t84 94.2753
R1168 VDDA.t38 VDDA.t76 91.936
R1169 VDDA.t74 VDDA.t41 91.936
R1170 VDDA.t24 VDDA.t53 84.2747
R1171 VDDA.t32 VDDA.t8 84.2747
R1172 VDDA.t9 VDDA.t20 84.2747
R1173 VDDA.t6 VDDA.t28 84.2747
R1174 VDDA.t80 VDDA.t66 84.2747
R1175 VDDA.t100 VDDA.t89 83.3974
R1176 VDDA.t12 VDDA.t29 83.3974
R1177 VDDA.n110 VDDA.n79 83.2005
R1178 VDDA.n90 VDDA.n79 83.2005
R1179 VDDA.n130 VDDA.n83 83.2005
R1180 VDDA.n130 VDDA.n129 83.2005
R1181 VDDA.t14 VDDA.t81 76.1455
R1182 VDDA.t96 VDDA.t86 76.1455
R1183 VDDA.n314 VDDA.n48 69.8479
R1184 VDDA.n314 VDDA.n47 69.8479
R1185 VDDA.n363 VDDA.n353 69.8479
R1186 VDDA.n363 VDDA.n344 69.8479
R1187 VDDA.n290 VDDA.n289 69.8479
R1188 VDDA.n291 VDDA.n290 69.8479
R1189 VDDA.n314 VDDA.n313 69.8479
R1190 VDDA.n314 VDDA.n46 69.8479
R1191 VDDA.n369 VDDA.n368 69.8479
R1192 VDDA.n370 VDDA.n369 69.8479
R1193 VDDA.n363 VDDA.n362 69.8479
R1194 VDDA.n363 VDDA.n315 69.8479
R1195 VDDA.n125 VDDA.n124 69.8479
R1196 VDDA.n125 VDDA.n88 69.8479
R1197 VDDA.n107 VDDA.n93 69.8479
R1198 VDDA.n107 VDDA.n94 69.8479
R1199 VDDA.n263 VDDA.n262 69.8479
R1200 VDDA.n263 VDDA.n178 69.8479
R1201 VDDA.n270 VDDA.n269 69.8479
R1202 VDDA.n269 VDDA.n268 69.8479
R1203 VDDA.n226 VDDA.n225 69.8479
R1204 VDDA.n131 VDDA.n130 69.3203
R1205 VDDA.t81 VDDA.t45 68.8936
R1206 VDDA.t86 VDDA.n107 68.8936
R1207 VDDA.n327 VDDA.n326 65.8183
R1208 VDDA.n327 VDDA.n319 65.8183
R1209 VDDA.n412 VDDA.n411 65.8183
R1210 VDDA.n411 VDDA.n410 65.8183
R1211 VDDA.n484 VDDA.n483 65.8183
R1212 VDDA.n483 VDDA.n475 65.8183
R1213 VDDA.n470 VDDA.n458 65.8183
R1214 VDDA.n470 VDDA.n447 65.8183
R1215 VDDA.n446 VDDA.n438 65.8183
R1216 VDDA.n446 VDDA.n431 65.8183
R1217 VDDA.n335 VDDA.n334 65.8183
R1218 VDDA.n335 VDDA.n318 65.8183
R1219 VDDA.n405 VDDA.n404 65.8183
R1220 VDDA.n405 VDDA.n27 65.8183
R1221 VDDA.n427 VDDA.n426 65.8183
R1222 VDDA.n427 VDDA.n19 65.8183
R1223 VDDA.n483 VDDA.n482 65.8183
R1224 VDDA.n483 VDDA.n428 65.8183
R1225 VDDA.n470 VDDA.n469 65.8183
R1226 VDDA.n470 VDDA.n429 65.8183
R1227 VDDA.n446 VDDA.n445 65.8183
R1228 VDDA.n446 VDDA.n430 65.8183
R1229 VDDA.n343 VDDA.n316 65.8183
R1230 VDDA.t89 VDDA.t16 61.6417
R1231 VDDA.t29 VDDA.t43 61.6417
R1232 VDDA.n516 VDDA.n1 58.0576
R1233 VDDA.n486 VDDA.n16 58.0576
R1234 VDDA.n421 VDDA.n420 58.0576
R1235 VDDA.n399 VDDA.n398 58.0576
R1236 VDDA.n389 VDDA.n35 58.0576
R1237 VDDA.n516 VDDA.n2 58.0576
R1238 VDDA.n486 VDDA.n485 58.0576
R1239 VDDA.n414 VDDA.n413 58.0576
R1240 VDDA.n397 VDDA.n31 58.0576
R1241 VDDA.n390 VDDA.n34 58.0576
R1242 VDDA.n356 VDDA.n38 57.2449
R1243 VDDA.n372 VDDA.n371 57.2449
R1244 VDDA.n307 VDDA.n306 57.2449
R1245 VDDA.n293 VDDA.n292 57.2449
R1246 VDDA.n352 VDDA.n38 57.2449
R1247 VDDA.n306 VDDA.n58 57.2449
R1248 VDDA.n503 VDDA.n7 54.4005
R1249 VDDA.n9 VDDA.n7 54.4005
R1250 VDDA.n9 VDDA.n8 54.4005
R1251 VDDA.n503 VDDA.n8 54.4005
R1252 VDDA.n432 VDDA.n431 53.3664
R1253 VDDA.n453 VDDA.n447 53.3664
R1254 VDDA.n475 VDDA.n474 53.3664
R1255 VDDA.n326 VDDA.n325 53.3664
R1256 VDDA.n320 VDDA.n319 53.3664
R1257 VDDA.n412 VDDA.n26 53.3664
R1258 VDDA.n410 VDDA.n409 53.3664
R1259 VDDA.n484 VDDA.n18 53.3664
R1260 VDDA.n458 VDDA.n448 53.3664
R1261 VDDA.n438 VDDA.n437 53.3664
R1262 VDDA.n334 VDDA.n328 53.3664
R1263 VDDA.n330 VDDA.n318 53.3664
R1264 VDDA.n404 VDDA.n28 53.3664
R1265 VDDA.n400 VDDA.n27 53.3664
R1266 VDDA.n426 VDDA.n20 53.3664
R1267 VDDA.n422 VDDA.n19 53.3664
R1268 VDDA.n482 VDDA.n476 53.3664
R1269 VDDA.n478 VDDA.n428 53.3664
R1270 VDDA.n469 VDDA.n459 53.3664
R1271 VDDA.n464 VDDA.n429 53.3664
R1272 VDDA.n445 VDDA.n439 53.3664
R1273 VDDA.n441 VDDA.n430 53.3664
R1274 VDDA.n341 VDDA.n316 53.3664
R1275 VDDA.n337 VDDA.n316 53.3664
R1276 VDDA.n108 VDDA.t22 50.7639
R1277 VDDA.t108 VDDA.n85 49.2505
R1278 VDDA.n85 VDDA.t63 49.2505
R1279 VDDA.n78 VDDA.t71 49.2505
R1280 VDDA.n78 VDDA.t82 49.2505
R1281 VDDA.n109 VDDA.t90 49.2505
R1282 VDDA.n109 VDDA.t50 49.2505
R1283 VDDA.n89 VDDA.t1 49.2505
R1284 VDDA.n89 VDDA.t93 49.2505
R1285 VDDA.n82 VDDA.t61 49.2505
R1286 VDDA.n82 VDDA.t59 49.2505
R1287 VDDA.n84 VDDA.t65 49.2505
R1288 VDDA.n84 VDDA.t114 49.2505
R1289 VDDA VDDA.n517 47.763
R1290 VDDA.n348 VDDA.n344 45.3071
R1291 VDDA.n55 VDDA.n47 45.3071
R1292 VDDA.n56 VDDA.n48 45.3071
R1293 VDDA.n353 VDDA.n345 45.3071
R1294 VDDA.n289 VDDA.n285 45.3071
R1295 VDDA.n291 VDDA.n284 45.3071
R1296 VDDA.n313 VDDA.n49 45.3071
R1297 VDDA.n308 VDDA.n46 45.3071
R1298 VDDA.n368 VDDA.n364 45.3071
R1299 VDDA.n370 VDDA.n45 45.3071
R1300 VDDA.n362 VDDA.n354 45.3071
R1301 VDDA.n357 VDDA.n315 45.3071
R1302 VDDA.n118 VDDA.n88 45.3071
R1303 VDDA.n124 VDDA.n115 45.3071
R1304 VDDA.n95 VDDA.n93 45.3071
R1305 VDDA.n100 VDDA.n94 45.3071
R1306 VDDA.n101 VDDA.n93 45.3071
R1307 VDDA.n262 VDDA.n179 45.3071
R1308 VDDA.n184 VDDA.n178 45.3071
R1309 VDDA.n270 VDDA.n177 45.3071
R1310 VDDA.n268 VDDA.n267 45.3071
R1311 VDDA.n227 VDDA.n226 45.3071
R1312 VDDA.n226 VDDA.n223 45.3071
R1313 VDDA.n137 VDDA.n79 41.6005
R1314 VDDA.t18 VDDA.t87 39.886
R1315 VDDA.n131 VDDA.n80 39.4988
R1316 VDDA.n279 VDDA.n278 38.1005
R1317 VDDA.n113 VDDA.t100 36.26
R1318 VDDA.t16 VDDA.t49 32.6341
R1319 VDDA.t43 VDDA.t85 32.6341
R1320 VDDA.n261 VDDA.n180 32.2291
R1321 VDDA.n294 VDDA.n62 32.0005
R1322 VDDA.n298 VDDA.n62 32.0005
R1323 VDDA.n299 VDDA.n298 32.0005
R1324 VDDA.n300 VDDA.n299 32.0005
R1325 VDDA.n300 VDDA.n59 32.0005
R1326 VDDA.n306 VDDA.n59 32.0005
R1327 VDDA.n306 VDDA.n60 32.0005
R1328 VDDA.n60 VDDA.n42 32.0005
R1329 VDDA.n373 VDDA.n42 32.0005
R1330 VDDA.n377 VDDA.n40 32.0005
R1331 VDDA.n378 VDDA.n377 32.0005
R1332 VDDA.n379 VDDA.n378 32.0005
R1333 VDDA.n383 VDDA.n382 32.0005
R1334 VDDA.n384 VDDA.n383 32.0005
R1335 VDDA.n384 VDDA.n36 32.0005
R1336 VDDA.n388 VDDA.n36 32.0005
R1337 VDDA.n392 VDDA.n391 32.0005
R1338 VDDA.n392 VDDA.n30 32.0005
R1339 VDDA.n396 VDDA.n32 32.0005
R1340 VDDA.n419 VDDA.n22 32.0005
R1341 VDDA.n487 VDDA.n15 32.0005
R1342 VDDA.n491 VDDA.n13 32.0005
R1343 VDDA.n492 VDDA.n491 32.0005
R1344 VDDA.n493 VDDA.n492 32.0005
R1345 VDDA.n493 VDDA.n11 32.0005
R1346 VDDA.n497 VDDA.n11 32.0005
R1347 VDDA.n498 VDDA.n497 32.0005
R1348 VDDA.n499 VDDA.n498 32.0005
R1349 VDDA.n505 VDDA.n504 32.0005
R1350 VDDA.n505 VDDA.n5 32.0005
R1351 VDDA.n509 VDDA.n5 32.0005
R1352 VDDA.n510 VDDA.n509 32.0005
R1353 VDDA.n511 VDDA.n510 32.0005
R1354 VDDA.n511 VDDA.n3 32.0005
R1355 VDDA.n515 VDDA.n3 32.0005
R1356 VDDA.n135 VDDA.n80 32.0005
R1357 VDDA.n136 VDDA.n135 32.0005
R1358 VDDA.n138 VDDA.n75 32.0005
R1359 VDDA.n143 VDDA.n75 32.0005
R1360 VDDA.n144 VDDA.n143 32.0005
R1361 VDDA.n145 VDDA.n144 32.0005
R1362 VDDA.n145 VDDA.n72 32.0005
R1363 VDDA.n150 VDDA.n72 32.0005
R1364 VDDA.n151 VDDA.n150 32.0005
R1365 VDDA.n152 VDDA.n151 32.0005
R1366 VDDA.n152 VDDA.n69 32.0005
R1367 VDDA.n157 VDDA.n69 32.0005
R1368 VDDA.n158 VDDA.n157 32.0005
R1369 VDDA.n159 VDDA.n158 32.0005
R1370 VDDA.n159 VDDA.n66 32.0005
R1371 VDDA.n164 VDDA.n66 32.0005
R1372 VDDA.n165 VDDA.n164 32.0005
R1373 VDDA.n165 VDDA.n64 32.0005
R1374 VDDA.n169 VDDA.n64 32.0005
R1375 VDDA.n170 VDDA.n169 32.0005
R1376 VDDA.n274 VDDA.n172 32.0005
R1377 VDDA.n278 VDDA.n172 32.0005
R1378 VDDA.n198 VDDA.n197 32.0005
R1379 VDDA.n197 VDDA.n196 32.0005
R1380 VDDA.n204 VDDA.n186 32.0005
R1381 VDDA.n204 VDDA.n203 32.0005
R1382 VDDA.n203 VDDA.n202 32.0005
R1383 VDDA.n253 VDDA.n208 32.0005
R1384 VDDA.n248 VDDA.n247 32.0005
R1385 VDDA.n241 VDDA.n240 32.0005
R1386 VDDA.n241 VDDA.n212 32.0005
R1387 VDDA.n245 VDDA.n212 32.0005
R1388 VDDA.n234 VDDA.n233 32.0005
R1389 VDDA.n234 VDDA.n215 32.0005
R1390 VDDA.n238 VDDA.n215 32.0005
R1391 VDDA.n128 VDDA.n127 30.754
R1392 VDDA.n92 VDDA.n91 30.754
R1393 VDDA.n112 VDDA.n111 30.186
R1394 VDDA.n87 VDDA.n86 30.186
R1395 VDDA.n373 VDDA.n372 28.8005
R1396 VDDA.n273 VDDA.n174 28.8005
R1397 VDDA.n198 VDDA.n189 28.8005
R1398 VDDA.n254 VDDA.n253 28.8005
R1399 VDDA.n294 VDDA.n293 25.6005
R1400 VDDA.n379 VDDA.n38 25.6005
R1401 VDDA.n391 VDDA.n390 25.6005
R1402 VDDA.n415 VDDA.n414 25.6005
R1403 VDDA.n420 VDDA.n15 25.6005
R1404 VDDA.n487 VDDA.n486 25.6005
R1405 VDDA.n502 VDDA.n9 25.6005
R1406 VDDA.n503 VDDA.n502 25.6005
R1407 VDDA.n517 VDDA.n516 25.6005
R1408 VDDA.n137 VDDA.n136 25.6005
R1409 VDDA VDDA.n170 25.6005
R1410 VDDA.t45 VDDA.t0 25.3822
R1411 VDDA.t92 VDDA.t36 25.3822
R1412 VDDA.n355 VDDA.t3 24.6255
R1413 VDDA.n44 VDDA.t128 24.6255
R1414 VDDA.n50 VDDA.t31 24.6255
R1415 VDDA.n283 VDDA.t124 24.6255
R1416 VDDA.n346 VDDA.t79 24.6255
R1417 VDDA.n51 VDDA.t55 24.6255
R1418 VDDA.n191 VDDA.t5 24.6255
R1419 VDDA.n191 VDDA.t121 24.6255
R1420 VDDA.n188 VDDA.t35 24.6255
R1421 VDDA.n188 VDDA.t27 24.6255
R1422 VDDA.t118 VDDA.n255 24.6255
R1423 VDDA.n255 VDDA.t11 24.6255
R1424 VDDA.n211 VDDA.t52 24.6255
R1425 VDDA.n211 VDDA.t104 24.6255
R1426 VDDA.n214 VDDA.t69 24.6255
R1427 VDDA.n214 VDDA.t57 24.6255
R1428 VDDA.n231 VDDA.t111 24.6255
R1429 VDDA.n231 VDDA.t73 24.6255
R1430 VDDA.t111 VDDA.n230 24.6255
R1431 VDDA.n175 VDDA.t122 24.6255
R1432 VDDA.n256 VDDA.t118 24.6255
R1433 VDDA.n260 VDDA.t105 24.6255
R1434 VDDA.n220 VDDA.n217 24.361
R1435 VDDA.n196 VDDA.n192 22.4005
R1436 VDDA.n247 VDDA.n246 22.4005
R1437 VDDA.n248 VDDA.n180 22.4005
R1438 VDDA.n105 VDDA.n96 22.0449
R1439 VDDA.n116 VDDA.t101 19.7005
R1440 VDDA.n97 VDDA.t98 19.7005
R1441 VDDA.n67 VDDA.t44 19.7005
R1442 VDDA.n67 VDDA.t97 19.7005
R1443 VDDA.n70 VDDA.t19 19.7005
R1444 VDDA.n70 VDDA.t13 19.7005
R1445 VDDA.n73 VDDA.t37 19.7005
R1446 VDDA.n73 VDDA.t23 19.7005
R1447 VDDA.n76 VDDA.t15 19.7005
R1448 VDDA.n76 VDDA.t46 19.7005
R1449 VDDA.t101 VDDA.n81 19.7005
R1450 VDDA.n81 VDDA.t17 19.7005
R1451 VDDA.n32 VDDA.n24 19.2005
R1452 VDDA.t70 VDDA.t14 18.1303
R1453 VDDA.t84 VDDA.t96 18.1303
R1454 VDDA.n273 VDDA.n272 17.6005
R1455 VDDA.n397 VDDA.n396 16.0005
R1456 VDDA.n129 VDDA.n128 16.0005
R1457 VDDA.n91 VDDA.n90 16.0005
R1458 VDDA.n111 VDDA.n110 16.0005
R1459 VDDA.n86 VDDA.n83 16.0005
R1460 VDDA.n192 VDDA.n174 16.0005
R1461 VDDA.n208 VDDA.n180 16.0005
R1462 VDDA.n246 VDDA.n245 16.0005
R1463 VDDA.n233 VDDA.n232 16.0005
R1464 VDDA.n171 VDDA 15.7005
R1465 VDDA.n272 VDDA.n271 15.6449
R1466 VDDA.n229 VDDA.n220 15.6449
R1467 VDDA.n293 VDDA.n281 13.8989
R1468 VDDA.n398 VDDA.n30 12.8005
R1469 VDDA.n415 VDDA.n24 12.8005
R1470 VDDA.n280 VDDA.n171 12.7493
R1471 VDDA.n281 VDDA.n280 12.3383
R1472 VDDA.n280 VDDA.n279 11.579
R1473 VDDA.n343 VDDA.t38 11.4924
R1474 VDDA.t76 VDDA.n335 11.4924
R1475 VDDA.n327 VDDA.t74 11.4924
R1476 VDDA.n405 VDDA.t41 11.4924
R1477 VDDA.n411 VDDA.t24 11.4924
R1478 VDDA.t127 VDDA.t12 10.8784
R1479 VDDA.n96 VDDA.n65 9.613
R1480 VDDA.n274 VDDA.n273 9.6005
R1481 VDDA.n254 VDDA.n186 9.6005
R1482 VDDA.n202 VDDA.n189 9.6005
R1483 VDDA.n170 VDDA.n63 9.3005
R1484 VDDA.n169 VDDA.n168 9.3005
R1485 VDDA.n167 VDDA.n64 9.3005
R1486 VDDA.n166 VDDA.n165 9.3005
R1487 VDDA.n164 VDDA.n163 9.3005
R1488 VDDA.n162 VDDA.n66 9.3005
R1489 VDDA.n160 VDDA.n159 9.3005
R1490 VDDA.n158 VDDA.n68 9.3005
R1491 VDDA.n157 VDDA.n156 9.3005
R1492 VDDA.n155 VDDA.n69 9.3005
R1493 VDDA.n153 VDDA.n152 9.3005
R1494 VDDA.n151 VDDA.n71 9.3005
R1495 VDDA.n150 VDDA.n149 9.3005
R1496 VDDA.n148 VDDA.n72 9.3005
R1497 VDDA.n146 VDDA.n145 9.3005
R1498 VDDA.n144 VDDA.n74 9.3005
R1499 VDDA.n143 VDDA.n142 9.3005
R1500 VDDA.n141 VDDA.n75 9.3005
R1501 VDDA.n139 VDDA.n138 9.3005
R1502 VDDA.n133 VDDA.n80 9.3005
R1503 VDDA.n135 VDDA.n134 9.3005
R1504 VDDA.n136 VDDA.n77 9.3005
R1505 VDDA.n233 VDDA.n216 9.3005
R1506 VDDA.n235 VDDA.n234 9.3005
R1507 VDDA.n236 VDDA.n215 9.3005
R1508 VDDA.n238 VDDA.n237 9.3005
R1509 VDDA.n240 VDDA.n213 9.3005
R1510 VDDA.n242 VDDA.n241 9.3005
R1511 VDDA.n243 VDDA.n212 9.3005
R1512 VDDA.n245 VDDA.n244 9.3005
R1513 VDDA.n246 VDDA.n210 9.3005
R1514 VDDA.n247 VDDA.n209 9.3005
R1515 VDDA.n249 VDDA.n248 9.3005
R1516 VDDA.n250 VDDA.n180 9.3005
R1517 VDDA.n251 VDDA.n208 9.3005
R1518 VDDA.n253 VDDA.n252 9.3005
R1519 VDDA.n254 VDDA.n207 9.3005
R1520 VDDA.n206 VDDA.n186 9.3005
R1521 VDDA.n205 VDDA.n204 9.3005
R1522 VDDA.n203 VDDA.n187 9.3005
R1523 VDDA.n202 VDDA.n201 9.3005
R1524 VDDA.n200 VDDA.n189 9.3005
R1525 VDDA.n199 VDDA.n198 9.3005
R1526 VDDA.n197 VDDA.n190 9.3005
R1527 VDDA.n196 VDDA.n195 9.3005
R1528 VDDA.n194 VDDA.n192 9.3005
R1529 VDDA.n193 VDDA.n174 9.3005
R1530 VDDA.n273 VDDA.n173 9.3005
R1531 VDDA.n275 VDDA.n274 9.3005
R1532 VDDA.n276 VDDA.n172 9.3005
R1533 VDDA.n278 VDDA.n277 9.3005
R1534 VDDA.n517 VDDA.n0 9.3005
R1535 VDDA.n295 VDDA.n294 9.3005
R1536 VDDA.n296 VDDA.n62 9.3005
R1537 VDDA.n298 VDDA.n297 9.3005
R1538 VDDA.n299 VDDA.n61 9.3005
R1539 VDDA.n301 VDDA.n300 9.3005
R1540 VDDA.n302 VDDA.n59 9.3005
R1541 VDDA.n306 VDDA.n305 9.3005
R1542 VDDA.n304 VDDA.n60 9.3005
R1543 VDDA.n303 VDDA.n42 9.3005
R1544 VDDA.n374 VDDA.n373 9.3005
R1545 VDDA.n375 VDDA.n40 9.3005
R1546 VDDA.n377 VDDA.n376 9.3005
R1547 VDDA.n378 VDDA.n39 9.3005
R1548 VDDA.n380 VDDA.n379 9.3005
R1549 VDDA.n382 VDDA.n381 9.3005
R1550 VDDA.n383 VDDA.n37 9.3005
R1551 VDDA.n385 VDDA.n384 9.3005
R1552 VDDA.n386 VDDA.n36 9.3005
R1553 VDDA.n388 VDDA.n387 9.3005
R1554 VDDA.n391 VDDA.n33 9.3005
R1555 VDDA.n393 VDDA.n392 9.3005
R1556 VDDA.n394 VDDA.n30 9.3005
R1557 VDDA.n396 VDDA.n395 9.3005
R1558 VDDA.n32 VDDA.n23 9.3005
R1559 VDDA.n416 VDDA.n415 9.3005
R1560 VDDA.n417 VDDA.n22 9.3005
R1561 VDDA.n419 VDDA.n418 9.3005
R1562 VDDA.n15 VDDA.n14 9.3005
R1563 VDDA.n488 VDDA.n487 9.3005
R1564 VDDA.n489 VDDA.n13 9.3005
R1565 VDDA.n491 VDDA.n490 9.3005
R1566 VDDA.n492 VDDA.n12 9.3005
R1567 VDDA.n494 VDDA.n493 9.3005
R1568 VDDA.n495 VDDA.n11 9.3005
R1569 VDDA.n497 VDDA.n496 9.3005
R1570 VDDA.n498 VDDA.n10 9.3005
R1571 VDDA.n500 VDDA.n499 9.3005
R1572 VDDA.n502 VDDA.n501 9.3005
R1573 VDDA.n504 VDDA.n6 9.3005
R1574 VDDA.n506 VDDA.n505 9.3005
R1575 VDDA.n507 VDDA.n5 9.3005
R1576 VDDA.n509 VDDA.n508 9.3005
R1577 VDDA.n510 VDDA.n4 9.3005
R1578 VDDA.n512 VDDA.n511 9.3005
R1579 VDDA.n513 VDDA.n3 9.3005
R1580 VDDA.n515 VDDA.n514 9.3005
R1581 VDDA.n442 VDDA.n440 9.14336
R1582 VDDA.n479 VDDA.n477 9.14336
R1583 VDDA.n423 VDDA.n21 9.14336
R1584 VDDA.n401 VDDA.n29 9.14336
R1585 VDDA.n331 VDDA.n329 9.14336
R1586 VDDA.n436 VDDA.n435 9.14336
R1587 VDDA.n473 VDDA.n472 9.14336
R1588 VDDA.n408 VDDA.n407 9.14336
R1589 VDDA.n324 VDDA.n323 9.14336
R1590 VDDA.n340 VDDA.n339 9.14336
R1591 VDDA.t53 VDDA.t47 7.66179
R1592 VDDA.n126 VDDA.n125 7.25241
R1593 VDDA.n361 VDDA.n360 7.11161
R1594 VDDA.n358 VDDA.n356 7.11161
R1595 VDDA.n367 VDDA.n366 7.11161
R1596 VDDA.n371 VDDA.n43 7.11161
R1597 VDDA.n312 VDDA.n311 7.11161
R1598 VDDA.n309 VDDA.n307 7.11161
R1599 VDDA.n288 VDDA.n287 7.11161
R1600 VDDA.n292 VDDA.n282 7.11161
R1601 VDDA.n352 VDDA.n351 7.11161
R1602 VDDA.n349 VDDA.n347 7.11161
R1603 VDDA.n58 VDDA.n57 7.11161
R1604 VDDA.n54 VDDA.n53 7.11161
R1605 VDDA.n123 VDDA.n122 7.11161
R1606 VDDA.n120 VDDA.n119 7.11161
R1607 VDDA.n105 VDDA.n104 7.11161
R1608 VDDA.n102 VDDA.n99 7.11161
R1609 VDDA.n271 VDDA.n176 7.11161
R1610 VDDA.n266 VDDA.n264 7.11161
R1611 VDDA.n229 VDDA.n228 7.11161
R1612 VDDA.n222 VDDA.n219 7.11161
R1613 VDDA.n232 VDDA.n217 6.54033
R1614 VDDA.n382 VDDA.n38 6.4005
R1615 VDDA.n414 VDDA.n22 6.4005
R1616 VDDA.n420 VDDA.n419 6.4005
R1617 VDDA.n486 VDDA.n13 6.4005
R1618 VDDA.n499 VDDA.n9 6.4005
R1619 VDDA.n504 VDDA.n503 6.4005
R1620 VDDA.n516 VDDA.n515 6.4005
R1621 VDDA.n138 VDDA.n137 6.4005
R1622 VDDA.n465 VDDA.n461 5.81868
R1623 VDDA.n454 VDDA.n450 5.81868
R1624 VDDA.n336 VDDA.n34 5.33286
R1625 VDDA.n443 VDDA.n1 5.33286
R1626 VDDA.n480 VDDA.n16 5.33286
R1627 VDDA.n424 VDDA.n421 5.33286
R1628 VDDA.n402 VDDA.n399 5.33286
R1629 VDDA.n332 VDDA.n35 5.33286
R1630 VDDA.n433 VDDA.n2 5.33286
R1631 VDDA.n485 VDDA.n17 5.33286
R1632 VDDA.n413 VDDA.n25 5.33286
R1633 VDDA.n321 VDDA.n31 5.33286
R1634 VDDA.n444 VDDA.n440 3.75335
R1635 VDDA.n443 VDDA.n442 3.75335
R1636 VDDA.n481 VDDA.n477 3.75335
R1637 VDDA.n480 VDDA.n479 3.75335
R1638 VDDA.n425 VDDA.n21 3.75335
R1639 VDDA.n424 VDDA.n423 3.75335
R1640 VDDA.n403 VDDA.n29 3.75335
R1641 VDDA.n402 VDDA.n401 3.75335
R1642 VDDA.n333 VDDA.n329 3.75335
R1643 VDDA.n332 VDDA.n331 3.75335
R1644 VDDA.n436 VDDA.n433 3.75335
R1645 VDDA.n435 VDDA.n434 3.75335
R1646 VDDA.n472 VDDA.n17 3.75335
R1647 VDDA.n473 VDDA.n471 3.75335
R1648 VDDA.n407 VDDA.n25 3.75335
R1649 VDDA.n408 VDDA.n406 3.75335
R1650 VDDA.n324 VDDA.n321 3.75335
R1651 VDDA.n323 VDDA.n322 3.75335
R1652 VDDA.n340 VDDA.n336 3.75335
R1653 VDDA.n339 VDDA.n338 3.75335
R1654 VDDA.n360 VDDA.n359 3.53508
R1655 VDDA.n359 VDDA.n358 3.53508
R1656 VDDA.n366 VDDA.n365 3.53508
R1657 VDDA.n365 VDDA.n43 3.53508
R1658 VDDA.n311 VDDA.n310 3.53508
R1659 VDDA.n310 VDDA.n309 3.53508
R1660 VDDA.n287 VDDA.n286 3.53508
R1661 VDDA.n286 VDDA.n282 3.53508
R1662 VDDA.n351 VDDA.n350 3.53508
R1663 VDDA.n350 VDDA.n349 3.53508
R1664 VDDA.n57 VDDA.n52 3.53508
R1665 VDDA.n54 VDDA.n52 3.53508
R1666 VDDA.n122 VDDA.n121 3.53508
R1667 VDDA.n119 VDDA.n117 3.53508
R1668 VDDA.n121 VDDA.n120 3.53508
R1669 VDDA.n104 VDDA.n103 3.53508
R1670 VDDA.n99 VDDA.n98 3.53508
R1671 VDDA.n103 VDDA.n102 3.53508
R1672 VDDA.n265 VDDA.n176 3.53508
R1673 VDDA.n266 VDDA.n265 3.53508
R1674 VDDA.n228 VDDA.n218 3.53508
R1675 VDDA.n222 VDDA.n218 3.53508
R1676 VDDA.n468 VDDA.n467 3.40194
R1677 VDDA.n466 VDDA.n462 3.40194
R1678 VDDA.n457 VDDA.n456 3.40194
R1679 VDDA.n455 VDDA.n451 3.40194
R1680 VDDA.n372 VDDA.n40 3.2005
R1681 VDDA.n389 VDDA.n388 3.2005
R1682 VDDA.n390 VDDA.n389 3.2005
R1683 VDDA.n398 VDDA.n397 3.2005
R1684 VDDA.n240 VDDA.n239 3.2005
R1685 VDDA.n239 VDDA.n238 3.2005
R1686 VDDA.n467 VDDA.n461 2.39444
R1687 VDDA.n466 VDDA.n465 2.39444
R1688 VDDA.n456 VDDA.n450 2.39444
R1689 VDDA.n455 VDDA.n454 2.39444
R1690 VDDA.n462 VDDA.n7 2.32777
R1691 VDDA.n457 VDDA.n8 2.32777
R1692 VDDA.n182 VDDA.n181 2.27782
R1693 VDDA.n183 VDDA.n182 2.27782
R1694 VDDA.n259 VDDA.n257 2.27782
R1695 VDDA.n185 VDDA.n183 2.27782
R1696 VDDA.n261 VDDA.n181 2.27782
R1697 VDDA.n257 VDDA.n185 2.27782
R1698 VDDA.n217 VDDA.n216 0.703395
R1699 VDDA.n295 VDDA.n281 0.193961
R1700 VDDA.n171 VDDA.n63 0.188
R1701 VDDA.n134 VDDA.n133 0.15675
R1702 VDDA.n134 VDDA.n77 0.15675
R1703 VDDA.n139 VDDA.n77 0.15675
R1704 VDDA.n142 VDDA.n141 0.15675
R1705 VDDA.n142 VDDA.n74 0.15675
R1706 VDDA.n146 VDDA.n74 0.15675
R1707 VDDA.n149 VDDA.n148 0.15675
R1708 VDDA.n149 VDDA.n71 0.15675
R1709 VDDA.n153 VDDA.n71 0.15675
R1710 VDDA.n156 VDDA.n155 0.15675
R1711 VDDA.n156 VDDA.n68 0.15675
R1712 VDDA.n160 VDDA.n68 0.15675
R1713 VDDA.n163 VDDA.n162 0.15675
R1714 VDDA.n167 VDDA.n166 0.15675
R1715 VDDA.n168 VDDA.n167 0.15675
R1716 VDDA.n168 VDDA.n63 0.15675
R1717 VDDA.n235 VDDA.n216 0.15675
R1718 VDDA.n236 VDDA.n235 0.15675
R1719 VDDA.n237 VDDA.n236 0.15675
R1720 VDDA.n237 VDDA.n213 0.15675
R1721 VDDA.n242 VDDA.n213 0.15675
R1722 VDDA.n243 VDDA.n242 0.15675
R1723 VDDA.n244 VDDA.n243 0.15675
R1724 VDDA.n244 VDDA.n210 0.15675
R1725 VDDA.n210 VDDA.n209 0.15675
R1726 VDDA.n249 VDDA.n209 0.15675
R1727 VDDA.n250 VDDA.n249 0.15675
R1728 VDDA.n251 VDDA.n250 0.15675
R1729 VDDA.n252 VDDA.n251 0.15675
R1730 VDDA.n252 VDDA.n207 0.15675
R1731 VDDA.n207 VDDA.n206 0.15675
R1732 VDDA.n206 VDDA.n205 0.15675
R1733 VDDA.n205 VDDA.n187 0.15675
R1734 VDDA.n201 VDDA.n187 0.15675
R1735 VDDA.n201 VDDA.n200 0.15675
R1736 VDDA.n200 VDDA.n199 0.15675
R1737 VDDA.n199 VDDA.n190 0.15675
R1738 VDDA.n195 VDDA.n190 0.15675
R1739 VDDA.n195 VDDA.n194 0.15675
R1740 VDDA.n194 VDDA.n193 0.15675
R1741 VDDA.n193 VDDA.n173 0.15675
R1742 VDDA.n275 VDDA.n173 0.15675
R1743 VDDA.n276 VDDA.n275 0.15675
R1744 VDDA.n277 VDDA.n276 0.15675
R1745 VDDA.n296 VDDA.n295 0.15675
R1746 VDDA.n297 VDDA.n296 0.15675
R1747 VDDA.n297 VDDA.n61 0.15675
R1748 VDDA.n301 VDDA.n61 0.15675
R1749 VDDA.n302 VDDA.n301 0.15675
R1750 VDDA.n305 VDDA.n302 0.15675
R1751 VDDA.n305 VDDA.n304 0.15675
R1752 VDDA.n304 VDDA.n303 0.15675
R1753 VDDA.n375 VDDA.n374 0.15675
R1754 VDDA.n376 VDDA.n375 0.15675
R1755 VDDA.n376 VDDA.n39 0.15675
R1756 VDDA.n380 VDDA.n39 0.15675
R1757 VDDA.n381 VDDA.n380 0.15675
R1758 VDDA.n381 VDDA.n37 0.15675
R1759 VDDA.n385 VDDA.n37 0.15675
R1760 VDDA.n386 VDDA.n385 0.15675
R1761 VDDA.n387 VDDA.n386 0.15675
R1762 VDDA.n387 VDDA.n33 0.15675
R1763 VDDA.n393 VDDA.n33 0.15675
R1764 VDDA.n394 VDDA.n393 0.15675
R1765 VDDA.n395 VDDA.n394 0.15675
R1766 VDDA.n395 VDDA.n23 0.15675
R1767 VDDA.n416 VDDA.n23 0.15675
R1768 VDDA.n417 VDDA.n416 0.15675
R1769 VDDA.n418 VDDA.n417 0.15675
R1770 VDDA.n418 VDDA.n14 0.15675
R1771 VDDA.n488 VDDA.n14 0.15675
R1772 VDDA.n489 VDDA.n488 0.15675
R1773 VDDA.n490 VDDA.n489 0.15675
R1774 VDDA.n490 VDDA.n12 0.15675
R1775 VDDA.n494 VDDA.n12 0.15675
R1776 VDDA.n495 VDDA.n494 0.15675
R1777 VDDA.n496 VDDA.n495 0.15675
R1778 VDDA.n496 VDDA.n10 0.15675
R1779 VDDA.n500 VDDA.n10 0.15675
R1780 VDDA.n501 VDDA.n500 0.15675
R1781 VDDA.n501 VDDA.n6 0.15675
R1782 VDDA.n506 VDDA.n6 0.15675
R1783 VDDA.n507 VDDA.n506 0.15675
R1784 VDDA.n508 VDDA.n507 0.15675
R1785 VDDA.n508 VDDA.n4 0.15675
R1786 VDDA.n512 VDDA.n4 0.15675
R1787 VDDA.n513 VDDA.n512 0.15675
R1788 VDDA.n514 VDDA.n513 0.15675
R1789 VDDA.n514 VDDA.n0 0.15675
R1790 VDDA VDDA.n0 0.1255
R1791 VDDA.n277 VDDA 0.122375
R1792 VDDA.n132 VDDA.n131 0.100307
R1793 VDDA.n133 VDDA.n132 0.09425
R1794 VDDA.n141 VDDA.n140 0.09425
R1795 VDDA.n148 VDDA.n147 0.09425
R1796 VDDA.n155 VDDA.n154 0.09425
R1797 VDDA.n162 VDDA.n161 0.09425
R1798 VDDA.n166 VDDA.n65 0.09425
R1799 VDDA.n303 VDDA.n41 0.078625
R1800 VDDA.n374 VDDA.n41 0.078625
R1801 VDDA.n140 VDDA.n139 0.063
R1802 VDDA.n147 VDDA.n146 0.063
R1803 VDDA.n154 VDDA.n153 0.063
R1804 VDDA.n161 VDDA.n160 0.063
R1805 VDDA.n163 VDDA.n65 0.063
R1806 VDDA.n279 VDDA 0.0505
R1807 pfd_8_0.DOWN_PFD_b.t1 pfd_8_0.DOWN_PFD_b.n1 203.528
R1808 pfd_8_0.DOWN_PFD_b.n0 pfd_8_0.DOWN_PFD_b.t2 203.528
R1809 pfd_8_0.DOWN_PFD_b.n1 pfd_8_0.DOWN_PFD_b.t0 183.935
R1810 pfd_8_0.DOWN_PFD_b.n0 pfd_8_0.DOWN_PFD_b.t3 183.935
R1811 pfd_8_0.DOWN_PFD_b.n1 pfd_8_0.DOWN_PFD_b.n0 83.2005
R1812 pfd_8_0.DOWN_b.n0 pfd_8_0.DOWN_b.t5 1028.27
R1813 pfd_8_0.DOWN_b.n2 pfd_8_0.DOWN_b.n1 569.734
R1814 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.n0 465.933
R1815 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.t3 401.668
R1816 pfd_8_0.DOWN_b.n0 pfd_8_0.DOWN_b.t4 385.601
R1817 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.t2 385.601
R1818 pfd_8_0.DOWN_b.t0 pfd_8_0.DOWN_b.n2 211.847
R1819 pfd_8_0.DOWN_b.n2 pfd_8_0.DOWN_b.t1 173.055
R1820 pfd_8_0.QA_b.t4 pfd_8_0.QA_b.t6 1188.93
R1821 pfd_8_0.QA_b pfd_8_0.QA_b.n2 837.38
R1822 pfd_8_0.QA_b.t6 pfd_8_0.QA_b.t3 835.467
R1823 pfd_8_0.QA_b.n0 pfd_8_0.QA_b.t5 562.333
R1824 pfd_8_0.QA_b pfd_8_0.QA_b.n0 482
R1825 pfd_8_0.QA_b.n2 pfd_8_0.QA_b.n1 247.917
R1826 pfd_8_0.QA_b.n0 pfd_8_0.QA_b.t4 224.934
R1827 pfd_8_0.QA_b.n2 pfd_8_0.QA_b.t1 221.411
R1828 pfd_8_0.QA_b.n1 pfd_8_0.QA_b.t2 24.0005
R1829 pfd_8_0.QA_b.n1 pfd_8_0.QA_b.t0 24.0005
R1830 a_870_1400.t0 a_870_1400.t1 39.4005
R1831 pfd_8_0.UP_input.n1 pfd_8_0.UP_input.t3 326.658
R1832 pfd_8_0.UP_input.n3 pfd_8_0.UP_input.t6 297.233
R1833 pfd_8_0.UP_input.t5 pfd_8_0.UP_input.n4 297.233
R1834 pfd_8_0.UP_input.n2 pfd_8_0.UP_input.n0 257.067
R1835 pfd_8_0.UP_input.n6 pfd_8_0.UP_input.n5 246.275
R1836 pfd_8_0.UP_input.t1 pfd_8_0.UP_input.n7 241.928
R1837 pfd_8_0.UP_input.n5 pfd_8_0.UP_input.n0 226.942
R1838 pfd_8_0.UP_input.n2 pfd_8_0.UP_input.n1 226.942
R1839 pfd_8_0.UP_input.n4 pfd_8_0.UP_input.n3 216.9
R1840 pfd_8_0.UP_input.n6 pfd_8_0.UP_input.t2 209.928
R1841 pfd_8_0.UP_input.n7 pfd_8_0.UP_input.t0 145.536
R1842 pfd_8_0.UP_input.n7 pfd_8_0.UP_input.n6 144
R1843 pfd_8_0.UP_input.n1 pfd_8_0.UP_input.t6 92.3838
R1844 pfd_8_0.UP_input.n5 pfd_8_0.UP_input.t5 92.3838
R1845 pfd_8_0.UP_input.n3 pfd_8_0.UP_input.t7 80.3338
R1846 pfd_8_0.UP_input.t7 pfd_8_0.UP_input.n2 80.3338
R1847 pfd_8_0.UP_input.n4 pfd_8_0.UP_input.t4 80.3338
R1848 pfd_8_0.UP_input.t4 pfd_8_0.UP_input.n0 80.3338
R1849 charge_pump_cell_6_0.UP_b pfd_8_0.UP_b.n1 507.072
R1850 pfd_8_0.UP_b.n1 pfd_8_0.UP_b.n0 409.067
R1851 pfd_8_0.UP_b.n1 pfd_8_0.UP_b.t3 369.534
R1852 pfd_8_0.UP_b.n0 pfd_8_0.UP_b.t0 209.928
R1853 pfd_8_0.UP_b.n0 pfd_8_0.UP_b.t2 177.536
R1854 charge_pump_cell_6_0.UP_b pfd_8_0.UP_b.t1 24.0223
R1855 pfd_8_0.DOWN.t3 pfd_8_0.DOWN.n0 605.311
R1856 charge_pump_cell_6_0.DOWN pfd_8_0.DOWN.t3 399.497
R1857 pfd_8_0.DOWN.n0 pfd_8_0.DOWN.t2 240.327
R1858 pfd_8_0.DOWN.n0 pfd_8_0.DOWN.t1 148.736
R1859 charge_pump_cell_6_0.DOWN pfd_8_0.DOWN.t0 24.487
R1860 pfd_8_0.opamp_out.n6 pfd_8_0.opamp_out.n5 424.447
R1861 pfd_8_0.opamp_out.n6 pfd_8_0.opamp_out.n4 354.048
R1862 pfd_8_0.opamp_out.n2 pfd_8_0.opamp_out.n1 313
R1863 pfd_8_0.opamp_out.n9 pfd_8_0.opamp_out.t14 297.233
R1864 pfd_8_0.opamp_out.n10 pfd_8_0.opamp_out.t14 297.233
R1865 pfd_8_0.opamp_out.t13 pfd_8_0.opamp_out.n11 297.233
R1866 pfd_8_0.opamp_out.n13 pfd_8_0.opamp_out.t1 281.596
R1867 pfd_8_0.opamp_out.n2 pfd_8_0.opamp_out.n0 242.601
R1868 pfd_8_0.opamp_out.n3 pfd_8_0.opamp_out.n2 220.8
R1869 pfd_8_0.opamp_out.n7 pfd_8_0.opamp_out.n6 220.8
R1870 pfd_8_0.opamp_out.n11 pfd_8_0.opamp_out.n10 216.9
R1871 pfd_8_0.opamp_out.n9 pfd_8_0.opamp_out.n8 216.9
R1872 pfd_8_0.opamp_out.n14 pfd_8_0.opamp_out.n12 215.107
R1873 pfd_8_0.opamp_out.n12 pfd_8_0.opamp_out.n8 184.768
R1874 pfd_8_0.opamp_out.n13 pfd_8_0.opamp_out.t0 118.666
R1875 pfd_8_0.opamp_out.n10 pfd_8_0.opamp_out.t15 80.3338
R1876 pfd_8_0.opamp_out.t15 pfd_8_0.opamp_out.n9 80.3338
R1877 pfd_8_0.opamp_out.n11 pfd_8_0.opamp_out.t10 80.3338
R1878 pfd_8_0.opamp_out.t10 pfd_8_0.opamp_out.n8 80.3338
R1879 pfd_8_0.opamp_out.n12 pfd_8_0.opamp_out.t13 80.3338
R1880 pfd_8_0.opamp_out.n15 pfd_8_0.opamp_out.n14 78.9255
R1881 pfd_8_0.opamp_out.n3 pfd_8_0.opamp_out.t12 70.0829
R1882 pfd_8_0.opamp_out.n7 pfd_8_0.opamp_out.t11 63.6829
R1883 opamp_cell_4_0.VOUT pfd_8_0.opamp_out.n3 62.4005
R1884 pfd_8_0.opamp_out.n15 pfd_8_0.opamp_out.n7 60.8005
R1885 pfd_8_0.opamp_out.n14 pfd_8_0.opamp_out.n13 60.2361
R1886 pfd_8_0.opamp_out.n0 pfd_8_0.opamp_out.t8 60.0005
R1887 pfd_8_0.opamp_out.n0 pfd_8_0.opamp_out.t7 60.0005
R1888 pfd_8_0.opamp_out.n1 pfd_8_0.opamp_out.t6 60.0005
R1889 pfd_8_0.opamp_out.n1 pfd_8_0.opamp_out.t9 60.0005
R1890 pfd_8_0.opamp_out.n5 pfd_8_0.opamp_out.t2 49.2505
R1891 pfd_8_0.opamp_out.n5 pfd_8_0.opamp_out.t5 49.2505
R1892 pfd_8_0.opamp_out.n4 pfd_8_0.opamp_out.t4 49.2505
R1893 pfd_8_0.opamp_out.n4 pfd_8_0.opamp_out.t3 49.2505
R1894 opamp_cell_4_0.VOUT pfd_8_0.opamp_out.n15 1.6005
R1895 opamp_cell_4_0.VIN+.n1 opamp_cell_4_0.VIN+.t8 377.567
R1896 opamp_cell_4_0.VIN+.n0 opamp_cell_4_0.VIN+.t6 321.334
R1897 opamp_cell_4_0.VIN+.n2 opamp_cell_4_0.VIN+.n1 233.476
R1898 opamp_cell_4_0.VIN+.n1 opamp_cell_4_0.VIN+.t7 216.9
R1899 opamp_cell_4_0.VIN+.n5 opamp_cell_4_0.VIN+.n4 199.462
R1900 opamp_cell_4_0.VIN+.n2 opamp_cell_4_0.VIN+.n0 189.898
R1901 opamp_cell_4_0.VIN+.n5 opamp_cell_4_0.VIN+.n3 172.502
R1902 opamp_cell_4_0.VIN+.n7 opamp_cell_4_0.VIN+.n6 172.5
R1903 opamp_cell_4_0.VIN+.n0 opamp_cell_4_0.VIN+.t9 112.468
R1904 opamp_cell_4_0.VIN+.n7 opamp_cell_4_0.VIN+.n5 70.4005
R1905 opamp_cell_4_0.VIN+ opamp_cell_4_0.VIN+.n7 50.088
R1906 opamp_cell_4_0.VIN+.n3 opamp_cell_4_0.VIN+.t2 24.6255
R1907 opamp_cell_4_0.VIN+.n3 opamp_cell_4_0.VIN+.t1 24.6255
R1908 opamp_cell_4_0.VIN+.n6 opamp_cell_4_0.VIN+.t4 24.6255
R1909 opamp_cell_4_0.VIN+.n6 opamp_cell_4_0.VIN+.t3 24.6255
R1910 opamp_cell_4_0.VIN+.n4 opamp_cell_4_0.VIN+.t5 15.0005
R1911 opamp_cell_4_0.VIN+.n4 opamp_cell_4_0.VIN+.t0 15.0005
R1912 opamp_cell_4_0.VIN+ opamp_cell_4_0.VIN+.n2 3.313
R1913 a_6320_5840.n7 a_6320_5840.n5 482.582
R1914 a_6320_5840.n10 a_6320_5840.t2 304.634
R1915 a_6320_5840.n3 a_6320_5840.t0 304.634
R1916 a_6320_5840.t4 a_6320_5840.n10 277.914
R1917 a_6320_5840.n3 a_6320_5840.t1 276.289
R1918 a_6320_5840.n8 a_6320_5840.n1 204.201
R1919 a_6320_5840.n4 a_6320_5840.n2 204.201
R1920 a_6320_5840.n9 a_6320_5840.n0 204.201
R1921 a_6320_5840.n7 a_6320_5840.n6 120.981
R1922 a_6320_5840.n8 a_6320_5840.n4 74.6672
R1923 a_6320_5840.n9 a_6320_5840.n8 74.6672
R1924 a_6320_5840.n1 a_6320_5840.t8 60.0005
R1925 a_6320_5840.n1 a_6320_5840.t10 60.0005
R1926 a_6320_5840.t1 a_6320_5840.n2 60.0005
R1927 a_6320_5840.n2 a_6320_5840.t9 60.0005
R1928 a_6320_5840.n0 a_6320_5840.t11 60.0005
R1929 a_6320_5840.n0 a_6320_5840.t3 60.0005
R1930 a_6320_5840.n8 a_6320_5840.n7 37.763
R1931 a_6320_5840.n5 a_6320_5840.t7 24.0005
R1932 a_6320_5840.n5 a_6320_5840.t6 24.0005
R1933 a_6320_5840.n6 a_6320_5840.t5 24.0005
R1934 a_6320_5840.n6 a_6320_5840.t12 24.0005
R1935 a_6320_5840.n4 a_6320_5840.n3 16.0005
R1936 a_6320_5840.n10 a_6320_5840.n9 16.0005
R1937 opamp_cell_4_0.n_right.t4 opamp_cell_4_0.n_right.n6 1010.36
R1938 opamp_cell_4_0.n_right.n3 opamp_cell_4_0.n_right.n2 404.8
R1939 opamp_cell_4_0.n_right.n2 opamp_cell_4_0.n_right.n1 322.048
R1940 opamp_cell_4_0.n_right.n2 opamp_cell_4_0.n_right.n0 316.2
R1941 opamp_cell_4_0.n_right.n4 opamp_cell_4_0.n_right.t8 289.2
R1942 opamp_cell_4_0.n_right.n5 opamp_cell_4_0.n_right.t7 289.2
R1943 opamp_cell_4_0.n_right.n6 opamp_cell_4_0.n_right.t6 289.2
R1944 opamp_cell_4_0.n_right.n3 opamp_cell_4_0.n_right.t5 232.968
R1945 opamp_cell_4_0.n_right.n6 opamp_cell_4_0.n_right.n5 208.868
R1946 opamp_cell_4_0.n_right.n5 opamp_cell_4_0.n_right.n4 208.868
R1947 opamp_cell_4_0.n_right.n4 opamp_cell_4_0.n_right.n3 199.829
R1948 opamp_cell_4_0.n_right.n0 opamp_cell_4_0.n_right.t0 60.0005
R1949 opamp_cell_4_0.n_right.n0 opamp_cell_4_0.n_right.t1 60.0005
R1950 opamp_cell_4_0.n_right.n1 opamp_cell_4_0.n_right.t2 49.2505
R1951 opamp_cell_4_0.n_right.n1 opamp_cell_4_0.n_right.t3 49.2505
R1952 opamp_cell_4_0.n_left.n1 opamp_cell_4_0.n_left.t7 359.894
R1953 opamp_cell_4_0.n_left.n5 opamp_cell_4_0.n_left.n4 325.248
R1954 opamp_cell_4_0.n_left.n4 opamp_cell_4_0.n_left.n0 313
R1955 opamp_cell_4_0.n_left.n3 opamp_cell_4_0.n_left.t0 252.248
R1956 opamp_cell_4_0.n_left.n2 opamp_cell_4_0.n_left.n1 208.868
R1957 opamp_cell_4_0.n_left.n2 opamp_cell_4_0.n_left.t2 192.8
R1958 opamp_cell_4_0.n_left.n1 opamp_cell_4_0.n_left.t6 192.8
R1959 opamp_cell_4_0.n_left.n4 opamp_cell_4_0.n_left.n3 152
R1960 opamp_cell_4_0.n_left.n0 opamp_cell_4_0.n_left.t5 60.0005
R1961 opamp_cell_4_0.n_left.n0 opamp_cell_4_0.n_left.t4 60.0005
R1962 opamp_cell_4_0.n_left.n3 opamp_cell_4_0.n_left.n2 59.4472
R1963 opamp_cell_4_0.n_left.t3 opamp_cell_4_0.n_left.n5 49.2505
R1964 opamp_cell_4_0.n_left.n5 opamp_cell_4_0.n_left.t1 49.2505
R1965 a_6490_4630.t0 a_6490_4630.n6 1112.76
R1966 a_6490_4630.n3 a_6490_4630.n2 441.433
R1967 a_6490_4630.n2 a_6490_4630.n1 379.647
R1968 a_6490_4630.n2 a_6490_4630.n0 258.601
R1969 a_6490_4630.n6 a_6490_4630.t6 208.868
R1970 a_6490_4630.n5 a_6490_4630.t7 208.868
R1971 a_6490_4630.n4 a_6490_4630.t8 208.868
R1972 a_6490_4630.n3 a_6490_4630.t5 208.868
R1973 a_6490_4630.n6 a_6490_4630.n5 208.868
R1974 a_6490_4630.n5 a_6490_4630.n4 208.868
R1975 a_6490_4630.n4 a_6490_4630.n3 208.868
R1976 a_6490_4630.n0 a_6490_4630.t4 60.0005
R1977 a_6490_4630.n0 a_6490_4630.t3 60.0005
R1978 a_6490_4630.n1 a_6490_4630.t2 49.2505
R1979 a_6490_4630.n1 a_6490_4630.t1 49.2505
R1980 pfd_8_0.before_Reset.n1 pfd_8_0.before_Reset.n0 481.334
R1981 pfd_8_0.before_Reset.n0 pfd_8_0.before_Reset.t4 465.933
R1982 pfd_8_0.before_Reset.n0 pfd_8_0.before_Reset.t3 321.334
R1983 pfd_8_0.before_Reset.n2 pfd_8_0.before_Reset.n1 226.889
R1984 pfd_8_0.before_Reset.n1 pfd_8_0.before_Reset.t1 172.458
R1985 pfd_8_0.before_Reset.t0 pfd_8_0.before_Reset.n2 19.7005
R1986 pfd_8_0.before_Reset.n2 pfd_8_0.before_Reset.t2 19.7005
R1987 a_2350_1400.t1 a_2350_1400.n2 500.086
R1988 a_2350_1400.n1 a_2350_1400.n0 473.334
R1989 a_2350_1400.n0 a_2350_1400.t3 465.933
R1990 a_2350_1400.t1 a_2350_1400.n2 461.389
R1991 a_2350_1400.n0 a_2350_1400.t2 321.334
R1992 a_2350_1400.n1 a_2350_1400.t0 177.577
R1993 a_2350_1400.n2 a_2350_1400.n1 48.3899
R1994 opamp_cell_4_0.p_bias opamp_cell_4_0.p_bias.t0 918.318
R1995 opamp_cell_4_0.p_bias opamp_cell_4_0.p_bias.n11 540.801
R1996 opamp_cell_4_0.p_bias.n8 opamp_cell_4_0.p_bias.t10 377.567
R1997 opamp_cell_4_0.p_bias.n3 opamp_cell_4_0.p_bias.t9 377.567
R1998 opamp_cell_4_0.p_bias.n9 opamp_cell_4_0.p_bias.n8 257.067
R1999 opamp_cell_4_0.p_bias.n7 opamp_cell_4_0.p_bias.n6 257.067
R2000 opamp_cell_4_0.p_bias.n4 opamp_cell_4_0.p_bias.n3 257.067
R2001 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n0 154.321
R2002 opamp_cell_4_0.p_bias.n2 opamp_cell_4_0.p_bias.n1 154.321
R2003 opamp_cell_4_0.p_bias.n5 opamp_cell_4_0.p_bias.n2 152
R2004 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n10 152
R2005 opamp_cell_4_0.p_bias.n8 opamp_cell_4_0.p_bias.t12 120.501
R2006 opamp_cell_4_0.p_bias.n9 opamp_cell_4_0.p_bias.t5 120.501
R2007 opamp_cell_4_0.p_bias.n7 opamp_cell_4_0.p_bias.t1 120.501
R2008 opamp_cell_4_0.p_bias.n6 opamp_cell_4_0.p_bias.t3 120.501
R2009 opamp_cell_4_0.p_bias.n3 opamp_cell_4_0.p_bias.t11 120.501
R2010 opamp_cell_4_0.p_bias.n4 opamp_cell_4_0.p_bias.t7 120.501
R2011 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n2 115.201
R2012 opamp_cell_4_0.p_bias.n10 opamp_cell_4_0.p_bias.n9 85.6894
R2013 opamp_cell_4_0.p_bias.n10 opamp_cell_4_0.p_bias.n7 85.6894
R2014 opamp_cell_4_0.p_bias.n6 opamp_cell_4_0.p_bias.n5 85.6894
R2015 opamp_cell_4_0.p_bias.n5 opamp_cell_4_0.p_bias.n4 85.6894
R2016 opamp_cell_4_0.p_bias.n0 opamp_cell_4_0.p_bias.t2 19.7005
R2017 opamp_cell_4_0.p_bias.n0 opamp_cell_4_0.p_bias.t6 19.7005
R2018 opamp_cell_4_0.p_bias.n1 opamp_cell_4_0.p_bias.t8 19.7005
R2019 opamp_cell_4_0.p_bias.n1 opamp_cell_4_0.p_bias.t4 19.7005
R2020 I_IN.n1 I_IN.n0 1269.42
R2021 I_IN.n1 I_IN.t1 275.325
R2022 I_IN.n5 I_IN.n2 248.4
R2023 I_IN.n4 I_IN.t0 238.892
R2024 I_IN.n4 I_IN.t5 161.371
R2025 I_IN.n0 I_IN.t6 151.792
R2026 I_IN I_IN.n4 149.153
R2027 I_IN.n2 I_IN.t3 140.583
R2028 I_IN.n2 I_IN.t1 140.583
R2029 I_IN.n5 I_IN.n3 98.6614
R2030 I_IN.t3 I_IN.n1 80.3338
R2031 I_IN.n0 I_IN.t7 44.2902
R2032 I_IN.n3 I_IN.t4 15.0005
R2033 I_IN.n3 I_IN.t2 15.0005
R2034 I_IN.n5 I_IN 11.488
R2035 I_IN I_IN.n5 3.2005
R2036 F_REF.n0 F_REF.t0 514.134
R2037 F_REF.n0 F_REF.t1 273.134
R2038 F_REF F_REF.n0 216.9
R2039 a_n30_1400.t0 a_n30_1400.t1 39.4005
R2040 pfd_8_0.QA.t5 pfd_8_0.QA.t7 835.467
R2041 pfd_8_0.QA.n2 pfd_8_0.QA.t4 517.347
R2042 pfd_8_0.QA.n0 pfd_8_0.QA.t8 465.933
R2043 pfd_8_0.QA.n1 pfd_8_0.QA.n0 454.031
R2044 pfd_8_0.QA.n1 pfd_8_0.QA.t5 394.267
R2045 pfd_8_0.QA.n0 pfd_8_0.QA.t6 321.334
R2046 pfd_8_0.QA.n4 pfd_8_0.QA.n3 244.715
R2047 pfd_8_0.QA.n2 pfd_8_0.QA.t3 228.148
R2048 pfd_8_0.QA.n4 pfd_8_0.QA.t1 221.411
R2049 pfd_8_0.QA.n5 pfd_8_0.QA.n2 216
R2050 pfd_8_0.QA.n5 pfd_8_0.QA.n4 201.573
R2051 pfd_8_0.QA pfd_8_0.QA.n5 60.8005
R2052 pfd_8_0.QA pfd_8_0.QA.n1 56.1505
R2053 pfd_8_0.QA.n3 pfd_8_0.QA.t0 24.0005
R2054 pfd_8_0.QA.n3 pfd_8_0.QA.t2 24.0005
R2055 pfd_8_0.DOWN_input.t5 pfd_8_0.DOWN_input.t4 377.567
R2056 pfd_8_0.DOWN_input.n2 pfd_8_0.DOWN_input.t3 326.658
R2057 pfd_8_0.DOWN_input pfd_8_0.DOWN_input.n3 237.65
R2058 pfd_8_0.DOWN_input.n0 pfd_8_0.DOWN_input.t1 229.127
R2059 pfd_8_0.DOWN_input.n3 pfd_8_0.DOWN_input.n2 196.817
R2060 pfd_8_0.DOWN_input.n0 pfd_8_0.DOWN_input.t0 158.335
R2061 pfd_8_0.DOWN_input.n1 pfd_8_0.DOWN_input.t2 158.335
R2062 pfd_8_0.DOWN_input.n1 pfd_8_0.DOWN_input.n0 121.6
R2063 pfd_8_0.DOWN_input.t4 pfd_8_0.DOWN_input.n2 92.3838
R2064 pfd_8_0.DOWN_input.n3 pfd_8_0.DOWN_input.t5 92.3838
R2065 pfd_8_0.DOWN_input pfd_8_0.DOWN_input.n1 3.2005
R2066 pfd_8_0.QB.t4 pfd_8_0.QB.t3 835.467
R2067 pfd_8_0.QB.n1 pfd_8_0.QB.t4 564.496
R2068 pfd_8_0.QB.n2 pfd_8_0.QB.t5 517.347
R2069 pfd_8_0.QB.n0 pfd_8_0.QB.t7 514.134
R2070 pfd_8_0.QB.n1 pfd_8_0.QB.n0 455.219
R2071 pfd_8_0.QB.n5 pfd_8_0.QB.n2 363.2
R2072 pfd_8_0.QB.n0 pfd_8_0.QB.t8 273.134
R2073 pfd_8_0.QB.n4 pfd_8_0.QB.n3 244.716
R2074 pfd_8_0.QB.n2 pfd_8_0.QB.t6 228.148
R2075 pfd_8_0.QB.n4 pfd_8_0.QB.t2 221.411
R2076 pfd_8_0.QB.n5 pfd_8_0.QB.n4 54.3734
R2077 pfd_8_0.QB pfd_8_0.QB.n1 26.7568
R2078 pfd_8_0.QB.n3 pfd_8_0.QB.t1 24.0005
R2079 pfd_8_0.QB.n3 pfd_8_0.QB.t0 24.0005
R2080 pfd_8_0.QB pfd_8_0.QB.n5 6.4005
R2081 a_1910_2020.t0 a_1910_2020.t1 48.0005
R2082 a_6220_5810.n4 a_6220_5810.t12 317.317
R2083 a_6220_5810.n2 a_6220_5810.t11 317.317
R2084 a_6220_5810.n5 a_6220_5810.n4 257.067
R2085 a_6220_5810.n3 a_6220_5810.n2 257.067
R2086 a_6220_5810.n10 a_6220_5810.n9 257.067
R2087 a_6220_5810.t0 a_6220_5810.n12 194.478
R2088 a_6220_5810.n8 a_6220_5810.n7 152
R2089 a_6220_5810.n12 a_6220_5810.n11 152
R2090 a_6220_5810.n1 a_6220_5810.n0 120.981
R2091 a_6220_5810.n7 a_6220_5810.n6 117.781
R2092 a_6220_5810.n7 a_6220_5810.n1 108.8
R2093 a_6220_5810.n8 a_6220_5810.n5 85.6894
R2094 a_6220_5810.n11 a_6220_5810.n3 85.6894
R2095 a_6220_5810.n11 a_6220_5810.n10 85.6894
R2096 a_6220_5810.n9 a_6220_5810.n8 85.6894
R2097 a_6220_5810.n4 a_6220_5810.t10 60.2505
R2098 a_6220_5810.n5 a_6220_5810.t1 60.2505
R2099 a_6220_5810.n2 a_6220_5810.t9 60.2505
R2100 a_6220_5810.n3 a_6220_5810.t3 60.2505
R2101 a_6220_5810.n10 a_6220_5810.t7 60.2505
R2102 a_6220_5810.n9 a_6220_5810.t5 60.2505
R2103 a_6220_5810.n6 a_6220_5810.t6 24.0005
R2104 a_6220_5810.n6 a_6220_5810.t2 24.0005
R2105 a_6220_5810.n0 a_6220_5810.t4 24.0005
R2106 a_6220_5810.n0 a_6220_5810.t8 24.0005
R2107 a_6220_5810.n12 a_6220_5810.n1 3.2005
R2108 pfd_8_0.UP_PFD_b.n0 pfd_8_0.UP_PFD_b.t2 441.834
R2109 pfd_8_0.UP_PFD_b.n0 pfd_8_0.UP_PFD_b.t3 313.3
R2110 pfd_8_0.UP_PFD_b.n1 pfd_8_0.UP_PFD_b.n0 235.201
R2111 pfd_8_0.UP_PFD_b.t1 pfd_8_0.UP_PFD_b.n1 219.528
R2112 pfd_8_0.UP_PFD_b.n1 pfd_8_0.UP_PFD_b.t0 167.935
R2113 pfd_8_0.UP.n0 pfd_8_0.UP.t5 1205
R2114 pfd_8_0.UP.n2 pfd_8_0.UP.t4 522.168
R2115 pfd_8_0.UP.n1 pfd_8_0.UP.n0 441.834
R2116 pfd_8_0.UP.n3 pfd_8_0.UP.n2 235.201
R2117 pfd_8_0.UP.t1 pfd_8_0.UP.n3 229.127
R2118 pfd_8_0.UP.n1 pfd_8_0.UP.t3 217.905
R2119 pfd_8_0.UP.n0 pfd_8_0.UP.t2 208.868
R2120 pfd_8_0.UP.n3 pfd_8_0.UP.t0 158.335
R2121 pfd_8_0.UP.n2 pfd_8_0.UP.n1 15.063
R2122 pfd_8_0.E.n4 pfd_8_0.E.n0 1319.38
R2123 pfd_8_0.E.n0 pfd_8_0.E.t3 562.333
R2124 pfd_8_0.E.n2 pfd_8_0.E.t5 388.813
R2125 pfd_8_0.E.n2 pfd_8_0.E.t4 356.68
R2126 pfd_8_0.E.n3 pfd_8_0.E.n2 232
R2127 pfd_8_0.E.n0 pfd_8_0.E.t6 224.934
R2128 pfd_8_0.E.t0 pfd_8_0.E.n4 221.411
R2129 pfd_8_0.E.n3 pfd_8_0.E.n1 157.278
R2130 pfd_8_0.E.n4 pfd_8_0.E.n3 90.64
R2131 pfd_8_0.E.n1 pfd_8_0.E.t2 24.0005
R2132 pfd_8_0.E.n1 pfd_8_0.E.t1 24.0005
R2133 pfd_8_0.E_b.n0 pfd_8_0.E_b.t4 517.347
R2134 pfd_8_0.E_b.n2 pfd_8_0.E_b.n0 417.574
R2135 pfd_8_0.E_b.n2 pfd_8_0.E_b.n1 244.716
R2136 pfd_8_0.E_b.n0 pfd_8_0.E_b.t3 228.148
R2137 pfd_8_0.E_b.t0 pfd_8_0.E_b.n2 221.411
R2138 pfd_8_0.E_b.n1 pfd_8_0.E_b.t2 24.0005
R2139 pfd_8_0.E_b.n1 pfd_8_0.E_b.t1 24.0005
R2140 a_1390_1400.t0 a_1390_1400.t1 39.4005
R2141 pfd_8_0.QB_b.t6 pfd_8_0.QB_b.t4 1188.93
R2142 pfd_8_0.QB_b pfd_8_0.QB_b.n2 899.734
R2143 pfd_8_0.QB_b.t4 pfd_8_0.QB_b.t3 835.467
R2144 pfd_8_0.QB_b.n2 pfd_8_0.QB_b.t5 562.333
R2145 pfd_8_0.QB_b pfd_8_0.QB_b.n1 419.647
R2146 pfd_8_0.QB_b.n1 pfd_8_0.QB_b.n0 247.917
R2147 pfd_8_0.QB_b.n2 pfd_8_0.QB_b.t6 224.934
R2148 pfd_8_0.QB_b.n1 pfd_8_0.QB_b.t1 221.411
R2149 pfd_8_0.QB_b.n0 pfd_8_0.QB_b.t2 24.0005
R2150 pfd_8_0.QB_b.n0 pfd_8_0.QB_b.t0 24.0005
R2151 a_870_640.t0 a_870_640.t1 39.4005
R2152 a_9360_3514.t1 a_9360_3514.t0 323.964
R2153 loop_filter_2_0.R1_C1.t0 loop_filter_2_0.R1_C1.t1 167.429
R2154 a_2530_190.t1 a_2530_190.n2 500.086
R2155 a_2530_190.n0 a_2530_190.t2 465.933
R2156 a_2530_190.t1 a_2530_190.n2 461.389
R2157 a_2530_190.n1 a_2530_190.n0 392.623
R2158 a_2530_190.n0 a_2530_190.t3 321.334
R2159 a_2530_190.n1 a_2530_190.t0 177.577
R2160 a_2530_190.n2 a_2530_190.n1 48.3899
R2161 a_2200_190.t1 a_2200_190.n2 500.086
R2162 a_2200_190.n1 a_2200_190.n0 473.334
R2163 a_2200_190.n0 a_2200_190.t2 465.933
R2164 a_2200_190.t1 a_2200_190.n2 461.389
R2165 a_2200_190.n0 a_2200_190.t3 321.334
R2166 a_2200_190.n1 a_2200_190.t0 177.577
R2167 a_2200_190.n2 a_2200_190.n1 48.3898
R2168 pfd_8_0.F.n4 pfd_8_0.F.n0 1319.38
R2169 pfd_8_0.F.n0 pfd_8_0.F.t3 562.333
R2170 pfd_8_0.F.n2 pfd_8_0.F.t5 388.813
R2171 pfd_8_0.F.n2 pfd_8_0.F.t6 356.68
R2172 pfd_8_0.F.n3 pfd_8_0.F.n2 232
R2173 pfd_8_0.F.n0 pfd_8_0.F.t4 224.934
R2174 pfd_8_0.F.t1 pfd_8_0.F.n4 221.411
R2175 pfd_8_0.F.n3 pfd_8_0.F.n1 157.278
R2176 pfd_8_0.F.n4 pfd_8_0.F.n3 90.64
R2177 pfd_8_0.F.n1 pfd_8_0.F.t2 24.0005
R2178 pfd_8_0.F.n1 pfd_8_0.F.t0 24.0005
R2179 a_9360_6440.t0 a_9360_6440.t1 245.883
R2180 pfd_8_0.F_b.n0 pfd_8_0.F_b.t3 517.347
R2181 pfd_8_0.F_b.n2 pfd_8_0.F_b.n0 417.574
R2182 pfd_8_0.F_b.n2 pfd_8_0.F_b.n1 244.716
R2183 pfd_8_0.F_b.n0 pfd_8_0.F_b.t4 228.148
R2184 pfd_8_0.F_b.t0 pfd_8_0.F_b.n2 221.411
R2185 pfd_8_0.F_b.n1 pfd_8_0.F_b.t2 24.0005
R2186 pfd_8_0.F_b.n1 pfd_8_0.F_b.t1 24.0005
R2187 a_1390_640.t0 a_1390_640.t1 39.4005
R2188 a_490_640.t0 a_490_640.t1 39.4005
R2189 a_490_1400.t0 a_490_1400.t1 39.4005
R2190 pfd_8_0.Reset.n1 pfd_8_0.Reset.t3 562.333
R2191 pfd_8_0.Reset.n2 pfd_8_0.Reset.n1 480.45
R2192 pfd_8_0.Reset.n0 pfd_8_0.Reset.t4 417.733
R2193 pfd_8_0.Reset.n0 pfd_8_0.Reset.t5 369.534
R2194 pfd_8_0.Reset.n3 pfd_8_0.Reset.n2 328.733
R2195 pfd_8_0.Reset.t1 pfd_8_0.Reset.n3 288.37
R2196 pfd_8_0.Reset.n1 pfd_8_0.Reset.t2 224.934
R2197 pfd_8_0.Reset.n3 pfd_8_0.Reset.t0 177.577
R2198 pfd_8_0.Reset.n2 pfd_8_0.Reset.n0 176.733
R2199 a_1870_190.t1 a_1870_190.n2 500.086
R2200 a_1870_190.n1 a_1870_190.n0 473.334
R2201 a_1870_190.n0 a_1870_190.t2 465.933
R2202 a_1870_190.t1 a_1870_190.n2 461.389
R2203 a_1870_190.n0 a_1870_190.t3 321.334
R2204 a_1870_190.n1 a_1870_190.t0 177.577
R2205 a_1870_190.n2 a_1870_190.n1 48.3898
R2206 a_n30_640.t0 a_n30_640.t1 39.4005
R2207 F_VCO.n0 F_VCO.t0 514.134
R2208 F_VCO.n0 F_VCO.t1 273.134
R2209 F_VCO F_VCO.n0 216.9
C0 pfd_8_0.QA pfd_8_0.QB 0.074487f
C1 VDDA pfd_8_0.DOWN_input 0.221484f
C2 F_VCO VDDA 0.12889f
C3 F_VCO pfd_8_0.QB_b 0.039516f
C4 opamp_cell_4_0.p_bias V_OUT 0.048995f
C5 F_VCO pfd_8_0.QB 0.058558f
C6 I_IN VDDA 0.541032f
C7 opamp_cell_4_0.VIN+ V_OUT 1.59847f
C8 pfd_8_0.QA F_REF 0.056f
C9 V_OUT pfd_8_0.DOWN_input 0.388147f
C10 pfd_8_0.QA_b pfd_8_0.QA 0.422694f
C11 pfd_8_0.QB_b VDDA 0.511838f
C12 pfd_8_0.QA_b F_REF 0.027208f
C13 opamp_cell_4_0.p_bias opamp_cell_4_0.VIN+ 0.100967f
C14 opamp_cell_4_0.VIN+ pfd_8_0.DOWN_input 0.080549f
C15 VDDA pfd_8_0.QB 2.7499f
C16 V_OUT VDDA 0.878147f
C17 pfd_8_0.QB_b pfd_8_0.QB 0.388258f
C18 pfd_8_0.QA VDDA 0.550605f
C19 I_IN opamp_cell_4_0.VIN+ 0.166322f
C20 I_IN pfd_8_0.DOWN_input 0.928029f
C21 VDDA F_REF 0.098433f
C22 opamp_cell_4_0.p_bias VDDA 2.86573f
C23 pfd_8_0.QA_b VDDA 0.52066f
C24 opamp_cell_4_0.VIN+ VDDA 0.832915f
C25 F_VCO GNDA 0.389374f
C26 I_IN GNDA 2.83598f
C27 F_REF GNDA 0.277742f
C28 V_OUT GNDA 24.468657f
C29 VDDA GNDA 44.497326f
C30 pfd_8_0.DOWN_input GNDA 3.03064f
C31 pfd_8_0.QB_b GNDA 1.05311f
C32 pfd_8_0.QB GNDA 1.307381f
C33 pfd_8_0.QA GNDA 3.10102f
C34 pfd_8_0.QA_b GNDA 1.05138f
C35 opamp_cell_4_0.VIN+ GNDA 2.37749f
C36 opamp_cell_4_0.p_bias GNDA 3.954681f
C37 loop_filter_2_0.R1_C1.t1 GNDA 2.39887f
C38 pfd_8_0.QB.t7 GNDA 0.066708f
C39 pfd_8_0.QB.t8 GNDA 0.031333f
C40 pfd_8_0.QB.n0 GNDA 0.096363f
C41 pfd_8_0.QB.t3 GNDA 0.066708f
C42 pfd_8_0.QB.t4 GNDA 0.100569f
C43 pfd_8_0.QB.n1 GNDA 1.20598f
C44 pfd_8_0.QB.t5 GNDA 0.067367f
C45 pfd_8_0.QB.t6 GNDA 0.029539f
C46 pfd_8_0.QB.n2 GNDA 0.170164f
C47 pfd_8_0.QB.t2 GNDA 0.14186f
C48 pfd_8_0.QB.t1 GNDA 0.026953f
C49 pfd_8_0.QB.t0 GNDA 0.026953f
C50 pfd_8_0.QB.n3 GNDA 0.143916f
C51 pfd_8_0.QB.n4 GNDA 0.255686f
C52 pfd_8_0.QB.n5 GNDA 0.218372f
C53 opamp_cell_4_0.p_bias.t0 GNDA 1.66267f
C54 opamp_cell_4_0.p_bias.t2 GNDA 0.019693f
C55 opamp_cell_4_0.p_bias.t6 GNDA 0.019693f
C56 opamp_cell_4_0.p_bias.n0 GNDA 0.054067f
C57 opamp_cell_4_0.p_bias.t8 GNDA 0.019693f
C58 opamp_cell_4_0.p_bias.t4 GNDA 0.019693f
C59 opamp_cell_4_0.p_bias.n1 GNDA 0.054067f
C60 opamp_cell_4_0.p_bias.n2 GNDA 0.068502f
C61 opamp_cell_4_0.p_bias.t1 GNDA 0.054353f
C62 opamp_cell_4_0.p_bias.t3 GNDA 0.054353f
C63 opamp_cell_4_0.p_bias.t7 GNDA 0.054353f
C64 opamp_cell_4_0.p_bias.t11 GNDA 0.054353f
C65 opamp_cell_4_0.p_bias.t9 GNDA 0.074733f
C66 opamp_cell_4_0.p_bias.n3 GNDA 0.04185f
C67 opamp_cell_4_0.p_bias.n4 GNDA 0.029697f
C68 opamp_cell_4_0.p_bias.n5 GNDA 0.012761f
C69 opamp_cell_4_0.p_bias.n6 GNDA 0.029697f
C70 opamp_cell_4_0.p_bias.n7 GNDA 0.029697f
C71 opamp_cell_4_0.p_bias.t5 GNDA 0.054353f
C72 opamp_cell_4_0.p_bias.t12 GNDA 0.054353f
C73 opamp_cell_4_0.p_bias.t10 GNDA 0.074733f
C74 opamp_cell_4_0.p_bias.n8 GNDA 0.04185f
C75 opamp_cell_4_0.p_bias.n9 GNDA 0.029697f
C76 opamp_cell_4_0.p_bias.n10 GNDA 0.012761f
C77 opamp_cell_4_0.p_bias.n11 GNDA 0.120625f
C78 pfd_8_0.opamp_out.t12 GNDA 0.957954f
C79 pfd_8_0.opamp_out.t11 GNDA 0.957546f
C80 pfd_8_0.opamp_out.n6 GNDA 0.012958f
C81 pfd_8_0.opamp_out.t14 GNDA 0.012873f
C82 pfd_8_0.opamp_out.t1 GNDA 0.012026f
C83 pfd_8_0.opamp_out.n13 GNDA 0.015342f
C84 pfd_8_0.opamp_out.n14 GNDA 0.081091f
C85 pfd_8_0.opamp_out.n15 GNDA 0.047633f
C86 VDDA.t47 GNDA 0.031725f
C87 VDDA.t25 GNDA 0.011505f
C88 VDDA.n24 GNDA 0.012601f
C89 VDDA.t41 GNDA 0.031725f
C90 VDDA.n41 GNDA 0.029191f
C91 VDDA.n44 GNDA 0.011371f
C92 VDDA.t30 GNDA 0.106924f
C93 VDDA.n50 GNDA 0.011371f
C94 VDDA.n51 GNDA 0.011371f
C95 VDDA.n79 GNDA 0.010592f
C96 VDDA.n87 GNDA 0.052094f
C97 VDDA.t107 GNDA 0.12759f
C98 VDDA.t62 GNDA 0.064549f
C99 VDDA.t60 GNDA 0.064549f
C100 VDDA.t58 GNDA 0.064549f
C101 VDDA.t64 GNDA 0.064549f
C102 VDDA.t113 GNDA 0.073238f
C103 VDDA.n92 GNDA 0.014257f
C104 VDDA.t95 GNDA 0.018775f
C105 VDDA.n97 GNDA 0.014214f
C106 VDDA.n107 GNDA 0.10303f
C107 VDDA.t86 GNDA 0.049653f
C108 VDDA.t96 GNDA 0.032274f
C109 VDDA.t84 GNDA 0.038481f
C110 VDDA.t85 GNDA 0.043446f
C111 VDDA.t43 GNDA 0.032274f
C112 VDDA.t29 GNDA 0.049653f
C113 VDDA.t12 GNDA 0.032274f
C114 VDDA.t127 GNDA 0.035998f
C115 VDDA.t87 GNDA 0.045929f
C116 VDDA.t18 GNDA 0.063308f
C117 VDDA.t22 GNDA 0.067032f
C118 VDDA.n108 GNDA 0.053501f
C119 VDDA.t36 GNDA 0.040964f
C120 VDDA.t92 GNDA 0.040964f
C121 VDDA.t0 GNDA 0.040964f
C122 VDDA.t45 GNDA 0.032274f
C123 VDDA.t81 GNDA 0.049653f
C124 VDDA.t14 GNDA 0.032274f
C125 VDDA.t70 GNDA 0.038481f
C126 VDDA.t49 GNDA 0.043446f
C127 VDDA.t16 GNDA 0.032274f
C128 VDDA.t89 GNDA 0.049653f
C129 VDDA.t100 GNDA 0.040964f
C130 VDDA.n112 GNDA 0.01694f
C131 VDDA.n113 GNDA 0.048391f
C132 VDDA.t99 GNDA 0.019159f
C133 VDDA.n116 GNDA 0.014214f
C134 VDDA.n123 GNDA 0.013387f
C135 VDDA.n125 GNDA 0.039154f
C136 VDDA.n126 GNDA 0.047295f
C137 VDDA.n127 GNDA 0.014257f
C138 VDDA.n130 GNDA 0.011731f
C139 VDDA.n131 GNDA 0.034084f
C140 VDDA.n132 GNDA 0.034247f
C141 VDDA.n140 GNDA 0.033211f
C142 VDDA.n147 GNDA 0.033211f
C143 VDDA.n154 GNDA 0.033211f
C144 VDDA.n161 GNDA 0.033211f
C145 VDDA.n171 GNDA 0.022301f
C146 VDDA.n175 GNDA 0.011371f
C147 VDDA.t103 GNDA 0.047265f
C148 VDDA.n182 GNDA 0.010613f
C149 VDDA.n185 GNDA 0.010613f
C150 VDDA.n188 GNDA 0.010959f
C151 VDDA.n189 GNDA 0.015421f
C152 VDDA.n191 GNDA 0.010959f
C153 VDDA.n192 GNDA 0.015421f
C154 VDDA.n211 GNDA 0.010959f
C155 VDDA.n214 GNDA 0.010959f
C156 VDDA.t109 GNDA 0.018893f
C157 VDDA.t51 GNDA 0.048364f
C158 VDDA.t56 GNDA 0.048364f
C159 VDDA.t68 GNDA 0.048364f
C160 VDDA.t72 GNDA 0.048364f
C161 VDDA.t110 GNDA 0.047265f
C162 VDDA.n225 GNDA 0.042868f
C163 VDDA.n230 GNDA 0.011371f
C164 VDDA.n231 GNDA 0.010959f
C165 VDDA.n232 GNDA 0.015617f
C166 VDDA.n239 GNDA 0.014663f
C167 VDDA.n246 GNDA 0.015421f
C168 VDDA.n254 GNDA 0.015421f
C169 VDDA.n255 GNDA 0.010959f
C170 VDDA.n256 GNDA 0.011371f
C171 VDDA.t102 GNDA 0.017827f
C172 VDDA.t116 GNDA 0.017827f
C173 VDDA.n259 GNDA 0.013686f
C174 VDDA.n260 GNDA 0.011371f
C175 VDDA.n261 GNDA 0.012894f
C176 VDDA.n263 GNDA 0.046166f
C177 VDDA.t117 GNDA 0.047265f
C178 VDDA.t10 GNDA 0.048364f
C179 VDDA.t34 GNDA 0.048364f
C180 VDDA.t26 GNDA 0.048364f
C181 VDDA.t4 GNDA 0.048364f
C182 VDDA.t120 GNDA 0.047265f
C183 VDDA.n269 GNDA 0.042868f
C184 VDDA.t119 GNDA 0.018893f
C185 VDDA.n279 GNDA 0.015519f
C186 VDDA.n280 GNDA 0.162393f
C187 VDDA.n281 GNDA 0.029102f
C188 VDDA.n283 GNDA 0.011371f
C189 VDDA.t123 GNDA 0.111624f
C190 VDDA.t40 GNDA 0.121024f
C191 VDDA.n290 GNDA 0.09165f
C192 VDDA.n314 GNDA 0.09165f
C193 VDDA.t83 GNDA 0.09165f
C194 VDDA.t74 GNDA 0.031725f
C195 VDDA.n327 GNDA 0.045825f
C196 VDDA.n335 GNDA 0.045825f
C197 VDDA.t76 GNDA 0.031725f
C198 VDDA.t38 GNDA 0.031725f
C199 VDDA.n343 GNDA 0.064625f
C200 VDDA.n346 GNDA 0.011371f
C201 VDDA.n355 GNDA 0.011371f
C202 VDDA.n363 GNDA 0.099874f
C203 VDDA.t2 GNDA 0.09165f
C204 VDDA.n369 GNDA 0.09165f
C205 VDDA.n405 GNDA 0.045825f
C206 VDDA.t53 GNDA 0.0282f
C207 VDDA.t24 GNDA 0.029375f
C208 VDDA.n411 GNDA 0.045825f
C209 VDDA.n427 GNDA 0.062275f
C210 VDDA.n446 GNDA 0.069325f
C211 VDDA.t66 GNDA 0.057575f
C212 VDDA.t80 GNDA 0.122199f
C213 VDDA.t28 GNDA 0.122199f
C214 VDDA.t6 GNDA 0.057575f
C215 VDDA.n470 GNDA 0.06345f
C216 VDDA.t20 GNDA 0.057575f
C217 VDDA.t9 GNDA 0.122199f
C218 VDDA.t8 GNDA 0.122199f
C219 VDDA.t32 GNDA 0.057575f
C220 VDDA.n483 GNDA 0.064625f
C221 a_5970_4630.t10 GNDA 0.030769f
C222 a_5970_4630.n0 GNDA 0.124795f
C223 a_5970_4630.t12 GNDA 0.020325f
C224 a_5970_4630.t3 GNDA 0.020325f
C225 a_5970_4630.t6 GNDA 0.020325f
C226 a_5970_4630.n1 GNDA 0.044943f
C227 a_5970_4630.t5 GNDA 0.020325f
C228 a_5970_4630.t8 GNDA 0.020325f
C229 a_5970_4630.n2 GNDA 0.044943f
C230 a_5970_4630.t9 GNDA 0.077457f
C231 a_5970_4630.t7 GNDA 0.030769f
C232 a_5970_4630.n3 GNDA 0.097952f
C233 a_5970_4630.n4 GNDA 0.087903f
C234 a_5970_4630.n5 GNDA 0.089425f
C235 a_5970_4630.t2 GNDA 0.050813f
C236 a_5970_4630.t1 GNDA 0.050813f
C237 a_5970_4630.n6 GNDA 0.295522f
C238 a_5970_4630.t0 GNDA 0.050813f
C239 a_5970_4630.t4 GNDA 0.050813f
C240 a_5970_4630.n7 GNDA 0.144587f
C241 a_5970_4630.n8 GNDA 0.360746f
C242 a_5970_4630.n9 GNDA 0.13437f
C243 a_5970_4630.n10 GNDA 0.085474f
C244 a_5970_4630.n11 GNDA 0.045257f
C245 a_5970_4630.t11 GNDA 0.100208f
C246 V_OUT.n2 GNDA 0.013587f
C247 V_OUT.n5 GNDA 0.011683f
C248 V_OUT.t7 GNDA 4.37553f
C249 V_OUT.n9 GNDA 0.09694f
C250 V_OUT.n10 GNDA 0.038187f
.ends

