magic
tech sky130A
magscale 1 2
timestamp 1751468147
<< nwell >>
rect 5200 6520 6640 7190
rect 6900 6520 9420 7190
rect 9680 6530 11120 7190
rect 5290 5400 6100 6060
rect 6360 5190 9960 6260
rect 10220 5400 11310 6060
rect 5260 4220 8020 4880
rect 8300 4220 11060 4880
<< pwell >>
rect 40 6840 2480 7330
rect 40 6310 2420 6800
rect 430 5890 2050 6270
rect 2610 6090 5020 7060
rect 430 5470 2050 5850
rect 2940 5680 4610 6050
rect 6150 3600 7650 4190
rect 8670 3600 10170 4190
rect -90 3370 260 3450
rect 5670 2650 8130 3540
rect 8190 2650 10650 3540
rect 5870 2100 10440 2610
rect 8599 2060 9202 2062
rect 5320 1460 7060 2060
rect 7110 1460 9210 2060
rect 9260 1460 11000 2060
<< nmos >>
rect 6340 3800 6380 3900
rect 6460 3800 6500 3900
rect 6580 3800 6620 3900
rect 6700 3800 6740 3900
rect 6820 3800 6860 3900
rect 6940 3800 6980 3900
rect 7060 3800 7100 3900
rect 7180 3800 7220 3900
rect 7300 3800 7340 3900
rect 7420 3800 7460 3900
rect 8860 3800 8900 3900
rect 8980 3800 9020 3900
rect 9100 3800 9140 3900
rect 9220 3800 9260 3900
rect 9340 3800 9380 3900
rect 9460 3800 9500 3900
rect 9580 3800 9620 3900
rect 9700 3800 9740 3900
rect 9820 3800 9860 3900
rect 9940 3800 9980 3900
rect 5860 2850 6860 3350
rect 6940 2850 7940 3350
rect 8380 2850 9380 3350
rect 9460 2850 10460 3350
rect 6120 2210 8120 2410
rect 8200 2210 10200 2410
rect 5510 1660 5610 1860
rect 5690 1660 5790 1860
rect 5870 1660 5970 1860
rect 6050 1660 6150 1860
rect 6230 1660 6330 1860
rect 6410 1660 6510 1860
rect 6590 1660 6690 1860
rect 6770 1660 6870 1860
rect 7300 1660 7400 1860
rect 7480 1660 7580 1860
rect 7660 1660 7760 1860
rect 7840 1660 7940 1860
rect 8020 1660 8120 1860
rect 8200 1660 8300 1860
rect 8380 1660 8480 1860
rect 8560 1660 8660 1860
rect 8740 1660 8840 1860
rect 8920 1660 9020 1860
rect 9450 1660 9550 1860
rect 9630 1660 9730 1860
rect 9810 1660 9910 1860
rect 9990 1660 10090 1860
rect 10170 1660 10270 1860
rect 10350 1660 10450 1860
rect 10530 1660 10630 1860
rect 10710 1660 10810 1860
<< pmos >>
rect 5420 6760 5520 6960
rect 5600 6760 5700 6960
rect 5780 6760 5880 6960
rect 5960 6760 6060 6960
rect 6140 6760 6240 6960
rect 6320 6760 6420 6960
rect 7120 6760 7220 6960
rect 7300 6760 7400 6960
rect 7480 6760 7580 6960
rect 7660 6760 7760 6960
rect 7840 6760 7940 6960
rect 8020 6760 8120 6960
rect 8200 6760 8300 6960
rect 8380 6760 8480 6960
rect 8560 6760 8660 6960
rect 8740 6760 8840 6960
rect 8920 6760 9020 6960
rect 9100 6760 9200 6960
rect 9900 6760 10000 6960
rect 10080 6760 10180 6960
rect 10260 6760 10360 6960
rect 10440 6760 10540 6960
rect 10620 6760 10720 6960
rect 10800 6760 10900 6960
rect 5510 5630 5540 5830
rect 5620 5630 5650 5830
rect 5730 5630 5760 5830
rect 5840 5630 5870 5830
rect 6580 5430 6680 6030
rect 6760 5430 6860 6030
rect 6940 5430 7040 6030
rect 7120 5430 7220 6030
rect 7300 5430 7400 6030
rect 7480 5430 7580 6030
rect 7660 5430 7760 6030
rect 7840 5430 7940 6030
rect 8020 5430 8120 6030
rect 8200 5430 8300 6030
rect 8380 5430 8480 6030
rect 8560 5430 8660 6030
rect 8740 5430 8840 6030
rect 8920 5430 9020 6030
rect 9100 5430 9200 6030
rect 9280 5430 9380 6030
rect 9460 5430 9560 6030
rect 9640 5430 9740 6030
rect 10440 5630 10540 5830
rect 10620 5630 10720 5830
rect 10800 5630 10900 5830
rect 10980 5630 11080 5830
rect 5480 4450 5520 4650
rect 5600 4450 5640 4650
rect 5720 4450 5760 4650
rect 5840 4450 5880 4650
rect 5960 4450 6000 4650
rect 6080 4450 6120 4650
rect 6200 4450 6240 4650
rect 6320 4450 6360 4650
rect 6440 4450 6480 4650
rect 6560 4450 6600 4650
rect 6680 4450 6720 4650
rect 6800 4450 6840 4650
rect 6920 4450 6960 4650
rect 7040 4450 7080 4650
rect 7160 4450 7200 4650
rect 7280 4450 7320 4650
rect 7400 4450 7440 4650
rect 7520 4450 7560 4650
rect 7640 4450 7680 4650
rect 7760 4450 7800 4650
rect 8520 4450 8560 4650
rect 8640 4450 8680 4650
rect 8760 4450 8800 4650
rect 8880 4450 8920 4650
rect 9000 4450 9040 4650
rect 9120 4450 9160 4650
rect 9240 4450 9280 4650
rect 9360 4450 9400 4650
rect 9480 4450 9520 4650
rect 9600 4450 9640 4650
rect 9720 4450 9760 4650
rect 9840 4450 9880 4650
rect 9960 4450 10000 4650
rect 10080 4450 10120 4650
rect 10200 4450 10240 4650
rect 10320 4450 10360 4650
rect 10440 4450 10480 4650
rect 10560 4450 10600 4650
rect 10680 4450 10720 4650
rect 10800 4450 10840 4650
<< ndiff >>
rect 6260 3870 6340 3900
rect 6260 3830 6280 3870
rect 6320 3830 6340 3870
rect 6260 3800 6340 3830
rect 6380 3870 6460 3900
rect 6380 3830 6400 3870
rect 6440 3830 6460 3870
rect 6380 3800 6460 3830
rect 6500 3870 6580 3900
rect 6500 3830 6520 3870
rect 6560 3830 6580 3870
rect 6500 3800 6580 3830
rect 6620 3870 6700 3900
rect 6620 3830 6640 3870
rect 6680 3830 6700 3870
rect 6620 3800 6700 3830
rect 6740 3870 6820 3900
rect 6740 3830 6760 3870
rect 6800 3830 6820 3870
rect 6740 3800 6820 3830
rect 6860 3870 6940 3900
rect 6860 3830 6880 3870
rect 6920 3830 6940 3870
rect 6860 3800 6940 3830
rect 6980 3870 7060 3900
rect 6980 3830 7000 3870
rect 7040 3830 7060 3870
rect 6980 3800 7060 3830
rect 7100 3870 7180 3900
rect 7100 3830 7120 3870
rect 7160 3830 7180 3870
rect 7100 3800 7180 3830
rect 7220 3870 7300 3900
rect 7220 3830 7240 3870
rect 7280 3830 7300 3870
rect 7220 3800 7300 3830
rect 7340 3870 7420 3900
rect 7340 3830 7360 3870
rect 7400 3830 7420 3870
rect 7340 3800 7420 3830
rect 7460 3870 7540 3900
rect 7460 3830 7480 3870
rect 7520 3830 7540 3870
rect 7460 3800 7540 3830
rect 8780 3870 8860 3900
rect 8780 3830 8800 3870
rect 8840 3830 8860 3870
rect 8780 3800 8860 3830
rect 8900 3870 8980 3900
rect 8900 3830 8920 3870
rect 8960 3830 8980 3870
rect 8900 3800 8980 3830
rect 9020 3870 9100 3900
rect 9020 3830 9040 3870
rect 9080 3830 9100 3870
rect 9020 3800 9100 3830
rect 9140 3870 9220 3900
rect 9140 3830 9160 3870
rect 9200 3830 9220 3870
rect 9140 3800 9220 3830
rect 9260 3870 9340 3900
rect 9260 3830 9280 3870
rect 9320 3830 9340 3870
rect 9260 3800 9340 3830
rect 9380 3870 9460 3900
rect 9380 3830 9400 3870
rect 9440 3830 9460 3870
rect 9380 3800 9460 3830
rect 9500 3870 9580 3900
rect 9500 3830 9520 3870
rect 9560 3830 9580 3870
rect 9500 3800 9580 3830
rect 9620 3870 9700 3900
rect 9620 3830 9640 3870
rect 9680 3830 9700 3870
rect 9620 3800 9700 3830
rect 9740 3870 9820 3900
rect 9740 3830 9760 3870
rect 9800 3830 9820 3870
rect 9740 3800 9820 3830
rect 9860 3870 9940 3900
rect 9860 3830 9880 3870
rect 9920 3830 9940 3870
rect 9860 3800 9940 3830
rect 9980 3870 10060 3900
rect 9980 3830 10000 3870
rect 10040 3830 10060 3870
rect 9980 3800 10060 3830
rect 5780 3320 5860 3350
rect 5780 3280 5800 3320
rect 5840 3280 5860 3320
rect 5780 3220 5860 3280
rect 5780 3180 5800 3220
rect 5840 3180 5860 3220
rect 5780 3120 5860 3180
rect 5780 3080 5800 3120
rect 5840 3080 5860 3120
rect 5780 3020 5860 3080
rect 5780 2980 5800 3020
rect 5840 2980 5860 3020
rect 5780 2920 5860 2980
rect 5780 2880 5800 2920
rect 5840 2880 5860 2920
rect 5780 2850 5860 2880
rect 6860 3320 6940 3350
rect 6860 3280 6880 3320
rect 6920 3280 6940 3320
rect 6860 3220 6940 3280
rect 6860 3180 6880 3220
rect 6920 3180 6940 3220
rect 6860 3120 6940 3180
rect 6860 3080 6880 3120
rect 6920 3080 6940 3120
rect 6860 3020 6940 3080
rect 6860 2980 6880 3020
rect 6920 2980 6940 3020
rect 6860 2920 6940 2980
rect 6860 2880 6880 2920
rect 6920 2880 6940 2920
rect 6860 2850 6940 2880
rect 7940 3320 8020 3350
rect 7940 3280 7960 3320
rect 8000 3280 8020 3320
rect 7940 3220 8020 3280
rect 7940 3180 7960 3220
rect 8000 3180 8020 3220
rect 7940 3120 8020 3180
rect 7940 3080 7960 3120
rect 8000 3080 8020 3120
rect 7940 3020 8020 3080
rect 7940 2980 7960 3020
rect 8000 2980 8020 3020
rect 7940 2920 8020 2980
rect 7940 2880 7960 2920
rect 8000 2880 8020 2920
rect 7940 2850 8020 2880
rect 8300 3320 8380 3350
rect 8300 3280 8320 3320
rect 8360 3280 8380 3320
rect 8300 3220 8380 3280
rect 8300 3180 8320 3220
rect 8360 3180 8380 3220
rect 8300 3120 8380 3180
rect 8300 3080 8320 3120
rect 8360 3080 8380 3120
rect 8300 3020 8380 3080
rect 8300 2980 8320 3020
rect 8360 2980 8380 3020
rect 8300 2920 8380 2980
rect 8300 2880 8320 2920
rect 8360 2880 8380 2920
rect 8300 2850 8380 2880
rect 9380 3320 9460 3350
rect 9380 3280 9400 3320
rect 9440 3280 9460 3320
rect 9380 3220 9460 3280
rect 9380 3180 9400 3220
rect 9440 3180 9460 3220
rect 9380 3120 9460 3180
rect 9380 3080 9400 3120
rect 9440 3080 9460 3120
rect 9380 3020 9460 3080
rect 9380 2980 9400 3020
rect 9440 2980 9460 3020
rect 9380 2920 9460 2980
rect 9380 2880 9400 2920
rect 9440 2880 9460 2920
rect 9380 2850 9460 2880
rect 10460 3320 10540 3350
rect 10460 3280 10480 3320
rect 10520 3280 10540 3320
rect 10460 3220 10540 3280
rect 10460 3180 10480 3220
rect 10520 3180 10540 3220
rect 10460 3120 10540 3180
rect 10460 3080 10480 3120
rect 10520 3080 10540 3120
rect 10460 3020 10540 3080
rect 10460 2980 10480 3020
rect 10520 2980 10540 3020
rect 10460 2920 10540 2980
rect 10460 2880 10480 2920
rect 10520 2880 10540 2920
rect 10460 2850 10540 2880
rect 6040 2380 6120 2410
rect 6040 2340 6060 2380
rect 6100 2340 6120 2380
rect 6040 2280 6120 2340
rect 6040 2240 6060 2280
rect 6100 2240 6120 2280
rect 6040 2210 6120 2240
rect 8120 2380 8200 2410
rect 8120 2340 8140 2380
rect 8180 2340 8200 2380
rect 8120 2280 8200 2340
rect 8120 2240 8140 2280
rect 8180 2240 8200 2280
rect 8120 2210 8200 2240
rect 10200 2380 10280 2410
rect 10200 2340 10220 2380
rect 10260 2340 10280 2380
rect 10200 2280 10280 2340
rect 10200 2240 10220 2280
rect 10260 2240 10280 2280
rect 10200 2210 10280 2240
rect 5430 1830 5510 1860
rect 5430 1790 5450 1830
rect 5490 1790 5510 1830
rect 5430 1730 5510 1790
rect 5430 1690 5450 1730
rect 5490 1690 5510 1730
rect 5430 1660 5510 1690
rect 5610 1830 5690 1860
rect 5610 1790 5630 1830
rect 5670 1790 5690 1830
rect 5610 1730 5690 1790
rect 5610 1690 5630 1730
rect 5670 1690 5690 1730
rect 5610 1660 5690 1690
rect 5790 1830 5870 1860
rect 5790 1790 5810 1830
rect 5850 1790 5870 1830
rect 5790 1730 5870 1790
rect 5790 1690 5810 1730
rect 5850 1690 5870 1730
rect 5790 1660 5870 1690
rect 5970 1830 6050 1860
rect 5970 1790 5990 1830
rect 6030 1790 6050 1830
rect 5970 1730 6050 1790
rect 5970 1690 5990 1730
rect 6030 1690 6050 1730
rect 5970 1660 6050 1690
rect 6150 1830 6230 1860
rect 6150 1790 6170 1830
rect 6210 1790 6230 1830
rect 6150 1730 6230 1790
rect 6150 1690 6170 1730
rect 6210 1690 6230 1730
rect 6150 1660 6230 1690
rect 6330 1830 6410 1860
rect 6330 1790 6350 1830
rect 6390 1790 6410 1830
rect 6330 1730 6410 1790
rect 6330 1690 6350 1730
rect 6390 1690 6410 1730
rect 6330 1660 6410 1690
rect 6510 1830 6590 1860
rect 6510 1790 6530 1830
rect 6570 1790 6590 1830
rect 6510 1730 6590 1790
rect 6510 1690 6530 1730
rect 6570 1690 6590 1730
rect 6510 1660 6590 1690
rect 6690 1830 6770 1860
rect 6690 1790 6710 1830
rect 6750 1790 6770 1830
rect 6690 1730 6770 1790
rect 6690 1690 6710 1730
rect 6750 1690 6770 1730
rect 6690 1660 6770 1690
rect 6870 1830 6950 1860
rect 6870 1790 6890 1830
rect 6930 1790 6950 1830
rect 6870 1730 6950 1790
rect 6870 1690 6890 1730
rect 6930 1690 6950 1730
rect 6870 1660 6950 1690
rect 7220 1830 7300 1860
rect 7220 1790 7240 1830
rect 7280 1790 7300 1830
rect 7220 1730 7300 1790
rect 7220 1690 7240 1730
rect 7280 1690 7300 1730
rect 7220 1660 7300 1690
rect 7400 1830 7480 1860
rect 7400 1790 7420 1830
rect 7460 1790 7480 1830
rect 7400 1730 7480 1790
rect 7400 1690 7420 1730
rect 7460 1690 7480 1730
rect 7400 1660 7480 1690
rect 7580 1830 7660 1860
rect 7580 1790 7600 1830
rect 7640 1790 7660 1830
rect 7580 1730 7660 1790
rect 7580 1690 7600 1730
rect 7640 1690 7660 1730
rect 7580 1660 7660 1690
rect 7760 1830 7840 1860
rect 7760 1790 7780 1830
rect 7820 1790 7840 1830
rect 7760 1730 7840 1790
rect 7760 1690 7780 1730
rect 7820 1690 7840 1730
rect 7760 1660 7840 1690
rect 7940 1830 8020 1860
rect 7940 1790 7960 1830
rect 8000 1790 8020 1830
rect 7940 1730 8020 1790
rect 7940 1690 7960 1730
rect 8000 1690 8020 1730
rect 7940 1660 8020 1690
rect 8120 1830 8200 1860
rect 8120 1790 8140 1830
rect 8180 1790 8200 1830
rect 8120 1730 8200 1790
rect 8120 1690 8140 1730
rect 8180 1690 8200 1730
rect 8120 1660 8200 1690
rect 8300 1830 8380 1860
rect 8300 1790 8320 1830
rect 8360 1790 8380 1830
rect 8300 1730 8380 1790
rect 8300 1690 8320 1730
rect 8360 1690 8380 1730
rect 8300 1660 8380 1690
rect 8480 1830 8560 1860
rect 8480 1790 8500 1830
rect 8540 1790 8560 1830
rect 8480 1730 8560 1790
rect 8480 1690 8500 1730
rect 8540 1690 8560 1730
rect 8480 1660 8560 1690
rect 8660 1830 8740 1860
rect 8660 1790 8680 1830
rect 8720 1790 8740 1830
rect 8660 1730 8740 1790
rect 8660 1690 8680 1730
rect 8720 1690 8740 1730
rect 8660 1660 8740 1690
rect 8840 1830 8920 1860
rect 8840 1790 8860 1830
rect 8900 1790 8920 1830
rect 8840 1730 8920 1790
rect 8840 1690 8860 1730
rect 8900 1690 8920 1730
rect 8840 1660 8920 1690
rect 9020 1830 9100 1860
rect 9020 1790 9040 1830
rect 9080 1790 9100 1830
rect 9020 1730 9100 1790
rect 9020 1690 9040 1730
rect 9080 1690 9100 1730
rect 9020 1660 9100 1690
rect 9370 1830 9450 1860
rect 9370 1790 9390 1830
rect 9430 1790 9450 1830
rect 9370 1730 9450 1790
rect 9370 1690 9390 1730
rect 9430 1690 9450 1730
rect 9370 1660 9450 1690
rect 9550 1830 9630 1860
rect 9550 1790 9570 1830
rect 9610 1790 9630 1830
rect 9550 1730 9630 1790
rect 9550 1690 9570 1730
rect 9610 1690 9630 1730
rect 9550 1660 9630 1690
rect 9730 1830 9810 1860
rect 9730 1790 9750 1830
rect 9790 1790 9810 1830
rect 9730 1730 9810 1790
rect 9730 1690 9750 1730
rect 9790 1690 9810 1730
rect 9730 1660 9810 1690
rect 9910 1830 9990 1860
rect 9910 1790 9930 1830
rect 9970 1790 9990 1830
rect 9910 1730 9990 1790
rect 9910 1690 9930 1730
rect 9970 1690 9990 1730
rect 9910 1660 9990 1690
rect 10090 1830 10170 1860
rect 10090 1790 10110 1830
rect 10150 1790 10170 1830
rect 10090 1730 10170 1790
rect 10090 1690 10110 1730
rect 10150 1690 10170 1730
rect 10090 1660 10170 1690
rect 10270 1830 10350 1860
rect 10270 1790 10290 1830
rect 10330 1790 10350 1830
rect 10270 1730 10350 1790
rect 10270 1690 10290 1730
rect 10330 1690 10350 1730
rect 10270 1660 10350 1690
rect 10450 1830 10530 1860
rect 10450 1790 10470 1830
rect 10510 1790 10530 1830
rect 10450 1730 10530 1790
rect 10450 1690 10470 1730
rect 10510 1690 10530 1730
rect 10450 1660 10530 1690
rect 10630 1830 10710 1860
rect 10630 1790 10650 1830
rect 10690 1790 10710 1830
rect 10630 1730 10710 1790
rect 10630 1690 10650 1730
rect 10690 1690 10710 1730
rect 10630 1660 10710 1690
rect 10810 1830 10890 1860
rect 10810 1790 10830 1830
rect 10870 1790 10890 1830
rect 10810 1730 10890 1790
rect 10810 1690 10830 1730
rect 10870 1690 10890 1730
rect 10810 1660 10890 1690
<< pdiff >>
rect 5340 6930 5420 6960
rect 5340 6786 5360 6930
rect 5400 6786 5420 6930
rect 5340 6760 5420 6786
rect 5520 6930 5600 6960
rect 5520 6786 5540 6930
rect 5580 6786 5600 6930
rect 5520 6760 5600 6786
rect 5700 6930 5780 6960
rect 5700 6786 5720 6930
rect 5760 6786 5780 6930
rect 5700 6760 5780 6786
rect 5880 6930 5960 6960
rect 5880 6786 5900 6930
rect 5940 6786 5960 6930
rect 5880 6760 5960 6786
rect 6060 6930 6140 6960
rect 6060 6786 6080 6930
rect 6120 6786 6140 6930
rect 6060 6760 6140 6786
rect 6240 6930 6320 6960
rect 6240 6786 6260 6930
rect 6300 6786 6320 6930
rect 6240 6760 6320 6786
rect 6420 6930 6500 6960
rect 6420 6786 6440 6930
rect 6480 6786 6500 6930
rect 6420 6760 6500 6786
rect 7040 6930 7120 6960
rect 7040 6890 7060 6930
rect 7100 6890 7120 6930
rect 7040 6830 7120 6890
rect 7040 6790 7060 6830
rect 7100 6790 7120 6830
rect 7040 6760 7120 6790
rect 7220 6930 7300 6960
rect 7220 6890 7240 6930
rect 7280 6890 7300 6930
rect 7220 6830 7300 6890
rect 7220 6790 7240 6830
rect 7280 6790 7300 6830
rect 7220 6760 7300 6790
rect 7400 6930 7480 6960
rect 7400 6890 7420 6930
rect 7460 6890 7480 6930
rect 7400 6830 7480 6890
rect 7400 6790 7420 6830
rect 7460 6790 7480 6830
rect 7400 6760 7480 6790
rect 7580 6930 7660 6960
rect 7580 6890 7600 6930
rect 7640 6890 7660 6930
rect 7580 6830 7660 6890
rect 7580 6790 7600 6830
rect 7640 6790 7660 6830
rect 7580 6760 7660 6790
rect 7760 6930 7840 6960
rect 7760 6890 7780 6930
rect 7820 6890 7840 6930
rect 7760 6830 7840 6890
rect 7760 6790 7780 6830
rect 7820 6790 7840 6830
rect 7760 6760 7840 6790
rect 7940 6930 8020 6960
rect 7940 6890 7960 6930
rect 8000 6890 8020 6930
rect 7940 6830 8020 6890
rect 7940 6790 7960 6830
rect 8000 6790 8020 6830
rect 7940 6760 8020 6790
rect 8120 6930 8200 6960
rect 8120 6890 8140 6930
rect 8180 6890 8200 6930
rect 8120 6830 8200 6890
rect 8120 6790 8140 6830
rect 8180 6790 8200 6830
rect 8120 6760 8200 6790
rect 8300 6930 8380 6960
rect 8300 6890 8320 6930
rect 8360 6890 8380 6930
rect 8300 6830 8380 6890
rect 8300 6790 8320 6830
rect 8360 6790 8380 6830
rect 8300 6760 8380 6790
rect 8480 6930 8560 6960
rect 8480 6890 8500 6930
rect 8540 6890 8560 6930
rect 8480 6830 8560 6890
rect 8480 6790 8500 6830
rect 8540 6790 8560 6830
rect 8480 6760 8560 6790
rect 8660 6930 8740 6960
rect 8660 6890 8680 6930
rect 8720 6890 8740 6930
rect 8660 6830 8740 6890
rect 8660 6790 8680 6830
rect 8720 6790 8740 6830
rect 8660 6760 8740 6790
rect 8840 6930 8920 6960
rect 8840 6890 8860 6930
rect 8900 6890 8920 6930
rect 8840 6830 8920 6890
rect 8840 6790 8860 6830
rect 8900 6790 8920 6830
rect 8840 6760 8920 6790
rect 9020 6930 9100 6960
rect 9020 6890 9040 6930
rect 9080 6890 9100 6930
rect 9020 6830 9100 6890
rect 9020 6790 9040 6830
rect 9080 6790 9100 6830
rect 9020 6760 9100 6790
rect 9200 6930 9280 6960
rect 9200 6890 9220 6930
rect 9260 6890 9280 6930
rect 9200 6830 9280 6890
rect 9200 6790 9220 6830
rect 9260 6790 9280 6830
rect 9200 6760 9280 6790
rect 9820 6930 9900 6960
rect 9820 6790 9840 6930
rect 9880 6790 9900 6930
rect 9820 6760 9900 6790
rect 10000 6930 10080 6960
rect 10000 6790 10020 6930
rect 10060 6790 10080 6930
rect 10000 6760 10080 6790
rect 10180 6930 10260 6960
rect 10180 6790 10200 6930
rect 10240 6790 10260 6930
rect 10180 6760 10260 6790
rect 10360 6930 10440 6960
rect 10360 6790 10380 6930
rect 10420 6790 10440 6930
rect 10360 6760 10440 6790
rect 10540 6930 10620 6960
rect 10540 6790 10560 6930
rect 10600 6790 10620 6930
rect 10540 6760 10620 6790
rect 10720 6930 10800 6960
rect 10720 6790 10740 6930
rect 10780 6790 10800 6930
rect 10720 6760 10800 6790
rect 10900 6930 10980 6960
rect 10900 6790 10920 6930
rect 10960 6790 10980 6930
rect 10900 6760 10980 6790
rect 5430 5800 5510 5830
rect 5430 5760 5450 5800
rect 5490 5760 5510 5800
rect 5430 5700 5510 5760
rect 5430 5660 5450 5700
rect 5490 5660 5510 5700
rect 5430 5630 5510 5660
rect 5540 5800 5620 5830
rect 5540 5760 5560 5800
rect 5600 5760 5620 5800
rect 5540 5700 5620 5760
rect 5540 5660 5560 5700
rect 5600 5660 5620 5700
rect 5540 5630 5620 5660
rect 5650 5800 5730 5830
rect 5650 5760 5670 5800
rect 5710 5760 5730 5800
rect 5650 5700 5730 5760
rect 5650 5660 5670 5700
rect 5710 5660 5730 5700
rect 5650 5630 5730 5660
rect 5760 5800 5840 5830
rect 5760 5760 5780 5800
rect 5820 5760 5840 5800
rect 5760 5700 5840 5760
rect 5760 5660 5780 5700
rect 5820 5660 5840 5700
rect 5760 5630 5840 5660
rect 5870 5800 5950 5830
rect 5870 5760 5890 5800
rect 5930 5760 5950 5800
rect 5870 5700 5950 5760
rect 5870 5660 5890 5700
rect 5930 5660 5950 5700
rect 5870 5630 5950 5660
rect 6500 6000 6580 6030
rect 6500 5960 6520 6000
rect 6560 5960 6580 6000
rect 6500 5900 6580 5960
rect 6500 5860 6520 5900
rect 6560 5860 6580 5900
rect 6500 5800 6580 5860
rect 6500 5760 6520 5800
rect 6560 5760 6580 5800
rect 6500 5700 6580 5760
rect 6500 5660 6520 5700
rect 6560 5660 6580 5700
rect 6500 5600 6580 5660
rect 6500 5560 6520 5600
rect 6560 5560 6580 5600
rect 6500 5500 6580 5560
rect 6500 5460 6520 5500
rect 6560 5460 6580 5500
rect 6500 5430 6580 5460
rect 6680 6000 6760 6030
rect 6680 5960 6700 6000
rect 6740 5960 6760 6000
rect 6680 5900 6760 5960
rect 6680 5860 6700 5900
rect 6740 5860 6760 5900
rect 6680 5800 6760 5860
rect 6680 5760 6700 5800
rect 6740 5760 6760 5800
rect 6680 5700 6760 5760
rect 6680 5660 6700 5700
rect 6740 5660 6760 5700
rect 6680 5600 6760 5660
rect 6680 5560 6700 5600
rect 6740 5560 6760 5600
rect 6680 5500 6760 5560
rect 6680 5460 6700 5500
rect 6740 5460 6760 5500
rect 6680 5430 6760 5460
rect 6860 6000 6940 6030
rect 6860 5960 6880 6000
rect 6920 5960 6940 6000
rect 6860 5900 6940 5960
rect 6860 5860 6880 5900
rect 6920 5860 6940 5900
rect 6860 5800 6940 5860
rect 6860 5760 6880 5800
rect 6920 5760 6940 5800
rect 6860 5700 6940 5760
rect 6860 5660 6880 5700
rect 6920 5660 6940 5700
rect 6860 5600 6940 5660
rect 6860 5560 6880 5600
rect 6920 5560 6940 5600
rect 6860 5500 6940 5560
rect 6860 5460 6880 5500
rect 6920 5460 6940 5500
rect 6860 5430 6940 5460
rect 7040 6000 7120 6030
rect 7040 5960 7060 6000
rect 7100 5960 7120 6000
rect 7040 5900 7120 5960
rect 7040 5860 7060 5900
rect 7100 5860 7120 5900
rect 7040 5800 7120 5860
rect 7040 5760 7060 5800
rect 7100 5760 7120 5800
rect 7040 5700 7120 5760
rect 7040 5660 7060 5700
rect 7100 5660 7120 5700
rect 7040 5600 7120 5660
rect 7040 5560 7060 5600
rect 7100 5560 7120 5600
rect 7040 5500 7120 5560
rect 7040 5460 7060 5500
rect 7100 5460 7120 5500
rect 7040 5430 7120 5460
rect 7220 6000 7300 6030
rect 7220 5960 7240 6000
rect 7280 5960 7300 6000
rect 7220 5900 7300 5960
rect 7220 5860 7240 5900
rect 7280 5860 7300 5900
rect 7220 5800 7300 5860
rect 7220 5760 7240 5800
rect 7280 5760 7300 5800
rect 7220 5700 7300 5760
rect 7220 5660 7240 5700
rect 7280 5660 7300 5700
rect 7220 5600 7300 5660
rect 7220 5560 7240 5600
rect 7280 5560 7300 5600
rect 7220 5500 7300 5560
rect 7220 5460 7240 5500
rect 7280 5460 7300 5500
rect 7220 5430 7300 5460
rect 7400 6000 7480 6030
rect 7400 5960 7420 6000
rect 7460 5960 7480 6000
rect 7400 5900 7480 5960
rect 7400 5860 7420 5900
rect 7460 5860 7480 5900
rect 7400 5800 7480 5860
rect 7400 5760 7420 5800
rect 7460 5760 7480 5800
rect 7400 5700 7480 5760
rect 7400 5660 7420 5700
rect 7460 5660 7480 5700
rect 7400 5600 7480 5660
rect 7400 5560 7420 5600
rect 7460 5560 7480 5600
rect 7400 5500 7480 5560
rect 7400 5460 7420 5500
rect 7460 5460 7480 5500
rect 7400 5430 7480 5460
rect 7580 6000 7660 6030
rect 7580 5960 7600 6000
rect 7640 5960 7660 6000
rect 7580 5900 7660 5960
rect 7580 5860 7600 5900
rect 7640 5860 7660 5900
rect 7580 5800 7660 5860
rect 7580 5760 7600 5800
rect 7640 5760 7660 5800
rect 7580 5700 7660 5760
rect 7580 5660 7600 5700
rect 7640 5660 7660 5700
rect 7580 5600 7660 5660
rect 7580 5560 7600 5600
rect 7640 5560 7660 5600
rect 7580 5500 7660 5560
rect 7580 5460 7600 5500
rect 7640 5460 7660 5500
rect 7580 5430 7660 5460
rect 7760 6000 7840 6030
rect 7760 5960 7780 6000
rect 7820 5960 7840 6000
rect 7760 5900 7840 5960
rect 7760 5860 7780 5900
rect 7820 5860 7840 5900
rect 7760 5800 7840 5860
rect 7760 5760 7780 5800
rect 7820 5760 7840 5800
rect 7760 5700 7840 5760
rect 7760 5660 7780 5700
rect 7820 5660 7840 5700
rect 7760 5600 7840 5660
rect 7760 5560 7780 5600
rect 7820 5560 7840 5600
rect 7760 5500 7840 5560
rect 7760 5460 7780 5500
rect 7820 5460 7840 5500
rect 7760 5430 7840 5460
rect 7940 6000 8020 6030
rect 7940 5960 7960 6000
rect 8000 5960 8020 6000
rect 7940 5900 8020 5960
rect 7940 5860 7960 5900
rect 8000 5860 8020 5900
rect 7940 5800 8020 5860
rect 7940 5760 7960 5800
rect 8000 5760 8020 5800
rect 7940 5700 8020 5760
rect 7940 5660 7960 5700
rect 8000 5660 8020 5700
rect 7940 5600 8020 5660
rect 7940 5560 7960 5600
rect 8000 5560 8020 5600
rect 7940 5500 8020 5560
rect 7940 5460 7960 5500
rect 8000 5460 8020 5500
rect 7940 5430 8020 5460
rect 8120 6000 8200 6030
rect 8120 5960 8140 6000
rect 8180 5960 8200 6000
rect 8120 5900 8200 5960
rect 8120 5860 8140 5900
rect 8180 5860 8200 5900
rect 8120 5800 8200 5860
rect 8120 5760 8140 5800
rect 8180 5760 8200 5800
rect 8120 5700 8200 5760
rect 8120 5660 8140 5700
rect 8180 5660 8200 5700
rect 8120 5600 8200 5660
rect 8120 5560 8140 5600
rect 8180 5560 8200 5600
rect 8120 5500 8200 5560
rect 8120 5460 8140 5500
rect 8180 5460 8200 5500
rect 8120 5430 8200 5460
rect 8300 6000 8380 6030
rect 8300 5960 8320 6000
rect 8360 5960 8380 6000
rect 8300 5900 8380 5960
rect 8300 5860 8320 5900
rect 8360 5860 8380 5900
rect 8300 5800 8380 5860
rect 8300 5760 8320 5800
rect 8360 5760 8380 5800
rect 8300 5700 8380 5760
rect 8300 5660 8320 5700
rect 8360 5660 8380 5700
rect 8300 5600 8380 5660
rect 8300 5560 8320 5600
rect 8360 5560 8380 5600
rect 8300 5500 8380 5560
rect 8300 5460 8320 5500
rect 8360 5460 8380 5500
rect 8300 5430 8380 5460
rect 8480 6000 8560 6030
rect 8480 5960 8500 6000
rect 8540 5960 8560 6000
rect 8480 5900 8560 5960
rect 8480 5860 8500 5900
rect 8540 5860 8560 5900
rect 8480 5800 8560 5860
rect 8480 5760 8500 5800
rect 8540 5760 8560 5800
rect 8480 5700 8560 5760
rect 8480 5660 8500 5700
rect 8540 5660 8560 5700
rect 8480 5600 8560 5660
rect 8480 5560 8500 5600
rect 8540 5560 8560 5600
rect 8480 5500 8560 5560
rect 8480 5460 8500 5500
rect 8540 5460 8560 5500
rect 8480 5430 8560 5460
rect 8660 6000 8740 6030
rect 8660 5960 8680 6000
rect 8720 5960 8740 6000
rect 8660 5900 8740 5960
rect 8660 5860 8680 5900
rect 8720 5860 8740 5900
rect 8660 5800 8740 5860
rect 8660 5760 8680 5800
rect 8720 5760 8740 5800
rect 8660 5700 8740 5760
rect 8660 5660 8680 5700
rect 8720 5660 8740 5700
rect 8660 5600 8740 5660
rect 8660 5560 8680 5600
rect 8720 5560 8740 5600
rect 8660 5500 8740 5560
rect 8660 5460 8680 5500
rect 8720 5460 8740 5500
rect 8660 5430 8740 5460
rect 8840 6000 8920 6030
rect 8840 5960 8860 6000
rect 8900 5960 8920 6000
rect 8840 5900 8920 5960
rect 8840 5860 8860 5900
rect 8900 5860 8920 5900
rect 8840 5800 8920 5860
rect 8840 5760 8860 5800
rect 8900 5760 8920 5800
rect 8840 5700 8920 5760
rect 8840 5660 8860 5700
rect 8900 5660 8920 5700
rect 8840 5600 8920 5660
rect 8840 5560 8860 5600
rect 8900 5560 8920 5600
rect 8840 5500 8920 5560
rect 8840 5460 8860 5500
rect 8900 5460 8920 5500
rect 8840 5430 8920 5460
rect 9020 6000 9100 6030
rect 9020 5960 9040 6000
rect 9080 5960 9100 6000
rect 9020 5900 9100 5960
rect 9020 5860 9040 5900
rect 9080 5860 9100 5900
rect 9020 5800 9100 5860
rect 9020 5760 9040 5800
rect 9080 5760 9100 5800
rect 9020 5700 9100 5760
rect 9020 5660 9040 5700
rect 9080 5660 9100 5700
rect 9020 5600 9100 5660
rect 9020 5560 9040 5600
rect 9080 5560 9100 5600
rect 9020 5500 9100 5560
rect 9020 5460 9040 5500
rect 9080 5460 9100 5500
rect 9020 5430 9100 5460
rect 9200 6000 9280 6030
rect 9200 5960 9220 6000
rect 9260 5960 9280 6000
rect 9200 5900 9280 5960
rect 9200 5860 9220 5900
rect 9260 5860 9280 5900
rect 9200 5800 9280 5860
rect 9200 5760 9220 5800
rect 9260 5760 9280 5800
rect 9200 5700 9280 5760
rect 9200 5660 9220 5700
rect 9260 5660 9280 5700
rect 9200 5600 9280 5660
rect 9200 5560 9220 5600
rect 9260 5560 9280 5600
rect 9200 5500 9280 5560
rect 9200 5460 9220 5500
rect 9260 5460 9280 5500
rect 9200 5430 9280 5460
rect 9380 6000 9460 6030
rect 9380 5960 9400 6000
rect 9440 5960 9460 6000
rect 9380 5900 9460 5960
rect 9380 5860 9400 5900
rect 9440 5860 9460 5900
rect 9380 5800 9460 5860
rect 9380 5760 9400 5800
rect 9440 5760 9460 5800
rect 9380 5700 9460 5760
rect 9380 5660 9400 5700
rect 9440 5660 9460 5700
rect 9380 5600 9460 5660
rect 9380 5560 9400 5600
rect 9440 5560 9460 5600
rect 9380 5500 9460 5560
rect 9380 5460 9400 5500
rect 9440 5460 9460 5500
rect 9380 5430 9460 5460
rect 9560 6000 9640 6030
rect 9560 5960 9580 6000
rect 9620 5960 9640 6000
rect 9560 5900 9640 5960
rect 9560 5860 9580 5900
rect 9620 5860 9640 5900
rect 9560 5800 9640 5860
rect 9560 5760 9580 5800
rect 9620 5760 9640 5800
rect 9560 5700 9640 5760
rect 9560 5660 9580 5700
rect 9620 5660 9640 5700
rect 9560 5600 9640 5660
rect 9560 5560 9580 5600
rect 9620 5560 9640 5600
rect 9560 5500 9640 5560
rect 9560 5460 9580 5500
rect 9620 5460 9640 5500
rect 9560 5430 9640 5460
rect 9740 6000 9820 6030
rect 9740 5960 9760 6000
rect 9800 5960 9820 6000
rect 9740 5900 9820 5960
rect 9740 5860 9760 5900
rect 9800 5860 9820 5900
rect 9740 5800 9820 5860
rect 9740 5760 9760 5800
rect 9800 5760 9820 5800
rect 9740 5700 9820 5760
rect 9740 5660 9760 5700
rect 9800 5660 9820 5700
rect 9740 5600 9820 5660
rect 9740 5560 9760 5600
rect 9800 5560 9820 5600
rect 9740 5500 9820 5560
rect 9740 5460 9760 5500
rect 9800 5460 9820 5500
rect 9740 5430 9820 5460
rect 10360 5800 10440 5830
rect 10360 5760 10380 5800
rect 10420 5760 10440 5800
rect 10360 5700 10440 5760
rect 10360 5660 10380 5700
rect 10420 5660 10440 5700
rect 10360 5630 10440 5660
rect 10540 5800 10620 5830
rect 10540 5760 10560 5800
rect 10600 5760 10620 5800
rect 10540 5700 10620 5760
rect 10540 5660 10560 5700
rect 10600 5660 10620 5700
rect 10540 5630 10620 5660
rect 10720 5800 10800 5830
rect 10720 5760 10740 5800
rect 10780 5760 10800 5800
rect 10720 5700 10800 5760
rect 10720 5660 10740 5700
rect 10780 5660 10800 5700
rect 10720 5630 10800 5660
rect 10900 5800 10980 5830
rect 10900 5760 10920 5800
rect 10960 5760 10980 5800
rect 10900 5700 10980 5760
rect 10900 5660 10920 5700
rect 10960 5660 10980 5700
rect 10900 5630 10980 5660
rect 11080 5800 11160 5830
rect 11080 5760 11100 5800
rect 11140 5760 11160 5800
rect 11080 5700 11160 5760
rect 11080 5660 11100 5700
rect 11140 5660 11160 5700
rect 11080 5630 11160 5660
rect 5400 4620 5480 4650
rect 5400 4580 5420 4620
rect 5460 4580 5480 4620
rect 5400 4520 5480 4580
rect 5400 4480 5420 4520
rect 5460 4480 5480 4520
rect 5400 4450 5480 4480
rect 5520 4620 5600 4650
rect 5520 4580 5540 4620
rect 5580 4580 5600 4620
rect 5520 4520 5600 4580
rect 5520 4480 5540 4520
rect 5580 4480 5600 4520
rect 5520 4450 5600 4480
rect 5640 4620 5720 4650
rect 5640 4580 5660 4620
rect 5700 4580 5720 4620
rect 5640 4520 5720 4580
rect 5640 4480 5660 4520
rect 5700 4480 5720 4520
rect 5640 4450 5720 4480
rect 5760 4620 5840 4650
rect 5760 4580 5780 4620
rect 5820 4580 5840 4620
rect 5760 4520 5840 4580
rect 5760 4480 5780 4520
rect 5820 4480 5840 4520
rect 5760 4450 5840 4480
rect 5880 4620 5960 4650
rect 5880 4580 5900 4620
rect 5940 4580 5960 4620
rect 5880 4520 5960 4580
rect 5880 4480 5900 4520
rect 5940 4480 5960 4520
rect 5880 4450 5960 4480
rect 6000 4620 6080 4650
rect 6000 4580 6020 4620
rect 6060 4580 6080 4620
rect 6000 4520 6080 4580
rect 6000 4480 6020 4520
rect 6060 4480 6080 4520
rect 6000 4450 6080 4480
rect 6120 4620 6200 4650
rect 6120 4580 6140 4620
rect 6180 4580 6200 4620
rect 6120 4520 6200 4580
rect 6120 4480 6140 4520
rect 6180 4480 6200 4520
rect 6120 4450 6200 4480
rect 6240 4620 6320 4650
rect 6240 4580 6260 4620
rect 6300 4580 6320 4620
rect 6240 4520 6320 4580
rect 6240 4480 6260 4520
rect 6300 4480 6320 4520
rect 6240 4450 6320 4480
rect 6360 4620 6440 4650
rect 6360 4580 6380 4620
rect 6420 4580 6440 4620
rect 6360 4520 6440 4580
rect 6360 4480 6380 4520
rect 6420 4480 6440 4520
rect 6360 4450 6440 4480
rect 6480 4620 6560 4650
rect 6480 4580 6500 4620
rect 6540 4580 6560 4620
rect 6480 4520 6560 4580
rect 6480 4480 6500 4520
rect 6540 4480 6560 4520
rect 6480 4450 6560 4480
rect 6600 4620 6680 4650
rect 6600 4580 6620 4620
rect 6660 4580 6680 4620
rect 6600 4520 6680 4580
rect 6600 4480 6620 4520
rect 6660 4480 6680 4520
rect 6600 4450 6680 4480
rect 6720 4620 6800 4650
rect 6720 4580 6740 4620
rect 6780 4580 6800 4620
rect 6720 4520 6800 4580
rect 6720 4480 6740 4520
rect 6780 4480 6800 4520
rect 6720 4450 6800 4480
rect 6840 4620 6920 4650
rect 6840 4580 6860 4620
rect 6900 4580 6920 4620
rect 6840 4520 6920 4580
rect 6840 4480 6860 4520
rect 6900 4480 6920 4520
rect 6840 4450 6920 4480
rect 6960 4620 7040 4650
rect 6960 4580 6980 4620
rect 7020 4580 7040 4620
rect 6960 4520 7040 4580
rect 6960 4480 6980 4520
rect 7020 4480 7040 4520
rect 6960 4450 7040 4480
rect 7080 4620 7160 4650
rect 7080 4580 7100 4620
rect 7140 4580 7160 4620
rect 7080 4520 7160 4580
rect 7080 4480 7100 4520
rect 7140 4480 7160 4520
rect 7080 4450 7160 4480
rect 7200 4620 7280 4650
rect 7200 4580 7220 4620
rect 7260 4580 7280 4620
rect 7200 4520 7280 4580
rect 7200 4480 7220 4520
rect 7260 4480 7280 4520
rect 7200 4450 7280 4480
rect 7320 4620 7400 4650
rect 7320 4580 7340 4620
rect 7380 4580 7400 4620
rect 7320 4520 7400 4580
rect 7320 4480 7340 4520
rect 7380 4480 7400 4520
rect 7320 4450 7400 4480
rect 7440 4620 7520 4650
rect 7440 4580 7460 4620
rect 7500 4580 7520 4620
rect 7440 4520 7520 4580
rect 7440 4480 7460 4520
rect 7500 4480 7520 4520
rect 7440 4450 7520 4480
rect 7560 4620 7640 4650
rect 7560 4580 7580 4620
rect 7620 4580 7640 4620
rect 7560 4520 7640 4580
rect 7560 4480 7580 4520
rect 7620 4480 7640 4520
rect 7560 4450 7640 4480
rect 7680 4620 7760 4650
rect 7680 4580 7700 4620
rect 7740 4580 7760 4620
rect 7680 4520 7760 4580
rect 7680 4480 7700 4520
rect 7740 4480 7760 4520
rect 7680 4450 7760 4480
rect 7800 4620 7880 4650
rect 7800 4580 7820 4620
rect 7860 4580 7880 4620
rect 7800 4520 7880 4580
rect 7800 4480 7820 4520
rect 7860 4480 7880 4520
rect 7800 4450 7880 4480
rect 8440 4620 8520 4650
rect 8440 4580 8460 4620
rect 8500 4580 8520 4620
rect 8440 4520 8520 4580
rect 8440 4480 8460 4520
rect 8500 4480 8520 4520
rect 8440 4450 8520 4480
rect 8560 4620 8640 4650
rect 8560 4580 8580 4620
rect 8620 4580 8640 4620
rect 8560 4520 8640 4580
rect 8560 4480 8580 4520
rect 8620 4480 8640 4520
rect 8560 4450 8640 4480
rect 8680 4620 8760 4650
rect 8680 4580 8700 4620
rect 8740 4580 8760 4620
rect 8680 4520 8760 4580
rect 8680 4480 8700 4520
rect 8740 4480 8760 4520
rect 8680 4450 8760 4480
rect 8800 4620 8880 4650
rect 8800 4580 8820 4620
rect 8860 4580 8880 4620
rect 8800 4520 8880 4580
rect 8800 4480 8820 4520
rect 8860 4480 8880 4520
rect 8800 4450 8880 4480
rect 8920 4620 9000 4650
rect 8920 4580 8940 4620
rect 8980 4580 9000 4620
rect 8920 4520 9000 4580
rect 8920 4480 8940 4520
rect 8980 4480 9000 4520
rect 8920 4450 9000 4480
rect 9040 4620 9120 4650
rect 9040 4580 9060 4620
rect 9100 4580 9120 4620
rect 9040 4520 9120 4580
rect 9040 4480 9060 4520
rect 9100 4480 9120 4520
rect 9040 4450 9120 4480
rect 9160 4620 9240 4650
rect 9160 4580 9180 4620
rect 9220 4580 9240 4620
rect 9160 4520 9240 4580
rect 9160 4480 9180 4520
rect 9220 4480 9240 4520
rect 9160 4450 9240 4480
rect 9280 4620 9360 4650
rect 9280 4580 9300 4620
rect 9340 4580 9360 4620
rect 9280 4520 9360 4580
rect 9280 4480 9300 4520
rect 9340 4480 9360 4520
rect 9280 4450 9360 4480
rect 9400 4620 9480 4650
rect 9400 4580 9420 4620
rect 9460 4580 9480 4620
rect 9400 4520 9480 4580
rect 9400 4480 9420 4520
rect 9460 4480 9480 4520
rect 9400 4450 9480 4480
rect 9520 4620 9600 4650
rect 9520 4580 9540 4620
rect 9580 4580 9600 4620
rect 9520 4520 9600 4580
rect 9520 4480 9540 4520
rect 9580 4480 9600 4520
rect 9520 4450 9600 4480
rect 9640 4620 9720 4650
rect 9640 4580 9660 4620
rect 9700 4580 9720 4620
rect 9640 4520 9720 4580
rect 9640 4480 9660 4520
rect 9700 4480 9720 4520
rect 9640 4450 9720 4480
rect 9760 4620 9840 4650
rect 9760 4580 9780 4620
rect 9820 4580 9840 4620
rect 9760 4520 9840 4580
rect 9760 4480 9780 4520
rect 9820 4480 9840 4520
rect 9760 4450 9840 4480
rect 9880 4620 9960 4650
rect 9880 4580 9900 4620
rect 9940 4580 9960 4620
rect 9880 4520 9960 4580
rect 9880 4480 9900 4520
rect 9940 4480 9960 4520
rect 9880 4450 9960 4480
rect 10000 4620 10080 4650
rect 10000 4580 10020 4620
rect 10060 4580 10080 4620
rect 10000 4520 10080 4580
rect 10000 4480 10020 4520
rect 10060 4480 10080 4520
rect 10000 4450 10080 4480
rect 10120 4620 10200 4650
rect 10120 4580 10140 4620
rect 10180 4580 10200 4620
rect 10120 4520 10200 4580
rect 10120 4480 10140 4520
rect 10180 4480 10200 4520
rect 10120 4450 10200 4480
rect 10240 4620 10320 4650
rect 10240 4580 10260 4620
rect 10300 4580 10320 4620
rect 10240 4520 10320 4580
rect 10240 4480 10260 4520
rect 10300 4480 10320 4520
rect 10240 4450 10320 4480
rect 10360 4620 10440 4650
rect 10360 4580 10380 4620
rect 10420 4580 10440 4620
rect 10360 4520 10440 4580
rect 10360 4480 10380 4520
rect 10420 4480 10440 4520
rect 10360 4450 10440 4480
rect 10480 4620 10560 4650
rect 10480 4580 10500 4620
rect 10540 4580 10560 4620
rect 10480 4520 10560 4580
rect 10480 4480 10500 4520
rect 10540 4480 10560 4520
rect 10480 4450 10560 4480
rect 10600 4620 10680 4650
rect 10600 4580 10620 4620
rect 10660 4580 10680 4620
rect 10600 4520 10680 4580
rect 10600 4480 10620 4520
rect 10660 4480 10680 4520
rect 10600 4450 10680 4480
rect 10720 4620 10800 4650
rect 10720 4580 10740 4620
rect 10780 4580 10800 4620
rect 10720 4520 10800 4580
rect 10720 4480 10740 4520
rect 10780 4480 10800 4520
rect 10720 4450 10800 4480
rect 10840 4620 10920 4650
rect 10840 4580 10860 4620
rect 10900 4580 10920 4620
rect 10840 4520 10920 4580
rect 10840 4480 10860 4520
rect 10900 4480 10920 4520
rect 10840 4450 10920 4480
<< ndiffc >>
rect 6280 3830 6320 3870
rect 6400 3830 6440 3870
rect 6520 3830 6560 3870
rect 6640 3830 6680 3870
rect 6760 3830 6800 3870
rect 6880 3830 6920 3870
rect 7000 3830 7040 3870
rect 7120 3830 7160 3870
rect 7240 3830 7280 3870
rect 7360 3830 7400 3870
rect 7480 3830 7520 3870
rect 8800 3830 8840 3870
rect 8920 3830 8960 3870
rect 9040 3830 9080 3870
rect 9160 3830 9200 3870
rect 9280 3830 9320 3870
rect 9400 3830 9440 3870
rect 9520 3830 9560 3870
rect 9640 3830 9680 3870
rect 9760 3830 9800 3870
rect 9880 3830 9920 3870
rect 10000 3830 10040 3870
rect 5800 3280 5840 3320
rect 5800 3180 5840 3220
rect 5800 3080 5840 3120
rect 5800 2980 5840 3020
rect 5800 2880 5840 2920
rect 6880 3280 6920 3320
rect 6880 3180 6920 3220
rect 6880 3080 6920 3120
rect 6880 2980 6920 3020
rect 6880 2880 6920 2920
rect 7960 3280 8000 3320
rect 7960 3180 8000 3220
rect 7960 3080 8000 3120
rect 7960 2980 8000 3020
rect 7960 2880 8000 2920
rect 8320 3280 8360 3320
rect 8320 3180 8360 3220
rect 8320 3080 8360 3120
rect 8320 2980 8360 3020
rect 8320 2880 8360 2920
rect 9400 3280 9440 3320
rect 9400 3180 9440 3220
rect 9400 3080 9440 3120
rect 9400 2980 9440 3020
rect 9400 2880 9440 2920
rect 10480 3280 10520 3320
rect 10480 3180 10520 3220
rect 10480 3080 10520 3120
rect 10480 2980 10520 3020
rect 10480 2880 10520 2920
rect 6060 2340 6100 2380
rect 6060 2240 6100 2280
rect 8140 2340 8180 2380
rect 8140 2240 8180 2280
rect 10220 2340 10260 2380
rect 10220 2240 10260 2280
rect 5450 1790 5490 1830
rect 5450 1690 5490 1730
rect 5630 1790 5670 1830
rect 5630 1690 5670 1730
rect 5810 1790 5850 1830
rect 5810 1690 5850 1730
rect 5990 1790 6030 1830
rect 5990 1690 6030 1730
rect 6170 1790 6210 1830
rect 6170 1690 6210 1730
rect 6350 1790 6390 1830
rect 6350 1690 6390 1730
rect 6530 1790 6570 1830
rect 6530 1690 6570 1730
rect 6710 1790 6750 1830
rect 6710 1690 6750 1730
rect 6890 1790 6930 1830
rect 6890 1690 6930 1730
rect 7240 1790 7280 1830
rect 7240 1690 7280 1730
rect 7420 1790 7460 1830
rect 7420 1690 7460 1730
rect 7600 1790 7640 1830
rect 7600 1690 7640 1730
rect 7780 1790 7820 1830
rect 7780 1690 7820 1730
rect 7960 1790 8000 1830
rect 7960 1690 8000 1730
rect 8140 1790 8180 1830
rect 8140 1690 8180 1730
rect 8320 1790 8360 1830
rect 8320 1690 8360 1730
rect 8500 1790 8540 1830
rect 8500 1690 8540 1730
rect 8680 1790 8720 1830
rect 8680 1690 8720 1730
rect 8860 1790 8900 1830
rect 8860 1690 8900 1730
rect 9040 1790 9080 1830
rect 9040 1690 9080 1730
rect 9390 1790 9430 1830
rect 9390 1690 9430 1730
rect 9570 1790 9610 1830
rect 9570 1690 9610 1730
rect 9750 1790 9790 1830
rect 9750 1690 9790 1730
rect 9930 1790 9970 1830
rect 9930 1690 9970 1730
rect 10110 1790 10150 1830
rect 10110 1690 10150 1730
rect 10290 1790 10330 1830
rect 10290 1690 10330 1730
rect 10470 1790 10510 1830
rect 10470 1690 10510 1730
rect 10650 1790 10690 1830
rect 10650 1690 10690 1730
rect 10830 1790 10870 1830
rect 10830 1690 10870 1730
<< pdiffc >>
rect 5360 6786 5400 6930
rect 5540 6786 5580 6930
rect 5720 6786 5760 6930
rect 5900 6786 5940 6930
rect 6080 6786 6120 6930
rect 6260 6786 6300 6930
rect 6440 6786 6480 6930
rect 7060 6890 7100 6930
rect 7060 6790 7100 6830
rect 7240 6890 7280 6930
rect 7240 6790 7280 6830
rect 7420 6890 7460 6930
rect 7420 6790 7460 6830
rect 7600 6890 7640 6930
rect 7600 6790 7640 6830
rect 7780 6890 7820 6930
rect 7780 6790 7820 6830
rect 7960 6890 8000 6930
rect 7960 6790 8000 6830
rect 8140 6890 8180 6930
rect 8140 6790 8180 6830
rect 8320 6890 8360 6930
rect 8320 6790 8360 6830
rect 8500 6890 8540 6930
rect 8500 6790 8540 6830
rect 8680 6890 8720 6930
rect 8680 6790 8720 6830
rect 8860 6890 8900 6930
rect 8860 6790 8900 6830
rect 9040 6890 9080 6930
rect 9040 6790 9080 6830
rect 9220 6890 9260 6930
rect 9220 6790 9260 6830
rect 9840 6790 9880 6930
rect 10020 6790 10060 6930
rect 10200 6790 10240 6930
rect 10380 6790 10420 6930
rect 10560 6790 10600 6930
rect 10740 6790 10780 6930
rect 10920 6790 10960 6930
rect 5450 5760 5490 5800
rect 5450 5660 5490 5700
rect 5560 5760 5600 5800
rect 5560 5660 5600 5700
rect 5670 5760 5710 5800
rect 5670 5660 5710 5700
rect 5780 5760 5820 5800
rect 5780 5660 5820 5700
rect 5890 5760 5930 5800
rect 5890 5660 5930 5700
rect 6520 5960 6560 6000
rect 6520 5860 6560 5900
rect 6520 5760 6560 5800
rect 6520 5660 6560 5700
rect 6520 5560 6560 5600
rect 6520 5460 6560 5500
rect 6700 5960 6740 6000
rect 6700 5860 6740 5900
rect 6700 5760 6740 5800
rect 6700 5660 6740 5700
rect 6700 5560 6740 5600
rect 6700 5460 6740 5500
rect 6880 5960 6920 6000
rect 6880 5860 6920 5900
rect 6880 5760 6920 5800
rect 6880 5660 6920 5700
rect 6880 5560 6920 5600
rect 6880 5460 6920 5500
rect 7060 5960 7100 6000
rect 7060 5860 7100 5900
rect 7060 5760 7100 5800
rect 7060 5660 7100 5700
rect 7060 5560 7100 5600
rect 7060 5460 7100 5500
rect 7240 5960 7280 6000
rect 7240 5860 7280 5900
rect 7240 5760 7280 5800
rect 7240 5660 7280 5700
rect 7240 5560 7280 5600
rect 7240 5460 7280 5500
rect 7420 5960 7460 6000
rect 7420 5860 7460 5900
rect 7420 5760 7460 5800
rect 7420 5660 7460 5700
rect 7420 5560 7460 5600
rect 7420 5460 7460 5500
rect 7600 5960 7640 6000
rect 7600 5860 7640 5900
rect 7600 5760 7640 5800
rect 7600 5660 7640 5700
rect 7600 5560 7640 5600
rect 7600 5460 7640 5500
rect 7780 5960 7820 6000
rect 7780 5860 7820 5900
rect 7780 5760 7820 5800
rect 7780 5660 7820 5700
rect 7780 5560 7820 5600
rect 7780 5460 7820 5500
rect 7960 5960 8000 6000
rect 7960 5860 8000 5900
rect 7960 5760 8000 5800
rect 7960 5660 8000 5700
rect 7960 5560 8000 5600
rect 7960 5460 8000 5500
rect 8140 5960 8180 6000
rect 8140 5860 8180 5900
rect 8140 5760 8180 5800
rect 8140 5660 8180 5700
rect 8140 5560 8180 5600
rect 8140 5460 8180 5500
rect 8320 5960 8360 6000
rect 8320 5860 8360 5900
rect 8320 5760 8360 5800
rect 8320 5660 8360 5700
rect 8320 5560 8360 5600
rect 8320 5460 8360 5500
rect 8500 5960 8540 6000
rect 8500 5860 8540 5900
rect 8500 5760 8540 5800
rect 8500 5660 8540 5700
rect 8500 5560 8540 5600
rect 8500 5460 8540 5500
rect 8680 5960 8720 6000
rect 8680 5860 8720 5900
rect 8680 5760 8720 5800
rect 8680 5660 8720 5700
rect 8680 5560 8720 5600
rect 8680 5460 8720 5500
rect 8860 5960 8900 6000
rect 8860 5860 8900 5900
rect 8860 5760 8900 5800
rect 8860 5660 8900 5700
rect 8860 5560 8900 5600
rect 8860 5460 8900 5500
rect 9040 5960 9080 6000
rect 9040 5860 9080 5900
rect 9040 5760 9080 5800
rect 9040 5660 9080 5700
rect 9040 5560 9080 5600
rect 9040 5460 9080 5500
rect 9220 5960 9260 6000
rect 9220 5860 9260 5900
rect 9220 5760 9260 5800
rect 9220 5660 9260 5700
rect 9220 5560 9260 5600
rect 9220 5460 9260 5500
rect 9400 5960 9440 6000
rect 9400 5860 9440 5900
rect 9400 5760 9440 5800
rect 9400 5660 9440 5700
rect 9400 5560 9440 5600
rect 9400 5460 9440 5500
rect 9580 5960 9620 6000
rect 9580 5860 9620 5900
rect 9580 5760 9620 5800
rect 9580 5660 9620 5700
rect 9580 5560 9620 5600
rect 9580 5460 9620 5500
rect 9760 5960 9800 6000
rect 9760 5860 9800 5900
rect 9760 5760 9800 5800
rect 9760 5660 9800 5700
rect 9760 5560 9800 5600
rect 9760 5460 9800 5500
rect 10380 5760 10420 5800
rect 10380 5660 10420 5700
rect 10560 5760 10600 5800
rect 10560 5660 10600 5700
rect 10740 5760 10780 5800
rect 10740 5660 10780 5700
rect 10920 5760 10960 5800
rect 10920 5660 10960 5700
rect 11100 5760 11140 5800
rect 11100 5660 11140 5700
rect 5420 4580 5460 4620
rect 5420 4480 5460 4520
rect 5540 4580 5580 4620
rect 5540 4480 5580 4520
rect 5660 4580 5700 4620
rect 5660 4480 5700 4520
rect 5780 4580 5820 4620
rect 5780 4480 5820 4520
rect 5900 4580 5940 4620
rect 5900 4480 5940 4520
rect 6020 4580 6060 4620
rect 6020 4480 6060 4520
rect 6140 4580 6180 4620
rect 6140 4480 6180 4520
rect 6260 4580 6300 4620
rect 6260 4480 6300 4520
rect 6380 4580 6420 4620
rect 6380 4480 6420 4520
rect 6500 4580 6540 4620
rect 6500 4480 6540 4520
rect 6620 4580 6660 4620
rect 6620 4480 6660 4520
rect 6740 4580 6780 4620
rect 6740 4480 6780 4520
rect 6860 4580 6900 4620
rect 6860 4480 6900 4520
rect 6980 4580 7020 4620
rect 6980 4480 7020 4520
rect 7100 4580 7140 4620
rect 7100 4480 7140 4520
rect 7220 4580 7260 4620
rect 7220 4480 7260 4520
rect 7340 4580 7380 4620
rect 7340 4480 7380 4520
rect 7460 4580 7500 4620
rect 7460 4480 7500 4520
rect 7580 4580 7620 4620
rect 7580 4480 7620 4520
rect 7700 4580 7740 4620
rect 7700 4480 7740 4520
rect 7820 4580 7860 4620
rect 7820 4480 7860 4520
rect 8460 4580 8500 4620
rect 8460 4480 8500 4520
rect 8580 4580 8620 4620
rect 8580 4480 8620 4520
rect 8700 4580 8740 4620
rect 8700 4480 8740 4520
rect 8820 4580 8860 4620
rect 8820 4480 8860 4520
rect 8940 4580 8980 4620
rect 8940 4480 8980 4520
rect 9060 4580 9100 4620
rect 9060 4480 9100 4520
rect 9180 4580 9220 4620
rect 9180 4480 9220 4520
rect 9300 4580 9340 4620
rect 9300 4480 9340 4520
rect 9420 4580 9460 4620
rect 9420 4480 9460 4520
rect 9540 4580 9580 4620
rect 9540 4480 9580 4520
rect 9660 4580 9700 4620
rect 9660 4480 9700 4520
rect 9780 4580 9820 4620
rect 9780 4480 9820 4520
rect 9900 4580 9940 4620
rect 9900 4480 9940 4520
rect 10020 4580 10060 4620
rect 10020 4480 10060 4520
rect 10140 4580 10180 4620
rect 10140 4480 10180 4520
rect 10260 4580 10300 4620
rect 10260 4480 10300 4520
rect 10380 4580 10420 4620
rect 10380 4480 10420 4520
rect 10500 4580 10540 4620
rect 10500 4480 10540 4520
rect 10620 4580 10660 4620
rect 10620 4480 10660 4520
rect 10740 4580 10780 4620
rect 10740 4480 10780 4520
rect 10860 4580 10900 4620
rect 10860 4480 10900 4520
<< psubdiff >>
rect 50 7280 1180 7320
rect 1340 7280 2470 7320
rect 50 7160 90 7280
rect 2430 7160 2470 7280
rect 50 6890 90 7000
rect 2430 6890 2470 7000
rect 50 6850 1180 6890
rect 1340 6850 2470 6890
rect 2620 7010 3690 7050
rect 3850 7010 5010 7050
rect 50 6750 1150 6790
rect 1310 6750 2410 6790
rect 50 6630 90 6750
rect 2370 6630 2410 6750
rect 50 6360 90 6470
rect 2370 6360 2410 6470
rect 50 6320 1150 6360
rect 1310 6320 2410 6360
rect 2620 6650 2660 7010
rect 4970 6650 5010 7010
rect 440 6220 1150 6260
rect 1310 6220 2040 6260
rect 440 6160 480 6220
rect 2000 6160 2040 6220
rect 440 5940 480 6000
rect 2620 6140 2660 6490
rect 4970 6140 5010 6490
rect 2620 6100 3690 6140
rect 3850 6100 5010 6140
rect 2000 5940 2040 6000
rect 440 5900 1150 5940
rect 1310 5900 2040 5940
rect 2950 6000 3690 6040
rect 3850 6000 4600 6040
rect 2950 5940 2990 6000
rect 440 5800 1150 5840
rect 1310 5800 2040 5840
rect 440 5740 480 5800
rect 2000 5740 2040 5800
rect 440 5520 480 5580
rect 4560 5940 4600 6000
rect 2950 5730 2990 5780
rect 4560 5730 4600 5780
rect 2950 5690 3690 5730
rect 3850 5690 4600 5730
rect 2000 5520 2040 5580
rect 440 5480 1150 5520
rect 1310 5480 2040 5520
rect 6160 4140 6820 4180
rect 6980 4140 7640 4180
rect 6160 3930 6200 4140
rect 7600 3930 7640 4140
rect 6160 3650 6200 3770
rect 7600 3650 7640 3770
rect 6160 3610 6820 3650
rect 6980 3610 7640 3650
rect 8680 4140 9340 4180
rect 9500 4140 10160 4180
rect 8680 3930 8720 4140
rect 10120 3930 10160 4140
rect 8680 3650 8720 3770
rect 10120 3650 10160 3770
rect 8680 3610 10160 3650
rect 5680 3490 6820 3530
rect 6980 3490 8120 3530
rect -100 3430 200 3460
rect -100 3390 -70 3430
rect -30 3390 30 3430
rect 70 3390 130 3430
rect 170 3390 200 3430
rect -100 3360 200 3390
rect 5680 3180 5720 3490
rect 5680 2700 5720 3020
rect 8080 3180 8120 3490
rect 8080 2700 8120 3020
rect 5680 2660 6820 2700
rect 6980 2660 8120 2700
rect 8200 3490 9340 3530
rect 9500 3490 10640 3530
rect 8200 3180 8240 3490
rect 8200 2700 8240 3020
rect 10600 3180 10640 3490
rect 10600 2700 10640 3020
rect 8200 2660 9340 2700
rect 9500 2660 10640 2700
rect 5880 2560 8080 2600
rect 8240 2560 10430 2600
rect 5880 2390 5920 2560
rect 5880 2150 5920 2230
rect 10390 2390 10430 2560
rect 10390 2150 10430 2230
rect 5880 2110 8080 2150
rect 8240 2110 10430 2150
rect 5330 2010 6110 2050
rect 6270 2010 7050 2050
rect 5330 1840 5370 2010
rect 5330 1510 5370 1680
rect 7010 1840 7050 2010
rect 7010 1510 7050 1680
rect 5330 1470 6110 1510
rect 6270 1470 7050 1510
rect 7120 2010 8080 2050
rect 8240 2010 9200 2050
rect 7120 1840 7160 2010
rect 7120 1510 7160 1680
rect 9160 1840 9200 2010
rect 9160 1510 9200 1680
rect 7120 1470 8080 1510
rect 8240 1470 9200 1510
rect 9270 2010 10050 2050
rect 10210 2010 10990 2050
rect 9270 1840 9310 2010
rect 9270 1510 9310 1680
rect 10950 1840 10990 2010
rect 10950 1510 10990 1680
rect 9270 1470 10050 1510
rect 10210 1470 10990 1510
<< nsubdiff >>
rect 5240 7110 5840 7150
rect 6000 7110 6600 7150
rect 5240 6940 5280 7110
rect 5240 6610 5280 6780
rect 6560 6940 6600 7110
rect 6560 6610 6600 6780
rect 5240 6570 5840 6610
rect 6000 6570 6600 6610
rect 6940 7110 8080 7150
rect 8240 7110 9380 7150
rect 6940 6940 6980 7110
rect 6940 6610 6980 6780
rect 9340 6940 9380 7110
rect 9340 6610 9380 6780
rect 6940 6570 8080 6610
rect 8240 6570 9380 6610
rect 9720 7110 10320 7150
rect 10480 7110 11080 7150
rect 9720 6940 9760 7110
rect 9720 6610 9760 6780
rect 11040 6940 11080 7110
rect 11040 6610 11080 6780
rect 9720 6570 10320 6610
rect 10480 6570 11080 6610
rect 6400 6180 8080 6220
rect 8240 6180 9920 6220
rect 5330 5980 5610 6020
rect 5770 5980 6050 6020
rect 5330 5810 5370 5980
rect 5330 5480 5370 5650
rect 6010 5810 6050 5980
rect 6010 5480 6050 5650
rect 5330 5440 5610 5480
rect 5770 5440 6050 5480
rect 6400 5810 6440 6180
rect 6400 5270 6440 5650
rect 9880 5810 9920 6180
rect 9880 5270 9920 5650
rect 10260 5980 10610 6020
rect 10910 5980 11260 6020
rect 10260 5810 10300 5980
rect 10260 5480 10300 5650
rect 11220 5810 11260 5980
rect 11220 5480 11260 5650
rect 10260 5440 10610 5480
rect 10910 5440 11260 5480
rect 6400 5230 8080 5270
rect 8240 5230 9920 5270
rect 5300 4800 6560 4840
rect 6720 4800 7980 4840
rect 5300 4630 5340 4800
rect 5300 4300 5340 4470
rect 7940 4630 7980 4800
rect 7940 4300 7980 4470
rect 5300 4260 6560 4300
rect 6720 4260 7980 4300
rect 8340 4800 9600 4840
rect 9760 4800 11020 4840
rect 8340 4630 8380 4800
rect 8340 4300 8380 4470
rect 10980 4630 11020 4800
rect 10980 4300 11020 4470
rect 8340 4260 9600 4300
rect 9760 4260 11020 4300
<< psubdiffcont >>
rect 1180 7280 1340 7320
rect 50 7000 90 7160
rect 2430 7000 2470 7160
rect 1180 6850 1340 6890
rect 3690 7010 3850 7050
rect 1150 6750 1310 6790
rect 50 6470 90 6630
rect 2370 6470 2410 6630
rect 1150 6320 1310 6360
rect 2620 6490 2660 6650
rect 1150 6220 1310 6260
rect 440 6000 480 6160
rect 2000 6000 2040 6160
rect 4970 6490 5010 6650
rect 3690 6100 3850 6140
rect 1150 5900 1310 5940
rect 3690 6000 3850 6040
rect 1150 5800 1310 5840
rect 440 5580 480 5740
rect 2000 5580 2040 5740
rect 2950 5780 2990 5940
rect 4560 5780 4600 5940
rect 3690 5690 3850 5730
rect 1150 5480 1310 5520
rect 6820 4140 6980 4180
rect 6160 3770 6200 3930
rect 7600 3770 7640 3930
rect 6820 3610 6980 3650
rect 9340 4140 9500 4180
rect 8680 3770 8720 3930
rect 10120 3770 10160 3930
rect 6820 3490 6980 3530
rect -70 3390 -30 3430
rect 30 3390 70 3430
rect 130 3390 170 3430
rect 5680 3020 5720 3180
rect 8080 3020 8120 3180
rect 6820 2660 6980 2700
rect 9340 3490 9500 3530
rect 8200 3020 8240 3180
rect 10600 3020 10640 3180
rect 9340 2660 9500 2700
rect 8080 2560 8240 2600
rect 5880 2230 5920 2390
rect 10390 2230 10430 2390
rect 8080 2110 8240 2150
rect 6110 2010 6270 2050
rect 5330 1680 5370 1840
rect 7010 1680 7050 1840
rect 6110 1470 6270 1510
rect 8080 2010 8240 2050
rect 7120 1680 7160 1840
rect 9160 1680 9200 1840
rect 8080 1470 8240 1510
rect 10050 2010 10210 2050
rect 9270 1680 9310 1840
rect 10950 1680 10990 1840
rect 10050 1470 10210 1510
<< nsubdiffcont >>
rect 5840 7110 6000 7150
rect 5240 6780 5280 6940
rect 6560 6780 6600 6940
rect 5840 6570 6000 6610
rect 8080 7110 8240 7150
rect 6940 6780 6980 6940
rect 9340 6780 9380 6940
rect 8080 6570 8240 6610
rect 10320 7110 10480 7150
rect 9720 6780 9760 6940
rect 11040 6780 11080 6940
rect 10320 6570 10480 6610
rect 8080 6180 8240 6220
rect 5610 5980 5770 6020
rect 5330 5650 5370 5810
rect 6010 5650 6050 5810
rect 5610 5440 5770 5480
rect 6400 5650 6440 5810
rect 9880 5650 9920 5810
rect 10610 5980 10910 6020
rect 10260 5650 10300 5810
rect 11220 5650 11260 5810
rect 10610 5440 10910 5480
rect 8080 5230 8240 5270
rect 6560 4800 6720 4840
rect 5300 4470 5340 4630
rect 7940 4470 7980 4630
rect 6560 4260 6720 4300
rect 9600 4800 9760 4840
rect 8340 4470 8380 4630
rect 10980 4470 11020 4630
rect 9600 4260 9760 4300
<< poly >>
rect 5340 7050 5420 7070
rect 5340 7010 5360 7050
rect 5400 7020 5420 7050
rect 5880 7050 5960 7070
rect 5400 7010 5520 7020
rect 5880 7010 5900 7050
rect 5940 7010 5960 7050
rect 6420 7050 6500 7070
rect 6420 7020 6440 7050
rect 6320 7010 6440 7020
rect 6480 7010 6500 7050
rect 5340 6990 5520 7010
rect 5420 6960 5520 6990
rect 5600 6980 6240 7010
rect 5600 6960 5700 6980
rect 5780 6960 5880 6980
rect 5960 6960 6060 6980
rect 6140 6960 6240 6980
rect 6320 6990 6500 7010
rect 6320 6960 6420 6990
rect 5420 6730 5520 6760
rect 5600 6730 5700 6760
rect 5780 6730 5880 6760
rect 5960 6730 6060 6760
rect 6140 6730 6240 6760
rect 6320 6730 6420 6760
rect 7040 7050 7120 7070
rect 7040 7010 7060 7050
rect 7100 7020 7120 7050
rect 7940 7050 8020 7070
rect 7100 7010 7220 7020
rect 7940 7010 7960 7050
rect 8000 7010 8020 7050
rect 8300 7050 8380 7070
rect 8300 7010 8320 7050
rect 8360 7010 8380 7050
rect 9200 7050 9280 7070
rect 9200 7020 9220 7050
rect 9100 7010 9220 7020
rect 9260 7010 9280 7050
rect 7040 6990 7220 7010
rect 7120 6960 7220 6990
rect 7300 6980 9020 7010
rect 7300 6960 7400 6980
rect 7480 6960 7580 6980
rect 7660 6960 7760 6980
rect 7840 6960 7940 6980
rect 8020 6960 8120 6980
rect 8200 6960 8300 6980
rect 8380 6960 8480 6980
rect 8560 6960 8660 6980
rect 8740 6960 8840 6980
rect 8920 6960 9020 6980
rect 9100 6990 9280 7010
rect 9100 6960 9200 6990
rect 7120 6730 7220 6760
rect 7300 6730 7400 6760
rect 7480 6730 7580 6760
rect 7660 6730 7760 6760
rect 7840 6730 7940 6760
rect 8020 6730 8120 6760
rect 8200 6730 8300 6760
rect 8380 6730 8480 6760
rect 8560 6730 8660 6760
rect 8740 6730 8840 6760
rect 8920 6730 9020 6760
rect 9100 6730 9200 6760
rect 9820 7050 9900 7070
rect 9820 7010 9840 7050
rect 9880 7020 9900 7050
rect 10360 7050 10440 7070
rect 9880 7010 10000 7020
rect 10360 7010 10380 7050
rect 10420 7010 10440 7050
rect 10900 7050 10980 7070
rect 10900 7020 10920 7050
rect 10800 7010 10920 7020
rect 10960 7010 10980 7050
rect 9820 6990 10000 7010
rect 9900 6960 10000 6990
rect 10080 6980 10720 7010
rect 10080 6960 10180 6980
rect 10260 6960 10360 6980
rect 10440 6960 10540 6980
rect 10620 6960 10720 6980
rect 10800 6990 10980 7010
rect 10800 6960 10900 6990
rect 9900 6730 10000 6760
rect 10080 6730 10180 6760
rect 10260 6730 10360 6760
rect 10440 6730 10540 6760
rect 10620 6730 10720 6760
rect 10800 6730 10900 6760
rect 5440 5920 5500 5940
rect 5440 5880 5450 5920
rect 5490 5880 5500 5920
rect 5880 5920 5940 5940
rect 5880 5880 5890 5920
rect 5930 5880 5940 5920
rect 5440 5850 5540 5880
rect 5510 5830 5540 5850
rect 5620 5830 5650 5860
rect 5730 5830 5760 5860
rect 5840 5850 5940 5880
rect 5840 5830 5870 5850
rect 5510 5600 5540 5630
rect 5620 5610 5650 5630
rect 5730 5610 5760 5630
rect 5620 5580 5760 5610
rect 5840 5600 5870 5630
rect 5650 5540 5670 5580
rect 5710 5540 5730 5580
rect 5650 5520 5730 5540
rect 6500 6120 6580 6140
rect 6500 6080 6520 6120
rect 6560 6090 6580 6120
rect 9740 6120 9820 6140
rect 9740 6090 9760 6120
rect 6560 6080 6680 6090
rect 6500 6060 6680 6080
rect 9640 6080 9760 6090
rect 9800 6080 9820 6120
rect 9640 6060 9820 6080
rect 6580 6030 6680 6060
rect 6760 6030 6860 6060
rect 6940 6030 7040 6060
rect 7120 6030 7220 6060
rect 7300 6030 7400 6060
rect 7480 6030 7580 6060
rect 7660 6030 7760 6060
rect 7840 6030 7940 6060
rect 8020 6030 8120 6060
rect 8200 6030 8300 6060
rect 8380 6030 8480 6060
rect 8560 6030 8660 6060
rect 8740 6030 8840 6060
rect 8920 6030 9020 6060
rect 9100 6030 9200 6060
rect 9280 6030 9380 6060
rect 9460 6030 9560 6060
rect 9640 6030 9740 6060
rect 6580 5400 6680 5430
rect 6760 5410 6860 5430
rect 6940 5410 7040 5430
rect 7120 5410 7220 5430
rect 7300 5410 7400 5430
rect 7480 5410 7580 5430
rect 7660 5410 7760 5430
rect 7840 5410 7940 5430
rect 8020 5410 8120 5430
rect 8200 5410 8300 5430
rect 8380 5410 8480 5430
rect 8560 5410 8660 5430
rect 8740 5410 8840 5430
rect 8920 5410 9020 5430
rect 9100 5410 9200 5430
rect 9280 5410 9380 5430
rect 9460 5410 9560 5430
rect 6760 5380 9560 5410
rect 9640 5400 9740 5430
rect 7940 5340 7960 5380
rect 8000 5340 8020 5380
rect 7940 5320 8020 5340
rect 9380 5340 9400 5380
rect 9440 5340 9460 5380
rect 9380 5320 9460 5340
rect 10370 5920 10430 5940
rect 10370 5880 10380 5920
rect 10420 5890 10430 5920
rect 11090 5920 11150 5940
rect 11090 5890 11100 5920
rect 10420 5880 10540 5890
rect 10370 5860 10540 5880
rect 10980 5880 11100 5890
rect 11140 5880 11150 5920
rect 10980 5860 11150 5880
rect 10440 5830 10540 5860
rect 10620 5830 10720 5860
rect 10800 5830 10900 5860
rect 10980 5830 11080 5860
rect 10440 5600 10540 5630
rect 10620 5610 10720 5630
rect 10800 5610 10900 5630
rect 10620 5580 10900 5610
rect 10980 5600 11080 5630
rect 10720 5540 10740 5580
rect 10780 5540 10800 5580
rect 10720 5520 10800 5540
rect 5480 4650 5520 4680
rect 5600 4650 5640 4680
rect 5720 4650 5760 4680
rect 5840 4650 5880 4680
rect 5960 4650 6000 4680
rect 6080 4650 6120 4680
rect 6200 4650 6240 4680
rect 6320 4650 6360 4680
rect 6440 4650 6480 4680
rect 6560 4650 6600 4680
rect 6680 4650 6720 4680
rect 6800 4650 6840 4680
rect 6920 4650 6960 4680
rect 7040 4650 7080 4680
rect 7160 4650 7200 4680
rect 7280 4650 7320 4680
rect 7400 4650 7440 4680
rect 7520 4650 7560 4680
rect 7640 4650 7680 4680
rect 7760 4650 7800 4680
rect 5480 4430 5520 4450
rect 5410 4400 5520 4430
rect 5600 4420 5640 4450
rect 5720 4430 5760 4450
rect 5840 4430 5880 4450
rect 5960 4430 6000 4450
rect 6080 4430 6120 4450
rect 5580 4400 5660 4420
rect 5720 4400 6120 4430
rect 6200 4430 6240 4450
rect 6320 4430 6360 4450
rect 6200 4400 6360 4430
rect 6440 4430 6480 4450
rect 6560 4430 6600 4450
rect 6680 4430 6720 4450
rect 6800 4430 6840 4450
rect 6440 4400 6840 4430
rect 6920 4430 6960 4450
rect 7040 4430 7080 4450
rect 6920 4400 7080 4430
rect 7160 4430 7200 4450
rect 7280 4430 7320 4450
rect 7400 4430 7440 4450
rect 7520 4430 7560 4450
rect 7160 4400 7560 4430
rect 7640 4420 7680 4450
rect 7760 4430 7800 4450
rect 7630 4400 7690 4420
rect 7760 4400 7870 4430
rect 5410 4360 5420 4400
rect 5460 4360 5470 4400
rect 5410 4340 5470 4360
rect 5580 4360 5600 4400
rect 5640 4360 5660 4400
rect 5580 4340 5660 4360
rect 5760 4360 5780 4400
rect 5820 4360 5840 4400
rect 5760 4340 5840 4360
rect 6240 4360 6260 4400
rect 6300 4360 6320 4400
rect 6240 4340 6320 4360
rect 6480 4360 6500 4400
rect 6540 4360 6560 4400
rect 6480 4340 6560 4360
rect 6960 4360 6980 4400
rect 7020 4360 7040 4400
rect 6960 4340 7040 4360
rect 7200 4360 7220 4400
rect 7260 4360 7280 4400
rect 7200 4340 7280 4360
rect 7630 4360 7640 4400
rect 7680 4360 7690 4400
rect 7630 4340 7690 4360
rect 7810 4360 7820 4400
rect 7860 4360 7870 4400
rect 7810 4340 7870 4360
rect 8520 4650 8560 4680
rect 8640 4650 8680 4680
rect 8760 4650 8800 4680
rect 8880 4650 8920 4680
rect 9000 4650 9040 4680
rect 9120 4650 9160 4680
rect 9240 4650 9280 4680
rect 9360 4650 9400 4680
rect 9480 4650 9520 4680
rect 9600 4650 9640 4680
rect 9720 4650 9760 4680
rect 9840 4650 9880 4680
rect 9960 4650 10000 4680
rect 10080 4650 10120 4680
rect 10200 4650 10240 4680
rect 10320 4650 10360 4680
rect 10440 4650 10480 4680
rect 10560 4650 10600 4680
rect 10680 4650 10720 4680
rect 10800 4650 10840 4680
rect 8520 4430 8560 4450
rect 8450 4400 8560 4430
rect 8640 4420 8680 4450
rect 8760 4430 8800 4450
rect 8880 4430 8920 4450
rect 9000 4430 9040 4450
rect 9120 4430 9160 4450
rect 8630 4400 8690 4420
rect 8760 4400 9160 4430
rect 9240 4430 9280 4450
rect 9360 4430 9400 4450
rect 9240 4400 9400 4430
rect 9480 4430 9520 4450
rect 9600 4430 9640 4450
rect 9720 4430 9760 4450
rect 9840 4430 9880 4450
rect 9480 4400 9880 4430
rect 9960 4430 10000 4450
rect 10080 4430 10120 4450
rect 9960 4400 10120 4430
rect 10200 4430 10240 4450
rect 10320 4430 10360 4450
rect 10440 4430 10480 4450
rect 10560 4430 10600 4450
rect 10200 4400 10600 4430
rect 10680 4420 10720 4450
rect 10800 4430 10840 4450
rect 10660 4400 10740 4420
rect 10800 4400 10910 4430
rect 8450 4360 8460 4400
rect 8500 4360 8510 4400
rect 8450 4340 8510 4360
rect 8630 4360 8640 4400
rect 8680 4360 8690 4400
rect 8630 4340 8690 4360
rect 9040 4360 9060 4400
rect 9100 4360 9120 4400
rect 9040 4340 9120 4360
rect 9280 4360 9300 4400
rect 9340 4360 9360 4400
rect 9280 4340 9360 4360
rect 9760 4360 9780 4400
rect 9820 4360 9840 4400
rect 9760 4340 9840 4360
rect 10000 4360 10020 4400
rect 10060 4360 10080 4400
rect 10000 4340 10080 4360
rect 10480 4360 10500 4400
rect 10540 4360 10560 4400
rect 10480 4340 10560 4360
rect 10660 4360 10680 4400
rect 10720 4360 10740 4400
rect 10660 4340 10740 4360
rect 10850 4360 10860 4400
rect 10900 4360 10910 4400
rect 10850 4340 10910 4360
rect 6380 4080 6460 4100
rect 6380 4040 6400 4080
rect 6440 4040 6460 4080
rect 6380 4010 6460 4040
rect 6380 3980 7460 4010
rect 6340 3900 6380 3930
rect 6460 3900 6500 3980
rect 6580 3900 6620 3980
rect 6700 3900 6740 3930
rect 6820 3900 6860 3930
rect 6940 3900 6980 3980
rect 7060 3900 7100 3980
rect 7180 3900 7220 3930
rect 7300 3900 7340 3930
rect 7420 3900 7460 3980
rect 6340 3770 6380 3800
rect 6460 3770 6500 3800
rect 6580 3770 6620 3800
rect 6260 3750 6380 3770
rect 6260 3710 6280 3750
rect 6320 3720 6380 3750
rect 6700 3720 6740 3800
rect 6820 3720 6860 3800
rect 6940 3770 6980 3800
rect 7060 3770 7100 3800
rect 7180 3720 7220 3800
rect 7300 3720 7340 3800
rect 7420 3770 7460 3800
rect 6320 3710 7340 3720
rect 6260 3690 7340 3710
rect 9860 4080 9940 4100
rect 9860 4040 9880 4080
rect 9920 4040 9940 4080
rect 9860 4010 9940 4040
rect 8860 3980 9940 4010
rect 8860 3900 8900 3980
rect 8980 3900 9020 3930
rect 9100 3900 9140 3930
rect 9220 3900 9260 3980
rect 9340 3900 9380 3980
rect 9460 3900 9500 3930
rect 9580 3900 9620 3930
rect 9700 3900 9740 3980
rect 9820 3900 9860 3980
rect 9940 3900 9980 3930
rect 8860 3770 8900 3800
rect 8980 3720 9020 3800
rect 9100 3720 9140 3800
rect 9220 3770 9260 3800
rect 9340 3770 9380 3800
rect 9460 3720 9500 3800
rect 9580 3720 9620 3800
rect 9700 3770 9740 3800
rect 9820 3770 9860 3800
rect 9940 3770 9980 3800
rect 9940 3750 10060 3770
rect 9940 3720 10000 3750
rect 8980 3710 10000 3720
rect 10040 3710 10060 3750
rect 8980 3690 10060 3710
rect 5960 3430 6040 3450
rect 5960 3390 5980 3430
rect 6020 3390 6040 3430
rect 5960 3380 6040 3390
rect 6200 3430 6280 3450
rect 6200 3390 6220 3430
rect 6260 3390 6280 3430
rect 6200 3380 6280 3390
rect 6440 3430 6520 3450
rect 6440 3390 6460 3430
rect 6500 3390 6520 3430
rect 6440 3380 6520 3390
rect 6680 3430 6760 3450
rect 6680 3390 6700 3430
rect 6740 3390 6760 3430
rect 6680 3380 6760 3390
rect 7160 3430 7240 3450
rect 7160 3390 7180 3430
rect 7220 3390 7240 3430
rect 7160 3380 7240 3390
rect 7400 3430 7480 3450
rect 7400 3390 7420 3430
rect 7460 3390 7480 3430
rect 7400 3380 7480 3390
rect 7640 3430 7720 3450
rect 7640 3390 7660 3430
rect 7700 3390 7720 3430
rect 7640 3380 7720 3390
rect 5860 3350 6860 3380
rect 6940 3350 7940 3380
rect 5860 2820 6860 2850
rect 6940 2820 7940 2850
rect 8600 3430 8680 3450
rect 8600 3390 8620 3430
rect 8660 3390 8680 3430
rect 8600 3380 8680 3390
rect 8840 3430 8920 3450
rect 8840 3390 8860 3430
rect 8900 3390 8920 3430
rect 8840 3380 8920 3390
rect 9080 3430 9160 3450
rect 9080 3390 9100 3430
rect 9140 3390 9160 3430
rect 9080 3380 9160 3390
rect 9560 3430 9640 3450
rect 9560 3390 9580 3430
rect 9620 3390 9640 3430
rect 9560 3380 9640 3390
rect 9800 3430 9880 3450
rect 9800 3390 9820 3430
rect 9860 3390 9880 3430
rect 9800 3380 9880 3390
rect 10040 3430 10120 3450
rect 10040 3390 10060 3430
rect 10100 3390 10120 3430
rect 10040 3380 10120 3390
rect 10280 3430 10360 3450
rect 10280 3390 10300 3430
rect 10340 3390 10360 3430
rect 10280 3380 10360 3390
rect 8380 3350 9380 3380
rect 9460 3350 10460 3380
rect 8380 2820 9380 2850
rect 9460 2820 10460 2850
rect 6200 2500 6280 2520
rect 6200 2460 6220 2500
rect 6260 2460 6280 2500
rect 6200 2440 6280 2460
rect 6360 2500 6440 2520
rect 6360 2460 6380 2500
rect 6420 2460 6440 2500
rect 6360 2440 6440 2460
rect 6520 2500 6600 2520
rect 6520 2460 6540 2500
rect 6580 2460 6600 2500
rect 6520 2440 6600 2460
rect 6680 2500 6760 2520
rect 6680 2460 6700 2500
rect 6740 2460 6760 2500
rect 6680 2440 6760 2460
rect 6840 2500 6920 2520
rect 6840 2460 6860 2500
rect 6900 2460 6920 2500
rect 6840 2440 6920 2460
rect 7000 2500 7080 2520
rect 7000 2460 7020 2500
rect 7060 2460 7080 2500
rect 7000 2440 7080 2460
rect 7160 2500 7240 2520
rect 7160 2460 7180 2500
rect 7220 2460 7240 2500
rect 7160 2440 7240 2460
rect 7320 2500 7400 2520
rect 7320 2460 7340 2500
rect 7380 2460 7400 2500
rect 7320 2440 7400 2460
rect 7480 2500 7560 2520
rect 7480 2460 7500 2500
rect 7540 2460 7560 2500
rect 7480 2440 7560 2460
rect 7640 2500 7720 2520
rect 7640 2460 7660 2500
rect 7700 2460 7720 2500
rect 7640 2440 7720 2460
rect 7800 2500 7880 2520
rect 7800 2460 7820 2500
rect 7860 2460 7880 2500
rect 7800 2440 7880 2460
rect 7960 2500 8040 2520
rect 7960 2460 7980 2500
rect 8020 2460 8040 2500
rect 7960 2440 8040 2460
rect 8280 2500 8360 2520
rect 8280 2460 8300 2500
rect 8340 2460 8360 2500
rect 8280 2440 8360 2460
rect 8440 2500 8520 2520
rect 8440 2460 8460 2500
rect 8500 2460 8520 2500
rect 8440 2440 8520 2460
rect 8600 2500 8680 2520
rect 8600 2460 8620 2500
rect 8660 2460 8680 2500
rect 8600 2440 8680 2460
rect 8760 2500 8840 2520
rect 8760 2460 8780 2500
rect 8820 2460 8840 2500
rect 8760 2440 8840 2460
rect 8920 2500 9000 2520
rect 8920 2460 8940 2500
rect 8980 2460 9000 2500
rect 8920 2440 9000 2460
rect 9080 2500 9160 2520
rect 9080 2460 9100 2500
rect 9140 2460 9160 2500
rect 9080 2440 9160 2460
rect 9240 2500 9320 2520
rect 9240 2460 9260 2500
rect 9300 2460 9320 2500
rect 9240 2440 9320 2460
rect 9400 2500 9480 2520
rect 9400 2460 9420 2500
rect 9460 2460 9480 2500
rect 9400 2440 9480 2460
rect 9560 2500 9640 2520
rect 9560 2460 9580 2500
rect 9620 2460 9640 2500
rect 9560 2440 9640 2460
rect 9720 2500 9800 2520
rect 9720 2460 9740 2500
rect 9780 2460 9800 2500
rect 9720 2440 9800 2460
rect 9880 2500 9960 2520
rect 9880 2460 9900 2500
rect 9940 2460 9960 2500
rect 9880 2440 9960 2460
rect 10040 2500 10120 2520
rect 10040 2460 10060 2500
rect 10100 2460 10120 2500
rect 10040 2440 10120 2460
rect 6120 2410 8120 2440
rect 8200 2410 10200 2440
rect 6120 2180 8120 2210
rect 8200 2180 10200 2210
rect 6330 1950 6410 1970
rect 6330 1910 6350 1950
rect 6390 1910 6410 1950
rect 5510 1860 5610 1890
rect 5690 1880 6690 1910
rect 5690 1860 5790 1880
rect 5870 1860 5970 1880
rect 6050 1860 6150 1880
rect 6230 1860 6330 1880
rect 6410 1860 6510 1880
rect 6590 1860 6690 1880
rect 6770 1860 6870 1890
rect 5510 1640 5610 1660
rect 5440 1610 5610 1640
rect 5690 1630 5790 1660
rect 5870 1630 5970 1660
rect 6050 1630 6150 1660
rect 6230 1630 6330 1660
rect 6410 1630 6510 1660
rect 6590 1630 6690 1660
rect 6770 1640 6870 1660
rect 6770 1610 6940 1640
rect 5440 1570 5450 1610
rect 5490 1570 5500 1610
rect 5440 1550 5500 1570
rect 6880 1570 6890 1610
rect 6930 1570 6940 1610
rect 6880 1550 6940 1570
rect 8120 1950 8200 1970
rect 8120 1910 8140 1950
rect 8180 1910 8200 1950
rect 7300 1860 7400 1890
rect 7480 1880 8840 1910
rect 7480 1860 7580 1880
rect 7660 1860 7760 1880
rect 7840 1860 7940 1880
rect 8020 1860 8120 1880
rect 8200 1860 8300 1880
rect 8380 1860 8480 1880
rect 8560 1860 8660 1880
rect 8740 1860 8840 1880
rect 8920 1860 9020 1890
rect 7300 1640 7400 1660
rect 7230 1610 7400 1640
rect 7480 1630 7580 1660
rect 7660 1630 7760 1660
rect 7840 1630 7940 1660
rect 8020 1630 8120 1660
rect 8200 1630 8300 1660
rect 8380 1630 8480 1660
rect 8560 1630 8660 1660
rect 8740 1630 8840 1660
rect 8920 1640 9020 1660
rect 7490 1610 7570 1630
rect 8920 1610 9090 1640
rect 7230 1570 7240 1610
rect 7280 1570 7290 1610
rect 7230 1550 7290 1570
rect 7490 1570 7510 1610
rect 7550 1570 7570 1610
rect 7490 1550 7570 1570
rect 9030 1570 9040 1610
rect 9080 1570 9090 1610
rect 9030 1550 9090 1570
rect 9910 1950 9990 1970
rect 9910 1910 9930 1950
rect 9970 1910 9990 1950
rect 9450 1860 9550 1890
rect 9630 1880 10630 1910
rect 9630 1860 9730 1880
rect 9810 1860 9910 1880
rect 9990 1860 10090 1880
rect 10170 1860 10270 1880
rect 10350 1860 10450 1880
rect 10530 1860 10630 1880
rect 10710 1860 10810 1890
rect 9450 1640 9550 1660
rect 9380 1610 9550 1640
rect 9630 1630 9730 1660
rect 9810 1630 9910 1660
rect 9990 1630 10090 1660
rect 10170 1630 10270 1660
rect 10350 1630 10450 1660
rect 10530 1630 10630 1660
rect 10710 1640 10810 1660
rect 10710 1610 10880 1640
rect 9380 1570 9390 1610
rect 9430 1570 9440 1610
rect 9380 1550 9440 1570
rect 10820 1570 10830 1610
rect 10870 1570 10880 1610
rect 10820 1550 10880 1570
<< polycont >>
rect 5360 7010 5400 7050
rect 5900 7010 5940 7050
rect 6440 7010 6480 7050
rect 7060 7010 7100 7050
rect 7960 7010 8000 7050
rect 8320 7010 8360 7050
rect 9220 7010 9260 7050
rect 9840 7010 9880 7050
rect 10380 7010 10420 7050
rect 10920 7010 10960 7050
rect 5450 5880 5490 5920
rect 5890 5880 5930 5920
rect 5670 5540 5710 5580
rect 6520 6080 6560 6120
rect 9760 6080 9800 6120
rect 7960 5340 8000 5380
rect 9400 5340 9440 5380
rect 10380 5880 10420 5920
rect 11100 5880 11140 5920
rect 10740 5540 10780 5580
rect 5420 4360 5460 4400
rect 5600 4360 5640 4400
rect 5780 4360 5820 4400
rect 6260 4360 6300 4400
rect 6500 4360 6540 4400
rect 6980 4360 7020 4400
rect 7220 4360 7260 4400
rect 7640 4360 7680 4400
rect 7820 4360 7860 4400
rect 8460 4360 8500 4400
rect 8640 4360 8680 4400
rect 9060 4360 9100 4400
rect 9300 4360 9340 4400
rect 9780 4360 9820 4400
rect 10020 4360 10060 4400
rect 10500 4360 10540 4400
rect 10680 4360 10720 4400
rect 10860 4360 10900 4400
rect 6400 4040 6440 4080
rect 6280 3710 6320 3750
rect 9880 4040 9920 4080
rect 10000 3710 10040 3750
rect 5980 3390 6020 3430
rect 6220 3390 6260 3430
rect 6460 3390 6500 3430
rect 6700 3390 6740 3430
rect 7180 3390 7220 3430
rect 7420 3390 7460 3430
rect 7660 3390 7700 3430
rect 8620 3390 8660 3430
rect 8860 3390 8900 3430
rect 9100 3390 9140 3430
rect 9580 3390 9620 3430
rect 9820 3390 9860 3430
rect 10060 3390 10100 3430
rect 10300 3390 10340 3430
rect 6220 2460 6260 2500
rect 6380 2460 6420 2500
rect 6540 2460 6580 2500
rect 6700 2460 6740 2500
rect 6860 2460 6900 2500
rect 7020 2460 7060 2500
rect 7180 2460 7220 2500
rect 7340 2460 7380 2500
rect 7500 2460 7540 2500
rect 7660 2460 7700 2500
rect 7820 2460 7860 2500
rect 7980 2460 8020 2500
rect 8300 2460 8340 2500
rect 8460 2460 8500 2500
rect 8620 2460 8660 2500
rect 8780 2460 8820 2500
rect 8940 2460 8980 2500
rect 9100 2460 9140 2500
rect 9260 2460 9300 2500
rect 9420 2460 9460 2500
rect 9580 2460 9620 2500
rect 9740 2460 9780 2500
rect 9900 2460 9940 2500
rect 10060 2460 10100 2500
rect 6350 1910 6390 1950
rect 5450 1570 5490 1610
rect 6890 1570 6930 1610
rect 8140 1910 8180 1950
rect 7240 1570 7280 1610
rect 7510 1570 7550 1610
rect 9040 1570 9080 1610
rect 9930 1910 9970 1950
rect 9390 1570 9430 1610
rect 10830 1570 10870 1610
<< xpolycontact >>
rect 222 7110 662 7180
rect 1890 7110 2330 7180
rect 222 6990 662 7060
rect 1890 6990 2330 7060
rect 222 6580 662 6650
rect 1830 6580 2270 6650
rect 222 6460 662 6530
rect 1830 6460 2270 6530
rect 2792 6840 3232 6910
rect 4400 6840 4840 6910
rect 2792 6720 3232 6790
rect 4400 6720 4840 6790
rect 2792 6600 3232 6670
rect 4400 6600 4840 6670
rect 612 6050 1050 6120
rect 1428 6050 1868 6120
rect 2792 6480 3232 6550
rect 4400 6480 4840 6550
rect 2792 6360 3232 6430
rect 4400 6360 4840 6430
rect 2792 6240 3232 6310
rect 4400 6240 4840 6310
rect 612 5630 1050 5700
rect 1428 5630 1868 5700
rect 3122 5830 3562 5900
rect 3990 5830 4430 5900
<< ppolyres >>
rect 1050 6050 1428 6120
rect 1050 5630 1428 5700
<< xpolyres >>
rect 662 7110 1890 7180
rect 662 6990 1890 7060
rect 662 6580 1830 6650
rect 662 6460 1830 6530
rect 3232 6840 4400 6910
rect 3232 6720 4400 6790
rect 3232 6600 4400 6670
rect 3232 6480 4400 6550
rect 3232 6360 4400 6430
rect 3232 6240 4400 6310
rect 3562 5830 3990 5900
<< locali >>
rect 8890 7630 8950 7690
rect 1890 7530 1950 7590
rect 3290 7530 3350 7590
rect 10290 7530 10350 7590
rect 5390 7420 5450 7480
rect 6790 7420 6850 7480
rect 50 7280 1180 7320
rect 1340 7280 2470 7320
rect 50 7160 90 7280
rect 132 7170 222 7180
rect 132 7120 152 7170
rect 202 7120 222 7170
rect 132 7110 222 7120
rect 2260 7060 2330 7110
rect 50 6890 90 7000
rect 132 7050 222 7060
rect 132 7000 152 7050
rect 202 7000 222 7050
rect 132 6990 222 7000
rect 2430 7160 2470 7280
rect 5240 7110 5840 7150
rect 6000 7110 6600 7150
rect 2430 6890 2470 7000
rect 50 6850 1180 6890
rect 1340 6850 2470 6890
rect 2620 7010 3690 7050
rect 3850 7010 5010 7050
rect 1230 6790 1270 6850
rect 50 6750 1150 6790
rect 1310 6750 2410 6790
rect 50 6630 90 6750
rect 132 6640 222 6650
rect 132 6590 152 6640
rect 202 6590 222 6640
rect 132 6580 222 6590
rect 2200 6530 2270 6580
rect 50 6360 90 6470
rect 132 6520 222 6530
rect 132 6470 152 6520
rect 202 6470 222 6520
rect 132 6460 222 6470
rect 2370 6630 2410 6750
rect 2620 6650 2660 7010
rect 2702 6900 2792 6910
rect 2702 6850 2722 6900
rect 2772 6850 2792 6900
rect 2702 6840 2792 6850
rect 4840 6840 4920 6910
rect 2702 6780 2792 6790
rect 2702 6730 2722 6780
rect 2772 6730 2792 6780
rect 2702 6720 2792 6730
rect 4770 6670 4840 6720
rect 2410 6570 2450 6590
rect 2430 6530 2450 6570
rect 2410 6510 2450 6530
rect 2580 6570 2620 6590
rect 2580 6530 2600 6570
rect 2580 6510 2620 6530
rect 1190 6380 1270 6400
rect 1190 6360 1210 6380
rect 1250 6360 1270 6380
rect 2370 6360 2410 6470
rect 50 6320 1150 6360
rect 1310 6320 2410 6360
rect 1210 6260 1250 6320
rect 440 6220 1150 6260
rect 1310 6220 2040 6260
rect 440 6160 480 6220
rect 2000 6160 2040 6220
rect 522 6110 612 6120
rect 522 6060 542 6110
rect 592 6060 612 6110
rect 522 6050 612 6060
rect 1868 6110 1958 6120
rect 1868 6060 1888 6110
rect 1938 6060 1958 6110
rect 1868 6050 1958 6060
rect 440 5940 480 6000
rect 2620 6140 2660 6490
rect 2712 6600 2792 6670
rect 2712 6310 2752 6600
rect 4880 6550 4920 6840
rect 4840 6480 4920 6550
rect 4970 6650 5010 7010
rect 5240 6940 5280 7110
rect 5360 7070 5400 7110
rect 6440 7070 6480 7110
rect 5340 7050 5420 7070
rect 5340 7010 5360 7050
rect 5400 7010 5420 7050
rect 5340 6990 5420 7010
rect 5700 7050 5780 7070
rect 5700 7010 5720 7050
rect 5760 7010 5780 7050
rect 5700 6990 5780 7010
rect 5880 7050 5960 7070
rect 5880 7010 5900 7050
rect 5940 7010 5960 7050
rect 5880 6990 5960 7010
rect 6060 7050 6140 7070
rect 6060 7010 6080 7050
rect 6120 7010 6140 7050
rect 6060 6990 6140 7010
rect 6240 7050 6320 7070
rect 6240 7010 6260 7050
rect 6300 7010 6320 7050
rect 6240 6990 6320 7010
rect 6420 7050 6500 7070
rect 6420 7010 6440 7050
rect 6480 7010 6500 7050
rect 6420 6990 6500 7010
rect 5360 6950 5400 6990
rect 5720 6950 5760 6990
rect 6080 6950 6120 6990
rect 6260 6950 6300 6990
rect 6440 6950 6480 6990
rect 5240 6610 5280 6780
rect 5350 6930 5410 6950
rect 5350 6786 5360 6930
rect 5400 6786 5410 6930
rect 5350 6770 5410 6786
rect 5530 6930 5590 6950
rect 5530 6786 5540 6930
rect 5580 6786 5590 6930
rect 5530 6770 5590 6786
rect 5710 6930 5770 6950
rect 5710 6786 5720 6930
rect 5760 6786 5770 6930
rect 5710 6770 5770 6786
rect 5890 6930 5950 6950
rect 5890 6786 5900 6930
rect 5940 6786 5950 6930
rect 5890 6770 5950 6786
rect 6070 6930 6130 6950
rect 6070 6786 6080 6930
rect 6120 6786 6130 6930
rect 6070 6770 6130 6786
rect 6250 6930 6310 6950
rect 6250 6786 6260 6930
rect 6300 6786 6310 6930
rect 6250 6770 6310 6786
rect 6430 6930 6490 6950
rect 6430 6786 6440 6930
rect 6480 6786 6490 6930
rect 6430 6770 6490 6786
rect 6560 6940 6600 7110
rect 5540 6730 5580 6770
rect 5900 6730 5940 6770
rect 6260 6730 6300 6770
rect 5520 6710 5600 6730
rect 5520 6670 5540 6710
rect 5580 6670 5600 6710
rect 5520 6650 5600 6670
rect 5880 6710 5960 6730
rect 5880 6670 5900 6710
rect 5940 6670 5960 6710
rect 5880 6650 5960 6670
rect 6240 6710 6320 6730
rect 6240 6670 6260 6710
rect 6300 6670 6320 6710
rect 6240 6650 6320 6670
rect 6560 6610 6600 6780
rect 5240 6570 5840 6610
rect 6000 6570 6600 6610
rect 6940 7110 8080 7150
rect 8240 7110 9380 7150
rect 6940 6940 6980 7110
rect 7060 7070 7100 7110
rect 9220 7070 9260 7110
rect 7040 7050 7120 7070
rect 7040 7010 7060 7050
rect 7100 7010 7120 7050
rect 7040 6990 7120 7010
rect 7400 7050 7480 7070
rect 7400 7010 7420 7050
rect 7460 7010 7480 7050
rect 7400 6990 7480 7010
rect 7760 7050 7840 7070
rect 7760 7010 7780 7050
rect 7820 7010 7840 7050
rect 7760 6990 7840 7010
rect 7940 7050 8020 7070
rect 7940 7010 7960 7050
rect 8000 7010 8020 7050
rect 7940 6990 8020 7010
rect 8120 7050 8200 7070
rect 8120 7010 8140 7050
rect 8180 7010 8200 7050
rect 8120 6990 8200 7010
rect 8300 7050 8380 7070
rect 8300 7010 8320 7050
rect 8360 7010 8380 7050
rect 8300 6990 8380 7010
rect 8480 7050 8560 7070
rect 8480 7010 8500 7050
rect 8540 7010 8560 7050
rect 8480 6990 8560 7010
rect 8840 7050 8920 7070
rect 8840 7010 8860 7050
rect 8900 7010 8920 7050
rect 8840 6990 8920 7010
rect 9020 7050 9100 7070
rect 9020 7010 9040 7050
rect 9080 7010 9100 7050
rect 9020 6990 9100 7010
rect 9200 7050 9280 7070
rect 9200 7010 9220 7050
rect 9260 7010 9280 7050
rect 9200 6990 9280 7010
rect 7060 6950 7100 6990
rect 7420 6950 7460 6990
rect 7780 6950 7820 6990
rect 8140 6950 8180 6990
rect 8500 6950 8540 6990
rect 8860 6950 8900 6990
rect 9040 6950 9080 6990
rect 9220 6950 9260 6990
rect 6940 6610 6980 6780
rect 7050 6930 7110 6950
rect 7050 6890 7060 6930
rect 7100 6890 7110 6930
rect 7050 6830 7110 6890
rect 7050 6790 7060 6830
rect 7100 6790 7110 6830
rect 7050 6770 7110 6790
rect 7230 6930 7290 6950
rect 7230 6890 7240 6930
rect 7280 6890 7290 6930
rect 7230 6830 7290 6890
rect 7230 6790 7240 6830
rect 7280 6790 7290 6830
rect 7230 6770 7290 6790
rect 7410 6930 7470 6950
rect 7410 6890 7420 6930
rect 7460 6890 7470 6930
rect 7410 6830 7470 6890
rect 7410 6790 7420 6830
rect 7460 6790 7470 6830
rect 7410 6770 7470 6790
rect 7590 6930 7650 6950
rect 7590 6890 7600 6930
rect 7640 6890 7650 6930
rect 7590 6830 7650 6890
rect 7590 6790 7600 6830
rect 7640 6790 7650 6830
rect 7590 6770 7650 6790
rect 7770 6930 7830 6950
rect 7770 6890 7780 6930
rect 7820 6890 7830 6930
rect 7770 6830 7830 6890
rect 7770 6790 7780 6830
rect 7820 6790 7830 6830
rect 7770 6770 7830 6790
rect 7950 6930 8010 6950
rect 7950 6890 7960 6930
rect 8000 6890 8010 6930
rect 7950 6830 8010 6890
rect 7950 6790 7960 6830
rect 8000 6790 8010 6830
rect 7950 6770 8010 6790
rect 8130 6930 8190 6950
rect 8130 6890 8140 6930
rect 8180 6890 8190 6930
rect 8130 6830 8190 6890
rect 8130 6790 8140 6830
rect 8180 6790 8190 6830
rect 8130 6770 8190 6790
rect 8310 6930 8370 6950
rect 8310 6890 8320 6930
rect 8360 6890 8370 6930
rect 8310 6830 8370 6890
rect 8310 6790 8320 6830
rect 8360 6790 8370 6830
rect 8310 6770 8370 6790
rect 8490 6930 8550 6950
rect 8490 6890 8500 6930
rect 8540 6890 8550 6930
rect 8490 6830 8550 6890
rect 8490 6790 8500 6830
rect 8540 6790 8550 6830
rect 8490 6770 8550 6790
rect 8670 6930 8730 6950
rect 8670 6890 8680 6930
rect 8720 6890 8730 6930
rect 8670 6830 8730 6890
rect 8670 6790 8680 6830
rect 8720 6790 8730 6830
rect 8670 6770 8730 6790
rect 8850 6930 8910 6950
rect 8850 6890 8860 6930
rect 8900 6890 8910 6930
rect 8850 6830 8910 6890
rect 8850 6790 8860 6830
rect 8900 6790 8910 6830
rect 8850 6770 8910 6790
rect 9030 6930 9090 6950
rect 9030 6890 9040 6930
rect 9080 6890 9090 6930
rect 9030 6830 9090 6890
rect 9030 6790 9040 6830
rect 9080 6790 9090 6830
rect 9030 6770 9090 6790
rect 9210 6930 9270 6950
rect 9210 6890 9220 6930
rect 9260 6890 9270 6930
rect 9210 6830 9270 6890
rect 9210 6790 9220 6830
rect 9260 6790 9270 6830
rect 9210 6770 9270 6790
rect 9340 6940 9380 7110
rect 7240 6730 7280 6770
rect 7600 6730 7640 6770
rect 7960 6730 8000 6770
rect 8320 6730 8360 6770
rect 8680 6730 8720 6770
rect 9040 6730 9080 6770
rect 7220 6710 7300 6730
rect 7220 6670 7240 6710
rect 7280 6670 7300 6710
rect 7220 6650 7300 6670
rect 7580 6710 7660 6730
rect 7580 6670 7600 6710
rect 7640 6670 7660 6710
rect 7580 6650 7660 6670
rect 7940 6710 8020 6730
rect 7940 6670 7960 6710
rect 8000 6670 8020 6710
rect 7940 6650 8020 6670
rect 8300 6710 8380 6730
rect 8300 6670 8320 6710
rect 8360 6670 8380 6710
rect 8300 6650 8380 6670
rect 8660 6710 8740 6730
rect 8660 6670 8680 6710
rect 8720 6670 8740 6710
rect 8660 6650 8740 6670
rect 9020 6710 9100 6730
rect 9020 6670 9040 6710
rect 9080 6670 9100 6710
rect 9020 6650 9100 6670
rect 9340 6610 9380 6780
rect 6940 6570 8080 6610
rect 8240 6570 9380 6610
rect 9720 7110 10320 7150
rect 10480 7110 11080 7150
rect 9720 6940 9760 7110
rect 9840 7070 9880 7110
rect 10920 7070 10960 7110
rect 9820 7050 9900 7070
rect 9820 7010 9840 7050
rect 9880 7010 9900 7050
rect 9820 6990 9900 7010
rect 10180 7050 10260 7070
rect 10180 7010 10200 7050
rect 10240 7010 10260 7050
rect 10180 6990 10260 7010
rect 10360 7050 10440 7070
rect 10360 7010 10380 7050
rect 10420 7010 10440 7050
rect 10360 6990 10440 7010
rect 10540 7050 10620 7070
rect 10540 7010 10560 7050
rect 10600 7010 10620 7050
rect 10540 6990 10620 7010
rect 10900 7050 10980 7070
rect 10900 7010 10920 7050
rect 10960 7010 10980 7050
rect 10900 6990 10980 7010
rect 9840 6950 9880 6990
rect 10200 6950 10240 6990
rect 10560 6950 10600 6990
rect 10920 6950 10960 6990
rect 9720 6610 9760 6780
rect 9830 6930 9890 6950
rect 9830 6790 9840 6930
rect 9880 6790 9890 6930
rect 9830 6770 9890 6790
rect 10010 6930 10070 6950
rect 10010 6790 10020 6930
rect 10060 6790 10070 6930
rect 10010 6770 10070 6790
rect 10190 6930 10250 6950
rect 10190 6790 10200 6930
rect 10240 6790 10250 6930
rect 10190 6770 10250 6790
rect 10370 6930 10430 6950
rect 10370 6790 10380 6930
rect 10420 6790 10430 6930
rect 10370 6770 10430 6790
rect 10550 6930 10610 6950
rect 10550 6790 10560 6930
rect 10600 6790 10610 6930
rect 10550 6770 10610 6790
rect 10730 6930 10790 6950
rect 10730 6790 10740 6930
rect 10780 6790 10790 6930
rect 10730 6770 10790 6790
rect 10910 6930 10970 6950
rect 10910 6790 10920 6930
rect 10960 6790 10970 6930
rect 10910 6770 10970 6790
rect 11040 6940 11080 7110
rect 10020 6730 10060 6770
rect 10380 6730 10420 6770
rect 10740 6730 10780 6770
rect 10000 6710 10080 6730
rect 10000 6670 10020 6710
rect 10060 6670 10080 6710
rect 10000 6650 10080 6670
rect 10360 6710 10440 6730
rect 10360 6670 10380 6710
rect 10420 6670 10440 6710
rect 10360 6650 10440 6670
rect 10720 6710 10800 6730
rect 10720 6670 10740 6710
rect 10780 6670 10800 6710
rect 10720 6650 10800 6670
rect 11040 6610 11080 6780
rect 9720 6570 10320 6610
rect 10480 6570 11080 6610
rect 2792 6430 2862 6480
rect 4840 6420 4930 6430
rect 4840 6370 4860 6420
rect 4910 6370 4930 6420
rect 4840 6360 4930 6370
rect 2712 6240 2792 6310
rect 4840 6300 4930 6320
rect 4840 6250 4860 6300
rect 4910 6250 4930 6300
rect 4840 6230 4930 6250
rect 4970 6140 5010 6490
rect 2620 6100 3690 6140
rect 3850 6100 5010 6140
rect 6400 6180 8080 6220
rect 8240 6180 9920 6220
rect 3750 6040 3790 6100
rect 5650 6040 5730 6060
rect 2000 5940 2040 6000
rect 440 5900 1150 5940
rect 1310 5900 2040 5940
rect 2950 6000 3690 6040
rect 3850 6000 4600 6040
rect 5650 6020 5670 6040
rect 5710 6020 5730 6040
rect 2950 5940 2990 6000
rect 1210 5840 1250 5900
rect 440 5800 1150 5840
rect 1310 5800 2040 5840
rect 440 5740 480 5800
rect 2000 5740 2040 5800
rect 522 5690 612 5700
rect 522 5640 542 5690
rect 592 5640 612 5690
rect 522 5630 612 5640
rect 1868 5690 1958 5700
rect 1868 5640 1888 5690
rect 1938 5640 1958 5690
rect 1868 5630 1958 5640
rect 440 5520 480 5580
rect 4560 5940 4600 6000
rect 3032 5890 3122 5900
rect 3032 5840 3052 5890
rect 3102 5840 3122 5890
rect 3032 5830 3122 5840
rect 4430 5890 4520 5900
rect 4430 5840 4450 5890
rect 4500 5840 4520 5890
rect 4430 5830 4520 5840
rect 2950 5730 2990 5780
rect 4560 5730 4600 5780
rect 2950 5690 3690 5730
rect 3850 5690 4600 5730
rect 5330 5980 5610 6020
rect 5770 5980 6050 6020
rect 5330 5810 5370 5980
rect 5450 5940 5490 5980
rect 5890 5940 5930 5980
rect 2000 5520 2040 5580
rect 440 5480 1150 5520
rect 1310 5480 2040 5520
rect 5330 5480 5370 5650
rect 5440 5920 5500 5940
rect 5440 5880 5450 5920
rect 5490 5880 5500 5920
rect 5440 5800 5500 5880
rect 5650 5920 5730 5940
rect 5650 5880 5670 5920
rect 5710 5880 5730 5920
rect 5650 5860 5730 5880
rect 5880 5920 5940 5940
rect 5880 5880 5890 5920
rect 5930 5880 5940 5920
rect 5670 5820 5710 5860
rect 5440 5760 5450 5800
rect 5490 5760 5500 5800
rect 5440 5700 5500 5760
rect 5440 5660 5450 5700
rect 5490 5660 5500 5700
rect 5440 5640 5500 5660
rect 5550 5800 5610 5820
rect 5550 5760 5560 5800
rect 5600 5760 5610 5800
rect 5550 5700 5610 5760
rect 5550 5660 5560 5700
rect 5600 5660 5610 5700
rect 5550 5640 5610 5660
rect 5660 5800 5720 5820
rect 5660 5760 5670 5800
rect 5710 5760 5720 5800
rect 5660 5700 5720 5760
rect 5660 5660 5670 5700
rect 5710 5660 5720 5700
rect 5660 5640 5720 5660
rect 5770 5800 5830 5820
rect 5770 5760 5780 5800
rect 5820 5760 5830 5800
rect 5770 5700 5830 5760
rect 5770 5660 5780 5700
rect 5820 5660 5830 5700
rect 5770 5640 5830 5660
rect 5880 5800 5940 5880
rect 5880 5760 5890 5800
rect 5930 5760 5940 5800
rect 5880 5700 5940 5760
rect 5880 5660 5890 5700
rect 5930 5660 5940 5700
rect 5880 5640 5940 5660
rect 6010 5810 6050 5980
rect 5560 5600 5600 5640
rect 5780 5600 5820 5640
rect 5520 5580 5600 5600
rect 5520 5540 5540 5580
rect 5580 5540 5600 5580
rect 5520 5520 5600 5540
rect 5650 5580 5730 5600
rect 5650 5540 5670 5580
rect 5710 5540 5730 5580
rect 5650 5520 5730 5540
rect 5780 5580 5860 5600
rect 5780 5540 5800 5580
rect 5840 5540 5860 5580
rect 5780 5520 5860 5540
rect 6010 5480 6050 5650
rect 5330 5440 5610 5480
rect 5770 5440 6050 5480
rect 6400 5810 6440 6180
rect 6520 6140 6560 6180
rect 9760 6140 9800 6180
rect 6500 6120 6580 6140
rect 6500 6080 6520 6120
rect 6560 6080 6580 6120
rect 6500 6060 6580 6080
rect 6860 6120 6940 6140
rect 6860 6080 6880 6120
rect 6920 6080 6940 6120
rect 6860 6060 6940 6080
rect 7220 6120 7300 6140
rect 7220 6080 7240 6120
rect 7280 6080 7300 6120
rect 7220 6060 7300 6080
rect 7580 6120 7660 6140
rect 7580 6080 7600 6120
rect 7640 6080 7660 6120
rect 7580 6060 7660 6080
rect 7940 6120 8020 6140
rect 7940 6080 7960 6120
rect 8000 6080 8020 6120
rect 7940 6060 8020 6080
rect 8300 6120 8380 6140
rect 8300 6080 8320 6120
rect 8360 6080 8380 6120
rect 8300 6060 8380 6080
rect 8660 6120 8740 6140
rect 8660 6080 8680 6120
rect 8720 6080 8740 6120
rect 8660 6060 8740 6080
rect 9020 6120 9100 6140
rect 9020 6080 9040 6120
rect 9080 6080 9100 6120
rect 9020 6060 9100 6080
rect 9380 6120 9460 6140
rect 9380 6080 9400 6120
rect 9440 6080 9460 6120
rect 9380 6060 9460 6080
rect 9740 6120 9820 6140
rect 9740 6080 9760 6120
rect 9800 6080 9820 6120
rect 9740 6060 9820 6080
rect 6520 6020 6560 6060
rect 6880 6020 6920 6060
rect 7240 6020 7280 6060
rect 7600 6020 7640 6060
rect 7960 6020 8000 6060
rect 8320 6020 8360 6060
rect 8680 6020 8720 6060
rect 9040 6020 9080 6060
rect 9400 6020 9440 6060
rect 9760 6020 9800 6060
rect 1300 4110 1550 5400
rect 2660 4110 2910 5400
rect 4020 4110 4270 5400
rect 6400 5270 6440 5650
rect 6510 6000 6570 6020
rect 6510 5960 6520 6000
rect 6560 5960 6570 6000
rect 6510 5900 6570 5960
rect 6510 5860 6520 5900
rect 6560 5860 6570 5900
rect 6510 5800 6570 5860
rect 6510 5760 6520 5800
rect 6560 5760 6570 5800
rect 6510 5700 6570 5760
rect 6510 5660 6520 5700
rect 6560 5660 6570 5700
rect 6510 5600 6570 5660
rect 6510 5560 6520 5600
rect 6560 5560 6570 5600
rect 6510 5500 6570 5560
rect 6510 5460 6520 5500
rect 6560 5460 6570 5500
rect 6510 5440 6570 5460
rect 6690 6000 6750 6020
rect 6690 5960 6700 6000
rect 6740 5960 6750 6000
rect 6690 5900 6750 5960
rect 6690 5860 6700 5900
rect 6740 5860 6750 5900
rect 6690 5800 6750 5860
rect 6690 5760 6700 5800
rect 6740 5760 6750 5800
rect 6690 5700 6750 5760
rect 6690 5660 6700 5700
rect 6740 5660 6750 5700
rect 6690 5600 6750 5660
rect 6690 5560 6700 5600
rect 6740 5560 6750 5600
rect 6690 5500 6750 5560
rect 6690 5460 6700 5500
rect 6740 5460 6750 5500
rect 6690 5440 6750 5460
rect 6870 6000 6930 6020
rect 6870 5960 6880 6000
rect 6920 5960 6930 6000
rect 6870 5900 6930 5960
rect 6870 5860 6880 5900
rect 6920 5860 6930 5900
rect 6870 5800 6930 5860
rect 6870 5760 6880 5800
rect 6920 5760 6930 5800
rect 6870 5700 6930 5760
rect 6870 5660 6880 5700
rect 6920 5660 6930 5700
rect 6870 5600 6930 5660
rect 6870 5560 6880 5600
rect 6920 5560 6930 5600
rect 6870 5500 6930 5560
rect 6870 5460 6880 5500
rect 6920 5460 6930 5500
rect 6870 5440 6930 5460
rect 7050 6000 7110 6020
rect 7050 5960 7060 6000
rect 7100 5960 7110 6000
rect 7050 5900 7110 5960
rect 7050 5860 7060 5900
rect 7100 5860 7110 5900
rect 7050 5800 7110 5860
rect 7050 5760 7060 5800
rect 7100 5760 7110 5800
rect 7050 5700 7110 5760
rect 7050 5660 7060 5700
rect 7100 5660 7110 5700
rect 7050 5600 7110 5660
rect 7050 5560 7060 5600
rect 7100 5560 7110 5600
rect 7050 5500 7110 5560
rect 7050 5460 7060 5500
rect 7100 5460 7110 5500
rect 7050 5440 7110 5460
rect 7230 6000 7290 6020
rect 7230 5960 7240 6000
rect 7280 5960 7290 6000
rect 7230 5900 7290 5960
rect 7230 5860 7240 5900
rect 7280 5860 7290 5900
rect 7230 5800 7290 5860
rect 7230 5760 7240 5800
rect 7280 5760 7290 5800
rect 7230 5700 7290 5760
rect 7230 5660 7240 5700
rect 7280 5660 7290 5700
rect 7230 5600 7290 5660
rect 7230 5560 7240 5600
rect 7280 5560 7290 5600
rect 7230 5500 7290 5560
rect 7230 5460 7240 5500
rect 7280 5460 7290 5500
rect 7230 5440 7290 5460
rect 7410 6000 7470 6020
rect 7410 5960 7420 6000
rect 7460 5960 7470 6000
rect 7410 5900 7470 5960
rect 7410 5860 7420 5900
rect 7460 5860 7470 5900
rect 7410 5800 7470 5860
rect 7410 5760 7420 5800
rect 7460 5760 7470 5800
rect 7410 5700 7470 5760
rect 7410 5660 7420 5700
rect 7460 5660 7470 5700
rect 7410 5600 7470 5660
rect 7410 5560 7420 5600
rect 7460 5560 7470 5600
rect 7410 5500 7470 5560
rect 7410 5460 7420 5500
rect 7460 5460 7470 5500
rect 7410 5440 7470 5460
rect 7590 6000 7650 6020
rect 7590 5960 7600 6000
rect 7640 5960 7650 6000
rect 7590 5900 7650 5960
rect 7590 5860 7600 5900
rect 7640 5860 7650 5900
rect 7590 5800 7650 5860
rect 7590 5760 7600 5800
rect 7640 5760 7650 5800
rect 7590 5700 7650 5760
rect 7590 5660 7600 5700
rect 7640 5660 7650 5700
rect 7590 5600 7650 5660
rect 7590 5560 7600 5600
rect 7640 5560 7650 5600
rect 7590 5500 7650 5560
rect 7590 5460 7600 5500
rect 7640 5460 7650 5500
rect 7590 5440 7650 5460
rect 7770 6000 7830 6020
rect 7770 5960 7780 6000
rect 7820 5960 7830 6000
rect 7770 5900 7830 5960
rect 7770 5860 7780 5900
rect 7820 5860 7830 5900
rect 7770 5800 7830 5860
rect 7770 5760 7780 5800
rect 7820 5760 7830 5800
rect 7770 5700 7830 5760
rect 7770 5660 7780 5700
rect 7820 5660 7830 5700
rect 7770 5600 7830 5660
rect 7770 5560 7780 5600
rect 7820 5560 7830 5600
rect 7770 5500 7830 5560
rect 7770 5460 7780 5500
rect 7820 5460 7830 5500
rect 7770 5440 7830 5460
rect 7950 6000 8010 6020
rect 7950 5960 7960 6000
rect 8000 5960 8010 6000
rect 7950 5900 8010 5960
rect 7950 5860 7960 5900
rect 8000 5860 8010 5900
rect 7950 5800 8010 5860
rect 7950 5760 7960 5800
rect 8000 5760 8010 5800
rect 7950 5700 8010 5760
rect 7950 5660 7960 5700
rect 8000 5660 8010 5700
rect 7950 5600 8010 5660
rect 7950 5560 7960 5600
rect 8000 5560 8010 5600
rect 7950 5500 8010 5560
rect 7950 5460 7960 5500
rect 8000 5460 8010 5500
rect 7950 5440 8010 5460
rect 8130 6000 8190 6020
rect 8130 5960 8140 6000
rect 8180 5960 8190 6000
rect 8130 5900 8190 5960
rect 8130 5860 8140 5900
rect 8180 5860 8190 5900
rect 8130 5800 8190 5860
rect 8130 5760 8140 5800
rect 8180 5760 8190 5800
rect 8130 5700 8190 5760
rect 8130 5660 8140 5700
rect 8180 5660 8190 5700
rect 8130 5600 8190 5660
rect 8130 5560 8140 5600
rect 8180 5560 8190 5600
rect 8130 5500 8190 5560
rect 8130 5460 8140 5500
rect 8180 5460 8190 5500
rect 8130 5440 8190 5460
rect 8310 6000 8370 6020
rect 8310 5960 8320 6000
rect 8360 5960 8370 6000
rect 8310 5900 8370 5960
rect 8310 5860 8320 5900
rect 8360 5860 8370 5900
rect 8310 5800 8370 5860
rect 8310 5760 8320 5800
rect 8360 5760 8370 5800
rect 8310 5700 8370 5760
rect 8310 5660 8320 5700
rect 8360 5660 8370 5700
rect 8310 5600 8370 5660
rect 8310 5560 8320 5600
rect 8360 5560 8370 5600
rect 8310 5500 8370 5560
rect 8310 5460 8320 5500
rect 8360 5460 8370 5500
rect 8310 5440 8370 5460
rect 8490 6000 8550 6020
rect 8490 5960 8500 6000
rect 8540 5960 8550 6000
rect 8490 5900 8550 5960
rect 8490 5860 8500 5900
rect 8540 5860 8550 5900
rect 8490 5800 8550 5860
rect 8490 5760 8500 5800
rect 8540 5760 8550 5800
rect 8490 5700 8550 5760
rect 8490 5660 8500 5700
rect 8540 5660 8550 5700
rect 8490 5600 8550 5660
rect 8490 5560 8500 5600
rect 8540 5560 8550 5600
rect 8490 5500 8550 5560
rect 8490 5460 8500 5500
rect 8540 5460 8550 5500
rect 8490 5440 8550 5460
rect 8670 6000 8730 6020
rect 8670 5960 8680 6000
rect 8720 5960 8730 6000
rect 8670 5900 8730 5960
rect 8670 5860 8680 5900
rect 8720 5860 8730 5900
rect 8670 5800 8730 5860
rect 8670 5760 8680 5800
rect 8720 5760 8730 5800
rect 8670 5700 8730 5760
rect 8670 5660 8680 5700
rect 8720 5660 8730 5700
rect 8670 5600 8730 5660
rect 8670 5560 8680 5600
rect 8720 5560 8730 5600
rect 8670 5500 8730 5560
rect 8670 5460 8680 5500
rect 8720 5460 8730 5500
rect 8670 5440 8730 5460
rect 8850 6000 8910 6020
rect 8850 5960 8860 6000
rect 8900 5960 8910 6000
rect 8850 5900 8910 5960
rect 8850 5860 8860 5900
rect 8900 5860 8910 5900
rect 8850 5800 8910 5860
rect 8850 5760 8860 5800
rect 8900 5760 8910 5800
rect 8850 5700 8910 5760
rect 8850 5660 8860 5700
rect 8900 5660 8910 5700
rect 8850 5600 8910 5660
rect 8850 5560 8860 5600
rect 8900 5560 8910 5600
rect 8850 5500 8910 5560
rect 8850 5460 8860 5500
rect 8900 5460 8910 5500
rect 8850 5440 8910 5460
rect 9030 6000 9090 6020
rect 9030 5960 9040 6000
rect 9080 5960 9090 6000
rect 9030 5900 9090 5960
rect 9030 5860 9040 5900
rect 9080 5860 9090 5900
rect 9030 5800 9090 5860
rect 9030 5760 9040 5800
rect 9080 5760 9090 5800
rect 9030 5700 9090 5760
rect 9030 5660 9040 5700
rect 9080 5660 9090 5700
rect 9030 5600 9090 5660
rect 9030 5560 9040 5600
rect 9080 5560 9090 5600
rect 9030 5500 9090 5560
rect 9030 5460 9040 5500
rect 9080 5460 9090 5500
rect 9030 5440 9090 5460
rect 9210 6000 9270 6020
rect 9210 5960 9220 6000
rect 9260 5960 9270 6000
rect 9210 5900 9270 5960
rect 9210 5860 9220 5900
rect 9260 5860 9270 5900
rect 9210 5800 9270 5860
rect 9210 5760 9220 5800
rect 9260 5760 9270 5800
rect 9210 5700 9270 5760
rect 9210 5660 9220 5700
rect 9260 5660 9270 5700
rect 9210 5600 9270 5660
rect 9210 5560 9220 5600
rect 9260 5560 9270 5600
rect 9210 5500 9270 5560
rect 9210 5460 9220 5500
rect 9260 5460 9270 5500
rect 9210 5440 9270 5460
rect 9390 6000 9450 6020
rect 9390 5960 9400 6000
rect 9440 5960 9450 6000
rect 9390 5900 9450 5960
rect 9390 5860 9400 5900
rect 9440 5860 9450 5900
rect 9390 5800 9450 5860
rect 9390 5760 9400 5800
rect 9440 5760 9450 5800
rect 9390 5700 9450 5760
rect 9390 5660 9400 5700
rect 9440 5660 9450 5700
rect 9390 5600 9450 5660
rect 9390 5560 9400 5600
rect 9440 5560 9450 5600
rect 9390 5500 9450 5560
rect 9390 5460 9400 5500
rect 9440 5460 9450 5500
rect 9390 5440 9450 5460
rect 9570 6000 9630 6020
rect 9570 5960 9580 6000
rect 9620 5960 9630 6000
rect 9570 5900 9630 5960
rect 9570 5860 9580 5900
rect 9620 5860 9630 5900
rect 9570 5800 9630 5860
rect 9570 5760 9580 5800
rect 9620 5760 9630 5800
rect 9570 5700 9630 5760
rect 9570 5660 9580 5700
rect 9620 5660 9630 5700
rect 9570 5600 9630 5660
rect 9570 5560 9580 5600
rect 9620 5560 9630 5600
rect 9570 5500 9630 5560
rect 9570 5460 9580 5500
rect 9620 5460 9630 5500
rect 9570 5440 9630 5460
rect 9750 6000 9810 6020
rect 9750 5960 9760 6000
rect 9800 5960 9810 6000
rect 9750 5900 9810 5960
rect 9750 5860 9760 5900
rect 9800 5860 9810 5900
rect 9750 5800 9810 5860
rect 9750 5760 9760 5800
rect 9800 5760 9810 5800
rect 9750 5700 9810 5760
rect 9750 5660 9760 5700
rect 9800 5660 9810 5700
rect 9750 5600 9810 5660
rect 9750 5560 9760 5600
rect 9800 5560 9810 5600
rect 9750 5500 9810 5560
rect 9750 5460 9760 5500
rect 9800 5460 9810 5500
rect 9750 5440 9810 5460
rect 9880 5810 9920 6180
rect 10720 6040 10800 6080
rect 10720 6020 10740 6040
rect 10780 6020 10800 6040
rect 6700 5400 6740 5440
rect 7060 5400 7100 5440
rect 7420 5400 7460 5440
rect 7780 5400 7820 5440
rect 8140 5400 8180 5440
rect 8500 5400 8540 5440
rect 8860 5400 8900 5440
rect 9220 5400 9260 5440
rect 9580 5400 9620 5440
rect 6680 5380 6760 5400
rect 6680 5340 6700 5380
rect 6740 5340 6760 5380
rect 6680 5320 6760 5340
rect 7040 5380 7120 5400
rect 7040 5340 7060 5380
rect 7100 5340 7120 5380
rect 7040 5320 7120 5340
rect 7400 5380 7480 5400
rect 7400 5340 7420 5380
rect 7460 5340 7480 5380
rect 7400 5320 7480 5340
rect 7760 5380 7840 5400
rect 7760 5340 7780 5380
rect 7820 5340 7840 5380
rect 7760 5320 7840 5340
rect 7940 5380 8020 5400
rect 7940 5340 7960 5380
rect 8000 5340 8020 5380
rect 7940 5320 8020 5340
rect 8120 5380 8200 5400
rect 8120 5340 8140 5380
rect 8180 5340 8200 5380
rect 8120 5320 8200 5340
rect 8480 5380 8560 5400
rect 8480 5340 8500 5380
rect 8540 5340 8560 5380
rect 8480 5320 8560 5340
rect 8840 5380 8920 5400
rect 8840 5340 8860 5380
rect 8900 5340 8920 5380
rect 8840 5320 8920 5340
rect 9200 5380 9280 5400
rect 9200 5340 9220 5380
rect 9260 5340 9280 5380
rect 9200 5320 9280 5340
rect 9380 5380 9460 5400
rect 9380 5340 9400 5380
rect 9440 5340 9460 5380
rect 9380 5320 9460 5340
rect 9560 5380 9640 5400
rect 9560 5340 9580 5380
rect 9620 5340 9640 5380
rect 9560 5320 9640 5340
rect 9880 5270 9920 5650
rect 10260 5980 10610 6020
rect 10910 5980 11260 6020
rect 10260 5810 10300 5980
rect 10380 5940 10420 5980
rect 11100 5940 11140 5980
rect 10370 5920 10430 5940
rect 10370 5880 10380 5920
rect 10420 5880 10430 5920
rect 10370 5860 10430 5880
rect 10720 5920 10800 5940
rect 10720 5880 10740 5920
rect 10780 5880 10800 5920
rect 10720 5860 10800 5880
rect 11090 5920 11150 5940
rect 11090 5880 11100 5920
rect 11140 5880 11150 5920
rect 11090 5860 11150 5880
rect 10380 5820 10420 5860
rect 10740 5820 10780 5860
rect 11100 5820 11140 5860
rect 10260 5480 10300 5650
rect 10370 5800 10430 5820
rect 10370 5760 10380 5800
rect 10420 5760 10430 5800
rect 10370 5700 10430 5760
rect 10370 5660 10380 5700
rect 10420 5660 10430 5700
rect 10370 5640 10430 5660
rect 10550 5800 10610 5820
rect 10550 5760 10560 5800
rect 10600 5760 10610 5800
rect 10550 5700 10610 5760
rect 10550 5660 10560 5700
rect 10600 5660 10610 5700
rect 10550 5640 10610 5660
rect 10730 5800 10790 5820
rect 10730 5760 10740 5800
rect 10780 5760 10790 5800
rect 10730 5700 10790 5760
rect 10730 5660 10740 5700
rect 10780 5660 10790 5700
rect 10730 5640 10790 5660
rect 10910 5800 10970 5820
rect 10910 5760 10920 5800
rect 10960 5760 10970 5800
rect 10910 5700 10970 5760
rect 10910 5660 10920 5700
rect 10960 5660 10970 5700
rect 10910 5640 10970 5660
rect 11090 5800 11150 5820
rect 11090 5760 11100 5800
rect 11140 5760 11150 5800
rect 11090 5700 11150 5760
rect 11090 5660 11100 5700
rect 11140 5660 11150 5700
rect 11090 5640 11150 5660
rect 11220 5810 11260 5980
rect 10560 5600 10600 5640
rect 10920 5600 10960 5640
rect 10520 5580 10600 5600
rect 10520 5540 10540 5580
rect 10580 5540 10600 5580
rect 10520 5520 10600 5540
rect 10720 5580 10800 5600
rect 10720 5540 10740 5580
rect 10780 5540 10800 5580
rect 10720 5520 10800 5540
rect 10920 5580 11000 5600
rect 10920 5540 10940 5580
rect 10980 5540 11000 5580
rect 10920 5520 11000 5540
rect 11220 5480 11260 5650
rect 10260 5440 10610 5480
rect 10910 5440 11260 5480
rect 6400 5230 8080 5270
rect 8240 5230 9920 5270
rect 6600 4860 6680 4880
rect 6600 4840 6620 4860
rect 6660 4840 6680 4860
rect 8680 4860 8760 4880
rect 8680 4840 8700 4860
rect 5300 4800 6560 4840
rect 6720 4800 7980 4840
rect 5300 4630 5340 4800
rect 5520 4740 5600 4760
rect 5520 4700 5540 4740
rect 5580 4700 5600 4740
rect 5520 4680 5600 4700
rect 5650 4740 5710 4760
rect 5650 4700 5660 4740
rect 5700 4700 5710 4740
rect 5650 4680 5710 4700
rect 5890 4740 5950 4760
rect 5890 4700 5900 4740
rect 5940 4700 5950 4740
rect 5890 4680 5950 4700
rect 6130 4740 6190 4760
rect 6130 4700 6140 4740
rect 6180 4700 6190 4740
rect 6130 4680 6190 4700
rect 6240 4740 6320 4760
rect 6240 4700 6260 4740
rect 6300 4700 6320 4740
rect 6240 4680 6320 4700
rect 6370 4740 6430 4760
rect 6370 4700 6380 4740
rect 6420 4700 6430 4740
rect 6370 4680 6430 4700
rect 6610 4740 6670 4760
rect 6610 4700 6620 4740
rect 6660 4700 6670 4740
rect 6610 4680 6670 4700
rect 6850 4740 6910 4760
rect 6850 4700 6860 4740
rect 6900 4700 6910 4740
rect 6850 4680 6910 4700
rect 6960 4740 7040 4760
rect 6960 4700 6980 4740
rect 7020 4700 7040 4740
rect 6960 4680 7040 4700
rect 7090 4740 7150 4760
rect 7090 4700 7100 4740
rect 7140 4700 7150 4740
rect 7090 4680 7150 4700
rect 7330 4740 7390 4760
rect 7330 4700 7340 4740
rect 7380 4700 7390 4740
rect 7330 4680 7390 4700
rect 7570 4740 7630 4760
rect 7570 4700 7580 4740
rect 7620 4700 7630 4740
rect 7570 4680 7630 4700
rect 7680 4740 7760 4760
rect 7680 4700 7700 4740
rect 7740 4700 7760 4740
rect 7680 4680 7760 4700
rect 5540 4640 5580 4680
rect 5660 4640 5700 4680
rect 5900 4640 5940 4680
rect 6140 4640 6180 4680
rect 6260 4640 6300 4680
rect 6380 4640 6420 4680
rect 6620 4640 6660 4680
rect 6860 4640 6900 4680
rect 6980 4640 7020 4680
rect 7100 4640 7140 4680
rect 7340 4640 7380 4680
rect 7580 4640 7620 4680
rect 7700 4640 7740 4680
rect 5300 4300 5340 4470
rect 5410 4620 5470 4640
rect 5410 4580 5420 4620
rect 5460 4580 5470 4620
rect 5410 4520 5470 4580
rect 5410 4480 5420 4520
rect 5460 4480 5470 4520
rect 5410 4400 5470 4480
rect 5530 4620 5590 4640
rect 5530 4580 5540 4620
rect 5580 4580 5590 4620
rect 5530 4520 5590 4580
rect 5530 4480 5540 4520
rect 5580 4480 5590 4520
rect 5530 4460 5590 4480
rect 5650 4620 5710 4640
rect 5650 4580 5660 4620
rect 5700 4580 5710 4620
rect 5650 4520 5710 4580
rect 5650 4480 5660 4520
rect 5700 4480 5710 4520
rect 5650 4460 5710 4480
rect 5770 4620 5830 4640
rect 5770 4580 5780 4620
rect 5820 4580 5830 4620
rect 5770 4520 5830 4580
rect 5770 4480 5780 4520
rect 5820 4480 5830 4520
rect 5770 4460 5830 4480
rect 5890 4620 5950 4640
rect 5890 4580 5900 4620
rect 5940 4580 5950 4620
rect 5890 4520 5950 4580
rect 5890 4480 5900 4520
rect 5940 4480 5950 4520
rect 5890 4460 5950 4480
rect 6010 4620 6070 4640
rect 6010 4580 6020 4620
rect 6060 4580 6070 4620
rect 6010 4520 6070 4580
rect 6010 4480 6020 4520
rect 6060 4480 6070 4520
rect 6010 4460 6070 4480
rect 6130 4620 6190 4640
rect 6130 4580 6140 4620
rect 6180 4580 6190 4620
rect 6130 4520 6190 4580
rect 6130 4480 6140 4520
rect 6180 4480 6190 4520
rect 6130 4460 6190 4480
rect 6250 4620 6310 4640
rect 6250 4580 6260 4620
rect 6300 4580 6310 4620
rect 6250 4520 6310 4580
rect 6250 4480 6260 4520
rect 6300 4480 6310 4520
rect 6250 4460 6310 4480
rect 6370 4620 6430 4640
rect 6370 4580 6380 4620
rect 6420 4580 6430 4620
rect 6370 4520 6430 4580
rect 6370 4480 6380 4520
rect 6420 4480 6430 4520
rect 6370 4460 6430 4480
rect 6490 4620 6550 4640
rect 6490 4580 6500 4620
rect 6540 4580 6550 4620
rect 6490 4520 6550 4580
rect 6490 4480 6500 4520
rect 6540 4480 6550 4520
rect 6490 4460 6550 4480
rect 6610 4620 6670 4640
rect 6610 4580 6620 4620
rect 6660 4580 6670 4620
rect 6610 4520 6670 4580
rect 6610 4480 6620 4520
rect 6660 4480 6670 4520
rect 6610 4460 6670 4480
rect 6730 4620 6790 4640
rect 6730 4580 6740 4620
rect 6780 4580 6790 4620
rect 6730 4520 6790 4580
rect 6730 4480 6740 4520
rect 6780 4480 6790 4520
rect 6730 4460 6790 4480
rect 6850 4620 6910 4640
rect 6850 4580 6860 4620
rect 6900 4580 6910 4620
rect 6850 4520 6910 4580
rect 6850 4480 6860 4520
rect 6900 4480 6910 4520
rect 6850 4460 6910 4480
rect 6970 4620 7030 4640
rect 6970 4580 6980 4620
rect 7020 4580 7030 4620
rect 6970 4520 7030 4580
rect 6970 4480 6980 4520
rect 7020 4480 7030 4520
rect 6970 4460 7030 4480
rect 7090 4620 7150 4640
rect 7090 4580 7100 4620
rect 7140 4580 7150 4620
rect 7090 4520 7150 4580
rect 7090 4480 7100 4520
rect 7140 4480 7150 4520
rect 7090 4460 7150 4480
rect 7210 4620 7270 4640
rect 7210 4580 7220 4620
rect 7260 4580 7270 4620
rect 7210 4520 7270 4580
rect 7210 4480 7220 4520
rect 7260 4480 7270 4520
rect 7210 4460 7270 4480
rect 7330 4620 7390 4640
rect 7330 4580 7340 4620
rect 7380 4580 7390 4620
rect 7330 4520 7390 4580
rect 7330 4480 7340 4520
rect 7380 4480 7390 4520
rect 7330 4460 7390 4480
rect 7450 4620 7510 4640
rect 7450 4580 7460 4620
rect 7500 4580 7510 4620
rect 7450 4520 7510 4580
rect 7450 4480 7460 4520
rect 7500 4480 7510 4520
rect 7450 4460 7510 4480
rect 7570 4620 7630 4640
rect 7570 4580 7580 4620
rect 7620 4580 7630 4620
rect 7570 4520 7630 4580
rect 7570 4480 7580 4520
rect 7620 4480 7630 4520
rect 7570 4460 7630 4480
rect 7690 4620 7750 4640
rect 7690 4580 7700 4620
rect 7740 4580 7750 4620
rect 7690 4520 7750 4580
rect 7690 4480 7700 4520
rect 7740 4480 7750 4520
rect 7690 4460 7750 4480
rect 7810 4620 7870 4640
rect 7810 4580 7820 4620
rect 7860 4580 7870 4620
rect 7810 4520 7870 4580
rect 7810 4480 7820 4520
rect 7860 4480 7870 4520
rect 5780 4420 5820 4460
rect 6020 4420 6060 4460
rect 6500 4420 6540 4460
rect 6740 4420 6780 4460
rect 7220 4420 7260 4460
rect 7460 4420 7500 4460
rect 5410 4360 5420 4400
rect 5460 4360 5470 4400
rect 5410 4340 5470 4360
rect 5580 4400 5660 4420
rect 5580 4360 5600 4400
rect 5640 4360 5660 4400
rect 5580 4340 5660 4360
rect 5760 4400 5840 4420
rect 5760 4360 5780 4400
rect 5820 4360 5840 4400
rect 5760 4340 5840 4360
rect 6000 4400 6080 4420
rect 6000 4360 6020 4400
rect 6060 4360 6080 4400
rect 6000 4340 6080 4360
rect 6240 4400 6320 4420
rect 6240 4360 6260 4400
rect 6300 4360 6320 4400
rect 6240 4340 6320 4360
rect 6480 4400 6560 4420
rect 6480 4360 6500 4400
rect 6540 4360 6560 4400
rect 6480 4340 6560 4360
rect 6720 4400 6800 4420
rect 6720 4360 6740 4400
rect 6780 4360 6800 4400
rect 6720 4340 6800 4360
rect 6960 4400 7040 4420
rect 6960 4360 6980 4400
rect 7020 4360 7040 4400
rect 6960 4340 7040 4360
rect 7200 4400 7280 4420
rect 7200 4360 7220 4400
rect 7260 4360 7280 4400
rect 7200 4340 7280 4360
rect 7440 4400 7520 4420
rect 7440 4360 7460 4400
rect 7500 4360 7520 4400
rect 7440 4340 7520 4360
rect 7630 4400 7690 4420
rect 7630 4360 7640 4400
rect 7680 4360 7690 4400
rect 7630 4340 7690 4360
rect 7810 4400 7870 4480
rect 7810 4360 7820 4400
rect 7860 4360 7870 4400
rect 7810 4340 7870 4360
rect 7940 4630 7980 4800
rect 5420 4300 5460 4340
rect 7820 4300 7860 4340
rect 7940 4300 7980 4470
rect 5300 4260 6560 4300
rect 6720 4260 7980 4300
rect 8340 4820 8700 4840
rect 8740 4840 8760 4860
rect 8920 4860 9000 4880
rect 8920 4840 8940 4860
rect 8740 4820 8940 4840
rect 8980 4840 9000 4860
rect 9160 4860 9240 4880
rect 9160 4840 9180 4860
rect 8980 4820 9180 4840
rect 9220 4840 9240 4860
rect 9400 4860 9480 4880
rect 9400 4840 9420 4860
rect 9220 4820 9420 4840
rect 9460 4840 9480 4860
rect 9640 4860 9720 4880
rect 9640 4840 9660 4860
rect 9700 4840 9720 4860
rect 9880 4860 9960 4880
rect 9880 4840 9900 4860
rect 9460 4820 9600 4840
rect 9760 4820 9900 4840
rect 9940 4840 9960 4860
rect 10120 4860 10200 4880
rect 10120 4840 10140 4860
rect 9940 4820 10140 4840
rect 10180 4840 10200 4860
rect 10360 4860 10440 4880
rect 10360 4840 10380 4860
rect 10180 4820 10380 4840
rect 10420 4840 10440 4860
rect 10600 4860 10680 4880
rect 10600 4840 10620 4860
rect 10420 4820 10620 4840
rect 10660 4840 10680 4860
rect 10660 4820 11020 4840
rect 8340 4800 9600 4820
rect 9760 4800 11020 4820
rect 8340 4630 8380 4800
rect 8560 4740 8640 4760
rect 8560 4700 8580 4740
rect 8620 4700 8640 4740
rect 8560 4680 8640 4700
rect 8690 4740 8750 4760
rect 8690 4700 8700 4740
rect 8740 4700 8750 4740
rect 8690 4680 8750 4700
rect 8930 4740 8990 4760
rect 8930 4700 8940 4740
rect 8980 4700 8990 4740
rect 8930 4680 8990 4700
rect 9170 4740 9230 4760
rect 9170 4700 9180 4740
rect 9220 4700 9230 4740
rect 9170 4680 9230 4700
rect 9280 4740 9360 4760
rect 9280 4700 9300 4740
rect 9340 4700 9360 4740
rect 9280 4680 9360 4700
rect 9410 4740 9470 4760
rect 9410 4700 9420 4740
rect 9460 4700 9470 4740
rect 9410 4680 9470 4700
rect 9650 4740 9710 4760
rect 9650 4700 9660 4740
rect 9700 4700 9710 4740
rect 9650 4680 9710 4700
rect 9890 4740 9950 4760
rect 9890 4700 9900 4740
rect 9940 4700 9950 4740
rect 9890 4680 9950 4700
rect 10000 4740 10080 4760
rect 10000 4700 10020 4740
rect 10060 4700 10080 4740
rect 10000 4680 10080 4700
rect 10130 4740 10190 4760
rect 10130 4700 10140 4740
rect 10180 4700 10190 4740
rect 10130 4680 10190 4700
rect 10370 4740 10430 4760
rect 10370 4700 10380 4740
rect 10420 4700 10430 4740
rect 10370 4680 10430 4700
rect 10610 4740 10670 4760
rect 10610 4700 10620 4740
rect 10660 4700 10670 4740
rect 10610 4680 10670 4700
rect 10720 4740 10800 4760
rect 10720 4700 10740 4740
rect 10780 4700 10800 4740
rect 10720 4680 10800 4700
rect 8580 4640 8620 4680
rect 8700 4640 8740 4680
rect 8940 4640 8980 4680
rect 9180 4640 9220 4680
rect 9300 4640 9340 4680
rect 9420 4640 9460 4680
rect 9660 4640 9700 4680
rect 9900 4640 9940 4680
rect 10020 4640 10060 4680
rect 10140 4640 10180 4680
rect 10380 4640 10420 4680
rect 10620 4640 10660 4680
rect 10740 4640 10780 4680
rect 8340 4300 8380 4470
rect 8450 4620 8510 4640
rect 8450 4580 8460 4620
rect 8500 4580 8510 4620
rect 8450 4520 8510 4580
rect 8450 4480 8460 4520
rect 8500 4480 8510 4520
rect 8450 4400 8510 4480
rect 8570 4620 8630 4640
rect 8570 4580 8580 4620
rect 8620 4580 8630 4620
rect 8570 4520 8630 4580
rect 8570 4480 8580 4520
rect 8620 4480 8630 4520
rect 8570 4460 8630 4480
rect 8690 4620 8750 4640
rect 8690 4580 8700 4620
rect 8740 4580 8750 4620
rect 8690 4520 8750 4580
rect 8690 4480 8700 4520
rect 8740 4480 8750 4520
rect 8690 4460 8750 4480
rect 8810 4620 8870 4640
rect 8810 4580 8820 4620
rect 8860 4580 8870 4620
rect 8810 4520 8870 4580
rect 8810 4480 8820 4520
rect 8860 4480 8870 4520
rect 8810 4460 8870 4480
rect 8930 4620 8990 4640
rect 8930 4580 8940 4620
rect 8980 4580 8990 4620
rect 8930 4520 8990 4580
rect 8930 4480 8940 4520
rect 8980 4480 8990 4520
rect 8930 4460 8990 4480
rect 9050 4620 9110 4640
rect 9050 4580 9060 4620
rect 9100 4580 9110 4620
rect 9050 4520 9110 4580
rect 9050 4480 9060 4520
rect 9100 4480 9110 4520
rect 9050 4460 9110 4480
rect 9170 4620 9230 4640
rect 9170 4580 9180 4620
rect 9220 4580 9230 4620
rect 9170 4520 9230 4580
rect 9170 4480 9180 4520
rect 9220 4480 9230 4520
rect 9170 4460 9230 4480
rect 9290 4620 9350 4640
rect 9290 4580 9300 4620
rect 9340 4580 9350 4620
rect 9290 4520 9350 4580
rect 9290 4480 9300 4520
rect 9340 4480 9350 4520
rect 9290 4460 9350 4480
rect 9410 4620 9470 4640
rect 9410 4580 9420 4620
rect 9460 4580 9470 4620
rect 9410 4520 9470 4580
rect 9410 4480 9420 4520
rect 9460 4480 9470 4520
rect 9410 4460 9470 4480
rect 9530 4620 9590 4640
rect 9530 4580 9540 4620
rect 9580 4580 9590 4620
rect 9530 4520 9590 4580
rect 9530 4480 9540 4520
rect 9580 4480 9590 4520
rect 9530 4460 9590 4480
rect 9650 4620 9710 4640
rect 9650 4580 9660 4620
rect 9700 4580 9710 4620
rect 9650 4520 9710 4580
rect 9650 4480 9660 4520
rect 9700 4480 9710 4520
rect 9650 4460 9710 4480
rect 9770 4620 9830 4640
rect 9770 4580 9780 4620
rect 9820 4580 9830 4620
rect 9770 4520 9830 4580
rect 9770 4480 9780 4520
rect 9820 4480 9830 4520
rect 9770 4460 9830 4480
rect 9890 4620 9950 4640
rect 9890 4580 9900 4620
rect 9940 4580 9950 4620
rect 9890 4520 9950 4580
rect 9890 4480 9900 4520
rect 9940 4480 9950 4520
rect 9890 4460 9950 4480
rect 10010 4620 10070 4640
rect 10010 4580 10020 4620
rect 10060 4580 10070 4620
rect 10010 4520 10070 4580
rect 10010 4480 10020 4520
rect 10060 4480 10070 4520
rect 10010 4460 10070 4480
rect 10130 4620 10190 4640
rect 10130 4580 10140 4620
rect 10180 4580 10190 4620
rect 10130 4520 10190 4580
rect 10130 4480 10140 4520
rect 10180 4480 10190 4520
rect 10130 4460 10190 4480
rect 10250 4620 10310 4640
rect 10250 4580 10260 4620
rect 10300 4580 10310 4620
rect 10250 4520 10310 4580
rect 10250 4480 10260 4520
rect 10300 4480 10310 4520
rect 10250 4460 10310 4480
rect 10370 4620 10430 4640
rect 10370 4580 10380 4620
rect 10420 4580 10430 4620
rect 10370 4520 10430 4580
rect 10370 4480 10380 4520
rect 10420 4480 10430 4520
rect 10370 4460 10430 4480
rect 10490 4620 10550 4640
rect 10490 4580 10500 4620
rect 10540 4580 10550 4620
rect 10490 4520 10550 4580
rect 10490 4480 10500 4520
rect 10540 4480 10550 4520
rect 10490 4460 10550 4480
rect 10610 4620 10670 4640
rect 10610 4580 10620 4620
rect 10660 4580 10670 4620
rect 10610 4520 10670 4580
rect 10610 4480 10620 4520
rect 10660 4480 10670 4520
rect 10610 4460 10670 4480
rect 10730 4620 10790 4640
rect 10730 4580 10740 4620
rect 10780 4580 10790 4620
rect 10730 4520 10790 4580
rect 10730 4480 10740 4520
rect 10780 4480 10790 4520
rect 10730 4460 10790 4480
rect 10850 4620 10910 4640
rect 10850 4580 10860 4620
rect 10900 4580 10910 4620
rect 10850 4520 10910 4580
rect 10850 4480 10860 4520
rect 10900 4480 10910 4520
rect 8820 4420 8860 4460
rect 9060 4420 9100 4460
rect 9540 4420 9580 4460
rect 9780 4420 9820 4460
rect 10260 4420 10300 4460
rect 10500 4420 10540 4460
rect 8450 4360 8460 4400
rect 8500 4360 8510 4400
rect 8450 4340 8510 4360
rect 8630 4400 8690 4420
rect 8630 4360 8640 4400
rect 8680 4360 8690 4400
rect 8630 4340 8690 4360
rect 8800 4400 8880 4420
rect 8800 4360 8820 4400
rect 8860 4360 8880 4400
rect 8800 4340 8880 4360
rect 9040 4400 9120 4420
rect 9040 4360 9060 4400
rect 9100 4360 9120 4400
rect 9040 4340 9120 4360
rect 9280 4400 9360 4420
rect 9280 4360 9300 4400
rect 9340 4360 9360 4400
rect 9280 4340 9360 4360
rect 9520 4400 9600 4420
rect 9520 4360 9540 4400
rect 9580 4360 9600 4400
rect 9520 4340 9600 4360
rect 9760 4400 9840 4420
rect 9760 4360 9780 4400
rect 9820 4360 9840 4400
rect 9760 4340 9840 4360
rect 10000 4400 10080 4420
rect 10000 4360 10020 4400
rect 10060 4360 10080 4400
rect 10000 4340 10080 4360
rect 10240 4400 10320 4420
rect 10240 4360 10260 4400
rect 10300 4360 10320 4400
rect 10240 4340 10320 4360
rect 10480 4400 10560 4420
rect 10480 4360 10500 4400
rect 10540 4360 10560 4400
rect 10480 4340 10560 4360
rect 10660 4400 10740 4420
rect 10660 4360 10680 4400
rect 10720 4360 10740 4400
rect 10660 4340 10740 4360
rect 10850 4400 10910 4480
rect 10850 4360 10860 4400
rect 10900 4360 10910 4400
rect 10850 4340 10910 4360
rect 10980 4630 11020 4800
rect 8460 4300 8500 4340
rect 10860 4300 10900 4340
rect 10980 4300 11020 4470
rect 8340 4260 9600 4300
rect 9760 4260 11020 4300
rect 250 4030 4270 4110
rect -90 3430 260 3450
rect -90 3390 -70 3430
rect -30 3390 30 3430
rect 70 3390 130 3430
rect 170 3390 260 3430
rect -90 3370 260 3390
rect 1300 2750 1550 4030
rect 2660 2750 2910 4030
rect 4020 2750 4270 4030
rect 6160 4140 6820 4180
rect 6980 4140 7640 4180
rect 6160 3930 6200 4140
rect 6380 4080 6460 4100
rect 6380 4040 6400 4080
rect 6440 4040 6460 4080
rect 6380 4020 6460 4040
rect 6260 3990 6340 4010
rect 6260 3950 6280 3990
rect 6320 3950 6340 3990
rect 6260 3930 6340 3950
rect 6510 3990 6570 4010
rect 6510 3950 6520 3990
rect 6560 3950 6570 3990
rect 6510 3930 6570 3950
rect 6740 3990 6820 4010
rect 6740 3950 6760 3990
rect 6800 3950 6820 3990
rect 6740 3930 6820 3950
rect 6990 3990 7050 4010
rect 6990 3950 7000 3990
rect 7040 3950 7050 3990
rect 6990 3930 7050 3950
rect 7220 3990 7300 4010
rect 7220 3950 7240 3990
rect 7280 3950 7300 3990
rect 7220 3930 7300 3950
rect 7470 3990 7530 4010
rect 7470 3950 7480 3990
rect 7520 3950 7530 3990
rect 7470 3930 7530 3950
rect 7600 3930 7640 4140
rect 6280 3890 6320 3930
rect 6520 3890 6560 3930
rect 6760 3890 6800 3930
rect 7000 3890 7040 3930
rect 7240 3890 7280 3930
rect 7480 3890 7520 3930
rect 6270 3870 6330 3890
rect 6270 3830 6280 3870
rect 6320 3830 6330 3870
rect 6270 3810 6330 3830
rect 6390 3870 6450 3890
rect 6390 3830 6400 3870
rect 6440 3830 6450 3870
rect 6390 3810 6450 3830
rect 6510 3870 6570 3890
rect 6510 3830 6520 3870
rect 6560 3830 6570 3870
rect 6510 3810 6570 3830
rect 6630 3870 6690 3890
rect 6630 3830 6640 3870
rect 6680 3830 6690 3870
rect 6630 3810 6690 3830
rect 6750 3870 6810 3890
rect 6750 3830 6760 3870
rect 6800 3830 6810 3870
rect 6750 3810 6810 3830
rect 6870 3870 6930 3890
rect 6870 3830 6880 3870
rect 6920 3830 6930 3870
rect 6870 3810 6930 3830
rect 6990 3870 7050 3890
rect 6990 3830 7000 3870
rect 7040 3830 7050 3870
rect 6990 3810 7050 3830
rect 7110 3870 7170 3890
rect 7110 3830 7120 3870
rect 7160 3830 7170 3870
rect 7110 3810 7170 3830
rect 7230 3870 7290 3890
rect 7230 3830 7240 3870
rect 7280 3830 7290 3870
rect 7230 3810 7290 3830
rect 7350 3870 7410 3890
rect 7350 3830 7360 3870
rect 7400 3830 7410 3870
rect 7350 3810 7410 3830
rect 7470 3870 7530 3890
rect 7470 3830 7480 3870
rect 7520 3830 7530 3870
rect 7470 3810 7530 3830
rect 7580 3810 7600 3890
rect 8680 4140 9340 4180
rect 9500 4140 10160 4180
rect 8680 3930 8720 4140
rect 9860 4080 9940 4100
rect 9860 4040 9880 4080
rect 9920 4040 9940 4080
rect 9860 4020 9940 4040
rect 8790 3990 8850 4010
rect 8790 3950 8800 3990
rect 8840 3950 8850 3990
rect 8790 3930 8850 3950
rect 9020 3990 9100 4010
rect 9020 3950 9040 3990
rect 9080 3950 9100 3990
rect 9020 3930 9100 3950
rect 9270 3990 9330 4010
rect 9270 3950 9280 3990
rect 9320 3950 9330 3990
rect 9270 3930 9330 3950
rect 9500 3990 9580 4010
rect 9500 3950 9520 3990
rect 9560 3950 9580 3990
rect 9500 3930 9580 3950
rect 9750 3990 9810 4010
rect 9750 3950 9760 3990
rect 9800 3950 9810 3990
rect 9750 3930 9810 3950
rect 9980 3990 10060 4010
rect 9980 3950 10000 3990
rect 10040 3950 10060 3990
rect 9980 3930 10060 3950
rect 10120 3930 10160 4140
rect 6400 3770 6440 3810
rect 6640 3770 6680 3810
rect 6880 3770 6920 3810
rect 7120 3770 7160 3810
rect 7360 3770 7400 3810
rect 7640 3810 7660 3890
rect 8660 3810 8680 3890
rect 8800 3890 8840 3930
rect 9040 3890 9080 3930
rect 9280 3890 9320 3930
rect 9520 3890 9560 3930
rect 9760 3890 9800 3930
rect 10000 3890 10040 3930
rect 6160 3650 6200 3770
rect 6260 3750 6340 3770
rect 6260 3710 6280 3750
rect 6320 3710 6340 3750
rect 6260 3690 6340 3710
rect 6390 3750 6450 3770
rect 6390 3710 6400 3750
rect 6440 3710 6450 3750
rect 6390 3690 6450 3710
rect 6630 3750 6690 3770
rect 6630 3710 6640 3750
rect 6680 3710 6690 3750
rect 6630 3690 6690 3710
rect 6870 3750 6930 3770
rect 6870 3710 6880 3750
rect 6920 3710 6930 3750
rect 6870 3690 6930 3710
rect 7110 3750 7170 3770
rect 7110 3710 7120 3750
rect 7160 3710 7170 3750
rect 7110 3690 7170 3710
rect 7350 3750 7410 3770
rect 7350 3710 7360 3750
rect 7400 3710 7410 3750
rect 7350 3690 7410 3710
rect 7600 3650 7640 3770
rect 6160 3610 6820 3650
rect 6980 3610 7640 3650
rect 8720 3810 8740 3890
rect 8790 3870 8850 3890
rect 8790 3830 8800 3870
rect 8840 3830 8850 3870
rect 8790 3810 8850 3830
rect 8910 3870 8970 3890
rect 8910 3830 8920 3870
rect 8960 3830 8970 3870
rect 8910 3810 8970 3830
rect 9030 3870 9090 3890
rect 9030 3830 9040 3870
rect 9080 3830 9090 3870
rect 9030 3810 9090 3830
rect 9150 3870 9210 3890
rect 9150 3830 9160 3870
rect 9200 3830 9210 3870
rect 9150 3810 9210 3830
rect 9270 3870 9330 3890
rect 9270 3830 9280 3870
rect 9320 3830 9330 3870
rect 9270 3810 9330 3830
rect 9390 3870 9450 3890
rect 9390 3830 9400 3870
rect 9440 3830 9450 3870
rect 9390 3810 9450 3830
rect 9510 3870 9570 3890
rect 9510 3830 9520 3870
rect 9560 3830 9570 3870
rect 9510 3810 9570 3830
rect 9630 3870 9690 3890
rect 9630 3830 9640 3870
rect 9680 3830 9690 3870
rect 9630 3810 9690 3830
rect 9750 3870 9810 3890
rect 9750 3830 9760 3870
rect 9800 3830 9810 3870
rect 9750 3810 9810 3830
rect 9870 3870 9930 3890
rect 9870 3830 9880 3870
rect 9920 3830 9930 3870
rect 9870 3810 9930 3830
rect 9990 3870 10050 3890
rect 9990 3830 10000 3870
rect 10040 3830 10050 3870
rect 9990 3810 10050 3830
rect 8920 3770 8960 3810
rect 9160 3770 9200 3810
rect 9400 3770 9440 3810
rect 9640 3770 9680 3810
rect 9880 3770 9920 3810
rect 8680 3650 8720 3770
rect 8910 3750 8970 3770
rect 8910 3710 8920 3750
rect 8960 3710 8970 3750
rect 8910 3690 8970 3710
rect 9150 3750 9210 3770
rect 9150 3710 9160 3750
rect 9200 3710 9210 3750
rect 9150 3690 9210 3710
rect 9390 3750 9450 3770
rect 9390 3710 9400 3750
rect 9440 3710 9450 3750
rect 9390 3690 9450 3710
rect 9630 3750 9690 3770
rect 9630 3710 9640 3750
rect 9680 3710 9690 3750
rect 9630 3690 9690 3710
rect 9870 3750 9930 3770
rect 9870 3710 9880 3750
rect 9920 3710 9930 3750
rect 9870 3690 9930 3710
rect 9980 3750 10060 3770
rect 9980 3710 10000 3750
rect 10040 3710 10060 3750
rect 9980 3690 10060 3710
rect 10120 3650 10160 3770
rect 8680 3610 10160 3650
rect 9860 3570 9940 3610
rect 250 2670 4270 2750
rect 1300 1380 1550 2670
rect 2660 1380 2910 2670
rect 4020 1390 4270 2670
rect 5680 3490 6820 3530
rect 6980 3490 8120 3530
rect 5680 3180 5720 3490
rect 5960 3430 6040 3450
rect 5780 3400 5860 3420
rect 5780 3360 5800 3400
rect 5840 3360 5860 3400
rect 5960 3390 5980 3430
rect 6020 3390 6040 3430
rect 5960 3370 6040 3390
rect 6200 3430 6280 3450
rect 6200 3390 6220 3430
rect 6260 3390 6280 3430
rect 6200 3370 6280 3390
rect 6440 3430 6520 3450
rect 6440 3390 6460 3430
rect 6500 3390 6520 3430
rect 6440 3370 6520 3390
rect 6680 3430 6760 3450
rect 6680 3390 6700 3430
rect 6740 3390 6760 3430
rect 6680 3370 6760 3390
rect 7160 3430 7240 3450
rect 7160 3390 7180 3430
rect 7220 3390 7240 3430
rect 7160 3370 7240 3390
rect 7400 3430 7480 3450
rect 7400 3390 7420 3430
rect 7460 3390 7480 3430
rect 7400 3370 7480 3390
rect 7640 3430 7720 3450
rect 7640 3390 7660 3430
rect 7700 3390 7720 3430
rect 7640 3370 7720 3390
rect 7940 3400 8020 3420
rect 5780 3340 5860 3360
rect 7940 3360 7960 3400
rect 8000 3360 8020 3400
rect 7940 3340 8020 3360
rect 5680 2700 5720 3020
rect 5790 3320 5850 3340
rect 5790 3280 5800 3320
rect 5840 3280 5850 3320
rect 5790 3220 5850 3280
rect 5790 3180 5800 3220
rect 5840 3180 5850 3220
rect 5790 3120 5850 3180
rect 5790 3080 5800 3120
rect 5840 3080 5850 3120
rect 5790 3020 5850 3080
rect 5790 2980 5800 3020
rect 5840 2980 5850 3020
rect 5790 2920 5850 2980
rect 5790 2880 5800 2920
rect 5840 2880 5850 2920
rect 5790 2860 5850 2880
rect 6870 3320 6930 3340
rect 6870 3280 6880 3320
rect 6920 3280 6930 3320
rect 6870 3220 6930 3280
rect 6870 3180 6880 3220
rect 6920 3180 6930 3220
rect 6870 3120 6930 3180
rect 6870 3080 6880 3120
rect 6920 3080 6930 3120
rect 6870 3020 6930 3080
rect 6870 2980 6880 3020
rect 6920 2980 6930 3020
rect 6870 2920 6930 2980
rect 6870 2880 6880 2920
rect 6920 2880 6930 2920
rect 6870 2860 6930 2880
rect 7950 3320 8010 3340
rect 7950 3280 7960 3320
rect 8000 3280 8010 3320
rect 7950 3220 8010 3280
rect 7950 3180 7960 3220
rect 8000 3180 8010 3220
rect 7950 3120 8010 3180
rect 7950 3080 7960 3120
rect 8000 3080 8010 3120
rect 7950 3020 8010 3080
rect 7950 2980 7960 3020
rect 8000 2980 8010 3020
rect 7950 2920 8010 2980
rect 7950 2880 7960 2920
rect 8000 2880 8010 2920
rect 7950 2860 8010 2880
rect 8080 3180 8120 3490
rect 6880 2820 6920 2860
rect 6860 2800 6940 2820
rect 6860 2760 6880 2800
rect 6920 2760 6940 2800
rect 6860 2740 6940 2760
rect 6880 2700 6920 2740
rect 8080 2700 8120 3020
rect 5680 2660 6820 2700
rect 6980 2660 8120 2700
rect 8200 3490 9340 3530
rect 9500 3490 10640 3530
rect 8200 3180 8240 3490
rect 8600 3430 8680 3450
rect 8300 3400 8380 3420
rect 8300 3360 8320 3400
rect 8360 3360 8380 3400
rect 8600 3390 8620 3430
rect 8660 3390 8680 3430
rect 8600 3370 8680 3390
rect 8840 3430 8920 3450
rect 8840 3390 8860 3430
rect 8900 3390 8920 3430
rect 8840 3370 8920 3390
rect 9080 3430 9160 3450
rect 9080 3390 9100 3430
rect 9140 3390 9160 3430
rect 9080 3370 9160 3390
rect 9560 3430 9640 3450
rect 9560 3390 9580 3430
rect 9620 3390 9640 3430
rect 9560 3370 9640 3390
rect 9800 3430 9880 3450
rect 9800 3390 9820 3430
rect 9860 3390 9880 3430
rect 9800 3370 9880 3390
rect 10040 3430 10120 3450
rect 10040 3390 10060 3430
rect 10100 3390 10120 3430
rect 10040 3370 10120 3390
rect 10280 3430 10360 3450
rect 10280 3390 10300 3430
rect 10340 3390 10360 3430
rect 10280 3370 10360 3390
rect 10460 3400 10540 3420
rect 8300 3340 8380 3360
rect 10460 3360 10480 3400
rect 10520 3360 10540 3400
rect 10460 3340 10540 3360
rect 8200 2700 8240 3020
rect 8310 3320 8370 3340
rect 8310 3280 8320 3320
rect 8360 3280 8370 3320
rect 8310 3220 8370 3280
rect 8310 3180 8320 3220
rect 8360 3180 8370 3220
rect 8310 3120 8370 3180
rect 8310 3080 8320 3120
rect 8360 3080 8370 3120
rect 8310 3020 8370 3080
rect 8310 2980 8320 3020
rect 8360 2980 8370 3020
rect 8310 2920 8370 2980
rect 8310 2880 8320 2920
rect 8360 2880 8370 2920
rect 8310 2860 8370 2880
rect 9390 3320 9450 3340
rect 9390 3280 9400 3320
rect 9440 3280 9450 3320
rect 9390 3220 9450 3280
rect 9390 3180 9400 3220
rect 9440 3180 9450 3220
rect 9390 3120 9450 3180
rect 9390 3080 9400 3120
rect 9440 3080 9450 3120
rect 9390 3020 9450 3080
rect 9390 2980 9400 3020
rect 9440 2980 9450 3020
rect 9390 2920 9450 2980
rect 9390 2880 9400 2920
rect 9440 2880 9450 2920
rect 9390 2860 9450 2880
rect 10470 3320 10530 3340
rect 10470 3280 10480 3320
rect 10520 3280 10530 3320
rect 10470 3220 10530 3280
rect 10470 3180 10480 3220
rect 10520 3180 10530 3220
rect 10470 3120 10530 3180
rect 10470 3080 10480 3120
rect 10520 3080 10530 3120
rect 10470 3020 10530 3080
rect 10470 2980 10480 3020
rect 10520 2980 10530 3020
rect 10470 2920 10530 2980
rect 10470 2880 10480 2920
rect 10520 2880 10530 2920
rect 10470 2860 10530 2880
rect 10600 3180 10640 3490
rect 9400 2820 9440 2860
rect 9380 2800 9460 2820
rect 9380 2760 9400 2800
rect 9440 2760 9460 2800
rect 9380 2740 9460 2760
rect 9400 2700 9440 2740
rect 10600 2700 10640 3020
rect 8200 2660 9340 2700
rect 9500 2660 10640 2700
rect 5880 2560 8080 2600
rect 8240 2560 10430 2600
rect 5880 2390 5920 2560
rect 6040 2500 6120 2520
rect 6040 2460 6060 2500
rect 6100 2460 6120 2500
rect 6040 2440 6120 2460
rect 6200 2500 6280 2520
rect 6200 2460 6220 2500
rect 6260 2460 6280 2500
rect 6200 2440 6280 2460
rect 6360 2500 6440 2520
rect 6360 2460 6380 2500
rect 6420 2460 6440 2500
rect 6360 2440 6440 2460
rect 6520 2500 6600 2520
rect 6520 2460 6540 2500
rect 6580 2460 6600 2500
rect 6520 2440 6600 2460
rect 6680 2500 6760 2520
rect 6680 2460 6700 2500
rect 6740 2460 6760 2500
rect 6680 2440 6760 2460
rect 6840 2500 6920 2520
rect 6840 2460 6860 2500
rect 6900 2460 6920 2500
rect 6840 2440 6920 2460
rect 7000 2500 7080 2520
rect 7000 2460 7020 2500
rect 7060 2460 7080 2500
rect 7000 2440 7080 2460
rect 7160 2500 7240 2520
rect 7160 2460 7180 2500
rect 7220 2460 7240 2500
rect 7160 2440 7240 2460
rect 7320 2500 7400 2520
rect 7320 2460 7340 2500
rect 7380 2460 7400 2500
rect 7320 2440 7400 2460
rect 7480 2500 7560 2520
rect 7480 2460 7500 2500
rect 7540 2460 7560 2500
rect 7480 2440 7560 2460
rect 7640 2500 7720 2520
rect 7640 2460 7660 2500
rect 7700 2460 7720 2500
rect 7640 2440 7720 2460
rect 7800 2500 7880 2520
rect 7800 2460 7820 2500
rect 7860 2460 7880 2500
rect 7800 2440 7880 2460
rect 7960 2500 8040 2520
rect 7960 2460 7980 2500
rect 8020 2460 8040 2500
rect 7960 2440 8040 2460
rect 8120 2500 8200 2520
rect 8120 2460 8140 2500
rect 8180 2460 8200 2500
rect 8120 2440 8200 2460
rect 8280 2500 8360 2520
rect 8280 2460 8300 2500
rect 8340 2460 8360 2500
rect 8280 2440 8360 2460
rect 8440 2500 8520 2520
rect 8440 2460 8460 2500
rect 8500 2460 8520 2500
rect 8440 2440 8520 2460
rect 8600 2500 8680 2520
rect 8600 2460 8620 2500
rect 8660 2460 8680 2500
rect 8600 2440 8680 2460
rect 8760 2500 8840 2520
rect 8760 2460 8780 2500
rect 8820 2460 8840 2500
rect 8760 2440 8840 2460
rect 8920 2500 9000 2520
rect 8920 2460 8940 2500
rect 8980 2460 9000 2500
rect 8920 2440 9000 2460
rect 9080 2500 9160 2520
rect 9080 2460 9100 2500
rect 9140 2460 9160 2500
rect 9080 2440 9160 2460
rect 9240 2500 9320 2520
rect 9240 2460 9260 2500
rect 9300 2460 9320 2500
rect 9240 2440 9320 2460
rect 9400 2500 9480 2520
rect 9400 2460 9420 2500
rect 9460 2460 9480 2500
rect 9400 2440 9480 2460
rect 9560 2500 9640 2520
rect 9560 2460 9580 2500
rect 9620 2460 9640 2500
rect 9560 2440 9640 2460
rect 9720 2500 9800 2520
rect 9720 2460 9740 2500
rect 9780 2460 9800 2500
rect 9720 2440 9800 2460
rect 9880 2500 9960 2520
rect 9880 2460 9900 2500
rect 9940 2460 9960 2500
rect 9880 2440 9960 2460
rect 10040 2500 10120 2520
rect 10040 2460 10060 2500
rect 10100 2460 10120 2500
rect 10040 2440 10120 2460
rect 6060 2400 6100 2440
rect 8140 2400 8180 2440
rect 6050 2380 6110 2400
rect 6050 2350 6060 2380
rect 5960 2340 6060 2350
rect 6100 2340 6110 2380
rect 5960 2330 6110 2340
rect 5960 2290 5980 2330
rect 6020 2290 6110 2330
rect 5960 2280 6110 2290
rect 5960 2270 6060 2280
rect 5880 2150 5920 2230
rect 6050 2240 6060 2270
rect 6100 2240 6110 2280
rect 6050 2220 6110 2240
rect 8130 2380 8190 2400
rect 8130 2340 8140 2380
rect 8180 2340 8190 2380
rect 8130 2280 8190 2340
rect 8130 2240 8140 2280
rect 8180 2240 8190 2280
rect 8130 2220 8190 2240
rect 10210 2380 10270 2400
rect 10210 2340 10220 2380
rect 10260 2350 10270 2380
rect 10390 2390 10430 2560
rect 10260 2340 10350 2350
rect 10210 2330 10350 2340
rect 10210 2290 10290 2330
rect 10330 2290 10350 2330
rect 10210 2280 10350 2290
rect 10210 2240 10220 2280
rect 10260 2270 10350 2280
rect 10260 2240 10270 2270
rect 10210 2220 10270 2240
rect 10390 2150 10430 2230
rect 5880 2110 8080 2150
rect 8240 2110 10430 2150
rect 5330 2010 6110 2050
rect 6270 2010 7050 2050
rect 5330 1840 5370 2010
rect 5790 1950 5870 1970
rect 5790 1910 5810 1950
rect 5850 1910 5870 1950
rect 5790 1890 5870 1910
rect 6150 1950 6230 1970
rect 6150 1910 6170 1950
rect 6210 1910 6230 1950
rect 6150 1890 6230 1910
rect 6330 1950 6410 1970
rect 6330 1910 6350 1950
rect 6390 1910 6410 1950
rect 6330 1890 6410 1910
rect 6510 1950 6590 1970
rect 6510 1910 6530 1950
rect 6570 1910 6590 1950
rect 6510 1890 6590 1910
rect 5810 1850 5850 1890
rect 6170 1850 6210 1890
rect 6530 1850 6570 1890
rect 5330 1510 5370 1680
rect 5440 1830 5500 1850
rect 5440 1790 5450 1830
rect 5490 1790 5500 1830
rect 5440 1730 5500 1790
rect 5440 1690 5450 1730
rect 5490 1690 5500 1730
rect 5440 1610 5500 1690
rect 5620 1830 5680 1850
rect 5620 1790 5630 1830
rect 5670 1790 5680 1830
rect 5620 1730 5680 1790
rect 5620 1690 5630 1730
rect 5670 1690 5680 1730
rect 5620 1670 5680 1690
rect 5800 1830 5860 1850
rect 5800 1790 5810 1830
rect 5850 1790 5860 1830
rect 5800 1730 5860 1790
rect 5800 1690 5810 1730
rect 5850 1690 5860 1730
rect 5800 1670 5860 1690
rect 5980 1830 6040 1850
rect 5980 1790 5990 1830
rect 6030 1790 6040 1830
rect 5980 1730 6040 1790
rect 5980 1690 5990 1730
rect 6030 1690 6040 1730
rect 5980 1670 6040 1690
rect 6160 1830 6220 1850
rect 6160 1790 6170 1830
rect 6210 1790 6220 1830
rect 6160 1730 6220 1790
rect 6160 1690 6170 1730
rect 6210 1690 6220 1730
rect 6160 1670 6220 1690
rect 6340 1830 6400 1850
rect 6340 1790 6350 1830
rect 6390 1790 6400 1830
rect 6340 1730 6400 1790
rect 6340 1690 6350 1730
rect 6390 1690 6400 1730
rect 6340 1670 6400 1690
rect 6520 1830 6580 1850
rect 6520 1790 6530 1830
rect 6570 1790 6580 1830
rect 6520 1730 6580 1790
rect 6520 1690 6530 1730
rect 6570 1690 6580 1730
rect 6520 1670 6580 1690
rect 6700 1830 6760 1850
rect 6700 1790 6710 1830
rect 6750 1790 6760 1830
rect 6700 1730 6760 1790
rect 6700 1690 6710 1730
rect 6750 1690 6760 1730
rect 6700 1670 6760 1690
rect 6880 1830 6940 1850
rect 6880 1790 6890 1830
rect 6930 1790 6940 1830
rect 6880 1730 6940 1790
rect 6880 1690 6890 1730
rect 6930 1690 6940 1730
rect 5630 1630 5670 1670
rect 5990 1630 6030 1670
rect 6350 1630 6390 1670
rect 6710 1630 6750 1670
rect 5440 1570 5450 1610
rect 5490 1570 5500 1610
rect 5440 1550 5500 1570
rect 5610 1610 5690 1630
rect 5610 1570 5630 1610
rect 5670 1570 5690 1610
rect 5610 1550 5690 1570
rect 5970 1610 6050 1630
rect 5970 1570 5990 1610
rect 6030 1570 6050 1610
rect 5970 1550 6050 1570
rect 6330 1610 6410 1630
rect 6330 1570 6350 1610
rect 6390 1570 6410 1610
rect 6330 1550 6410 1570
rect 6690 1610 6770 1630
rect 6690 1570 6710 1610
rect 6750 1570 6770 1610
rect 6690 1550 6770 1570
rect 6880 1610 6940 1690
rect 6880 1570 6890 1610
rect 6930 1570 6940 1610
rect 6880 1550 6940 1570
rect 7010 1840 7050 2010
rect 5450 1510 5490 1550
rect 6890 1510 6930 1550
rect 7010 1510 7050 1680
rect 5330 1470 6110 1510
rect 6270 1470 7050 1510
rect 7120 2010 8080 2050
rect 8240 2010 9200 2050
rect 7120 1840 7160 2010
rect 7580 1950 7660 1970
rect 7580 1910 7600 1950
rect 7640 1910 7660 1950
rect 7580 1890 7660 1910
rect 7940 1950 8020 1970
rect 7940 1910 7960 1950
rect 8000 1910 8020 1950
rect 7940 1890 8020 1910
rect 8120 1950 8200 1970
rect 8120 1910 8140 1950
rect 8180 1910 8200 1950
rect 8120 1890 8200 1910
rect 8300 1950 8380 1970
rect 8300 1910 8320 1950
rect 8360 1910 8380 1950
rect 8300 1890 8380 1910
rect 8660 1950 8740 1970
rect 8660 1910 8680 1950
rect 8720 1910 8740 1950
rect 8660 1890 8740 1910
rect 7600 1850 7640 1890
rect 7960 1850 8000 1890
rect 8320 1850 8360 1890
rect 8680 1850 8720 1890
rect 7120 1510 7160 1680
rect 7230 1830 7290 1850
rect 7230 1790 7240 1830
rect 7280 1790 7290 1830
rect 7230 1730 7290 1790
rect 7230 1690 7240 1730
rect 7280 1690 7290 1730
rect 7230 1610 7290 1690
rect 7230 1570 7240 1610
rect 7280 1570 7290 1610
rect 7410 1830 7470 1850
rect 7410 1790 7420 1830
rect 7460 1790 7470 1830
rect 7410 1730 7470 1790
rect 7410 1690 7420 1730
rect 7460 1690 7470 1730
rect 7410 1670 7470 1690
rect 7590 1830 7650 1850
rect 7590 1790 7600 1830
rect 7640 1790 7650 1830
rect 7590 1730 7650 1790
rect 7590 1690 7600 1730
rect 7640 1690 7650 1730
rect 7590 1670 7650 1690
rect 7770 1830 7830 1850
rect 7770 1790 7780 1830
rect 7820 1790 7830 1830
rect 7770 1730 7830 1790
rect 7770 1690 7780 1730
rect 7820 1690 7830 1730
rect 7770 1670 7830 1690
rect 7950 1830 8010 1850
rect 7950 1790 7960 1830
rect 8000 1790 8010 1830
rect 7950 1730 8010 1790
rect 7950 1690 7960 1730
rect 8000 1690 8010 1730
rect 7950 1670 8010 1690
rect 8130 1830 8190 1850
rect 8130 1790 8140 1830
rect 8180 1790 8190 1830
rect 8130 1730 8190 1790
rect 8130 1690 8140 1730
rect 8180 1690 8190 1730
rect 8130 1670 8190 1690
rect 8310 1830 8370 1850
rect 8310 1790 8320 1830
rect 8360 1790 8370 1830
rect 8310 1730 8370 1790
rect 8310 1690 8320 1730
rect 8360 1690 8370 1730
rect 8310 1670 8370 1690
rect 8490 1830 8550 1850
rect 8490 1790 8500 1830
rect 8540 1790 8550 1830
rect 8490 1730 8550 1790
rect 8490 1690 8500 1730
rect 8540 1690 8550 1730
rect 8490 1670 8550 1690
rect 8670 1830 8730 1850
rect 8670 1790 8680 1830
rect 8720 1790 8730 1830
rect 8670 1730 8730 1790
rect 8670 1690 8680 1730
rect 8720 1690 8730 1730
rect 8670 1670 8730 1690
rect 8850 1830 8910 1850
rect 8850 1790 8860 1830
rect 8900 1790 8910 1830
rect 8850 1730 8910 1790
rect 8850 1690 8860 1730
rect 8900 1690 8910 1730
rect 8850 1670 8910 1690
rect 9030 1830 9090 1850
rect 9030 1790 9040 1830
rect 9080 1790 9090 1830
rect 9030 1730 9090 1790
rect 9030 1690 9040 1730
rect 9080 1690 9090 1730
rect 7410 1610 7450 1670
rect 7780 1630 7820 1670
rect 8140 1630 8180 1670
rect 8500 1630 8540 1670
rect 8860 1630 8900 1670
rect 7490 1610 7570 1630
rect 7410 1570 7510 1610
rect 7550 1570 7570 1610
rect 7230 1550 7290 1570
rect 7490 1550 7570 1570
rect 7760 1610 7840 1630
rect 7760 1570 7780 1610
rect 7820 1570 7840 1610
rect 7760 1550 7840 1570
rect 8120 1610 8200 1630
rect 8120 1570 8140 1610
rect 8180 1570 8200 1610
rect 8120 1550 8200 1570
rect 8480 1610 8560 1630
rect 8480 1570 8500 1610
rect 8540 1570 8560 1610
rect 8480 1550 8560 1570
rect 8840 1610 8920 1630
rect 8840 1570 8860 1610
rect 8900 1570 8920 1610
rect 8840 1550 8920 1570
rect 9030 1610 9090 1690
rect 9030 1570 9040 1610
rect 9080 1570 9090 1610
rect 9030 1550 9090 1570
rect 9160 1840 9200 2010
rect 7240 1510 7280 1550
rect 9040 1510 9080 1550
rect 9160 1510 9200 1680
rect 7120 1470 8080 1510
rect 8240 1470 9200 1510
rect 9270 2010 10050 2050
rect 10210 2010 10990 2050
rect 9270 1840 9310 2010
rect 9730 1950 9810 1970
rect 9730 1910 9750 1950
rect 9790 1910 9810 1950
rect 9730 1890 9810 1910
rect 9910 1950 9990 1970
rect 9910 1910 9930 1950
rect 9970 1910 9990 1950
rect 9910 1890 9990 1910
rect 10090 1950 10170 1970
rect 10090 1910 10110 1950
rect 10150 1910 10170 1950
rect 10090 1890 10170 1910
rect 10450 1950 10530 1970
rect 10450 1910 10470 1950
rect 10510 1910 10530 1950
rect 10450 1890 10530 1910
rect 9750 1850 9790 1890
rect 10110 1850 10150 1890
rect 10470 1850 10510 1890
rect 9270 1510 9310 1680
rect 9380 1830 9440 1850
rect 9380 1790 9390 1830
rect 9430 1790 9440 1830
rect 9380 1730 9440 1790
rect 9380 1690 9390 1730
rect 9430 1690 9440 1730
rect 9380 1610 9440 1690
rect 9560 1830 9620 1850
rect 9560 1790 9570 1830
rect 9610 1790 9620 1830
rect 9560 1730 9620 1790
rect 9560 1690 9570 1730
rect 9610 1690 9620 1730
rect 9560 1670 9620 1690
rect 9740 1830 9800 1850
rect 9740 1790 9750 1830
rect 9790 1790 9800 1830
rect 9740 1730 9800 1790
rect 9740 1690 9750 1730
rect 9790 1690 9800 1730
rect 9740 1670 9800 1690
rect 9920 1830 9980 1850
rect 9920 1790 9930 1830
rect 9970 1790 9980 1830
rect 9920 1730 9980 1790
rect 9920 1690 9930 1730
rect 9970 1690 9980 1730
rect 9920 1670 9980 1690
rect 10100 1830 10160 1850
rect 10100 1790 10110 1830
rect 10150 1790 10160 1830
rect 10100 1730 10160 1790
rect 10100 1690 10110 1730
rect 10150 1690 10160 1730
rect 10100 1670 10160 1690
rect 10280 1830 10340 1850
rect 10280 1790 10290 1830
rect 10330 1790 10340 1830
rect 10280 1730 10340 1790
rect 10280 1690 10290 1730
rect 10330 1690 10340 1730
rect 10280 1670 10340 1690
rect 10460 1830 10520 1850
rect 10460 1790 10470 1830
rect 10510 1790 10520 1830
rect 10460 1730 10520 1790
rect 10460 1690 10470 1730
rect 10510 1690 10520 1730
rect 10460 1670 10520 1690
rect 10640 1830 10700 1850
rect 10640 1790 10650 1830
rect 10690 1790 10700 1830
rect 10640 1730 10700 1790
rect 10640 1690 10650 1730
rect 10690 1690 10700 1730
rect 10640 1670 10700 1690
rect 10820 1830 10880 1850
rect 10820 1790 10830 1830
rect 10870 1790 10880 1830
rect 10820 1730 10880 1790
rect 10820 1690 10830 1730
rect 10870 1690 10880 1730
rect 9570 1630 9610 1670
rect 9930 1630 9970 1670
rect 10290 1630 10330 1670
rect 10650 1630 10690 1670
rect 9380 1570 9390 1610
rect 9430 1570 9440 1610
rect 9380 1550 9440 1570
rect 9550 1610 9630 1630
rect 9550 1570 9570 1610
rect 9610 1570 9630 1610
rect 9550 1550 9630 1570
rect 9910 1610 9990 1630
rect 9910 1570 9930 1610
rect 9970 1570 9990 1610
rect 9910 1550 9990 1570
rect 10270 1610 10350 1630
rect 10270 1570 10290 1610
rect 10330 1570 10350 1610
rect 10270 1550 10350 1570
rect 10630 1610 10710 1630
rect 10630 1570 10650 1610
rect 10690 1570 10710 1610
rect 10630 1550 10710 1570
rect 10820 1610 10880 1690
rect 10820 1570 10830 1610
rect 10870 1570 10880 1610
rect 10820 1550 10880 1570
rect 10950 1840 10990 2010
rect 9390 1510 9430 1550
rect 10830 1510 10870 1550
rect 10950 1510 10990 1680
rect 9270 1470 10050 1510
rect 10210 1470 10990 1510
rect 5980 1450 6040 1470
rect 6700 1450 6760 1470
rect 9560 1450 9620 1470
rect 10280 1450 10340 1470
<< viali >>
rect 152 7120 202 7170
rect 152 7000 202 7050
rect 152 6590 202 6640
rect 152 6470 202 6520
rect 2722 6850 2772 6900
rect 2722 6730 2772 6780
rect 2390 6530 2410 6570
rect 2410 6530 2430 6570
rect 2600 6530 2620 6570
rect 2620 6530 2640 6570
rect 1210 6360 1250 6380
rect 1210 6340 1250 6360
rect 542 6060 592 6110
rect 1888 6060 1938 6110
rect 5360 7010 5400 7050
rect 5720 7010 5760 7050
rect 5900 7010 5940 7050
rect 6080 7010 6120 7050
rect 6260 7010 6300 7050
rect 6440 7010 6480 7050
rect 5540 6670 5580 6710
rect 5900 6670 5940 6710
rect 6260 6670 6300 6710
rect 7060 7010 7100 7050
rect 7420 7010 7460 7050
rect 7780 7010 7820 7050
rect 7960 7010 8000 7050
rect 8140 7010 8180 7050
rect 8320 7010 8360 7050
rect 8500 7010 8540 7050
rect 8860 7010 8900 7050
rect 9040 7010 9080 7050
rect 9220 7010 9260 7050
rect 7240 6670 7280 6710
rect 7600 6670 7640 6710
rect 7960 6670 8000 6710
rect 8320 6670 8360 6710
rect 8680 6670 8720 6710
rect 9040 6670 9080 6710
rect 9840 7010 9880 7050
rect 10200 7010 10240 7050
rect 10380 7010 10420 7050
rect 10560 7010 10600 7050
rect 10920 7010 10960 7050
rect 10020 6670 10060 6710
rect 10380 6670 10420 6710
rect 10740 6670 10780 6710
rect 4860 6370 4910 6420
rect 4860 6250 4910 6300
rect 5670 6020 5710 6040
rect 542 5640 592 5690
rect 1888 5640 1938 5690
rect 3052 5840 3102 5890
rect 4450 5840 4500 5890
rect 5670 6000 5710 6020
rect 5670 5880 5710 5920
rect 5540 5540 5580 5580
rect 5670 5540 5710 5580
rect 5800 5540 5840 5580
rect 6520 6080 6560 6120
rect 6880 6080 6920 6120
rect 7240 6080 7280 6120
rect 7600 6080 7640 6120
rect 7960 6080 8000 6120
rect 8320 6080 8360 6120
rect 8680 6080 8720 6120
rect 9040 6080 9080 6120
rect 9400 6080 9440 6120
rect 9760 6080 9800 6120
rect 10740 6020 10780 6040
rect 6700 5340 6740 5380
rect 7060 5340 7100 5380
rect 7420 5340 7460 5380
rect 7780 5340 7820 5380
rect 7960 5340 8000 5380
rect 8140 5340 8180 5380
rect 8500 5340 8540 5380
rect 8860 5340 8900 5380
rect 9220 5340 9260 5380
rect 9400 5340 9440 5380
rect 9580 5340 9620 5380
rect 10740 6000 10780 6020
rect 10740 5880 10780 5920
rect 10540 5540 10580 5580
rect 10740 5540 10780 5580
rect 10940 5540 10980 5580
rect 6620 4840 6660 4860
rect 6620 4820 6660 4840
rect 5540 4700 5580 4740
rect 5660 4700 5700 4740
rect 5900 4700 5940 4740
rect 6140 4700 6180 4740
rect 6260 4700 6300 4740
rect 6380 4700 6420 4740
rect 6620 4700 6660 4740
rect 6860 4700 6900 4740
rect 6980 4700 7020 4740
rect 7100 4700 7140 4740
rect 7340 4700 7380 4740
rect 7580 4700 7620 4740
rect 7700 4700 7740 4740
rect 5600 4360 5640 4400
rect 5780 4360 5820 4400
rect 6020 4360 6060 4400
rect 6260 4360 6300 4400
rect 6500 4360 6540 4400
rect 6740 4360 6780 4400
rect 6980 4360 7020 4400
rect 7220 4360 7260 4400
rect 7460 4360 7500 4400
rect 7640 4360 7680 4400
rect 8700 4820 8740 4860
rect 8940 4820 8980 4860
rect 9180 4820 9220 4860
rect 9420 4820 9460 4860
rect 9660 4840 9700 4860
rect 9660 4820 9700 4840
rect 9900 4820 9940 4860
rect 10140 4820 10180 4860
rect 10380 4820 10420 4860
rect 10620 4820 10660 4860
rect 8580 4700 8620 4740
rect 8700 4700 8740 4740
rect 8940 4700 8980 4740
rect 9180 4700 9220 4740
rect 9300 4700 9340 4740
rect 9420 4700 9460 4740
rect 9660 4700 9700 4740
rect 9900 4700 9940 4740
rect 10020 4700 10060 4740
rect 10140 4700 10180 4740
rect 10380 4700 10420 4740
rect 10620 4700 10660 4740
rect 10740 4700 10780 4740
rect 8640 4360 8680 4400
rect 8820 4360 8860 4400
rect 9060 4360 9100 4400
rect 9300 4360 9340 4400
rect 9540 4360 9580 4400
rect 9780 4360 9820 4400
rect 10020 4360 10060 4400
rect 10260 4360 10300 4400
rect 10500 4360 10540 4400
rect 10680 4360 10720 4400
rect -70 3390 -30 3430
rect 6400 4040 6440 4080
rect 6280 3950 6320 3990
rect 6520 3950 6560 3990
rect 6760 3950 6800 3990
rect 7000 3950 7040 3990
rect 7240 3950 7280 3990
rect 7480 3950 7520 3990
rect 9880 4040 9920 4080
rect 8800 3950 8840 3990
rect 9040 3950 9080 3990
rect 9280 3950 9320 3990
rect 9520 3950 9560 3990
rect 9760 3950 9800 3990
rect 10000 3950 10040 3990
rect 7600 3830 7640 3870
rect 8680 3830 8720 3870
rect 6280 3710 6320 3750
rect 6400 3710 6440 3750
rect 6640 3710 6680 3750
rect 6880 3710 6920 3750
rect 7120 3710 7160 3750
rect 7360 3710 7400 3750
rect 8920 3710 8960 3750
rect 9160 3710 9200 3750
rect 9400 3710 9440 3750
rect 9640 3710 9680 3750
rect 9880 3710 9920 3750
rect 10000 3710 10040 3750
rect 5800 3360 5840 3400
rect 5980 3390 6020 3430
rect 6220 3390 6260 3430
rect 6460 3390 6500 3430
rect 6700 3390 6740 3430
rect 7180 3390 7220 3430
rect 7420 3390 7460 3430
rect 7660 3390 7700 3430
rect 7960 3360 8000 3400
rect 6880 2760 6920 2800
rect 8320 3360 8360 3400
rect 8620 3390 8660 3430
rect 8860 3390 8900 3430
rect 9100 3390 9140 3430
rect 9580 3390 9620 3430
rect 9820 3390 9860 3430
rect 10060 3390 10100 3430
rect 10300 3390 10340 3430
rect 10480 3360 10520 3400
rect 9400 2760 9440 2800
rect 8140 2560 8180 2600
rect 6060 2460 6100 2500
rect 6220 2460 6260 2500
rect 6380 2460 6420 2500
rect 6540 2460 6580 2500
rect 6700 2460 6740 2500
rect 6860 2460 6900 2500
rect 7020 2460 7060 2500
rect 7180 2460 7220 2500
rect 7340 2460 7380 2500
rect 7500 2460 7540 2500
rect 7660 2460 7700 2500
rect 7820 2460 7860 2500
rect 7980 2460 8020 2500
rect 8140 2460 8180 2500
rect 8300 2460 8340 2500
rect 8460 2460 8500 2500
rect 8620 2460 8660 2500
rect 8780 2460 8820 2500
rect 8940 2460 8980 2500
rect 9100 2460 9140 2500
rect 9260 2460 9300 2500
rect 9420 2460 9460 2500
rect 9580 2460 9620 2500
rect 9740 2460 9780 2500
rect 9900 2460 9940 2500
rect 10060 2460 10100 2500
rect 5980 2290 6020 2330
rect 10290 2290 10330 2330
rect 5810 1910 5850 1950
rect 6170 1910 6210 1950
rect 6350 1910 6390 1950
rect 6530 1910 6570 1950
rect 5630 1570 5670 1610
rect 5990 1570 6030 1610
rect 6350 1570 6390 1610
rect 6710 1570 6750 1610
rect 7010 1740 7050 1780
rect 7600 1910 7640 1950
rect 7960 1910 8000 1950
rect 8140 1910 8180 1950
rect 8320 1910 8360 1950
rect 8680 1910 8720 1950
rect 7120 1740 7160 1780
rect 7510 1570 7550 1610
rect 7780 1570 7820 1610
rect 8140 1570 8180 1610
rect 8500 1570 8540 1610
rect 8860 1570 8900 1610
rect 9160 1740 9200 1780
rect 9750 1910 9790 1950
rect 9930 1910 9970 1950
rect 10110 1910 10150 1950
rect 10470 1910 10510 1950
rect 9270 1740 9310 1780
rect 9570 1570 9610 1610
rect 9930 1570 9970 1610
rect 10290 1570 10330 1610
rect 10650 1570 10690 1610
rect 10950 1740 10990 1780
<< metal1 >>
rect 2700 7750 2780 7760
rect 2700 7690 2710 7750
rect 2770 7690 2780 7750
rect 2700 7680 2780 7690
rect 8880 7690 8960 7700
rect -30 7590 50 7600
rect -30 7530 -20 7590
rect 40 7530 50 7590
rect -30 7520 50 7530
rect 1880 7590 1960 7600
rect 1880 7530 1890 7590
rect 1950 7530 1960 7590
rect 1880 7520 1960 7530
rect -120 7480 -40 7490
rect -120 7420 -110 7480
rect -50 7420 -40 7480
rect -120 7410 -40 7420
rect -100 6120 -60 7410
rect -120 6110 -40 6120
rect -120 6050 -110 6110
rect -50 6050 -40 6110
rect -120 6040 -40 6050
rect -10 5710 30 7520
rect 2510 7380 2590 7390
rect 2510 7320 2520 7380
rect 2580 7320 2590 7380
rect 2510 7310 2590 7320
rect 140 7280 220 7290
rect 140 7220 150 7280
rect 210 7220 220 7280
rect 140 7210 220 7220
rect 150 7180 200 7210
rect 132 7110 142 7180
rect 212 7110 222 7180
rect 132 6990 142 7060
rect 212 6990 222 7060
rect 2530 6760 2570 7310
rect 2720 6910 2760 7680
rect 8880 7630 8890 7690
rect 8950 7630 8960 7690
rect 8880 7620 8960 7630
rect 3270 7590 3370 7610
rect 3270 7530 3290 7590
rect 3350 7530 3370 7590
rect 5020 7600 5100 7610
rect 5020 7540 5030 7600
rect 5090 7540 5100 7600
rect 5020 7530 5100 7540
rect 9600 7590 9680 7600
rect 9600 7530 9610 7590
rect 9670 7530 9680 7590
rect 3270 7510 3370 7530
rect 2702 6840 2712 6910
rect 2782 6840 2792 6910
rect 2722 6790 2762 6840
rect 140 6750 220 6760
rect 140 6690 150 6750
rect 210 6690 220 6750
rect 140 6680 220 6690
rect 2510 6750 2590 6760
rect 2510 6690 2520 6750
rect 2580 6690 2590 6750
rect 2702 6720 2712 6790
rect 2782 6720 2792 6790
rect 2510 6680 2590 6690
rect 150 6650 200 6680
rect 132 6580 142 6650
rect 212 6580 222 6650
rect 2370 6580 2450 6590
rect 132 6460 142 6530
rect 212 6460 222 6530
rect 2370 6520 2380 6580
rect 2440 6520 2450 6580
rect 2370 6510 2450 6520
rect 2580 6580 2660 6590
rect 2580 6520 2590 6580
rect 2650 6520 2660 6580
rect 2580 6510 2660 6520
rect 1190 6390 1270 6400
rect 1190 6330 1200 6390
rect 1260 6330 1270 6390
rect 4840 6360 4850 6430
rect 4920 6360 4930 6430
rect 1190 6320 1270 6330
rect 4840 6310 4930 6320
rect 4840 6240 4850 6310
rect 4920 6240 4930 6310
rect 4840 6230 4930 6240
rect 522 6050 532 6120
rect 602 6050 612 6120
rect 1868 6050 1878 6120
rect 1948 6050 1958 6120
rect 2420 6110 2500 6120
rect 2420 6050 2430 6110
rect 2490 6050 2500 6110
rect 2420 6040 2500 6050
rect 2210 5900 2290 5910
rect 2210 5840 2220 5900
rect 2280 5840 2290 5900
rect 2210 5830 2290 5840
rect -30 5700 50 5710
rect -30 5640 -20 5700
rect 40 5640 50 5700
rect -30 5630 50 5640
rect 522 5630 532 5700
rect 602 5630 612 5700
rect 1868 5630 1878 5700
rect 1948 5630 1958 5700
rect 2230 5100 2270 5830
rect 2440 5610 2480 6040
rect 4860 5900 4900 6230
rect 3032 5830 3042 5900
rect 3112 5830 3122 5900
rect 4430 5830 4440 5900
rect 4510 5830 4520 5900
rect 4840 5890 4920 5900
rect 4840 5830 4850 5890
rect 4910 5830 4920 5890
rect 4840 5820 4920 5830
rect 2420 5600 2500 5610
rect 2420 5540 2430 5600
rect 2490 5540 2500 5600
rect 2420 5530 2500 5540
rect 4750 5600 4830 5610
rect 4750 5540 4760 5600
rect 4820 5540 4830 5600
rect 4750 5530 4830 5540
rect 4660 5280 4740 5290
rect 4660 5220 4670 5280
rect 4730 5220 4740 5280
rect 4660 5210 4740 5220
rect 4550 5190 4630 5200
rect 4550 5130 4560 5190
rect 4620 5130 4630 5190
rect 4550 5120 4630 5130
rect 550 4400 3970 5100
rect -220 3440 -140 3450
rect -220 3380 -210 3440
rect -150 3430 -140 3440
rect -90 3440 -10 3450
rect -90 3430 -80 3440
rect -150 3390 -80 3430
rect -150 3380 -140 3390
rect -220 3370 -140 3380
rect -90 3380 -80 3390
rect -20 3380 -10 3440
rect -90 3370 -10 3380
rect 550 2380 1250 4400
rect 1904 3420 2604 3740
rect 1904 3360 2540 3420
rect 2594 3360 2604 3420
rect 1904 3040 2604 3360
rect 3270 2380 3970 4400
rect 550 1680 3970 2380
rect 4570 2350 4610 5120
rect 4680 4100 4720 5210
rect 4770 5010 4810 5530
rect 4860 5400 4900 5820
rect 4930 5690 5010 5700
rect 4930 5630 4940 5690
rect 5000 5630 5010 5690
rect 4930 5620 5010 5630
rect 4840 5390 4920 5400
rect 4840 5330 4850 5390
rect 4910 5330 4920 5390
rect 4840 5320 4920 5330
rect 4750 5000 4830 5010
rect 4750 4940 4760 5000
rect 4820 4940 4830 5000
rect 4750 4930 4830 4940
rect 4660 4090 4740 4100
rect 4660 4030 4670 4090
rect 4730 4030 4740 4090
rect 4660 4020 4740 4030
rect 4680 3430 4720 4020
rect 4860 3770 4900 5320
rect 4950 4760 4990 5620
rect 4930 4750 5010 4760
rect 4930 4690 4940 4750
rect 5000 4690 5010 4750
rect 4930 4680 5010 4690
rect 5040 4300 5080 7530
rect 9600 7520 9680 7530
rect 10270 7590 10370 7610
rect 10270 7530 10290 7590
rect 10350 7530 10370 7590
rect 5380 7480 5460 7490
rect 5380 7420 5390 7480
rect 5450 7420 5460 7480
rect 5380 7410 5460 7420
rect 6770 7480 6870 7500
rect 6770 7420 6790 7480
rect 6850 7420 6870 7480
rect 6770 7400 6870 7420
rect 9510 7480 9590 7490
rect 9510 7420 9520 7480
rect 9580 7420 9590 7480
rect 9510 7410 9590 7420
rect 9020 7380 9100 7390
rect 9020 7320 9030 7380
rect 9090 7320 9100 7380
rect 9020 7310 9100 7320
rect 5110 7280 5190 7290
rect 5110 7220 5120 7280
rect 5180 7220 5190 7280
rect 5110 7210 5190 7220
rect 6240 7270 6320 7280
rect 6240 7210 6250 7270
rect 6310 7210 6320 7270
rect 5130 6520 5170 7210
rect 6240 7200 6320 7210
rect 5880 7180 5960 7190
rect 5880 7120 5890 7180
rect 5950 7120 5960 7180
rect 5880 7110 5960 7120
rect 5900 7070 5940 7110
rect 6260 7070 6300 7200
rect 7940 7180 8020 7190
rect 7940 7120 7950 7180
rect 8010 7120 8020 7180
rect 7940 7110 8020 7120
rect 8300 7180 8380 7190
rect 8300 7120 8310 7180
rect 8370 7120 8380 7180
rect 8300 7110 8380 7120
rect 7960 7070 8000 7110
rect 8320 7070 8360 7110
rect 9040 7070 9080 7310
rect 9420 7180 9500 7190
rect 9420 7120 9430 7180
rect 9490 7120 9500 7180
rect 9420 7110 9500 7120
rect 5340 7060 5420 7070
rect 5340 7000 5350 7060
rect 5410 7000 5420 7060
rect 5340 6990 5420 7000
rect 5700 7060 5780 7070
rect 5700 7000 5710 7060
rect 5770 7000 5780 7060
rect 5700 6990 5780 7000
rect 5880 7050 5960 7070
rect 5880 7010 5900 7050
rect 5940 7010 5960 7050
rect 5880 6990 5960 7010
rect 6060 7060 6140 7070
rect 6060 7000 6070 7060
rect 6130 7000 6140 7060
rect 6060 6990 6140 7000
rect 6240 7050 6320 7070
rect 6240 7010 6260 7050
rect 6300 7010 6320 7050
rect 6240 6990 6320 7010
rect 6420 7060 6500 7070
rect 6420 7000 6430 7060
rect 6490 7000 6500 7060
rect 6420 6990 6500 7000
rect 7040 7060 7120 7070
rect 7040 7000 7050 7060
rect 7110 7000 7120 7060
rect 7040 6990 7120 7000
rect 7400 7060 7480 7070
rect 7400 7000 7410 7060
rect 7470 7000 7480 7060
rect 7400 6990 7480 7000
rect 7760 7060 7840 7070
rect 7760 7000 7770 7060
rect 7830 7000 7840 7060
rect 7760 6990 7840 7000
rect 7940 7050 8020 7070
rect 7940 7010 7960 7050
rect 8000 7010 8020 7050
rect 7940 6990 8020 7010
rect 8120 7060 8200 7070
rect 8120 7000 8130 7060
rect 8190 7000 8200 7060
rect 8120 6990 8200 7000
rect 8300 7050 8380 7070
rect 8300 7010 8320 7050
rect 8360 7010 8380 7050
rect 8300 6990 8380 7010
rect 8480 7060 8560 7070
rect 8480 7000 8490 7060
rect 8550 7000 8560 7060
rect 8480 6990 8560 7000
rect 8840 7060 8920 7070
rect 8840 7000 8850 7060
rect 8910 7000 8920 7060
rect 8840 6990 8920 7000
rect 9020 7050 9100 7070
rect 9020 7010 9040 7050
rect 9080 7010 9100 7050
rect 9020 6990 9100 7010
rect 9200 7060 9280 7070
rect 9200 7000 9210 7060
rect 9270 7000 9280 7060
rect 9200 6990 9280 7000
rect 5520 6720 5600 6730
rect 5520 6660 5530 6720
rect 5590 6660 5600 6720
rect 5520 6650 5600 6660
rect 5880 6720 5960 6730
rect 5880 6660 5890 6720
rect 5950 6660 5960 6720
rect 5880 6650 5960 6660
rect 6240 6720 6320 6730
rect 6240 6660 6250 6720
rect 6310 6660 6320 6720
rect 6240 6650 6320 6660
rect 7220 6710 7300 6730
rect 7220 6670 7240 6710
rect 7280 6670 7300 6710
rect 7220 6650 7300 6670
rect 7580 6720 7660 6730
rect 7580 6660 7590 6720
rect 7650 6660 7660 6720
rect 7580 6650 7660 6660
rect 7940 6720 8020 6730
rect 7940 6660 7950 6720
rect 8010 6660 8020 6720
rect 7940 6650 8020 6660
rect 8300 6720 8380 6730
rect 8300 6660 8310 6720
rect 8370 6660 8380 6720
rect 8300 6650 8380 6660
rect 8660 6720 8740 6730
rect 8660 6660 8670 6720
rect 8730 6660 8740 6720
rect 8660 6650 8740 6660
rect 9020 6710 9100 6730
rect 9020 6670 9040 6710
rect 9080 6670 9100 6710
rect 9020 6650 9100 6670
rect 5110 6510 5190 6520
rect 5110 6450 5120 6510
rect 5180 6450 5190 6510
rect 5110 6440 5190 6450
rect 5220 6510 5300 6520
rect 5220 6450 5230 6510
rect 5290 6450 5300 6510
rect 5220 6440 5300 6450
rect 5110 6330 5190 6340
rect 5110 6270 5120 6330
rect 5180 6270 5190 6330
rect 5110 6260 5190 6270
rect 5020 4290 5100 4300
rect 5020 4230 5030 4290
rect 5090 4230 5100 4290
rect 5020 4220 5100 4230
rect 4840 3760 4920 3770
rect 4840 3700 4850 3760
rect 4910 3700 4920 3760
rect 4840 3690 4920 3700
rect 4660 3420 4740 3430
rect 4660 3360 4670 3420
rect 4730 3360 4740 3420
rect 4660 3350 4740 3360
rect 4550 2340 4630 2350
rect 4550 2280 4560 2340
rect 4620 2280 4630 2340
rect 4550 2270 4630 2280
rect 5130 1430 5170 6260
rect 5240 5110 5280 6440
rect 6120 6420 6200 6430
rect 6120 6360 6130 6420
rect 6190 6360 6200 6420
rect 6120 6350 6200 6360
rect 5650 6050 5730 6060
rect 5650 5990 5660 6050
rect 5720 5990 5730 6050
rect 5650 5980 5730 5990
rect 6140 5940 6180 6350
rect 7240 6340 7280 6650
rect 7220 6330 7300 6340
rect 7220 6270 7230 6330
rect 7290 6270 7300 6330
rect 7220 6260 7300 6270
rect 8680 6260 8720 6650
rect 9040 6330 9080 6650
rect 9440 6640 9480 7110
rect 9420 6630 9500 6640
rect 9420 6570 9430 6630
rect 9490 6570 9500 6630
rect 9420 6560 9500 6570
rect 9530 6530 9570 7410
rect 9510 6520 9590 6530
rect 9510 6460 9520 6520
rect 9580 6460 9590 6520
rect 9510 6450 9590 6460
rect 9620 6420 9660 7520
rect 10270 7510 10370 7530
rect 10360 7180 10440 7190
rect 10360 7120 10370 7180
rect 10430 7120 10440 7180
rect 10360 7110 10440 7120
rect 10380 7070 10420 7110
rect 9820 7060 9900 7070
rect 9820 7000 9830 7060
rect 9890 7000 9900 7060
rect 9820 6990 9900 7000
rect 10180 7060 10260 7070
rect 10180 7000 10190 7060
rect 10250 7000 10260 7060
rect 10180 6990 10260 7000
rect 10360 7050 10440 7070
rect 10360 7010 10380 7050
rect 10420 7010 10440 7050
rect 10360 6990 10440 7010
rect 10540 7060 10620 7070
rect 10540 7000 10550 7060
rect 10610 7000 10620 7060
rect 10540 6990 10620 7000
rect 10900 7060 10980 7070
rect 10900 7000 10910 7060
rect 10970 7000 10980 7060
rect 10900 6990 10980 7000
rect 10000 6720 10080 6730
rect 10000 6660 10010 6720
rect 10070 6660 10080 6720
rect 10000 6650 10080 6660
rect 10360 6720 10440 6730
rect 10360 6660 10370 6720
rect 10430 6660 10440 6720
rect 10360 6650 10440 6660
rect 10720 6720 10800 6730
rect 10720 6660 10730 6720
rect 10790 6660 10800 6720
rect 10720 6650 10800 6660
rect 9940 6610 10020 6620
rect 9940 6550 9950 6610
rect 10010 6550 10020 6610
rect 9940 6540 10020 6550
rect 9600 6410 9680 6420
rect 9600 6350 9610 6410
rect 9670 6350 9680 6410
rect 9600 6340 9680 6350
rect 9020 6320 9100 6330
rect 9020 6260 9030 6320
rect 9090 6260 9100 6320
rect 8660 6250 8740 6260
rect 9020 6250 9100 6260
rect 8660 6190 8670 6250
rect 8730 6190 8740 6250
rect 8660 6180 8740 6190
rect 6500 6130 6580 6140
rect 6500 6070 6510 6130
rect 6570 6070 6580 6130
rect 6500 6060 6580 6070
rect 6860 6130 6940 6140
rect 6860 6070 6870 6130
rect 6930 6070 6940 6130
rect 6860 6060 6940 6070
rect 7220 6130 7300 6140
rect 7220 6070 7230 6130
rect 7290 6070 7300 6130
rect 7220 6060 7300 6070
rect 7580 6130 7660 6140
rect 7580 6070 7590 6130
rect 7650 6070 7660 6130
rect 7580 6060 7660 6070
rect 7940 6130 8020 6140
rect 7940 6070 7950 6130
rect 8010 6070 8020 6130
rect 7940 6060 8020 6070
rect 8300 6130 8380 6140
rect 8300 6070 8310 6130
rect 8370 6070 8380 6130
rect 8300 6060 8380 6070
rect 8660 6130 8740 6140
rect 8660 6070 8670 6130
rect 8730 6070 8740 6130
rect 8660 6060 8740 6070
rect 9020 6130 9100 6140
rect 9020 6070 9030 6130
rect 9090 6070 9100 6130
rect 9020 6060 9100 6070
rect 9380 6130 9460 6140
rect 9380 6070 9390 6130
rect 9450 6070 9460 6130
rect 9380 6060 9460 6070
rect 9740 6130 9820 6140
rect 9740 6070 9750 6130
rect 9810 6070 9820 6130
rect 9740 6060 9820 6070
rect 5650 5930 5730 5940
rect 5650 5870 5660 5930
rect 5720 5870 5730 5930
rect 5650 5860 5730 5870
rect 6120 5930 6200 5940
rect 6120 5870 6130 5930
rect 6190 5870 6200 5930
rect 6120 5860 6200 5870
rect 5520 5590 5600 5600
rect 5520 5530 5530 5590
rect 5590 5530 5600 5590
rect 5520 5520 5600 5530
rect 5650 5580 5730 5600
rect 5650 5540 5670 5580
rect 5710 5540 5730 5580
rect 5650 5520 5730 5540
rect 5780 5590 5860 5600
rect 5780 5530 5790 5590
rect 5850 5530 5860 5590
rect 5780 5520 5860 5530
rect 5670 5200 5710 5520
rect 6140 5290 6180 5860
rect 6240 5590 6320 5600
rect 6240 5530 6250 5590
rect 6310 5530 6320 5590
rect 6240 5520 6320 5530
rect 6120 5280 6200 5290
rect 6120 5220 6130 5280
rect 6190 5220 6200 5280
rect 6120 5210 6200 5220
rect 5650 5190 5730 5200
rect 5650 5130 5660 5190
rect 5720 5130 5730 5190
rect 5650 5120 5730 5130
rect 5220 5100 5300 5110
rect 5220 5040 5230 5100
rect 5290 5040 5300 5100
rect 5220 5030 5300 5040
rect 5640 4870 5720 4880
rect 5640 4810 5650 4870
rect 5710 4810 5720 4870
rect 5640 4800 5720 4810
rect 5880 4870 5960 4880
rect 5880 4810 5890 4870
rect 5950 4810 5960 4870
rect 5880 4800 5960 4810
rect 6120 4870 6200 4880
rect 6120 4810 6130 4870
rect 6190 4810 6200 4870
rect 6120 4800 6200 4810
rect 5660 4760 5700 4800
rect 5900 4760 5940 4800
rect 6140 4760 6180 4800
rect 6260 4760 6300 5520
rect 6680 5380 6760 5400
rect 6680 5340 6700 5380
rect 6740 5340 6760 5380
rect 6680 5320 6760 5340
rect 7040 5380 7120 5400
rect 7040 5340 7060 5380
rect 7100 5340 7120 5380
rect 7040 5320 7120 5340
rect 7400 5380 7480 5400
rect 7400 5340 7420 5380
rect 7460 5340 7480 5380
rect 7400 5320 7480 5340
rect 7760 5390 7840 5400
rect 7760 5330 7770 5390
rect 7830 5330 7840 5390
rect 7760 5320 7840 5330
rect 7940 5380 8020 5400
rect 7940 5340 7960 5380
rect 8000 5340 8020 5380
rect 7940 5320 8020 5340
rect 8120 5380 8200 5400
rect 8120 5340 8140 5380
rect 8180 5340 8200 5380
rect 8120 5320 8200 5340
rect 8480 5390 8560 5400
rect 8480 5330 8490 5390
rect 8550 5330 8560 5390
rect 8480 5320 8560 5330
rect 8840 5380 8920 5400
rect 8840 5340 8860 5380
rect 8900 5340 8920 5380
rect 8840 5320 8920 5340
rect 9200 5380 9280 5400
rect 9200 5340 9220 5380
rect 9260 5340 9280 5380
rect 9200 5320 9280 5340
rect 9380 5380 9460 5400
rect 9380 5340 9400 5380
rect 9440 5340 9460 5380
rect 9380 5320 9460 5340
rect 9560 5380 9640 5400
rect 9560 5340 9580 5380
rect 9620 5340 9640 5380
rect 9560 5320 9640 5340
rect 6700 5110 6740 5320
rect 7060 5200 7100 5320
rect 7420 5290 7460 5320
rect 7400 5280 7480 5290
rect 7400 5220 7410 5280
rect 7470 5220 7480 5280
rect 7400 5210 7480 5220
rect 7040 5190 7120 5200
rect 7040 5130 7050 5190
rect 7110 5130 7120 5190
rect 7040 5120 7120 5130
rect 6680 5100 6760 5110
rect 6680 5040 6690 5100
rect 6750 5040 6760 5100
rect 6680 5030 6760 5040
rect 6360 4870 6440 4880
rect 6360 4810 6370 4870
rect 6430 4810 6440 4870
rect 6360 4800 6440 4810
rect 6600 4870 6680 4880
rect 6600 4810 6610 4870
rect 6670 4810 6680 4870
rect 6600 4800 6680 4810
rect 6840 4870 6920 4880
rect 6840 4810 6850 4870
rect 6910 4810 6920 4870
rect 6840 4800 6920 4810
rect 7080 4870 7160 4880
rect 7080 4810 7090 4870
rect 7150 4810 7160 4870
rect 7080 4800 7160 4810
rect 7320 4870 7400 4880
rect 7320 4810 7330 4870
rect 7390 4810 7400 4870
rect 7320 4800 7400 4810
rect 7560 4870 7640 4880
rect 7560 4810 7570 4870
rect 7630 4810 7640 4870
rect 7560 4800 7640 4810
rect 6380 4760 6420 4800
rect 6620 4760 6660 4800
rect 6860 4760 6900 4800
rect 7100 4760 7140 4800
rect 7340 4760 7380 4800
rect 7580 4760 7620 4800
rect 7960 4760 8000 5320
rect 8140 5110 8180 5320
rect 8860 5290 8900 5320
rect 8840 5280 8920 5290
rect 8840 5220 8850 5280
rect 8910 5220 8920 5280
rect 8840 5210 8920 5220
rect 9220 5200 9260 5320
rect 9400 5200 9440 5320
rect 9200 5190 9280 5200
rect 9200 5130 9210 5190
rect 9270 5130 9280 5190
rect 9200 5120 9280 5130
rect 9380 5190 9460 5200
rect 9380 5130 9390 5190
rect 9450 5130 9460 5190
rect 9380 5120 9460 5130
rect 9580 5110 9620 5320
rect 8120 5100 8200 5110
rect 8120 5040 8130 5100
rect 8190 5040 8200 5100
rect 8120 5030 8200 5040
rect 9560 5100 9640 5110
rect 9560 5040 9570 5100
rect 9630 5040 9640 5100
rect 9560 5030 9640 5040
rect 9960 5010 10000 6540
rect 10120 6520 10200 6530
rect 10120 6460 10130 6520
rect 10190 6460 10200 6520
rect 10120 6450 10200 6460
rect 10030 6410 10110 6420
rect 10030 6350 10040 6410
rect 10100 6350 10110 6410
rect 10030 6340 10110 6350
rect 10050 5200 10090 6340
rect 10140 5310 10180 6450
rect 11230 6320 11310 6330
rect 11230 6260 11240 6320
rect 11300 6260 11310 6320
rect 11230 6250 11310 6260
rect 10720 6060 10800 6080
rect 10720 5990 10730 6060
rect 10790 5990 10800 6060
rect 10720 5980 10800 5990
rect 10740 5940 10780 5980
rect 10720 5930 10800 5940
rect 10720 5870 10730 5930
rect 10790 5870 10800 5930
rect 10720 5860 10800 5870
rect 10520 5590 10600 5600
rect 10520 5530 10530 5590
rect 10590 5530 10600 5590
rect 10520 5520 10600 5530
rect 10720 5580 10800 5600
rect 10720 5540 10740 5580
rect 10780 5540 10800 5580
rect 10720 5520 10800 5540
rect 10920 5590 11000 5600
rect 10920 5530 10930 5590
rect 10990 5530 11000 5590
rect 10920 5520 11000 5530
rect 10120 5300 10200 5310
rect 10120 5240 10130 5300
rect 10190 5240 10200 5300
rect 10120 5230 10200 5240
rect 10030 5190 10110 5200
rect 10030 5130 10040 5190
rect 10100 5130 10110 5190
rect 10030 5120 10110 5130
rect 10740 5010 10780 5520
rect 11050 5300 11130 5310
rect 11050 5240 11060 5300
rect 11120 5240 11130 5300
rect 11050 5230 11130 5240
rect 8560 5000 8640 5010
rect 8560 4940 8570 5000
rect 8630 4940 8640 5000
rect 8560 4930 8640 4940
rect 9940 5000 10020 5010
rect 9940 4940 9950 5000
rect 10010 4940 10020 5000
rect 9940 4930 10020 4940
rect 10720 5000 10800 5010
rect 10720 4940 10730 5000
rect 10790 4940 10800 5000
rect 10720 4930 10800 4940
rect 8580 4760 8620 4930
rect 8680 4870 8760 4880
rect 8680 4810 8690 4870
rect 8750 4810 8760 4870
rect 8680 4800 8760 4810
rect 8920 4870 9000 4880
rect 8920 4810 8930 4870
rect 8990 4810 9000 4870
rect 8920 4800 9000 4810
rect 9160 4870 9240 4880
rect 9160 4810 9170 4870
rect 9230 4810 9240 4870
rect 9160 4800 9240 4810
rect 9400 4870 9480 4880
rect 9400 4810 9410 4870
rect 9470 4810 9480 4870
rect 9400 4800 9480 4810
rect 9640 4870 9720 4880
rect 9640 4810 9650 4870
rect 9710 4810 9720 4870
rect 9640 4800 9720 4810
rect 9880 4870 9960 4880
rect 9880 4810 9890 4870
rect 9950 4810 9960 4870
rect 9880 4800 9960 4810
rect 10120 4870 10200 4880
rect 10120 4810 10130 4870
rect 10190 4810 10200 4870
rect 10120 4800 10200 4810
rect 10360 4870 10440 4880
rect 10360 4810 10370 4870
rect 10430 4810 10440 4870
rect 10360 4800 10440 4810
rect 10600 4870 10680 4880
rect 10600 4810 10610 4870
rect 10670 4810 10680 4870
rect 10600 4800 10680 4810
rect 8700 4760 8740 4800
rect 8940 4760 8980 4800
rect 9180 4760 9220 4800
rect 9420 4760 9460 4800
rect 9660 4760 9700 4800
rect 9900 4760 9940 4800
rect 10140 4760 10180 4800
rect 10380 4760 10420 4800
rect 10620 4760 10660 4800
rect 5520 4750 5600 4760
rect 5520 4690 5530 4750
rect 5590 4690 5600 4750
rect 5520 4680 5600 4690
rect 5650 4740 5710 4760
rect 5650 4700 5660 4740
rect 5700 4700 5710 4740
rect 5650 4680 5710 4700
rect 5890 4740 5950 4760
rect 5890 4700 5900 4740
rect 5940 4700 5950 4740
rect 5890 4680 5950 4700
rect 6130 4740 6190 4760
rect 6130 4700 6140 4740
rect 6180 4700 6190 4740
rect 6130 4680 6190 4700
rect 6240 4750 6320 4760
rect 6240 4690 6250 4750
rect 6310 4690 6320 4750
rect 6240 4680 6320 4690
rect 6370 4740 6430 4760
rect 6370 4700 6380 4740
rect 6420 4700 6430 4740
rect 6370 4680 6430 4700
rect 6610 4740 6670 4760
rect 6610 4700 6620 4740
rect 6660 4700 6670 4740
rect 6610 4680 6670 4700
rect 6850 4740 6910 4760
rect 6850 4700 6860 4740
rect 6900 4700 6910 4740
rect 6850 4680 6910 4700
rect 6960 4750 7040 4760
rect 6960 4690 6970 4750
rect 7030 4690 7040 4750
rect 6960 4680 7040 4690
rect 7090 4740 7150 4760
rect 7090 4700 7100 4740
rect 7140 4700 7150 4740
rect 7090 4680 7150 4700
rect 7330 4740 7390 4760
rect 7330 4700 7340 4740
rect 7380 4700 7390 4740
rect 7330 4680 7390 4700
rect 7570 4740 7630 4760
rect 7570 4700 7580 4740
rect 7620 4700 7630 4740
rect 7570 4680 7630 4700
rect 7680 4750 7760 4760
rect 7680 4690 7690 4750
rect 7750 4690 7760 4750
rect 7680 4680 7760 4690
rect 7940 4750 8020 4760
rect 7940 4690 7950 4750
rect 8010 4690 8020 4750
rect 7940 4680 8020 4690
rect 8300 4750 8380 4760
rect 8300 4690 8310 4750
rect 8370 4690 8380 4750
rect 8300 4680 8380 4690
rect 8560 4750 8640 4760
rect 8560 4690 8570 4750
rect 8630 4690 8640 4750
rect 8560 4680 8640 4690
rect 8690 4740 8750 4760
rect 8690 4700 8700 4740
rect 8740 4700 8750 4740
rect 8690 4680 8750 4700
rect 8930 4740 8990 4760
rect 8930 4700 8940 4740
rect 8980 4700 8990 4740
rect 8930 4680 8990 4700
rect 9170 4740 9230 4760
rect 9170 4700 9180 4740
rect 9220 4700 9230 4740
rect 9170 4680 9230 4700
rect 9280 4750 9360 4760
rect 9280 4690 9290 4750
rect 9350 4690 9360 4750
rect 9280 4680 9360 4690
rect 9410 4740 9470 4760
rect 9410 4700 9420 4740
rect 9460 4700 9470 4740
rect 9410 4680 9470 4700
rect 9650 4740 9710 4760
rect 9650 4700 9660 4740
rect 9700 4700 9710 4740
rect 9650 4680 9710 4700
rect 9890 4740 9950 4760
rect 9890 4700 9900 4740
rect 9940 4700 9950 4740
rect 9890 4680 9950 4700
rect 10000 4750 10080 4760
rect 10000 4690 10010 4750
rect 10070 4690 10080 4750
rect 10000 4680 10080 4690
rect 10130 4740 10190 4760
rect 10130 4700 10140 4740
rect 10180 4700 10190 4740
rect 10130 4680 10190 4700
rect 10370 4740 10430 4760
rect 10370 4700 10380 4740
rect 10420 4700 10430 4740
rect 10370 4680 10430 4700
rect 10610 4740 10670 4760
rect 10610 4700 10620 4740
rect 10660 4700 10670 4740
rect 10610 4680 10670 4700
rect 10720 4750 10800 4760
rect 10720 4690 10730 4750
rect 10790 4690 10800 4750
rect 10720 4680 10800 4690
rect 5580 4400 5660 4420
rect 5580 4360 5600 4400
rect 5640 4360 5660 4400
rect 5580 4340 5660 4360
rect 5760 4410 5840 4420
rect 5760 4350 5770 4410
rect 5830 4350 5840 4410
rect 5760 4340 5840 4350
rect 6000 4400 6080 4420
rect 6000 4360 6020 4400
rect 6060 4360 6080 4400
rect 6000 4340 6080 4360
rect 6240 4400 6320 4420
rect 6240 4360 6260 4400
rect 6300 4360 6320 4400
rect 6240 4340 6320 4360
rect 6480 4410 6560 4420
rect 6480 4350 6490 4410
rect 6550 4350 6560 4410
rect 6480 4340 6560 4350
rect 6720 4400 6800 4420
rect 6720 4360 6740 4400
rect 6780 4360 6800 4400
rect 6720 4340 6800 4360
rect 6960 4400 7040 4420
rect 6960 4360 6980 4400
rect 7020 4360 7040 4400
rect 6960 4340 7040 4360
rect 7200 4410 7280 4420
rect 7200 4350 7210 4410
rect 7270 4350 7280 4410
rect 7200 4340 7280 4350
rect 7440 4400 7520 4420
rect 7440 4360 7460 4400
rect 7500 4360 7520 4400
rect 7440 4340 7520 4360
rect 7630 4400 7690 4420
rect 7630 4360 7640 4400
rect 7680 4360 7690 4400
rect 7630 4340 7690 4360
rect 5600 4300 5640 4340
rect 6020 4300 6060 4340
rect 6260 4300 6300 4340
rect 5580 4290 5660 4300
rect 5580 4230 5590 4290
rect 5650 4230 5660 4290
rect 5580 4220 5660 4230
rect 6000 4290 6080 4300
rect 6000 4230 6010 4290
rect 6070 4230 6080 4290
rect 6000 4220 6080 4230
rect 6240 4290 6320 4300
rect 6240 4230 6250 4290
rect 6310 4230 6320 4290
rect 6240 4220 6320 4230
rect 6520 4130 6560 4340
rect 6740 4300 6780 4340
rect 6980 4300 7020 4340
rect 7460 4300 7500 4340
rect 7640 4300 7680 4340
rect 6720 4290 6800 4300
rect 6720 4230 6730 4290
rect 6790 4230 6800 4290
rect 6720 4220 6800 4230
rect 6960 4290 7040 4300
rect 6960 4230 6970 4290
rect 7030 4230 7040 4290
rect 6960 4220 7040 4230
rect 7440 4290 7520 4300
rect 7440 4230 7450 4290
rect 7510 4230 7520 4290
rect 7440 4220 7520 4230
rect 7620 4290 7700 4300
rect 7620 4230 7630 4290
rect 7690 4230 7700 4290
rect 7620 4220 7700 4230
rect 6500 4120 6580 4130
rect 6380 4090 6460 4100
rect 6380 4030 6390 4090
rect 6450 4030 6460 4090
rect 6500 4060 6510 4120
rect 6570 4060 6580 4120
rect 6500 4050 6580 4060
rect 6380 4020 6460 4030
rect 6520 4010 6560 4050
rect 6740 4010 6780 4220
rect 6980 4120 7060 4130
rect 6980 4060 6990 4120
rect 7050 4060 7060 4120
rect 6980 4050 7060 4060
rect 7460 4120 7540 4130
rect 7460 4060 7470 4120
rect 7530 4060 7540 4120
rect 7460 4050 7540 4060
rect 7000 4010 7040 4050
rect 7480 4010 7520 4050
rect 6260 4000 6340 4010
rect 6260 3940 6270 4000
rect 6330 3940 6340 4000
rect 6260 3930 6340 3940
rect 6510 3990 6570 4010
rect 6510 3950 6520 3990
rect 6560 3950 6570 3990
rect 6510 3930 6570 3950
rect 6740 4000 6820 4010
rect 6740 3940 6750 4000
rect 6810 3940 6820 4000
rect 6740 3930 6820 3940
rect 6990 3990 7050 4010
rect 6990 3950 7000 3990
rect 7040 3950 7050 3990
rect 6990 3930 7050 3950
rect 7220 4000 7300 4010
rect 7220 3940 7230 4000
rect 7290 3940 7300 4000
rect 7220 3930 7300 3940
rect 7470 3990 7530 4010
rect 7470 3950 7480 3990
rect 7520 3950 7530 3990
rect 7470 3930 7530 3950
rect 7580 3880 7660 3890
rect 7580 3820 7590 3880
rect 7650 3820 7660 3880
rect 7580 3810 7660 3820
rect 6260 3760 6340 3770
rect 6260 3700 6270 3760
rect 6330 3700 6340 3760
rect 6260 3690 6340 3700
rect 6390 3750 6450 3770
rect 6390 3710 6400 3750
rect 6440 3710 6450 3750
rect 6390 3690 6450 3710
rect 6630 3750 6690 3770
rect 6630 3710 6640 3750
rect 6680 3710 6690 3750
rect 6630 3690 6690 3710
rect 6870 3750 6930 3770
rect 6870 3710 6880 3750
rect 6920 3710 6930 3750
rect 6870 3690 6930 3710
rect 7110 3750 7170 3770
rect 7110 3710 7120 3750
rect 7160 3710 7170 3750
rect 7110 3690 7170 3710
rect 7350 3750 7410 3770
rect 7350 3710 7360 3750
rect 7400 3710 7410 3750
rect 7350 3690 7410 3710
rect 6400 3650 6440 3690
rect 6640 3650 6680 3690
rect 6880 3650 6920 3690
rect 7120 3650 7160 3690
rect 7360 3650 7400 3690
rect 5780 3640 5860 3650
rect 5780 3580 5790 3640
rect 5850 3580 5860 3640
rect 5780 3570 5860 3580
rect 6380 3640 6460 3650
rect 6380 3580 6390 3640
rect 6450 3580 6460 3640
rect 6380 3570 6460 3580
rect 6620 3640 6700 3650
rect 6620 3580 6630 3640
rect 6690 3580 6700 3640
rect 6620 3570 6700 3580
rect 6860 3640 6940 3650
rect 6860 3580 6870 3640
rect 6930 3580 6940 3640
rect 6860 3570 6940 3580
rect 7100 3640 7180 3650
rect 7100 3580 7110 3640
rect 7170 3580 7180 3640
rect 7100 3570 7180 3580
rect 7340 3640 7420 3650
rect 7340 3580 7350 3640
rect 7410 3580 7420 3640
rect 7340 3570 7420 3580
rect 5800 3420 5840 3570
rect 5960 3440 6040 3450
rect 5780 3400 5860 3420
rect 5780 3360 5800 3400
rect 5840 3360 5860 3400
rect 5960 3380 5970 3440
rect 6030 3380 6040 3440
rect 5960 3370 6040 3380
rect 6200 3440 6280 3450
rect 6200 3380 6210 3440
rect 6270 3380 6280 3440
rect 6200 3370 6280 3380
rect 6440 3440 6520 3450
rect 6440 3380 6450 3440
rect 6510 3380 6520 3440
rect 6440 3370 6520 3380
rect 6680 3440 6760 3450
rect 6680 3380 6690 3440
rect 6750 3380 6760 3440
rect 6680 3370 6760 3380
rect 7160 3440 7240 3450
rect 7160 3380 7170 3440
rect 7230 3380 7240 3440
rect 7160 3370 7240 3380
rect 7400 3440 7480 3450
rect 7400 3380 7410 3440
rect 7470 3380 7480 3440
rect 7400 3370 7480 3380
rect 7640 3440 7720 3450
rect 7640 3380 7650 3440
rect 7710 3380 7720 3440
rect 7960 3420 8000 4680
rect 8120 3880 8200 3890
rect 8120 3820 8130 3880
rect 8190 3820 8200 3880
rect 8120 3810 8200 3820
rect 7640 3370 7720 3380
rect 7940 3400 8020 3420
rect 5780 3340 5860 3360
rect 7940 3360 7960 3400
rect 8000 3360 8020 3400
rect 7940 3340 8020 3360
rect 8140 2820 8180 3810
rect 8320 3420 8360 4680
rect 8630 4400 8690 4420
rect 8630 4360 8640 4400
rect 8680 4360 8690 4400
rect 8630 4340 8690 4360
rect 8800 4400 8880 4420
rect 8800 4360 8820 4400
rect 8860 4360 8880 4400
rect 8800 4340 8880 4360
rect 9040 4410 9120 4420
rect 9040 4350 9050 4410
rect 9110 4350 9120 4410
rect 9040 4340 9120 4350
rect 9280 4400 9360 4420
rect 9280 4360 9300 4400
rect 9340 4360 9360 4400
rect 9280 4340 9360 4360
rect 9520 4400 9600 4420
rect 9520 4360 9540 4400
rect 9580 4360 9600 4400
rect 9520 4340 9600 4360
rect 9760 4410 9840 4420
rect 9760 4350 9770 4410
rect 9830 4350 9840 4410
rect 9760 4340 9840 4350
rect 10000 4400 10080 4420
rect 10000 4360 10020 4400
rect 10060 4360 10080 4400
rect 10000 4340 10080 4360
rect 10240 4400 10320 4420
rect 10240 4360 10260 4400
rect 10300 4360 10320 4400
rect 10240 4340 10320 4360
rect 10480 4410 10560 4420
rect 10480 4350 10490 4410
rect 10550 4350 10560 4410
rect 10480 4340 10560 4350
rect 10660 4400 10740 4420
rect 10660 4360 10680 4400
rect 10720 4360 10740 4400
rect 10660 4340 10740 4360
rect 8640 4300 8680 4340
rect 8820 4300 8860 4340
rect 9300 4300 9340 4340
rect 9540 4300 9580 4340
rect 8620 4290 8700 4300
rect 8620 4230 8630 4290
rect 8690 4230 8700 4290
rect 8620 4220 8700 4230
rect 8800 4290 8880 4300
rect 8800 4230 8810 4290
rect 8870 4230 8880 4290
rect 8800 4220 8880 4230
rect 9280 4290 9360 4300
rect 9280 4230 9290 4290
rect 9350 4230 9360 4290
rect 9280 4220 9360 4230
rect 9520 4290 9600 4300
rect 9520 4230 9530 4290
rect 9590 4230 9600 4290
rect 9520 4220 9600 4230
rect 8780 4120 8860 4130
rect 8780 4060 8790 4120
rect 8850 4060 8860 4120
rect 8780 4050 8860 4060
rect 9260 4120 9340 4130
rect 9260 4060 9270 4120
rect 9330 4060 9340 4120
rect 9260 4050 9340 4060
rect 8800 4010 8840 4050
rect 9280 4010 9320 4050
rect 9520 4010 9560 4220
rect 9760 4130 9800 4340
rect 10020 4300 10060 4340
rect 10260 4300 10300 4340
rect 10680 4300 10720 4340
rect 11070 4300 11110 5230
rect 11140 5100 11220 5110
rect 11140 5040 11150 5100
rect 11210 5040 11220 5100
rect 11140 5030 11220 5040
rect 10000 4290 10080 4300
rect 10000 4230 10010 4290
rect 10070 4230 10080 4290
rect 10000 4220 10080 4230
rect 10240 4290 10320 4300
rect 10240 4230 10250 4290
rect 10310 4230 10320 4290
rect 10240 4220 10320 4230
rect 10660 4290 10740 4300
rect 10660 4230 10670 4290
rect 10730 4230 10740 4290
rect 10660 4220 10740 4230
rect 11050 4290 11130 4300
rect 11050 4230 11060 4290
rect 11120 4230 11130 4290
rect 11050 4220 11130 4230
rect 9740 4120 9820 4130
rect 9740 4060 9750 4120
rect 9810 4060 9820 4120
rect 11160 4100 11200 5030
rect 9740 4050 9820 4060
rect 9860 4090 9940 4100
rect 9760 4010 9800 4050
rect 9860 4030 9870 4090
rect 9930 4030 9940 4090
rect 9860 4020 9940 4030
rect 11140 4090 11220 4100
rect 11140 4030 11150 4090
rect 11210 4030 11220 4090
rect 11140 4020 11220 4030
rect 8790 3990 8850 4010
rect 8790 3950 8800 3990
rect 8840 3950 8850 3990
rect 8790 3930 8850 3950
rect 9020 4000 9100 4010
rect 9020 3940 9030 4000
rect 9090 3940 9100 4000
rect 9020 3930 9100 3940
rect 9270 3990 9330 4010
rect 9270 3950 9280 3990
rect 9320 3950 9330 3990
rect 9270 3930 9330 3950
rect 9500 4000 9580 4010
rect 9500 3940 9510 4000
rect 9570 3940 9580 4000
rect 9500 3930 9580 3940
rect 9750 3990 9810 4010
rect 9750 3950 9760 3990
rect 9800 3950 9810 3990
rect 9750 3930 9810 3950
rect 9980 4000 10060 4010
rect 9980 3940 9990 4000
rect 10050 3940 10060 4000
rect 9980 3930 10060 3940
rect 8660 3880 8740 3890
rect 8660 3820 8670 3880
rect 8730 3820 8740 3880
rect 8660 3810 8740 3820
rect 11250 3770 11290 6250
rect 8910 3750 8970 3770
rect 8910 3710 8920 3750
rect 8960 3710 8970 3750
rect 8910 3690 8970 3710
rect 9150 3750 9210 3770
rect 9150 3710 9160 3750
rect 9200 3710 9210 3750
rect 9150 3690 9210 3710
rect 9390 3750 9450 3770
rect 9390 3710 9400 3750
rect 9440 3710 9450 3750
rect 9390 3690 9450 3710
rect 9630 3750 9690 3770
rect 9630 3710 9640 3750
rect 9680 3710 9690 3750
rect 9630 3690 9690 3710
rect 9870 3750 9930 3770
rect 9870 3710 9880 3750
rect 9920 3710 9930 3750
rect 9870 3690 9930 3710
rect 9980 3760 10060 3770
rect 9980 3700 9990 3760
rect 10050 3700 10060 3760
rect 9980 3690 10060 3700
rect 11230 3760 11310 3770
rect 11230 3700 11240 3760
rect 11300 3700 11310 3760
rect 11230 3690 11310 3700
rect 8920 3650 8960 3690
rect 9160 3650 9200 3690
rect 9400 3650 9440 3690
rect 9640 3650 9680 3690
rect 9880 3650 9920 3690
rect 8900 3640 8980 3650
rect 8900 3580 8910 3640
rect 8970 3580 8980 3640
rect 8900 3570 8980 3580
rect 9140 3640 9220 3650
rect 9140 3580 9150 3640
rect 9210 3580 9220 3640
rect 9140 3570 9220 3580
rect 9380 3640 9460 3650
rect 9380 3580 9390 3640
rect 9450 3580 9460 3640
rect 9380 3570 9460 3580
rect 9620 3640 9700 3650
rect 9620 3580 9630 3640
rect 9690 3580 9700 3640
rect 9620 3570 9700 3580
rect 9860 3640 9940 3650
rect 9860 3580 9870 3640
rect 9930 3580 9940 3640
rect 9860 3570 9940 3580
rect 10460 3640 10540 3650
rect 10460 3580 10470 3640
rect 10530 3580 10540 3640
rect 10460 3570 10540 3580
rect 8600 3440 8680 3450
rect 8300 3400 8380 3420
rect 8300 3360 8320 3400
rect 8360 3360 8380 3400
rect 8600 3380 8610 3440
rect 8670 3380 8680 3440
rect 8600 3370 8680 3380
rect 8840 3440 8920 3450
rect 8840 3380 8850 3440
rect 8910 3380 8920 3440
rect 8840 3370 8920 3380
rect 9080 3440 9160 3450
rect 9080 3380 9090 3440
rect 9150 3380 9160 3440
rect 9080 3370 9160 3380
rect 9560 3440 9640 3450
rect 9560 3380 9570 3440
rect 9630 3380 9640 3440
rect 9560 3370 9640 3380
rect 9800 3440 9880 3450
rect 9800 3380 9810 3440
rect 9870 3380 9880 3440
rect 9800 3370 9880 3380
rect 10040 3440 10120 3450
rect 10040 3380 10050 3440
rect 10110 3380 10120 3440
rect 10040 3370 10120 3380
rect 10280 3440 10360 3450
rect 10280 3380 10290 3440
rect 10350 3380 10360 3440
rect 10480 3420 10520 3570
rect 10280 3370 10360 3380
rect 10460 3400 10540 3420
rect 8300 3340 8380 3360
rect 10460 3360 10480 3400
rect 10520 3360 10540 3400
rect 10460 3340 10540 3360
rect 6860 2810 6940 2820
rect 6860 2750 6870 2810
rect 6930 2750 6940 2810
rect 6860 2740 6940 2750
rect 8120 2810 8200 2820
rect 8120 2750 8130 2810
rect 8190 2750 8200 2810
rect 8120 2740 8200 2750
rect 9380 2810 9460 2820
rect 9380 2750 9390 2810
rect 9450 2750 9460 2810
rect 9380 2740 9460 2750
rect 8140 2630 8180 2740
rect 8120 2620 8200 2630
rect 8120 2560 8130 2620
rect 8190 2560 8200 2620
rect 8120 2550 8200 2560
rect 6040 2510 6120 2520
rect 6040 2450 6050 2510
rect 6110 2450 6120 2510
rect 6040 2440 6120 2450
rect 6200 2510 6280 2520
rect 6200 2450 6210 2510
rect 6270 2450 6280 2510
rect 6200 2440 6280 2450
rect 6360 2510 6440 2520
rect 6360 2450 6370 2510
rect 6430 2450 6440 2510
rect 6360 2440 6440 2450
rect 6520 2510 6600 2520
rect 6520 2450 6530 2510
rect 6590 2450 6600 2510
rect 6520 2440 6600 2450
rect 6680 2510 6760 2520
rect 6680 2450 6690 2510
rect 6750 2450 6760 2510
rect 6680 2440 6760 2450
rect 6840 2510 6920 2520
rect 6840 2450 6850 2510
rect 6910 2450 6920 2510
rect 6840 2440 6920 2450
rect 7000 2510 7080 2520
rect 7000 2450 7010 2510
rect 7070 2450 7080 2510
rect 7000 2440 7080 2450
rect 7160 2510 7240 2520
rect 7160 2450 7170 2510
rect 7230 2450 7240 2510
rect 7160 2440 7240 2450
rect 7320 2510 7400 2520
rect 7320 2450 7330 2510
rect 7390 2450 7400 2510
rect 7320 2440 7400 2450
rect 7480 2510 7560 2520
rect 7480 2450 7490 2510
rect 7550 2450 7560 2510
rect 7480 2440 7560 2450
rect 7640 2510 7720 2520
rect 7640 2450 7650 2510
rect 7710 2450 7720 2510
rect 7640 2440 7720 2450
rect 7800 2510 7880 2520
rect 7800 2450 7810 2510
rect 7870 2450 7880 2510
rect 7800 2440 7880 2450
rect 7960 2510 8040 2520
rect 7960 2450 7970 2510
rect 8030 2450 8040 2510
rect 7960 2440 8040 2450
rect 8120 2510 8200 2520
rect 8120 2450 8130 2510
rect 8190 2450 8200 2510
rect 8120 2440 8200 2450
rect 8280 2510 8360 2520
rect 8280 2450 8290 2510
rect 8350 2450 8360 2510
rect 8280 2440 8360 2450
rect 8440 2510 8520 2520
rect 8440 2450 8450 2510
rect 8510 2450 8520 2510
rect 8440 2440 8520 2450
rect 8600 2510 8680 2520
rect 8600 2450 8610 2510
rect 8670 2450 8680 2510
rect 8600 2440 8680 2450
rect 8760 2510 8840 2520
rect 8760 2450 8770 2510
rect 8830 2450 8840 2510
rect 8760 2440 8840 2450
rect 8920 2510 9000 2520
rect 8920 2450 8930 2510
rect 8990 2450 9000 2510
rect 8920 2440 9000 2450
rect 9080 2510 9160 2520
rect 9080 2450 9090 2510
rect 9150 2450 9160 2510
rect 9080 2440 9160 2450
rect 9240 2510 9320 2520
rect 9240 2450 9250 2510
rect 9310 2450 9320 2510
rect 9240 2440 9320 2450
rect 9400 2510 9480 2520
rect 9400 2450 9410 2510
rect 9470 2450 9480 2510
rect 9400 2440 9480 2450
rect 9560 2510 9640 2520
rect 9560 2450 9570 2510
rect 9630 2450 9640 2510
rect 9560 2440 9640 2450
rect 9720 2510 9800 2520
rect 9720 2450 9730 2510
rect 9790 2450 9800 2510
rect 9720 2440 9800 2450
rect 9880 2510 9960 2520
rect 9880 2450 9890 2510
rect 9950 2450 9960 2510
rect 9880 2440 9960 2450
rect 10040 2510 10120 2520
rect 10040 2450 10050 2510
rect 10110 2450 10120 2510
rect 10040 2440 10120 2450
rect 5960 2340 6040 2350
rect 5960 2280 5970 2340
rect 6030 2280 6040 2340
rect 5960 2270 6040 2280
rect 10270 2340 10350 2350
rect 10270 2280 10280 2340
rect 10340 2280 10350 2340
rect 10270 2270 10350 2280
rect 6330 2100 6410 2110
rect 6330 2040 6340 2100
rect 6400 2040 6410 2100
rect 6330 2030 6410 2040
rect 8120 2100 8200 2110
rect 8120 2040 8130 2100
rect 8190 2040 8200 2100
rect 8120 2030 8200 2040
rect 9910 2100 9990 2110
rect 9910 2040 9920 2100
rect 9980 2040 9990 2100
rect 9910 2030 9990 2040
rect 6350 1970 6390 2030
rect 8140 1970 8180 2030
rect 9930 1970 9970 2030
rect 5790 1960 5870 1970
rect 5790 1900 5800 1960
rect 5860 1900 5870 1960
rect 5790 1890 5870 1900
rect 6150 1960 6230 1970
rect 6150 1900 6160 1960
rect 6220 1900 6230 1960
rect 6150 1890 6230 1900
rect 6330 1950 6410 1970
rect 6330 1910 6350 1950
rect 6390 1910 6410 1950
rect 6330 1890 6410 1910
rect 6510 1960 6590 1970
rect 6510 1900 6520 1960
rect 6580 1900 6590 1960
rect 6510 1890 6590 1900
rect 7580 1960 7660 1970
rect 7580 1900 7590 1960
rect 7650 1900 7660 1960
rect 7580 1890 7660 1900
rect 7940 1960 8020 1970
rect 7940 1900 7950 1960
rect 8010 1900 8020 1960
rect 7940 1890 8020 1900
rect 8120 1950 8200 1970
rect 8120 1910 8140 1950
rect 8180 1910 8200 1950
rect 8120 1890 8200 1910
rect 8300 1960 8380 1970
rect 8300 1900 8310 1960
rect 8370 1900 8380 1960
rect 8300 1890 8380 1900
rect 8660 1960 8740 1970
rect 8660 1900 8670 1960
rect 8730 1900 8740 1960
rect 8660 1890 8740 1900
rect 9730 1960 9810 1970
rect 9730 1900 9740 1960
rect 9800 1900 9810 1960
rect 9730 1890 9810 1900
rect 9910 1950 9990 1970
rect 9910 1910 9930 1950
rect 9970 1910 9990 1950
rect 9910 1890 9990 1910
rect 10090 1960 10170 1970
rect 10090 1900 10100 1960
rect 10160 1900 10170 1960
rect 10090 1890 10170 1900
rect 10450 1960 10530 1970
rect 10450 1900 10460 1960
rect 10520 1900 10530 1960
rect 10450 1890 10530 1900
rect 6990 1790 7070 1800
rect 6990 1730 7000 1790
rect 7060 1730 7070 1790
rect 6990 1720 7070 1730
rect 7100 1790 7180 1800
rect 7100 1730 7110 1790
rect 7170 1730 7180 1790
rect 7100 1720 7180 1730
rect 9140 1790 9220 1800
rect 9140 1730 9150 1790
rect 9210 1730 9220 1790
rect 9140 1720 9220 1730
rect 9250 1790 9330 1800
rect 9250 1730 9260 1790
rect 9320 1730 9330 1790
rect 9250 1720 9330 1730
rect 10930 1790 11010 1800
rect 10930 1730 10940 1790
rect 11000 1730 11010 1790
rect 10930 1720 11010 1730
rect 5610 1620 5690 1630
rect 5610 1560 5620 1620
rect 5680 1560 5690 1620
rect 5610 1550 5690 1560
rect 5970 1610 6050 1630
rect 5970 1570 5990 1610
rect 6030 1570 6050 1610
rect 5970 1550 6050 1570
rect 6330 1620 6410 1630
rect 6330 1560 6340 1620
rect 6400 1560 6410 1620
rect 6330 1550 6410 1560
rect 6690 1610 6770 1630
rect 6690 1570 6710 1610
rect 6750 1570 6770 1610
rect 6690 1550 6770 1570
rect 7490 1610 7570 1630
rect 7490 1570 7510 1610
rect 7550 1570 7570 1610
rect 7490 1550 7570 1570
rect 7760 1610 7840 1630
rect 7760 1570 7780 1610
rect 7820 1570 7840 1610
rect 7760 1550 7840 1570
rect 8120 1620 8200 1630
rect 8120 1560 8130 1620
rect 8190 1560 8200 1620
rect 8120 1550 8200 1560
rect 8480 1620 8560 1630
rect 8480 1560 8490 1620
rect 8550 1560 8560 1620
rect 8480 1550 8560 1560
rect 8840 1620 8920 1630
rect 8840 1560 8850 1620
rect 8910 1560 8920 1620
rect 8840 1550 8920 1560
rect 9550 1610 9630 1630
rect 9550 1570 9570 1610
rect 9610 1570 9630 1610
rect 9550 1550 9630 1570
rect 9910 1620 9990 1630
rect 9910 1560 9920 1620
rect 9980 1560 9990 1620
rect 9910 1550 9990 1560
rect 10270 1610 10350 1630
rect 10270 1570 10290 1610
rect 10330 1570 10350 1610
rect 10270 1550 10350 1570
rect 10630 1620 10710 1630
rect 10630 1560 10640 1620
rect 10700 1560 10710 1620
rect 10630 1550 10710 1560
rect 5110 1420 5190 1430
rect 5110 1360 5120 1420
rect 5180 1360 5190 1420
rect 5110 1350 5190 1360
rect 5630 1140 5670 1550
rect 5990 1520 6030 1550
rect 6710 1520 6750 1550
rect 5970 1510 6050 1520
rect 5970 1450 5980 1510
rect 6040 1450 6050 1510
rect 5970 1440 6050 1450
rect 6690 1510 6770 1520
rect 6690 1450 6700 1510
rect 6760 1450 6770 1510
rect 6690 1440 6770 1450
rect 7510 1430 7550 1550
rect 7490 1420 7570 1430
rect 7490 1360 7500 1420
rect 7560 1360 7570 1420
rect 7490 1350 7570 1360
rect 7780 1140 7820 1550
rect 8120 1510 8200 1520
rect 8120 1450 8130 1510
rect 8190 1450 8200 1510
rect 8120 1440 8200 1450
rect 8140 1140 8180 1440
rect 8500 1140 8540 1550
rect 9570 1520 9610 1550
rect 10290 1520 10330 1550
rect 9550 1510 9630 1520
rect 9550 1450 9560 1510
rect 9620 1450 9630 1510
rect 9550 1440 9630 1450
rect 10270 1510 10350 1520
rect 10270 1450 10280 1510
rect 10340 1450 10350 1510
rect 10270 1440 10350 1450
rect 10650 1140 10690 1550
<< via1 >>
rect 2710 7690 2770 7750
rect -20 7530 40 7590
rect 1890 7530 1950 7590
rect -110 7420 -50 7480
rect -110 6050 -50 6110
rect 2520 7320 2580 7380
rect 150 7220 210 7280
rect 142 7170 212 7180
rect 142 7120 152 7170
rect 152 7120 202 7170
rect 202 7120 212 7170
rect 142 7110 212 7120
rect 142 7050 212 7060
rect 142 7000 152 7050
rect 152 7000 202 7050
rect 202 7000 212 7050
rect 142 6990 212 7000
rect 8890 7630 8950 7690
rect 3290 7530 3350 7590
rect 5030 7540 5090 7600
rect 9610 7530 9670 7590
rect 2712 6900 2782 6910
rect 2712 6850 2722 6900
rect 2722 6850 2772 6900
rect 2772 6850 2782 6900
rect 2712 6840 2782 6850
rect 150 6690 210 6750
rect 2520 6690 2580 6750
rect 2712 6780 2782 6790
rect 2712 6730 2722 6780
rect 2722 6730 2772 6780
rect 2772 6730 2782 6780
rect 2712 6720 2782 6730
rect 142 6640 212 6650
rect 142 6590 152 6640
rect 152 6590 202 6640
rect 202 6590 212 6640
rect 142 6580 212 6590
rect 142 6520 212 6530
rect 142 6470 152 6520
rect 152 6470 202 6520
rect 202 6470 212 6520
rect 142 6460 212 6470
rect 2380 6570 2440 6580
rect 2380 6530 2390 6570
rect 2390 6530 2430 6570
rect 2430 6530 2440 6570
rect 2380 6520 2440 6530
rect 2590 6570 2650 6580
rect 2590 6530 2600 6570
rect 2600 6530 2640 6570
rect 2640 6530 2650 6570
rect 2590 6520 2650 6530
rect 1200 6380 1260 6390
rect 1200 6340 1210 6380
rect 1210 6340 1250 6380
rect 1250 6340 1260 6380
rect 1200 6330 1260 6340
rect 4850 6420 4920 6430
rect 4850 6370 4860 6420
rect 4860 6370 4910 6420
rect 4910 6370 4920 6420
rect 4850 6360 4920 6370
rect 4850 6300 4920 6310
rect 4850 6250 4860 6300
rect 4860 6250 4910 6300
rect 4910 6250 4920 6300
rect 4850 6240 4920 6250
rect 532 6110 602 6120
rect 532 6060 542 6110
rect 542 6060 592 6110
rect 592 6060 602 6110
rect 532 6050 602 6060
rect 1878 6110 1948 6120
rect 1878 6060 1888 6110
rect 1888 6060 1938 6110
rect 1938 6060 1948 6110
rect 1878 6050 1948 6060
rect 2430 6050 2490 6110
rect 2220 5840 2280 5900
rect -20 5640 40 5700
rect 532 5690 602 5700
rect 532 5640 542 5690
rect 542 5640 592 5690
rect 592 5640 602 5690
rect 532 5630 602 5640
rect 1878 5690 1948 5700
rect 1878 5640 1888 5690
rect 1888 5640 1938 5690
rect 1938 5640 1948 5690
rect 1878 5630 1948 5640
rect 3042 5890 3112 5900
rect 3042 5840 3052 5890
rect 3052 5840 3102 5890
rect 3102 5840 3112 5890
rect 3042 5830 3112 5840
rect 4440 5890 4510 5900
rect 4440 5840 4450 5890
rect 4450 5840 4500 5890
rect 4500 5840 4510 5890
rect 4440 5830 4510 5840
rect 4850 5830 4910 5890
rect 2430 5540 2490 5600
rect 4760 5540 4820 5600
rect 4670 5220 4730 5280
rect 4560 5130 4620 5190
rect -210 3380 -150 3440
rect -80 3430 -20 3440
rect -80 3390 -70 3430
rect -70 3390 -30 3430
rect -30 3390 -20 3430
rect -80 3380 -20 3390
rect 2540 3360 2594 3420
rect 4940 5630 5000 5690
rect 4850 5330 4910 5390
rect 4760 4940 4820 5000
rect 4670 4030 4730 4090
rect 4940 4690 5000 4750
rect 10290 7530 10350 7590
rect 5390 7420 5450 7480
rect 6790 7420 6850 7480
rect 9520 7420 9580 7480
rect 9030 7320 9090 7380
rect 5120 7220 5180 7280
rect 6250 7210 6310 7270
rect 5890 7120 5950 7180
rect 7950 7120 8010 7180
rect 8310 7120 8370 7180
rect 9430 7120 9490 7180
rect 5350 7050 5410 7060
rect 5350 7010 5360 7050
rect 5360 7010 5400 7050
rect 5400 7010 5410 7050
rect 5350 7000 5410 7010
rect 5710 7050 5770 7060
rect 5710 7010 5720 7050
rect 5720 7010 5760 7050
rect 5760 7010 5770 7050
rect 5710 7000 5770 7010
rect 6070 7050 6130 7060
rect 6070 7010 6080 7050
rect 6080 7010 6120 7050
rect 6120 7010 6130 7050
rect 6070 7000 6130 7010
rect 6430 7050 6490 7060
rect 6430 7010 6440 7050
rect 6440 7010 6480 7050
rect 6480 7010 6490 7050
rect 6430 7000 6490 7010
rect 7050 7050 7110 7060
rect 7050 7010 7060 7050
rect 7060 7010 7100 7050
rect 7100 7010 7110 7050
rect 7050 7000 7110 7010
rect 7410 7050 7470 7060
rect 7410 7010 7420 7050
rect 7420 7010 7460 7050
rect 7460 7010 7470 7050
rect 7410 7000 7470 7010
rect 7770 7050 7830 7060
rect 7770 7010 7780 7050
rect 7780 7010 7820 7050
rect 7820 7010 7830 7050
rect 7770 7000 7830 7010
rect 8130 7050 8190 7060
rect 8130 7010 8140 7050
rect 8140 7010 8180 7050
rect 8180 7010 8190 7050
rect 8130 7000 8190 7010
rect 8490 7050 8550 7060
rect 8490 7010 8500 7050
rect 8500 7010 8540 7050
rect 8540 7010 8550 7050
rect 8490 7000 8550 7010
rect 8850 7050 8910 7060
rect 8850 7010 8860 7050
rect 8860 7010 8900 7050
rect 8900 7010 8910 7050
rect 8850 7000 8910 7010
rect 9210 7050 9270 7060
rect 9210 7010 9220 7050
rect 9220 7010 9260 7050
rect 9260 7010 9270 7050
rect 9210 7000 9270 7010
rect 5530 6710 5590 6720
rect 5530 6670 5540 6710
rect 5540 6670 5580 6710
rect 5580 6670 5590 6710
rect 5530 6660 5590 6670
rect 5890 6710 5950 6720
rect 5890 6670 5900 6710
rect 5900 6670 5940 6710
rect 5940 6670 5950 6710
rect 5890 6660 5950 6670
rect 6250 6710 6310 6720
rect 6250 6670 6260 6710
rect 6260 6670 6300 6710
rect 6300 6670 6310 6710
rect 6250 6660 6310 6670
rect 7590 6710 7650 6720
rect 7590 6670 7600 6710
rect 7600 6670 7640 6710
rect 7640 6670 7650 6710
rect 7590 6660 7650 6670
rect 7950 6710 8010 6720
rect 7950 6670 7960 6710
rect 7960 6670 8000 6710
rect 8000 6670 8010 6710
rect 7950 6660 8010 6670
rect 8310 6710 8370 6720
rect 8310 6670 8320 6710
rect 8320 6670 8360 6710
rect 8360 6670 8370 6710
rect 8310 6660 8370 6670
rect 8670 6710 8730 6720
rect 8670 6670 8680 6710
rect 8680 6670 8720 6710
rect 8720 6670 8730 6710
rect 8670 6660 8730 6670
rect 5120 6450 5180 6510
rect 5230 6450 5290 6510
rect 5120 6270 5180 6330
rect 5030 4230 5090 4290
rect 4850 3700 4910 3760
rect 4670 3360 4730 3420
rect 4560 2280 4620 2340
rect 6130 6360 6190 6420
rect 5660 6040 5720 6050
rect 5660 6000 5670 6040
rect 5670 6000 5710 6040
rect 5710 6000 5720 6040
rect 5660 5990 5720 6000
rect 7230 6270 7290 6330
rect 9430 6570 9490 6630
rect 9520 6460 9580 6520
rect 10370 7120 10430 7180
rect 9830 7050 9890 7060
rect 9830 7010 9840 7050
rect 9840 7010 9880 7050
rect 9880 7010 9890 7050
rect 9830 7000 9890 7010
rect 10190 7050 10250 7060
rect 10190 7010 10200 7050
rect 10200 7010 10240 7050
rect 10240 7010 10250 7050
rect 10190 7000 10250 7010
rect 10550 7050 10610 7060
rect 10550 7010 10560 7050
rect 10560 7010 10600 7050
rect 10600 7010 10610 7050
rect 10550 7000 10610 7010
rect 10910 7050 10970 7060
rect 10910 7010 10920 7050
rect 10920 7010 10960 7050
rect 10960 7010 10970 7050
rect 10910 7000 10970 7010
rect 10010 6710 10070 6720
rect 10010 6670 10020 6710
rect 10020 6670 10060 6710
rect 10060 6670 10070 6710
rect 10010 6660 10070 6670
rect 10370 6710 10430 6720
rect 10370 6670 10380 6710
rect 10380 6670 10420 6710
rect 10420 6670 10430 6710
rect 10370 6660 10430 6670
rect 10730 6710 10790 6720
rect 10730 6670 10740 6710
rect 10740 6670 10780 6710
rect 10780 6670 10790 6710
rect 10730 6660 10790 6670
rect 9950 6550 10010 6610
rect 9610 6350 9670 6410
rect 9030 6260 9090 6320
rect 8670 6190 8730 6250
rect 6510 6120 6570 6130
rect 6510 6080 6520 6120
rect 6520 6080 6560 6120
rect 6560 6080 6570 6120
rect 6510 6070 6570 6080
rect 6870 6120 6930 6130
rect 6870 6080 6880 6120
rect 6880 6080 6920 6120
rect 6920 6080 6930 6120
rect 6870 6070 6930 6080
rect 7230 6120 7290 6130
rect 7230 6080 7240 6120
rect 7240 6080 7280 6120
rect 7280 6080 7290 6120
rect 7230 6070 7290 6080
rect 7590 6120 7650 6130
rect 7590 6080 7600 6120
rect 7600 6080 7640 6120
rect 7640 6080 7650 6120
rect 7590 6070 7650 6080
rect 7950 6120 8010 6130
rect 7950 6080 7960 6120
rect 7960 6080 8000 6120
rect 8000 6080 8010 6120
rect 7950 6070 8010 6080
rect 8310 6120 8370 6130
rect 8310 6080 8320 6120
rect 8320 6080 8360 6120
rect 8360 6080 8370 6120
rect 8310 6070 8370 6080
rect 8670 6120 8730 6130
rect 8670 6080 8680 6120
rect 8680 6080 8720 6120
rect 8720 6080 8730 6120
rect 8670 6070 8730 6080
rect 9030 6120 9090 6130
rect 9030 6080 9040 6120
rect 9040 6080 9080 6120
rect 9080 6080 9090 6120
rect 9030 6070 9090 6080
rect 9390 6120 9450 6130
rect 9390 6080 9400 6120
rect 9400 6080 9440 6120
rect 9440 6080 9450 6120
rect 9390 6070 9450 6080
rect 9750 6120 9810 6130
rect 9750 6080 9760 6120
rect 9760 6080 9800 6120
rect 9800 6080 9810 6120
rect 9750 6070 9810 6080
rect 5660 5920 5720 5930
rect 5660 5880 5670 5920
rect 5670 5880 5710 5920
rect 5710 5880 5720 5920
rect 5660 5870 5720 5880
rect 6130 5870 6190 5930
rect 5530 5580 5590 5590
rect 5530 5540 5540 5580
rect 5540 5540 5580 5580
rect 5580 5540 5590 5580
rect 5530 5530 5590 5540
rect 5790 5580 5850 5590
rect 5790 5540 5800 5580
rect 5800 5540 5840 5580
rect 5840 5540 5850 5580
rect 5790 5530 5850 5540
rect 6250 5530 6310 5590
rect 6130 5220 6190 5280
rect 5660 5130 5720 5190
rect 5230 5040 5290 5100
rect 5650 4810 5710 4870
rect 5890 4810 5950 4870
rect 6130 4810 6190 4870
rect 7770 5380 7830 5390
rect 7770 5340 7780 5380
rect 7780 5340 7820 5380
rect 7820 5340 7830 5380
rect 7770 5330 7830 5340
rect 8490 5380 8550 5390
rect 8490 5340 8500 5380
rect 8500 5340 8540 5380
rect 8540 5340 8550 5380
rect 8490 5330 8550 5340
rect 7410 5220 7470 5280
rect 7050 5130 7110 5190
rect 6690 5040 6750 5100
rect 6370 4810 6430 4870
rect 6610 4860 6670 4870
rect 6610 4820 6620 4860
rect 6620 4820 6660 4860
rect 6660 4820 6670 4860
rect 6610 4810 6670 4820
rect 6850 4810 6910 4870
rect 7090 4810 7150 4870
rect 7330 4810 7390 4870
rect 7570 4810 7630 4870
rect 8850 5220 8910 5280
rect 9210 5130 9270 5190
rect 9390 5130 9450 5190
rect 8130 5040 8190 5100
rect 9570 5040 9630 5100
rect 10130 6460 10190 6520
rect 10040 6350 10100 6410
rect 11240 6260 11300 6320
rect 10730 6040 10790 6060
rect 10730 6000 10740 6040
rect 10740 6000 10780 6040
rect 10780 6000 10790 6040
rect 10730 5990 10790 6000
rect 10730 5920 10790 5930
rect 10730 5880 10740 5920
rect 10740 5880 10780 5920
rect 10780 5880 10790 5920
rect 10730 5870 10790 5880
rect 10530 5580 10590 5590
rect 10530 5540 10540 5580
rect 10540 5540 10580 5580
rect 10580 5540 10590 5580
rect 10530 5530 10590 5540
rect 10930 5580 10990 5590
rect 10930 5540 10940 5580
rect 10940 5540 10980 5580
rect 10980 5540 10990 5580
rect 10930 5530 10990 5540
rect 10130 5240 10190 5300
rect 10040 5130 10100 5190
rect 11060 5240 11120 5300
rect 8570 4940 8630 5000
rect 9950 4940 10010 5000
rect 10730 4940 10790 5000
rect 8690 4860 8750 4870
rect 8690 4820 8700 4860
rect 8700 4820 8740 4860
rect 8740 4820 8750 4860
rect 8690 4810 8750 4820
rect 8930 4860 8990 4870
rect 8930 4820 8940 4860
rect 8940 4820 8980 4860
rect 8980 4820 8990 4860
rect 8930 4810 8990 4820
rect 9170 4860 9230 4870
rect 9170 4820 9180 4860
rect 9180 4820 9220 4860
rect 9220 4820 9230 4860
rect 9170 4810 9230 4820
rect 9410 4860 9470 4870
rect 9410 4820 9420 4860
rect 9420 4820 9460 4860
rect 9460 4820 9470 4860
rect 9410 4810 9470 4820
rect 9650 4860 9710 4870
rect 9650 4820 9660 4860
rect 9660 4820 9700 4860
rect 9700 4820 9710 4860
rect 9650 4810 9710 4820
rect 9890 4860 9950 4870
rect 9890 4820 9900 4860
rect 9900 4820 9940 4860
rect 9940 4820 9950 4860
rect 9890 4810 9950 4820
rect 10130 4860 10190 4870
rect 10130 4820 10140 4860
rect 10140 4820 10180 4860
rect 10180 4820 10190 4860
rect 10130 4810 10190 4820
rect 10370 4860 10430 4870
rect 10370 4820 10380 4860
rect 10380 4820 10420 4860
rect 10420 4820 10430 4860
rect 10370 4810 10430 4820
rect 10610 4860 10670 4870
rect 10610 4820 10620 4860
rect 10620 4820 10660 4860
rect 10660 4820 10670 4860
rect 10610 4810 10670 4820
rect 5530 4740 5590 4750
rect 5530 4700 5540 4740
rect 5540 4700 5580 4740
rect 5580 4700 5590 4740
rect 5530 4690 5590 4700
rect 6250 4740 6310 4750
rect 6250 4700 6260 4740
rect 6260 4700 6300 4740
rect 6300 4700 6310 4740
rect 6250 4690 6310 4700
rect 6970 4740 7030 4750
rect 6970 4700 6980 4740
rect 6980 4700 7020 4740
rect 7020 4700 7030 4740
rect 6970 4690 7030 4700
rect 7690 4740 7750 4750
rect 7690 4700 7700 4740
rect 7700 4700 7740 4740
rect 7740 4700 7750 4740
rect 7690 4690 7750 4700
rect 7950 4690 8010 4750
rect 8310 4690 8370 4750
rect 8570 4740 8630 4750
rect 8570 4700 8580 4740
rect 8580 4700 8620 4740
rect 8620 4700 8630 4740
rect 8570 4690 8630 4700
rect 9290 4740 9350 4750
rect 9290 4700 9300 4740
rect 9300 4700 9340 4740
rect 9340 4700 9350 4740
rect 9290 4690 9350 4700
rect 10010 4740 10070 4750
rect 10010 4700 10020 4740
rect 10020 4700 10060 4740
rect 10060 4700 10070 4740
rect 10010 4690 10070 4700
rect 10730 4740 10790 4750
rect 10730 4700 10740 4740
rect 10740 4700 10780 4740
rect 10780 4700 10790 4740
rect 10730 4690 10790 4700
rect 5770 4400 5830 4410
rect 5770 4360 5780 4400
rect 5780 4360 5820 4400
rect 5820 4360 5830 4400
rect 5770 4350 5830 4360
rect 6490 4400 6550 4410
rect 6490 4360 6500 4400
rect 6500 4360 6540 4400
rect 6540 4360 6550 4400
rect 6490 4350 6550 4360
rect 7210 4400 7270 4410
rect 7210 4360 7220 4400
rect 7220 4360 7260 4400
rect 7260 4360 7270 4400
rect 7210 4350 7270 4360
rect 5590 4230 5650 4290
rect 6010 4230 6070 4290
rect 6250 4230 6310 4290
rect 6730 4230 6790 4290
rect 6970 4230 7030 4290
rect 7450 4230 7510 4290
rect 7630 4230 7690 4290
rect 6390 4080 6450 4090
rect 6390 4040 6400 4080
rect 6400 4040 6440 4080
rect 6440 4040 6450 4080
rect 6390 4030 6450 4040
rect 6510 4060 6570 4120
rect 6990 4060 7050 4120
rect 7470 4060 7530 4120
rect 6270 3990 6330 4000
rect 6270 3950 6280 3990
rect 6280 3950 6320 3990
rect 6320 3950 6330 3990
rect 6270 3940 6330 3950
rect 6750 3990 6810 4000
rect 6750 3950 6760 3990
rect 6760 3950 6800 3990
rect 6800 3950 6810 3990
rect 6750 3940 6810 3950
rect 7230 3990 7290 4000
rect 7230 3950 7240 3990
rect 7240 3950 7280 3990
rect 7280 3950 7290 3990
rect 7230 3940 7290 3950
rect 7590 3870 7650 3880
rect 7590 3830 7600 3870
rect 7600 3830 7640 3870
rect 7640 3830 7650 3870
rect 7590 3820 7650 3830
rect 6270 3750 6330 3760
rect 6270 3710 6280 3750
rect 6280 3710 6320 3750
rect 6320 3710 6330 3750
rect 6270 3700 6330 3710
rect 5790 3580 5850 3640
rect 6390 3580 6450 3640
rect 6630 3580 6690 3640
rect 6870 3580 6930 3640
rect 7110 3580 7170 3640
rect 7350 3580 7410 3640
rect 5970 3430 6030 3440
rect 5970 3390 5980 3430
rect 5980 3390 6020 3430
rect 6020 3390 6030 3430
rect 5970 3380 6030 3390
rect 6210 3430 6270 3440
rect 6210 3390 6220 3430
rect 6220 3390 6260 3430
rect 6260 3390 6270 3430
rect 6210 3380 6270 3390
rect 6450 3430 6510 3440
rect 6450 3390 6460 3430
rect 6460 3390 6500 3430
rect 6500 3390 6510 3430
rect 6450 3380 6510 3390
rect 6690 3430 6750 3440
rect 6690 3390 6700 3430
rect 6700 3390 6740 3430
rect 6740 3390 6750 3430
rect 6690 3380 6750 3390
rect 7170 3430 7230 3440
rect 7170 3390 7180 3430
rect 7180 3390 7220 3430
rect 7220 3390 7230 3430
rect 7170 3380 7230 3390
rect 7410 3430 7470 3440
rect 7410 3390 7420 3430
rect 7420 3390 7460 3430
rect 7460 3390 7470 3430
rect 7410 3380 7470 3390
rect 7650 3430 7710 3440
rect 7650 3390 7660 3430
rect 7660 3390 7700 3430
rect 7700 3390 7710 3430
rect 7650 3380 7710 3390
rect 8130 3820 8190 3880
rect 9050 4400 9110 4410
rect 9050 4360 9060 4400
rect 9060 4360 9100 4400
rect 9100 4360 9110 4400
rect 9050 4350 9110 4360
rect 9770 4400 9830 4410
rect 9770 4360 9780 4400
rect 9780 4360 9820 4400
rect 9820 4360 9830 4400
rect 9770 4350 9830 4360
rect 10490 4400 10550 4410
rect 10490 4360 10500 4400
rect 10500 4360 10540 4400
rect 10540 4360 10550 4400
rect 10490 4350 10550 4360
rect 8630 4230 8690 4290
rect 8810 4230 8870 4290
rect 9290 4230 9350 4290
rect 9530 4230 9590 4290
rect 8790 4060 8850 4120
rect 9270 4060 9330 4120
rect 11150 5040 11210 5100
rect 10010 4230 10070 4290
rect 10250 4230 10310 4290
rect 10670 4230 10730 4290
rect 11060 4230 11120 4290
rect 9750 4060 9810 4120
rect 9870 4080 9930 4090
rect 9870 4040 9880 4080
rect 9880 4040 9920 4080
rect 9920 4040 9930 4080
rect 9870 4030 9930 4040
rect 11150 4030 11210 4090
rect 9030 3990 9090 4000
rect 9030 3950 9040 3990
rect 9040 3950 9080 3990
rect 9080 3950 9090 3990
rect 9030 3940 9090 3950
rect 9510 3990 9570 4000
rect 9510 3950 9520 3990
rect 9520 3950 9560 3990
rect 9560 3950 9570 3990
rect 9510 3940 9570 3950
rect 9990 3990 10050 4000
rect 9990 3950 10000 3990
rect 10000 3950 10040 3990
rect 10040 3950 10050 3990
rect 9990 3940 10050 3950
rect 8670 3870 8730 3880
rect 8670 3830 8680 3870
rect 8680 3830 8720 3870
rect 8720 3830 8730 3870
rect 8670 3820 8730 3830
rect 9990 3750 10050 3760
rect 9990 3710 10000 3750
rect 10000 3710 10040 3750
rect 10040 3710 10050 3750
rect 9990 3700 10050 3710
rect 11240 3700 11300 3760
rect 8910 3580 8970 3640
rect 9150 3580 9210 3640
rect 9390 3580 9450 3640
rect 9630 3580 9690 3640
rect 9870 3580 9930 3640
rect 10470 3580 10530 3640
rect 8610 3430 8670 3440
rect 8610 3390 8620 3430
rect 8620 3390 8660 3430
rect 8660 3390 8670 3430
rect 8610 3380 8670 3390
rect 8850 3430 8910 3440
rect 8850 3390 8860 3430
rect 8860 3390 8900 3430
rect 8900 3390 8910 3430
rect 8850 3380 8910 3390
rect 9090 3430 9150 3440
rect 9090 3390 9100 3430
rect 9100 3390 9140 3430
rect 9140 3390 9150 3430
rect 9090 3380 9150 3390
rect 9570 3430 9630 3440
rect 9570 3390 9580 3430
rect 9580 3390 9620 3430
rect 9620 3390 9630 3430
rect 9570 3380 9630 3390
rect 9810 3430 9870 3440
rect 9810 3390 9820 3430
rect 9820 3390 9860 3430
rect 9860 3390 9870 3430
rect 9810 3380 9870 3390
rect 10050 3430 10110 3440
rect 10050 3390 10060 3430
rect 10060 3390 10100 3430
rect 10100 3390 10110 3430
rect 10050 3380 10110 3390
rect 10290 3430 10350 3440
rect 10290 3390 10300 3430
rect 10300 3390 10340 3430
rect 10340 3390 10350 3430
rect 10290 3380 10350 3390
rect 6870 2800 6930 2810
rect 6870 2760 6880 2800
rect 6880 2760 6920 2800
rect 6920 2760 6930 2800
rect 6870 2750 6930 2760
rect 8130 2750 8190 2810
rect 9390 2800 9450 2810
rect 9390 2760 9400 2800
rect 9400 2760 9440 2800
rect 9440 2760 9450 2800
rect 9390 2750 9450 2760
rect 8130 2600 8190 2620
rect 8130 2560 8140 2600
rect 8140 2560 8180 2600
rect 8180 2560 8190 2600
rect 6050 2500 6110 2510
rect 6050 2460 6060 2500
rect 6060 2460 6100 2500
rect 6100 2460 6110 2500
rect 6050 2450 6110 2460
rect 6210 2500 6270 2510
rect 6210 2460 6220 2500
rect 6220 2460 6260 2500
rect 6260 2460 6270 2500
rect 6210 2450 6270 2460
rect 6370 2500 6430 2510
rect 6370 2460 6380 2500
rect 6380 2460 6420 2500
rect 6420 2460 6430 2500
rect 6370 2450 6430 2460
rect 6530 2500 6590 2510
rect 6530 2460 6540 2500
rect 6540 2460 6580 2500
rect 6580 2460 6590 2500
rect 6530 2450 6590 2460
rect 6690 2500 6750 2510
rect 6690 2460 6700 2500
rect 6700 2460 6740 2500
rect 6740 2460 6750 2500
rect 6690 2450 6750 2460
rect 6850 2500 6910 2510
rect 6850 2460 6860 2500
rect 6860 2460 6900 2500
rect 6900 2460 6910 2500
rect 6850 2450 6910 2460
rect 7010 2500 7070 2510
rect 7010 2460 7020 2500
rect 7020 2460 7060 2500
rect 7060 2460 7070 2500
rect 7010 2450 7070 2460
rect 7170 2500 7230 2510
rect 7170 2460 7180 2500
rect 7180 2460 7220 2500
rect 7220 2460 7230 2500
rect 7170 2450 7230 2460
rect 7330 2500 7390 2510
rect 7330 2460 7340 2500
rect 7340 2460 7380 2500
rect 7380 2460 7390 2500
rect 7330 2450 7390 2460
rect 7490 2500 7550 2510
rect 7490 2460 7500 2500
rect 7500 2460 7540 2500
rect 7540 2460 7550 2500
rect 7490 2450 7550 2460
rect 7650 2500 7710 2510
rect 7650 2460 7660 2500
rect 7660 2460 7700 2500
rect 7700 2460 7710 2500
rect 7650 2450 7710 2460
rect 7810 2500 7870 2510
rect 7810 2460 7820 2500
rect 7820 2460 7860 2500
rect 7860 2460 7870 2500
rect 7810 2450 7870 2460
rect 7970 2500 8030 2510
rect 7970 2460 7980 2500
rect 7980 2460 8020 2500
rect 8020 2460 8030 2500
rect 7970 2450 8030 2460
rect 8130 2500 8190 2510
rect 8130 2460 8140 2500
rect 8140 2460 8180 2500
rect 8180 2460 8190 2500
rect 8130 2450 8190 2460
rect 8290 2500 8350 2510
rect 8290 2460 8300 2500
rect 8300 2460 8340 2500
rect 8340 2460 8350 2500
rect 8290 2450 8350 2460
rect 8450 2500 8510 2510
rect 8450 2460 8460 2500
rect 8460 2460 8500 2500
rect 8500 2460 8510 2500
rect 8450 2450 8510 2460
rect 8610 2500 8670 2510
rect 8610 2460 8620 2500
rect 8620 2460 8660 2500
rect 8660 2460 8670 2500
rect 8610 2450 8670 2460
rect 8770 2500 8830 2510
rect 8770 2460 8780 2500
rect 8780 2460 8820 2500
rect 8820 2460 8830 2500
rect 8770 2450 8830 2460
rect 8930 2500 8990 2510
rect 8930 2460 8940 2500
rect 8940 2460 8980 2500
rect 8980 2460 8990 2500
rect 8930 2450 8990 2460
rect 9090 2500 9150 2510
rect 9090 2460 9100 2500
rect 9100 2460 9140 2500
rect 9140 2460 9150 2500
rect 9090 2450 9150 2460
rect 9250 2500 9310 2510
rect 9250 2460 9260 2500
rect 9260 2460 9300 2500
rect 9300 2460 9310 2500
rect 9250 2450 9310 2460
rect 9410 2500 9470 2510
rect 9410 2460 9420 2500
rect 9420 2460 9460 2500
rect 9460 2460 9470 2500
rect 9410 2450 9470 2460
rect 9570 2500 9630 2510
rect 9570 2460 9580 2500
rect 9580 2460 9620 2500
rect 9620 2460 9630 2500
rect 9570 2450 9630 2460
rect 9730 2500 9790 2510
rect 9730 2460 9740 2500
rect 9740 2460 9780 2500
rect 9780 2460 9790 2500
rect 9730 2450 9790 2460
rect 9890 2500 9950 2510
rect 9890 2460 9900 2500
rect 9900 2460 9940 2500
rect 9940 2460 9950 2500
rect 9890 2450 9950 2460
rect 10050 2500 10110 2510
rect 10050 2460 10060 2500
rect 10060 2460 10100 2500
rect 10100 2460 10110 2500
rect 10050 2450 10110 2460
rect 5970 2330 6030 2340
rect 5970 2290 5980 2330
rect 5980 2290 6020 2330
rect 6020 2290 6030 2330
rect 5970 2280 6030 2290
rect 10280 2330 10340 2340
rect 10280 2290 10290 2330
rect 10290 2290 10330 2330
rect 10330 2290 10340 2330
rect 10280 2280 10340 2290
rect 6340 2040 6400 2100
rect 8130 2040 8190 2100
rect 9920 2040 9980 2100
rect 5800 1950 5860 1960
rect 5800 1910 5810 1950
rect 5810 1910 5850 1950
rect 5850 1910 5860 1950
rect 5800 1900 5860 1910
rect 6160 1950 6220 1960
rect 6160 1910 6170 1950
rect 6170 1910 6210 1950
rect 6210 1910 6220 1950
rect 6160 1900 6220 1910
rect 6520 1950 6580 1960
rect 6520 1910 6530 1950
rect 6530 1910 6570 1950
rect 6570 1910 6580 1950
rect 6520 1900 6580 1910
rect 7590 1950 7650 1960
rect 7590 1910 7600 1950
rect 7600 1910 7640 1950
rect 7640 1910 7650 1950
rect 7590 1900 7650 1910
rect 7950 1950 8010 1960
rect 7950 1910 7960 1950
rect 7960 1910 8000 1950
rect 8000 1910 8010 1950
rect 7950 1900 8010 1910
rect 8310 1950 8370 1960
rect 8310 1910 8320 1950
rect 8320 1910 8360 1950
rect 8360 1910 8370 1950
rect 8310 1900 8370 1910
rect 8670 1950 8730 1960
rect 8670 1910 8680 1950
rect 8680 1910 8720 1950
rect 8720 1910 8730 1950
rect 8670 1900 8730 1910
rect 9740 1950 9800 1960
rect 9740 1910 9750 1950
rect 9750 1910 9790 1950
rect 9790 1910 9800 1950
rect 9740 1900 9800 1910
rect 10100 1950 10160 1960
rect 10100 1910 10110 1950
rect 10110 1910 10150 1950
rect 10150 1910 10160 1950
rect 10100 1900 10160 1910
rect 10460 1950 10520 1960
rect 10460 1910 10470 1950
rect 10470 1910 10510 1950
rect 10510 1910 10520 1950
rect 10460 1900 10520 1910
rect 7000 1780 7060 1790
rect 7000 1740 7010 1780
rect 7010 1740 7050 1780
rect 7050 1740 7060 1780
rect 7000 1730 7060 1740
rect 7110 1780 7170 1790
rect 7110 1740 7120 1780
rect 7120 1740 7160 1780
rect 7160 1740 7170 1780
rect 7110 1730 7170 1740
rect 9150 1780 9210 1790
rect 9150 1740 9160 1780
rect 9160 1740 9200 1780
rect 9200 1740 9210 1780
rect 9150 1730 9210 1740
rect 9260 1780 9320 1790
rect 9260 1740 9270 1780
rect 9270 1740 9310 1780
rect 9310 1740 9320 1780
rect 9260 1730 9320 1740
rect 10940 1780 11000 1790
rect 10940 1740 10950 1780
rect 10950 1740 10990 1780
rect 10990 1740 11000 1780
rect 10940 1730 11000 1740
rect 5620 1610 5680 1620
rect 5620 1570 5630 1610
rect 5630 1570 5670 1610
rect 5670 1570 5680 1610
rect 5620 1560 5680 1570
rect 6340 1610 6400 1620
rect 6340 1570 6350 1610
rect 6350 1570 6390 1610
rect 6390 1570 6400 1610
rect 6340 1560 6400 1570
rect 8130 1610 8190 1620
rect 8130 1570 8140 1610
rect 8140 1570 8180 1610
rect 8180 1570 8190 1610
rect 8130 1560 8190 1570
rect 8490 1610 8550 1620
rect 8490 1570 8500 1610
rect 8500 1570 8540 1610
rect 8540 1570 8550 1610
rect 8490 1560 8550 1570
rect 8850 1610 8910 1620
rect 8850 1570 8860 1610
rect 8860 1570 8900 1610
rect 8900 1570 8910 1610
rect 8850 1560 8910 1570
rect 9920 1610 9980 1620
rect 9920 1570 9930 1610
rect 9930 1570 9970 1610
rect 9970 1570 9980 1610
rect 9920 1560 9980 1570
rect 10640 1610 10700 1620
rect 10640 1570 10650 1610
rect 10650 1570 10690 1610
rect 10690 1570 10700 1610
rect 10640 1560 10700 1570
rect 5120 1360 5180 1420
rect 5980 1450 6040 1510
rect 6700 1450 6760 1510
rect 7500 1360 7560 1420
rect 8130 1450 8190 1510
rect 9560 1450 9620 1510
rect 10280 1450 10340 1510
<< metal2 >>
rect -390 10680 -310 10690
rect -390 10620 -380 10680
rect -320 10620 -310 10680
rect -390 10610 -310 10620
rect 11500 10680 11580 10690
rect 11500 10620 11510 10680
rect 11570 10620 11580 10680
rect 11500 10610 11580 10620
rect -220 7750 -140 7760
rect -220 7690 -210 7750
rect -150 7740 -140 7750
rect 2700 7750 2780 7760
rect 2700 7740 2710 7750
rect -150 7700 2710 7740
rect -150 7690 -140 7700
rect -220 7680 -140 7690
rect 2700 7690 2710 7700
rect 2770 7690 2780 7750
rect 2700 7680 2780 7690
rect 8880 7690 8960 7700
rect 8880 7630 8890 7690
rect 8950 7680 8960 7690
rect 11500 7690 11580 7700
rect 11500 7680 11510 7690
rect 8950 7640 11510 7680
rect 8950 7630 8960 7640
rect 8880 7620 8960 7630
rect 11500 7630 11510 7640
rect 11570 7630 11580 7690
rect 11500 7620 11580 7630
rect -30 7590 50 7600
rect -30 7530 -20 7590
rect 40 7580 50 7590
rect 1880 7590 1960 7600
rect 1880 7580 1890 7590
rect 40 7540 1890 7580
rect 40 7530 50 7540
rect -30 7520 50 7530
rect 1880 7530 1890 7540
rect 1950 7530 1960 7590
rect 1880 7520 1960 7530
rect 3270 7590 3370 7610
rect 5020 7600 5100 7610
rect 5020 7590 5030 7600
rect 3270 7530 3290 7590
rect 3350 7550 5030 7590
rect 3350 7530 3370 7550
rect 5020 7540 5030 7550
rect 5090 7540 5100 7600
rect 5020 7530 5100 7540
rect 9600 7590 9680 7600
rect 9600 7530 9610 7590
rect 9670 7580 9680 7590
rect 10270 7590 10370 7610
rect 10270 7580 10290 7590
rect 9670 7540 10290 7580
rect 9670 7530 9680 7540
rect 3270 7510 3370 7530
rect 9600 7520 9680 7530
rect 10270 7530 10290 7540
rect 10350 7530 10370 7590
rect 10270 7510 10370 7530
rect -120 7480 -40 7490
rect -120 7420 -110 7480
rect -50 7470 -40 7480
rect 5380 7480 5460 7490
rect 5380 7470 5390 7480
rect -50 7430 5390 7470
rect -50 7420 -40 7430
rect -120 7410 -40 7420
rect 5380 7420 5390 7430
rect 5450 7420 5460 7480
rect 5380 7410 5460 7420
rect 6770 7480 6870 7500
rect 6770 7420 6790 7480
rect 6850 7470 6870 7480
rect 9510 7480 9590 7490
rect 9510 7470 9520 7480
rect 6850 7430 9520 7470
rect 6850 7420 6870 7430
rect 6770 7400 6870 7420
rect 9510 7420 9520 7430
rect 9580 7420 9590 7480
rect 9510 7410 9590 7420
rect 2510 7380 2590 7390
rect 2510 7320 2520 7380
rect 2580 7370 2590 7380
rect 9020 7380 9100 7390
rect 9020 7370 9030 7380
rect 2580 7330 9030 7370
rect 2580 7320 2590 7330
rect 2510 7310 2590 7320
rect 9020 7320 9030 7330
rect 9090 7320 9100 7380
rect 9020 7310 9100 7320
rect 140 7280 220 7290
rect 140 7220 150 7280
rect 210 7270 220 7280
rect 5110 7280 5190 7290
rect 5110 7270 5120 7280
rect 210 7230 5120 7270
rect 210 7220 220 7230
rect 140 7210 220 7220
rect 5110 7220 5120 7230
rect 5180 7220 5190 7280
rect 5110 7210 5190 7220
rect 6240 7270 6320 7280
rect 6240 7210 6250 7270
rect 6310 7260 6320 7270
rect 6310 7220 12200 7260
rect 6310 7210 6320 7220
rect 6240 7200 6320 7210
rect 5880 7180 5960 7190
rect 132 7110 142 7180
rect 212 7110 222 7180
rect 5880 7120 5890 7180
rect 5950 7170 5960 7180
rect 7940 7180 8020 7190
rect 7940 7170 7950 7180
rect 5950 7130 7950 7170
rect 5950 7120 5960 7130
rect 5880 7110 5960 7120
rect 7940 7120 7950 7130
rect 8010 7170 8020 7180
rect 8300 7180 8380 7190
rect 8300 7170 8310 7180
rect 8010 7130 8310 7170
rect 8010 7120 8020 7130
rect 7940 7110 8020 7120
rect 8300 7120 8310 7130
rect 8370 7170 8380 7180
rect 9420 7180 9500 7190
rect 9420 7170 9430 7180
rect 8370 7130 9430 7170
rect 8370 7120 8380 7130
rect 8300 7110 8380 7120
rect 9420 7120 9430 7130
rect 9490 7170 9500 7180
rect 10360 7180 10440 7190
rect 10360 7170 10370 7180
rect 9490 7130 10370 7170
rect 9490 7120 9500 7130
rect 9420 7110 9500 7120
rect 10360 7120 10370 7130
rect 10430 7120 10440 7180
rect 10360 7110 10440 7120
rect 5340 7060 5420 7070
rect -220 7050 -140 7060
rect -220 6990 -210 7050
rect -150 7040 -140 7050
rect 132 7040 142 7060
rect -150 7000 142 7040
rect -150 6990 -140 7000
rect 132 6990 142 7000
rect 212 6990 222 7060
rect 5340 7000 5350 7060
rect 5410 7050 5420 7060
rect 5700 7060 5780 7070
rect 5700 7050 5710 7060
rect 5410 7010 5710 7050
rect 5410 7000 5420 7010
rect 5340 6990 5420 7000
rect 5700 7000 5710 7010
rect 5770 7050 5780 7060
rect 6060 7060 6140 7070
rect 6060 7050 6070 7060
rect 5770 7010 6070 7050
rect 5770 7000 5780 7010
rect 5700 6990 5780 7000
rect 6060 7000 6070 7010
rect 6130 7050 6140 7060
rect 6420 7060 6500 7070
rect 6420 7050 6430 7060
rect 6130 7010 6430 7050
rect 6130 7000 6140 7010
rect 6060 6990 6140 7000
rect 6420 7000 6430 7010
rect 6490 7050 6500 7060
rect 7040 7060 7120 7070
rect 7040 7050 7050 7060
rect 6490 7010 7050 7050
rect 6490 7000 6500 7010
rect 6420 6990 6500 7000
rect 7040 7000 7050 7010
rect 7110 7050 7120 7060
rect 7400 7060 7480 7070
rect 7400 7050 7410 7060
rect 7110 7010 7410 7050
rect 7110 7000 7120 7010
rect 7040 6990 7120 7000
rect 7400 7000 7410 7010
rect 7470 7050 7480 7060
rect 7760 7060 7840 7070
rect 7760 7050 7770 7060
rect 7470 7010 7770 7050
rect 7470 7000 7480 7010
rect 7400 6990 7480 7000
rect 7760 7000 7770 7010
rect 7830 7050 7840 7060
rect 8120 7060 8200 7070
rect 8120 7050 8130 7060
rect 7830 7010 8130 7050
rect 7830 7000 7840 7010
rect 7760 6990 7840 7000
rect 8120 7000 8130 7010
rect 8190 7050 8200 7060
rect 8480 7060 8560 7070
rect 8480 7050 8490 7060
rect 8190 7010 8490 7050
rect 8190 7000 8200 7010
rect 8120 6990 8200 7000
rect 8480 7000 8490 7010
rect 8550 7050 8560 7060
rect 8840 7060 8920 7070
rect 8840 7050 8850 7060
rect 8550 7010 8850 7050
rect 8550 7000 8560 7010
rect 8480 6990 8560 7000
rect 8840 7000 8850 7010
rect 8910 7050 8920 7060
rect 9200 7060 9280 7070
rect 9200 7050 9210 7060
rect 8910 7010 9210 7050
rect 8910 7000 8920 7010
rect 8840 6990 8920 7000
rect 9200 7000 9210 7010
rect 9270 7050 9280 7060
rect 9820 7060 9900 7070
rect 9820 7050 9830 7060
rect 9270 7010 9830 7050
rect 9270 7000 9280 7010
rect 9200 6990 9280 7000
rect 9820 7000 9830 7010
rect 9890 7050 9900 7060
rect 10180 7060 10260 7070
rect 10180 7050 10190 7060
rect 9890 7010 10190 7050
rect 9890 7000 9900 7010
rect 9820 6990 9900 7000
rect 10180 7000 10190 7010
rect 10250 7050 10260 7060
rect 10540 7060 10620 7070
rect 10540 7050 10550 7060
rect 10250 7010 10550 7050
rect 10250 7000 10260 7010
rect 10180 6990 10260 7000
rect 10540 7000 10550 7010
rect 10610 7050 10620 7060
rect 10900 7060 10980 7070
rect 10900 7050 10910 7060
rect 10610 7010 10910 7050
rect 10610 7000 10620 7010
rect 10540 6990 10620 7000
rect 10900 7000 10910 7010
rect 10970 7050 10980 7060
rect 11500 7060 11580 7070
rect 11500 7050 11510 7060
rect 10970 7010 11510 7050
rect 10970 7000 10980 7010
rect 10900 6990 10980 7000
rect 11500 7000 11510 7010
rect 11570 7000 11580 7060
rect 11500 6990 11580 7000
rect -220 6980 -140 6990
rect 2702 6840 2712 6910
rect 2782 6840 2792 6910
rect 140 6750 220 6760
rect 140 6690 150 6750
rect 210 6740 220 6750
rect 2510 6750 2590 6760
rect 2510 6740 2520 6750
rect 210 6700 2520 6740
rect 210 6690 220 6700
rect 140 6680 220 6690
rect 2510 6690 2520 6700
rect 2580 6690 2590 6750
rect 2702 6720 2712 6790
rect 2782 6720 2792 6790
rect 5520 6720 5600 6730
rect 2510 6680 2590 6690
rect 5520 6660 5530 6720
rect 5590 6710 5600 6720
rect 5880 6720 5960 6730
rect 5880 6710 5890 6720
rect 5590 6670 5890 6710
rect 5590 6660 5600 6670
rect 5520 6650 5600 6660
rect 5880 6660 5890 6670
rect 5950 6710 5960 6720
rect 6240 6720 6320 6730
rect 6240 6710 6250 6720
rect 5950 6670 6250 6710
rect 5950 6660 5960 6670
rect 5880 6650 5960 6660
rect 6240 6660 6250 6670
rect 6310 6660 6320 6720
rect 6240 6650 6320 6660
rect 7580 6720 7660 6730
rect 7580 6660 7590 6720
rect 7650 6710 7660 6720
rect 7940 6720 8020 6730
rect 7940 6710 7950 6720
rect 7650 6670 7950 6710
rect 7650 6660 7660 6670
rect 7580 6650 7660 6660
rect 7940 6660 7950 6670
rect 8010 6710 8020 6720
rect 8300 6720 8380 6730
rect 8300 6710 8310 6720
rect 8010 6670 8310 6710
rect 8010 6660 8020 6670
rect 7940 6650 8020 6660
rect 8300 6660 8310 6670
rect 8370 6710 8380 6720
rect 8660 6720 8740 6730
rect 8660 6710 8670 6720
rect 8370 6670 8670 6710
rect 8370 6660 8380 6670
rect 8300 6650 8380 6660
rect 8660 6660 8670 6670
rect 8730 6660 8740 6720
rect 8660 6650 8740 6660
rect 10000 6720 10080 6730
rect 10000 6660 10010 6720
rect 10070 6710 10080 6720
rect 10360 6720 10440 6730
rect 10360 6710 10370 6720
rect 10070 6670 10370 6710
rect 10070 6660 10080 6670
rect 10000 6650 10080 6660
rect 10360 6660 10370 6670
rect 10430 6710 10440 6720
rect 10720 6720 10800 6730
rect 10720 6710 10730 6720
rect 10430 6670 10730 6710
rect 10430 6660 10440 6670
rect 10360 6650 10440 6660
rect 10720 6660 10730 6670
rect 10790 6710 10800 6720
rect 10790 6670 12200 6710
rect 10790 6660 10800 6670
rect 10720 6650 10800 6660
rect 132 6580 142 6650
rect 212 6580 222 6650
rect 9420 6630 9500 6640
rect 2370 6580 2450 6590
rect -220 6520 -140 6530
rect -220 6460 -210 6520
rect -150 6510 -140 6520
rect 132 6510 142 6530
rect -150 6470 142 6510
rect -150 6460 -140 6470
rect 132 6460 142 6470
rect 212 6460 222 6530
rect 2370 6520 2380 6580
rect 2440 6570 2450 6580
rect 2580 6580 2660 6590
rect 2580 6570 2590 6580
rect 2440 6530 2590 6570
rect 2440 6520 2450 6530
rect 2370 6510 2450 6520
rect 2580 6520 2590 6530
rect 2650 6520 2660 6580
rect 9420 6570 9430 6630
rect 9490 6620 9500 6630
rect 9490 6610 10020 6620
rect 9490 6580 9950 6610
rect 9490 6570 9500 6580
rect 9420 6560 9500 6570
rect 9940 6550 9950 6580
rect 10010 6550 10020 6610
rect 9940 6540 10020 6550
rect 9510 6520 9590 6530
rect 2580 6510 2660 6520
rect 5110 6510 5190 6520
rect -220 6450 -140 6460
rect 5110 6450 5120 6510
rect 5180 6500 5190 6510
rect 5220 6510 5300 6520
rect 5220 6500 5230 6510
rect 5180 6460 5230 6500
rect 5180 6450 5190 6460
rect 5110 6440 5190 6450
rect 5220 6450 5230 6460
rect 5290 6450 5300 6510
rect 9510 6460 9520 6520
rect 9580 6510 9590 6520
rect 10120 6520 10200 6530
rect 10120 6510 10130 6520
rect 9580 6470 10130 6510
rect 9580 6460 9590 6470
rect 9510 6450 9590 6460
rect 10120 6460 10130 6470
rect 10190 6460 10200 6520
rect 10120 6450 10200 6460
rect 5220 6440 5300 6450
rect -220 6390 -140 6400
rect -220 6330 -210 6390
rect -150 6380 -140 6390
rect 1190 6390 1270 6400
rect 1190 6380 1200 6390
rect -150 6340 1200 6380
rect -150 6330 -140 6340
rect -220 6320 -140 6330
rect 1190 6330 1200 6340
rect 1260 6330 1270 6390
rect 4840 6360 4850 6430
rect 4920 6410 4930 6430
rect 6120 6420 6200 6430
rect 6120 6410 6130 6420
rect 4920 6370 6130 6410
rect 4920 6360 4930 6370
rect 6120 6360 6130 6370
rect 6190 6360 6200 6420
rect 6120 6350 6200 6360
rect 9600 6410 9680 6420
rect 9600 6350 9610 6410
rect 9670 6400 9680 6410
rect 10030 6410 10110 6420
rect 10030 6400 10040 6410
rect 9670 6360 10040 6400
rect 9670 6350 9680 6360
rect 9600 6340 9680 6350
rect 10030 6350 10040 6360
rect 10100 6350 10110 6410
rect 10030 6340 10110 6350
rect 1190 6320 1270 6330
rect 5110 6330 5190 6340
rect 4840 6310 4930 6320
rect 4840 6240 4850 6310
rect 4920 6240 4930 6310
rect 5110 6270 5120 6330
rect 5180 6320 5190 6330
rect 7220 6330 7300 6340
rect 7220 6320 7230 6330
rect 5180 6280 7230 6320
rect 5180 6270 5190 6280
rect 5110 6260 5190 6270
rect 7220 6270 7230 6280
rect 7290 6270 7300 6330
rect 7220 6260 7300 6270
rect 9020 6320 9100 6330
rect 9020 6260 9030 6320
rect 9090 6310 9100 6320
rect 11230 6320 11310 6330
rect 11230 6310 11240 6320
rect 9090 6270 11240 6310
rect 9090 6260 9100 6270
rect 4840 6230 4930 6240
rect 8660 6250 8740 6260
rect 9020 6250 9100 6260
rect 11230 6260 11240 6270
rect 11300 6260 11310 6320
rect 11230 6250 11310 6260
rect 8660 6190 8670 6250
rect 8730 6220 8740 6250
rect 8730 6190 12200 6220
rect 8660 6180 12200 6190
rect 6500 6130 6580 6140
rect -120 6110 -40 6120
rect -120 6050 -110 6110
rect -50 6100 -40 6110
rect 522 6100 532 6120
rect -50 6060 532 6100
rect -50 6050 -40 6060
rect 522 6050 532 6060
rect 602 6050 612 6120
rect 1868 6050 1878 6120
rect 1948 6100 1958 6120
rect 2420 6110 2500 6120
rect 2420 6100 2430 6110
rect 1948 6060 2430 6100
rect 1948 6050 1958 6060
rect 2420 6050 2430 6060
rect 2490 6050 2500 6110
rect 6500 6100 6510 6130
rect -120 6040 -40 6050
rect 2420 6040 2500 6050
rect 5650 6070 6510 6100
rect 6570 6120 6580 6130
rect 6860 6130 6940 6140
rect 6860 6120 6870 6130
rect 6570 6080 6870 6120
rect 6570 6070 6580 6080
rect 5650 6060 6580 6070
rect 6860 6070 6870 6080
rect 6930 6120 6940 6130
rect 7220 6130 7300 6140
rect 7220 6120 7230 6130
rect 6930 6080 7230 6120
rect 6930 6070 6940 6080
rect 6860 6060 6940 6070
rect 7220 6070 7230 6080
rect 7290 6120 7300 6130
rect 7580 6130 7660 6140
rect 7580 6120 7590 6130
rect 7290 6080 7590 6120
rect 7290 6070 7300 6080
rect 7220 6060 7300 6070
rect 7580 6070 7590 6080
rect 7650 6120 7660 6130
rect 7940 6130 8020 6140
rect 7940 6120 7950 6130
rect 7650 6080 7950 6120
rect 7650 6070 7660 6080
rect 7580 6060 7660 6070
rect 7940 6070 7950 6080
rect 8010 6120 8020 6130
rect 8300 6130 8380 6140
rect 8300 6120 8310 6130
rect 8010 6080 8310 6120
rect 8010 6070 8020 6080
rect 7940 6060 8020 6070
rect 8300 6070 8310 6080
rect 8370 6120 8380 6130
rect 8660 6130 8740 6140
rect 8660 6120 8670 6130
rect 8370 6080 8670 6120
rect 8370 6070 8380 6080
rect 8300 6060 8380 6070
rect 8660 6070 8670 6080
rect 8730 6120 8740 6130
rect 9020 6130 9100 6140
rect 9020 6120 9030 6130
rect 8730 6080 9030 6120
rect 8730 6070 8740 6080
rect 8660 6060 8740 6070
rect 9020 6070 9030 6080
rect 9090 6120 9100 6130
rect 9380 6130 9460 6140
rect 9380 6120 9390 6130
rect 9090 6080 9390 6120
rect 9090 6070 9100 6080
rect 9020 6060 9100 6070
rect 9380 6070 9390 6080
rect 9450 6120 9460 6130
rect 9740 6130 9820 6140
rect 9740 6120 9750 6130
rect 9450 6080 9750 6120
rect 9450 6070 9460 6080
rect 9380 6060 9460 6070
rect 9740 6070 9750 6080
rect 9810 6120 9820 6130
rect 11500 6130 11580 6140
rect 11500 6120 11510 6130
rect 9810 6080 11510 6120
rect 9810 6070 9820 6080
rect 9740 6060 9820 6070
rect 10720 6060 10800 6080
rect 11500 6070 11510 6080
rect 11570 6070 11580 6130
rect 11500 6060 11580 6070
rect 5650 6050 5730 6060
rect 5650 5990 5660 6050
rect 5720 5990 5730 6050
rect 5650 5980 5730 5990
rect 10720 5990 10730 6060
rect 10790 5990 10800 6060
rect 10720 5980 10800 5990
rect 5650 5930 5730 5940
rect 2210 5900 2290 5910
rect 2210 5840 2220 5900
rect 2280 5890 2290 5900
rect 3032 5890 3042 5900
rect 2280 5850 3042 5890
rect 2280 5840 2290 5850
rect 2210 5830 2290 5840
rect 3032 5830 3042 5850
rect 3112 5830 3122 5900
rect 4430 5830 4440 5900
rect 4510 5880 4520 5900
rect 4840 5890 4920 5900
rect 4840 5880 4850 5890
rect 4510 5840 4850 5880
rect 4510 5830 4520 5840
rect 4840 5830 4850 5840
rect 4910 5830 4920 5890
rect 5650 5870 5660 5930
rect 5720 5920 5730 5930
rect 6120 5930 6200 5940
rect 6120 5920 6130 5930
rect 5720 5880 6130 5920
rect 5720 5870 5730 5880
rect 5650 5860 5730 5870
rect 6120 5870 6130 5880
rect 6190 5870 6200 5930
rect 6120 5860 6200 5870
rect 10720 5930 10800 5940
rect 10720 5870 10730 5930
rect 10790 5870 10800 5930
rect 10720 5860 10800 5870
rect 4840 5820 4920 5830
rect -30 5700 50 5710
rect -30 5640 -20 5700
rect 40 5680 50 5700
rect 522 5680 532 5700
rect 40 5640 532 5680
rect -30 5630 50 5640
rect 522 5630 532 5640
rect 602 5630 612 5700
rect 1868 5630 1878 5700
rect 1948 5680 1958 5700
rect 4930 5690 5010 5700
rect 4930 5680 4940 5690
rect 1948 5640 4940 5680
rect 1948 5630 1958 5640
rect 4930 5630 4940 5640
rect 5000 5630 5010 5690
rect 4930 5620 5010 5630
rect 2420 5600 2500 5610
rect 2420 5540 2430 5600
rect 2490 5590 2500 5600
rect 4750 5600 4830 5610
rect 4750 5590 4760 5600
rect 2490 5550 4760 5590
rect 2490 5540 2500 5550
rect 2420 5530 2500 5540
rect 4750 5540 4760 5550
rect 4820 5540 4830 5600
rect 4750 5530 4830 5540
rect 5520 5590 5600 5600
rect 5520 5530 5530 5590
rect 5590 5580 5600 5590
rect 5780 5590 5860 5600
rect 5780 5580 5790 5590
rect 5590 5540 5790 5580
rect 5590 5530 5600 5540
rect 5520 5520 5600 5530
rect 5780 5530 5790 5540
rect 5850 5580 5860 5590
rect 6240 5590 6320 5600
rect 6240 5580 6250 5590
rect 5850 5540 6250 5580
rect 5850 5530 5860 5540
rect 5780 5520 5860 5530
rect 6240 5530 6250 5540
rect 6310 5530 6320 5590
rect 6240 5520 6320 5530
rect 10520 5590 10600 5600
rect 10520 5530 10530 5590
rect 10590 5580 10600 5590
rect 10920 5590 11000 5600
rect 10920 5580 10930 5590
rect 10590 5540 10930 5580
rect 10590 5530 10600 5540
rect 10520 5520 10600 5530
rect 10920 5530 10930 5540
rect 10990 5580 11000 5590
rect 10990 5540 12200 5580
rect 10990 5530 11000 5540
rect 10920 5520 11000 5530
rect 4840 5390 4920 5400
rect 4840 5330 4850 5390
rect 4910 5380 4920 5390
rect 7760 5390 7840 5400
rect 7760 5380 7770 5390
rect 4910 5340 7770 5380
rect 4910 5330 4920 5340
rect 4840 5320 4920 5330
rect 7760 5330 7770 5340
rect 7830 5380 7840 5390
rect 8480 5390 8560 5400
rect 8480 5380 8490 5390
rect 7830 5340 8490 5380
rect 7830 5330 7840 5340
rect 7760 5320 7840 5330
rect 8480 5330 8490 5340
rect 8550 5330 8560 5390
rect 8480 5320 8560 5330
rect 10120 5300 10200 5310
rect 4660 5280 4740 5290
rect 4660 5220 4670 5280
rect 4730 5270 4740 5280
rect 6120 5280 6200 5290
rect 6120 5270 6130 5280
rect 4730 5230 6130 5270
rect 4730 5220 4740 5230
rect 4660 5210 4740 5220
rect 6120 5220 6130 5230
rect 6190 5270 6200 5280
rect 7400 5280 7480 5290
rect 7400 5270 7410 5280
rect 6190 5230 7410 5270
rect 6190 5220 6200 5230
rect 6120 5210 6200 5220
rect 7400 5220 7410 5230
rect 7470 5270 7480 5280
rect 8840 5280 8920 5290
rect 8840 5270 8850 5280
rect 7470 5230 8850 5270
rect 7470 5220 7480 5230
rect 7400 5210 7480 5220
rect 8840 5220 8850 5230
rect 8910 5220 8920 5280
rect 10120 5240 10130 5300
rect 10190 5290 10200 5300
rect 11050 5300 11130 5310
rect 11050 5290 11060 5300
rect 10190 5250 11060 5290
rect 10190 5240 10200 5250
rect 10120 5230 10200 5240
rect 11050 5240 11060 5250
rect 11120 5240 11130 5300
rect 11050 5230 11130 5240
rect 8840 5210 8920 5220
rect 4550 5190 4630 5200
rect 4550 5130 4560 5190
rect 4620 5180 4630 5190
rect 5650 5190 5730 5200
rect 5650 5180 5660 5190
rect 4620 5140 5660 5180
rect 4620 5130 4630 5140
rect 4550 5120 4630 5130
rect 5650 5130 5660 5140
rect 5720 5180 5730 5190
rect 7040 5190 7120 5200
rect 7040 5180 7050 5190
rect 5720 5140 7050 5180
rect 5720 5130 5730 5140
rect 5650 5120 5730 5130
rect 7040 5130 7050 5140
rect 7110 5180 7120 5190
rect 9200 5190 9280 5200
rect 9200 5180 9210 5190
rect 7110 5140 9210 5180
rect 7110 5130 7120 5140
rect 7040 5120 7120 5130
rect 9200 5130 9210 5140
rect 9270 5130 9280 5190
rect 9200 5120 9280 5130
rect 9380 5190 9460 5200
rect 9380 5130 9390 5190
rect 9450 5180 9460 5190
rect 10030 5190 10110 5200
rect 10030 5180 10040 5190
rect 9450 5140 10040 5180
rect 9450 5130 9460 5140
rect 9380 5120 9460 5130
rect 10030 5130 10040 5140
rect 10100 5130 10110 5190
rect 10030 5120 10110 5130
rect 5220 5100 5300 5110
rect 5220 5040 5230 5100
rect 5290 5090 5300 5100
rect 6680 5100 6760 5110
rect 6680 5090 6690 5100
rect 5290 5050 6690 5090
rect 5290 5040 5300 5050
rect 5220 5030 5300 5040
rect 6680 5040 6690 5050
rect 6750 5090 6760 5100
rect 8120 5100 8200 5110
rect 8120 5090 8130 5100
rect 6750 5050 8130 5090
rect 6750 5040 6760 5050
rect 6680 5030 6760 5040
rect 8120 5040 8130 5050
rect 8190 5090 8200 5100
rect 9560 5100 9640 5110
rect 9560 5090 9570 5100
rect 8190 5050 9570 5090
rect 8190 5040 8200 5050
rect 8120 5030 8200 5040
rect 9560 5040 9570 5050
rect 9630 5090 9640 5100
rect 11140 5100 11220 5110
rect 11140 5090 11150 5100
rect 9630 5050 11150 5090
rect 9630 5040 9640 5050
rect 9560 5030 9640 5040
rect 11140 5040 11150 5050
rect 11210 5040 11220 5100
rect 11140 5030 11220 5040
rect 4750 5000 4830 5010
rect 4750 4940 4760 5000
rect 4820 4990 4830 5000
rect 8560 5000 8640 5010
rect 8560 4990 8570 5000
rect 4820 4950 8570 4990
rect 4820 4940 4830 4950
rect 4750 4930 4830 4940
rect 8560 4940 8570 4950
rect 8630 4990 8640 5000
rect 9940 5000 10020 5010
rect 9940 4990 9950 5000
rect 8630 4950 9950 4990
rect 8630 4940 8640 4950
rect 8560 4930 8640 4940
rect 9940 4940 9950 4950
rect 10010 4990 10020 5000
rect 10720 5000 10800 5010
rect 10720 4990 10730 5000
rect 10010 4950 10730 4990
rect 10010 4940 10020 4950
rect 9940 4930 10020 4940
rect 10720 4940 10730 4950
rect 10790 4940 10800 5000
rect 10720 4930 10800 4940
rect 5640 4870 5720 4880
rect 5640 4810 5650 4870
rect 5710 4860 5720 4870
rect 5880 4870 5960 4880
rect 5880 4860 5890 4870
rect 5710 4820 5890 4860
rect 5710 4810 5720 4820
rect 5640 4800 5720 4810
rect 5880 4810 5890 4820
rect 5950 4860 5960 4870
rect 6120 4870 6200 4880
rect 6120 4860 6130 4870
rect 5950 4820 6130 4860
rect 5950 4810 5960 4820
rect 5880 4800 5960 4810
rect 6120 4810 6130 4820
rect 6190 4860 6200 4870
rect 6360 4870 6440 4880
rect 6360 4860 6370 4870
rect 6190 4820 6370 4860
rect 6190 4810 6200 4820
rect 6120 4800 6200 4810
rect 6360 4810 6370 4820
rect 6430 4860 6440 4870
rect 6600 4870 6680 4880
rect 6600 4860 6610 4870
rect 6430 4820 6610 4860
rect 6430 4810 6440 4820
rect 6360 4800 6440 4810
rect 6600 4810 6610 4820
rect 6670 4860 6680 4870
rect 6840 4870 6920 4880
rect 6840 4860 6850 4870
rect 6670 4820 6850 4860
rect 6670 4810 6680 4820
rect 6600 4800 6680 4810
rect 6840 4810 6850 4820
rect 6910 4860 6920 4870
rect 7080 4870 7160 4880
rect 7080 4860 7090 4870
rect 6910 4820 7090 4860
rect 6910 4810 6920 4820
rect 6840 4800 6920 4810
rect 7080 4810 7090 4820
rect 7150 4860 7160 4870
rect 7320 4870 7400 4880
rect 7320 4860 7330 4870
rect 7150 4820 7330 4860
rect 7150 4810 7160 4820
rect 7080 4800 7160 4810
rect 7320 4810 7330 4820
rect 7390 4860 7400 4870
rect 7560 4870 7640 4880
rect 7560 4860 7570 4870
rect 7390 4820 7570 4860
rect 7390 4810 7400 4820
rect 7320 4800 7400 4810
rect 7560 4810 7570 4820
rect 7630 4860 7640 4870
rect 8680 4870 8760 4880
rect 8680 4860 8690 4870
rect 7630 4820 8690 4860
rect 7630 4810 7640 4820
rect 7560 4800 7640 4810
rect 8680 4810 8690 4820
rect 8750 4860 8760 4870
rect 8920 4870 9000 4880
rect 8920 4860 8930 4870
rect 8750 4820 8930 4860
rect 8750 4810 8760 4820
rect 8680 4800 8760 4810
rect 8920 4810 8930 4820
rect 8990 4860 9000 4870
rect 9160 4870 9240 4880
rect 9160 4860 9170 4870
rect 8990 4820 9170 4860
rect 8990 4810 9000 4820
rect 8920 4800 9000 4810
rect 9160 4810 9170 4820
rect 9230 4860 9240 4870
rect 9400 4870 9480 4880
rect 9400 4860 9410 4870
rect 9230 4820 9410 4860
rect 9230 4810 9240 4820
rect 9160 4800 9240 4810
rect 9400 4810 9410 4820
rect 9470 4860 9480 4870
rect 9640 4870 9720 4880
rect 9640 4860 9650 4870
rect 9470 4820 9650 4860
rect 9470 4810 9480 4820
rect 9400 4800 9480 4810
rect 9640 4810 9650 4820
rect 9710 4860 9720 4870
rect 9880 4870 9960 4880
rect 9880 4860 9890 4870
rect 9710 4820 9890 4860
rect 9710 4810 9720 4820
rect 9640 4800 9720 4810
rect 9880 4810 9890 4820
rect 9950 4860 9960 4870
rect 10120 4870 10200 4880
rect 10120 4860 10130 4870
rect 9950 4820 10130 4860
rect 9950 4810 9960 4820
rect 9880 4800 9960 4810
rect 10120 4810 10130 4820
rect 10190 4860 10200 4870
rect 10360 4870 10440 4880
rect 10360 4860 10370 4870
rect 10190 4820 10370 4860
rect 10190 4810 10200 4820
rect 10120 4800 10200 4810
rect 10360 4810 10370 4820
rect 10430 4860 10440 4870
rect 10600 4870 10680 4880
rect 10600 4860 10610 4870
rect 10430 4820 10610 4860
rect 10430 4810 10440 4820
rect 10360 4800 10440 4810
rect 10600 4810 10610 4820
rect 10670 4860 10680 4870
rect 11500 4870 11580 4880
rect 11500 4860 11510 4870
rect 10670 4820 11510 4860
rect 10670 4810 10680 4820
rect 10600 4800 10680 4810
rect 11500 4810 11510 4820
rect 11570 4810 11580 4870
rect 11500 4800 11580 4810
rect 4930 4750 5010 4760
rect 4930 4690 4940 4750
rect 5000 4740 5010 4750
rect 5520 4750 5600 4760
rect 5520 4740 5530 4750
rect 5000 4700 5530 4740
rect 5000 4690 5010 4700
rect 4930 4680 5010 4690
rect 5520 4690 5530 4700
rect 5590 4740 5600 4750
rect 6240 4750 6320 4760
rect 6240 4740 6250 4750
rect 5590 4700 6250 4740
rect 5590 4690 5600 4700
rect 5520 4680 5600 4690
rect 6240 4690 6250 4700
rect 6310 4740 6320 4750
rect 6960 4750 7040 4760
rect 6960 4740 6970 4750
rect 6310 4700 6970 4740
rect 6310 4690 6320 4700
rect 6240 4680 6320 4690
rect 6960 4690 6970 4700
rect 7030 4740 7040 4750
rect 7680 4750 7760 4760
rect 7680 4740 7690 4750
rect 7030 4700 7690 4740
rect 7030 4690 7040 4700
rect 6960 4680 7040 4690
rect 7680 4690 7690 4700
rect 7750 4740 7760 4750
rect 7940 4750 8020 4760
rect 7940 4740 7950 4750
rect 7750 4700 7950 4740
rect 7750 4690 7760 4700
rect 7680 4680 7760 4690
rect 7940 4690 7950 4700
rect 8010 4690 8020 4750
rect 7940 4680 8020 4690
rect 8300 4750 8380 4760
rect 8300 4690 8310 4750
rect 8370 4740 8380 4750
rect 8560 4750 8640 4760
rect 8560 4740 8570 4750
rect 8370 4700 8570 4740
rect 8370 4690 8380 4700
rect 8300 4680 8380 4690
rect 8560 4690 8570 4700
rect 8630 4740 8640 4750
rect 9280 4750 9360 4760
rect 9280 4740 9290 4750
rect 8630 4700 9290 4740
rect 8630 4690 8640 4700
rect 8560 4680 8640 4690
rect 9280 4690 9290 4700
rect 9350 4740 9360 4750
rect 10000 4750 10080 4760
rect 10000 4740 10010 4750
rect 9350 4700 10010 4740
rect 9350 4690 9360 4700
rect 9280 4680 9360 4690
rect 10000 4690 10010 4700
rect 10070 4740 10080 4750
rect 10720 4750 10800 4760
rect 10720 4740 10730 4750
rect 10070 4700 10730 4740
rect 10070 4690 10080 4700
rect 10000 4680 10080 4690
rect 10720 4690 10730 4700
rect 10790 4690 10800 4750
rect 10720 4680 10800 4690
rect 5760 4410 5840 4420
rect 5760 4350 5770 4410
rect 5830 4400 5840 4410
rect 6000 4400 6080 4420
rect 6480 4410 6560 4420
rect 6480 4400 6490 4410
rect 5830 4360 6490 4400
rect 5830 4350 5840 4360
rect 5760 4340 5840 4350
rect 6000 4340 6080 4360
rect 6480 4350 6490 4360
rect 6550 4400 6560 4410
rect 6720 4400 6800 4420
rect 7200 4410 7280 4420
rect 7200 4400 7210 4410
rect 6550 4360 7210 4400
rect 6550 4350 6560 4360
rect 6480 4340 6560 4350
rect 6720 4340 6800 4360
rect 7200 4350 7210 4360
rect 7270 4350 7280 4410
rect 7200 4340 7280 4350
rect 7440 4340 7520 4420
rect 8800 4340 8880 4420
rect 9040 4410 9120 4420
rect 9040 4350 9050 4410
rect 9110 4400 9120 4410
rect 9520 4400 9600 4420
rect 9760 4410 9840 4420
rect 9760 4400 9770 4410
rect 9110 4360 9770 4400
rect 9110 4350 9120 4360
rect 9040 4340 9120 4350
rect 9520 4340 9600 4360
rect 9760 4350 9770 4360
rect 9830 4400 9840 4410
rect 10240 4400 10320 4420
rect 10480 4410 10560 4420
rect 10480 4400 10490 4410
rect 9830 4360 10490 4400
rect 9830 4350 9840 4360
rect 9760 4340 9840 4350
rect 10240 4340 10320 4360
rect 10480 4350 10490 4360
rect 10550 4350 10560 4410
rect 10480 4340 10560 4350
rect 5020 4290 5100 4300
rect 5020 4230 5030 4290
rect 5090 4280 5100 4290
rect 5580 4290 5660 4300
rect 5580 4280 5590 4290
rect 5090 4240 5590 4280
rect 5090 4230 5100 4240
rect 5020 4220 5100 4230
rect 5580 4230 5590 4240
rect 5650 4280 5660 4290
rect 6000 4290 6080 4300
rect 6000 4280 6010 4290
rect 5650 4240 6010 4280
rect 5650 4230 5660 4240
rect 5580 4220 5660 4230
rect 6000 4230 6010 4240
rect 6070 4280 6080 4290
rect 6240 4290 6320 4300
rect 6240 4280 6250 4290
rect 6070 4240 6250 4280
rect 6070 4230 6080 4240
rect 6000 4220 6080 4230
rect 6240 4230 6250 4240
rect 6310 4280 6320 4290
rect 6720 4290 6800 4300
rect 6720 4280 6730 4290
rect 6310 4240 6730 4280
rect 6310 4230 6320 4240
rect 6240 4220 6320 4230
rect 6720 4230 6730 4240
rect 6790 4280 6800 4290
rect 6960 4290 7040 4300
rect 6960 4280 6970 4290
rect 6790 4240 6970 4280
rect 6790 4230 6800 4240
rect 6720 4220 6800 4230
rect 6960 4230 6970 4240
rect 7030 4280 7040 4290
rect 7440 4290 7520 4300
rect 7440 4280 7450 4290
rect 7030 4240 7450 4280
rect 7030 4230 7040 4240
rect 6960 4220 7040 4230
rect 7440 4230 7450 4240
rect 7510 4280 7520 4290
rect 7620 4290 7700 4300
rect 7620 4280 7630 4290
rect 7510 4240 7630 4280
rect 7510 4230 7520 4240
rect 7440 4220 7520 4230
rect 7620 4230 7630 4240
rect 7690 4230 7700 4290
rect 7620 4220 7700 4230
rect 8620 4290 8700 4300
rect 8620 4230 8630 4290
rect 8690 4280 8700 4290
rect 8800 4290 8880 4300
rect 8800 4280 8810 4290
rect 8690 4240 8810 4280
rect 8690 4230 8700 4240
rect 8620 4220 8700 4230
rect 8800 4230 8810 4240
rect 8870 4280 8880 4290
rect 9280 4290 9360 4300
rect 9280 4280 9290 4290
rect 8870 4240 9290 4280
rect 8870 4230 8880 4240
rect 8800 4220 8880 4230
rect 9280 4230 9290 4240
rect 9350 4280 9360 4290
rect 9520 4290 9600 4300
rect 9520 4280 9530 4290
rect 9350 4240 9530 4280
rect 9350 4230 9360 4240
rect 9280 4220 9360 4230
rect 9520 4230 9530 4240
rect 9590 4280 9600 4290
rect 10000 4290 10080 4300
rect 10000 4280 10010 4290
rect 9590 4240 10010 4280
rect 9590 4230 9600 4240
rect 9520 4220 9600 4230
rect 10000 4230 10010 4240
rect 10070 4280 10080 4290
rect 10240 4290 10320 4300
rect 10240 4280 10250 4290
rect 10070 4240 10250 4280
rect 10070 4230 10080 4240
rect 10000 4220 10080 4230
rect 10240 4230 10250 4240
rect 10310 4280 10320 4290
rect 10660 4290 10740 4300
rect 10660 4280 10670 4290
rect 10310 4240 10670 4280
rect 10310 4230 10320 4240
rect 10240 4220 10320 4230
rect 10660 4230 10670 4240
rect 10730 4280 10740 4290
rect 11050 4290 11130 4300
rect 11050 4280 11060 4290
rect 10730 4240 11060 4280
rect 10730 4230 10740 4240
rect 10660 4220 10740 4230
rect 11050 4230 11060 4240
rect 11120 4230 11130 4290
rect 11050 4220 11130 4230
rect 6500 4120 6580 4130
rect 4660 4090 4740 4100
rect 4660 4030 4670 4090
rect 4730 4080 4740 4090
rect 6380 4090 6460 4100
rect 6380 4080 6390 4090
rect 4730 4040 6390 4080
rect 4730 4030 4740 4040
rect 4660 4020 4740 4030
rect 6380 4030 6390 4040
rect 6450 4030 6460 4090
rect 6500 4060 6510 4120
rect 6570 4110 6580 4120
rect 6980 4120 7060 4130
rect 6980 4110 6990 4120
rect 6570 4070 6990 4110
rect 6570 4060 6580 4070
rect 6500 4050 6580 4060
rect 6980 4060 6990 4070
rect 7050 4110 7060 4120
rect 7460 4120 7540 4130
rect 7460 4110 7470 4120
rect 7050 4070 7470 4110
rect 7050 4060 7060 4070
rect 6980 4050 7060 4060
rect 7460 4060 7470 4070
rect 7530 4060 7540 4120
rect 7460 4050 7540 4060
rect 8780 4120 8860 4130
rect 8780 4060 8790 4120
rect 8850 4110 8860 4120
rect 9260 4120 9340 4130
rect 9260 4110 9270 4120
rect 8850 4070 9270 4110
rect 8850 4060 8860 4070
rect 8780 4050 8860 4060
rect 9260 4060 9270 4070
rect 9330 4110 9340 4120
rect 9740 4120 9820 4130
rect 9740 4110 9750 4120
rect 9330 4070 9750 4110
rect 9330 4060 9340 4070
rect 9260 4050 9340 4060
rect 9740 4060 9750 4070
rect 9810 4060 9820 4120
rect 9740 4050 9820 4060
rect 9860 4090 9940 4100
rect 6380 4020 6460 4030
rect 9860 4030 9870 4090
rect 9930 4080 9940 4090
rect 11140 4090 11220 4100
rect 11140 4080 11150 4090
rect 9930 4040 11150 4080
rect 9930 4030 9940 4040
rect 9860 4020 9940 4030
rect 11140 4030 11150 4040
rect 11210 4080 11220 4090
rect 11210 4040 12200 4080
rect 11210 4030 11220 4040
rect 11140 4020 11220 4030
rect 6260 4000 6340 4010
rect 6260 3940 6270 4000
rect 6330 3990 6340 4000
rect 6740 4000 6820 4010
rect 6740 3990 6750 4000
rect 6330 3950 6750 3990
rect 6330 3940 6340 3950
rect 6260 3930 6340 3940
rect 6740 3940 6750 3950
rect 6810 3990 6820 4000
rect 7220 4000 7300 4010
rect 7220 3990 7230 4000
rect 6810 3950 7230 3990
rect 6810 3940 6820 3950
rect 6740 3930 6820 3940
rect 7220 3940 7230 3950
rect 7290 3940 7300 4000
rect 7220 3930 7300 3940
rect 9020 4000 9100 4010
rect 9020 3940 9030 4000
rect 9090 3990 9100 4000
rect 9500 4000 9580 4010
rect 9500 3990 9510 4000
rect 9090 3950 9510 3990
rect 9090 3940 9100 3950
rect 9020 3930 9100 3940
rect 9500 3940 9510 3950
rect 9570 3990 9580 4000
rect 9980 4000 10060 4010
rect 9980 3990 9990 4000
rect 9570 3950 9990 3990
rect 9570 3940 9580 3950
rect 9500 3930 9580 3940
rect 9980 3940 9990 3950
rect 10050 3940 10060 4000
rect 9980 3930 10060 3940
rect 7580 3880 7660 3890
rect 7580 3820 7590 3880
rect 7650 3870 7660 3880
rect 8120 3880 8200 3890
rect 8120 3870 8130 3880
rect 7650 3830 8130 3870
rect 7650 3820 7660 3830
rect 7580 3810 7660 3820
rect 8120 3820 8130 3830
rect 8190 3870 8200 3880
rect 8660 3880 8740 3890
rect 8660 3870 8670 3880
rect 8190 3830 8670 3870
rect 8190 3820 8200 3830
rect 8120 3810 8200 3820
rect 8660 3820 8670 3830
rect 8730 3820 8740 3880
rect 8660 3810 8740 3820
rect 4840 3760 4920 3770
rect 4840 3700 4850 3760
rect 4910 3750 4920 3760
rect 6260 3760 6340 3770
rect 6260 3750 6270 3760
rect 4910 3710 6270 3750
rect 4910 3700 4920 3710
rect 4840 3690 4920 3700
rect 6260 3700 6270 3710
rect 6330 3700 6340 3760
rect 6260 3690 6340 3700
rect 9980 3760 10060 3770
rect 9980 3700 9990 3760
rect 10050 3750 10060 3760
rect 11230 3760 11310 3770
rect 11230 3750 11240 3760
rect 10050 3710 11240 3750
rect 10050 3700 10060 3710
rect 9980 3690 10060 3700
rect 11230 3700 11240 3710
rect 11300 3700 11310 3760
rect 11230 3690 11310 3700
rect 5780 3640 5860 3650
rect 5780 3580 5790 3640
rect 5850 3630 5860 3640
rect 6380 3640 6460 3650
rect 6380 3630 6390 3640
rect 5850 3590 6390 3630
rect 5850 3580 5860 3590
rect 5780 3570 5860 3580
rect 6380 3580 6390 3590
rect 6450 3630 6460 3640
rect 6620 3640 6700 3650
rect 6620 3630 6630 3640
rect 6450 3590 6630 3630
rect 6450 3580 6460 3590
rect 6380 3570 6460 3580
rect 6620 3580 6630 3590
rect 6690 3630 6700 3640
rect 6860 3640 6940 3650
rect 6860 3630 6870 3640
rect 6690 3590 6870 3630
rect 6690 3580 6700 3590
rect 6620 3570 6700 3580
rect 6860 3580 6870 3590
rect 6930 3630 6940 3640
rect 7100 3640 7180 3650
rect 7100 3630 7110 3640
rect 6930 3590 7110 3630
rect 6930 3580 6940 3590
rect 6860 3570 6940 3580
rect 7100 3580 7110 3590
rect 7170 3630 7180 3640
rect 7340 3640 7420 3650
rect 7340 3630 7350 3640
rect 7170 3590 7350 3630
rect 7170 3580 7180 3590
rect 7100 3570 7180 3580
rect 7340 3580 7350 3590
rect 7410 3580 7420 3640
rect 7340 3570 7420 3580
rect 8900 3640 8980 3650
rect 8900 3580 8910 3640
rect 8970 3630 8980 3640
rect 9140 3640 9220 3650
rect 9140 3630 9150 3640
rect 8970 3590 9150 3630
rect 8970 3580 8980 3590
rect 8900 3570 8980 3580
rect 9140 3580 9150 3590
rect 9210 3630 9220 3640
rect 9380 3640 9460 3650
rect 9380 3630 9390 3640
rect 9210 3590 9390 3630
rect 9210 3580 9220 3590
rect 9140 3570 9220 3580
rect 9380 3580 9390 3590
rect 9450 3630 9460 3640
rect 9620 3640 9700 3650
rect 9620 3630 9630 3640
rect 9450 3590 9630 3630
rect 9450 3580 9460 3590
rect 9380 3570 9460 3580
rect 9620 3580 9630 3590
rect 9690 3630 9700 3640
rect 9860 3640 9940 3650
rect 9860 3630 9870 3640
rect 9690 3590 9870 3630
rect 9690 3580 9700 3590
rect 9620 3570 9700 3580
rect 9860 3580 9870 3590
rect 9930 3630 9940 3640
rect 10460 3640 10540 3650
rect 10460 3630 10470 3640
rect 9930 3590 10470 3630
rect 9930 3580 9940 3590
rect 9860 3570 9940 3580
rect 10460 3580 10470 3590
rect 10530 3580 10540 3640
rect 10460 3570 10540 3580
rect -220 3440 -140 3450
rect -220 3380 -210 3440
rect -150 3380 -140 3440
rect -220 3370 -140 3380
rect -90 3440 -10 3450
rect -90 3380 -80 3440
rect -20 3380 -10 3440
rect 5960 3440 6040 3450
rect -90 3370 -10 3380
rect 2524 3420 2604 3430
rect 2524 3360 2540 3420
rect 2594 3410 2604 3420
rect 4660 3420 4740 3430
rect 4660 3410 4670 3420
rect 2594 3370 4670 3410
rect 2594 3360 2604 3370
rect 2524 3350 2604 3360
rect 4660 3360 4670 3370
rect 4730 3360 4740 3420
rect 5960 3380 5970 3440
rect 6030 3430 6040 3440
rect 6200 3440 6280 3450
rect 6200 3430 6210 3440
rect 6030 3390 6210 3430
rect 6030 3380 6040 3390
rect 5960 3370 6040 3380
rect 6200 3380 6210 3390
rect 6270 3430 6280 3440
rect 6440 3440 6520 3450
rect 6440 3430 6450 3440
rect 6270 3390 6450 3430
rect 6270 3380 6280 3390
rect 6200 3370 6280 3380
rect 6440 3380 6450 3390
rect 6510 3430 6520 3440
rect 6680 3440 6760 3450
rect 6680 3430 6690 3440
rect 6510 3390 6690 3430
rect 6510 3380 6520 3390
rect 6440 3370 6520 3380
rect 6680 3380 6690 3390
rect 6750 3430 6760 3440
rect 7160 3440 7240 3450
rect 7160 3430 7170 3440
rect 6750 3390 7170 3430
rect 6750 3380 6760 3390
rect 6680 3370 6760 3380
rect 7160 3380 7170 3390
rect 7230 3430 7240 3440
rect 7400 3440 7480 3450
rect 7400 3430 7410 3440
rect 7230 3390 7410 3430
rect 7230 3380 7240 3390
rect 7160 3370 7240 3380
rect 7400 3380 7410 3390
rect 7470 3430 7480 3440
rect 7640 3440 7720 3450
rect 7640 3430 7650 3440
rect 7470 3390 7650 3430
rect 7470 3380 7480 3390
rect 7400 3370 7480 3380
rect 7640 3380 7650 3390
rect 7710 3430 7720 3440
rect 8600 3440 8680 3450
rect 8600 3430 8610 3440
rect 7710 3390 8610 3430
rect 7710 3380 7720 3390
rect 7640 3370 7720 3380
rect 8600 3380 8610 3390
rect 8670 3430 8680 3440
rect 8840 3440 8920 3450
rect 8840 3430 8850 3440
rect 8670 3390 8850 3430
rect 8670 3380 8680 3390
rect 8600 3370 8680 3380
rect 8840 3380 8850 3390
rect 8910 3430 8920 3440
rect 9080 3440 9160 3450
rect 9080 3430 9090 3440
rect 8910 3390 9090 3430
rect 8910 3380 8920 3390
rect 8840 3370 8920 3380
rect 9080 3380 9090 3390
rect 9150 3430 9160 3440
rect 9560 3440 9640 3450
rect 9560 3430 9570 3440
rect 9150 3390 9570 3430
rect 9150 3380 9160 3390
rect 9080 3370 9160 3380
rect 9560 3380 9570 3390
rect 9630 3430 9640 3440
rect 9800 3440 9880 3450
rect 9800 3430 9810 3440
rect 9630 3390 9810 3430
rect 9630 3380 9640 3390
rect 9560 3370 9640 3380
rect 9800 3380 9810 3390
rect 9870 3430 9880 3440
rect 10040 3440 10120 3450
rect 10040 3430 10050 3440
rect 9870 3390 10050 3430
rect 9870 3380 9880 3390
rect 9800 3370 9880 3380
rect 10040 3380 10050 3390
rect 10110 3430 10120 3440
rect 10280 3440 10360 3450
rect 10280 3430 10290 3440
rect 10110 3390 10290 3430
rect 10110 3380 10120 3390
rect 10040 3370 10120 3380
rect 10280 3380 10290 3390
rect 10350 3430 10360 3440
rect 11500 3440 11580 3450
rect 11500 3430 11510 3440
rect 10350 3390 11510 3430
rect 10350 3380 10360 3390
rect 10280 3370 10360 3380
rect 11500 3380 11510 3390
rect 11570 3380 11580 3440
rect 11500 3370 11580 3380
rect 4660 3350 4740 3360
rect 6860 2810 6940 2820
rect 6860 2750 6870 2810
rect 6930 2800 6940 2810
rect 8120 2810 8200 2820
rect 8120 2800 8130 2810
rect 6930 2760 8130 2800
rect 6930 2750 6940 2760
rect 6860 2740 6940 2750
rect 8120 2750 8130 2760
rect 8190 2800 8200 2810
rect 9380 2810 9460 2820
rect 9380 2800 9390 2810
rect 8190 2760 9390 2800
rect 8190 2750 8200 2760
rect 8120 2740 8200 2750
rect 9380 2750 9390 2760
rect 9450 2800 9460 2810
rect 11330 2810 11410 2820
rect 11330 2800 11340 2810
rect 9450 2760 11340 2800
rect 9450 2750 9460 2760
rect 9380 2740 9460 2750
rect 11330 2750 11340 2760
rect 11400 2750 11410 2810
rect 11330 2740 11410 2750
rect 8120 2620 8200 2630
rect 8120 2560 8130 2620
rect 8190 2560 8200 2620
rect 8120 2550 8200 2560
rect 6040 2510 6120 2520
rect 6040 2450 6050 2510
rect 6110 2500 6120 2510
rect 6200 2510 6280 2520
rect 6200 2500 6210 2510
rect 6110 2460 6210 2500
rect 6110 2450 6120 2460
rect 6040 2440 6120 2450
rect 6200 2450 6210 2460
rect 6270 2500 6280 2510
rect 6360 2510 6440 2520
rect 6360 2500 6370 2510
rect 6270 2460 6370 2500
rect 6270 2450 6280 2460
rect 6200 2440 6280 2450
rect 6360 2450 6370 2460
rect 6430 2500 6440 2510
rect 6520 2510 6600 2520
rect 6520 2500 6530 2510
rect 6430 2460 6530 2500
rect 6430 2450 6440 2460
rect 6360 2440 6440 2450
rect 6520 2450 6530 2460
rect 6590 2500 6600 2510
rect 6680 2510 6760 2520
rect 6680 2500 6690 2510
rect 6590 2460 6690 2500
rect 6590 2450 6600 2460
rect 6520 2440 6600 2450
rect 6680 2450 6690 2460
rect 6750 2500 6760 2510
rect 6840 2510 6920 2520
rect 6840 2500 6850 2510
rect 6750 2460 6850 2500
rect 6750 2450 6760 2460
rect 6680 2440 6760 2450
rect 6840 2450 6850 2460
rect 6910 2500 6920 2510
rect 7000 2510 7080 2520
rect 7000 2500 7010 2510
rect 6910 2460 7010 2500
rect 6910 2450 6920 2460
rect 6840 2440 6920 2450
rect 7000 2450 7010 2460
rect 7070 2500 7080 2510
rect 7160 2510 7240 2520
rect 7160 2500 7170 2510
rect 7070 2460 7170 2500
rect 7070 2450 7080 2460
rect 7000 2440 7080 2450
rect 7160 2450 7170 2460
rect 7230 2500 7240 2510
rect 7320 2510 7400 2520
rect 7320 2500 7330 2510
rect 7230 2460 7330 2500
rect 7230 2450 7240 2460
rect 7160 2440 7240 2450
rect 7320 2450 7330 2460
rect 7390 2500 7400 2510
rect 7480 2510 7560 2520
rect 7480 2500 7490 2510
rect 7390 2460 7490 2500
rect 7390 2450 7400 2460
rect 7320 2440 7400 2450
rect 7480 2450 7490 2460
rect 7550 2500 7560 2510
rect 7640 2510 7720 2520
rect 7640 2500 7650 2510
rect 7550 2460 7650 2500
rect 7550 2450 7560 2460
rect 7480 2440 7560 2450
rect 7640 2450 7650 2460
rect 7710 2500 7720 2510
rect 7800 2510 7880 2520
rect 7800 2500 7810 2510
rect 7710 2460 7810 2500
rect 7710 2450 7720 2460
rect 7640 2440 7720 2450
rect 7800 2450 7810 2460
rect 7870 2500 7880 2510
rect 7960 2510 8040 2520
rect 7960 2500 7970 2510
rect 7870 2460 7970 2500
rect 7870 2450 7880 2460
rect 7800 2440 7880 2450
rect 7960 2450 7970 2460
rect 8030 2450 8040 2510
rect 7960 2440 8040 2450
rect 8120 2510 8200 2520
rect 8120 2450 8130 2510
rect 8190 2500 8200 2510
rect 8280 2510 8360 2520
rect 8280 2500 8290 2510
rect 8190 2460 8290 2500
rect 8190 2450 8200 2460
rect 8120 2440 8200 2450
rect 8280 2450 8290 2460
rect 8350 2500 8360 2510
rect 8440 2510 8520 2520
rect 8440 2500 8450 2510
rect 8350 2460 8450 2500
rect 8350 2450 8360 2460
rect 8280 2440 8360 2450
rect 8440 2450 8450 2460
rect 8510 2500 8520 2510
rect 8600 2510 8680 2520
rect 8600 2500 8610 2510
rect 8510 2460 8610 2500
rect 8510 2450 8520 2460
rect 8440 2440 8520 2450
rect 8600 2450 8610 2460
rect 8670 2500 8680 2510
rect 8760 2510 8840 2520
rect 8760 2500 8770 2510
rect 8670 2460 8770 2500
rect 8670 2450 8680 2460
rect 8600 2440 8680 2450
rect 8760 2450 8770 2460
rect 8830 2500 8840 2510
rect 8920 2510 9000 2520
rect 8920 2500 8930 2510
rect 8830 2460 8930 2500
rect 8830 2450 8840 2460
rect 8760 2440 8840 2450
rect 8920 2450 8930 2460
rect 8990 2500 9000 2510
rect 9080 2510 9160 2520
rect 9080 2500 9090 2510
rect 8990 2460 9090 2500
rect 8990 2450 9000 2460
rect 8920 2440 9000 2450
rect 9080 2450 9090 2460
rect 9150 2500 9160 2510
rect 9240 2510 9320 2520
rect 9240 2500 9250 2510
rect 9150 2460 9250 2500
rect 9150 2450 9160 2460
rect 9080 2440 9160 2450
rect 9240 2450 9250 2460
rect 9310 2500 9320 2510
rect 9400 2510 9480 2520
rect 9400 2500 9410 2510
rect 9310 2460 9410 2500
rect 9310 2450 9320 2460
rect 9240 2440 9320 2450
rect 9400 2450 9410 2460
rect 9470 2500 9480 2510
rect 9560 2510 9640 2520
rect 9560 2500 9570 2510
rect 9470 2460 9570 2500
rect 9470 2450 9480 2460
rect 9400 2440 9480 2450
rect 9560 2450 9570 2460
rect 9630 2500 9640 2510
rect 9720 2510 9800 2520
rect 9720 2500 9730 2510
rect 9630 2460 9730 2500
rect 9630 2450 9640 2460
rect 9560 2440 9640 2450
rect 9720 2450 9730 2460
rect 9790 2500 9800 2510
rect 9880 2510 9960 2520
rect 9880 2500 9890 2510
rect 9790 2460 9890 2500
rect 9790 2450 9800 2460
rect 9720 2440 9800 2450
rect 9880 2450 9890 2460
rect 9950 2500 9960 2510
rect 10040 2510 10120 2520
rect 10040 2500 10050 2510
rect 9950 2460 10050 2500
rect 9950 2450 9960 2460
rect 9880 2440 9960 2450
rect 10040 2450 10050 2460
rect 10110 2450 10120 2510
rect 10040 2440 10120 2450
rect 4550 2340 4630 2350
rect 4550 2280 4560 2340
rect 4620 2330 4630 2340
rect 5960 2340 6040 2350
rect 5960 2330 5970 2340
rect 4620 2290 5970 2330
rect 4620 2280 4630 2290
rect 4550 2270 4630 2280
rect 5960 2280 5970 2290
rect 6030 2280 6040 2340
rect 5960 2270 6040 2280
rect 10270 2340 10350 2350
rect 10270 2280 10280 2340
rect 10340 2330 10350 2340
rect 11330 2340 11410 2350
rect 11330 2330 11340 2340
rect 10340 2290 11340 2330
rect 10340 2280 10350 2290
rect 10270 2270 10350 2280
rect 11330 2280 11340 2290
rect 11400 2280 11410 2340
rect 11330 2270 11410 2280
rect 6330 2100 6410 2110
rect 6330 2040 6340 2100
rect 6400 2090 6410 2100
rect 8120 2100 8200 2110
rect 8120 2090 8130 2100
rect 6400 2050 8130 2090
rect 6400 2040 6410 2050
rect 6330 2030 6410 2040
rect 8120 2040 8130 2050
rect 8190 2090 8200 2100
rect 9910 2100 9990 2110
rect 9910 2090 9920 2100
rect 8190 2050 9920 2090
rect 8190 2040 8200 2050
rect 8120 2030 8200 2040
rect 9910 2040 9920 2050
rect 9980 2040 9990 2100
rect 9910 2030 9990 2040
rect 5790 1960 5870 1970
rect 5790 1900 5800 1960
rect 5860 1950 5870 1960
rect 6150 1960 6230 1970
rect 6150 1950 6160 1960
rect 5860 1910 6160 1950
rect 5860 1900 5870 1910
rect 5790 1890 5870 1900
rect 6150 1900 6160 1910
rect 6220 1950 6230 1960
rect 6510 1960 6590 1970
rect 6510 1950 6520 1960
rect 6220 1910 6520 1950
rect 6220 1900 6230 1910
rect 6150 1890 6230 1900
rect 6510 1900 6520 1910
rect 6580 1950 6590 1960
rect 7580 1960 7660 1970
rect 7580 1950 7590 1960
rect 6580 1910 7590 1950
rect 6580 1900 6590 1910
rect 6510 1890 6590 1900
rect 7580 1900 7590 1910
rect 7650 1950 7660 1960
rect 7940 1960 8020 1970
rect 7940 1950 7950 1960
rect 7650 1910 7950 1950
rect 7650 1900 7660 1910
rect 7580 1890 7660 1900
rect 7940 1900 7950 1910
rect 8010 1950 8020 1960
rect 8300 1960 8380 1970
rect 8300 1950 8310 1960
rect 8010 1910 8310 1950
rect 8010 1900 8020 1910
rect 7940 1890 8020 1900
rect 8300 1900 8310 1910
rect 8370 1950 8380 1960
rect 8660 1960 8740 1970
rect 8660 1950 8670 1960
rect 8370 1910 8670 1950
rect 8370 1900 8380 1910
rect 8300 1890 8380 1900
rect 8660 1900 8670 1910
rect 8730 1950 8740 1960
rect 9730 1960 9810 1970
rect 9730 1950 9740 1960
rect 8730 1910 9740 1950
rect 8730 1900 8740 1910
rect 8660 1890 8740 1900
rect 9730 1900 9740 1910
rect 9800 1950 9810 1960
rect 10090 1960 10170 1970
rect 10090 1950 10100 1960
rect 9800 1910 10100 1950
rect 9800 1900 9810 1910
rect 9730 1890 9810 1900
rect 10090 1900 10100 1910
rect 10160 1950 10170 1960
rect 10450 1960 10530 1970
rect 10450 1950 10460 1960
rect 10160 1910 10460 1950
rect 10160 1900 10170 1910
rect 10090 1890 10170 1900
rect 10450 1900 10460 1910
rect 10520 1950 10530 1960
rect 11330 1960 11410 1970
rect 11330 1950 11340 1960
rect 10520 1910 11340 1950
rect 10520 1900 10530 1910
rect 10450 1890 10530 1900
rect 11330 1900 11340 1910
rect 11400 1900 11410 1960
rect 11330 1890 11410 1900
rect 6990 1790 7070 1800
rect 6990 1730 7000 1790
rect 7060 1780 7070 1790
rect 7100 1790 7180 1800
rect 7100 1780 7110 1790
rect 7060 1740 7110 1780
rect 7060 1730 7070 1740
rect 6990 1720 7070 1730
rect 7100 1730 7110 1740
rect 7170 1730 7180 1790
rect 7100 1720 7180 1730
rect 9140 1790 9220 1800
rect 9140 1730 9150 1790
rect 9210 1780 9220 1790
rect 9250 1790 9330 1800
rect 9250 1780 9260 1790
rect 9210 1740 9260 1780
rect 9210 1730 9220 1740
rect 9140 1720 9220 1730
rect 9250 1730 9260 1740
rect 9320 1730 9330 1790
rect 9250 1720 9330 1730
rect 10930 1790 11010 1800
rect 10930 1730 10940 1790
rect 11000 1780 11010 1790
rect 11330 1790 11410 1800
rect 11330 1780 11340 1790
rect 11000 1740 11340 1780
rect 11000 1730 11010 1740
rect 10930 1720 11010 1730
rect 11330 1730 11340 1740
rect 11400 1730 11410 1790
rect 11330 1720 11410 1730
rect 5610 1620 5690 1630
rect 5610 1560 5620 1620
rect 5680 1610 5690 1620
rect 6330 1620 6410 1630
rect 6330 1610 6340 1620
rect 5680 1570 6340 1610
rect 5680 1560 5690 1570
rect 5610 1550 5690 1560
rect 6330 1560 6340 1570
rect 6400 1560 6410 1620
rect 6330 1550 6410 1560
rect 8120 1620 8200 1630
rect 8120 1560 8130 1620
rect 8190 1610 8200 1620
rect 8480 1620 8560 1630
rect 8480 1610 8490 1620
rect 8190 1570 8490 1610
rect 8190 1560 8200 1570
rect 8120 1550 8200 1560
rect 8480 1560 8490 1570
rect 8550 1610 8560 1620
rect 8840 1620 8920 1630
rect 8840 1610 8850 1620
rect 8550 1570 8850 1610
rect 8550 1560 8560 1570
rect 8480 1550 8560 1560
rect 8840 1560 8850 1570
rect 8910 1560 8920 1620
rect 8840 1550 8920 1560
rect 9910 1620 9990 1630
rect 9910 1560 9920 1620
rect 9980 1610 9990 1620
rect 10630 1620 10710 1630
rect 10630 1610 10640 1620
rect 9980 1570 10640 1610
rect 9980 1560 9990 1570
rect 9910 1550 9990 1560
rect 10630 1560 10640 1570
rect 10700 1560 10710 1620
rect 10630 1550 10710 1560
rect 5970 1510 6050 1520
rect 5970 1450 5980 1510
rect 6040 1500 6050 1510
rect 6690 1510 6770 1520
rect 6690 1500 6700 1510
rect 6040 1460 6700 1500
rect 6040 1450 6050 1460
rect 5970 1440 6050 1450
rect 6690 1450 6700 1460
rect 6760 1500 6770 1510
rect 8120 1510 8200 1520
rect 8120 1500 8130 1510
rect 6760 1460 8130 1500
rect 6760 1450 6770 1460
rect 6690 1440 6770 1450
rect 8120 1450 8130 1460
rect 8190 1500 8200 1510
rect 9550 1510 9630 1520
rect 9550 1500 9560 1510
rect 8190 1460 9560 1500
rect 8190 1450 8200 1460
rect 8120 1440 8200 1450
rect 9550 1450 9560 1460
rect 9620 1500 9630 1510
rect 10270 1510 10350 1520
rect 10270 1500 10280 1510
rect 9620 1460 10280 1500
rect 9620 1450 9630 1460
rect 9550 1440 9630 1450
rect 10270 1450 10280 1460
rect 10340 1450 10350 1510
rect 10270 1440 10350 1450
rect 5110 1420 5190 1430
rect 5110 1360 5120 1420
rect 5180 1410 5190 1420
rect 7490 1420 7570 1430
rect 7490 1410 7500 1420
rect 5180 1370 7500 1410
rect 5180 1360 5190 1370
rect 5110 1350 5190 1360
rect 7490 1360 7500 1370
rect 7560 1360 7570 1420
rect 7490 1350 7570 1360
rect -390 1150 -310 1160
rect -390 1090 -380 1150
rect -320 1090 -310 1150
rect -390 1080 -310 1090
<< via2 >>
rect -380 10620 -320 10680
rect 11510 10620 11570 10680
rect -210 7690 -150 7750
rect 8890 7630 8950 7690
rect 11510 7630 11570 7690
rect 1890 7530 1950 7590
rect 3290 7530 3350 7590
rect 10290 7530 10350 7590
rect 5390 7420 5450 7480
rect 6790 7420 6850 7480
rect -210 6990 -150 7050
rect 11510 7000 11570 7060
rect -210 6460 -150 6520
rect -210 6330 -150 6390
rect 11510 6070 11570 6130
rect 11510 4810 11570 4870
rect -210 3380 -150 3440
rect 11510 3380 11570 3440
rect 11340 2750 11400 2810
rect 11340 2280 11400 2340
rect 11340 1900 11400 1960
rect 11340 1730 11400 1790
rect -380 1090 -320 1150
<< metal3 >>
rect -400 10690 -300 10700
rect -400 10610 -390 10690
rect -310 10610 -300 10690
rect -400 10600 -300 10610
rect 11490 10690 11590 10700
rect 11490 10610 11500 10690
rect 11580 10610 11590 10690
rect 11490 10600 11590 10610
rect -390 1170 -310 10600
rect -230 10520 -130 10530
rect -230 10440 -220 10520
rect -140 10440 -130 10520
rect -230 10430 -130 10440
rect 11320 10520 11420 10530
rect 11320 10440 11330 10520
rect 11410 10440 11420 10520
rect 11320 10430 11420 10440
rect -220 7750 -140 10430
rect 290 10240 750 10410
rect 990 10240 1450 10410
rect 1690 10240 2150 10410
rect 2390 10240 2850 10410
rect 3090 10240 3550 10410
rect 290 10140 3550 10240
rect 290 9950 750 10140
rect 990 9950 1450 10140
rect 1690 9950 2150 10140
rect 2390 9950 2850 10140
rect 3090 9950 3550 10140
rect 3790 10240 4250 10410
rect 4490 10240 4950 10410
rect 5190 10240 5650 10410
rect 5890 10240 6350 10410
rect 6590 10240 7050 10410
rect 3790 10140 7050 10240
rect 3790 9950 4250 10140
rect 4490 9950 4950 10140
rect 5190 9950 5650 10140
rect 5890 9950 6350 10140
rect 6590 9950 7050 10140
rect 7290 10240 7750 10410
rect 7990 10240 8450 10410
rect 8690 10240 9150 10410
rect 9390 10240 9850 10410
rect 10090 10240 10550 10410
rect 7290 10140 10550 10240
rect 7290 9950 7750 10140
rect 7990 9950 8450 10140
rect 8690 9950 9150 10140
rect 9390 9950 9850 10140
rect 10090 9950 10550 10140
rect 1870 9710 1970 9950
rect 5370 9710 5470 9950
rect 8870 9710 8970 9950
rect 290 9540 750 9710
rect 990 9540 1450 9710
rect 1690 9540 2150 9710
rect 2390 9540 2850 9710
rect 3090 9540 3550 9710
rect 290 9440 3550 9540
rect 290 9250 750 9440
rect 990 9250 1450 9440
rect 1690 9250 2150 9440
rect 2390 9250 2850 9440
rect 3090 9250 3550 9440
rect 3790 9540 4250 9710
rect 4490 9540 4950 9710
rect 5190 9540 5650 9710
rect 5890 9540 6350 9710
rect 6590 9540 7050 9710
rect 3790 9440 7050 9540
rect 3790 9250 4250 9440
rect 4490 9250 4950 9440
rect 5190 9250 5650 9440
rect 5890 9250 6350 9440
rect 6590 9250 7050 9440
rect 7290 9540 7750 9710
rect 7990 9540 8450 9710
rect 8690 9540 9150 9710
rect 9390 9540 9850 9710
rect 10090 9540 10550 9710
rect 7290 9440 10550 9540
rect 7290 9250 7750 9440
rect 7990 9250 8450 9440
rect 8690 9250 9150 9440
rect 9390 9250 9850 9440
rect 10090 9250 10550 9440
rect 1870 9010 1970 9250
rect 5370 9010 5470 9250
rect 8870 9010 8970 9250
rect 290 8840 750 9010
rect 990 8840 1450 9010
rect 1690 8840 2150 9010
rect 2390 8840 2850 9010
rect 3090 8840 3550 9010
rect 290 8740 3550 8840
rect 290 8550 750 8740
rect 990 8550 1450 8740
rect 1690 8550 2150 8740
rect 2390 8550 2850 8740
rect 3090 8550 3550 8740
rect 3790 8840 4250 9010
rect 4490 8840 4950 9010
rect 5190 8840 5650 9010
rect 5890 8840 6350 9010
rect 6590 8840 7050 9010
rect 3790 8740 7050 8840
rect 3790 8550 4250 8740
rect 4490 8550 4950 8740
rect 5190 8550 5650 8740
rect 5890 8550 6350 8740
rect 6590 8550 7050 8740
rect 7290 8840 7750 9010
rect 7990 8840 8450 9010
rect 8690 8840 9150 9010
rect 9390 8840 9850 9010
rect 10090 8840 10550 9010
rect 7290 8740 10550 8840
rect 7290 8550 7750 8740
rect 7990 8550 8450 8740
rect 8690 8550 9150 8740
rect 9390 8550 9850 8740
rect 10090 8550 10550 8740
rect 1870 8310 1970 8550
rect 5370 8310 5470 8550
rect 8870 8310 8970 8550
rect 290 8140 750 8310
rect 990 8140 1450 8310
rect 1690 8140 2150 8310
rect 2390 8140 2850 8310
rect 3090 8140 3550 8310
rect 290 8040 3550 8140
rect 290 7850 750 8040
rect 990 7850 1450 8040
rect 1690 7850 2150 8040
rect 2390 7850 2850 8040
rect 3090 7850 3550 8040
rect 3790 8140 4250 8310
rect 4490 8140 4950 8310
rect 5190 8140 5650 8310
rect 5890 8140 6350 8310
rect 6590 8140 7050 8310
rect 3790 8040 7050 8140
rect 3790 7850 4250 8040
rect 4490 7850 4950 8040
rect 5190 7850 5650 8040
rect 5890 7850 6350 8040
rect 6590 7850 7050 8040
rect 7290 8140 7750 8310
rect 7990 8140 8450 8310
rect 8690 8140 9150 8310
rect 9390 8140 9850 8310
rect 10090 8140 10550 8310
rect 7290 8040 10550 8140
rect 7290 7850 7750 8040
rect 7990 7850 8450 8040
rect 8690 7850 9150 8040
rect 9390 7850 9850 8040
rect 10090 7850 10550 8040
rect -220 7690 -210 7750
rect -150 7690 -140 7750
rect -220 7050 -140 7690
rect 1880 7590 1960 7850
rect 1880 7530 1890 7590
rect 1950 7530 1960 7590
rect 1880 7520 1960 7530
rect 3270 7600 3370 7610
rect 3270 7520 3280 7600
rect 3360 7520 3370 7600
rect 3270 7510 3370 7520
rect 5380 7480 5460 7850
rect 8880 7690 8960 7850
rect 8880 7630 8890 7690
rect 8950 7630 8960 7690
rect 8880 7620 8960 7630
rect 10270 7600 10370 7610
rect 10270 7520 10280 7600
rect 10360 7520 10370 7600
rect 10270 7510 10370 7520
rect 5380 7420 5390 7480
rect 5450 7420 5460 7480
rect 5380 7410 5460 7420
rect 6770 7490 6870 7500
rect 6770 7410 6780 7490
rect 6860 7410 6870 7490
rect 6770 7400 6870 7410
rect -220 6990 -210 7050
rect -150 6990 -140 7050
rect -220 6520 -140 6990
rect -220 6460 -210 6520
rect -150 6460 -140 6520
rect -220 6390 -140 6460
rect -220 6330 -210 6390
rect -150 6330 -140 6390
rect -220 3440 -140 6330
rect -220 3380 -210 3440
rect -150 3380 -140 3440
rect -220 1330 -140 3380
rect 11330 2810 11410 10430
rect 11330 2750 11340 2810
rect 11400 2750 11410 2810
rect 11330 2340 11410 2750
rect 11330 2280 11340 2340
rect 11400 2280 11410 2340
rect 11330 1960 11410 2280
rect 11330 1900 11340 1960
rect 11400 1900 11410 1960
rect 11330 1790 11410 1900
rect 11330 1730 11340 1790
rect 11400 1730 11410 1790
rect 11330 1330 11410 1730
rect 11500 7690 11580 10600
rect 11500 7630 11510 7690
rect 11570 7630 11580 7690
rect 11500 7060 11580 7630
rect 11500 7000 11510 7060
rect 11570 7000 11580 7060
rect 11500 6130 11580 7000
rect 11500 6070 11510 6130
rect 11570 6070 11580 6130
rect 11500 4870 11580 6070
rect 11500 4810 11510 4870
rect 11570 4810 11580 4870
rect 11500 3440 11580 4810
rect 11500 3380 11510 3440
rect 11570 3380 11580 3440
rect -230 1320 -130 1330
rect -230 1240 -220 1320
rect -140 1240 -130 1320
rect -230 1230 -130 1240
rect 11320 1320 11420 1330
rect 11320 1240 11330 1320
rect 11410 1240 11420 1320
rect 11320 1230 11420 1240
rect 11500 1170 11580 3380
rect -400 1160 -300 1170
rect -400 1080 -390 1160
rect -310 1080 -300 1160
rect -400 1070 -300 1080
rect 11490 1160 11590 1170
rect 11490 1080 11500 1160
rect 11580 1080 11590 1160
rect 11490 1070 11590 1080
<< via3 >>
rect -390 10680 -310 10690
rect -390 10620 -380 10680
rect -380 10620 -320 10680
rect -320 10620 -310 10680
rect -390 10610 -310 10620
rect 11500 10680 11580 10690
rect 11500 10620 11510 10680
rect 11510 10620 11570 10680
rect 11570 10620 11580 10680
rect 11500 10610 11580 10620
rect -220 10440 -140 10520
rect 11330 10440 11410 10520
rect 3280 7590 3360 7600
rect 3280 7530 3290 7590
rect 3290 7530 3350 7590
rect 3350 7530 3360 7590
rect 3280 7520 3360 7530
rect 10280 7590 10360 7600
rect 10280 7530 10290 7590
rect 10290 7530 10350 7590
rect 10350 7530 10360 7590
rect 10280 7520 10360 7530
rect 6780 7480 6860 7490
rect 6780 7420 6790 7480
rect 6790 7420 6850 7480
rect 6850 7420 6860 7480
rect 6780 7410 6860 7420
rect -220 1240 -140 1320
rect 11330 1240 11410 1320
rect -390 1150 -310 1160
rect -390 1090 -380 1150
rect -380 1090 -320 1150
rect -320 1090 -310 1150
rect -390 1080 -310 1090
rect 11500 1080 11580 1160
<< mimcap >>
rect 320 10230 720 10380
rect 320 10150 480 10230
rect 560 10150 720 10230
rect 320 9980 720 10150
rect 1020 10230 1420 10380
rect 1020 10150 1180 10230
rect 1260 10150 1420 10230
rect 1020 9980 1420 10150
rect 1720 10230 2120 10380
rect 1720 10150 1880 10230
rect 1960 10150 2120 10230
rect 1720 9980 2120 10150
rect 2420 10230 2820 10380
rect 2420 10150 2580 10230
rect 2660 10150 2820 10230
rect 2420 9980 2820 10150
rect 3120 10230 3520 10380
rect 3120 10150 3280 10230
rect 3360 10150 3520 10230
rect 3120 9980 3520 10150
rect 3820 10230 4220 10380
rect 3820 10150 3980 10230
rect 4060 10150 4220 10230
rect 3820 9980 4220 10150
rect 4520 10230 4920 10380
rect 4520 10150 4680 10230
rect 4760 10150 4920 10230
rect 4520 9980 4920 10150
rect 5220 10230 5620 10380
rect 5220 10150 5380 10230
rect 5460 10150 5620 10230
rect 5220 9980 5620 10150
rect 5920 10230 6320 10380
rect 5920 10150 6080 10230
rect 6160 10150 6320 10230
rect 5920 9980 6320 10150
rect 6620 10230 7020 10380
rect 6620 10150 6780 10230
rect 6860 10150 7020 10230
rect 6620 9980 7020 10150
rect 7320 10230 7720 10380
rect 7320 10150 7480 10230
rect 7560 10150 7720 10230
rect 7320 9980 7720 10150
rect 8020 10230 8420 10380
rect 8020 10150 8180 10230
rect 8260 10150 8420 10230
rect 8020 9980 8420 10150
rect 8720 10230 9120 10380
rect 8720 10150 8880 10230
rect 8960 10150 9120 10230
rect 8720 9980 9120 10150
rect 9420 10230 9820 10380
rect 9420 10150 9580 10230
rect 9660 10150 9820 10230
rect 9420 9980 9820 10150
rect 10120 10230 10520 10380
rect 10120 10150 10280 10230
rect 10360 10150 10520 10230
rect 10120 9980 10520 10150
rect 320 9530 720 9680
rect 320 9450 480 9530
rect 560 9450 720 9530
rect 320 9280 720 9450
rect 1020 9530 1420 9680
rect 1020 9450 1180 9530
rect 1260 9450 1420 9530
rect 1020 9280 1420 9450
rect 1720 9530 2120 9680
rect 1720 9450 1880 9530
rect 1960 9450 2120 9530
rect 1720 9280 2120 9450
rect 2420 9530 2820 9680
rect 2420 9450 2580 9530
rect 2660 9450 2820 9530
rect 2420 9280 2820 9450
rect 3120 9530 3520 9680
rect 3120 9450 3280 9530
rect 3360 9450 3520 9530
rect 3120 9280 3520 9450
rect 3820 9530 4220 9680
rect 3820 9450 3980 9530
rect 4060 9450 4220 9530
rect 3820 9280 4220 9450
rect 4520 9530 4920 9680
rect 4520 9450 4680 9530
rect 4760 9450 4920 9530
rect 4520 9280 4920 9450
rect 5220 9530 5620 9680
rect 5220 9450 5380 9530
rect 5460 9450 5620 9530
rect 5220 9280 5620 9450
rect 5920 9530 6320 9680
rect 5920 9450 6080 9530
rect 6160 9450 6320 9530
rect 5920 9280 6320 9450
rect 6620 9530 7020 9680
rect 6620 9450 6780 9530
rect 6860 9450 7020 9530
rect 6620 9280 7020 9450
rect 7320 9530 7720 9680
rect 7320 9450 7480 9530
rect 7560 9450 7720 9530
rect 7320 9280 7720 9450
rect 8020 9530 8420 9680
rect 8020 9450 8180 9530
rect 8260 9450 8420 9530
rect 8020 9280 8420 9450
rect 8720 9530 9120 9680
rect 8720 9450 8880 9530
rect 8960 9450 9120 9530
rect 8720 9280 9120 9450
rect 9420 9530 9820 9680
rect 9420 9450 9580 9530
rect 9660 9450 9820 9530
rect 9420 9280 9820 9450
rect 10120 9530 10520 9680
rect 10120 9450 10280 9530
rect 10360 9450 10520 9530
rect 10120 9280 10520 9450
rect 320 8830 720 8980
rect 320 8750 480 8830
rect 560 8750 720 8830
rect 320 8580 720 8750
rect 1020 8830 1420 8980
rect 1020 8750 1180 8830
rect 1260 8750 1420 8830
rect 1020 8580 1420 8750
rect 1720 8830 2120 8980
rect 1720 8750 1880 8830
rect 1960 8750 2120 8830
rect 1720 8580 2120 8750
rect 2420 8830 2820 8980
rect 2420 8750 2580 8830
rect 2660 8750 2820 8830
rect 2420 8580 2820 8750
rect 3120 8830 3520 8980
rect 3120 8750 3280 8830
rect 3360 8750 3520 8830
rect 3120 8580 3520 8750
rect 3820 8830 4220 8980
rect 3820 8750 3980 8830
rect 4060 8750 4220 8830
rect 3820 8580 4220 8750
rect 4520 8830 4920 8980
rect 4520 8750 4680 8830
rect 4760 8750 4920 8830
rect 4520 8580 4920 8750
rect 5220 8830 5620 8980
rect 5220 8750 5380 8830
rect 5460 8750 5620 8830
rect 5220 8580 5620 8750
rect 5920 8830 6320 8980
rect 5920 8750 6080 8830
rect 6160 8750 6320 8830
rect 5920 8580 6320 8750
rect 6620 8830 7020 8980
rect 6620 8750 6780 8830
rect 6860 8750 7020 8830
rect 6620 8580 7020 8750
rect 7320 8830 7720 8980
rect 7320 8750 7480 8830
rect 7560 8750 7720 8830
rect 7320 8580 7720 8750
rect 8020 8830 8420 8980
rect 8020 8750 8180 8830
rect 8260 8750 8420 8830
rect 8020 8580 8420 8750
rect 8720 8830 9120 8980
rect 8720 8750 8880 8830
rect 8960 8750 9120 8830
rect 8720 8580 9120 8750
rect 9420 8830 9820 8980
rect 9420 8750 9580 8830
rect 9660 8750 9820 8830
rect 9420 8580 9820 8750
rect 10120 8830 10520 8980
rect 10120 8750 10280 8830
rect 10360 8750 10520 8830
rect 10120 8580 10520 8750
rect 320 8130 720 8280
rect 320 8050 480 8130
rect 560 8050 720 8130
rect 320 7880 720 8050
rect 1020 8130 1420 8280
rect 1020 8050 1180 8130
rect 1260 8050 1420 8130
rect 1020 7880 1420 8050
rect 1720 8130 2120 8280
rect 1720 8050 1880 8130
rect 1960 8050 2120 8130
rect 1720 7880 2120 8050
rect 2420 8130 2820 8280
rect 2420 8050 2580 8130
rect 2660 8050 2820 8130
rect 2420 7880 2820 8050
rect 3120 8130 3520 8280
rect 3120 8050 3280 8130
rect 3360 8050 3520 8130
rect 3120 7880 3520 8050
rect 3820 8130 4220 8280
rect 3820 8050 3980 8130
rect 4060 8050 4220 8130
rect 3820 7880 4220 8050
rect 4520 8130 4920 8280
rect 4520 8050 4680 8130
rect 4760 8050 4920 8130
rect 4520 7880 4920 8050
rect 5220 8130 5620 8280
rect 5220 8050 5380 8130
rect 5460 8050 5620 8130
rect 5220 7880 5620 8050
rect 5920 8130 6320 8280
rect 5920 8050 6080 8130
rect 6160 8050 6320 8130
rect 5920 7880 6320 8050
rect 6620 8130 7020 8280
rect 6620 8050 6780 8130
rect 6860 8050 7020 8130
rect 6620 7880 7020 8050
rect 7320 8130 7720 8280
rect 7320 8050 7480 8130
rect 7560 8050 7720 8130
rect 7320 7880 7720 8050
rect 8020 8130 8420 8280
rect 8020 8050 8180 8130
rect 8260 8050 8420 8130
rect 8020 7880 8420 8050
rect 8720 8130 9120 8280
rect 8720 8050 8880 8130
rect 8960 8050 9120 8130
rect 8720 7880 9120 8050
rect 9420 8130 9820 8280
rect 9420 8050 9580 8130
rect 9660 8050 9820 8130
rect 9420 7880 9820 8050
rect 10120 8130 10520 8280
rect 10120 8050 10280 8130
rect 10360 8050 10520 8130
rect 10120 7880 10520 8050
<< mimcapcontact >>
rect 480 10150 560 10230
rect 1180 10150 1260 10230
rect 1880 10150 1960 10230
rect 2580 10150 2660 10230
rect 3280 10150 3360 10230
rect 3980 10150 4060 10230
rect 4680 10150 4760 10230
rect 5380 10150 5460 10230
rect 6080 10150 6160 10230
rect 6780 10150 6860 10230
rect 7480 10150 7560 10230
rect 8180 10150 8260 10230
rect 8880 10150 8960 10230
rect 9580 10150 9660 10230
rect 10280 10150 10360 10230
rect 480 9450 560 9530
rect 1180 9450 1260 9530
rect 1880 9450 1960 9530
rect 2580 9450 2660 9530
rect 3280 9450 3360 9530
rect 3980 9450 4060 9530
rect 4680 9450 4760 9530
rect 5380 9450 5460 9530
rect 6080 9450 6160 9530
rect 6780 9450 6860 9530
rect 7480 9450 7560 9530
rect 8180 9450 8260 9530
rect 8880 9450 8960 9530
rect 9580 9450 9660 9530
rect 10280 9450 10360 9530
rect 480 8750 560 8830
rect 1180 8750 1260 8830
rect 1880 8750 1960 8830
rect 2580 8750 2660 8830
rect 3280 8750 3360 8830
rect 3980 8750 4060 8830
rect 4680 8750 4760 8830
rect 5380 8750 5460 8830
rect 6080 8750 6160 8830
rect 6780 8750 6860 8830
rect 7480 8750 7560 8830
rect 8180 8750 8260 8830
rect 8880 8750 8960 8830
rect 9580 8750 9660 8830
rect 10280 8750 10360 8830
rect 480 8050 560 8130
rect 1180 8050 1260 8130
rect 1880 8050 1960 8130
rect 2580 8050 2660 8130
rect 3280 8050 3360 8130
rect 3980 8050 4060 8130
rect 4680 8050 4760 8130
rect 5380 8050 5460 8130
rect 6080 8050 6160 8130
rect 6780 8050 6860 8130
rect 7480 8050 7560 8130
rect 8180 8050 8260 8130
rect 8880 8050 8960 8130
rect 9580 8050 9660 8130
rect 10280 8050 10360 8130
<< metal4 >>
rect -400 10690 11590 10700
rect -400 10610 -390 10690
rect -310 10610 11500 10690
rect 11580 10610 11590 10690
rect -400 10600 11590 10610
rect -230 10520 11420 10530
rect -230 10440 -220 10520
rect -140 10440 11330 10520
rect 11410 10440 11420 10520
rect -230 10430 11420 10440
rect 470 10230 3370 10240
rect 470 10150 480 10230
rect 560 10150 1180 10230
rect 1260 10150 1880 10230
rect 1960 10150 2580 10230
rect 2660 10150 3280 10230
rect 3360 10150 3370 10230
rect 470 10140 3370 10150
rect 3970 10230 6870 10240
rect 3970 10150 3980 10230
rect 4060 10150 4680 10230
rect 4760 10150 5380 10230
rect 5460 10150 6080 10230
rect 6160 10150 6780 10230
rect 6860 10150 6870 10230
rect 3970 10140 6870 10150
rect 7470 10230 10370 10240
rect 7470 10150 7480 10230
rect 7560 10150 8180 10230
rect 8260 10150 8880 10230
rect 8960 10150 9580 10230
rect 9660 10150 10280 10230
rect 10360 10150 10370 10230
rect 7470 10140 10370 10150
rect 1870 9540 1970 10140
rect 5370 9540 5470 10140
rect 8870 9540 8970 10140
rect 470 9530 3370 9540
rect 470 9450 480 9530
rect 560 9450 1180 9530
rect 1260 9450 1880 9530
rect 1960 9450 2580 9530
rect 2660 9450 3280 9530
rect 3360 9450 3370 9530
rect 470 9440 3370 9450
rect 3970 9530 6870 9540
rect 3970 9450 3980 9530
rect 4060 9450 4680 9530
rect 4760 9450 5380 9530
rect 5460 9450 6080 9530
rect 6160 9450 6780 9530
rect 6860 9450 6870 9530
rect 3970 9440 6870 9450
rect 7470 9530 10370 9540
rect 7470 9450 7480 9530
rect 7560 9450 8180 9530
rect 8260 9450 8880 9530
rect 8960 9450 9580 9530
rect 9660 9450 10280 9530
rect 10360 9450 10370 9530
rect 7470 9440 10370 9450
rect 1870 8840 1970 9440
rect 5370 8840 5470 9440
rect 8870 8840 8970 9440
rect 470 8830 3370 8840
rect 470 8750 480 8830
rect 560 8750 1180 8830
rect 1260 8750 1880 8830
rect 1960 8750 2580 8830
rect 2660 8750 3280 8830
rect 3360 8750 3370 8830
rect 470 8740 3370 8750
rect 3970 8830 6870 8840
rect 3970 8750 3980 8830
rect 4060 8750 4680 8830
rect 4760 8750 5380 8830
rect 5460 8750 6080 8830
rect 6160 8750 6780 8830
rect 6860 8750 6870 8830
rect 3970 8740 6870 8750
rect 7470 8830 10370 8840
rect 7470 8750 7480 8830
rect 7560 8750 8180 8830
rect 8260 8750 8880 8830
rect 8960 8750 9580 8830
rect 9660 8750 10280 8830
rect 10360 8750 10370 8830
rect 7470 8740 10370 8750
rect 1870 8140 1970 8740
rect 5370 8140 5470 8740
rect 8870 8140 8970 8740
rect 470 8130 3370 8140
rect 470 8050 480 8130
rect 560 8050 1180 8130
rect 1260 8050 1880 8130
rect 1960 8050 2580 8130
rect 2660 8050 3280 8130
rect 3360 8050 3370 8130
rect 470 8040 3370 8050
rect 3970 8130 6870 8140
rect 3970 8050 3980 8130
rect 4060 8050 4680 8130
rect 4760 8050 5380 8130
rect 5460 8050 6080 8130
rect 6160 8050 6780 8130
rect 6860 8050 6870 8130
rect 3970 8040 6870 8050
rect 7470 8130 10370 8140
rect 7470 8050 7480 8130
rect 7560 8050 8180 8130
rect 8260 8050 8880 8130
rect 8960 8050 9580 8130
rect 9660 8050 10280 8130
rect 10360 8050 10370 8130
rect 7470 8040 10370 8050
rect 3270 7600 3370 8040
rect 3270 7520 3280 7600
rect 3360 7520 3370 7600
rect 3270 7510 3370 7520
rect 6770 7490 6870 8040
rect 10270 7600 10370 8040
rect 10270 7520 10280 7600
rect 10360 7520 10370 7600
rect 10270 7510 10370 7520
rect 6770 7410 6780 7490
rect 6860 7410 6870 7490
rect 6770 7400 6870 7410
rect -230 1320 11420 1330
rect -230 1240 -220 1320
rect -140 1240 11330 1320
rect 11410 1240 11420 1320
rect -230 1230 11420 1240
rect -400 1160 11590 1170
rect -400 1080 -390 1160
rect -310 1080 11500 1160
rect 11580 1080 11590 1160
rect -400 1070 11590 1080
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_9 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 2950 0 1 2720
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_10
timestamp 1723858470
transform 1 0 2950 0 1 1360
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_11
timestamp 1723858470
transform 1 0 2950 0 1 4080
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_12
timestamp 1723858470
transform 1 0 230 0 1 1360
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_13
timestamp 1723858470
transform 1 0 230 0 1 2720
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_14
timestamp 1723858470
transform 1 0 230 0 1 4080
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_15
timestamp 1723858470
transform 1 0 1590 0 1 1360
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_16
timestamp 1723858470
transform 1 0 1590 0 1 4080
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17
timestamp 1723858470
transform 1 0 1590 0 1 2720
box 0 0 1340 1340
<< labels >>
flabel metal2 910 7580 910 7580 1 FreeSans 800 0 0 80 cap_res1
flabel metal3 5460 7450 5460 7450 3 FreeSans 800 0 80 0 cap_res2
flabel metal1 3970 4740 3970 4740 3 FreeSans 800 0 80 0 Vbe2
flabel poly 9420 5380 9420 5380 5 FreeSans 800 0 0 -80 V_TOP
flabel metal1 10120 2480 10120 2480 3 FreeSans 800 0 400 0 START_UP_NFET1
flabel metal2 10420 3750 10420 3750 1 FreeSans 800 0 0 160 V_CUR_REF_REG
flabel metal2 10520 4340 10520 4340 5 FreeSans 800 0 0 -80 V_mir2
flabel metal1 5170 1990 5170 1990 3 FreeSans 800 0 80 0 NFET_GATE_10uA
flabel metal2 8160 7170 8160 7170 1 FreeSans 800 0 0 400 PFET_GATE_10uA
flabel metal2 12200 6200 12200 6200 3 FreeSans 800 0 400 0 TAIL_CUR_MIR_BIAS
port 9 e
flabel metal2 12200 7240 12200 7240 3 FreeSans 800 0 400 0 V_CMFB_S1
port 10 e
flabel metal2 12200 4060 12200 4060 3 FreeSans 800 0 400 0 ERR_AMP_REF
port 3 e
flabel metal3 11580 9500 11580 9500 3 FreeSans 800 0 400 0 VDDA
port 4 e
flabel metal3 11410 9050 11410 9050 3 FreeSans 800 0 400 0 GNDA
port 2 e
flabel metal2 5900 3750 5900 3750 1 FreeSans 800 0 0 160 Vin+
flabel metal2 5890 4040 5890 4040 5 FreeSans 800 0 0 -160 Vin-
flabel metal1 4610 2910 4610 2910 3 FreeSans 800 0 400 0 START_UP
flabel metal2 8620 4260 8620 4260 7 FreeSans 480 0 -240 0 1st_Vout_2
flabel metal2 8900 3570 8900 3570 7 FreeSans 800 0 -400 0 V_p_2
flabel metal2 7420 3570 7420 3570 3 FreeSans 800 0 400 0 V_p_1
flabel metal2 5800 4340 5800 4340 5 FreeSans 800 0 0 -80 V_mir1
flabel metal2 7700 4260 7700 4260 3 FreeSans 480 0 240 0 1st_Vout_1
flabel metal2 12200 5560 12200 5560 3 FreeSans 800 0 400 0 VB1_CUR_BIAS
port 1 e
flabel metal2 12200 6690 12200 6690 3 FreeSans 800 0 400 0 V_CMFB_S3
port 12 e
flabel metal1 8540 1210 8540 1210 3 FreeSans 800 0 400 0 VB3_CUR_BIAS
port 6 e
flabel metal1 7780 1210 7780 1210 7 FreeSans 800 0 -400 0 ERR_AMP_CUR_BIAS
port 7 w
flabel metal1 10670 1140 10670 1140 5 FreeSans 800 0 0 -400 V_CMFB_S4
port 11 s
flabel metal1 5650 1140 5650 1140 5 FreeSans 800 0 0 -400 V_CMFB_S2
port 8 s
flabel metal1 8160 1140 8160 1140 5 FreeSans 800 0 0 -400 VB2_CUR_BIAS
port 5 s
<< end >>
