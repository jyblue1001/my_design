* PEX produced on Sun Jul 27 05:06:34 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic_16.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic_16 VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 VOUT+.t12 two_stage_opamp_dummy_magic_23_0.Y.t25 VDDA.t308 VDDA.t307 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X1 VDDA.t469 GNDA.t398 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2 VDDA.t470 GNDA.t397 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 VDDA.t471 GNDA.t396 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4 bgr_11_0.1st_Vout_2.t11 bgr_11_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5 VDDA.t472 GNDA.t395 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 VOUT-.t19 two_stage_opamp_dummy_magic_23_0.cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 VDDA.t473 GNDA.t394 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8 two_stage_opamp_dummy_magic_23_0.VD1.t21 two_stage_opamp_dummy_magic_23_0.Vb1.t14 two_stage_opamp_dummy_magic_23_0.X.t16 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X9 two_stage_opamp_dummy_magic_23_0.X.t10 two_stage_opamp_dummy_magic_23_0.Vb2.t11 two_stage_opamp_dummy_magic_23_0.VD3.t34 two_stage_opamp_dummy_magic_23_0.VD3.t33 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X10 VOUT-.t15 VDDA.t421 VDDA.t423 VDDA.t422 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X11 GNDA.t154 bgr_11_0.NFET_GATE_10uA.t5 two_stage_opamp_dummy_magic_23_0.V_err_gate.t4 GNDA.t153 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X12 VOUT+.t19 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 GNDA.t573 GNDA.t571 VDDA.t440 GNDA.t572 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X14 VDDA.t474 GNDA.t393 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 VDDA.t475 GNDA.t392 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 bgr_11_0.1st_Vout_1.t11 bgr_11_0.cap_res1.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 VDDA.t476 GNDA.t391 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 GNDA.t570 GNDA.t567 GNDA.t569 GNDA.t568 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X19 VDDA.t477 GNDA.t390 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 two_stage_opamp_dummy_magic_23_0.VD2.t21 two_stage_opamp_dummy_magic_23_0.Vb1.t15 two_stage_opamp_dummy_magic_23_0.Y.t9 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X21 GNDA.t77 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t12 two_stage_opamp_dummy_magic_23_0.V_source.t25 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X22 VDDA.t478 GNDA.t389 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X23 bgr_11_0.V_mir2.t14 bgr_11_0.V_mir2.t13 VDDA.t84 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X24 VDDA.t145 bgr_11_0.V_TOP.t14 bgr_11_0.Vin-.t7 VDDA.t144 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X25 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t13 VDDA.t418 VDDA.t420 VDDA.t419 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X26 bgr_11_0.1st_Vout_1.t12 bgr_11_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t15 bgr_11_0.PFET_GATE_10uA.t10 VDDA.t450 VDDA.t449 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X28 two_stage_opamp_dummy_magic_23_0.VD1.t20 two_stage_opamp_dummy_magic_23_0.Vb1.t16 two_stage_opamp_dummy_magic_23_0.X.t15 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X29 VOUT-.t20 two_stage_opamp_dummy_magic_23_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 two_stage_opamp_dummy_magic_23_0.VD4.t9 two_stage_opamp_dummy_magic_23_0.Vb3.t8 VDDA.t23 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X31 VDDA.t479 GNDA.t388 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t16 two_stage_opamp_dummy_magic_23_0.X.t25 GNDA.t150 VDDA.t215 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X33 two_stage_opamp_dummy_magic_23_0.Vb2_2.t5 two_stage_opamp_dummy_magic_23_0.Vb2_2.t3 two_stage_opamp_dummy_magic_23_0.Vb2_2.t5 two_stage_opamp_dummy_magic_23_0.Vb2_2.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X34 VOUT-.t21 two_stage_opamp_dummy_magic_23_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 VDDA.t480 GNDA.t387 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 bgr_11_0.V_mir2.t15 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t7 bgr_11_0.V_p_2.t7 GNDA.t114 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X37 VDDA.t481 GNDA.t386 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 GNDA.t100 a_6470_23450.t0 GNDA.t35 sky130_fd_pr__res_xhigh_po_0p35 l=6
X39 VDDA.t482 GNDA.t385 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 VOUT+.t20 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X41 VDDA.t483 GNDA.t384 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 VOUT-.t22 two_stage_opamp_dummy_magic_23_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 VDDA.t484 GNDA.t383 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 VOUT-.t23 two_stage_opamp_dummy_magic_23_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 two_stage_opamp_dummy_magic_23_0.err_amp_out.t6 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t8 two_stage_opamp_dummy_magic_23_0.V_err_p.t16 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X46 VDDA.t305 two_stage_opamp_dummy_magic_23_0.Y.t26 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t13 GNDA.t202 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X47 VOUT+.t21 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X48 VOUT+.t22 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 VDDA.t485 GNDA.t382 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 VDDA.t486 GNDA.t381 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 VOUT+.t23 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 GNDA.t66 bgr_11_0.NFET_GATE_10uA.t6 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t3 GNDA.t65 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X53 bgr_11_0.V_TOP.t15 VDDA.t146 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X54 two_stage_opamp_dummy_magic_23_0.Vb2.t8 GNDA.t564 GNDA.t566 GNDA.t565 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X55 bgr_11_0.PFET_GATE_10uA.t8 bgr_11_0.1st_Vout_2.t12 VDDA.t71 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X56 VDDA.t212 two_stage_opamp_dummy_magic_23_0.V_err_gate.t14 two_stage_opamp_dummy_magic_23_0.V_err_p.t12 VDDA.t211 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X57 VDDA.t487 GNDA.t380 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X58 VDDA.t488 GNDA.t379 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 GNDA.t112 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t17 two_stage_opamp_dummy_magic_23_0.err_amp_out.t1 GNDA.t111 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X60 VOUT-.t24 two_stage_opamp_dummy_magic_23_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 VDDA.t217 bgr_11_0.V_TOP.t16 bgr_11_0.Vin+.t5 VDDA.t216 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X62 VDDA.t214 two_stage_opamp_dummy_magic_23_0.V_err_gate.t15 a_7460_6300.t10 VDDA.t213 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X63 GNDA.t200 two_stage_opamp_dummy_magic_23_0.Y.t27 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t11 VDDA.t306 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X64 VOUT-.t25 two_stage_opamp_dummy_magic_23_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X65 two_stage_opamp_dummy_magic_23_0.V_source.t26 VIN-.t0 two_stage_opamp_dummy_magic_23_0.VD1.t4 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X66 VDDA.t489 GNDA.t378 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 VDDA.t490 GNDA.t377 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 two_stage_opamp_dummy_magic_23_0.err_amp_out.t5 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t9 two_stage_opamp_dummy_magic_23_0.V_err_p.t13 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X69 bgr_11_0.V_TOP.t17 VDDA.t218 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X70 VOUT+.t24 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X71 VOUT-.t26 two_stage_opamp_dummy_magic_23_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 VDDA.t491 GNDA.t376 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X73 VDDA.t492 GNDA.t375 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 VDDA.t493 GNDA.t374 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 VOUT-.t27 two_stage_opamp_dummy_magic_23_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 VOUT-.t28 two_stage_opamp_dummy_magic_23_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X77 VDDA.t16 two_stage_opamp_dummy_magic_23_0.Vb3.t9 two_stage_opamp_dummy_magic_23_0.VD3.t6 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X78 two_stage_opamp_dummy_magic_23_0.V_err_p.t11 two_stage_opamp_dummy_magic_23_0.V_err_gate.t16 VDDA.t76 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X79 VDDA.t494 GNDA.t373 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X80 VOUT-.t29 two_stage_opamp_dummy_magic_23_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X81 VDDA.t156 two_stage_opamp_dummy_magic_23_0.Vb3.t10 two_stage_opamp_dummy_magic_23_0.VD4.t8 VDDA.t155 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X82 VOUT+.t11 two_stage_opamp_dummy_magic_23_0.Y.t28 VDDA.t304 VDDA.t303 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X83 bgr_11_0.V_TOP.t18 VDDA.t141 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 VOUT-.t30 two_stage_opamp_dummy_magic_23_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 two_stage_opamp_dummy_magic_23_0.VD1.t6 VIN-.t1 two_stage_opamp_dummy_magic_23_0.V_source.t31 GNDA.t113 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X86 VOUT-.t31 two_stage_opamp_dummy_magic_23_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X87 VOUT+.t25 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 VOUT-.t32 two_stage_opamp_dummy_magic_23_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 two_stage_opamp_dummy_magic_23_0.Y.t23 two_stage_opamp_dummy_magic_23_0.Vb2.t12 two_stage_opamp_dummy_magic_23_0.VD4.t37 two_stage_opamp_dummy_magic_23_0.VD4.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X90 VDDA.t417 VDDA.t415 two_stage_opamp_dummy_magic_23_0.err_amp_out.t9 VDDA.t416 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X91 VDDA.t495 GNDA.t372 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X92 VOUT+.t26 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X93 VOUT-.t33 two_stage_opamp_dummy_magic_23_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X94 bgr_11_0.V_mir2.t0 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t10 bgr_11_0.V_p_2.t6 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X95 VOUT+.t27 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X96 VDDA.t496 GNDA.t371 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 VDDA.t497 GNDA.t370 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X98 VDDA.t498 GNDA.t369 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X99 bgr_11_0.Vin+.t4 bgr_11_0.V_TOP.t19 VDDA.t143 VDDA.t142 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X100 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t14 two_stage_opamp_dummy_magic_23_0.X.t26 VDDA.t189 GNDA.t148 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X101 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t10 two_stage_opamp_dummy_magic_23_0.Y.t29 GNDA.t201 VDDA.t302 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X102 two_stage_opamp_dummy_magic_23_0.VD2.t4 VIN+.t0 two_stage_opamp_dummy_magic_23_0.V_source.t29 GNDA.t109 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X103 VDDA.t499 GNDA.t368 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X104 bgr_11_0.NFET_GATE_10uA.t4 bgr_11_0.PFET_GATE_10uA.t11 VDDA.t465 VDDA.t464 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X105 VDDA.t500 GNDA.t367 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X106 VOUT-.t34 two_stage_opamp_dummy_magic_23_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 VDDA.t121 bgr_11_0.PFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t3 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X108 VDDA.t414 VDDA.t412 two_stage_opamp_dummy_magic_23_0.V_err_gate.t11 VDDA.t413 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X109 bgr_11_0.V_TOP.t20 VDDA.t429 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X110 VOUT-.t35 two_stage_opamp_dummy_magic_23_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 VOUT+.t28 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X112 bgr_11_0.1st_Vout_2.t5 bgr_11_0.V_mir2.t17 VDDA.t220 VDDA.t219 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X113 GNDA.t64 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t13 two_stage_opamp_dummy_magic_23_0.V_source.t24 GNDA.t63 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X114 VOUT-.t36 two_stage_opamp_dummy_magic_23_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 VOUT-.t37 two_stage_opamp_dummy_magic_23_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X116 VOUT+.t29 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X117 GNDA.t563 GNDA.t561 two_stage_opamp_dummy_magic_23_0.Vb1.t5 GNDA.t562 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X118 VDDA.t501 GNDA.t366 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 two_stage_opamp_dummy_magic_23_0.VD1.t19 two_stage_opamp_dummy_magic_23_0.Vb1.t17 two_stage_opamp_dummy_magic_23_0.X.t20 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X120 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t15 two_stage_opamp_dummy_magic_23_0.X.t27 GNDA.t149 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X121 VOUT-.t38 two_stage_opamp_dummy_magic_23_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t14 two_stage_opamp_dummy_magic_23_0.X.t28 GNDA.t145 VDDA.t180 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X123 VDDA.t502 GNDA.t365 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 VDDA.t503 GNDA.t364 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 VDDA.t504 GNDA.t363 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 VDDA.t505 GNDA.t362 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X127 bgr_11_0.V_TOP.t21 VDDA.t430 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 bgr_11_0.V_mir2.t2 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t11 bgr_11_0.V_p_2.t5 GNDA.t101 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X129 VOUT+.t30 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 a_12070_24908.t1 bgr_11_0.V_CUR_REF_REG.t1 GNDA.t89 sky130_fd_pr__res_xhigh_po_0p35 l=4
X131 two_stage_opamp_dummy_magic_23_0.Vb3.t6 GNDA.t558 GNDA.t560 GNDA.t559 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X132 VDDA.t459 two_stage_opamp_dummy_magic_23_0.Vb3.t11 two_stage_opamp_dummy_magic_23_0.VD4.t7 VDDA.t458 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X133 VOUT+.t31 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 VOUT-.t39 two_stage_opamp_dummy_magic_23_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X135 VDDA.t506 GNDA.t361 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X136 VOUT+.t32 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X137 VOUT+.t33 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 two_stage_opamp_dummy_magic_23_0.Vb3.t4 bgr_11_0.NFET_GATE_10uA.t7 GNDA.t68 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X139 bgr_11_0.1st_Vout_2.t13 bgr_11_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 VDDA.t507 GNDA.t360 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X141 VDDA.t508 GNDA.t359 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X142 bgr_11_0.V_mir1.t11 bgr_11_0.V_mir1.t10 VDDA.t246 VDDA.t245 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X143 two_stage_opamp_dummy_magic_23_0.X.t19 two_stage_opamp_dummy_magic_23_0.Vb1.t18 two_stage_opamp_dummy_magic_23_0.VD1.t18 GNDA.t113 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X144 VDDA.t411 VDDA.t409 VOUT-.t14 VDDA.t410 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X145 VDDA.t509 GNDA.t358 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X146 VDDA.t510 GNDA.t357 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 VOUT+.t34 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 bgr_11_0.1st_Vout_1.t13 bgr_11_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 VOUT+.t35 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 VDDA.t78 two_stage_opamp_dummy_magic_23_0.V_err_gate.t17 a_7460_6300.t9 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X151 GNDA.t39 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t11 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t12 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X152 bgr_11_0.1st_Vout_2.t14 bgr_11_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X153 VDDA.t511 GNDA.t356 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 VOUT-.t40 two_stage_opamp_dummy_magic_23_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X155 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t4 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0 ps=0 w=3.5 l=0.2
X156 VDDA.t512 GNDA.t355 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 VOUT-.t41 two_stage_opamp_dummy_magic_23_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 VOUT+.t36 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 GNDA.t477 VDDA.t403 VDDA.t405 VDDA.t404 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X160 two_stage_opamp_dummy_magic_23_0.Y.t19 two_stage_opamp_dummy_magic_23_0.Vb1.t19 two_stage_opamp_dummy_magic_23_0.VD2.t20 GNDA.t109 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X161 two_stage_opamp_dummy_magic_23_0.V_source.t23 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t14 GNDA.t152 GNDA.t151 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X162 two_stage_opamp_dummy_magic_23_0.V_source.t22 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t15 GNDA.t168 GNDA.t167 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X163 VDDA.t152 bgr_11_0.PFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_23_0.Vb1.t1 VDDA.t151 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X164 VDDA.t88 two_stage_opamp_dummy_magic_23_0.Vb3.t12 two_stage_opamp_dummy_magic_23_0.VD4.t6 VDDA.t87 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X165 VOUT-.t42 two_stage_opamp_dummy_magic_23_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 VOUT-.t43 two_stage_opamp_dummy_magic_23_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X167 VOUT+.t37 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X168 VDDA.t513 GNDA.t354 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X169 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t13 VDDA.t406 VDDA.t408 VDDA.t407 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X170 VDDA.t514 GNDA.t353 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 VOUT+.t38 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X172 VDDA.t402 VDDA.t400 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t6 VDDA.t401 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X173 VDDA.t515 GNDA.t352 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t3 bgr_11_0.PFET_GATE_10uA.t14 VDDA.t48 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X175 VOUT+.t39 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 two_stage_opamp_dummy_magic_23_0.X.t4 two_stage_opamp_dummy_magic_23_0.VD3.t3 two_stage_opamp_dummy_magic_23_0.VD3.t5 two_stage_opamp_dummy_magic_23_0.VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X177 VDDA.t516 GNDA.t351 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X178 VOUT+.t40 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X179 VOUT+.t41 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X180 VOUT-.t44 two_stage_opamp_dummy_magic_23_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 VOUT+.t42 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 VDDA.t517 GNDA.t350 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 VDDA.t518 GNDA.t349 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X184 VDDA.t519 GNDA.t348 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 two_stage_opamp_dummy_magic_23_0.VD3.t32 two_stage_opamp_dummy_magic_23_0.Vb2.t13 two_stage_opamp_dummy_magic_23_0.X.t12 two_stage_opamp_dummy_magic_23_0.VD3.t31 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X186 VOUT+.t10 two_stage_opamp_dummy_magic_23_0.Y.t30 VDDA.t301 VDDA.t300 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X187 VOUT-.t45 two_stage_opamp_dummy_magic_23_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 bgr_11_0.START_UP_NFET1.t0 bgr_11_0.START_UP_NFET1 GNDA.t166 GNDA.t165 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X189 bgr_11_0.1st_Vout_2.t15 bgr_11_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X190 VOUT-.t46 two_stage_opamp_dummy_magic_23_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 VOUT+.t43 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 VDDA.t520 GNDA.t347 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X193 bgr_11_0.PFET_GATE_10uA.t7 bgr_11_0.1st_Vout_2.t16 VDDA.t66 VDDA.t65 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X194 VDDA.t521 GNDA.t346 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 two_stage_opamp_dummy_magic_23_0.VD2.t6 VIN+.t1 two_stage_opamp_dummy_magic_23_0.V_source.t33 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X196 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t13 two_stage_opamp_dummy_magic_23_0.X.t29 VDDA.t181 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X197 bgr_11_0.V_TOP.t22 VDDA.t427 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t9 two_stage_opamp_dummy_magic_23_0.Y.t31 GNDA.t199 VDDA.t299 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X199 two_stage_opamp_dummy_magic_23_0.VD2.t5 VIN+.t2 two_stage_opamp_dummy_magic_23_0.V_source.t30 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X200 two_stage_opamp_dummy_magic_23_0.V_p_mir.t3 VIN+.t3 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t6 GNDA.t151 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X201 VOUT+.t44 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 VOUT+.t45 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X203 VDDA.t522 GNDA.t345 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X204 VDDA.t399 VDDA.t397 two_stage_opamp_dummy_magic_23_0.VD4.t17 VDDA.t398 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X205 a_7460_6300.t16 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t12 two_stage_opamp_dummy_magic_23_0.V_err_gate.t5 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X206 VDDA.t523 GNDA.t344 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 VOUT-.t47 two_stage_opamp_dummy_magic_23_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 VDDA.t524 GNDA.t343 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 VOUT+.t46 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 GNDA.t18 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t16 two_stage_opamp_dummy_magic_23_0.V_source.t21 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X211 VDDA.t525 GNDA.t342 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 a_6350_25058.t0 bgr_11_0.Vin+.t1 GNDA.t35 sky130_fd_pr__res_xhigh_po_0p35 l=6
X213 bgr_11_0.1st_Vout_2.t7 bgr_11_0.V_CUR_REF_REG.t3 bgr_11_0.V_p_2.t10 GNDA.t574 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X214 a_8260_1600.t4 two_stage_opamp_dummy_magic_23_0.Vb1.t10 two_stage_opamp_dummy_magic_23_0.Vb1.t11 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X215 VDDA.t526 GNDA.t341 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t13 two_stage_opamp_dummy_magic_23_0.X.t30 GNDA.t180 VDDA.t260 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X217 VOUT-.t48 two_stage_opamp_dummy_magic_23_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X218 VOUT+.t47 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X219 VOUT-.t49 two_stage_opamp_dummy_magic_23_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X220 two_stage_opamp_dummy_magic_23_0.VD3.t14 VDDA.t394 VDDA.t396 VDDA.t395 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X221 VDDA.t527 GNDA.t340 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 VDDA.t528 GNDA.t339 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 VOUT-.t50 two_stage_opamp_dummy_magic_23_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X224 VDDA.t529 GNDA.t338 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X225 bgr_11_0.1st_Vout_2.t10 bgr_11_0.V_mir2.t18 VDDA.t461 VDDA.t460 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X226 bgr_11_0.V_TOP.t13 bgr_11_0.1st_Vout_1.t14 VDDA.t62 VDDA.t61 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X227 VDDA.t289 two_stage_opamp_dummy_magic_23_0.Y.t32 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t12 GNDA.t198 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X228 VOUT-.t51 two_stage_opamp_dummy_magic_23_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 bgr_11_0.V_CUR_REF_REG.t2 VDDA.t391 VDDA.t393 VDDA.t392 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X230 VDDA.t110 bgr_11_0.PFET_GATE_10uA.t15 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t2 VDDA.t109 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X231 VDDA.t530 GNDA.t337 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 VOUT-.t52 two_stage_opamp_dummy_magic_23_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X233 VOUT-.t53 two_stage_opamp_dummy_magic_23_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X234 VOUT-.t54 two_stage_opamp_dummy_magic_23_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X235 VDDA.t531 GNDA.t336 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 VDDA.t262 two_stage_opamp_dummy_magic_23_0.X.t31 VOUT-.t13 VDDA.t261 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X237 bgr_11_0.1st_Vout_1.t8 bgr_11_0.Vin+.t6 bgr_11_0.V_p_1.t4 GNDA.t575 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X238 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t10 bgr_11_0.PFET_GATE_10uA.t16 VDDA.t448 VDDA.t447 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X239 bgr_11_0.V_TOP.t23 VDDA.t428 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 VDDA.t532 GNDA.t335 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 bgr_11_0.1st_Vout_1.t5 bgr_11_0.V_mir1.t17 VDDA.t135 VDDA.t134 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X242 GNDA.t43 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t9 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t10 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X243 VOUT-.t55 two_stage_opamp_dummy_magic_23_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 VOUT+.t48 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 VOUT+.t49 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 VOUT+.t50 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 VOUT+.t51 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X248 bgr_11_0.START_UP.t5 bgr_11_0.V_TOP.t24 VDDA.t33 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X249 VDDA.t204 two_stage_opamp_dummy_magic_23_0.V_err_gate.t18 two_stage_opamp_dummy_magic_23_0.V_err_p.t10 VDDA.t203 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X250 two_stage_opamp_dummy_magic_23_0.Y.t7 two_stage_opamp_dummy_magic_23_0.Vb1.t20 two_stage_opamp_dummy_magic_23_0.VD2.t19 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X251 VDDA.t533 GNDA.t334 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X252 VDDA.t534 GNDA.t333 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 two_stage_opamp_dummy_magic_23_0.Y.t8 two_stage_opamp_dummy_magic_23_0.Vb1.t21 two_stage_opamp_dummy_magic_23_0.VD2.t18 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X254 VDDA.t535 GNDA.t332 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X255 VOUT+.t52 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 two_stage_opamp_dummy_magic_23_0.V_source.t20 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t17 GNDA.t120 GNDA.t119 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X257 two_stage_opamp_dummy_magic_23_0.VD3.t30 two_stage_opamp_dummy_magic_23_0.Vb2.t14 two_stage_opamp_dummy_magic_23_0.X.t0 two_stage_opamp_dummy_magic_23_0.VD3.t29 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X258 GNDA.t557 GNDA.t555 VOUT+.t16 GNDA.t556 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X259 GNDA.t485 GNDA.t486 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X260 bgr_11_0.Vin+.t0 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 GNDA.t16 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X261 VDDA.t536 GNDA.t331 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 VOUT-.t56 two_stage_opamp_dummy_magic_23_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 two_stage_opamp_dummy_magic_23_0.VD3.t9 two_stage_opamp_dummy_magic_23_0.Vb3.t13 VDDA.t97 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X264 VDDA.t537 GNDA.t330 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 two_stage_opamp_dummy_magic_23_0.VD4.t5 two_stage_opamp_dummy_magic_23_0.Vb3.t14 VDDA.t103 VDDA.t102 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X266 bgr_11_0.1st_Vout_2.t17 bgr_11_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X267 VDDA.t538 GNDA.t329 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X268 VOUT-.t57 two_stage_opamp_dummy_magic_23_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 VDDA.t390 VDDA.t388 bgr_11_0.PFET_GATE_10uA.t1 VDDA.t389 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X270 bgr_11_0.1st_Vout_1.t4 bgr_11_0.Vin+.t7 bgr_11_0.V_p_1.t3 GNDA.t88 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X271 VOUT-.t58 two_stage_opamp_dummy_magic_23_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X272 VDDA.t539 GNDA.t328 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X273 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t11 two_stage_opamp_dummy_magic_23_0.Y.t33 VDDA.t298 GNDA.t197 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X274 VDDA.t540 GNDA.t327 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X275 VDDA.t541 GNDA.t326 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X276 VOUT+.t53 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 VDDA.t542 GNDA.t325 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X278 bgr_11_0.V_TOP.t2 bgr_11_0.START_UP.t6 bgr_11_0.Vin-.t2 VDDA.t247 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X279 VOUT+.t54 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X280 bgr_11_0.cap_res1.t0 bgr_11_0.V_TOP.t0 GNDA.t57 sky130_fd_pr__res_high_po_0p35 l=2.05
X281 bgr_11_0.V_mir2.t12 bgr_11_0.V_mir2.t11 VDDA.t127 VDDA.t126 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X282 VOUT+.t55 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X283 VOUT+.t56 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t12 two_stage_opamp_dummy_magic_23_0.X.t32 VDDA.t241 GNDA.t161 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X285 VDDA.t543 GNDA.t324 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 VDDA.t387 VDDA.t385 bgr_11_0.V_TOP.t6 VDDA.t386 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X287 a_7460_6300.t8 two_stage_opamp_dummy_magic_23_0.V_err_gate.t19 VDDA.t206 VDDA.t205 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X288 a_7460_6300.t7 two_stage_opamp_dummy_magic_23_0.V_err_gate.t20 VDDA.t183 VDDA.t182 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X289 two_stage_opamp_dummy_magic_23_0.VD2.t10 VIN+.t4 two_stage_opamp_dummy_magic_23_0.V_source.t38 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X290 VDDA.t544 GNDA.t323 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X291 a_7460_6300.t15 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t13 two_stage_opamp_dummy_magic_23_0.V_err_gate.t2 VDDA.t69 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X292 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t8 two_stage_opamp_dummy_magic_23_0.Y.t34 GNDA.t194 VDDA.t297 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X293 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t11 two_stage_opamp_dummy_magic_23_0.X.t33 VDDA.t242 GNDA.t162 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X294 VOUT+.t57 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 VDDA.t384 VDDA.t382 GNDA.t476 VDDA.t383 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X296 VDDA.t545 GNDA.t322 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X297 VDDA.t546 GNDA.t321 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X298 VDDA.t547 GNDA.t320 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X299 GNDA.t70 bgr_11_0.NFET_GATE_10uA.t8 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t2 GNDA.t69 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X300 bgr_11_0.1st_Vout_2.t3 bgr_11_0.V_CUR_REF_REG.t4 bgr_11_0.V_p_2.t1 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X301 bgr_11_0.1st_Vout_2.t18 bgr_11_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 two_stage_opamp_dummy_magic_23_0.Vb2.t6 bgr_11_0.NFET_GATE_10uA.t9 GNDA.t129 GNDA.t128 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X303 VOUT-.t59 two_stage_opamp_dummy_magic_23_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 VDDA.t548 GNDA.t319 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X305 a_8260_1600.t3 two_stage_opamp_dummy_magic_23_0.Vb1.t12 two_stage_opamp_dummy_magic_23_0.Vb1.t13 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X306 VOUT+.t58 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X307 bgr_11_0.1st_Vout_1.t1 bgr_11_0.V_mir1.t18 VDDA.t39 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X308 VOUT-.t10 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t2 GNDA.t164 GNDA.t163 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X309 VOUT-.t60 two_stage_opamp_dummy_magic_23_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 VDDA.t549 GNDA.t318 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X311 VDDA.t550 GNDA.t317 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X312 VOUT+.t59 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 VDDA.t551 GNDA.t316 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 VDDA.t552 GNDA.t315 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 VDDA.t35 bgr_11_0.V_TOP.t25 bgr_11_0.Vin+.t3 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X316 VDDA.t441 GNDA.t552 GNDA.t554 GNDA.t553 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X317 bgr_11_0.1st_Vout_1.t15 bgr_11_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 VOUT+.t60 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 VOUT-.t61 two_stage_opamp_dummy_magic_23_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 VOUT+.t61 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X321 VDDA.t553 GNDA.t314 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X322 VDDA.t554 GNDA.t313 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 VDDA.t555 GNDA.t312 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X324 two_stage_opamp_dummy_magic_23_0.Vb3.t7 two_stage_opamp_dummy_magic_23_0.Vb2.t15 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t10 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t9 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X325 VDDA.t187 two_stage_opamp_dummy_magic_23_0.X.t34 VOUT-.t6 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X326 a_4200_4468.t0 two_stage_opamp_dummy_magic_23_0.V_tot.t2 GNDA.t136 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X327 VOUT+.t62 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 two_stage_opamp_dummy_magic_23_0.VD4.t4 two_stage_opamp_dummy_magic_23_0.Vb3.t15 VDDA.t73 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X329 GNDA.t20 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t18 two_stage_opamp_dummy_magic_23_0.err_amp_out.t0 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X330 VDDA.t556 GNDA.t311 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X331 VDDA.t185 two_stage_opamp_dummy_magic_23_0.V_err_gate.t21 a_7460_6300.t6 VDDA.t184 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X332 two_stage_opamp_dummy_magic_23_0.Y.t5 two_stage_opamp_dummy_magic_23_0.Vb1.t22 two_stage_opamp_dummy_magic_23_0.VD2.t17 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X333 bgr_11_0.1st_Vout_1.t16 bgr_11_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X334 VOUT-.t0 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t3 GNDA.t80 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X335 VOUT+.t63 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X336 VDDA.t557 GNDA.t310 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X337 bgr_11_0.V_TOP.t12 bgr_11_0.1st_Vout_1.t17 VDDA.t31 VDDA.t30 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X338 two_stage_opamp_dummy_magic_23_0.VD3.t28 two_stage_opamp_dummy_magic_23_0.Vb2.t16 two_stage_opamp_dummy_magic_23_0.X.t8 two_stage_opamp_dummy_magic_23_0.VD3.t27 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X339 two_stage_opamp_dummy_magic_23_0.V_source.t19 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t18 GNDA.t172 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X340 GNDA.t135 a_5820_23634.t0 GNDA.t73 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X341 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t6 bgr_11_0.V_TOP.t26 VDDA.t28 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X342 VDDA.t558 GNDA.t309 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X343 two_stage_opamp_dummy_magic_23_0.X.t9 two_stage_opamp_dummy_magic_23_0.Vb2.t17 two_stage_opamp_dummy_magic_23_0.VD3.t26 two_stage_opamp_dummy_magic_23_0.VD3.t25 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X344 VOUT+.t0 GNDA.t549 GNDA.t551 GNDA.t550 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X345 VDDA.t559 GNDA.t308 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X346 VOUT-.t62 two_stage_opamp_dummy_magic_23_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X347 VDDA.t560 GNDA.t307 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X348 VOUT-.t63 two_stage_opamp_dummy_magic_23_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X349 VOUT+.t9 two_stage_opamp_dummy_magic_23_0.Y.t35 VDDA.t296 VDDA.t295 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X350 VOUT+.t64 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 VOUT-.t64 two_stage_opamp_dummy_magic_23_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X352 two_stage_opamp_dummy_magic_23_0.VD4.t35 two_stage_opamp_dummy_magic_23_0.Vb2.t18 two_stage_opamp_dummy_magic_23_0.Y.t22 two_stage_opamp_dummy_magic_23_0.VD4.t34 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X353 bgr_11_0.V_TOP.t11 bgr_11_0.1st_Vout_1.t18 VDDA.t6 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X354 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t10 two_stage_opamp_dummy_magic_23_0.Y.t36 VDDA.t294 GNDA.t196 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X355 VDDA.t561 GNDA.t306 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X356 VOUT+.t65 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X357 VOUT+.t66 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X358 a_11420_25058.t1 bgr_11_0.Vin-.t0 GNDA.t2 sky130_fd_pr__res_xhigh_po_0p35 l=6
X359 bgr_11_0.V_TOP.t27 VDDA.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X360 VOUT+.t67 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X361 VDDA.t562 GNDA.t305 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X362 GNDA.t548 GNDA.t546 bgr_11_0.NFET_GATE_10uA.t3 GNDA.t547 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X363 two_stage_opamp_dummy_magic_23_0.V_err_gate.t3 bgr_11_0.NFET_GATE_10uA.t10 GNDA.t131 GNDA.t130 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X364 VDDA.t563 GNDA.t304 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X365 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t10 two_stage_opamp_dummy_magic_23_0.X.t35 VDDA.t188 GNDA.t147 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X366 bgr_11_0.1st_Vout_1.t19 bgr_11_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X367 two_stage_opamp_dummy_magic_23_0.V_err_p.t9 two_stage_opamp_dummy_magic_23_0.V_err_gate.t22 VDDA.t167 VDDA.t166 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X368 two_stage_opamp_dummy_magic_23_0.VD2.t7 VIN+.t5 two_stage_opamp_dummy_magic_23_0.V_source.t35 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X369 VDDA.t564 GNDA.t303 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X370 a_7460_6300.t0 two_stage_opamp_dummy_magic_23_0.V_tot.t4 two_stage_opamp_dummy_magic_23_0.V_err_gate.t0 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X371 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t7 two_stage_opamp_dummy_magic_23_0.Y.t37 GNDA.t195 VDDA.t293 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X372 VOUT+.t15 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t4 GNDA.t581 GNDA.t580 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X373 GNDA.t37 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t19 two_stage_opamp_dummy_magic_23_0.V_source.t18 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X374 bgr_11_0.V_TOP.t28 VDDA.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 VOUT+.t68 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X376 VOUT-.t65 two_stage_opamp_dummy_magic_23_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X377 VDDA.t68 two_stage_opamp_dummy_magic_23_0.Vb3.t16 two_stage_opamp_dummy_magic_23_0.VD3.t7 VDDA.t67 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X378 VOUT-.t66 two_stage_opamp_dummy_magic_23_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 VDDA.t60 bgr_11_0.V_TOP.t29 bgr_11_0.START_UP.t4 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X380 VDDA.t565 GNDA.t302 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X381 VDDA.t457 bgr_11_0.PFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t16 VDDA.t456 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X382 VOUT-.t67 two_stage_opamp_dummy_magic_23_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 bgr_11_0.Vin-.t6 bgr_11_0.V_TOP.t30 VDDA.t94 VDDA.t93 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X384 VDDA.t566 GNDA.t301 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X385 VOUT-.t68 two_stage_opamp_dummy_magic_23_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X386 VDDA.t567 GNDA.t300 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X387 VDDA.t568 GNDA.t299 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 bgr_11_0.V_mir1.t9 bgr_11_0.V_mir1.t8 VDDA.t113 VDDA.t112 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X389 bgr_11_0.V_mir1.t14 bgr_11_0.Vin-.t8 bgr_11_0.V_p_1.t10 GNDA.t132 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X390 VDDA.t292 two_stage_opamp_dummy_magic_23_0.Y.t38 VOUT+.t8 VDDA.t291 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X391 VOUT-.t69 two_stage_opamp_dummy_magic_23_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X392 VDDA.t569 GNDA.t298 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X393 VDDA.t570 GNDA.t297 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 bgr_11_0.V_TOP.t5 VDDA.t379 VDDA.t381 VDDA.t380 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X395 bgr_11_0.V_TOP.t31 VDDA.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X396 VOUT+.t69 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X397 VDDA.t571 GNDA.t296 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X398 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t8 VDDA.t376 VDDA.t378 VDDA.t377 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X399 VOUT+.t70 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 VDDA.t208 two_stage_opamp_dummy_magic_23_0.X.t36 VOUT-.t7 VDDA.t207 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X401 VDDA.t572 GNDA.t295 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X402 GNDA.t53 bgr_11_0.NFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_23_0.Vb2.t3 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X403 two_stage_opamp_dummy_magic_23_0.Y.t17 two_stage_opamp_dummy_magic_23_0.VD4.t13 two_stage_opamp_dummy_magic_23_0.VD4.t15 two_stage_opamp_dummy_magic_23_0.VD4.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X404 VDDA.t210 two_stage_opamp_dummy_magic_23_0.X.t37 VOUT-.t8 VDDA.t209 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X405 VDDA.t573 GNDA.t294 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 VDDA.t574 GNDA.t293 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X407 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t2 bgr_11_0.NFET_GATE_10uA.t12 GNDA.t55 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X408 bgr_11_0.V_TOP.t32 VDDA.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X409 GNDA.t589 a_11950_23700.t1 GNDA.t588 sky130_fd_pr__res_xhigh_po_0p35 l=4
X410 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t1 bgr_11_0.NFET_GATE_10uA.t13 GNDA.t97 GNDA.t96 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X411 two_stage_opamp_dummy_magic_23_0.X.t11 two_stage_opamp_dummy_magic_23_0.Vb2.t19 two_stage_opamp_dummy_magic_23_0.VD3.t24 two_stage_opamp_dummy_magic_23_0.VD3.t23 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X412 VOUT-.t70 two_stage_opamp_dummy_magic_23_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X413 VOUT+.t71 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 two_stage_opamp_dummy_magic_23_0.Y.t6 two_stage_opamp_dummy_magic_23_0.Vb1.t23 two_stage_opamp_dummy_magic_23_0.VD2.t16 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X415 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t0 a_4600_1446.t0 GNDA.t74 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X416 VDDA.t575 GNDA.t292 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 VDDA.t154 two_stage_opamp_dummy_magic_23_0.Vb3.t17 two_stage_opamp_dummy_magic_23_0.VD3.t12 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X418 a_4080_4468.t1 two_stage_opamp_dummy_magic_23_0.V_tot.t1 GNDA.t110 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X419 VDDA.t576 GNDA.t291 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X420 VDDA.t444 bgr_11_0.V_mir2.t19 bgr_11_0.1st_Vout_2.t9 VDDA.t443 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X421 VOUT-.t9 a_13130_1456.t1 GNDA.t156 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X422 bgr_11_0.1st_Vout_2.t19 bgr_11_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 VOUT-.t71 two_stage_opamp_dummy_magic_23_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X424 two_stage_opamp_dummy_magic_23_0.V_source.t17 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t20 GNDA.t601 GNDA.t482 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X425 VDDA.t577 GNDA.t290 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X426 VDDA.t578 GNDA.t289 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 VOUT+.t72 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 VOUT-.t72 two_stage_opamp_dummy_magic_23_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X429 bgr_11_0.V_mir1.t16 bgr_11_0.Vin-.t9 bgr_11_0.V_p_1.t9 GNDA.t133 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X430 GNDA.t485 GNDA.t539 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X431 GNDA.t144 two_stage_opamp_dummy_magic_23_0.X.t38 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t12 VDDA.t177 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X432 bgr_11_0.V_mir1.t7 bgr_11_0.V_mir1.t6 VDDA.t26 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X433 VOUT-.t73 two_stage_opamp_dummy_magic_23_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 VDDA.t579 GNDA.t288 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 VOUT+.t73 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 bgr_11_0.1st_Vout_1.t20 bgr_11_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 VDDA.t580 GNDA.t287 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 VOUT+.t74 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 bgr_11_0.START_UP.t1 bgr_11_0.START_UP.t0 bgr_11_0.START_UP_NFET1.t0 GNDA.t591 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X440 bgr_11_0.1st_Vout_2.t20 bgr_11_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 bgr_11_0.PFET_GATE_10uA.t0 VDDA.t373 VDDA.t375 VDDA.t374 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X442 VDDA.t581 GNDA.t286 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X443 VOUT+.t75 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X444 VDDA.t582 GNDA.t285 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 VOUT+.t14 VDDA.t370 VDDA.t372 VDDA.t371 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X446 two_stage_opamp_dummy_magic_23_0.cap_res_X.t0 two_stage_opamp_dummy_magic_23_0.X.t7 GNDA.t155 sky130_fd_pr__res_high_po_1p41 l=1.41
X447 VOUT+.t76 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X448 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t9 two_stage_opamp_dummy_magic_23_0.Y.t39 VDDA.t290 GNDA.t193 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X449 two_stage_opamp_dummy_magic_23_0.VD1.t8 VIN-.t2 two_stage_opamp_dummy_magic_23_0.V_source.t34 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X450 GNDA.t545 GNDA.t543 two_stage_opamp_dummy_magic_23_0.V_source.t36 GNDA.t544 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X451 GNDA.t542 GNDA.t540 VDDA.t40 GNDA.t541 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X452 VDDA.t583 GNDA.t284 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X453 two_stage_opamp_dummy_magic_23_0.V_err_p.t0 two_stage_opamp_dummy_magic_23_0.V_tot.t5 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t0 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X454 VDDA.t584 GNDA.t283 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X455 bgr_11_0.1st_Vout_1.t21 bgr_11_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 bgr_11_0.1st_Vout_2.t21 bgr_11_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X457 VOUT+.t77 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X458 two_stage_opamp_dummy_magic_23_0.err_amp_out.t11 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t19 GNDA.t577 GNDA.t576 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X459 VDDA.t585 GNDA.t282 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 VOUT-.t74 two_stage_opamp_dummy_magic_23_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 GNDA.t170 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t5 VOUT-.t11 GNDA.t169 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X462 VOUT-.t75 two_stage_opamp_dummy_magic_23_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 two_stage_opamp_dummy_magic_23_0.VD2.t9 GNDA.t537 GNDA.t538 GNDA.t535 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X464 VOUT-.t76 two_stage_opamp_dummy_magic_23_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X465 VOUT+.t78 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X466 VDDA.t101 bgr_11_0.PFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t1 VDDA.t100 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X467 a_7460_6300.t5 two_stage_opamp_dummy_magic_23_0.V_err_gate.t23 VDDA.t169 VDDA.t168 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X468 VDDA.t586 GNDA.t281 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X469 VDDA.t587 GNDA.t280 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t9 bgr_11_0.PFET_GATE_10uA.t19 VDDA.t437 VDDA.t436 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X471 a_7460_6300.t14 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t14 two_stage_opamp_dummy_magic_23_0.V_err_gate.t6 VDDA.t111 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X472 VDDA.t588 GNDA.t279 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X473 GNDA.t483 GNDA.t481 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t8 GNDA.t482 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X474 two_stage_opamp_dummy_magic_23_0.VD1.t0 VIN-.t3 two_stage_opamp_dummy_magic_23_0.V_source.t0 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X475 GNDA.t485 GNDA.t484 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X476 two_stage_opamp_dummy_magic_23_0.V_err_p.t21 two_stage_opamp_dummy_magic_23_0.V_tot.t6 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t16 VDDA.t431 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X477 bgr_11_0.1st_Vout_1.t3 bgr_11_0.Vin+.t8 bgr_11_0.V_p_1.t2 GNDA.t78 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X478 VOUT+.t79 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X479 VOUT-.t77 two_stage_opamp_dummy_magic_23_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X480 VOUT+.t80 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X481 VOUT-.t78 two_stage_opamp_dummy_magic_23_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 VDDA.t589 GNDA.t278 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 VDDA.t1 bgr_11_0.V_mir2.t9 bgr_11_0.V_mir2.t10 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X484 bgr_11_0.1st_Vout_2.t22 bgr_11_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X485 VDDA.t590 GNDA.t277 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X486 VDDA.t591 GNDA.t276 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X487 VDDA.t592 GNDA.t275 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 two_stage_opamp_dummy_magic_23_0.Y.t18 two_stage_opamp_dummy_magic_23_0.Vb2.t20 two_stage_opamp_dummy_magic_23_0.VD4.t33 two_stage_opamp_dummy_magic_23_0.VD4.t32 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X489 VOUT+.t81 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 two_stage_opamp_dummy_magic_23_0.Vb3.t3 bgr_11_0.NFET_GATE_10uA.t14 GNDA.t99 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X491 VDDA.t288 two_stage_opamp_dummy_magic_23_0.Y.t40 VOUT+.t7 VDDA.t287 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X492 VOUT+.t82 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 VDDA.t593 GNDA.t274 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X494 VDDA.t594 GNDA.t273 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X495 GNDA.t93 bgr_11_0.NFET_GATE_10uA.t15 two_stage_opamp_dummy_magic_23_0.Vb3.t2 GNDA.t92 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X496 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t0 two_stage_opamp_dummy_magic_23_0.Vb3.t5 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t1 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X497 bgr_11_0.1st_Vout_1.t22 bgr_11_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 a_4200_4468.t1 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t14 GNDA.t582 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X499 bgr_11_0.1st_Vout_2.t23 bgr_11_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X500 VOUT-.t79 two_stage_opamp_dummy_magic_23_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X501 two_stage_opamp_dummy_magic_23_0.X.t18 two_stage_opamp_dummy_magic_23_0.Vb1.t24 two_stage_opamp_dummy_magic_23_0.VD1.t17 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X502 VDDA.t595 GNDA.t272 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X503 VOUT-.t80 two_stage_opamp_dummy_magic_23_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X504 VDDA.t50 two_stage_opamp_dummy_magic_23_0.Vb3.t18 two_stage_opamp_dummy_magic_23_0.VD4.t3 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X505 VDDA.t179 two_stage_opamp_dummy_magic_23_0.X.t39 VOUT-.t5 VDDA.t178 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X506 bgr_11_0.V_TOP.t33 VDDA.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X507 VDDA.t596 GNDA.t271 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X508 VOUT-.t81 two_stage_opamp_dummy_magic_23_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X509 VOUT-.t82 two_stage_opamp_dummy_magic_23_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 VOUT-.t83 two_stage_opamp_dummy_magic_23_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 VOUT-.t84 two_stage_opamp_dummy_magic_23_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X512 a_5700_24908.t0 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t0 GNDA.t73 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X513 VDDA.t252 two_stage_opamp_dummy_magic_23_0.V_err_gate.t24 a_7460_6300.t4 VDDA.t251 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X514 VDDA.t597 GNDA.t270 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X515 VDDA.t598 GNDA.t269 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X516 VOUT-.t85 two_stage_opamp_dummy_magic_23_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X517 VOUT+.t83 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X518 two_stage_opamp_dummy_magic_23_0.X.t5 two_stage_opamp_dummy_magic_23_0.Vb2.t21 two_stage_opamp_dummy_magic_23_0.VD3.t22 two_stage_opamp_dummy_magic_23_0.VD3.t21 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X519 VDDA.t599 GNDA.t268 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X520 VOUT+.t84 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X521 VDDA.t64 bgr_11_0.1st_Vout_2.t24 bgr_11_0.PFET_GATE_10uA.t6 VDDA.t63 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X522 VDDA.t369 VDDA.t367 two_stage_opamp_dummy_magic_23_0.Vb1.t3 VDDA.t368 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X523 two_stage_opamp_dummy_magic_23_0.Y.t15 GNDA.t534 GNDA.t536 GNDA.t535 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X524 two_stage_opamp_dummy_magic_23_0.V_p_mir.t2 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t21 GNDA.t107 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X525 two_stage_opamp_dummy_magic_23_0.V_source.t16 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t22 GNDA.t32 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X526 two_stage_opamp_dummy_magic_23_0.Vb1.t2 VDDA.t364 VDDA.t366 VDDA.t365 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X527 VDDA.t600 GNDA.t267 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 VOUT+.t85 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X529 GNDA.t485 GNDA.t497 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X530 two_stage_opamp_dummy_magic_23_0.X.t17 two_stage_opamp_dummy_magic_23_0.Vb1.t25 two_stage_opamp_dummy_magic_23_0.VD1.t16 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X531 VDDA.t601 GNDA.t266 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 VDDA.t602 GNDA.t460 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X533 VOUT-.t86 two_stage_opamp_dummy_magic_23_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X534 VOUT-.t87 two_stage_opamp_dummy_magic_23_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X535 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t2 bgr_11_0.PFET_GATE_10uA.t20 VDDA.t12 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X536 GNDA.t178 two_stage_opamp_dummy_magic_23_0.X.t40 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t11 VDDA.t258 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X537 VDDA.t46 bgr_11_0.PFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t1 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X538 GNDA.t600 a_11300_23450.t1 GNDA.t599 sky130_fd_pr__res_xhigh_po_0p35 l=6
X539 two_stage_opamp_dummy_magic_23_0.Y.t20 two_stage_opamp_dummy_magic_23_0.Vb2.t22 two_stage_opamp_dummy_magic_23_0.VD4.t31 two_stage_opamp_dummy_magic_23_0.VD4.t30 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X540 VOUT-.t88 two_stage_opamp_dummy_magic_23_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X541 VOUT+.t86 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X542 VDDA.t603 GNDA.t459 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X543 VDDA.t604 GNDA.t458 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X544 VOUT-.t89 two_stage_opamp_dummy_magic_23_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X545 VDDA.t605 GNDA.t457 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X546 VDDA.t606 GNDA.t456 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 two_stage_opamp_dummy_magic_23_0.VD1.t1 VIN-.t4 two_stage_opamp_dummy_magic_23_0.V_source.t5 GNDA.t72 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X548 bgr_11_0.V_TOP.t34 VDDA.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X549 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t8 two_stage_opamp_dummy_magic_23_0.Y.t41 VDDA.t286 GNDA.t192 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X550 two_stage_opamp_dummy_magic_23_0.V_err_p.t14 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t15 two_stage_opamp_dummy_magic_23_0.err_amp_out.t4 VDDA.t91 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X551 VOUT-.t90 two_stage_opamp_dummy_magic_23_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X552 VOUT+.t87 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X553 VDDA.t607 GNDA.t455 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X554 VDDA.t608 GNDA.t454 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X555 VOUT+.t88 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X556 bgr_11_0.V_TOP.t35 VDDA.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X557 VOUT-.t91 two_stage_opamp_dummy_magic_23_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X558 VDDA.t609 GNDA.t453 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X559 two_stage_opamp_dummy_magic_23_0.VD3.t11 two_stage_opamp_dummy_magic_23_0.Vb3.t19 VDDA.t131 VDDA.t130 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X560 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t8 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t7 GNDA.t597 GNDA.t596 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X561 VOUT+.t89 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X562 two_stage_opamp_dummy_magic_23_0.V_err_p.t8 two_stage_opamp_dummy_magic_23_0.V_err_gate.t25 VDDA.t254 VDDA.t253 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X563 bgr_11_0.1st_Vout_1.t6 bgr_11_0.V_mir1.t19 VDDA.t244 VDDA.t243 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X564 VDDA.t610 GNDA.t452 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X565 VDDA.t611 GNDA.t451 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X566 VDDA.t612 GNDA.t450 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X567 a_7460_6300.t11 two_stage_opamp_dummy_magic_23_0.V_tot.t7 two_stage_opamp_dummy_magic_23_0.V_err_gate.t7 VDDA.t140 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X568 two_stage_opamp_dummy_magic_23_0.VD1.t11 VIN-.t5 two_stage_opamp_dummy_magic_23_0.V_source.t37 GNDA.t82 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X569 VDDA.t613 GNDA.t449 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 two_stage_opamp_dummy_magic_23_0.V_err_p.t17 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t16 two_stage_opamp_dummy_magic_23_0.err_amp_out.t3 VDDA.t455 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X571 VOUT-.t92 two_stage_opamp_dummy_magic_23_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X572 VOUT+.t90 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X573 VDDA.t232 bgr_11_0.V_TOP.t36 bgr_11_0.START_UP.t3 VDDA.t231 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X574 VOUT+.t91 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X575 VOUT-.t93 two_stage_opamp_dummy_magic_23_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X576 VOUT-.t94 two_stage_opamp_dummy_magic_23_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X577 VDDA.t614 GNDA.t448 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X578 VDDA.t230 two_stage_opamp_dummy_magic_23_0.Vb3.t20 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t7 VDDA.t229 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X579 VDDA.t615 GNDA.t447 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X580 VDDA.t285 two_stage_opamp_dummy_magic_23_0.Y.t42 VOUT+.t6 VDDA.t284 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X581 VDDA.t363 VDDA.t361 two_stage_opamp_dummy_magic_23_0.V_err_p.t19 VDDA.t362 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X582 two_stage_opamp_dummy_magic_23_0.X.t6 two_stage_opamp_dummy_magic_23_0.Vb2.t23 two_stage_opamp_dummy_magic_23_0.VD3.t20 two_stage_opamp_dummy_magic_23_0.VD3.t19 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X583 VDDA.t360 VDDA.t358 VOUT+.t13 VDDA.t359 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X584 VOUT+.t92 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X585 bgr_11_0.V_p_2.t4 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t17 bgr_11_0.V_mir2.t16 GNDA.t593 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X586 GNDA.t533 GNDA.t532 two_stage_opamp_dummy_magic_23_0.VD1.t10 GNDA.t528 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X587 VDDA.t616 GNDA.t446 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X588 two_stage_opamp_dummy_magic_23_0.VD4.t29 two_stage_opamp_dummy_magic_23_0.Vb2.t24 two_stage_opamp_dummy_magic_23_0.Y.t1 two_stage_opamp_dummy_magic_23_0.VD4.t28 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X589 VOUT-.t95 two_stage_opamp_dummy_magic_23_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X590 VDDA.t617 GNDA.t445 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X591 VOUT+.t93 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X592 VOUT+.t94 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X593 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t4 bgr_11_0.PFET_GATE_10uA.t22 VDDA.t129 VDDA.t128 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X594 VOUT+.t95 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X595 VDDA.t618 GNDA.t444 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X596 VDDA.t619 GNDA.t443 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X597 two_stage_opamp_dummy_magic_23_0.VD3.t2 two_stage_opamp_dummy_magic_23_0.VD3.t0 two_stage_opamp_dummy_magic_23_0.X.t3 two_stage_opamp_dummy_magic_23_0.VD3.t1 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X598 two_stage_opamp_dummy_magic_23_0.X.t24 two_stage_opamp_dummy_magic_23_0.Vb1.t26 two_stage_opamp_dummy_magic_23_0.VD1.t15 GNDA.t72 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X599 VDDA.t620 GNDA.t442 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X600 VOUT+.t96 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X601 VDDA.t228 bgr_11_0.V_mir2.t7 bgr_11_0.V_mir2.t8 VDDA.t227 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X602 VOUT+.t97 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X603 VDDA.t425 bgr_11_0.V_mir1.t4 bgr_11_0.V_mir1.t5 VDDA.t424 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X604 VOUT+.t17 a_4600_1446.t1 GNDA.t592 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X605 VOUT+.t98 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X606 two_stage_opamp_dummy_magic_23_0.VD3.t36 two_stage_opamp_dummy_magic_23_0.Vb3.t21 VDDA.t454 VDDA.t453 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X607 VDDA.t259 two_stage_opamp_dummy_magic_23_0.X.t41 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t9 GNDA.t179 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X608 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t1 a_13130_1456.t0 GNDA.t134 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X609 GNDA.t531 GNDA.t530 two_stage_opamp_dummy_magic_23_0.VD2.t8 GNDA.t525 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X610 VDDA.t621 GNDA.t441 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X611 VDDA.t622 GNDA.t440 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X612 VOUT+.t99 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X613 VDDA.t623 GNDA.t439 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X614 two_stage_opamp_dummy_magic_23_0.V_source.t15 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t23 GNDA.t585 GNDA.t584 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X615 two_stage_opamp_dummy_magic_23_0.X.t23 two_stage_opamp_dummy_magic_23_0.Vb1.t27 two_stage_opamp_dummy_magic_23_0.VD1.t14 GNDA.t82 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X616 VOUT+.t100 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X617 two_stage_opamp_dummy_magic_23_0.V_source.t40 two_stage_opamp_dummy_magic_23_0.Vb1.t28 a_8260_1600.t0 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.6 ps=3.8 w=1.5 l=3
X618 VOUT-.t96 two_stage_opamp_dummy_magic_23_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X619 VDDA.t624 GNDA.t438 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X620 GNDA.t142 two_stage_opamp_dummy_magic_23_0.X.t42 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t10 VDDA.t175 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X621 VDDA.t625 GNDA.t437 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X622 VOUT-.t97 two_stage_opamp_dummy_magic_23_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X623 VDDA.t626 GNDA.t436 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X624 VOUT-.t98 two_stage_opamp_dummy_magic_23_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X625 VOUT-.t99 two_stage_opamp_dummy_magic_23_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X626 bgr_11_0.1st_Vout_1.t23 bgr_11_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X627 VOUT+.t101 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X628 VOUT+.t102 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X629 VDDA.t627 GNDA.t435 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X630 VDDA.t628 GNDA.t434 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X631 VDDA.t629 GNDA.t433 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X632 GNDA.t529 GNDA.t527 two_stage_opamp_dummy_magic_23_0.X.t14 GNDA.t528 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X633 VOUT+.t103 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X634 VOUT+.t104 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X635 VOUT+.t105 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X636 bgr_11_0.Vin-.t1 bgr_11_0.START_UP.t7 bgr_11_0.V_TOP.t1 VDDA.t157 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X637 VDDA.t630 GNDA.t432 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X638 VDDA.t631 GNDA.t431 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X639 bgr_11_0.1st_Vout_1.t24 bgr_11_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X640 VDDA.t632 GNDA.t430 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X641 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t5 bgr_11_0.V_TOP.t37 VDDA.t234 VDDA.t233 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X642 two_stage_opamp_dummy_magic_23_0.V_err_p.t18 VDDA.t355 VDDA.t357 VDDA.t356 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X643 two_stage_opamp_dummy_magic_23_0.V_err_p.t7 two_stage_opamp_dummy_magic_23_0.V_err_gate.t26 VDDA.t264 VDDA.t263 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X644 two_stage_opamp_dummy_magic_23_0.err_amp_out.t7 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t20 GNDA.t159 GNDA.t158 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X645 VDDA.t42 bgr_11_0.1st_Vout_2.t25 bgr_11_0.PFET_GATE_10uA.t5 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X646 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t6 two_stage_opamp_dummy_magic_23_0.Y.t43 GNDA.t185 VDDA.t283 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X647 GNDA.t526 GNDA.t524 two_stage_opamp_dummy_magic_23_0.Y.t24 GNDA.t525 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X648 VOUT-.t100 two_stage_opamp_dummy_magic_23_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X649 GNDA.t523 GNDA.t521 two_stage_opamp_dummy_magic_23_0.Vb2.t7 GNDA.t522 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X650 two_stage_opamp_dummy_magic_23_0.VD4.t16 VDDA.t352 VDDA.t354 VDDA.t353 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X651 two_stage_opamp_dummy_magic_23_0.VD1.t9 GNDA.t519 GNDA.t520 GNDA.t515 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X652 VOUT-.t101 two_stage_opamp_dummy_magic_23_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X653 VOUT-.t102 two_stage_opamp_dummy_magic_23_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X654 VOUT+.t106 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X655 GNDA.t485 GNDA.t513 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X656 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t1 bgr_11_0.NFET_GATE_10uA.t16 GNDA.t95 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X657 GNDA.t6 bgr_11_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t0 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X658 two_stage_opamp_dummy_magic_23_0.VD4.t27 two_stage_opamp_dummy_magic_23_0.Vb2.t25 two_stage_opamp_dummy_magic_23_0.Y.t2 two_stage_opamp_dummy_magic_23_0.VD4.t26 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X659 two_stage_opamp_dummy_magic_23_0.V_err_p.t20 two_stage_opamp_dummy_magic_23_0.V_tot.t8 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t15 VDDA.t426 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X660 VOUT+.t107 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X661 VDDA.t633 GNDA.t429 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X662 bgr_11_0.V_p_2.t2 bgr_11_0.V_CUR_REF_REG.t5 bgr_11_0.1st_Vout_2.t4 GNDA.t121 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X663 VDDA.t634 GNDA.t428 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X664 a_6350_25058.t1 a_6470_23450.t1 GNDA.t35 sky130_fd_pr__res_xhigh_po_0p35 l=6
X665 VOUT+.t108 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X666 bgr_11_0.1st_Vout_1.t25 bgr_11_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X667 a_4080_4468.t0 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t0 GNDA.t0 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X668 VDDA.t635 GNDA.t475 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X669 VDDA.t636 GNDA.t474 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X670 two_stage_opamp_dummy_magic_23_0.VD3.t37 two_stage_opamp_dummy_magic_23_0.Vb3.t22 VDDA.t467 VDDA.t466 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X671 a_13450_4368.t0 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t4 GNDA.t579 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X672 VDDA.t637 GNDA.t473 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X673 VDDA.t282 two_stage_opamp_dummy_magic_23_0.Y.t44 VOUT+.t5 VDDA.t281 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X674 bgr_11_0.V_TOP.t38 VDDA.t434 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X675 VOUT+.t109 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X676 VDDA.t351 VDDA.t349 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t2 VDDA.t350 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X677 two_stage_opamp_dummy_magic_23_0.err_amp_out.t2 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t18 two_stage_opamp_dummy_magic_23_0.V_err_p.t15 VDDA.t104 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X678 VDDA.t638 GNDA.t472 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X679 VDDA.t8 bgr_11_0.V_mir2.t20 bgr_11_0.1st_Vout_2.t1 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X680 bgr_11_0.1st_Vout_1.t26 bgr_11_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X681 two_stage_opamp_dummy_magic_23_0.VD3.t18 two_stage_opamp_dummy_magic_23_0.Vb2.t26 two_stage_opamp_dummy_magic_23_0.X.t1 two_stage_opamp_dummy_magic_23_0.VD3.t17 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X682 VDDA.t639 GNDA.t471 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X683 VDDA.t640 GNDA.t470 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X684 GNDA.t184 two_stage_opamp_dummy_magic_23_0.Y.t45 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t5 VDDA.t280 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X685 VDDA.t176 two_stage_opamp_dummy_magic_23_0.X.t43 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t8 GNDA.t143 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X686 bgr_11_0.cap_res2.t20 bgr_11_0.PFET_GATE_10uA.t9 GNDA.t578 sky130_fd_pr__res_high_po_0p35 l=2.05
X687 two_stage_opamp_dummy_magic_23_0.V_source.t27 VIN+.t6 two_stage_opamp_dummy_magic_23_0.VD2.t3 GNDA.t50 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X688 VOUT-.t103 two_stage_opamp_dummy_magic_23_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X689 VOUT+.t110 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X690 VDDA.t641 GNDA.t469 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X691 two_stage_opamp_dummy_magic_23_0.V_err_gate.t13 two_stage_opamp_dummy_magic_23_0.V_tot.t9 a_7460_6300.t19 VDDA.t468 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X692 VOUT-.t104 two_stage_opamp_dummy_magic_23_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X693 VOUT-.t105 two_stage_opamp_dummy_magic_23_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X694 VDDA.t642 GNDA.t468 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X695 GNDA.t485 GNDA.t518 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X696 two_stage_opamp_dummy_magic_23_0.VD4.t25 two_stage_opamp_dummy_magic_23_0.Vb2.t27 two_stage_opamp_dummy_magic_23_0.Y.t13 two_stage_opamp_dummy_magic_23_0.VD4.t24 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X697 two_stage_opamp_dummy_magic_23_0.V_source.t14 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t24 GNDA.t30 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X698 GNDA.t485 GNDA.t517 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X699 two_stage_opamp_dummy_magic_23_0.X.t13 GNDA.t514 GNDA.t516 GNDA.t515 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X700 two_stage_opamp_dummy_magic_23_0.Vb1.t9 two_stage_opamp_dummy_magic_23_0.Vb1.t8 a_8260_1600.t2 GNDA.t75 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X701 GNDA.t140 two_stage_opamp_dummy_magic_23_0.X.t44 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t9 VDDA.t173 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X702 VOUT+.t111 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X703 GNDA.t141 two_stage_opamp_dummy_magic_23_0.X.t45 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t8 VDDA.t174 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X704 VDDA.t643 GNDA.t467 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X705 VDDA.t644 GNDA.t466 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X706 VDDA.t645 GNDA.t465 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X707 bgr_11_0.V_TOP.t39 VDDA.t435 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X708 VDDA.t646 GNDA.t464 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X709 VOUT-.t106 two_stage_opamp_dummy_magic_23_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X710 VOUT+.t112 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X711 bgr_11_0.V_p_2.t8 bgr_11_0.V_CUR_REF_REG.t6 bgr_11_0.1st_Vout_2.t6 GNDA.t157 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X712 VDDA.t647 GNDA.t463 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X713 VDDA.t222 bgr_11_0.V_TOP.t40 bgr_11_0.Vin-.t5 VDDA.t221 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X714 bgr_11_0.1st_Vout_2.t26 bgr_11_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X715 GNDA.t462 VDDA.t648 bgr_11_0.V_TOP.t7 GNDA.t461 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X716 VDDA.t649 GNDA.t427 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X717 VDDA.t348 VDDA.t345 VDDA.t347 VDDA.t346 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0 ps=0 w=1.8 l=0.2
X718 VDDA.t125 two_stage_opamp_dummy_magic_23_0.Vb3.t23 two_stage_opamp_dummy_magic_23_0.VD3.t10 VDDA.t124 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X719 VOUT-.t4 two_stage_opamp_dummy_magic_23_0.X.t46 VDDA.t171 VDDA.t170 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X720 bgr_11_0.NFET_GATE_10uA.t1 bgr_11_0.NFET_GATE_10uA.t0 GNDA.t86 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X721 GNDA.t8 bgr_11_0.NFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_23_0.Vb3.t1 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X722 bgr_11_0.V_p_1.t8 bgr_11_0.Vin-.t10 bgr_11_0.V_mir1.t12 GNDA.t461 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X723 VDDA.t650 GNDA.t426 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X724 VOUT-.t107 two_stage_opamp_dummy_magic_23_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X725 VDDA.t99 bgr_11_0.V_mir2.t5 bgr_11_0.V_mir2.t6 VDDA.t98 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X726 a_7460_6300.t3 two_stage_opamp_dummy_magic_23_0.V_err_gate.t27 VDDA.t266 VDDA.t265 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X727 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t6 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t5 GNDA.t174 GNDA.t173 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X728 bgr_11_0.1st_Vout_2.t27 bgr_11_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X729 VDDA.t651 GNDA.t425 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X730 VOUT-.t108 two_stage_opamp_dummy_magic_23_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X731 VDDA.t652 GNDA.t424 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X732 two_stage_opamp_dummy_magic_23_0.VD2.t15 two_stage_opamp_dummy_magic_23_0.Vb1.t29 two_stage_opamp_dummy_magic_23_0.Y.t10 GNDA.t50 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X733 GNDA.t62 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t25 two_stage_opamp_dummy_magic_23_0.V_source.t13 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X734 GNDA.t118 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t26 two_stage_opamp_dummy_magic_23_0.V_source.t12 GNDA.t117 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X735 bgr_11_0.V_p_1.t5 VDDA.t653 GNDA.t423 GNDA.t422 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X736 VDDA.t119 bgr_11_0.PFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t0 VDDA.t118 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X737 VDDA.t344 VDDA.t342 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t12 VDDA.t343 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X738 VDDA.t654 GNDA.t265 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X739 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t1 bgr_11_0.PFET_GATE_10uA.t24 VDDA.t226 VDDA.t225 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X740 VDDA.t341 VDDA.t339 VDDA.t341 VDDA.t340 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X741 bgr_11_0.1st_Vout_1.t27 bgr_11_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X742 VDDA.t655 GNDA.t264 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X743 bgr_11_0.V_p_2.t0 bgr_11_0.V_CUR_REF_REG.t7 bgr_11_0.1st_Vout_2.t0 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X744 bgr_11_0.1st_Vout_2.t28 bgr_11_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X745 VOUT+.t113 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X746 VDDA.t656 GNDA.t263 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X747 a_12070_24908.t0 a_11950_23700.t0 GNDA.t84 sky130_fd_pr__res_xhigh_po_0p35 l=4
X748 two_stage_opamp_dummy_magic_23_0.VD3.t16 two_stage_opamp_dummy_magic_23_0.Vb2.t28 two_stage_opamp_dummy_magic_23_0.X.t2 two_stage_opamp_dummy_magic_23_0.VD3.t15 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X749 VOUT-.t109 two_stage_opamp_dummy_magic_23_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X750 VOUT+.t114 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X751 VOUT+.t115 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X752 VDDA.t657 GNDA.t262 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X753 VDDA.t250 bgr_11_0.V_mir1.t20 bgr_11_0.1st_Vout_1.t7 VDDA.t249 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X754 VDDA.t658 GNDA.t261 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X755 bgr_11_0.1st_Vout_1.t28 bgr_11_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X756 VDDA.t86 two_stage_opamp_dummy_magic_23_0.Vb3.t24 two_stage_opamp_dummy_magic_23_0.VD3.t8 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X757 VDDA.t659 GNDA.t260 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X758 VOUT-.t110 two_stage_opamp_dummy_magic_23_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X759 VDDA.t660 GNDA.t259 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X760 VOUT-.t111 two_stage_opamp_dummy_magic_23_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X761 two_stage_opamp_dummy_magic_23_0.Vb2.t2 two_stage_opamp_dummy_magic_23_0.Vb2_2.t0 two_stage_opamp_dummy_magic_23_0.Vb2_2.t2 two_stage_opamp_dummy_magic_23_0.Vb2_2.t1 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X762 VOUT-.t112 two_stage_opamp_dummy_magic_23_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X763 two_stage_opamp_dummy_magic_23_0.Vb2.t0 bgr_11_0.NFET_GATE_10uA.t19 GNDA.t11 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X764 VOUT+.t2 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t6 GNDA.t182 GNDA.t181 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X765 bgr_11_0.1st_Vout_2.t29 bgr_11_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X766 VDDA.t661 GNDA.t258 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X767 VOUT-.t113 two_stage_opamp_dummy_magic_23_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X768 VOUT-.t114 two_stage_opamp_dummy_magic_23_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X769 GNDA.t13 bgr_11_0.NFET_GATE_10uA.t20 two_stage_opamp_dummy_magic_23_0.Vb2.t1 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X770 bgr_11_0.Vin-.t4 bgr_11_0.V_TOP.t41 VDDA.t224 VDDA.t223 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X771 two_stage_opamp_dummy_magic_23_0.V_source.t4 VIN+.t7 two_stage_opamp_dummy_magic_23_0.VD2.t2 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X772 VDDA.t172 two_stage_opamp_dummy_magic_23_0.X.t47 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t7 GNDA.t139 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X773 VOUT-.t115 two_stage_opamp_dummy_magic_23_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X774 two_stage_opamp_dummy_magic_23_0.V_err_gate.t8 two_stage_opamp_dummy_magic_23_0.V_tot.t10 a_7460_6300.t17 VDDA.t240 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X775 GNDA.t191 two_stage_opamp_dummy_magic_23_0.Y.t46 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t4 VDDA.t279 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X776 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t7 GNDA.t511 GNDA.t512 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X777 VOUT+.t116 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X778 VOUT+.t117 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X779 two_stage_opamp_dummy_magic_23_0.V_err_gate.t12 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t19 a_7460_6300.t13 VDDA.t442 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X780 VDDA.t662 GNDA.t257 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X781 VDDA.t663 GNDA.t256 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X782 VOUT+.t118 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X783 bgr_11_0.1st_Vout_1.t29 bgr_11_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X784 VDDA.t664 GNDA.t255 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X785 two_stage_opamp_dummy_magic_23_0.V_source.t11 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t27 GNDA.t60 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X786 bgr_11_0.1st_Vout_2.t30 bgr_11_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X787 VDDA.t665 GNDA.t254 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X788 two_stage_opamp_dummy_magic_23_0.Vb1.t7 two_stage_opamp_dummy_magic_23_0.Vb1.t6 a_8260_1600.t1 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X789 VDDA.t666 GNDA.t253 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X790 GNDA.t421 VDDA.t336 VDDA.t338 VDDA.t337 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X791 VOUT+.t119 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X792 VOUT-.t116 two_stage_opamp_dummy_magic_23_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X793 VDDA.t335 VDDA.t333 bgr_11_0.V_TOP.t4 VDDA.t334 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X794 VDDA.t332 VDDA.t330 two_stage_opamp_dummy_magic_23_0.Vb2_2.t6 VDDA.t331 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.36 ps=2.2 w=1.8 l=0.2
X795 VOUT-.t117 two_stage_opamp_dummy_magic_23_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X796 VDDA.t667 GNDA.t420 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X797 VDDA.t668 GNDA.t419 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X798 bgr_11_0.1st_Vout_1.t30 bgr_11_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X799 VDDA.t669 GNDA.t418 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X800 VOUT-.t118 two_stage_opamp_dummy_magic_23_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X801 VDDA.t670 GNDA.t417 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X802 VDDA.t671 GNDA.t416 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X803 VDDA.t672 GNDA.t415 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X804 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t7 two_stage_opamp_dummy_magic_23_0.Y.t47 VDDA.t277 GNDA.t190 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X805 VOUT-.t119 two_stage_opamp_dummy_magic_23_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X806 VDDA.t673 GNDA.t414 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X807 VDDA.t674 GNDA.t413 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X808 VOUT-.t120 two_stage_opamp_dummy_magic_23_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X809 VDDA.t115 bgr_11_0.1st_Vout_1.t31 bgr_11_0.V_TOP.t10 VDDA.t114 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X810 VOUT-.t3 two_stage_opamp_dummy_magic_23_0.X.t48 VDDA.t164 VDDA.t163 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X811 VOUT+.t120 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X812 VOUT+.t121 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X813 VOUT+.t122 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X814 VDDA.t90 two_stage_opamp_dummy_magic_23_0.Vb3.t25 two_stage_opamp_dummy_magic_23_0.VD4.t2 VDDA.t89 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X815 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t4 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t3 GNDA.t116 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X816 VDDA.t329 VDDA.t327 bgr_11_0.NFET_GATE_10uA.t2 VDDA.t328 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X817 VDDA.t675 GNDA.t412 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X818 VOUT+.t123 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X819 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t5 bgr_11_0.PFET_GATE_10uA.t25 VDDA.t150 VDDA.t149 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X820 two_stage_opamp_dummy_magic_23_0.Y.t14 two_stage_opamp_dummy_magic_23_0.Vb2.t29 two_stage_opamp_dummy_magic_23_0.VD4.t23 two_stage_opamp_dummy_magic_23_0.VD4.t22 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X821 two_stage_opamp_dummy_magic_23_0.V_err_p.t6 two_stage_opamp_dummy_magic_23_0.V_err_gate.t28 VDDA.t200 VDDA.t199 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X822 two_stage_opamp_dummy_magic_23_0.VD2.t14 two_stage_opamp_dummy_magic_23_0.Vb1.t30 two_stage_opamp_dummy_magic_23_0.Y.t11 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X823 VOUT-.t121 two_stage_opamp_dummy_magic_23_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X824 VDDA.t676 GNDA.t411 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X825 VDDA.t677 GNDA.t410 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X826 VDDA.t678 GNDA.t409 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X827 VDDA.t679 GNDA.t408 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X828 GNDA.t4 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t28 two_stage_opamp_dummy_magic_23_0.V_source.t10 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X829 VOUT-.t122 two_stage_opamp_dummy_magic_23_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X830 VOUT-.t123 two_stage_opamp_dummy_magic_23_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X831 VOUT+.t124 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X832 VDDA.t680 GNDA.t407 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X833 VDDA.t681 GNDA.t406 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X834 VDDA.t326 VDDA.t324 two_stage_opamp_dummy_magic_23_0.VD3.t13 VDDA.t325 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X835 a_13570_4368.t1 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t4 GNDA.t160 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X836 bgr_11_0.V_TOP.t42 VDDA.t237 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X837 VDDA.t682 GNDA.t405 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X838 VOUT-.t124 two_stage_opamp_dummy_magic_23_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X839 VOUT-.t125 two_stage_opamp_dummy_magic_23_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X840 VDDA.t683 GNDA.t404 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X841 VOUT-.t126 two_stage_opamp_dummy_magic_23_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X842 GNDA.t125 bgr_11_0.NFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_23_0.Vb3.t0 GNDA.t124 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X843 VDDA.t268 bgr_11_0.V_mir1.t2 bgr_11_0.V_mir1.t3 VDDA.t267 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X844 VDDA.t239 bgr_11_0.V_TOP.t43 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t4 VDDA.t238 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X845 VOUT+.t125 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X846 VDDA.t278 two_stage_opamp_dummy_magic_23_0.Y.t48 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t6 GNDA.t189 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X847 VDDA.t684 GNDA.t403 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X848 VOUT-.t127 two_stage_opamp_dummy_magic_23_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X849 VDDA.t685 GNDA.t402 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X850 bgr_11_0.V_p_1.t7 bgr_11_0.Vin-.t11 bgr_11_0.V_mir1.t13 GNDA.t587 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X851 VDDA.t686 GNDA.t401 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X852 bgr_11_0.V_TOP.t44 VDDA.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X853 VDDA.t108 bgr_11_0.1st_Vout_1.t32 bgr_11_0.V_TOP.t9 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X854 GNDA.t603 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t7 VOUT-.t18 GNDA.t602 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X855 VOUT+.t126 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X856 VOUT+.t127 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X857 VOUT+.t128 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X858 bgr_11_0.PFET_GATE_10uA.t2 VDDA.t687 GNDA.t400 GNDA.t114 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X859 VDDA.t688 GNDA.t252 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X860 VOUT+.t129 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X861 VOUT-.t128 two_stage_opamp_dummy_magic_23_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X862 VDDA.t165 two_stage_opamp_dummy_magic_23_0.X.t49 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t6 GNDA.t138 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X863 VOUT+.t130 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X864 VDDA.t202 two_stage_opamp_dummy_magic_23_0.V_err_gate.t29 two_stage_opamp_dummy_magic_23_0.V_err_p.t5 VDDA.t201 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X865 two_stage_opamp_dummy_magic_23_0.V_source.t39 VIN+.t8 two_stage_opamp_dummy_magic_23_0.VD2.t11 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X866 VDDA.t689 GNDA.t251 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X867 VDDA.t690 GNDA.t250 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X868 VDDA.t196 two_stage_opamp_dummy_magic_23_0.V_err_gate.t30 two_stage_opamp_dummy_magic_23_0.V_err_p.t4 VDDA.t195 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X869 VDDA.t255 two_stage_opamp_dummy_magic_23_0.X.t50 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t5 GNDA.t177 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X870 VOUT-.t129 two_stage_opamp_dummy_magic_23_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X871 two_stage_opamp_dummy_magic_23_0.Y.t0 two_stage_opamp_dummy_magic_23_0.Vb2.t30 two_stage_opamp_dummy_magic_23_0.VD4.t21 two_stage_opamp_dummy_magic_23_0.VD4.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X872 two_stage_opamp_dummy_magic_23_0.V_err_gate.t1 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t20 a_7460_6300.t12 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X873 GNDA.t188 two_stage_opamp_dummy_magic_23_0.Y.t49 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t3 VDDA.t276 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X874 VOUT-.t130 two_stage_opamp_dummy_magic_23_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X875 two_stage_opamp_dummy_magic_23_0.Vb1.t0 bgr_11_0.PFET_GATE_10uA.t26 VDDA.t10 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X876 VDDA.t691 GNDA.t249 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X877 VOUT-.t131 two_stage_opamp_dummy_magic_23_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X878 VOUT+.t131 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X879 bgr_11_0.PFET_GATE_10uA.t4 bgr_11_0.1st_Vout_2.t31 VDDA.t80 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X880 two_stage_opamp_dummy_magic_23_0.Vb1.t4 GNDA.t508 GNDA.t510 GNDA.t509 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X881 VOUT-.t132 two_stage_opamp_dummy_magic_23_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X882 VDDA.t692 GNDA.t248 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X883 VDDA.t148 bgr_11_0.PFET_GATE_10uA.t27 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t0 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X884 VDDA.t693 GNDA.t247 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X885 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t5 VDDA.t321 VDDA.t323 VDDA.t322 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X886 VDDA.t694 GNDA.t246 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X887 VOUT+.t132 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X888 bgr_11_0.V_p_1.t6 bgr_11_0.Vin-.t12 bgr_11_0.V_mir1.t15 GNDA.t598 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X889 GNDA.t507 GNDA.t505 VOUT-.t17 GNDA.t506 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X890 VOUT-.t133 two_stage_opamp_dummy_magic_23_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X891 VDDA.t236 bgr_11_0.V_mir1.t0 bgr_11_0.V_mir1.t1 VDDA.t235 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X892 VDDA.t695 GNDA.t245 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X893 VOUT-.t134 two_stage_opamp_dummy_magic_23_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X894 VOUT-.t135 two_stage_opamp_dummy_magic_23_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X895 VDDA.t696 GNDA.t244 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X896 two_stage_opamp_dummy_magic_23_0.Vb2_2.t9 two_stage_opamp_dummy_magic_23_0.Vb2.t31 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.36 ps=2.2 w=1.8 l=0.2
X897 VOUT+.t133 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X898 two_stage_opamp_dummy_magic_23_0.VD3.t35 two_stage_opamp_dummy_magic_23_0.Vb3.t26 VDDA.t452 VDDA.t451 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X899 bgr_11_0.V_TOP.t45 VDDA.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X900 VDDA.t697 GNDA.t243 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X901 VOUT+.t134 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X902 VDDA.t82 bgr_11_0.1st_Vout_2.t32 bgr_11_0.PFET_GATE_10uA.t3 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X903 VOUT+.t135 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X904 GNDA.t595 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t8 VOUT+.t18 GNDA.t594 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X905 VOUT+.t136 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X906 VOUT+.t137 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X907 VOUT-.t136 two_stage_opamp_dummy_magic_23_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X908 VDDA.t698 GNDA.t242 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X909 VOUT-.t12 two_stage_opamp_dummy_magic_23_0.X.t51 VDDA.t257 VDDA.t256 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X910 VDDA.t699 GNDA.t241 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X911 VDDA.t700 GNDA.t240 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X912 a_13450_4368.t1 two_stage_opamp_dummy_magic_23_0.V_tot.t3 GNDA.t583 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X913 two_stage_opamp_dummy_magic_23_0.err_amp_out.t10 GNDA.t502 GNDA.t504 GNDA.t503 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X914 bgr_11_0.V_p_2.t3 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t21 bgr_11_0.V_mir2.t1 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X915 VOUT-.t137 two_stage_opamp_dummy_magic_23_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X916 a_7460_6300.t2 two_stage_opamp_dummy_magic_23_0.V_err_gate.t31 VDDA.t198 VDDA.t197 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X917 two_stage_opamp_dummy_magic_23_0.VD2.t13 two_stage_opamp_dummy_magic_23_0.Vb1.t31 two_stage_opamp_dummy_magic_23_0.Y.t12 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X918 GNDA.t485 GNDA.t501 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X919 VOUT-.t138 two_stage_opamp_dummy_magic_23_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X920 VDDA.t701 GNDA.t239 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X921 GNDA.t105 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t29 two_stage_opamp_dummy_magic_23_0.V_source.t9 GNDA.t104 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X922 bgr_11_0.1st_Vout_2.t33 bgr_11_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X923 VDDA.t702 GNDA.t238 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X924 VOUT-.t139 two_stage_opamp_dummy_magic_23_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X925 VOUT-.t140 two_stage_opamp_dummy_magic_23_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X926 VOUT-.t141 two_stage_opamp_dummy_magic_23_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X927 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t3 GNDA.t498 GNDA.t500 GNDA.t499 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X928 VDDA.t320 VDDA.t318 GNDA.t399 VDDA.t319 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X929 VDDA.t703 GNDA.t237 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X930 bgr_11_0.V_p_1.t1 bgr_11_0.Vin+.t9 bgr_11_0.1st_Vout_1.t2 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X931 VDDA.t704 GNDA.t236 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X932 GNDA.t47 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t9 VOUT+.t1 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X933 bgr_11_0.1st_Vout_1.t33 bgr_11_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X934 VDDA.t705 GNDA.t235 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X935 VOUT+.t138 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X936 VDDA.t439 bgr_11_0.V_mir2.t21 bgr_11_0.1st_Vout_2.t8 VDDA.t438 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X937 VDDA.t706 GNDA.t234 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X938 VDDA.t707 GNDA.t233 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X939 VOUT-.t142 two_stage_opamp_dummy_magic_23_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X940 VOUT+.t139 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X941 VDDA.t275 two_stage_opamp_dummy_magic_23_0.Y.t50 VOUT+.t4 VDDA.t274 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X942 two_stage_opamp_dummy_magic_23_0.Vb2_2.t8 two_stage_opamp_dummy_magic_23_0.Vb2.t9 two_stage_opamp_dummy_magic_23_0.Vb2.t10 two_stage_opamp_dummy_magic_23_0.Vb2_2.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X943 VDDA.t273 two_stage_opamp_dummy_magic_23_0.Y.t51 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t5 GNDA.t187 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X944 two_stage_opamp_dummy_magic_23_0.V_source.t6 VIN-.t6 two_stage_opamp_dummy_magic_23_0.VD1.t2 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X945 VOUT+.t140 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X946 VDDA.t708 GNDA.t232 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X947 VDDA.t446 bgr_11_0.PFET_GATE_10uA.t28 bgr_11_0.V_CUR_REF_REG.t0 VDDA.t445 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X948 VDDA.t709 GNDA.t231 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X949 VDDA.t463 bgr_11_0.PFET_GATE_10uA.t29 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t11 VDDA.t462 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X950 GNDA.t176 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t21 two_stage_opamp_dummy_magic_23_0.err_amp_out.t8 GNDA.t175 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X951 VOUT-.t143 two_stage_opamp_dummy_magic_23_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X952 VDDA.t44 GNDA.t494 GNDA.t496 GNDA.t495 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X953 VOUT-.t144 two_stage_opamp_dummy_magic_23_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X954 VDDA.t192 two_stage_opamp_dummy_magic_23_0.V_err_gate.t32 a_7460_6300.t1 VDDA.t191 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X955 two_stage_opamp_dummy_magic_23_0.V_source.t3 VIN+.t9 two_stage_opamp_dummy_magic_23_0.VD2.t1 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X956 VOUT-.t145 two_stage_opamp_dummy_magic_23_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X957 VOUT+.t141 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X958 VDDA.t710 GNDA.t230 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X959 a_5700_24908.t1 a_5820_23634.t1 GNDA.t73 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X960 two_stage_opamp_dummy_magic_23_0.V_err_gate.t9 two_stage_opamp_dummy_magic_23_0.V_tot.t11 a_7460_6300.t18 VDDA.t248 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X961 VDDA.t711 GNDA.t229 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X962 GNDA.t186 two_stage_opamp_dummy_magic_23_0.Y.t52 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t2 VDDA.t272 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X963 two_stage_opamp_dummy_magic_23_0.V_source.t7 VIN-.t7 two_stage_opamp_dummy_magic_23_0.VD1.t3 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X964 bgr_11_0.V_TOP.t46 VDDA.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X965 GNDA.t485 GNDA.t493 bgr_11_0.Vin-.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X966 VDDA.t712 GNDA.t228 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X967 bgr_11_0.V_mir2.t4 bgr_11_0.V_mir2.t3 VDDA.t117 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X968 VOUT+.t142 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X969 bgr_11_0.1st_Vout_1.t34 bgr_11_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X970 VOUT+.t143 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X971 VOUT+.t144 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X972 VDDA.t713 GNDA.t227 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X973 VDDA.t714 GNDA.t226 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X974 VDDA.t715 GNDA.t225 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X975 VDDA.t716 GNDA.t224 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X976 VDDA.t717 GNDA.t223 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X977 VOUT+.t145 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X978 VOUT+.t3 two_stage_opamp_dummy_magic_23_0.Y.t53 VDDA.t271 VDDA.t270 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X979 VOUT+.t146 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X980 VOUT+.t147 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X981 VOUT+.t148 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X982 a_11420_25058.t0 a_11300_23450.t0 GNDA.t1 sky130_fd_pr__res_xhigh_po_0p35 l=6
X983 VDDA.t718 GNDA.t222 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X984 VDDA.t719 GNDA.t221 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X985 VOUT-.t16 GNDA.t490 GNDA.t492 GNDA.t491 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X986 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_23_0.Y.t16 GNDA.t90 sky130_fd_pr__res_high_po_1p41 l=1.41
X987 VDDA.t720 GNDA.t220 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X988 VDDA.t55 bgr_11_0.V_TOP.t47 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t3 VDDA.t54 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X989 two_stage_opamp_dummy_magic_23_0.VD4.t1 two_stage_opamp_dummy_magic_23_0.Vb3.t27 VDDA.t14 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X990 two_stage_opamp_dummy_magic_23_0.VD1.t13 two_stage_opamp_dummy_magic_23_0.Vb1.t32 two_stage_opamp_dummy_magic_23_0.X.t22 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X991 VOUT-.t1 two_stage_opamp_dummy_magic_23_0.X.t52 VDDA.t160 VDDA.t159 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X992 VOUT+.t149 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X993 VOUT-.t146 two_stage_opamp_dummy_magic_23_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X994 bgr_11_0.V_TOP.t3 VDDA.t315 VDDA.t317 VDDA.t316 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.45 ps=2.9 w=1 l=0.15
X995 two_stage_opamp_dummy_magic_23_0.VD4.t19 two_stage_opamp_dummy_magic_23_0.Vb2.t32 two_stage_opamp_dummy_magic_23_0.Y.t21 two_stage_opamp_dummy_magic_23_0.VD4.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X996 VOUT-.t2 two_stage_opamp_dummy_magic_23_0.X.t53 VDDA.t162 VDDA.t161 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X997 VOUT-.t147 two_stage_opamp_dummy_magic_23_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X998 VOUT-.t148 two_stage_opamp_dummy_magic_23_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X999 VDDA.t721 GNDA.t219 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1000 VOUT-.t149 two_stage_opamp_dummy_magic_23_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1001 VDDA.t722 GNDA.t218 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1002 VOUT-.t150 two_stage_opamp_dummy_magic_23_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1003 VDDA.t723 GNDA.t217 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1004 two_stage_opamp_dummy_magic_23_0.VD2.t12 two_stage_opamp_dummy_magic_23_0.Vb1.t33 two_stage_opamp_dummy_magic_23_0.Y.t4 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1005 GNDA.t103 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t30 two_stage_opamp_dummy_magic_23_0.V_p_mir.t1 GNDA.t102 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X1006 a_13570_4368.t0 two_stage_opamp_dummy_magic_23_0.V_tot.t0 GNDA.t48 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X1007 VOUT+.t150 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1008 two_stage_opamp_dummy_magic_23_0.Vb2.t5 bgr_11_0.NFET_GATE_10uA.t22 GNDA.t127 GNDA.t126 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1009 two_stage_opamp_dummy_magic_23_0.VD1.t12 two_stage_opamp_dummy_magic_23_0.Vb1.t34 two_stage_opamp_dummy_magic_23_0.X.t21 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1010 GNDA.t123 bgr_11_0.NFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_23_0.Vb2.t4 GNDA.t122 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1011 VDDA.t433 bgr_11_0.V_mir1.t21 bgr_11_0.1st_Vout_1.t9 VDDA.t432 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X1012 GNDA.t586 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t31 two_stage_opamp_dummy_magic_23_0.V_source.t8 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X1013 VDDA.t724 GNDA.t216 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1014 VOUT-.t151 two_stage_opamp_dummy_magic_23_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1015 VDDA.t725 GNDA.t215 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1016 GNDA.t489 GNDA.t487 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t14 GNDA.t488 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X1017 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t7 two_stage_opamp_dummy_magic_23_0.X.t54 GNDA.t137 VDDA.t158 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X1018 VDDA.t726 GNDA.t214 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1019 VOUT+.t151 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1020 VDDA.t727 GNDA.t213 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1021 bgr_11_0.1st_Vout_2.t34 bgr_11_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1022 VDDA.t728 GNDA.t212 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1023 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t1 VDDA.t312 VDDA.t314 VDDA.t313 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X1024 two_stage_opamp_dummy_magic_23_0.V_source.t2 two_stage_opamp_dummy_magic_23_0.err_amp_out.t12 GNDA.t41 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X1025 two_stage_opamp_dummy_magic_23_0.VD4.t0 two_stage_opamp_dummy_magic_23_0.Vb3.t28 VDDA.t123 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X1026 VDDA.t269 two_stage_opamp_dummy_magic_23_0.Y.t54 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t4 GNDA.t183 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X1027 two_stage_opamp_dummy_magic_23_0.V_source.t32 VIN-.t8 two_stage_opamp_dummy_magic_23_0.VD1.t7 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1028 VOUT-.t152 two_stage_opamp_dummy_magic_23_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1029 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t2 two_stage_opamp_dummy_magic_23_0.V_tot.t12 two_stage_opamp_dummy_magic_23_0.V_err_p.t2 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X1030 VOUT-.t153 two_stage_opamp_dummy_magic_23_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1031 VDDA.t729 GNDA.t211 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1032 two_stage_opamp_dummy_magic_23_0.VD4.t12 two_stage_opamp_dummy_magic_23_0.VD4.t10 two_stage_opamp_dummy_magic_23_0.Y.t3 two_stage_opamp_dummy_magic_23_0.VD4.t11 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X1033 bgr_11_0.1st_Vout_2.t35 bgr_11_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1034 VOUT-.t154 two_stage_opamp_dummy_magic_23_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1035 VDDA.t730 GNDA.t210 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1036 bgr_11_0.START_UP.t2 bgr_11_0.V_TOP.t48 VDDA.t137 VDDA.t136 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X1037 GNDA.t480 GNDA.t478 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t14 GNDA.t479 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X1038 bgr_11_0.1st_Vout_2.t2 bgr_11_0.V_mir2.t22 VDDA.t52 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X1039 VDDA.t106 bgr_11_0.1st_Vout_1.t35 bgr_11_0.V_TOP.t8 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X1040 VOUT+.t152 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1041 VOUT+.t153 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1042 VOUT+.t154 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1043 VDDA.t194 two_stage_opamp_dummy_magic_23_0.V_err_gate.t33 two_stage_opamp_dummy_magic_23_0.V_err_p.t3 VDDA.t193 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X1044 VOUT+.t155 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1045 two_stage_opamp_dummy_magic_23_0.V_err_gate.t10 VDDA.t309 VDDA.t311 VDDA.t310 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X1046 two_stage_opamp_dummy_magic_23_0.V_source.t1 VIN+.t10 two_stage_opamp_dummy_magic_23_0.VD2.t0 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1047 VDDA.t731 GNDA.t209 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1048 VDDA.t732 GNDA.t208 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1049 GNDA.t207 VDDA.t733 bgr_11_0.V_p_2.t9 GNDA.t206 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X1050 bgr_11_0.V_p_1.t0 bgr_11_0.Vin+.t10 bgr_11_0.1st_Vout_1.t10 GNDA.t590 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X1051 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t0 VIN-.t9 two_stage_opamp_dummy_magic_23_0.V_p_mir.t0 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1052 two_stage_opamp_dummy_magic_23_0.V_source.t28 VIN-.t10 two_stage_opamp_dummy_magic_23_0.VD1.t5 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X1053 bgr_11_0.1st_Vout_1.t36 bgr_11_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1054 VDDA.t734 GNDA.t205 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1055 VDDA.t735 GNDA.t204 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1056 VDDA.t21 bgr_11_0.V_mir1.t22 bgr_11_0.1st_Vout_1.t0 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X1057 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t1 two_stage_opamp_dummy_magic_23_0.V_tot.t13 two_stage_opamp_dummy_magic_23_0.V_err_p.t1 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X1058 VOUT-.t155 two_stage_opamp_dummy_magic_23_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1059 VDDA.t736 GNDA.t203 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1060 VOUT+.t156 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1061 bgr_11_0.1st_Vout_2.t36 bgr_11_0.cap_res2.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1062 bgr_11_0.Vin+.t2 bgr_11_0.V_TOP.t49 VDDA.t139 VDDA.t138 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X1063 VOUT-.t156 two_stage_opamp_dummy_magic_23_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 two_stage_opamp_dummy_magic_23_0.Y.n65 two_stage_opamp_dummy_magic_23_0.Y.t28 1172.87
R1 two_stage_opamp_dummy_magic_23_0.Y.n63 two_stage_opamp_dummy_magic_23_0.Y.t50 1172.87
R2 two_stage_opamp_dummy_magic_23_0.Y.n65 two_stage_opamp_dummy_magic_23_0.Y.t44 996.134
R3 two_stage_opamp_dummy_magic_23_0.Y.n66 two_stage_opamp_dummy_magic_23_0.Y.t30 996.134
R4 two_stage_opamp_dummy_magic_23_0.Y.n67 two_stage_opamp_dummy_magic_23_0.Y.t38 996.134
R5 two_stage_opamp_dummy_magic_23_0.Y.n68 two_stage_opamp_dummy_magic_23_0.Y.t53 996.134
R6 two_stage_opamp_dummy_magic_23_0.Y.n69 two_stage_opamp_dummy_magic_23_0.Y.t40 996.134
R7 two_stage_opamp_dummy_magic_23_0.Y.n70 two_stage_opamp_dummy_magic_23_0.Y.t25 996.134
R8 two_stage_opamp_dummy_magic_23_0.Y.n64 two_stage_opamp_dummy_magic_23_0.Y.t42 996.134
R9 two_stage_opamp_dummy_magic_23_0.Y.n63 two_stage_opamp_dummy_magic_23_0.Y.t35 996.134
R10 two_stage_opamp_dummy_magic_23_0.Y.n58 two_stage_opamp_dummy_magic_23_0.Y.t54 690.867
R11 two_stage_opamp_dummy_magic_23_0.Y.n51 two_stage_opamp_dummy_magic_23_0.Y.t47 690.867
R12 two_stage_opamp_dummy_magic_23_0.Y.n49 two_stage_opamp_dummy_magic_23_0.Y.t49 530.201
R13 two_stage_opamp_dummy_magic_23_0.Y.n42 two_stage_opamp_dummy_magic_23_0.Y.t43 530.201
R14 two_stage_opamp_dummy_magic_23_0.Y.n58 two_stage_opamp_dummy_magic_23_0.Y.t41 514.134
R15 two_stage_opamp_dummy_magic_23_0.Y.n51 two_stage_opamp_dummy_magic_23_0.Y.t32 514.134
R16 two_stage_opamp_dummy_magic_23_0.Y.n52 two_stage_opamp_dummy_magic_23_0.Y.t39 514.134
R17 two_stage_opamp_dummy_magic_23_0.Y.n53 two_stage_opamp_dummy_magic_23_0.Y.t51 514.134
R18 two_stage_opamp_dummy_magic_23_0.Y.n54 two_stage_opamp_dummy_magic_23_0.Y.t36 514.134
R19 two_stage_opamp_dummy_magic_23_0.Y.n55 two_stage_opamp_dummy_magic_23_0.Y.t48 514.134
R20 two_stage_opamp_dummy_magic_23_0.Y.n56 two_stage_opamp_dummy_magic_23_0.Y.t33 514.134
R21 two_stage_opamp_dummy_magic_23_0.Y.n57 two_stage_opamp_dummy_magic_23_0.Y.t26 514.134
R22 two_stage_opamp_dummy_magic_23_0.Y.n49 two_stage_opamp_dummy_magic_23_0.Y.t37 353.467
R23 two_stage_opamp_dummy_magic_23_0.Y.n48 two_stage_opamp_dummy_magic_23_0.Y.t52 353.467
R24 two_stage_opamp_dummy_magic_23_0.Y.n47 two_stage_opamp_dummy_magic_23_0.Y.t29 353.467
R25 two_stage_opamp_dummy_magic_23_0.Y.n46 two_stage_opamp_dummy_magic_23_0.Y.t45 353.467
R26 two_stage_opamp_dummy_magic_23_0.Y.n45 two_stage_opamp_dummy_magic_23_0.Y.t31 353.467
R27 two_stage_opamp_dummy_magic_23_0.Y.n44 two_stage_opamp_dummy_magic_23_0.Y.t46 353.467
R28 two_stage_opamp_dummy_magic_23_0.Y.n43 two_stage_opamp_dummy_magic_23_0.Y.t34 353.467
R29 two_stage_opamp_dummy_magic_23_0.Y.n42 two_stage_opamp_dummy_magic_23_0.Y.t27 353.467
R30 two_stage_opamp_dummy_magic_23_0.Y.n72 two_stage_opamp_dummy_magic_23_0.Y.n71 304.375
R31 two_stage_opamp_dummy_magic_23_0.Y.n60 two_stage_opamp_dummy_magic_23_0.Y.n50 216.9
R32 two_stage_opamp_dummy_magic_23_0.Y.n60 two_stage_opamp_dummy_magic_23_0.Y.n59 216.9
R33 two_stage_opamp_dummy_magic_23_0.Y.n64 two_stage_opamp_dummy_magic_23_0.Y.n63 176.733
R34 two_stage_opamp_dummy_magic_23_0.Y.n66 two_stage_opamp_dummy_magic_23_0.Y.n65 176.733
R35 two_stage_opamp_dummy_magic_23_0.Y.n67 two_stage_opamp_dummy_magic_23_0.Y.n66 176.733
R36 two_stage_opamp_dummy_magic_23_0.Y.n68 two_stage_opamp_dummy_magic_23_0.Y.n67 176.733
R37 two_stage_opamp_dummy_magic_23_0.Y.n69 two_stage_opamp_dummy_magic_23_0.Y.n68 176.733
R38 two_stage_opamp_dummy_magic_23_0.Y.n70 two_stage_opamp_dummy_magic_23_0.Y.n69 176.733
R39 two_stage_opamp_dummy_magic_23_0.Y.n48 two_stage_opamp_dummy_magic_23_0.Y.n47 176.733
R40 two_stage_opamp_dummy_magic_23_0.Y.n47 two_stage_opamp_dummy_magic_23_0.Y.n46 176.733
R41 two_stage_opamp_dummy_magic_23_0.Y.n46 two_stage_opamp_dummy_magic_23_0.Y.n45 176.733
R42 two_stage_opamp_dummy_magic_23_0.Y.n45 two_stage_opamp_dummy_magic_23_0.Y.n44 176.733
R43 two_stage_opamp_dummy_magic_23_0.Y.n44 two_stage_opamp_dummy_magic_23_0.Y.n43 176.733
R44 two_stage_opamp_dummy_magic_23_0.Y.n43 two_stage_opamp_dummy_magic_23_0.Y.n42 176.733
R45 two_stage_opamp_dummy_magic_23_0.Y.n57 two_stage_opamp_dummy_magic_23_0.Y.n56 176.733
R46 two_stage_opamp_dummy_magic_23_0.Y.n56 two_stage_opamp_dummy_magic_23_0.Y.n55 176.733
R47 two_stage_opamp_dummy_magic_23_0.Y.n55 two_stage_opamp_dummy_magic_23_0.Y.n54 176.733
R48 two_stage_opamp_dummy_magic_23_0.Y.n54 two_stage_opamp_dummy_magic_23_0.Y.n53 176.733
R49 two_stage_opamp_dummy_magic_23_0.Y.n53 two_stage_opamp_dummy_magic_23_0.Y.n52 176.733
R50 two_stage_opamp_dummy_magic_23_0.Y.n52 two_stage_opamp_dummy_magic_23_0.Y.n51 176.733
R51 two_stage_opamp_dummy_magic_23_0.Y.n61 two_stage_opamp_dummy_magic_23_0.Y.n60 175.05
R52 two_stage_opamp_dummy_magic_23_0.Y.n22 two_stage_opamp_dummy_magic_23_0.Y.n21 66.0338
R53 two_stage_opamp_dummy_magic_23_0.Y.n26 two_stage_opamp_dummy_magic_23_0.Y.n25 66.0338
R54 two_stage_opamp_dummy_magic_23_0.Y.n28 two_stage_opamp_dummy_magic_23_0.Y.n27 66.0338
R55 two_stage_opamp_dummy_magic_23_0.Y.n32 two_stage_opamp_dummy_magic_23_0.Y.n31 66.0338
R56 two_stage_opamp_dummy_magic_23_0.Y.n35 two_stage_opamp_dummy_magic_23_0.Y.n34 66.0338
R57 two_stage_opamp_dummy_magic_23_0.Y.n39 two_stage_opamp_dummy_magic_23_0.Y.n38 66.0338
R58 two_stage_opamp_dummy_magic_23_0.Y.t16 two_stage_opamp_dummy_magic_23_0.Y.n72 49.4802
R59 two_stage_opamp_dummy_magic_23_0.Y.n1 two_stage_opamp_dummy_magic_23_0.Y.n0 49.3505
R60 two_stage_opamp_dummy_magic_23_0.Y.n6 two_stage_opamp_dummy_magic_23_0.Y.n5 49.3505
R61 two_stage_opamp_dummy_magic_23_0.Y.n9 two_stage_opamp_dummy_magic_23_0.Y.n8 49.3505
R62 two_stage_opamp_dummy_magic_23_0.Y.n12 two_stage_opamp_dummy_magic_23_0.Y.n11 49.3505
R63 two_stage_opamp_dummy_magic_23_0.Y.n4 two_stage_opamp_dummy_magic_23_0.Y.n3 49.3505
R64 two_stage_opamp_dummy_magic_23_0.Y.n17 two_stage_opamp_dummy_magic_23_0.Y.n16 49.3505
R65 two_stage_opamp_dummy_magic_23_0.Y.n71 two_stage_opamp_dummy_magic_23_0.Y.n64 40.1672
R66 two_stage_opamp_dummy_magic_23_0.Y.n71 two_stage_opamp_dummy_magic_23_0.Y.n70 40.1672
R67 two_stage_opamp_dummy_magic_23_0.Y.n50 two_stage_opamp_dummy_magic_23_0.Y.n48 40.1672
R68 two_stage_opamp_dummy_magic_23_0.Y.n50 two_stage_opamp_dummy_magic_23_0.Y.n49 40.1672
R69 two_stage_opamp_dummy_magic_23_0.Y.n59 two_stage_opamp_dummy_magic_23_0.Y.n57 40.1672
R70 two_stage_opamp_dummy_magic_23_0.Y.n59 two_stage_opamp_dummy_magic_23_0.Y.n58 40.1672
R71 two_stage_opamp_dummy_magic_23_0.Y.n61 two_stage_opamp_dummy_magic_23_0.Y.n41 17.6567
R72 two_stage_opamp_dummy_magic_23_0.Y.n0 two_stage_opamp_dummy_magic_23_0.Y.t11 16.0005
R73 two_stage_opamp_dummy_magic_23_0.Y.n0 two_stage_opamp_dummy_magic_23_0.Y.t5 16.0005
R74 two_stage_opamp_dummy_magic_23_0.Y.n5 two_stage_opamp_dummy_magic_23_0.Y.t24 16.0005
R75 two_stage_opamp_dummy_magic_23_0.Y.n5 two_stage_opamp_dummy_magic_23_0.Y.t19 16.0005
R76 two_stage_opamp_dummy_magic_23_0.Y.n8 two_stage_opamp_dummy_magic_23_0.Y.t10 16.0005
R77 two_stage_opamp_dummy_magic_23_0.Y.n8 two_stage_opamp_dummy_magic_23_0.Y.t8 16.0005
R78 two_stage_opamp_dummy_magic_23_0.Y.n11 two_stage_opamp_dummy_magic_23_0.Y.t9 16.0005
R79 two_stage_opamp_dummy_magic_23_0.Y.n11 two_stage_opamp_dummy_magic_23_0.Y.t7 16.0005
R80 two_stage_opamp_dummy_magic_23_0.Y.n3 two_stage_opamp_dummy_magic_23_0.Y.t4 16.0005
R81 two_stage_opamp_dummy_magic_23_0.Y.n3 two_stage_opamp_dummy_magic_23_0.Y.t15 16.0005
R82 two_stage_opamp_dummy_magic_23_0.Y.n16 two_stage_opamp_dummy_magic_23_0.Y.t12 16.0005
R83 two_stage_opamp_dummy_magic_23_0.Y.n16 two_stage_opamp_dummy_magic_23_0.Y.t6 16.0005
R84 two_stage_opamp_dummy_magic_23_0.Y.n21 two_stage_opamp_dummy_magic_23_0.Y.t1 11.2576
R85 two_stage_opamp_dummy_magic_23_0.Y.n21 two_stage_opamp_dummy_magic_23_0.Y.t17 11.2576
R86 two_stage_opamp_dummy_magic_23_0.Y.n25 two_stage_opamp_dummy_magic_23_0.Y.t3 11.2576
R87 two_stage_opamp_dummy_magic_23_0.Y.n25 two_stage_opamp_dummy_magic_23_0.Y.t0 11.2576
R88 two_stage_opamp_dummy_magic_23_0.Y.n27 two_stage_opamp_dummy_magic_23_0.Y.t13 11.2576
R89 two_stage_opamp_dummy_magic_23_0.Y.n27 two_stage_opamp_dummy_magic_23_0.Y.t20 11.2576
R90 two_stage_opamp_dummy_magic_23_0.Y.n31 two_stage_opamp_dummy_magic_23_0.Y.t22 11.2576
R91 two_stage_opamp_dummy_magic_23_0.Y.n31 two_stage_opamp_dummy_magic_23_0.Y.t23 11.2576
R92 two_stage_opamp_dummy_magic_23_0.Y.n34 two_stage_opamp_dummy_magic_23_0.Y.t21 11.2576
R93 two_stage_opamp_dummy_magic_23_0.Y.n34 two_stage_opamp_dummy_magic_23_0.Y.t14 11.2576
R94 two_stage_opamp_dummy_magic_23_0.Y.n38 two_stage_opamp_dummy_magic_23_0.Y.t2 11.2576
R95 two_stage_opamp_dummy_magic_23_0.Y.n38 two_stage_opamp_dummy_magic_23_0.Y.t18 11.2576
R96 two_stage_opamp_dummy_magic_23_0.Y.n62 two_stage_opamp_dummy_magic_23_0.Y.n20 10.2817
R97 two_stage_opamp_dummy_magic_23_0.Y.n29 two_stage_opamp_dummy_magic_23_0.Y.n26 5.91717
R98 two_stage_opamp_dummy_magic_23_0.Y.n26 two_stage_opamp_dummy_magic_23_0.Y.n24 5.91717
R99 two_stage_opamp_dummy_magic_23_0.Y.n37 two_stage_opamp_dummy_magic_23_0.Y.n22 5.91717
R100 two_stage_opamp_dummy_magic_23_0.Y.n15 two_stage_opamp_dummy_magic_23_0.Y.n4 5.6255
R101 two_stage_opamp_dummy_magic_23_0.Y.n10 two_stage_opamp_dummy_magic_23_0.Y.n6 5.6255
R102 two_stage_opamp_dummy_magic_23_0.Y.n18 two_stage_opamp_dummy_magic_23_0.Y.n4 5.438
R103 two_stage_opamp_dummy_magic_23_0.Y.n7 two_stage_opamp_dummy_magic_23_0.Y.n6 5.438
R104 two_stage_opamp_dummy_magic_23_0.Y.n28 two_stage_opamp_dummy_magic_23_0.Y.n24 5.29217
R105 two_stage_opamp_dummy_magic_23_0.Y.n29 two_stage_opamp_dummy_magic_23_0.Y.n28 5.29217
R106 two_stage_opamp_dummy_magic_23_0.Y.n33 two_stage_opamp_dummy_magic_23_0.Y.n32 5.29217
R107 two_stage_opamp_dummy_magic_23_0.Y.n32 two_stage_opamp_dummy_magic_23_0.Y.n30 5.29217
R108 two_stage_opamp_dummy_magic_23_0.Y.n36 two_stage_opamp_dummy_magic_23_0.Y.n35 5.29217
R109 two_stage_opamp_dummy_magic_23_0.Y.n35 two_stage_opamp_dummy_magic_23_0.Y.n23 5.29217
R110 two_stage_opamp_dummy_magic_23_0.Y.n39 two_stage_opamp_dummy_magic_23_0.Y.n37 5.29217
R111 two_stage_opamp_dummy_magic_23_0.Y.n40 two_stage_opamp_dummy_magic_23_0.Y.n39 5.29217
R112 two_stage_opamp_dummy_magic_23_0.Y.n41 two_stage_opamp_dummy_magic_23_0.Y.n40 5.1255
R113 two_stage_opamp_dummy_magic_23_0.Y.n10 two_stage_opamp_dummy_magic_23_0.Y.n9 5.063
R114 two_stage_opamp_dummy_magic_23_0.Y.n13 two_stage_opamp_dummy_magic_23_0.Y.n12 5.063
R115 two_stage_opamp_dummy_magic_23_0.Y.n17 two_stage_opamp_dummy_magic_23_0.Y.n15 5.063
R116 two_stage_opamp_dummy_magic_23_0.Y.n14 two_stage_opamp_dummy_magic_23_0.Y.n1 5.063
R117 two_stage_opamp_dummy_magic_23_0.Y.n9 two_stage_opamp_dummy_magic_23_0.Y.n7 4.8755
R118 two_stage_opamp_dummy_magic_23_0.Y.n12 two_stage_opamp_dummy_magic_23_0.Y.n2 4.8755
R119 two_stage_opamp_dummy_magic_23_0.Y.n18 two_stage_opamp_dummy_magic_23_0.Y.n17 4.8755
R120 two_stage_opamp_dummy_magic_23_0.Y.n20 two_stage_opamp_dummy_magic_23_0.Y.n19 4.5005
R121 two_stage_opamp_dummy_magic_23_0.Y.n62 two_stage_opamp_dummy_magic_23_0.Y.n61 4.5005
R122 two_stage_opamp_dummy_magic_23_0.Y.n72 two_stage_opamp_dummy_magic_23_0.Y.n62 3.27133
R123 two_stage_opamp_dummy_magic_23_0.Y.n41 two_stage_opamp_dummy_magic_23_0.Y.n22 0.792167
R124 two_stage_opamp_dummy_magic_23_0.Y.n40 two_stage_opamp_dummy_magic_23_0.Y.n23 0.6255
R125 two_stage_opamp_dummy_magic_23_0.Y.n30 two_stage_opamp_dummy_magic_23_0.Y.n23 0.6255
R126 two_stage_opamp_dummy_magic_23_0.Y.n30 two_stage_opamp_dummy_magic_23_0.Y.n29 0.6255
R127 two_stage_opamp_dummy_magic_23_0.Y.n33 two_stage_opamp_dummy_magic_23_0.Y.n24 0.6255
R128 two_stage_opamp_dummy_magic_23_0.Y.n36 two_stage_opamp_dummy_magic_23_0.Y.n33 0.6255
R129 two_stage_opamp_dummy_magic_23_0.Y.n37 two_stage_opamp_dummy_magic_23_0.Y.n36 0.6255
R130 two_stage_opamp_dummy_magic_23_0.Y.n15 two_stage_opamp_dummy_magic_23_0.Y.n14 0.563
R131 two_stage_opamp_dummy_magic_23_0.Y.n19 two_stage_opamp_dummy_magic_23_0.Y.n18 0.563
R132 two_stage_opamp_dummy_magic_23_0.Y.n19 two_stage_opamp_dummy_magic_23_0.Y.n2 0.563
R133 two_stage_opamp_dummy_magic_23_0.Y.n7 two_stage_opamp_dummy_magic_23_0.Y.n2 0.563
R134 two_stage_opamp_dummy_magic_23_0.Y.n13 two_stage_opamp_dummy_magic_23_0.Y.n10 0.563
R135 two_stage_opamp_dummy_magic_23_0.Y.n14 two_stage_opamp_dummy_magic_23_0.Y.n13 0.563
R136 two_stage_opamp_dummy_magic_23_0.Y.n20 two_stage_opamp_dummy_magic_23_0.Y.n1 0.3755
R137 VDDA.n500 VDDA.t370 1231.74
R138 VDDA.n503 VDDA.t358 1231.74
R139 VDDA.n419 VDDA.t409 1231.74
R140 VDDA.n422 VDDA.t421 1231.74
R141 VDDA.t413 VDDA.n485 1095.3
R142 VDDA.n486 VDDA.t310 1095.3
R143 VDDA.n446 VDDA.t362 1095.3
R144 VDDA.t356 VDDA.n445 1095.3
R145 VDDA.n405 VDDA.t416 1095.3
R146 VDDA.t407 VDDA.n404 1095.3
R147 VDDA.n557 VDDA.t316 676.966
R148 VDDA.n457 VDDA.t397 672.293
R149 VDDA.n460 VDDA.t352 672.293
R150 VDDA.n376 VDDA.t324 672.293
R151 VDDA.n379 VDDA.t394 672.293
R152 VDDA.n485 VDDA.t414 663.801
R153 VDDA.n486 VDDA.t311 663.801
R154 VDDA.n446 VDDA.t363 663.801
R155 VDDA.n445 VDDA.t357 663.801
R156 VDDA.n405 VDDA.t417 663.801
R157 VDDA.n404 VDDA.t408 663.801
R158 VDDA.n518 VDDA.t339 661.375
R159 VDDA.n521 VDDA.t376 661.375
R160 VDDA.t380 VDDA.n302 660.001
R161 VDDA.t328 VDDA.n350 645.231
R162 VDDA.n351 VDDA.t392 645.231
R163 VDDA.t386 VDDA.n556 643.038
R164 VDDA.t368 VDDA.n536 643.038
R165 VDDA.n537 VDDA.t365 643.038
R166 VDDA.n334 VDDA.t343 643.037
R167 VDDA.t419 VDDA.n333 643.037
R168 VDDA.t401 VDDA.n342 643.037
R169 VDDA.n343 VDDA.t322 643.037
R170 VDDA.n425 VDDA.n424 599.342
R171 VDDA.n427 VDDA.n426 599.342
R172 VDDA.n429 VDDA.n428 599.342
R173 VDDA.n431 VDDA.n430 599.342
R174 VDDA.n433 VDDA.n432 599.342
R175 VDDA.n435 VDDA.n434 599.342
R176 VDDA.n437 VDDA.n436 599.342
R177 VDDA.n439 VDDA.n438 599.342
R178 VDDA.n441 VDDA.n440 599.342
R179 VDDA.n443 VDDA.n442 599.342
R180 VDDA.n478 VDDA.t403 589.076
R181 VDDA.n481 VDDA.t382 589.076
R182 VDDA.n397 VDDA.t318 589.076
R183 VDDA.n400 VDDA.t336 589.076
R184 VDDA.n582 VDDA.n550 587.407
R185 VDDA.n578 VDDA.n577 587.407
R186 VDDA.n595 VDDA.n594 587.407
R187 VDDA.n589 VDDA.n544 587.407
R188 VDDA.n594 VDDA.n593 585
R189 VDDA.n592 VDDA.n589 585
R190 VDDA.n580 VDDA.n550 585
R191 VDDA.n579 VDDA.n578 585
R192 VDDA.t468 VDDA.t413 580.557
R193 VDDA.t74 VDDA.t468 580.557
R194 VDDA.t442 VDDA.t74 580.557
R195 VDDA.t140 VDDA.t442 580.557
R196 VDDA.t240 VDDA.t140 580.557
R197 VDDA.t69 VDDA.t240 580.557
R198 VDDA.t17 VDDA.t69 580.557
R199 VDDA.t4 VDDA.t17 580.557
R200 VDDA.t248 VDDA.t4 580.557
R201 VDDA.t111 VDDA.t248 580.557
R202 VDDA.t310 VDDA.t111 580.557
R203 VDDA.t362 VDDA.t75 580.557
R204 VDDA.t75 VDDA.t251 580.557
R205 VDDA.t251 VDDA.t182 580.557
R206 VDDA.t182 VDDA.t195 580.557
R207 VDDA.t195 VDDA.t166 580.557
R208 VDDA.t166 VDDA.t191 580.557
R209 VDDA.t191 VDDA.t168 580.557
R210 VDDA.t168 VDDA.t193 580.557
R211 VDDA.t193 VDDA.t253 580.557
R212 VDDA.t253 VDDA.t213 580.557
R213 VDDA.t213 VDDA.t205 580.557
R214 VDDA.t205 VDDA.t201 580.557
R215 VDDA.t201 VDDA.t263 580.557
R216 VDDA.t263 VDDA.t77 580.557
R217 VDDA.t77 VDDA.t265 580.557
R218 VDDA.t265 VDDA.t203 580.557
R219 VDDA.t203 VDDA.t199 580.557
R220 VDDA.t199 VDDA.t184 580.557
R221 VDDA.t184 VDDA.t197 580.557
R222 VDDA.t197 VDDA.t211 580.557
R223 VDDA.t211 VDDA.t356 580.557
R224 VDDA.t416 VDDA.t104 580.557
R225 VDDA.t104 VDDA.t18 580.557
R226 VDDA.t18 VDDA.t24 580.557
R227 VDDA.t24 VDDA.t91 580.557
R228 VDDA.t91 VDDA.t92 580.557
R229 VDDA.t92 VDDA.t431 580.557
R230 VDDA.t431 VDDA.t19 580.557
R231 VDDA.t19 VDDA.t455 580.557
R232 VDDA.t455 VDDA.t43 580.557
R233 VDDA.t43 VDDA.t426 580.557
R234 VDDA.t426 VDDA.t407 580.557
R235 VDDA.n303 VDDA.t334 540.818
R236 VDDA.n296 VDDA.t389 540.818
R237 VDDA.t374 VDDA.n295 540.818
R238 VDDA.n510 VDDA.t345 456.526
R239 VDDA.n513 VDDA.t330 456.526
R240 VDDA.n535 VDDA.t367 419.108
R241 VDDA.n538 VDDA.t364 419.108
R242 VDDA.n555 VDDA.t385 413.084
R243 VDDA.n558 VDDA.t315 413.084
R244 VDDA.n349 VDDA.t327 409.067
R245 VDDA.n352 VDDA.t391 409.067
R246 VDDA.n332 VDDA.t418 409.067
R247 VDDA.n335 VDDA.t342 409.067
R248 VDDA.n341 VDDA.t400 409.067
R249 VDDA.t334 VDDA.t30 407.144
R250 VDDA.t30 VDDA.t424 407.144
R251 VDDA.t424 VDDA.t245 407.144
R252 VDDA.t245 VDDA.t249 407.144
R253 VDDA.t249 VDDA.t38 407.144
R254 VDDA.t38 VDDA.t105 407.144
R255 VDDA.t105 VDDA.t61 407.144
R256 VDDA.t61 VDDA.t267 407.144
R257 VDDA.t267 VDDA.t112 407.144
R258 VDDA.t112 VDDA.t432 407.144
R259 VDDA.t432 VDDA.t243 407.144
R260 VDDA.t243 VDDA.t114 407.144
R261 VDDA.t114 VDDA.t5 407.144
R262 VDDA.t5 VDDA.t235 407.144
R263 VDDA.t235 VDDA.t25 407.144
R264 VDDA.t25 VDDA.t20 407.144
R265 VDDA.t20 VDDA.t134 407.144
R266 VDDA.t134 VDDA.t107 407.144
R267 VDDA.t107 VDDA.t380 407.144
R268 VDDA.t389 VDDA.t79 407.144
R269 VDDA.t79 VDDA.t443 407.144
R270 VDDA.t443 VDDA.t51 407.144
R271 VDDA.t51 VDDA.t227 407.144
R272 VDDA.t227 VDDA.t116 407.144
R273 VDDA.t116 VDDA.t63 407.144
R274 VDDA.t63 VDDA.t70 407.144
R275 VDDA.t70 VDDA.t7 407.144
R276 VDDA.t7 VDDA.t460 407.144
R277 VDDA.t460 VDDA.t0 407.144
R278 VDDA.t0 VDDA.t83 407.144
R279 VDDA.t83 VDDA.t41 407.144
R280 VDDA.t41 VDDA.t65 407.144
R281 VDDA.t65 VDDA.t438 407.144
R282 VDDA.t438 VDDA.t219 407.144
R283 VDDA.t219 VDDA.t98 407.144
R284 VDDA.t98 VDDA.t126 407.144
R285 VDDA.t126 VDDA.t81 407.144
R286 VDDA.t81 VDDA.t374 407.144
R287 VDDA.n512 VDDA.t331 397.784
R288 VDDA.t346 VDDA.n511 397.784
R289 VDDA.n344 VDDA.t321 390.322
R290 VDDA.t333 VDDA.n304 379.582
R291 VDDA.t388 VDDA.n297 379.582
R292 VDDA.n294 VDDA.t373 379.277
R293 VDDA.t247 VDDA.t386 373.214
R294 VDDA.t157 VDDA.t247 373.214
R295 VDDA.t316 VDDA.t157 373.214
R296 VDDA.t9 VDDA.t368 373.214
R297 VDDA.t151 VDDA.t9 373.214
R298 VDDA.t365 VDDA.t151 373.214
R299 VDDA.t343 VDDA.t449 373.214
R300 VDDA.t449 VDDA.t456 373.214
R301 VDDA.t456 VDDA.t225 373.214
R302 VDDA.t225 VDDA.t118 373.214
R303 VDDA.t118 VDDA.t419 373.214
R304 VDDA.t464 VDDA.t328 373.214
R305 VDDA.t100 VDDA.t464 373.214
R306 VDDA.t149 VDDA.t100 373.214
R307 VDDA.t120 VDDA.t149 373.214
R308 VDDA.t436 VDDA.t120 373.214
R309 VDDA.t462 VDDA.t436 373.214
R310 VDDA.t447 VDDA.t462 373.214
R311 VDDA.t109 VDDA.t447 373.214
R312 VDDA.t128 VDDA.t109 373.214
R313 VDDA.t445 VDDA.t128 373.214
R314 VDDA.t392 VDDA.t445 373.214
R315 VDDA.t11 VDDA.t401 373.214
R316 VDDA.t147 VDDA.t11 373.214
R317 VDDA.t47 VDDA.t147 373.214
R318 VDDA.t45 VDDA.t47 373.214
R319 VDDA.t322 VDDA.t45 373.214
R320 VDDA.n575 VDDA.t349 360.868
R321 VDDA.n600 VDDA.t312 360.868
R322 VDDA.n301 VDDA.t379 358.858
R323 VDDA.n305 VDDA.t333 358.858
R324 VDDA.n298 VDDA.t388 358.858
R325 VDDA.t373 VDDA.n292 358.858
R326 VDDA.n350 VDDA.t329 354.154
R327 VDDA.n351 VDDA.t393 354.154
R328 VDDA.n537 VDDA.t366 354.065
R329 VDDA.n302 VDDA.t381 354.065
R330 VDDA.n556 VDDA.t387 354.063
R331 VDDA.n536 VDDA.t369 354.063
R332 VDDA.n254 VDDA.t335 351.793
R333 VDDA.n274 VDDA.t390 351.793
R334 VDDA.n293 VDDA.t375 351.793
R335 VDDA.n444 VDDA.t355 348.325
R336 VDDA.n447 VDDA.t361 348.325
R337 VDDA.n484 VDDA.t412 348.075
R338 VDDA.n487 VDDA.t309 348.075
R339 VDDA.n403 VDDA.t406 348.075
R340 VDDA.n406 VDDA.t415 348.075
R341 VDDA.n557 VDDA.t317 347.224
R342 VDDA.n338 VDDA.n337 345.127
R343 VDDA.n340 VDDA.n339 345.127
R344 VDDA.n329 VDDA.n328 344.7
R345 VDDA.n331 VDDA.n330 344.7
R346 VDDA.n480 VDDA.t383 343.882
R347 VDDA.t404 VDDA.n479 343.882
R348 VDDA.t319 VDDA.n398 343.882
R349 VDDA.n399 VDDA.t337 343.882
R350 VDDA.n252 VDDA.n251 341.675
R351 VDDA.n256 VDDA.n255 341.675
R352 VDDA.n258 VDDA.n257 341.675
R353 VDDA.n260 VDDA.n259 341.675
R354 VDDA.n262 VDDA.n261 341.675
R355 VDDA.n264 VDDA.n263 341.675
R356 VDDA.n266 VDDA.n265 341.675
R357 VDDA.n268 VDDA.n267 341.675
R358 VDDA.n270 VDDA.n269 341.675
R359 VDDA.n272 VDDA.n271 341.675
R360 VDDA.n277 VDDA.n276 341.675
R361 VDDA.n279 VDDA.n278 341.675
R362 VDDA.n281 VDDA.n280 341.675
R363 VDDA.n283 VDDA.n282 341.675
R364 VDDA.n285 VDDA.n284 341.675
R365 VDDA.n287 VDDA.n286 341.675
R366 VDDA.n289 VDDA.n288 341.675
R367 VDDA.n291 VDDA.n290 341.675
R368 VDDA.n327 VDDA.n326 339.272
R369 VDDA.n347 VDDA.n346 339.272
R370 VDDA.n355 VDDA.n354 339.272
R371 VDDA.n357 VDDA.n356 339.272
R372 VDDA.n541 VDDA.n540 334.772
R373 VDDA.n360 VDDA.n359 334.772
R374 VDDA.n342 VDDA.t402 332.267
R375 VDDA.n343 VDDA.t323 332.267
R376 VDDA.n334 VDDA.t344 332.084
R377 VDDA.n333 VDDA.t420 332.084
R378 VDDA.t331 VDDA.t2 259.091
R379 VDDA.t2 VDDA.t346 259.091
R380 VDDA.t27 VDDA.t350 251.471
R381 VDDA.t59 VDDA.t27 251.471
R382 VDDA.t136 VDDA.t59 251.471
R383 VDDA.t221 VDDA.t136 251.471
R384 VDDA.t93 VDDA.t221 251.471
R385 VDDA.t216 VDDA.t93 251.471
R386 VDDA.t142 VDDA.t216 251.471
R387 VDDA.t238 VDDA.t142 251.471
R388 VDDA.t233 VDDA.t238 251.471
R389 VDDA.t34 VDDA.t233 251.471
R390 VDDA.t138 VDDA.t34 251.471
R391 VDDA.t144 VDDA.t138 251.471
R392 VDDA.t223 VDDA.t144 251.471
R393 VDDA.t231 VDDA.t223 251.471
R394 VDDA.t32 VDDA.t231 251.471
R395 VDDA.t54 VDDA.t32 251.471
R396 VDDA.t313 VDDA.t54 251.471
R397 VDDA.n596 VDDA.n595 243.698
R398 VDDA.n304 VDDA.n303 238.367
R399 VDDA.n303 VDDA.n253 238.367
R400 VDDA.n297 VDDA.n296 238.367
R401 VDDA.n296 VDDA.n273 238.367
R402 VDDA.n295 VDDA.n275 238.367
R403 VDDA.n295 VDDA.n294 238.367
R404 VDDA.t350 VDDA.n584 237.5
R405 VDDA.n597 VDDA.t313 237.5
R406 VDDA.t383 VDDA.t276 217.708
R407 VDDA.t276 VDDA.t293 217.708
R408 VDDA.t293 VDDA.t272 217.708
R409 VDDA.t272 VDDA.t302 217.708
R410 VDDA.t302 VDDA.t280 217.708
R411 VDDA.t280 VDDA.t299 217.708
R412 VDDA.t299 VDDA.t279 217.708
R413 VDDA.t279 VDDA.t297 217.708
R414 VDDA.t297 VDDA.t306 217.708
R415 VDDA.t306 VDDA.t283 217.708
R416 VDDA.t283 VDDA.t404 217.708
R417 VDDA.t177 VDDA.t319 217.708
R418 VDDA.t158 VDDA.t177 217.708
R419 VDDA.t258 VDDA.t158 217.708
R420 VDDA.t215 VDDA.t258 217.708
R421 VDDA.t175 VDDA.t215 217.708
R422 VDDA.t180 VDDA.t175 217.708
R423 VDDA.t174 VDDA.t180 217.708
R424 VDDA.t190 VDDA.t174 217.708
R425 VDDA.t173 VDDA.t190 217.708
R426 VDDA.t260 VDDA.t173 217.708
R427 VDDA.t337 VDDA.t260 217.708
R428 VDDA.t340 VDDA.n519 213.131
R429 VDDA.n520 VDDA.t377 213.131
R430 VDDA.t398 VDDA.n458 213.131
R431 VDDA.n459 VDDA.t353 213.131
R432 VDDA.t325 VDDA.n377 213.131
R433 VDDA.n378 VDDA.t395 213.131
R434 VDDA.n583 VDDA.n582 190.333
R435 VDDA.n588 VDDA.n587 185
R436 VDDA.n593 VDDA.n586 185
R437 VDDA.n597 VDDA.n586 185
R438 VDDA.n592 VDDA.n591 185
R439 VDDA.n590 VDDA.n545 185
R440 VDDA.n599 VDDA.n598 185
R441 VDDA.n598 VDDA.n597 185
R442 VDDA.n584 VDDA.n583 185
R443 VDDA.n581 VDDA.n549 185
R444 VDDA.n580 VDDA.n551 185
R445 VDDA.n579 VDDA.n552 185
R446 VDDA.n554 VDDA.n553 185
R447 VDDA.n576 VDDA.n548 185
R448 VDDA.n584 VDDA.n548 185
R449 VDDA.n543 VDDA.n542 168.435
R450 VDDA.n561 VDDA.n560 168.435
R451 VDDA.n563 VDDA.n562 168.435
R452 VDDA.n565 VDDA.n564 168.435
R453 VDDA.n567 VDDA.n566 168.435
R454 VDDA.n569 VDDA.n568 168.435
R455 VDDA.n571 VDDA.n570 168.435
R456 VDDA.n573 VDDA.n572 168.435
R457 VDDA.n512 VDDA.t332 168.139
R458 VDDA.n511 VDDA.t348 168.139
R459 VDDA.n509 VDDA.n508 153.576
R460 VDDA.n587 VDDA.n586 150
R461 VDDA.n591 VDDA.n586 150
R462 VDDA.n598 VDDA.n545 150
R463 VDDA.n583 VDDA.n549 150
R464 VDDA.n552 VDDA.n551 150
R465 VDDA.n553 VDDA.n548 150
R466 VDDA.t229 VDDA.t340 146.155
R467 VDDA.t377 VDDA.t229 146.155
R468 VDDA.t22 VDDA.t398 146.155
R469 VDDA.t458 VDDA.t22 146.155
R470 VDDA.t122 VDDA.t458 146.155
R471 VDDA.t49 VDDA.t122 146.155
R472 VDDA.t72 VDDA.t49 146.155
R473 VDDA.t87 VDDA.t72 146.155
R474 VDDA.t102 VDDA.t87 146.155
R475 VDDA.t155 VDDA.t102 146.155
R476 VDDA.t13 VDDA.t155 146.155
R477 VDDA.t89 VDDA.t13 146.155
R478 VDDA.t353 VDDA.t89 146.155
R479 VDDA.t466 VDDA.t325 146.155
R480 VDDA.t85 VDDA.t466 146.155
R481 VDDA.t453 VDDA.t85 146.155
R482 VDDA.t153 VDDA.t453 146.155
R483 VDDA.t96 VDDA.t153 146.155
R484 VDDA.t15 VDDA.t96 146.155
R485 VDDA.t451 VDDA.t15 146.155
R486 VDDA.t124 VDDA.t451 146.155
R487 VDDA.t130 VDDA.t124 146.155
R488 VDDA.t67 VDDA.t130 146.155
R489 VDDA.t395 VDDA.t67 146.155
R490 VDDA.n480 VDDA.t384 136.701
R491 VDDA.n479 VDDA.t405 136.701
R492 VDDA.n398 VDDA.t320 136.701
R493 VDDA.n399 VDDA.t338 136.701
R494 VDDA.t351 VDDA.n550 123.126
R495 VDDA.n578 VDDA.t351 123.126
R496 VDDA.n594 VDDA.t314 123.126
R497 VDDA.n589 VDDA.t314 123.126
R498 VDDA.n502 VDDA.t359 122.829
R499 VDDA.t371 VDDA.n501 122.829
R500 VDDA.t410 VDDA.n420 122.829
R501 VDDA.n421 VDDA.t422 122.829
R502 VDDA.t359 VDDA.t303 81.6411
R503 VDDA.t303 VDDA.t281 81.6411
R504 VDDA.t281 VDDA.t300 81.6411
R505 VDDA.t300 VDDA.t291 81.6411
R506 VDDA.t291 VDDA.t270 81.6411
R507 VDDA.t270 VDDA.t287 81.6411
R508 VDDA.t287 VDDA.t307 81.6411
R509 VDDA.t307 VDDA.t284 81.6411
R510 VDDA.t284 VDDA.t295 81.6411
R511 VDDA.t295 VDDA.t274 81.6411
R512 VDDA.t274 VDDA.t371 81.6411
R513 VDDA.t170 VDDA.t410 81.6411
R514 VDDA.t261 VDDA.t170 81.6411
R515 VDDA.t163 VDDA.t261 81.6411
R516 VDDA.t186 VDDA.t163 81.6411
R517 VDDA.t256 VDDA.t186 81.6411
R518 VDDA.t209 VDDA.t256 81.6411
R519 VDDA.t161 VDDA.t209 81.6411
R520 VDDA.t207 VDDA.t161 81.6411
R521 VDDA.t159 VDDA.t207 81.6411
R522 VDDA.t178 VDDA.t159 81.6411
R523 VDDA.t422 VDDA.t178 81.6411
R524 VDDA.n424 VDDA.t76 78.8005
R525 VDDA.n424 VDDA.t252 78.8005
R526 VDDA.n426 VDDA.t183 78.8005
R527 VDDA.n426 VDDA.t196 78.8005
R528 VDDA.n428 VDDA.t167 78.8005
R529 VDDA.n428 VDDA.t192 78.8005
R530 VDDA.n430 VDDA.t169 78.8005
R531 VDDA.n430 VDDA.t194 78.8005
R532 VDDA.n432 VDDA.t254 78.8005
R533 VDDA.n432 VDDA.t214 78.8005
R534 VDDA.n434 VDDA.t206 78.8005
R535 VDDA.n434 VDDA.t202 78.8005
R536 VDDA.n436 VDDA.t264 78.8005
R537 VDDA.n436 VDDA.t78 78.8005
R538 VDDA.n438 VDDA.t266 78.8005
R539 VDDA.n438 VDDA.t204 78.8005
R540 VDDA.n440 VDDA.t200 78.8005
R541 VDDA.n440 VDDA.t185 78.8005
R542 VDDA.n442 VDDA.t198 78.8005
R543 VDDA.n442 VDDA.t212 78.8005
R544 VDDA.n519 VDDA.t341 76.2576
R545 VDDA.n520 VDDA.t378 76.2576
R546 VDDA.n458 VDDA.t399 76.2576
R547 VDDA.n459 VDDA.t354 76.2576
R548 VDDA.n377 VDDA.t326 76.2576
R549 VDDA.n378 VDDA.t396 76.2576
R550 VDDA.n454 VDDA.n453 71.513
R551 VDDA.n456 VDDA.n455 71.513
R552 VDDA.n462 VDDA.n461 71.513
R553 VDDA.n464 VDDA.n463 71.513
R554 VDDA.n373 VDDA.n372 71.513
R555 VDDA.n375 VDDA.n374 71.513
R556 VDDA.n381 VDDA.n380 71.513
R557 VDDA.n383 VDDA.n382 71.513
R558 VDDA.n517 VDDA.n516 71.388
R559 VDDA.n466 VDDA.n452 67.013
R560 VDDA.n385 VDDA.n371 67.013
R561 VDDA.n597 VDDA.n596 65.8183
R562 VDDA.n597 VDDA.n585 65.8183
R563 VDDA.n584 VDDA.n546 65.8183
R564 VDDA.n584 VDDA.n547 65.8183
R565 VDDA.n229 VDDA.t687 59.5681
R566 VDDA.n230 VDDA.t648 59.5681
R567 VDDA.n591 VDDA.n585 53.3664
R568 VDDA.n596 VDDA.n587 53.3664
R569 VDDA.n585 VDDA.n545 53.3664
R570 VDDA.n549 VDDA.n546 53.3664
R571 VDDA.n552 VDDA.n547 53.3664
R572 VDDA.n551 VDDA.n546 53.3664
R573 VDDA.n553 VDDA.n547 53.3664
R574 VDDA.n229 VDDA.t733 52.3877
R575 VDDA.n231 VDDA.t653 48.9557
R576 VDDA.n491 VDDA.n490 41.1393
R577 VDDA.n493 VDDA.n492 41.1393
R578 VDDA.n495 VDDA.n494 41.1393
R579 VDDA.n497 VDDA.n496 41.1393
R580 VDDA.n499 VDDA.n498 41.1393
R581 VDDA.n410 VDDA.n409 41.1393
R582 VDDA.n412 VDDA.n411 41.1393
R583 VDDA.n414 VDDA.n413 41.1393
R584 VDDA.n416 VDDA.n415 41.1393
R585 VDDA.n418 VDDA.n417 41.1393
R586 VDDA.n502 VDDA.t360 40.9789
R587 VDDA.n501 VDDA.t372 40.9789
R588 VDDA.n420 VDDA.t411 40.9789
R589 VDDA.n421 VDDA.t423 40.9789
R590 VDDA.n627 VDDA.t237 39.4831
R591 VDDA.n540 VDDA.t10 39.4005
R592 VDDA.n540 VDDA.t152 39.4005
R593 VDDA.n359 VDDA.t437 39.4005
R594 VDDA.n359 VDDA.t463 39.4005
R595 VDDA.n326 VDDA.t150 39.4005
R596 VDDA.n326 VDDA.t121 39.4005
R597 VDDA.n346 VDDA.t465 39.4005
R598 VDDA.n346 VDDA.t101 39.4005
R599 VDDA.n328 VDDA.t450 39.4005
R600 VDDA.n328 VDDA.t457 39.4005
R601 VDDA.n330 VDDA.t226 39.4005
R602 VDDA.n330 VDDA.t119 39.4005
R603 VDDA.n354 VDDA.t129 39.4005
R604 VDDA.n354 VDDA.t446 39.4005
R605 VDDA.n356 VDDA.t448 39.4005
R606 VDDA.n356 VDDA.t110 39.4005
R607 VDDA.n337 VDDA.t48 39.4005
R608 VDDA.n337 VDDA.t46 39.4005
R609 VDDA.n339 VDDA.t12 39.4005
R610 VDDA.n339 VDDA.t148 39.4005
R611 VDDA.n251 VDDA.t31 39.4005
R612 VDDA.n251 VDDA.t425 39.4005
R613 VDDA.n255 VDDA.t246 39.4005
R614 VDDA.n255 VDDA.t250 39.4005
R615 VDDA.n257 VDDA.t39 39.4005
R616 VDDA.n257 VDDA.t106 39.4005
R617 VDDA.n259 VDDA.t62 39.4005
R618 VDDA.n259 VDDA.t268 39.4005
R619 VDDA.n261 VDDA.t113 39.4005
R620 VDDA.n261 VDDA.t433 39.4005
R621 VDDA.n263 VDDA.t244 39.4005
R622 VDDA.n263 VDDA.t115 39.4005
R623 VDDA.n265 VDDA.t6 39.4005
R624 VDDA.n265 VDDA.t236 39.4005
R625 VDDA.n267 VDDA.t26 39.4005
R626 VDDA.n267 VDDA.t21 39.4005
R627 VDDA.n269 VDDA.t135 39.4005
R628 VDDA.n269 VDDA.t108 39.4005
R629 VDDA.n271 VDDA.t80 39.4005
R630 VDDA.n271 VDDA.t444 39.4005
R631 VDDA.n276 VDDA.t52 39.4005
R632 VDDA.n276 VDDA.t228 39.4005
R633 VDDA.n278 VDDA.t117 39.4005
R634 VDDA.n278 VDDA.t64 39.4005
R635 VDDA.n280 VDDA.t71 39.4005
R636 VDDA.n280 VDDA.t8 39.4005
R637 VDDA.n282 VDDA.t461 39.4005
R638 VDDA.n282 VDDA.t1 39.4005
R639 VDDA.n284 VDDA.t84 39.4005
R640 VDDA.n284 VDDA.t42 39.4005
R641 VDDA.n286 VDDA.t66 39.4005
R642 VDDA.n286 VDDA.t439 39.4005
R643 VDDA.n288 VDDA.t220 39.4005
R644 VDDA.n288 VDDA.t99 39.4005
R645 VDDA.n290 VDDA.t127 39.4005
R646 VDDA.n290 VDDA.t82 39.4005
R647 VDDA.n469 VDDA.n467 30.2255
R648 VDDA.n388 VDDA.n386 30.2255
R649 VDDA.n477 VDDA.n476 29.663
R650 VDDA.n475 VDDA.n474 29.663
R651 VDDA.n473 VDDA.n472 29.663
R652 VDDA.n471 VDDA.n470 29.663
R653 VDDA.n469 VDDA.n468 29.663
R654 VDDA.n396 VDDA.n395 29.663
R655 VDDA.n394 VDDA.n393 29.663
R656 VDDA.n392 VDDA.n391 29.663
R657 VDDA.n390 VDDA.n389 29.663
R658 VDDA.n388 VDDA.n387 29.663
R659 VDDA.n335 VDDA.n334 27.2462
R660 VDDA.n333 VDDA.n332 27.2462
R661 VDDA.n344 VDDA.n343 27.2462
R662 VDDA.n342 VDDA.n341 27.2462
R663 VDDA.n536 VDDA.n535 25.087
R664 VDDA.n538 VDDA.n537 25.087
R665 VDDA.n352 VDDA.n351 25.0384
R666 VDDA.n350 VDDA.n349 25.0384
R667 VDDA.n556 VDDA.n555 22.9536
R668 VDDA.n302 VDDA.n301 22.9536
R669 VDDA.n600 VDDA.n599 22.8576
R670 VDDA.n576 VDDA.n575 22.8576
R671 VDDA.n508 VDDA.t3 21.8894
R672 VDDA.n508 VDDA.t347 21.8894
R673 VDDA.n305 VDDA.n253 20.7243
R674 VDDA.n298 VDDA.n273 20.7243
R675 VDDA.n292 VDDA.n275 20.7243
R676 VDDA.n558 VDDA.n557 20.4312
R677 VDDA.n232 VDDA.n231 18.8097
R678 VDDA.n559 VDDA.n555 15.488
R679 VDDA.n292 VDDA.n291 14.6963
R680 VDDA.n539 VDDA.n538 14.363
R681 VDDA.n539 VDDA.n535 14.363
R682 VDDA.n332 VDDA.n331 14.363
R683 VDDA.n341 VDDA.n340 14.363
R684 VDDA.n559 VDDA.n558 14.238
R685 VDDA.n301 VDDA.n300 14.0713
R686 VDDA.n306 VDDA.n305 14.0713
R687 VDDA.n299 VDDA.n298 14.0713
R688 VDDA.n575 VDDA.n574 13.8005
R689 VDDA.n601 VDDA.n600 13.8005
R690 VDDA.n336 VDDA.n335 13.8005
R691 VDDA.n353 VDDA.n352 13.8005
R692 VDDA.n349 VDDA.n348 13.8005
R693 VDDA.n345 VDDA.n344 13.8005
R694 VDDA.n542 VDDA.t33 13.1338
R695 VDDA.n542 VDDA.t55 13.1338
R696 VDDA.n560 VDDA.t224 13.1338
R697 VDDA.n560 VDDA.t232 13.1338
R698 VDDA.n562 VDDA.t139 13.1338
R699 VDDA.n562 VDDA.t145 13.1338
R700 VDDA.n564 VDDA.t234 13.1338
R701 VDDA.n564 VDDA.t35 13.1338
R702 VDDA.n566 VDDA.t143 13.1338
R703 VDDA.n566 VDDA.t239 13.1338
R704 VDDA.n568 VDDA.t94 13.1338
R705 VDDA.n568 VDDA.t217 13.1338
R706 VDDA.n570 VDDA.t137 13.1338
R707 VDDA.n570 VDDA.t222 13.1338
R708 VDDA.n572 VDDA.t28 13.1338
R709 VDDA.n572 VDDA.t60 13.1338
R710 VDDA.n307 VDDA.n306 12.5786
R711 VDDA.n483 VDDA.n477 11.3443
R712 VDDA.n402 VDDA.n396 11.3443
R713 VDDA.t341 VDDA.n517 11.2576
R714 VDDA.n517 VDDA.t230 11.2576
R715 VDDA.n453 VDDA.t123 11.2576
R716 VDDA.n453 VDDA.t50 11.2576
R717 VDDA.n455 VDDA.t23 11.2576
R718 VDDA.n455 VDDA.t459 11.2576
R719 VDDA.n461 VDDA.t14 11.2576
R720 VDDA.n461 VDDA.t90 11.2576
R721 VDDA.n463 VDDA.t103 11.2576
R722 VDDA.n463 VDDA.t156 11.2576
R723 VDDA.n452 VDDA.t73 11.2576
R724 VDDA.n452 VDDA.t88 11.2576
R725 VDDA.n372 VDDA.t454 11.2576
R726 VDDA.n372 VDDA.t154 11.2576
R727 VDDA.n374 VDDA.t467 11.2576
R728 VDDA.n374 VDDA.t86 11.2576
R729 VDDA.n380 VDDA.t131 11.2576
R730 VDDA.n380 VDDA.t68 11.2576
R731 VDDA.n382 VDDA.t452 11.2576
R732 VDDA.n382 VDDA.t125 11.2576
R733 VDDA.n371 VDDA.t97 11.2576
R734 VDDA.n371 VDDA.t16 11.2576
R735 VDDA.n524 VDDA.n523 9.7005
R736 VDDA.n487 VDDA.n486 9.5505
R737 VDDA.n485 VDDA.n484 9.5505
R738 VDDA.n406 VDDA.n405 9.5505
R739 VDDA.n404 VDDA.n403 9.5505
R740 VDDA.n506 VDDA.n505 9.5005
R741 VDDA.n451 VDDA.n450 9.5005
R742 VDDA.n447 VDDA.n446 9.3005
R743 VDDA.n445 VDDA.n444 9.3005
R744 VDDA.n593 VDDA.n588 9.14336
R745 VDDA.n593 VDDA.n592 9.14336
R746 VDDA.n592 VDDA.n590 9.14336
R747 VDDA.n581 VDDA.n580 9.14336
R748 VDDA.n580 VDDA.n579 9.14336
R749 VDDA.n579 VDDA.n554 9.14336
R750 VDDA.n488 VDDA.n484 9.02133
R751 VDDA.n407 VDDA.n403 9.02133
R752 VDDA.n482 VDDA.n478 8.79217
R753 VDDA.n401 VDDA.n397 8.79217
R754 VDDA.n476 VDDA.t40 8.0005
R755 VDDA.n476 VDDA.t269 8.0005
R756 VDDA.n474 VDDA.t286 8.0005
R757 VDDA.n474 VDDA.t305 8.0005
R758 VDDA.n472 VDDA.t298 8.0005
R759 VDDA.n472 VDDA.t278 8.0005
R760 VDDA.n470 VDDA.t294 8.0005
R761 VDDA.n470 VDDA.t273 8.0005
R762 VDDA.n468 VDDA.t290 8.0005
R763 VDDA.n468 VDDA.t289 8.0005
R764 VDDA.n467 VDDA.t277 8.0005
R765 VDDA.n467 VDDA.t441 8.0005
R766 VDDA.n395 VDDA.t188 8.0005
R767 VDDA.n395 VDDA.t44 8.0005
R768 VDDA.n393 VDDA.t241 8.0005
R769 VDDA.n393 VDDA.t165 8.0005
R770 VDDA.n391 VDDA.t242 8.0005
R771 VDDA.n391 VDDA.t255 8.0005
R772 VDDA.n389 VDDA.t181 8.0005
R773 VDDA.n389 VDDA.t172 8.0005
R774 VDDA.n387 VDDA.t189 8.0005
R775 VDDA.n387 VDDA.t176 8.0005
R776 VDDA.n386 VDDA.t440 8.0005
R777 VDDA.n386 VDDA.t259 8.0005
R778 VDDA.n506 VDDA.n466 7.71925
R779 VDDA.n451 VDDA.n385 7.71925
R780 VDDA.n602 VDDA.n601 7.0005
R781 VDDA.n507 VDDA.n451 6.90675
R782 VDDA.n507 VDDA.n506 6.8755
R783 VDDA.n515 VDDA.n507 6.813
R784 VDDA.n490 VDDA.t304 6.56717
R785 VDDA.n490 VDDA.t282 6.56717
R786 VDDA.n492 VDDA.t301 6.56717
R787 VDDA.n492 VDDA.t292 6.56717
R788 VDDA.n494 VDDA.t271 6.56717
R789 VDDA.n494 VDDA.t288 6.56717
R790 VDDA.n496 VDDA.t308 6.56717
R791 VDDA.n496 VDDA.t285 6.56717
R792 VDDA.n498 VDDA.t296 6.56717
R793 VDDA.n498 VDDA.t275 6.56717
R794 VDDA.n409 VDDA.t160 6.56717
R795 VDDA.n409 VDDA.t179 6.56717
R796 VDDA.n411 VDDA.t162 6.56717
R797 VDDA.n411 VDDA.t208 6.56717
R798 VDDA.n413 VDDA.t257 6.56717
R799 VDDA.n413 VDDA.t210 6.56717
R800 VDDA.n415 VDDA.t164 6.56717
R801 VDDA.n415 VDDA.t187 6.56717
R802 VDDA.n417 VDDA.t171 6.56717
R803 VDDA.n417 VDDA.t262 6.56717
R804 VDDA.n462 VDDA.n460 6.10467
R805 VDDA.n457 VDDA.n456 6.10467
R806 VDDA.n381 VDDA.n379 6.10467
R807 VDDA.n376 VDDA.n375 6.10467
R808 VDDA.n408 VDDA.n407 6.09425
R809 VDDA.n489 VDDA.n488 6.063
R810 VDDA.n444 VDDA.n443 5.60467
R811 VDDA.n599 VDDA.n544 5.33286
R812 VDDA.n577 VDDA.n576 5.33286
R813 VDDA.n500 VDDA.n499 5.313
R814 VDDA.n419 VDDA.n418 5.313
R815 VDDA.n523 VDDA.n522 5.28175
R816 VDDA.n515 VDDA.n514 5.28175
R817 VDDA.n505 VDDA.n504 5.28175
R818 VDDA.n483 VDDA.n482 5.28175
R819 VDDA.n402 VDDA.n401 5.28175
R820 VDDA.n448 VDDA.n447 5.04217
R821 VDDA.n488 VDDA.n487 5.02133
R822 VDDA.n407 VDDA.n406 5.02133
R823 VDDA.n5 VDDA.t480 4.8295
R824 VDDA.n9 VDDA.t474 4.8295
R825 VDDA.n14 VDDA.t670 4.8295
R826 VDDA.n18 VDDA.t662 4.8295
R827 VDDA.n23 VDDA.t469 4.8295
R828 VDDA.n27 VDDA.t734 4.8295
R829 VDDA.n32 VDDA.t659 4.8295
R830 VDDA.n36 VDDA.t655 4.8295
R831 VDDA.n41 VDDA.t585 4.8295
R832 VDDA.n45 VDDA.t580 4.8295
R833 VDDA.n50 VDDA.t512 4.8295
R834 VDDA.n54 VDDA.t506 4.8295
R835 VDDA.n59 VDDA.t575 4.8295
R836 VDDA.n63 VDDA.t569 4.8295
R837 VDDA.n68 VDDA.t501 4.8295
R838 VDDA.n72 VDDA.t495 4.8295
R839 VDDA.n77 VDDA.t694 4.8295
R840 VDDA.n81 VDDA.t688 4.8295
R841 VDDA.n86 VDDA.t491 4.8295
R842 VDDA.n90 VDDA.t486 4.8295
R843 VDDA.n95 VDDA.t683 4.8295
R844 VDDA.n99 VDDA.t675 4.8295
R845 VDDA.n104 VDDA.t606 4.8295
R846 VDDA.n108 VDDA.t600 4.8295
R847 VDDA.n113 VDDA.t671 4.8295
R848 VDDA.n117 VDDA.t664 4.8295
R849 VDDA.n122 VDDA.t596 4.8295
R850 VDDA.n126 VDDA.t589 4.8295
R851 VDDA.n131 VDDA.t532 4.8295
R852 VDDA.n135 VDDA.t528 4.8295
R853 VDDA.n140 VDDA.t723 4.8295
R854 VDDA.n144 VDDA.t719 4.8295
R855 VDDA.n149 VDDA.t522 4.8295
R856 VDDA.n153 VDDA.t519 4.8295
R857 VDDA.n158 VDDA.t712 4.8295
R858 VDDA.n162 VDDA.t708 4.8295
R859 VDDA.n167 VDDA.t634 4.8295
R860 VDDA.n171 VDDA.t631 4.8295
R861 VDDA.n176 VDDA.t703 4.8295
R862 VDDA.n180 VDDA.t700 4.8295
R863 VDDA.n185 VDDA.t626 4.8295
R864 VDDA.n189 VDDA.t622 4.8295
R865 VDDA.n194 VDDA.t552 4.8295
R866 VDDA.n198 VDDA.t547 4.8295
R867 VDDA.n203 VDDA.t616 4.8295
R868 VDDA.n207 VDDA.t613 4.8295
R869 VDDA.n212 VDDA.t542 4.8295
R870 VDDA.n482 VDDA.n481 4.79217
R871 VDDA.n401 VDDA.n400 4.79217
R872 VDDA.n518 VDDA.n516 4.7505
R873 VDDA.n510 VDDA.n509 4.7505
R874 VDDA.n504 VDDA.n503 4.7505
R875 VDDA.n423 VDDA.n422 4.7505
R876 VDDA.n254 VDDA.n253 4.54311
R877 VDDA.n304 VDDA.n254 4.54311
R878 VDDA.n274 VDDA.n273 4.54311
R879 VDDA.n297 VDDA.n274 4.54311
R880 VDDA.n293 VDDA.n275 4.54311
R881 VDDA.n294 VDDA.n293 4.54311
R882 VDDA.n541 VDDA.n539 4.5005
R883 VDDA.n603 VDDA.n534 4.5005
R884 VDDA.n606 VDDA.n604 4.5005
R885 VDDA.n607 VDDA.n533 4.5005
R886 VDDA.n611 VDDA.n610 4.5005
R887 VDDA.n360 VDDA.n358 4.5005
R888 VDDA.n522 VDDA.n521 4.5005
R889 VDDA.n514 VDDA.n513 4.5005
R890 VDDA.n466 VDDA.n465 4.5005
R891 VDDA.n450 VDDA.n449 4.5005
R892 VDDA.n385 VDDA.n384 4.5005
R893 VDDA.n361 VDDA.n325 4.5005
R894 VDDA.n364 VDDA.n362 4.5005
R895 VDDA.n365 VDDA.n324 4.5005
R896 VDDA.n369 VDDA.n368 4.5005
R897 VDDA.n370 VDDA.n323 4.5005
R898 VDDA.n525 VDDA.n524 4.5005
R899 VDDA.n627 VDDA.n621 4.5005
R900 VDDA.n630 VDDA.n628 4.5005
R901 VDDA.n631 VDDA.n620 4.5005
R902 VDDA.n635 VDDA.n634 4.5005
R903 VDDA.n232 VDDA.n228 4.5005
R904 VDDA.n235 VDDA.n233 4.5005
R905 VDDA.n236 VDDA.n227 4.5005
R906 VDDA.n240 VDDA.n239 4.5005
R907 VDDA.n307 VDDA.n250 4.5005
R908 VDDA.n310 VDDA.n308 4.5005
R909 VDDA.n311 VDDA.n249 4.5005
R910 VDDA.n315 VDDA.n314 4.5005
R911 VDDA.n5 VDDA.t526 4.5005
R912 VDDA.n6 VDDA.t559 4.5005
R913 VDDA.n7 VDDA.t487 4.5005
R914 VDDA.n8 VDDA.t682 4.5005
R915 VDDA.n13 VDDA.t724 4.5005
R916 VDDA.n12 VDDA.t649 4.5005
R917 VDDA.n11 VDDA.t577 4.5005
R918 VDDA.n10 VDDA.t621 4.5005
R919 VDDA.n9 VDDA.t549 4.5005
R920 VDDA.n14 VDDA.t716 4.5005
R921 VDDA.n15 VDDA.t482 4.5005
R922 VDDA.n16 VDDA.t677 4.5005
R923 VDDA.n17 VDDA.t603 4.5005
R924 VDDA.n22 VDDA.t643 4.5005
R925 VDDA.n21 VDDA.t573 4.5005
R926 VDDA.n20 VDDA.t502 4.5005
R927 VDDA.n19 VDDA.t545 4.5005
R928 VDDA.n18 VDDA.t470 4.5005
R929 VDDA.n23 VDDA.t516 4.5005
R930 VDDA.n24 VDDA.t550 4.5005
R931 VDDA.n25 VDDA.t476 4.5005
R932 VDDA.n26 VDDA.t669 4.5005
R933 VDDA.n31 VDDA.t713 4.5005
R934 VDDA.n30 VDDA.t639 4.5005
R935 VDDA.n29 VDDA.t568 4.5005
R936 VDDA.n28 VDDA.t610 4.5005
R937 VDDA.n27 VDDA.t540 4.5005
R938 VDDA.n32 VDDA.t707 4.5005
R939 VDDA.n33 VDDA.t472 4.5005
R940 VDDA.n34 VDDA.t665 4.5005
R941 VDDA.n35 VDDA.t595 4.5005
R942 VDDA.n40 VDDA.t635 4.5005
R943 VDDA.n39 VDDA.t564 4.5005
R944 VDDA.n38 VDDA.t494 4.5005
R945 VDDA.n37 VDDA.t536 4.5005
R946 VDDA.n36 VDDA.t729 4.5005
R947 VDDA.n41 VDDA.t628 4.5005
R948 VDDA.n42 VDDA.t661 4.5005
R949 VDDA.n43 VDDA.t590 4.5005
R950 VDDA.n44 VDDA.t521 4.5005
R951 VDDA.n49 VDDA.t561 4.5005
R952 VDDA.n48 VDDA.t489 4.5005
R953 VDDA.n47 VDDA.t686 4.5005
R954 VDDA.n46 VDDA.t727 4.5005
R955 VDDA.n45 VDDA.t650 4.5005
R956 VDDA.n50 VDDA.t553 4.5005
R957 VDDA.n51 VDDA.t586 4.5005
R958 VDDA.n52 VDDA.t517 4.5005
R959 VDDA.n53 VDDA.t711 4.5005
R960 VDDA.n58 VDDA.t485 4.5005
R961 VDDA.n57 VDDA.t680 4.5005
R962 VDDA.n56 VDDA.t608 4.5005
R963 VDDA.n55 VDDA.t647 4.5005
R964 VDDA.n54 VDDA.t576 4.5005
R965 VDDA.n59 VDDA.t620 4.5005
R966 VDDA.n60 VDDA.t651 4.5005
R967 VDDA.n61 VDDA.t581 4.5005
R968 VDDA.n62 VDDA.t511 4.5005
R969 VDDA.n67 VDDA.t554 4.5005
R970 VDDA.n66 VDDA.t479 4.5005
R971 VDDA.n65 VDDA.t673 4.5005
R972 VDDA.n64 VDDA.t718 4.5005
R973 VDDA.n63 VDDA.t641 4.5005
R974 VDDA.n68 VDDA.t544 4.5005
R975 VDDA.n69 VDDA.t578 4.5005
R976 VDDA.n70 VDDA.t508 4.5005
R977 VDDA.n71 VDDA.t702 4.5005
R978 VDDA.n76 VDDA.t475 4.5005
R979 VDDA.n75 VDDA.t668 4.5005
R980 VDDA.n74 VDDA.t597 4.5005
R981 VDDA.n73 VDDA.t638 4.5005
R982 VDDA.n72 VDDA.t565 4.5005
R983 VDDA.n77 VDDA.t735 4.5005
R984 VDDA.n78 VDDA.t503 4.5005
R985 VDDA.n79 VDDA.t699 4.5005
R986 VDDA.n80 VDDA.t625 4.5005
R987 VDDA.n85 VDDA.t663 4.5005
R988 VDDA.n84 VDDA.t594 4.5005
R989 VDDA.n83 VDDA.t523 4.5005
R990 VDDA.n82 VDDA.t563 4.5005
R991 VDDA.n81 VDDA.t492 4.5005
R992 VDDA.n86 VDDA.t535 4.5005
R993 VDDA.n87 VDDA.t566 4.5005
R994 VDDA.n88 VDDA.t496 4.5005
R995 VDDA.n89 VDDA.t693 4.5005
R996 VDDA.n94 VDDA.t731 4.5005
R997 VDDA.n93 VDDA.t658 4.5005
R998 VDDA.n92 VDDA.t588 4.5005
R999 VDDA.n91 VDDA.t630 4.5005
R1000 VDDA.n90 VDDA.t558 4.5005
R1001 VDDA.n95 VDDA.t726 4.5005
R1002 VDDA.n96 VDDA.t493 4.5005
R1003 VDDA.n97 VDDA.t689 4.5005
R1004 VDDA.n98 VDDA.t615 4.5005
R1005 VDDA.n103 VDDA.t654 4.5005
R1006 VDDA.n102 VDDA.t584 4.5005
R1007 VDDA.n101 VDDA.t514 4.5005
R1008 VDDA.n100 VDDA.t556 4.5005
R1009 VDDA.n99 VDDA.t481 4.5005
R1010 VDDA.n104 VDDA.t646 4.5005
R1011 VDDA.n105 VDDA.t684 4.5005
R1012 VDDA.n106 VDDA.t611 4.5005
R1013 VDDA.n107 VDDA.t541 4.5005
R1014 VDDA.n112 VDDA.t579 4.5005
R1015 VDDA.n111 VDDA.t510 4.5005
R1016 VDDA.n110 VDDA.t705 4.5005
R1017 VDDA.n109 VDDA.t478 4.5005
R1018 VDDA.n108 VDDA.t672 4.5005
R1019 VDDA.n113 VDDA.t717 4.5005
R1020 VDDA.n114 VDDA.t483 4.5005
R1021 VDDA.n115 VDDA.t678 4.5005
R1022 VDDA.n116 VDDA.t604 4.5005
R1023 VDDA.n121 VDDA.t644 4.5005
R1024 VDDA.n120 VDDA.t574 4.5005
R1025 VDDA.n119 VDDA.t504 4.5005
R1026 VDDA.n118 VDDA.t546 4.5005
R1027 VDDA.n117 VDDA.t471 4.5005
R1028 VDDA.n122 VDDA.t637 4.5005
R1029 VDDA.n123 VDDA.t674 4.5005
R1030 VDDA.n124 VDDA.t602 4.5005
R1031 VDDA.n125 VDDA.t530 4.5005
R1032 VDDA.n130 VDDA.t570 4.5005
R1033 VDDA.n129 VDDA.t500 4.5005
R1034 VDDA.n128 VDDA.t695 4.5005
R1035 VDDA.n127 VDDA.t736 4.5005
R1036 VDDA.n126 VDDA.t660 4.5005
R1037 VDDA.n131 VDDA.t571 4.5005
R1038 VDDA.n132 VDDA.t609 4.5005
R1039 VDDA.n133 VDDA.t538 4.5005
R1040 VDDA.n134 VDDA.t730 4.5005
R1041 VDDA.n139 VDDA.t507 4.5005
R1042 VDDA.n138 VDDA.t701 4.5005
R1043 VDDA.n137 VDDA.t629 4.5005
R1044 VDDA.n136 VDDA.t667 4.5005
R1045 VDDA.n135 VDDA.t598 4.5005
R1046 VDDA.n140 VDDA.t498 4.5005
R1047 VDDA.n141 VDDA.t533 4.5005
R1048 VDDA.n142 VDDA.t728 4.5005
R1049 VDDA.n143 VDDA.t652 4.5005
R1050 VDDA.n148 VDDA.t698 4.5005
R1051 VDDA.n147 VDDA.t624 4.5005
R1052 VDDA.n146 VDDA.t555 4.5005
R1053 VDDA.n145 VDDA.t593 4.5005
R1054 VDDA.n144 VDDA.t524 4.5005
R1055 VDDA.n149 VDDA.t562 4.5005
R1056 VDDA.n150 VDDA.t599 4.5005
R1057 VDDA.n151 VDDA.t529 4.5005
R1058 VDDA.n152 VDDA.t722 4.5005
R1059 VDDA.n157 VDDA.t497 4.5005
R1060 VDDA.n156 VDDA.t692 4.5005
R1061 VDDA.n155 VDDA.t619 4.5005
R1062 VDDA.n154 VDDA.t657 4.5005
R1063 VDDA.n153 VDDA.t587 4.5005
R1064 VDDA.n158 VDDA.t488 4.5005
R1065 VDDA.n159 VDDA.t525 4.5005
R1066 VDDA.n160 VDDA.t720 4.5005
R1067 VDDA.n161 VDDA.t642 4.5005
R1068 VDDA.n166 VDDA.t690 4.5005
R1069 VDDA.n165 VDDA.t614 4.5005
R1070 VDDA.n164 VDDA.t543 4.5005
R1071 VDDA.n163 VDDA.t583 4.5005
R1072 VDDA.n162 VDDA.t513 4.5005
R1073 VDDA.n167 VDDA.t679 4.5005
R1074 VDDA.n168 VDDA.t715 4.5005
R1075 VDDA.n169 VDDA.t640 4.5005
R1076 VDDA.n170 VDDA.t567 4.5005
R1077 VDDA.n175 VDDA.t612 4.5005
R1078 VDDA.n174 VDDA.t539 4.5005
R1079 VDDA.n173 VDDA.t732 4.5005
R1080 VDDA.n172 VDDA.t509 4.5005
R1081 VDDA.n171 VDDA.t704 4.5005
R1082 VDDA.n176 VDDA.t477 4.5005
R1083 VDDA.n177 VDDA.t515 4.5005
R1084 VDDA.n178 VDDA.t709 4.5005
R1085 VDDA.n179 VDDA.t633 4.5005
R1086 VDDA.n184 VDDA.t676 4.5005
R1087 VDDA.n183 VDDA.t605 4.5005
R1088 VDDA.n182 VDDA.t534 4.5005
R1089 VDDA.n181 VDDA.t572 4.5005
R1090 VDDA.n180 VDDA.t505 4.5005
R1091 VDDA.n185 VDDA.t666 4.5005
R1092 VDDA.n186 VDDA.t706 4.5005
R1093 VDDA.n187 VDDA.t632 4.5005
R1094 VDDA.n188 VDDA.t560 4.5005
R1095 VDDA.n193 VDDA.t601 4.5005
R1096 VDDA.n192 VDDA.t531 4.5005
R1097 VDDA.n191 VDDA.t725 4.5005
R1098 VDDA.n190 VDDA.t499 4.5005
R1099 VDDA.n189 VDDA.t696 4.5005
R1100 VDDA.n194 VDDA.t592 4.5005
R1101 VDDA.n195 VDDA.t627 4.5005
R1102 VDDA.n196 VDDA.t557 4.5005
R1103 VDDA.n197 VDDA.t484 4.5005
R1104 VDDA.n202 VDDA.t527 4.5005
R1105 VDDA.n201 VDDA.t721 4.5005
R1106 VDDA.n200 VDDA.t645 4.5005
R1107 VDDA.n199 VDDA.t691 4.5005
R1108 VDDA.n198 VDDA.t617 4.5005
R1109 VDDA.n203 VDDA.t656 4.5005
R1110 VDDA.n204 VDDA.t697 4.5005
R1111 VDDA.n205 VDDA.t623 4.5005
R1112 VDDA.n206 VDDA.t551 4.5005
R1113 VDDA.n211 VDDA.t591 4.5005
R1114 VDDA.n210 VDDA.t520 4.5005
R1115 VDDA.n209 VDDA.t714 4.5005
R1116 VDDA.n208 VDDA.t490 4.5005
R1117 VDDA.n207 VDDA.t685 4.5005
R1118 VDDA.n212 VDDA.t582 4.5005
R1119 VDDA.n213 VDDA.t618 4.5005
R1120 VDDA.n214 VDDA.t548 4.5005
R1121 VDDA.n215 VDDA.t473 4.5005
R1122 VDDA.n216 VDDA.t518 4.5005
R1123 VDDA.n217 VDDA.t710 4.5005
R1124 VDDA.n218 VDDA.t636 4.5005
R1125 VDDA.n219 VDDA.t681 4.5005
R1126 VDDA.n220 VDDA.t607 4.5005
R1127 VDDA.n221 VDDA.t537 4.5005
R1128 VDDA.n230 VDDA.n229 4.12334
R1129 VDDA.n505 VDDA.n489 3.84425
R1130 VDDA.n450 VDDA.n408 3.84425
R1131 VDDA.n595 VDDA.n588 3.75335
R1132 VDDA.n590 VDDA.n544 3.75335
R1133 VDDA.n582 VDDA.n581 3.75335
R1134 VDDA.n577 VDDA.n554 3.75335
R1135 VDDA.n613 VDDA.n612 3.47871
R1136 VDDA.n637 VDDA.n636 3.47871
R1137 VDDA.n242 VDDA.n241 3.47871
R1138 VDDA.n317 VDDA.n316 3.47871
R1139 VDDA.n231 VDDA.n230 3.43377
R1140 VDDA.n532 VDDA.n531 3.4105
R1141 VDDA.n610 VDDA.n609 3.4105
R1142 VDDA.n608 VDDA.n607 3.4105
R1143 VDDA.n606 VDDA.n605 3.4105
R1144 VDDA.n534 VDDA.n528 3.4105
R1145 VDDA.n323 VDDA.n322 3.4105
R1146 VDDA.n368 VDDA.n367 3.4105
R1147 VDDA.n366 VDDA.n365 3.4105
R1148 VDDA.n364 VDDA.n363 3.4105
R1149 VDDA.n325 VDDA.n319 3.4105
R1150 VDDA.n526 VDDA.n525 3.4105
R1151 VDDA.n619 VDDA.n618 3.4105
R1152 VDDA.n634 VDDA.n633 3.4105
R1153 VDDA.n632 VDDA.n631 3.4105
R1154 VDDA.n630 VDDA.n629 3.4105
R1155 VDDA.n621 VDDA.n615 3.4105
R1156 VDDA.n226 VDDA.n225 3.4105
R1157 VDDA.n239 VDDA.n238 3.4105
R1158 VDDA.n237 VDDA.n236 3.4105
R1159 VDDA.n235 VDDA.n234 3.4105
R1160 VDDA.n228 VDDA.n222 3.4105
R1161 VDDA.n248 VDDA.n247 3.4105
R1162 VDDA.n314 VDDA.n313 3.4105
R1163 VDDA.n312 VDDA.n311 3.4105
R1164 VDDA.n310 VDDA.n309 3.4105
R1165 VDDA.n250 VDDA.n244 3.4105
R1166 VDDA.n318 VDDA.n244 3.4105
R1167 VDDA.n318 VDDA.n317 3.4105
R1168 VDDA.n243 VDDA.n222 3.4105
R1169 VDDA.n243 VDDA.n242 3.4105
R1170 VDDA.n638 VDDA.n615 3.4105
R1171 VDDA.n638 VDDA.n637 3.4105
R1172 VDDA.n527 VDDA.n319 3.4105
R1173 VDDA.n527 VDDA.n526 3.4105
R1174 VDDA.n614 VDDA.n528 3.4105
R1175 VDDA.n614 VDDA.n613 3.4105
R1176 VDDA.n653 VDDA.n3 3.4105
R1177 VDDA.n653 VDDA.n4 3.4105
R1178 VDDA.n653 VDDA.n652 3.4105
R1179 VDDA.n647 VDDA.n642 3.4105
R1180 VDDA.n652 VDDA.n642 3.4105
R1181 VDDA.n647 VDDA.n639 3.4105
R1182 VDDA.n646 VDDA.n639 3.4105
R1183 VDDA.n650 VDDA.n639 3.4105
R1184 VDDA.n645 VDDA.n639 3.4105
R1185 VDDA.n639 VDDA.n4 3.4105
R1186 VDDA.n652 VDDA.n639 3.4105
R1187 VDDA.n651 VDDA.n646 3.4105
R1188 VDDA.n651 VDDA.n650 3.4105
R1189 VDDA.n651 VDDA.n645 3.4105
R1190 VDDA.n651 VDDA.n4 3.4105
R1191 VDDA.n652 VDDA.n651 3.4105
R1192 VDDA.n603 VDDA.n602 3.29738
R1193 VDDA.n449 VDDA.n448 3.1255
R1194 VDDA.n513 VDDA.n512 2.8255
R1195 VDDA.n511 VDDA.n510 2.8255
R1196 VDDA.n481 VDDA.n480 2.423
R1197 VDDA.n479 VDDA.n478 2.423
R1198 VDDA.n400 VDDA.n399 2.423
R1199 VDDA.n398 VDDA.n397 2.423
R1200 VDDA.n612 VDDA.n611 2.39683
R1201 VDDA.n636 VDDA.n635 2.39683
R1202 VDDA.n241 VDDA.n240 2.39683
R1203 VDDA.n316 VDDA.n315 2.39683
R1204 VDDA.n503 VDDA.n502 1.97758
R1205 VDDA.n501 VDDA.n500 1.97758
R1206 VDDA.n422 VDDA.n421 1.97758
R1207 VDDA.n420 VDDA.n419 1.97758
R1208 VDDA.n521 VDDA.n520 1.888
R1209 VDDA.n519 VDDA.n518 1.888
R1210 VDDA.n300 VDDA.n299 1.8755
R1211 VDDA.n361 VDDA.n360 1.85675
R1212 VDDA.n574 VDDA.n559 1.84425
R1213 VDDA.n353 VDDA.n336 1.813
R1214 VDDA.n348 VDDA.n345 1.813
R1215 VDDA.n640 VDDA.n0 1.70468
R1216 VDDA.n643 VDDA.n640 1.70468
R1217 VDDA.n641 VDDA.n3 1.70453
R1218 VDDA.n653 VDDA.n2 1.70321
R1219 VDDA.n651 VDDA.n648 1.70321
R1220 VDDA.n653 VDDA.n1 1.70307
R1221 VDDA.n649 VDDA.n642 1.70307
R1222 VDDA.n644 VDDA.n642 1.70307
R1223 VDDA.n318 VDDA.n246 1.6924
R1224 VDDA.n318 VDDA.n245 1.6924
R1225 VDDA.n243 VDDA.n224 1.6924
R1226 VDDA.n243 VDDA.n223 1.6924
R1227 VDDA.n638 VDDA.n617 1.6924
R1228 VDDA.n638 VDDA.n616 1.6924
R1229 VDDA.n614 VDDA.n530 1.6924
R1230 VDDA.n614 VDDA.n529 1.6924
R1231 VDDA.n527 VDDA.n321 1.68971
R1232 VDDA.n527 VDDA.n320 1.68971
R1233 VDDA.n489 VDDA.n483 1.438
R1234 VDDA.n408 VDDA.n402 1.438
R1235 VDDA.n460 VDDA.n459 1.03383
R1236 VDDA.n458 VDDA.n457 1.03383
R1237 VDDA.n379 VDDA.n378 1.03383
R1238 VDDA.n377 VDDA.n376 1.03383
R1239 VDDA.n574 VDDA.n573 1.0005
R1240 VDDA.n573 VDDA.n571 1.0005
R1241 VDDA.n571 VDDA.n569 1.0005
R1242 VDDA.n569 VDDA.n567 1.0005
R1243 VDDA.n567 VDDA.n565 1.0005
R1244 VDDA.n565 VDDA.n563 1.0005
R1245 VDDA.n563 VDDA.n561 1.0005
R1246 VDDA.n561 VDDA.n543 1.0005
R1247 VDDA.n601 VDDA.n543 1.0005
R1248 VDDA.n523 VDDA.n515 0.938
R1249 VDDA.n449 VDDA.n423 0.78175
R1250 VDDA.n522 VDDA.n516 0.6255
R1251 VDDA.n514 VDDA.n509 0.6255
R1252 VDDA.n465 VDDA.n464 0.6255
R1253 VDDA.n464 VDDA.n462 0.6255
R1254 VDDA.n456 VDDA.n454 0.6255
R1255 VDDA.n465 VDDA.n454 0.6255
R1256 VDDA.n384 VDDA.n383 0.6255
R1257 VDDA.n383 VDDA.n381 0.6255
R1258 VDDA.n375 VDDA.n373 0.6255
R1259 VDDA.n384 VDDA.n373 0.6255
R1260 VDDA.n291 VDDA.n289 0.6255
R1261 VDDA.n289 VDDA.n287 0.6255
R1262 VDDA.n287 VDDA.n285 0.6255
R1263 VDDA.n285 VDDA.n283 0.6255
R1264 VDDA.n283 VDDA.n281 0.6255
R1265 VDDA.n281 VDDA.n279 0.6255
R1266 VDDA.n279 VDDA.n277 0.6255
R1267 VDDA.n277 VDDA.n272 0.6255
R1268 VDDA.n299 VDDA.n272 0.6255
R1269 VDDA.n300 VDDA.n270 0.6255
R1270 VDDA.n270 VDDA.n268 0.6255
R1271 VDDA.n268 VDDA.n266 0.6255
R1272 VDDA.n266 VDDA.n264 0.6255
R1273 VDDA.n264 VDDA.n262 0.6255
R1274 VDDA.n262 VDDA.n260 0.6255
R1275 VDDA.n260 VDDA.n258 0.6255
R1276 VDDA.n258 VDDA.n256 0.6255
R1277 VDDA.n256 VDDA.n252 0.6255
R1278 VDDA.n306 VDDA.n252 0.6255
R1279 VDDA.n331 VDDA.n329 0.563
R1280 VDDA.n336 VDDA.n329 0.563
R1281 VDDA.n358 VDDA.n357 0.563
R1282 VDDA.n357 VDDA.n355 0.563
R1283 VDDA.n355 VDDA.n353 0.563
R1284 VDDA.n340 VDDA.n338 0.563
R1285 VDDA.n345 VDDA.n338 0.563
R1286 VDDA.n348 VDDA.n347 0.563
R1287 VDDA.n347 VDDA.n327 0.563
R1288 VDDA.n358 VDDA.n327 0.563
R1289 VDDA.n499 VDDA.n497 0.563
R1290 VDDA.n497 VDDA.n495 0.563
R1291 VDDA.n495 VDDA.n493 0.563
R1292 VDDA.n493 VDDA.n491 0.563
R1293 VDDA.n504 VDDA.n491 0.563
R1294 VDDA.n471 VDDA.n469 0.563
R1295 VDDA.n473 VDDA.n471 0.563
R1296 VDDA.n475 VDDA.n473 0.563
R1297 VDDA.n477 VDDA.n475 0.563
R1298 VDDA.n443 VDDA.n441 0.563
R1299 VDDA.n441 VDDA.n439 0.563
R1300 VDDA.n439 VDDA.n437 0.563
R1301 VDDA.n437 VDDA.n435 0.563
R1302 VDDA.n435 VDDA.n433 0.563
R1303 VDDA.n433 VDDA.n431 0.563
R1304 VDDA.n431 VDDA.n429 0.563
R1305 VDDA.n429 VDDA.n427 0.563
R1306 VDDA.n427 VDDA.n425 0.563
R1307 VDDA.n448 VDDA.n425 0.563
R1308 VDDA.n418 VDDA.n416 0.563
R1309 VDDA.n416 VDDA.n414 0.563
R1310 VDDA.n414 VDDA.n412 0.563
R1311 VDDA.n412 VDDA.n410 0.563
R1312 VDDA.n423 VDDA.n410 0.563
R1313 VDDA.n390 VDDA.n388 0.563
R1314 VDDA.n392 VDDA.n390 0.563
R1315 VDDA.n394 VDDA.n392 0.563
R1316 VDDA.n396 VDDA.n394 0.563
R1317 VDDA.n602 VDDA.n541 0.5005
R1318 VDDA.n652 VDDA.n638 0.482838
R1319 VDDA.n6 VDDA.n5 0.3295
R1320 VDDA.n7 VDDA.n6 0.3295
R1321 VDDA.n8 VDDA.n7 0.3295
R1322 VDDA.n13 VDDA.n8 0.3295
R1323 VDDA.n13 VDDA.n12 0.3295
R1324 VDDA.n12 VDDA.n11 0.3295
R1325 VDDA.n11 VDDA.n10 0.3295
R1326 VDDA.n10 VDDA.n9 0.3295
R1327 VDDA.n15 VDDA.n14 0.3295
R1328 VDDA.n16 VDDA.n15 0.3295
R1329 VDDA.n17 VDDA.n16 0.3295
R1330 VDDA.n22 VDDA.n17 0.3295
R1331 VDDA.n22 VDDA.n21 0.3295
R1332 VDDA.n21 VDDA.n20 0.3295
R1333 VDDA.n20 VDDA.n19 0.3295
R1334 VDDA.n19 VDDA.n18 0.3295
R1335 VDDA.n24 VDDA.n23 0.3295
R1336 VDDA.n25 VDDA.n24 0.3295
R1337 VDDA.n26 VDDA.n25 0.3295
R1338 VDDA.n31 VDDA.n26 0.3295
R1339 VDDA.n31 VDDA.n30 0.3295
R1340 VDDA.n30 VDDA.n29 0.3295
R1341 VDDA.n29 VDDA.n28 0.3295
R1342 VDDA.n28 VDDA.n27 0.3295
R1343 VDDA.n33 VDDA.n32 0.3295
R1344 VDDA.n34 VDDA.n33 0.3295
R1345 VDDA.n35 VDDA.n34 0.3295
R1346 VDDA.n40 VDDA.n35 0.3295
R1347 VDDA.n40 VDDA.n39 0.3295
R1348 VDDA.n39 VDDA.n38 0.3295
R1349 VDDA.n38 VDDA.n37 0.3295
R1350 VDDA.n37 VDDA.n36 0.3295
R1351 VDDA.n42 VDDA.n41 0.3295
R1352 VDDA.n43 VDDA.n42 0.3295
R1353 VDDA.n44 VDDA.n43 0.3295
R1354 VDDA.n49 VDDA.n44 0.3295
R1355 VDDA.n49 VDDA.n48 0.3295
R1356 VDDA.n48 VDDA.n47 0.3295
R1357 VDDA.n47 VDDA.n46 0.3295
R1358 VDDA.n46 VDDA.n45 0.3295
R1359 VDDA.n51 VDDA.n50 0.3295
R1360 VDDA.n52 VDDA.n51 0.3295
R1361 VDDA.n53 VDDA.n52 0.3295
R1362 VDDA.n58 VDDA.n53 0.3295
R1363 VDDA.n58 VDDA.n57 0.3295
R1364 VDDA.n57 VDDA.n56 0.3295
R1365 VDDA.n56 VDDA.n55 0.3295
R1366 VDDA.n55 VDDA.n54 0.3295
R1367 VDDA.n60 VDDA.n59 0.3295
R1368 VDDA.n61 VDDA.n60 0.3295
R1369 VDDA.n62 VDDA.n61 0.3295
R1370 VDDA.n67 VDDA.n62 0.3295
R1371 VDDA.n67 VDDA.n66 0.3295
R1372 VDDA.n66 VDDA.n65 0.3295
R1373 VDDA.n65 VDDA.n64 0.3295
R1374 VDDA.n64 VDDA.n63 0.3295
R1375 VDDA.n69 VDDA.n68 0.3295
R1376 VDDA.n70 VDDA.n69 0.3295
R1377 VDDA.n71 VDDA.n70 0.3295
R1378 VDDA.n76 VDDA.n71 0.3295
R1379 VDDA.n76 VDDA.n75 0.3295
R1380 VDDA.n75 VDDA.n74 0.3295
R1381 VDDA.n74 VDDA.n73 0.3295
R1382 VDDA.n73 VDDA.n72 0.3295
R1383 VDDA.n78 VDDA.n77 0.3295
R1384 VDDA.n79 VDDA.n78 0.3295
R1385 VDDA.n80 VDDA.n79 0.3295
R1386 VDDA.n85 VDDA.n80 0.3295
R1387 VDDA.n85 VDDA.n84 0.3295
R1388 VDDA.n84 VDDA.n83 0.3295
R1389 VDDA.n83 VDDA.n82 0.3295
R1390 VDDA.n82 VDDA.n81 0.3295
R1391 VDDA.n87 VDDA.n86 0.3295
R1392 VDDA.n88 VDDA.n87 0.3295
R1393 VDDA.n89 VDDA.n88 0.3295
R1394 VDDA.n94 VDDA.n89 0.3295
R1395 VDDA.n94 VDDA.n93 0.3295
R1396 VDDA.n93 VDDA.n92 0.3295
R1397 VDDA.n92 VDDA.n91 0.3295
R1398 VDDA.n91 VDDA.n90 0.3295
R1399 VDDA.n96 VDDA.n95 0.3295
R1400 VDDA.n97 VDDA.n96 0.3295
R1401 VDDA.n98 VDDA.n97 0.3295
R1402 VDDA.n103 VDDA.n98 0.3295
R1403 VDDA.n103 VDDA.n102 0.3295
R1404 VDDA.n102 VDDA.n101 0.3295
R1405 VDDA.n101 VDDA.n100 0.3295
R1406 VDDA.n100 VDDA.n99 0.3295
R1407 VDDA.n105 VDDA.n104 0.3295
R1408 VDDA.n106 VDDA.n105 0.3295
R1409 VDDA.n107 VDDA.n106 0.3295
R1410 VDDA.n112 VDDA.n107 0.3295
R1411 VDDA.n112 VDDA.n111 0.3295
R1412 VDDA.n111 VDDA.n110 0.3295
R1413 VDDA.n110 VDDA.n109 0.3295
R1414 VDDA.n109 VDDA.n108 0.3295
R1415 VDDA.n114 VDDA.n113 0.3295
R1416 VDDA.n115 VDDA.n114 0.3295
R1417 VDDA.n116 VDDA.n115 0.3295
R1418 VDDA.n121 VDDA.n116 0.3295
R1419 VDDA.n121 VDDA.n120 0.3295
R1420 VDDA.n120 VDDA.n119 0.3295
R1421 VDDA.n119 VDDA.n118 0.3295
R1422 VDDA.n118 VDDA.n117 0.3295
R1423 VDDA.n123 VDDA.n122 0.3295
R1424 VDDA.n124 VDDA.n123 0.3295
R1425 VDDA.n125 VDDA.n124 0.3295
R1426 VDDA.n130 VDDA.n125 0.3295
R1427 VDDA.n130 VDDA.n129 0.3295
R1428 VDDA.n129 VDDA.n128 0.3295
R1429 VDDA.n128 VDDA.n127 0.3295
R1430 VDDA.n127 VDDA.n126 0.3295
R1431 VDDA.n132 VDDA.n131 0.3295
R1432 VDDA.n133 VDDA.n132 0.3295
R1433 VDDA.n134 VDDA.n133 0.3295
R1434 VDDA.n139 VDDA.n134 0.3295
R1435 VDDA.n139 VDDA.n138 0.3295
R1436 VDDA.n138 VDDA.n137 0.3295
R1437 VDDA.n137 VDDA.n136 0.3295
R1438 VDDA.n136 VDDA.n135 0.3295
R1439 VDDA.n141 VDDA.n140 0.3295
R1440 VDDA.n142 VDDA.n141 0.3295
R1441 VDDA.n143 VDDA.n142 0.3295
R1442 VDDA.n148 VDDA.n143 0.3295
R1443 VDDA.n148 VDDA.n147 0.3295
R1444 VDDA.n147 VDDA.n146 0.3295
R1445 VDDA.n146 VDDA.n145 0.3295
R1446 VDDA.n145 VDDA.n144 0.3295
R1447 VDDA.n150 VDDA.n149 0.3295
R1448 VDDA.n151 VDDA.n150 0.3295
R1449 VDDA.n152 VDDA.n151 0.3295
R1450 VDDA.n157 VDDA.n152 0.3295
R1451 VDDA.n157 VDDA.n156 0.3295
R1452 VDDA.n156 VDDA.n155 0.3295
R1453 VDDA.n155 VDDA.n154 0.3295
R1454 VDDA.n154 VDDA.n153 0.3295
R1455 VDDA.n159 VDDA.n158 0.3295
R1456 VDDA.n160 VDDA.n159 0.3295
R1457 VDDA.n161 VDDA.n160 0.3295
R1458 VDDA.n166 VDDA.n161 0.3295
R1459 VDDA.n166 VDDA.n165 0.3295
R1460 VDDA.n165 VDDA.n164 0.3295
R1461 VDDA.n164 VDDA.n163 0.3295
R1462 VDDA.n163 VDDA.n162 0.3295
R1463 VDDA.n168 VDDA.n167 0.3295
R1464 VDDA.n169 VDDA.n168 0.3295
R1465 VDDA.n170 VDDA.n169 0.3295
R1466 VDDA.n175 VDDA.n170 0.3295
R1467 VDDA.n175 VDDA.n174 0.3295
R1468 VDDA.n174 VDDA.n173 0.3295
R1469 VDDA.n173 VDDA.n172 0.3295
R1470 VDDA.n172 VDDA.n171 0.3295
R1471 VDDA.n177 VDDA.n176 0.3295
R1472 VDDA.n178 VDDA.n177 0.3295
R1473 VDDA.n179 VDDA.n178 0.3295
R1474 VDDA.n184 VDDA.n179 0.3295
R1475 VDDA.n184 VDDA.n183 0.3295
R1476 VDDA.n183 VDDA.n182 0.3295
R1477 VDDA.n182 VDDA.n181 0.3295
R1478 VDDA.n181 VDDA.n180 0.3295
R1479 VDDA.n186 VDDA.n185 0.3295
R1480 VDDA.n187 VDDA.n186 0.3295
R1481 VDDA.n188 VDDA.n187 0.3295
R1482 VDDA.n193 VDDA.n188 0.3295
R1483 VDDA.n193 VDDA.n192 0.3295
R1484 VDDA.n192 VDDA.n191 0.3295
R1485 VDDA.n191 VDDA.n190 0.3295
R1486 VDDA.n190 VDDA.n189 0.3295
R1487 VDDA.n195 VDDA.n194 0.3295
R1488 VDDA.n196 VDDA.n195 0.3295
R1489 VDDA.n197 VDDA.n196 0.3295
R1490 VDDA.n202 VDDA.n197 0.3295
R1491 VDDA.n202 VDDA.n201 0.3295
R1492 VDDA.n201 VDDA.n200 0.3295
R1493 VDDA.n200 VDDA.n199 0.3295
R1494 VDDA.n199 VDDA.n198 0.3295
R1495 VDDA.n204 VDDA.n203 0.3295
R1496 VDDA.n205 VDDA.n204 0.3295
R1497 VDDA.n206 VDDA.n205 0.3295
R1498 VDDA.n211 VDDA.n206 0.3295
R1499 VDDA.n211 VDDA.n210 0.3295
R1500 VDDA.n210 VDDA.n209 0.3295
R1501 VDDA.n209 VDDA.n208 0.3295
R1502 VDDA.n208 VDDA.n207 0.3295
R1503 VDDA.n213 VDDA.n212 0.3295
R1504 VDDA.n214 VDDA.n213 0.3295
R1505 VDDA.n215 VDDA.n214 0.3295
R1506 VDDA.n216 VDDA.n215 0.3295
R1507 VDDA.n217 VDDA.n216 0.3295
R1508 VDDA.n218 VDDA.n217 0.3295
R1509 VDDA.n219 VDDA.n218 0.3295
R1510 VDDA.n220 VDDA.n219 0.3295
R1511 VDDA.n221 VDDA.n220 0.3295
R1512 VDDA.n243 VDDA.n221 0.318925
R1513 VDDA.n22 VDDA.n13 0.2825
R1514 VDDA.n31 VDDA.n22 0.2825
R1515 VDDA.n40 VDDA.n31 0.2825
R1516 VDDA.n49 VDDA.n40 0.2825
R1517 VDDA.n58 VDDA.n49 0.2825
R1518 VDDA.n67 VDDA.n58 0.2825
R1519 VDDA.n76 VDDA.n67 0.2825
R1520 VDDA.n85 VDDA.n76 0.2825
R1521 VDDA.n94 VDDA.n85 0.2825
R1522 VDDA.n103 VDDA.n94 0.2825
R1523 VDDA.n112 VDDA.n103 0.2825
R1524 VDDA.n121 VDDA.n112 0.2825
R1525 VDDA.n130 VDDA.n121 0.2825
R1526 VDDA.n139 VDDA.n130 0.2825
R1527 VDDA.n148 VDDA.n139 0.2825
R1528 VDDA.n157 VDDA.n148 0.2825
R1529 VDDA.n166 VDDA.n157 0.2825
R1530 VDDA.n175 VDDA.n166 0.2825
R1531 VDDA.n184 VDDA.n175 0.2825
R1532 VDDA.n193 VDDA.n184 0.2825
R1533 VDDA.n202 VDDA.n193 0.2825
R1534 VDDA.n211 VDDA.n202 0.2825
R1535 VDDA.n216 VDDA.n211 0.2825
R1536 VDDA.n527 VDDA.n318 0.215525
R1537 VDDA.n362 VDDA.n324 0.1755
R1538 VDDA.n369 VDDA.n324 0.1755
R1539 VDDA.n370 VDDA.n369 0.1755
R1540 VDDA.n365 VDDA.n364 0.1755
R1541 VDDA.n368 VDDA.n365 0.1755
R1542 VDDA.n368 VDDA.n323 0.1755
R1543 VDDA.n362 VDDA.n361 0.163
R1544 VDDA.n524 VDDA.n370 0.163
R1545 VDDA.n364 VDDA.n325 0.163
R1546 VDDA.n525 VDDA.n323 0.163
R1547 VDDA.t146 VDDA.t53 0.1603
R1548 VDDA.t29 VDDA.t427 0.1603
R1549 VDDA.t434 VDDA.t133 0.1603
R1550 VDDA.t95 VDDA.t428 0.1603
R1551 VDDA.t435 VDDA.t56 0.1603
R1552 VDDA.n623 VDDA.t132 0.159278
R1553 VDDA.n624 VDDA.t429 0.159278
R1554 VDDA.n625 VDDA.t58 0.159278
R1555 VDDA.n626 VDDA.t218 0.159278
R1556 VDDA.n604 VDDA.n533 0.146333
R1557 VDDA.n611 VDDA.n533 0.146333
R1558 VDDA.n607 VDDA.n606 0.146333
R1559 VDDA.n610 VDDA.n607 0.146333
R1560 VDDA.n610 VDDA.n532 0.146333
R1561 VDDA.n628 VDDA.n620 0.146333
R1562 VDDA.n635 VDDA.n620 0.146333
R1563 VDDA.n631 VDDA.n630 0.146333
R1564 VDDA.n634 VDDA.n631 0.146333
R1565 VDDA.n634 VDDA.n619 0.146333
R1566 VDDA.n233 VDDA.n227 0.146333
R1567 VDDA.n240 VDDA.n227 0.146333
R1568 VDDA.n236 VDDA.n235 0.146333
R1569 VDDA.n239 VDDA.n236 0.146333
R1570 VDDA.n239 VDDA.n226 0.146333
R1571 VDDA.n308 VDDA.n249 0.146333
R1572 VDDA.n315 VDDA.n249 0.146333
R1573 VDDA.n311 VDDA.n310 0.146333
R1574 VDDA.n314 VDDA.n311 0.146333
R1575 VDDA.n314 VDDA.n248 0.146333
R1576 VDDA.n614 VDDA.n527 0.145025
R1577 VDDA.n626 VDDA.t57 0.1368
R1578 VDDA.n626 VDDA.t146 0.1368
R1579 VDDA.n625 VDDA.t36 0.1368
R1580 VDDA.n625 VDDA.t29 0.1368
R1581 VDDA.n624 VDDA.t141 0.1368
R1582 VDDA.n624 VDDA.t434 0.1368
R1583 VDDA.n623 VDDA.t37 0.1368
R1584 VDDA.n623 VDDA.t95 0.1368
R1585 VDDA.n622 VDDA.t430 0.1368
R1586 VDDA.n622 VDDA.t435 0.1368
R1587 VDDA.n604 VDDA.n603 0.135917
R1588 VDDA.n606 VDDA.n534 0.135917
R1589 VDDA.n628 VDDA.n627 0.135917
R1590 VDDA.n630 VDDA.n621 0.135917
R1591 VDDA.n233 VDDA.n232 0.135917
R1592 VDDA.n235 VDDA.n228 0.135917
R1593 VDDA.n308 VDDA.n307 0.135917
R1594 VDDA.n310 VDDA.n250 0.135917
R1595 VDDA.n638 VDDA.n614 0.100963
R1596 VDDA VDDA.n653 0.0806938
R1597 VDDA.n612 VDDA.n532 0.0667303
R1598 VDDA.n636 VDDA.n619 0.0667303
R1599 VDDA.n241 VDDA.n226 0.0667303
R1600 VDDA.n316 VDDA.n248 0.0667303
R1601 VDDA.n367 VDDA.n366 0.0663
R1602 VDDA.n363 VDDA.n319 0.0616
R1603 VDDA.n526 VDDA.n322 0.0616
R1604 VDDA.n609 VDDA.n608 0.0553333
R1605 VDDA.n633 VDDA.n632 0.0553333
R1606 VDDA.n238 VDDA.n237 0.0553333
R1607 VDDA.n313 VDDA.n312 0.0553333
R1608 VDDA.n605 VDDA.n528 0.0514167
R1609 VDDA.n613 VDDA.n531 0.0514167
R1610 VDDA.n629 VDDA.n615 0.0514167
R1611 VDDA.n637 VDDA.n618 0.0514167
R1612 VDDA.n234 VDDA.n222 0.0514167
R1613 VDDA.n242 VDDA.n225 0.0514167
R1614 VDDA.n309 VDDA.n244 0.0514167
R1615 VDDA.n317 VDDA.n247 0.0514167
R1616 VDDA.n318 VDDA.n243 0.034575
R1617 VDDA.n366 VDDA.n320 0.0335856
R1618 VDDA.n322 VDDA.n321 0.0335856
R1619 VDDA.n367 VDDA.n321 0.0335856
R1620 VDDA.n363 VDDA.n320 0.0335856
R1621 VDDA.n608 VDDA.n529 0.028198
R1622 VDDA.n531 VDDA.n530 0.028198
R1623 VDDA.n632 VDDA.n616 0.028198
R1624 VDDA.n618 VDDA.n617 0.028198
R1625 VDDA.n237 VDDA.n223 0.028198
R1626 VDDA.n225 VDDA.n224 0.028198
R1627 VDDA.n312 VDDA.n245 0.028198
R1628 VDDA.n247 VDDA.n246 0.028198
R1629 VDDA.n313 VDDA.n246 0.028198
R1630 VDDA.n309 VDDA.n245 0.028198
R1631 VDDA.n238 VDDA.n224 0.028198
R1632 VDDA.n234 VDDA.n223 0.028198
R1633 VDDA.n633 VDDA.n617 0.028198
R1634 VDDA.n629 VDDA.n616 0.028198
R1635 VDDA.n609 VDDA.n530 0.028198
R1636 VDDA.n605 VDDA.n529 0.028198
R1637 VDDA.n652 VDDA.n640 0.0116625
R1638 VDDA.n640 VDDA.n4 0.0116625
R1639 VDDA.n645 VDDA.n644 0.0068649
R1640 VDDA.n645 VDDA.n1 0.0068649
R1641 VDDA.n649 VDDA.n646 0.0068649
R1642 VDDA.n650 VDDA.n1 0.0068649
R1643 VDDA.n650 VDDA.n649 0.0068649
R1644 VDDA.n644 VDDA.n4 0.0068649
R1645 VDDA.n646 VDDA.n2 0.00657213
R1646 VDDA.n648 VDDA.n3 0.00657213
R1647 VDDA.n647 VDDA.n2 0.00657213
R1648 VDDA.n648 VDDA.n647 0.00657213
R1649 VDDA.n641 VDDA.n639 0.00393497
R1650 VDDA.n642 VDDA.n641 0.00393497
R1651 VDDA.n642 VDDA.n0 0.0036417
R1652 VDDA.n651 VDDA.n643 0.0036417
R1653 VDDA.n653 VDDA.n0 0.0036417
R1654 VDDA.n643 VDDA.n639 0.0036417
R1655 VDDA.t132 VDDA.n622 0.00152174
R1656 VDDA.t429 VDDA.n623 0.00152174
R1657 VDDA.t58 VDDA.n624 0.00152174
R1658 VDDA.t218 VDDA.n625 0.00152174
R1659 VDDA.t237 VDDA.n626 0.00152174
R1660 VOUT+.n9 VOUT+.t17 113.192
R1661 VOUT+.n11 VOUT+.n10 34.9935
R1662 VOUT+.n13 VOUT+.n12 34.9935
R1663 VOUT+.n17 VOUT+.n16 34.9935
R1664 VOUT+.n20 VOUT+.n19 34.9935
R1665 VOUT+.n23 VOUT+.n22 34.9935
R1666 VOUT+.n27 VOUT+.n26 34.9935
R1667 VOUT+.n110 VOUT+.n30 20.5005
R1668 VOUT+.n110 VOUT+.n109 11.6871
R1669 VOUT+.n2 VOUT+.n1 9.73997
R1670 VOUT+.n4 VOUT+.n3 9.73997
R1671 VOUT+.n7 VOUT+.n6 9.73997
R1672 VOUT+ VOUT+.n110 9.34425
R1673 VOUT+.n7 VOUT+.n5 7.14633
R1674 VOUT+.n5 VOUT+.n2 7.14633
R1675 VOUT+.n2 VOUT+.n0 7.14633
R1676 VOUT+.n10 VOUT+.t5 6.56717
R1677 VOUT+.n10 VOUT+.t10 6.56717
R1678 VOUT+.n12 VOUT+.t13 6.56717
R1679 VOUT+.n12 VOUT+.t11 6.56717
R1680 VOUT+.n16 VOUT+.t4 6.56717
R1681 VOUT+.n16 VOUT+.t14 6.56717
R1682 VOUT+.n19 VOUT+.t6 6.56717
R1683 VOUT+.n19 VOUT+.t9 6.56717
R1684 VOUT+.n22 VOUT+.t7 6.56717
R1685 VOUT+.n22 VOUT+.t12 6.56717
R1686 VOUT+.n26 VOUT+.t8 6.56717
R1687 VOUT+.n26 VOUT+.t3 6.56717
R1688 VOUT+.n21 VOUT+.n17 6.3755
R1689 VOUT+.n18 VOUT+.n17 6.3755
R1690 VOUT+.n29 VOUT+.n13 6.3755
R1691 VOUT+.n15 VOUT+.n13 6.3755
R1692 VOUT+.n4 VOUT+.n0 6.02133
R1693 VOUT+.n5 VOUT+.n4 6.02133
R1694 VOUT+.n8 VOUT+.n7 6.02133
R1695 VOUT+.n20 VOUT+.n18 5.813
R1696 VOUT+.n21 VOUT+.n20 5.813
R1697 VOUT+.n23 VOUT+.n14 5.813
R1698 VOUT+.n24 VOUT+.n23 5.813
R1699 VOUT+.n28 VOUT+.n27 5.813
R1700 VOUT+.n27 VOUT+.n25 5.813
R1701 VOUT+.n15 VOUT+.n11 5.813
R1702 VOUT+.n57 VOUT+.t66 4.8295
R1703 VOUT+.n59 VOUT+.t137 4.8295
R1704 VOUT+.n61 VOUT+.t27 4.8295
R1705 VOUT+.n63 VOUT+.t81 4.8295
R1706 VOUT+.n65 VOUT+.t114 4.8295
R1707 VOUT+.n77 VOUT+.t105 4.8295
R1708 VOUT+.n79 VOUT+.t48 4.8295
R1709 VOUT+.n80 VOUT+.t62 4.8295
R1710 VOUT+.n82 VOUT+.t139 4.8295
R1711 VOUT+.n83 VOUT+.t26 4.8295
R1712 VOUT+.n85 VOUT+.t104 4.8295
R1713 VOUT+.n86 VOUT+.t129 4.8295
R1714 VOUT+.n88 VOUT+.t135 4.8295
R1715 VOUT+.n89 VOUT+.t23 4.8295
R1716 VOUT+.n91 VOUT+.t97 4.8295
R1717 VOUT+.n92 VOUT+.t123 4.8295
R1718 VOUT+.n94 VOUT+.t57 4.8295
R1719 VOUT+.n95 VOUT+.t85 4.8295
R1720 VOUT+.n97 VOUT+.t89 4.8295
R1721 VOUT+.n98 VOUT+.t118 4.8295
R1722 VOUT+.n100 VOUT+.t52 4.8295
R1723 VOUT+.n101 VOUT+.t80 4.8295
R1724 VOUT+.n103 VOUT+.t151 4.8295
R1725 VOUT+.n104 VOUT+.t41 4.8295
R1726 VOUT+.n31 VOUT+.t35 4.8295
R1727 VOUT+.n43 VOUT+.t58 4.8295
R1728 VOUT+.n45 VOUT+.t103 4.8295
R1729 VOUT+.n46 VOUT+.t130 4.8295
R1730 VOUT+.n48 VOUT+.t67 4.8295
R1731 VOUT+.n49 VOUT+.t98 4.8295
R1732 VOUT+.n51 VOUT+.t109 4.8295
R1733 VOUT+.n52 VOUT+.t136 4.8295
R1734 VOUT+.n54 VOUT+.t145 4.8295
R1735 VOUT+.n55 VOUT+.t32 4.8295
R1736 VOUT+.n106 VOUT+.t74 4.8295
R1737 VOUT+.n70 VOUT+.t37 4.8154
R1738 VOUT+.n69 VOUT+.t76 4.8154
R1739 VOUT+.n68 VOUT+.t56 4.8154
R1740 VOUT+.n67 VOUT+.t91 4.8154
R1741 VOUT+.n76 VOUT+.t75 4.806
R1742 VOUT+.n75 VOUT+.t53 4.806
R1743 VOUT+.n74 VOUT+.t90 4.806
R1744 VOUT+.n73 VOUT+.t126 4.806
R1745 VOUT+.n72 VOUT+.t110 4.806
R1746 VOUT+.n71 VOUT+.t148 4.806
R1747 VOUT+.n70 VOUT+.t44 4.806
R1748 VOUT+.n69 VOUT+.t82 4.806
R1749 VOUT+.n68 VOUT+.t61 4.806
R1750 VOUT+.n67 VOUT+.t100 4.806
R1751 VOUT+.n42 VOUT+.t99 4.806
R1752 VOUT+.n41 VOUT+.t149 4.806
R1753 VOUT+.n40 VOUT+.t43 4.806
R1754 VOUT+.n39 VOUT+.t77 4.806
R1755 VOUT+.n38 VOUT+.t125 4.806
R1756 VOUT+.n37 VOUT+.t20 4.806
R1757 VOUT+.n36 VOUT+.t59 4.806
R1758 VOUT+.n35 VOUT+.t92 4.806
R1759 VOUT+.n34 VOUT+.t143 4.806
R1760 VOUT+.n33 VOUT+.t39 4.806
R1761 VOUT+.n58 VOUT+.t36 4.5005
R1762 VOUT+.n57 VOUT+.t28 4.5005
R1763 VOUT+.n59 VOUT+.t33 4.5005
R1764 VOUT+.n60 VOUT+.t86 4.5005
R1765 VOUT+.n61 VOUT+.t69 4.5005
R1766 VOUT+.n62 VOUT+.t122 4.5005
R1767 VOUT+.n63 VOUT+.t119 4.5005
R1768 VOUT+.n64 VOUT+.t106 4.5005
R1769 VOUT+.n65 VOUT+.t156 4.5005
R1770 VOUT+.n66 VOUT+.t140 4.5005
R1771 VOUT+.n67 VOUT+.t131 4.5005
R1772 VOUT+.n68 VOUT+.t94 4.5005
R1773 VOUT+.n69 VOUT+.t115 4.5005
R1774 VOUT+.n70 VOUT+.t78 4.5005
R1775 VOUT+.n71 VOUT+.t42 4.5005
R1776 VOUT+.n72 VOUT+.t141 4.5005
R1777 VOUT+.n73 VOUT+.t22 4.5005
R1778 VOUT+.n74 VOUT+.t124 4.5005
R1779 VOUT+.n75 VOUT+.t87 4.5005
R1780 VOUT+.n76 VOUT+.t112 4.5005
R1781 VOUT+.n78 VOUT+.t71 4.5005
R1782 VOUT+.n77 VOUT+.t68 4.5005
R1783 VOUT+.n79 VOUT+.t70 4.5005
R1784 VOUT+.n81 VOUT+.t29 4.5005
R1785 VOUT+.n80 VOUT+.t24 4.5005
R1786 VOUT+.n82 VOUT+.t88 4.5005
R1787 VOUT+.n84 VOUT+.t54 4.5005
R1788 VOUT+.n83 VOUT+.t25 4.5005
R1789 VOUT+.n85 VOUT+.t51 4.5005
R1790 VOUT+.n87 VOUT+.t154 4.5005
R1791 VOUT+.n86 VOUT+.t128 4.5005
R1792 VOUT+.n88 VOUT+.t83 4.5005
R1793 VOUT+.n90 VOUT+.t50 4.5005
R1794 VOUT+.n89 VOUT+.t21 4.5005
R1795 VOUT+.n91 VOUT+.t46 4.5005
R1796 VOUT+.n93 VOUT+.t150 4.5005
R1797 VOUT+.n92 VOUT+.t121 4.5005
R1798 VOUT+.n94 VOUT+.t144 4.5005
R1799 VOUT+.n96 VOUT+.t111 4.5005
R1800 VOUT+.n95 VOUT+.t84 4.5005
R1801 VOUT+.n97 VOUT+.t38 4.5005
R1802 VOUT+.n99 VOUT+.t142 4.5005
R1803 VOUT+.n98 VOUT+.t117 4.5005
R1804 VOUT+.n100 VOUT+.t138 4.5005
R1805 VOUT+.n102 VOUT+.t108 4.5005
R1806 VOUT+.n101 VOUT+.t79 4.5005
R1807 VOUT+.n103 VOUT+.t102 4.5005
R1808 VOUT+.n105 VOUT+.t64 4.5005
R1809 VOUT+.n104 VOUT+.t40 4.5005
R1810 VOUT+.n32 VOUT+.t63 4.5005
R1811 VOUT+.n31 VOUT+.t34 4.5005
R1812 VOUT+.n33 VOUT+.t95 4.5005
R1813 VOUT+.n34 VOUT+.t146 4.5005
R1814 VOUT+.n35 VOUT+.t107 4.5005
R1815 VOUT+.n36 VOUT+.t153 4.5005
R1816 VOUT+.n37 VOUT+.t65 4.5005
R1817 VOUT+.n38 VOUT+.t113 4.5005
R1818 VOUT+.n39 VOUT+.t72 4.5005
R1819 VOUT+.n40 VOUT+.t120 4.5005
R1820 VOUT+.n41 VOUT+.t31 4.5005
R1821 VOUT+.n42 VOUT+.t132 4.5005
R1822 VOUT+.n44 VOUT+.t45 4.5005
R1823 VOUT+.n43 VOUT+.t147 4.5005
R1824 VOUT+.n45 VOUT+.t49 4.5005
R1825 VOUT+.n47 VOUT+.t152 4.5005
R1826 VOUT+.n46 VOUT+.t127 4.5005
R1827 VOUT+.n48 VOUT+.t155 4.5005
R1828 VOUT+.n50 VOUT+.t116 4.5005
R1829 VOUT+.n49 VOUT+.t96 4.5005
R1830 VOUT+.n51 VOUT+.t55 4.5005
R1831 VOUT+.n53 VOUT+.t19 4.5005
R1832 VOUT+.n52 VOUT+.t134 4.5005
R1833 VOUT+.n54 VOUT+.t93 4.5005
R1834 VOUT+.n56 VOUT+.t60 4.5005
R1835 VOUT+.n55 VOUT+.t30 4.5005
R1836 VOUT+.n109 VOUT+.t47 4.5005
R1837 VOUT+.n108 VOUT+.t133 4.5005
R1838 VOUT+.n107 VOUT+.t101 4.5005
R1839 VOUT+.n106 VOUT+.t73 4.5005
R1840 VOUT+.n30 VOUT+.n29 4.5005
R1841 VOUT+.n1 VOUT+.t16 3.42907
R1842 VOUT+.n1 VOUT+.t2 3.42907
R1843 VOUT+.n3 VOUT+.t1 3.42907
R1844 VOUT+.n3 VOUT+.t15 3.42907
R1845 VOUT+.n6 VOUT+.t18 3.42907
R1846 VOUT+.n6 VOUT+.t0 3.42907
R1847 VOUT+ VOUT+.n9 1.938
R1848 VOUT+.n9 VOUT+.n8 1.84425
R1849 VOUT+.n30 VOUT+.n11 1.313
R1850 VOUT+.n8 VOUT+.n0 1.1255
R1851 VOUT+.n25 VOUT+.n15 0.563
R1852 VOUT+.n25 VOUT+.n24 0.563
R1853 VOUT+.n24 VOUT+.n21 0.563
R1854 VOUT+.n18 VOUT+.n14 0.563
R1855 VOUT+.n28 VOUT+.n14 0.563
R1856 VOUT+.n29 VOUT+.n28 0.563
R1857 VOUT+.n58 VOUT+.n57 0.3295
R1858 VOUT+.n60 VOUT+.n59 0.3295
R1859 VOUT+.n62 VOUT+.n61 0.3295
R1860 VOUT+.n64 VOUT+.n63 0.3295
R1861 VOUT+.n66 VOUT+.n65 0.3295
R1862 VOUT+.n68 VOUT+.n67 0.3295
R1863 VOUT+.n69 VOUT+.n68 0.3295
R1864 VOUT+.n70 VOUT+.n69 0.3295
R1865 VOUT+.n71 VOUT+.n70 0.3295
R1866 VOUT+.n72 VOUT+.n71 0.3295
R1867 VOUT+.n73 VOUT+.n72 0.3295
R1868 VOUT+.n74 VOUT+.n73 0.3295
R1869 VOUT+.n75 VOUT+.n74 0.3295
R1870 VOUT+.n76 VOUT+.n75 0.3295
R1871 VOUT+.n78 VOUT+.n76 0.3295
R1872 VOUT+.n78 VOUT+.n77 0.3295
R1873 VOUT+.n81 VOUT+.n79 0.3295
R1874 VOUT+.n81 VOUT+.n80 0.3295
R1875 VOUT+.n84 VOUT+.n82 0.3295
R1876 VOUT+.n84 VOUT+.n83 0.3295
R1877 VOUT+.n87 VOUT+.n85 0.3295
R1878 VOUT+.n87 VOUT+.n86 0.3295
R1879 VOUT+.n90 VOUT+.n88 0.3295
R1880 VOUT+.n90 VOUT+.n89 0.3295
R1881 VOUT+.n93 VOUT+.n91 0.3295
R1882 VOUT+.n93 VOUT+.n92 0.3295
R1883 VOUT+.n96 VOUT+.n94 0.3295
R1884 VOUT+.n96 VOUT+.n95 0.3295
R1885 VOUT+.n99 VOUT+.n97 0.3295
R1886 VOUT+.n99 VOUT+.n98 0.3295
R1887 VOUT+.n102 VOUT+.n100 0.3295
R1888 VOUT+.n102 VOUT+.n101 0.3295
R1889 VOUT+.n105 VOUT+.n103 0.3295
R1890 VOUT+.n105 VOUT+.n104 0.3295
R1891 VOUT+.n32 VOUT+.n31 0.3295
R1892 VOUT+.n34 VOUT+.n33 0.3295
R1893 VOUT+.n35 VOUT+.n34 0.3295
R1894 VOUT+.n36 VOUT+.n35 0.3295
R1895 VOUT+.n37 VOUT+.n36 0.3295
R1896 VOUT+.n38 VOUT+.n37 0.3295
R1897 VOUT+.n39 VOUT+.n38 0.3295
R1898 VOUT+.n40 VOUT+.n39 0.3295
R1899 VOUT+.n41 VOUT+.n40 0.3295
R1900 VOUT+.n42 VOUT+.n41 0.3295
R1901 VOUT+.n44 VOUT+.n42 0.3295
R1902 VOUT+.n44 VOUT+.n43 0.3295
R1903 VOUT+.n47 VOUT+.n45 0.3295
R1904 VOUT+.n47 VOUT+.n46 0.3295
R1905 VOUT+.n50 VOUT+.n48 0.3295
R1906 VOUT+.n50 VOUT+.n49 0.3295
R1907 VOUT+.n53 VOUT+.n51 0.3295
R1908 VOUT+.n53 VOUT+.n52 0.3295
R1909 VOUT+.n56 VOUT+.n54 0.3295
R1910 VOUT+.n56 VOUT+.n55 0.3295
R1911 VOUT+.n109 VOUT+.n108 0.3295
R1912 VOUT+.n108 VOUT+.n107 0.3295
R1913 VOUT+.n107 VOUT+.n106 0.3295
R1914 VOUT+.n74 VOUT+.n60 0.306
R1915 VOUT+.n73 VOUT+.n62 0.306
R1916 VOUT+.n72 VOUT+.n64 0.306
R1917 VOUT+.n71 VOUT+.n66 0.306
R1918 VOUT+.n78 VOUT+.n58 0.2825
R1919 VOUT+.n81 VOUT+.n78 0.2825
R1920 VOUT+.n84 VOUT+.n81 0.2825
R1921 VOUT+.n87 VOUT+.n84 0.2825
R1922 VOUT+.n90 VOUT+.n87 0.2825
R1923 VOUT+.n93 VOUT+.n90 0.2825
R1924 VOUT+.n96 VOUT+.n93 0.2825
R1925 VOUT+.n99 VOUT+.n96 0.2825
R1926 VOUT+.n102 VOUT+.n99 0.2825
R1927 VOUT+.n105 VOUT+.n102 0.2825
R1928 VOUT+.n44 VOUT+.n32 0.2825
R1929 VOUT+.n47 VOUT+.n44 0.2825
R1930 VOUT+.n50 VOUT+.n47 0.2825
R1931 VOUT+.n53 VOUT+.n50 0.2825
R1932 VOUT+.n56 VOUT+.n53 0.2825
R1933 VOUT+.n107 VOUT+.n56 0.2825
R1934 VOUT+.n107 VOUT+.n105 0.2825
R1935 GNDA.n1266 GNDA.n443 580164
R1936 GNDA.n2007 GNDA.n158 289300
R1937 GNDA.n2006 GNDA.n160 162800
R1938 GNDA.n1898 GNDA.n1897 162800
R1939 GNDA.n1898 GNDA.n189 150171
R1940 GNDA.n1287 GNDA.n160 150171
R1941 GNDA.n1294 GNDA.n158 146899
R1942 GNDA.n2007 GNDA.n159 127050
R1943 GNDA.n1897 GNDA.n1896 111525
R1944 GNDA.n2006 GNDA.n2005 111525
R1945 GNDA.n1268 GNDA.n1266 86533.3
R1946 GNDA.n1900 GNDA.n187 58614.3
R1947 GNDA.n1268 GNDA.n1267 19712
R1948 GNDA.n1278 GNDA.n1270 15280.4
R1949 GNDA.n1284 GNDA.n160 14922.8
R1950 GNDA.n1279 GNDA.n189 14221.4
R1951 GNDA.n1283 GNDA.n1282 14173
R1952 GNDA.n1899 GNDA.n1898 14149
R1953 GNDA.n1285 GNDA.n1283 13700
R1954 GNDA.n1290 GNDA.n1289 13528.5
R1955 GNDA.n1278 GNDA.n1269 13062.1
R1956 GNDA.n1899 GNDA.n188 12650
R1957 GNDA.n1295 GNDA.n443 11953.3
R1958 GNDA.n1295 GNDA.n1294 11890.5
R1959 GNDA.n1288 GNDA.n159 11867.9
R1960 GNDA.n1272 GNDA.n1271 11440
R1961 GNDA.n1280 GNDA.n1279 11412.4
R1962 GNDA.n1288 GNDA.n1287 11404.3
R1963 GNDA.n1292 GNDA.n1291 10293.6
R1964 GNDA.n1294 GNDA.n1293 9950.42
R1965 GNDA.n1267 GNDA.n443 9950.42
R1966 GNDA.n1267 GNDA.n444 9384.59
R1967 GNDA.n1293 GNDA.n444 9384.59
R1968 GNDA.n1291 GNDA.n1269 8422.86
R1969 GNDA.n1280 GNDA.n1272 7648.95
R1970 GNDA.n1286 GNDA.n1272 7630.38
R1971 GNDA.n1289 GNDA.n1271 7385.71
R1972 GNDA.n1289 GNDA.n1288 6364.29
R1973 GNDA.n1290 GNDA.n1270 5234.66
R1974 GNDA.t57 GNDA.t583 5225.11
R1975 GNDA.n1281 GNDA.n189 5028.57
R1976 GNDA.n1279 GNDA.n1278 4435.89
R1977 GNDA.n1291 GNDA.n444 3995.79
R1978 GNDA.n1595 GNDA.n1295 3974.19
R1979 GNDA.n2007 GNDA.t110 3588.39
R1980 GNDA.n1286 GNDA.n1285 3498
R1981 GNDA.n1269 GNDA.n1268 3314.67
R1982 GNDA.n1291 GNDA.n1290 3205.71
R1983 GNDA.n1271 GNDA.n1270 2928.92
R1984 GNDA.n1291 GNDA.n159 2704.59
R1985 GNDA.n1285 GNDA.n1284 2520.94
R1986 GNDA.t206 GNDA.n2007 2346.41
R1987 GNDA.n1282 GNDA.n188 2021.46
R1988 GNDA.n1282 GNDA.n1281 1985.64
R1989 GNDA.n1281 GNDA.n1280 1868.49
R1990 GNDA.n1283 GNDA.n1277 1800
R1991 GNDA.n1901 GNDA.n188 1650
R1992 GNDA.n1293 GNDA.n1292 1440.71
R1993 GNDA.n1292 GNDA.n158 1440.71
R1994 GNDA.n1284 GNDA.t535 1426.21
R1995 GNDA.n2068 GNDA.n140 1214.72
R1996 GNDA.n2068 GNDA.n2067 1214.72
R1997 GNDA.n2067 GNDA.n2066 1214.72
R1998 GNDA.n2066 GNDA.n2038 1214.72
R1999 GNDA.n2060 GNDA.n2038 1214.72
R2000 GNDA.n2058 GNDA.n2057 1214.72
R2001 GNDA.n2057 GNDA.n2056 1214.72
R2002 GNDA.n2056 GNDA.n2048 1214.72
R2003 GNDA.n2048 GNDA.n114 1214.72
R2004 GNDA.n2201 GNDA.n114 1214.72
R2005 GNDA.n1214 GNDA.n1213 1214.72
R2006 GNDA.n1213 GNDA.n1212 1214.72
R2007 GNDA.n1212 GNDA.n1181 1214.72
R2008 GNDA.n1206 GNDA.n1181 1214.72
R2009 GNDA.n1206 GNDA.n1205 1214.72
R2010 GNDA.n1202 GNDA.n1189 1214.72
R2011 GNDA.n1194 GNDA.n1189 1214.72
R2012 GNDA.n1195 GNDA.n1194 1214.72
R2013 GNDA.n1195 GNDA.n87 1214.72
R2014 GNDA.n2301 GNDA.n87 1214.72
R2015 GNDA.n1569 GNDA.n1568 1185.07
R2016 GNDA.n1568 GNDA.n1536 1185.07
R2017 GNDA.n1926 GNDA.n1925 1182.8
R2018 GNDA.n1911 GNDA.n166 1182.8
R2019 GNDA.t528 GNDA.n1901 1016.55
R2020 GNDA.n2101 GNDA.n2100 970.366
R2021 GNDA.n2060 GNDA.t485 823.313
R2022 GNDA.n1205 GNDA.t485 823.313
R2023 GNDA.n2009 GNDA.n156 760.444
R2024 GNDA.n2001 GNDA.t540 749.742
R2025 GNDA.n2003 GNDA.t552 749.742
R2026 GNDA.n1894 GNDA.t571 749.742
R2027 GNDA.n1879 GNDA.t494 749.742
R2028 GNDA.n402 GNDA.n401 686.717
R2029 GNDA.n1566 GNDA.n1565 686.717
R2030 GNDA.n2010 GNDA.n2009 686.717
R2031 GNDA.n2010 GNDA.n155 686.717
R2032 GNDA.n1558 GNDA.n1542 686.717
R2033 GNDA.n398 GNDA.n387 686.717
R2034 GNDA.n2016 GNDA.n152 669.307
R2035 GNDA.n1966 GNDA.t567 659.367
R2036 GNDA.n1941 GNDA.t543 659.367
R2037 GNDA.n1823 GNDA.n1822 585.001
R2038 GNDA.n1742 GNDA.n1741 585.001
R2039 GNDA.n1736 GNDA.n1735 585.001
R2040 GNDA.n1633 GNDA.n1632 585.001
R2041 GNDA.n1647 GNDA.n1646 585.001
R2042 GNDA.n1636 GNDA.n157 585.001
R2043 GNDA.n1455 GNDA.n1454 585
R2044 GNDA.n1395 GNDA.n1394 585
R2045 GNDA.n1453 GNDA.n1395 585
R2046 GNDA.n1451 GNDA.n1450 585
R2047 GNDA.n1452 GNDA.n1451 585
R2048 GNDA.n1449 GNDA.n1397 585
R2049 GNDA.n1397 GNDA.n1396 585
R2050 GNDA.n1448 GNDA.n1447 585
R2051 GNDA.n1447 GNDA.n1446 585
R2052 GNDA.n1445 GNDA.n1398 585
R2053 GNDA.n1445 GNDA.n386 585
R2054 GNDA.n1444 GNDA.n1443 585
R2055 GNDA.n1444 GNDA.n385 585
R2056 GNDA.n1442 GNDA.n1399 585
R2057 GNDA.n1438 GNDA.n1399 585
R2058 GNDA.n1441 GNDA.n1440 585
R2059 GNDA.n1440 GNDA.n1439 585
R2060 GNDA.n1401 GNDA.n1400 585
R2061 GNDA.n1437 GNDA.n1401 585
R2062 GNDA.n1435 GNDA.n1434 585
R2063 GNDA.n1436 GNDA.n1435 585
R2064 GNDA.n1433 GNDA.n1403 585
R2065 GNDA.n1403 GNDA.n1402 585
R2066 GNDA.n1393 GNDA.n156 585
R2067 GNDA.n841 GNDA.n840 585
R2068 GNDA.n835 GNDA.n778 585
R2069 GNDA.n839 GNDA.n778 585
R2070 GNDA.n837 GNDA.n836 585
R2071 GNDA.n838 GNDA.n837 585
R2072 GNDA.n834 GNDA.n780 585
R2073 GNDA.n780 GNDA.n779 585
R2074 GNDA.n833 GNDA.n832 585
R2075 GNDA.n832 GNDA.n831 585
R2076 GNDA.n829 GNDA.n781 585
R2077 GNDA.n830 GNDA.n829 585
R2078 GNDA.n828 GNDA.n783 585
R2079 GNDA.n828 GNDA.n827 585
R2080 GNDA.n822 GNDA.n782 585
R2081 GNDA.n826 GNDA.n782 585
R2082 GNDA.n824 GNDA.n823 585
R2083 GNDA.n825 GNDA.n824 585
R2084 GNDA.n821 GNDA.n785 585
R2085 GNDA.n785 GNDA.n784 585
R2086 GNDA.n820 GNDA.n819 585
R2087 GNDA.n819 GNDA.n818 585
R2088 GNDA.n816 GNDA.n786 585
R2089 GNDA.n817 GNDA.n816 585
R2090 GNDA.n843 GNDA.n777 585
R2091 GNDA.n2125 GNDA.n2124 585
R2092 GNDA.n2127 GNDA.n117 585
R2093 GNDA.n2119 GNDA.n118 585
R2094 GNDA.n2123 GNDA.n118 585
R2095 GNDA.n2121 GNDA.n2120 585
R2096 GNDA.n2122 GNDA.n2121 585
R2097 GNDA.n2118 GNDA.n120 585
R2098 GNDA.n120 GNDA.n119 585
R2099 GNDA.n2117 GNDA.n2116 585
R2100 GNDA.n2116 GNDA.n2115 585
R2101 GNDA.n2113 GNDA.n121 585
R2102 GNDA.n2114 GNDA.n2113 585
R2103 GNDA.n2112 GNDA.n123 585
R2104 GNDA.n2112 GNDA.n2111 585
R2105 GNDA.n2106 GNDA.n122 585
R2106 GNDA.n2110 GNDA.n122 585
R2107 GNDA.n2108 GNDA.n2107 585
R2108 GNDA.n2109 GNDA.n2108 585
R2109 GNDA.n2105 GNDA.n125 585
R2110 GNDA.n125 GNDA.n124 585
R2111 GNDA.n2104 GNDA.n2103 585
R2112 GNDA.n2103 GNDA.n2102 585
R2113 GNDA.n127 GNDA.n126 585
R2114 GNDA.n2101 GNDA.n127 585
R2115 GNDA.n2202 GNDA.n113 585
R2116 GNDA.n2202 GNDA.n2201 585
R2117 GNDA.n2052 GNDA.n112 585
R2118 GNDA.n114 GNDA.n112 585
R2119 GNDA.n2053 GNDA.n2051 585
R2120 GNDA.n2051 GNDA.n2048 585
R2121 GNDA.n2054 GNDA.n2047 585
R2122 GNDA.n2056 GNDA.n2047 585
R2123 GNDA.n2050 GNDA.n2046 585
R2124 GNDA.n2057 GNDA.n2046 585
R2125 GNDA.n2045 GNDA.n2043 585
R2126 GNDA.n2058 GNDA.n2045 585
R2127 GNDA.n2062 GNDA.n2042 585
R2128 GNDA.n2060 GNDA.n2042 585
R2129 GNDA.n2063 GNDA.n2041 585
R2130 GNDA.n2041 GNDA.n2038 585
R2131 GNDA.n2064 GNDA.n2037 585
R2132 GNDA.n2066 GNDA.n2037 585
R2133 GNDA.n2040 GNDA.n2036 585
R2134 GNDA.n2067 GNDA.n2036 585
R2135 GNDA.n2035 GNDA.n2033 585
R2136 GNDA.n2068 GNDA.n2035 585
R2137 GNDA.n2071 GNDA.n143 585
R2138 GNDA.n143 GNDA.n140 585
R2139 GNDA.n2071 GNDA.n2070 585
R2140 GNDA.n2070 GNDA.n140 585
R2141 GNDA.n2069 GNDA.n2033 585
R2142 GNDA.n2069 GNDA.n2068 585
R2143 GNDA.n2040 GNDA.n2034 585
R2144 GNDA.n2067 GNDA.n2034 585
R2145 GNDA.n2065 GNDA.n2064 585
R2146 GNDA.n2066 GNDA.n2065 585
R2147 GNDA.n2063 GNDA.n2039 585
R2148 GNDA.n2039 GNDA.n2038 585
R2149 GNDA.n2062 GNDA.n2061 585
R2150 GNDA.n2061 GNDA.n2060 585
R2151 GNDA.n2059 GNDA.n2043 585
R2152 GNDA.n2059 GNDA.n2058 585
R2153 GNDA.n2050 GNDA.n2044 585
R2154 GNDA.n2057 GNDA.n2044 585
R2155 GNDA.n2055 GNDA.n2054 585
R2156 GNDA.n2056 GNDA.n2055 585
R2157 GNDA.n2053 GNDA.n2049 585
R2158 GNDA.n2049 GNDA.n2048 585
R2159 GNDA.n2052 GNDA.n115 585
R2160 GNDA.n115 GNDA.n114 585
R2161 GNDA.n2200 GNDA.n113 585
R2162 GNDA.n2201 GNDA.n2200 585
R2163 GNDA.n944 GNDA.n636 585
R2164 GNDA.n946 GNDA.n629 585
R2165 GNDA.n947 GNDA.n628 585
R2166 GNDA.n950 GNDA.n627 585
R2167 GNDA.n951 GNDA.n626 585
R2168 GNDA.n954 GNDA.n625 585
R2169 GNDA.n955 GNDA.n624 585
R2170 GNDA.n958 GNDA.n623 585
R2171 GNDA.n959 GNDA.n622 585
R2172 GNDA.n960 GNDA.n621 585
R2173 GNDA.n620 GNDA.n611 585
R2174 GNDA.n966 GNDA.n965 585
R2175 GNDA.n965 GNDA.n964 585
R2176 GNDA.n613 GNDA.n611 585
R2177 GNDA.n961 GNDA.n960 585
R2178 GNDA.n962 GNDA.n961 585
R2179 GNDA.n959 GNDA.n619 585
R2180 GNDA.n958 GNDA.n957 585
R2181 GNDA.n956 GNDA.n955 585
R2182 GNDA.n954 GNDA.n953 585
R2183 GNDA.n952 GNDA.n951 585
R2184 GNDA.n950 GNDA.n949 585
R2185 GNDA.n948 GNDA.n947 585
R2186 GNDA.n946 GNDA.n945 585
R2187 GNDA.n944 GNDA.n618 585
R2188 GNDA.n962 GNDA.n618 585
R2189 GNDA.n1629 GNDA.n441 585
R2190 GNDA.n1621 GNDA.n442 585
R2191 GNDA.n1625 GNDA.n1624 585
R2192 GNDA.n1620 GNDA.n1599 585
R2193 GNDA.n1617 GNDA.n1616 585
R2194 GNDA.n1615 GNDA.n1612 585
R2195 GNDA.n1611 GNDA.n1610 585
R2196 GNDA.n1609 GNDA.n1606 585
R2197 GNDA.n1605 GNDA.n1604 585
R2198 GNDA.n1603 GNDA.n1601 585
R2199 GNDA.n1600 GNDA.n377 585
R2200 GNDA.n1680 GNDA.n1679 585
R2201 GNDA.n1679 GNDA.n1678 585
R2202 GNDA.n379 GNDA.n377 585
R2203 GNDA.n1603 GNDA.n1602 585
R2204 GNDA.n1607 GNDA.n1604 585
R2205 GNDA.n1609 GNDA.n1608 585
R2206 GNDA.n1613 GNDA.n1610 585
R2207 GNDA.n1615 GNDA.n1614 585
R2208 GNDA.n1618 GNDA.n1617 585
R2209 GNDA.n1620 GNDA.n1619 585
R2210 GNDA.n1624 GNDA.n1623 585
R2211 GNDA.n1622 GNDA.n1621 585
R2212 GNDA.n441 GNDA.n440 585
R2213 GNDA.n1730 GNDA.n344 585
R2214 GNDA.n352 GNDA.n345 585
R2215 GNDA.n1726 GNDA.n1725 585
R2216 GNDA.n351 GNDA.n350 585
R2217 GNDA.n357 GNDA.n356 585
R2218 GNDA.n1718 GNDA.n1717 585
R2219 GNDA.n1716 GNDA.n1715 585
R2220 GNDA.n1714 GNDA.n361 585
R2221 GNDA.n360 GNDA.n359 585
R2222 GNDA.n1708 GNDA.n1707 585
R2223 GNDA.n1706 GNDA.n1705 585
R2224 GNDA.n1704 GNDA.n364 585
R2225 GNDA.n1704 GNDA.n1703 585
R2226 GNDA.n1705 GNDA.n362 585
R2227 GNDA.n1709 GNDA.n1708 585
R2228 GNDA.n1711 GNDA.n359 585
R2229 GNDA.n1714 GNDA.n1713 585
R2230 GNDA.n1715 GNDA.n358 585
R2231 GNDA.n1719 GNDA.n1718 585
R2232 GNDA.n1721 GNDA.n357 585
R2233 GNDA.n1722 GNDA.n351 585
R2234 GNDA.n1725 GNDA.n1724 585
R2235 GNDA.n353 GNDA.n352 585
R2236 GNDA.n344 GNDA.n340 585
R2237 GNDA.n1016 GNDA.n527 585
R2238 GNDA.n536 GNDA.n528 585
R2239 GNDA.n1012 GNDA.n1011 585
R2240 GNDA.n535 GNDA.n534 585
R2241 GNDA.n540 GNDA.n539 585
R2242 GNDA.n1004 GNDA.n1003 585
R2243 GNDA.n1002 GNDA.n1001 585
R2244 GNDA.n1000 GNDA.n544 585
R2245 GNDA.n543 GNDA.n542 585
R2246 GNDA.n994 GNDA.n993 585
R2247 GNDA.n992 GNDA.n991 585
R2248 GNDA.n990 GNDA.n547 585
R2249 GNDA.n990 GNDA.n989 585
R2250 GNDA.n991 GNDA.n545 585
R2251 GNDA.n995 GNDA.n994 585
R2252 GNDA.n997 GNDA.n542 585
R2253 GNDA.n1000 GNDA.n999 585
R2254 GNDA.n1001 GNDA.n541 585
R2255 GNDA.n1005 GNDA.n1004 585
R2256 GNDA.n1007 GNDA.n540 585
R2257 GNDA.n1008 GNDA.n535 585
R2258 GNDA.n1011 GNDA.n1010 585
R2259 GNDA.n537 GNDA.n536 585
R2260 GNDA.n713 GNDA.n527 585
R2261 GNDA.n2302 GNDA.n86 585
R2262 GNDA.n2302 GNDA.n2301 585
R2263 GNDA.n1193 GNDA.n85 585
R2264 GNDA.n87 GNDA.n85 585
R2265 GNDA.n1197 GNDA.n1192 585
R2266 GNDA.n1195 GNDA.n1192 585
R2267 GNDA.n1198 GNDA.n1191 585
R2268 GNDA.n1194 GNDA.n1191 585
R2269 GNDA.n1199 GNDA.n1187 585
R2270 GNDA.n1189 GNDA.n1187 585
R2271 GNDA.n1203 GNDA.n1188 585
R2272 GNDA.n1203 GNDA.n1202 585
R2273 GNDA.n1204 GNDA.n1185 585
R2274 GNDA.n1205 GNDA.n1204 585
R2275 GNDA.n1208 GNDA.n1184 585
R2276 GNDA.n1206 GNDA.n1184 585
R2277 GNDA.n1209 GNDA.n1183 585
R2278 GNDA.n1183 GNDA.n1181 585
R2279 GNDA.n1210 GNDA.n1180 585
R2280 GNDA.n1212 GNDA.n1180 585
R2281 GNDA.n1179 GNDA.n1166 585
R2282 GNDA.n1213 GNDA.n1179 585
R2283 GNDA.n1216 GNDA.n1164 585
R2284 GNDA.n1214 GNDA.n1164 585
R2285 GNDA.n1216 GNDA.n1215 585
R2286 GNDA.n1215 GNDA.n1214 585
R2287 GNDA.n1178 GNDA.n1166 585
R2288 GNDA.n1213 GNDA.n1178 585
R2289 GNDA.n1211 GNDA.n1210 585
R2290 GNDA.n1212 GNDA.n1211 585
R2291 GNDA.n1209 GNDA.n1182 585
R2292 GNDA.n1182 GNDA.n1181 585
R2293 GNDA.n1208 GNDA.n1207 585
R2294 GNDA.n1207 GNDA.n1206 585
R2295 GNDA.n1186 GNDA.n1185 585
R2296 GNDA.n1205 GNDA.n1186 585
R2297 GNDA.n1201 GNDA.n1188 585
R2298 GNDA.n1202 GNDA.n1201 585
R2299 GNDA.n1200 GNDA.n1199 585
R2300 GNDA.n1200 GNDA.n1189 585
R2301 GNDA.n1198 GNDA.n1190 585
R2302 GNDA.n1194 GNDA.n1190 585
R2303 GNDA.n1197 GNDA.n1196 585
R2304 GNDA.n1196 GNDA.n1195 585
R2305 GNDA.n1193 GNDA.n88 585
R2306 GNDA.n88 GNDA.n87 585
R2307 GNDA.n2300 GNDA.n86 585
R2308 GNDA.n2301 GNDA.n2300 585
R2309 GNDA.n1219 GNDA.n1218 585
R2310 GNDA.n1220 GNDA.n1219 585
R2311 GNDA.n1162 GNDA.n1161 585
R2312 GNDA.n1221 GNDA.n1162 585
R2313 GNDA.n1224 GNDA.n1223 585
R2314 GNDA.n1223 GNDA.n1222 585
R2315 GNDA.n1225 GNDA.n1160 585
R2316 GNDA.n1160 GNDA.n1159 585
R2317 GNDA.n1227 GNDA.n1226 585
R2318 GNDA.n1228 GNDA.n1227 585
R2319 GNDA.n1158 GNDA.n1157 585
R2320 GNDA.n1229 GNDA.n1158 585
R2321 GNDA.n1232 GNDA.n1231 585
R2322 GNDA.n1231 GNDA.n1230 585
R2323 GNDA.n1233 GNDA.n1156 585
R2324 GNDA.n1156 GNDA.n1155 585
R2325 GNDA.n1235 GNDA.n1234 585
R2326 GNDA.n1236 GNDA.n1235 585
R2327 GNDA.n1153 GNDA.n1152 585
R2328 GNDA.n1237 GNDA.n1153 585
R2329 GNDA.n1240 GNDA.n1239 585
R2330 GNDA.n1239 GNDA.n1238 585
R2331 GNDA.n1241 GNDA.n1151 585
R2332 GNDA.n1154 GNDA.n1151 585
R2333 GNDA.n2074 GNDA.n2073 585
R2334 GNDA.n2075 GNDA.n2074 585
R2335 GNDA.n2032 GNDA.n142 585
R2336 GNDA.n142 GNDA.n141 585
R2337 GNDA.n2031 GNDA.n2030 585
R2338 GNDA.n2030 GNDA.n2029 585
R2339 GNDA.n145 GNDA.n144 585
R2340 GNDA.n2028 GNDA.n145 585
R2341 GNDA.n2026 GNDA.n2025 585
R2342 GNDA.n2027 GNDA.n2026 585
R2343 GNDA.n2024 GNDA.n147 585
R2344 GNDA.n147 GNDA.n146 585
R2345 GNDA.n2022 GNDA.n2021 585
R2346 GNDA.n2021 GNDA.n2020 585
R2347 GNDA.n150 GNDA.n149 585
R2348 GNDA.n151 GNDA.n150 585
R2349 GNDA.n1171 GNDA.n1169 585
R2350 GNDA.n1169 GNDA.n1168 585
R2351 GNDA.n1173 GNDA.n1172 585
R2352 GNDA.n1174 GNDA.n1173 585
R2353 GNDA.n1170 GNDA.n1167 585
R2354 GNDA.n1175 GNDA.n1167 585
R2355 GNDA.n1177 GNDA.n1165 585
R2356 GNDA.n1177 GNDA.n1176 585
R2357 GNDA.n2099 GNDA.n2098 585
R2358 GNDA.n2100 GNDA.n2099 585
R2359 GNDA.n2097 GNDA.n129 585
R2360 GNDA.n129 GNDA.n128 585
R2361 GNDA.n2096 GNDA.n2095 585
R2362 GNDA.n2095 GNDA.n2094 585
R2363 GNDA.n131 GNDA.n130 585
R2364 GNDA.n2093 GNDA.n131 585
R2365 GNDA.n2091 GNDA.n2090 585
R2366 GNDA.n2092 GNDA.n2091 585
R2367 GNDA.n2089 GNDA.n133 585
R2368 GNDA.n133 GNDA.n132 585
R2369 GNDA.n2088 GNDA.n2087 585
R2370 GNDA.n2087 GNDA.n2086 585
R2371 GNDA.n135 GNDA.n134 585
R2372 GNDA.n2085 GNDA.n135 585
R2373 GNDA.n2083 GNDA.n2082 585
R2374 GNDA.n2084 GNDA.n2083 585
R2375 GNDA.n2081 GNDA.n137 585
R2376 GNDA.n137 GNDA.n136 585
R2377 GNDA.n2080 GNDA.n2079 585
R2378 GNDA.n2079 GNDA.n2078 585
R2379 GNDA.n139 GNDA.n138 585
R2380 GNDA.n2077 GNDA.n139 585
R2381 GNDA.n2018 GNDA.n2017 585
R2382 GNDA.n2019 GNDA.n148 585
R2383 GNDA.t485 GNDA.n2019 585
R2384 GNDA.n598 GNDA.n597 585
R2385 GNDA.n596 GNDA.n554 585
R2386 GNDA.n595 GNDA.n594 585
R2387 GNDA.n593 GNDA.n592 585
R2388 GNDA.n591 GNDA.n590 585
R2389 GNDA.n589 GNDA.n588 585
R2390 GNDA.n587 GNDA.n586 585
R2391 GNDA.n585 GNDA.n584 585
R2392 GNDA.n583 GNDA.n582 585
R2393 GNDA.n581 GNDA.n580 585
R2394 GNDA.n579 GNDA.n578 585
R2395 GNDA.n577 GNDA.n576 585
R2396 GNDA.n968 GNDA.n967 585
R2397 GNDA.n969 GNDA.n607 585
R2398 GNDA.n971 GNDA.n970 585
R2399 GNDA.n973 GNDA.n605 585
R2400 GNDA.n975 GNDA.n974 585
R2401 GNDA.n976 GNDA.n604 585
R2402 GNDA.n978 GNDA.n977 585
R2403 GNDA.n980 GNDA.n602 585
R2404 GNDA.n982 GNDA.n981 585
R2405 GNDA.n983 GNDA.n601 585
R2406 GNDA.n985 GNDA.n984 585
R2407 GNDA.n987 GNDA.n548 585
R2408 GNDA.n815 GNDA.n814 585
R2409 GNDA.n813 GNDA.n812 585
R2410 GNDA.n811 GNDA.n788 585
R2411 GNDA.n809 GNDA.n808 585
R2412 GNDA.n807 GNDA.n789 585
R2413 GNDA.n806 GNDA.n805 585
R2414 GNDA.n803 GNDA.n790 585
R2415 GNDA.n801 GNDA.n800 585
R2416 GNDA.n799 GNDA.n791 585
R2417 GNDA.n798 GNDA.n797 585
R2418 GNDA.n795 GNDA.n793 585
R2419 GNDA.n792 GNDA.n612 585
R2420 GNDA.n2303 GNDA.n84 585
R2421 GNDA.n2303 GNDA.n83 585
R2422 GNDA.n2393 GNDA.n2392 585
R2423 GNDA.n2390 GNDA.n54 585
R2424 GNDA.n59 GNDA.n58 585
R2425 GNDA.n2385 GNDA.n2384 585
R2426 GNDA.n2383 GNDA.n2382 585
R2427 GNDA.n2309 GNDA.n63 585
R2428 GNDA.n2311 GNDA.n2310 585
R2429 GNDA.n2316 GNDA.n2315 585
R2430 GNDA.n2314 GNDA.n2307 585
R2431 GNDA.n2322 GNDA.n2321 585
R2432 GNDA.n2324 GNDA.n2323 585
R2433 GNDA.n2305 GNDA.n2304 585
R2434 GNDA.n2203 GNDA.n111 585
R2435 GNDA.n2203 GNDA.n83 585
R2436 GNDA.n2299 GNDA.n84 585
R2437 GNDA.n2299 GNDA.n83 585
R2438 GNDA.n2298 GNDA.n2297 585
R2439 GNDA.n2295 GNDA.n2294 585
R2440 GNDA.n2293 GNDA.n2292 585
R2441 GNDA.n2209 GNDA.n91 585
R2442 GNDA.n2211 GNDA.n2210 585
R2443 GNDA.n2215 GNDA.n2214 585
R2444 GNDA.n2217 GNDA.n2216 585
R2445 GNDA.n2224 GNDA.n2223 585
R2446 GNDA.n2222 GNDA.n2207 585
R2447 GNDA.n2230 GNDA.n2229 585
R2448 GNDA.n2232 GNDA.n2231 585
R2449 GNDA.n2205 GNDA.n2204 585
R2450 GNDA.n2199 GNDA.n111 585
R2451 GNDA.n2199 GNDA.n83 585
R2452 GNDA.n2198 GNDA.n2197 585
R2453 GNDA.n24 GNDA.n22 585
R2454 GNDA.n2398 GNDA.n2397 585
R2455 GNDA.n32 GNDA.n25 585
R2456 GNDA.n40 GNDA.n39 585
R2457 GNDA.n35 GNDA.n31 585
R2458 GNDA.n30 GNDA.n0 585
R2459 GNDA.n2132 GNDA.n1 585
R2460 GNDA.n2134 GNDA.n2133 585
R2461 GNDA.n2138 GNDA.n2137 585
R2462 GNDA.n2140 GNDA.n2139 585
R2463 GNDA.n2129 GNDA.n2128 585
R2464 GNDA.n1107 GNDA.n1106 585
R2465 GNDA.n1109 GNDA.n1104 585
R2466 GNDA.n1111 GNDA.n1110 585
R2467 GNDA.n1112 GNDA.n1103 585
R2468 GNDA.n1114 GNDA.n1113 585
R2469 GNDA.n1116 GNDA.n1101 585
R2470 GNDA.n1118 GNDA.n1117 585
R2471 GNDA.n1119 GNDA.n1100 585
R2472 GNDA.n1121 GNDA.n1120 585
R2473 GNDA.n1123 GNDA.n1098 585
R2474 GNDA.n1125 GNDA.n1124 585
R2475 GNDA.n1126 GNDA.n1097 585
R2476 GNDA.n1682 GNDA.n1681 585
R2477 GNDA.n1683 GNDA.n373 585
R2478 GNDA.n1685 GNDA.n1684 585
R2479 GNDA.n1687 GNDA.n371 585
R2480 GNDA.n1689 GNDA.n1688 585
R2481 GNDA.n1690 GNDA.n370 585
R2482 GNDA.n1692 GNDA.n1691 585
R2483 GNDA.n1694 GNDA.n368 585
R2484 GNDA.n1696 GNDA.n1695 585
R2485 GNDA.n1697 GNDA.n367 585
R2486 GNDA.n1699 GNDA.n1698 585
R2487 GNDA.n1701 GNDA.n365 585
R2488 GNDA.n1432 GNDA.n1431 585
R2489 GNDA.n1429 GNDA.n1404 585
R2490 GNDA.n1428 GNDA.n1427 585
R2491 GNDA.n1426 GNDA.n1425 585
R2492 GNDA.n1424 GNDA.n1406 585
R2493 GNDA.n1422 GNDA.n1421 585
R2494 GNDA.n1420 GNDA.n1407 585
R2495 GNDA.n1419 GNDA.n1418 585
R2496 GNDA.n1416 GNDA.n1408 585
R2497 GNDA.n1414 GNDA.n1413 585
R2498 GNDA.n1412 GNDA.n1410 585
R2499 GNDA.n1411 GNDA.n378 585
R2500 GNDA.n1017 GNDA.n526 585
R2501 GNDA.n1017 GNDA.n525 585
R2502 GNDA.n1086 GNDA.n456 585
R2503 GNDA.n1084 GNDA.n1083 585
R2504 GNDA.n479 GNDA.n460 585
R2505 GNDA.n1079 GNDA.n1078 585
R2506 GNDA.n481 GNDA.n478 585
R2507 GNDA.n507 GNDA.n506 585
R2508 GNDA.n509 GNDA.n508 585
R2509 GNDA.n512 GNDA.n511 585
R2510 GNDA.n510 GNDA.n500 585
R2511 GNDA.n521 GNDA.n520 585
R2512 GNDA.n523 GNDA.n522 585
R2513 GNDA.n1019 GNDA.n1018 585
R2514 GNDA.n942 GNDA.n939 585
R2515 GNDA.n939 GNDA.n525 585
R2516 GNDA.n714 GNDA.n526 585
R2517 GNDA.n714 GNDA.n525 585
R2518 GNDA.n716 GNDA.n715 585
R2519 GNDA.n740 GNDA.n718 585
R2520 GNDA.n742 GNDA.n741 585
R2521 GNDA.n738 GNDA.n737 585
R2522 GNDA.n736 GNDA.n735 585
R2523 GNDA.n731 GNDA.n730 585
R2524 GNDA.n729 GNDA.n728 585
R2525 GNDA.n724 GNDA.n723 585
R2526 GNDA.n722 GNDA.n639 585
R2527 GNDA.n750 GNDA.n749 585
R2528 GNDA.n752 GNDA.n751 585
R2529 GNDA.n938 GNDA.n754 585
R2530 GNDA.n942 GNDA.n941 585
R2531 GNDA.n941 GNDA.n525 585
R2532 GNDA.n940 GNDA.n937 585
R2533 GNDA.n935 GNDA.n934 585
R2534 GNDA.n933 GNDA.n932 585
R2535 GNDA.n849 GNDA.n757 585
R2536 GNDA.n851 GNDA.n850 585
R2537 GNDA.n855 GNDA.n854 585
R2538 GNDA.n857 GNDA.n856 585
R2539 GNDA.n864 GNDA.n863 585
R2540 GNDA.n862 GNDA.n847 585
R2541 GNDA.n870 GNDA.n869 585
R2542 GNDA.n872 GNDA.n871 585
R2543 GNDA.n845 GNDA.n844 585
R2544 GNDA.n1147 GNDA.n1146 585
R2545 GNDA.n1145 GNDA.n1096 585
R2546 GNDA.n1144 GNDA.n1143 585
R2547 GNDA.n1142 GNDA.n1141 585
R2548 GNDA.n1140 GNDA.n1139 585
R2549 GNDA.n1138 GNDA.n1137 585
R2550 GNDA.n1136 GNDA.n1135 585
R2551 GNDA.n1134 GNDA.n1133 585
R2552 GNDA.n1132 GNDA.n1131 585
R2553 GNDA.n1130 GNDA.n1129 585
R2554 GNDA.n1128 GNDA.n1127 585
R2555 GNDA.n1264 GNDA.n296 585
R2556 GNDA.n575 GNDA.n574 585
R2557 GNDA.n573 GNDA.n572 585
R2558 GNDA.n571 GNDA.n570 585
R2559 GNDA.n569 GNDA.n568 585
R2560 GNDA.n567 GNDA.n566 585
R2561 GNDA.n565 GNDA.n564 585
R2562 GNDA.n563 GNDA.n562 585
R2563 GNDA.n561 GNDA.n560 585
R2564 GNDA.n559 GNDA.n558 585
R2565 GNDA.n557 GNDA.n556 585
R2566 GNDA.n555 GNDA.n457 585
R2567 GNDA.n1264 GNDA.n1089 585
R2568 GNDA.n1262 GNDA.n1261 585
R2569 GNDA.n1260 GNDA.n1150 585
R2570 GNDA.n1259 GNDA.n1149 585
R2571 GNDA.n1264 GNDA.n1149 585
R2572 GNDA.n1258 GNDA.n1257 585
R2573 GNDA.n1256 GNDA.n1255 585
R2574 GNDA.n1254 GNDA.n1253 585
R2575 GNDA.n1252 GNDA.n1251 585
R2576 GNDA.n1250 GNDA.n1249 585
R2577 GNDA.n1248 GNDA.n1247 585
R2578 GNDA.n1246 GNDA.n1245 585
R2579 GNDA.n1244 GNDA.n1243 585
R2580 GNDA.n1242 GNDA.n56 585
R2581 GNDA.n56 GNDA.n55 585
R2582 GNDA.n1541 GNDA.n1538 585
R2583 GNDA.n1563 GNDA.n1562 585
R2584 GNDA.n1564 GNDA.n1563 585
R2585 GNDA.n1560 GNDA.n1557 585
R2586 GNDA.n391 GNDA.n389 585
R2587 GNDA.n395 GNDA.n388 585
R2588 GNDA.n403 GNDA.n388 585
R2589 GNDA.n394 GNDA.n393 585
R2590 GNDA.n1732 GNDA.n1731 585
R2591 GNDA.n1731 GNDA.n332 585
R2592 GNDA.n1820 GNDA.n1819 585
R2593 GNDA.n1821 GNDA.n1820 585
R2594 GNDA.n1817 GNDA.n297 585
R2595 GNDA.n306 GNDA.n297 585
R2596 GNDA.n304 GNDA.n300 585
R2597 GNDA.n307 GNDA.n304 585
R2598 GNDA.n1812 GNDA.n1811 585
R2599 GNDA.n1811 GNDA.n1810 585
R2600 GNDA.n309 GNDA.n305 585
R2601 GNDA.n1809 GNDA.n305 585
R2602 GNDA.n1807 GNDA.n1806 585
R2603 GNDA.n1808 GNDA.n1807 585
R2604 GNDA.n1546 GNDA.n308 585
R2605 GNDA.n1556 GNDA.n308 585
R2606 GNDA.n1554 GNDA.n1553 585
R2607 GNDA.n1555 GNDA.n1554 585
R2608 GNDA.n1548 GNDA.n1545 585
R2609 GNDA.n1545 GNDA.n1544 585
R2610 GNDA.n330 GNDA.n329 585
R2611 GNDA.n1543 GNDA.n330 585
R2612 GNDA.n1746 GNDA.n1745 585
R2613 GNDA.n1745 GNDA.n1744 585
R2614 GNDA.n342 GNDA.n331 585
R2615 GNDA.n1743 GNDA.n331 585
R2616 GNDA.n1630 GNDA.n438 585
R2617 GNDA.n1631 GNDA.n1630 585
R2618 GNDA.n1733 GNDA.n1732 585
R2619 GNDA.n1734 GNDA.n1733 585
R2620 GNDA.n1334 GNDA.n341 585
R2621 GNDA.n341 GNDA.n339 585
R2622 GNDA.n1321 GNDA.n1319 585
R2623 GNDA.n1570 GNDA.n1321 585
R2624 GNDA.n1585 GNDA.n1584 585
R2625 GNDA.n1584 GNDA.n1583 585
R2626 GNDA.n1572 GNDA.n1322 585
R2627 GNDA.n1582 GNDA.n1322 585
R2628 GNDA.n1580 GNDA.n1579 585
R2629 GNDA.n1581 GNDA.n1580 585
R2630 GNDA.n1575 GNDA.n1296 585
R2631 GNDA.n1571 GNDA.n1296 585
R2632 GNDA.n1593 GNDA.n1592 585
R2633 GNDA.n1594 GNDA.n1593 585
R2634 GNDA.n1298 GNDA.n1297 585
R2635 GNDA.n1325 GNDA.n1297 585
R2636 GNDA.n1329 GNDA.n1328 585
R2637 GNDA.n1328 GNDA.n1327 585
R2638 GNDA.n1332 GNDA.n1323 585
R2639 GNDA.n1326 GNDA.n1323 585
R2640 GNDA.n1533 GNDA.n1532 585
R2641 GNDA.n1534 GNDA.n1533 585
R2642 GNDA.n1530 GNDA.n437 585
R2643 GNDA.n1535 GNDA.n437 585
R2644 GNDA.n439 GNDA.n438 585
R2645 GNDA.n439 GNDA.n430 585
R2646 GNDA.n1528 GNDA.n429 585
R2647 GNDA.n1648 GNDA.n429 585
R2648 GNDA.n1650 GNDA.n427 585
R2649 GNDA.n1650 GNDA.n1649 585
R2650 GNDA.n1666 GNDA.n1665 585
R2651 GNDA.n1665 GNDA.n1664 585
R2652 GNDA.n1653 GNDA.n1651 585
R2653 GNDA.n1663 GNDA.n1651 585
R2654 GNDA.n1661 GNDA.n1660 585
R2655 GNDA.n1662 GNDA.n1661 585
R2656 GNDA.n1656 GNDA.n404 585
R2657 GNDA.n1652 GNDA.n404 585
R2658 GNDA.n1674 GNDA.n1673 585
R2659 GNDA.n1675 GNDA.n1674 585
R2660 GNDA.n406 GNDA.n405 585
R2661 GNDA.n1460 GNDA.n405 585
R2662 GNDA.n1465 GNDA.n1464 585
R2663 GNDA.n1466 GNDA.n1465 585
R2664 GNDA.n1392 GNDA.n1391 585
R2665 GNDA.n1467 GNDA.n1392 585
R2666 GNDA.n1471 GNDA.n1470 585
R2667 GNDA.n1470 GNDA.n1469 585
R2668 GNDA.n1459 GNDA.n1458 585
R2669 GNDA.n1468 GNDA.n1459 585
R2670 GNDA.n1996 GNDA.t555 524.808
R2671 GNDA.n1989 GNDA.t549 524.808
R2672 GNDA.n1891 GNDA.t505 524.808
R2673 GNDA.n1884 GNDA.t490 524.808
R2674 GNDA.n2201 GNDA.t485 512.884
R2675 GNDA.n2301 GNDA.t485 512.884
R2676 GNDA.n1932 GNDA.t514 508.743
R2677 GNDA.n1929 GNDA.t524 508.743
R2678 GNDA.n1273 GNDA.t561 508.743
R2679 GNDA.n1974 GNDA.t508 508.743
R2680 GNDA.n1902 GNDA.t527 499.442
R2681 GNDA.n170 GNDA.t534 499.442
R2682 GNDA.n1906 GNDA.t532 499.442
R2683 GNDA.n174 GNDA.t537 499.442
R2684 GNDA.n1999 GNDA.n163 490.517
R2685 GNDA.n184 GNDA.t481 475.976
R2686 GNDA.n184 GNDA.t519 475.976
R2687 GNDA.n178 GNDA.t530 475.976
R2688 GNDA.n178 GNDA.t511 475.976
R2689 GNDA.n1637 GNDA.t564 409.067
R2690 GNDA.n1645 GNDA.t487 409.067
R2691 GNDA.n1634 GNDA.t558 409.067
R2692 GNDA.n1737 GNDA.t546 409.067
R2693 GNDA.n1740 GNDA.t498 409.067
R2694 GNDA.n1824 GNDA.t521 409.067
R2695 GNDA.n2058 GNDA.t485 391.411
R2696 GNDA.n1202 GNDA.t485 391.411
R2697 GNDA.n1901 GNDA.n1900 364.139
R2698 GNDA.n1912 GNDA.t478 338.034
R2699 GNDA.n1924 GNDA.t502 338.034
R2700 GNDA.t158 GNDA.t111 333.793
R2701 GNDA.t38 GNDA.t158 333.793
R2702 GNDA.t173 GNDA.t38 333.793
R2703 GNDA.t576 GNDA.t42 333.793
R2704 GNDA.t42 GNDA.t115 333.793
R2705 GNDA.t26 GNDA.t15 333.793
R2706 GNDA.t25 GNDA.t15 333.793
R2707 GNDA.n1728 GNDA.t485 172.876
R2708 GNDA.n1627 GNDA.t485 172.876
R2709 GNDA.t485 GNDA.n355 172.615
R2710 GNDA.n1676 GNDA.t485 172.615
R2711 GNDA.n1934 GNDA.n1933 296.158
R2712 GNDA.n1928 GNDA.n1927 296.158
R2713 GNDA.n1275 GNDA.n1274 296.158
R2714 GNDA.n1973 GNDA.n1972 296.158
R2715 GNDA.n1905 GNDA.n1904 292.5
R2716 GNDA.n1934 GNDA.n167 292.5
R2717 GNDA.n1927 GNDA.n171 292.5
R2718 GNDA.n173 GNDA.n163 292.5
R2719 GNDA.n1904 GNDA.n1903 292.5
R2720 GNDA.n169 GNDA.n163 292.5
R2721 GNDA.t591 GNDA.t485 279.212
R2722 GNDA.t206 GNDA.n155 271.719
R2723 GNDA.n1264 GNDA.n449 264.301
R2724 GNDA.n1457 GNDA.n1456 264.301
R2725 GNDA.n842 GNDA.n776 264.301
R2726 GNDA.n2126 GNDA.n116 264.301
R2727 GNDA.n1090 GNDA.n298 264.301
R2728 GNDA.n1088 GNDA.n1087 264.301
R2729 GNDA.n1219 GNDA.n1164 259.416
R2730 GNDA.n598 GNDA.n547 259.416
R2731 GNDA.n1107 GNDA.n364 259.416
R2732 GNDA.n1681 GNDA.n1680 259.416
R2733 GNDA.n967 GNDA.n966 259.416
R2734 GNDA.n2074 GNDA.n143 259.416
R2735 GNDA.n816 GNDA.n815 259.416
R2736 GNDA.n1431 GNDA.n1403 259.416
R2737 GNDA.n2099 GNDA.n127 259.416
R2738 GNDA.n2361 GNDA.n80 258.334
R2739 GNDA.n1056 GNDA.n1054 258.334
R2740 GNDA.n1783 GNDA.n326 258.334
R2741 GNDA.n1353 GNDA.n1352 258.334
R2742 GNDA.n695 GNDA.n694 258.334
R2743 GNDA.n2271 GNDA.n2270 258.334
R2744 GNDA.n911 GNDA.n910 258.334
R2745 GNDA.n1510 GNDA.n1509 258.334
R2746 GNDA.n2179 GNDA.n2178 258.334
R2747 GNDA.t82 GNDA.n166 257.932
R2748 GNDA.t50 GNDA.n1926 257.932
R2749 GNDA.n635 GNDA.n634 254.34
R2750 GNDA.n634 GNDA.n633 254.34
R2751 GNDA.n634 GNDA.n632 254.34
R2752 GNDA.n634 GNDA.n631 254.34
R2753 GNDA.n634 GNDA.n630 254.34
R2754 GNDA.n634 GNDA.n610 254.34
R2755 GNDA.n963 GNDA.n962 254.34
R2756 GNDA.n962 GNDA.n614 254.34
R2757 GNDA.n962 GNDA.n615 254.34
R2758 GNDA.n962 GNDA.n616 254.34
R2759 GNDA.n962 GNDA.n617 254.34
R2760 GNDA.n1628 GNDA.n1627 254.34
R2761 GNDA.n1627 GNDA.n1626 254.34
R2762 GNDA.n1627 GNDA.n1598 254.34
R2763 GNDA.n1627 GNDA.n1597 254.34
R2764 GNDA.n1627 GNDA.n1596 254.34
R2765 GNDA.n1627 GNDA.n376 254.34
R2766 GNDA.n1677 GNDA.n1676 254.34
R2767 GNDA.n1676 GNDA.n384 254.34
R2768 GNDA.n1676 GNDA.n383 254.34
R2769 GNDA.n1676 GNDA.n382 254.34
R2770 GNDA.n1676 GNDA.n381 254.34
R2771 GNDA.n1676 GNDA.n380 254.34
R2772 GNDA.n1729 GNDA.n1728 254.34
R2773 GNDA.n1728 GNDA.n1727 254.34
R2774 GNDA.n1728 GNDA.n349 254.34
R2775 GNDA.n1728 GNDA.n348 254.34
R2776 GNDA.n1728 GNDA.n347 254.34
R2777 GNDA.n1728 GNDA.n346 254.34
R2778 GNDA.n1702 GNDA.n355 254.34
R2779 GNDA.n1710 GNDA.n355 254.34
R2780 GNDA.n1712 GNDA.n355 254.34
R2781 GNDA.n1720 GNDA.n355 254.34
R2782 GNDA.n1723 GNDA.n355 254.34
R2783 GNDA.n355 GNDA.n354 254.34
R2784 GNDA.n1015 GNDA.n1014 254.34
R2785 GNDA.n1014 GNDA.n1013 254.34
R2786 GNDA.n1014 GNDA.n533 254.34
R2787 GNDA.n1014 GNDA.n532 254.34
R2788 GNDA.n1014 GNDA.n531 254.34
R2789 GNDA.n1014 GNDA.n530 254.34
R2790 GNDA.n988 GNDA.n538 254.34
R2791 GNDA.n996 GNDA.n538 254.34
R2792 GNDA.n998 GNDA.n538 254.34
R2793 GNDA.n1006 GNDA.n538 254.34
R2794 GNDA.n1009 GNDA.n538 254.34
R2795 GNDA.n712 GNDA.n538 254.34
R2796 GNDA.n600 GNDA.n599 254.34
R2797 GNDA.n600 GNDA.n553 254.34
R2798 GNDA.n600 GNDA.n552 254.34
R2799 GNDA.n600 GNDA.n551 254.34
R2800 GNDA.n600 GNDA.n550 254.34
R2801 GNDA.n600 GNDA.n549 254.34
R2802 GNDA.n609 GNDA.n600 254.34
R2803 GNDA.n972 GNDA.n600 254.34
R2804 GNDA.n606 GNDA.n600 254.34
R2805 GNDA.n979 GNDA.n600 254.34
R2806 GNDA.n603 GNDA.n600 254.34
R2807 GNDA.n986 GNDA.n600 254.34
R2808 GNDA.n787 GNDA.n600 254.34
R2809 GNDA.n810 GNDA.n600 254.34
R2810 GNDA.n804 GNDA.n600 254.34
R2811 GNDA.n802 GNDA.n600 254.34
R2812 GNDA.n796 GNDA.n600 254.34
R2813 GNDA.n794 GNDA.n600 254.34
R2814 GNDA.n2395 GNDA.n2394 254.34
R2815 GNDA.n2395 GNDA.n53 254.34
R2816 GNDA.n2395 GNDA.n52 254.34
R2817 GNDA.n2395 GNDA.n51 254.34
R2818 GNDA.n2395 GNDA.n50 254.34
R2819 GNDA.n2395 GNDA.n49 254.34
R2820 GNDA.n2395 GNDA.n48 254.34
R2821 GNDA.n2395 GNDA.n47 254.34
R2822 GNDA.n2395 GNDA.n46 254.34
R2823 GNDA.n2395 GNDA.n45 254.34
R2824 GNDA.n2395 GNDA.n44 254.34
R2825 GNDA.n2395 GNDA.n43 254.34
R2826 GNDA.n2395 GNDA.n42 254.34
R2827 GNDA.n2396 GNDA.n2395 254.34
R2828 GNDA.n2395 GNDA.n41 254.34
R2829 GNDA.n2395 GNDA.n29 254.34
R2830 GNDA.n2395 GNDA.n28 254.34
R2831 GNDA.n2395 GNDA.n27 254.34
R2832 GNDA.n1108 GNDA.n366 254.34
R2833 GNDA.n1105 GNDA.n366 254.34
R2834 GNDA.n1115 GNDA.n366 254.34
R2835 GNDA.n1102 GNDA.n366 254.34
R2836 GNDA.n1122 GNDA.n366 254.34
R2837 GNDA.n1099 GNDA.n366 254.34
R2838 GNDA.n375 GNDA.n366 254.34
R2839 GNDA.n1686 GNDA.n366 254.34
R2840 GNDA.n372 GNDA.n366 254.34
R2841 GNDA.n1693 GNDA.n366 254.34
R2842 GNDA.n369 GNDA.n366 254.34
R2843 GNDA.n1700 GNDA.n366 254.34
R2844 GNDA.n1430 GNDA.n366 254.34
R2845 GNDA.n1405 GNDA.n366 254.34
R2846 GNDA.n1423 GNDA.n366 254.34
R2847 GNDA.n1417 GNDA.n366 254.34
R2848 GNDA.n1415 GNDA.n366 254.34
R2849 GNDA.n1409 GNDA.n366 254.34
R2850 GNDA.n1082 GNDA.n1081 254.34
R2851 GNDA.n1081 GNDA.n1080 254.34
R2852 GNDA.n1081 GNDA.n477 254.34
R2853 GNDA.n1081 GNDA.n476 254.34
R2854 GNDA.n1081 GNDA.n475 254.34
R2855 GNDA.n1081 GNDA.n474 254.34
R2856 GNDA.n1081 GNDA.n473 254.34
R2857 GNDA.n1081 GNDA.n472 254.34
R2858 GNDA.n1081 GNDA.n471 254.34
R2859 GNDA.n1081 GNDA.n470 254.34
R2860 GNDA.n1081 GNDA.n469 254.34
R2861 GNDA.n1081 GNDA.n468 254.34
R2862 GNDA.n1081 GNDA.n467 254.34
R2863 GNDA.n1081 GNDA.n466 254.34
R2864 GNDA.n1081 GNDA.n465 254.34
R2865 GNDA.n1081 GNDA.n464 254.34
R2866 GNDA.n1081 GNDA.n463 254.34
R2867 GNDA.n1081 GNDA.n462 254.34
R2868 GNDA.n1264 GNDA.n1148 254.34
R2869 GNDA.n1264 GNDA.n1095 254.34
R2870 GNDA.n1264 GNDA.n1094 254.34
R2871 GNDA.n1264 GNDA.n1093 254.34
R2872 GNDA.n1264 GNDA.n1092 254.34
R2873 GNDA.n1264 GNDA.n1091 254.34
R2874 GNDA.n1264 GNDA.n450 254.34
R2875 GNDA.n1264 GNDA.n451 254.34
R2876 GNDA.n1264 GNDA.n452 254.34
R2877 GNDA.n1264 GNDA.n453 254.34
R2878 GNDA.n1264 GNDA.n454 254.34
R2879 GNDA.n1264 GNDA.n455 254.34
R2880 GNDA.n1264 GNDA.n1263 254.34
R2881 GNDA.n1264 GNDA.n445 254.34
R2882 GNDA.n1264 GNDA.n446 254.34
R2883 GNDA.n1264 GNDA.n447 254.34
R2884 GNDA.n1264 GNDA.n448 254.34
R2885 GNDA.t485 GNDA.n152 250.349
R2886 GNDA.n1262 GNDA.n1151 249.663
R2887 GNDA.n576 GNDA.n575 249.663
R2888 GNDA.n1147 GNDA.n1097 249.663
R2889 GNDA.n1703 GNDA.n1701 249.663
R2890 GNDA.n989 GNDA.n987 249.663
R2891 GNDA.n1215 GNDA.n1177 249.663
R2892 GNDA.n964 GNDA.n612 249.663
R2893 GNDA.n1678 GNDA.n378 249.663
R2894 GNDA.n2070 GNDA.n139 249.663
R2895 GNDA.n389 GNDA.n388 246.25
R2896 GNDA.n393 GNDA.n388 246.25
R2897 GNDA.n1563 GNDA.n1541 246.25
R2898 GNDA.n1563 GNDA.n1557 246.25
R2899 GNDA.t175 GNDA.n1276 242.76
R2900 GNDA.n2011 GNDA.n2010 241.643
R2901 GNDA.n1565 GNDA.n1564 241.643
R2902 GNDA.n1564 GNDA.n1542 241.643
R2903 GNDA.n403 GNDA.n402 241.643
R2904 GNDA.n403 GNDA.n387 241.643
R2905 GNDA.n1904 GNDA.n187 234.276
R2906 GNDA.n1911 GNDA.t480 233
R2907 GNDA.n1925 GNDA.t504 233
R2908 GNDA.n1940 GNDA.n1939 199.883
R2909 GNDA.n1968 GNDA.n1967 199.883
R2910 GNDA.n1915 GNDA.n1914 199.03
R2911 GNDA.n1917 GNDA.n1916 199.03
R2912 GNDA.n1919 GNDA.n1918 199.03
R2913 GNDA.n1921 GNDA.n1920 199.03
R2914 GNDA.n1923 GNDA.n1922 199.03
R2915 GNDA.n2019 GNDA.n2018 197
R2916 GNDA.n2304 GNDA.n2303 197
R2917 GNDA.n1018 GNDA.n1017 197
R2918 GNDA.n1731 GNDA.n331 197
R2919 GNDA.n1630 GNDA.n437 197
R2920 GNDA.n939 GNDA.n938 197
R2921 GNDA.n2204 GNDA.n2203 197
R2922 GNDA.n844 GNDA.n843 197
R2923 GNDA.n1459 GNDA.n1393 197
R2924 GNDA.n2128 GNDA.n2127 197
R2925 GNDA.n2393 GNDA.n55 187.249
R2926 GNDA.n1089 GNDA.n456 187.249
R2927 GNDA.n1820 GNDA.n296 187.249
R2928 GNDA.n1733 GNDA.n341 187.249
R2929 GNDA.n715 GNDA.n714 187.249
R2930 GNDA.n2299 GNDA.n2298 187.249
R2931 GNDA.n941 GNDA.n940 187.249
R2932 GNDA.n439 GNDA.n429 187.249
R2933 GNDA.n2199 GNDA.n2198 187.249
R2934 GNDA.n2363 GNDA.n80 185
R2935 GNDA.n2377 GNDA.n2376 185
R2936 GNDA.n2375 GNDA.n81 185
R2937 GNDA.n2374 GNDA.n2373 185
R2938 GNDA.n2372 GNDA.n2371 185
R2939 GNDA.n2370 GNDA.n2369 185
R2940 GNDA.n2368 GNDA.n2367 185
R2941 GNDA.n2366 GNDA.n2365 185
R2942 GNDA.n2364 GNDA.n57 185
R2943 GNDA.n2346 GNDA.n2345 185
R2944 GNDA.n2348 GNDA.n2347 185
R2945 GNDA.n2350 GNDA.n2349 185
R2946 GNDA.n2352 GNDA.n2351 185
R2947 GNDA.n2354 GNDA.n2353 185
R2948 GNDA.n2356 GNDA.n2355 185
R2949 GNDA.n2358 GNDA.n2357 185
R2950 GNDA.n2360 GNDA.n2359 185
R2951 GNDA.n2362 GNDA.n2361 185
R2952 GNDA.n2328 GNDA.n2327 185
R2953 GNDA.n2330 GNDA.n2329 185
R2954 GNDA.n2332 GNDA.n2331 185
R2955 GNDA.n2334 GNDA.n2333 185
R2956 GNDA.n2336 GNDA.n2335 185
R2957 GNDA.n2338 GNDA.n2337 185
R2958 GNDA.n2340 GNDA.n2339 185
R2959 GNDA.n2342 GNDA.n2341 185
R2960 GNDA.n2344 GNDA.n2343 185
R2961 GNDA.n2326 GNDA.n2325 185
R2962 GNDA.n2320 GNDA.n2319 185
R2963 GNDA.n2318 GNDA.n2317 185
R2964 GNDA.n2313 GNDA.n2312 185
R2965 GNDA.n2308 GNDA.n65 185
R2966 GNDA.n2381 GNDA.n2380 185
R2967 GNDA.n64 GNDA.n62 185
R2968 GNDA.n2387 GNDA.n2386 185
R2969 GNDA.n2389 GNDA.n2388 185
R2970 GNDA.n1057 GNDA.n1056 185
R2971 GNDA.n1058 GNDA.n486 185
R2972 GNDA.n1060 GNDA.n1059 185
R2973 GNDA.n1062 GNDA.n485 185
R2974 GNDA.n1065 GNDA.n1064 185
R2975 GNDA.n1066 GNDA.n484 185
R2976 GNDA.n1068 GNDA.n1067 185
R2977 GNDA.n1070 GNDA.n483 185
R2978 GNDA.n1071 GNDA.n458 185
R2979 GNDA.n1038 GNDA.n491 185
R2980 GNDA.n1041 GNDA.n1040 185
R2981 GNDA.n1042 GNDA.n490 185
R2982 GNDA.n1044 GNDA.n1043 185
R2983 GNDA.n1046 GNDA.n489 185
R2984 GNDA.n1049 GNDA.n1048 185
R2985 GNDA.n1050 GNDA.n488 185
R2986 GNDA.n1052 GNDA.n1051 185
R2987 GNDA.n1054 GNDA.n487 185
R2988 GNDA.n1022 GNDA.n1021 185
R2989 GNDA.n1024 GNDA.n496 185
R2990 GNDA.n1026 GNDA.n1025 185
R2991 GNDA.n1027 GNDA.n495 185
R2992 GNDA.n1029 GNDA.n1028 185
R2993 GNDA.n1031 GNDA.n493 185
R2994 GNDA.n1033 GNDA.n1032 185
R2995 GNDA.n1034 GNDA.n492 185
R2996 GNDA.n1036 GNDA.n1035 185
R2997 GNDA.n499 GNDA.n498 185
R2998 GNDA.n519 GNDA.n518 185
R2999 GNDA.n516 GNDA.n501 185
R3000 GNDA.n514 GNDA.n513 185
R3001 GNDA.n505 GNDA.n503 185
R3002 GNDA.n504 GNDA.n482 185
R3003 GNDA.n1077 GNDA.n1076 185
R3004 GNDA.n1074 GNDA.n480 185
R3005 GNDA.n1073 GNDA.n459 185
R3006 GNDA.n1785 GNDA.n326 185
R3007 GNDA.n1799 GNDA.n1798 185
R3008 GNDA.n1797 GNDA.n327 185
R3009 GNDA.n1796 GNDA.n1795 185
R3010 GNDA.n1794 GNDA.n1793 185
R3011 GNDA.n1792 GNDA.n1791 185
R3012 GNDA.n1790 GNDA.n1789 185
R3013 GNDA.n1788 GNDA.n1787 185
R3014 GNDA.n1786 GNDA.n299 185
R3015 GNDA.n1768 GNDA.n1767 185
R3016 GNDA.n1770 GNDA.n1769 185
R3017 GNDA.n1772 GNDA.n1771 185
R3018 GNDA.n1774 GNDA.n1773 185
R3019 GNDA.n1776 GNDA.n1775 185
R3020 GNDA.n1778 GNDA.n1777 185
R3021 GNDA.n1780 GNDA.n1779 185
R3022 GNDA.n1782 GNDA.n1781 185
R3023 GNDA.n1784 GNDA.n1783 185
R3024 GNDA.n1750 GNDA.n1749 185
R3025 GNDA.n1752 GNDA.n1751 185
R3026 GNDA.n1754 GNDA.n1753 185
R3027 GNDA.n1756 GNDA.n1755 185
R3028 GNDA.n1758 GNDA.n1757 185
R3029 GNDA.n1760 GNDA.n1759 185
R3030 GNDA.n1762 GNDA.n1761 185
R3031 GNDA.n1764 GNDA.n1763 185
R3032 GNDA.n1766 GNDA.n1765 185
R3033 GNDA.n1748 GNDA.n1747 185
R3034 GNDA.n1550 GNDA.n1549 185
R3035 GNDA.n1552 GNDA.n1551 185
R3036 GNDA.n1547 GNDA.n311 185
R3037 GNDA.n1805 GNDA.n1804 185
R3038 GNDA.n1802 GNDA.n310 185
R3039 GNDA.n1801 GNDA.n303 185
R3040 GNDA.n1814 GNDA.n1813 185
R3041 GNDA.n1816 GNDA.n1815 185
R3042 GNDA.n1352 GNDA.n1351 185
R3043 GNDA.n1350 GNDA.n1349 185
R3044 GNDA.n1348 GNDA.n1347 185
R3045 GNDA.n1346 GNDA.n1345 185
R3046 GNDA.n1344 GNDA.n1343 185
R3047 GNDA.n1342 GNDA.n1341 185
R3048 GNDA.n1340 GNDA.n1339 185
R3049 GNDA.n1338 GNDA.n1337 185
R3050 GNDA.n1336 GNDA.n1317 185
R3051 GNDA.n1370 GNDA.n1369 185
R3052 GNDA.n1368 GNDA.n1367 185
R3053 GNDA.n1366 GNDA.n1365 185
R3054 GNDA.n1364 GNDA.n1363 185
R3055 GNDA.n1362 GNDA.n1361 185
R3056 GNDA.n1360 GNDA.n1359 185
R3057 GNDA.n1358 GNDA.n1357 185
R3058 GNDA.n1356 GNDA.n1355 185
R3059 GNDA.n1354 GNDA.n1353 185
R3060 GNDA.n1389 GNDA.n1388 185
R3061 GNDA.n1386 GNDA.n1385 185
R3062 GNDA.n1384 GNDA.n1383 185
R3063 GNDA.n1382 GNDA.n1381 185
R3064 GNDA.n1380 GNDA.n1379 185
R3065 GNDA.n1378 GNDA.n1377 185
R3066 GNDA.n1376 GNDA.n1375 185
R3067 GNDA.n1374 GNDA.n1373 185
R3068 GNDA.n1372 GNDA.n1371 185
R3069 GNDA.n1387 GNDA.n1333 185
R3070 GNDA.n1331 GNDA.n1330 185
R3071 GNDA.n1324 GNDA.n1300 185
R3072 GNDA.n1591 GNDA.n1590 185
R3073 GNDA.n1574 GNDA.n1299 185
R3074 GNDA.n1578 GNDA.n1577 185
R3075 GNDA.n1576 GNDA.n1573 185
R3076 GNDA.n1320 GNDA.n1318 185
R3077 GNDA.n1587 GNDA.n1586 185
R3078 GNDA.n696 GNDA.n695 185
R3079 GNDA.n698 GNDA.n697 185
R3080 GNDA.n700 GNDA.n699 185
R3081 GNDA.n702 GNDA.n701 185
R3082 GNDA.n704 GNDA.n703 185
R3083 GNDA.n706 GNDA.n705 185
R3084 GNDA.n708 GNDA.n707 185
R3085 GNDA.n710 GNDA.n709 185
R3086 GNDA.n711 GNDA.n659 185
R3087 GNDA.n678 GNDA.n677 185
R3088 GNDA.n680 GNDA.n679 185
R3089 GNDA.n682 GNDA.n681 185
R3090 GNDA.n684 GNDA.n683 185
R3091 GNDA.n686 GNDA.n685 185
R3092 GNDA.n688 GNDA.n687 185
R3093 GNDA.n690 GNDA.n689 185
R3094 GNDA.n692 GNDA.n691 185
R3095 GNDA.n694 GNDA.n693 185
R3096 GNDA.n651 GNDA.n637 185
R3097 GNDA.n662 GNDA.n661 185
R3098 GNDA.n664 GNDA.n663 185
R3099 GNDA.n666 GNDA.n665 185
R3100 GNDA.n668 GNDA.n667 185
R3101 GNDA.n670 GNDA.n669 185
R3102 GNDA.n672 GNDA.n671 185
R3103 GNDA.n674 GNDA.n673 185
R3104 GNDA.n676 GNDA.n675 185
R3105 GNDA.n641 GNDA.n638 185
R3106 GNDA.n748 GNDA.n747 185
R3107 GNDA.n721 GNDA.n640 185
R3108 GNDA.n727 GNDA.n726 185
R3109 GNDA.n725 GNDA.n720 185
R3110 GNDA.n734 GNDA.n733 185
R3111 GNDA.n732 GNDA.n719 185
R3112 GNDA.n739 GNDA.n660 185
R3113 GNDA.n744 GNDA.n743 185
R3114 GNDA.n2272 GNDA.n2271 185
R3115 GNDA.n2274 GNDA.n2273 185
R3116 GNDA.n2276 GNDA.n2275 185
R3117 GNDA.n2278 GNDA.n2277 185
R3118 GNDA.n2280 GNDA.n2279 185
R3119 GNDA.n2282 GNDA.n2281 185
R3120 GNDA.n2284 GNDA.n2283 185
R3121 GNDA.n2286 GNDA.n2285 185
R3122 GNDA.n2287 GNDA.n89 185
R3123 GNDA.n2254 GNDA.n2253 185
R3124 GNDA.n2256 GNDA.n2255 185
R3125 GNDA.n2258 GNDA.n2257 185
R3126 GNDA.n2260 GNDA.n2259 185
R3127 GNDA.n2262 GNDA.n2261 185
R3128 GNDA.n2264 GNDA.n2263 185
R3129 GNDA.n2266 GNDA.n2265 185
R3130 GNDA.n2268 GNDA.n2267 185
R3131 GNDA.n2270 GNDA.n2269 185
R3132 GNDA.n2236 GNDA.n2235 185
R3133 GNDA.n2238 GNDA.n2237 185
R3134 GNDA.n2240 GNDA.n2239 185
R3135 GNDA.n2242 GNDA.n2241 185
R3136 GNDA.n2244 GNDA.n2243 185
R3137 GNDA.n2246 GNDA.n2245 185
R3138 GNDA.n2248 GNDA.n2247 185
R3139 GNDA.n2250 GNDA.n2249 185
R3140 GNDA.n2252 GNDA.n2251 185
R3141 GNDA.n2234 GNDA.n2233 185
R3142 GNDA.n2228 GNDA.n2227 185
R3143 GNDA.n2226 GNDA.n2225 185
R3144 GNDA.n2221 GNDA.n2220 185
R3145 GNDA.n2219 GNDA.n2218 185
R3146 GNDA.n2213 GNDA.n2212 185
R3147 GNDA.n2208 GNDA.n93 185
R3148 GNDA.n2291 GNDA.n2290 185
R3149 GNDA.n92 GNDA.n90 185
R3150 GNDA.n912 GNDA.n911 185
R3151 GNDA.n914 GNDA.n913 185
R3152 GNDA.n916 GNDA.n915 185
R3153 GNDA.n918 GNDA.n917 185
R3154 GNDA.n920 GNDA.n919 185
R3155 GNDA.n922 GNDA.n921 185
R3156 GNDA.n924 GNDA.n923 185
R3157 GNDA.n926 GNDA.n925 185
R3158 GNDA.n927 GNDA.n755 185
R3159 GNDA.n894 GNDA.n893 185
R3160 GNDA.n896 GNDA.n895 185
R3161 GNDA.n898 GNDA.n897 185
R3162 GNDA.n900 GNDA.n899 185
R3163 GNDA.n902 GNDA.n901 185
R3164 GNDA.n904 GNDA.n903 185
R3165 GNDA.n906 GNDA.n905 185
R3166 GNDA.n908 GNDA.n907 185
R3167 GNDA.n910 GNDA.n909 185
R3168 GNDA.n876 GNDA.n875 185
R3169 GNDA.n878 GNDA.n877 185
R3170 GNDA.n880 GNDA.n879 185
R3171 GNDA.n882 GNDA.n881 185
R3172 GNDA.n884 GNDA.n883 185
R3173 GNDA.n886 GNDA.n885 185
R3174 GNDA.n888 GNDA.n887 185
R3175 GNDA.n890 GNDA.n889 185
R3176 GNDA.n892 GNDA.n891 185
R3177 GNDA.n874 GNDA.n873 185
R3178 GNDA.n868 GNDA.n867 185
R3179 GNDA.n866 GNDA.n865 185
R3180 GNDA.n861 GNDA.n860 185
R3181 GNDA.n859 GNDA.n858 185
R3182 GNDA.n853 GNDA.n852 185
R3183 GNDA.n848 GNDA.n759 185
R3184 GNDA.n931 GNDA.n930 185
R3185 GNDA.n758 GNDA.n756 185
R3186 GNDA.n1511 GNDA.n1510 185
R3187 GNDA.n1513 GNDA.n1512 185
R3188 GNDA.n1515 GNDA.n1514 185
R3189 GNDA.n1517 GNDA.n1516 185
R3190 GNDA.n1519 GNDA.n1518 185
R3191 GNDA.n1521 GNDA.n1520 185
R3192 GNDA.n1523 GNDA.n1522 185
R3193 GNDA.n1525 GNDA.n1524 185
R3194 GNDA.n1526 GNDA.n425 185
R3195 GNDA.n1493 GNDA.n1492 185
R3196 GNDA.n1495 GNDA.n1494 185
R3197 GNDA.n1497 GNDA.n1496 185
R3198 GNDA.n1499 GNDA.n1498 185
R3199 GNDA.n1501 GNDA.n1500 185
R3200 GNDA.n1503 GNDA.n1502 185
R3201 GNDA.n1505 GNDA.n1504 185
R3202 GNDA.n1507 GNDA.n1506 185
R3203 GNDA.n1509 GNDA.n1508 185
R3204 GNDA.n1475 GNDA.n1474 185
R3205 GNDA.n1477 GNDA.n1476 185
R3206 GNDA.n1479 GNDA.n1478 185
R3207 GNDA.n1481 GNDA.n1480 185
R3208 GNDA.n1483 GNDA.n1482 185
R3209 GNDA.n1485 GNDA.n1484 185
R3210 GNDA.n1487 GNDA.n1486 185
R3211 GNDA.n1489 GNDA.n1488 185
R3212 GNDA.n1491 GNDA.n1490 185
R3213 GNDA.n1473 GNDA.n1472 185
R3214 GNDA.n1463 GNDA.n1462 185
R3215 GNDA.n1461 GNDA.n408 185
R3216 GNDA.n1672 GNDA.n1671 185
R3217 GNDA.n1655 GNDA.n407 185
R3218 GNDA.n1659 GNDA.n1658 185
R3219 GNDA.n1657 GNDA.n1654 185
R3220 GNDA.n428 GNDA.n426 185
R3221 GNDA.n1668 GNDA.n1667 185
R3222 GNDA.n401 GNDA.n400 185
R3223 GNDA.n398 GNDA.n397 185
R3224 GNDA.n1566 GNDA.n1540 185
R3225 GNDA.n1562 GNDA.n1540 185
R3226 GNDA.n1566 GNDA.n1537 185
R3227 GNDA.n1558 GNDA.n1537 185
R3228 GNDA.n2180 GNDA.n2179 185
R3229 GNDA.n2182 GNDA.n2181 185
R3230 GNDA.n2184 GNDA.n2183 185
R3231 GNDA.n2186 GNDA.n2185 185
R3232 GNDA.n2188 GNDA.n2187 185
R3233 GNDA.n2190 GNDA.n2189 185
R3234 GNDA.n2192 GNDA.n2191 185
R3235 GNDA.n2194 GNDA.n2193 185
R3236 GNDA.n2195 GNDA.n20 185
R3237 GNDA.n2162 GNDA.n2161 185
R3238 GNDA.n2164 GNDA.n2163 185
R3239 GNDA.n2166 GNDA.n2165 185
R3240 GNDA.n2168 GNDA.n2167 185
R3241 GNDA.n2170 GNDA.n2169 185
R3242 GNDA.n2172 GNDA.n2171 185
R3243 GNDA.n2174 GNDA.n2173 185
R3244 GNDA.n2176 GNDA.n2175 185
R3245 GNDA.n2178 GNDA.n2177 185
R3246 GNDA.n2144 GNDA.n2143 185
R3247 GNDA.n2146 GNDA.n2145 185
R3248 GNDA.n2148 GNDA.n2147 185
R3249 GNDA.n2150 GNDA.n2149 185
R3250 GNDA.n2152 GNDA.n2151 185
R3251 GNDA.n2154 GNDA.n2153 185
R3252 GNDA.n2156 GNDA.n2155 185
R3253 GNDA.n2158 GNDA.n2157 185
R3254 GNDA.n2160 GNDA.n2159 185
R3255 GNDA.n2142 GNDA.n2141 185
R3256 GNDA.n2136 GNDA.n2135 185
R3257 GNDA.n2131 GNDA.n3 185
R3258 GNDA.n2404 GNDA.n2403 185
R3259 GNDA.n34 GNDA.n2 185
R3260 GNDA.n38 GNDA.n37 185
R3261 GNDA.n36 GNDA.n33 185
R3262 GNDA.n23 GNDA.n21 185
R3263 GNDA.n2400 GNDA.n2399 185
R3264 GNDA.t87 GNDA.t479 182.07
R3265 GNDA.t515 GNDA.t596 182.07
R3266 GNDA.t525 GNDA.t19 182.07
R3267 GNDA.t109 GNDA.t503 182.07
R3268 GNDA.n1150 GNDA.n1149 175.546
R3269 GNDA.n1257 GNDA.n1149 175.546
R3270 GNDA.n1255 GNDA.n1254 175.546
R3271 GNDA.n1251 GNDA.n1250 175.546
R3272 GNDA.n1247 GNDA.n1246 175.546
R3273 GNDA.n1243 GNDA.n1242 175.546
R3274 GNDA.n1239 GNDA.n1151 175.546
R3275 GNDA.n1239 GNDA.n1153 175.546
R3276 GNDA.n1235 GNDA.n1153 175.546
R3277 GNDA.n1235 GNDA.n1156 175.546
R3278 GNDA.n1231 GNDA.n1156 175.546
R3279 GNDA.n1231 GNDA.n1158 175.546
R3280 GNDA.n1227 GNDA.n1158 175.546
R3281 GNDA.n1227 GNDA.n1160 175.546
R3282 GNDA.n1223 GNDA.n1160 175.546
R3283 GNDA.n1223 GNDA.n1162 175.546
R3284 GNDA.n1219 GNDA.n1162 175.546
R3285 GNDA.n58 GNDA.n54 175.546
R3286 GNDA.n2384 GNDA.n2383 175.546
R3287 GNDA.n2310 GNDA.n2309 175.546
R3288 GNDA.n2315 GNDA.n2314 175.546
R3289 GNDA.n2323 GNDA.n2322 175.546
R3290 GNDA.n1179 GNDA.n1164 175.546
R3291 GNDA.n1180 GNDA.n1179 175.546
R3292 GNDA.n1183 GNDA.n1180 175.546
R3293 GNDA.n1184 GNDA.n1183 175.546
R3294 GNDA.n1204 GNDA.n1184 175.546
R3295 GNDA.n1204 GNDA.n1203 175.546
R3296 GNDA.n1203 GNDA.n1187 175.546
R3297 GNDA.n1191 GNDA.n1187 175.546
R3298 GNDA.n1192 GNDA.n1191 175.546
R3299 GNDA.n1192 GNDA.n85 175.546
R3300 GNDA.n2302 GNDA.n85 175.546
R3301 GNDA.n572 GNDA.n571 175.546
R3302 GNDA.n568 GNDA.n567 175.546
R3303 GNDA.n564 GNDA.n563 175.546
R3304 GNDA.n560 GNDA.n559 175.546
R3305 GNDA.n556 GNDA.n555 175.546
R3306 GNDA.n580 GNDA.n579 175.546
R3307 GNDA.n584 GNDA.n583 175.546
R3308 GNDA.n588 GNDA.n587 175.546
R3309 GNDA.n592 GNDA.n591 175.546
R3310 GNDA.n594 GNDA.n554 175.546
R3311 GNDA.n1083 GNDA.n460 175.546
R3312 GNDA.n1079 GNDA.n478 175.546
R3313 GNDA.n508 GNDA.n507 175.546
R3314 GNDA.n511 GNDA.n510 175.546
R3315 GNDA.n522 GNDA.n521 175.546
R3316 GNDA.n993 GNDA.n992 175.546
R3317 GNDA.n544 GNDA.n543 175.546
R3318 GNDA.n1003 GNDA.n1002 175.546
R3319 GNDA.n539 GNDA.n534 175.546
R3320 GNDA.n1012 GNDA.n528 175.546
R3321 GNDA.n1143 GNDA.n1096 175.546
R3322 GNDA.n1141 GNDA.n1140 175.546
R3323 GNDA.n1137 GNDA.n1136 175.546
R3324 GNDA.n1133 GNDA.n1132 175.546
R3325 GNDA.n1129 GNDA.n1128 175.546
R3326 GNDA.n1124 GNDA.n1123 175.546
R3327 GNDA.n1121 GNDA.n1100 175.546
R3328 GNDA.n1117 GNDA.n1116 175.546
R3329 GNDA.n1114 GNDA.n1103 175.546
R3330 GNDA.n1110 GNDA.n1109 175.546
R3331 GNDA.n1820 GNDA.n297 175.546
R3332 GNDA.n304 GNDA.n297 175.546
R3333 GNDA.n1811 GNDA.n304 175.546
R3334 GNDA.n1811 GNDA.n305 175.546
R3335 GNDA.n1807 GNDA.n305 175.546
R3336 GNDA.n1807 GNDA.n308 175.546
R3337 GNDA.n1554 GNDA.n308 175.546
R3338 GNDA.n1554 GNDA.n1545 175.546
R3339 GNDA.n1545 GNDA.n330 175.546
R3340 GNDA.n1745 GNDA.n330 175.546
R3341 GNDA.n1745 GNDA.n331 175.546
R3342 GNDA.n1707 GNDA.n1706 175.546
R3343 GNDA.n361 GNDA.n360 175.546
R3344 GNDA.n1717 GNDA.n1716 175.546
R3345 GNDA.n356 GNDA.n350 175.546
R3346 GNDA.n1726 GNDA.n345 175.546
R3347 GNDA.n1709 GNDA.n362 175.546
R3348 GNDA.n1713 GNDA.n1711 175.546
R3349 GNDA.n1719 GNDA.n358 175.546
R3350 GNDA.n1722 GNDA.n1721 175.546
R3351 GNDA.n1724 GNDA.n353 175.546
R3352 GNDA.n1699 GNDA.n367 175.546
R3353 GNDA.n1695 GNDA.n1694 175.546
R3354 GNDA.n1692 GNDA.n370 175.546
R3355 GNDA.n1688 GNDA.n1687 175.546
R3356 GNDA.n1685 GNDA.n373 175.546
R3357 GNDA.n1321 GNDA.n341 175.546
R3358 GNDA.n1584 GNDA.n1321 175.546
R3359 GNDA.n1584 GNDA.n1322 175.546
R3360 GNDA.n1580 GNDA.n1322 175.546
R3361 GNDA.n1580 GNDA.n1296 175.546
R3362 GNDA.n1593 GNDA.n1296 175.546
R3363 GNDA.n1593 GNDA.n1297 175.546
R3364 GNDA.n1328 GNDA.n1297 175.546
R3365 GNDA.n1328 GNDA.n1323 175.546
R3366 GNDA.n1533 GNDA.n1323 175.546
R3367 GNDA.n1533 GNDA.n437 175.546
R3368 GNDA.n1601 GNDA.n1600 175.546
R3369 GNDA.n1606 GNDA.n1605 175.546
R3370 GNDA.n1612 GNDA.n1611 175.546
R3371 GNDA.n1616 GNDA.n1599 175.546
R3372 GNDA.n1625 GNDA.n442 175.546
R3373 GNDA.n995 GNDA.n545 175.546
R3374 GNDA.n999 GNDA.n997 175.546
R3375 GNDA.n1005 GNDA.n541 175.546
R3376 GNDA.n1008 GNDA.n1007 175.546
R3377 GNDA.n1010 GNDA.n537 175.546
R3378 GNDA.n985 GNDA.n601 175.546
R3379 GNDA.n981 GNDA.n980 175.546
R3380 GNDA.n978 GNDA.n604 175.546
R3381 GNDA.n974 GNDA.n973 175.546
R3382 GNDA.n971 GNDA.n607 175.546
R3383 GNDA.n741 GNDA.n740 175.546
R3384 GNDA.n737 GNDA.n736 175.546
R3385 GNDA.n730 GNDA.n729 175.546
R3386 GNDA.n723 GNDA.n722 175.546
R3387 GNDA.n751 GNDA.n750 175.546
R3388 GNDA.n621 GNDA.n620 175.546
R3389 GNDA.n623 GNDA.n622 175.546
R3390 GNDA.n625 GNDA.n624 175.546
R3391 GNDA.n627 GNDA.n626 175.546
R3392 GNDA.n629 GNDA.n628 175.546
R3393 GNDA.n1215 GNDA.n1178 175.546
R3394 GNDA.n1211 GNDA.n1178 175.546
R3395 GNDA.n1211 GNDA.n1182 175.546
R3396 GNDA.n1207 GNDA.n1182 175.546
R3397 GNDA.n1207 GNDA.n1186 175.546
R3398 GNDA.n1201 GNDA.n1186 175.546
R3399 GNDA.n1201 GNDA.n1200 175.546
R3400 GNDA.n1200 GNDA.n1190 175.546
R3401 GNDA.n1196 GNDA.n1190 175.546
R3402 GNDA.n1196 GNDA.n88 175.546
R3403 GNDA.n2300 GNDA.n88 175.546
R3404 GNDA.n1177 GNDA.n1167 175.546
R3405 GNDA.n1173 GNDA.n1167 175.546
R3406 GNDA.n1173 GNDA.n1169 175.546
R3407 GNDA.n1169 GNDA.n150 175.546
R3408 GNDA.n2021 GNDA.n150 175.546
R3409 GNDA.n2021 GNDA.n147 175.546
R3410 GNDA.n2026 GNDA.n147 175.546
R3411 GNDA.n2026 GNDA.n145 175.546
R3412 GNDA.n2030 GNDA.n145 175.546
R3413 GNDA.n2030 GNDA.n142 175.546
R3414 GNDA.n2074 GNDA.n142 175.546
R3415 GNDA.n2294 GNDA.n2293 175.546
R3416 GNDA.n2210 GNDA.n2209 175.546
R3417 GNDA.n2216 GNDA.n2215 175.546
R3418 GNDA.n2223 GNDA.n2222 175.546
R3419 GNDA.n2231 GNDA.n2230 175.546
R3420 GNDA.n2035 GNDA.n143 175.546
R3421 GNDA.n2036 GNDA.n2035 175.546
R3422 GNDA.n2037 GNDA.n2036 175.546
R3423 GNDA.n2041 GNDA.n2037 175.546
R3424 GNDA.n2042 GNDA.n2041 175.546
R3425 GNDA.n2045 GNDA.n2042 175.546
R3426 GNDA.n2046 GNDA.n2045 175.546
R3427 GNDA.n2047 GNDA.n2046 175.546
R3428 GNDA.n2051 GNDA.n2047 175.546
R3429 GNDA.n2051 GNDA.n112 175.546
R3430 GNDA.n2202 GNDA.n112 175.546
R3431 GNDA.n961 GNDA.n613 175.546
R3432 GNDA.n961 GNDA.n619 175.546
R3433 GNDA.n957 GNDA.n956 175.546
R3434 GNDA.n953 GNDA.n952 175.546
R3435 GNDA.n949 GNDA.n948 175.546
R3436 GNDA.n945 GNDA.n618 175.546
R3437 GNDA.n797 GNDA.n795 175.546
R3438 GNDA.n801 GNDA.n791 175.546
R3439 GNDA.n805 GNDA.n803 175.546
R3440 GNDA.n809 GNDA.n789 175.546
R3441 GNDA.n812 GNDA.n811 175.546
R3442 GNDA.n934 GNDA.n933 175.546
R3443 GNDA.n850 GNDA.n849 175.546
R3444 GNDA.n856 GNDA.n855 175.546
R3445 GNDA.n863 GNDA.n862 175.546
R3446 GNDA.n871 GNDA.n870 175.546
R3447 GNDA.n819 GNDA.n816 175.546
R3448 GNDA.n819 GNDA.n785 175.546
R3449 GNDA.n824 GNDA.n785 175.546
R3450 GNDA.n824 GNDA.n782 175.546
R3451 GNDA.n828 GNDA.n782 175.546
R3452 GNDA.n829 GNDA.n828 175.546
R3453 GNDA.n832 GNDA.n829 175.546
R3454 GNDA.n832 GNDA.n780 175.546
R3455 GNDA.n837 GNDA.n780 175.546
R3456 GNDA.n837 GNDA.n778 175.546
R3457 GNDA.n841 GNDA.n778 175.546
R3458 GNDA.n1602 GNDA.n379 175.546
R3459 GNDA.n1608 GNDA.n1607 175.546
R3460 GNDA.n1614 GNDA.n1613 175.546
R3461 GNDA.n1619 GNDA.n1618 175.546
R3462 GNDA.n1623 GNDA.n1622 175.546
R3463 GNDA.n1414 GNDA.n1410 175.546
R3464 GNDA.n1418 GNDA.n1416 175.546
R3465 GNDA.n1422 GNDA.n1407 175.546
R3466 GNDA.n1425 GNDA.n1424 175.546
R3467 GNDA.n1429 GNDA.n1428 175.546
R3468 GNDA.n1650 GNDA.n429 175.546
R3469 GNDA.n1665 GNDA.n1650 175.546
R3470 GNDA.n1665 GNDA.n1651 175.546
R3471 GNDA.n1661 GNDA.n1651 175.546
R3472 GNDA.n1661 GNDA.n404 175.546
R3473 GNDA.n1674 GNDA.n404 175.546
R3474 GNDA.n1674 GNDA.n405 175.546
R3475 GNDA.n1465 GNDA.n405 175.546
R3476 GNDA.n1465 GNDA.n1392 175.546
R3477 GNDA.n1470 GNDA.n1392 175.546
R3478 GNDA.n1470 GNDA.n1459 175.546
R3479 GNDA.n1435 GNDA.n1403 175.546
R3480 GNDA.n1435 GNDA.n1401 175.546
R3481 GNDA.n1440 GNDA.n1401 175.546
R3482 GNDA.n1440 GNDA.n1399 175.546
R3483 GNDA.n1444 GNDA.n1399 175.546
R3484 GNDA.n1445 GNDA.n1444 175.546
R3485 GNDA.n1447 GNDA.n1445 175.546
R3486 GNDA.n1447 GNDA.n1397 175.546
R3487 GNDA.n1451 GNDA.n1397 175.546
R3488 GNDA.n1451 GNDA.n1395 175.546
R3489 GNDA.n1455 GNDA.n1395 175.546
R3490 GNDA.n2070 GNDA.n2069 175.546
R3491 GNDA.n2069 GNDA.n2034 175.546
R3492 GNDA.n2065 GNDA.n2034 175.546
R3493 GNDA.n2065 GNDA.n2039 175.546
R3494 GNDA.n2061 GNDA.n2039 175.546
R3495 GNDA.n2061 GNDA.n2059 175.546
R3496 GNDA.n2059 GNDA.n2044 175.546
R3497 GNDA.n2055 GNDA.n2044 175.546
R3498 GNDA.n2055 GNDA.n2049 175.546
R3499 GNDA.n2049 GNDA.n115 175.546
R3500 GNDA.n2200 GNDA.n115 175.546
R3501 GNDA.n2079 GNDA.n139 175.546
R3502 GNDA.n2079 GNDA.n137 175.546
R3503 GNDA.n2083 GNDA.n137 175.546
R3504 GNDA.n2083 GNDA.n135 175.546
R3505 GNDA.n2087 GNDA.n135 175.546
R3506 GNDA.n2087 GNDA.n133 175.546
R3507 GNDA.n2091 GNDA.n133 175.546
R3508 GNDA.n2091 GNDA.n131 175.546
R3509 GNDA.n2095 GNDA.n131 175.546
R3510 GNDA.n2095 GNDA.n129 175.546
R3511 GNDA.n2099 GNDA.n129 175.546
R3512 GNDA.n2397 GNDA.n24 175.546
R3513 GNDA.n40 GNDA.n25 175.546
R3514 GNDA.n31 GNDA.n30 175.546
R3515 GNDA.n2133 GNDA.n2132 175.546
R3516 GNDA.n2139 GNDA.n2138 175.546
R3517 GNDA.n2103 GNDA.n127 175.546
R3518 GNDA.n2103 GNDA.n125 175.546
R3519 GNDA.n2108 GNDA.n125 175.546
R3520 GNDA.n2108 GNDA.n122 175.546
R3521 GNDA.n2112 GNDA.n122 175.546
R3522 GNDA.n2113 GNDA.n2112 175.546
R3523 GNDA.n2116 GNDA.n2113 175.546
R3524 GNDA.n2116 GNDA.n120 175.546
R3525 GNDA.n2121 GNDA.n120 175.546
R3526 GNDA.n2121 GNDA.n118 175.546
R3527 GNDA.n2125 GNDA.n118 175.546
R3528 GNDA.n1014 GNDA.n529 173.881
R3529 GNDA.n634 GNDA.t485 172.876
R3530 GNDA.n962 GNDA.t485 172.615
R3531 GNDA.n538 GNDA.n529 171.624
R3532 GNDA.n1277 GNDA.t173 166.898
R3533 GNDA.n1277 GNDA.t175 166.898
R3534 GNDA.n2327 GNDA.n2326 163.333
R3535 GNDA.n1022 GNDA.n498 163.333
R3536 GNDA.n1749 GNDA.n1748 163.333
R3537 GNDA.n1388 GNDA.n1387 163.333
R3538 GNDA.n651 GNDA.n641 163.333
R3539 GNDA.n2235 GNDA.n2234 163.333
R3540 GNDA.n875 GNDA.n874 163.333
R3541 GNDA.n1474 GNDA.n1473 163.333
R3542 GNDA.n2143 GNDA.n2142 163.333
R3543 GNDA.n185 GNDA.n184 161.3
R3544 GNDA.n179 GNDA.n178 161.3
R3545 GNDA.n1220 GNDA.n1163 159.365
R3546 GNDA.n2076 GNDA.n2075 159.365
R3547 GNDA.n1900 GNDA.n1899 157.143
R3548 GNDA.n1176 GNDA.n1163 155.957
R3549 GNDA.n2077 GNDA.n2076 155.957
R3550 GNDA.t82 GNDA.t479 151.725
R3551 GNDA.t87 GNDA.t596 151.725
R3552 GNDA.t515 GNDA.t111 151.725
R3553 GNDA.t525 GNDA.t115 151.725
R3554 GNDA.t109 GNDA.t19 151.725
R3555 GNDA.t50 GNDA.t503 151.725
R3556 GNDA.n2359 GNDA.n2358 150
R3557 GNDA.n2355 GNDA.n2354 150
R3558 GNDA.n2351 GNDA.n2350 150
R3559 GNDA.n2347 GNDA.n2346 150
R3560 GNDA.n2343 GNDA.n2342 150
R3561 GNDA.n2339 GNDA.n2338 150
R3562 GNDA.n2335 GNDA.n2334 150
R3563 GNDA.n2331 GNDA.n2330 150
R3564 GNDA.n2388 GNDA.n2387 150
R3565 GNDA.n2380 GNDA.n64 150
R3566 GNDA.n2312 GNDA.n65 150
R3567 GNDA.n2319 GNDA.n2318 150
R3568 GNDA.n2377 GNDA.n81 150
R3569 GNDA.n2373 GNDA.n2372 150
R3570 GNDA.n2369 GNDA.n2368 150
R3571 GNDA.n2365 GNDA.n2364 150
R3572 GNDA.n1052 GNDA.n488 150
R3573 GNDA.n1048 GNDA.n1046 150
R3574 GNDA.n1044 GNDA.n490 150
R3575 GNDA.n1040 GNDA.n1038 150
R3576 GNDA.n1036 GNDA.n492 150
R3577 GNDA.n1032 GNDA.n1031 150
R3578 GNDA.n1029 GNDA.n495 150
R3579 GNDA.n1025 GNDA.n1024 150
R3580 GNDA.n1074 GNDA.n1073 150
R3581 GNDA.n1076 GNDA.n482 150
R3582 GNDA.n514 GNDA.n503 150
R3583 GNDA.n518 GNDA.n516 150
R3584 GNDA.n1060 GNDA.n486 150
R3585 GNDA.n1064 GNDA.n1062 150
R3586 GNDA.n1068 GNDA.n484 150
R3587 GNDA.n1071 GNDA.n1070 150
R3588 GNDA.n1781 GNDA.n1780 150
R3589 GNDA.n1777 GNDA.n1776 150
R3590 GNDA.n1773 GNDA.n1772 150
R3591 GNDA.n1769 GNDA.n1768 150
R3592 GNDA.n1765 GNDA.n1764 150
R3593 GNDA.n1761 GNDA.n1760 150
R3594 GNDA.n1757 GNDA.n1756 150
R3595 GNDA.n1753 GNDA.n1752 150
R3596 GNDA.n1815 GNDA.n1814 150
R3597 GNDA.n1802 GNDA.n1801 150
R3598 GNDA.n1804 GNDA.n311 150
R3599 GNDA.n1551 GNDA.n1550 150
R3600 GNDA.n1799 GNDA.n327 150
R3601 GNDA.n1795 GNDA.n1794 150
R3602 GNDA.n1791 GNDA.n1790 150
R3603 GNDA.n1787 GNDA.n1786 150
R3604 GNDA.n1357 GNDA.n1356 150
R3605 GNDA.n1361 GNDA.n1360 150
R3606 GNDA.n1365 GNDA.n1364 150
R3607 GNDA.n1369 GNDA.n1368 150
R3608 GNDA.n1373 GNDA.n1372 150
R3609 GNDA.n1377 GNDA.n1376 150
R3610 GNDA.n1381 GNDA.n1380 150
R3611 GNDA.n1385 GNDA.n1384 150
R3612 GNDA.n1587 GNDA.n1318 150
R3613 GNDA.n1577 GNDA.n1576 150
R3614 GNDA.n1590 GNDA.n1299 150
R3615 GNDA.n1330 GNDA.n1300 150
R3616 GNDA.n1349 GNDA.n1348 150
R3617 GNDA.n1345 GNDA.n1344 150
R3618 GNDA.n1341 GNDA.n1340 150
R3619 GNDA.n1337 GNDA.n1317 150
R3620 GNDA.n691 GNDA.n690 150
R3621 GNDA.n687 GNDA.n686 150
R3622 GNDA.n683 GNDA.n682 150
R3623 GNDA.n679 GNDA.n678 150
R3624 GNDA.n675 GNDA.n674 150
R3625 GNDA.n671 GNDA.n670 150
R3626 GNDA.n667 GNDA.n666 150
R3627 GNDA.n663 GNDA.n662 150
R3628 GNDA.n744 GNDA.n660 150
R3629 GNDA.n733 GNDA.n732 150
R3630 GNDA.n726 GNDA.n725 150
R3631 GNDA.n747 GNDA.n640 150
R3632 GNDA.n699 GNDA.n698 150
R3633 GNDA.n703 GNDA.n702 150
R3634 GNDA.n707 GNDA.n706 150
R3635 GNDA.n709 GNDA.n659 150
R3636 GNDA.n2267 GNDA.n2266 150
R3637 GNDA.n2263 GNDA.n2262 150
R3638 GNDA.n2259 GNDA.n2258 150
R3639 GNDA.n2255 GNDA.n2254 150
R3640 GNDA.n2251 GNDA.n2250 150
R3641 GNDA.n2247 GNDA.n2246 150
R3642 GNDA.n2243 GNDA.n2242 150
R3643 GNDA.n2239 GNDA.n2238 150
R3644 GNDA.n2290 GNDA.n92 150
R3645 GNDA.n2212 GNDA.n93 150
R3646 GNDA.n2220 GNDA.n2219 150
R3647 GNDA.n2227 GNDA.n2226 150
R3648 GNDA.n2275 GNDA.n2274 150
R3649 GNDA.n2279 GNDA.n2278 150
R3650 GNDA.n2283 GNDA.n2282 150
R3651 GNDA.n2287 GNDA.n2286 150
R3652 GNDA.n907 GNDA.n906 150
R3653 GNDA.n903 GNDA.n902 150
R3654 GNDA.n899 GNDA.n898 150
R3655 GNDA.n895 GNDA.n894 150
R3656 GNDA.n891 GNDA.n890 150
R3657 GNDA.n887 GNDA.n886 150
R3658 GNDA.n883 GNDA.n882 150
R3659 GNDA.n879 GNDA.n878 150
R3660 GNDA.n930 GNDA.n758 150
R3661 GNDA.n852 GNDA.n759 150
R3662 GNDA.n860 GNDA.n859 150
R3663 GNDA.n867 GNDA.n866 150
R3664 GNDA.n915 GNDA.n914 150
R3665 GNDA.n919 GNDA.n918 150
R3666 GNDA.n923 GNDA.n922 150
R3667 GNDA.n927 GNDA.n926 150
R3668 GNDA.n1506 GNDA.n1505 150
R3669 GNDA.n1502 GNDA.n1501 150
R3670 GNDA.n1498 GNDA.n1497 150
R3671 GNDA.n1494 GNDA.n1493 150
R3672 GNDA.n1490 GNDA.n1489 150
R3673 GNDA.n1486 GNDA.n1485 150
R3674 GNDA.n1482 GNDA.n1481 150
R3675 GNDA.n1478 GNDA.n1477 150
R3676 GNDA.n1668 GNDA.n426 150
R3677 GNDA.n1658 GNDA.n1657 150
R3678 GNDA.n1671 GNDA.n407 150
R3679 GNDA.n1462 GNDA.n408 150
R3680 GNDA.n1514 GNDA.n1513 150
R3681 GNDA.n1518 GNDA.n1517 150
R3682 GNDA.n1522 GNDA.n1521 150
R3683 GNDA.n1524 GNDA.n425 150
R3684 GNDA.n2175 GNDA.n2174 150
R3685 GNDA.n2171 GNDA.n2170 150
R3686 GNDA.n2167 GNDA.n2166 150
R3687 GNDA.n2163 GNDA.n2162 150
R3688 GNDA.n2159 GNDA.n2158 150
R3689 GNDA.n2155 GNDA.n2154 150
R3690 GNDA.n2151 GNDA.n2150 150
R3691 GNDA.n2147 GNDA.n2146 150
R3692 GNDA.n2400 GNDA.n21 150
R3693 GNDA.n37 GNDA.n36 150
R3694 GNDA.n2403 GNDA.n2 150
R3695 GNDA.n2135 GNDA.n3 150
R3696 GNDA.n2183 GNDA.n2182 150
R3697 GNDA.n2187 GNDA.n2186 150
R3698 GNDA.n2191 GNDA.n2190 150
R3699 GNDA.n2193 GNDA.n20 150
R3700 GNDA.n2000 GNDA.n1999 148.017
R3701 GNDA.n2005 GNDA.n2004 148.017
R3702 GNDA.n1881 GNDA.n1880 148.017
R3703 GNDA.n1896 GNDA.n1895 148.017
R3704 GNDA.n295 GNDA.n294 139.077
R3705 GNDA.n334 GNDA.n333 139.077
R3706 GNDA.n336 GNDA.n335 139.077
R3707 GNDA.n338 GNDA.n337 139.077
R3708 GNDA.n432 GNDA.n431 139.077
R3709 GNDA.n434 GNDA.n433 139.077
R3710 GNDA.n436 GNDA.n435 139.077
R3711 GNDA.n1643 GNDA.n1642 139.077
R3712 GNDA.n1641 GNDA.n1640 139.077
R3713 GNDA.n1639 GNDA.n1638 139.077
R3714 GNDA.n2011 GNDA.t166 135.69
R3715 GNDA.n1540 GNDA.n1539 134.268
R3716 GNDA.n1539 GNDA.n1537 134.268
R3717 GNDA.n1088 GNDA.n455 132.721
R3718 GNDA.n1091 GNDA.n1090 132.721
R3719 GNDA.t599 GNDA.t422 131.767
R3720 GNDA.n1646 GNDA.t489 130.001
R3721 GNDA.n1633 GNDA.t560 130.001
R3722 GNDA.n1736 GNDA.t548 130.001
R3723 GNDA.n1741 GNDA.t500 130.001
R3724 GNDA.n1823 GNDA.t523 130.001
R3725 GNDA.n1636 GNDA.t566 130.001
R3726 GNDA.n2303 GNDA.n2302 124.832
R3727 GNDA.n1017 GNDA.n1016 124.832
R3728 GNDA.n1731 GNDA.n1730 124.832
R3729 GNDA.n1733 GNDA.n340 124.832
R3730 GNDA.n1630 GNDA.n1629 124.832
R3731 GNDA.n714 GNDA.n713 124.832
R3732 GNDA.n939 GNDA.n636 124.832
R3733 GNDA.n2300 GNDA.n2299 124.832
R3734 GNDA.n2203 GNDA.n2202 124.832
R3735 GNDA.n941 GNDA.n618 124.832
R3736 GNDA.n440 GNDA.n439 124.832
R3737 GNDA.n2200 GNDA.n2199 124.832
R3738 GNDA.n1979 GNDA.n1977 124.59
R3739 GNDA.n192 GNDA.n190 124.59
R3740 GNDA.n1987 GNDA.n1986 124.028
R3741 GNDA.n1985 GNDA.n1984 124.028
R3742 GNDA.n1983 GNDA.n1982 124.028
R3743 GNDA.n1981 GNDA.n1980 124.028
R3744 GNDA.n1979 GNDA.n1978 124.028
R3745 GNDA.n200 GNDA.n199 124.028
R3746 GNDA.n198 GNDA.n197 124.028
R3747 GNDA.n196 GNDA.n195 124.028
R3748 GNDA.n194 GNDA.n193 124.028
R3749 GNDA.n192 GNDA.n191 124.028
R3750 GNDA.n1826 GNDA.t600 116.073
R3751 GNDA.n2014 GNDA.t135 115.105
R3752 GNDA.n2015 GNDA.t100 114.635
R3753 GNDA.n1826 GNDA.t589 114.635
R3754 GNDA.n1631 GNDA.t559 101.942
R3755 GNDA.n393 GNDA.n387 101.718
R3756 GNDA.n1557 GNDA.n1542 101.718
R3757 GNDA.n1565 GNDA.n1541 101.718
R3758 GNDA.n402 GNDA.n389 101.718
R3759 GNDA.n366 GNDA.t485 47.6748
R3760 GNDA.n1734 GNDA.n339 98.8538
R3761 GNDA.n1904 GNDA.t528 98.8358
R3762 GNDA.t535 GNDA.n163 98.8358
R3763 GNDA.n1266 GNDA.t2 95.0725
R3764 GNDA.n1649 GNDA.n1648 92.6754
R3765 GNDA.n400 GNDA.n392 91.069
R3766 GNDA.n400 GNDA.n399 91.069
R3767 GNDA.n397 GNDA.n390 91.069
R3768 GNDA.n397 GNDA.n396 91.069
R3769 GNDA.n1559 GNDA.n1540 91.069
R3770 GNDA.n1561 GNDA.n1537 91.069
R3771 GNDA.n1276 GNDA.t576 91.035
R3772 GNDA.t499 GNDA.n1743 90.616
R3773 GNDA.t579 GNDA.t134 89.5224
R3774 GNDA.n2008 GNDA.t206 85.4674
R3775 GNDA.n1581 GNDA.t7 84.4377
R3776 GNDA.n2018 GNDA.n152 84.306
R3777 GNDA.t89 GNDA.t57 83.1688
R3778 GNDA.t591 GNDA.t71 82.3782
R3779 GNDA.t574 GNDA.t165 82.3782
R3780 GNDA.n2076 GNDA.n140 80.9821
R3781 GNDA.n1214 GNDA.n1163 80.9821
R3782 GNDA.t148 GNDA.t179 80.5329
R3783 GNDA.t146 GNDA.t143 80.5329
R3784 GNDA.t162 GNDA.t139 80.5329
R3785 GNDA.t161 GNDA.t177 80.5329
R3786 GNDA.t147 GNDA.t138 80.5329
R3787 GNDA.t482 GNDA.t104 80.5329
R3788 GNDA.t56 GNDA.t482 80.5329
R3789 GNDA.t151 GNDA.t56 80.5329
R3790 GNDA.t61 GNDA.t31 80.5329
R3791 GNDA.t183 GNDA.t192 80.5329
R3792 GNDA.t202 GNDA.t197 80.5329
R3793 GNDA.t189 GNDA.t196 80.5329
R3794 GNDA.t187 GNDA.t193 80.5329
R3795 GNDA.t198 GNDA.t190 80.5329
R3796 GNDA.n1325 GNDA.t67 80.3188
R3797 GNDA.t506 GNDA.t572 76.8724
R3798 GNDA.t495 GNDA.t491 76.8724
R3799 GNDA.t541 GNDA.t556 76.8724
R3800 GNDA.t550 GNDA.t553 76.8724
R3801 GNDA.n1238 GNDA.n1154 76.7001
R3802 GNDA.n1238 GNDA.n1237 76.7001
R3803 GNDA.n1237 GNDA.n1236 76.7001
R3804 GNDA.n1236 GNDA.n1155 76.7001
R3805 GNDA.n1230 GNDA.n1155 76.7001
R3806 GNDA.n1229 GNDA.n1228 76.7001
R3807 GNDA.n1228 GNDA.n1159 76.7001
R3808 GNDA.n1222 GNDA.n1159 76.7001
R3809 GNDA.n1222 GNDA.n1221 76.7001
R3810 GNDA.n1221 GNDA.n1220 76.7001
R3811 GNDA.n1176 GNDA.n1175 76.7001
R3812 GNDA.n1175 GNDA.n1174 76.7001
R3813 GNDA.n1174 GNDA.n1168 76.7001
R3814 GNDA.n1168 GNDA.n151 76.7001
R3815 GNDA.n2020 GNDA.n151 76.7001
R3816 GNDA.n2027 GNDA.n146 76.7001
R3817 GNDA.n2028 GNDA.n2027 76.7001
R3818 GNDA.n2029 GNDA.n2028 76.7001
R3819 GNDA.n2029 GNDA.n141 76.7001
R3820 GNDA.n2075 GNDA.n141 76.7001
R3821 GNDA.n2078 GNDA.n2077 76.7001
R3822 GNDA.n2078 GNDA.n136 76.7001
R3823 GNDA.n2084 GNDA.n136 76.7001
R3824 GNDA.n2085 GNDA.n2084 76.7001
R3825 GNDA.n2086 GNDA.n2085 76.7001
R3826 GNDA.n2092 GNDA.n132 76.7001
R3827 GNDA.n2093 GNDA.n2092 76.7001
R3828 GNDA.n2094 GNDA.n2093 76.7001
R3829 GNDA.n2094 GNDA.n128 76.7001
R3830 GNDA.n2100 GNDA.n128 76.7001
R3831 GNDA.n529 GNDA.t485 76.3879
R3832 GNDA.n1263 GNDA.n1262 76.3222
R3833 GNDA.n1257 GNDA.n445 76.3222
R3834 GNDA.n1254 GNDA.n446 76.3222
R3835 GNDA.n1250 GNDA.n447 76.3222
R3836 GNDA.n1246 GNDA.n448 76.3222
R3837 GNDA.n2394 GNDA.n2393 76.3222
R3838 GNDA.n58 GNDA.n53 76.3222
R3839 GNDA.n2383 GNDA.n52 76.3222
R3840 GNDA.n2310 GNDA.n51 76.3222
R3841 GNDA.n2314 GNDA.n50 76.3222
R3842 GNDA.n2323 GNDA.n49 76.3222
R3843 GNDA.n575 GNDA.n450 76.3222
R3844 GNDA.n571 GNDA.n451 76.3222
R3845 GNDA.n567 GNDA.n452 76.3222
R3846 GNDA.n563 GNDA.n453 76.3222
R3847 GNDA.n559 GNDA.n454 76.3222
R3848 GNDA.n555 GNDA.n455 76.3222
R3849 GNDA.n579 GNDA.n549 76.3222
R3850 GNDA.n583 GNDA.n550 76.3222
R3851 GNDA.n587 GNDA.n551 76.3222
R3852 GNDA.n591 GNDA.n552 76.3222
R3853 GNDA.n594 GNDA.n553 76.3222
R3854 GNDA.n599 GNDA.n598 76.3222
R3855 GNDA.n1082 GNDA.n456 76.3222
R3856 GNDA.n1080 GNDA.n460 76.3222
R3857 GNDA.n478 GNDA.n477 76.3222
R3858 GNDA.n508 GNDA.n476 76.3222
R3859 GNDA.n510 GNDA.n475 76.3222
R3860 GNDA.n522 GNDA.n474 76.3222
R3861 GNDA.n547 GNDA.n530 76.3222
R3862 GNDA.n993 GNDA.n531 76.3222
R3863 GNDA.n544 GNDA.n532 76.3222
R3864 GNDA.n1003 GNDA.n533 76.3222
R3865 GNDA.n1013 GNDA.n534 76.3222
R3866 GNDA.n1015 GNDA.n528 76.3222
R3867 GNDA.n1148 GNDA.n1147 76.3222
R3868 GNDA.n1143 GNDA.n1095 76.3222
R3869 GNDA.n1140 GNDA.n1094 76.3222
R3870 GNDA.n1136 GNDA.n1093 76.3222
R3871 GNDA.n1132 GNDA.n1092 76.3222
R3872 GNDA.n1128 GNDA.n1091 76.3222
R3873 GNDA.n1124 GNDA.n1099 76.3222
R3874 GNDA.n1122 GNDA.n1121 76.3222
R3875 GNDA.n1117 GNDA.n1102 76.3222
R3876 GNDA.n1115 GNDA.n1114 76.3222
R3877 GNDA.n1110 GNDA.n1105 76.3222
R3878 GNDA.n1108 GNDA.n1107 76.3222
R3879 GNDA.n364 GNDA.n346 76.3222
R3880 GNDA.n1707 GNDA.n347 76.3222
R3881 GNDA.n361 GNDA.n348 76.3222
R3882 GNDA.n1717 GNDA.n349 76.3222
R3883 GNDA.n1727 GNDA.n350 76.3222
R3884 GNDA.n1729 GNDA.n345 76.3222
R3885 GNDA.n1703 GNDA.n1702 76.3222
R3886 GNDA.n1710 GNDA.n1709 76.3222
R3887 GNDA.n1713 GNDA.n1712 76.3222
R3888 GNDA.n1720 GNDA.n1719 76.3222
R3889 GNDA.n1723 GNDA.n1722 76.3222
R3890 GNDA.n354 GNDA.n353 76.3222
R3891 GNDA.n1700 GNDA.n1699 76.3222
R3892 GNDA.n1695 GNDA.n369 76.3222
R3893 GNDA.n1693 GNDA.n1692 76.3222
R3894 GNDA.n1688 GNDA.n372 76.3222
R3895 GNDA.n1686 GNDA.n1685 76.3222
R3896 GNDA.n1681 GNDA.n375 76.3222
R3897 GNDA.n1680 GNDA.n376 76.3222
R3898 GNDA.n1601 GNDA.n1596 76.3222
R3899 GNDA.n1606 GNDA.n1597 76.3222
R3900 GNDA.n1612 GNDA.n1598 76.3222
R3901 GNDA.n1626 GNDA.n1599 76.3222
R3902 GNDA.n1628 GNDA.n442 76.3222
R3903 GNDA.n989 GNDA.n988 76.3222
R3904 GNDA.n996 GNDA.n995 76.3222
R3905 GNDA.n999 GNDA.n998 76.3222
R3906 GNDA.n1006 GNDA.n1005 76.3222
R3907 GNDA.n1009 GNDA.n1008 76.3222
R3908 GNDA.n712 GNDA.n537 76.3222
R3909 GNDA.n986 GNDA.n985 76.3222
R3910 GNDA.n981 GNDA.n603 76.3222
R3911 GNDA.n979 GNDA.n978 76.3222
R3912 GNDA.n974 GNDA.n606 76.3222
R3913 GNDA.n972 GNDA.n971 76.3222
R3914 GNDA.n967 GNDA.n609 76.3222
R3915 GNDA.n715 GNDA.n473 76.3222
R3916 GNDA.n741 GNDA.n472 76.3222
R3917 GNDA.n736 GNDA.n471 76.3222
R3918 GNDA.n729 GNDA.n470 76.3222
R3919 GNDA.n722 GNDA.n469 76.3222
R3920 GNDA.n751 GNDA.n468 76.3222
R3921 GNDA.n966 GNDA.n610 76.3222
R3922 GNDA.n630 GNDA.n621 76.3222
R3923 GNDA.n631 GNDA.n623 76.3222
R3924 GNDA.n632 GNDA.n625 76.3222
R3925 GNDA.n633 GNDA.n627 76.3222
R3926 GNDA.n635 GNDA.n629 76.3222
R3927 GNDA.n2298 GNDA.n48 76.3222
R3928 GNDA.n2293 GNDA.n47 76.3222
R3929 GNDA.n2210 GNDA.n46 76.3222
R3930 GNDA.n2216 GNDA.n45 76.3222
R3931 GNDA.n2222 GNDA.n44 76.3222
R3932 GNDA.n2231 GNDA.n43 76.3222
R3933 GNDA.n964 GNDA.n963 76.3222
R3934 GNDA.n619 GNDA.n614 76.3222
R3935 GNDA.n956 GNDA.n615 76.3222
R3936 GNDA.n952 GNDA.n616 76.3222
R3937 GNDA.n948 GNDA.n617 76.3222
R3938 GNDA.n795 GNDA.n794 76.3222
R3939 GNDA.n796 GNDA.n791 76.3222
R3940 GNDA.n803 GNDA.n802 76.3222
R3941 GNDA.n804 GNDA.n789 76.3222
R3942 GNDA.n811 GNDA.n810 76.3222
R3943 GNDA.n815 GNDA.n787 76.3222
R3944 GNDA.n940 GNDA.n467 76.3222
R3945 GNDA.n933 GNDA.n466 76.3222
R3946 GNDA.n850 GNDA.n465 76.3222
R3947 GNDA.n856 GNDA.n464 76.3222
R3948 GNDA.n862 GNDA.n463 76.3222
R3949 GNDA.n871 GNDA.n462 76.3222
R3950 GNDA.n1678 GNDA.n1677 76.3222
R3951 GNDA.n1602 GNDA.n384 76.3222
R3952 GNDA.n1608 GNDA.n383 76.3222
R3953 GNDA.n1614 GNDA.n382 76.3222
R3954 GNDA.n1619 GNDA.n381 76.3222
R3955 GNDA.n1622 GNDA.n380 76.3222
R3956 GNDA.n1410 GNDA.n1409 76.3222
R3957 GNDA.n1416 GNDA.n1415 76.3222
R3958 GNDA.n1417 GNDA.n1407 76.3222
R3959 GNDA.n1424 GNDA.n1423 76.3222
R3960 GNDA.n1428 GNDA.n1405 76.3222
R3961 GNDA.n1431 GNDA.n1430 76.3222
R3962 GNDA.n2198 GNDA.n42 76.3222
R3963 GNDA.n2397 GNDA.n2396 76.3222
R3964 GNDA.n41 GNDA.n40 76.3222
R3965 GNDA.n30 GNDA.n29 76.3222
R3966 GNDA.n2133 GNDA.n28 76.3222
R3967 GNDA.n2139 GNDA.n27 76.3222
R3968 GNDA.n636 GNDA.n635 76.3222
R3969 GNDA.n633 GNDA.n628 76.3222
R3970 GNDA.n632 GNDA.n626 76.3222
R3971 GNDA.n631 GNDA.n624 76.3222
R3972 GNDA.n630 GNDA.n622 76.3222
R3973 GNDA.n620 GNDA.n610 76.3222
R3974 GNDA.n963 GNDA.n613 76.3222
R3975 GNDA.n957 GNDA.n614 76.3222
R3976 GNDA.n953 GNDA.n615 76.3222
R3977 GNDA.n949 GNDA.n616 76.3222
R3978 GNDA.n945 GNDA.n617 76.3222
R3979 GNDA.n1629 GNDA.n1628 76.3222
R3980 GNDA.n1626 GNDA.n1625 76.3222
R3981 GNDA.n1616 GNDA.n1598 76.3222
R3982 GNDA.n1611 GNDA.n1597 76.3222
R3983 GNDA.n1605 GNDA.n1596 76.3222
R3984 GNDA.n1600 GNDA.n376 76.3222
R3985 GNDA.n1677 GNDA.n379 76.3222
R3986 GNDA.n1607 GNDA.n384 76.3222
R3987 GNDA.n1613 GNDA.n383 76.3222
R3988 GNDA.n1618 GNDA.n382 76.3222
R3989 GNDA.n1623 GNDA.n381 76.3222
R3990 GNDA.n440 GNDA.n380 76.3222
R3991 GNDA.n1730 GNDA.n1729 76.3222
R3992 GNDA.n1727 GNDA.n1726 76.3222
R3993 GNDA.n356 GNDA.n349 76.3222
R3994 GNDA.n1716 GNDA.n348 76.3222
R3995 GNDA.n360 GNDA.n347 76.3222
R3996 GNDA.n1706 GNDA.n346 76.3222
R3997 GNDA.n1702 GNDA.n362 76.3222
R3998 GNDA.n1711 GNDA.n1710 76.3222
R3999 GNDA.n1712 GNDA.n358 76.3222
R4000 GNDA.n1721 GNDA.n1720 76.3222
R4001 GNDA.n1724 GNDA.n1723 76.3222
R4002 GNDA.n354 GNDA.n340 76.3222
R4003 GNDA.n1016 GNDA.n1015 76.3222
R4004 GNDA.n1013 GNDA.n1012 76.3222
R4005 GNDA.n539 GNDA.n533 76.3222
R4006 GNDA.n1002 GNDA.n532 76.3222
R4007 GNDA.n543 GNDA.n531 76.3222
R4008 GNDA.n992 GNDA.n530 76.3222
R4009 GNDA.n988 GNDA.n545 76.3222
R4010 GNDA.n997 GNDA.n996 76.3222
R4011 GNDA.n998 GNDA.n541 76.3222
R4012 GNDA.n1007 GNDA.n1006 76.3222
R4013 GNDA.n1010 GNDA.n1009 76.3222
R4014 GNDA.n713 GNDA.n712 76.3222
R4015 GNDA.n599 GNDA.n554 76.3222
R4016 GNDA.n592 GNDA.n553 76.3222
R4017 GNDA.n588 GNDA.n552 76.3222
R4018 GNDA.n584 GNDA.n551 76.3222
R4019 GNDA.n580 GNDA.n550 76.3222
R4020 GNDA.n576 GNDA.n549 76.3222
R4021 GNDA.n609 GNDA.n607 76.3222
R4022 GNDA.n973 GNDA.n972 76.3222
R4023 GNDA.n606 GNDA.n604 76.3222
R4024 GNDA.n980 GNDA.n979 76.3222
R4025 GNDA.n603 GNDA.n601 76.3222
R4026 GNDA.n987 GNDA.n986 76.3222
R4027 GNDA.n812 GNDA.n787 76.3222
R4028 GNDA.n810 GNDA.n809 76.3222
R4029 GNDA.n805 GNDA.n804 76.3222
R4030 GNDA.n802 GNDA.n801 76.3222
R4031 GNDA.n797 GNDA.n796 76.3222
R4032 GNDA.n794 GNDA.n612 76.3222
R4033 GNDA.n2394 GNDA.n54 76.3222
R4034 GNDA.n2384 GNDA.n53 76.3222
R4035 GNDA.n2309 GNDA.n52 76.3222
R4036 GNDA.n2315 GNDA.n51 76.3222
R4037 GNDA.n2322 GNDA.n50 76.3222
R4038 GNDA.n2304 GNDA.n49 76.3222
R4039 GNDA.n2294 GNDA.n48 76.3222
R4040 GNDA.n2209 GNDA.n47 76.3222
R4041 GNDA.n2215 GNDA.n46 76.3222
R4042 GNDA.n2223 GNDA.n45 76.3222
R4043 GNDA.n2230 GNDA.n44 76.3222
R4044 GNDA.n2204 GNDA.n43 76.3222
R4045 GNDA.n42 GNDA.n24 76.3222
R4046 GNDA.n2396 GNDA.n25 76.3222
R4047 GNDA.n41 GNDA.n31 76.3222
R4048 GNDA.n2132 GNDA.n29 76.3222
R4049 GNDA.n2138 GNDA.n28 76.3222
R4050 GNDA.n2128 GNDA.n27 76.3222
R4051 GNDA.n1109 GNDA.n1108 76.3222
R4052 GNDA.n1105 GNDA.n1103 76.3222
R4053 GNDA.n1116 GNDA.n1115 76.3222
R4054 GNDA.n1102 GNDA.n1100 76.3222
R4055 GNDA.n1123 GNDA.n1122 76.3222
R4056 GNDA.n1099 GNDA.n1097 76.3222
R4057 GNDA.n375 GNDA.n373 76.3222
R4058 GNDA.n1687 GNDA.n1686 76.3222
R4059 GNDA.n372 GNDA.n370 76.3222
R4060 GNDA.n1694 GNDA.n1693 76.3222
R4061 GNDA.n369 GNDA.n367 76.3222
R4062 GNDA.n1701 GNDA.n1700 76.3222
R4063 GNDA.n1430 GNDA.n1429 76.3222
R4064 GNDA.n1425 GNDA.n1405 76.3222
R4065 GNDA.n1423 GNDA.n1422 76.3222
R4066 GNDA.n1418 GNDA.n1417 76.3222
R4067 GNDA.n1415 GNDA.n1414 76.3222
R4068 GNDA.n1409 GNDA.n378 76.3222
R4069 GNDA.n1083 GNDA.n1082 76.3222
R4070 GNDA.n1080 GNDA.n1079 76.3222
R4071 GNDA.n507 GNDA.n477 76.3222
R4072 GNDA.n511 GNDA.n476 76.3222
R4073 GNDA.n521 GNDA.n475 76.3222
R4074 GNDA.n1018 GNDA.n474 76.3222
R4075 GNDA.n740 GNDA.n473 76.3222
R4076 GNDA.n737 GNDA.n472 76.3222
R4077 GNDA.n730 GNDA.n471 76.3222
R4078 GNDA.n723 GNDA.n470 76.3222
R4079 GNDA.n750 GNDA.n469 76.3222
R4080 GNDA.n938 GNDA.n468 76.3222
R4081 GNDA.n934 GNDA.n467 76.3222
R4082 GNDA.n849 GNDA.n466 76.3222
R4083 GNDA.n855 GNDA.n465 76.3222
R4084 GNDA.n863 GNDA.n464 76.3222
R4085 GNDA.n870 GNDA.n463 76.3222
R4086 GNDA.n844 GNDA.n462 76.3222
R4087 GNDA.n1148 GNDA.n1096 76.3222
R4088 GNDA.n1141 GNDA.n1095 76.3222
R4089 GNDA.n1137 GNDA.n1094 76.3222
R4090 GNDA.n1133 GNDA.n1093 76.3222
R4091 GNDA.n1129 GNDA.n1092 76.3222
R4092 GNDA.n572 GNDA.n450 76.3222
R4093 GNDA.n568 GNDA.n451 76.3222
R4094 GNDA.n564 GNDA.n452 76.3222
R4095 GNDA.n560 GNDA.n453 76.3222
R4096 GNDA.n556 GNDA.n454 76.3222
R4097 GNDA.n1263 GNDA.n1150 76.3222
R4098 GNDA.n1255 GNDA.n445 76.3222
R4099 GNDA.n1251 GNDA.n446 76.3222
R4100 GNDA.n1247 GNDA.n447 76.3222
R4101 GNDA.n1243 GNDA.n448 76.3222
R4102 GNDA.t108 GNDA.n166 75.8626
R4103 GNDA.t26 GNDA.n1926 75.8626
R4104 GNDA.n2346 GNDA.n70 74.5978
R4105 GNDA.n2343 GNDA.n70 74.5978
R4106 GNDA.n1038 GNDA.n1037 74.5978
R4107 GNDA.n1037 GNDA.n1036 74.5978
R4108 GNDA.n1768 GNDA.n316 74.5978
R4109 GNDA.n1765 GNDA.n316 74.5978
R4110 GNDA.n1369 GNDA.n1306 74.5978
R4111 GNDA.n1372 GNDA.n1306 74.5978
R4112 GNDA.n678 GNDA.n647 74.5978
R4113 GNDA.n675 GNDA.n647 74.5978
R4114 GNDA.n2254 GNDA.n99 74.5978
R4115 GNDA.n2251 GNDA.n99 74.5978
R4116 GNDA.n894 GNDA.n765 74.5978
R4117 GNDA.n891 GNDA.n765 74.5978
R4118 GNDA.n1493 GNDA.n414 74.5978
R4119 GNDA.n1490 GNDA.n414 74.5978
R4120 GNDA.n2162 GNDA.n9 74.5978
R4121 GNDA.n2159 GNDA.n9 74.5978
R4122 GNDA.n1326 GNDA.t124 74.1404
R4123 GNDA.t0 GNDA.t74 71.618
R4124 GNDA.n1583 GNDA.t85 70.0216
R4125 GNDA.t592 GNDA.n2006 69.38
R4126 GNDA.n2388 GNDA.n60 69.3109
R4127 GNDA.n2364 GNDA.n60 69.3109
R4128 GNDA.n1073 GNDA.n1072 69.3109
R4129 GNDA.n1072 GNDA.n1071 69.3109
R4130 GNDA.n1815 GNDA.n301 69.3109
R4131 GNDA.n1786 GNDA.n301 69.3109
R4132 GNDA.n1588 GNDA.n1587 69.3109
R4133 GNDA.n1588 GNDA.n1317 69.3109
R4134 GNDA.n745 GNDA.n744 69.3109
R4135 GNDA.n745 GNDA.n659 69.3109
R4136 GNDA.n2288 GNDA.n92 69.3109
R4137 GNDA.n2288 GNDA.n2287 69.3109
R4138 GNDA.n928 GNDA.n758 69.3109
R4139 GNDA.n928 GNDA.n927 69.3109
R4140 GNDA.n1669 GNDA.n1668 69.3109
R4141 GNDA.n1669 GNDA.n425 69.3109
R4142 GNDA.n2401 GNDA.n2400 69.3109
R4143 GNDA.n2401 GNDA.n20 69.3109
R4144 GNDA.t484 GNDA.n2378 65.8183
R4145 GNDA.t484 GNDA.n79 65.8183
R4146 GNDA.t484 GNDA.n78 65.8183
R4147 GNDA.t484 GNDA.n77 65.8183
R4148 GNDA.t484 GNDA.n68 65.8183
R4149 GNDA.t484 GNDA.n75 65.8183
R4150 GNDA.t484 GNDA.n66 65.8183
R4151 GNDA.t484 GNDA.n76 65.8183
R4152 GNDA.t484 GNDA.n74 65.8183
R4153 GNDA.t484 GNDA.n73 65.8183
R4154 GNDA.t484 GNDA.n72 65.8183
R4155 GNDA.t484 GNDA.n71 65.8183
R4156 GNDA.t484 GNDA.n69 65.8183
R4157 GNDA.t484 GNDA.n67 65.8183
R4158 GNDA.n2379 GNDA.t484 65.8183
R4159 GNDA.t484 GNDA.n61 65.8183
R4160 GNDA.n1055 GNDA.t497 65.8183
R4161 GNDA.n1061 GNDA.t497 65.8183
R4162 GNDA.n1063 GNDA.t497 65.8183
R4163 GNDA.n1069 GNDA.t497 65.8183
R4164 GNDA.n1039 GNDA.t497 65.8183
R4165 GNDA.n1045 GNDA.t497 65.8183
R4166 GNDA.n1047 GNDA.t497 65.8183
R4167 GNDA.n1053 GNDA.t497 65.8183
R4168 GNDA.n1023 GNDA.t497 65.8183
R4169 GNDA.n497 GNDA.t497 65.8183
R4170 GNDA.n1030 GNDA.t497 65.8183
R4171 GNDA.n494 GNDA.t497 65.8183
R4172 GNDA.n517 GNDA.t497 65.8183
R4173 GNDA.n515 GNDA.t497 65.8183
R4174 GNDA.n502 GNDA.t497 65.8183
R4175 GNDA.n1075 GNDA.t497 65.8183
R4176 GNDA.t486 GNDA.n1800 65.8183
R4177 GNDA.t486 GNDA.n325 65.8183
R4178 GNDA.t486 GNDA.n324 65.8183
R4179 GNDA.t486 GNDA.n323 65.8183
R4180 GNDA.t486 GNDA.n314 65.8183
R4181 GNDA.t486 GNDA.n321 65.8183
R4182 GNDA.t486 GNDA.n312 65.8183
R4183 GNDA.t486 GNDA.n322 65.8183
R4184 GNDA.t486 GNDA.n320 65.8183
R4185 GNDA.t486 GNDA.n319 65.8183
R4186 GNDA.t486 GNDA.n318 65.8183
R4187 GNDA.t486 GNDA.n317 65.8183
R4188 GNDA.t486 GNDA.n315 65.8183
R4189 GNDA.t486 GNDA.n313 65.8183
R4190 GNDA.n1803 GNDA.t486 65.8183
R4191 GNDA.t486 GNDA.n302 65.8183
R4192 GNDA.t518 GNDA.n1316 65.8183
R4193 GNDA.t518 GNDA.n1315 65.8183
R4194 GNDA.t518 GNDA.n1314 65.8183
R4195 GNDA.t518 GNDA.n1313 65.8183
R4196 GNDA.t518 GNDA.n1304 65.8183
R4197 GNDA.t518 GNDA.n1311 65.8183
R4198 GNDA.t518 GNDA.n1302 65.8183
R4199 GNDA.t518 GNDA.n1312 65.8183
R4200 GNDA.t518 GNDA.n1310 65.8183
R4201 GNDA.t518 GNDA.n1309 65.8183
R4202 GNDA.t518 GNDA.n1308 65.8183
R4203 GNDA.t518 GNDA.n1307 65.8183
R4204 GNDA.t518 GNDA.n1305 65.8183
R4205 GNDA.n1589 GNDA.t518 65.8183
R4206 GNDA.t518 GNDA.n1303 65.8183
R4207 GNDA.t518 GNDA.n1301 65.8183
R4208 GNDA.t493 GNDA.n658 65.8183
R4209 GNDA.t493 GNDA.n657 65.8183
R4210 GNDA.t493 GNDA.n656 65.8183
R4211 GNDA.t493 GNDA.n655 65.8183
R4212 GNDA.t493 GNDA.n646 65.8183
R4213 GNDA.t493 GNDA.n653 65.8183
R4214 GNDA.t493 GNDA.n643 65.8183
R4215 GNDA.t493 GNDA.n654 65.8183
R4216 GNDA.t493 GNDA.n652 65.8183
R4217 GNDA.t493 GNDA.n650 65.8183
R4218 GNDA.t493 GNDA.n649 65.8183
R4219 GNDA.t493 GNDA.n648 65.8183
R4220 GNDA.n746 GNDA.t493 65.8183
R4221 GNDA.t493 GNDA.n645 65.8183
R4222 GNDA.t493 GNDA.n644 65.8183
R4223 GNDA.t493 GNDA.n642 65.8183
R4224 GNDA.t501 GNDA.n109 65.8183
R4225 GNDA.t501 GNDA.n108 65.8183
R4226 GNDA.t501 GNDA.n107 65.8183
R4227 GNDA.t501 GNDA.n106 65.8183
R4228 GNDA.t501 GNDA.n97 65.8183
R4229 GNDA.t501 GNDA.n104 65.8183
R4230 GNDA.t501 GNDA.n94 65.8183
R4231 GNDA.t501 GNDA.n105 65.8183
R4232 GNDA.t501 GNDA.n103 65.8183
R4233 GNDA.t501 GNDA.n102 65.8183
R4234 GNDA.t501 GNDA.n101 65.8183
R4235 GNDA.t501 GNDA.n100 65.8183
R4236 GNDA.t501 GNDA.n98 65.8183
R4237 GNDA.t501 GNDA.n96 65.8183
R4238 GNDA.t501 GNDA.n95 65.8183
R4239 GNDA.n2289 GNDA.t501 65.8183
R4240 GNDA.t517 GNDA.n775 65.8183
R4241 GNDA.t517 GNDA.n774 65.8183
R4242 GNDA.t517 GNDA.n773 65.8183
R4243 GNDA.t517 GNDA.n772 65.8183
R4244 GNDA.t517 GNDA.n763 65.8183
R4245 GNDA.t517 GNDA.n770 65.8183
R4246 GNDA.t517 GNDA.n760 65.8183
R4247 GNDA.t517 GNDA.n771 65.8183
R4248 GNDA.t517 GNDA.n769 65.8183
R4249 GNDA.t517 GNDA.n768 65.8183
R4250 GNDA.t517 GNDA.n767 65.8183
R4251 GNDA.t517 GNDA.n766 65.8183
R4252 GNDA.t517 GNDA.n764 65.8183
R4253 GNDA.t517 GNDA.n762 65.8183
R4254 GNDA.t517 GNDA.n761 65.8183
R4255 GNDA.n929 GNDA.t517 65.8183
R4256 GNDA.t539 GNDA.n424 65.8183
R4257 GNDA.t539 GNDA.n423 65.8183
R4258 GNDA.t539 GNDA.n422 65.8183
R4259 GNDA.t539 GNDA.n421 65.8183
R4260 GNDA.t539 GNDA.n412 65.8183
R4261 GNDA.t539 GNDA.n419 65.8183
R4262 GNDA.t539 GNDA.n410 65.8183
R4263 GNDA.t539 GNDA.n420 65.8183
R4264 GNDA.t539 GNDA.n418 65.8183
R4265 GNDA.t539 GNDA.n417 65.8183
R4266 GNDA.t539 GNDA.n416 65.8183
R4267 GNDA.t539 GNDA.n415 65.8183
R4268 GNDA.t539 GNDA.n413 65.8183
R4269 GNDA.n1670 GNDA.t539 65.8183
R4270 GNDA.t539 GNDA.n411 65.8183
R4271 GNDA.t539 GNDA.n409 65.8183
R4272 GNDA.t513 GNDA.n19 65.8183
R4273 GNDA.t513 GNDA.n18 65.8183
R4274 GNDA.t513 GNDA.n17 65.8183
R4275 GNDA.t513 GNDA.n16 65.8183
R4276 GNDA.t513 GNDA.n7 65.8183
R4277 GNDA.t513 GNDA.n14 65.8183
R4278 GNDA.t513 GNDA.n5 65.8183
R4279 GNDA.t513 GNDA.n15 65.8183
R4280 GNDA.t513 GNDA.n13 65.8183
R4281 GNDA.t513 GNDA.n12 65.8183
R4282 GNDA.t513 GNDA.n11 65.8183
R4283 GNDA.t513 GNDA.n10 65.8183
R4284 GNDA.t513 GNDA.n8 65.8183
R4285 GNDA.n2402 GNDA.t513 65.8183
R4286 GNDA.t513 GNDA.n6 65.8183
R4287 GNDA.t513 GNDA.n4 65.8183
R4288 GNDA.t528 GNDA.t113 64.8799
R4289 GNDA.t113 GNDA.t21 64.8799
R4290 GNDA.t21 GNDA.t45 64.8799
R4291 GNDA.t22 GNDA.t24 64.8799
R4292 GNDA.t535 GNDA.t22 64.8799
R4293 GNDA.t126 GNDA.n307 63.8432
R4294 GNDA.n1582 GNDA.t130 63.8432
R4295 GNDA.n1662 GNDA.t10 63.8432
R4296 GNDA.n1903 GNDA.t529 62.2505
R4297 GNDA.n1933 GNDA.t516 62.2505
R4298 GNDA.n1928 GNDA.t526 62.2505
R4299 GNDA.n169 GNDA.t536 62.2505
R4300 GNDA.n1274 GNDA.t563 62.2505
R4301 GNDA.n1973 GNDA.t510 62.2505
R4302 GNDA.n1905 GNDA.t533 62.2505
R4303 GNDA.n182 GNDA.t483 62.2505
R4304 GNDA.n181 GNDA.t520 62.2505
R4305 GNDA.n176 GNDA.t531 62.2505
R4306 GNDA.n175 GNDA.t512 62.2505
R4307 GNDA.n173 GNDA.t538 62.2505
R4308 GNDA.t79 GNDA.t148 62.2301
R4309 GNDA.t138 GNDA.t169 62.2301
R4310 GNDA.n1927 GNDA.t76 62.2301
R4311 GNDA.t192 GNDA.t181 62.2301
R4312 GNDA.t594 GNDA.t198 62.2301
R4313 GNDA.n1402 GNDA.t485 62.0551
R4314 GNDA.t122 GNDA.n1555 59.7243
R4315 GNDA.n1327 GNDA.t92 59.7243
R4316 GNDA.n1467 GNDA.t12 59.7243
R4317 GNDA.n1998 GNDA.n1997 59.2425
R4318 GNDA.n1988 GNDA.n161 59.2425
R4319 GNDA.n1883 GNDA.n1882 59.2425
R4320 GNDA.n1893 GNDA.n1892 59.2425
R4321 GNDA.n1821 GNDA.t88 58.6946
R4322 GNDA.n1809 GNDA.t590 58.6946
R4323 GNDA.n1544 GNDA.t132 58.6946
R4324 GNDA.n1881 GNDA.n187 58.5695
R4325 GNDA.n1276 GNDA.t151 58.5695
R4326 GNDA.t484 GNDA.n60 57.8461
R4327 GNDA.n1072 GNDA.t497 57.8461
R4328 GNDA.t486 GNDA.n301 57.8461
R4329 GNDA.t518 GNDA.n1588 57.8461
R4330 GNDA.t493 GNDA.n745 57.8461
R4331 GNDA.t501 GNDA.n2288 57.8461
R4332 GNDA.t517 GNDA.n928 57.8461
R4333 GNDA.t539 GNDA.n1669 57.8461
R4334 GNDA.t513 GNDA.n2401 57.8461
R4335 GNDA.t133 GNDA.t69 56.6352
R4336 GNDA.n1569 GNDA.t547 56.6352
R4337 GNDA.t58 GNDA.t54 56.6352
R4338 GNDA.n1242 GNDA.n449 56.3995
R4339 GNDA.n449 GNDA.n55 56.3995
R4340 GNDA.n842 GNDA.n841 56.3995
R4341 GNDA.n1456 GNDA.n1455 56.3995
R4342 GNDA.n1456 GNDA.n1393 56.3995
R4343 GNDA.n843 GNDA.n842 56.3995
R4344 GNDA.n2126 GNDA.n2125 56.3995
R4345 GNDA.n2127 GNDA.n2126 56.3995
R4346 GNDA.n1090 GNDA.n296 56.3995
R4347 GNDA.n1089 GNDA.n1088 56.3995
R4348 GNDA.n817 GNDA.t35 56.1801
R4349 GNDA.n1742 GNDA.n332 55.6055
R4350 GNDA.t484 GNDA.n70 55.2026
R4351 GNDA.n1037 GNDA.t497 55.2026
R4352 GNDA.t486 GNDA.n316 55.2026
R4353 GNDA.t518 GNDA.n1306 55.2026
R4354 GNDA.t493 GNDA.n647 55.2026
R4355 GNDA.t501 GNDA.n99 55.2026
R4356 GNDA.t517 GNDA.n765 55.2026
R4357 GNDA.t539 GNDA.n414 55.2026
R4358 GNDA.t513 GNDA.n9 55.2026
R4359 GNDA.n1893 GNDA.t572 54.909
R4360 GNDA.n1882 GNDA.t495 54.909
R4361 GNDA.n1998 GNDA.t541 54.909
R4362 GNDA.t553 GNDA.n161 54.909
R4363 GNDA.n1536 GNDA.n1535 54.5757
R4364 GNDA.n1647 GNDA.n430 54.5757
R4365 GNDA.t593 GNDA.n1663 54.5757
R4366 GNDA.n1460 GNDA.t91 54.5757
R4367 GNDA.t157 GNDA.n1468 54.5757
R4368 GNDA.t74 GNDA.t592 53.7136
R4369 GNDA.t136 GNDA.t582 53.7136
R4370 GNDA.t110 GNDA.t136 53.7136
R4371 GNDA.t583 GNDA.t48 53.7136
R4372 GNDA.t48 GNDA.t160 53.7136
R4373 GNDA.t134 GNDA.t156 53.7136
R4374 GNDA.n1327 GNDA.t98 53.546
R4375 GNDA.n2361 GNDA.n76 53.3664
R4376 GNDA.n2358 GNDA.n66 53.3664
R4377 GNDA.n2354 GNDA.n75 53.3664
R4378 GNDA.n2350 GNDA.n68 53.3664
R4379 GNDA.n2339 GNDA.n71 53.3664
R4380 GNDA.n2335 GNDA.n72 53.3664
R4381 GNDA.n2331 GNDA.n73 53.3664
R4382 GNDA.n2327 GNDA.n74 53.3664
R4383 GNDA.n2387 GNDA.n61 53.3664
R4384 GNDA.n2380 GNDA.n2379 53.3664
R4385 GNDA.n2312 GNDA.n67 53.3664
R4386 GNDA.n2319 GNDA.n69 53.3664
R4387 GNDA.n2378 GNDA.n2377 53.3664
R4388 GNDA.n81 GNDA.n79 53.3664
R4389 GNDA.n2372 GNDA.n78 53.3664
R4390 GNDA.n2368 GNDA.n77 53.3664
R4391 GNDA.n2378 GNDA.n80 53.3664
R4392 GNDA.n2373 GNDA.n79 53.3664
R4393 GNDA.n2369 GNDA.n78 53.3664
R4394 GNDA.n2365 GNDA.n77 53.3664
R4395 GNDA.n2347 GNDA.n68 53.3664
R4396 GNDA.n2351 GNDA.n75 53.3664
R4397 GNDA.n2355 GNDA.n66 53.3664
R4398 GNDA.n2359 GNDA.n76 53.3664
R4399 GNDA.n2330 GNDA.n74 53.3664
R4400 GNDA.n2334 GNDA.n73 53.3664
R4401 GNDA.n2338 GNDA.n72 53.3664
R4402 GNDA.n2342 GNDA.n71 53.3664
R4403 GNDA.n2326 GNDA.n69 53.3664
R4404 GNDA.n2318 GNDA.n67 53.3664
R4405 GNDA.n2379 GNDA.n65 53.3664
R4406 GNDA.n64 GNDA.n61 53.3664
R4407 GNDA.n1054 GNDA.n1053 53.3664
R4408 GNDA.n1047 GNDA.n488 53.3664
R4409 GNDA.n1046 GNDA.n1045 53.3664
R4410 GNDA.n1039 GNDA.n490 53.3664
R4411 GNDA.n1032 GNDA.n494 53.3664
R4412 GNDA.n1030 GNDA.n1029 53.3664
R4413 GNDA.n1025 GNDA.n497 53.3664
R4414 GNDA.n1023 GNDA.n1022 53.3664
R4415 GNDA.n1075 GNDA.n1074 53.3664
R4416 GNDA.n502 GNDA.n482 53.3664
R4417 GNDA.n515 GNDA.n514 53.3664
R4418 GNDA.n518 GNDA.n517 53.3664
R4419 GNDA.n1055 GNDA.n486 53.3664
R4420 GNDA.n1061 GNDA.n1060 53.3664
R4421 GNDA.n1064 GNDA.n1063 53.3664
R4422 GNDA.n1069 GNDA.n1068 53.3664
R4423 GNDA.n1056 GNDA.n1055 53.3664
R4424 GNDA.n1062 GNDA.n1061 53.3664
R4425 GNDA.n1063 GNDA.n484 53.3664
R4426 GNDA.n1070 GNDA.n1069 53.3664
R4427 GNDA.n1040 GNDA.n1039 53.3664
R4428 GNDA.n1045 GNDA.n1044 53.3664
R4429 GNDA.n1048 GNDA.n1047 53.3664
R4430 GNDA.n1053 GNDA.n1052 53.3664
R4431 GNDA.n1024 GNDA.n1023 53.3664
R4432 GNDA.n497 GNDA.n495 53.3664
R4433 GNDA.n1031 GNDA.n1030 53.3664
R4434 GNDA.n494 GNDA.n492 53.3664
R4435 GNDA.n517 GNDA.n498 53.3664
R4436 GNDA.n516 GNDA.n515 53.3664
R4437 GNDA.n503 GNDA.n502 53.3664
R4438 GNDA.n1076 GNDA.n1075 53.3664
R4439 GNDA.n1783 GNDA.n322 53.3664
R4440 GNDA.n1780 GNDA.n312 53.3664
R4441 GNDA.n1776 GNDA.n321 53.3664
R4442 GNDA.n1772 GNDA.n314 53.3664
R4443 GNDA.n1761 GNDA.n317 53.3664
R4444 GNDA.n1757 GNDA.n318 53.3664
R4445 GNDA.n1753 GNDA.n319 53.3664
R4446 GNDA.n1749 GNDA.n320 53.3664
R4447 GNDA.n1814 GNDA.n302 53.3664
R4448 GNDA.n1803 GNDA.n1802 53.3664
R4449 GNDA.n313 GNDA.n311 53.3664
R4450 GNDA.n1550 GNDA.n315 53.3664
R4451 GNDA.n1800 GNDA.n1799 53.3664
R4452 GNDA.n327 GNDA.n325 53.3664
R4453 GNDA.n1794 GNDA.n324 53.3664
R4454 GNDA.n1790 GNDA.n323 53.3664
R4455 GNDA.n1800 GNDA.n326 53.3664
R4456 GNDA.n1795 GNDA.n325 53.3664
R4457 GNDA.n1791 GNDA.n324 53.3664
R4458 GNDA.n1787 GNDA.n323 53.3664
R4459 GNDA.n1769 GNDA.n314 53.3664
R4460 GNDA.n1773 GNDA.n321 53.3664
R4461 GNDA.n1777 GNDA.n312 53.3664
R4462 GNDA.n1781 GNDA.n322 53.3664
R4463 GNDA.n1752 GNDA.n320 53.3664
R4464 GNDA.n1756 GNDA.n319 53.3664
R4465 GNDA.n1760 GNDA.n318 53.3664
R4466 GNDA.n1764 GNDA.n317 53.3664
R4467 GNDA.n1748 GNDA.n315 53.3664
R4468 GNDA.n1551 GNDA.n313 53.3664
R4469 GNDA.n1804 GNDA.n1803 53.3664
R4470 GNDA.n1801 GNDA.n302 53.3664
R4471 GNDA.n1353 GNDA.n1312 53.3664
R4472 GNDA.n1357 GNDA.n1302 53.3664
R4473 GNDA.n1361 GNDA.n1311 53.3664
R4474 GNDA.n1365 GNDA.n1304 53.3664
R4475 GNDA.n1376 GNDA.n1307 53.3664
R4476 GNDA.n1380 GNDA.n1308 53.3664
R4477 GNDA.n1384 GNDA.n1309 53.3664
R4478 GNDA.n1388 GNDA.n1310 53.3664
R4479 GNDA.n1318 GNDA.n1301 53.3664
R4480 GNDA.n1577 GNDA.n1303 53.3664
R4481 GNDA.n1590 GNDA.n1589 53.3664
R4482 GNDA.n1330 GNDA.n1305 53.3664
R4483 GNDA.n1349 GNDA.n1316 53.3664
R4484 GNDA.n1348 GNDA.n1315 53.3664
R4485 GNDA.n1344 GNDA.n1314 53.3664
R4486 GNDA.n1340 GNDA.n1313 53.3664
R4487 GNDA.n1352 GNDA.n1316 53.3664
R4488 GNDA.n1345 GNDA.n1315 53.3664
R4489 GNDA.n1341 GNDA.n1314 53.3664
R4490 GNDA.n1337 GNDA.n1313 53.3664
R4491 GNDA.n1368 GNDA.n1304 53.3664
R4492 GNDA.n1364 GNDA.n1311 53.3664
R4493 GNDA.n1360 GNDA.n1302 53.3664
R4494 GNDA.n1356 GNDA.n1312 53.3664
R4495 GNDA.n1385 GNDA.n1310 53.3664
R4496 GNDA.n1381 GNDA.n1309 53.3664
R4497 GNDA.n1377 GNDA.n1308 53.3664
R4498 GNDA.n1373 GNDA.n1307 53.3664
R4499 GNDA.n1387 GNDA.n1305 53.3664
R4500 GNDA.n1589 GNDA.n1300 53.3664
R4501 GNDA.n1303 GNDA.n1299 53.3664
R4502 GNDA.n1576 GNDA.n1301 53.3664
R4503 GNDA.n694 GNDA.n654 53.3664
R4504 GNDA.n690 GNDA.n643 53.3664
R4505 GNDA.n686 GNDA.n653 53.3664
R4506 GNDA.n682 GNDA.n646 53.3664
R4507 GNDA.n671 GNDA.n648 53.3664
R4508 GNDA.n667 GNDA.n649 53.3664
R4509 GNDA.n663 GNDA.n650 53.3664
R4510 GNDA.n652 GNDA.n651 53.3664
R4511 GNDA.n660 GNDA.n642 53.3664
R4512 GNDA.n733 GNDA.n644 53.3664
R4513 GNDA.n726 GNDA.n645 53.3664
R4514 GNDA.n747 GNDA.n746 53.3664
R4515 GNDA.n698 GNDA.n658 53.3664
R4516 GNDA.n699 GNDA.n657 53.3664
R4517 GNDA.n703 GNDA.n656 53.3664
R4518 GNDA.n707 GNDA.n655 53.3664
R4519 GNDA.n695 GNDA.n658 53.3664
R4520 GNDA.n702 GNDA.n657 53.3664
R4521 GNDA.n706 GNDA.n656 53.3664
R4522 GNDA.n709 GNDA.n655 53.3664
R4523 GNDA.n679 GNDA.n646 53.3664
R4524 GNDA.n683 GNDA.n653 53.3664
R4525 GNDA.n687 GNDA.n643 53.3664
R4526 GNDA.n691 GNDA.n654 53.3664
R4527 GNDA.n662 GNDA.n652 53.3664
R4528 GNDA.n666 GNDA.n650 53.3664
R4529 GNDA.n670 GNDA.n649 53.3664
R4530 GNDA.n674 GNDA.n648 53.3664
R4531 GNDA.n746 GNDA.n641 53.3664
R4532 GNDA.n645 GNDA.n640 53.3664
R4533 GNDA.n725 GNDA.n644 53.3664
R4534 GNDA.n732 GNDA.n642 53.3664
R4535 GNDA.n2270 GNDA.n105 53.3664
R4536 GNDA.n2266 GNDA.n94 53.3664
R4537 GNDA.n2262 GNDA.n104 53.3664
R4538 GNDA.n2258 GNDA.n97 53.3664
R4539 GNDA.n2247 GNDA.n100 53.3664
R4540 GNDA.n2243 GNDA.n101 53.3664
R4541 GNDA.n2239 GNDA.n102 53.3664
R4542 GNDA.n2235 GNDA.n103 53.3664
R4543 GNDA.n2290 GNDA.n2289 53.3664
R4544 GNDA.n2212 GNDA.n95 53.3664
R4545 GNDA.n2220 GNDA.n96 53.3664
R4546 GNDA.n2227 GNDA.n98 53.3664
R4547 GNDA.n2274 GNDA.n109 53.3664
R4548 GNDA.n2275 GNDA.n108 53.3664
R4549 GNDA.n2279 GNDA.n107 53.3664
R4550 GNDA.n2283 GNDA.n106 53.3664
R4551 GNDA.n2271 GNDA.n109 53.3664
R4552 GNDA.n2278 GNDA.n108 53.3664
R4553 GNDA.n2282 GNDA.n107 53.3664
R4554 GNDA.n2286 GNDA.n106 53.3664
R4555 GNDA.n2255 GNDA.n97 53.3664
R4556 GNDA.n2259 GNDA.n104 53.3664
R4557 GNDA.n2263 GNDA.n94 53.3664
R4558 GNDA.n2267 GNDA.n105 53.3664
R4559 GNDA.n2238 GNDA.n103 53.3664
R4560 GNDA.n2242 GNDA.n102 53.3664
R4561 GNDA.n2246 GNDA.n101 53.3664
R4562 GNDA.n2250 GNDA.n100 53.3664
R4563 GNDA.n2234 GNDA.n98 53.3664
R4564 GNDA.n2226 GNDA.n96 53.3664
R4565 GNDA.n2219 GNDA.n95 53.3664
R4566 GNDA.n2289 GNDA.n93 53.3664
R4567 GNDA.n910 GNDA.n771 53.3664
R4568 GNDA.n906 GNDA.n760 53.3664
R4569 GNDA.n902 GNDA.n770 53.3664
R4570 GNDA.n898 GNDA.n763 53.3664
R4571 GNDA.n887 GNDA.n766 53.3664
R4572 GNDA.n883 GNDA.n767 53.3664
R4573 GNDA.n879 GNDA.n768 53.3664
R4574 GNDA.n875 GNDA.n769 53.3664
R4575 GNDA.n930 GNDA.n929 53.3664
R4576 GNDA.n852 GNDA.n761 53.3664
R4577 GNDA.n860 GNDA.n762 53.3664
R4578 GNDA.n867 GNDA.n764 53.3664
R4579 GNDA.n914 GNDA.n775 53.3664
R4580 GNDA.n915 GNDA.n774 53.3664
R4581 GNDA.n919 GNDA.n773 53.3664
R4582 GNDA.n923 GNDA.n772 53.3664
R4583 GNDA.n911 GNDA.n775 53.3664
R4584 GNDA.n918 GNDA.n774 53.3664
R4585 GNDA.n922 GNDA.n773 53.3664
R4586 GNDA.n926 GNDA.n772 53.3664
R4587 GNDA.n895 GNDA.n763 53.3664
R4588 GNDA.n899 GNDA.n770 53.3664
R4589 GNDA.n903 GNDA.n760 53.3664
R4590 GNDA.n907 GNDA.n771 53.3664
R4591 GNDA.n878 GNDA.n769 53.3664
R4592 GNDA.n882 GNDA.n768 53.3664
R4593 GNDA.n886 GNDA.n767 53.3664
R4594 GNDA.n890 GNDA.n766 53.3664
R4595 GNDA.n874 GNDA.n764 53.3664
R4596 GNDA.n866 GNDA.n762 53.3664
R4597 GNDA.n859 GNDA.n761 53.3664
R4598 GNDA.n929 GNDA.n759 53.3664
R4599 GNDA.n1509 GNDA.n420 53.3664
R4600 GNDA.n1505 GNDA.n410 53.3664
R4601 GNDA.n1501 GNDA.n419 53.3664
R4602 GNDA.n1497 GNDA.n412 53.3664
R4603 GNDA.n1486 GNDA.n415 53.3664
R4604 GNDA.n1482 GNDA.n416 53.3664
R4605 GNDA.n1478 GNDA.n417 53.3664
R4606 GNDA.n1474 GNDA.n418 53.3664
R4607 GNDA.n426 GNDA.n409 53.3664
R4608 GNDA.n1658 GNDA.n411 53.3664
R4609 GNDA.n1671 GNDA.n1670 53.3664
R4610 GNDA.n1462 GNDA.n413 53.3664
R4611 GNDA.n1513 GNDA.n424 53.3664
R4612 GNDA.n1514 GNDA.n423 53.3664
R4613 GNDA.n1518 GNDA.n422 53.3664
R4614 GNDA.n1522 GNDA.n421 53.3664
R4615 GNDA.n1510 GNDA.n424 53.3664
R4616 GNDA.n1517 GNDA.n423 53.3664
R4617 GNDA.n1521 GNDA.n422 53.3664
R4618 GNDA.n1524 GNDA.n421 53.3664
R4619 GNDA.n1494 GNDA.n412 53.3664
R4620 GNDA.n1498 GNDA.n419 53.3664
R4621 GNDA.n1502 GNDA.n410 53.3664
R4622 GNDA.n1506 GNDA.n420 53.3664
R4623 GNDA.n1477 GNDA.n418 53.3664
R4624 GNDA.n1481 GNDA.n417 53.3664
R4625 GNDA.n1485 GNDA.n416 53.3664
R4626 GNDA.n1489 GNDA.n415 53.3664
R4627 GNDA.n1473 GNDA.n413 53.3664
R4628 GNDA.n1670 GNDA.n408 53.3664
R4629 GNDA.n411 GNDA.n407 53.3664
R4630 GNDA.n1657 GNDA.n409 53.3664
R4631 GNDA.n2178 GNDA.n15 53.3664
R4632 GNDA.n2174 GNDA.n5 53.3664
R4633 GNDA.n2170 GNDA.n14 53.3664
R4634 GNDA.n2166 GNDA.n7 53.3664
R4635 GNDA.n2155 GNDA.n10 53.3664
R4636 GNDA.n2151 GNDA.n11 53.3664
R4637 GNDA.n2147 GNDA.n12 53.3664
R4638 GNDA.n2143 GNDA.n13 53.3664
R4639 GNDA.n21 GNDA.n4 53.3664
R4640 GNDA.n37 GNDA.n6 53.3664
R4641 GNDA.n2403 GNDA.n2402 53.3664
R4642 GNDA.n2135 GNDA.n8 53.3664
R4643 GNDA.n2182 GNDA.n19 53.3664
R4644 GNDA.n2183 GNDA.n18 53.3664
R4645 GNDA.n2187 GNDA.n17 53.3664
R4646 GNDA.n2191 GNDA.n16 53.3664
R4647 GNDA.n2179 GNDA.n19 53.3664
R4648 GNDA.n2186 GNDA.n18 53.3664
R4649 GNDA.n2190 GNDA.n17 53.3664
R4650 GNDA.n2193 GNDA.n16 53.3664
R4651 GNDA.n2163 GNDA.n7 53.3664
R4652 GNDA.n2167 GNDA.n14 53.3664
R4653 GNDA.n2171 GNDA.n5 53.3664
R4654 GNDA.n2175 GNDA.n15 53.3664
R4655 GNDA.n2146 GNDA.n13 53.3664
R4656 GNDA.n2150 GNDA.n12 53.3664
R4657 GNDA.n2154 GNDA.n11 53.3664
R4658 GNDA.n2158 GNDA.n10 53.3664
R4659 GNDA.n2142 GNDA.n8 53.3664
R4660 GNDA.n2402 GNDA.n3 53.3664
R4661 GNDA.n6 GNDA.n2 53.3664
R4662 GNDA.n36 GNDA.n4 53.3664
R4663 GNDA.n1735 GNDA.t485 51.4866
R4664 GNDA.n1632 GNDA.t485 51.4866
R4665 GNDA.t83 GNDA.n1968 50.135
R4666 GNDA.n1939 GNDA.t27 50.135
R4667 GNDA.t153 GNDA.n1582 49.4271
R4668 GNDA.n430 GNDA.t114 48.3974
R4669 GNDA.n1914 GNDA.t597 48.0005
R4670 GNDA.n1914 GNDA.t112 48.0005
R4671 GNDA.n1916 GNDA.t159 48.0005
R4672 GNDA.n1916 GNDA.t39 48.0005
R4673 GNDA.n1918 GNDA.t174 48.0005
R4674 GNDA.n1918 GNDA.t176 48.0005
R4675 GNDA.n1920 GNDA.t577 48.0005
R4676 GNDA.n1920 GNDA.t43 48.0005
R4677 GNDA.n1922 GNDA.t116 48.0005
R4678 GNDA.n1922 GNDA.t20 48.0005
R4679 GNDA.n600 GNDA.t485 47.6748
R4680 GNDA.t602 GNDA.t146 47.5879
R4681 GNDA.t177 GNDA.t163 47.5879
R4682 GNDA.t171 GNDA.t49 47.5879
R4683 GNDA.t197 GNDA.t46 47.5879
R4684 GNDA.t580 GNDA.t187 47.5879
R4685 GNDA.t461 GNDA.n332 47.3677
R4686 GNDA.n1897 GNDA.t156 46.9995
R4687 GNDA.t598 GNDA.t522 46.338
R4688 GNDA.t565 GNDA.t33 46.338
R4689 GNDA.n1287 GNDA.n1286 44.0005
R4690 GNDA.n1896 GNDA.n1893 43.9273
R4691 GNDA.n1882 GNDA.n1881 43.9273
R4692 GNDA.t117 GNDA.t82 43.9273
R4693 GNDA.t119 GNDA.t87 43.9273
R4694 GNDA.t3 GNDA.t515 43.9273
R4695 GNDA.t525 GNDA.t584 43.9273
R4696 GNDA.t109 GNDA.t63 43.9273
R4697 GNDA.t50 GNDA.t29 43.9273
R4698 GNDA.t26 GNDA.t17 43.9273
R4699 GNDA.t15 GNDA.t59 43.9273
R4700 GNDA.n1999 GNDA.n1998 43.9273
R4701 GNDA.n2005 GNDA.n161 43.9273
R4702 GNDA.t522 GNDA.n306 43.2488
R4703 GNDA.n1583 GNDA.t153 43.2488
R4704 GNDA.n1663 GNDA.t52 43.2488
R4705 GNDA.n1571 GNDA.t16 42.2191
R4706 GNDA.t485 GNDA.t461 41.1894
R4707 GNDA.t114 GNDA.t485 41.1894
R4708 GNDA.n777 GNDA.t485 40.7582
R4709 GNDA.n1967 GNDA.t570 40.4338
R4710 GNDA.n1940 GNDA.t545 40.4338
R4711 GNDA.n1230 GNDA.t485 40.0547
R4712 GNDA.n2020 GNDA.t485 40.0547
R4713 GNDA.n2086 GNDA.t485 40.0547
R4714 GNDA.t2 GNDA.t1 40.0308
R4715 GNDA.t1 GNDA.t599 40.0308
R4716 GNDA.n1567 GNDA.n1566 39.3903
R4717 GNDA.n1544 GNDA.t128 39.1299
R4718 GNDA.n1595 GNDA.n1594 39.1299
R4719 GNDA.t98 GNDA.n1326 39.1299
R4720 GNDA.n1469 GNDA.t565 39.1299
R4721 GNDA.n1735 GNDA.n1734 38.1002
R4722 GNDA.n1536 GNDA.n1534 38.1002
R4723 GNDA.n1675 GNDA.t91 38.1002
R4724 GNDA.n1469 GNDA.t157 38.1002
R4725 GNDA.n1964 GNDA.n1963 37.5297
R4726 GNDA.n1962 GNDA.n1961 37.5297
R4727 GNDA.n1960 GNDA.n1959 37.5297
R4728 GNDA.n1958 GNDA.n1957 37.5297
R4729 GNDA.n1956 GNDA.n1955 37.5297
R4730 GNDA.n1954 GNDA.n1953 37.5297
R4731 GNDA.n1952 GNDA.n1951 37.5297
R4732 GNDA.n1950 GNDA.n1949 37.5297
R4733 GNDA.n1948 GNDA.n1947 37.5297
R4734 GNDA.n1946 GNDA.n1945 37.5297
R4735 GNDA.n1944 GNDA.n1943 37.5297
R4736 GNDA.n1632 GNDA.n1631 37.0705
R4737 GNDA.t485 GNDA.n1229 36.6459
R4738 GNDA.t485 GNDA.n146 36.6459
R4739 GNDA.t485 GNDA.n132 36.6459
R4740 GNDA.t108 GNDA.t117 36.6062
R4741 GNDA.t82 GNDA.t119 36.6062
R4742 GNDA.t87 GNDA.t3 36.6062
R4743 GNDA.t515 GNDA.t171 36.6062
R4744 GNDA.t94 GNDA.t485 36.0408
R4745 GNDA.t485 GNDA.t65 36.0408
R4746 GNDA.n1938 GNDA.t72 35.3897
R4747 GNDA.n1937 GNDA.t81 35.3897
R4748 GNDA.n1936 GNDA.t14 35.3897
R4749 GNDA.n1935 GNDA.t108 35.3897
R4750 GNDA.t25 GNDA.n1971 35.3897
R4751 GNDA.t44 GNDA.n1970 35.3897
R4752 GNDA.t23 GNDA.n1969 35.3897
R4753 GNDA.n401 GNDA.n154 35.3278
R4754 GNDA.n306 GNDA.t88 33.9813
R4755 GNDA.t590 GNDA.n1808 33.9813
R4756 GNDA.n1570 GNDA.n1569 33.9813
R4757 GNDA.t582 GNDA.t90 33.1236
R4758 GNDA.t160 GNDA.t155 33.1236
R4759 GNDA.n2012 GNDA.n2011 33.1151
R4760 GNDA.n2102 GNDA.n2101 33.0473
R4761 GNDA.n2102 GNDA.n124 33.0473
R4762 GNDA.n2109 GNDA.n124 33.0473
R4763 GNDA.n2110 GNDA.n2109 33.0473
R4764 GNDA.n2111 GNDA.n2110 33.0473
R4765 GNDA.n2115 GNDA.n2114 33.0473
R4766 GNDA.n2115 GNDA.n119 33.0473
R4767 GNDA.n2122 GNDA.n119 33.0473
R4768 GNDA.n2123 GNDA.n2122 33.0473
R4769 GNDA.n2124 GNDA.n2123 33.0473
R4770 GNDA.n2124 GNDA.n117 33.0473
R4771 GNDA.t578 GNDA.n117 33.0473
R4772 GNDA.n818 GNDA.n817 33.0473
R4773 GNDA.n818 GNDA.n784 33.0473
R4774 GNDA.n825 GNDA.n784 33.0473
R4775 GNDA.n826 GNDA.n825 33.0473
R4776 GNDA.n827 GNDA.n826 33.0473
R4777 GNDA.n831 GNDA.n830 33.0473
R4778 GNDA.n831 GNDA.n779 33.0473
R4779 GNDA.n838 GNDA.n779 33.0473
R4780 GNDA.n839 GNDA.n838 33.0473
R4781 GNDA.n840 GNDA.n839 33.0473
R4782 GNDA.n840 GNDA.n777 33.0473
R4783 GNDA.n1436 GNDA.n1402 33.0473
R4784 GNDA.n1437 GNDA.n1436 33.0473
R4785 GNDA.n1439 GNDA.n1437 33.0473
R4786 GNDA.n1439 GNDA.n1438 33.0473
R4787 GNDA.n1438 GNDA.n385 33.0473
R4788 GNDA.n1446 GNDA.n386 33.0473
R4789 GNDA.n1446 GNDA.n1396 33.0473
R4790 GNDA.n1452 GNDA.n1396 33.0473
R4791 GNDA.n1453 GNDA.n1452 33.0473
R4792 GNDA.n1454 GNDA.n1453 33.0473
R4793 GNDA.n1454 GNDA.n156 33.0473
R4794 GNDA.n1556 GNDA.t122 32.9516
R4795 GNDA.t92 GNDA.n1325 32.9516
R4796 GNDA.t12 GNDA.n1466 32.9516
R4797 GNDA.t139 GNDA.t602 32.9456
R4798 GNDA.t163 GNDA.t162 32.9456
R4799 GNDA.n1972 GNDA.t59 32.9456
R4800 GNDA.t46 GNDA.t189 32.9456
R4801 GNDA.t196 GNDA.t580 32.9456
R4802 GNDA.t485 GNDA.n26 32.9056
R4803 GNDA.n461 GNDA.t485 32.9056
R4804 GNDA.n174 GNDA.n173 31.5738
R4805 GNDA.n2000 GNDA.t542 31.1255
R4806 GNDA.n2004 GNDA.t554 31.1255
R4807 GNDA.n1895 GNDA.t573 31.1255
R4808 GNDA.n1880 GNDA.t496 31.1255
R4809 GNDA.n1990 GNDA.n1987 30.8755
R4810 GNDA.n1890 GNDA.n200 30.813
R4811 GNDA.n1903 GNDA.n1902 29.8672
R4812 GNDA.n170 GNDA.n169 29.8672
R4813 GNDA.n1906 GNDA.n1905 29.8672
R4814 GNDA.t27 GNDA.n1938 29.4916
R4815 GNDA.t72 GNDA.n1937 29.4916
R4816 GNDA.t81 GNDA.n1936 29.4916
R4817 GNDA.t14 GNDA.n1935 29.4916
R4818 GNDA.n1971 GNDA.t44 29.4916
R4819 GNDA.n1970 GNDA.t23 29.4916
R4820 GNDA.n1969 GNDA.t83 29.4916
R4821 GNDA.n1810 GNDA.t126 28.8327
R4822 GNDA.t130 GNDA.n1581 28.8327
R4823 GNDA.t10 GNDA.n1652 28.8327
R4824 GNDA.n1810 GNDA.t133 27.803
R4825 GNDA.n1555 GNDA.t587 27.803
R4826 GNDA.n1743 GNDA.t78 27.803
R4827 GNDA.n2363 GNDA.n2362 27.5561
R4828 GNDA.n1057 GNDA.n487 27.5561
R4829 GNDA.n1785 GNDA.n1784 27.5561
R4830 GNDA.n1354 GNDA.n1351 27.5561
R4831 GNDA.n696 GNDA.n693 27.5561
R4832 GNDA.n2272 GNDA.n2269 27.5561
R4833 GNDA.n912 GNDA.n909 27.5561
R4834 GNDA.n1511 GNDA.n1508 27.5561
R4835 GNDA.n2180 GNDA.n2177 27.5561
R4836 GNDA.n2345 GNDA.n2344 26.6672
R4837 GNDA.n1035 GNDA.n491 26.6672
R4838 GNDA.n1767 GNDA.n1766 26.6672
R4839 GNDA.n1371 GNDA.n1370 26.6672
R4840 GNDA.n677 GNDA.n676 26.6672
R4841 GNDA.n2253 GNDA.n2252 26.6672
R4842 GNDA.n893 GNDA.n892 26.6672
R4843 GNDA.n1492 GNDA.n1491 26.6672
R4844 GNDA.n2161 GNDA.n2160 26.6672
R4845 GNDA.t128 GNDA.t587 25.7435
R4846 GNDA.t52 GNDA.t101 25.7435
R4847 GNDA.n1539 GNDA.n1538 25.3679
R4848 GNDA.n1266 GNDA.t588 24.753
R4849 GNDA.n294 GNDA.t127 24.0005
R4850 GNDA.n294 GNDA.t70 24.0005
R4851 GNDA.n333 GNDA.t95 24.0005
R4852 GNDA.n333 GNDA.t123 24.0005
R4853 GNDA.n335 GNDA.t129 24.0005
R4854 GNDA.n335 GNDA.t6 24.0005
R4855 GNDA.n337 GNDA.t86 24.0005
R4856 GNDA.n337 GNDA.t154 24.0005
R4857 GNDA.n431 GNDA.t131 24.0005
R4858 GNDA.n431 GNDA.t8 24.0005
R4859 GNDA.n433 GNDA.t68 24.0005
R4860 GNDA.n433 GNDA.t93 24.0005
R4861 GNDA.n435 GNDA.t99 24.0005
R4862 GNDA.n435 GNDA.t125 24.0005
R4863 GNDA.n1642 GNDA.t97 24.0005
R4864 GNDA.n1642 GNDA.t53 24.0005
R4865 GNDA.n1640 GNDA.t11 24.0005
R4866 GNDA.n1640 GNDA.t66 24.0005
R4867 GNDA.n1638 GNDA.t55 24.0005
R4868 GNDA.n1638 GNDA.t13 24.0005
R4869 GNDA.t84 GNDA.t89 23.7629
R4870 GNDA.t588 GNDA.t84 23.7629
R4871 GNDA.n1648 GNDA.t121 23.6841
R4872 GNDA.t101 GNDA.n1662 23.6841
R4873 GNDA.n1466 GNDA.t58 23.6841
R4874 GNDA.t85 GNDA.n1570 22.6544
R4875 GNDA.n1664 GNDA.t96 22.6544
R4876 GNDA.n2111 GNDA.t485 22.3989
R4877 GNDA.n827 GNDA.t485 22.3989
R4878 GNDA.t485 GNDA.n385 22.3989
R4879 GNDA.t75 GNDA.t525 21.9639
R4880 GNDA.t28 GNDA.t109 21.9639
R4881 GNDA.t34 GNDA.t50 21.9639
R4882 GNDA.t51 GNDA.t26 21.9639
R4883 GNDA.t509 GNDA.t15 21.9639
R4884 GNDA.n1827 GNDA.n1825 21.8755
R4885 GNDA.n2016 GNDA.n2015 21.0192
R4886 GNDA.n1646 GNDA.n1645 20.8233
R4887 GNDA.n1634 GNDA.n1633 20.8233
R4888 GNDA.n1737 GNDA.n1736 20.8233
R4889 GNDA.n1741 GNDA.n1740 20.8233
R4890 GNDA.n1824 GNDA.n1823 20.8233
R4891 GNDA.n1637 GNDA.n1636 20.8233
R4892 GNDA.n1564 GNDA.t485 20.5949
R4893 GNDA.n1564 GNDA.t575 20.5949
R4894 GNDA.t78 GNDA.n1742 20.5949
R4895 GNDA.t121 GNDA.n1647 20.5949
R4896 GNDA.t9 GNDA.n403 20.5949
R4897 GNDA.t485 GNDA.n403 20.5949
R4898 GNDA.t90 GNDA.t0 20.5905
R4899 GNDA.t155 GNDA.t579 20.5905
R4900 GNDA.n1986 GNDA.t185 19.7005
R4901 GNDA.n1986 GNDA.t477 19.7005
R4902 GNDA.n1984 GNDA.t194 19.7005
R4903 GNDA.n1984 GNDA.t200 19.7005
R4904 GNDA.n1982 GNDA.t199 19.7005
R4905 GNDA.n1982 GNDA.t191 19.7005
R4906 GNDA.n1980 GNDA.t201 19.7005
R4907 GNDA.n1980 GNDA.t184 19.7005
R4908 GNDA.n1978 GNDA.t195 19.7005
R4909 GNDA.n1978 GNDA.t186 19.7005
R4910 GNDA.n1977 GNDA.t476 19.7005
R4911 GNDA.n1977 GNDA.t188 19.7005
R4912 GNDA.n199 GNDA.t399 19.7005
R4913 GNDA.n199 GNDA.t144 19.7005
R4914 GNDA.n197 GNDA.t137 19.7005
R4915 GNDA.n197 GNDA.t178 19.7005
R4916 GNDA.n195 GNDA.t150 19.7005
R4917 GNDA.n195 GNDA.t142 19.7005
R4918 GNDA.n193 GNDA.t145 19.7005
R4919 GNDA.n193 GNDA.t141 19.7005
R4920 GNDA.n191 GNDA.t149 19.7005
R4921 GNDA.n191 GNDA.t140 19.7005
R4922 GNDA.n190 GNDA.t180 19.7005
R4923 GNDA.n190 GNDA.t421 19.7005
R4924 GNDA.n1265 GNDA.t485 19.1501
R4925 GNDA.n2023 GNDA.n148 18.5605
R4926 GNDA.t5 GNDA.n1543 18.5355
R4927 GNDA.n1534 GNDA.t124 18.5355
R4928 GNDA.n180 GNDA.n174 18.4151
R4929 GNDA.t165 GNDA.n155 18.3598
R4930 GNDA.t143 GNDA.t79 18.3033
R4931 GNDA.t169 GNDA.t161 18.3033
R4932 GNDA.n1934 GNDA.t104 18.3033
R4933 GNDA.n1276 GNDA.n1275 18.3033
R4934 GNDA.t181 GNDA.t202 18.3033
R4935 GNDA.t193 GNDA.t594 18.3033
R4936 GNDA.n1930 GNDA.n170 18.0922
R4937 GNDA.n814 GNDA.n786 17.5843
R4938 GNDA.n1433 GNDA.n1432 17.5843
R4939 GNDA.n2098 GNDA.n126 17.5843
R4940 GNDA.n1822 GNDA.t485 17.5058
R4941 GNDA.n2008 GNDA.n157 17.5058
R4942 GNDA.n1154 GNDA.t485 17.0449
R4943 GNDA.n1261 GNDA.n1241 16.9379
R4944 GNDA.n577 GNDA.n574 16.9379
R4945 GNDA.n1146 GNDA.n1126 16.9379
R4946 GNDA.n608 GNDA.n111 16.7709
R4947 GNDA.n942 GNDA.n374 16.7709
R4948 GNDA.n526 GNDA.n363 16.7709
R4949 GNDA.n546 GNDA.n84 16.7709
R4950 GNDA.n1994 GNDA.n1993 16.2608
R4951 GNDA.n1992 GNDA.n1991 16.2608
R4952 GNDA.n1887 GNDA.n1886 16.2608
R4953 GNDA.n1889 GNDA.n1888 16.2608
R4954 GNDA.n2376 GNDA.n2363 16.0005
R4955 GNDA.n2376 GNDA.n2375 16.0005
R4956 GNDA.n2375 GNDA.n2374 16.0005
R4957 GNDA.n2374 GNDA.n2371 16.0005
R4958 GNDA.n2371 GNDA.n2370 16.0005
R4959 GNDA.n2370 GNDA.n2367 16.0005
R4960 GNDA.n2367 GNDA.n2366 16.0005
R4961 GNDA.n2366 GNDA.n57 16.0005
R4962 GNDA.n2362 GNDA.n2360 16.0005
R4963 GNDA.n2360 GNDA.n2357 16.0005
R4964 GNDA.n2357 GNDA.n2356 16.0005
R4965 GNDA.n2356 GNDA.n2353 16.0005
R4966 GNDA.n2353 GNDA.n2352 16.0005
R4967 GNDA.n2352 GNDA.n2349 16.0005
R4968 GNDA.n2349 GNDA.n2348 16.0005
R4969 GNDA.n2348 GNDA.n2345 16.0005
R4970 GNDA.n2344 GNDA.n2341 16.0005
R4971 GNDA.n2341 GNDA.n2340 16.0005
R4972 GNDA.n2340 GNDA.n2337 16.0005
R4973 GNDA.n2337 GNDA.n2336 16.0005
R4974 GNDA.n2336 GNDA.n2333 16.0005
R4975 GNDA.n2333 GNDA.n2332 16.0005
R4976 GNDA.n2332 GNDA.n2329 16.0005
R4977 GNDA.n2329 GNDA.n2328 16.0005
R4978 GNDA.n1058 GNDA.n1057 16.0005
R4979 GNDA.n1059 GNDA.n1058 16.0005
R4980 GNDA.n1059 GNDA.n485 16.0005
R4981 GNDA.n1065 GNDA.n485 16.0005
R4982 GNDA.n1066 GNDA.n1065 16.0005
R4983 GNDA.n1067 GNDA.n1066 16.0005
R4984 GNDA.n1067 GNDA.n483 16.0005
R4985 GNDA.n483 GNDA.n458 16.0005
R4986 GNDA.n1051 GNDA.n487 16.0005
R4987 GNDA.n1051 GNDA.n1050 16.0005
R4988 GNDA.n1050 GNDA.n1049 16.0005
R4989 GNDA.n1049 GNDA.n489 16.0005
R4990 GNDA.n1043 GNDA.n489 16.0005
R4991 GNDA.n1043 GNDA.n1042 16.0005
R4992 GNDA.n1042 GNDA.n1041 16.0005
R4993 GNDA.n1041 GNDA.n491 16.0005
R4994 GNDA.n1035 GNDA.n1034 16.0005
R4995 GNDA.n1034 GNDA.n1033 16.0005
R4996 GNDA.n1033 GNDA.n493 16.0005
R4997 GNDA.n1028 GNDA.n493 16.0005
R4998 GNDA.n1028 GNDA.n1027 16.0005
R4999 GNDA.n1027 GNDA.n1026 16.0005
R5000 GNDA.n1026 GNDA.n496 16.0005
R5001 GNDA.n1021 GNDA.n496 16.0005
R5002 GNDA.n1798 GNDA.n1785 16.0005
R5003 GNDA.n1798 GNDA.n1797 16.0005
R5004 GNDA.n1797 GNDA.n1796 16.0005
R5005 GNDA.n1796 GNDA.n1793 16.0005
R5006 GNDA.n1793 GNDA.n1792 16.0005
R5007 GNDA.n1792 GNDA.n1789 16.0005
R5008 GNDA.n1789 GNDA.n1788 16.0005
R5009 GNDA.n1788 GNDA.n299 16.0005
R5010 GNDA.n1784 GNDA.n1782 16.0005
R5011 GNDA.n1782 GNDA.n1779 16.0005
R5012 GNDA.n1779 GNDA.n1778 16.0005
R5013 GNDA.n1778 GNDA.n1775 16.0005
R5014 GNDA.n1775 GNDA.n1774 16.0005
R5015 GNDA.n1774 GNDA.n1771 16.0005
R5016 GNDA.n1771 GNDA.n1770 16.0005
R5017 GNDA.n1770 GNDA.n1767 16.0005
R5018 GNDA.n1766 GNDA.n1763 16.0005
R5019 GNDA.n1763 GNDA.n1762 16.0005
R5020 GNDA.n1762 GNDA.n1759 16.0005
R5021 GNDA.n1759 GNDA.n1758 16.0005
R5022 GNDA.n1758 GNDA.n1755 16.0005
R5023 GNDA.n1755 GNDA.n1754 16.0005
R5024 GNDA.n1754 GNDA.n1751 16.0005
R5025 GNDA.n1751 GNDA.n1750 16.0005
R5026 GNDA.n1351 GNDA.n1350 16.0005
R5027 GNDA.n1350 GNDA.n1347 16.0005
R5028 GNDA.n1347 GNDA.n1346 16.0005
R5029 GNDA.n1346 GNDA.n1343 16.0005
R5030 GNDA.n1343 GNDA.n1342 16.0005
R5031 GNDA.n1342 GNDA.n1339 16.0005
R5032 GNDA.n1339 GNDA.n1338 16.0005
R5033 GNDA.n1338 GNDA.n1336 16.0005
R5034 GNDA.n1355 GNDA.n1354 16.0005
R5035 GNDA.n1358 GNDA.n1355 16.0005
R5036 GNDA.n1359 GNDA.n1358 16.0005
R5037 GNDA.n1362 GNDA.n1359 16.0005
R5038 GNDA.n1363 GNDA.n1362 16.0005
R5039 GNDA.n1366 GNDA.n1363 16.0005
R5040 GNDA.n1367 GNDA.n1366 16.0005
R5041 GNDA.n1370 GNDA.n1367 16.0005
R5042 GNDA.n1374 GNDA.n1371 16.0005
R5043 GNDA.n1375 GNDA.n1374 16.0005
R5044 GNDA.n1378 GNDA.n1375 16.0005
R5045 GNDA.n1379 GNDA.n1378 16.0005
R5046 GNDA.n1382 GNDA.n1379 16.0005
R5047 GNDA.n1383 GNDA.n1382 16.0005
R5048 GNDA.n1386 GNDA.n1383 16.0005
R5049 GNDA.n1389 GNDA.n1386 16.0005
R5050 GNDA.n697 GNDA.n696 16.0005
R5051 GNDA.n700 GNDA.n697 16.0005
R5052 GNDA.n701 GNDA.n700 16.0005
R5053 GNDA.n704 GNDA.n701 16.0005
R5054 GNDA.n705 GNDA.n704 16.0005
R5055 GNDA.n708 GNDA.n705 16.0005
R5056 GNDA.n710 GNDA.n708 16.0005
R5057 GNDA.n711 GNDA.n710 16.0005
R5058 GNDA.n693 GNDA.n692 16.0005
R5059 GNDA.n692 GNDA.n689 16.0005
R5060 GNDA.n689 GNDA.n688 16.0005
R5061 GNDA.n688 GNDA.n685 16.0005
R5062 GNDA.n685 GNDA.n684 16.0005
R5063 GNDA.n684 GNDA.n681 16.0005
R5064 GNDA.n681 GNDA.n680 16.0005
R5065 GNDA.n680 GNDA.n677 16.0005
R5066 GNDA.n676 GNDA.n673 16.0005
R5067 GNDA.n673 GNDA.n672 16.0005
R5068 GNDA.n672 GNDA.n669 16.0005
R5069 GNDA.n669 GNDA.n668 16.0005
R5070 GNDA.n668 GNDA.n665 16.0005
R5071 GNDA.n665 GNDA.n664 16.0005
R5072 GNDA.n664 GNDA.n661 16.0005
R5073 GNDA.n661 GNDA.n637 16.0005
R5074 GNDA.n2273 GNDA.n2272 16.0005
R5075 GNDA.n2276 GNDA.n2273 16.0005
R5076 GNDA.n2277 GNDA.n2276 16.0005
R5077 GNDA.n2280 GNDA.n2277 16.0005
R5078 GNDA.n2281 GNDA.n2280 16.0005
R5079 GNDA.n2284 GNDA.n2281 16.0005
R5080 GNDA.n2285 GNDA.n2284 16.0005
R5081 GNDA.n2285 GNDA.n89 16.0005
R5082 GNDA.n2269 GNDA.n2268 16.0005
R5083 GNDA.n2268 GNDA.n2265 16.0005
R5084 GNDA.n2265 GNDA.n2264 16.0005
R5085 GNDA.n2264 GNDA.n2261 16.0005
R5086 GNDA.n2261 GNDA.n2260 16.0005
R5087 GNDA.n2260 GNDA.n2257 16.0005
R5088 GNDA.n2257 GNDA.n2256 16.0005
R5089 GNDA.n2256 GNDA.n2253 16.0005
R5090 GNDA.n2252 GNDA.n2249 16.0005
R5091 GNDA.n2249 GNDA.n2248 16.0005
R5092 GNDA.n2248 GNDA.n2245 16.0005
R5093 GNDA.n2245 GNDA.n2244 16.0005
R5094 GNDA.n2244 GNDA.n2241 16.0005
R5095 GNDA.n2241 GNDA.n2240 16.0005
R5096 GNDA.n2240 GNDA.n2237 16.0005
R5097 GNDA.n2237 GNDA.n2236 16.0005
R5098 GNDA.n913 GNDA.n912 16.0005
R5099 GNDA.n916 GNDA.n913 16.0005
R5100 GNDA.n917 GNDA.n916 16.0005
R5101 GNDA.n920 GNDA.n917 16.0005
R5102 GNDA.n921 GNDA.n920 16.0005
R5103 GNDA.n924 GNDA.n921 16.0005
R5104 GNDA.n925 GNDA.n924 16.0005
R5105 GNDA.n925 GNDA.n755 16.0005
R5106 GNDA.n909 GNDA.n908 16.0005
R5107 GNDA.n908 GNDA.n905 16.0005
R5108 GNDA.n905 GNDA.n904 16.0005
R5109 GNDA.n904 GNDA.n901 16.0005
R5110 GNDA.n901 GNDA.n900 16.0005
R5111 GNDA.n900 GNDA.n897 16.0005
R5112 GNDA.n897 GNDA.n896 16.0005
R5113 GNDA.n896 GNDA.n893 16.0005
R5114 GNDA.n892 GNDA.n889 16.0005
R5115 GNDA.n889 GNDA.n888 16.0005
R5116 GNDA.n888 GNDA.n885 16.0005
R5117 GNDA.n885 GNDA.n884 16.0005
R5118 GNDA.n884 GNDA.n881 16.0005
R5119 GNDA.n881 GNDA.n880 16.0005
R5120 GNDA.n880 GNDA.n877 16.0005
R5121 GNDA.n877 GNDA.n876 16.0005
R5122 GNDA.n1512 GNDA.n1511 16.0005
R5123 GNDA.n1515 GNDA.n1512 16.0005
R5124 GNDA.n1516 GNDA.n1515 16.0005
R5125 GNDA.n1519 GNDA.n1516 16.0005
R5126 GNDA.n1520 GNDA.n1519 16.0005
R5127 GNDA.n1523 GNDA.n1520 16.0005
R5128 GNDA.n1525 GNDA.n1523 16.0005
R5129 GNDA.n1526 GNDA.n1525 16.0005
R5130 GNDA.n1508 GNDA.n1507 16.0005
R5131 GNDA.n1507 GNDA.n1504 16.0005
R5132 GNDA.n1504 GNDA.n1503 16.0005
R5133 GNDA.n1503 GNDA.n1500 16.0005
R5134 GNDA.n1500 GNDA.n1499 16.0005
R5135 GNDA.n1499 GNDA.n1496 16.0005
R5136 GNDA.n1496 GNDA.n1495 16.0005
R5137 GNDA.n1495 GNDA.n1492 16.0005
R5138 GNDA.n1491 GNDA.n1488 16.0005
R5139 GNDA.n1488 GNDA.n1487 16.0005
R5140 GNDA.n1487 GNDA.n1484 16.0005
R5141 GNDA.n1484 GNDA.n1483 16.0005
R5142 GNDA.n1483 GNDA.n1480 16.0005
R5143 GNDA.n1480 GNDA.n1479 16.0005
R5144 GNDA.n1479 GNDA.n1476 16.0005
R5145 GNDA.n1476 GNDA.n1475 16.0005
R5146 GNDA.n2017 GNDA.n2016 16.0005
R5147 GNDA.n2017 GNDA.n148 16.0005
R5148 GNDA.n2181 GNDA.n2180 16.0005
R5149 GNDA.n2184 GNDA.n2181 16.0005
R5150 GNDA.n2185 GNDA.n2184 16.0005
R5151 GNDA.n2188 GNDA.n2185 16.0005
R5152 GNDA.n2189 GNDA.n2188 16.0005
R5153 GNDA.n2192 GNDA.n2189 16.0005
R5154 GNDA.n2194 GNDA.n2192 16.0005
R5155 GNDA.n2195 GNDA.n2194 16.0005
R5156 GNDA.n2177 GNDA.n2176 16.0005
R5157 GNDA.n2176 GNDA.n2173 16.0005
R5158 GNDA.n2173 GNDA.n2172 16.0005
R5159 GNDA.n2172 GNDA.n2169 16.0005
R5160 GNDA.n2169 GNDA.n2168 16.0005
R5161 GNDA.n2168 GNDA.n2165 16.0005
R5162 GNDA.n2165 GNDA.n2164 16.0005
R5163 GNDA.n2164 GNDA.n2161 16.0005
R5164 GNDA.n2160 GNDA.n2157 16.0005
R5165 GNDA.n2157 GNDA.n2156 16.0005
R5166 GNDA.n2156 GNDA.n2153 16.0005
R5167 GNDA.n2153 GNDA.n2152 16.0005
R5168 GNDA.n2152 GNDA.n2149 16.0005
R5169 GNDA.n2149 GNDA.n2148 16.0005
R5170 GNDA.n2148 GNDA.n2145 16.0005
R5171 GNDA.n2145 GNDA.n2144 16.0005
R5172 GNDA.t132 GNDA.t5 15.4463
R5173 GNDA.t96 GNDA.t593 15.4463
R5174 GNDA.n1939 GNDA.t45 14.7463
R5175 GNDA.n1968 GNDA.t24 14.7463
R5176 GNDA.t49 GNDA.n1934 14.6428
R5177 GNDA.t31 GNDA.t562 14.6428
R5178 GNDA.t76 GNDA.t75 14.6428
R5179 GNDA.t584 GNDA.t28 14.6428
R5180 GNDA.t63 GNDA.t34 14.6428
R5181 GNDA.t29 GNDA.t51 14.6428
R5182 GNDA.t17 GNDA.t509 14.6428
R5183 GNDA.n2395 GNDA.n26 14.555
R5184 GNDA.n1081 GNDA.n461 14.555
R5185 GNDA.n1639 GNDA.n1637 14.363
R5186 GNDA.n2012 GNDA.n154 14.2974
R5187 GNDA.n1907 GNDA.n1906 14.1651
R5188 GNDA.n1902 GNDA.n168 14.0922
R5189 GNDA.n1645 GNDA.n1644 13.8005
R5190 GNDA.n1635 GNDA.n1634 13.8005
R5191 GNDA.n1738 GNDA.n1737 13.8005
R5192 GNDA.n1740 GNDA.n1739 13.8005
R5193 GNDA.n1825 GNDA.n1824 13.8005
R5194 GNDA.n2008 GNDA.t165 13.2192
R5195 GNDA.n1997 GNDA.t557 12.6791
R5196 GNDA.n1988 GNDA.t551 12.6791
R5197 GNDA.n1892 GNDA.t507 12.6791
R5198 GNDA.n1883 GNDA.t492 12.6791
R5199 GNDA.n1808 GNDA.t94 12.3572
R5200 GNDA.n1594 GNDA.t67 12.3572
R5201 GNDA.t54 GNDA.n1460 12.3572
R5202 GNDA.n1913 GNDA.n1910 12.2505
R5203 GNDA.n1568 GNDA.n1567 12.2193
R5204 GNDA.n1261 GNDA.n1260 11.6369
R5205 GNDA.n1260 GNDA.n1259 11.6369
R5206 GNDA.n1259 GNDA.n1258 11.6369
R5207 GNDA.n1258 GNDA.n1256 11.6369
R5208 GNDA.n1256 GNDA.n1253 11.6369
R5209 GNDA.n1253 GNDA.n1252 11.6369
R5210 GNDA.n1252 GNDA.n1249 11.6369
R5211 GNDA.n1249 GNDA.n1248 11.6369
R5212 GNDA.n1248 GNDA.n1245 11.6369
R5213 GNDA.n1245 GNDA.n1244 11.6369
R5214 GNDA.n1241 GNDA.n1240 11.6369
R5215 GNDA.n1240 GNDA.n1152 11.6369
R5216 GNDA.n1234 GNDA.n1152 11.6369
R5217 GNDA.n1234 GNDA.n1233 11.6369
R5218 GNDA.n1233 GNDA.n1232 11.6369
R5219 GNDA.n1232 GNDA.n1157 11.6369
R5220 GNDA.n1226 GNDA.n1157 11.6369
R5221 GNDA.n1226 GNDA.n1225 11.6369
R5222 GNDA.n1225 GNDA.n1224 11.6369
R5223 GNDA.n1224 GNDA.n1161 11.6369
R5224 GNDA.n1218 GNDA.n1161 11.6369
R5225 GNDA.n574 GNDA.n573 11.6369
R5226 GNDA.n573 GNDA.n570 11.6369
R5227 GNDA.n570 GNDA.n569 11.6369
R5228 GNDA.n569 GNDA.n566 11.6369
R5229 GNDA.n566 GNDA.n565 11.6369
R5230 GNDA.n565 GNDA.n562 11.6369
R5231 GNDA.n562 GNDA.n561 11.6369
R5232 GNDA.n561 GNDA.n558 11.6369
R5233 GNDA.n558 GNDA.n557 11.6369
R5234 GNDA.n557 GNDA.n457 11.6369
R5235 GNDA.n578 GNDA.n577 11.6369
R5236 GNDA.n581 GNDA.n578 11.6369
R5237 GNDA.n582 GNDA.n581 11.6369
R5238 GNDA.n585 GNDA.n582 11.6369
R5239 GNDA.n586 GNDA.n585 11.6369
R5240 GNDA.n589 GNDA.n586 11.6369
R5241 GNDA.n590 GNDA.n589 11.6369
R5242 GNDA.n593 GNDA.n590 11.6369
R5243 GNDA.n595 GNDA.n593 11.6369
R5244 GNDA.n596 GNDA.n595 11.6369
R5245 GNDA.n597 GNDA.n596 11.6369
R5246 GNDA.n1146 GNDA.n1145 11.6369
R5247 GNDA.n1145 GNDA.n1144 11.6369
R5248 GNDA.n1144 GNDA.n1142 11.6369
R5249 GNDA.n1142 GNDA.n1139 11.6369
R5250 GNDA.n1139 GNDA.n1138 11.6369
R5251 GNDA.n1138 GNDA.n1135 11.6369
R5252 GNDA.n1135 GNDA.n1134 11.6369
R5253 GNDA.n1134 GNDA.n1131 11.6369
R5254 GNDA.n1131 GNDA.n1130 11.6369
R5255 GNDA.n1130 GNDA.n1127 11.6369
R5256 GNDA.n984 GNDA.n548 11.6369
R5257 GNDA.n984 GNDA.n983 11.6369
R5258 GNDA.n983 GNDA.n982 11.6369
R5259 GNDA.n982 GNDA.n602 11.6369
R5260 GNDA.n977 GNDA.n602 11.6369
R5261 GNDA.n977 GNDA.n976 11.6369
R5262 GNDA.n976 GNDA.n975 11.6369
R5263 GNDA.n975 GNDA.n605 11.6369
R5264 GNDA.n970 GNDA.n605 11.6369
R5265 GNDA.n970 GNDA.n969 11.6369
R5266 GNDA.n969 GNDA.n968 11.6369
R5267 GNDA.n793 GNDA.n792 11.6369
R5268 GNDA.n798 GNDA.n793 11.6369
R5269 GNDA.n799 GNDA.n798 11.6369
R5270 GNDA.n800 GNDA.n799 11.6369
R5271 GNDA.n800 GNDA.n790 11.6369
R5272 GNDA.n806 GNDA.n790 11.6369
R5273 GNDA.n807 GNDA.n806 11.6369
R5274 GNDA.n808 GNDA.n807 11.6369
R5275 GNDA.n808 GNDA.n788 11.6369
R5276 GNDA.n813 GNDA.n788 11.6369
R5277 GNDA.n814 GNDA.n813 11.6369
R5278 GNDA.n820 GNDA.n786 11.6369
R5279 GNDA.n821 GNDA.n820 11.6369
R5280 GNDA.n823 GNDA.n821 11.6369
R5281 GNDA.n823 GNDA.n822 11.6369
R5282 GNDA.n822 GNDA.n783 11.6369
R5283 GNDA.n783 GNDA.n781 11.6369
R5284 GNDA.n833 GNDA.n781 11.6369
R5285 GNDA.n834 GNDA.n833 11.6369
R5286 GNDA.n836 GNDA.n834 11.6369
R5287 GNDA.n836 GNDA.n835 11.6369
R5288 GNDA.n1412 GNDA.n1411 11.6369
R5289 GNDA.n1413 GNDA.n1412 11.6369
R5290 GNDA.n1413 GNDA.n1408 11.6369
R5291 GNDA.n1419 GNDA.n1408 11.6369
R5292 GNDA.n1420 GNDA.n1419 11.6369
R5293 GNDA.n1421 GNDA.n1420 11.6369
R5294 GNDA.n1421 GNDA.n1406 11.6369
R5295 GNDA.n1426 GNDA.n1406 11.6369
R5296 GNDA.n1427 GNDA.n1426 11.6369
R5297 GNDA.n1427 GNDA.n1404 11.6369
R5298 GNDA.n1432 GNDA.n1404 11.6369
R5299 GNDA.n1434 GNDA.n1433 11.6369
R5300 GNDA.n1434 GNDA.n1400 11.6369
R5301 GNDA.n1441 GNDA.n1400 11.6369
R5302 GNDA.n1442 GNDA.n1441 11.6369
R5303 GNDA.n1443 GNDA.n1442 11.6369
R5304 GNDA.n1443 GNDA.n1398 11.6369
R5305 GNDA.n1448 GNDA.n1398 11.6369
R5306 GNDA.n1449 GNDA.n1448 11.6369
R5307 GNDA.n1450 GNDA.n1449 11.6369
R5308 GNDA.n1450 GNDA.n1394 11.6369
R5309 GNDA.n2104 GNDA.n126 11.6369
R5310 GNDA.n2105 GNDA.n2104 11.6369
R5311 GNDA.n2107 GNDA.n2105 11.6369
R5312 GNDA.n2107 GNDA.n2106 11.6369
R5313 GNDA.n2106 GNDA.n123 11.6369
R5314 GNDA.n123 GNDA.n121 11.6369
R5315 GNDA.n2117 GNDA.n121 11.6369
R5316 GNDA.n2118 GNDA.n2117 11.6369
R5317 GNDA.n2120 GNDA.n2118 11.6369
R5318 GNDA.n2120 GNDA.n2119 11.6369
R5319 GNDA.n2080 GNDA.n138 11.6369
R5320 GNDA.n2081 GNDA.n2080 11.6369
R5321 GNDA.n2082 GNDA.n2081 11.6369
R5322 GNDA.n2082 GNDA.n134 11.6369
R5323 GNDA.n2088 GNDA.n134 11.6369
R5324 GNDA.n2089 GNDA.n2088 11.6369
R5325 GNDA.n2090 GNDA.n2089 11.6369
R5326 GNDA.n2090 GNDA.n130 11.6369
R5327 GNDA.n2096 GNDA.n130 11.6369
R5328 GNDA.n2097 GNDA.n2096 11.6369
R5329 GNDA.n2098 GNDA.n2097 11.6369
R5330 GNDA.n1170 GNDA.n1165 11.6369
R5331 GNDA.n1172 GNDA.n1170 11.6369
R5332 GNDA.n1172 GNDA.n1171 11.6369
R5333 GNDA.n1171 GNDA.n149 11.6369
R5334 GNDA.n2022 GNDA.n149 11.6369
R5335 GNDA.n2025 GNDA.n2024 11.6369
R5336 GNDA.n2025 GNDA.n144 11.6369
R5337 GNDA.n2031 GNDA.n144 11.6369
R5338 GNDA.n2032 GNDA.n2031 11.6369
R5339 GNDA.n2073 GNDA.n2032 11.6369
R5340 GNDA.n1698 GNDA.n365 11.6369
R5341 GNDA.n1698 GNDA.n1697 11.6369
R5342 GNDA.n1697 GNDA.n1696 11.6369
R5343 GNDA.n1696 GNDA.n368 11.6369
R5344 GNDA.n1691 GNDA.n368 11.6369
R5345 GNDA.n1691 GNDA.n1690 11.6369
R5346 GNDA.n1690 GNDA.n1689 11.6369
R5347 GNDA.n1689 GNDA.n371 11.6369
R5348 GNDA.n1684 GNDA.n371 11.6369
R5349 GNDA.n1684 GNDA.n1683 11.6369
R5350 GNDA.n1683 GNDA.n1682 11.6369
R5351 GNDA.n1126 GNDA.n1125 11.6369
R5352 GNDA.n1125 GNDA.n1098 11.6369
R5353 GNDA.n1120 GNDA.n1098 11.6369
R5354 GNDA.n1120 GNDA.n1119 11.6369
R5355 GNDA.n1119 GNDA.n1118 11.6369
R5356 GNDA.n1118 GNDA.n1101 11.6369
R5357 GNDA.n1113 GNDA.n1101 11.6369
R5358 GNDA.n1113 GNDA.n1112 11.6369
R5359 GNDA.n1112 GNDA.n1111 11.6369
R5360 GNDA.n1111 GNDA.n1104 11.6369
R5361 GNDA.n1106 GNDA.n1104 11.6369
R5362 GNDA.n2114 GNDA.t485 10.6489
R5363 GNDA.n830 GNDA.t485 10.6489
R5364 GNDA.t485 GNDA.n386 10.6489
R5365 GNDA.n2013 GNDA.n2012 9.95362
R5366 GNDA.n1877 GNDA.n1876 9.71925
R5367 GNDA.n397 GNDA.t207 9.6005
R5368 GNDA.n400 GNDA.t400 9.6005
R5369 GNDA.n1537 GNDA.t423 9.6005
R5370 GNDA.n1540 GNDA.t462 9.6005
R5371 GNDA.n1963 GNDA.t107 9.6005
R5372 GNDA.n1963 GNDA.t569 9.6005
R5373 GNDA.n1961 GNDA.t60 9.6005
R5374 GNDA.n1961 GNDA.t103 9.6005
R5375 GNDA.n1959 GNDA.t30 9.6005
R5376 GNDA.n1959 GNDA.t18 9.6005
R5377 GNDA.n1957 GNDA.t585 9.6005
R5378 GNDA.n1957 GNDA.t64 9.6005
R5379 GNDA.n1955 GNDA.t32 9.6005
R5380 GNDA.n1955 GNDA.t77 9.6005
R5381 GNDA.n1953 GNDA.t152 9.6005
R5382 GNDA.n1953 GNDA.t62 9.6005
R5383 GNDA.n1951 GNDA.t601 9.6005
R5384 GNDA.n1951 GNDA.t586 9.6005
R5385 GNDA.n1949 GNDA.t172 9.6005
R5386 GNDA.n1949 GNDA.t105 9.6005
R5387 GNDA.n1947 GNDA.t120 9.6005
R5388 GNDA.n1947 GNDA.t4 9.6005
R5389 GNDA.n1945 GNDA.t168 9.6005
R5390 GNDA.n1945 GNDA.t118 9.6005
R5391 GNDA.n1943 GNDA.t41 9.6005
R5392 GNDA.n1943 GNDA.t37 9.6005
R5393 GNDA.n1925 GNDA.n1924 9.52967
R5394 GNDA.n1912 GNDA.n1911 9.52967
R5395 GNDA.n2003 GNDA.n2002 9.0005
R5396 GNDA.n1894 GNDA.n172 9.0005
R5397 GNDA.n1827 GNDA.n1826 8.938
R5398 GNDA.n2002 GNDA.n162 8.90675
R5399 GNDA.n83 GNDA.n26 8.60107
R5400 GNDA.n525 GNDA.n461 8.60107
R5401 GNDA.n2014 GNDA.n2013 8.3755
R5402 GNDA.t69 GNDA.n1809 8.23827
R5403 GNDA.t7 GNDA.n1571 8.23827
R5404 GNDA.t65 GNDA.n1675 8.23827
R5405 GNDA.n1976 GNDA.n162 7.46925
R5406 GNDA.n1878 GNDA.n165 7.40675
R5407 GNDA.t73 GNDA.t578 7.34424
R5408 GNDA.n1543 GNDA.t591 7.20855
R5409 GNDA.n1652 GNDA.t9 7.20855
R5410 GNDA.t33 GNDA.n1467 7.20855
R5411 GNDA.n1468 GNDA.n157 7.20855
R5412 GNDA.n1965 GNDA.n162 7.09425
R5413 GNDA.n1942 GNDA.n165 7.03175
R5414 GNDA.n1218 GNDA.n1217 6.72373
R5415 GNDA.n597 GNDA.n546 6.72373
R5416 GNDA.n968 GNDA.n608 6.72373
R5417 GNDA.n2073 GNDA.n2072 6.72373
R5418 GNDA.n1682 GNDA.n374 6.72373
R5419 GNDA.n1106 GNDA.n363 6.72373
R5420 GNDA.n1828 GNDA.n1827 6.42238
R5421 GNDA.n1878 GNDA.n1877 6.313
R5422 GNDA.t35 GNDA.t73 6.24268
R5423 GNDA.n548 GNDA.n546 6.20656
R5424 GNDA.n792 GNDA.n608 6.20656
R5425 GNDA.n1411 GNDA.n374 6.20656
R5426 GNDA.n2072 GNDA.n138 6.20656
R5427 GNDA.n1217 GNDA.n1165 6.20656
R5428 GNDA.n365 GNDA.n363 6.20656
R5429 GNDA.n2013 GNDA.n153 6.188
R5430 GNDA.t485 GNDA.t16 6.17883
R5431 GNDA.n2023 GNDA.n2022 6.07727
R5432 GNDA.n1566 GNDA.n1538 5.81868
R5433 GNDA.n1562 GNDA.n1538 5.81868
R5434 GNDA.n2024 GNDA.n2023 5.5601
R5435 GNDA.n2328 GNDA.n2306 5.51161
R5436 GNDA.n1021 GNDA.n1020 5.51161
R5437 GNDA.n1750 GNDA.n328 5.51161
R5438 GNDA.n1531 GNDA.n1389 5.51161
R5439 GNDA.n753 GNDA.n637 5.51161
R5440 GNDA.n2236 GNDA.n2206 5.51161
R5441 GNDA.n876 GNDA.n846 5.51161
R5442 GNDA.n1475 GNDA.n1390 5.51161
R5443 GNDA.n2144 GNDA.n2130 5.51161
R5444 GNDA.n1910 GNDA.n168 5.5005
R5445 GNDA.n845 GNDA.n776 5.1717
R5446 GNDA.n1458 GNDA.n1457 5.1717
R5447 GNDA.n2129 GNDA.n116 5.1717
R5448 GNDA.t485 GNDA.n1595 5.14911
R5449 GNDA.t488 GNDA.t574 5.14911
R5450 GNDA.n2009 GNDA.n2008 5.14112
R5451 GNDA.n1924 GNDA.n1923 5.063
R5452 GNDA.n1273 GNDA.n164 5.02133
R5453 GNDA.n1975 GNDA.n1974 5.02133
R5454 GNDA.n2002 GNDA.n2001 5.0005
R5455 GNDA.n1879 GNDA.n172 5.0005
R5456 GNDA.n1996 GNDA.n1995 4.91717
R5457 GNDA.n1990 GNDA.n1989 4.91717
R5458 GNDA.n1885 GNDA.n1884 4.91717
R5459 GNDA.n1891 GNDA.n1890 4.91717
R5460 GNDA.n2392 GNDA.n56 4.9157
R5461 GNDA.n1087 GNDA.n1086 4.9157
R5462 GNDA.n1819 GNDA.n298 4.9157
R5463 GNDA.n186 GNDA.n185 4.86508
R5464 GNDA.n180 GNDA.n179 4.86508
R5465 GNDA.n1932 GNDA.n1931 4.79217
R5466 GNDA.n1930 GNDA.n1929 4.79217
R5467 GNDA.n275 GNDA.n274 4.5005
R5468 GNDA.n276 GNDA.n268 4.5005
R5469 GNDA.n278 GNDA.n277 4.5005
R5470 GNDA.n279 GNDA.n153 4.5005
R5471 GNDA.n1876 GNDA.n1875 4.5005
R5472 GNDA.n1874 GNDA.n201 4.5005
R5473 GNDA.n1873 GNDA.n1872 4.5005
R5474 GNDA.n1871 GNDA.n205 4.5005
R5475 GNDA.n1942 GNDA.n1941 4.5005
R5476 GNDA.n1966 GNDA.n1965 4.5005
R5477 GNDA.n1909 GNDA.n1908 4.5005
R5478 GNDA.n1913 GNDA.n1912 4.5005
R5479 GNDA.n288 GNDA.n284 4.5005
R5480 GNDA.n292 GNDA.n291 4.5005
R5481 GNDA.n293 GNDA.n283 4.5005
R5482 GNDA.n1829 GNDA.n1828 4.5005
R5483 GNDA.n2071 GNDA.n2033 4.26717
R5484 GNDA.n2040 GNDA.n2033 4.26717
R5485 GNDA.n2064 GNDA.n2040 4.26717
R5486 GNDA.n2064 GNDA.n2063 4.26717
R5487 GNDA.n2063 GNDA.n2062 4.26717
R5488 GNDA.n2062 GNDA.n2043 4.26717
R5489 GNDA.n2050 GNDA.n2043 4.26717
R5490 GNDA.n2054 GNDA.n2050 4.26717
R5491 GNDA.n2054 GNDA.n2053 4.26717
R5492 GNDA.n2053 GNDA.n2052 4.26717
R5493 GNDA.n2052 GNDA.n113 4.26717
R5494 GNDA.n965 GNDA.n611 4.26717
R5495 GNDA.n960 GNDA.n611 4.26717
R5496 GNDA.n960 GNDA.n959 4.26717
R5497 GNDA.n959 GNDA.n958 4.26717
R5498 GNDA.n958 GNDA.n955 4.26717
R5499 GNDA.n955 GNDA.n954 4.26717
R5500 GNDA.n954 GNDA.n951 4.26717
R5501 GNDA.n951 GNDA.n950 4.26717
R5502 GNDA.n950 GNDA.n947 4.26717
R5503 GNDA.n947 GNDA.n946 4.26717
R5504 GNDA.n946 GNDA.n944 4.26717
R5505 GNDA.n1679 GNDA.n377 4.26717
R5506 GNDA.n1603 GNDA.n377 4.26717
R5507 GNDA.n1604 GNDA.n1603 4.26717
R5508 GNDA.n1609 GNDA.n1604 4.26717
R5509 GNDA.n1610 GNDA.n1609 4.26717
R5510 GNDA.n1615 GNDA.n1610 4.26717
R5511 GNDA.n1617 GNDA.n1615 4.26717
R5512 GNDA.n1620 GNDA.n1617 4.26717
R5513 GNDA.n1624 GNDA.n1620 4.26717
R5514 GNDA.n1624 GNDA.n1621 4.26717
R5515 GNDA.n1621 GNDA.n441 4.26717
R5516 GNDA.n1705 GNDA.n1704 4.26717
R5517 GNDA.n1708 GNDA.n1705 4.26717
R5518 GNDA.n1708 GNDA.n359 4.26717
R5519 GNDA.n1714 GNDA.n359 4.26717
R5520 GNDA.n1715 GNDA.n1714 4.26717
R5521 GNDA.n1718 GNDA.n1715 4.26717
R5522 GNDA.n1718 GNDA.n357 4.26717
R5523 GNDA.n357 GNDA.n351 4.26717
R5524 GNDA.n1725 GNDA.n351 4.26717
R5525 GNDA.n1725 GNDA.n352 4.26717
R5526 GNDA.n352 GNDA.n344 4.26717
R5527 GNDA.n991 GNDA.n990 4.26717
R5528 GNDA.n994 GNDA.n991 4.26717
R5529 GNDA.n994 GNDA.n542 4.26717
R5530 GNDA.n1000 GNDA.n542 4.26717
R5531 GNDA.n1001 GNDA.n1000 4.26717
R5532 GNDA.n1004 GNDA.n1001 4.26717
R5533 GNDA.n1004 GNDA.n540 4.26717
R5534 GNDA.n540 GNDA.n535 4.26717
R5535 GNDA.n1011 GNDA.n535 4.26717
R5536 GNDA.n1011 GNDA.n536 4.26717
R5537 GNDA.n536 GNDA.n527 4.26717
R5538 GNDA.n1216 GNDA.n1166 4.26717
R5539 GNDA.n1210 GNDA.n1166 4.26717
R5540 GNDA.n1210 GNDA.n1209 4.26717
R5541 GNDA.n1209 GNDA.n1208 4.26717
R5542 GNDA.n1208 GNDA.n1185 4.26717
R5543 GNDA.n1188 GNDA.n1185 4.26717
R5544 GNDA.n1199 GNDA.n1188 4.26717
R5545 GNDA.n1199 GNDA.n1198 4.26717
R5546 GNDA.n1198 GNDA.n1197 4.26717
R5547 GNDA.n1197 GNDA.n1193 4.26717
R5548 GNDA.n1193 GNDA.n86 4.26717
R5549 GNDA.n1907 GNDA.n186 4.2505
R5550 GNDA.n1567 GNDA.n154 4.063
R5551 GNDA.n1931 GNDA.n168 4.0005
R5552 GNDA.n2072 GNDA.n2071 3.93531
R5553 GNDA.n965 GNDA.n608 3.93531
R5554 GNDA.n1679 GNDA.n374 3.93531
R5555 GNDA.n1704 GNDA.n363 3.93531
R5556 GNDA.n990 GNDA.n546 3.93531
R5557 GNDA.n1217 GNDA.n1216 3.93531
R5558 GNDA.n1976 GNDA.n1975 3.90675
R5559 GNDA.n1938 GNDA.t544 3.88193
R5560 GNDA.n1937 GNDA.t40 3.88193
R5561 GNDA.n1936 GNDA.t36 3.88193
R5562 GNDA.n1935 GNDA.t167 3.88193
R5563 GNDA.n1971 GNDA.t102 3.88193
R5564 GNDA.n1970 GNDA.t106 3.88193
R5565 GNDA.n1969 GNDA.t568 3.88193
R5566 GNDA.n2390 GNDA.n2389 3.7893
R5567 GNDA.n2386 GNDA.n59 3.7893
R5568 GNDA.n2385 GNDA.n62 3.7893
R5569 GNDA.n2382 GNDA.n2381 3.7893
R5570 GNDA.n2308 GNDA.n63 3.7893
R5571 GNDA.n2317 GNDA.n2316 3.7893
R5572 GNDA.n2320 GNDA.n2307 3.7893
R5573 GNDA.n2325 GNDA.n2321 3.7893
R5574 GNDA.n1084 GNDA.n459 3.7893
R5575 GNDA.n480 GNDA.n479 3.7893
R5576 GNDA.n1078 GNDA.n1077 3.7893
R5577 GNDA.n504 GNDA.n481 3.7893
R5578 GNDA.n506 GNDA.n505 3.7893
R5579 GNDA.n512 GNDA.n501 3.7893
R5580 GNDA.n519 GNDA.n500 3.7893
R5581 GNDA.n520 GNDA.n499 3.7893
R5582 GNDA.n1817 GNDA.n1816 3.7893
R5583 GNDA.n1813 GNDA.n300 3.7893
R5584 GNDA.n1812 GNDA.n303 3.7893
R5585 GNDA.n310 GNDA.n309 3.7893
R5586 GNDA.n1806 GNDA.n1805 3.7893
R5587 GNDA.n1553 GNDA.n1552 3.7893
R5588 GNDA.n1549 GNDA.n1548 3.7893
R5589 GNDA.n1747 GNDA.n329 3.7893
R5590 GNDA.n1586 GNDA.n1319 3.7893
R5591 GNDA.n1585 GNDA.n1320 3.7893
R5592 GNDA.n1573 GNDA.n1572 3.7893
R5593 GNDA.n1579 GNDA.n1578 3.7893
R5594 GNDA.n1575 GNDA.n1574 3.7893
R5595 GNDA.n1324 GNDA.n1298 3.7893
R5596 GNDA.n1331 GNDA.n1329 3.7893
R5597 GNDA.n1333 GNDA.n1332 3.7893
R5598 GNDA.n743 GNDA.n718 3.7893
R5599 GNDA.n742 GNDA.n739 3.7893
R5600 GNDA.n738 GNDA.n719 3.7893
R5601 GNDA.n735 GNDA.n734 3.7893
R5602 GNDA.n731 GNDA.n720 3.7893
R5603 GNDA.n724 GNDA.n721 3.7893
R5604 GNDA.n748 GNDA.n639 3.7893
R5605 GNDA.n749 GNDA.n638 3.7893
R5606 GNDA.n2295 GNDA.n90 3.7893
R5607 GNDA.n2292 GNDA.n2291 3.7893
R5608 GNDA.n2208 GNDA.n91 3.7893
R5609 GNDA.n2213 GNDA.n2211 3.7893
R5610 GNDA.n2218 GNDA.n2214 3.7893
R5611 GNDA.n2225 GNDA.n2224 3.7893
R5612 GNDA.n2228 GNDA.n2207 3.7893
R5613 GNDA.n2233 GNDA.n2229 3.7893
R5614 GNDA.n935 GNDA.n756 3.7893
R5615 GNDA.n932 GNDA.n931 3.7893
R5616 GNDA.n848 GNDA.n757 3.7893
R5617 GNDA.n853 GNDA.n851 3.7893
R5618 GNDA.n858 GNDA.n854 3.7893
R5619 GNDA.n865 GNDA.n864 3.7893
R5620 GNDA.n868 GNDA.n847 3.7893
R5621 GNDA.n873 GNDA.n869 3.7893
R5622 GNDA.n1667 GNDA.n427 3.7893
R5623 GNDA.n1666 GNDA.n428 3.7893
R5624 GNDA.n1654 GNDA.n1653 3.7893
R5625 GNDA.n1660 GNDA.n1659 3.7893
R5626 GNDA.n1656 GNDA.n1655 3.7893
R5627 GNDA.n1461 GNDA.n406 3.7893
R5628 GNDA.n1464 GNDA.n1463 3.7893
R5629 GNDA.n1472 GNDA.n1391 3.7893
R5630 GNDA.n2399 GNDA.n22 3.7893
R5631 GNDA.n2398 GNDA.n23 3.7893
R5632 GNDA.n33 GNDA.n32 3.7893
R5633 GNDA.n39 GNDA.n38 3.7893
R5634 GNDA.n35 GNDA.n34 3.7893
R5635 GNDA.n2131 GNDA.n1 3.7893
R5636 GNDA.n2136 GNDA.n2134 3.7893
R5637 GNDA.n2141 GNDA.n2137 3.7893
R5638 GNDA.n2313 GNDA 3.7381
R5639 GNDA.n513 GNDA 3.7381
R5640 GNDA.n1547 GNDA 3.7381
R5641 GNDA GNDA.n1591 3.7381
R5642 GNDA GNDA.n727 3.7381
R5643 GNDA.n2221 GNDA 3.7381
R5644 GNDA.n861 GNDA 3.7381
R5645 GNDA GNDA.n1672 3.7381
R5646 GNDA GNDA.n2404 3.7381
R5647 GNDA.t179 GNDA.t506 3.66107
R5648 GNDA.t491 GNDA.t147 3.66107
R5649 GNDA.n1275 GNDA.t61 3.66107
R5650 GNDA.n1927 GNDA.t562 3.66107
R5651 GNDA.n1972 GNDA.t25 3.66107
R5652 GNDA.t556 GNDA.t183 3.66107
R5653 GNDA.t190 GNDA.t550 3.66107
R5654 GNDA.n181 GNDA.n167 3.65764
R5655 GNDA.n182 GNDA.n167 3.65764
R5656 GNDA.n175 GNDA.n171 3.65764
R5657 GNDA.n176 GNDA.n171 3.65764
R5658 GNDA.n1909 GNDA.n165 3.53175
R5659 GNDA.n1870 GNDA.n206 3.50448
R5660 GNDA.n269 GNDA.n264 3.47871
R5661 GNDA.n285 GNDA.n261 3.47871
R5662 GNDA.n1875 GNDA.n202 3.43627
R5663 GNDA.n1993 GNDA.t182 3.42907
R5664 GNDA.n1993 GNDA.t47 3.42907
R5665 GNDA.n1991 GNDA.t581 3.42907
R5666 GNDA.n1991 GNDA.t595 3.42907
R5667 GNDA.n1886 GNDA.t164 3.42907
R5668 GNDA.n1886 GNDA.t170 3.42907
R5669 GNDA.n1888 GNDA.t80 3.42907
R5670 GNDA.n1888 GNDA.t603 3.42907
R5671 GNDA.n278 GNDA.n267 3.4105
R5672 GNDA.n272 GNDA.n268 3.4105
R5673 GNDA.n274 GNDA.n273 3.4105
R5674 GNDA.n271 GNDA.n270 3.4105
R5675 GNDA.n280 GNDA.n279 3.4105
R5676 GNDA.n1869 GNDA.n1868 3.4105
R5677 GNDA.n1867 GNDA.n205 3.4105
R5678 GNDA.n1873 GNDA.n204 3.4105
R5679 GNDA.n1874 GNDA.n203 3.4105
R5680 GNDA.n283 GNDA.n282 3.4105
R5681 GNDA.n291 GNDA.n290 3.4105
R5682 GNDA.n289 GNDA.n288 3.4105
R5683 GNDA.n287 GNDA.n286 3.4105
R5684 GNDA.n1830 GNDA.n1829 3.4105
R5685 GNDA.n1831 GNDA.n261 3.4105
R5686 GNDA.n1831 GNDA.n1830 3.4105
R5687 GNDA.n281 GNDA.n264 3.4105
R5688 GNDA.n281 GNDA.n280 3.4105
R5689 GNDA.n1832 GNDA.n256 3.4105
R5690 GNDA.n256 GNDA.n253 3.4105
R5691 GNDA.n1837 GNDA.n256 3.4105
R5692 GNDA.n1836 GNDA.n1835 3.4105
R5693 GNDA.n1837 GNDA.n1836 3.4105
R5694 GNDA.n1835 GNDA.n254 3.4105
R5695 GNDA.n254 GNDA.n250 3.4105
R5696 GNDA.n254 GNDA.n252 3.4105
R5697 GNDA.n254 GNDA.n249 3.4105
R5698 GNDA.n254 GNDA.n253 3.4105
R5699 GNDA.n1837 GNDA.n254 3.4105
R5700 GNDA.n1838 GNDA.n250 3.4105
R5701 GNDA.n1838 GNDA.n252 3.4105
R5702 GNDA.n1838 GNDA.n249 3.4105
R5703 GNDA.n1838 GNDA.n253 3.4105
R5704 GNDA.n1838 GNDA.n1837 3.4105
R5705 GNDA.n1864 GNDA.n1847 3.4105
R5706 GNDA.n1860 GNDA.n1847 3.4105
R5707 GNDA.n1862 GNDA.n1847 3.4105
R5708 GNDA.n1861 GNDA.n1860 3.4105
R5709 GNDA.n1862 GNDA.n1861 3.4105
R5710 GNDA.n1864 GNDA.n208 3.4105
R5711 GNDA.n1852 GNDA.n208 3.4105
R5712 GNDA.n1850 GNDA.n208 3.4105
R5713 GNDA.n1853 GNDA.n208 3.4105
R5714 GNDA.n1860 GNDA.n208 3.4105
R5715 GNDA.n1862 GNDA.n208 3.4105
R5716 GNDA.n1864 GNDA.n1863 3.4105
R5717 GNDA.n1863 GNDA.n1852 3.4105
R5718 GNDA.n1863 GNDA.n1850 3.4105
R5719 GNDA.n1863 GNDA.n1853 3.4105
R5720 GNDA.n1863 GNDA.n1862 3.4105
R5721 GNDA.n1841 GNDA.n222 3.4105
R5722 GNDA.n1844 GNDA.n222 3.4105
R5723 GNDA.n1844 GNDA.n210 3.4105
R5724 GNDA.n1844 GNDA.n1843 3.4105
R5725 GNDA.n1845 GNDA.n1844 3.4105
R5726 GNDA.n222 GNDA.n214 3.4105
R5727 GNDA.n214 GNDA.n212 3.4105
R5728 GNDA.n1843 GNDA.n214 3.4105
R5729 GNDA.n1845 GNDA.n214 3.4105
R5730 GNDA.n1846 GNDA.n210 3.4105
R5731 GNDA.n1846 GNDA.n212 3.4105
R5732 GNDA.n1846 GNDA.n1845 3.4105
R5733 GNDA.n1933 GNDA.n1932 3.39217
R5734 GNDA.n1929 GNDA.n1928 3.39217
R5735 GNDA.n1274 GNDA.n1273 3.39217
R5736 GNDA.n1974 GNDA.n1973 3.39217
R5737 GNDA.n183 GNDA.n181 3.13621
R5738 GNDA.n183 GNDA.n182 3.13621
R5739 GNDA.n177 GNDA.n175 3.13621
R5740 GNDA.n177 GNDA.n176 3.13621
R5741 GNDA.n1822 GNDA.n1821 3.08966
R5742 GNDA.n307 GNDA.t598 3.08966
R5743 GNDA.t575 GNDA.n1556 3.08966
R5744 GNDA.n1744 GNDA.t71 3.08966
R5745 GNDA.n1664 GNDA.t165 3.08966
R5746 GNDA.n391 GNDA.n390 2.86505
R5747 GNDA.n392 GNDA.n391 2.86505
R5748 GNDA.n396 GNDA.n394 2.86505
R5749 GNDA.n399 GNDA.n394 2.86505
R5750 GNDA.n395 GNDA.n392 2.86505
R5751 GNDA.n399 GNDA.n398 2.86505
R5752 GNDA.n401 GNDA.n390 2.86505
R5753 GNDA.n396 GNDA.n395 2.86505
R5754 GNDA.n1561 GNDA.n1560 2.86505
R5755 GNDA.n1560 GNDA.n1559 2.86505
R5756 GNDA.n1559 GNDA.n1558 2.86505
R5757 GNDA.n1562 GNDA.n1561 2.86505
R5758 GNDA.n1910 GNDA.n1909 2.813
R5759 GNDA.n2392 GNDA.n2391 2.6629
R5760 GNDA.n2305 GNDA.n82 2.6629
R5761 GNDA.n1086 GNDA.n1085 2.6629
R5762 GNDA.n1019 GNDA.n524 2.6629
R5763 GNDA.n1819 GNDA.n1818 2.6629
R5764 GNDA.n343 GNDA.n342 2.6629
R5765 GNDA.n1335 GNDA.n1334 2.6629
R5766 GNDA.n1530 GNDA.n1529 2.6629
R5767 GNDA.n717 GNDA.n716 2.6629
R5768 GNDA.n943 GNDA.n754 2.6629
R5769 GNDA.n2297 GNDA.n2296 2.6629
R5770 GNDA.n2205 GNDA.n110 2.6629
R5771 GNDA.n937 GNDA.n936 2.6629
R5772 GNDA.n1528 GNDA.n1527 2.6629
R5773 GNDA.n2197 GNDA.n2196 2.6629
R5774 GNDA.n2306 GNDA.n2305 2.4581
R5775 GNDA.n1020 GNDA.n1019 2.4581
R5776 GNDA.n342 GNDA.n328 2.4581
R5777 GNDA.n1334 GNDA.n343 2.4581
R5778 GNDA.n1531 GNDA.n1530 2.4581
R5779 GNDA.n716 GNDA.n524 2.4581
R5780 GNDA.n754 GNDA.n753 2.4581
R5781 GNDA.n2297 GNDA.n82 2.4581
R5782 GNDA.n2206 GNDA.n2205 2.4581
R5783 GNDA.n943 GNDA.n937 2.4581
R5784 GNDA.n846 GNDA.n845 2.4581
R5785 GNDA.n1529 GNDA.n1528 2.4581
R5786 GNDA.n1458 GNDA.n1390 2.4581
R5787 GNDA.n2197 GNDA.n110 2.4581
R5788 GNDA.n2130 GNDA.n2129 2.4581
R5789 GNDA.n275 GNDA.n269 2.39683
R5790 GNDA.n1871 GNDA.n1870 2.39683
R5791 GNDA.n285 GNDA.n284 2.39683
R5792 GNDA.n1931 GNDA.n1930 2.2505
R5793 GNDA.n1941 GNDA.n1940 2.19633
R5794 GNDA.n113 GNDA.n110 2.18124
R5795 GNDA.n944 GNDA.n943 2.18124
R5796 GNDA.n1529 GNDA.n441 2.18124
R5797 GNDA.n344 GNDA.n343 2.18124
R5798 GNDA.n527 GNDA.n524 2.18124
R5799 GNDA.n86 GNDA.n82 2.18124
R5800 GNDA.n2324 GNDA.n2306 2.1509
R5801 GNDA.n1020 GNDA.n523 2.1509
R5802 GNDA.n1746 GNDA.n328 2.1509
R5803 GNDA.n1532 GNDA.n1531 2.1509
R5804 GNDA.n753 GNDA.n752 2.1509
R5805 GNDA.n2232 GNDA.n2206 2.1509
R5806 GNDA.n872 GNDA.n846 2.1509
R5807 GNDA.n1471 GNDA.n1390 2.1509
R5808 GNDA.n2140 GNDA.n2130 2.1509
R5809 GNDA.n2391 GNDA.n57 2.13383
R5810 GNDA.n1085 GNDA.n458 2.13383
R5811 GNDA.n1818 GNDA.n299 2.13383
R5812 GNDA.n1336 GNDA.n1335 2.13383
R5813 GNDA.n717 GNDA.n711 2.13383
R5814 GNDA.n2296 GNDA.n89 2.13383
R5815 GNDA.n936 GNDA.n755 2.13383
R5816 GNDA.n1527 GNDA.n1526 2.13383
R5817 GNDA.n2196 GNDA.n2195 2.13383
R5818 GNDA.n1997 GNDA.n1996 2.09414
R5819 GNDA.n1989 GNDA.n1988 2.09414
R5820 GNDA.n1884 GNDA.n1883 2.09414
R5821 GNDA.n1892 GNDA.n1891 2.09414
R5822 GNDA.n111 GNDA.n110 2.08643
R5823 GNDA.n943 GNDA.n942 2.08643
R5824 GNDA.n1529 GNDA.n438 2.08643
R5825 GNDA.n1732 GNDA.n343 2.08643
R5826 GNDA.n526 GNDA.n524 2.08643
R5827 GNDA.n84 GNDA.n82 2.08643
R5828 GNDA.n1744 GNDA.t499 2.05994
R5829 GNDA.t547 GNDA.n339 2.05994
R5830 GNDA.n1535 GNDA.t559 2.05994
R5831 GNDA.n1649 GNDA.t488 2.05994
R5832 GNDA.n2391 GNDA.n2390 1.9461
R5833 GNDA.n1085 GNDA.n1084 1.9461
R5834 GNDA.n1818 GNDA.n1817 1.9461
R5835 GNDA.n1335 GNDA.n1319 1.9461
R5836 GNDA.n718 GNDA.n717 1.9461
R5837 GNDA.n2296 GNDA.n2295 1.9461
R5838 GNDA.n936 GNDA.n935 1.9461
R5839 GNDA.n1527 GNDA.n427 1.9461
R5840 GNDA.n2196 GNDA.n22 1.9461
R5841 GNDA.n1975 GNDA.n164 1.938
R5842 GNDA.n2001 GNDA.n2000 1.93383
R5843 GNDA.n2004 GNDA.n2003 1.93383
R5844 GNDA.n1880 GNDA.n1879 1.93383
R5845 GNDA.n1895 GNDA.n1894 1.93383
R5846 GNDA.n1967 GNDA.n1966 1.91062
R5847 GNDA.n2015 GNDA.n2014 1.90675
R5848 GNDA.t422 GNDA.n1265 1.76473
R5849 GNDA.n186 GNDA.n180 1.7505
R5850 GNDA.n258 GNDA.n257 1.70468
R5851 GNDA.n257 GNDA.n248 1.70468
R5852 GNDA.n1855 GNDA.n1854 1.70468
R5853 GNDA.n1854 GNDA.n1848 1.70468
R5854 GNDA.n218 GNDA.n217 1.70468
R5855 GNDA.n223 GNDA.n209 1.70468
R5856 GNDA.n1833 GNDA.n1832 1.70453
R5857 GNDA.n1858 GNDA.n1857 1.70453
R5858 GNDA.n220 GNDA.n219 1.70453
R5859 GNDA.n1834 GNDA.n256 1.70321
R5860 GNDA.n1838 GNDA.n251 1.70321
R5861 GNDA.n1851 GNDA.n1847 1.70321
R5862 GNDA.n1861 GNDA.n207 1.70321
R5863 GNDA.n1841 GNDA.n215 1.70321
R5864 GNDA.n216 GNDA.n214 1.70321
R5865 GNDA.n1846 GNDA.n211 1.70321
R5866 GNDA.n1846 GNDA.n213 1.70321
R5867 GNDA.n256 GNDA.n255 1.70307
R5868 GNDA.n1836 GNDA.n260 1.70307
R5869 GNDA.n1836 GNDA.n259 1.70307
R5870 GNDA.n1856 GNDA.n1847 1.70307
R5871 GNDA.n1861 GNDA.n1859 1.70307
R5872 GNDA.n1863 GNDA.n1849 1.70307
R5873 GNDA.n1841 GNDA.n1840 1.70307
R5874 GNDA.n1842 GNDA.n1841 1.70307
R5875 GNDA.n1844 GNDA.n221 1.70307
R5876 GNDA.n1865 GNDA.n202 1.69337
R5877 GNDA.n1865 GNDA.n206 1.69337
R5878 GNDA.n1831 GNDA.n263 1.6924
R5879 GNDA.n1831 GNDA.n262 1.6924
R5880 GNDA.n281 GNDA.n266 1.6924
R5881 GNDA.n281 GNDA.n265 1.6924
R5882 GNDA.n1866 GNDA.n1865 1.6924
R5883 GNDA.n1885 GNDA.n1878 1.563
R5884 GNDA.n1244 GNDA.n56 1.47392
R5885 GNDA.n1087 GNDA.n457 1.47392
R5886 GNDA.n1127 GNDA.n298 1.47392
R5887 GNDA.n835 GNDA.n776 1.47392
R5888 GNDA.n1457 GNDA.n1394 1.47392
R5889 GNDA.n2119 GNDA.n116 1.47392
R5890 GNDA.n1908 GNDA.n172 1.3755
R5891 GNDA.n1992 GNDA.n1990 1.1255
R5892 GNDA.n1994 GNDA.n1992 1.1255
R5893 GNDA.n1995 GNDA.n1994 1.1255
R5894 GNDA.n1995 GNDA.n1976 1.1255
R5895 GNDA.n1890 GNDA.n1889 1.1255
R5896 GNDA.n1889 GNDA.n1887 1.1255
R5897 GNDA.n1887 GNDA.n1885 1.1255
R5898 GNDA.n1908 GNDA.n1907 1.0005
R5899 GNDA.n1644 GNDA.n1635 0.96925
R5900 GNDA.n1739 GNDA.n1738 0.96925
R5901 GNDA.n2389 GNDA.n59 0.8197
R5902 GNDA.n2386 GNDA.n2385 0.8197
R5903 GNDA.n2382 GNDA.n62 0.8197
R5904 GNDA.n2381 GNDA.n63 0.8197
R5905 GNDA.n2316 GNDA.n2313 0.8197
R5906 GNDA.n2317 GNDA.n2307 0.8197
R5907 GNDA.n2321 GNDA.n2320 0.8197
R5908 GNDA.n2325 GNDA.n2324 0.8197
R5909 GNDA.n479 GNDA.n459 0.8197
R5910 GNDA.n1078 GNDA.n480 0.8197
R5911 GNDA.n1077 GNDA.n481 0.8197
R5912 GNDA.n506 GNDA.n504 0.8197
R5913 GNDA.n513 GNDA.n512 0.8197
R5914 GNDA.n501 GNDA.n500 0.8197
R5915 GNDA.n520 GNDA.n519 0.8197
R5916 GNDA.n523 GNDA.n499 0.8197
R5917 GNDA.n1816 GNDA.n300 0.8197
R5918 GNDA.n1813 GNDA.n1812 0.8197
R5919 GNDA.n309 GNDA.n303 0.8197
R5920 GNDA.n1806 GNDA.n310 0.8197
R5921 GNDA.n1553 GNDA.n1547 0.8197
R5922 GNDA.n1552 GNDA.n1548 0.8197
R5923 GNDA.n1549 GNDA.n329 0.8197
R5924 GNDA.n1747 GNDA.n1746 0.8197
R5925 GNDA.n1586 GNDA.n1585 0.8197
R5926 GNDA.n1572 GNDA.n1320 0.8197
R5927 GNDA.n1579 GNDA.n1573 0.8197
R5928 GNDA.n1578 GNDA.n1575 0.8197
R5929 GNDA.n1591 GNDA.n1298 0.8197
R5930 GNDA.n1329 GNDA.n1324 0.8197
R5931 GNDA.n1332 GNDA.n1331 0.8197
R5932 GNDA.n1532 GNDA.n1333 0.8197
R5933 GNDA.n743 GNDA.n742 0.8197
R5934 GNDA.n739 GNDA.n738 0.8197
R5935 GNDA.n735 GNDA.n719 0.8197
R5936 GNDA.n734 GNDA.n731 0.8197
R5937 GNDA.n727 GNDA.n724 0.8197
R5938 GNDA.n721 GNDA.n639 0.8197
R5939 GNDA.n749 GNDA.n748 0.8197
R5940 GNDA.n752 GNDA.n638 0.8197
R5941 GNDA.n2292 GNDA.n90 0.8197
R5942 GNDA.n2291 GNDA.n91 0.8197
R5943 GNDA.n2211 GNDA.n2208 0.8197
R5944 GNDA.n2214 GNDA.n2213 0.8197
R5945 GNDA.n2224 GNDA.n2221 0.8197
R5946 GNDA.n2225 GNDA.n2207 0.8197
R5947 GNDA.n2229 GNDA.n2228 0.8197
R5948 GNDA.n2233 GNDA.n2232 0.8197
R5949 GNDA.n932 GNDA.n756 0.8197
R5950 GNDA.n931 GNDA.n757 0.8197
R5951 GNDA.n851 GNDA.n848 0.8197
R5952 GNDA.n854 GNDA.n853 0.8197
R5953 GNDA.n864 GNDA.n861 0.8197
R5954 GNDA.n865 GNDA.n847 0.8197
R5955 GNDA.n869 GNDA.n868 0.8197
R5956 GNDA.n873 GNDA.n872 0.8197
R5957 GNDA.n1667 GNDA.n1666 0.8197
R5958 GNDA.n1653 GNDA.n428 0.8197
R5959 GNDA.n1660 GNDA.n1654 0.8197
R5960 GNDA.n1659 GNDA.n1656 0.8197
R5961 GNDA.n1672 GNDA.n406 0.8197
R5962 GNDA.n1464 GNDA.n1461 0.8197
R5963 GNDA.n1463 GNDA.n1391 0.8197
R5964 GNDA.n1472 GNDA.n1471 0.8197
R5965 GNDA.n2399 GNDA.n2398 0.8197
R5966 GNDA.n32 GNDA.n23 0.8197
R5967 GNDA.n39 GNDA.n33 0.8197
R5968 GNDA.n38 GNDA.n35 0.8197
R5969 GNDA.n2404 GNDA.n1 0.8197
R5970 GNDA.n2134 GNDA.n2131 0.8197
R5971 GNDA.n2137 GNDA.n2136 0.8197
R5972 GNDA.n2141 GNDA.n2140 0.8197
R5973 GNDA.n1865 GNDA.n1864 0.7384
R5974 GNDA.n1877 GNDA.n164 0.6255
R5975 GNDA GNDA.n2308 0.5637
R5976 GNDA.n505 GNDA 0.5637
R5977 GNDA.n1805 GNDA 0.5637
R5978 GNDA.n1574 GNDA 0.5637
R5979 GNDA GNDA.n720 0.5637
R5980 GNDA.n2218 GNDA 0.5637
R5981 GNDA.n858 GNDA 0.5637
R5982 GNDA.n1655 GNDA 0.5637
R5983 GNDA.n34 GNDA 0.5637
R5984 GNDA.n1923 GNDA.n1921 0.563
R5985 GNDA.n1921 GNDA.n1919 0.563
R5986 GNDA.n1919 GNDA.n1917 0.563
R5987 GNDA.n1917 GNDA.n1915 0.563
R5988 GNDA.n1915 GNDA.n1913 0.563
R5989 GNDA.n1944 GNDA.n1942 0.563
R5990 GNDA.n1946 GNDA.n1944 0.563
R5991 GNDA.n1948 GNDA.n1946 0.563
R5992 GNDA.n1950 GNDA.n1948 0.563
R5993 GNDA.n1952 GNDA.n1950 0.563
R5994 GNDA.n1954 GNDA.n1952 0.563
R5995 GNDA.n1956 GNDA.n1954 0.563
R5996 GNDA.n1958 GNDA.n1956 0.563
R5997 GNDA.n1960 GNDA.n1958 0.563
R5998 GNDA.n1962 GNDA.n1960 0.563
R5999 GNDA.n1964 GNDA.n1962 0.563
R6000 GNDA.n1981 GNDA.n1979 0.563
R6001 GNDA.n1983 GNDA.n1981 0.563
R6002 GNDA.n1985 GNDA.n1983 0.563
R6003 GNDA.n1987 GNDA.n1985 0.563
R6004 GNDA.n194 GNDA.n192 0.563
R6005 GNDA.n196 GNDA.n194 0.563
R6006 GNDA.n198 GNDA.n196 0.563
R6007 GNDA.n200 GNDA.n198 0.563
R6008 GNDA.n1641 GNDA.n1639 0.563
R6009 GNDA.n1643 GNDA.n1641 0.563
R6010 GNDA.n1644 GNDA.n1643 0.563
R6011 GNDA.n1635 GNDA.n436 0.563
R6012 GNDA.n436 GNDA.n434 0.563
R6013 GNDA.n434 GNDA.n432 0.563
R6014 GNDA.n432 GNDA.n338 0.563
R6015 GNDA.n1738 GNDA.n338 0.563
R6016 GNDA.n1739 GNDA.n336 0.563
R6017 GNDA.n336 GNDA.n334 0.563
R6018 GNDA.n334 GNDA.n295 0.563
R6019 GNDA.n1825 GNDA.n295 0.563
R6020 GNDA.n1265 GNDA.n1264 0.524185
R6021 GNDA.n1831 GNDA.n281 0.513975
R6022 GNDA.n1832 GNDA.n1831 0.476375
R6023 GNDA.n1841 GNDA.n1839 0.466681
R6024 GNDA.n1845 GNDA 0.422325
R6025 GNDA.n1847 GNDA.n1846 0.404112
R6026 GNDA.n2311 GNDA 0.2565
R6027 GNDA.n509 GNDA 0.2565
R6028 GNDA.n1546 GNDA 0.2565
R6029 GNDA.n1592 GNDA 0.2565
R6030 GNDA.n728 GNDA 0.2565
R6031 GNDA GNDA.n2217 0.2565
R6032 GNDA GNDA.n857 0.2565
R6033 GNDA.n1673 GNDA 0.2565
R6034 GNDA GNDA.n0 0.2565
R6035 GNDA.n1965 GNDA.n1964 0.21925
R6036 GNDA.n185 GNDA.n183 0.208833
R6037 GNDA.n179 GNDA.n177 0.208833
R6038 GNDA.t318 GNDA.t393 0.1603
R6039 GNDA.t441 GNDA.t318 0.1603
R6040 GNDA.t290 GNDA.t441 0.1603
R6041 GNDA.t427 GNDA.t290 0.1603
R6042 GNDA.t397 GNDA.t257 0.1603
R6043 GNDA.t322 GNDA.t397 0.1603
R6044 GNDA.t365 GNDA.t322 0.1603
R6045 GNDA.t294 GNDA.t365 0.1603
R6046 GNDA.t224 GNDA.t417 0.1603
R6047 GNDA.t385 GNDA.t224 0.1603
R6048 GNDA.t410 GNDA.t385 0.1603
R6049 GNDA.t459 GNDA.t410 0.1603
R6050 GNDA.t327 GNDA.t205 0.1603
R6051 GNDA.t452 GNDA.t327 0.1603
R6052 GNDA.t299 GNDA.t452 0.1603
R6053 GNDA.t471 GNDA.t299 0.1603
R6054 GNDA.t351 GNDA.t398 0.1603
R6055 GNDA.t317 GNDA.t351 0.1603
R6056 GNDA.t391 GNDA.t317 0.1603
R6057 GNDA.t418 GNDA.t391 0.1603
R6058 GNDA.t211 GNDA.t264 0.1603
R6059 GNDA.t331 GNDA.t211 0.1603
R6060 GNDA.t373 GNDA.t331 0.1603
R6061 GNDA.t303 GNDA.t373 0.1603
R6062 GNDA.t233 GNDA.t260 0.1603
R6063 GNDA.t395 GNDA.t233 0.1603
R6064 GNDA.t254 GNDA.t395 0.1603
R6065 GNDA.t272 GNDA.t254 0.1603
R6066 GNDA.t426 GNDA.t287 0.1603
R6067 GNDA.t213 GNDA.t426 0.1603
R6068 GNDA.t401 GNDA.t213 0.1603
R6069 GNDA.t378 GNDA.t401 0.1603
R6070 GNDA.t434 GNDA.t282 0.1603
R6071 GNDA.t258 GNDA.t434 0.1603
R6072 GNDA.t277 GNDA.t258 0.1603
R6073 GNDA.t346 GNDA.t277 0.1603
R6074 GNDA.t291 GNDA.t361 0.1603
R6075 GNDA.t463 GNDA.t291 0.1603
R6076 GNDA.t454 GNDA.t463 0.1603
R6077 GNDA.t407 GNDA.t454 0.1603
R6078 GNDA.t314 GNDA.t355 0.1603
R6079 GNDA.t281 GNDA.t314 0.1603
R6080 GNDA.t350 GNDA.t281 0.1603
R6081 GNDA.t229 GNDA.t350 0.1603
R6082 GNDA.t469 GNDA.t298 0.1603
R6083 GNDA.t222 GNDA.t469 0.1603
R6084 GNDA.t414 GNDA.t222 0.1603
R6085 GNDA.t388 GNDA.t414 0.1603
R6086 GNDA.t442 GNDA.t292 0.1603
R6087 GNDA.t425 GNDA.t442 0.1603
R6088 GNDA.t286 GNDA.t425 0.1603
R6089 GNDA.t356 GNDA.t286 0.1603
R6090 GNDA.t302 GNDA.t372 0.1603
R6091 GNDA.t472 GNDA.t302 0.1603
R6092 GNDA.t270 GNDA.t472 0.1603
R6093 GNDA.t419 GNDA.t270 0.1603
R6094 GNDA.t323 GNDA.t366 0.1603
R6095 GNDA.t289 GNDA.t323 0.1603
R6096 GNDA.t359 GNDA.t289 0.1603
R6097 GNDA.t238 GNDA.t359 0.1603
R6098 GNDA.t375 GNDA.t252 0.1603
R6099 GNDA.t304 GNDA.t375 0.1603
R6100 GNDA.t344 GNDA.t304 0.1603
R6101 GNDA.t273 GNDA.t344 0.1603
R6102 GNDA.t204 GNDA.t246 0.1603
R6103 GNDA.t364 GNDA.t204 0.1603
R6104 GNDA.t241 GNDA.t364 0.1603
R6105 GNDA.t437 GNDA.t241 0.1603
R6106 GNDA.t309 GNDA.t381 0.1603
R6107 GNDA.t432 GNDA.t309 0.1603
R6108 GNDA.t279 GNDA.t432 0.1603
R6109 GNDA.t261 GNDA.t279 0.1603
R6110 GNDA.t332 GNDA.t376 0.1603
R6111 GNDA.t301 GNDA.t332 0.1603
R6112 GNDA.t371 GNDA.t301 0.1603
R6113 GNDA.t247 GNDA.t371 0.1603
R6114 GNDA.t386 GNDA.t412 0.1603
R6115 GNDA.t311 GNDA.t386 0.1603
R6116 GNDA.t353 GNDA.t311 0.1603
R6117 GNDA.t283 GNDA.t353 0.1603
R6118 GNDA.t214 GNDA.t404 0.1603
R6119 GNDA.t374 GNDA.t214 0.1603
R6120 GNDA.t251 GNDA.t374 0.1603
R6121 GNDA.t447 GNDA.t251 0.1603
R6122 GNDA.t415 GNDA.t267 0.1603
R6123 GNDA.t389 GNDA.t415 0.1603
R6124 GNDA.t235 GNDA.t389 0.1603
R6125 GNDA.t357 GNDA.t235 0.1603
R6126 GNDA.t464 GNDA.t456 0.1603
R6127 GNDA.t403 GNDA.t464 0.1603
R6128 GNDA.t451 GNDA.t403 0.1603
R6129 GNDA.t326 GNDA.t451 0.1603
R6130 GNDA.t396 GNDA.t255 0.1603
R6131 GNDA.t321 GNDA.t396 0.1603
R6132 GNDA.t363 GNDA.t321 0.1603
R6133 GNDA.t293 GNDA.t363 0.1603
R6134 GNDA.t223 GNDA.t416 0.1603
R6135 GNDA.t384 GNDA.t223 0.1603
R6136 GNDA.t409 GNDA.t384 0.1603
R6137 GNDA.t458 GNDA.t409 0.1603
R6138 GNDA.t259 GNDA.t278 0.1603
R6139 GNDA.t203 GNDA.t259 0.1603
R6140 GNDA.t245 GNDA.t203 0.1603
R6141 GNDA.t367 GNDA.t245 0.1603
R6142 GNDA.t473 GNDA.t271 0.1603
R6143 GNDA.t413 GNDA.t473 0.1603
R6144 GNDA.t460 GNDA.t413 0.1603
R6145 GNDA.t337 GNDA.t460 0.1603
R6146 GNDA.t269 GNDA.t339 0.1603
R6147 GNDA.t420 GNDA.t269 0.1603
R6148 GNDA.t433 GNDA.t420 0.1603
R6149 GNDA.t239 GNDA.t433 0.1603
R6150 GNDA.t296 GNDA.t335 0.1603
R6151 GNDA.t453 GNDA.t296 0.1603
R6152 GNDA.t329 GNDA.t453 0.1603
R6153 GNDA.t210 GNDA.t329 0.1603
R6154 GNDA.t343 GNDA.t221 0.1603
R6155 GNDA.t274 GNDA.t343 0.1603
R6156 GNDA.t312 GNDA.t274 0.1603
R6157 GNDA.t438 GNDA.t312 0.1603
R6158 GNDA.t369 GNDA.t217 0.1603
R6159 GNDA.t334 GNDA.t369 0.1603
R6160 GNDA.t212 GNDA.t334 0.1603
R6161 GNDA.t424 GNDA.t212 0.1603
R6162 GNDA.t280 GNDA.t348 0.1603
R6163 GNDA.t262 GNDA.t280 0.1603
R6164 GNDA.t443 GNDA.t262 0.1603
R6165 GNDA.t248 GNDA.t443 0.1603
R6166 GNDA.t305 GNDA.t345 0.1603
R6167 GNDA.t268 GNDA.t305 0.1603
R6168 GNDA.t338 GNDA.t268 0.1603
R6169 GNDA.t218 GNDA.t338 0.1603
R6170 GNDA.t354 GNDA.t232 0.1603
R6171 GNDA.t284 GNDA.t354 0.1603
R6172 GNDA.t324 GNDA.t284 0.1603
R6173 GNDA.t448 GNDA.t324 0.1603
R6174 GNDA.t379 GNDA.t228 0.1603
R6175 GNDA.t342 GNDA.t379 0.1603
R6176 GNDA.t220 GNDA.t342 0.1603
R6177 GNDA.t468 GNDA.t220 0.1603
R6178 GNDA.t236 GNDA.t431 0.1603
R6179 GNDA.t358 GNDA.t236 0.1603
R6180 GNDA.t208 GNDA.t358 0.1603
R6181 GNDA.t328 GNDA.t208 0.1603
R6182 GNDA.t408 GNDA.t428 0.1603
R6183 GNDA.t225 GNDA.t408 0.1603
R6184 GNDA.t470 GNDA.t225 0.1603
R6185 GNDA.t300 GNDA.t470 0.1603
R6186 GNDA.t362 GNDA.t240 0.1603
R6187 GNDA.t295 GNDA.t362 0.1603
R6188 GNDA.t333 GNDA.t295 0.1603
R6189 GNDA.t457 GNDA.t333 0.1603
R6190 GNDA.t390 GNDA.t237 0.1603
R6191 GNDA.t352 GNDA.t390 0.1603
R6192 GNDA.t231 GNDA.t352 0.1603
R6193 GNDA.t429 GNDA.t231 0.1603
R6194 GNDA.t244 GNDA.t440 0.1603
R6195 GNDA.t368 GNDA.t244 0.1603
R6196 GNDA.t215 GNDA.t368 0.1603
R6197 GNDA.t336 GNDA.t215 0.1603
R6198 GNDA.t253 GNDA.t436 0.1603
R6199 GNDA.t234 GNDA.t253 0.1603
R6200 GNDA.t430 GNDA.t234 0.1603
R6201 GNDA.t307 GNDA.t430 0.1603
R6202 GNDA.t445 GNDA.t320 0.1603
R6203 GNDA.t249 GNDA.t445 0.1603
R6204 GNDA.t465 GNDA.t249 0.1603
R6205 GNDA.t219 GNDA.t465 0.1603
R6206 GNDA.t275 GNDA.t315 0.1603
R6207 GNDA.t435 GNDA.t275 0.1603
R6208 GNDA.t310 GNDA.t435 0.1603
R6209 GNDA.t383 GNDA.t310 0.1603
R6210 GNDA.t402 GNDA.t449 0.1603
R6211 GNDA.t377 GNDA.t402 0.1603
R6212 GNDA.t226 GNDA.t377 0.1603
R6213 GNDA.t347 GNDA.t226 0.1603
R6214 GNDA.t263 GNDA.t446 0.1603
R6215 GNDA.t243 GNDA.t263 0.1603
R6216 GNDA.t439 GNDA.t243 0.1603
R6217 GNDA.t316 GNDA.t439 0.1603
R6218 GNDA.t455 GNDA.t330 0.1603
R6219 GNDA.t406 GNDA.t455 0.1603
R6220 GNDA.t474 GNDA.t406 0.1603
R6221 GNDA.t230 GNDA.t474 0.1603
R6222 GNDA.t285 GNDA.t325 0.1603
R6223 GNDA.t444 GNDA.t285 0.1603
R6224 GNDA.t319 GNDA.t444 0.1603
R6225 GNDA.t394 GNDA.t319 0.1603
R6226 GNDA.t380 GNDA.t405 0.1603
R6227 GNDA.t308 GNDA.t380 0.1603
R6228 GNDA.t341 GNDA.t308 0.1603
R6229 GNDA.t387 GNDA.t341 0.1603
R6230 GNDA.t276 GNDA.n224 0.159278
R6231 GNDA.t340 GNDA.n225 0.159278
R6232 GNDA.t266 GNDA.n226 0.159278
R6233 GNDA.t411 GNDA.n227 0.159278
R6234 GNDA.t450 GNDA.n228 0.159278
R6235 GNDA.t250 GNDA.n229 0.159278
R6236 GNDA.t370 GNDA.n230 0.159278
R6237 GNDA.t242 GNDA.n231 0.159278
R6238 GNDA.t360 GNDA.n232 0.159278
R6239 GNDA.t297 GNDA.n233 0.159278
R6240 GNDA.t466 GNDA.n234 0.159278
R6241 GNDA.t288 GNDA.n235 0.159278
R6242 GNDA.t265 GNDA.n236 0.159278
R6243 GNDA.t209 GNDA.n237 0.159278
R6244 GNDA.t256 GNDA.n238 0.159278
R6245 GNDA.t392 GNDA.n239 0.159278
R6246 GNDA.t313 GNDA.n240 0.159278
R6247 GNDA.t382 GNDA.n241 0.159278
R6248 GNDA.t306 GNDA.n242 0.159278
R6249 GNDA.t475 GNDA.n243 0.159278
R6250 GNDA.t227 GNDA.n244 0.159278
R6251 GNDA.t467 GNDA.n245 0.159278
R6252 GNDA.t216 GNDA.n246 0.159278
R6253 GNDA.n274 GNDA.n271 0.146333
R6254 GNDA.n274 GNDA.n268 0.146333
R6255 GNDA.n278 GNDA.n268 0.146333
R6256 GNDA.n276 GNDA.n275 0.146333
R6257 GNDA.n277 GNDA.n276 0.146333
R6258 GNDA.n1874 GNDA.n1873 0.146333
R6259 GNDA.n1873 GNDA.n205 0.146333
R6260 GNDA.n1869 GNDA.n205 0.146333
R6261 GNDA.n1872 GNDA.n201 0.146333
R6262 GNDA.n1872 GNDA.n1871 0.146333
R6263 GNDA.n292 GNDA.n284 0.146333
R6264 GNDA.n293 GNDA.n292 0.146333
R6265 GNDA.n288 GNDA.n287 0.146333
R6266 GNDA.n291 GNDA.n288 0.146333
R6267 GNDA.n291 GNDA.n283 0.146333
R6268 GNDA.n247 GNDA.t427 0.1368
R6269 GNDA.n246 GNDA.t294 0.1368
R6270 GNDA.n246 GNDA.t459 0.1368
R6271 GNDA.n245 GNDA.t471 0.1368
R6272 GNDA.n245 GNDA.t418 0.1368
R6273 GNDA.n244 GNDA.t303 0.1368
R6274 GNDA.n244 GNDA.t272 0.1368
R6275 GNDA.n243 GNDA.t378 0.1368
R6276 GNDA.n243 GNDA.t346 0.1368
R6277 GNDA.n242 GNDA.t407 0.1368
R6278 GNDA.n242 GNDA.t229 0.1368
R6279 GNDA.n241 GNDA.t388 0.1368
R6280 GNDA.n241 GNDA.t356 0.1368
R6281 GNDA.n240 GNDA.t419 0.1368
R6282 GNDA.n240 GNDA.t238 0.1368
R6283 GNDA.n239 GNDA.t273 0.1368
R6284 GNDA.n239 GNDA.t437 0.1368
R6285 GNDA.n238 GNDA.t261 0.1368
R6286 GNDA.n238 GNDA.t247 0.1368
R6287 GNDA.n237 GNDA.t283 0.1368
R6288 GNDA.n237 GNDA.t447 0.1368
R6289 GNDA.n236 GNDA.t357 0.1368
R6290 GNDA.n236 GNDA.t326 0.1368
R6291 GNDA.n235 GNDA.t293 0.1368
R6292 GNDA.n235 GNDA.t458 0.1368
R6293 GNDA.n234 GNDA.t367 0.1368
R6294 GNDA.n234 GNDA.t337 0.1368
R6295 GNDA.n233 GNDA.t239 0.1368
R6296 GNDA.n233 GNDA.t210 0.1368
R6297 GNDA.n232 GNDA.t438 0.1368
R6298 GNDA.n232 GNDA.t424 0.1368
R6299 GNDA.n231 GNDA.t248 0.1368
R6300 GNDA.n231 GNDA.t218 0.1368
R6301 GNDA.n230 GNDA.t448 0.1368
R6302 GNDA.n230 GNDA.t468 0.1368
R6303 GNDA.n229 GNDA.t328 0.1368
R6304 GNDA.n229 GNDA.t300 0.1368
R6305 GNDA.n228 GNDA.t457 0.1368
R6306 GNDA.n228 GNDA.t429 0.1368
R6307 GNDA.n227 GNDA.t336 0.1368
R6308 GNDA.n227 GNDA.t307 0.1368
R6309 GNDA.n226 GNDA.t219 0.1368
R6310 GNDA.n226 GNDA.t383 0.1368
R6311 GNDA.n225 GNDA.t347 0.1368
R6312 GNDA.n225 GNDA.t316 0.1368
R6313 GNDA.n224 GNDA.t230 0.1368
R6314 GNDA.n224 GNDA.t394 0.1368
R6315 GNDA.t405 GNDA.n247 0.1368
R6316 GNDA.n1839 GNDA.t387 0.1368
R6317 GNDA.n279 GNDA.n278 0.135917
R6318 GNDA.n277 GNDA.n153 0.135917
R6319 GNDA.n1875 GNDA.n1874 0.135917
R6320 GNDA.n1876 GNDA.n201 0.135917
R6321 GNDA.n1828 GNDA.n293 0.135917
R6322 GNDA.n1829 GNDA.n283 0.135917
R6323 GNDA.n271 GNDA.n269 0.0667303
R6324 GNDA.n1870 GNDA.n1869 0.0667303
R6325 GNDA.n287 GNDA.n285 0.0667303
R6326 GNDA.n273 GNDA.n272 0.0553333
R6327 GNDA.n204 GNDA.n203 0.0553333
R6328 GNDA.n1868 GNDA.n1867 0.0553333
R6329 GNDA.n290 GNDA.n289 0.0553333
R6330 GNDA GNDA.n2311 0.0517
R6331 GNDA GNDA.n509 0.0517
R6332 GNDA GNDA.n1546 0.0517
R6333 GNDA.n1592 GNDA 0.0517
R6334 GNDA.n728 GNDA 0.0517
R6335 GNDA.n2217 GNDA 0.0517
R6336 GNDA.n857 GNDA 0.0517
R6337 GNDA.n1673 GNDA 0.0517
R6338 GNDA GNDA.n0 0.0517
R6339 GNDA.n270 GNDA.n264 0.0514167
R6340 GNDA.n280 GNDA.n267 0.0514167
R6341 GNDA.n286 GNDA.n261 0.0514167
R6342 GNDA.n1830 GNDA.n282 0.0514167
R6343 GNDA.n273 GNDA.n265 0.028198
R6344 GNDA.n267 GNDA.n266 0.028198
R6345 GNDA.n289 GNDA.n262 0.028198
R6346 GNDA.n282 GNDA.n263 0.028198
R6347 GNDA.n290 GNDA.n263 0.028198
R6348 GNDA.n286 GNDA.n262 0.028198
R6349 GNDA.n272 GNDA.n266 0.028198
R6350 GNDA.n270 GNDA.n265 0.028198
R6351 GNDA.n1866 GNDA.n204 0.028198
R6352 GNDA.n1867 GNDA.n1866 0.028198
R6353 GNDA.n1868 GNDA.n206 0.0262697
R6354 GNDA.n203 GNDA.n202 0.0262697
R6355 GNDA.n1839 GNDA.n1838 0.015775
R6356 GNDA.n1862 GNDA.n1854 0.0116625
R6357 GNDA.n1860 GNDA.n1854 0.0116625
R6358 GNDA.n1837 GNDA.n257 0.0116625
R6359 GNDA.n257 GNDA.n253 0.0116625
R6360 GNDA.n1857 GNDA.n1849 0.0068649
R6361 GNDA.n1857 GNDA.n1856 0.0068649
R6362 GNDA.n1859 GNDA.n1850 0.0068649
R6363 GNDA.n259 GNDA.n249 0.0068649
R6364 GNDA.n255 GNDA.n249 0.0068649
R6365 GNDA.n260 GNDA.n250 0.0068649
R6366 GNDA.n255 GNDA.n252 0.0068649
R6367 GNDA.n260 GNDA.n252 0.0068649
R6368 GNDA.n259 GNDA.n253 0.0068649
R6369 GNDA.n1856 GNDA.n1853 0.0068649
R6370 GNDA.n1859 GNDA.n1853 0.0068649
R6371 GNDA.n1860 GNDA.n1849 0.0068649
R6372 GNDA.n1843 GNDA.n1842 0.0068649
R6373 GNDA.n223 GNDA.n221 0.0068649
R6374 GNDA.n1840 GNDA.n212 0.0068649
R6375 GNDA.n1840 GNDA.n210 0.0068649
R6376 GNDA.n1842 GNDA.n223 0.0068649
R6377 GNDA.n221 GNDA.n212 0.0068649
R6378 GNDA.n1851 GNDA.n1850 0.00657213
R6379 GNDA.n1864 GNDA.n207 0.00657213
R6380 GNDA.n1834 GNDA.n250 0.00657213
R6381 GNDA.n1832 GNDA.n251 0.00657213
R6382 GNDA.n1835 GNDA.n1834 0.00657213
R6383 GNDA.n1835 GNDA.n251 0.00657213
R6384 GNDA.n1852 GNDA.n1851 0.00657213
R6385 GNDA.n1852 GNDA.n207 0.00657213
R6386 GNDA.n1845 GNDA.n215 0.00657213
R6387 GNDA.n1843 GNDA.n213 0.00657213
R6388 GNDA.n216 GNDA.n210 0.00657213
R6389 GNDA.n222 GNDA.n211 0.00657213
R6390 GNDA.n219 GNDA.n215 0.00657213
R6391 GNDA.n217 GNDA.n216 0.00657213
R6392 GNDA.n217 GNDA.n211 0.00657213
R6393 GNDA.n219 GNDA.n213 0.00657213
R6394 GNDA.n1833 GNDA.n254 0.00393497
R6395 GNDA.n220 GNDA.n214 0.00393497
R6396 GNDA.n1858 GNDA.n208 0.00393497
R6397 GNDA.n1836 GNDA.n1833 0.00393497
R6398 GNDA.n1861 GNDA.n1858 0.00393497
R6399 GNDA.n1844 GNDA.n220 0.00393497
R6400 GNDA.n1836 GNDA.n258 0.0036417
R6401 GNDA.n1838 GNDA.n248 0.0036417
R6402 GNDA.n1844 GNDA.n218 0.0036417
R6403 GNDA.n1846 GNDA.n209 0.0036417
R6404 GNDA.n1861 GNDA.n1855 0.0036417
R6405 GNDA.n1863 GNDA.n1848 0.0036417
R6406 GNDA.n258 GNDA.n256 0.0036417
R6407 GNDA.n254 GNDA.n248 0.0036417
R6408 GNDA.n1855 GNDA.n1847 0.0036417
R6409 GNDA.n1848 GNDA.n208 0.0036417
R6410 GNDA.n1841 GNDA.n218 0.0036417
R6411 GNDA.n214 GNDA.n209 0.0036417
R6412 GNDA.n224 GNDA.t349 0.00152174
R6413 GNDA.n225 GNDA.t276 0.00152174
R6414 GNDA.n226 GNDA.t340 0.00152174
R6415 GNDA.n227 GNDA.t266 0.00152174
R6416 GNDA.n228 GNDA.t411 0.00152174
R6417 GNDA.n229 GNDA.t450 0.00152174
R6418 GNDA.n230 GNDA.t250 0.00152174
R6419 GNDA.n231 GNDA.t370 0.00152174
R6420 GNDA.n232 GNDA.t242 0.00152174
R6421 GNDA.n233 GNDA.t360 0.00152174
R6422 GNDA.n234 GNDA.t297 0.00152174
R6423 GNDA.n235 GNDA.t466 0.00152174
R6424 GNDA.n236 GNDA.t288 0.00152174
R6425 GNDA.n237 GNDA.t265 0.00152174
R6426 GNDA.n238 GNDA.t209 0.00152174
R6427 GNDA.n239 GNDA.t256 0.00152174
R6428 GNDA.n240 GNDA.t392 0.00152174
R6429 GNDA.n241 GNDA.t313 0.00152174
R6430 GNDA.n242 GNDA.t382 0.00152174
R6431 GNDA.n243 GNDA.t306 0.00152174
R6432 GNDA.n244 GNDA.t475 0.00152174
R6433 GNDA.n245 GNDA.t227 0.00152174
R6434 GNDA.n246 GNDA.t467 0.00152174
R6435 GNDA.n247 GNDA.t216 0.00152174
R6436 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t31 355.293
R6437 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t32 346.8
R6438 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.n10 339.522
R6439 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.n8 339.522
R6440 bgr_11_0.1st_Vout_2.n12 bgr_11_0.1st_Vout_2.n3 335.022
R6441 bgr_11_0.1st_Vout_2.n6 bgr_11_0.1st_Vout_2.t6 275.909
R6442 bgr_11_0.1st_Vout_2.n6 bgr_11_0.1st_Vout_2.n5 227.909
R6443 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.n7 222.034
R6444 bgr_11_0.1st_Vout_2.n11 bgr_11_0.1st_Vout_2.t16 184.097
R6445 bgr_11_0.1st_Vout_2.n11 bgr_11_0.1st_Vout_2.t25 184.097
R6446 bgr_11_0.1st_Vout_2.n9 bgr_11_0.1st_Vout_2.t12 184.097
R6447 bgr_11_0.1st_Vout_2.n9 bgr_11_0.1st_Vout_2.t24 184.097
R6448 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.n11 166.05
R6449 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.n9 166.05
R6450 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.n4 52.9634
R6451 bgr_11_0.1st_Vout_2.n7 bgr_11_0.1st_Vout_2.t0 48.0005
R6452 bgr_11_0.1st_Vout_2.n7 bgr_11_0.1st_Vout_2.t3 48.0005
R6453 bgr_11_0.1st_Vout_2.n5 bgr_11_0.1st_Vout_2.t4 48.0005
R6454 bgr_11_0.1st_Vout_2.n5 bgr_11_0.1st_Vout_2.t7 48.0005
R6455 bgr_11_0.1st_Vout_2.n10 bgr_11_0.1st_Vout_2.t8 39.4005
R6456 bgr_11_0.1st_Vout_2.n10 bgr_11_0.1st_Vout_2.t5 39.4005
R6457 bgr_11_0.1st_Vout_2.n8 bgr_11_0.1st_Vout_2.t9 39.4005
R6458 bgr_11_0.1st_Vout_2.n8 bgr_11_0.1st_Vout_2.t2 39.4005
R6459 bgr_11_0.1st_Vout_2.t1 bgr_11_0.1st_Vout_2.n12 39.4005
R6460 bgr_11_0.1st_Vout_2.n12 bgr_11_0.1st_Vout_2.t10 39.4005
R6461 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.n1 5.28175
R6462 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.n0 5.188
R6463 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t18 4.8295
R6464 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t23 4.8295
R6465 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t36 4.8295
R6466 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t15 4.8295
R6467 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t17 4.8295
R6468 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t21 4.8295
R6469 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.t34 4.8295
R6470 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.t14 4.8295
R6471 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.t33 4.8295
R6472 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t11 4.5005
R6473 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t30 4.5005
R6474 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t29 4.5005
R6475 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t22 4.5005
R6476 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t35 4.5005
R6477 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t28 4.5005
R6478 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.t27 4.5005
R6479 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.t20 4.5005
R6480 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.t26 4.5005
R6481 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.t19 4.5005
R6482 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.t13 4.5005
R6483 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.n6 4.5005
R6484 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.n2 3.1025
R6485 bgr_11_0.cap_res2.t20 bgr_11_0.cap_res2.t18 121.245
R6486 bgr_11_0.cap_res2.t13 bgr_11_0.cap_res2.t8 0.1603
R6487 bgr_11_0.cap_res2.t7 bgr_11_0.cap_res2.t2 0.1603
R6488 bgr_11_0.cap_res2.t1 bgr_11_0.cap_res2.t15 0.1603
R6489 bgr_11_0.cap_res2.t5 bgr_11_0.cap_res2.t0 0.1603
R6490 bgr_11_0.cap_res2.t19 bgr_11_0.cap_res2.t14 0.1603
R6491 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t4 0.159278
R6492 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t10 0.159278
R6493 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t6 0.159278
R6494 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t12 0.159278
R6495 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t3 0.1368
R6496 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t13 0.1368
R6497 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t17 0.1368
R6498 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t7 0.1368
R6499 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t11 0.1368
R6500 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t1 0.1368
R6501 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t16 0.1368
R6502 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t5 0.1368
R6503 bgr_11_0.cap_res2.n0 bgr_11_0.cap_res2.t9 0.1368
R6504 bgr_11_0.cap_res2.n0 bgr_11_0.cap_res2.t19 0.1368
R6505 bgr_11_0.cap_res2.t4 bgr_11_0.cap_res2.n0 0.00152174
R6506 bgr_11_0.cap_res2.t10 bgr_11_0.cap_res2.n1 0.00152174
R6507 bgr_11_0.cap_res2.t6 bgr_11_0.cap_res2.n2 0.00152174
R6508 bgr_11_0.cap_res2.t12 bgr_11_0.cap_res2.n3 0.00152174
R6509 bgr_11_0.cap_res2.t18 bgr_11_0.cap_res2.n4 0.00152174
R6510 VOUT-.n110 VOUT-.t9 113.16
R6511 VOUT-.n1 VOUT-.n0 34.9935
R6512 VOUT-.n5 VOUT-.n4 34.9935
R6513 VOUT-.n7 VOUT-.n6 34.9935
R6514 VOUT-.n11 VOUT-.n10 34.9935
R6515 VOUT-.n14 VOUT-.n13 34.9935
R6516 VOUT-.n18 VOUT-.n17 34.9935
R6517 VOUT-.n100 VOUT-.n20 20.4693
R6518 VOUT-.n100 VOUT-.n99 11.6871
R6519 VOUT-.n103 VOUT-.n102 9.73997
R6520 VOUT-.n105 VOUT-.n104 9.73997
R6521 VOUT-.n108 VOUT-.n107 9.73997
R6522 VOUT- VOUT-.n100 9.6255
R6523 VOUT-.n108 VOUT-.n106 7.14633
R6524 VOUT-.n106 VOUT-.n103 7.14633
R6525 VOUT-.n103 VOUT-.n101 7.14633
R6526 VOUT-.n0 VOUT-.t7 6.56717
R6527 VOUT-.n0 VOUT-.t1 6.56717
R6528 VOUT-.n4 VOUT-.t14 6.56717
R6529 VOUT-.n4 VOUT-.t4 6.56717
R6530 VOUT-.n6 VOUT-.t13 6.56717
R6531 VOUT-.n6 VOUT-.t3 6.56717
R6532 VOUT-.n10 VOUT-.t6 6.56717
R6533 VOUT-.n10 VOUT-.t12 6.56717
R6534 VOUT-.n13 VOUT-.t8 6.56717
R6535 VOUT-.n13 VOUT-.t2 6.56717
R6536 VOUT-.n17 VOUT-.t5 6.56717
R6537 VOUT-.n17 VOUT-.t15 6.56717
R6538 VOUT-.n18 VOUT-.n16 6.3755
R6539 VOUT-.n19 VOUT-.n18 6.3755
R6540 VOUT-.n8 VOUT-.n5 6.3755
R6541 VOUT-.n5 VOUT-.n3 6.3755
R6542 VOUT-.n105 VOUT-.n101 6.02133
R6543 VOUT-.n106 VOUT-.n105 6.02133
R6544 VOUT-.n109 VOUT-.n108 6.02133
R6545 VOUT-.n7 VOUT-.n3 5.813
R6546 VOUT-.n8 VOUT-.n7 5.813
R6547 VOUT-.n12 VOUT-.n11 5.813
R6548 VOUT-.n11 VOUT-.n9 5.813
R6549 VOUT-.n15 VOUT-.n14 5.813
R6550 VOUT-.n14 VOUT-.n2 5.813
R6551 VOUT-.n16 VOUT-.n1 5.813
R6552 VOUT-.n47 VOUT-.t56 4.8295
R6553 VOUT-.n56 VOUT-.t88 4.8295
R6554 VOUT-.n54 VOUT-.t117 4.8295
R6555 VOUT-.n52 VOUT-.t156 4.8295
R6556 VOUT-.n50 VOUT-.t57 4.8295
R6557 VOUT-.n49 VOUT-.t87 4.8295
R6558 VOUT-.n69 VOUT-.t50 4.8295
R6559 VOUT-.n70 VOUT-.t95 4.8295
R6560 VOUT-.n72 VOUT-.t19 4.8295
R6561 VOUT-.n73 VOUT-.t144 4.8295
R6562 VOUT-.n75 VOUT-.t114 4.8295
R6563 VOUT-.n76 VOUT-.t100 4.8295
R6564 VOUT-.n78 VOUT-.t154 4.8295
R6565 VOUT-.n79 VOUT-.t138 4.8295
R6566 VOUT-.n81 VOUT-.t108 4.8295
R6567 VOUT-.n82 VOUT-.t96 4.8295
R6568 VOUT-.n84 VOUT-.t72 4.8295
R6569 VOUT-.n85 VOUT-.t60 4.8295
R6570 VOUT-.n87 VOUT-.t105 4.8295
R6571 VOUT-.n88 VOUT-.t93 4.8295
R6572 VOUT-.n90 VOUT-.t68 4.8295
R6573 VOUT-.n91 VOUT-.t58 4.8295
R6574 VOUT-.n93 VOUT-.t28 4.8295
R6575 VOUT-.n94 VOUT-.t152 4.8295
R6576 VOUT-.n21 VOUT-.t24 4.8295
R6577 VOUT-.n23 VOUT-.t61 4.8295
R6578 VOUT-.n35 VOUT-.t113 4.8295
R6579 VOUT-.n36 VOUT-.t102 4.8295
R6580 VOUT-.n38 VOUT-.t85 4.8295
R6581 VOUT-.n39 VOUT-.t66 4.8295
R6582 VOUT-.n41 VOUT-.t120 4.8295
R6583 VOUT-.n42 VOUT-.t103 4.8295
R6584 VOUT-.n44 VOUT-.t22 4.8295
R6585 VOUT-.n45 VOUT-.t147 4.8295
R6586 VOUT-.n96 VOUT-.t62 4.8295
R6587 VOUT-.n58 VOUT-.t128 4.8154
R6588 VOUT-.n59 VOUT-.t104 4.8154
R6589 VOUT-.n60 VOUT-.t122 4.8154
R6590 VOUT-.n61 VOUT-.t23 4.8154
R6591 VOUT-.n58 VOUT-.t136 4.806
R6592 VOUT-.n59 VOUT-.t107 4.806
R6593 VOUT-.n60 VOUT-.t130 4.806
R6594 VOUT-.n61 VOUT-.t30 4.806
R6595 VOUT-.n62 VOUT-.t146 4.806
R6596 VOUT-.n63 VOUT-.t49 4.806
R6597 VOUT-.n64 VOUT-.t82 4.806
R6598 VOUT-.n65 VOUT-.t116 4.806
R6599 VOUT-.n66 VOUT-.t99 4.806
R6600 VOUT-.n67 VOUT-.t137 4.806
R6601 VOUT-.n24 VOUT-.t73 4.806
R6602 VOUT-.n25 VOUT-.t121 4.806
R6603 VOUT-.n26 VOUT-.t52 4.806
R6604 VOUT-.n27 VOUT-.t81 4.806
R6605 VOUT-.n28 VOUT-.t134 4.806
R6606 VOUT-.n29 VOUT-.t29 4.806
R6607 VOUT-.n30 VOUT-.t63 4.806
R6608 VOUT-.n31 VOUT-.t98 4.806
R6609 VOUT-.n32 VOUT-.t151 4.806
R6610 VOUT-.n33 VOUT-.t48 4.806
R6611 VOUT-.n47 VOUT-.t153 4.5005
R6612 VOUT-.n48 VOUT-.t39 4.5005
R6613 VOUT-.n56 VOUT-.t123 4.5005
R6614 VOUT-.n57 VOUT-.t143 4.5005
R6615 VOUT-.n54 VOUT-.t20 4.5005
R6616 VOUT-.n55 VOUT-.t44 4.5005
R6617 VOUT-.n52 VOUT-.t59 4.5005
R6618 VOUT-.n53 VOUT-.t75 4.5005
R6619 VOUT-.n50 VOUT-.t92 4.5005
R6620 VOUT-.n51 VOUT-.t109 4.5005
R6621 VOUT-.n49 VOUT-.t54 4.5005
R6622 VOUT-.n68 VOUT-.t69 4.5005
R6623 VOUT-.n67 VOUT-.t34 4.5005
R6624 VOUT-.n66 VOUT-.t135 4.5005
R6625 VOUT-.n65 VOUT-.t155 4.5005
R6626 VOUT-.n64 VOUT-.t111 4.5005
R6627 VOUT-.n63 VOUT-.t78 4.5005
R6628 VOUT-.n62 VOUT-.t45 4.5005
R6629 VOUT-.n61 VOUT-.t64 4.5005
R6630 VOUT-.n60 VOUT-.t25 4.5005
R6631 VOUT-.n59 VOUT-.t149 4.5005
R6632 VOUT-.n58 VOUT-.t33 4.5005
R6633 VOUT-.n69 VOUT-.t148 4.5005
R6634 VOUT-.n71 VOUT-.t32 4.5005
R6635 VOUT-.n70 VOUT-.t131 4.5005
R6636 VOUT-.n72 VOUT-.t119 4.5005
R6637 VOUT-.n74 VOUT-.t70 4.5005
R6638 VOUT-.n73 VOUT-.t40 4.5005
R6639 VOUT-.n75 VOUT-.t84 4.5005
R6640 VOUT-.n77 VOUT-.t37 4.5005
R6641 VOUT-.n76 VOUT-.t140 4.5005
R6642 VOUT-.n78 VOUT-.t112 4.5005
R6643 VOUT-.n80 VOUT-.t65 4.5005
R6644 VOUT-.n79 VOUT-.t35 4.5005
R6645 VOUT-.n81 VOUT-.t76 4.5005
R6646 VOUT-.n83 VOUT-.t26 4.5005
R6647 VOUT-.n82 VOUT-.t132 4.5005
R6648 VOUT-.n84 VOUT-.t43 4.5005
R6649 VOUT-.n86 VOUT-.t125 4.5005
R6650 VOUT-.n85 VOUT-.t94 4.5005
R6651 VOUT-.n87 VOUT-.t71 4.5005
R6652 VOUT-.n89 VOUT-.t21 4.5005
R6653 VOUT-.n88 VOUT-.t124 4.5005
R6654 VOUT-.n90 VOUT-.t38 4.5005
R6655 VOUT-.n92 VOUT-.t118 4.5005
R6656 VOUT-.n91 VOUT-.t89 4.5005
R6657 VOUT-.n93 VOUT-.t133 4.5005
R6658 VOUT-.n95 VOUT-.t80 4.5005
R6659 VOUT-.n94 VOUT-.t53 4.5005
R6660 VOUT-.n21 VOUT-.t129 4.5005
R6661 VOUT-.n22 VOUT-.t77 4.5005
R6662 VOUT-.n23 VOUT-.t106 4.5005
R6663 VOUT-.n34 VOUT-.t67 4.5005
R6664 VOUT-.n33 VOUT-.t115 4.5005
R6665 VOUT-.n32 VOUT-.t31 4.5005
R6666 VOUT-.n31 VOUT-.t126 4.5005
R6667 VOUT-.n30 VOUT-.t42 4.5005
R6668 VOUT-.n29 VOUT-.t91 4.5005
R6669 VOUT-.n28 VOUT-.t142 4.5005
R6670 VOUT-.n27 VOUT-.t97 4.5005
R6671 VOUT-.n26 VOUT-.t150 4.5005
R6672 VOUT-.n25 VOUT-.t86 4.5005
R6673 VOUT-.n24 VOUT-.t47 4.5005
R6674 VOUT-.n35 VOUT-.t83 4.5005
R6675 VOUT-.n37 VOUT-.t36 4.5005
R6676 VOUT-.n36 VOUT-.t139 4.5005
R6677 VOUT-.n38 VOUT-.t55 4.5005
R6678 VOUT-.n40 VOUT-.t141 4.5005
R6679 VOUT-.n39 VOUT-.t101 4.5005
R6680 VOUT-.n41 VOUT-.t90 4.5005
R6681 VOUT-.n43 VOUT-.t41 4.5005
R6682 VOUT-.n42 VOUT-.t145 4.5005
R6683 VOUT-.n44 VOUT-.t127 4.5005
R6684 VOUT-.n46 VOUT-.t74 4.5005
R6685 VOUT-.n45 VOUT-.t46 4.5005
R6686 VOUT-.n96 VOUT-.t27 4.5005
R6687 VOUT-.n97 VOUT-.t110 4.5005
R6688 VOUT-.n98 VOUT-.t79 4.5005
R6689 VOUT-.n99 VOUT-.t51 4.5005
R6690 VOUT-.n20 VOUT-.n19 4.5005
R6691 VOUT-.n102 VOUT-.t11 3.42907
R6692 VOUT-.n102 VOUT-.t16 3.42907
R6693 VOUT-.n104 VOUT-.t18 3.42907
R6694 VOUT-.n104 VOUT-.t10 3.42907
R6695 VOUT-.n107 VOUT-.t17 3.42907
R6696 VOUT-.n107 VOUT-.t0 3.42907
R6697 VOUT- VOUT-.n110 1.78175
R6698 VOUT-.n110 VOUT-.n109 1.69693
R6699 VOUT-.n20 VOUT-.n1 1.313
R6700 VOUT-.n109 VOUT-.n101 1.13443
R6701 VOUT-.n19 VOUT-.n2 0.563
R6702 VOUT-.n9 VOUT-.n2 0.563
R6703 VOUT-.n9 VOUT-.n8 0.563
R6704 VOUT-.n12 VOUT-.n3 0.563
R6705 VOUT-.n15 VOUT-.n12 0.563
R6706 VOUT-.n16 VOUT-.n15 0.563
R6707 VOUT-.n48 VOUT-.n47 0.3295
R6708 VOUT-.n57 VOUT-.n56 0.3295
R6709 VOUT-.n55 VOUT-.n54 0.3295
R6710 VOUT-.n53 VOUT-.n52 0.3295
R6711 VOUT-.n51 VOUT-.n50 0.3295
R6712 VOUT-.n68 VOUT-.n49 0.3295
R6713 VOUT-.n68 VOUT-.n67 0.3295
R6714 VOUT-.n67 VOUT-.n66 0.3295
R6715 VOUT-.n66 VOUT-.n65 0.3295
R6716 VOUT-.n65 VOUT-.n64 0.3295
R6717 VOUT-.n64 VOUT-.n63 0.3295
R6718 VOUT-.n63 VOUT-.n62 0.3295
R6719 VOUT-.n62 VOUT-.n61 0.3295
R6720 VOUT-.n61 VOUT-.n60 0.3295
R6721 VOUT-.n60 VOUT-.n59 0.3295
R6722 VOUT-.n59 VOUT-.n58 0.3295
R6723 VOUT-.n71 VOUT-.n69 0.3295
R6724 VOUT-.n71 VOUT-.n70 0.3295
R6725 VOUT-.n74 VOUT-.n72 0.3295
R6726 VOUT-.n74 VOUT-.n73 0.3295
R6727 VOUT-.n77 VOUT-.n75 0.3295
R6728 VOUT-.n77 VOUT-.n76 0.3295
R6729 VOUT-.n80 VOUT-.n78 0.3295
R6730 VOUT-.n80 VOUT-.n79 0.3295
R6731 VOUT-.n83 VOUT-.n81 0.3295
R6732 VOUT-.n83 VOUT-.n82 0.3295
R6733 VOUT-.n86 VOUT-.n84 0.3295
R6734 VOUT-.n86 VOUT-.n85 0.3295
R6735 VOUT-.n89 VOUT-.n87 0.3295
R6736 VOUT-.n89 VOUT-.n88 0.3295
R6737 VOUT-.n92 VOUT-.n90 0.3295
R6738 VOUT-.n92 VOUT-.n91 0.3295
R6739 VOUT-.n95 VOUT-.n93 0.3295
R6740 VOUT-.n95 VOUT-.n94 0.3295
R6741 VOUT-.n22 VOUT-.n21 0.3295
R6742 VOUT-.n34 VOUT-.n23 0.3295
R6743 VOUT-.n34 VOUT-.n33 0.3295
R6744 VOUT-.n33 VOUT-.n32 0.3295
R6745 VOUT-.n32 VOUT-.n31 0.3295
R6746 VOUT-.n31 VOUT-.n30 0.3295
R6747 VOUT-.n30 VOUT-.n29 0.3295
R6748 VOUT-.n29 VOUT-.n28 0.3295
R6749 VOUT-.n28 VOUT-.n27 0.3295
R6750 VOUT-.n27 VOUT-.n26 0.3295
R6751 VOUT-.n26 VOUT-.n25 0.3295
R6752 VOUT-.n25 VOUT-.n24 0.3295
R6753 VOUT-.n37 VOUT-.n35 0.3295
R6754 VOUT-.n37 VOUT-.n36 0.3295
R6755 VOUT-.n40 VOUT-.n38 0.3295
R6756 VOUT-.n40 VOUT-.n39 0.3295
R6757 VOUT-.n43 VOUT-.n41 0.3295
R6758 VOUT-.n43 VOUT-.n42 0.3295
R6759 VOUT-.n46 VOUT-.n44 0.3295
R6760 VOUT-.n46 VOUT-.n45 0.3295
R6761 VOUT-.n97 VOUT-.n96 0.3295
R6762 VOUT-.n98 VOUT-.n97 0.3295
R6763 VOUT-.n99 VOUT-.n98 0.3295
R6764 VOUT-.n62 VOUT-.n57 0.306
R6765 VOUT-.n63 VOUT-.n55 0.306
R6766 VOUT-.n64 VOUT-.n53 0.306
R6767 VOUT-.n65 VOUT-.n51 0.306
R6768 VOUT-.n68 VOUT-.n48 0.2825
R6769 VOUT-.n71 VOUT-.n68 0.2825
R6770 VOUT-.n74 VOUT-.n71 0.2825
R6771 VOUT-.n77 VOUT-.n74 0.2825
R6772 VOUT-.n80 VOUT-.n77 0.2825
R6773 VOUT-.n83 VOUT-.n80 0.2825
R6774 VOUT-.n86 VOUT-.n83 0.2825
R6775 VOUT-.n89 VOUT-.n86 0.2825
R6776 VOUT-.n92 VOUT-.n89 0.2825
R6777 VOUT-.n95 VOUT-.n92 0.2825
R6778 VOUT-.n34 VOUT-.n22 0.2825
R6779 VOUT-.n37 VOUT-.n34 0.2825
R6780 VOUT-.n40 VOUT-.n37 0.2825
R6781 VOUT-.n43 VOUT-.n40 0.2825
R6782 VOUT-.n46 VOUT-.n43 0.2825
R6783 VOUT-.n97 VOUT-.n46 0.2825
R6784 VOUT-.n97 VOUT-.n95 0.2825
R6785 two_stage_opamp_dummy_magic_23_0.cap_res_X.t0 two_stage_opamp_dummy_magic_23_0.cap_res_X.t1 50.1603
R6786 two_stage_opamp_dummy_magic_23_0.cap_res_X.t124 two_stage_opamp_dummy_magic_23_0.cap_res_X.t29 0.1603
R6787 two_stage_opamp_dummy_magic_23_0.cap_res_X.t8 two_stage_opamp_dummy_magic_23_0.cap_res_X.t53 0.1603
R6788 two_stage_opamp_dummy_magic_23_0.cap_res_X.t132 two_stage_opamp_dummy_magic_23_0.cap_res_X.t35 0.1603
R6789 two_stage_opamp_dummy_magic_23_0.cap_res_X.t93 two_stage_opamp_dummy_magic_23_0.cap_res_X.t134 0.1603
R6790 two_stage_opamp_dummy_magic_23_0.cap_res_X.t34 two_stage_opamp_dummy_magic_23_0.cap_res_X.t69 0.1603
R6791 two_stage_opamp_dummy_magic_23_0.cap_res_X.t14 two_stage_opamp_dummy_magic_23_0.cap_res_X.t34 0.1603
R6792 two_stage_opamp_dummy_magic_23_0.cap_res_X.t112 two_stage_opamp_dummy_magic_23_0.cap_res_X.t14 0.1603
R6793 two_stage_opamp_dummy_magic_23_0.cap_res_X.t137 two_stage_opamp_dummy_magic_23_0.cap_res_X.t40 0.1603
R6794 two_stage_opamp_dummy_magic_23_0.cap_res_X.t113 two_stage_opamp_dummy_magic_23_0.cap_res_X.t137 0.1603
R6795 two_stage_opamp_dummy_magic_23_0.cap_res_X.t79 two_stage_opamp_dummy_magic_23_0.cap_res_X.t113 0.1603
R6796 two_stage_opamp_dummy_magic_23_0.cap_res_X.t103 two_stage_opamp_dummy_magic_23_0.cap_res_X.t70 0.1603
R6797 two_stage_opamp_dummy_magic_23_0.cap_res_X.t4 two_stage_opamp_dummy_magic_23_0.cap_res_X.t101 0.1603
R6798 two_stage_opamp_dummy_magic_23_0.cap_res_X.t26 two_stage_opamp_dummy_magic_23_0.cap_res_X.t62 0.1603
R6799 two_stage_opamp_dummy_magic_23_0.cap_res_X.t9 two_stage_opamp_dummy_magic_23_0.cap_res_X.t107 0.1603
R6800 two_stage_opamp_dummy_magic_23_0.cap_res_X.t117 two_stage_opamp_dummy_magic_23_0.cap_res_X.t13 0.1603
R6801 two_stage_opamp_dummy_magic_23_0.cap_res_X.t38 two_stage_opamp_dummy_magic_23_0.cap_res_X.t138 0.1603
R6802 two_stage_opamp_dummy_magic_23_0.cap_res_X.t17 two_stage_opamp_dummy_magic_23_0.cap_res_X.t57 0.1603
R6803 two_stage_opamp_dummy_magic_23_0.cap_res_X.t73 two_stage_opamp_dummy_magic_23_0.cap_res_X.t43 0.1603
R6804 two_stage_opamp_dummy_magic_23_0.cap_res_X.t122 two_stage_opamp_dummy_magic_23_0.cap_res_X.t19 0.1603
R6805 two_stage_opamp_dummy_magic_23_0.cap_res_X.t45 two_stage_opamp_dummy_magic_23_0.cap_res_X.t3 0.1603
R6806 two_stage_opamp_dummy_magic_23_0.cap_res_X.t25 two_stage_opamp_dummy_magic_23_0.cap_res_X.t61 0.1603
R6807 two_stage_opamp_dummy_magic_23_0.cap_res_X.t81 two_stage_opamp_dummy_magic_23_0.cap_res_X.t49 0.1603
R6808 two_stage_opamp_dummy_magic_23_0.cap_res_X.t63 two_stage_opamp_dummy_magic_23_0.cap_res_X.t97 0.1603
R6809 two_stage_opamp_dummy_magic_23_0.cap_res_X.t114 two_stage_opamp_dummy_magic_23_0.cap_res_X.t85 0.1603
R6810 two_stage_opamp_dummy_magic_23_0.cap_res_X.t33 two_stage_opamp_dummy_magic_23_0.cap_res_X.t64 0.1603
R6811 two_stage_opamp_dummy_magic_23_0.cap_res_X.t86 two_stage_opamp_dummy_magic_23_0.cap_res_X.t52 0.1603
R6812 two_stage_opamp_dummy_magic_23_0.cap_res_X.t68 two_stage_opamp_dummy_magic_23_0.cap_res_X.t99 0.1603
R6813 two_stage_opamp_dummy_magic_23_0.cap_res_X.t119 two_stage_opamp_dummy_magic_23_0.cap_res_X.t89 0.1603
R6814 two_stage_opamp_dummy_magic_23_0.cap_res_X.t104 two_stage_opamp_dummy_magic_23_0.cap_res_X.t5 0.1603
R6815 two_stage_opamp_dummy_magic_23_0.cap_res_X.t24 two_stage_opamp_dummy_magic_23_0.cap_res_X.t129 0.1603
R6816 two_stage_opamp_dummy_magic_23_0.cap_res_X.t78 two_stage_opamp_dummy_magic_23_0.cap_res_X.t106 0.1603
R6817 two_stage_opamp_dummy_magic_23_0.cap_res_X.t130 two_stage_opamp_dummy_magic_23_0.cap_res_X.t95 0.1603
R6818 two_stage_opamp_dummy_magic_23_0.cap_res_X.t111 two_stage_opamp_dummy_magic_23_0.cap_res_X.t10 0.1603
R6819 two_stage_opamp_dummy_magic_23_0.cap_res_X.t30 two_stage_opamp_dummy_magic_23_0.cap_res_X.t135 0.1603
R6820 two_stage_opamp_dummy_magic_23_0.cap_res_X.t12 two_stage_opamp_dummy_magic_23_0.cap_res_X.t54 0.1603
R6821 two_stage_opamp_dummy_magic_23_0.cap_res_X.t67 two_stage_opamp_dummy_magic_23_0.cap_res_X.t37 0.1603
R6822 two_stage_opamp_dummy_magic_23_0.cap_res_X.t56 two_stage_opamp_dummy_magic_23_0.cap_res_X.t91 0.1603
R6823 two_stage_opamp_dummy_magic_23_0.cap_res_X.t102 two_stage_opamp_dummy_magic_23_0.cap_res_X.t72 0.1603
R6824 two_stage_opamp_dummy_magic_23_0.cap_res_X.t18 two_stage_opamp_dummy_magic_23_0.cap_res_X.t55 0.1603
R6825 two_stage_opamp_dummy_magic_23_0.cap_res_X.t74 two_stage_opamp_dummy_magic_23_0.cap_res_X.t44 0.1603
R6826 two_stage_opamp_dummy_magic_23_0.cap_res_X.t110 two_stage_opamp_dummy_magic_23_0.cap_res_X.t84 0.1603
R6827 two_stage_opamp_dummy_magic_23_0.cap_res_X.t71 two_stage_opamp_dummy_magic_23_0.cap_res_X.t36 0.1603
R6828 two_stage_opamp_dummy_magic_23_0.cap_res_X.t7 two_stage_opamp_dummy_magic_23_0.cap_res_X.t105 0.1603
R6829 two_stage_opamp_dummy_magic_23_0.cap_res_X.t60 two_stage_opamp_dummy_magic_23_0.cap_res_X.t76 0.1603
R6830 two_stage_opamp_dummy_magic_23_0.cap_res_X.t15 two_stage_opamp_dummy_magic_23_0.cap_res_X.t23 0.1603
R6831 two_stage_opamp_dummy_magic_23_0.cap_res_X.t66 two_stage_opamp_dummy_magic_23_0.cap_res_X.t128 0.1603
R6832 two_stage_opamp_dummy_magic_23_0.cap_res_X.t115 two_stage_opamp_dummy_magic_23_0.cap_res_X.t94 0.1603
R6833 two_stage_opamp_dummy_magic_23_0.cap_res_X.t31 two_stage_opamp_dummy_magic_23_0.cap_res_X.t59 0.1603
R6834 two_stage_opamp_dummy_magic_23_0.cap_res_X.t126 two_stage_opamp_dummy_magic_23_0.cap_res_X.t6 0.1603
R6835 two_stage_opamp_dummy_magic_23_0.cap_res_X.t42 two_stage_opamp_dummy_magic_23_0.cap_res_X.t109 0.1603
R6836 two_stage_opamp_dummy_magic_23_0.cap_res_X.t51 two_stage_opamp_dummy_magic_23_0.cap_res_X.t96 0.1603
R6837 two_stage_opamp_dummy_magic_23_0.cap_res_X.t28 two_stage_opamp_dummy_magic_23_0.cap_res_X.t133 0.1603
R6838 two_stage_opamp_dummy_magic_23_0.cap_res_X.t65 two_stage_opamp_dummy_magic_23_0.cap_res_X.t100 0.1603
R6839 two_stage_opamp_dummy_magic_23_0.cap_res_X.t48 two_stage_opamp_dummy_magic_23_0.cap_res_X.t65 0.1603
R6840 two_stage_opamp_dummy_magic_23_0.cap_res_X.t2 two_stage_opamp_dummy_magic_23_0.cap_res_X.t48 0.1603
R6841 two_stage_opamp_dummy_magic_23_0.cap_res_X.t82 two_stage_opamp_dummy_magic_23_0.cap_res_X.t46 0.1603
R6842 two_stage_opamp_dummy_magic_23_0.cap_res_X.t98 two_stage_opamp_dummy_magic_23_0.cap_res_X.t82 0.1603
R6843 two_stage_opamp_dummy_magic_23_0.cap_res_X.t1 two_stage_opamp_dummy_magic_23_0.cap_res_X.t98 0.1603
R6844 two_stage_opamp_dummy_magic_23_0.cap_res_X.n29 two_stage_opamp_dummy_magic_23_0.cap_res_X.t21 0.159278
R6845 two_stage_opamp_dummy_magic_23_0.cap_res_X.n30 two_stage_opamp_dummy_magic_23_0.cap_res_X.t50 0.159278
R6846 two_stage_opamp_dummy_magic_23_0.cap_res_X.n31 two_stage_opamp_dummy_magic_23_0.cap_res_X.t27 0.159278
R6847 two_stage_opamp_dummy_magic_23_0.cap_res_X.n32 two_stage_opamp_dummy_magic_23_0.cap_res_X.t127 0.159278
R6848 two_stage_opamp_dummy_magic_23_0.cap_res_X.n33 two_stage_opamp_dummy_magic_23_0.cap_res_X.t11 0.159278
R6849 two_stage_opamp_dummy_magic_23_0.cap_res_X.n34 two_stage_opamp_dummy_magic_23_0.cap_res_X.t108 0.159278
R6850 two_stage_opamp_dummy_magic_23_0.cap_res_X.n25 two_stage_opamp_dummy_magic_23_0.cap_res_X.t118 0.159278
R6851 two_stage_opamp_dummy_magic_23_0.cap_res_X.t90 two_stage_opamp_dummy_magic_23_0.cap_res_X.n9 0.159278
R6852 two_stage_opamp_dummy_magic_23_0.cap_res_X.t121 two_stage_opamp_dummy_magic_23_0.cap_res_X.n10 0.159278
R6853 two_stage_opamp_dummy_magic_23_0.cap_res_X.t16 two_stage_opamp_dummy_magic_23_0.cap_res_X.n11 0.159278
R6854 two_stage_opamp_dummy_magic_23_0.cap_res_X.t116 two_stage_opamp_dummy_magic_23_0.cap_res_X.n12 0.159278
R6855 two_stage_opamp_dummy_magic_23_0.cap_res_X.t83 two_stage_opamp_dummy_magic_23_0.cap_res_X.n13 0.159278
R6856 two_stage_opamp_dummy_magic_23_0.cap_res_X.t47 two_stage_opamp_dummy_magic_23_0.cap_res_X.n14 0.159278
R6857 two_stage_opamp_dummy_magic_23_0.cap_res_X.t77 two_stage_opamp_dummy_magic_23_0.cap_res_X.n15 0.159278
R6858 two_stage_opamp_dummy_magic_23_0.cap_res_X.t39 two_stage_opamp_dummy_magic_23_0.cap_res_X.n16 0.159278
R6859 two_stage_opamp_dummy_magic_23_0.cap_res_X.t136 two_stage_opamp_dummy_magic_23_0.cap_res_X.n17 0.159278
R6860 two_stage_opamp_dummy_magic_23_0.cap_res_X.t32 two_stage_opamp_dummy_magic_23_0.cap_res_X.n18 0.159278
R6861 two_stage_opamp_dummy_magic_23_0.cap_res_X.t131 two_stage_opamp_dummy_magic_23_0.cap_res_X.n19 0.159278
R6862 two_stage_opamp_dummy_magic_23_0.cap_res_X.t92 two_stage_opamp_dummy_magic_23_0.cap_res_X.n20 0.159278
R6863 two_stage_opamp_dummy_magic_23_0.cap_res_X.t120 two_stage_opamp_dummy_magic_23_0.cap_res_X.n21 0.159278
R6864 two_stage_opamp_dummy_magic_23_0.cap_res_X.t87 two_stage_opamp_dummy_magic_23_0.cap_res_X.n22 0.159278
R6865 two_stage_opamp_dummy_magic_23_0.cap_res_X.t125 two_stage_opamp_dummy_magic_23_0.cap_res_X.n23 0.159278
R6866 two_stage_opamp_dummy_magic_23_0.cap_res_X.t88 two_stage_opamp_dummy_magic_23_0.cap_res_X.n24 0.159278
R6867 two_stage_opamp_dummy_magic_23_0.cap_res_X.n26 two_stage_opamp_dummy_magic_23_0.cap_res_X.t20 0.159278
R6868 two_stage_opamp_dummy_magic_23_0.cap_res_X.n27 two_stage_opamp_dummy_magic_23_0.cap_res_X.t58 0.159278
R6869 two_stage_opamp_dummy_magic_23_0.cap_res_X.n28 two_stage_opamp_dummy_magic_23_0.cap_res_X.t41 0.159278
R6870 two_stage_opamp_dummy_magic_23_0.cap_res_X.n35 two_stage_opamp_dummy_magic_23_0.cap_res_X.t75 0.159278
R6871 two_stage_opamp_dummy_magic_23_0.cap_res_X.t118 two_stage_opamp_dummy_magic_23_0.cap_res_X.t4 0.137822
R6872 two_stage_opamp_dummy_magic_23_0.cap_res_X.n25 two_stage_opamp_dummy_magic_23_0.cap_res_X.t103 0.1368
R6873 two_stage_opamp_dummy_magic_23_0.cap_res_X.n24 two_stage_opamp_dummy_magic_23_0.cap_res_X.t26 0.1368
R6874 two_stage_opamp_dummy_magic_23_0.cap_res_X.n24 two_stage_opamp_dummy_magic_23_0.cap_res_X.t9 0.1368
R6875 two_stage_opamp_dummy_magic_23_0.cap_res_X.n23 two_stage_opamp_dummy_magic_23_0.cap_res_X.t117 0.1368
R6876 two_stage_opamp_dummy_magic_23_0.cap_res_X.n23 two_stage_opamp_dummy_magic_23_0.cap_res_X.t38 0.1368
R6877 two_stage_opamp_dummy_magic_23_0.cap_res_X.n22 two_stage_opamp_dummy_magic_23_0.cap_res_X.t17 0.1368
R6878 two_stage_opamp_dummy_magic_23_0.cap_res_X.n22 two_stage_opamp_dummy_magic_23_0.cap_res_X.t73 0.1368
R6879 two_stage_opamp_dummy_magic_23_0.cap_res_X.n21 two_stage_opamp_dummy_magic_23_0.cap_res_X.t122 0.1368
R6880 two_stage_opamp_dummy_magic_23_0.cap_res_X.n21 two_stage_opamp_dummy_magic_23_0.cap_res_X.t45 0.1368
R6881 two_stage_opamp_dummy_magic_23_0.cap_res_X.n20 two_stage_opamp_dummy_magic_23_0.cap_res_X.t25 0.1368
R6882 two_stage_opamp_dummy_magic_23_0.cap_res_X.n20 two_stage_opamp_dummy_magic_23_0.cap_res_X.t81 0.1368
R6883 two_stage_opamp_dummy_magic_23_0.cap_res_X.n19 two_stage_opamp_dummy_magic_23_0.cap_res_X.t63 0.1368
R6884 two_stage_opamp_dummy_magic_23_0.cap_res_X.n19 two_stage_opamp_dummy_magic_23_0.cap_res_X.t114 0.1368
R6885 two_stage_opamp_dummy_magic_23_0.cap_res_X.n18 two_stage_opamp_dummy_magic_23_0.cap_res_X.t33 0.1368
R6886 two_stage_opamp_dummy_magic_23_0.cap_res_X.n18 two_stage_opamp_dummy_magic_23_0.cap_res_X.t86 0.1368
R6887 two_stage_opamp_dummy_magic_23_0.cap_res_X.n17 two_stage_opamp_dummy_magic_23_0.cap_res_X.t68 0.1368
R6888 two_stage_opamp_dummy_magic_23_0.cap_res_X.n17 two_stage_opamp_dummy_magic_23_0.cap_res_X.t119 0.1368
R6889 two_stage_opamp_dummy_magic_23_0.cap_res_X.n16 two_stage_opamp_dummy_magic_23_0.cap_res_X.t104 0.1368
R6890 two_stage_opamp_dummy_magic_23_0.cap_res_X.n16 two_stage_opamp_dummy_magic_23_0.cap_res_X.t24 0.1368
R6891 two_stage_opamp_dummy_magic_23_0.cap_res_X.n15 two_stage_opamp_dummy_magic_23_0.cap_res_X.t78 0.1368
R6892 two_stage_opamp_dummy_magic_23_0.cap_res_X.n15 two_stage_opamp_dummy_magic_23_0.cap_res_X.t130 0.1368
R6893 two_stage_opamp_dummy_magic_23_0.cap_res_X.n14 two_stage_opamp_dummy_magic_23_0.cap_res_X.t111 0.1368
R6894 two_stage_opamp_dummy_magic_23_0.cap_res_X.n14 two_stage_opamp_dummy_magic_23_0.cap_res_X.t30 0.1368
R6895 two_stage_opamp_dummy_magic_23_0.cap_res_X.n13 two_stage_opamp_dummy_magic_23_0.cap_res_X.t12 0.1368
R6896 two_stage_opamp_dummy_magic_23_0.cap_res_X.n13 two_stage_opamp_dummy_magic_23_0.cap_res_X.t67 0.1368
R6897 two_stage_opamp_dummy_magic_23_0.cap_res_X.n12 two_stage_opamp_dummy_magic_23_0.cap_res_X.t56 0.1368
R6898 two_stage_opamp_dummy_magic_23_0.cap_res_X.n12 two_stage_opamp_dummy_magic_23_0.cap_res_X.t102 0.1368
R6899 two_stage_opamp_dummy_magic_23_0.cap_res_X.n11 two_stage_opamp_dummy_magic_23_0.cap_res_X.t18 0.1368
R6900 two_stage_opamp_dummy_magic_23_0.cap_res_X.n11 two_stage_opamp_dummy_magic_23_0.cap_res_X.t74 0.1368
R6901 two_stage_opamp_dummy_magic_23_0.cap_res_X.n10 two_stage_opamp_dummy_magic_23_0.cap_res_X.t51 0.1368
R6902 two_stage_opamp_dummy_magic_23_0.cap_res_X.n9 two_stage_opamp_dummy_magic_23_0.cap_res_X.t28 0.1368
R6903 two_stage_opamp_dummy_magic_23_0.cap_res_X.n0 two_stage_opamp_dummy_magic_23_0.cap_res_X.t110 0.114322
R6904 two_stage_opamp_dummy_magic_23_0.cap_res_X.n30 two_stage_opamp_dummy_magic_23_0.cap_res_X.n29 0.1133
R6905 two_stage_opamp_dummy_magic_23_0.cap_res_X.n31 two_stage_opamp_dummy_magic_23_0.cap_res_X.n30 0.1133
R6906 two_stage_opamp_dummy_magic_23_0.cap_res_X.n32 two_stage_opamp_dummy_magic_23_0.cap_res_X.n31 0.1133
R6907 two_stage_opamp_dummy_magic_23_0.cap_res_X.n33 two_stage_opamp_dummy_magic_23_0.cap_res_X.n32 0.1133
R6908 two_stage_opamp_dummy_magic_23_0.cap_res_X.n34 two_stage_opamp_dummy_magic_23_0.cap_res_X.n33 0.1133
R6909 two_stage_opamp_dummy_magic_23_0.cap_res_X.n1 two_stage_opamp_dummy_magic_23_0.cap_res_X.n0 0.1133
R6910 two_stage_opamp_dummy_magic_23_0.cap_res_X.n2 two_stage_opamp_dummy_magic_23_0.cap_res_X.n1 0.1133
R6911 two_stage_opamp_dummy_magic_23_0.cap_res_X.n3 two_stage_opamp_dummy_magic_23_0.cap_res_X.n2 0.1133
R6912 two_stage_opamp_dummy_magic_23_0.cap_res_X.n4 two_stage_opamp_dummy_magic_23_0.cap_res_X.n3 0.1133
R6913 two_stage_opamp_dummy_magic_23_0.cap_res_X.n5 two_stage_opamp_dummy_magic_23_0.cap_res_X.n4 0.1133
R6914 two_stage_opamp_dummy_magic_23_0.cap_res_X.n6 two_stage_opamp_dummy_magic_23_0.cap_res_X.n5 0.1133
R6915 two_stage_opamp_dummy_magic_23_0.cap_res_X.n7 two_stage_opamp_dummy_magic_23_0.cap_res_X.n6 0.1133
R6916 two_stage_opamp_dummy_magic_23_0.cap_res_X.n8 two_stage_opamp_dummy_magic_23_0.cap_res_X.n7 0.1133
R6917 two_stage_opamp_dummy_magic_23_0.cap_res_X.n10 two_stage_opamp_dummy_magic_23_0.cap_res_X.n8 0.1133
R6918 two_stage_opamp_dummy_magic_23_0.cap_res_X.n26 two_stage_opamp_dummy_magic_23_0.cap_res_X.n25 0.1133
R6919 two_stage_opamp_dummy_magic_23_0.cap_res_X.n27 two_stage_opamp_dummy_magic_23_0.cap_res_X.n26 0.1133
R6920 two_stage_opamp_dummy_magic_23_0.cap_res_X.n28 two_stage_opamp_dummy_magic_23_0.cap_res_X.n27 0.1133
R6921 two_stage_opamp_dummy_magic_23_0.cap_res_X.n35 two_stage_opamp_dummy_magic_23_0.cap_res_X.n28 0.1133
R6922 two_stage_opamp_dummy_magic_23_0.cap_res_X.n35 two_stage_opamp_dummy_magic_23_0.cap_res_X.n34 0.1133
R6923 two_stage_opamp_dummy_magic_23_0.cap_res_X.n29 two_stage_opamp_dummy_magic_23_0.cap_res_X.t124 0.00152174
R6924 two_stage_opamp_dummy_magic_23_0.cap_res_X.n30 two_stage_opamp_dummy_magic_23_0.cap_res_X.t8 0.00152174
R6925 two_stage_opamp_dummy_magic_23_0.cap_res_X.n31 two_stage_opamp_dummy_magic_23_0.cap_res_X.t132 0.00152174
R6926 two_stage_opamp_dummy_magic_23_0.cap_res_X.n32 two_stage_opamp_dummy_magic_23_0.cap_res_X.t93 0.00152174
R6927 two_stage_opamp_dummy_magic_23_0.cap_res_X.n33 two_stage_opamp_dummy_magic_23_0.cap_res_X.t112 0.00152174
R6928 two_stage_opamp_dummy_magic_23_0.cap_res_X.n34 two_stage_opamp_dummy_magic_23_0.cap_res_X.t79 0.00152174
R6929 two_stage_opamp_dummy_magic_23_0.cap_res_X.n0 two_stage_opamp_dummy_magic_23_0.cap_res_X.t71 0.00152174
R6930 two_stage_opamp_dummy_magic_23_0.cap_res_X.n1 two_stage_opamp_dummy_magic_23_0.cap_res_X.t7 0.00152174
R6931 two_stage_opamp_dummy_magic_23_0.cap_res_X.n2 two_stage_opamp_dummy_magic_23_0.cap_res_X.t60 0.00152174
R6932 two_stage_opamp_dummy_magic_23_0.cap_res_X.n3 two_stage_opamp_dummy_magic_23_0.cap_res_X.t15 0.00152174
R6933 two_stage_opamp_dummy_magic_23_0.cap_res_X.n4 two_stage_opamp_dummy_magic_23_0.cap_res_X.t66 0.00152174
R6934 two_stage_opamp_dummy_magic_23_0.cap_res_X.n5 two_stage_opamp_dummy_magic_23_0.cap_res_X.t115 0.00152174
R6935 two_stage_opamp_dummy_magic_23_0.cap_res_X.n6 two_stage_opamp_dummy_magic_23_0.cap_res_X.t31 0.00152174
R6936 two_stage_opamp_dummy_magic_23_0.cap_res_X.n7 two_stage_opamp_dummy_magic_23_0.cap_res_X.t126 0.00152174
R6937 two_stage_opamp_dummy_magic_23_0.cap_res_X.n8 two_stage_opamp_dummy_magic_23_0.cap_res_X.t42 0.00152174
R6938 two_stage_opamp_dummy_magic_23_0.cap_res_X.n9 two_stage_opamp_dummy_magic_23_0.cap_res_X.t80 0.00152174
R6939 two_stage_opamp_dummy_magic_23_0.cap_res_X.n10 two_stage_opamp_dummy_magic_23_0.cap_res_X.t90 0.00152174
R6940 two_stage_opamp_dummy_magic_23_0.cap_res_X.n11 two_stage_opamp_dummy_magic_23_0.cap_res_X.t121 0.00152174
R6941 two_stage_opamp_dummy_magic_23_0.cap_res_X.n12 two_stage_opamp_dummy_magic_23_0.cap_res_X.t16 0.00152174
R6942 two_stage_opamp_dummy_magic_23_0.cap_res_X.n13 two_stage_opamp_dummy_magic_23_0.cap_res_X.t116 0.00152174
R6943 two_stage_opamp_dummy_magic_23_0.cap_res_X.n14 two_stage_opamp_dummy_magic_23_0.cap_res_X.t83 0.00152174
R6944 two_stage_opamp_dummy_magic_23_0.cap_res_X.n15 two_stage_opamp_dummy_magic_23_0.cap_res_X.t47 0.00152174
R6945 two_stage_opamp_dummy_magic_23_0.cap_res_X.n16 two_stage_opamp_dummy_magic_23_0.cap_res_X.t77 0.00152174
R6946 two_stage_opamp_dummy_magic_23_0.cap_res_X.n17 two_stage_opamp_dummy_magic_23_0.cap_res_X.t39 0.00152174
R6947 two_stage_opamp_dummy_magic_23_0.cap_res_X.n18 two_stage_opamp_dummy_magic_23_0.cap_res_X.t136 0.00152174
R6948 two_stage_opamp_dummy_magic_23_0.cap_res_X.n19 two_stage_opamp_dummy_magic_23_0.cap_res_X.t32 0.00152174
R6949 two_stage_opamp_dummy_magic_23_0.cap_res_X.n20 two_stage_opamp_dummy_magic_23_0.cap_res_X.t131 0.00152174
R6950 two_stage_opamp_dummy_magic_23_0.cap_res_X.n21 two_stage_opamp_dummy_magic_23_0.cap_res_X.t92 0.00152174
R6951 two_stage_opamp_dummy_magic_23_0.cap_res_X.n22 two_stage_opamp_dummy_magic_23_0.cap_res_X.t120 0.00152174
R6952 two_stage_opamp_dummy_magic_23_0.cap_res_X.n23 two_stage_opamp_dummy_magic_23_0.cap_res_X.t87 0.00152174
R6953 two_stage_opamp_dummy_magic_23_0.cap_res_X.n24 two_stage_opamp_dummy_magic_23_0.cap_res_X.t125 0.00152174
R6954 two_stage_opamp_dummy_magic_23_0.cap_res_X.n25 two_stage_opamp_dummy_magic_23_0.cap_res_X.t88 0.00152174
R6955 two_stage_opamp_dummy_magic_23_0.cap_res_X.n26 two_stage_opamp_dummy_magic_23_0.cap_res_X.t123 0.00152174
R6956 two_stage_opamp_dummy_magic_23_0.cap_res_X.n27 two_stage_opamp_dummy_magic_23_0.cap_res_X.t22 0.00152174
R6957 two_stage_opamp_dummy_magic_23_0.cap_res_X.n28 two_stage_opamp_dummy_magic_23_0.cap_res_X.t2 0.00152174
R6958 two_stage_opamp_dummy_magic_23_0.cap_res_X.t46 two_stage_opamp_dummy_magic_23_0.cap_res_X.n35 0.00152174
R6959 two_stage_opamp_dummy_magic_23_0.Vb1.n25 two_stage_opamp_dummy_magic_23_0.Vb1.n24 611.782
R6960 two_stage_opamp_dummy_magic_23_0.Vb1.n16 two_stage_opamp_dummy_magic_23_0.Vb1.t18 449.868
R6961 two_stage_opamp_dummy_magic_23_0.Vb1.n9 two_stage_opamp_dummy_magic_23_0.Vb1.t12 449.868
R6962 two_stage_opamp_dummy_magic_23_0.Vb1.n8 two_stage_opamp_dummy_magic_23_0.Vb1.t8 449.868
R6963 two_stage_opamp_dummy_magic_23_0.Vb1.n4 two_stage_opamp_dummy_magic_23_0.Vb1.n2 339.961
R6964 two_stage_opamp_dummy_magic_23_0.Vb1.n4 two_stage_opamp_dummy_magic_23_0.Vb1.n3 339.272
R6965 two_stage_opamp_dummy_magic_23_0.Vb1.n35 two_stage_opamp_dummy_magic_23_0.Vb1.n34 310.392
R6966 two_stage_opamp_dummy_magic_23_0.Vb1.n34 two_stage_opamp_dummy_magic_23_0.Vb1.t33 273.134
R6967 two_stage_opamp_dummy_magic_23_0.Vb1.n25 two_stage_opamp_dummy_magic_23_0.Vb1.t19 273.134
R6968 two_stage_opamp_dummy_magic_23_0.Vb1.n24 two_stage_opamp_dummy_magic_23_0.Vb1.t17 273.134
R6969 two_stage_opamp_dummy_magic_23_0.Vb1.n23 two_stage_opamp_dummy_magic_23_0.Vb1.t27 273.134
R6970 two_stage_opamp_dummy_magic_23_0.Vb1.n22 two_stage_opamp_dummy_magic_23_0.Vb1.t16 273.134
R6971 two_stage_opamp_dummy_magic_23_0.Vb1.n21 two_stage_opamp_dummy_magic_23_0.Vb1.t25 273.134
R6972 two_stage_opamp_dummy_magic_23_0.Vb1.n20 two_stage_opamp_dummy_magic_23_0.Vb1.t34 273.134
R6973 two_stage_opamp_dummy_magic_23_0.Vb1.n19 two_stage_opamp_dummy_magic_23_0.Vb1.t26 273.134
R6974 two_stage_opamp_dummy_magic_23_0.Vb1.n18 two_stage_opamp_dummy_magic_23_0.Vb1.t14 273.134
R6975 two_stage_opamp_dummy_magic_23_0.Vb1.n17 two_stage_opamp_dummy_magic_23_0.Vb1.t24 273.134
R6976 two_stage_opamp_dummy_magic_23_0.Vb1.n16 two_stage_opamp_dummy_magic_23_0.Vb1.t32 273.134
R6977 two_stage_opamp_dummy_magic_23_0.Vb1.n33 two_stage_opamp_dummy_magic_23_0.Vb1.t23 273.134
R6978 two_stage_opamp_dummy_magic_23_0.Vb1.n32 two_stage_opamp_dummy_magic_23_0.Vb1.t31 273.134
R6979 two_stage_opamp_dummy_magic_23_0.Vb1.n31 two_stage_opamp_dummy_magic_23_0.Vb1.t22 273.134
R6980 two_stage_opamp_dummy_magic_23_0.Vb1.n30 two_stage_opamp_dummy_magic_23_0.Vb1.t30 273.134
R6981 two_stage_opamp_dummy_magic_23_0.Vb1.n29 two_stage_opamp_dummy_magic_23_0.Vb1.t20 273.134
R6982 two_stage_opamp_dummy_magic_23_0.Vb1.n28 two_stage_opamp_dummy_magic_23_0.Vb1.t15 273.134
R6983 two_stage_opamp_dummy_magic_23_0.Vb1.n27 two_stage_opamp_dummy_magic_23_0.Vb1.t21 273.134
R6984 two_stage_opamp_dummy_magic_23_0.Vb1.n26 two_stage_opamp_dummy_magic_23_0.Vb1.t29 273.134
R6985 two_stage_opamp_dummy_magic_23_0.Vb1.n9 two_stage_opamp_dummy_magic_23_0.Vb1.t6 273.134
R6986 two_stage_opamp_dummy_magic_23_0.Vb1.n8 two_stage_opamp_dummy_magic_23_0.Vb1.t10 273.134
R6987 two_stage_opamp_dummy_magic_23_0.Vb1.n17 two_stage_opamp_dummy_magic_23_0.Vb1.n16 176.733
R6988 two_stage_opamp_dummy_magic_23_0.Vb1.n18 two_stage_opamp_dummy_magic_23_0.Vb1.n17 176.733
R6989 two_stage_opamp_dummy_magic_23_0.Vb1.n19 two_stage_opamp_dummy_magic_23_0.Vb1.n18 176.733
R6990 two_stage_opamp_dummy_magic_23_0.Vb1.n20 two_stage_opamp_dummy_magic_23_0.Vb1.n19 176.733
R6991 two_stage_opamp_dummy_magic_23_0.Vb1.n21 two_stage_opamp_dummy_magic_23_0.Vb1.n20 176.733
R6992 two_stage_opamp_dummy_magic_23_0.Vb1.n22 two_stage_opamp_dummy_magic_23_0.Vb1.n21 176.733
R6993 two_stage_opamp_dummy_magic_23_0.Vb1.n23 two_stage_opamp_dummy_magic_23_0.Vb1.n22 176.733
R6994 two_stage_opamp_dummy_magic_23_0.Vb1.n24 two_stage_opamp_dummy_magic_23_0.Vb1.n23 176.733
R6995 two_stage_opamp_dummy_magic_23_0.Vb1.n26 two_stage_opamp_dummy_magic_23_0.Vb1.n25 176.733
R6996 two_stage_opamp_dummy_magic_23_0.Vb1.n27 two_stage_opamp_dummy_magic_23_0.Vb1.n26 176.733
R6997 two_stage_opamp_dummy_magic_23_0.Vb1.n28 two_stage_opamp_dummy_magic_23_0.Vb1.n27 176.733
R6998 two_stage_opamp_dummy_magic_23_0.Vb1.n29 two_stage_opamp_dummy_magic_23_0.Vb1.n28 176.733
R6999 two_stage_opamp_dummy_magic_23_0.Vb1.n30 two_stage_opamp_dummy_magic_23_0.Vb1.n29 176.733
R7000 two_stage_opamp_dummy_magic_23_0.Vb1.n31 two_stage_opamp_dummy_magic_23_0.Vb1.n30 176.733
R7001 two_stage_opamp_dummy_magic_23_0.Vb1.n32 two_stage_opamp_dummy_magic_23_0.Vb1.n31 176.733
R7002 two_stage_opamp_dummy_magic_23_0.Vb1.n33 two_stage_opamp_dummy_magic_23_0.Vb1.n32 176.733
R7003 two_stage_opamp_dummy_magic_23_0.Vb1.n34 two_stage_opamp_dummy_magic_23_0.Vb1.n33 176.733
R7004 two_stage_opamp_dummy_magic_23_0.Vb1.n5 two_stage_opamp_dummy_magic_23_0.Vb1.t28 167.769
R7005 two_stage_opamp_dummy_magic_23_0.Vb1.n1 two_stage_opamp_dummy_magic_23_0.Vb1.n10 161.3
R7006 two_stage_opamp_dummy_magic_23_0.Vb1.n14 two_stage_opamp_dummy_magic_23_0.Vb1.n13 49.3505
R7007 two_stage_opamp_dummy_magic_23_0.Vb1.n1 two_stage_opamp_dummy_magic_23_0.Vb1.n11 49.3505
R7008 two_stage_opamp_dummy_magic_23_0.Vb1.n7 two_stage_opamp_dummy_magic_23_0.Vb1.n6 49.3505
R7009 two_stage_opamp_dummy_magic_23_0.Vb1.n10 two_stage_opamp_dummy_magic_23_0.Vb1.n9 45.5227
R7010 two_stage_opamp_dummy_magic_23_0.Vb1.n10 two_stage_opamp_dummy_magic_23_0.Vb1.n8 45.5227
R7011 bgr_11_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_23_0.Vb1.n35 40.7922
R7012 two_stage_opamp_dummy_magic_23_0.Vb1.n3 two_stage_opamp_dummy_magic_23_0.Vb1.t1 39.4005
R7013 two_stage_opamp_dummy_magic_23_0.Vb1.n3 two_stage_opamp_dummy_magic_23_0.Vb1.t2 39.4005
R7014 two_stage_opamp_dummy_magic_23_0.Vb1.n2 two_stage_opamp_dummy_magic_23_0.Vb1.t3 39.4005
R7015 two_stage_opamp_dummy_magic_23_0.Vb1.n2 two_stage_opamp_dummy_magic_23_0.Vb1.t0 39.4005
R7016 two_stage_opamp_dummy_magic_23_0.Vb1.n35 two_stage_opamp_dummy_magic_23_0.Vb1.n15 17.8547
R7017 two_stage_opamp_dummy_magic_23_0.Vb1.n13 two_stage_opamp_dummy_magic_23_0.Vb1.t13 16.0005
R7018 two_stage_opamp_dummy_magic_23_0.Vb1.n13 two_stage_opamp_dummy_magic_23_0.Vb1.t4 16.0005
R7019 two_stage_opamp_dummy_magic_23_0.Vb1.n11 two_stage_opamp_dummy_magic_23_0.Vb1.t11 16.0005
R7020 two_stage_opamp_dummy_magic_23_0.Vb1.n11 two_stage_opamp_dummy_magic_23_0.Vb1.t7 16.0005
R7021 two_stage_opamp_dummy_magic_23_0.Vb1.n6 two_stage_opamp_dummy_magic_23_0.Vb1.t5 16.0005
R7022 two_stage_opamp_dummy_magic_23_0.Vb1.n6 two_stage_opamp_dummy_magic_23_0.Vb1.t9 16.0005
R7023 bgr_11_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_23_0.Vb1.n4 12.1255
R7024 two_stage_opamp_dummy_magic_23_0.Vb1.n14 two_stage_opamp_dummy_magic_23_0.Vb1.n12 5.6255
R7025 two_stage_opamp_dummy_magic_23_0.Vb1.n12 two_stage_opamp_dummy_magic_23_0.Vb1.n7 5.6255
R7026 two_stage_opamp_dummy_magic_23_0.Vb1.n12 two_stage_opamp_dummy_magic_23_0.Vb1.n1 5.063
R7027 two_stage_opamp_dummy_magic_23_0.Vb1.n7 two_stage_opamp_dummy_magic_23_0.Vb1.n5 4.938
R7028 two_stage_opamp_dummy_magic_23_0.Vb1.n15 two_stage_opamp_dummy_magic_23_0.Vb1.n14 4.938
R7029 two_stage_opamp_dummy_magic_23_0.Vb1.n1 two_stage_opamp_dummy_magic_23_0.Vb1.n0 4.938
R7030 two_stage_opamp_dummy_magic_23_0.Vb1.n5 two_stage_opamp_dummy_magic_23_0.Vb1.n0 0.563
R7031 two_stage_opamp_dummy_magic_23_0.Vb1.n15 two_stage_opamp_dummy_magic_23_0.Vb1.n0 0.563
R7032 two_stage_opamp_dummy_magic_23_0.X.n27 two_stage_opamp_dummy_magic_23_0.X.t46 1172.87
R7033 two_stage_opamp_dummy_magic_23_0.X.n21 two_stage_opamp_dummy_magic_23_0.X.t39 1172.87
R7034 two_stage_opamp_dummy_magic_23_0.X.n27 two_stage_opamp_dummy_magic_23_0.X.t31 996.134
R7035 two_stage_opamp_dummy_magic_23_0.X.n28 two_stage_opamp_dummy_magic_23_0.X.t48 996.134
R7036 two_stage_opamp_dummy_magic_23_0.X.n26 two_stage_opamp_dummy_magic_23_0.X.t34 996.134
R7037 two_stage_opamp_dummy_magic_23_0.X.n25 two_stage_opamp_dummy_magic_23_0.X.t51 996.134
R7038 two_stage_opamp_dummy_magic_23_0.X.n24 two_stage_opamp_dummy_magic_23_0.X.t37 996.134
R7039 two_stage_opamp_dummy_magic_23_0.X.n23 two_stage_opamp_dummy_magic_23_0.X.t53 996.134
R7040 two_stage_opamp_dummy_magic_23_0.X.n22 two_stage_opamp_dummy_magic_23_0.X.t36 996.134
R7041 two_stage_opamp_dummy_magic_23_0.X.n21 two_stage_opamp_dummy_magic_23_0.X.t52 996.134
R7042 two_stage_opamp_dummy_magic_23_0.X.n62 two_stage_opamp_dummy_magic_23_0.X.t41 690.867
R7043 two_stage_opamp_dummy_magic_23_0.X.n61 two_stage_opamp_dummy_magic_23_0.X.t35 690.867
R7044 two_stage_opamp_dummy_magic_23_0.X.n53 two_stage_opamp_dummy_magic_23_0.X.t38 530.201
R7045 two_stage_opamp_dummy_magic_23_0.X.n52 two_stage_opamp_dummy_magic_23_0.X.t30 530.201
R7046 two_stage_opamp_dummy_magic_23_0.X.n68 two_stage_opamp_dummy_magic_23_0.X.t32 514.134
R7047 two_stage_opamp_dummy_magic_23_0.X.n67 two_stage_opamp_dummy_magic_23_0.X.t50 514.134
R7048 two_stage_opamp_dummy_magic_23_0.X.n66 two_stage_opamp_dummy_magic_23_0.X.t33 514.134
R7049 two_stage_opamp_dummy_magic_23_0.X.n65 two_stage_opamp_dummy_magic_23_0.X.t47 514.134
R7050 two_stage_opamp_dummy_magic_23_0.X.n64 two_stage_opamp_dummy_magic_23_0.X.t29 514.134
R7051 two_stage_opamp_dummy_magic_23_0.X.n63 two_stage_opamp_dummy_magic_23_0.X.t43 514.134
R7052 two_stage_opamp_dummy_magic_23_0.X.n62 two_stage_opamp_dummy_magic_23_0.X.t26 514.134
R7053 two_stage_opamp_dummy_magic_23_0.X.n61 two_stage_opamp_dummy_magic_23_0.X.t49 514.134
R7054 two_stage_opamp_dummy_magic_23_0.X.n53 two_stage_opamp_dummy_magic_23_0.X.t54 353.467
R7055 two_stage_opamp_dummy_magic_23_0.X.n54 two_stage_opamp_dummy_magic_23_0.X.t40 353.467
R7056 two_stage_opamp_dummy_magic_23_0.X.n55 two_stage_opamp_dummy_magic_23_0.X.t25 353.467
R7057 two_stage_opamp_dummy_magic_23_0.X.n56 two_stage_opamp_dummy_magic_23_0.X.t42 353.467
R7058 two_stage_opamp_dummy_magic_23_0.X.n57 two_stage_opamp_dummy_magic_23_0.X.t28 353.467
R7059 two_stage_opamp_dummy_magic_23_0.X.n58 two_stage_opamp_dummy_magic_23_0.X.t45 353.467
R7060 two_stage_opamp_dummy_magic_23_0.X.n59 two_stage_opamp_dummy_magic_23_0.X.t27 353.467
R7061 two_stage_opamp_dummy_magic_23_0.X.n52 two_stage_opamp_dummy_magic_23_0.X.t44 353.467
R7062 two_stage_opamp_dummy_magic_23_0.X.n30 two_stage_opamp_dummy_magic_23_0.X.n29 304.375
R7063 two_stage_opamp_dummy_magic_23_0.X.n70 two_stage_opamp_dummy_magic_23_0.X.n60 216.9
R7064 two_stage_opamp_dummy_magic_23_0.X.n70 two_stage_opamp_dummy_magic_23_0.X.n69 216.9
R7065 two_stage_opamp_dummy_magic_23_0.X.n26 two_stage_opamp_dummy_magic_23_0.X.n25 176.733
R7066 two_stage_opamp_dummy_magic_23_0.X.n25 two_stage_opamp_dummy_magic_23_0.X.n24 176.733
R7067 two_stage_opamp_dummy_magic_23_0.X.n24 two_stage_opamp_dummy_magic_23_0.X.n23 176.733
R7068 two_stage_opamp_dummy_magic_23_0.X.n23 two_stage_opamp_dummy_magic_23_0.X.n22 176.733
R7069 two_stage_opamp_dummy_magic_23_0.X.n22 two_stage_opamp_dummy_magic_23_0.X.n21 176.733
R7070 two_stage_opamp_dummy_magic_23_0.X.n28 two_stage_opamp_dummy_magic_23_0.X.n27 176.733
R7071 two_stage_opamp_dummy_magic_23_0.X.n54 two_stage_opamp_dummy_magic_23_0.X.n53 176.733
R7072 two_stage_opamp_dummy_magic_23_0.X.n55 two_stage_opamp_dummy_magic_23_0.X.n54 176.733
R7073 two_stage_opamp_dummy_magic_23_0.X.n56 two_stage_opamp_dummy_magic_23_0.X.n55 176.733
R7074 two_stage_opamp_dummy_magic_23_0.X.n57 two_stage_opamp_dummy_magic_23_0.X.n56 176.733
R7075 two_stage_opamp_dummy_magic_23_0.X.n58 two_stage_opamp_dummy_magic_23_0.X.n57 176.733
R7076 two_stage_opamp_dummy_magic_23_0.X.n59 two_stage_opamp_dummy_magic_23_0.X.n58 176.733
R7077 two_stage_opamp_dummy_magic_23_0.X.n63 two_stage_opamp_dummy_magic_23_0.X.n62 176.733
R7078 two_stage_opamp_dummy_magic_23_0.X.n64 two_stage_opamp_dummy_magic_23_0.X.n63 176.733
R7079 two_stage_opamp_dummy_magic_23_0.X.n65 two_stage_opamp_dummy_magic_23_0.X.n64 176.733
R7080 two_stage_opamp_dummy_magic_23_0.X.n66 two_stage_opamp_dummy_magic_23_0.X.n65 176.733
R7081 two_stage_opamp_dummy_magic_23_0.X.n67 two_stage_opamp_dummy_magic_23_0.X.n66 176.733
R7082 two_stage_opamp_dummy_magic_23_0.X.n68 two_stage_opamp_dummy_magic_23_0.X.n67 176.733
R7083 two_stage_opamp_dummy_magic_23_0.X.n71 two_stage_opamp_dummy_magic_23_0.X.n70 175.05
R7084 two_stage_opamp_dummy_magic_23_0.X.n32 two_stage_opamp_dummy_magic_23_0.X.n31 66.0338
R7085 two_stage_opamp_dummy_magic_23_0.X.n36 two_stage_opamp_dummy_magic_23_0.X.n35 66.0338
R7086 two_stage_opamp_dummy_magic_23_0.X.n38 two_stage_opamp_dummy_magic_23_0.X.n37 66.0338
R7087 two_stage_opamp_dummy_magic_23_0.X.n42 two_stage_opamp_dummy_magic_23_0.X.n41 66.0338
R7088 two_stage_opamp_dummy_magic_23_0.X.n45 two_stage_opamp_dummy_magic_23_0.X.n44 66.0338
R7089 two_stage_opamp_dummy_magic_23_0.X.n49 two_stage_opamp_dummy_magic_23_0.X.n48 66.0338
R7090 two_stage_opamp_dummy_magic_23_0.X.n30 two_stage_opamp_dummy_magic_23_0.X.t7 49.4481
R7091 two_stage_opamp_dummy_magic_23_0.X.n1 two_stage_opamp_dummy_magic_23_0.X.n0 49.3505
R7092 two_stage_opamp_dummy_magic_23_0.X.n5 two_stage_opamp_dummy_magic_23_0.X.n4 49.3505
R7093 two_stage_opamp_dummy_magic_23_0.X.n7 two_stage_opamp_dummy_magic_23_0.X.n6 49.3505
R7094 two_stage_opamp_dummy_magic_23_0.X.n11 two_stage_opamp_dummy_magic_23_0.X.n10 49.3505
R7095 two_stage_opamp_dummy_magic_23_0.X.n13 two_stage_opamp_dummy_magic_23_0.X.n12 49.3505
R7096 two_stage_opamp_dummy_magic_23_0.X.n17 two_stage_opamp_dummy_magic_23_0.X.n16 49.3505
R7097 two_stage_opamp_dummy_magic_23_0.X.n29 two_stage_opamp_dummy_magic_23_0.X.n26 40.1672
R7098 two_stage_opamp_dummy_magic_23_0.X.n29 two_stage_opamp_dummy_magic_23_0.X.n28 40.1672
R7099 two_stage_opamp_dummy_magic_23_0.X.n60 two_stage_opamp_dummy_magic_23_0.X.n52 40.1672
R7100 two_stage_opamp_dummy_magic_23_0.X.n60 two_stage_opamp_dummy_magic_23_0.X.n59 40.1672
R7101 two_stage_opamp_dummy_magic_23_0.X.n69 two_stage_opamp_dummy_magic_23_0.X.n61 40.1672
R7102 two_stage_opamp_dummy_magic_23_0.X.n69 two_stage_opamp_dummy_magic_23_0.X.n68 40.1672
R7103 two_stage_opamp_dummy_magic_23_0.X.n71 two_stage_opamp_dummy_magic_23_0.X.n51 17.688
R7104 two_stage_opamp_dummy_magic_23_0.X.n0 two_stage_opamp_dummy_magic_23_0.X.t16 16.0005
R7105 two_stage_opamp_dummy_magic_23_0.X.n0 two_stage_opamp_dummy_magic_23_0.X.t24 16.0005
R7106 two_stage_opamp_dummy_magic_23_0.X.n4 two_stage_opamp_dummy_magic_23_0.X.t14 16.0005
R7107 two_stage_opamp_dummy_magic_23_0.X.n4 two_stage_opamp_dummy_magic_23_0.X.t19 16.0005
R7108 two_stage_opamp_dummy_magic_23_0.X.n6 two_stage_opamp_dummy_magic_23_0.X.t22 16.0005
R7109 two_stage_opamp_dummy_magic_23_0.X.n6 two_stage_opamp_dummy_magic_23_0.X.t18 16.0005
R7110 two_stage_opamp_dummy_magic_23_0.X.n10 two_stage_opamp_dummy_magic_23_0.X.t20 16.0005
R7111 two_stage_opamp_dummy_magic_23_0.X.n10 two_stage_opamp_dummy_magic_23_0.X.t13 16.0005
R7112 two_stage_opamp_dummy_magic_23_0.X.n12 two_stage_opamp_dummy_magic_23_0.X.t15 16.0005
R7113 two_stage_opamp_dummy_magic_23_0.X.n12 two_stage_opamp_dummy_magic_23_0.X.t23 16.0005
R7114 two_stage_opamp_dummy_magic_23_0.X.n16 two_stage_opamp_dummy_magic_23_0.X.t21 16.0005
R7115 two_stage_opamp_dummy_magic_23_0.X.n16 two_stage_opamp_dummy_magic_23_0.X.t17 16.0005
R7116 two_stage_opamp_dummy_magic_23_0.X.n31 two_stage_opamp_dummy_magic_23_0.X.t3 11.2576
R7117 two_stage_opamp_dummy_magic_23_0.X.n31 two_stage_opamp_dummy_magic_23_0.X.t11 11.2576
R7118 two_stage_opamp_dummy_magic_23_0.X.n35 two_stage_opamp_dummy_magic_23_0.X.t8 11.2576
R7119 two_stage_opamp_dummy_magic_23_0.X.n35 two_stage_opamp_dummy_magic_23_0.X.t4 11.2576
R7120 two_stage_opamp_dummy_magic_23_0.X.n37 two_stage_opamp_dummy_magic_23_0.X.t1 11.2576
R7121 two_stage_opamp_dummy_magic_23_0.X.n37 two_stage_opamp_dummy_magic_23_0.X.t5 11.2576
R7122 two_stage_opamp_dummy_magic_23_0.X.n41 two_stage_opamp_dummy_magic_23_0.X.t2 11.2576
R7123 two_stage_opamp_dummy_magic_23_0.X.n41 two_stage_opamp_dummy_magic_23_0.X.t6 11.2576
R7124 two_stage_opamp_dummy_magic_23_0.X.n44 two_stage_opamp_dummy_magic_23_0.X.t12 11.2576
R7125 two_stage_opamp_dummy_magic_23_0.X.n44 two_stage_opamp_dummy_magic_23_0.X.t10 11.2576
R7126 two_stage_opamp_dummy_magic_23_0.X.n48 two_stage_opamp_dummy_magic_23_0.X.t0 11.2576
R7127 two_stage_opamp_dummy_magic_23_0.X.n48 two_stage_opamp_dummy_magic_23_0.X.t9 11.2576
R7128 two_stage_opamp_dummy_magic_23_0.X.n73 two_stage_opamp_dummy_magic_23_0.X.n72 8.09425
R7129 two_stage_opamp_dummy_magic_23_0.X.n39 two_stage_opamp_dummy_magic_23_0.X.n36 5.91717
R7130 two_stage_opamp_dummy_magic_23_0.X.n36 two_stage_opamp_dummy_magic_23_0.X.n34 5.91717
R7131 two_stage_opamp_dummy_magic_23_0.X.n47 two_stage_opamp_dummy_magic_23_0.X.n32 5.91717
R7132 two_stage_opamp_dummy_magic_23_0.X.n14 two_stage_opamp_dummy_magic_23_0.X.n11 5.6255
R7133 two_stage_opamp_dummy_magic_23_0.X.n8 two_stage_opamp_dummy_magic_23_0.X.n5 5.6255
R7134 two_stage_opamp_dummy_magic_23_0.X.n11 two_stage_opamp_dummy_magic_23_0.X.n3 5.438
R7135 two_stage_opamp_dummy_magic_23_0.X.n5 two_stage_opamp_dummy_magic_23_0.X.n2 5.438
R7136 two_stage_opamp_dummy_magic_23_0.X.n38 two_stage_opamp_dummy_magic_23_0.X.n34 5.29217
R7137 two_stage_opamp_dummy_magic_23_0.X.n39 two_stage_opamp_dummy_magic_23_0.X.n38 5.29217
R7138 two_stage_opamp_dummy_magic_23_0.X.n43 two_stage_opamp_dummy_magic_23_0.X.n42 5.29217
R7139 two_stage_opamp_dummy_magic_23_0.X.n42 two_stage_opamp_dummy_magic_23_0.X.n40 5.29217
R7140 two_stage_opamp_dummy_magic_23_0.X.n46 two_stage_opamp_dummy_magic_23_0.X.n45 5.29217
R7141 two_stage_opamp_dummy_magic_23_0.X.n45 two_stage_opamp_dummy_magic_23_0.X.n33 5.29217
R7142 two_stage_opamp_dummy_magic_23_0.X.n49 two_stage_opamp_dummy_magic_23_0.X.n47 5.29217
R7143 two_stage_opamp_dummy_magic_23_0.X.n50 two_stage_opamp_dummy_magic_23_0.X.n49 5.29217
R7144 two_stage_opamp_dummy_magic_23_0.X.n51 two_stage_opamp_dummy_magic_23_0.X.n50 5.1255
R7145 two_stage_opamp_dummy_magic_23_0.X.n8 two_stage_opamp_dummy_magic_23_0.X.n7 5.063
R7146 two_stage_opamp_dummy_magic_23_0.X.n14 two_stage_opamp_dummy_magic_23_0.X.n13 5.063
R7147 two_stage_opamp_dummy_magic_23_0.X.n17 two_stage_opamp_dummy_magic_23_0.X.n15 5.063
R7148 two_stage_opamp_dummy_magic_23_0.X.n9 two_stage_opamp_dummy_magic_23_0.X.n1 5.063
R7149 two_stage_opamp_dummy_magic_23_0.X.n7 two_stage_opamp_dummy_magic_23_0.X.n2 4.8755
R7150 two_stage_opamp_dummy_magic_23_0.X.n13 two_stage_opamp_dummy_magic_23_0.X.n3 4.8755
R7151 two_stage_opamp_dummy_magic_23_0.X.n18 two_stage_opamp_dummy_magic_23_0.X.n17 4.8755
R7152 two_stage_opamp_dummy_magic_23_0.X.n20 two_stage_opamp_dummy_magic_23_0.X.n19 4.5005
R7153 two_stage_opamp_dummy_magic_23_0.X.n72 two_stage_opamp_dummy_magic_23_0.X.n71 4.5005
R7154 two_stage_opamp_dummy_magic_23_0.X.n72 two_stage_opamp_dummy_magic_23_0.X.n30 3.27133
R7155 two_stage_opamp_dummy_magic_23_0.X.n73 two_stage_opamp_dummy_magic_23_0.X.n20 2.15675
R7156 two_stage_opamp_dummy_magic_23_0.X.n51 two_stage_opamp_dummy_magic_23_0.X.n32 0.792167
R7157 two_stage_opamp_dummy_magic_23_0.X.n50 two_stage_opamp_dummy_magic_23_0.X.n33 0.6255
R7158 two_stage_opamp_dummy_magic_23_0.X.n40 two_stage_opamp_dummy_magic_23_0.X.n33 0.6255
R7159 two_stage_opamp_dummy_magic_23_0.X.n40 two_stage_opamp_dummy_magic_23_0.X.n39 0.6255
R7160 two_stage_opamp_dummy_magic_23_0.X.n43 two_stage_opamp_dummy_magic_23_0.X.n34 0.6255
R7161 two_stage_opamp_dummy_magic_23_0.X.n46 two_stage_opamp_dummy_magic_23_0.X.n43 0.6255
R7162 two_stage_opamp_dummy_magic_23_0.X.n47 two_stage_opamp_dummy_magic_23_0.X.n46 0.6255
R7163 two_stage_opamp_dummy_magic_23_0.X.n15 two_stage_opamp_dummy_magic_23_0.X.n9 0.563
R7164 two_stage_opamp_dummy_magic_23_0.X.n15 two_stage_opamp_dummy_magic_23_0.X.n14 0.563
R7165 two_stage_opamp_dummy_magic_23_0.X.n18 two_stage_opamp_dummy_magic_23_0.X.n3 0.563
R7166 two_stage_opamp_dummy_magic_23_0.X.n19 two_stage_opamp_dummy_magic_23_0.X.n18 0.563
R7167 two_stage_opamp_dummy_magic_23_0.X.n19 two_stage_opamp_dummy_magic_23_0.X.n2 0.563
R7168 two_stage_opamp_dummy_magic_23_0.X.n9 two_stage_opamp_dummy_magic_23_0.X.n8 0.563
R7169 two_stage_opamp_dummy_magic_23_0.X.n20 two_stage_opamp_dummy_magic_23_0.X.n1 0.3755
R7170 two_stage_opamp_dummy_magic_23_0.X two_stage_opamp_dummy_magic_23_0.X.n73 0.063
R7171 two_stage_opamp_dummy_magic_23_0.VD1.n3 two_stage_opamp_dummy_magic_23_0.VD1.n2 49.3505
R7172 two_stage_opamp_dummy_magic_23_0.VD1.n5 two_stage_opamp_dummy_magic_23_0.VD1.n4 49.3505
R7173 two_stage_opamp_dummy_magic_23_0.VD1.n9 two_stage_opamp_dummy_magic_23_0.VD1.n8 49.3505
R7174 two_stage_opamp_dummy_magic_23_0.VD1.n13 two_stage_opamp_dummy_magic_23_0.VD1.n12 49.3505
R7175 two_stage_opamp_dummy_magic_23_0.VD1.n16 two_stage_opamp_dummy_magic_23_0.VD1.n15 49.3505
R7176 two_stage_opamp_dummy_magic_23_0.VD1.n19 two_stage_opamp_dummy_magic_23_0.VD1.n18 49.3505
R7177 two_stage_opamp_dummy_magic_23_0.VD1.n22 two_stage_opamp_dummy_magic_23_0.VD1.n21 49.3505
R7178 two_stage_opamp_dummy_magic_23_0.VD1.n24 two_stage_opamp_dummy_magic_23_0.VD1.n23 49.3505
R7179 two_stage_opamp_dummy_magic_23_0.VD1.n28 two_stage_opamp_dummy_magic_23_0.VD1.n27 49.3505
R7180 two_stage_opamp_dummy_magic_23_0.VD1.n34 two_stage_opamp_dummy_magic_23_0.VD1.n33 49.3505
R7181 two_stage_opamp_dummy_magic_23_0.VD1.n37 two_stage_opamp_dummy_magic_23_0.VD1.n36 49.3505
R7182 two_stage_opamp_dummy_magic_23_0.VD1.n2 two_stage_opamp_dummy_magic_23_0.VD1.t18 16.0005
R7183 two_stage_opamp_dummy_magic_23_0.VD1.n2 two_stage_opamp_dummy_magic_23_0.VD1.t13 16.0005
R7184 two_stage_opamp_dummy_magic_23_0.VD1.n4 two_stage_opamp_dummy_magic_23_0.VD1.t17 16.0005
R7185 two_stage_opamp_dummy_magic_23_0.VD1.n4 two_stage_opamp_dummy_magic_23_0.VD1.t21 16.0005
R7186 two_stage_opamp_dummy_magic_23_0.VD1.n8 two_stage_opamp_dummy_magic_23_0.VD1.t15 16.0005
R7187 two_stage_opamp_dummy_magic_23_0.VD1.n8 two_stage_opamp_dummy_magic_23_0.VD1.t12 16.0005
R7188 two_stage_opamp_dummy_magic_23_0.VD1.n12 two_stage_opamp_dummy_magic_23_0.VD1.t10 16.0005
R7189 two_stage_opamp_dummy_magic_23_0.VD1.n12 two_stage_opamp_dummy_magic_23_0.VD1.t6 16.0005
R7190 two_stage_opamp_dummy_magic_23_0.VD1.n15 two_stage_opamp_dummy_magic_23_0.VD1.t2 16.0005
R7191 two_stage_opamp_dummy_magic_23_0.VD1.n15 two_stage_opamp_dummy_magic_23_0.VD1.t8 16.0005
R7192 two_stage_opamp_dummy_magic_23_0.VD1.n18 two_stage_opamp_dummy_magic_23_0.VD1.t7 16.0005
R7193 two_stage_opamp_dummy_magic_23_0.VD1.n18 two_stage_opamp_dummy_magic_23_0.VD1.t1 16.0005
R7194 two_stage_opamp_dummy_magic_23_0.VD1.n21 two_stage_opamp_dummy_magic_23_0.VD1.t4 16.0005
R7195 two_stage_opamp_dummy_magic_23_0.VD1.n21 two_stage_opamp_dummy_magic_23_0.VD1.t9 16.0005
R7196 two_stage_opamp_dummy_magic_23_0.VD1.n23 two_stage_opamp_dummy_magic_23_0.VD1.t5 16.0005
R7197 two_stage_opamp_dummy_magic_23_0.VD1.n23 two_stage_opamp_dummy_magic_23_0.VD1.t11 16.0005
R7198 two_stage_opamp_dummy_magic_23_0.VD1.n27 two_stage_opamp_dummy_magic_23_0.VD1.t3 16.0005
R7199 two_stage_opamp_dummy_magic_23_0.VD1.n27 two_stage_opamp_dummy_magic_23_0.VD1.t0 16.0005
R7200 two_stage_opamp_dummy_magic_23_0.VD1.n33 two_stage_opamp_dummy_magic_23_0.VD1.t14 16.0005
R7201 two_stage_opamp_dummy_magic_23_0.VD1.n33 two_stage_opamp_dummy_magic_23_0.VD1.t19 16.0005
R7202 two_stage_opamp_dummy_magic_23_0.VD1.n37 two_stage_opamp_dummy_magic_23_0.VD1.t16 16.0005
R7203 two_stage_opamp_dummy_magic_23_0.VD1.t20 two_stage_opamp_dummy_magic_23_0.VD1.n37 16.0005
R7204 two_stage_opamp_dummy_magic_23_0.VD1.n31 two_stage_opamp_dummy_magic_23_0.VD1.n30 5.77133
R7205 two_stage_opamp_dummy_magic_23_0.VD1.n22 two_stage_opamp_dummy_magic_23_0.VD1.n11 5.64633
R7206 two_stage_opamp_dummy_magic_23_0.VD1.n14 two_stage_opamp_dummy_magic_23_0.VD1.n13 5.64633
R7207 two_stage_opamp_dummy_magic_23_0.VD1.n34 two_stage_opamp_dummy_magic_23_0.VD1.n0 5.6255
R7208 two_stage_opamp_dummy_magic_23_0.VD1.n6 two_stage_opamp_dummy_magic_23_0.VD1.n3 5.6255
R7209 two_stage_opamp_dummy_magic_23_0.VD1.n25 two_stage_opamp_dummy_magic_23_0.VD1.n22 5.438
R7210 two_stage_opamp_dummy_magic_23_0.VD1.n17 two_stage_opamp_dummy_magic_23_0.VD1.n13 5.438
R7211 two_stage_opamp_dummy_magic_23_0.VD1.n35 two_stage_opamp_dummy_magic_23_0.VD1.n34 5.438
R7212 two_stage_opamp_dummy_magic_23_0.VD1.n3 two_stage_opamp_dummy_magic_23_0.VD1.n1 5.438
R7213 two_stage_opamp_dummy_magic_23_0.VD1.n16 two_stage_opamp_dummy_magic_23_0.VD1.n14 5.08383
R7214 two_stage_opamp_dummy_magic_23_0.VD1.n19 two_stage_opamp_dummy_magic_23_0.VD1.n10 5.08383
R7215 two_stage_opamp_dummy_magic_23_0.VD1.n24 two_stage_opamp_dummy_magic_23_0.VD1.n11 5.08383
R7216 two_stage_opamp_dummy_magic_23_0.VD1.n29 two_stage_opamp_dummy_magic_23_0.VD1.n28 5.08383
R7217 two_stage_opamp_dummy_magic_23_0.VD1.n6 two_stage_opamp_dummy_magic_23_0.VD1.n5 5.063
R7218 two_stage_opamp_dummy_magic_23_0.VD1.n9 two_stage_opamp_dummy_magic_23_0.VD1.n7 5.063
R7219 two_stage_opamp_dummy_magic_23_0.VD1.n36 two_stage_opamp_dummy_magic_23_0.VD1.n0 5.063
R7220 two_stage_opamp_dummy_magic_23_0.VD1.n5 two_stage_opamp_dummy_magic_23_0.VD1.n1 4.8755
R7221 two_stage_opamp_dummy_magic_23_0.VD1.n17 two_stage_opamp_dummy_magic_23_0.VD1.n16 4.8755
R7222 two_stage_opamp_dummy_magic_23_0.VD1.n20 two_stage_opamp_dummy_magic_23_0.VD1.n19 4.8755
R7223 two_stage_opamp_dummy_magic_23_0.VD1.n25 two_stage_opamp_dummy_magic_23_0.VD1.n24 4.8755
R7224 two_stage_opamp_dummy_magic_23_0.VD1.n28 two_stage_opamp_dummy_magic_23_0.VD1.n26 4.8755
R7225 two_stage_opamp_dummy_magic_23_0.VD1.n36 two_stage_opamp_dummy_magic_23_0.VD1.n35 4.8755
R7226 two_stage_opamp_dummy_magic_23_0.VD1.n32 two_stage_opamp_dummy_magic_23_0.VD1.n31 4.5005
R7227 two_stage_opamp_dummy_magic_23_0.VD1.n29 two_stage_opamp_dummy_magic_23_0.VD1.n11 0.563
R7228 two_stage_opamp_dummy_magic_23_0.VD1.n26 two_stage_opamp_dummy_magic_23_0.VD1.n25 0.563
R7229 two_stage_opamp_dummy_magic_23_0.VD1.n26 two_stage_opamp_dummy_magic_23_0.VD1.n20 0.563
R7230 two_stage_opamp_dummy_magic_23_0.VD1.n20 two_stage_opamp_dummy_magic_23_0.VD1.n17 0.563
R7231 two_stage_opamp_dummy_magic_23_0.VD1.n14 two_stage_opamp_dummy_magic_23_0.VD1.n10 0.563
R7232 two_stage_opamp_dummy_magic_23_0.VD1.n7 two_stage_opamp_dummy_magic_23_0.VD1.n0 0.563
R7233 two_stage_opamp_dummy_magic_23_0.VD1.n7 two_stage_opamp_dummy_magic_23_0.VD1.n6 0.563
R7234 two_stage_opamp_dummy_magic_23_0.VD1.n32 two_stage_opamp_dummy_magic_23_0.VD1.n1 0.563
R7235 two_stage_opamp_dummy_magic_23_0.VD1.n35 two_stage_opamp_dummy_magic_23_0.VD1.n32 0.563
R7236 two_stage_opamp_dummy_magic_23_0.VD1.n31 two_stage_opamp_dummy_magic_23_0.VD1.n9 0.3755
R7237 two_stage_opamp_dummy_magic_23_0.VD1.n30 two_stage_opamp_dummy_magic_23_0.VD1.n29 0.234875
R7238 two_stage_opamp_dummy_magic_23_0.VD1.n30 two_stage_opamp_dummy_magic_23_0.VD1.n10 0.234875
R7239 two_stage_opamp_dummy_magic_23_0.Vb2.n7 two_stage_opamp_dummy_magic_23_0.Vb2.t15 746.673
R7240 two_stage_opamp_dummy_magic_23_0.Vb2.n29 two_stage_opamp_dummy_magic_23_0.Vb2.t9 721.625
R7241 two_stage_opamp_dummy_magic_23_0.Vb2.n21 two_stage_opamp_dummy_magic_23_0.Vb2.t30 611.739
R7242 two_stage_opamp_dummy_magic_23_0.Vb2.n17 two_stage_opamp_dummy_magic_23_0.Vb2.t24 611.739
R7243 two_stage_opamp_dummy_magic_23_0.Vb2.n12 two_stage_opamp_dummy_magic_23_0.Vb2.t19 611.739
R7244 two_stage_opamp_dummy_magic_23_0.Vb2.n8 two_stage_opamp_dummy_magic_23_0.Vb2.t16 611.739
R7245 two_stage_opamp_dummy_magic_23_0.Vb2.n28 two_stage_opamp_dummy_magic_23_0.Vb2.t31 563.451
R7246 two_stage_opamp_dummy_magic_23_0.Vb2.n21 two_stage_opamp_dummy_magic_23_0.Vb2.t27 421.75
R7247 two_stage_opamp_dummy_magic_23_0.Vb2.n22 two_stage_opamp_dummy_magic_23_0.Vb2.t22 421.75
R7248 two_stage_opamp_dummy_magic_23_0.Vb2.n23 two_stage_opamp_dummy_magic_23_0.Vb2.t18 421.75
R7249 two_stage_opamp_dummy_magic_23_0.Vb2.n24 two_stage_opamp_dummy_magic_23_0.Vb2.t12 421.75
R7250 two_stage_opamp_dummy_magic_23_0.Vb2.n17 two_stage_opamp_dummy_magic_23_0.Vb2.t20 421.75
R7251 two_stage_opamp_dummy_magic_23_0.Vb2.n18 two_stage_opamp_dummy_magic_23_0.Vb2.t25 421.75
R7252 two_stage_opamp_dummy_magic_23_0.Vb2.n19 two_stage_opamp_dummy_magic_23_0.Vb2.t29 421.75
R7253 two_stage_opamp_dummy_magic_23_0.Vb2.n20 two_stage_opamp_dummy_magic_23_0.Vb2.t32 421.75
R7254 two_stage_opamp_dummy_magic_23_0.Vb2.n12 two_stage_opamp_dummy_magic_23_0.Vb2.t14 421.75
R7255 two_stage_opamp_dummy_magic_23_0.Vb2.n13 two_stage_opamp_dummy_magic_23_0.Vb2.t17 421.75
R7256 two_stage_opamp_dummy_magic_23_0.Vb2.n14 two_stage_opamp_dummy_magic_23_0.Vb2.t13 421.75
R7257 two_stage_opamp_dummy_magic_23_0.Vb2.n15 two_stage_opamp_dummy_magic_23_0.Vb2.t11 421.75
R7258 two_stage_opamp_dummy_magic_23_0.Vb2.n8 two_stage_opamp_dummy_magic_23_0.Vb2.t21 421.75
R7259 two_stage_opamp_dummy_magic_23_0.Vb2.n9 two_stage_opamp_dummy_magic_23_0.Vb2.t26 421.75
R7260 two_stage_opamp_dummy_magic_23_0.Vb2.n10 two_stage_opamp_dummy_magic_23_0.Vb2.t23 421.75
R7261 two_stage_opamp_dummy_magic_23_0.Vb2.n11 two_stage_opamp_dummy_magic_23_0.Vb2.t28 421.75
R7262 two_stage_opamp_dummy_magic_23_0.Vb2.n26 two_stage_opamp_dummy_magic_23_0.Vb2.n16 313.776
R7263 two_stage_opamp_dummy_magic_23_0.Vb2.n26 two_stage_opamp_dummy_magic_23_0.Vb2.n25 313.212
R7264 two_stage_opamp_dummy_magic_23_0.Vb2.n22 two_stage_opamp_dummy_magic_23_0.Vb2.n21 167.094
R7265 two_stage_opamp_dummy_magic_23_0.Vb2.n23 two_stage_opamp_dummy_magic_23_0.Vb2.n22 167.094
R7266 two_stage_opamp_dummy_magic_23_0.Vb2.n24 two_stage_opamp_dummy_magic_23_0.Vb2.n23 167.094
R7267 two_stage_opamp_dummy_magic_23_0.Vb2.n18 two_stage_opamp_dummy_magic_23_0.Vb2.n17 167.094
R7268 two_stage_opamp_dummy_magic_23_0.Vb2.n19 two_stage_opamp_dummy_magic_23_0.Vb2.n18 167.094
R7269 two_stage_opamp_dummy_magic_23_0.Vb2.n20 two_stage_opamp_dummy_magic_23_0.Vb2.n19 167.094
R7270 two_stage_opamp_dummy_magic_23_0.Vb2.n13 two_stage_opamp_dummy_magic_23_0.Vb2.n12 167.094
R7271 two_stage_opamp_dummy_magic_23_0.Vb2.n14 two_stage_opamp_dummy_magic_23_0.Vb2.n13 167.094
R7272 two_stage_opamp_dummy_magic_23_0.Vb2.n15 two_stage_opamp_dummy_magic_23_0.Vb2.n14 167.094
R7273 two_stage_opamp_dummy_magic_23_0.Vb2.n9 two_stage_opamp_dummy_magic_23_0.Vb2.n8 167.094
R7274 two_stage_opamp_dummy_magic_23_0.Vb2.n10 two_stage_opamp_dummy_magic_23_0.Vb2.n9 167.094
R7275 two_stage_opamp_dummy_magic_23_0.Vb2.n11 two_stage_opamp_dummy_magic_23_0.Vb2.n10 167.094
R7276 two_stage_opamp_dummy_magic_23_0.Vb2.n2 two_stage_opamp_dummy_magic_23_0.Vb2.n0 140.857
R7277 two_stage_opamp_dummy_magic_23_0.Vb2.n6 two_stage_opamp_dummy_magic_23_0.Vb2.n5 139.608
R7278 two_stage_opamp_dummy_magic_23_0.Vb2.n4 two_stage_opamp_dummy_magic_23_0.Vb2.n3 139.608
R7279 two_stage_opamp_dummy_magic_23_0.Vb2.n2 two_stage_opamp_dummy_magic_23_0.Vb2.n1 139.608
R7280 two_stage_opamp_dummy_magic_23_0.Vb2.n30 two_stage_opamp_dummy_magic_23_0.Vb2.n29 67.013
R7281 two_stage_opamp_dummy_magic_23_0.Vb2.n7 two_stage_opamp_dummy_magic_23_0.Vb2.n6 65.9474
R7282 two_stage_opamp_dummy_magic_23_0.Vb2.n25 two_stage_opamp_dummy_magic_23_0.Vb2.n24 35.3472
R7283 two_stage_opamp_dummy_magic_23_0.Vb2.n25 two_stage_opamp_dummy_magic_23_0.Vb2.n20 35.3472
R7284 two_stage_opamp_dummy_magic_23_0.Vb2.n16 two_stage_opamp_dummy_magic_23_0.Vb2.n15 35.3472
R7285 two_stage_opamp_dummy_magic_23_0.Vb2.n16 two_stage_opamp_dummy_magic_23_0.Vb2.n11 35.3472
R7286 two_stage_opamp_dummy_magic_23_0.Vb2.n5 two_stage_opamp_dummy_magic_23_0.Vb2.t7 24.0005
R7287 two_stage_opamp_dummy_magic_23_0.Vb2.n5 two_stage_opamp_dummy_magic_23_0.Vb2.t5 24.0005
R7288 two_stage_opamp_dummy_magic_23_0.Vb2.n3 two_stage_opamp_dummy_magic_23_0.Vb2.t4 24.0005
R7289 two_stage_opamp_dummy_magic_23_0.Vb2.n3 two_stage_opamp_dummy_magic_23_0.Vb2.t6 24.0005
R7290 two_stage_opamp_dummy_magic_23_0.Vb2.n1 two_stage_opamp_dummy_magic_23_0.Vb2.t3 24.0005
R7291 two_stage_opamp_dummy_magic_23_0.Vb2.n1 two_stage_opamp_dummy_magic_23_0.Vb2.t0 24.0005
R7292 two_stage_opamp_dummy_magic_23_0.Vb2.n0 two_stage_opamp_dummy_magic_23_0.Vb2.t1 24.0005
R7293 two_stage_opamp_dummy_magic_23_0.Vb2.n0 two_stage_opamp_dummy_magic_23_0.Vb2.t8 24.0005
R7294 two_stage_opamp_dummy_magic_23_0.Vb2.n27 two_stage_opamp_dummy_magic_23_0.Vb2.n26 13.2817
R7295 two_stage_opamp_dummy_magic_23_0.Vb2.n30 two_stage_opamp_dummy_magic_23_0.Vb2.t10 11.2576
R7296 two_stage_opamp_dummy_magic_23_0.Vb2.t2 two_stage_opamp_dummy_magic_23_0.Vb2.n30 11.2576
R7297 two_stage_opamp_dummy_magic_23_0.Vb2.n4 two_stage_opamp_dummy_magic_23_0.Vb2.n2 7.563
R7298 two_stage_opamp_dummy_magic_23_0.Vb2.n29 two_stage_opamp_dummy_magic_23_0.Vb2.n28 7.35988
R7299 two_stage_opamp_dummy_magic_23_0.Vb2.n27 two_stage_opamp_dummy_magic_23_0.Vb2.n7 4.55362
R7300 two_stage_opamp_dummy_magic_23_0.Vb2.n6 two_stage_opamp_dummy_magic_23_0.Vb2.n4 1.2505
R7301 two_stage_opamp_dummy_magic_23_0.Vb2.n28 two_stage_opamp_dummy_magic_23_0.Vb2.n27 1.14112
R7302 two_stage_opamp_dummy_magic_23_0.VD3.n26 two_stage_opamp_dummy_magic_23_0.VD3.t0 672.293
R7303 two_stage_opamp_dummy_magic_23_0.VD3.n29 two_stage_opamp_dummy_magic_23_0.VD3.t3 672.293
R7304 two_stage_opamp_dummy_magic_23_0.VD3.t1 two_stage_opamp_dummy_magic_23_0.VD3.n27 213.131
R7305 two_stage_opamp_dummy_magic_23_0.VD3.n28 two_stage_opamp_dummy_magic_23_0.VD3.t4 213.131
R7306 two_stage_opamp_dummy_magic_23_0.VD3.t23 two_stage_opamp_dummy_magic_23_0.VD3.t1 146.155
R7307 two_stage_opamp_dummy_magic_23_0.VD3.t29 two_stage_opamp_dummy_magic_23_0.VD3.t23 146.155
R7308 two_stage_opamp_dummy_magic_23_0.VD3.t25 two_stage_opamp_dummy_magic_23_0.VD3.t29 146.155
R7309 two_stage_opamp_dummy_magic_23_0.VD3.t31 two_stage_opamp_dummy_magic_23_0.VD3.t25 146.155
R7310 two_stage_opamp_dummy_magic_23_0.VD3.t33 two_stage_opamp_dummy_magic_23_0.VD3.t31 146.155
R7311 two_stage_opamp_dummy_magic_23_0.VD3.t15 two_stage_opamp_dummy_magic_23_0.VD3.t33 146.155
R7312 two_stage_opamp_dummy_magic_23_0.VD3.t19 two_stage_opamp_dummy_magic_23_0.VD3.t15 146.155
R7313 two_stage_opamp_dummy_magic_23_0.VD3.t17 two_stage_opamp_dummy_magic_23_0.VD3.t19 146.155
R7314 two_stage_opamp_dummy_magic_23_0.VD3.t21 two_stage_opamp_dummy_magic_23_0.VD3.t17 146.155
R7315 two_stage_opamp_dummy_magic_23_0.VD3.t27 two_stage_opamp_dummy_magic_23_0.VD3.t21 146.155
R7316 two_stage_opamp_dummy_magic_23_0.VD3.t4 two_stage_opamp_dummy_magic_23_0.VD3.t27 146.155
R7317 two_stage_opamp_dummy_magic_23_0.VD3.n27 two_stage_opamp_dummy_magic_23_0.VD3.t2 76.2576
R7318 two_stage_opamp_dummy_magic_23_0.VD3.n28 two_stage_opamp_dummy_magic_23_0.VD3.t5 76.2576
R7319 two_stage_opamp_dummy_magic_23_0.VD3.n1 two_stage_opamp_dummy_magic_23_0.VD3.n0 71.513
R7320 two_stage_opamp_dummy_magic_23_0.VD3.n24 two_stage_opamp_dummy_magic_23_0.VD3.n23 71.513
R7321 two_stage_opamp_dummy_magic_23_0.VD3.n31 two_stage_opamp_dummy_magic_23_0.VD3.n30 71.513
R7322 two_stage_opamp_dummy_magic_23_0.VD3.n33 two_stage_opamp_dummy_magic_23_0.VD3.n32 71.513
R7323 two_stage_opamp_dummy_magic_23_0.VD3.n35 two_stage_opamp_dummy_magic_23_0.VD3.n34 71.513
R7324 two_stage_opamp_dummy_magic_23_0.VD3.n5 two_stage_opamp_dummy_magic_23_0.VD3.n4 66.0338
R7325 two_stage_opamp_dummy_magic_23_0.VD3.n8 two_stage_opamp_dummy_magic_23_0.VD3.n7 66.0338
R7326 two_stage_opamp_dummy_magic_23_0.VD3.n11 two_stage_opamp_dummy_magic_23_0.VD3.n10 66.0338
R7327 two_stage_opamp_dummy_magic_23_0.VD3.n15 two_stage_opamp_dummy_magic_23_0.VD3.n14 66.0338
R7328 two_stage_opamp_dummy_magic_23_0.VD3.n18 two_stage_opamp_dummy_magic_23_0.VD3.n17 66.0338
R7329 two_stage_opamp_dummy_magic_23_0.VD3.n21 two_stage_opamp_dummy_magic_23_0.VD3.n20 66.0338
R7330 two_stage_opamp_dummy_magic_23_0.VD3.n25 two_stage_opamp_dummy_magic_23_0.VD3.n22 14.0005
R7331 two_stage_opamp_dummy_magic_23_0.VD3.n0 two_stage_opamp_dummy_magic_23_0.VD3.t26 11.2576
R7332 two_stage_opamp_dummy_magic_23_0.VD3.n0 two_stage_opamp_dummy_magic_23_0.VD3.t32 11.2576
R7333 two_stage_opamp_dummy_magic_23_0.VD3.n23 two_stage_opamp_dummy_magic_23_0.VD3.t24 11.2576
R7334 two_stage_opamp_dummy_magic_23_0.VD3.n23 two_stage_opamp_dummy_magic_23_0.VD3.t30 11.2576
R7335 two_stage_opamp_dummy_magic_23_0.VD3.n30 two_stage_opamp_dummy_magic_23_0.VD3.t22 11.2576
R7336 two_stage_opamp_dummy_magic_23_0.VD3.n30 two_stage_opamp_dummy_magic_23_0.VD3.t28 11.2576
R7337 two_stage_opamp_dummy_magic_23_0.VD3.n32 two_stage_opamp_dummy_magic_23_0.VD3.t20 11.2576
R7338 two_stage_opamp_dummy_magic_23_0.VD3.n32 two_stage_opamp_dummy_magic_23_0.VD3.t18 11.2576
R7339 two_stage_opamp_dummy_magic_23_0.VD3.n4 two_stage_opamp_dummy_magic_23_0.VD3.t13 11.2576
R7340 two_stage_opamp_dummy_magic_23_0.VD3.n4 two_stage_opamp_dummy_magic_23_0.VD3.t37 11.2576
R7341 two_stage_opamp_dummy_magic_23_0.VD3.n7 two_stage_opamp_dummy_magic_23_0.VD3.t8 11.2576
R7342 two_stage_opamp_dummy_magic_23_0.VD3.n7 two_stage_opamp_dummy_magic_23_0.VD3.t36 11.2576
R7343 two_stage_opamp_dummy_magic_23_0.VD3.n10 two_stage_opamp_dummy_magic_23_0.VD3.t12 11.2576
R7344 two_stage_opamp_dummy_magic_23_0.VD3.n10 two_stage_opamp_dummy_magic_23_0.VD3.t9 11.2576
R7345 two_stage_opamp_dummy_magic_23_0.VD3.n14 two_stage_opamp_dummy_magic_23_0.VD3.t6 11.2576
R7346 two_stage_opamp_dummy_magic_23_0.VD3.n14 two_stage_opamp_dummy_magic_23_0.VD3.t35 11.2576
R7347 two_stage_opamp_dummy_magic_23_0.VD3.n17 two_stage_opamp_dummy_magic_23_0.VD3.t10 11.2576
R7348 two_stage_opamp_dummy_magic_23_0.VD3.n17 two_stage_opamp_dummy_magic_23_0.VD3.t11 11.2576
R7349 two_stage_opamp_dummy_magic_23_0.VD3.n20 two_stage_opamp_dummy_magic_23_0.VD3.t7 11.2576
R7350 two_stage_opamp_dummy_magic_23_0.VD3.n20 two_stage_opamp_dummy_magic_23_0.VD3.t14 11.2576
R7351 two_stage_opamp_dummy_magic_23_0.VD3.t34 two_stage_opamp_dummy_magic_23_0.VD3.n35 11.2576
R7352 two_stage_opamp_dummy_magic_23_0.VD3.n35 two_stage_opamp_dummy_magic_23_0.VD3.t16 11.2576
R7353 two_stage_opamp_dummy_magic_23_0.VD3.n31 two_stage_opamp_dummy_magic_23_0.VD3.n29 6.10467
R7354 two_stage_opamp_dummy_magic_23_0.VD3.n21 two_stage_opamp_dummy_magic_23_0.VD3.n19 5.91717
R7355 two_stage_opamp_dummy_magic_23_0.VD3.n6 two_stage_opamp_dummy_magic_23_0.VD3.n5 5.91717
R7356 two_stage_opamp_dummy_magic_23_0.VD3.n9 two_stage_opamp_dummy_magic_23_0.VD3.n5 5.91717
R7357 two_stage_opamp_dummy_magic_23_0.VD3.n26 two_stage_opamp_dummy_magic_23_0.VD3.n25 5.47967
R7358 two_stage_opamp_dummy_magic_23_0.VD3.n9 two_stage_opamp_dummy_magic_23_0.VD3.n8 5.29217
R7359 two_stage_opamp_dummy_magic_23_0.VD3.n8 two_stage_opamp_dummy_magic_23_0.VD3.n6 5.29217
R7360 two_stage_opamp_dummy_magic_23_0.VD3.n12 two_stage_opamp_dummy_magic_23_0.VD3.n11 5.29217
R7361 two_stage_opamp_dummy_magic_23_0.VD3.n11 two_stage_opamp_dummy_magic_23_0.VD3.n3 5.29217
R7362 two_stage_opamp_dummy_magic_23_0.VD3.n15 two_stage_opamp_dummy_magic_23_0.VD3.n13 5.29217
R7363 two_stage_opamp_dummy_magic_23_0.VD3.n16 two_stage_opamp_dummy_magic_23_0.VD3.n15 5.29217
R7364 two_stage_opamp_dummy_magic_23_0.VD3.n18 two_stage_opamp_dummy_magic_23_0.VD3.n2 5.29217
R7365 two_stage_opamp_dummy_magic_23_0.VD3.n19 two_stage_opamp_dummy_magic_23_0.VD3.n18 5.29217
R7366 two_stage_opamp_dummy_magic_23_0.VD3.n22 two_stage_opamp_dummy_magic_23_0.VD3.n21 5.29217
R7367 two_stage_opamp_dummy_magic_23_0.VD3.n29 two_stage_opamp_dummy_magic_23_0.VD3.n28 1.03383
R7368 two_stage_opamp_dummy_magic_23_0.VD3.n27 two_stage_opamp_dummy_magic_23_0.VD3.n26 1.03383
R7369 two_stage_opamp_dummy_magic_23_0.VD3.n34 two_stage_opamp_dummy_magic_23_0.VD3.n33 0.6255
R7370 two_stage_opamp_dummy_magic_23_0.VD3.n33 two_stage_opamp_dummy_magic_23_0.VD3.n31 0.6255
R7371 two_stage_opamp_dummy_magic_23_0.VD3.n19 two_stage_opamp_dummy_magic_23_0.VD3.n16 0.6255
R7372 two_stage_opamp_dummy_magic_23_0.VD3.n16 two_stage_opamp_dummy_magic_23_0.VD3.n3 0.6255
R7373 two_stage_opamp_dummy_magic_23_0.VD3.n6 two_stage_opamp_dummy_magic_23_0.VD3.n3 0.6255
R7374 two_stage_opamp_dummy_magic_23_0.VD3.n12 two_stage_opamp_dummy_magic_23_0.VD3.n9 0.6255
R7375 two_stage_opamp_dummy_magic_23_0.VD3.n13 two_stage_opamp_dummy_magic_23_0.VD3.n12 0.6255
R7376 two_stage_opamp_dummy_magic_23_0.VD3.n13 two_stage_opamp_dummy_magic_23_0.VD3.n2 0.6255
R7377 two_stage_opamp_dummy_magic_23_0.VD3.n22 two_stage_opamp_dummy_magic_23_0.VD3.n2 0.6255
R7378 two_stage_opamp_dummy_magic_23_0.VD3.n25 two_stage_opamp_dummy_magic_23_0.VD3.n24 0.6255
R7379 two_stage_opamp_dummy_magic_23_0.VD3.n24 two_stage_opamp_dummy_magic_23_0.VD3.n1 0.6255
R7380 two_stage_opamp_dummy_magic_23_0.VD3.n34 two_stage_opamp_dummy_magic_23_0.VD3.n1 0.6255
R7381 bgr_11_0.NFET_GATE_10uA.n19 bgr_11_0.NFET_GATE_10uA.t0 384.967
R7382 bgr_11_0.NFET_GATE_10uA.n10 bgr_11_0.NFET_GATE_10uA.t20 369.534
R7383 bgr_11_0.NFET_GATE_10uA.n9 bgr_11_0.NFET_GATE_10uA.t13 369.534
R7384 bgr_11_0.NFET_GATE_10uA.n7 bgr_11_0.NFET_GATE_10uA.t17 369.534
R7385 bgr_11_0.NFET_GATE_10uA.n4 bgr_11_0.NFET_GATE_10uA.t22 369.534
R7386 bgr_11_0.NFET_GATE_10uA.n1 bgr_11_0.NFET_GATE_10uA.t21 369.534
R7387 bgr_11_0.NFET_GATE_10uA.t0 bgr_11_0.NFET_GATE_10uA.n18 369.534
R7388 bgr_11_0.NFET_GATE_10uA bgr_11_0.NFET_GATE_10uA.n20 366.553
R7389 bgr_11_0.NFET_GATE_10uA.n12 bgr_11_0.NFET_GATE_10uA.t19 192.8
R7390 bgr_11_0.NFET_GATE_10uA.n11 bgr_11_0.NFET_GATE_10uA.t6 192.8
R7391 bgr_11_0.NFET_GATE_10uA.n10 bgr_11_0.NFET_GATE_10uA.t12 192.8
R7392 bgr_11_0.NFET_GATE_10uA.n9 bgr_11_0.NFET_GATE_10uA.t11 192.8
R7393 bgr_11_0.NFET_GATE_10uA.n7 bgr_11_0.NFET_GATE_10uA.t9 192.8
R7394 bgr_11_0.NFET_GATE_10uA.n4 bgr_11_0.NFET_GATE_10uA.t8 192.8
R7395 bgr_11_0.NFET_GATE_10uA.n5 bgr_11_0.NFET_GATE_10uA.t16 192.8
R7396 bgr_11_0.NFET_GATE_10uA.n6 bgr_11_0.NFET_GATE_10uA.t23 192.8
R7397 bgr_11_0.NFET_GATE_10uA.n3 bgr_11_0.NFET_GATE_10uA.t7 192.8
R7398 bgr_11_0.NFET_GATE_10uA.n2 bgr_11_0.NFET_GATE_10uA.t15 192.8
R7399 bgr_11_0.NFET_GATE_10uA.n1 bgr_11_0.NFET_GATE_10uA.t14 192.8
R7400 bgr_11_0.NFET_GATE_10uA.n18 bgr_11_0.NFET_GATE_10uA.t5 192.8
R7401 bgr_11_0.NFET_GATE_10uA.n17 bgr_11_0.NFET_GATE_10uA.t10 192.8
R7402 bgr_11_0.NFET_GATE_10uA.n16 bgr_11_0.NFET_GATE_10uA.t18 192.8
R7403 bgr_11_0.NFET_GATE_10uA.n12 bgr_11_0.NFET_GATE_10uA.n11 176.733
R7404 bgr_11_0.NFET_GATE_10uA.n11 bgr_11_0.NFET_GATE_10uA.n10 176.733
R7405 bgr_11_0.NFET_GATE_10uA.n5 bgr_11_0.NFET_GATE_10uA.n4 176.733
R7406 bgr_11_0.NFET_GATE_10uA.n6 bgr_11_0.NFET_GATE_10uA.n5 176.733
R7407 bgr_11_0.NFET_GATE_10uA.n3 bgr_11_0.NFET_GATE_10uA.n2 176.733
R7408 bgr_11_0.NFET_GATE_10uA.n2 bgr_11_0.NFET_GATE_10uA.n1 176.733
R7409 bgr_11_0.NFET_GATE_10uA.n18 bgr_11_0.NFET_GATE_10uA.n17 176.733
R7410 bgr_11_0.NFET_GATE_10uA.n17 bgr_11_0.NFET_GATE_10uA.n16 176.733
R7411 bgr_11_0.NFET_GATE_10uA.n14 bgr_11_0.NFET_GATE_10uA.n13 169.852
R7412 bgr_11_0.NFET_GATE_10uA.n14 bgr_11_0.NFET_GATE_10uA.n8 169.852
R7413 bgr_11_0.NFET_GATE_10uA.n15 bgr_11_0.NFET_GATE_10uA.n14 166.133
R7414 bgr_11_0.NFET_GATE_10uA.n19 bgr_11_0.NFET_GATE_10uA.n0 126.877
R7415 bgr_11_0.NFET_GATE_10uA.n13 bgr_11_0.NFET_GATE_10uA.n12 56.2338
R7416 bgr_11_0.NFET_GATE_10uA.n13 bgr_11_0.NFET_GATE_10uA.n9 56.2338
R7417 bgr_11_0.NFET_GATE_10uA.n8 bgr_11_0.NFET_GATE_10uA.n7 56.2338
R7418 bgr_11_0.NFET_GATE_10uA.n8 bgr_11_0.NFET_GATE_10uA.n6 56.2338
R7419 bgr_11_0.NFET_GATE_10uA.n15 bgr_11_0.NFET_GATE_10uA.n3 56.2338
R7420 bgr_11_0.NFET_GATE_10uA.n16 bgr_11_0.NFET_GATE_10uA.n15 56.2338
R7421 bgr_11_0.NFET_GATE_10uA.n20 bgr_11_0.NFET_GATE_10uA.t2 39.4005
R7422 bgr_11_0.NFET_GATE_10uA.n20 bgr_11_0.NFET_GATE_10uA.t4 39.4005
R7423 bgr_11_0.NFET_GATE_10uA bgr_11_0.NFET_GATE_10uA.n19 30.6442
R7424 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.t3 24.0005
R7425 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.t1 24.0005
R7426 two_stage_opamp_dummy_magic_23_0.V_err_gate.n2 two_stage_opamp_dummy_magic_23_0.V_err_gate.n26 594.301
R7427 two_stage_opamp_dummy_magic_23_0.V_err_gate.n28 two_stage_opamp_dummy_magic_23_0.V_err_gate.n27 594.301
R7428 two_stage_opamp_dummy_magic_23_0.V_err_gate.n30 two_stage_opamp_dummy_magic_23_0.V_err_gate.n29 594.301
R7429 two_stage_opamp_dummy_magic_23_0.V_err_gate.n32 two_stage_opamp_dummy_magic_23_0.V_err_gate.n31 594.301
R7430 two_stage_opamp_dummy_magic_23_0.V_err_gate.n34 two_stage_opamp_dummy_magic_23_0.V_err_gate.n33 594.301
R7431 two_stage_opamp_dummy_magic_23_0.V_err_gate.n36 two_stage_opamp_dummy_magic_23_0.V_err_gate.n35 594.301
R7432 two_stage_opamp_dummy_magic_23_0.V_err_gate.n7 two_stage_opamp_dummy_magic_23_0.V_err_gate.t16 289.2
R7433 two_stage_opamp_dummy_magic_23_0.V_err_gate.n17 two_stage_opamp_dummy_magic_23_0.V_err_gate.t14 224.934
R7434 two_stage_opamp_dummy_magic_23_0.V_err_gate.n24 two_stage_opamp_dummy_magic_23_0.V_err_gate.n23 176.733
R7435 two_stage_opamp_dummy_magic_23_0.V_err_gate.n23 two_stage_opamp_dummy_magic_23_0.V_err_gate.n22 176.733
R7436 two_stage_opamp_dummy_magic_23_0.V_err_gate.n22 two_stage_opamp_dummy_magic_23_0.V_err_gate.n21 176.733
R7437 two_stage_opamp_dummy_magic_23_0.V_err_gate.n21 two_stage_opamp_dummy_magic_23_0.V_err_gate.n20 176.733
R7438 two_stage_opamp_dummy_magic_23_0.V_err_gate.n20 two_stage_opamp_dummy_magic_23_0.V_err_gate.n19 176.733
R7439 two_stage_opamp_dummy_magic_23_0.V_err_gate.n19 two_stage_opamp_dummy_magic_23_0.V_err_gate.n18 176.733
R7440 two_stage_opamp_dummy_magic_23_0.V_err_gate.n18 two_stage_opamp_dummy_magic_23_0.V_err_gate.n17 176.733
R7441 two_stage_opamp_dummy_magic_23_0.V_err_gate.n8 two_stage_opamp_dummy_magic_23_0.V_err_gate.n7 176.733
R7442 two_stage_opamp_dummy_magic_23_0.V_err_gate.n9 two_stage_opamp_dummy_magic_23_0.V_err_gate.n8 176.733
R7443 two_stage_opamp_dummy_magic_23_0.V_err_gate.n10 two_stage_opamp_dummy_magic_23_0.V_err_gate.n9 176.733
R7444 two_stage_opamp_dummy_magic_23_0.V_err_gate.n11 two_stage_opamp_dummy_magic_23_0.V_err_gate.n10 176.733
R7445 two_stage_opamp_dummy_magic_23_0.V_err_gate.n12 two_stage_opamp_dummy_magic_23_0.V_err_gate.n11 176.733
R7446 two_stage_opamp_dummy_magic_23_0.V_err_gate.n13 two_stage_opamp_dummy_magic_23_0.V_err_gate.n12 176.733
R7447 two_stage_opamp_dummy_magic_23_0.V_err_gate.n14 two_stage_opamp_dummy_magic_23_0.V_err_gate.n13 176.733
R7448 two_stage_opamp_dummy_magic_23_0.V_err_gate.n15 two_stage_opamp_dummy_magic_23_0.V_err_gate.n14 176.733
R7449 two_stage_opamp_dummy_magic_23_0.V_err_gate.n16 two_stage_opamp_dummy_magic_23_0.V_err_gate.n15 176.733
R7450 two_stage_opamp_dummy_magic_23_0.V_err_gate two_stage_opamp_dummy_magic_23_0.V_err_gate.n6 175.171
R7451 two_stage_opamp_dummy_magic_23_0.V_err_gate two_stage_opamp_dummy_magic_23_0.V_err_gate.n25 161.869
R7452 two_stage_opamp_dummy_magic_23_0.V_err_gate.n24 two_stage_opamp_dummy_magic_23_0.V_err_gate.t29 112.468
R7453 two_stage_opamp_dummy_magic_23_0.V_err_gate.n23 two_stage_opamp_dummy_magic_23_0.V_err_gate.t26 112.468
R7454 two_stage_opamp_dummy_magic_23_0.V_err_gate.n22 two_stage_opamp_dummy_magic_23_0.V_err_gate.t17 112.468
R7455 two_stage_opamp_dummy_magic_23_0.V_err_gate.n21 two_stage_opamp_dummy_magic_23_0.V_err_gate.t27 112.468
R7456 two_stage_opamp_dummy_magic_23_0.V_err_gate.n20 two_stage_opamp_dummy_magic_23_0.V_err_gate.t18 112.468
R7457 two_stage_opamp_dummy_magic_23_0.V_err_gate.n19 two_stage_opamp_dummy_magic_23_0.V_err_gate.t28 112.468
R7458 two_stage_opamp_dummy_magic_23_0.V_err_gate.n18 two_stage_opamp_dummy_magic_23_0.V_err_gate.t21 112.468
R7459 two_stage_opamp_dummy_magic_23_0.V_err_gate.n17 two_stage_opamp_dummy_magic_23_0.V_err_gate.t31 112.468
R7460 two_stage_opamp_dummy_magic_23_0.V_err_gate.n7 two_stage_opamp_dummy_magic_23_0.V_err_gate.t24 112.468
R7461 two_stage_opamp_dummy_magic_23_0.V_err_gate.n8 two_stage_opamp_dummy_magic_23_0.V_err_gate.t20 112.468
R7462 two_stage_opamp_dummy_magic_23_0.V_err_gate.n9 two_stage_opamp_dummy_magic_23_0.V_err_gate.t30 112.468
R7463 two_stage_opamp_dummy_magic_23_0.V_err_gate.n10 two_stage_opamp_dummy_magic_23_0.V_err_gate.t22 112.468
R7464 two_stage_opamp_dummy_magic_23_0.V_err_gate.n11 two_stage_opamp_dummy_magic_23_0.V_err_gate.t32 112.468
R7465 two_stage_opamp_dummy_magic_23_0.V_err_gate.n12 two_stage_opamp_dummy_magic_23_0.V_err_gate.t23 112.468
R7466 two_stage_opamp_dummy_magic_23_0.V_err_gate.n13 two_stage_opamp_dummy_magic_23_0.V_err_gate.t33 112.468
R7467 two_stage_opamp_dummy_magic_23_0.V_err_gate.n14 two_stage_opamp_dummy_magic_23_0.V_err_gate.t25 112.468
R7468 two_stage_opamp_dummy_magic_23_0.V_err_gate.n15 two_stage_opamp_dummy_magic_23_0.V_err_gate.t15 112.468
R7469 two_stage_opamp_dummy_magic_23_0.V_err_gate.n16 two_stage_opamp_dummy_magic_23_0.V_err_gate.t19 112.468
R7470 two_stage_opamp_dummy_magic_23_0.V_err_gate.n26 two_stage_opamp_dummy_magic_23_0.V_err_gate.t6 78.8005
R7471 two_stage_opamp_dummy_magic_23_0.V_err_gate.n26 two_stage_opamp_dummy_magic_23_0.V_err_gate.t10 78.8005
R7472 two_stage_opamp_dummy_magic_23_0.V_err_gate.n27 two_stage_opamp_dummy_magic_23_0.V_err_gate.t0 78.8005
R7473 two_stage_opamp_dummy_magic_23_0.V_err_gate.n27 two_stage_opamp_dummy_magic_23_0.V_err_gate.t9 78.8005
R7474 two_stage_opamp_dummy_magic_23_0.V_err_gate.n29 two_stage_opamp_dummy_magic_23_0.V_err_gate.t2 78.8005
R7475 two_stage_opamp_dummy_magic_23_0.V_err_gate.n29 two_stage_opamp_dummy_magic_23_0.V_err_gate.t1 78.8005
R7476 two_stage_opamp_dummy_magic_23_0.V_err_gate.n31 two_stage_opamp_dummy_magic_23_0.V_err_gate.t7 78.8005
R7477 two_stage_opamp_dummy_magic_23_0.V_err_gate.n31 two_stage_opamp_dummy_magic_23_0.V_err_gate.t8 78.8005
R7478 two_stage_opamp_dummy_magic_23_0.V_err_gate.n33 two_stage_opamp_dummy_magic_23_0.V_err_gate.t5 78.8005
R7479 two_stage_opamp_dummy_magic_23_0.V_err_gate.n33 two_stage_opamp_dummy_magic_23_0.V_err_gate.t12 78.8005
R7480 two_stage_opamp_dummy_magic_23_0.V_err_gate.n35 two_stage_opamp_dummy_magic_23_0.V_err_gate.t11 78.8005
R7481 two_stage_opamp_dummy_magic_23_0.V_err_gate.n35 two_stage_opamp_dummy_magic_23_0.V_err_gate.t13 78.8005
R7482 two_stage_opamp_dummy_magic_23_0.V_err_gate.n25 two_stage_opamp_dummy_magic_23_0.V_err_gate.n24 56.2338
R7483 two_stage_opamp_dummy_magic_23_0.V_err_gate.n25 two_stage_opamp_dummy_magic_23_0.V_err_gate.n16 56.2338
R7484 two_stage_opamp_dummy_magic_23_0.V_err_gate.n6 two_stage_opamp_dummy_magic_23_0.V_err_gate.t4 24.0005
R7485 two_stage_opamp_dummy_magic_23_0.V_err_gate.n6 two_stage_opamp_dummy_magic_23_0.V_err_gate.t3 24.0005
R7486 two_stage_opamp_dummy_magic_23_0.V_err_gate two_stage_opamp_dummy_magic_23_0.V_err_gate.n3 6.89112
R7487 two_stage_opamp_dummy_magic_23_0.V_err_gate.n4 two_stage_opamp_dummy_magic_23_0.V_err_gate.n2 5.41717
R7488 two_stage_opamp_dummy_magic_23_0.V_err_gate.n36 two_stage_opamp_dummy_magic_23_0.V_err_gate.n1 5.22967
R7489 two_stage_opamp_dummy_magic_23_0.V_err_gate.n0 two_stage_opamp_dummy_magic_23_0.V_err_gate.n2 5.22967
R7490 two_stage_opamp_dummy_magic_23_0.V_err_gate.n4 two_stage_opamp_dummy_magic_23_0.V_err_gate.n28 4.85467
R7491 two_stage_opamp_dummy_magic_23_0.V_err_gate.n5 two_stage_opamp_dummy_magic_23_0.V_err_gate.n30 4.85467
R7492 two_stage_opamp_dummy_magic_23_0.V_err_gate.n32 two_stage_opamp_dummy_magic_23_0.V_err_gate.n5 4.85467
R7493 two_stage_opamp_dummy_magic_23_0.V_err_gate.n34 two_stage_opamp_dummy_magic_23_0.V_err_gate.n3 4.85467
R7494 two_stage_opamp_dummy_magic_23_0.V_err_gate.n3 two_stage_opamp_dummy_magic_23_0.V_err_gate.n36 4.85467
R7495 two_stage_opamp_dummy_magic_23_0.V_err_gate.n28 two_stage_opamp_dummy_magic_23_0.V_err_gate.n0 4.66717
R7496 two_stage_opamp_dummy_magic_23_0.V_err_gate.n30 two_stage_opamp_dummy_magic_23_0.V_err_gate.n0 4.66717
R7497 two_stage_opamp_dummy_magic_23_0.V_err_gate.n1 two_stage_opamp_dummy_magic_23_0.V_err_gate.n32 4.66717
R7498 two_stage_opamp_dummy_magic_23_0.V_err_gate.n1 two_stage_opamp_dummy_magic_23_0.V_err_gate.n34 4.66717
R7499 two_stage_opamp_dummy_magic_23_0.V_err_gate.n1 two_stage_opamp_dummy_magic_23_0.V_err_gate.n0 1.688
R7500 two_stage_opamp_dummy_magic_23_0.V_err_gate.n5 two_stage_opamp_dummy_magic_23_0.V_err_gate.n3 1.1255
R7501 two_stage_opamp_dummy_magic_23_0.V_err_gate.n5 two_stage_opamp_dummy_magic_23_0.V_err_gate.n4 1.1255
R7502 two_stage_opamp_dummy_magic_23_0.cap_res_Y two_stage_opamp_dummy_magic_23_0.cap_res_Y.t0 49.2388
R7503 two_stage_opamp_dummy_magic_23_0.cap_res_Y two_stage_opamp_dummy_magic_23_0.cap_res_Y.t130 0.922875
R7504 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t89 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t52 0.1603
R7505 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t129 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t91 0.1603
R7506 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t133 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t95 0.1603
R7507 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t87 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t109 0.1603
R7508 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t132 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t131 0.1603
R7509 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t69 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t18 0.1603
R7510 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t29 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t28 0.1603
R7511 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t106 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t53 0.1603
R7512 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t136 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t134 0.1603
R7513 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t74 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t22 0.1603
R7514 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t36 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t34 0.1603
R7515 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t111 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t60 0.1603
R7516 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t73 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t72 0.1603
R7517 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t13 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t100 0.1603
R7518 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t40 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t39 0.1603
R7519 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t119 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t68 0.1603
R7520 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t78 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t77 0.1603
R7521 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t19 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t105 0.1603
R7522 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t117 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t116 0.1603
R7523 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t55 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t6 0.1603
R7524 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t84 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t83 0.1603
R7525 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t24 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t110 0.1603
R7526 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t127 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t125 0.1603
R7527 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t64 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t12 0.1603
R7528 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t23 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t21 0.1603
R7529 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t102 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t48 0.1603
R7530 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t61 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t59 0.1603
R7531 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t2 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t90 0.1603
R7532 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t30 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t27 0.1603
R7533 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t108 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t54 0.1603
R7534 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t10 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t99 0.1603
R7535 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t62 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t118 0.1603
R7536 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t11 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t14 0.1603
R7537 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t50 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t65 0.1603
R7538 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t4 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t98 0.1603
R7539 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t92 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t137 0.1603
R7540 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t32 0.1603
R7541 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t85 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t80 0.1603
R7542 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t37 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t114 0.1603
R7543 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t126 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t8 0.1603
R7544 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t25 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t58 0.1603
R7545 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t123 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t122 0.1603
R7546 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t124 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t20 0.1603
R7547 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t71 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t124 0.1603
R7548 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t33 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t71 0.1603
R7549 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t26 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t66 0.1603
R7550 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t63 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t101 0.1603
R7551 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t42 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t81 0.1603
R7552 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t79 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t120 0.1603
R7553 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t1 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t43 0.1603
R7554 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t17 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t1 0.1603
R7555 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t115 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t17 0.1603
R7556 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t38 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t76 0.1603
R7557 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t51 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t38 0.1603
R7558 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t51 0.1603
R7559 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t35 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t135 0.1603
R7560 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t88 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t35 0.1603
R7561 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t130 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t88 0.1603
R7562 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t121 0.159278
R7563 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t112 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n15 0.159278
R7564 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t5 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n16 0.159278
R7565 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t41 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n17 0.159278
R7566 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n18 0.159278
R7567 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t97 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n19 0.159278
R7568 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t56 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n20 0.159278
R7569 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t93 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n21 0.159278
R7570 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t49 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n22 0.159278
R7571 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t15 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n23 0.159278
R7572 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t46 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n24 0.159278
R7573 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t7 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n25 0.159278
R7574 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t107 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n26 0.159278
R7575 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t3 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n27 0.159278
R7576 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t103 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n28 0.159278
R7577 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t128 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n29 0.159278
R7578 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t86 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n30 0.159278
R7579 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t82 0.159278
R7580 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t104 0.159278
R7581 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t67 0.159278
R7582 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t57 0.159278
R7583 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t96 0.159278
R7584 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t75 0.159278
R7585 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t113 0.159278
R7586 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t9 0.159278
R7587 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t47 0.159278
R7588 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t31 0.159278
R7589 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t121 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t129 0.137822
R7590 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t89 0.1368
R7591 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t133 0.1368
R7592 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t87 0.1368
R7593 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t132 0.1368
R7594 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t69 0.1368
R7595 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t29 0.1368
R7596 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t106 0.1368
R7597 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t136 0.1368
R7598 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t74 0.1368
R7599 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t36 0.1368
R7600 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t111 0.1368
R7601 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t73 0.1368
R7602 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t13 0.1368
R7603 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t40 0.1368
R7604 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t119 0.1368
R7605 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t78 0.1368
R7606 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t19 0.1368
R7607 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t117 0.1368
R7608 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t55 0.1368
R7609 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t84 0.1368
R7610 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t24 0.1368
R7611 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t127 0.1368
R7612 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t64 0.1368
R7613 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t23 0.1368
R7614 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t102 0.1368
R7615 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t61 0.1368
R7616 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t2 0.1368
R7617 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t30 0.1368
R7618 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t108 0.1368
R7619 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t10 0.1368
R7620 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t123 0.1368
R7621 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t62 0.114322
R7622 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n6 0.1133
R7623 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n7 0.1133
R7624 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n8 0.1133
R7625 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n9 0.1133
R7626 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n10 0.1133
R7627 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n11 0.1133
R7628 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n12 0.1133
R7629 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n13 0.1133
R7630 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n14 0.1133
R7631 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n31 0.1133
R7632 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n32 0.1133
R7633 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n33 0.1133
R7634 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n0 0.1133
R7635 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n1 0.1133
R7636 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n2 0.1133
R7637 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n3 0.1133
R7638 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n4 0.1133
R7639 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n5 0.1133
R7640 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n34 0.1133
R7641 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t11 0.00152174
R7642 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t50 0.00152174
R7643 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t4 0.00152174
R7644 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t92 0.00152174
R7645 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t44 0.00152174
R7646 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t85 0.00152174
R7647 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t37 0.00152174
R7648 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t126 0.00152174
R7649 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t25 0.00152174
R7650 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t94 0.00152174
R7651 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t112 0.00152174
R7652 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t5 0.00152174
R7653 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t41 0.00152174
R7654 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t138 0.00152174
R7655 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t97 0.00152174
R7656 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t56 0.00152174
R7657 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t93 0.00152174
R7658 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t49 0.00152174
R7659 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t15 0.00152174
R7660 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t46 0.00152174
R7661 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t7 0.00152174
R7662 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t107 0.00152174
R7663 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t3 0.00152174
R7664 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t103 0.00152174
R7665 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t128 0.00152174
R7666 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t86 0.00152174
R7667 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t45 0.00152174
R7668 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t70 0.00152174
R7669 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t33 0.00152174
R7670 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t26 0.00152174
R7671 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t63 0.00152174
R7672 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t42 0.00152174
R7673 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t79 0.00152174
R7674 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t115 0.00152174
R7675 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t16 0.00152174
R7676 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t135 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n35 0.00152174
R7677 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.t32 354.854
R7678 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.t17 346.8
R7679 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.n11 339.522
R7680 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.n4 339.522
R7681 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.n9 335.022
R7682 bgr_11_0.1st_Vout_1.n7 bgr_11_0.1st_Vout_1.t4 275.909
R7683 bgr_11_0.1st_Vout_1.n7 bgr_11_0.1st_Vout_1.n6 227.909
R7684 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.n8 222.034
R7685 bgr_11_0.1st_Vout_1.n10 bgr_11_0.1st_Vout_1.t18 184.097
R7686 bgr_11_0.1st_Vout_1.n10 bgr_11_0.1st_Vout_1.t31 184.097
R7687 bgr_11_0.1st_Vout_1.n5 bgr_11_0.1st_Vout_1.t14 184.097
R7688 bgr_11_0.1st_Vout_1.n5 bgr_11_0.1st_Vout_1.t35 184.097
R7689 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.n10 166.05
R7690 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.n5 166.05
R7691 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.n3 54.2759
R7692 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.t10 48.0005
R7693 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.t8 48.0005
R7694 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.t2 48.0005
R7695 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.t3 48.0005
R7696 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.t9 39.4005
R7697 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.t6 39.4005
R7698 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.t7 39.4005
R7699 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.t1 39.4005
R7700 bgr_11_0.1st_Vout_1.n11 bgr_11_0.1st_Vout_1.t0 39.4005
R7701 bgr_11_0.1st_Vout_1.n11 bgr_11_0.1st_Vout_1.t5 39.4005
R7702 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.n0 5.6255
R7703 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.n2 5.28175
R7704 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t11 4.8295
R7705 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t26 4.8295
R7706 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t29 4.8295
R7707 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t19 4.8295
R7708 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t36 4.8295
R7709 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t24 4.8295
R7710 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t27 4.8295
R7711 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t16 4.8295
R7712 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t20 4.8295
R7713 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.n7 4.5005
R7714 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t30 4.5005
R7715 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t34 4.5005
R7716 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t22 4.5005
R7717 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t25 4.5005
R7718 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t28 4.5005
R7719 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t33 4.5005
R7720 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t21 4.5005
R7721 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t23 4.5005
R7722 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t13 4.5005
R7723 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t15 4.5005
R7724 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t12 4.5005
R7725 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.n1 3.1025
R7726 bgr_11_0.cap_res1.t0 bgr_11_0.cap_res1.t18 121.245
R7727 bgr_11_0.cap_res1.t17 bgr_11_0.cap_res1.t19 0.1603
R7728 bgr_11_0.cap_res1.t11 bgr_11_0.cap_res1.t16 0.1603
R7729 bgr_11_0.cap_res1.t3 bgr_11_0.cap_res1.t10 0.1603
R7730 bgr_11_0.cap_res1.t9 bgr_11_0.cap_res1.t15 0.1603
R7731 bgr_11_0.cap_res1.t2 bgr_11_0.cap_res1.t8 0.1603
R7732 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t4 0.159278
R7733 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t12 0.159278
R7734 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t6 0.159278
R7735 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t13 0.159278
R7736 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t17 0.1368
R7737 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t14 0.1368
R7738 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t11 0.1368
R7739 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t7 0.1368
R7740 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t3 0.1368
R7741 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t1 0.1368
R7742 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t9 0.1368
R7743 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t5 0.1368
R7744 bgr_11_0.cap_res1.n0 bgr_11_0.cap_res1.t2 0.1368
R7745 bgr_11_0.cap_res1.n0 bgr_11_0.cap_res1.t20 0.1368
R7746 bgr_11_0.cap_res1.t4 bgr_11_0.cap_res1.n0 0.00152174
R7747 bgr_11_0.cap_res1.t12 bgr_11_0.cap_res1.n1 0.00152174
R7748 bgr_11_0.cap_res1.t6 bgr_11_0.cap_res1.n2 0.00152174
R7749 bgr_11_0.cap_res1.t13 bgr_11_0.cap_res1.n3 0.00152174
R7750 bgr_11_0.cap_res1.t18 bgr_11_0.cap_res1.n4 0.00152174
R7751 two_stage_opamp_dummy_magic_23_0.VD2.n4 two_stage_opamp_dummy_magic_23_0.VD2.n3 49.3505
R7752 two_stage_opamp_dummy_magic_23_0.VD2.n13 two_stage_opamp_dummy_magic_23_0.VD2.n12 49.3505
R7753 two_stage_opamp_dummy_magic_23_0.VD2.n1 two_stage_opamp_dummy_magic_23_0.VD2.n0 49.3505
R7754 two_stage_opamp_dummy_magic_23_0.VD2.n20 two_stage_opamp_dummy_magic_23_0.VD2.n19 49.3505
R7755 two_stage_opamp_dummy_magic_23_0.VD2.n23 two_stage_opamp_dummy_magic_23_0.VD2.n22 49.3505
R7756 two_stage_opamp_dummy_magic_23_0.VD2.n26 two_stage_opamp_dummy_magic_23_0.VD2.n25 49.3505
R7757 two_stage_opamp_dummy_magic_23_0.VD2.n29 two_stage_opamp_dummy_magic_23_0.VD2.n28 49.3505
R7758 two_stage_opamp_dummy_magic_23_0.VD2.n31 two_stage_opamp_dummy_magic_23_0.VD2.n30 49.3505
R7759 two_stage_opamp_dummy_magic_23_0.VD2.n35 two_stage_opamp_dummy_magic_23_0.VD2.n34 49.3505
R7760 two_stage_opamp_dummy_magic_23_0.VD2.n8 two_stage_opamp_dummy_magic_23_0.VD2.n7 49.3505
R7761 two_stage_opamp_dummy_magic_23_0.VD2.n6 two_stage_opamp_dummy_magic_23_0.VD2.n5 49.3505
R7762 two_stage_opamp_dummy_magic_23_0.VD2.n3 two_stage_opamp_dummy_magic_23_0.VD2.t16 16.0005
R7763 two_stage_opamp_dummy_magic_23_0.VD2.n3 two_stage_opamp_dummy_magic_23_0.VD2.t12 16.0005
R7764 two_stage_opamp_dummy_magic_23_0.VD2.n12 two_stage_opamp_dummy_magic_23_0.VD2.t17 16.0005
R7765 two_stage_opamp_dummy_magic_23_0.VD2.n12 two_stage_opamp_dummy_magic_23_0.VD2.t13 16.0005
R7766 two_stage_opamp_dummy_magic_23_0.VD2.n0 two_stage_opamp_dummy_magic_23_0.VD2.t19 16.0005
R7767 two_stage_opamp_dummy_magic_23_0.VD2.n0 two_stage_opamp_dummy_magic_23_0.VD2.t14 16.0005
R7768 two_stage_opamp_dummy_magic_23_0.VD2.n19 two_stage_opamp_dummy_magic_23_0.VD2.t8 16.0005
R7769 two_stage_opamp_dummy_magic_23_0.VD2.n19 two_stage_opamp_dummy_magic_23_0.VD2.t4 16.0005
R7770 two_stage_opamp_dummy_magic_23_0.VD2.n22 two_stage_opamp_dummy_magic_23_0.VD2.t3 16.0005
R7771 two_stage_opamp_dummy_magic_23_0.VD2.n22 two_stage_opamp_dummy_magic_23_0.VD2.t5 16.0005
R7772 two_stage_opamp_dummy_magic_23_0.VD2.n25 two_stage_opamp_dummy_magic_23_0.VD2.t0 16.0005
R7773 two_stage_opamp_dummy_magic_23_0.VD2.n25 two_stage_opamp_dummy_magic_23_0.VD2.t6 16.0005
R7774 two_stage_opamp_dummy_magic_23_0.VD2.n28 two_stage_opamp_dummy_magic_23_0.VD2.t1 16.0005
R7775 two_stage_opamp_dummy_magic_23_0.VD2.n28 two_stage_opamp_dummy_magic_23_0.VD2.t9 16.0005
R7776 two_stage_opamp_dummy_magic_23_0.VD2.n30 two_stage_opamp_dummy_magic_23_0.VD2.t11 16.0005
R7777 two_stage_opamp_dummy_magic_23_0.VD2.n30 two_stage_opamp_dummy_magic_23_0.VD2.t7 16.0005
R7778 two_stage_opamp_dummy_magic_23_0.VD2.n34 two_stage_opamp_dummy_magic_23_0.VD2.t2 16.0005
R7779 two_stage_opamp_dummy_magic_23_0.VD2.n34 two_stage_opamp_dummy_magic_23_0.VD2.t10 16.0005
R7780 two_stage_opamp_dummy_magic_23_0.VD2.n7 two_stage_opamp_dummy_magic_23_0.VD2.t18 16.0005
R7781 two_stage_opamp_dummy_magic_23_0.VD2.n7 two_stage_opamp_dummy_magic_23_0.VD2.t21 16.0005
R7782 two_stage_opamp_dummy_magic_23_0.VD2.n5 two_stage_opamp_dummy_magic_23_0.VD2.t20 16.0005
R7783 two_stage_opamp_dummy_magic_23_0.VD2.n5 two_stage_opamp_dummy_magic_23_0.VD2.t15 16.0005
R7784 two_stage_opamp_dummy_magic_23_0.VD2.n29 two_stage_opamp_dummy_magic_23_0.VD2.n18 5.64633
R7785 two_stage_opamp_dummy_magic_23_0.VD2.n21 two_stage_opamp_dummy_magic_23_0.VD2.n20 5.64633
R7786 two_stage_opamp_dummy_magic_23_0.VD2.n9 two_stage_opamp_dummy_magic_23_0.VD2.n6 5.6255
R7787 two_stage_opamp_dummy_magic_23_0.VD2.n11 two_stage_opamp_dummy_magic_23_0.VD2.n4 5.6255
R7788 two_stage_opamp_dummy_magic_23_0.VD2.n32 two_stage_opamp_dummy_magic_23_0.VD2.n29 5.438
R7789 two_stage_opamp_dummy_magic_23_0.VD2.n24 two_stage_opamp_dummy_magic_23_0.VD2.n20 5.438
R7790 two_stage_opamp_dummy_magic_23_0.VD2.n14 two_stage_opamp_dummy_magic_23_0.VD2.n4 5.438
R7791 two_stage_opamp_dummy_magic_23_0.VD2.n6 two_stage_opamp_dummy_magic_23_0.VD2.n2 5.438
R7792 two_stage_opamp_dummy_magic_23_0.VD2.n23 two_stage_opamp_dummy_magic_23_0.VD2.n21 5.08383
R7793 two_stage_opamp_dummy_magic_23_0.VD2.n26 two_stage_opamp_dummy_magic_23_0.VD2.n17 5.08383
R7794 two_stage_opamp_dummy_magic_23_0.VD2.n31 two_stage_opamp_dummy_magic_23_0.VD2.n18 5.08383
R7795 two_stage_opamp_dummy_magic_23_0.VD2.n36 two_stage_opamp_dummy_magic_23_0.VD2.n35 5.08383
R7796 two_stage_opamp_dummy_magic_23_0.VD2.n13 two_stage_opamp_dummy_magic_23_0.VD2.n11 5.063
R7797 two_stage_opamp_dummy_magic_23_0.VD2.n10 two_stage_opamp_dummy_magic_23_0.VD2.n1 5.063
R7798 two_stage_opamp_dummy_magic_23_0.VD2.n9 two_stage_opamp_dummy_magic_23_0.VD2.n8 5.063
R7799 two_stage_opamp_dummy_magic_23_0.VD2 two_stage_opamp_dummy_magic_23_0.VD2.n37 5.02133
R7800 two_stage_opamp_dummy_magic_23_0.VD2.n14 two_stage_opamp_dummy_magic_23_0.VD2.n13 4.8755
R7801 two_stage_opamp_dummy_magic_23_0.VD2.n24 two_stage_opamp_dummy_magic_23_0.VD2.n23 4.8755
R7802 two_stage_opamp_dummy_magic_23_0.VD2.n27 two_stage_opamp_dummy_magic_23_0.VD2.n26 4.8755
R7803 two_stage_opamp_dummy_magic_23_0.VD2.n32 two_stage_opamp_dummy_magic_23_0.VD2.n31 4.8755
R7804 two_stage_opamp_dummy_magic_23_0.VD2.n35 two_stage_opamp_dummy_magic_23_0.VD2.n33 4.8755
R7805 two_stage_opamp_dummy_magic_23_0.VD2.n8 two_stage_opamp_dummy_magic_23_0.VD2.n2 4.8755
R7806 two_stage_opamp_dummy_magic_23_0.VD2.n16 two_stage_opamp_dummy_magic_23_0.VD2.n15 4.5005
R7807 two_stage_opamp_dummy_magic_23_0.VD2 two_stage_opamp_dummy_magic_23_0.VD2.n16 0.7505
R7808 two_stage_opamp_dummy_magic_23_0.VD2.n36 two_stage_opamp_dummy_magic_23_0.VD2.n18 0.563
R7809 two_stage_opamp_dummy_magic_23_0.VD2.n33 two_stage_opamp_dummy_magic_23_0.VD2.n32 0.563
R7810 two_stage_opamp_dummy_magic_23_0.VD2.n33 two_stage_opamp_dummy_magic_23_0.VD2.n27 0.563
R7811 two_stage_opamp_dummy_magic_23_0.VD2.n27 two_stage_opamp_dummy_magic_23_0.VD2.n24 0.563
R7812 two_stage_opamp_dummy_magic_23_0.VD2.n21 two_stage_opamp_dummy_magic_23_0.VD2.n17 0.563
R7813 two_stage_opamp_dummy_magic_23_0.VD2.n10 two_stage_opamp_dummy_magic_23_0.VD2.n9 0.563
R7814 two_stage_opamp_dummy_magic_23_0.VD2.n11 two_stage_opamp_dummy_magic_23_0.VD2.n10 0.563
R7815 two_stage_opamp_dummy_magic_23_0.VD2.n15 two_stage_opamp_dummy_magic_23_0.VD2.n14 0.563
R7816 two_stage_opamp_dummy_magic_23_0.VD2.n15 two_stage_opamp_dummy_magic_23_0.VD2.n2 0.563
R7817 two_stage_opamp_dummy_magic_23_0.VD2.n16 two_stage_opamp_dummy_magic_23_0.VD2.n1 0.3755
R7818 two_stage_opamp_dummy_magic_23_0.VD2.n37 two_stage_opamp_dummy_magic_23_0.VD2.n36 0.234875
R7819 two_stage_opamp_dummy_magic_23_0.VD2.n37 two_stage_opamp_dummy_magic_23_0.VD2.n17 0.234875
R7820 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t21 610.534
R7821 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t19 610.534
R7822 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t30 433.8
R7823 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t27 433.8
R7824 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t16 433.8
R7825 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t24 433.8
R7826 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t13 433.8
R7827 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t23 433.8
R7828 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t12 433.8
R7829 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t22 433.8
R7830 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t25 433.8
R7831 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t14 433.8
R7832 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t31 433.8
R7833 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t20 433.8
R7834 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t29 433.8
R7835 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t18 433.8
R7836 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t28 433.8
R7837 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t17 433.8
R7838 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t26 433.8
R7839 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t15 433.8
R7840 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n0 339.836
R7841 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n1 339.834
R7842 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n2 339.272
R7843 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n5 287.264
R7844 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n24 176.733
R7845 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n23 176.733
R7846 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n22 176.733
R7847 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n21 176.733
R7848 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n20 176.733
R7849 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n19 176.733
R7850 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n18 176.733
R7851 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n17 176.733
R7852 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n8 176.733
R7853 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n9 176.733
R7854 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n10 176.733
R7855 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n11 176.733
R7856 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n12 176.733
R7857 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n13 176.733
R7858 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n14 176.733
R7859 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n15 176.733
R7860 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n26 162.508
R7861 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n25 56.2338
R7862 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n16 56.2338
R7863 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n4 52.01
R7864 two_stage_opamp_dummy_magic_23_0.V_tail_gate two_stage_opamp_dummy_magic_23_0.V_tail_gate.n6 51.6642
R7865 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n7 50.5797
R7866 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n28 49.3505
R7867 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t3 39.4005
R7868 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t9 39.4005
R7869 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t11 39.4005
R7870 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t10 39.4005
R7871 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t2 39.4005
R7872 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t4 39.4005
R7873 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t1 39.4005
R7874 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t5 39.4005
R7875 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t6 16.0005
R7876 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t7 16.0005
R7877 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t8 16.0005
R7878 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t0 16.0005
R7879 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n27 10.7922
R7880 two_stage_opamp_dummy_magic_23_0.V_tail_gate two_stage_opamp_dummy_magic_23_0.V_tail_gate.n29 1.04217
R7881 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n3 0.563
R7882 two_stage_opamp_dummy_magic_23_0.V_source.n48 two_stage_opamp_dummy_magic_23_0.V_source.t40 66.2047
R7883 two_stage_opamp_dummy_magic_23_0.V_source.n5 two_stage_opamp_dummy_magic_23_0.V_source.n4 49.3505
R7884 two_stage_opamp_dummy_magic_23_0.V_source.n8 two_stage_opamp_dummy_magic_23_0.V_source.n7 49.3505
R7885 two_stage_opamp_dummy_magic_23_0.V_source.n11 two_stage_opamp_dummy_magic_23_0.V_source.n10 49.3505
R7886 two_stage_opamp_dummy_magic_23_0.V_source.n14 two_stage_opamp_dummy_magic_23_0.V_source.n13 49.3505
R7887 two_stage_opamp_dummy_magic_23_0.V_source.n18 two_stage_opamp_dummy_magic_23_0.V_source.n17 49.3505
R7888 two_stage_opamp_dummy_magic_23_0.V_source.n23 two_stage_opamp_dummy_magic_23_0.V_source.n22 49.3505
R7889 two_stage_opamp_dummy_magic_23_0.V_source.n25 two_stage_opamp_dummy_magic_23_0.V_source.n24 49.3505
R7890 two_stage_opamp_dummy_magic_23_0.V_source.n29 two_stage_opamp_dummy_magic_23_0.V_source.n28 49.3505
R7891 two_stage_opamp_dummy_magic_23_0.V_source.n32 two_stage_opamp_dummy_magic_23_0.V_source.n31 49.3505
R7892 two_stage_opamp_dummy_magic_23_0.V_source.n35 two_stage_opamp_dummy_magic_23_0.V_source.n34 49.3505
R7893 two_stage_opamp_dummy_magic_23_0.V_source.n40 two_stage_opamp_dummy_magic_23_0.V_source.n39 32.3838
R7894 two_stage_opamp_dummy_magic_23_0.V_source.n42 two_stage_opamp_dummy_magic_23_0.V_source.n41 32.3838
R7895 two_stage_opamp_dummy_magic_23_0.V_source.n47 two_stage_opamp_dummy_magic_23_0.V_source.n46 32.3838
R7896 two_stage_opamp_dummy_magic_23_0.V_source.n51 two_stage_opamp_dummy_magic_23_0.V_source.n50 32.3838
R7897 two_stage_opamp_dummy_magic_23_0.V_source.n55 two_stage_opamp_dummy_magic_23_0.V_source.n54 32.3838
R7898 two_stage_opamp_dummy_magic_23_0.V_source.n58 two_stage_opamp_dummy_magic_23_0.V_source.n57 32.3838
R7899 two_stage_opamp_dummy_magic_23_0.V_source.n62 two_stage_opamp_dummy_magic_23_0.V_source.n61 32.3838
R7900 two_stage_opamp_dummy_magic_23_0.V_source.n65 two_stage_opamp_dummy_magic_23_0.V_source.n64 32.3838
R7901 two_stage_opamp_dummy_magic_23_0.V_source.n68 two_stage_opamp_dummy_magic_23_0.V_source.n67 32.3838
R7902 two_stage_opamp_dummy_magic_23_0.V_source.n72 two_stage_opamp_dummy_magic_23_0.V_source.n71 32.3838
R7903 two_stage_opamp_dummy_magic_23_0.V_source.n4 two_stage_opamp_dummy_magic_23_0.V_source.t37 16.0005
R7904 two_stage_opamp_dummy_magic_23_0.V_source.n4 two_stage_opamp_dummy_magic_23_0.V_source.t26 16.0005
R7905 two_stage_opamp_dummy_magic_23_0.V_source.n7 two_stage_opamp_dummy_magic_23_0.V_source.t31 16.0005
R7906 two_stage_opamp_dummy_magic_23_0.V_source.n7 two_stage_opamp_dummy_magic_23_0.V_source.t6 16.0005
R7907 two_stage_opamp_dummy_magic_23_0.V_source.n10 two_stage_opamp_dummy_magic_23_0.V_source.t34 16.0005
R7908 two_stage_opamp_dummy_magic_23_0.V_source.n10 two_stage_opamp_dummy_magic_23_0.V_source.t32 16.0005
R7909 two_stage_opamp_dummy_magic_23_0.V_source.n13 two_stage_opamp_dummy_magic_23_0.V_source.t5 16.0005
R7910 two_stage_opamp_dummy_magic_23_0.V_source.n13 two_stage_opamp_dummy_magic_23_0.V_source.t7 16.0005
R7911 two_stage_opamp_dummy_magic_23_0.V_source.n17 two_stage_opamp_dummy_magic_23_0.V_source.t0 16.0005
R7912 two_stage_opamp_dummy_magic_23_0.V_source.n17 two_stage_opamp_dummy_magic_23_0.V_source.t28 16.0005
R7913 two_stage_opamp_dummy_magic_23_0.V_source.n22 two_stage_opamp_dummy_magic_23_0.V_source.t35 16.0005
R7914 two_stage_opamp_dummy_magic_23_0.V_source.n22 two_stage_opamp_dummy_magic_23_0.V_source.t3 16.0005
R7915 two_stage_opamp_dummy_magic_23_0.V_source.n24 two_stage_opamp_dummy_magic_23_0.V_source.t38 16.0005
R7916 two_stage_opamp_dummy_magic_23_0.V_source.n24 two_stage_opamp_dummy_magic_23_0.V_source.t39 16.0005
R7917 two_stage_opamp_dummy_magic_23_0.V_source.n28 two_stage_opamp_dummy_magic_23_0.V_source.t33 16.0005
R7918 two_stage_opamp_dummy_magic_23_0.V_source.n28 two_stage_opamp_dummy_magic_23_0.V_source.t4 16.0005
R7919 two_stage_opamp_dummy_magic_23_0.V_source.n31 two_stage_opamp_dummy_magic_23_0.V_source.t30 16.0005
R7920 two_stage_opamp_dummy_magic_23_0.V_source.n31 two_stage_opamp_dummy_magic_23_0.V_source.t1 16.0005
R7921 two_stage_opamp_dummy_magic_23_0.V_source.n34 two_stage_opamp_dummy_magic_23_0.V_source.t29 16.0005
R7922 two_stage_opamp_dummy_magic_23_0.V_source.n34 two_stage_opamp_dummy_magic_23_0.V_source.t27 16.0005
R7923 two_stage_opamp_dummy_magic_23_0.V_source.n39 two_stage_opamp_dummy_magic_23_0.V_source.t36 9.6005
R7924 two_stage_opamp_dummy_magic_23_0.V_source.n39 two_stage_opamp_dummy_magic_23_0.V_source.t2 9.6005
R7925 two_stage_opamp_dummy_magic_23_0.V_source.n41 two_stage_opamp_dummy_magic_23_0.V_source.t18 9.6005
R7926 two_stage_opamp_dummy_magic_23_0.V_source.n41 two_stage_opamp_dummy_magic_23_0.V_source.t22 9.6005
R7927 two_stage_opamp_dummy_magic_23_0.V_source.n46 two_stage_opamp_dummy_magic_23_0.V_source.t12 9.6005
R7928 two_stage_opamp_dummy_magic_23_0.V_source.n46 two_stage_opamp_dummy_magic_23_0.V_source.t20 9.6005
R7929 two_stage_opamp_dummy_magic_23_0.V_source.n50 two_stage_opamp_dummy_magic_23_0.V_source.t10 9.6005
R7930 two_stage_opamp_dummy_magic_23_0.V_source.n50 two_stage_opamp_dummy_magic_23_0.V_source.t19 9.6005
R7931 two_stage_opamp_dummy_magic_23_0.V_source.n54 two_stage_opamp_dummy_magic_23_0.V_source.t9 9.6005
R7932 two_stage_opamp_dummy_magic_23_0.V_source.n54 two_stage_opamp_dummy_magic_23_0.V_source.t17 9.6005
R7933 two_stage_opamp_dummy_magic_23_0.V_source.n57 two_stage_opamp_dummy_magic_23_0.V_source.t8 9.6005
R7934 two_stage_opamp_dummy_magic_23_0.V_source.n57 two_stage_opamp_dummy_magic_23_0.V_source.t23 9.6005
R7935 two_stage_opamp_dummy_magic_23_0.V_source.n61 two_stage_opamp_dummy_magic_23_0.V_source.t13 9.6005
R7936 two_stage_opamp_dummy_magic_23_0.V_source.n61 two_stage_opamp_dummy_magic_23_0.V_source.t16 9.6005
R7937 two_stage_opamp_dummy_magic_23_0.V_source.n64 two_stage_opamp_dummy_magic_23_0.V_source.t21 9.6005
R7938 two_stage_opamp_dummy_magic_23_0.V_source.n64 two_stage_opamp_dummy_magic_23_0.V_source.t11 9.6005
R7939 two_stage_opamp_dummy_magic_23_0.V_source.n67 two_stage_opamp_dummy_magic_23_0.V_source.t24 9.6005
R7940 two_stage_opamp_dummy_magic_23_0.V_source.n67 two_stage_opamp_dummy_magic_23_0.V_source.t14 9.6005
R7941 two_stage_opamp_dummy_magic_23_0.V_source.t25 two_stage_opamp_dummy_magic_23_0.V_source.n72 9.6005
R7942 two_stage_opamp_dummy_magic_23_0.V_source.n72 two_stage_opamp_dummy_magic_23_0.V_source.t15 9.6005
R7943 two_stage_opamp_dummy_magic_23_0.V_source.n69 two_stage_opamp_dummy_magic_23_0.V_source.n65 5.89633
R7944 two_stage_opamp_dummy_magic_23_0.V_source.n40 two_stage_opamp_dummy_magic_23_0.V_source.n3 5.89633
R7945 two_stage_opamp_dummy_magic_23_0.V_source.n66 two_stage_opamp_dummy_magic_23_0.V_source.n65 5.70883
R7946 two_stage_opamp_dummy_magic_23_0.V_source.n43 two_stage_opamp_dummy_magic_23_0.V_source.n40 5.70883
R7947 two_stage_opamp_dummy_magic_23_0.V_source.n26 two_stage_opamp_dummy_magic_23_0.V_source.n23 5.6255
R7948 two_stage_opamp_dummy_magic_23_0.V_source.n9 two_stage_opamp_dummy_magic_23_0.V_source.n8 5.6255
R7949 two_stage_opamp_dummy_magic_23_0.V_source.n35 two_stage_opamp_dummy_magic_23_0.V_source.n33 5.45883
R7950 two_stage_opamp_dummy_magic_23_0.V_source.n23 two_stage_opamp_dummy_magic_23_0.V_source.n21 5.45883
R7951 two_stage_opamp_dummy_magic_23_0.V_source.n12 two_stage_opamp_dummy_magic_23_0.V_source.n8 5.45883
R7952 two_stage_opamp_dummy_magic_23_0.V_source.n16 two_stage_opamp_dummy_magic_23_0.V_source.n5 5.45883
R7953 two_stage_opamp_dummy_magic_23_0.V_source.n42 two_stage_opamp_dummy_magic_23_0.V_source.n3 5.33383
R7954 two_stage_opamp_dummy_magic_23_0.V_source.n52 two_stage_opamp_dummy_magic_23_0.V_source.n51 5.33383
R7955 two_stage_opamp_dummy_magic_23_0.V_source.n55 two_stage_opamp_dummy_magic_23_0.V_source.n53 5.33383
R7956 two_stage_opamp_dummy_magic_23_0.V_source.n58 two_stage_opamp_dummy_magic_23_0.V_source.n1 5.33383
R7957 two_stage_opamp_dummy_magic_23_0.V_source.n63 two_stage_opamp_dummy_magic_23_0.V_source.n62 5.33383
R7958 two_stage_opamp_dummy_magic_23_0.V_source.n69 two_stage_opamp_dummy_magic_23_0.V_source.n68 5.33383
R7959 two_stage_opamp_dummy_magic_23_0.V_source.n71 two_stage_opamp_dummy_magic_23_0.V_source.n70 5.33383
R7960 two_stage_opamp_dummy_magic_23_0.V_source.n43 two_stage_opamp_dummy_magic_23_0.V_source.n42 5.14633
R7961 two_stage_opamp_dummy_magic_23_0.V_source.n51 two_stage_opamp_dummy_magic_23_0.V_source.n2 5.14633
R7962 two_stage_opamp_dummy_magic_23_0.V_source.n56 two_stage_opamp_dummy_magic_23_0.V_source.n55 5.14633
R7963 two_stage_opamp_dummy_magic_23_0.V_source.n59 two_stage_opamp_dummy_magic_23_0.V_source.n58 5.14633
R7964 two_stage_opamp_dummy_magic_23_0.V_source.n62 two_stage_opamp_dummy_magic_23_0.V_source.n60 5.14633
R7965 two_stage_opamp_dummy_magic_23_0.V_source.n71 two_stage_opamp_dummy_magic_23_0.V_source.n0 5.14633
R7966 two_stage_opamp_dummy_magic_23_0.V_source.n68 two_stage_opamp_dummy_magic_23_0.V_source.n66 5.14633
R7967 two_stage_opamp_dummy_magic_23_0.V_source.n11 two_stage_opamp_dummy_magic_23_0.V_source.n9 5.063
R7968 two_stage_opamp_dummy_magic_23_0.V_source.n14 two_stage_opamp_dummy_magic_23_0.V_source.n6 5.063
R7969 two_stage_opamp_dummy_magic_23_0.V_source.n19 two_stage_opamp_dummy_magic_23_0.V_source.n18 5.063
R7970 two_stage_opamp_dummy_magic_23_0.V_source.n26 two_stage_opamp_dummy_magic_23_0.V_source.n25 5.063
R7971 two_stage_opamp_dummy_magic_23_0.V_source.n29 two_stage_opamp_dummy_magic_23_0.V_source.n27 5.063
R7972 two_stage_opamp_dummy_magic_23_0.V_source.n32 two_stage_opamp_dummy_magic_23_0.V_source.n20 5.063
R7973 two_stage_opamp_dummy_magic_23_0.V_source.n36 two_stage_opamp_dummy_magic_23_0.V_source.n35 5.063
R7974 two_stage_opamp_dummy_magic_23_0.V_source.n12 two_stage_opamp_dummy_magic_23_0.V_source.n11 4.89633
R7975 two_stage_opamp_dummy_magic_23_0.V_source.n15 two_stage_opamp_dummy_magic_23_0.V_source.n14 4.89633
R7976 two_stage_opamp_dummy_magic_23_0.V_source.n18 two_stage_opamp_dummy_magic_23_0.V_source.n16 4.89633
R7977 two_stage_opamp_dummy_magic_23_0.V_source.n25 two_stage_opamp_dummy_magic_23_0.V_source.n21 4.89633
R7978 two_stage_opamp_dummy_magic_23_0.V_source.n30 two_stage_opamp_dummy_magic_23_0.V_source.n29 4.89633
R7979 two_stage_opamp_dummy_magic_23_0.V_source.n33 two_stage_opamp_dummy_magic_23_0.V_source.n32 4.89633
R7980 two_stage_opamp_dummy_magic_23_0.V_source.n38 two_stage_opamp_dummy_magic_23_0.V_source.n37 4.5005
R7981 two_stage_opamp_dummy_magic_23_0.V_source.n45 two_stage_opamp_dummy_magic_23_0.V_source.n44 4.5005
R7982 two_stage_opamp_dummy_magic_23_0.V_source.n49 two_stage_opamp_dummy_magic_23_0.V_source.n48 4.5005
R7983 two_stage_opamp_dummy_magic_23_0.V_source.n37 two_stage_opamp_dummy_magic_23_0.V_source.n36 3.6255
R7984 two_stage_opamp_dummy_magic_23_0.V_source.n45 two_stage_opamp_dummy_magic_23_0.V_source.n38 1.738
R7985 two_stage_opamp_dummy_magic_23_0.V_source.n48 two_stage_opamp_dummy_magic_23_0.V_source.n47 0.833833
R7986 two_stage_opamp_dummy_magic_23_0.V_source.n47 two_stage_opamp_dummy_magic_23_0.V_source.n45 0.633833
R7987 two_stage_opamp_dummy_magic_23_0.V_source.n33 two_stage_opamp_dummy_magic_23_0.V_source.n30 0.563
R7988 two_stage_opamp_dummy_magic_23_0.V_source.n30 two_stage_opamp_dummy_magic_23_0.V_source.n21 0.563
R7989 two_stage_opamp_dummy_magic_23_0.V_source.n27 two_stage_opamp_dummy_magic_23_0.V_source.n26 0.563
R7990 two_stage_opamp_dummy_magic_23_0.V_source.n27 two_stage_opamp_dummy_magic_23_0.V_source.n20 0.563
R7991 two_stage_opamp_dummy_magic_23_0.V_source.n36 two_stage_opamp_dummy_magic_23_0.V_source.n20 0.563
R7992 two_stage_opamp_dummy_magic_23_0.V_source.n37 two_stage_opamp_dummy_magic_23_0.V_source.n19 0.563
R7993 two_stage_opamp_dummy_magic_23_0.V_source.n19 two_stage_opamp_dummy_magic_23_0.V_source.n6 0.563
R7994 two_stage_opamp_dummy_magic_23_0.V_source.n9 two_stage_opamp_dummy_magic_23_0.V_source.n6 0.563
R7995 two_stage_opamp_dummy_magic_23_0.V_source.n15 two_stage_opamp_dummy_magic_23_0.V_source.n12 0.563
R7996 two_stage_opamp_dummy_magic_23_0.V_source.n16 two_stage_opamp_dummy_magic_23_0.V_source.n15 0.563
R7997 two_stage_opamp_dummy_magic_23_0.V_source.n38 two_stage_opamp_dummy_magic_23_0.V_source.n5 0.563
R7998 two_stage_opamp_dummy_magic_23_0.V_source.n70 two_stage_opamp_dummy_magic_23_0.V_source.n69 0.563
R7999 two_stage_opamp_dummy_magic_23_0.V_source.n66 two_stage_opamp_dummy_magic_23_0.V_source.n0 0.563
R8000 two_stage_opamp_dummy_magic_23_0.V_source.n60 two_stage_opamp_dummy_magic_23_0.V_source.n0 0.563
R8001 two_stage_opamp_dummy_magic_23_0.V_source.n60 two_stage_opamp_dummy_magic_23_0.V_source.n59 0.563
R8002 two_stage_opamp_dummy_magic_23_0.V_source.n59 two_stage_opamp_dummy_magic_23_0.V_source.n56 0.563
R8003 two_stage_opamp_dummy_magic_23_0.V_source.n56 two_stage_opamp_dummy_magic_23_0.V_source.n2 0.563
R8004 two_stage_opamp_dummy_magic_23_0.V_source.n44 two_stage_opamp_dummy_magic_23_0.V_source.n2 0.563
R8005 two_stage_opamp_dummy_magic_23_0.V_source.n44 two_stage_opamp_dummy_magic_23_0.V_source.n43 0.563
R8006 two_stage_opamp_dummy_magic_23_0.V_source.n49 two_stage_opamp_dummy_magic_23_0.V_source.n3 0.563
R8007 two_stage_opamp_dummy_magic_23_0.V_source.n52 two_stage_opamp_dummy_magic_23_0.V_source.n49 0.563
R8008 two_stage_opamp_dummy_magic_23_0.V_source.n53 two_stage_opamp_dummy_magic_23_0.V_source.n52 0.563
R8009 two_stage_opamp_dummy_magic_23_0.V_source.n53 two_stage_opamp_dummy_magic_23_0.V_source.n1 0.563
R8010 two_stage_opamp_dummy_magic_23_0.V_source.n63 two_stage_opamp_dummy_magic_23_0.V_source.n1 0.563
R8011 two_stage_opamp_dummy_magic_23_0.V_source.n70 two_stage_opamp_dummy_magic_23_0.V_source.n63 0.563
R8012 bgr_11_0.V_mir2.n20 bgr_11_0.V_mir2.n19 325.473
R8013 bgr_11_0.V_mir2.n13 bgr_11_0.V_mir2.n12 325.473
R8014 bgr_11_0.V_mir2.n8 bgr_11_0.V_mir2.n7 325.473
R8015 bgr_11_0.V_mir2.n16 bgr_11_0.V_mir2.t20 310.488
R8016 bgr_11_0.V_mir2.n9 bgr_11_0.V_mir2.t21 310.488
R8017 bgr_11_0.V_mir2.n4 bgr_11_0.V_mir2.t19 310.488
R8018 bgr_11_0.V_mir2.n2 bgr_11_0.V_mir2.t15 278.312
R8019 bgr_11_0.V_mir2.n2 bgr_11_0.V_mir2.n1 228.939
R8020 bgr_11_0.V_mir2.n3 bgr_11_0.V_mir2.n0 224.439
R8021 bgr_11_0.V_mir2.n18 bgr_11_0.V_mir2.t13 184.097
R8022 bgr_11_0.V_mir2.n11 bgr_11_0.V_mir2.t11 184.097
R8023 bgr_11_0.V_mir2.n6 bgr_11_0.V_mir2.t3 184.097
R8024 bgr_11_0.V_mir2.n17 bgr_11_0.V_mir2.n16 167.094
R8025 bgr_11_0.V_mir2.n10 bgr_11_0.V_mir2.n9 167.094
R8026 bgr_11_0.V_mir2.n5 bgr_11_0.V_mir2.n4 167.094
R8027 bgr_11_0.V_mir2.n13 bgr_11_0.V_mir2.n11 152
R8028 bgr_11_0.V_mir2.n8 bgr_11_0.V_mir2.n6 152
R8029 bgr_11_0.V_mir2.n19 bgr_11_0.V_mir2.n18 152
R8030 bgr_11_0.V_mir2.n16 bgr_11_0.V_mir2.t18 120.501
R8031 bgr_11_0.V_mir2.n17 bgr_11_0.V_mir2.t9 120.501
R8032 bgr_11_0.V_mir2.n9 bgr_11_0.V_mir2.t17 120.501
R8033 bgr_11_0.V_mir2.n10 bgr_11_0.V_mir2.t5 120.501
R8034 bgr_11_0.V_mir2.n4 bgr_11_0.V_mir2.t22 120.501
R8035 bgr_11_0.V_mir2.n5 bgr_11_0.V_mir2.t7 120.501
R8036 bgr_11_0.V_mir2.n1 bgr_11_0.V_mir2.t16 48.0005
R8037 bgr_11_0.V_mir2.n1 bgr_11_0.V_mir2.t2 48.0005
R8038 bgr_11_0.V_mir2.n0 bgr_11_0.V_mir2.t1 48.0005
R8039 bgr_11_0.V_mir2.n0 bgr_11_0.V_mir2.t0 48.0005
R8040 bgr_11_0.V_mir2.n18 bgr_11_0.V_mir2.n17 40.7027
R8041 bgr_11_0.V_mir2.n11 bgr_11_0.V_mir2.n10 40.7027
R8042 bgr_11_0.V_mir2.n6 bgr_11_0.V_mir2.n5 40.7027
R8043 bgr_11_0.V_mir2.n12 bgr_11_0.V_mir2.t6 39.4005
R8044 bgr_11_0.V_mir2.n12 bgr_11_0.V_mir2.t12 39.4005
R8045 bgr_11_0.V_mir2.n7 bgr_11_0.V_mir2.t8 39.4005
R8046 bgr_11_0.V_mir2.n7 bgr_11_0.V_mir2.t4 39.4005
R8047 bgr_11_0.V_mir2.n20 bgr_11_0.V_mir2.t10 39.4005
R8048 bgr_11_0.V_mir2.t14 bgr_11_0.V_mir2.n20 39.4005
R8049 bgr_11_0.V_mir2.n14 bgr_11_0.V_mir2.n13 15.9255
R8050 bgr_11_0.V_mir2.n14 bgr_11_0.V_mir2.n8 15.9255
R8051 bgr_11_0.V_mir2.n19 bgr_11_0.V_mir2.n15 9.3005
R8052 bgr_11_0.V_mir2.n3 bgr_11_0.V_mir2.n2 5.8755
R8053 bgr_11_0.V_mir2.n15 bgr_11_0.V_mir2.n14 4.5005
R8054 bgr_11_0.V_mir2.n15 bgr_11_0.V_mir2.n3 0.78175
R8055 bgr_11_0.V_TOP.n0 bgr_11_0.V_TOP.t26 369.534
R8056 bgr_11_0.V_TOP.n23 bgr_11_0.V_TOP.n21 339.961
R8057 bgr_11_0.V_TOP.n23 bgr_11_0.V_TOP.n22 339.272
R8058 bgr_11_0.V_TOP.n19 bgr_11_0.V_TOP.n18 339.272
R8059 bgr_11_0.V_TOP.n27 bgr_11_0.V_TOP.n26 339.272
R8060 bgr_11_0.V_TOP.n29 bgr_11_0.V_TOP.n28 339.272
R8061 bgr_11_0.V_TOP.n24 bgr_11_0.V_TOP.n20 334.772
R8062 bgr_11_0.V_TOP.n39 bgr_11_0.V_TOP.n38 224.934
R8063 bgr_11_0.V_TOP.n38 bgr_11_0.V_TOP.n37 224.934
R8064 bgr_11_0.V_TOP.n37 bgr_11_0.V_TOP.n36 224.934
R8065 bgr_11_0.V_TOP.n36 bgr_11_0.V_TOP.n35 224.934
R8066 bgr_11_0.V_TOP.n35 bgr_11_0.V_TOP.n34 224.934
R8067 bgr_11_0.V_TOP.n34 bgr_11_0.V_TOP.n33 224.934
R8068 bgr_11_0.V_TOP.n33 bgr_11_0.V_TOP.n32 224.934
R8069 bgr_11_0.V_TOP.n1 bgr_11_0.V_TOP.n0 224.934
R8070 bgr_11_0.V_TOP.n2 bgr_11_0.V_TOP.n1 224.934
R8071 bgr_11_0.V_TOP.n3 bgr_11_0.V_TOP.n2 224.934
R8072 bgr_11_0.V_TOP.n4 bgr_11_0.V_TOP.n3 224.934
R8073 bgr_11_0.V_TOP.n5 bgr_11_0.V_TOP.n4 224.934
R8074 bgr_11_0.V_TOP bgr_11_0.V_TOP.t47 214.222
R8075 bgr_11_0.V_TOP.n31 bgr_11_0.V_TOP.n30 163.175
R8076 bgr_11_0.V_TOP.n39 bgr_11_0.V_TOP.t24 144.601
R8077 bgr_11_0.V_TOP.n38 bgr_11_0.V_TOP.t36 144.601
R8078 bgr_11_0.V_TOP.n37 bgr_11_0.V_TOP.t41 144.601
R8079 bgr_11_0.V_TOP.n36 bgr_11_0.V_TOP.t14 144.601
R8080 bgr_11_0.V_TOP.n35 bgr_11_0.V_TOP.t49 144.601
R8081 bgr_11_0.V_TOP.n34 bgr_11_0.V_TOP.t25 144.601
R8082 bgr_11_0.V_TOP.n33 bgr_11_0.V_TOP.t37 144.601
R8083 bgr_11_0.V_TOP.n32 bgr_11_0.V_TOP.t43 144.601
R8084 bgr_11_0.V_TOP.n0 bgr_11_0.V_TOP.t29 144.601
R8085 bgr_11_0.V_TOP.n1 bgr_11_0.V_TOP.t48 144.601
R8086 bgr_11_0.V_TOP.n2 bgr_11_0.V_TOP.t40 144.601
R8087 bgr_11_0.V_TOP.n3 bgr_11_0.V_TOP.t30 144.601
R8088 bgr_11_0.V_TOP.n4 bgr_11_0.V_TOP.t16 144.601
R8089 bgr_11_0.V_TOP.n5 bgr_11_0.V_TOP.t19 144.601
R8090 bgr_11_0.V_TOP.n17 bgr_11_0.V_TOP.t0 108.424
R8091 bgr_11_0.V_TOP.n30 bgr_11_0.V_TOP.t7 95.4467
R8092 bgr_11_0.V_TOP bgr_11_0.V_TOP.n39 69.6227
R8093 bgr_11_0.V_TOP.n32 bgr_11_0.V_TOP.n31 69.6227
R8094 bgr_11_0.V_TOP.n31 bgr_11_0.V_TOP.n5 69.6227
R8095 bgr_11_0.V_TOP.n18 bgr_11_0.V_TOP.t4 39.4005
R8096 bgr_11_0.V_TOP.n18 bgr_11_0.V_TOP.t12 39.4005
R8097 bgr_11_0.V_TOP.n20 bgr_11_0.V_TOP.t8 39.4005
R8098 bgr_11_0.V_TOP.n20 bgr_11_0.V_TOP.t13 39.4005
R8099 bgr_11_0.V_TOP.n22 bgr_11_0.V_TOP.t1 39.4005
R8100 bgr_11_0.V_TOP.n22 bgr_11_0.V_TOP.t3 39.4005
R8101 bgr_11_0.V_TOP.n21 bgr_11_0.V_TOP.t6 39.4005
R8102 bgr_11_0.V_TOP.n21 bgr_11_0.V_TOP.t2 39.4005
R8103 bgr_11_0.V_TOP.n26 bgr_11_0.V_TOP.t10 39.4005
R8104 bgr_11_0.V_TOP.n26 bgr_11_0.V_TOP.t11 39.4005
R8105 bgr_11_0.V_TOP.n28 bgr_11_0.V_TOP.t9 39.4005
R8106 bgr_11_0.V_TOP.n28 bgr_11_0.V_TOP.t5 39.4005
R8107 bgr_11_0.V_TOP.n17 bgr_11_0.V_TOP.n16 37.1479
R8108 bgr_11_0.V_TOP.n19 bgr_11_0.V_TOP.n17 27.8371
R8109 bgr_11_0.V_TOP.n24 bgr_11_0.V_TOP.n23 8.313
R8110 bgr_11_0.V_TOP.n30 bgr_11_0.V_TOP.n29 5.188
R8111 bgr_11_0.V_TOP.n6 bgr_11_0.V_TOP.t34 4.8295
R8112 bgr_11_0.V_TOP.n7 bgr_11_0.V_TOP.t21 4.8295
R8113 bgr_11_0.V_TOP.n8 bgr_11_0.V_TOP.t23 4.8295
R8114 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.t45 4.8295
R8115 bgr_11_0.V_TOP.n10 bgr_11_0.V_TOP.t33 4.8295
R8116 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.t18 4.8295
R8117 bgr_11_0.V_TOP.n12 bgr_11_0.V_TOP.t22 4.8295
R8118 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.t44 4.8295
R8119 bgr_11_0.V_TOP.n14 bgr_11_0.V_TOP.t35 4.8295
R8120 bgr_11_0.V_TOP.n6 bgr_11_0.V_TOP.t39 4.5005
R8121 bgr_11_0.V_TOP.n7 bgr_11_0.V_TOP.t32 4.5005
R8122 bgr_11_0.V_TOP.n8 bgr_11_0.V_TOP.t31 4.5005
R8123 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.t20 4.5005
R8124 bgr_11_0.V_TOP.n10 bgr_11_0.V_TOP.t38 4.5005
R8125 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.t28 4.5005
R8126 bgr_11_0.V_TOP.n12 bgr_11_0.V_TOP.t27 4.5005
R8127 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.t17 4.5005
R8128 bgr_11_0.V_TOP.n16 bgr_11_0.V_TOP.t46 4.5005
R8129 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.t15 4.5005
R8130 bgr_11_0.V_TOP.n14 bgr_11_0.V_TOP.t42 4.5005
R8131 bgr_11_0.V_TOP.n25 bgr_11_0.V_TOP.n24 4.5005
R8132 bgr_11_0.V_TOP.n29 bgr_11_0.V_TOP.n27 2.1255
R8133 bgr_11_0.V_TOP.n27 bgr_11_0.V_TOP.n25 2.1255
R8134 bgr_11_0.V_TOP.n25 bgr_11_0.V_TOP.n19 2.1255
R8135 bgr_11_0.V_TOP.n7 bgr_11_0.V_TOP.n6 0.3295
R8136 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.n8 0.3295
R8137 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.n10 0.3295
R8138 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.n12 0.3295
R8139 bgr_11_0.V_TOP.n16 bgr_11_0.V_TOP.n15 0.3295
R8140 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.n14 0.3295
R8141 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.n7 0.2825
R8142 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.n9 0.2825
R8143 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.n11 0.2825
R8144 bgr_11_0.V_TOP.n14 bgr_11_0.V_TOP.n13 0.2825
R8145 bgr_11_0.Vin-.n7 bgr_11_0.Vin-.t10 688.859
R8146 bgr_11_0.Vin-.n9 bgr_11_0.Vin-.n8 514.134
R8147 bgr_11_0.Vin-.n6 bgr_11_0.Vin-.n5 351.522
R8148 bgr_11_0.Vin-.n11 bgr_11_0.Vin-.n10 213.4
R8149 bgr_11_0.Vin-.n7 bgr_11_0.Vin-.t8 174.726
R8150 bgr_11_0.Vin-.n8 bgr_11_0.Vin-.t11 174.726
R8151 bgr_11_0.Vin-.n9 bgr_11_0.Vin-.t9 174.726
R8152 bgr_11_0.Vin-.n10 bgr_11_0.Vin-.t12 174.726
R8153 bgr_11_0.Vin-.n4 bgr_11_0.Vin-.n2 173.029
R8154 bgr_11_0.Vin-.n4 bgr_11_0.Vin-.n3 168.654
R8155 bgr_11_0.Vin-.n8 bgr_11_0.Vin-.n7 128.534
R8156 bgr_11_0.Vin-.n10 bgr_11_0.Vin-.n9 128.534
R8157 bgr_11_0.Vin-.n12 bgr_11_0.Vin-.t0 119.099
R8158 bgr_11_0.Vin-.n16 bgr_11_0.Vin-.n15 83.5719
R8159 bgr_11_0.Vin-.n1 bgr_11_0.Vin-.n0 83.5719
R8160 bgr_11_0.Vin-.n19 bgr_11_0.Vin-.n1 73.8495
R8161 bgr_11_0.Vin-.t3 bgr_11_0.Vin-.n14 65.0341
R8162 bgr_11_0.Vin-.n5 bgr_11_0.Vin-.t2 39.4005
R8163 bgr_11_0.Vin-.n5 bgr_11_0.Vin-.t1 39.4005
R8164 bgr_11_0.Vin-.n13 bgr_11_0.Vin-.n12 28.813
R8165 bgr_11_0.Vin-.n15 bgr_11_0.Vin-.n1 26.074
R8166 bgr_11_0.Vin-.n12 bgr_11_0.Vin-.n11 16.188
R8167 bgr_11_0.Vin-.n3 bgr_11_0.Vin-.t5 13.1338
R8168 bgr_11_0.Vin-.n3 bgr_11_0.Vin-.t6 13.1338
R8169 bgr_11_0.Vin-.n2 bgr_11_0.Vin-.t7 13.1338
R8170 bgr_11_0.Vin-.n2 bgr_11_0.Vin-.t4 13.1338
R8171 bgr_11_0.Vin-.n11 bgr_11_0.Vin-.n6 11.2193
R8172 bgr_11_0.Vin-.n6 bgr_11_0.Vin-.n4 3.8755
R8173 bgr_11_0.Vin-.n16 bgr_11_0.Vin-.n14 1.56483
R8174 bgr_11_0.Vin-.n18 bgr_11_0.Vin-.n17 1.5505
R8175 bgr_11_0.Vin-.n17 bgr_11_0.Vin-.n0 0.885803
R8176 bgr_11_0.Vin-.n17 bgr_11_0.Vin-.n16 0.77514
R8177 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_11_0.Vin-.n0 0.756696
R8178 bgr_11_0.Vin-.n19 bgr_11_0.Vin-.n18 0.711459
R8179 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_11_0.Vin-.n19 0.576566
R8180 bgr_11_0.Vin-.n14 bgr_11_0.Vin-.n13 0.531499
R8181 bgr_11_0.Vin-.n15 bgr_11_0.Vin-.t3 0.290206
R8182 bgr_11_0.Vin-.n18 bgr_11_0.Vin-.n13 0.00817857
R8183 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n0 345.264
R8184 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n1 344.7
R8185 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n3 292.5
R8186 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n22 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t14 122.442
R8187 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n7 118.861
R8188 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n9 118.861
R8189 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n13 118.861
R8190 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n17 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n16 118.861
R8191 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n20 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n19 118.861
R8192 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n2 52.763
R8193 bgr_11_0.V_CMFB_S3 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n4 51.7297
R8194 bgr_11_0.V_CMFB_S3 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n22 47.5943
R8195 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t12 39.4005
R8196 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t15 39.4005
R8197 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t16 39.4005
R8198 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t1 39.4005
R8199 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t0 39.4005
R8200 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t13 39.4005
R8201 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t3 19.7005
R8202 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t7 19.7005
R8203 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t2 19.7005
R8204 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t10 19.7005
R8205 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t5 19.7005
R8206 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t9 19.7005
R8207 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t4 19.7005
R8208 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t8 19.7005
R8209 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n19 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t11 19.7005
R8210 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n19 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t6 19.7005
R8211 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n22 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n21 6.28175
R8212 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n8 5.60467
R8213 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n20 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n18 5.54217
R8214 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n6 5.54217
R8215 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n10 5.04217
R8216 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n12 5.04217
R8217 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n17 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n5 5.04217
R8218 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n21 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n20 5.04217
R8219 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n6 4.97967
R8220 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n14 4.97967
R8221 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n18 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n17 4.97967
R8222 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n18 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n15 0.563
R8223 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n6 0.563
R8224 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n11 0.563
R8225 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n5 0.563
R8226 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n21 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n5 0.563
R8227 bgr_11_0.PFET_GATE_10uA.n4 bgr_11_0.PFET_GATE_10uA.t23 369.534
R8228 bgr_11_0.PFET_GATE_10uA.n3 bgr_11_0.PFET_GATE_10uA.t10 369.534
R8229 bgr_11_0.PFET_GATE_10uA.n23 bgr_11_0.PFET_GATE_10uA.t28 369.534
R8230 bgr_11_0.PFET_GATE_10uA.n18 bgr_11_0.PFET_GATE_10uA.t11 369.534
R8231 bgr_11_0.PFET_GATE_10uA.n1 bgr_11_0.PFET_GATE_10uA.t21 369.534
R8232 bgr_11_0.PFET_GATE_10uA.n0 bgr_11_0.PFET_GATE_10uA.t20 369.534
R8233 bgr_11_0.PFET_GATE_10uA.n8 bgr_11_0.PFET_GATE_10uA.n6 341.397
R8234 bgr_11_0.PFET_GATE_10uA.n10 bgr_11_0.PFET_GATE_10uA.n9 339.272
R8235 bgr_11_0.PFET_GATE_10uA.n8 bgr_11_0.PFET_GATE_10uA.n7 339.272
R8236 bgr_11_0.PFET_GATE_10uA.n13 bgr_11_0.PFET_GATE_10uA.n12 334.772
R8237 bgr_11_0.PFET_GATE_10uA.n14 bgr_11_0.PFET_GATE_10uA.t13 238.322
R8238 bgr_11_0.PFET_GATE_10uA.n14 bgr_11_0.PFET_GATE_10uA.t26 238.322
R8239 bgr_11_0.PFET_GATE_10uA.n4 bgr_11_0.PFET_GATE_10uA.t24 192.8
R8240 bgr_11_0.PFET_GATE_10uA.n3 bgr_11_0.PFET_GATE_10uA.t17 192.8
R8241 bgr_11_0.PFET_GATE_10uA.n25 bgr_11_0.PFET_GATE_10uA.t16 192.8
R8242 bgr_11_0.PFET_GATE_10uA.n24 bgr_11_0.PFET_GATE_10uA.t15 192.8
R8243 bgr_11_0.PFET_GATE_10uA.n23 bgr_11_0.PFET_GATE_10uA.t22 192.8
R8244 bgr_11_0.PFET_GATE_10uA.n18 bgr_11_0.PFET_GATE_10uA.t18 192.8
R8245 bgr_11_0.PFET_GATE_10uA.n19 bgr_11_0.PFET_GATE_10uA.t25 192.8
R8246 bgr_11_0.PFET_GATE_10uA.n20 bgr_11_0.PFET_GATE_10uA.t12 192.8
R8247 bgr_11_0.PFET_GATE_10uA.n21 bgr_11_0.PFET_GATE_10uA.t19 192.8
R8248 bgr_11_0.PFET_GATE_10uA.n22 bgr_11_0.PFET_GATE_10uA.t29 192.8
R8249 bgr_11_0.PFET_GATE_10uA.n1 bgr_11_0.PFET_GATE_10uA.t14 192.8
R8250 bgr_11_0.PFET_GATE_10uA.n0 bgr_11_0.PFET_GATE_10uA.t27 192.8
R8251 bgr_11_0.PFET_GATE_10uA.n25 bgr_11_0.PFET_GATE_10uA.n24 176.733
R8252 bgr_11_0.PFET_GATE_10uA.n24 bgr_11_0.PFET_GATE_10uA.n23 176.733
R8253 bgr_11_0.PFET_GATE_10uA.n19 bgr_11_0.PFET_GATE_10uA.n18 176.733
R8254 bgr_11_0.PFET_GATE_10uA.n20 bgr_11_0.PFET_GATE_10uA.n19 176.733
R8255 bgr_11_0.PFET_GATE_10uA.n21 bgr_11_0.PFET_GATE_10uA.n20 176.733
R8256 bgr_11_0.PFET_GATE_10uA.n22 bgr_11_0.PFET_GATE_10uA.n21 176.733
R8257 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n2 171.321
R8258 bgr_11_0.PFET_GATE_10uA.n17 bgr_11_0.PFET_GATE_10uA.n5 168.166
R8259 bgr_11_0.PFET_GATE_10uA.n15 bgr_11_0.PFET_GATE_10uA.n14 167.519
R8260 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n26 166.071
R8261 bgr_11_0.PFET_GATE_10uA.n15 bgr_11_0.PFET_GATE_10uA.t9 137.48
R8262 bgr_11_0.PFET_GATE_10uA.n11 bgr_11_0.PFET_GATE_10uA.t2 100.635
R8263 bgr_11_0.PFET_GATE_10uA.n5 bgr_11_0.PFET_GATE_10uA.n4 56.2338
R8264 bgr_11_0.PFET_GATE_10uA.n5 bgr_11_0.PFET_GATE_10uA.n3 56.2338
R8265 bgr_11_0.PFET_GATE_10uA.n26 bgr_11_0.PFET_GATE_10uA.n25 56.2338
R8266 bgr_11_0.PFET_GATE_10uA.n26 bgr_11_0.PFET_GATE_10uA.n22 56.2338
R8267 bgr_11_0.PFET_GATE_10uA.n2 bgr_11_0.PFET_GATE_10uA.n1 56.2338
R8268 bgr_11_0.PFET_GATE_10uA.n2 bgr_11_0.PFET_GATE_10uA.n0 56.2338
R8269 bgr_11_0.PFET_GATE_10uA.n12 bgr_11_0.PFET_GATE_10uA.t1 39.4005
R8270 bgr_11_0.PFET_GATE_10uA.n12 bgr_11_0.PFET_GATE_10uA.t4 39.4005
R8271 bgr_11_0.PFET_GATE_10uA.n9 bgr_11_0.PFET_GATE_10uA.t6 39.4005
R8272 bgr_11_0.PFET_GATE_10uA.n9 bgr_11_0.PFET_GATE_10uA.t8 39.4005
R8273 bgr_11_0.PFET_GATE_10uA.n7 bgr_11_0.PFET_GATE_10uA.t5 39.4005
R8274 bgr_11_0.PFET_GATE_10uA.n7 bgr_11_0.PFET_GATE_10uA.t7 39.4005
R8275 bgr_11_0.PFET_GATE_10uA.n6 bgr_11_0.PFET_GATE_10uA.t3 39.4005
R8276 bgr_11_0.PFET_GATE_10uA.n6 bgr_11_0.PFET_GATE_10uA.t0 39.4005
R8277 bgr_11_0.PFET_GATE_10uA.n17 bgr_11_0.PFET_GATE_10uA.n16 27.5005
R8278 bgr_11_0.PFET_GATE_10uA.n16 bgr_11_0.PFET_GATE_10uA.n13 9.53175
R8279 bgr_11_0.PFET_GATE_10uA.n13 bgr_11_0.PFET_GATE_10uA.n11 4.5005
R8280 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n17 2.34425
R8281 bgr_11_0.PFET_GATE_10uA.n10 bgr_11_0.PFET_GATE_10uA.n8 2.1255
R8282 bgr_11_0.PFET_GATE_10uA.n11 bgr_11_0.PFET_GATE_10uA.n10 2.1255
R8283 bgr_11_0.PFET_GATE_10uA.n16 bgr_11_0.PFET_GATE_10uA.n15 1.688
R8284 two_stage_opamp_dummy_magic_23_0.Vb3.n25 two_stage_opamp_dummy_magic_23_0.Vb3.t20 768.551
R8285 two_stage_opamp_dummy_magic_23_0.Vb3.n19 two_stage_opamp_dummy_magic_23_0.Vb3.t8 611.739
R8286 two_stage_opamp_dummy_magic_23_0.Vb3.n15 two_stage_opamp_dummy_magic_23_0.Vb3.t25 611.739
R8287 two_stage_opamp_dummy_magic_23_0.Vb3.n10 two_stage_opamp_dummy_magic_23_0.Vb3.t22 611.739
R8288 two_stage_opamp_dummy_magic_23_0.Vb3.n6 two_stage_opamp_dummy_magic_23_0.Vb3.t16 611.739
R8289 two_stage_opamp_dummy_magic_23_0.Vb3.n24 two_stage_opamp_dummy_magic_23_0.Vb3.n23 428.976
R8290 two_stage_opamp_dummy_magic_23_0.Vb3.n24 two_stage_opamp_dummy_magic_23_0.Vb3.n14 428.445
R8291 two_stage_opamp_dummy_magic_23_0.Vb3.n19 two_stage_opamp_dummy_magic_23_0.Vb3.t11 421.75
R8292 two_stage_opamp_dummy_magic_23_0.Vb3.n20 two_stage_opamp_dummy_magic_23_0.Vb3.t28 421.75
R8293 two_stage_opamp_dummy_magic_23_0.Vb3.n21 two_stage_opamp_dummy_magic_23_0.Vb3.t18 421.75
R8294 two_stage_opamp_dummy_magic_23_0.Vb3.n22 two_stage_opamp_dummy_magic_23_0.Vb3.t15 421.75
R8295 two_stage_opamp_dummy_magic_23_0.Vb3.n15 two_stage_opamp_dummy_magic_23_0.Vb3.t27 421.75
R8296 two_stage_opamp_dummy_magic_23_0.Vb3.n16 two_stage_opamp_dummy_magic_23_0.Vb3.t10 421.75
R8297 two_stage_opamp_dummy_magic_23_0.Vb3.n17 two_stage_opamp_dummy_magic_23_0.Vb3.t14 421.75
R8298 two_stage_opamp_dummy_magic_23_0.Vb3.n18 two_stage_opamp_dummy_magic_23_0.Vb3.t12 421.75
R8299 two_stage_opamp_dummy_magic_23_0.Vb3.n10 two_stage_opamp_dummy_magic_23_0.Vb3.t24 421.75
R8300 two_stage_opamp_dummy_magic_23_0.Vb3.n11 two_stage_opamp_dummy_magic_23_0.Vb3.t21 421.75
R8301 two_stage_opamp_dummy_magic_23_0.Vb3.n12 two_stage_opamp_dummy_magic_23_0.Vb3.t17 421.75
R8302 two_stage_opamp_dummy_magic_23_0.Vb3.n13 two_stage_opamp_dummy_magic_23_0.Vb3.t13 421.75
R8303 two_stage_opamp_dummy_magic_23_0.Vb3.n6 two_stage_opamp_dummy_magic_23_0.Vb3.t19 421.75
R8304 two_stage_opamp_dummy_magic_23_0.Vb3.n7 two_stage_opamp_dummy_magic_23_0.Vb3.t23 421.75
R8305 two_stage_opamp_dummy_magic_23_0.Vb3.n8 two_stage_opamp_dummy_magic_23_0.Vb3.t26 421.75
R8306 two_stage_opamp_dummy_magic_23_0.Vb3.n9 two_stage_opamp_dummy_magic_23_0.Vb3.t9 421.75
R8307 two_stage_opamp_dummy_magic_23_0.Vb3.n20 two_stage_opamp_dummy_magic_23_0.Vb3.n19 167.094
R8308 two_stage_opamp_dummy_magic_23_0.Vb3.n21 two_stage_opamp_dummy_magic_23_0.Vb3.n20 167.094
R8309 two_stage_opamp_dummy_magic_23_0.Vb3.n22 two_stage_opamp_dummy_magic_23_0.Vb3.n21 167.094
R8310 two_stage_opamp_dummy_magic_23_0.Vb3.n16 two_stage_opamp_dummy_magic_23_0.Vb3.n15 167.094
R8311 two_stage_opamp_dummy_magic_23_0.Vb3.n17 two_stage_opamp_dummy_magic_23_0.Vb3.n16 167.094
R8312 two_stage_opamp_dummy_magic_23_0.Vb3.n18 two_stage_opamp_dummy_magic_23_0.Vb3.n17 167.094
R8313 two_stage_opamp_dummy_magic_23_0.Vb3.n11 two_stage_opamp_dummy_magic_23_0.Vb3.n10 167.094
R8314 two_stage_opamp_dummy_magic_23_0.Vb3.n12 two_stage_opamp_dummy_magic_23_0.Vb3.n11 167.094
R8315 two_stage_opamp_dummy_magic_23_0.Vb3.n13 two_stage_opamp_dummy_magic_23_0.Vb3.n12 167.094
R8316 two_stage_opamp_dummy_magic_23_0.Vb3.n7 two_stage_opamp_dummy_magic_23_0.Vb3.n6 167.094
R8317 two_stage_opamp_dummy_magic_23_0.Vb3.n8 two_stage_opamp_dummy_magic_23_0.Vb3.n7 167.094
R8318 two_stage_opamp_dummy_magic_23_0.Vb3.n9 two_stage_opamp_dummy_magic_23_0.Vb3.n8 167.094
R8319 two_stage_opamp_dummy_magic_23_0.Vb3.n3 two_stage_opamp_dummy_magic_23_0.Vb3.n1 139.639
R8320 two_stage_opamp_dummy_magic_23_0.Vb3.n3 two_stage_opamp_dummy_magic_23_0.Vb3.n2 139.638
R8321 two_stage_opamp_dummy_magic_23_0.Vb3.n4 two_stage_opamp_dummy_magic_23_0.Vb3.n0 134.577
R8322 two_stage_opamp_dummy_magic_23_0.Vb3.n26 two_stage_opamp_dummy_magic_23_0.Vb3.n5 73.3151
R8323 bgr_11_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_23_0.Vb3.n26 52.6818
R8324 bgr_11_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_23_0.Vb3.n4 41.063
R8325 two_stage_opamp_dummy_magic_23_0.Vb3.n23 two_stage_opamp_dummy_magic_23_0.Vb3.n22 35.3472
R8326 two_stage_opamp_dummy_magic_23_0.Vb3.n23 two_stage_opamp_dummy_magic_23_0.Vb3.n18 35.3472
R8327 two_stage_opamp_dummy_magic_23_0.Vb3.n14 two_stage_opamp_dummy_magic_23_0.Vb3.n13 35.3472
R8328 two_stage_opamp_dummy_magic_23_0.Vb3.n14 two_stage_opamp_dummy_magic_23_0.Vb3.n9 35.3472
R8329 two_stage_opamp_dummy_magic_23_0.Vb3.n0 two_stage_opamp_dummy_magic_23_0.Vb3.t2 24.0005
R8330 two_stage_opamp_dummy_magic_23_0.Vb3.n0 two_stage_opamp_dummy_magic_23_0.Vb3.t3 24.0005
R8331 two_stage_opamp_dummy_magic_23_0.Vb3.n2 two_stage_opamp_dummy_magic_23_0.Vb3.t0 24.0005
R8332 two_stage_opamp_dummy_magic_23_0.Vb3.n2 two_stage_opamp_dummy_magic_23_0.Vb3.t6 24.0005
R8333 two_stage_opamp_dummy_magic_23_0.Vb3.n1 two_stage_opamp_dummy_magic_23_0.Vb3.t1 24.0005
R8334 two_stage_opamp_dummy_magic_23_0.Vb3.n1 two_stage_opamp_dummy_magic_23_0.Vb3.t4 24.0005
R8335 two_stage_opamp_dummy_magic_23_0.Vb3.n25 two_stage_opamp_dummy_magic_23_0.Vb3.n24 14.3443
R8336 two_stage_opamp_dummy_magic_23_0.Vb3.n5 two_stage_opamp_dummy_magic_23_0.Vb3.t5 11.2576
R8337 two_stage_opamp_dummy_magic_23_0.Vb3.n5 two_stage_opamp_dummy_magic_23_0.Vb3.t7 11.2576
R8338 two_stage_opamp_dummy_magic_23_0.Vb3.n4 two_stage_opamp_dummy_magic_23_0.Vb3.n3 4.5005
R8339 two_stage_opamp_dummy_magic_23_0.Vb3.n26 two_stage_opamp_dummy_magic_23_0.Vb3.n25 1.21925
R8340 two_stage_opamp_dummy_magic_23_0.VD4.n10 two_stage_opamp_dummy_magic_23_0.VD4.t10 672.293
R8341 two_stage_opamp_dummy_magic_23_0.VD4.n13 two_stage_opamp_dummy_magic_23_0.VD4.t13 672.293
R8342 two_stage_opamp_dummy_magic_23_0.VD4.t11 two_stage_opamp_dummy_magic_23_0.VD4.n11 213.131
R8343 two_stage_opamp_dummy_magic_23_0.VD4.n12 two_stage_opamp_dummy_magic_23_0.VD4.t14 213.131
R8344 two_stage_opamp_dummy_magic_23_0.VD4.t20 two_stage_opamp_dummy_magic_23_0.VD4.t11 146.155
R8345 two_stage_opamp_dummy_magic_23_0.VD4.t24 two_stage_opamp_dummy_magic_23_0.VD4.t20 146.155
R8346 two_stage_opamp_dummy_magic_23_0.VD4.t30 two_stage_opamp_dummy_magic_23_0.VD4.t24 146.155
R8347 two_stage_opamp_dummy_magic_23_0.VD4.t34 two_stage_opamp_dummy_magic_23_0.VD4.t30 146.155
R8348 two_stage_opamp_dummy_magic_23_0.VD4.t36 two_stage_opamp_dummy_magic_23_0.VD4.t34 146.155
R8349 two_stage_opamp_dummy_magic_23_0.VD4.t18 two_stage_opamp_dummy_magic_23_0.VD4.t36 146.155
R8350 two_stage_opamp_dummy_magic_23_0.VD4.t22 two_stage_opamp_dummy_magic_23_0.VD4.t18 146.155
R8351 two_stage_opamp_dummy_magic_23_0.VD4.t26 two_stage_opamp_dummy_magic_23_0.VD4.t22 146.155
R8352 two_stage_opamp_dummy_magic_23_0.VD4.t32 two_stage_opamp_dummy_magic_23_0.VD4.t26 146.155
R8353 two_stage_opamp_dummy_magic_23_0.VD4.t28 two_stage_opamp_dummy_magic_23_0.VD4.t32 146.155
R8354 two_stage_opamp_dummy_magic_23_0.VD4.t14 two_stage_opamp_dummy_magic_23_0.VD4.t28 146.155
R8355 two_stage_opamp_dummy_magic_23_0.VD4.n11 two_stage_opamp_dummy_magic_23_0.VD4.t12 76.2576
R8356 two_stage_opamp_dummy_magic_23_0.VD4.n12 two_stage_opamp_dummy_magic_23_0.VD4.t15 76.2576
R8357 two_stage_opamp_dummy_magic_23_0.VD4.n7 two_stage_opamp_dummy_magic_23_0.VD4.n6 71.513
R8358 two_stage_opamp_dummy_magic_23_0.VD4.n9 two_stage_opamp_dummy_magic_23_0.VD4.n8 71.513
R8359 two_stage_opamp_dummy_magic_23_0.VD4.n1 two_stage_opamp_dummy_magic_23_0.VD4.n0 71.513
R8360 two_stage_opamp_dummy_magic_23_0.VD4.n3 two_stage_opamp_dummy_magic_23_0.VD4.n2 71.513
R8361 two_stage_opamp_dummy_magic_23_0.VD4.n5 two_stage_opamp_dummy_magic_23_0.VD4.n4 71.513
R8362 two_stage_opamp_dummy_magic_23_0.VD4.n18 two_stage_opamp_dummy_magic_23_0.VD4.n17 66.0338
R8363 two_stage_opamp_dummy_magic_23_0.VD4.n21 two_stage_opamp_dummy_magic_23_0.VD4.n20 66.0338
R8364 two_stage_opamp_dummy_magic_23_0.VD4.n24 two_stage_opamp_dummy_magic_23_0.VD4.n23 66.0338
R8365 two_stage_opamp_dummy_magic_23_0.VD4.n28 two_stage_opamp_dummy_magic_23_0.VD4.n27 66.0338
R8366 two_stage_opamp_dummy_magic_23_0.VD4.n31 two_stage_opamp_dummy_magic_23_0.VD4.n30 66.0338
R8367 two_stage_opamp_dummy_magic_23_0.VD4.n34 two_stage_opamp_dummy_magic_23_0.VD4.n33 66.0338
R8368 two_stage_opamp_dummy_magic_23_0.VD4.n6 two_stage_opamp_dummy_magic_23_0.VD4.t31 11.2576
R8369 two_stage_opamp_dummy_magic_23_0.VD4.n6 two_stage_opamp_dummy_magic_23_0.VD4.t35 11.2576
R8370 two_stage_opamp_dummy_magic_23_0.VD4.n8 two_stage_opamp_dummy_magic_23_0.VD4.t21 11.2576
R8371 two_stage_opamp_dummy_magic_23_0.VD4.n8 two_stage_opamp_dummy_magic_23_0.VD4.t25 11.2576
R8372 two_stage_opamp_dummy_magic_23_0.VD4.n17 two_stage_opamp_dummy_magic_23_0.VD4.t2 11.2576
R8373 two_stage_opamp_dummy_magic_23_0.VD4.n17 two_stage_opamp_dummy_magic_23_0.VD4.t16 11.2576
R8374 two_stage_opamp_dummy_magic_23_0.VD4.n20 two_stage_opamp_dummy_magic_23_0.VD4.t8 11.2576
R8375 two_stage_opamp_dummy_magic_23_0.VD4.n20 two_stage_opamp_dummy_magic_23_0.VD4.t1 11.2576
R8376 two_stage_opamp_dummy_magic_23_0.VD4.n23 two_stage_opamp_dummy_magic_23_0.VD4.t6 11.2576
R8377 two_stage_opamp_dummy_magic_23_0.VD4.n23 two_stage_opamp_dummy_magic_23_0.VD4.t5 11.2576
R8378 two_stage_opamp_dummy_magic_23_0.VD4.n27 two_stage_opamp_dummy_magic_23_0.VD4.t3 11.2576
R8379 two_stage_opamp_dummy_magic_23_0.VD4.n27 two_stage_opamp_dummy_magic_23_0.VD4.t4 11.2576
R8380 two_stage_opamp_dummy_magic_23_0.VD4.n30 two_stage_opamp_dummy_magic_23_0.VD4.t7 11.2576
R8381 two_stage_opamp_dummy_magic_23_0.VD4.n30 two_stage_opamp_dummy_magic_23_0.VD4.t0 11.2576
R8382 two_stage_opamp_dummy_magic_23_0.VD4.n33 two_stage_opamp_dummy_magic_23_0.VD4.t17 11.2576
R8383 two_stage_opamp_dummy_magic_23_0.VD4.n33 two_stage_opamp_dummy_magic_23_0.VD4.t9 11.2576
R8384 two_stage_opamp_dummy_magic_23_0.VD4.n0 two_stage_opamp_dummy_magic_23_0.VD4.t33 11.2576
R8385 two_stage_opamp_dummy_magic_23_0.VD4.n0 two_stage_opamp_dummy_magic_23_0.VD4.t29 11.2576
R8386 two_stage_opamp_dummy_magic_23_0.VD4.n2 two_stage_opamp_dummy_magic_23_0.VD4.t23 11.2576
R8387 two_stage_opamp_dummy_magic_23_0.VD4.n2 two_stage_opamp_dummy_magic_23_0.VD4.t27 11.2576
R8388 two_stage_opamp_dummy_magic_23_0.VD4.n4 two_stage_opamp_dummy_magic_23_0.VD4.t37 11.2576
R8389 two_stage_opamp_dummy_magic_23_0.VD4.n4 two_stage_opamp_dummy_magic_23_0.VD4.t19 11.2576
R8390 two_stage_opamp_dummy_magic_23_0.VD4 two_stage_opamp_dummy_magic_23_0.VD4.n35 8.59425
R8391 two_stage_opamp_dummy_magic_23_0.VD4.n10 two_stage_opamp_dummy_magic_23_0.VD4.n9 6.10467
R8392 two_stage_opamp_dummy_magic_23_0.VD4.n34 two_stage_opamp_dummy_magic_23_0.VD4.n32 5.91717
R8393 two_stage_opamp_dummy_magic_23_0.VD4.n19 two_stage_opamp_dummy_magic_23_0.VD4.n18 5.91717
R8394 two_stage_opamp_dummy_magic_23_0.VD4.n22 two_stage_opamp_dummy_magic_23_0.VD4.n18 5.91717
R8395 two_stage_opamp_dummy_magic_23_0.VD4.n14 two_stage_opamp_dummy_magic_23_0.VD4.n13 5.47967
R8396 two_stage_opamp_dummy_magic_23_0.VD4 two_stage_opamp_dummy_magic_23_0.VD4.n14 5.3755
R8397 two_stage_opamp_dummy_magic_23_0.VD4.n22 two_stage_opamp_dummy_magic_23_0.VD4.n21 5.29217
R8398 two_stage_opamp_dummy_magic_23_0.VD4.n21 two_stage_opamp_dummy_magic_23_0.VD4.n19 5.29217
R8399 two_stage_opamp_dummy_magic_23_0.VD4.n25 two_stage_opamp_dummy_magic_23_0.VD4.n24 5.29217
R8400 two_stage_opamp_dummy_magic_23_0.VD4.n24 two_stage_opamp_dummy_magic_23_0.VD4.n16 5.29217
R8401 two_stage_opamp_dummy_magic_23_0.VD4.n28 two_stage_opamp_dummy_magic_23_0.VD4.n26 5.29217
R8402 two_stage_opamp_dummy_magic_23_0.VD4.n29 two_stage_opamp_dummy_magic_23_0.VD4.n28 5.29217
R8403 two_stage_opamp_dummy_magic_23_0.VD4.n31 two_stage_opamp_dummy_magic_23_0.VD4.n15 5.29217
R8404 two_stage_opamp_dummy_magic_23_0.VD4.n32 two_stage_opamp_dummy_magic_23_0.VD4.n31 5.29217
R8405 two_stage_opamp_dummy_magic_23_0.VD4.n35 two_stage_opamp_dummy_magic_23_0.VD4.n34 5.29217
R8406 two_stage_opamp_dummy_magic_23_0.VD4.n13 two_stage_opamp_dummy_magic_23_0.VD4.n12 1.03383
R8407 two_stage_opamp_dummy_magic_23_0.VD4.n11 two_stage_opamp_dummy_magic_23_0.VD4.n10 1.03383
R8408 two_stage_opamp_dummy_magic_23_0.VD4.n32 two_stage_opamp_dummy_magic_23_0.VD4.n29 0.6255
R8409 two_stage_opamp_dummy_magic_23_0.VD4.n29 two_stage_opamp_dummy_magic_23_0.VD4.n16 0.6255
R8410 two_stage_opamp_dummy_magic_23_0.VD4.n19 two_stage_opamp_dummy_magic_23_0.VD4.n16 0.6255
R8411 two_stage_opamp_dummy_magic_23_0.VD4.n25 two_stage_opamp_dummy_magic_23_0.VD4.n22 0.6255
R8412 two_stage_opamp_dummy_magic_23_0.VD4.n26 two_stage_opamp_dummy_magic_23_0.VD4.n25 0.6255
R8413 two_stage_opamp_dummy_magic_23_0.VD4.n26 two_stage_opamp_dummy_magic_23_0.VD4.n15 0.6255
R8414 two_stage_opamp_dummy_magic_23_0.VD4.n35 two_stage_opamp_dummy_magic_23_0.VD4.n15 0.6255
R8415 two_stage_opamp_dummy_magic_23_0.VD4.n5 two_stage_opamp_dummy_magic_23_0.VD4.n3 0.6255
R8416 two_stage_opamp_dummy_magic_23_0.VD4.n3 two_stage_opamp_dummy_magic_23_0.VD4.n1 0.6255
R8417 two_stage_opamp_dummy_magic_23_0.VD4.n14 two_stage_opamp_dummy_magic_23_0.VD4.n1 0.6255
R8418 two_stage_opamp_dummy_magic_23_0.VD4.n9 two_stage_opamp_dummy_magic_23_0.VD4.n7 0.6255
R8419 two_stage_opamp_dummy_magic_23_0.VD4.n7 two_stage_opamp_dummy_magic_23_0.VD4.n5 0.6255
R8420 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n0 344.837
R8421 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n1 344.274
R8422 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n3 292.5
R8423 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n22 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t4 122.754
R8424 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n7 118.861
R8425 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n9 118.861
R8426 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n13 118.861
R8427 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n17 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n16 118.861
R8428 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n20 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n19 118.861
R8429 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n2 52.3363
R8430 bgr_11_0.V_CMFB_S1 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n4 52.1563
R8431 bgr_11_0.V_CMFB_S1 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n22 47.5943
R8432 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t1 39.4005
R8433 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t5 39.4005
R8434 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t0 39.4005
R8435 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t3 39.4005
R8436 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t6 39.4005
R8437 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t2 39.4005
R8438 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t9 19.7005
R8439 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t13 19.7005
R8440 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t8 19.7005
R8441 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t15 19.7005
R8442 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t10 19.7005
R8443 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t14 19.7005
R8444 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t11 19.7005
R8445 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t16 19.7005
R8446 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n19 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t12 19.7005
R8447 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n19 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t7 19.7005
R8448 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n22 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n21 6.2505
R8449 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n8 5.60467
R8450 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n20 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n18 5.54217
R8451 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n6 5.54217
R8452 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n10 5.04217
R8453 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n12 5.04217
R8454 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n17 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n5 5.04217
R8455 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n21 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n20 5.04217
R8456 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n6 4.97967
R8457 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n14 4.97967
R8458 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n18 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n17 4.97967
R8459 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n18 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n15 0.563
R8460 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n6 0.563
R8461 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n11 0.563
R8462 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n5 0.563
R8463 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n21 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n5 0.563
R8464 two_stage_opamp_dummy_magic_23_0.Vb2_2.n2 two_stage_opamp_dummy_magic_23_0.Vb2_2.t3 661.375
R8465 two_stage_opamp_dummy_magic_23_0.Vb2_2.n4 two_stage_opamp_dummy_magic_23_0.Vb2_2.t0 661.375
R8466 two_stage_opamp_dummy_magic_23_0.Vb2_2.t4 two_stage_opamp_dummy_magic_23_0.Vb2_2.n0 213.131
R8467 two_stage_opamp_dummy_magic_23_0.Vb2_2.n3 two_stage_opamp_dummy_magic_23_0.Vb2_2.t1 213.131
R8468 two_stage_opamp_dummy_magic_23_0.Vb2_2.n6 two_stage_opamp_dummy_magic_23_0.Vb2_2.n1 154.983
R8469 two_stage_opamp_dummy_magic_23_0.Vb2_2.t7 two_stage_opamp_dummy_magic_23_0.Vb2_2.t4 146.155
R8470 two_stage_opamp_dummy_magic_23_0.Vb2_2.t1 two_stage_opamp_dummy_magic_23_0.Vb2_2.t7 146.155
R8471 two_stage_opamp_dummy_magic_23_0.Vb2_2.t5 two_stage_opamp_dummy_magic_23_0.Vb2_2.n0 76.2576
R8472 two_stage_opamp_dummy_magic_23_0.Vb2_2.n3 two_stage_opamp_dummy_magic_23_0.Vb2_2.t2 76.2576
R8473 two_stage_opamp_dummy_magic_23_0.Vb2_2.n7 two_stage_opamp_dummy_magic_23_0.Vb2_2.n6 66.4421
R8474 two_stage_opamp_dummy_magic_23_0.Vb2_2.n1 two_stage_opamp_dummy_magic_23_0.Vb2_2.t6 21.8894
R8475 two_stage_opamp_dummy_magic_23_0.Vb2_2.n1 two_stage_opamp_dummy_magic_23_0.Vb2_2.t9 21.8894
R8476 two_stage_opamp_dummy_magic_23_0.Vb2_2.t5 two_stage_opamp_dummy_magic_23_0.Vb2_2.n7 11.2576
R8477 two_stage_opamp_dummy_magic_23_0.Vb2_2.n7 two_stage_opamp_dummy_magic_23_0.Vb2_2.t8 11.2576
R8478 two_stage_opamp_dummy_magic_23_0.Vb2_2.n5 two_stage_opamp_dummy_magic_23_0.Vb2_2.n4 5.1255
R8479 two_stage_opamp_dummy_magic_23_0.Vb2_2.n6 two_stage_opamp_dummy_magic_23_0.Vb2_2.n5 4.92067
R8480 two_stage_opamp_dummy_magic_23_0.Vb2_2.n5 two_stage_opamp_dummy_magic_23_0.Vb2_2.n2 4.7505
R8481 two_stage_opamp_dummy_magic_23_0.Vb2_2.n4 two_stage_opamp_dummy_magic_23_0.Vb2_2.n3 1.888
R8482 two_stage_opamp_dummy_magic_23_0.Vb2_2.n2 two_stage_opamp_dummy_magic_23_0.Vb2_2.n0 1.888
R8483 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t18 739.067
R8484 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n3 724.936
R8485 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t7 688.859
R8486 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n1 530.201
R8487 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n5 530.201
R8488 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n7 530.201
R8489 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n10 514.134
R8490 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n8 361.5
R8491 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n12 214.056
R8492 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t14 208.868
R8493 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t9 208.868
R8494 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t15 208.868
R8495 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t8 208.868
R8496 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t16 208.868
R8497 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t12 208.868
R8498 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t19 208.868
R8499 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t13 208.868
R8500 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t20 208.868
R8501 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n0 176.733
R8502 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n2 176.733
R8503 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n4 176.733
R8504 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n6 176.733
R8505 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t17 174.726
R8506 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t11 174.726
R8507 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t21 174.726
R8508 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t10 174.726
R8509 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n14 173.591
R8510 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n17 169.216
R8511 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n15 169.216
R8512 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n9 128.534
R8513 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n11 128.534
R8514 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t0 125.736
R8515 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n19 51.4693
R8516 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t3 13.1338
R8517 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t1 13.1338
R8518 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t4 13.1338
R8519 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t5 13.1338
R8520 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t2 13.1338
R8521 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t6 13.1338
R8522 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n18 10.0317
R8523 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n16 4.3755
R8524 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n13 3.03175
R8525 bgr_11_0.V_p_2.n6 bgr_11_0.V_p_2.n1 229.562
R8526 bgr_11_0.V_p_2.n1 bgr_11_0.V_p_2.n5 228.939
R8527 bgr_11_0.V_p_2.n1 bgr_11_0.V_p_2.n4 228.939
R8528 bgr_11_0.V_p_2.n0 bgr_11_0.V_p_2.n3 228.939
R8529 bgr_11_0.V_p_2.n0 bgr_11_0.V_p_2.n2 228.939
R8530 bgr_11_0.V_p_2.n0 bgr_11_0.V_p_2.t9 98.7279
R8531 bgr_11_0.V_p_2.n5 bgr_11_0.V_p_2.t10 48.0005
R8532 bgr_11_0.V_p_2.n5 bgr_11_0.V_p_2.t4 48.0005
R8533 bgr_11_0.V_p_2.n4 bgr_11_0.V_p_2.t5 48.0005
R8534 bgr_11_0.V_p_2.n4 bgr_11_0.V_p_2.t0 48.0005
R8535 bgr_11_0.V_p_2.n3 bgr_11_0.V_p_2.t1 48.0005
R8536 bgr_11_0.V_p_2.n3 bgr_11_0.V_p_2.t3 48.0005
R8537 bgr_11_0.V_p_2.n2 bgr_11_0.V_p_2.t6 48.0005
R8538 bgr_11_0.V_p_2.n2 bgr_11_0.V_p_2.t8 48.0005
R8539 bgr_11_0.V_p_2.t7 bgr_11_0.V_p_2.n6 48.0005
R8540 bgr_11_0.V_p_2.n6 bgr_11_0.V_p_2.t2 48.0005
R8541 bgr_11_0.V_p_2.n1 bgr_11_0.V_p_2.n0 1.8755
R8542 a_6470_23450.t0 a_6470_23450.t1 178.133
R8543 two_stage_opamp_dummy_magic_23_0.V_err_p.n4 two_stage_opamp_dummy_magic_23_0.V_err_p.n3 594.301
R8544 two_stage_opamp_dummy_magic_23_0.V_err_p.n0 two_stage_opamp_dummy_magic_23_0.V_err_p.n23 594.301
R8545 two_stage_opamp_dummy_magic_23_0.V_err_p.n6 two_stage_opamp_dummy_magic_23_0.V_err_p.n5 594.301
R8546 two_stage_opamp_dummy_magic_23_0.V_err_p.n9 two_stage_opamp_dummy_magic_23_0.V_err_p.n8 594.301
R8547 two_stage_opamp_dummy_magic_23_0.V_err_p.n12 two_stage_opamp_dummy_magic_23_0.V_err_p.n11 594.301
R8548 two_stage_opamp_dummy_magic_23_0.V_err_p.n15 two_stage_opamp_dummy_magic_23_0.V_err_p.n14 594.301
R8549 two_stage_opamp_dummy_magic_23_0.V_err_p.n19 two_stage_opamp_dummy_magic_23_0.V_err_p.n18 594.301
R8550 two_stage_opamp_dummy_magic_23_0.V_err_p.n26 two_stage_opamp_dummy_magic_23_0.V_err_p.n25 594.301
R8551 two_stage_opamp_dummy_magic_23_0.V_err_p.n30 two_stage_opamp_dummy_magic_23_0.V_err_p.n29 594.301
R8552 two_stage_opamp_dummy_magic_23_0.V_err_p.n33 two_stage_opamp_dummy_magic_23_0.V_err_p.n32 594.301
R8553 two_stage_opamp_dummy_magic_23_0.V_err_p.n36 two_stage_opamp_dummy_magic_23_0.V_err_p.n35 594.301
R8554 two_stage_opamp_dummy_magic_23_0.V_err_p.n3 two_stage_opamp_dummy_magic_23_0.V_err_p.t19 78.8005
R8555 two_stage_opamp_dummy_magic_23_0.V_err_p.n3 two_stage_opamp_dummy_magic_23_0.V_err_p.t11 78.8005
R8556 two_stage_opamp_dummy_magic_23_0.V_err_p.n23 two_stage_opamp_dummy_magic_23_0.V_err_p.t4 78.8005
R8557 two_stage_opamp_dummy_magic_23_0.V_err_p.n23 two_stage_opamp_dummy_magic_23_0.V_err_p.t9 78.8005
R8558 two_stage_opamp_dummy_magic_23_0.V_err_p.n5 two_stage_opamp_dummy_magic_23_0.V_err_p.t13 78.8005
R8559 two_stage_opamp_dummy_magic_23_0.V_err_p.n5 two_stage_opamp_dummy_magic_23_0.V_err_p.t20 78.8005
R8560 two_stage_opamp_dummy_magic_23_0.V_err_p.n8 two_stage_opamp_dummy_magic_23_0.V_err_p.t15 78.8005
R8561 two_stage_opamp_dummy_magic_23_0.V_err_p.n8 two_stage_opamp_dummy_magic_23_0.V_err_p.t0 78.8005
R8562 two_stage_opamp_dummy_magic_23_0.V_err_p.n11 two_stage_opamp_dummy_magic_23_0.V_err_p.t2 78.8005
R8563 two_stage_opamp_dummy_magic_23_0.V_err_p.n11 two_stage_opamp_dummy_magic_23_0.V_err_p.t14 78.8005
R8564 two_stage_opamp_dummy_magic_23_0.V_err_p.n14 two_stage_opamp_dummy_magic_23_0.V_err_p.t16 78.8005
R8565 two_stage_opamp_dummy_magic_23_0.V_err_p.n14 two_stage_opamp_dummy_magic_23_0.V_err_p.t21 78.8005
R8566 two_stage_opamp_dummy_magic_23_0.V_err_p.n18 two_stage_opamp_dummy_magic_23_0.V_err_p.t1 78.8005
R8567 two_stage_opamp_dummy_magic_23_0.V_err_p.n18 two_stage_opamp_dummy_magic_23_0.V_err_p.t17 78.8005
R8568 two_stage_opamp_dummy_magic_23_0.V_err_p.n25 two_stage_opamp_dummy_magic_23_0.V_err_p.t3 78.8005
R8569 two_stage_opamp_dummy_magic_23_0.V_err_p.n25 two_stage_opamp_dummy_magic_23_0.V_err_p.t8 78.8005
R8570 two_stage_opamp_dummy_magic_23_0.V_err_p.n29 two_stage_opamp_dummy_magic_23_0.V_err_p.t5 78.8005
R8571 two_stage_opamp_dummy_magic_23_0.V_err_p.n29 two_stage_opamp_dummy_magic_23_0.V_err_p.t7 78.8005
R8572 two_stage_opamp_dummy_magic_23_0.V_err_p.n32 two_stage_opamp_dummy_magic_23_0.V_err_p.t10 78.8005
R8573 two_stage_opamp_dummy_magic_23_0.V_err_p.n32 two_stage_opamp_dummy_magic_23_0.V_err_p.t6 78.8005
R8574 two_stage_opamp_dummy_magic_23_0.V_err_p.t12 two_stage_opamp_dummy_magic_23_0.V_err_p.n36 78.8005
R8575 two_stage_opamp_dummy_magic_23_0.V_err_p.n36 two_stage_opamp_dummy_magic_23_0.V_err_p.t18 78.8005
R8576 two_stage_opamp_dummy_magic_23_0.V_err_p.n35 two_stage_opamp_dummy_magic_23_0.V_err_p.n1 6.10467
R8577 two_stage_opamp_dummy_magic_23_0.V_err_p.n24 two_stage_opamp_dummy_magic_23_0.V_err_p.n4 6.10467
R8578 two_stage_opamp_dummy_magic_23_0.V_err_p.n22 two_stage_opamp_dummy_magic_23_0.V_err_p.n4 5.91717
R8579 two_stage_opamp_dummy_magic_23_0.V_err_p.n35 two_stage_opamp_dummy_magic_23_0.V_err_p.n34 5.91717
R8580 two_stage_opamp_dummy_magic_23_0.V_err_p.n10 two_stage_opamp_dummy_magic_23_0.V_err_p.n9 5.41717
R8581 two_stage_opamp_dummy_magic_23_0.V_err_p.n13 two_stage_opamp_dummy_magic_23_0.V_err_p.n9 5.22967
R8582 two_stage_opamp_dummy_magic_23_0.V_err_p.n17 two_stage_opamp_dummy_magic_23_0.V_err_p.n6 5.22967
R8583 two_stage_opamp_dummy_magic_23_0.V_err_p.n21 two_stage_opamp_dummy_magic_23_0.V_err_p.n20 5.063
R8584 two_stage_opamp_dummy_magic_23_0.V_err_p.n12 two_stage_opamp_dummy_magic_23_0.V_err_p.n10 4.85467
R8585 two_stage_opamp_dummy_magic_23_0.V_err_p.n15 two_stage_opamp_dummy_magic_23_0.V_err_p.n7 4.85467
R8586 two_stage_opamp_dummy_magic_23_0.V_err_p.n20 two_stage_opamp_dummy_magic_23_0.V_err_p.n19 4.85467
R8587 two_stage_opamp_dummy_magic_23_0.V_err_p.n24 two_stage_opamp_dummy_magic_23_0.V_err_p.n0 4.85467
R8588 two_stage_opamp_dummy_magic_23_0.V_err_p.n27 two_stage_opamp_dummy_magic_23_0.V_err_p.n26 4.85467
R8589 two_stage_opamp_dummy_magic_23_0.V_err_p.n30 two_stage_opamp_dummy_magic_23_0.V_err_p.n28 4.85467
R8590 two_stage_opamp_dummy_magic_23_0.V_err_p.n33 two_stage_opamp_dummy_magic_23_0.V_err_p.n1 4.85467
R8591 two_stage_opamp_dummy_magic_23_0.V_err_p.n13 two_stage_opamp_dummy_magic_23_0.V_err_p.n12 4.66717
R8592 two_stage_opamp_dummy_magic_23_0.V_err_p.n16 two_stage_opamp_dummy_magic_23_0.V_err_p.n15 4.66717
R8593 two_stage_opamp_dummy_magic_23_0.V_err_p.n19 two_stage_opamp_dummy_magic_23_0.V_err_p.n17 4.66717
R8594 two_stage_opamp_dummy_magic_23_0.V_err_p.n26 two_stage_opamp_dummy_magic_23_0.V_err_p.n2 4.66717
R8595 two_stage_opamp_dummy_magic_23_0.V_err_p.n31 two_stage_opamp_dummy_magic_23_0.V_err_p.n30 4.66717
R8596 two_stage_opamp_dummy_magic_23_0.V_err_p.n34 two_stage_opamp_dummy_magic_23_0.V_err_p.n33 4.66717
R8597 two_stage_opamp_dummy_magic_23_0.V_err_p.n0 two_stage_opamp_dummy_magic_23_0.V_err_p.n22 4.5005
R8598 two_stage_opamp_dummy_magic_23_0.V_err_p.n28 two_stage_opamp_dummy_magic_23_0.V_err_p.n1 1.2505
R8599 two_stage_opamp_dummy_magic_23_0.V_err_p.n28 two_stage_opamp_dummy_magic_23_0.V_err_p.n27 1.2505
R8600 two_stage_opamp_dummy_magic_23_0.V_err_p.n27 two_stage_opamp_dummy_magic_23_0.V_err_p.n24 1.2505
R8601 two_stage_opamp_dummy_magic_23_0.V_err_p.n22 two_stage_opamp_dummy_magic_23_0.V_err_p.n2 1.2505
R8602 two_stage_opamp_dummy_magic_23_0.V_err_p.n31 two_stage_opamp_dummy_magic_23_0.V_err_p.n2 1.2505
R8603 two_stage_opamp_dummy_magic_23_0.V_err_p.n34 two_stage_opamp_dummy_magic_23_0.V_err_p.n31 1.2505
R8604 two_stage_opamp_dummy_magic_23_0.V_err_p.n0 two_stage_opamp_dummy_magic_23_0.V_err_p.n21 1.11508
R8605 two_stage_opamp_dummy_magic_23_0.V_err_p.n20 two_stage_opamp_dummy_magic_23_0.V_err_p.n7 0.563
R8606 two_stage_opamp_dummy_magic_23_0.V_err_p.n10 two_stage_opamp_dummy_magic_23_0.V_err_p.n7 0.563
R8607 two_stage_opamp_dummy_magic_23_0.V_err_p.n16 two_stage_opamp_dummy_magic_23_0.V_err_p.n13 0.563
R8608 two_stage_opamp_dummy_magic_23_0.V_err_p.n17 two_stage_opamp_dummy_magic_23_0.V_err_p.n16 0.563
R8609 two_stage_opamp_dummy_magic_23_0.V_err_p.n21 two_stage_opamp_dummy_magic_23_0.V_err_p.n6 0.333833
R8610 two_stage_opamp_dummy_magic_23_0.err_amp_out.n6 two_stage_opamp_dummy_magic_23_0.err_amp_out.t12 840.595
R8611 two_stage_opamp_dummy_magic_23_0.err_amp_out.n12 two_stage_opamp_dummy_magic_23_0.err_amp_out.n10 601.051
R8612 two_stage_opamp_dummy_magic_23_0.err_amp_out two_stage_opamp_dummy_magic_23_0.err_amp_out.n13 599.801
R8613 two_stage_opamp_dummy_magic_23_0.err_amp_out.n12 two_stage_opamp_dummy_magic_23_0.err_amp_out.n11 599.801
R8614 two_stage_opamp_dummy_magic_23_0.err_amp_out.n2 two_stage_opamp_dummy_magic_23_0.err_amp_out.n1 194.3
R8615 two_stage_opamp_dummy_magic_23_0.err_amp_out.n4 two_stage_opamp_dummy_magic_23_0.err_amp_out.n3 194.3
R8616 two_stage_opamp_dummy_magic_23_0.err_amp_out.n8 two_stage_opamp_dummy_magic_23_0.err_amp_out.n7 194.3
R8617 two_stage_opamp_dummy_magic_23_0.err_amp_out.n13 two_stage_opamp_dummy_magic_23_0.err_amp_out.t3 78.8005
R8618 two_stage_opamp_dummy_magic_23_0.err_amp_out.n13 two_stage_opamp_dummy_magic_23_0.err_amp_out.t5 78.8005
R8619 two_stage_opamp_dummy_magic_23_0.err_amp_out.n10 two_stage_opamp_dummy_magic_23_0.err_amp_out.t9 78.8005
R8620 two_stage_opamp_dummy_magic_23_0.err_amp_out.n10 two_stage_opamp_dummy_magic_23_0.err_amp_out.t2 78.8005
R8621 two_stage_opamp_dummy_magic_23_0.err_amp_out.n11 two_stage_opamp_dummy_magic_23_0.err_amp_out.t4 78.8005
R8622 two_stage_opamp_dummy_magic_23_0.err_amp_out.n11 two_stage_opamp_dummy_magic_23_0.err_amp_out.t6 78.8005
R8623 two_stage_opamp_dummy_magic_23_0.err_amp_out.n1 two_stage_opamp_dummy_magic_23_0.err_amp_out.t0 48.0005
R8624 two_stage_opamp_dummy_magic_23_0.err_amp_out.n1 two_stage_opamp_dummy_magic_23_0.err_amp_out.t10 48.0005
R8625 two_stage_opamp_dummy_magic_23_0.err_amp_out.n3 two_stage_opamp_dummy_magic_23_0.err_amp_out.t8 48.0005
R8626 two_stage_opamp_dummy_magic_23_0.err_amp_out.n3 two_stage_opamp_dummy_magic_23_0.err_amp_out.t11 48.0005
R8627 two_stage_opamp_dummy_magic_23_0.err_amp_out.n7 two_stage_opamp_dummy_magic_23_0.err_amp_out.t1 48.0005
R8628 two_stage_opamp_dummy_magic_23_0.err_amp_out.n7 two_stage_opamp_dummy_magic_23_0.err_amp_out.t7 48.0005
R8629 two_stage_opamp_dummy_magic_23_0.err_amp_out.n5 two_stage_opamp_dummy_magic_23_0.err_amp_out.n2 6.20883
R8630 two_stage_opamp_dummy_magic_23_0.err_amp_out.n2 two_stage_opamp_dummy_magic_23_0.err_amp_out.n0 6.20883
R8631 two_stage_opamp_dummy_magic_23_0.err_amp_out.n4 two_stage_opamp_dummy_magic_23_0.err_amp_out.n0 4.95883
R8632 two_stage_opamp_dummy_magic_23_0.err_amp_out.n5 two_stage_opamp_dummy_magic_23_0.err_amp_out.n4 4.95883
R8633 two_stage_opamp_dummy_magic_23_0.err_amp_out.n9 two_stage_opamp_dummy_magic_23_0.err_amp_out.n8 4.95883
R8634 two_stage_opamp_dummy_magic_23_0.err_amp_out.n8 two_stage_opamp_dummy_magic_23_0.err_amp_out.n6 4.95883
R8635 two_stage_opamp_dummy_magic_23_0.err_amp_out.n6 two_stage_opamp_dummy_magic_23_0.err_amp_out.n5 1.2505
R8636 two_stage_opamp_dummy_magic_23_0.err_amp_out.n9 two_stage_opamp_dummy_magic_23_0.err_amp_out.n0 1.2505
R8637 two_stage_opamp_dummy_magic_23_0.err_amp_out two_stage_opamp_dummy_magic_23_0.err_amp_out.n12 1.2505
R8638 two_stage_opamp_dummy_magic_23_0.err_amp_out two_stage_opamp_dummy_magic_23_0.err_amp_out.n9 1.063
R8639 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n0 144.827
R8640 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n1 134.577
R8641 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t0 120.504
R8642 bgr_11_0.V_CMFB_S4 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n20 40.4693
R8643 bgr_11_0.V_CMFB_S4 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n2 37.563
R8644 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n5 24.288
R8645 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n7 24.288
R8646 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n11 24.288
R8647 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n14 24.288
R8648 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n17 24.288
R8649 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t3 24.0005
R8650 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t2 24.0005
R8651 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t14 24.0005
R8652 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t1 24.0005
R8653 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t4 8.0005
R8654 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t8 8.0005
R8655 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t13 8.0005
R8656 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t11 8.0005
R8657 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t6 8.0005
R8658 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t10 8.0005
R8659 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t5 8.0005
R8660 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t9 8.0005
R8661 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t12 8.0005
R8662 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t7 8.0005
R8663 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n19 6.0005
R8664 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n16 5.7505
R8665 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n4 5.7505
R8666 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n6 5.7505
R8667 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n8 5.188
R8668 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n4 5.188
R8669 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n10 5.188
R8670 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n12 5.188
R8671 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n3 5.188
R8672 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n15 5.188
R8673 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n18 5.188
R8674 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n13 0.563
R8675 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n4 0.563
R8676 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n9 0.563
R8677 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n3 0.563
R8678 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n3 0.563
R8679 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n15 594.301
R8680 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n16 594.301
R8681 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n19 594.301
R8682 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t18 289.2
R8683 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t7 289.2
R8684 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n3 194.3
R8685 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n24 194.3
R8686 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n26 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n1 194.3
R8687 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n5 176.733
R8688 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n6 176.733
R8689 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n9 176.733
R8690 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n10 176.733
R8691 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n11 176.733
R8692 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n1 161.3
R8693 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n14 161.3
R8694 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t3 112.468
R8695 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t11 112.468
R8696 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t20 112.468
R8697 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t17 112.468
R8698 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t9 112.468
R8699 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t19 112.468
R8700 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t21 112.468
R8701 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t5 112.468
R8702 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t16 78.8005
R8703 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t1 78.8005
R8704 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t0 78.8005
R8705 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t2 78.8005
R8706 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t15 78.8005
R8707 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t13 78.8005
R8708 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t14 48.0005
R8709 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t8 48.0005
R8710 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n24 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t10 48.0005
R8711 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n24 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t4 48.0005
R8712 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t12 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n26 48.0005
R8713 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n26 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t6 48.0005
R8714 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n13 45.5227
R8715 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n7 45.5227
R8716 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n8 45.5227
R8717 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n12 45.5227
R8718 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n25 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n2 6.39633
R8719 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n22 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n0 6.39633
R8720 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n25 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n4 6.39633
R8721 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n20 6.10467
R8722 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n17 6.10467
R8723 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n23 5.97967
R8724 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n18 5.91717
R8725 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n17 5.91717
R8726 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n25 5.14633
R8727 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n21 4.85467
R8728 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n22 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n4 4.72967
R8729 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n23 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n1 4.72967
R8730 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n0 4.66717
R8731 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n23 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n22 1.2505
R8732 bgr_11_0.Vin+.n3 bgr_11_0.Vin+.n2 526.183
R8733 bgr_11_0.Vin+.n1 bgr_11_0.Vin+.n0 514.134
R8734 bgr_11_0.Vin+.n0 bgr_11_0.Vin+.t8 303.259
R8735 bgr_11_0.Vin+.n5 bgr_11_0.Vin+.n3 227.169
R8736 bgr_11_0.Vin+.n0 bgr_11_0.Vin+.t9 174.726
R8737 bgr_11_0.Vin+.n1 bgr_11_0.Vin+.t6 174.726
R8738 bgr_11_0.Vin+.n2 bgr_11_0.Vin+.t10 174.726
R8739 bgr_11_0.Vin+.n7 bgr_11_0.Vin+.n6 168.435
R8740 bgr_11_0.Vin+.n5 bgr_11_0.Vin+.n4 168.435
R8741 bgr_11_0.Vin+.t0 bgr_11_0.Vin+.n8 158.989
R8742 bgr_11_0.Vin+.n2 bgr_11_0.Vin+.n1 128.534
R8743 bgr_11_0.Vin+.n8 bgr_11_0.Vin+.t1 119.067
R8744 bgr_11_0.Vin+.n3 bgr_11_0.Vin+.t7 96.4005
R8745 bgr_11_0.Vin+.n8 bgr_11_0.Vin+.n7 35.0317
R8746 bgr_11_0.Vin+.n6 bgr_11_0.Vin+.t3 13.1338
R8747 bgr_11_0.Vin+.n6 bgr_11_0.Vin+.t2 13.1338
R8748 bgr_11_0.Vin+.n4 bgr_11_0.Vin+.t5 13.1338
R8749 bgr_11_0.Vin+.n4 bgr_11_0.Vin+.t4 13.1338
R8750 bgr_11_0.Vin+.n7 bgr_11_0.Vin+.n5 2.1255
R8751 a_7460_6300.n2 a_7460_6300.n1 594.301
R8752 a_7460_6300.n5 a_7460_6300.n4 594.301
R8753 a_7460_6300.n26 a_7460_6300.n25 594.301
R8754 a_7460_6300.n29 a_7460_6300.n28 594.301
R8755 a_7460_6300.n8 a_7460_6300.n7 594.301
R8756 a_7460_6300.n10 a_7460_6300.n9 594.301
R8757 a_7460_6300.n14 a_7460_6300.n13 594.301
R8758 a_7460_6300.n16 a_7460_6300.n15 594.301
R8759 a_7460_6300.n20 a_7460_6300.n19 594.301
R8760 a_7460_6300.n33 a_7460_6300.n32 594.301
R8761 a_7460_6300.n1 a_7460_6300.t4 78.8005
R8762 a_7460_6300.n1 a_7460_6300.t7 78.8005
R8763 a_7460_6300.n4 a_7460_6300.t1 78.8005
R8764 a_7460_6300.n4 a_7460_6300.t5 78.8005
R8765 a_7460_6300.n25 a_7460_6300.t6 78.8005
R8766 a_7460_6300.n25 a_7460_6300.t2 78.8005
R8767 a_7460_6300.n28 a_7460_6300.t9 78.8005
R8768 a_7460_6300.n28 a_7460_6300.t3 78.8005
R8769 a_7460_6300.n7 a_7460_6300.t13 78.8005
R8770 a_7460_6300.n7 a_7460_6300.t11 78.8005
R8771 a_7460_6300.n9 a_7460_6300.t19 78.8005
R8772 a_7460_6300.n9 a_7460_6300.t16 78.8005
R8773 a_7460_6300.n13 a_7460_6300.t18 78.8005
R8774 a_7460_6300.n13 a_7460_6300.t14 78.8005
R8775 a_7460_6300.n15 a_7460_6300.t12 78.8005
R8776 a_7460_6300.n15 a_7460_6300.t0 78.8005
R8777 a_7460_6300.n19 a_7460_6300.t17 78.8005
R8778 a_7460_6300.n19 a_7460_6300.t15 78.8005
R8779 a_7460_6300.t10 a_7460_6300.n33 78.8005
R8780 a_7460_6300.n33 a_7460_6300.t8 78.8005
R8781 a_7460_6300.n6 a_7460_6300.n2 6.20883
R8782 a_7460_6300.n27 a_7460_6300.n26 5.91717
R8783 a_7460_6300.n3 a_7460_6300.n2 5.91717
R8784 a_7460_6300.n30 a_7460_6300.n24 5.7505
R8785 a_7460_6300.n14 a_7460_6300.n11 5.41717
R8786 a_7460_6300.n22 a_7460_6300.n10 5.41717
R8787 a_7460_6300.n17 a_7460_6300.n14 5.22967
R8788 a_7460_6300.n12 a_7460_6300.n10 5.22967
R8789 a_7460_6300.n6 a_7460_6300.n5 4.95883
R8790 a_7460_6300.n30 a_7460_6300.n29 4.95883
R8791 a_7460_6300.n32 a_7460_6300.n31 4.95883
R8792 a_7460_6300.n16 a_7460_6300.n11 4.85467
R8793 a_7460_6300.n21 a_7460_6300.n20 4.85467
R8794 a_7460_6300.n5 a_7460_6300.n3 4.66717
R8795 a_7460_6300.n32 a_7460_6300.n0 4.66717
R8796 a_7460_6300.n29 a_7460_6300.n27 4.66717
R8797 a_7460_6300.n17 a_7460_6300.n16 4.66717
R8798 a_7460_6300.n20 a_7460_6300.n18 4.66717
R8799 a_7460_6300.n12 a_7460_6300.n8 4.66717
R8800 a_7460_6300.n23 a_7460_6300.n22 4.5005
R8801 a_7460_6300.n31 a_7460_6300.n30 1.2505
R8802 a_7460_6300.n27 a_7460_6300.n0 1.2505
R8803 a_7460_6300.n3 a_7460_6300.n0 1.2505
R8804 a_7460_6300.n31 a_7460_6300.n6 1.2505
R8805 a_7460_6300.n18 a_7460_6300.n12 0.563
R8806 a_7460_6300.n18 a_7460_6300.n17 0.563
R8807 a_7460_6300.n21 a_7460_6300.n11 0.563
R8808 a_7460_6300.n22 a_7460_6300.n21 0.563
R8809 a_7460_6300.n24 a_7460_6300.n23 0.51925
R8810 a_7460_6300.n26 a_7460_6300.n24 0.446333
R8811 a_7460_6300.n23 a_7460_6300.n8 0.354667
R8812 VIN-.n0 VIN-.t9 1000.38
R8813 VIN- VIN-.n9 433.019
R8814 VIN-.n9 VIN-.t1 273.134
R8815 VIN-.n0 VIN-.t0 273.134
R8816 VIN-.n1 VIN-.t5 273.134
R8817 VIN-.n2 VIN-.t10 273.134
R8818 VIN-.n3 VIN-.t3 273.134
R8819 VIN-.n4 VIN-.t7 273.134
R8820 VIN-.n5 VIN-.t4 273.134
R8821 VIN-.n6 VIN-.t8 273.134
R8822 VIN-.n7 VIN-.t2 273.134
R8823 VIN-.n8 VIN-.t6 273.134
R8824 VIN-.n9 VIN-.n8 176.733
R8825 VIN-.n8 VIN-.n7 176.733
R8826 VIN-.n7 VIN-.n6 176.733
R8827 VIN-.n6 VIN-.n5 176.733
R8828 VIN-.n5 VIN-.n4 176.733
R8829 VIN-.n4 VIN-.n3 176.733
R8830 VIN-.n3 VIN-.n2 176.733
R8831 VIN-.n2 VIN-.n1 176.733
R8832 VIN-.n1 VIN-.n0 176.733
R8833 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n0 144.827
R8834 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n1 134.577
R8835 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t4 120.817
R8836 bgr_11_0.V_CMFB_S2 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n20 40.4693
R8837 bgr_11_0.V_CMFB_S2 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n2 37.563
R8838 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n5 24.288
R8839 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n7 24.288
R8840 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n11 24.288
R8841 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n14 24.288
R8842 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n17 24.288
R8843 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t2 24.0005
R8844 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t1 24.0005
R8845 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t0 24.0005
R8846 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t3 24.0005
R8847 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t6 8.0005
R8848 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t10 8.0005
R8849 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t5 8.0005
R8850 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t12 8.0005
R8851 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t7 8.0005
R8852 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t11 8.0005
R8853 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t8 8.0005
R8854 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t13 8.0005
R8855 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t9 8.0005
R8856 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t14 8.0005
R8857 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n19 5.96925
R8858 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n16 5.7505
R8859 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n4 5.7505
R8860 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n6 5.7505
R8861 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n8 5.188
R8862 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n4 5.188
R8863 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n10 5.188
R8864 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n12 5.188
R8865 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n3 5.188
R8866 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n15 5.188
R8867 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n18 5.188
R8868 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n13 0.563
R8869 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n4 0.563
R8870 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n9 0.563
R8871 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n3 0.563
R8872 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n3 0.563
R8873 VIN+.n0 VIN+.t3 1001.28
R8874 VIN+ VIN+.n9 433.019
R8875 VIN+.n9 VIN+.t9 273.134
R8876 VIN+.n0 VIN+.t0 273.134
R8877 VIN+.n8 VIN+.t5 273.134
R8878 VIN+.n7 VIN+.t8 273.134
R8879 VIN+.n6 VIN+.t4 273.134
R8880 VIN+.n5 VIN+.t7 273.134
R8881 VIN+.n4 VIN+.t1 273.134
R8882 VIN+.n3 VIN+.t10 273.134
R8883 VIN+.n2 VIN+.t2 273.134
R8884 VIN+.n1 VIN+.t6 273.134
R8885 VIN+.n1 VIN+.n0 176.733
R8886 VIN+.n2 VIN+.n1 176.733
R8887 VIN+.n3 VIN+.n2 176.733
R8888 VIN+.n4 VIN+.n3 176.733
R8889 VIN+.n5 VIN+.n4 176.733
R8890 VIN+.n6 VIN+.n5 176.733
R8891 VIN+.n7 VIN+.n6 176.733
R8892 VIN+.n8 VIN+.n7 176.733
R8893 VIN+.n9 VIN+.n8 176.733
R8894 a_12070_24908.t0 a_12070_24908.t1 178.133
R8895 bgr_11_0.V_CUR_REF_REG.n4 bgr_11_0.V_CUR_REF_REG.n3 526.183
R8896 bgr_11_0.V_CUR_REF_REG.n2 bgr_11_0.V_CUR_REF_REG.n1 514.134
R8897 bgr_11_0.V_CUR_REF_REG.n5 bgr_11_0.V_CUR_REF_REG.n0 360.586
R8898 bgr_11_0.V_CUR_REF_REG.n1 bgr_11_0.V_CUR_REF_REG.t5 303.259
R8899 bgr_11_0.V_CUR_REF_REG.n5 bgr_11_0.V_CUR_REF_REG.n4 210.169
R8900 bgr_11_0.V_CUR_REF_REG.n1 bgr_11_0.V_CUR_REF_REG.t3 174.726
R8901 bgr_11_0.V_CUR_REF_REG.n2 bgr_11_0.V_CUR_REF_REG.t7 174.726
R8902 bgr_11_0.V_CUR_REF_REG.n3 bgr_11_0.V_CUR_REF_REG.t4 174.726
R8903 bgr_11_0.V_CUR_REF_REG.t1 bgr_11_0.V_CUR_REF_REG.n5 153.474
R8904 bgr_11_0.V_CUR_REF_REG.n3 bgr_11_0.V_CUR_REF_REG.n2 128.534
R8905 bgr_11_0.V_CUR_REF_REG.n4 bgr_11_0.V_CUR_REF_REG.t6 96.4005
R8906 bgr_11_0.V_CUR_REF_REG.n0 bgr_11_0.V_CUR_REF_REG.t0 39.4005
R8907 bgr_11_0.V_CUR_REF_REG.n0 bgr_11_0.V_CUR_REF_REG.t2 39.4005
R8908 bgr_11_0.V_mir1.n20 bgr_11_0.V_mir1.n19 325.473
R8909 bgr_11_0.V_mir1.n13 bgr_11_0.V_mir1.n12 325.473
R8910 bgr_11_0.V_mir1.n4 bgr_11_0.V_mir1.n3 325.473
R8911 bgr_11_0.V_mir1.n16 bgr_11_0.V_mir1.t18 310.488
R8912 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.t19 310.488
R8913 bgr_11_0.V_mir1.n0 bgr_11_0.V_mir1.t17 310.488
R8914 bgr_11_0.V_mir1.n7 bgr_11_0.V_mir1.t12 278.312
R8915 bgr_11_0.V_mir1.n7 bgr_11_0.V_mir1.n6 228.939
R8916 bgr_11_0.V_mir1.n8 bgr_11_0.V_mir1.n5 224.439
R8917 bgr_11_0.V_mir1.n18 bgr_11_0.V_mir1.t4 184.097
R8918 bgr_11_0.V_mir1.n11 bgr_11_0.V_mir1.t2 184.097
R8919 bgr_11_0.V_mir1.n2 bgr_11_0.V_mir1.t0 184.097
R8920 bgr_11_0.V_mir1.n17 bgr_11_0.V_mir1.n16 167.094
R8921 bgr_11_0.V_mir1.n10 bgr_11_0.V_mir1.n9 167.094
R8922 bgr_11_0.V_mir1.n1 bgr_11_0.V_mir1.n0 167.094
R8923 bgr_11_0.V_mir1.n13 bgr_11_0.V_mir1.n11 152
R8924 bgr_11_0.V_mir1.n4 bgr_11_0.V_mir1.n2 152
R8925 bgr_11_0.V_mir1.n19 bgr_11_0.V_mir1.n18 152
R8926 bgr_11_0.V_mir1.n16 bgr_11_0.V_mir1.t20 120.501
R8927 bgr_11_0.V_mir1.n17 bgr_11_0.V_mir1.t10 120.501
R8928 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.t21 120.501
R8929 bgr_11_0.V_mir1.n10 bgr_11_0.V_mir1.t8 120.501
R8930 bgr_11_0.V_mir1.n0 bgr_11_0.V_mir1.t22 120.501
R8931 bgr_11_0.V_mir1.n1 bgr_11_0.V_mir1.t6 120.501
R8932 bgr_11_0.V_mir1.n6 bgr_11_0.V_mir1.t13 48.0005
R8933 bgr_11_0.V_mir1.n6 bgr_11_0.V_mir1.t14 48.0005
R8934 bgr_11_0.V_mir1.n5 bgr_11_0.V_mir1.t15 48.0005
R8935 bgr_11_0.V_mir1.n5 bgr_11_0.V_mir1.t16 48.0005
R8936 bgr_11_0.V_mir1.n18 bgr_11_0.V_mir1.n17 40.7027
R8937 bgr_11_0.V_mir1.n11 bgr_11_0.V_mir1.n10 40.7027
R8938 bgr_11_0.V_mir1.n2 bgr_11_0.V_mir1.n1 40.7027
R8939 bgr_11_0.V_mir1.n12 bgr_11_0.V_mir1.t3 39.4005
R8940 bgr_11_0.V_mir1.n12 bgr_11_0.V_mir1.t9 39.4005
R8941 bgr_11_0.V_mir1.n3 bgr_11_0.V_mir1.t1 39.4005
R8942 bgr_11_0.V_mir1.n3 bgr_11_0.V_mir1.t7 39.4005
R8943 bgr_11_0.V_mir1.n20 bgr_11_0.V_mir1.t5 39.4005
R8944 bgr_11_0.V_mir1.t11 bgr_11_0.V_mir1.n20 39.4005
R8945 bgr_11_0.V_mir1.n15 bgr_11_0.V_mir1.n4 15.9255
R8946 bgr_11_0.V_mir1.n19 bgr_11_0.V_mir1.n15 15.9255
R8947 bgr_11_0.V_mir1.n14 bgr_11_0.V_mir1.n13 9.3005
R8948 bgr_11_0.V_mir1.n8 bgr_11_0.V_mir1.n7 5.8755
R8949 bgr_11_0.V_mir1.n15 bgr_11_0.V_mir1.n14 4.5005
R8950 bgr_11_0.V_mir1.n14 bgr_11_0.V_mir1.n8 0.78175
R8951 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t3 661.375
R8952 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t0 661.375
R8953 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n6 213.131
R8954 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t4 213.131
R8955 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t9 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t1 146.155
R8956 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t9 146.155
R8957 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t2 76.2576
R8958 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n7 76.2576
R8959 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n1 72.4424
R8960 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n2 66.4532
R8961 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t10 11.2576
R8962 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t5 11.2576
R8963 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t7 11.2576
R8964 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.t8 11.2576
R8965 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n4 5.1255
R8966 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n3 4.9096
R8967 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n0 4.7505
R8968 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n5 1.888
R8969 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_23_0.Vb2_Vb3.n0 1.888
R8970 bgr_11_0.START_UP_NFET1 bgr_11_0.START_UP_NFET1.t0 141.653
R8971 two_stage_opamp_dummy_magic_23_0.V_p_mir.n1 two_stage_opamp_dummy_magic_23_0.V_p_mir.n0 97.1193
R8972 two_stage_opamp_dummy_magic_23_0.V_p_mir.n0 two_stage_opamp_dummy_magic_23_0.V_p_mir.t0 16.0005
R8973 two_stage_opamp_dummy_magic_23_0.V_p_mir.n0 two_stage_opamp_dummy_magic_23_0.V_p_mir.t3 16.0005
R8974 two_stage_opamp_dummy_magic_23_0.V_p_mir.n1 two_stage_opamp_dummy_magic_23_0.V_p_mir.t1 9.6005
R8975 two_stage_opamp_dummy_magic_23_0.V_p_mir.t2 two_stage_opamp_dummy_magic_23_0.V_p_mir.n1 9.6005
R8976 a_6350_25058.t0 a_6350_25058.t1 178.133
R8977 a_8260_1600.n1 a_8260_1600.t0 65.3505
R8978 a_8260_1600.n3 a_8260_1600.n2 49.3505
R8979 a_8260_1600.n6 a_8260_1600.n5 49.3505
R8980 a_8260_1600.n2 a_8260_1600.t2 16.0005
R8981 a_8260_1600.n2 a_8260_1600.t4 16.0005
R8982 a_8260_1600.n6 a_8260_1600.t1 16.0005
R8983 a_8260_1600.t3 a_8260_1600.n6 16.0005
R8984 a_8260_1600.n1 a_8260_1600.n0 6.3755
R8985 a_8260_1600.n4 a_8260_1600.n1 6.1255
R8986 a_8260_1600.n5 a_8260_1600.n0 5.688
R8987 a_8260_1600.n5 a_8260_1600.n4 5.438
R8988 a_8260_1600.n3 a_8260_1600.n0 5.1255
R8989 a_8260_1600.n4 a_8260_1600.n3 4.8755
R8990 bgr_11_0.V_p_1.n1 bgr_11_0.V_p_1.n4 229.562
R8991 bgr_11_0.V_p_1.n1 bgr_11_0.V_p_1.n5 228.939
R8992 bgr_11_0.V_p_1.n0 bgr_11_0.V_p_1.n3 228.939
R8993 bgr_11_0.V_p_1.n0 bgr_11_0.V_p_1.n2 228.939
R8994 bgr_11_0.V_p_1.n6 bgr_11_0.V_p_1.n0 228.938
R8995 bgr_11_0.V_p_1.n0 bgr_11_0.V_p_1.t5 98.7279
R8996 bgr_11_0.V_p_1.n5 bgr_11_0.V_p_1.t10 48.0005
R8997 bgr_11_0.V_p_1.n5 bgr_11_0.V_p_1.t1 48.0005
R8998 bgr_11_0.V_p_1.n4 bgr_11_0.V_p_1.t2 48.0005
R8999 bgr_11_0.V_p_1.n4 bgr_11_0.V_p_1.t8 48.0005
R9000 bgr_11_0.V_p_1.n3 bgr_11_0.V_p_1.t9 48.0005
R9001 bgr_11_0.V_p_1.n3 bgr_11_0.V_p_1.t0 48.0005
R9002 bgr_11_0.V_p_1.n2 bgr_11_0.V_p_1.t3 48.0005
R9003 bgr_11_0.V_p_1.n2 bgr_11_0.V_p_1.t6 48.0005
R9004 bgr_11_0.V_p_1.t4 bgr_11_0.V_p_1.n6 48.0005
R9005 bgr_11_0.V_p_1.n6 bgr_11_0.V_p_1.t7 48.0005
R9006 bgr_11_0.V_p_1.n0 bgr_11_0.V_p_1.n1 1.8755
R9007 bgr_11_0.START_UP.n4 bgr_11_0.START_UP.t7 238.322
R9008 bgr_11_0.START_UP.n4 bgr_11_0.START_UP.t6 238.322
R9009 bgr_11_0.START_UP.n3 bgr_11_0.START_UP.n1 175.561
R9010 bgr_11_0.START_UP.n3 bgr_11_0.START_UP.n2 168.935
R9011 bgr_11_0.START_UP.n5 bgr_11_0.START_UP.n4 166.925
R9012 bgr_11_0.START_UP.n0 bgr_11_0.START_UP.t1 130.001
R9013 bgr_11_0.START_UP.n0 bgr_11_0.START_UP.t0 81.7074
R9014 bgr_11_0.START_UP bgr_11_0.START_UP.n0 36.9489
R9015 bgr_11_0.START_UP bgr_11_0.START_UP.n5 13.4693
R9016 bgr_11_0.START_UP.n2 bgr_11_0.START_UP.t4 13.1338
R9017 bgr_11_0.START_UP.n2 bgr_11_0.START_UP.t2 13.1338
R9018 bgr_11_0.START_UP.n1 bgr_11_0.START_UP.t3 13.1338
R9019 bgr_11_0.START_UP.n1 bgr_11_0.START_UP.t5 13.1338
R9020 bgr_11_0.START_UP.n5 bgr_11_0.START_UP.n3 4.21925
R9021 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 195.608
R9022 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 83.5719
R9023 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 83.5719
R9024 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 83.5719
R9025 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 83.5719
R9026 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 83.5719
R9027 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 83.5719
R9028 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 83.5719
R9029 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 83.5719
R9030 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 83.5719
R9031 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 83.5719
R9032 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 83.5719
R9033 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 83.5719
R9034 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 83.5719
R9035 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 83.5719
R9036 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 83.5719
R9037 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 83.5719
R9038 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 83.5719
R9039 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 83.5719
R9040 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 83.5719
R9041 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 83.5719
R9042 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R9043 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 83.5719
R9044 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 73.8495
R9045 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 73.8495
R9046 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 73.3165
R9047 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 73.3165
R9048 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 73.3165
R9049 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 73.3165
R9050 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 73.3165
R9051 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 73.3165
R9052 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 73.19
R9053 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 73.19
R9054 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 73.19
R9055 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 73.19
R9056 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 73.19
R9057 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 73.19
R9058 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 65.0299
R9059 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 65.0299
R9060 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 26.074
R9061 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 26.074
R9062 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 26.074
R9063 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 26.074
R9064 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 26.074
R9065 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 26.074
R9066 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 26.074
R9067 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 26.074
R9068 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 25.7843
R9069 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 25.7843
R9070 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 25.7843
R9071 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 25.7843
R9072 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 25.7843
R9073 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 25.7843
R9074 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R9075 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R9076 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R9077 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R9078 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R9079 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R9080 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R9081 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 9.3005
R9082 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R9083 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R9084 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R9085 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R9086 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 9.3005
R9087 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 9.3005
R9088 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R9089 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R9090 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R9091 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R9092 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R9093 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R9094 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R9095 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R9096 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R9097 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R9098 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R9099 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 9.3005
R9100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 9.3005
R9101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 9.3005
R9102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R9103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R9104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R9105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 9.3005
R9106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R9107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R9108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R9109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 9.3005
R9110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R9111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R9112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R9113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R9114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R9115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R9116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R9117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R9118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R9119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R9120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R9121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R9122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 9.3005
R9123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 9.3005
R9124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R9125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R9126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R9127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R9128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 4.64654
R9129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 4.64654
R9130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 4.64654
R9131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 4.64654
R9132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 4.64654
R9133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 4.64654
R9134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 4.64654
R9135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 4.64654
R9136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 4.64654
R9137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 2.36206
R9138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 2.36206
R9139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 2.36206
R9140 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 2.36206
R9141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 2.19742
R9142 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 2.19742
R9143 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 2.19742
R9144 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 2.19742
R9145 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 1.56363
R9146 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.56363
R9147 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 1.5505
R9148 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R9149 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 1.5505
R9150 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 1.5505
R9151 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 1.5505
R9152 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 1.5505
R9153 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 1.5505
R9154 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 1.5505
R9155 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 1.5505
R9156 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 1.5505
R9157 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 1.5505
R9158 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 1.5505
R9159 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 1.5505
R9160 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 1.5505
R9161 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 1.5505
R9162 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 1.5505
R9163 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 1.5505
R9164 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 1.5505
R9165 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.25468
R9166 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 1.25468
R9167 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.25468
R9168 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.25468
R9169 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 1.25468
R9170 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 1.25468
R9171 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 1.19225
R9172 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 1.19225
R9173 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 1.19225
R9174 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 1.19225
R9175 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 1.19225
R9176 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.19225
R9177 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 1.07024
R9178 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 1.07024
R9179 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 1.07024
R9180 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 1.07024
R9181 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 1.07024
R9182 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.07024
R9183 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.0237
R9184 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 1.0237
R9185 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.0237
R9186 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.0237
R9187 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 1.0237
R9188 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 1.0237
R9189 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.885803
R9190 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 0.885803
R9191 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 0.885803
R9192 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 0.885803
R9193 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.885803
R9194 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.885803
R9195 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 0.885803
R9196 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.885803
R9197 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 0.812055
R9198 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 0.812055
R9199 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.77514
R9200 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.77514
R9201 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 0.77514
R9202 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.77514
R9203 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.77514
R9204 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 0.77514
R9205 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 0.77514
R9206 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 0.77514
R9207 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.756696
R9208 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R9209 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.756696
R9210 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 0.756696
R9211 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R9212 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.756696
R9213 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R9214 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.756696
R9215 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 0.711459
R9216 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.711459
R9217 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.647417
R9218 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 0.647417
R9219 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.590702
R9220 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 0.590702
R9221 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.590702
R9222 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 0.590702
R9223 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.590702
R9224 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 0.590702
R9225 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.576566
R9226 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.576566
R9227 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 0.530034
R9228 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 0.530034
R9229 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 0.290206
R9230 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 0.290206
R9231 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 0.290206
R9232 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 0.290206
R9233 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 0.290206
R9234 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 0.290206
R9235 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 0.290206
R9236 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 0.290206
R9237 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R9238 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R9239 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R9240 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.203382
R9241 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R9242 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 0.203382
R9243 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 0.154071
R9244 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 0.154071
R9245 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 0.154071
R9246 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 0.154071
R9247 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 0.137464
R9248 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 0.137464
R9249 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 0.134964
R9250 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 0.134964
R9251 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R9252 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 0.0183571
R9253 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R9254 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R9255 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 0.0183571
R9256 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R9257 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R9258 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 0.0183571
R9259 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0183571
R9260 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R9261 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R9262 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R9263 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R9264 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 0.0183571
R9265 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R9266 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R9267 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 0.0183571
R9268 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0183571
R9269 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0106786
R9270 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0106786
R9271 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.0106786
R9272 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 0.00992001
R9273 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 0.00992001
R9274 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R9275 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 0.00992001
R9276 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R9277 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R9278 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R9279 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 0.00992001
R9280 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 0.00992001
R9281 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 0.00992001
R9282 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R9283 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 0.00992001
R9284 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R9285 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R9286 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R9287 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R9288 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 0.00992001
R9289 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R9290 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.00817857
R9291 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00817857
R9292 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 0.00817857
R9293 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 0.00817857
R9294 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.00817857
R9295 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t8 525.38
R9296 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t3 525.38
R9297 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t5 483.608
R9298 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t6 360.43
R9299 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t2 291.209
R9300 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t4 281.168
R9301 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t9 281.168
R9302 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t7 281.168
R9303 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n3 244.214
R9304 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n0 202.44
R9305 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n1 202.159
R9306 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n5 165.972
R9307 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t0 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n6 117.754
R9308 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t1 117.254
R9309 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n4 79.2627
R9310 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n2 18.9067
R9311 a_4200_4468.t0 a_4200_4468.t1 169.905
R9312 two_stage_opamp_dummy_magic_23_0.V_tot.n6 two_stage_opamp_dummy_magic_23_0.V_tot.n5 771.76
R9313 two_stage_opamp_dummy_magic_23_0.V_tot.n1 two_stage_opamp_dummy_magic_23_0.V_tot.n0 595.444
R9314 two_stage_opamp_dummy_magic_23_0.V_tot.n11 two_stage_opamp_dummy_magic_23_0.V_tot.n10 595.131
R9315 two_stage_opamp_dummy_magic_23_0.V_tot.n5 two_stage_opamp_dummy_magic_23_0.V_tot.n4 530.201
R9316 two_stage_opamp_dummy_magic_23_0.V_tot.n3 two_stage_opamp_dummy_magic_23_0.V_tot.n2 530.201
R9317 two_stage_opamp_dummy_magic_23_0.V_tot.n9 two_stage_opamp_dummy_magic_23_0.V_tot.n8 530.201
R9318 two_stage_opamp_dummy_magic_23_0.V_tot.n7 two_stage_opamp_dummy_magic_23_0.V_tot.n6 530.201
R9319 two_stage_opamp_dummy_magic_23_0.V_tot.n1 two_stage_opamp_dummy_magic_23_0.V_tot.t11 208.868
R9320 two_stage_opamp_dummy_magic_23_0.V_tot.n2 two_stage_opamp_dummy_magic_23_0.V_tot.t4 208.868
R9321 two_stage_opamp_dummy_magic_23_0.V_tot.n3 two_stage_opamp_dummy_magic_23_0.V_tot.t10 208.868
R9322 two_stage_opamp_dummy_magic_23_0.V_tot.n4 two_stage_opamp_dummy_magic_23_0.V_tot.t7 208.868
R9323 two_stage_opamp_dummy_magic_23_0.V_tot.n5 two_stage_opamp_dummy_magic_23_0.V_tot.t9 208.868
R9324 two_stage_opamp_dummy_magic_23_0.V_tot.n6 two_stage_opamp_dummy_magic_23_0.V_tot.t8 208.868
R9325 two_stage_opamp_dummy_magic_23_0.V_tot.n7 two_stage_opamp_dummy_magic_23_0.V_tot.t13 208.868
R9326 two_stage_opamp_dummy_magic_23_0.V_tot.n8 two_stage_opamp_dummy_magic_23_0.V_tot.t6 208.868
R9327 two_stage_opamp_dummy_magic_23_0.V_tot.n9 two_stage_opamp_dummy_magic_23_0.V_tot.t12 208.868
R9328 two_stage_opamp_dummy_magic_23_0.V_tot.n10 two_stage_opamp_dummy_magic_23_0.V_tot.t5 208.868
R9329 two_stage_opamp_dummy_magic_23_0.V_tot.n4 two_stage_opamp_dummy_magic_23_0.V_tot.n3 176.733
R9330 two_stage_opamp_dummy_magic_23_0.V_tot.n2 two_stage_opamp_dummy_magic_23_0.V_tot.n1 176.733
R9331 two_stage_opamp_dummy_magic_23_0.V_tot.n10 two_stage_opamp_dummy_magic_23_0.V_tot.n9 176.733
R9332 two_stage_opamp_dummy_magic_23_0.V_tot.n8 two_stage_opamp_dummy_magic_23_0.V_tot.n7 176.733
R9333 two_stage_opamp_dummy_magic_23_0.V_tot.n0 two_stage_opamp_dummy_magic_23_0.V_tot.t2 117.591
R9334 two_stage_opamp_dummy_magic_23_0.V_tot.t0 two_stage_opamp_dummy_magic_23_0.V_tot.n11 117.591
R9335 two_stage_opamp_dummy_magic_23_0.V_tot.n11 two_stage_opamp_dummy_magic_23_0.V_tot.t3 108.424
R9336 two_stage_opamp_dummy_magic_23_0.V_tot.n0 two_stage_opamp_dummy_magic_23_0.V_tot.t1 108.424
R9337 a_5820_23634.t0 a_5820_23634.t1 178.133
R9338 a_11420_25058.t0 a_11420_25058.t1 178.133
R9339 a_11950_23700.t0 a_11950_23700.t1 178.133
R9340 a_4600_1446.t0 a_4600_1446.t1 169.905
R9341 a_4080_4468.t0 a_4080_4468.t1 294.339
R9342 a_13130_1456.t0 a_13130_1456.t1 169.905
R9343 a_5700_24908.t0 a_5700_24908.t1 178.133
R9344 a_11300_23450.t0 a_11300_23450.t1 178.133
R9345 a_13450_4368.t0 a_13450_4368.t1 294.339
R9346 a_13570_4368.t0 a_13570_4368.t1 169.905
C0 bgr_11_0.START_UP bgr_11_0.NFET_GATE_10uA 1.64177f
C1 VDDA two_stage_opamp_dummy_magic_23_0.V_err_gate 2.31861f
C2 two_stage_opamp_dummy_magic_23_0.V_err_gate two_stage_opamp_dummy_magic_23_0.V_tail_gate 1.43091f
C3 two_stage_opamp_dummy_magic_23_0.X two_stage_opamp_dummy_magic_23_0.err_amp_out 0.20522f
C4 VDDA bgr_11_0.START_UP 1.26407f
C5 VOUT+ two_stage_opamp_dummy_magic_23_0.VD4 0.028865f
C6 VDDA two_stage_opamp_dummy_magic_23_0.err_amp_out 1.0994f
C7 two_stage_opamp_dummy_magic_23_0.V_tail_gate two_stage_opamp_dummy_magic_23_0.err_amp_out 0.343731f
C8 bgr_11_0.PFET_GATE_10uA bgr_11_0.START_UP_NFET1 0.0108f
C9 bgr_11_0.1st_Vout_1 bgr_11_0.V_TOP 2.48406f
C10 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref two_stage_opamp_dummy_magic_23_0.V_err_gate 0.492517f
C11 bgr_11_0.PFET_GATE_10uA bgr_11_0.V_TOP 0.221314f
C12 bgr_11_0.1st_Vout_1 bgr_11_0.NFET_GATE_10uA 0.038363f
C13 two_stage_opamp_dummy_magic_23_0.VD4 two_stage_opamp_dummy_magic_23_0.cap_res_Y 0.054393f
C14 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref bgr_11_0.START_UP 1.36583f
C15 VDDA bgr_11_0.1st_Vout_1 1.3286f
C16 bgr_11_0.PFET_GATE_10uA bgr_11_0.NFET_GATE_10uA 0.012365f
C17 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref two_stage_opamp_dummy_magic_23_0.err_amp_out 0.289292f
C18 VDDA two_stage_opamp_dummy_magic_23_0.VD4 8.479321f
C19 VDDA bgr_11_0.PFET_GATE_10uA 7.75313f
C20 VOUT+ VOUT- 0.305434f
C21 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_23_0.V_tail_gate 0.24038f
C22 two_stage_opamp_dummy_magic_23_0.V_err_gate two_stage_opamp_dummy_magic_23_0.err_amp_out 0.026461f
C23 VIN+ two_stage_opamp_dummy_magic_23_0.VD2 0.510937f
C24 VOUT+ two_stage_opamp_dummy_magic_23_0.cap_res_Y 50.8462f
C25 VDDA two_stage_opamp_dummy_magic_23_0.VD2 0.027746f
C26 bgr_11_0.START_UP_NFET1 bgr_11_0.NFET_GATE_10uA 0.351171f
C27 two_stage_opamp_dummy_magic_23_0.VD2 two_stage_opamp_dummy_magic_23_0.V_tail_gate 0.02379f
C28 VDDA VOUT+ 13.4377f
C29 two_stage_opamp_dummy_magic_23_0.VD4 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref 0.04352f
C30 VOUT- two_stage_opamp_dummy_magic_23_0.cap_res_Y 0.028842f
C31 VOUT+ two_stage_opamp_dummy_magic_23_0.V_tail_gate 0.010408f
C32 VDDA bgr_11_0.START_UP_NFET1 0.167059f
C33 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.V_TOP 0.055802f
C34 VOUT- two_stage_opamp_dummy_magic_23_0.X 2.33193f
C35 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_23_0.V_err_amp_ref 1.67528f
C36 two_stage_opamp_dummy_magic_23_0.V_err_gate bgr_11_0.1st_Vout_1 0.040732f
C37 bgr_11_0.V_TOP bgr_11_0.NFET_GATE_10uA 0.043918f
C38 bgr_11_0.START_UP bgr_11_0.1st_Vout_1 0.043153f
C39 VDDA VOUT- 13.403299f
C40 VOUT- two_stage_opamp_dummy_magic_23_0.V_tail_gate 0.02527f
C41 VDDA bgr_11_0.V_TOP 13.6718f
C42 VDDA bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.046803f
C43 VDDA two_stage_opamp_dummy_magic_23_0.cap_res_Y 0.533063f
C44 two_stage_opamp_dummy_magic_23_0.V_tail_gate two_stage_opamp_dummy_magic_23_0.cap_res_Y 0.03128f
C45 VIN+ VIN- 0.151796f
C46 VIN+ two_stage_opamp_dummy_magic_23_0.V_tail_gate 0.056847f
C47 VDDA two_stage_opamp_dummy_magic_23_0.X 5.01789f
C48 VDDA bgr_11_0.NFET_GATE_10uA 0.893844f
C49 VOUT+ two_stage_opamp_dummy_magic_23_0.V_err_amp_ref 0.039549f
C50 two_stage_opamp_dummy_magic_23_0.V_tail_gate two_stage_opamp_dummy_magic_23_0.X 0.18001f
C51 two_stage_opamp_dummy_magic_23_0.V_tail_gate bgr_11_0.NFET_GATE_10uA 0.038519f
C52 VDDA two_stage_opamp_dummy_magic_23_0.V_tail_gate 5.00585f
C53 VIN- two_stage_opamp_dummy_magic_23_0.V_tail_gate 0.135101f
C54 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref bgr_11_0.V_TOP 0.583702f
C55 bgr_11_0.START_UP_NFET1 bgr_11_0.START_UP 0.145663f
C56 VOUT- two_stage_opamp_dummy_magic_23_0.V_err_gate 0.038404f
C57 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref two_stage_opamp_dummy_magic_23_0.cap_res_Y 0.243261f
C58 two_stage_opamp_dummy_magic_23_0.V_err_gate bgr_11_0.V_TOP 0.075936f
C59 bgr_11_0.START_UP bgr_11_0.V_TOP 0.740874f
C60 VDDA two_stage_opamp_dummy_magic_23_0.V_err_amp_ref 4.03349f
C61 two_stage_opamp_dummy_magic_23_0.V_err_gate two_stage_opamp_dummy_magic_23_0.X 0.161254f
C62 two_stage_opamp_dummy_magic_23_0.V_err_gate bgr_11_0.NFET_GATE_10uA 3.46607f
C63 VIN- GNDA 1.92317f
C64 VIN+ GNDA 1.90963f
C65 VOUT- GNDA 20.532288f
C66 VOUT+ GNDA 20.582405f
C67 VDDA GNDA 0.228872p
C68 two_stage_opamp_dummy_magic_23_0.VD2 GNDA 2.003606f
C69 two_stage_opamp_dummy_magic_23_0.err_amp_out GNDA 5.194764f
C70 two_stage_opamp_dummy_magic_23_0.cap_res_Y GNDA 33.372776f
C71 two_stage_opamp_dummy_magic_23_0.X GNDA 7.15177f
C72 two_stage_opamp_dummy_magic_23_0.V_tail_gate GNDA 9.812429f
C73 bgr_11_0.1st_Vout_1 GNDA 7.474261f
C74 bgr_11_0.START_UP GNDA 5.955617f
C75 bgr_11_0.START_UP_NFET1 GNDA 4.27813f
C76 two_stage_opamp_dummy_magic_23_0.V_err_gate GNDA 13.4333f
C77 bgr_11_0.NFET_GATE_10uA GNDA 8.00746f
C78 bgr_11_0.V_TOP GNDA 9.658216f
C79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA 17.8988f
C80 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref GNDA 9.053741f
C81 bgr_11_0.PFET_GATE_10uA GNDA 6.62186f
C82 two_stage_opamp_dummy_magic_23_0.VD4 GNDA 5.12103f
C83 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t1 GNDA 0.124526f
C84 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t5 GNDA 0.365905f
C85 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t7 GNDA 0.313782f
C86 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t3 GNDA 0.37241f
C87 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n0 GNDA 0.195093f
C88 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t2 GNDA 0.317627f
C89 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n1 GNDA 0.210094f
C90 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n2 GNDA 0.585951f
C91 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t6 GNDA 0.340499f
C92 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t9 GNDA 0.313782f
C93 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t4 GNDA 0.313782f
C94 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t8 GNDA 0.37241f
C95 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n3 GNDA 0.196704f
C96 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n4 GNDA 0.124569f
C97 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n5 GNDA 0.118809f
C98 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.n6 GNDA 0.608541f
C99 two_stage_opamp_dummy_magic_23_0.V_b_2nd_stage.t0 GNDA 0.125517f
C100 bgr_11_0.START_UP.t0 GNDA 1.06745f
C101 bgr_11_0.START_UP.t1 GNDA 0.02806f
C102 bgr_11_0.START_UP.n0 GNDA 0.714928f
C103 bgr_11_0.START_UP.t3 GNDA 0.026778f
C104 bgr_11_0.START_UP.t5 GNDA 0.026778f
C105 bgr_11_0.START_UP.n1 GNDA 0.097147f
C106 bgr_11_0.START_UP.t4 GNDA 0.026778f
C107 bgr_11_0.START_UP.t2 GNDA 0.026778f
C108 bgr_11_0.START_UP.n2 GNDA 0.08937f
C109 bgr_11_0.START_UP.n3 GNDA 0.462855f
C110 bgr_11_0.START_UP.t6 GNDA 0.010062f
C111 bgr_11_0.START_UP.t7 GNDA 0.010062f
C112 bgr_11_0.START_UP.n4 GNDA 0.028407f
C113 bgr_11_0.START_UP.n5 GNDA 0.260836f
C114 a_8260_1600.t1 GNDA 0.047649f
C115 a_8260_1600.n0 GNDA 0.318351f
C116 a_8260_1600.t0 GNDA 0.161927f
C117 a_8260_1600.n1 GNDA 0.491746f
C118 a_8260_1600.t2 GNDA 0.047649f
C119 a_8260_1600.t4 GNDA 0.047649f
C120 a_8260_1600.n2 GNDA 0.103679f
C121 a_8260_1600.n3 GNDA 0.407675f
C122 a_8260_1600.n4 GNDA 0.297965f
C123 a_8260_1600.n5 GNDA 0.42438f
C124 a_8260_1600.n6 GNDA 0.103679f
C125 a_8260_1600.t3 GNDA 0.047649f
C126 bgr_11_0.V_mir1.t5 GNDA 0.019544f
C127 bgr_11_0.V_mir1.t0 GNDA 0.029773f
C128 bgr_11_0.V_mir1.t6 GNDA 0.023453f
C129 bgr_11_0.V_mir1.t22 GNDA 0.023453f
C130 bgr_11_0.V_mir1.t17 GNDA 0.037856f
C131 bgr_11_0.V_mir1.n0 GNDA 0.042274f
C132 bgr_11_0.V_mir1.n1 GNDA 0.028879f
C133 bgr_11_0.V_mir1.n2 GNDA 0.044932f
C134 bgr_11_0.V_mir1.t1 GNDA 0.019544f
C135 bgr_11_0.V_mir1.t7 GNDA 0.019544f
C136 bgr_11_0.V_mir1.n3 GNDA 0.044741f
C137 bgr_11_0.V_mir1.n4 GNDA 0.11173f
C138 bgr_11_0.V_mir1.n5 GNDA 0.025551f
C139 bgr_11_0.V_mir1.t12 GNDA 0.041699f
C140 bgr_11_0.V_mir1.n6 GNDA 0.027738f
C141 bgr_11_0.V_mir1.n7 GNDA 0.457418f
C142 bgr_11_0.V_mir1.n8 GNDA 0.148244f
C143 bgr_11_0.V_mir1.t2 GNDA 0.029773f
C144 bgr_11_0.V_mir1.t8 GNDA 0.023453f
C145 bgr_11_0.V_mir1.t21 GNDA 0.023453f
C146 bgr_11_0.V_mir1.t19 GNDA 0.037856f
C147 bgr_11_0.V_mir1.n9 GNDA 0.042274f
C148 bgr_11_0.V_mir1.n10 GNDA 0.028879f
C149 bgr_11_0.V_mir1.n11 GNDA 0.044932f
C150 bgr_11_0.V_mir1.t3 GNDA 0.019544f
C151 bgr_11_0.V_mir1.t9 GNDA 0.019544f
C152 bgr_11_0.V_mir1.n12 GNDA 0.044741f
C153 bgr_11_0.V_mir1.n13 GNDA 0.086204f
C154 bgr_11_0.V_mir1.n14 GNDA 0.051792f
C155 bgr_11_0.V_mir1.n15 GNDA 0.355461f
C156 bgr_11_0.V_mir1.t4 GNDA 0.029773f
C157 bgr_11_0.V_mir1.t10 GNDA 0.023453f
C158 bgr_11_0.V_mir1.t20 GNDA 0.023453f
C159 bgr_11_0.V_mir1.t18 GNDA 0.037856f
C160 bgr_11_0.V_mir1.n16 GNDA 0.042274f
C161 bgr_11_0.V_mir1.n17 GNDA 0.028879f
C162 bgr_11_0.V_mir1.n18 GNDA 0.044932f
C163 bgr_11_0.V_mir1.n19 GNDA 0.11173f
C164 bgr_11_0.V_mir1.n20 GNDA 0.044741f
C165 bgr_11_0.V_mir1.t11 GNDA 0.019544f
C166 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t0 GNDA 0.028527f
C167 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t3 GNDA 0.028527f
C168 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n0 GNDA 0.103686f
C169 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t2 GNDA 0.028527f
C170 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t1 GNDA 0.028527f
C171 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n1 GNDA 0.086163f
C172 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n2 GNDA 1.68702f
C173 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t4 GNDA 0.355774f
C174 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n3 GNDA 0.099225f
C175 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n4 GNDA 0.170727f
C176 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t6 GNDA 0.08558f
C177 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t10 GNDA 0.08558f
C178 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n5 GNDA 0.183039f
C179 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n6 GNDA 0.572546f
C180 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t5 GNDA 0.08558f
C181 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t12 GNDA 0.08558f
C182 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n7 GNDA 0.183039f
C183 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n8 GNDA 0.557039f
C184 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n9 GNDA 0.170727f
C185 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n10 GNDA 0.099225f
C186 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t7 GNDA 0.08558f
C187 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t11 GNDA 0.08558f
C188 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n11 GNDA 0.183039f
C189 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n12 GNDA 0.557039f
C190 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n13 GNDA 0.099225f
C191 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t8 GNDA 0.08558f
C192 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t13 GNDA 0.08558f
C193 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n14 GNDA 0.183039f
C194 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n15 GNDA 0.557039f
C195 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n16 GNDA 0.170727f
C196 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t9 GNDA 0.08558f
C197 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.t14 GNDA 0.08558f
C198 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n17 GNDA 0.183039f
C199 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n18 GNDA 0.564792f
C200 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n19 GNDA 0.22124f
C201 two_stage_opamp_dummy_magic_23_0.V_CMFB_S2.n20 GNDA 2.35028f
C202 bgr_11_0.V_CMFB_S2 GNDA 2.89243f
C203 a_7460_6300.t8 GNDA 0.020006f
C204 a_7460_6300.n0 GNDA 0.210468f
C205 a_7460_6300.t4 GNDA 0.020006f
C206 a_7460_6300.t7 GNDA 0.020006f
C207 a_7460_6300.n1 GNDA 0.040763f
C208 a_7460_6300.n2 GNDA 0.365375f
C209 a_7460_6300.n3 GNDA 0.319666f
C210 a_7460_6300.t1 GNDA 0.020006f
C211 a_7460_6300.t5 GNDA 0.020006f
C212 a_7460_6300.n4 GNDA 0.040763f
C213 a_7460_6300.n5 GNDA 0.306668f
C214 a_7460_6300.n6 GNDA 0.335179f
C215 a_7460_6300.t13 GNDA 0.020006f
C216 a_7460_6300.t11 GNDA 0.020006f
C217 a_7460_6300.n7 GNDA 0.040763f
C218 a_7460_6300.n8 GNDA 0.191134f
C219 a_7460_6300.t19 GNDA 0.020006f
C220 a_7460_6300.t16 GNDA 0.020006f
C221 a_7460_6300.n9 GNDA 0.040763f
C222 a_7460_6300.n10 GNDA 0.300378f
C223 a_7460_6300.n11 GNDA 0.215758f
C224 a_7460_6300.n12 GNDA 0.206718f
C225 a_7460_6300.t18 GNDA 0.020006f
C226 a_7460_6300.t14 GNDA 0.020006f
C227 a_7460_6300.n13 GNDA 0.040763f
C228 a_7460_6300.n14 GNDA 0.300378f
C229 a_7460_6300.t12 GNDA 0.020006f
C230 a_7460_6300.t0 GNDA 0.020006f
C231 a_7460_6300.n15 GNDA 0.040763f
C232 a_7460_6300.n16 GNDA 0.279938f
C233 a_7460_6300.n17 GNDA 0.206718f
C234 a_7460_6300.n18 GNDA 0.122442f
C235 a_7460_6300.t17 GNDA 0.020006f
C236 a_7460_6300.t15 GNDA 0.020006f
C237 a_7460_6300.n19 GNDA 0.040763f
C238 a_7460_6300.n20 GNDA 0.279938f
C239 a_7460_6300.n21 GNDA 0.127024f
C240 a_7460_6300.n22 GNDA 0.208769f
C241 a_7460_6300.n23 GNDA 0.121174f
C242 a_7460_6300.n24 GNDA 0.18461f
C243 a_7460_6300.t6 GNDA 0.020006f
C244 a_7460_6300.t2 GNDA 0.020006f
C245 a_7460_6300.n25 GNDA 0.040763f
C246 a_7460_6300.n26 GNDA 0.233788f
C247 a_7460_6300.n27 GNDA 0.319666f
C248 a_7460_6300.t9 GNDA 0.020006f
C249 a_7460_6300.t3 GNDA 0.020006f
C250 a_7460_6300.n28 GNDA 0.040763f
C251 a_7460_6300.n29 GNDA 0.306668f
C252 a_7460_6300.n30 GNDA 0.324795f
C253 a_7460_6300.n31 GNDA 0.218329f
C254 a_7460_6300.n32 GNDA 0.306668f
C255 a_7460_6300.n33 GNDA 0.040763f
C256 a_7460_6300.t10 GNDA 0.020006f
C257 bgr_11_0.Vin+.t7 GNDA 0.010696f
C258 bgr_11_0.Vin+.t8 GNDA 0.025367f
C259 bgr_11_0.Vin+.t9 GNDA 0.01649f
C260 bgr_11_0.Vin+.n0 GNDA 0.054406f
C261 bgr_11_0.Vin+.t6 GNDA 0.01649f
C262 bgr_11_0.Vin+.n1 GNDA 0.042338f
C263 bgr_11_0.Vin+.t10 GNDA 0.01649f
C264 bgr_11_0.Vin+.n2 GNDA 0.042909f
C265 bgr_11_0.Vin+.n3 GNDA 0.130793f
C266 bgr_11_0.Vin+.t5 GNDA 0.05348f
C267 bgr_11_0.Vin+.t4 GNDA 0.05348f
C268 bgr_11_0.Vin+.n4 GNDA 0.17668f
C269 bgr_11_0.Vin+.n5 GNDA 1.27851f
C270 bgr_11_0.Vin+.t3 GNDA 0.05348f
C271 bgr_11_0.Vin+.t2 GNDA 0.05348f
C272 bgr_11_0.Vin+.n6 GNDA 0.17668f
C273 bgr_11_0.Vin+.n7 GNDA 1.06526f
C274 bgr_11_0.Vin+.t1 GNDA 0.232527f
C275 bgr_11_0.Vin+.n8 GNDA 1.7265f
C276 bgr_11_0.Vin+.t0 GNDA 0.173951f
C277 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n0 GNDA 0.408216f
C278 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n1 GNDA 0.318908f
C279 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n2 GNDA 0.362794f
C280 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t6 GNDA 0.014742f
C281 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t14 GNDA 0.014742f
C282 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t8 GNDA 0.014742f
C283 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n3 GNDA 0.031178f
C284 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n4 GNDA 0.293793f
C285 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t9 GNDA 0.012162f
C286 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t19 GNDA 0.012162f
C287 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t21 GNDA 0.012162f
C288 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t5 GNDA 0.012162f
C289 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t11 GNDA 0.012162f
C290 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t20 GNDA 0.012162f
C291 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t17 GNDA 0.012162f
C292 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t7 GNDA 0.026351f
C293 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n5 GNDA 0.041093f
C294 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n6 GNDA 0.032064f
C295 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n7 GNDA 0.028584f
C296 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n8 GNDA 0.04506f
C297 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n9 GNDA 0.028584f
C298 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n10 GNDA 0.032064f
C299 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n11 GNDA 0.032064f
C300 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n12 GNDA 0.028584f
C301 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t3 GNDA 0.012162f
C302 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t18 GNDA 0.026351f
C303 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n13 GNDA 0.037614f
C304 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n14 GNDA 0.04506f
C305 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t16 GNDA 0.014742f
C306 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t1 GNDA 0.014742f
C307 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n15 GNDA 0.030038f
C308 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t0 GNDA 0.014742f
C309 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t2 GNDA 0.014742f
C310 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n16 GNDA 0.030038f
C311 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n17 GNDA 0.249418f
C312 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n18 GNDA 0.316023f
C313 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t15 GNDA 0.014742f
C314 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t13 GNDA 0.014742f
C315 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n19 GNDA 0.030038f
C316 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n20 GNDA 0.249418f
C317 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n21 GNDA 0.320943f
C318 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n22 GNDA 0.239385f
C319 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n23 GNDA 0.23177f
C320 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t10 GNDA 0.014742f
C321 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t4 GNDA 0.014742f
C322 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n24 GNDA 0.031178f
C323 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n25 GNDA 0.348011f
C324 two_stage_opamp_dummy_magic_23_0.err_amp_mir.n26 GNDA 0.031178f
C325 two_stage_opamp_dummy_magic_23_0.err_amp_mir.t12 GNDA 0.014742f
C326 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t14 GNDA 0.029652f
C327 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t1 GNDA 0.029652f
C328 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n0 GNDA 0.107777f
C329 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t3 GNDA 0.029652f
C330 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t2 GNDA 0.029652f
C331 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n1 GNDA 0.089562f
C332 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n2 GNDA 1.75357f
C333 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t0 GNDA 0.368222f
C334 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n3 GNDA 0.103139f
C335 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n4 GNDA 0.177463f
C336 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t4 GNDA 0.088956f
C337 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t8 GNDA 0.088956f
C338 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n5 GNDA 0.19026f
C339 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n6 GNDA 0.595133f
C340 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t13 GNDA 0.088956f
C341 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t11 GNDA 0.088956f
C342 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n7 GNDA 0.19026f
C343 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n8 GNDA 0.579015f
C344 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n9 GNDA 0.177463f
C345 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n10 GNDA 0.103139f
C346 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t6 GNDA 0.088956f
C347 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t10 GNDA 0.088956f
C348 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n11 GNDA 0.19026f
C349 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n12 GNDA 0.579015f
C350 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n13 GNDA 0.103139f
C351 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t5 GNDA 0.088956f
C352 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t9 GNDA 0.088956f
C353 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n14 GNDA 0.19026f
C354 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n15 GNDA 0.579015f
C355 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n16 GNDA 0.177463f
C356 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t12 GNDA 0.088956f
C357 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.t7 GNDA 0.088956f
C358 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n17 GNDA 0.19026f
C359 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n18 GNDA 0.587074f
C360 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n19 GNDA 0.232126f
C361 two_stage_opamp_dummy_magic_23_0.V_CMFB_S4.n20 GNDA 2.41715f
C362 bgr_11_0.V_CMFB_S4 GNDA 3.01107f
C363 two_stage_opamp_dummy_magic_23_0.err_amp_out.n0 GNDA 0.095072f
C364 two_stage_opamp_dummy_magic_23_0.err_amp_out.t12 GNDA 0.054088f
C365 two_stage_opamp_dummy_magic_23_0.err_amp_out.n1 GNDA 0.012001f
C366 two_stage_opamp_dummy_magic_23_0.err_amp_out.n2 GNDA 0.124861f
C367 two_stage_opamp_dummy_magic_23_0.err_amp_out.n3 GNDA 0.012001f
C368 two_stage_opamp_dummy_magic_23_0.err_amp_out.n4 GNDA 0.10815f
C369 two_stage_opamp_dummy_magic_23_0.err_amp_out.n5 GNDA 0.095072f
C370 two_stage_opamp_dummy_magic_23_0.err_amp_out.n6 GNDA 0.719147f
C371 two_stage_opamp_dummy_magic_23_0.err_amp_out.n7 GNDA 0.012001f
C372 two_stage_opamp_dummy_magic_23_0.err_amp_out.n8 GNDA 0.10815f
C373 two_stage_opamp_dummy_magic_23_0.err_amp_out.n9 GNDA 0.057175f
C374 two_stage_opamp_dummy_magic_23_0.err_amp_out.n10 GNDA 0.012844f
C375 two_stage_opamp_dummy_magic_23_0.err_amp_out.n11 GNDA 0.012527f
C376 two_stage_opamp_dummy_magic_23_0.err_amp_out.n12 GNDA 0.325317f
C377 two_stage_opamp_dummy_magic_23_0.err_amp_out.n13 GNDA 0.012527f
C378 two_stage_opamp_dummy_magic_23_0.V_err_p.n0 GNDA 0.388376f
C379 two_stage_opamp_dummy_magic_23_0.V_err_p.t18 GNDA 0.023181f
C380 two_stage_opamp_dummy_magic_23_0.V_err_p.n1 GNDA 0.38098f
C381 two_stage_opamp_dummy_magic_23_0.V_err_p.n2 GNDA 0.243876f
C382 two_stage_opamp_dummy_magic_23_0.V_err_p.t19 GNDA 0.023181f
C383 two_stage_opamp_dummy_magic_23_0.V_err_p.t11 GNDA 0.023181f
C384 two_stage_opamp_dummy_magic_23_0.V_err_p.n3 GNDA 0.047234f
C385 two_stage_opamp_dummy_magic_23_0.V_err_p.n4 GNDA 0.392203f
C386 two_stage_opamp_dummy_magic_23_0.V_err_p.t13 GNDA 0.023181f
C387 two_stage_opamp_dummy_magic_23_0.V_err_p.t20 GNDA 0.023181f
C388 two_stage_opamp_dummy_magic_23_0.V_err_p.n5 GNDA 0.047234f
C389 two_stage_opamp_dummy_magic_23_0.V_err_p.n6 GNDA 0.230943f
C390 two_stage_opamp_dummy_magic_23_0.V_err_p.n7 GNDA 0.147187f
C391 two_stage_opamp_dummy_magic_23_0.V_err_p.t15 GNDA 0.023181f
C392 two_stage_opamp_dummy_magic_23_0.V_err_p.t0 GNDA 0.023181f
C393 two_stage_opamp_dummy_magic_23_0.V_err_p.n8 GNDA 0.047234f
C394 two_stage_opamp_dummy_magic_23_0.V_err_p.n9 GNDA 0.348058f
C395 two_stage_opamp_dummy_magic_23_0.V_err_p.n10 GNDA 0.250006f
C396 two_stage_opamp_dummy_magic_23_0.V_err_p.t2 GNDA 0.023181f
C397 two_stage_opamp_dummy_magic_23_0.V_err_p.t14 GNDA 0.023181f
C398 two_stage_opamp_dummy_magic_23_0.V_err_p.n11 GNDA 0.047234f
C399 two_stage_opamp_dummy_magic_23_0.V_err_p.n12 GNDA 0.324373f
C400 two_stage_opamp_dummy_magic_23_0.V_err_p.n13 GNDA 0.239531f
C401 two_stage_opamp_dummy_magic_23_0.V_err_p.t16 GNDA 0.023181f
C402 two_stage_opamp_dummy_magic_23_0.V_err_p.t21 GNDA 0.023181f
C403 two_stage_opamp_dummy_magic_23_0.V_err_p.n14 GNDA 0.047234f
C404 two_stage_opamp_dummy_magic_23_0.V_err_p.n15 GNDA 0.324373f
C405 two_stage_opamp_dummy_magic_23_0.V_err_p.n16 GNDA 0.141878f
C406 two_stage_opamp_dummy_magic_23_0.V_err_p.n17 GNDA 0.239531f
C407 two_stage_opamp_dummy_magic_23_0.V_err_p.t1 GNDA 0.023181f
C408 two_stage_opamp_dummy_magic_23_0.V_err_p.t17 GNDA 0.023181f
C409 two_stage_opamp_dummy_magic_23_0.V_err_p.n18 GNDA 0.047234f
C410 two_stage_opamp_dummy_magic_23_0.V_err_p.n19 GNDA 0.324373f
C411 two_stage_opamp_dummy_magic_23_0.V_err_p.n20 GNDA 0.241974f
C412 two_stage_opamp_dummy_magic_23_0.V_err_p.n21 GNDA 0.226203f
C413 two_stage_opamp_dummy_magic_23_0.V_err_p.n22 GNDA 0.367618f
C414 two_stage_opamp_dummy_magic_23_0.V_err_p.t4 GNDA 0.023181f
C415 two_stage_opamp_dummy_magic_23_0.V_err_p.t9 GNDA 0.023181f
C416 two_stage_opamp_dummy_magic_23_0.V_err_p.n23 GNDA 0.047234f
C417 two_stage_opamp_dummy_magic_23_0.V_err_p.n24 GNDA 0.38098f
C418 two_stage_opamp_dummy_magic_23_0.V_err_p.t3 GNDA 0.023181f
C419 two_stage_opamp_dummy_magic_23_0.V_err_p.t8 GNDA 0.023181f
C420 two_stage_opamp_dummy_magic_23_0.V_err_p.n25 GNDA 0.047234f
C421 two_stage_opamp_dummy_magic_23_0.V_err_p.n26 GNDA 0.324373f
C422 two_stage_opamp_dummy_magic_23_0.V_err_p.n27 GNDA 0.249186f
C423 two_stage_opamp_dummy_magic_23_0.V_err_p.n28 GNDA 0.249186f
C424 two_stage_opamp_dummy_magic_23_0.V_err_p.t5 GNDA 0.023181f
C425 two_stage_opamp_dummy_magic_23_0.V_err_p.t7 GNDA 0.023181f
C426 two_stage_opamp_dummy_magic_23_0.V_err_p.n29 GNDA 0.047234f
C427 two_stage_opamp_dummy_magic_23_0.V_err_p.n30 GNDA 0.324373f
C428 two_stage_opamp_dummy_magic_23_0.V_err_p.n31 GNDA 0.243876f
C429 two_stage_opamp_dummy_magic_23_0.V_err_p.t10 GNDA 0.023181f
C430 two_stage_opamp_dummy_magic_23_0.V_err_p.t6 GNDA 0.023181f
C431 two_stage_opamp_dummy_magic_23_0.V_err_p.n32 GNDA 0.047234f
C432 two_stage_opamp_dummy_magic_23_0.V_err_p.n33 GNDA 0.324373f
C433 two_stage_opamp_dummy_magic_23_0.V_err_p.n34 GNDA 0.370407f
C434 two_stage_opamp_dummy_magic_23_0.V_err_p.n35 GNDA 0.392203f
C435 two_stage_opamp_dummy_magic_23_0.V_err_p.n36 GNDA 0.047234f
C436 two_stage_opamp_dummy_magic_23_0.V_err_p.t12 GNDA 0.023181f
C437 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t14 GNDA 0.014089f
C438 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t20 GNDA 0.014089f
C439 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t13 GNDA 0.014089f
C440 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t19 GNDA 0.014089f
C441 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t12 GNDA 0.014089f
C442 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t9 GNDA 0.014089f
C443 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t16 GNDA 0.014089f
C444 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t8 GNDA 0.014089f
C445 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t15 GNDA 0.014089f
C446 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t18 GNDA 0.043221f
C447 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n0 GNDA 0.058715f
C448 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n1 GNDA 0.047239f
C449 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n2 GNDA 0.047239f
C450 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n3 GNDA 0.278183f
C451 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n4 GNDA 0.278183f
C452 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n5 GNDA 0.047239f
C453 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n6 GNDA 0.047239f
C454 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n7 GNDA 0.047239f
C455 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n8 GNDA 0.070246f
C456 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t0 GNDA 0.34959f
C457 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t7 GNDA 0.054668f
C458 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t17 GNDA 0.020442f
C459 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n9 GNDA 0.064119f
C460 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t11 GNDA 0.020442f
C461 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n10 GNDA 0.052487f
C462 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t21 GNDA 0.020442f
C463 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n11 GNDA 0.052487f
C464 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t10 GNDA 0.020442f
C465 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n12 GNDA 0.090979f
C466 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n13 GNDA 1.81893f
C467 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t2 GNDA 0.0663f
C468 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t6 GNDA 0.0663f
C469 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n14 GNDA 0.233505f
C470 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t4 GNDA 0.0663f
C471 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t5 GNDA 0.0663f
C472 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n15 GNDA 0.222172f
C473 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n16 GNDA 1.03828f
C474 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t3 GNDA 0.0663f
C475 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.t1 GNDA 0.0663f
C476 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n17 GNDA 0.222172f
C477 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n18 GNDA 0.74245f
C478 two_stage_opamp_dummy_magic_23_0.V_err_amp_ref.n19 GNDA 1.74622f
C479 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t6 GNDA 0.013923f
C480 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t2 GNDA 0.013923f
C481 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n0 GNDA 0.0349f
C482 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t0 GNDA 0.013923f
C483 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t3 GNDA 0.013923f
C484 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n1 GNDA 0.034715f
C485 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n2 GNDA 0.308549f
C486 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t1 GNDA 0.013923f
C487 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t5 GNDA 0.013923f
C488 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n3 GNDA 0.027846f
C489 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n4 GNDA 0.051784f
C490 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t4 GNDA 0.178969f
C491 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n5 GNDA 0.043982f
C492 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n6 GNDA 0.077795f
C493 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t9 GNDA 0.027846f
C494 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t13 GNDA 0.027846f
C495 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n7 GNDA 0.056933f
C496 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n8 GNDA 0.191235f
C497 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t8 GNDA 0.027846f
C498 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t15 GNDA 0.027846f
C499 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n9 GNDA 0.056933f
C500 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n10 GNDA 0.184161f
C501 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n11 GNDA 0.074781f
C502 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n12 GNDA 0.043982f
C503 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t10 GNDA 0.027846f
C504 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t14 GNDA 0.027846f
C505 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n13 GNDA 0.056933f
C506 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n14 GNDA 0.184161f
C507 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n15 GNDA 0.04559f
C508 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t11 GNDA 0.027846f
C509 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t16 GNDA 0.027846f
C510 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n16 GNDA 0.056933f
C511 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n17 GNDA 0.184161f
C512 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n18 GNDA 0.077795f
C513 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t12 GNDA 0.027846f
C514 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.t7 GNDA 0.027846f
C515 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n19 GNDA 0.056933f
C516 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n20 GNDA 0.187799f
C517 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n21 GNDA 0.112537f
C518 two_stage_opamp_dummy_magic_23_0.V_CMFB_S1.n22 GNDA 1.36338f
C519 bgr_11_0.V_CMFB_S1 GNDA 0.945225f
C520 two_stage_opamp_dummy_magic_23_0.VD4.t33 GNDA 0.060801f
C521 two_stage_opamp_dummy_magic_23_0.VD4.t29 GNDA 0.060801f
C522 two_stage_opamp_dummy_magic_23_0.VD4.n0 GNDA 0.154331f
C523 two_stage_opamp_dummy_magic_23_0.VD4.n1 GNDA 0.431096f
C524 two_stage_opamp_dummy_magic_23_0.VD4.t13 GNDA 0.106612f
C525 two_stage_opamp_dummy_magic_23_0.VD4.t12 GNDA 0.216278f
C526 two_stage_opamp_dummy_magic_23_0.VD4.t23 GNDA 0.060801f
C527 two_stage_opamp_dummy_magic_23_0.VD4.t27 GNDA 0.060801f
C528 two_stage_opamp_dummy_magic_23_0.VD4.n2 GNDA 0.154331f
C529 two_stage_opamp_dummy_magic_23_0.VD4.n3 GNDA 0.431096f
C530 two_stage_opamp_dummy_magic_23_0.VD4.t37 GNDA 0.060801f
C531 two_stage_opamp_dummy_magic_23_0.VD4.t19 GNDA 0.060801f
C532 two_stage_opamp_dummy_magic_23_0.VD4.n4 GNDA 0.154331f
C533 two_stage_opamp_dummy_magic_23_0.VD4.n5 GNDA 0.431096f
C534 two_stage_opamp_dummy_magic_23_0.VD4.t31 GNDA 0.060801f
C535 two_stage_opamp_dummy_magic_23_0.VD4.t35 GNDA 0.060801f
C536 two_stage_opamp_dummy_magic_23_0.VD4.n6 GNDA 0.154331f
C537 two_stage_opamp_dummy_magic_23_0.VD4.n7 GNDA 0.431096f
C538 two_stage_opamp_dummy_magic_23_0.VD4.t21 GNDA 0.060801f
C539 two_stage_opamp_dummy_magic_23_0.VD4.t25 GNDA 0.060801f
C540 two_stage_opamp_dummy_magic_23_0.VD4.n8 GNDA 0.154331f
C541 two_stage_opamp_dummy_magic_23_0.VD4.n9 GNDA 0.481515f
C542 two_stage_opamp_dummy_magic_23_0.VD4.t10 GNDA 0.106612f
C543 two_stage_opamp_dummy_magic_23_0.VD4.n10 GNDA 0.316782f
C544 two_stage_opamp_dummy_magic_23_0.VD4.n11 GNDA 0.627403f
C545 two_stage_opamp_dummy_magic_23_0.VD4.t11 GNDA 0.518263f
C546 two_stage_opamp_dummy_magic_23_0.VD4.t20 GNDA 0.406498f
C547 two_stage_opamp_dummy_magic_23_0.VD4.t24 GNDA 0.406498f
C548 two_stage_opamp_dummy_magic_23_0.VD4.t30 GNDA 0.406498f
C549 two_stage_opamp_dummy_magic_23_0.VD4.t34 GNDA 0.406498f
C550 two_stage_opamp_dummy_magic_23_0.VD4.t36 GNDA 0.406498f
C551 two_stage_opamp_dummy_magic_23_0.VD4.t18 GNDA 0.406498f
C552 two_stage_opamp_dummy_magic_23_0.VD4.t22 GNDA 0.406498f
C553 two_stage_opamp_dummy_magic_23_0.VD4.t26 GNDA 0.406498f
C554 two_stage_opamp_dummy_magic_23_0.VD4.t32 GNDA 0.406498f
C555 two_stage_opamp_dummy_magic_23_0.VD4.t28 GNDA 0.406498f
C556 two_stage_opamp_dummy_magic_23_0.VD4.t14 GNDA 0.518263f
C557 two_stage_opamp_dummy_magic_23_0.VD4.t15 GNDA 0.216278f
C558 two_stage_opamp_dummy_magic_23_0.VD4.n12 GNDA 0.627403f
C559 two_stage_opamp_dummy_magic_23_0.VD4.n13 GNDA 0.311031f
C560 two_stage_opamp_dummy_magic_23_0.VD4.n14 GNDA 0.102448f
C561 two_stage_opamp_dummy_magic_23_0.VD4.n15 GNDA 0.065949f
C562 two_stage_opamp_dummy_magic_23_0.VD4.n16 GNDA 0.065949f
C563 two_stage_opamp_dummy_magic_23_0.VD4.t2 GNDA 0.060801f
C564 two_stage_opamp_dummy_magic_23_0.VD4.t16 GNDA 0.060801f
C565 two_stage_opamp_dummy_magic_23_0.VD4.n17 GNDA 0.124375f
C566 two_stage_opamp_dummy_magic_23_0.VD4.n18 GNDA 0.402689f
C567 two_stage_opamp_dummy_magic_23_0.VD4.n19 GNDA 0.112503f
C568 two_stage_opamp_dummy_magic_23_0.VD4.t8 GNDA 0.060801f
C569 two_stage_opamp_dummy_magic_23_0.VD4.t1 GNDA 0.060801f
C570 two_stage_opamp_dummy_magic_23_0.VD4.n20 GNDA 0.124375f
C571 two_stage_opamp_dummy_magic_23_0.VD4.n21 GNDA 0.391692f
C572 two_stage_opamp_dummy_magic_23_0.VD4.n22 GNDA 0.112503f
C573 two_stage_opamp_dummy_magic_23_0.VD4.t6 GNDA 0.060801f
C574 two_stage_opamp_dummy_magic_23_0.VD4.t5 GNDA 0.060801f
C575 two_stage_opamp_dummy_magic_23_0.VD4.n23 GNDA 0.124375f
C576 two_stage_opamp_dummy_magic_23_0.VD4.n24 GNDA 0.391692f
C577 two_stage_opamp_dummy_magic_23_0.VD4.n25 GNDA 0.065949f
C578 two_stage_opamp_dummy_magic_23_0.VD4.n26 GNDA 0.065949f
C579 two_stage_opamp_dummy_magic_23_0.VD4.t3 GNDA 0.060801f
C580 two_stage_opamp_dummy_magic_23_0.VD4.t4 GNDA 0.060801f
C581 two_stage_opamp_dummy_magic_23_0.VD4.n27 GNDA 0.124375f
C582 two_stage_opamp_dummy_magic_23_0.VD4.n28 GNDA 0.391692f
C583 two_stage_opamp_dummy_magic_23_0.VD4.n29 GNDA 0.065949f
C584 two_stage_opamp_dummy_magic_23_0.VD4.t7 GNDA 0.060801f
C585 two_stage_opamp_dummy_magic_23_0.VD4.t0 GNDA 0.060801f
C586 two_stage_opamp_dummy_magic_23_0.VD4.n30 GNDA 0.124375f
C587 two_stage_opamp_dummy_magic_23_0.VD4.n31 GNDA 0.391692f
C588 two_stage_opamp_dummy_magic_23_0.VD4.n32 GNDA 0.112503f
C589 two_stage_opamp_dummy_magic_23_0.VD4.t17 GNDA 0.060801f
C590 two_stage_opamp_dummy_magic_23_0.VD4.t9 GNDA 0.060801f
C591 two_stage_opamp_dummy_magic_23_0.VD4.n33 GNDA 0.124375f
C592 two_stage_opamp_dummy_magic_23_0.VD4.n34 GNDA 0.39719f
C593 two_stage_opamp_dummy_magic_23_0.VD4.n35 GNDA 0.183347f
C594 two_stage_opamp_dummy_magic_23_0.Vb3.t2 GNDA 0.0123f
C595 two_stage_opamp_dummy_magic_23_0.Vb3.t3 GNDA 0.0123f
C596 two_stage_opamp_dummy_magic_23_0.Vb3.n0 GNDA 0.037152f
C597 two_stage_opamp_dummy_magic_23_0.Vb3.t1 GNDA 0.0123f
C598 two_stage_opamp_dummy_magic_23_0.Vb3.t4 GNDA 0.0123f
C599 two_stage_opamp_dummy_magic_23_0.Vb3.n1 GNDA 0.03962f
C600 two_stage_opamp_dummy_magic_23_0.Vb3.t0 GNDA 0.0123f
C601 two_stage_opamp_dummy_magic_23_0.Vb3.t6 GNDA 0.0123f
C602 two_stage_opamp_dummy_magic_23_0.Vb3.n2 GNDA 0.03962f
C603 two_stage_opamp_dummy_magic_23_0.Vb3.n3 GNDA 0.218425f
C604 two_stage_opamp_dummy_magic_23_0.Vb3.n4 GNDA 0.66157f
C605 two_stage_opamp_dummy_magic_23_0.Vb3.t5 GNDA 0.043051f
C606 two_stage_opamp_dummy_magic_23_0.Vb3.t7 GNDA 0.043051f
C607 two_stage_opamp_dummy_magic_23_0.Vb3.n5 GNDA 0.118766f
C608 two_stage_opamp_dummy_magic_23_0.Vb3.t9 GNDA 0.060886f
C609 two_stage_opamp_dummy_magic_23_0.Vb3.t26 GNDA 0.060886f
C610 two_stage_opamp_dummy_magic_23_0.Vb3.t23 GNDA 0.060886f
C611 two_stage_opamp_dummy_magic_23_0.Vb3.t19 GNDA 0.060886f
C612 two_stage_opamp_dummy_magic_23_0.Vb3.t16 GNDA 0.070262f
C613 two_stage_opamp_dummy_magic_23_0.Vb3.n6 GNDA 0.057045f
C614 two_stage_opamp_dummy_magic_23_0.Vb3.n7 GNDA 0.035056f
C615 two_stage_opamp_dummy_magic_23_0.Vb3.n8 GNDA 0.035056f
C616 two_stage_opamp_dummy_magic_23_0.Vb3.n9 GNDA 0.030737f
C617 two_stage_opamp_dummy_magic_23_0.Vb3.t13 GNDA 0.060886f
C618 two_stage_opamp_dummy_magic_23_0.Vb3.t17 GNDA 0.060886f
C619 two_stage_opamp_dummy_magic_23_0.Vb3.t21 GNDA 0.060886f
C620 two_stage_opamp_dummy_magic_23_0.Vb3.t24 GNDA 0.060886f
C621 two_stage_opamp_dummy_magic_23_0.Vb3.t22 GNDA 0.070262f
C622 two_stage_opamp_dummy_magic_23_0.Vb3.n10 GNDA 0.057045f
C623 two_stage_opamp_dummy_magic_23_0.Vb3.n11 GNDA 0.035056f
C624 two_stage_opamp_dummy_magic_23_0.Vb3.n12 GNDA 0.035056f
C625 two_stage_opamp_dummy_magic_23_0.Vb3.n13 GNDA 0.030737f
C626 two_stage_opamp_dummy_magic_23_0.Vb3.n14 GNDA 0.031021f
C627 two_stage_opamp_dummy_magic_23_0.Vb3.t12 GNDA 0.060886f
C628 two_stage_opamp_dummy_magic_23_0.Vb3.t14 GNDA 0.060886f
C629 two_stage_opamp_dummy_magic_23_0.Vb3.t10 GNDA 0.060886f
C630 two_stage_opamp_dummy_magic_23_0.Vb3.t27 GNDA 0.060886f
C631 two_stage_opamp_dummy_magic_23_0.Vb3.t25 GNDA 0.070262f
C632 two_stage_opamp_dummy_magic_23_0.Vb3.n15 GNDA 0.057045f
C633 two_stage_opamp_dummy_magic_23_0.Vb3.n16 GNDA 0.035056f
C634 two_stage_opamp_dummy_magic_23_0.Vb3.n17 GNDA 0.035056f
C635 two_stage_opamp_dummy_magic_23_0.Vb3.n18 GNDA 0.030737f
C636 two_stage_opamp_dummy_magic_23_0.Vb3.t15 GNDA 0.060886f
C637 two_stage_opamp_dummy_magic_23_0.Vb3.t18 GNDA 0.060886f
C638 two_stage_opamp_dummy_magic_23_0.Vb3.t28 GNDA 0.060886f
C639 two_stage_opamp_dummy_magic_23_0.Vb3.t11 GNDA 0.060886f
C640 two_stage_opamp_dummy_magic_23_0.Vb3.t8 GNDA 0.070262f
C641 two_stage_opamp_dummy_magic_23_0.Vb3.n19 GNDA 0.057045f
C642 two_stage_opamp_dummy_magic_23_0.Vb3.n20 GNDA 0.035056f
C643 two_stage_opamp_dummy_magic_23_0.Vb3.n21 GNDA 0.035056f
C644 two_stage_opamp_dummy_magic_23_0.Vb3.n22 GNDA 0.030737f
C645 two_stage_opamp_dummy_magic_23_0.Vb3.n23 GNDA 0.031585f
C646 two_stage_opamp_dummy_magic_23_0.Vb3.n24 GNDA 1.03635f
C647 two_stage_opamp_dummy_magic_23_0.Vb3.t20 GNDA 0.079537f
C648 two_stage_opamp_dummy_magic_23_0.Vb3.n25 GNDA 0.279443f
C649 two_stage_opamp_dummy_magic_23_0.Vb3.n26 GNDA 0.978365f
C650 bgr_11_0.VB3_CUR_BIAS GNDA 1.50184f
C651 bgr_11_0.PFET_GATE_10uA.t27 GNDA 0.020335f
C652 bgr_11_0.PFET_GATE_10uA.t20 GNDA 0.03006f
C653 bgr_11_0.PFET_GATE_10uA.n0 GNDA 0.033123f
C654 bgr_11_0.PFET_GATE_10uA.t14 GNDA 0.020335f
C655 bgr_11_0.PFET_GATE_10uA.t21 GNDA 0.03006f
C656 bgr_11_0.PFET_GATE_10uA.n1 GNDA 0.033123f
C657 bgr_11_0.PFET_GATE_10uA.n2 GNDA 0.039856f
C658 bgr_11_0.PFET_GATE_10uA.t17 GNDA 0.020335f
C659 bgr_11_0.PFET_GATE_10uA.t10 GNDA 0.03006f
C660 bgr_11_0.PFET_GATE_10uA.n3 GNDA 0.033123f
C661 bgr_11_0.PFET_GATE_10uA.t24 GNDA 0.020335f
C662 bgr_11_0.PFET_GATE_10uA.t23 GNDA 0.03006f
C663 bgr_11_0.PFET_GATE_10uA.n4 GNDA 0.033123f
C664 bgr_11_0.PFET_GATE_10uA.n5 GNDA 0.033229f
C665 bgr_11_0.PFET_GATE_10uA.t2 GNDA 0.304654f
C666 bgr_11_0.PFET_GATE_10uA.t3 GNDA 0.020856f
C667 bgr_11_0.PFET_GATE_10uA.t0 GNDA 0.020856f
C668 bgr_11_0.PFET_GATE_10uA.n6 GNDA 0.053306f
C669 bgr_11_0.PFET_GATE_10uA.t5 GNDA 0.020856f
C670 bgr_11_0.PFET_GATE_10uA.t7 GNDA 0.020856f
C671 bgr_11_0.PFET_GATE_10uA.n7 GNDA 0.051929f
C672 bgr_11_0.PFET_GATE_10uA.n8 GNDA 0.507929f
C673 bgr_11_0.PFET_GATE_10uA.t6 GNDA 0.020856f
C674 bgr_11_0.PFET_GATE_10uA.t8 GNDA 0.020856f
C675 bgr_11_0.PFET_GATE_10uA.n9 GNDA 0.051929f
C676 bgr_11_0.PFET_GATE_10uA.n10 GNDA 0.288022f
C677 bgr_11_0.PFET_GATE_10uA.n11 GNDA 0.587978f
C678 bgr_11_0.PFET_GATE_10uA.t1 GNDA 0.020856f
C679 bgr_11_0.PFET_GATE_10uA.t4 GNDA 0.020856f
C680 bgr_11_0.PFET_GATE_10uA.n12 GNDA 0.0503f
C681 bgr_11_0.PFET_GATE_10uA.n13 GNDA 0.268525f
C682 bgr_11_0.PFET_GATE_10uA.t9 GNDA 0.453343f
C683 bgr_11_0.PFET_GATE_10uA.t26 GNDA 0.023511f
C684 bgr_11_0.PFET_GATE_10uA.t13 GNDA 0.023511f
C685 bgr_11_0.PFET_GATE_10uA.n14 GNDA 0.067972f
C686 bgr_11_0.PFET_GATE_10uA.n15 GNDA 1.8717f
C687 bgr_11_0.PFET_GATE_10uA.n16 GNDA 0.75222f
C688 bgr_11_0.PFET_GATE_10uA.n17 GNDA 0.740244f
C689 bgr_11_0.PFET_GATE_10uA.t29 GNDA 0.020335f
C690 bgr_11_0.PFET_GATE_10uA.t19 GNDA 0.020335f
C691 bgr_11_0.PFET_GATE_10uA.t12 GNDA 0.020335f
C692 bgr_11_0.PFET_GATE_10uA.t25 GNDA 0.020335f
C693 bgr_11_0.PFET_GATE_10uA.t18 GNDA 0.020335f
C694 bgr_11_0.PFET_GATE_10uA.t11 GNDA 0.03006f
C695 bgr_11_0.PFET_GATE_10uA.n18 GNDA 0.037201f
C696 bgr_11_0.PFET_GATE_10uA.n19 GNDA 0.026591f
C697 bgr_11_0.PFET_GATE_10uA.n20 GNDA 0.026591f
C698 bgr_11_0.PFET_GATE_10uA.n21 GNDA 0.026591f
C699 bgr_11_0.PFET_GATE_10uA.n22 GNDA 0.022513f
C700 bgr_11_0.PFET_GATE_10uA.t16 GNDA 0.020335f
C701 bgr_11_0.PFET_GATE_10uA.t15 GNDA 0.020335f
C702 bgr_11_0.PFET_GATE_10uA.t22 GNDA 0.020335f
C703 bgr_11_0.PFET_GATE_10uA.t28 GNDA 0.03006f
C704 bgr_11_0.PFET_GATE_10uA.n23 GNDA 0.037201f
C705 bgr_11_0.PFET_GATE_10uA.n24 GNDA 0.026591f
C706 bgr_11_0.PFET_GATE_10uA.n25 GNDA 0.022513f
C707 bgr_11_0.PFET_GATE_10uA.n26 GNDA 0.030903f
C708 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t0 GNDA 0.013958f
C709 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t13 GNDA 0.013958f
C710 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n0 GNDA 0.035002f
C711 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t16 GNDA 0.013958f
C712 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t1 GNDA 0.013958f
C713 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n1 GNDA 0.034818f
C714 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n2 GNDA 0.309517f
C715 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t12 GNDA 0.013958f
C716 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t15 GNDA 0.013958f
C717 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n3 GNDA 0.027915f
C718 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n4 GNDA 0.051892f
C719 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t14 GNDA 0.178492f
C720 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n5 GNDA 0.044092f
C721 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n6 GNDA 0.077991f
C722 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t3 GNDA 0.027915f
C723 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t7 GNDA 0.027915f
C724 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n7 GNDA 0.057076f
C725 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n8 GNDA 0.191716f
C726 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t2 GNDA 0.027915f
C727 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t10 GNDA 0.027915f
C728 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n9 GNDA 0.057076f
C729 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n10 GNDA 0.184623f
C730 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n11 GNDA 0.074969f
C731 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n12 GNDA 0.044092f
C732 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t5 GNDA 0.027915f
C733 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t9 GNDA 0.027915f
C734 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n13 GNDA 0.057076f
C735 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n14 GNDA 0.184623f
C736 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n15 GNDA 0.045704f
C737 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t4 GNDA 0.027915f
C738 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t8 GNDA 0.027915f
C739 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n16 GNDA 0.057076f
C740 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n17 GNDA 0.184623f
C741 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n18 GNDA 0.077991f
C742 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t11 GNDA 0.027915f
C743 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.t6 GNDA 0.027915f
C744 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n19 GNDA 0.057076f
C745 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n20 GNDA 0.188271f
C746 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n21 GNDA 0.113808f
C747 two_stage_opamp_dummy_magic_23_0.V_CMFB_S3.n22 GNDA 1.35418f
C748 bgr_11_0.V_CMFB_S3 GNDA 0.947399f
C749 bgr_11_0.Vin-.n0 GNDA 0.069747f
C750 bgr_11_0.Vin-.n1 GNDA 0.316148f
C751 bgr_11_0.Vin-.t7 GNDA 0.027101f
C752 bgr_11_0.Vin-.t4 GNDA 0.027101f
C753 bgr_11_0.Vin-.n2 GNDA 0.094346f
C754 bgr_11_0.Vin-.t5 GNDA 0.027101f
C755 bgr_11_0.Vin-.t6 GNDA 0.027101f
C756 bgr_11_0.Vin-.n3 GNDA 0.090091f
C757 bgr_11_0.Vin-.n4 GNDA 0.386489f
C758 bgr_11_0.Vin-.n5 GNDA 0.027681f
C759 bgr_11_0.Vin-.n6 GNDA 0.366254f
C760 bgr_11_0.Vin-.t10 GNDA 0.022346f
C761 bgr_11_0.Vin-.n7 GNDA 0.026209f
C762 bgr_11_0.Vin-.n8 GNDA 0.021455f
C763 bgr_11_0.Vin-.n9 GNDA 0.021455f
C764 bgr_11_0.Vin-.n10 GNDA 0.036491f
C765 bgr_11_0.Vin-.n11 GNDA 0.497932f
C766 bgr_11_0.Vin-.t0 GNDA 0.117924f
C767 bgr_11_0.Vin-.n12 GNDA 0.655831f
C768 bgr_11_0.Vin-.n13 GNDA 1.07297f
C769 bgr_11_0.Vin-.n14 GNDA 0.471323f
C770 bgr_11_0.Vin-.t3 GNDA 0.261631f
C771 bgr_11_0.Vin-.n15 GNDA 0.069875f
C772 bgr_11_0.Vin-.n16 GNDA 0.119593f
C773 bgr_11_0.Vin-.n17 GNDA 0.07053f
C774 bgr_11_0.Vin-.n18 GNDA 0.579028f
C775 bgr_11_0.Vin-.n19 GNDA 0.358216f
C776 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter GNDA 0.086538f
C777 bgr_11_0.V_TOP.t24 GNDA 0.098487f
C778 bgr_11_0.V_TOP.t36 GNDA 0.098487f
C779 bgr_11_0.V_TOP.t41 GNDA 0.098487f
C780 bgr_11_0.V_TOP.t14 GNDA 0.098487f
C781 bgr_11_0.V_TOP.t49 GNDA 0.098487f
C782 bgr_11_0.V_TOP.t25 GNDA 0.098487f
C783 bgr_11_0.V_TOP.t37 GNDA 0.098487f
C784 bgr_11_0.V_TOP.t43 GNDA 0.098487f
C785 bgr_11_0.V_TOP.t19 GNDA 0.098487f
C786 bgr_11_0.V_TOP.t16 GNDA 0.098487f
C787 bgr_11_0.V_TOP.t30 GNDA 0.098487f
C788 bgr_11_0.V_TOP.t40 GNDA 0.098487f
C789 bgr_11_0.V_TOP.t48 GNDA 0.098487f
C790 bgr_11_0.V_TOP.t29 GNDA 0.098487f
C791 bgr_11_0.V_TOP.t26 GNDA 0.128747f
C792 bgr_11_0.V_TOP.n0 GNDA 0.071979f
C793 bgr_11_0.V_TOP.n1 GNDA 0.052527f
C794 bgr_11_0.V_TOP.n2 GNDA 0.052527f
C795 bgr_11_0.V_TOP.n3 GNDA 0.052527f
C796 bgr_11_0.V_TOP.n4 GNDA 0.052527f
C797 bgr_11_0.V_TOP.n5 GNDA 0.048982f
C798 bgr_11_0.V_TOP.t7 GNDA 0.126654f
C799 bgr_11_0.V_TOP.t46 GNDA 0.37519f
C800 bgr_11_0.V_TOP.t34 GNDA 0.38158f
C801 bgr_11_0.V_TOP.t39 GNDA 0.37519f
C802 bgr_11_0.V_TOP.n6 GNDA 0.251553f
C803 bgr_11_0.V_TOP.t32 GNDA 0.37519f
C804 bgr_11_0.V_TOP.t21 GNDA 0.38158f
C805 bgr_11_0.V_TOP.n7 GNDA 0.321901f
C806 bgr_11_0.V_TOP.t23 GNDA 0.38158f
C807 bgr_11_0.V_TOP.t31 GNDA 0.37519f
C808 bgr_11_0.V_TOP.n8 GNDA 0.251553f
C809 bgr_11_0.V_TOP.t20 GNDA 0.37519f
C810 bgr_11_0.V_TOP.t45 GNDA 0.38158f
C811 bgr_11_0.V_TOP.n9 GNDA 0.392249f
C812 bgr_11_0.V_TOP.t33 GNDA 0.38158f
C813 bgr_11_0.V_TOP.t38 GNDA 0.37519f
C814 bgr_11_0.V_TOP.n10 GNDA 0.251553f
C815 bgr_11_0.V_TOP.t28 GNDA 0.37519f
C816 bgr_11_0.V_TOP.t18 GNDA 0.38158f
C817 bgr_11_0.V_TOP.n11 GNDA 0.392249f
C818 bgr_11_0.V_TOP.t22 GNDA 0.38158f
C819 bgr_11_0.V_TOP.t27 GNDA 0.37519f
C820 bgr_11_0.V_TOP.n12 GNDA 0.251553f
C821 bgr_11_0.V_TOP.t17 GNDA 0.37519f
C822 bgr_11_0.V_TOP.t44 GNDA 0.38158f
C823 bgr_11_0.V_TOP.n13 GNDA 0.392249f
C824 bgr_11_0.V_TOP.t35 GNDA 0.38158f
C825 bgr_11_0.V_TOP.t42 GNDA 0.37519f
C826 bgr_11_0.V_TOP.n14 GNDA 0.321901f
C827 bgr_11_0.V_TOP.t15 GNDA 0.37519f
C828 bgr_11_0.V_TOP.n15 GNDA 0.164146f
C829 bgr_11_0.V_TOP.n16 GNDA 0.561746f
C830 bgr_11_0.V_TOP.t0 GNDA 0.105546f
C831 bgr_11_0.V_TOP.n17 GNDA 0.747366f
C832 bgr_11_0.V_TOP.n18 GNDA 0.023355f
C833 bgr_11_0.V_TOP.n19 GNDA 0.427854f
C834 bgr_11_0.V_TOP.n20 GNDA 0.022622f
C835 bgr_11_0.V_TOP.n21 GNDA 0.023512f
C836 bgr_11_0.V_TOP.n22 GNDA 0.023355f
C837 bgr_11_0.V_TOP.n23 GNDA 0.216436f
C838 bgr_11_0.V_TOP.n24 GNDA 0.131474f
C839 bgr_11_0.V_TOP.n25 GNDA 0.075038f
C840 bgr_11_0.V_TOP.n26 GNDA 0.023355f
C841 bgr_11_0.V_TOP.n27 GNDA 0.129535f
C842 bgr_11_0.V_TOP.n28 GNDA 0.023355f
C843 bgr_11_0.V_TOP.n29 GNDA 0.128304f
C844 bgr_11_0.V_TOP.n30 GNDA 0.282032f
C845 bgr_11_0.V_TOP.n31 GNDA 0.019847f
C846 bgr_11_0.V_TOP.n32 GNDA 0.048982f
C847 bgr_11_0.V_TOP.n33 GNDA 0.052527f
C848 bgr_11_0.V_TOP.n34 GNDA 0.052527f
C849 bgr_11_0.V_TOP.n35 GNDA 0.052527f
C850 bgr_11_0.V_TOP.n36 GNDA 0.052527f
C851 bgr_11_0.V_TOP.n37 GNDA 0.052527f
C852 bgr_11_0.V_TOP.n38 GNDA 0.052527f
C853 bgr_11_0.V_TOP.n39 GNDA 0.048982f
C854 bgr_11_0.V_TOP.t47 GNDA 0.113492f
C855 bgr_11_0.V_mir2.t10 GNDA 0.019544f
C856 bgr_11_0.V_mir2.n0 GNDA 0.025551f
C857 bgr_11_0.V_mir2.t15 GNDA 0.041699f
C858 bgr_11_0.V_mir2.n1 GNDA 0.027738f
C859 bgr_11_0.V_mir2.n2 GNDA 0.457418f
C860 bgr_11_0.V_mir2.n3 GNDA 0.148244f
C861 bgr_11_0.V_mir2.t7 GNDA 0.023453f
C862 bgr_11_0.V_mir2.t22 GNDA 0.023453f
C863 bgr_11_0.V_mir2.t19 GNDA 0.037856f
C864 bgr_11_0.V_mir2.n4 GNDA 0.042274f
C865 bgr_11_0.V_mir2.n5 GNDA 0.028879f
C866 bgr_11_0.V_mir2.t3 GNDA 0.029773f
C867 bgr_11_0.V_mir2.n6 GNDA 0.044932f
C868 bgr_11_0.V_mir2.t8 GNDA 0.019544f
C869 bgr_11_0.V_mir2.t4 GNDA 0.019544f
C870 bgr_11_0.V_mir2.n7 GNDA 0.044741f
C871 bgr_11_0.V_mir2.n8 GNDA 0.11173f
C872 bgr_11_0.V_mir2.t5 GNDA 0.023453f
C873 bgr_11_0.V_mir2.t17 GNDA 0.023453f
C874 bgr_11_0.V_mir2.t21 GNDA 0.037856f
C875 bgr_11_0.V_mir2.n9 GNDA 0.042274f
C876 bgr_11_0.V_mir2.n10 GNDA 0.028879f
C877 bgr_11_0.V_mir2.t11 GNDA 0.029773f
C878 bgr_11_0.V_mir2.n11 GNDA 0.044932f
C879 bgr_11_0.V_mir2.t6 GNDA 0.019544f
C880 bgr_11_0.V_mir2.t12 GNDA 0.019544f
C881 bgr_11_0.V_mir2.n12 GNDA 0.044741f
C882 bgr_11_0.V_mir2.n13 GNDA 0.11173f
C883 bgr_11_0.V_mir2.n14 GNDA 0.355461f
C884 bgr_11_0.V_mir2.n15 GNDA 0.051792f
C885 bgr_11_0.V_mir2.t9 GNDA 0.023453f
C886 bgr_11_0.V_mir2.t18 GNDA 0.023453f
C887 bgr_11_0.V_mir2.t20 GNDA 0.037856f
C888 bgr_11_0.V_mir2.n16 GNDA 0.042274f
C889 bgr_11_0.V_mir2.n17 GNDA 0.028879f
C890 bgr_11_0.V_mir2.t13 GNDA 0.029773f
C891 bgr_11_0.V_mir2.n18 GNDA 0.044932f
C892 bgr_11_0.V_mir2.n19 GNDA 0.086204f
C893 bgr_11_0.V_mir2.n20 GNDA 0.044741f
C894 bgr_11_0.V_mir2.t14 GNDA 0.019544f
C895 two_stage_opamp_dummy_magic_23_0.V_source.t15 GNDA 0.038168f
C896 two_stage_opamp_dummy_magic_23_0.V_source.n0 GNDA 0.052428f
C897 two_stage_opamp_dummy_magic_23_0.V_source.n1 GNDA 0.05567f
C898 two_stage_opamp_dummy_magic_23_0.V_source.n2 GNDA 0.052428f
C899 two_stage_opamp_dummy_magic_23_0.V_source.n3 GNDA 0.096361f
C900 two_stage_opamp_dummy_magic_23_0.V_source.t37 GNDA 0.022901f
C901 two_stage_opamp_dummy_magic_23_0.V_source.t26 GNDA 0.022901f
C902 two_stage_opamp_dummy_magic_23_0.V_source.n4 GNDA 0.049829f
C903 two_stage_opamp_dummy_magic_23_0.V_source.n5 GNDA 0.153174f
C904 two_stage_opamp_dummy_magic_23_0.V_source.n6 GNDA 0.051154f
C905 two_stage_opamp_dummy_magic_23_0.V_source.t31 GNDA 0.022901f
C906 two_stage_opamp_dummy_magic_23_0.V_source.t6 GNDA 0.022901f
C907 two_stage_opamp_dummy_magic_23_0.V_source.n7 GNDA 0.049829f
C908 two_stage_opamp_dummy_magic_23_0.V_source.n8 GNDA 0.200044f
C909 two_stage_opamp_dummy_magic_23_0.V_source.n9 GNDA 0.087575f
C910 two_stage_opamp_dummy_magic_23_0.V_source.t34 GNDA 0.022901f
C911 two_stage_opamp_dummy_magic_23_0.V_source.t32 GNDA 0.022901f
C912 two_stage_opamp_dummy_magic_23_0.V_source.n10 GNDA 0.049829f
C913 two_stage_opamp_dummy_magic_23_0.V_source.n11 GNDA 0.192055f
C914 two_stage_opamp_dummy_magic_23_0.V_source.n12 GNDA 0.083262f
C915 two_stage_opamp_dummy_magic_23_0.V_source.t5 GNDA 0.022901f
C916 two_stage_opamp_dummy_magic_23_0.V_source.t7 GNDA 0.022901f
C917 two_stage_opamp_dummy_magic_23_0.V_source.n13 GNDA 0.049829f
C918 two_stage_opamp_dummy_magic_23_0.V_source.n14 GNDA 0.192055f
C919 two_stage_opamp_dummy_magic_23_0.V_source.n15 GNDA 0.048946f
C920 two_stage_opamp_dummy_magic_23_0.V_source.n16 GNDA 0.083262f
C921 two_stage_opamp_dummy_magic_23_0.V_source.t0 GNDA 0.022901f
C922 two_stage_opamp_dummy_magic_23_0.V_source.t28 GNDA 0.022901f
C923 two_stage_opamp_dummy_magic_23_0.V_source.n17 GNDA 0.049829f
C924 two_stage_opamp_dummy_magic_23_0.V_source.n18 GNDA 0.192055f
C925 two_stage_opamp_dummy_magic_23_0.V_source.n19 GNDA 0.051154f
C926 two_stage_opamp_dummy_magic_23_0.V_source.n20 GNDA 0.051154f
C927 two_stage_opamp_dummy_magic_23_0.V_source.n21 GNDA 0.083262f
C928 two_stage_opamp_dummy_magic_23_0.V_source.t35 GNDA 0.022901f
C929 two_stage_opamp_dummy_magic_23_0.V_source.t3 GNDA 0.022901f
C930 two_stage_opamp_dummy_magic_23_0.V_source.n22 GNDA 0.049829f
C931 two_stage_opamp_dummy_magic_23_0.V_source.n23 GNDA 0.200044f
C932 two_stage_opamp_dummy_magic_23_0.V_source.t38 GNDA 0.022901f
C933 two_stage_opamp_dummy_magic_23_0.V_source.t39 GNDA 0.022901f
C934 two_stage_opamp_dummy_magic_23_0.V_source.n24 GNDA 0.049829f
C935 two_stage_opamp_dummy_magic_23_0.V_source.n25 GNDA 0.192055f
C936 two_stage_opamp_dummy_magic_23_0.V_source.n26 GNDA 0.087575f
C937 two_stage_opamp_dummy_magic_23_0.V_source.n27 GNDA 0.051154f
C938 two_stage_opamp_dummy_magic_23_0.V_source.t33 GNDA 0.022901f
C939 two_stage_opamp_dummy_magic_23_0.V_source.t4 GNDA 0.022901f
C940 two_stage_opamp_dummy_magic_23_0.V_source.n28 GNDA 0.049829f
C941 two_stage_opamp_dummy_magic_23_0.V_source.n29 GNDA 0.192055f
C942 two_stage_opamp_dummy_magic_23_0.V_source.n30 GNDA 0.048946f
C943 two_stage_opamp_dummy_magic_23_0.V_source.t30 GNDA 0.022901f
C944 two_stage_opamp_dummy_magic_23_0.V_source.t1 GNDA 0.022901f
C945 two_stage_opamp_dummy_magic_23_0.V_source.n31 GNDA 0.049829f
C946 two_stage_opamp_dummy_magic_23_0.V_source.n32 GNDA 0.192055f
C947 two_stage_opamp_dummy_magic_23_0.V_source.n33 GNDA 0.083262f
C948 two_stage_opamp_dummy_magic_23_0.V_source.t29 GNDA 0.022901f
C949 two_stage_opamp_dummy_magic_23_0.V_source.t27 GNDA 0.022901f
C950 two_stage_opamp_dummy_magic_23_0.V_source.n34 GNDA 0.049829f
C951 two_stage_opamp_dummy_magic_23_0.V_source.n35 GNDA 0.195998f
C952 two_stage_opamp_dummy_magic_23_0.V_source.n36 GNDA 0.125964f
C953 two_stage_opamp_dummy_magic_23_0.V_source.n37 GNDA 0.120611f
C954 two_stage_opamp_dummy_magic_23_0.V_source.n38 GNDA 0.087586f
C955 two_stage_opamp_dummy_magic_23_0.V_source.t36 GNDA 0.038168f
C956 two_stage_opamp_dummy_magic_23_0.V_source.t2 GNDA 0.038168f
C957 two_stage_opamp_dummy_magic_23_0.V_source.n39 GNDA 0.081597f
C958 two_stage_opamp_dummy_magic_23_0.V_source.n40 GNDA 0.294282f
C959 two_stage_opamp_dummy_magic_23_0.V_source.t18 GNDA 0.038168f
C960 two_stage_opamp_dummy_magic_23_0.V_source.t22 GNDA 0.038168f
C961 two_stage_opamp_dummy_magic_23_0.V_source.n41 GNDA 0.081597f
C962 two_stage_opamp_dummy_magic_23_0.V_source.n42 GNDA 0.285878f
C963 two_stage_opamp_dummy_magic_23_0.V_source.n43 GNDA 0.090055f
C964 two_stage_opamp_dummy_magic_23_0.V_source.n44 GNDA 0.045802f
C965 two_stage_opamp_dummy_magic_23_0.V_source.n45 GNDA 0.099442f
C966 two_stage_opamp_dummy_magic_23_0.V_source.t12 GNDA 0.038168f
C967 two_stage_opamp_dummy_magic_23_0.V_source.t20 GNDA 0.038168f
C968 two_stage_opamp_dummy_magic_23_0.V_source.n46 GNDA 0.081597f
C969 two_stage_opamp_dummy_magic_23_0.V_source.n47 GNDA 0.185859f
C970 two_stage_opamp_dummy_magic_23_0.V_source.t40 GNDA 0.079851f
C971 two_stage_opamp_dummy_magic_23_0.V_source.n48 GNDA 0.258116f
C972 two_stage_opamp_dummy_magic_23_0.V_source.n49 GNDA 0.045802f
C973 two_stage_opamp_dummy_magic_23_0.V_source.t10 GNDA 0.038168f
C974 two_stage_opamp_dummy_magic_23_0.V_source.t19 GNDA 0.038168f
C975 two_stage_opamp_dummy_magic_23_0.V_source.n50 GNDA 0.081597f
C976 two_stage_opamp_dummy_magic_23_0.V_source.n51 GNDA 0.285878f
C977 two_stage_opamp_dummy_magic_23_0.V_source.n52 GNDA 0.05567f
C978 two_stage_opamp_dummy_magic_23_0.V_source.n53 GNDA 0.05567f
C979 two_stage_opamp_dummy_magic_23_0.V_source.t9 GNDA 0.038168f
C980 two_stage_opamp_dummy_magic_23_0.V_source.t17 GNDA 0.038168f
C981 two_stage_opamp_dummy_magic_23_0.V_source.n54 GNDA 0.081597f
C982 two_stage_opamp_dummy_magic_23_0.V_source.n55 GNDA 0.285878f
C983 two_stage_opamp_dummy_magic_23_0.V_source.n56 GNDA 0.052428f
C984 two_stage_opamp_dummy_magic_23_0.V_source.t8 GNDA 0.038168f
C985 two_stage_opamp_dummy_magic_23_0.V_source.t23 GNDA 0.038168f
C986 two_stage_opamp_dummy_magic_23_0.V_source.n57 GNDA 0.081597f
C987 two_stage_opamp_dummy_magic_23_0.V_source.n58 GNDA 0.285878f
C988 two_stage_opamp_dummy_magic_23_0.V_source.n59 GNDA 0.052428f
C989 two_stage_opamp_dummy_magic_23_0.V_source.n60 GNDA 0.052428f
C990 two_stage_opamp_dummy_magic_23_0.V_source.t13 GNDA 0.038168f
C991 two_stage_opamp_dummy_magic_23_0.V_source.t16 GNDA 0.038168f
C992 two_stage_opamp_dummy_magic_23_0.V_source.n61 GNDA 0.081597f
C993 two_stage_opamp_dummy_magic_23_0.V_source.n62 GNDA 0.285878f
C994 two_stage_opamp_dummy_magic_23_0.V_source.n63 GNDA 0.05567f
C995 two_stage_opamp_dummy_magic_23_0.V_source.t21 GNDA 0.038168f
C996 two_stage_opamp_dummy_magic_23_0.V_source.t11 GNDA 0.038168f
C997 two_stage_opamp_dummy_magic_23_0.V_source.n64 GNDA 0.081597f
C998 two_stage_opamp_dummy_magic_23_0.V_source.n65 GNDA 0.294282f
C999 two_stage_opamp_dummy_magic_23_0.V_source.n66 GNDA 0.090055f
C1000 two_stage_opamp_dummy_magic_23_0.V_source.t24 GNDA 0.038168f
C1001 two_stage_opamp_dummy_magic_23_0.V_source.t14 GNDA 0.038168f
C1002 two_stage_opamp_dummy_magic_23_0.V_source.n67 GNDA 0.081597f
C1003 two_stage_opamp_dummy_magic_23_0.V_source.n68 GNDA 0.285878f
C1004 two_stage_opamp_dummy_magic_23_0.V_source.n69 GNDA 0.096361f
C1005 two_stage_opamp_dummy_magic_23_0.V_source.n70 GNDA 0.05567f
C1006 two_stage_opamp_dummy_magic_23_0.V_source.n71 GNDA 0.285878f
C1007 two_stage_opamp_dummy_magic_23_0.V_source.n72 GNDA 0.081597f
C1008 two_stage_opamp_dummy_magic_23_0.V_source.t25 GNDA 0.038168f
C1009 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t1 GNDA 0.01412f
C1010 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t5 GNDA 0.01412f
C1011 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n0 GNDA 0.035347f
C1012 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t2 GNDA 0.01412f
C1013 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t4 GNDA 0.01412f
C1014 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n1 GNDA 0.035347f
C1015 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t11 GNDA 0.01412f
C1016 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t10 GNDA 0.01412f
C1017 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n2 GNDA 0.035158f
C1018 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n3 GNDA 0.238729f
C1019 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n4 GNDA 0.200523f
C1020 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t3 GNDA 0.01412f
C1021 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t9 GNDA 0.01412f
C1022 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n5 GNDA 0.028241f
C1023 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n6 GNDA 0.050138f
C1024 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t6 GNDA 0.021181f
C1025 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t7 GNDA 0.021181f
C1026 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n7 GNDA 0.04919f
C1027 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t14 GNDA 0.037595f
C1028 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t31 GNDA 0.037595f
C1029 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t20 GNDA 0.037595f
C1030 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t29 GNDA 0.037595f
C1031 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t18 GNDA 0.037595f
C1032 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t28 GNDA 0.037595f
C1033 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t17 GNDA 0.037595f
C1034 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t26 GNDA 0.037595f
C1035 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t15 GNDA 0.037595f
C1036 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t19 GNDA 0.04388f
C1037 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n8 GNDA 0.041372f
C1038 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n9 GNDA 0.025946f
C1039 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n10 GNDA 0.025946f
C1040 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n11 GNDA 0.025946f
C1041 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n12 GNDA 0.025946f
C1042 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n13 GNDA 0.025946f
C1043 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n14 GNDA 0.025946f
C1044 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n15 GNDA 0.025946f
C1045 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n16 GNDA 0.023185f
C1046 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t25 GNDA 0.037595f
C1047 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t22 GNDA 0.037595f
C1048 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t12 GNDA 0.037595f
C1049 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t23 GNDA 0.037595f
C1050 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t13 GNDA 0.037595f
C1051 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t24 GNDA 0.037595f
C1052 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t16 GNDA 0.037595f
C1053 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t27 GNDA 0.037595f
C1054 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t30 GNDA 0.037595f
C1055 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t21 GNDA 0.04388f
C1056 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n17 GNDA 0.041372f
C1057 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n18 GNDA 0.025946f
C1058 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n19 GNDA 0.025946f
C1059 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n20 GNDA 0.025946f
C1060 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n21 GNDA 0.025946f
C1061 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n22 GNDA 0.025946f
C1062 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n23 GNDA 0.025946f
C1063 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n24 GNDA 0.025946f
C1064 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n25 GNDA 0.023185f
C1065 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n26 GNDA 0.019627f
C1066 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n27 GNDA 0.296199f
C1067 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t8 GNDA 0.021181f
C1068 two_stage_opamp_dummy_magic_23_0.V_tail_gate.t0 GNDA 0.021181f
C1069 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n28 GNDA 0.046086f
C1070 two_stage_opamp_dummy_magic_23_0.V_tail_gate.n29 GNDA 0.208228f
C1071 two_stage_opamp_dummy_magic_23_0.VD2.t19 GNDA 0.053331f
C1072 two_stage_opamp_dummy_magic_23_0.VD2.t14 GNDA 0.053331f
C1073 two_stage_opamp_dummy_magic_23_0.VD2.n0 GNDA 0.116042f
C1074 two_stage_opamp_dummy_magic_23_0.VD2.n1 GNDA 0.361396f
C1075 two_stage_opamp_dummy_magic_23_0.VD2.n2 GNDA 0.192793f
C1076 two_stage_opamp_dummy_magic_23_0.VD2.t16 GNDA 0.053331f
C1077 two_stage_opamp_dummy_magic_23_0.VD2.t12 GNDA 0.053331f
C1078 two_stage_opamp_dummy_magic_23_0.VD2.n3 GNDA 0.116042f
C1079 two_stage_opamp_dummy_magic_23_0.VD2.n4 GNDA 0.461069f
C1080 two_stage_opamp_dummy_magic_23_0.VD2.t20 GNDA 0.053331f
C1081 two_stage_opamp_dummy_magic_23_0.VD2.t15 GNDA 0.053331f
C1082 two_stage_opamp_dummy_magic_23_0.VD2.n5 GNDA 0.116042f
C1083 two_stage_opamp_dummy_magic_23_0.VD2.n6 GNDA 0.461069f
C1084 two_stage_opamp_dummy_magic_23_0.VD2.t18 GNDA 0.053331f
C1085 two_stage_opamp_dummy_magic_23_0.VD2.t21 GNDA 0.053331f
C1086 two_stage_opamp_dummy_magic_23_0.VD2.n7 GNDA 0.116042f
C1087 two_stage_opamp_dummy_magic_23_0.VD2.n8 GNDA 0.442486f
C1088 two_stage_opamp_dummy_magic_23_0.VD2.n9 GNDA 0.203944f
C1089 two_stage_opamp_dummy_magic_23_0.VD2.n10 GNDA 0.119128f
C1090 two_stage_opamp_dummy_magic_23_0.VD2.n11 GNDA 0.203944f
C1091 two_stage_opamp_dummy_magic_23_0.VD2.t17 GNDA 0.053331f
C1092 two_stage_opamp_dummy_magic_23_0.VD2.t13 GNDA 0.053331f
C1093 two_stage_opamp_dummy_magic_23_0.VD2.n12 GNDA 0.116042f
C1094 two_stage_opamp_dummy_magic_23_0.VD2.n13 GNDA 0.442486f
C1095 two_stage_opamp_dummy_magic_23_0.VD2.n14 GNDA 0.192793f
C1096 two_stage_opamp_dummy_magic_23_0.VD2.n15 GNDA 0.106662f
C1097 two_stage_opamp_dummy_magic_23_0.VD2.n16 GNDA 0.122513f
C1098 two_stage_opamp_dummy_magic_23_0.VD2.n17 GNDA 0.099935f
C1099 two_stage_opamp_dummy_magic_23_0.VD2.n18 GNDA 0.205342f
C1100 two_stage_opamp_dummy_magic_23_0.VD2.t8 GNDA 0.053331f
C1101 two_stage_opamp_dummy_magic_23_0.VD2.t4 GNDA 0.053331f
C1102 two_stage_opamp_dummy_magic_23_0.VD2.n19 GNDA 0.116042f
C1103 two_stage_opamp_dummy_magic_23_0.VD2.n20 GNDA 0.465721f
C1104 two_stage_opamp_dummy_magic_23_0.VD2.n21 GNDA 0.205342f
C1105 two_stage_opamp_dummy_magic_23_0.VD2.t3 GNDA 0.053331f
C1106 two_stage_opamp_dummy_magic_23_0.VD2.t5 GNDA 0.053331f
C1107 two_stage_opamp_dummy_magic_23_0.VD2.n22 GNDA 0.116042f
C1108 two_stage_opamp_dummy_magic_23_0.VD2.n23 GNDA 0.447102f
C1109 two_stage_opamp_dummy_magic_23_0.VD2.n24 GNDA 0.192793f
C1110 two_stage_opamp_dummy_magic_23_0.VD2.t0 GNDA 0.053331f
C1111 two_stage_opamp_dummy_magic_23_0.VD2.t6 GNDA 0.053331f
C1112 two_stage_opamp_dummy_magic_23_0.VD2.n25 GNDA 0.116042f
C1113 two_stage_opamp_dummy_magic_23_0.VD2.n26 GNDA 0.447102f
C1114 two_stage_opamp_dummy_magic_23_0.VD2.n27 GNDA 0.113419f
C1115 two_stage_opamp_dummy_magic_23_0.VD2.t1 GNDA 0.053331f
C1116 two_stage_opamp_dummy_magic_23_0.VD2.t9 GNDA 0.053331f
C1117 two_stage_opamp_dummy_magic_23_0.VD2.n28 GNDA 0.116042f
C1118 two_stage_opamp_dummy_magic_23_0.VD2.n29 GNDA 0.465721f
C1119 two_stage_opamp_dummy_magic_23_0.VD2.t11 GNDA 0.053331f
C1120 two_stage_opamp_dummy_magic_23_0.VD2.t7 GNDA 0.053331f
C1121 two_stage_opamp_dummy_magic_23_0.VD2.n30 GNDA 0.116042f
C1122 two_stage_opamp_dummy_magic_23_0.VD2.n31 GNDA 0.447102f
C1123 two_stage_opamp_dummy_magic_23_0.VD2.n32 GNDA 0.192793f
C1124 two_stage_opamp_dummy_magic_23_0.VD2.n33 GNDA 0.113419f
C1125 two_stage_opamp_dummy_magic_23_0.VD2.t2 GNDA 0.053331f
C1126 two_stage_opamp_dummy_magic_23_0.VD2.t10 GNDA 0.053331f
C1127 two_stage_opamp_dummy_magic_23_0.VD2.n34 GNDA 0.116042f
C1128 two_stage_opamp_dummy_magic_23_0.VD2.n35 GNDA 0.447102f
C1129 two_stage_opamp_dummy_magic_23_0.VD2.n36 GNDA 0.099935f
C1130 two_stage_opamp_dummy_magic_23_0.VD2.n37 GNDA 0.06757f
C1131 bgr_11_0.cap_res1.t14 GNDA 0.331712f
C1132 bgr_11_0.cap_res1.t19 GNDA 0.349187f
C1133 bgr_11_0.cap_res1.t17 GNDA 0.350452f
C1134 bgr_11_0.cap_res1.t7 GNDA 0.331712f
C1135 bgr_11_0.cap_res1.t16 GNDA 0.349187f
C1136 bgr_11_0.cap_res1.t11 GNDA 0.350452f
C1137 bgr_11_0.cap_res1.t1 GNDA 0.331712f
C1138 bgr_11_0.cap_res1.t10 GNDA 0.349187f
C1139 bgr_11_0.cap_res1.t3 GNDA 0.350452f
C1140 bgr_11_0.cap_res1.t5 GNDA 0.331712f
C1141 bgr_11_0.cap_res1.t15 GNDA 0.349187f
C1142 bgr_11_0.cap_res1.t9 GNDA 0.350452f
C1143 bgr_11_0.cap_res1.t20 GNDA 0.331712f
C1144 bgr_11_0.cap_res1.t8 GNDA 0.349187f
C1145 bgr_11_0.cap_res1.t2 GNDA 0.350452f
C1146 bgr_11_0.cap_res1.n0 GNDA 0.23406f
C1147 bgr_11_0.cap_res1.t4 GNDA 0.186395f
C1148 bgr_11_0.cap_res1.n1 GNDA 0.253961f
C1149 bgr_11_0.cap_res1.t12 GNDA 0.186395f
C1150 bgr_11_0.cap_res1.n2 GNDA 0.253961f
C1151 bgr_11_0.cap_res1.t6 GNDA 0.186395f
C1152 bgr_11_0.cap_res1.n3 GNDA 0.253961f
C1153 bgr_11_0.cap_res1.t13 GNDA 0.186395f
C1154 bgr_11_0.cap_res1.n4 GNDA 0.253961f
C1155 bgr_11_0.cap_res1.t18 GNDA 0.363549f
C1156 bgr_11_0.cap_res1.t0 GNDA 0.08421f
C1157 bgr_11_0.1st_Vout_1.n0 GNDA 0.902643f
C1158 bgr_11_0.1st_Vout_1.n1 GNDA 1.74831f
C1159 bgr_11_0.1st_Vout_1.n2 GNDA 0.127561f
C1160 bgr_11_0.1st_Vout_1.n3 GNDA 1.79885f
C1161 bgr_11_0.1st_Vout_1.t11 GNDA 0.358464f
C1162 bgr_11_0.1st_Vout_1.t30 GNDA 0.35246f
C1163 bgr_11_0.1st_Vout_1.t26 GNDA 0.358464f
C1164 bgr_11_0.1st_Vout_1.t34 GNDA 0.35246f
C1165 bgr_11_0.1st_Vout_1.t29 GNDA 0.358464f
C1166 bgr_11_0.1st_Vout_1.t22 GNDA 0.35246f
C1167 bgr_11_0.1st_Vout_1.t19 GNDA 0.358464f
C1168 bgr_11_0.1st_Vout_1.t25 GNDA 0.35246f
C1169 bgr_11_0.1st_Vout_1.t36 GNDA 0.358464f
C1170 bgr_11_0.1st_Vout_1.t28 GNDA 0.35246f
C1171 bgr_11_0.1st_Vout_1.t24 GNDA 0.358464f
C1172 bgr_11_0.1st_Vout_1.t33 GNDA 0.35246f
C1173 bgr_11_0.1st_Vout_1.t27 GNDA 0.358464f
C1174 bgr_11_0.1st_Vout_1.t21 GNDA 0.35246f
C1175 bgr_11_0.1st_Vout_1.t16 GNDA 0.358464f
C1176 bgr_11_0.1st_Vout_1.t23 GNDA 0.35246f
C1177 bgr_11_0.1st_Vout_1.t20 GNDA 0.358464f
C1178 bgr_11_0.1st_Vout_1.t13 GNDA 0.35246f
C1179 bgr_11_0.1st_Vout_1.t15 GNDA 0.35246f
C1180 bgr_11_0.1st_Vout_1.t12 GNDA 0.35246f
C1181 bgr_11_0.1st_Vout_1.t17 GNDA 0.023025f
C1182 bgr_11_0.1st_Vout_1.n4 GNDA 0.022212f
C1183 bgr_11_0.1st_Vout_1.t35 GNDA 0.013423f
C1184 bgr_11_0.1st_Vout_1.t14 GNDA 0.013423f
C1185 bgr_11_0.1st_Vout_1.n5 GNDA 0.029862f
C1186 bgr_11_0.1st_Vout_1.t4 GNDA 0.018559f
C1187 bgr_11_0.1st_Vout_1.n6 GNDA 0.012728f
C1188 bgr_11_0.1st_Vout_1.n7 GNDA 0.192525f
C1189 bgr_11_0.1st_Vout_1.n8 GNDA 0.011517f
C1190 bgr_11_0.1st_Vout_1.n9 GNDA 0.021291f
C1191 bgr_11_0.1st_Vout_1.t31 GNDA 0.013423f
C1192 bgr_11_0.1st_Vout_1.t18 GNDA 0.013423f
C1193 bgr_11_0.1st_Vout_1.n10 GNDA 0.029862f
C1194 bgr_11_0.1st_Vout_1.n11 GNDA 0.022212f
C1195 bgr_11_0.1st_Vout_1.t32 GNDA 0.021069f
C1196 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t57 GNDA 0.343734f
C1197 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t66 GNDA 0.344881f
C1198 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t26 GNDA 0.185242f
C1199 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n0 GNDA 0.197802f
C1200 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t96 GNDA 0.343734f
C1201 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t101 GNDA 0.344881f
C1202 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t63 GNDA 0.185242f
C1203 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n1 GNDA 0.216311f
C1204 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t75 GNDA 0.343734f
C1205 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t81 GNDA 0.344881f
C1206 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t42 GNDA 0.185242f
C1207 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n2 GNDA 0.216311f
C1208 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t113 GNDA 0.343734f
C1209 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t120 GNDA 0.344881f
C1210 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t79 GNDA 0.185242f
C1211 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n3 GNDA 0.216311f
C1212 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t9 GNDA 0.343734f
C1213 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t43 GNDA 0.344881f
C1214 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t1 GNDA 0.36339f
C1215 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t17 GNDA 0.36339f
C1216 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t115 GNDA 0.185242f
C1217 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n4 GNDA 0.216311f
C1218 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t47 GNDA 0.343734f
C1219 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t76 GNDA 0.344881f
C1220 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t38 GNDA 0.36339f
C1221 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t51 GNDA 0.36339f
C1222 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t16 GNDA 0.185242f
C1223 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n5 GNDA 0.216311f
C1224 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t52 GNDA 0.344881f
C1225 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t89 GNDA 0.346131f
C1226 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t91 GNDA 0.344881f
C1227 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t129 GNDA 0.347585f
C1228 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t121 GNDA 0.378048f
C1229 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t109 GNDA 0.344881f
C1230 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t87 GNDA 0.346131f
C1231 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t95 GNDA 0.344881f
C1232 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t133 GNDA 0.346131f
C1233 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t18 GNDA 0.344881f
C1234 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t69 GNDA 0.346131f
C1235 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t131 GNDA 0.344881f
C1236 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t132 GNDA 0.346131f
C1237 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t53 GNDA 0.344881f
C1238 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t106 GNDA 0.346131f
C1239 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t28 GNDA 0.344881f
C1240 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t29 GNDA 0.346131f
C1241 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t22 GNDA 0.344881f
C1242 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t74 GNDA 0.346131f
C1243 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t134 GNDA 0.344881f
C1244 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t136 GNDA 0.346131f
C1245 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t60 GNDA 0.344881f
C1246 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t111 GNDA 0.346131f
C1247 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t34 GNDA 0.344881f
C1248 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t36 GNDA 0.346131f
C1249 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t100 GNDA 0.344881f
C1250 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t13 GNDA 0.346131f
C1251 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t72 GNDA 0.344881f
C1252 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t73 GNDA 0.346131f
C1253 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t68 GNDA 0.344881f
C1254 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t119 GNDA 0.346131f
C1255 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t39 GNDA 0.344881f
C1256 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t40 GNDA 0.346131f
C1257 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t105 GNDA 0.344881f
C1258 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t19 GNDA 0.346131f
C1259 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t77 GNDA 0.344881f
C1260 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t78 GNDA 0.346131f
C1261 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t6 GNDA 0.344881f
C1262 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t55 GNDA 0.346131f
C1263 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t116 GNDA 0.344881f
C1264 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t117 GNDA 0.346131f
C1265 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t110 GNDA 0.344881f
C1266 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t24 GNDA 0.346131f
C1267 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t83 GNDA 0.344881f
C1268 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t84 GNDA 0.346131f
C1269 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t12 GNDA 0.344881f
C1270 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t64 GNDA 0.346131f
C1271 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t125 GNDA 0.344881f
C1272 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t127 GNDA 0.346131f
C1273 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t48 GNDA 0.344881f
C1274 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t102 GNDA 0.346131f
C1275 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t21 GNDA 0.344881f
C1276 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t23 GNDA 0.346131f
C1277 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t90 GNDA 0.344881f
C1278 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t2 GNDA 0.346131f
C1279 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t59 GNDA 0.344881f
C1280 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t61 GNDA 0.346131f
C1281 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t54 GNDA 0.344881f
C1282 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t108 GNDA 0.346131f
C1283 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t27 GNDA 0.344881f
C1284 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t30 GNDA 0.346131f
C1285 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t118 GNDA 0.344881f
C1286 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t62 GNDA 0.36179f
C1287 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t14 GNDA 0.344881f
C1288 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t11 GNDA 0.185242f
C1289 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n6 GNDA 0.198255f
C1290 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t65 GNDA 0.344881f
C1291 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t50 GNDA 0.185242f
C1292 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n7 GNDA 0.196656f
C1293 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t98 GNDA 0.344881f
C1294 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t4 GNDA 0.185242f
C1295 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n8 GNDA 0.196656f
C1296 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t137 GNDA 0.344881f
C1297 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t92 GNDA 0.185242f
C1298 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n9 GNDA 0.196656f
C1299 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t32 GNDA 0.344881f
C1300 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t44 GNDA 0.185242f
C1301 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n10 GNDA 0.196656f
C1302 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t80 GNDA 0.344881f
C1303 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t85 GNDA 0.185242f
C1304 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n11 GNDA 0.196656f
C1305 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t114 GNDA 0.344881f
C1306 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t37 GNDA 0.185242f
C1307 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n12 GNDA 0.196656f
C1308 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t8 GNDA 0.344881f
C1309 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t126 GNDA 0.185242f
C1310 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n13 GNDA 0.196656f
C1311 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t58 GNDA 0.344881f
C1312 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t25 GNDA 0.185242f
C1313 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n14 GNDA 0.196656f
C1314 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t99 GNDA 0.344881f
C1315 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t10 GNDA 0.346131f
C1316 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t122 GNDA 0.344881f
C1317 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t123 GNDA 0.346131f
C1318 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t94 GNDA 0.166734f
C1319 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n15 GNDA 0.215061f
C1320 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t112 GNDA 0.184096f
C1321 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n16 GNDA 0.23357f
C1322 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t5 GNDA 0.184096f
C1323 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n17 GNDA 0.250829f
C1324 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t41 GNDA 0.184096f
C1325 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n18 GNDA 0.250829f
C1326 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t138 GNDA 0.184096f
C1327 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n19 GNDA 0.250829f
C1328 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t97 GNDA 0.184096f
C1329 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n20 GNDA 0.250829f
C1330 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t56 GNDA 0.184096f
C1331 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n21 GNDA 0.250829f
C1332 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t93 GNDA 0.184096f
C1333 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n22 GNDA 0.250829f
C1334 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t49 GNDA 0.184096f
C1335 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n23 GNDA 0.250829f
C1336 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t15 GNDA 0.184096f
C1337 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n24 GNDA 0.250829f
C1338 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t46 GNDA 0.184096f
C1339 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n25 GNDA 0.250829f
C1340 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t7 GNDA 0.184096f
C1341 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n26 GNDA 0.250829f
C1342 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t107 GNDA 0.184096f
C1343 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n27 GNDA 0.250829f
C1344 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t3 GNDA 0.184096f
C1345 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n28 GNDA 0.250829f
C1346 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t103 GNDA 0.184096f
C1347 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n29 GNDA 0.250829f
C1348 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t128 GNDA 0.184096f
C1349 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n30 GNDA 0.250829f
C1350 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t86 GNDA 0.184096f
C1351 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n31 GNDA 0.23357f
C1352 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t82 GNDA 0.343734f
C1353 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t45 GNDA 0.166734f
C1354 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n32 GNDA 0.216311f
C1355 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t104 GNDA 0.343734f
C1356 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t70 GNDA 0.166734f
C1357 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n33 GNDA 0.216311f
C1358 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t67 GNDA 0.343734f
C1359 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t20 GNDA 0.344881f
C1360 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t124 GNDA 0.36339f
C1361 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t71 GNDA 0.36339f
C1362 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t33 GNDA 0.185242f
C1363 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n34 GNDA 0.216311f
C1364 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t31 GNDA 0.343734f
C1365 two_stage_opamp_dummy_magic_23_0.cap_res_Y.n35 GNDA 0.216311f
C1366 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t135 GNDA 0.185242f
C1367 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t35 GNDA 0.36339f
C1368 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t88 GNDA 0.36339f
C1369 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t130 GNDA 0.434792f
C1370 two_stage_opamp_dummy_magic_23_0.cap_res_Y.t0 GNDA 0.291879f
C1371 two_stage_opamp_dummy_magic_23_0.V_err_gate.n0 GNDA 0.273851f
C1372 two_stage_opamp_dummy_magic_23_0.V_err_gate.n1 GNDA 0.273851f
C1373 two_stage_opamp_dummy_magic_23_0.V_err_gate.n2 GNDA 0.249906f
C1374 two_stage_opamp_dummy_magic_23_0.V_err_gate.n3 GNDA 0.347481f
C1375 two_stage_opamp_dummy_magic_23_0.V_err_gate.n4 GNDA 0.179504f
C1376 two_stage_opamp_dummy_magic_23_0.V_err_gate.n5 GNDA 0.211361f
C1377 two_stage_opamp_dummy_magic_23_0.V_err_gate.t4 GNDA 0.033289f
C1378 two_stage_opamp_dummy_magic_23_0.V_err_gate.t3 GNDA 0.033289f
C1379 two_stage_opamp_dummy_magic_23_0.V_err_gate.n6 GNDA 0.509125f
C1380 two_stage_opamp_dummy_magic_23_0.V_err_gate.t19 GNDA 0.013731f
C1381 two_stage_opamp_dummy_magic_23_0.V_err_gate.t15 GNDA 0.013731f
C1382 two_stage_opamp_dummy_magic_23_0.V_err_gate.t25 GNDA 0.013731f
C1383 two_stage_opamp_dummy_magic_23_0.V_err_gate.t33 GNDA 0.013731f
C1384 two_stage_opamp_dummy_magic_23_0.V_err_gate.t23 GNDA 0.013731f
C1385 two_stage_opamp_dummy_magic_23_0.V_err_gate.t32 GNDA 0.013731f
C1386 two_stage_opamp_dummy_magic_23_0.V_err_gate.t22 GNDA 0.013731f
C1387 two_stage_opamp_dummy_magic_23_0.V_err_gate.t30 GNDA 0.013731f
C1388 two_stage_opamp_dummy_magic_23_0.V_err_gate.t20 GNDA 0.013731f
C1389 two_stage_opamp_dummy_magic_23_0.V_err_gate.t24 GNDA 0.013731f
C1390 two_stage_opamp_dummy_magic_23_0.V_err_gate.t16 GNDA 0.029752f
C1391 two_stage_opamp_dummy_magic_23_0.V_err_gate.n7 GNDA 0.046396f
C1392 two_stage_opamp_dummy_magic_23_0.V_err_gate.n8 GNDA 0.036201f
C1393 two_stage_opamp_dummy_magic_23_0.V_err_gate.n9 GNDA 0.036201f
C1394 two_stage_opamp_dummy_magic_23_0.V_err_gate.n10 GNDA 0.036201f
C1395 two_stage_opamp_dummy_magic_23_0.V_err_gate.n11 GNDA 0.036201f
C1396 two_stage_opamp_dummy_magic_23_0.V_err_gate.n12 GNDA 0.036201f
C1397 two_stage_opamp_dummy_magic_23_0.V_err_gate.n13 GNDA 0.036201f
C1398 two_stage_opamp_dummy_magic_23_0.V_err_gate.n14 GNDA 0.036201f
C1399 two_stage_opamp_dummy_magic_23_0.V_err_gate.n15 GNDA 0.036201f
C1400 two_stage_opamp_dummy_magic_23_0.V_err_gate.n16 GNDA 0.029692f
C1401 two_stage_opamp_dummy_magic_23_0.V_err_gate.t29 GNDA 0.013731f
C1402 two_stage_opamp_dummy_magic_23_0.V_err_gate.t26 GNDA 0.013731f
C1403 two_stage_opamp_dummy_magic_23_0.V_err_gate.t17 GNDA 0.013731f
C1404 two_stage_opamp_dummy_magic_23_0.V_err_gate.t27 GNDA 0.013731f
C1405 two_stage_opamp_dummy_magic_23_0.V_err_gate.t18 GNDA 0.013731f
C1406 two_stage_opamp_dummy_magic_23_0.V_err_gate.t28 GNDA 0.013731f
C1407 two_stage_opamp_dummy_magic_23_0.V_err_gate.t21 GNDA 0.013731f
C1408 two_stage_opamp_dummy_magic_23_0.V_err_gate.t31 GNDA 0.013731f
C1409 two_stage_opamp_dummy_magic_23_0.V_err_gate.t14 GNDA 0.034329f
C1410 two_stage_opamp_dummy_magic_23_0.V_err_gate.n17 GNDA 0.071779f
C1411 two_stage_opamp_dummy_magic_23_0.V_err_gate.n18 GNDA 0.036201f
C1412 two_stage_opamp_dummy_magic_23_0.V_err_gate.n19 GNDA 0.036201f
C1413 two_stage_opamp_dummy_magic_23_0.V_err_gate.n20 GNDA 0.036201f
C1414 two_stage_opamp_dummy_magic_23_0.V_err_gate.n21 GNDA 0.036201f
C1415 two_stage_opamp_dummy_magic_23_0.V_err_gate.n22 GNDA 0.036201f
C1416 two_stage_opamp_dummy_magic_23_0.V_err_gate.n23 GNDA 0.036201f
C1417 two_stage_opamp_dummy_magic_23_0.V_err_gate.n24 GNDA 0.029692f
C1418 two_stage_opamp_dummy_magic_23_0.V_err_gate.n25 GNDA 0.045627f
C1419 two_stage_opamp_dummy_magic_23_0.V_err_gate.t6 GNDA 0.016644f
C1420 two_stage_opamp_dummy_magic_23_0.V_err_gate.t10 GNDA 0.016644f
C1421 two_stage_opamp_dummy_magic_23_0.V_err_gate.n26 GNDA 0.033914f
C1422 two_stage_opamp_dummy_magic_23_0.V_err_gate.t0 GNDA 0.016644f
C1423 two_stage_opamp_dummy_magic_23_0.V_err_gate.t9 GNDA 0.016644f
C1424 two_stage_opamp_dummy_magic_23_0.V_err_gate.n27 GNDA 0.033914f
C1425 two_stage_opamp_dummy_magic_23_0.V_err_gate.n28 GNDA 0.2329f
C1426 two_stage_opamp_dummy_magic_23_0.V_err_gate.t2 GNDA 0.016644f
C1427 two_stage_opamp_dummy_magic_23_0.V_err_gate.t1 GNDA 0.016644f
C1428 two_stage_opamp_dummy_magic_23_0.V_err_gate.n29 GNDA 0.033914f
C1429 two_stage_opamp_dummy_magic_23_0.V_err_gate.n30 GNDA 0.2329f
C1430 two_stage_opamp_dummy_magic_23_0.V_err_gate.t7 GNDA 0.016644f
C1431 two_stage_opamp_dummy_magic_23_0.V_err_gate.t8 GNDA 0.016644f
C1432 two_stage_opamp_dummy_magic_23_0.V_err_gate.n31 GNDA 0.033914f
C1433 two_stage_opamp_dummy_magic_23_0.V_err_gate.n32 GNDA 0.2329f
C1434 two_stage_opamp_dummy_magic_23_0.V_err_gate.t5 GNDA 0.016644f
C1435 two_stage_opamp_dummy_magic_23_0.V_err_gate.t12 GNDA 0.016644f
C1436 two_stage_opamp_dummy_magic_23_0.V_err_gate.n33 GNDA 0.033914f
C1437 two_stage_opamp_dummy_magic_23_0.V_err_gate.n34 GNDA 0.2329f
C1438 two_stage_opamp_dummy_magic_23_0.V_err_gate.t11 GNDA 0.016644f
C1439 two_stage_opamp_dummy_magic_23_0.V_err_gate.t13 GNDA 0.016644f
C1440 two_stage_opamp_dummy_magic_23_0.V_err_gate.n35 GNDA 0.033914f
C1441 two_stage_opamp_dummy_magic_23_0.V_err_gate.n36 GNDA 0.241351f
C1442 bgr_11_0.NFET_GATE_10uA.t3 GNDA 0.01496f
C1443 bgr_11_0.NFET_GATE_10uA.t1 GNDA 0.01496f
C1444 bgr_11_0.NFET_GATE_10uA.n0 GNDA 0.042091f
C1445 bgr_11_0.NFET_GATE_10uA.t5 GNDA 0.014586f
C1446 bgr_11_0.NFET_GATE_10uA.t10 GNDA 0.014586f
C1447 bgr_11_0.NFET_GATE_10uA.t18 GNDA 0.014586f
C1448 bgr_11_0.NFET_GATE_10uA.t7 GNDA 0.014586f
C1449 bgr_11_0.NFET_GATE_10uA.t15 GNDA 0.014586f
C1450 bgr_11_0.NFET_GATE_10uA.t14 GNDA 0.014586f
C1451 bgr_11_0.NFET_GATE_10uA.t21 GNDA 0.021563f
C1452 bgr_11_0.NFET_GATE_10uA.n1 GNDA 0.026685f
C1453 bgr_11_0.NFET_GATE_10uA.n2 GNDA 0.019075f
C1454 bgr_11_0.NFET_GATE_10uA.n3 GNDA 0.016149f
C1455 bgr_11_0.NFET_GATE_10uA.t23 GNDA 0.014586f
C1456 bgr_11_0.NFET_GATE_10uA.t16 GNDA 0.014586f
C1457 bgr_11_0.NFET_GATE_10uA.t8 GNDA 0.014586f
C1458 bgr_11_0.NFET_GATE_10uA.t22 GNDA 0.021563f
C1459 bgr_11_0.NFET_GATE_10uA.n4 GNDA 0.026685f
C1460 bgr_11_0.NFET_GATE_10uA.n5 GNDA 0.019075f
C1461 bgr_11_0.NFET_GATE_10uA.n6 GNDA 0.016149f
C1462 bgr_11_0.NFET_GATE_10uA.t9 GNDA 0.014586f
C1463 bgr_11_0.NFET_GATE_10uA.t17 GNDA 0.021563f
C1464 bgr_11_0.NFET_GATE_10uA.n7 GNDA 0.02376f
C1465 bgr_11_0.NFET_GATE_10uA.n8 GNDA 0.026114f
C1466 bgr_11_0.NFET_GATE_10uA.t11 GNDA 0.014586f
C1467 bgr_11_0.NFET_GATE_10uA.t13 GNDA 0.021563f
C1468 bgr_11_0.NFET_GATE_10uA.n9 GNDA 0.02376f
C1469 bgr_11_0.NFET_GATE_10uA.t19 GNDA 0.014586f
C1470 bgr_11_0.NFET_GATE_10uA.t6 GNDA 0.014586f
C1471 bgr_11_0.NFET_GATE_10uA.t12 GNDA 0.014586f
C1472 bgr_11_0.NFET_GATE_10uA.t20 GNDA 0.021563f
C1473 bgr_11_0.NFET_GATE_10uA.n10 GNDA 0.026685f
C1474 bgr_11_0.NFET_GATE_10uA.n11 GNDA 0.019075f
C1475 bgr_11_0.NFET_GATE_10uA.n12 GNDA 0.016149f
C1476 bgr_11_0.NFET_GATE_10uA.n13 GNDA 0.026114f
C1477 bgr_11_0.NFET_GATE_10uA.n14 GNDA 0.605807f
C1478 bgr_11_0.NFET_GATE_10uA.n15 GNDA 0.022264f
C1479 bgr_11_0.NFET_GATE_10uA.n16 GNDA 0.016149f
C1480 bgr_11_0.NFET_GATE_10uA.n17 GNDA 0.019075f
C1481 bgr_11_0.NFET_GATE_10uA.n18 GNDA 0.026685f
C1482 bgr_11_0.NFET_GATE_10uA.t0 GNDA 0.034164f
C1483 bgr_11_0.NFET_GATE_10uA.n19 GNDA 0.327308f
C1484 bgr_11_0.NFET_GATE_10uA.t2 GNDA 0.01496f
C1485 bgr_11_0.NFET_GATE_10uA.t4 GNDA 0.01496f
C1486 bgr_11_0.NFET_GATE_10uA.n20 GNDA 0.088541f
C1487 two_stage_opamp_dummy_magic_23_0.VD3.t16 GNDA 0.060837f
C1488 two_stage_opamp_dummy_magic_23_0.VD3.t26 GNDA 0.060837f
C1489 two_stage_opamp_dummy_magic_23_0.VD3.t32 GNDA 0.060837f
C1490 two_stage_opamp_dummy_magic_23_0.VD3.n0 GNDA 0.154422f
C1491 two_stage_opamp_dummy_magic_23_0.VD3.n1 GNDA 0.43135f
C1492 two_stage_opamp_dummy_magic_23_0.VD3.t3 GNDA 0.106675f
C1493 two_stage_opamp_dummy_magic_23_0.VD3.t2 GNDA 0.216405f
C1494 two_stage_opamp_dummy_magic_23_0.VD3.n2 GNDA 0.065988f
C1495 two_stage_opamp_dummy_magic_23_0.VD3.n3 GNDA 0.065988f
C1496 two_stage_opamp_dummy_magic_23_0.VD3.t13 GNDA 0.060837f
C1497 two_stage_opamp_dummy_magic_23_0.VD3.t37 GNDA 0.060837f
C1498 two_stage_opamp_dummy_magic_23_0.VD3.n4 GNDA 0.124448f
C1499 two_stage_opamp_dummy_magic_23_0.VD3.n5 GNDA 0.402926f
C1500 two_stage_opamp_dummy_magic_23_0.VD3.n6 GNDA 0.112569f
C1501 two_stage_opamp_dummy_magic_23_0.VD3.t8 GNDA 0.060837f
C1502 two_stage_opamp_dummy_magic_23_0.VD3.t36 GNDA 0.060837f
C1503 two_stage_opamp_dummy_magic_23_0.VD3.n7 GNDA 0.124448f
C1504 two_stage_opamp_dummy_magic_23_0.VD3.n8 GNDA 0.391923f
C1505 two_stage_opamp_dummy_magic_23_0.VD3.n9 GNDA 0.112569f
C1506 two_stage_opamp_dummy_magic_23_0.VD3.t12 GNDA 0.060837f
C1507 two_stage_opamp_dummy_magic_23_0.VD3.t9 GNDA 0.060837f
C1508 two_stage_opamp_dummy_magic_23_0.VD3.n10 GNDA 0.124448f
C1509 two_stage_opamp_dummy_magic_23_0.VD3.n11 GNDA 0.391923f
C1510 two_stage_opamp_dummy_magic_23_0.VD3.n12 GNDA 0.065988f
C1511 two_stage_opamp_dummy_magic_23_0.VD3.n13 GNDA 0.065988f
C1512 two_stage_opamp_dummy_magic_23_0.VD3.t6 GNDA 0.060837f
C1513 two_stage_opamp_dummy_magic_23_0.VD3.t35 GNDA 0.060837f
C1514 two_stage_opamp_dummy_magic_23_0.VD3.n14 GNDA 0.124448f
C1515 two_stage_opamp_dummy_magic_23_0.VD3.n15 GNDA 0.391923f
C1516 two_stage_opamp_dummy_magic_23_0.VD3.n16 GNDA 0.065988f
C1517 two_stage_opamp_dummy_magic_23_0.VD3.t10 GNDA 0.060837f
C1518 two_stage_opamp_dummy_magic_23_0.VD3.t11 GNDA 0.060837f
C1519 two_stage_opamp_dummy_magic_23_0.VD3.n17 GNDA 0.124448f
C1520 two_stage_opamp_dummy_magic_23_0.VD3.n18 GNDA 0.391923f
C1521 two_stage_opamp_dummy_magic_23_0.VD3.n19 GNDA 0.112569f
C1522 two_stage_opamp_dummy_magic_23_0.VD3.t7 GNDA 0.060837f
C1523 two_stage_opamp_dummy_magic_23_0.VD3.t14 GNDA 0.060837f
C1524 two_stage_opamp_dummy_magic_23_0.VD3.n20 GNDA 0.124448f
C1525 two_stage_opamp_dummy_magic_23_0.VD3.n21 GNDA 0.397425f
C1526 two_stage_opamp_dummy_magic_23_0.VD3.n22 GNDA 0.257485f
C1527 two_stage_opamp_dummy_magic_23_0.VD3.t24 GNDA 0.060837f
C1528 two_stage_opamp_dummy_magic_23_0.VD3.t30 GNDA 0.060837f
C1529 two_stage_opamp_dummy_magic_23_0.VD3.n23 GNDA 0.154422f
C1530 two_stage_opamp_dummy_magic_23_0.VD3.n24 GNDA 0.43135f
C1531 two_stage_opamp_dummy_magic_23_0.VD3.n25 GNDA 0.2193f
C1532 two_stage_opamp_dummy_magic_23_0.VD3.t0 GNDA 0.106675f
C1533 two_stage_opamp_dummy_magic_23_0.VD3.n26 GNDA 0.311214f
C1534 two_stage_opamp_dummy_magic_23_0.VD3.n27 GNDA 0.627773f
C1535 two_stage_opamp_dummy_magic_23_0.VD3.t1 GNDA 0.518568f
C1536 two_stage_opamp_dummy_magic_23_0.VD3.t23 GNDA 0.406738f
C1537 two_stage_opamp_dummy_magic_23_0.VD3.t29 GNDA 0.406738f
C1538 two_stage_opamp_dummy_magic_23_0.VD3.t25 GNDA 0.406738f
C1539 two_stage_opamp_dummy_magic_23_0.VD3.t31 GNDA 0.402972f
C1540 two_stage_opamp_dummy_magic_23_0.VD3.t33 GNDA 0.399206f
C1541 two_stage_opamp_dummy_magic_23_0.VD3.t15 GNDA 0.406738f
C1542 two_stage_opamp_dummy_magic_23_0.VD3.t19 GNDA 0.406738f
C1543 two_stage_opamp_dummy_magic_23_0.VD3.t17 GNDA 0.406738f
C1544 two_stage_opamp_dummy_magic_23_0.VD3.t21 GNDA 0.406738f
C1545 two_stage_opamp_dummy_magic_23_0.VD3.t27 GNDA 0.406738f
C1546 two_stage_opamp_dummy_magic_23_0.VD3.t4 GNDA 0.518568f
C1547 two_stage_opamp_dummy_magic_23_0.VD3.t5 GNDA 0.216405f
C1548 two_stage_opamp_dummy_magic_23_0.VD3.n28 GNDA 0.627773f
C1549 two_stage_opamp_dummy_magic_23_0.VD3.n29 GNDA 0.316969f
C1550 two_stage_opamp_dummy_magic_23_0.VD3.t22 GNDA 0.060837f
C1551 two_stage_opamp_dummy_magic_23_0.VD3.t28 GNDA 0.060837f
C1552 two_stage_opamp_dummy_magic_23_0.VD3.n30 GNDA 0.154422f
C1553 two_stage_opamp_dummy_magic_23_0.VD3.n31 GNDA 0.481799f
C1554 two_stage_opamp_dummy_magic_23_0.VD3.t20 GNDA 0.060837f
C1555 two_stage_opamp_dummy_magic_23_0.VD3.t18 GNDA 0.060837f
C1556 two_stage_opamp_dummy_magic_23_0.VD3.n32 GNDA 0.154422f
C1557 two_stage_opamp_dummy_magic_23_0.VD3.n33 GNDA 0.43135f
C1558 two_stage_opamp_dummy_magic_23_0.VD3.n34 GNDA 0.43135f
C1559 two_stage_opamp_dummy_magic_23_0.VD3.n35 GNDA 0.154422f
C1560 two_stage_opamp_dummy_magic_23_0.VD3.t34 GNDA 0.060837f
C1561 two_stage_opamp_dummy_magic_23_0.Vb2.t10 GNDA 0.047503f
C1562 two_stage_opamp_dummy_magic_23_0.Vb2.t1 GNDA 0.013572f
C1563 two_stage_opamp_dummy_magic_23_0.Vb2.t8 GNDA 0.013572f
C1564 two_stage_opamp_dummy_magic_23_0.Vb2.n0 GNDA 0.046239f
C1565 two_stage_opamp_dummy_magic_23_0.Vb2.t3 GNDA 0.013572f
C1566 two_stage_opamp_dummy_magic_23_0.Vb2.t0 GNDA 0.013572f
C1567 two_stage_opamp_dummy_magic_23_0.Vb2.n1 GNDA 0.044879f
C1568 two_stage_opamp_dummy_magic_23_0.Vb2.n2 GNDA 0.466707f
C1569 two_stage_opamp_dummy_magic_23_0.Vb2.t4 GNDA 0.013572f
C1570 two_stage_opamp_dummy_magic_23_0.Vb2.t6 GNDA 0.013572f
C1571 two_stage_opamp_dummy_magic_23_0.Vb2.n3 GNDA 0.044879f
C1572 two_stage_opamp_dummy_magic_23_0.Vb2.n4 GNDA 0.314789f
C1573 two_stage_opamp_dummy_magic_23_0.Vb2.t7 GNDA 0.013572f
C1574 two_stage_opamp_dummy_magic_23_0.Vb2.t5 GNDA 0.013572f
C1575 two_stage_opamp_dummy_magic_23_0.Vb2.n5 GNDA 0.044879f
C1576 two_stage_opamp_dummy_magic_23_0.Vb2.n6 GNDA 1.3433f
C1577 two_stage_opamp_dummy_magic_23_0.Vb2.t15 GNDA 0.087308f
C1578 two_stage_opamp_dummy_magic_23_0.Vb2.n7 GNDA 1.22205f
C1579 two_stage_opamp_dummy_magic_23_0.Vb2.t28 GNDA 0.067183f
C1580 two_stage_opamp_dummy_magic_23_0.Vb2.t23 GNDA 0.067183f
C1581 two_stage_opamp_dummy_magic_23_0.Vb2.t26 GNDA 0.067183f
C1582 two_stage_opamp_dummy_magic_23_0.Vb2.t21 GNDA 0.067183f
C1583 two_stage_opamp_dummy_magic_23_0.Vb2.t16 GNDA 0.077529f
C1584 two_stage_opamp_dummy_magic_23_0.Vb2.n8 GNDA 0.062945f
C1585 two_stage_opamp_dummy_magic_23_0.Vb2.n9 GNDA 0.038681f
C1586 two_stage_opamp_dummy_magic_23_0.Vb2.n10 GNDA 0.038681f
C1587 two_stage_opamp_dummy_magic_23_0.Vb2.n11 GNDA 0.033916f
C1588 two_stage_opamp_dummy_magic_23_0.Vb2.t11 GNDA 0.067183f
C1589 two_stage_opamp_dummy_magic_23_0.Vb2.t13 GNDA 0.067183f
C1590 two_stage_opamp_dummy_magic_23_0.Vb2.t17 GNDA 0.067183f
C1591 two_stage_opamp_dummy_magic_23_0.Vb2.t14 GNDA 0.067183f
C1592 two_stage_opamp_dummy_magic_23_0.Vb2.t19 GNDA 0.077529f
C1593 two_stage_opamp_dummy_magic_23_0.Vb2.n12 GNDA 0.062945f
C1594 two_stage_opamp_dummy_magic_23_0.Vb2.n13 GNDA 0.038681f
C1595 two_stage_opamp_dummy_magic_23_0.Vb2.n14 GNDA 0.038681f
C1596 two_stage_opamp_dummy_magic_23_0.Vb2.n15 GNDA 0.033916f
C1597 two_stage_opamp_dummy_magic_23_0.Vb2.n16 GNDA 0.025137f
C1598 two_stage_opamp_dummy_magic_23_0.Vb2.t32 GNDA 0.067183f
C1599 two_stage_opamp_dummy_magic_23_0.Vb2.t29 GNDA 0.067183f
C1600 two_stage_opamp_dummy_magic_23_0.Vb2.t25 GNDA 0.067183f
C1601 two_stage_opamp_dummy_magic_23_0.Vb2.t20 GNDA 0.067183f
C1602 two_stage_opamp_dummy_magic_23_0.Vb2.t24 GNDA 0.077529f
C1603 two_stage_opamp_dummy_magic_23_0.Vb2.n17 GNDA 0.062945f
C1604 two_stage_opamp_dummy_magic_23_0.Vb2.n18 GNDA 0.038681f
C1605 two_stage_opamp_dummy_magic_23_0.Vb2.n19 GNDA 0.038681f
C1606 two_stage_opamp_dummy_magic_23_0.Vb2.n20 GNDA 0.033916f
C1607 two_stage_opamp_dummy_magic_23_0.Vb2.t12 GNDA 0.067183f
C1608 two_stage_opamp_dummy_magic_23_0.Vb2.t18 GNDA 0.067183f
C1609 two_stage_opamp_dummy_magic_23_0.Vb2.t22 GNDA 0.067183f
C1610 two_stage_opamp_dummy_magic_23_0.Vb2.t27 GNDA 0.067183f
C1611 two_stage_opamp_dummy_magic_23_0.Vb2.t30 GNDA 0.077529f
C1612 two_stage_opamp_dummy_magic_23_0.Vb2.n21 GNDA 0.062945f
C1613 two_stage_opamp_dummy_magic_23_0.Vb2.n22 GNDA 0.038681f
C1614 two_stage_opamp_dummy_magic_23_0.Vb2.n23 GNDA 0.038681f
C1615 two_stage_opamp_dummy_magic_23_0.Vb2.n24 GNDA 0.033916f
C1616 two_stage_opamp_dummy_magic_23_0.Vb2.n25 GNDA 0.024767f
C1617 two_stage_opamp_dummy_magic_23_0.Vb2.n26 GNDA 0.539878f
C1618 two_stage_opamp_dummy_magic_23_0.Vb2.n27 GNDA 0.251782f
C1619 two_stage_opamp_dummy_magic_23_0.Vb2.t31 GNDA 0.053254f
C1620 two_stage_opamp_dummy_magic_23_0.Vb2.n28 GNDA 0.204443f
C1621 two_stage_opamp_dummy_magic_23_0.Vb2.t9 GNDA 0.088676f
C1622 two_stage_opamp_dummy_magic_23_0.Vb2.n29 GNDA 0.410624f
C1623 two_stage_opamp_dummy_magic_23_0.Vb2.n30 GNDA 0.100877f
C1624 two_stage_opamp_dummy_magic_23_0.Vb2.t2 GNDA 0.047503f
C1625 two_stage_opamp_dummy_magic_23_0.VD1.t16 GNDA 0.053331f
C1626 two_stage_opamp_dummy_magic_23_0.VD1.n0 GNDA 0.203944f
C1627 two_stage_opamp_dummy_magic_23_0.VD1.n1 GNDA 0.192793f
C1628 two_stage_opamp_dummy_magic_23_0.VD1.t18 GNDA 0.053331f
C1629 two_stage_opamp_dummy_magic_23_0.VD1.t13 GNDA 0.053331f
C1630 two_stage_opamp_dummy_magic_23_0.VD1.n2 GNDA 0.116042f
C1631 two_stage_opamp_dummy_magic_23_0.VD1.n3 GNDA 0.461069f
C1632 two_stage_opamp_dummy_magic_23_0.VD1.t17 GNDA 0.053331f
C1633 two_stage_opamp_dummy_magic_23_0.VD1.t21 GNDA 0.053331f
C1634 two_stage_opamp_dummy_magic_23_0.VD1.n4 GNDA 0.116042f
C1635 two_stage_opamp_dummy_magic_23_0.VD1.n5 GNDA 0.442486f
C1636 two_stage_opamp_dummy_magic_23_0.VD1.n6 GNDA 0.203944f
C1637 two_stage_opamp_dummy_magic_23_0.VD1.n7 GNDA 0.119128f
C1638 two_stage_opamp_dummy_magic_23_0.VD1.t15 GNDA 0.053331f
C1639 two_stage_opamp_dummy_magic_23_0.VD1.t12 GNDA 0.053331f
C1640 two_stage_opamp_dummy_magic_23_0.VD1.n8 GNDA 0.116042f
C1641 two_stage_opamp_dummy_magic_23_0.VD1.n9 GNDA 0.361396f
C1642 two_stage_opamp_dummy_magic_23_0.VD1.n10 GNDA 0.099935f
C1643 two_stage_opamp_dummy_magic_23_0.VD1.n11 GNDA 0.205342f
C1644 two_stage_opamp_dummy_magic_23_0.VD1.t10 GNDA 0.053331f
C1645 two_stage_opamp_dummy_magic_23_0.VD1.t6 GNDA 0.053331f
C1646 two_stage_opamp_dummy_magic_23_0.VD1.n12 GNDA 0.116042f
C1647 two_stage_opamp_dummy_magic_23_0.VD1.n13 GNDA 0.465721f
C1648 two_stage_opamp_dummy_magic_23_0.VD1.n14 GNDA 0.205342f
C1649 two_stage_opamp_dummy_magic_23_0.VD1.t2 GNDA 0.053331f
C1650 two_stage_opamp_dummy_magic_23_0.VD1.t8 GNDA 0.053331f
C1651 two_stage_opamp_dummy_magic_23_0.VD1.n15 GNDA 0.116042f
C1652 two_stage_opamp_dummy_magic_23_0.VD1.n16 GNDA 0.447102f
C1653 two_stage_opamp_dummy_magic_23_0.VD1.n17 GNDA 0.192793f
C1654 two_stage_opamp_dummy_magic_23_0.VD1.t7 GNDA 0.053331f
C1655 two_stage_opamp_dummy_magic_23_0.VD1.t1 GNDA 0.053331f
C1656 two_stage_opamp_dummy_magic_23_0.VD1.n18 GNDA 0.116042f
C1657 two_stage_opamp_dummy_magic_23_0.VD1.n19 GNDA 0.447102f
C1658 two_stage_opamp_dummy_magic_23_0.VD1.n20 GNDA 0.113419f
C1659 two_stage_opamp_dummy_magic_23_0.VD1.t4 GNDA 0.053331f
C1660 two_stage_opamp_dummy_magic_23_0.VD1.t9 GNDA 0.053331f
C1661 two_stage_opamp_dummy_magic_23_0.VD1.n21 GNDA 0.116042f
C1662 two_stage_opamp_dummy_magic_23_0.VD1.n22 GNDA 0.465721f
C1663 two_stage_opamp_dummy_magic_23_0.VD1.t5 GNDA 0.053331f
C1664 two_stage_opamp_dummy_magic_23_0.VD1.t11 GNDA 0.053331f
C1665 two_stage_opamp_dummy_magic_23_0.VD1.n23 GNDA 0.116042f
C1666 two_stage_opamp_dummy_magic_23_0.VD1.n24 GNDA 0.447102f
C1667 two_stage_opamp_dummy_magic_23_0.VD1.n25 GNDA 0.192793f
C1668 two_stage_opamp_dummy_magic_23_0.VD1.n26 GNDA 0.113419f
C1669 two_stage_opamp_dummy_magic_23_0.VD1.t3 GNDA 0.053331f
C1670 two_stage_opamp_dummy_magic_23_0.VD1.t0 GNDA 0.053331f
C1671 two_stage_opamp_dummy_magic_23_0.VD1.n27 GNDA 0.116042f
C1672 two_stage_opamp_dummy_magic_23_0.VD1.n28 GNDA 0.447102f
C1673 two_stage_opamp_dummy_magic_23_0.VD1.n29 GNDA 0.099935f
C1674 two_stage_opamp_dummy_magic_23_0.VD1.n30 GNDA 0.08441f
C1675 two_stage_opamp_dummy_magic_23_0.VD1.n31 GNDA 0.235249f
C1676 two_stage_opamp_dummy_magic_23_0.VD1.n32 GNDA 0.106662f
C1677 two_stage_opamp_dummy_magic_23_0.VD1.t14 GNDA 0.053331f
C1678 two_stage_opamp_dummy_magic_23_0.VD1.t19 GNDA 0.053331f
C1679 two_stage_opamp_dummy_magic_23_0.VD1.n33 GNDA 0.116042f
C1680 two_stage_opamp_dummy_magic_23_0.VD1.n34 GNDA 0.461069f
C1681 two_stage_opamp_dummy_magic_23_0.VD1.n35 GNDA 0.192793f
C1682 two_stage_opamp_dummy_magic_23_0.VD1.n36 GNDA 0.442486f
C1683 two_stage_opamp_dummy_magic_23_0.VD1.n37 GNDA 0.116042f
C1684 two_stage_opamp_dummy_magic_23_0.VD1.t20 GNDA 0.053331f
C1685 two_stage_opamp_dummy_magic_23_0.X.t16 GNDA 0.038289f
C1686 two_stage_opamp_dummy_magic_23_0.X.t24 GNDA 0.038289f
C1687 two_stage_opamp_dummy_magic_23_0.X.n0 GNDA 0.083312f
C1688 two_stage_opamp_dummy_magic_23_0.X.n1 GNDA 0.259463f
C1689 two_stage_opamp_dummy_magic_23_0.X.n2 GNDA 0.138415f
C1690 two_stage_opamp_dummy_magic_23_0.X.n3 GNDA 0.138415f
C1691 two_stage_opamp_dummy_magic_23_0.X.t14 GNDA 0.038289f
C1692 two_stage_opamp_dummy_magic_23_0.X.t19 GNDA 0.038289f
C1693 two_stage_opamp_dummy_magic_23_0.X.n4 GNDA 0.083312f
C1694 two_stage_opamp_dummy_magic_23_0.X.n5 GNDA 0.331023f
C1695 two_stage_opamp_dummy_magic_23_0.X.t22 GNDA 0.038289f
C1696 two_stage_opamp_dummy_magic_23_0.X.t18 GNDA 0.038289f
C1697 two_stage_opamp_dummy_magic_23_0.X.n6 GNDA 0.083312f
C1698 two_stage_opamp_dummy_magic_23_0.X.n7 GNDA 0.317681f
C1699 two_stage_opamp_dummy_magic_23_0.X.n8 GNDA 0.146421f
C1700 two_stage_opamp_dummy_magic_23_0.X.n9 GNDA 0.085527f
C1701 two_stage_opamp_dummy_magic_23_0.X.t20 GNDA 0.038289f
C1702 two_stage_opamp_dummy_magic_23_0.X.t13 GNDA 0.038289f
C1703 two_stage_opamp_dummy_magic_23_0.X.n10 GNDA 0.083312f
C1704 two_stage_opamp_dummy_magic_23_0.X.n11 GNDA 0.331023f
C1705 two_stage_opamp_dummy_magic_23_0.X.t15 GNDA 0.038289f
C1706 two_stage_opamp_dummy_magic_23_0.X.t23 GNDA 0.038289f
C1707 two_stage_opamp_dummy_magic_23_0.X.n12 GNDA 0.083312f
C1708 two_stage_opamp_dummy_magic_23_0.X.n13 GNDA 0.317681f
C1709 two_stage_opamp_dummy_magic_23_0.X.n14 GNDA 0.146421f
C1710 two_stage_opamp_dummy_magic_23_0.X.n15 GNDA 0.085527f
C1711 two_stage_opamp_dummy_magic_23_0.X.t21 GNDA 0.038289f
C1712 two_stage_opamp_dummy_magic_23_0.X.t17 GNDA 0.038289f
C1713 two_stage_opamp_dummy_magic_23_0.X.n16 GNDA 0.083312f
C1714 two_stage_opamp_dummy_magic_23_0.X.n17 GNDA 0.317681f
C1715 two_stage_opamp_dummy_magic_23_0.X.n18 GNDA 0.081429f
C1716 two_stage_opamp_dummy_magic_23_0.X.n19 GNDA 0.076577f
C1717 two_stage_opamp_dummy_magic_23_0.X.n20 GNDA 0.145807f
C1718 two_stage_opamp_dummy_magic_23_0.X.t7 GNDA 1.22341f
C1719 two_stage_opamp_dummy_magic_23_0.X.t34 GNDA 0.16847f
C1720 two_stage_opamp_dummy_magic_23_0.X.t51 GNDA 0.16847f
C1721 two_stage_opamp_dummy_magic_23_0.X.t37 GNDA 0.16847f
C1722 two_stage_opamp_dummy_magic_23_0.X.t53 GNDA 0.16847f
C1723 two_stage_opamp_dummy_magic_23_0.X.t36 GNDA 0.16847f
C1724 two_stage_opamp_dummy_magic_23_0.X.t52 GNDA 0.16847f
C1725 two_stage_opamp_dummy_magic_23_0.X.t39 GNDA 0.179433f
C1726 two_stage_opamp_dummy_magic_23_0.X.n21 GNDA 0.142193f
C1727 two_stage_opamp_dummy_magic_23_0.X.n22 GNDA 0.080406f
C1728 two_stage_opamp_dummy_magic_23_0.X.n23 GNDA 0.080406f
C1729 two_stage_opamp_dummy_magic_23_0.X.n24 GNDA 0.080406f
C1730 two_stage_opamp_dummy_magic_23_0.X.n25 GNDA 0.080406f
C1731 two_stage_opamp_dummy_magic_23_0.X.n26 GNDA 0.07227f
C1732 two_stage_opamp_dummy_magic_23_0.X.t48 GNDA 0.16847f
C1733 two_stage_opamp_dummy_magic_23_0.X.t31 GNDA 0.16847f
C1734 two_stage_opamp_dummy_magic_23_0.X.t46 GNDA 0.179433f
C1735 two_stage_opamp_dummy_magic_23_0.X.n27 GNDA 0.142193f
C1736 two_stage_opamp_dummy_magic_23_0.X.n28 GNDA 0.07227f
C1737 two_stage_opamp_dummy_magic_23_0.X.n29 GNDA 0.036557f
C1738 two_stage_opamp_dummy_magic_23_0.X.n30 GNDA 1.2754f
C1739 two_stage_opamp_dummy_magic_23_0.X.t3 GNDA 0.08934f
C1740 two_stage_opamp_dummy_magic_23_0.X.t11 GNDA 0.08934f
C1741 two_stage_opamp_dummy_magic_23_0.X.n31 GNDA 0.182755f
C1742 two_stage_opamp_dummy_magic_23_0.X.n32 GNDA 0.497099f
C1743 two_stage_opamp_dummy_magic_23_0.X.n33 GNDA 0.096905f
C1744 two_stage_opamp_dummy_magic_23_0.X.n34 GNDA 0.16531f
C1745 two_stage_opamp_dummy_magic_23_0.X.t8 GNDA 0.08934f
C1746 two_stage_opamp_dummy_magic_23_0.X.t4 GNDA 0.08934f
C1747 two_stage_opamp_dummy_magic_23_0.X.n35 GNDA 0.182755f
C1748 two_stage_opamp_dummy_magic_23_0.X.n36 GNDA 0.591707f
C1749 two_stage_opamp_dummy_magic_23_0.X.t1 GNDA 0.08934f
C1750 two_stage_opamp_dummy_magic_23_0.X.t5 GNDA 0.08934f
C1751 two_stage_opamp_dummy_magic_23_0.X.n37 GNDA 0.182755f
C1752 two_stage_opamp_dummy_magic_23_0.X.n38 GNDA 0.575548f
C1753 two_stage_opamp_dummy_magic_23_0.X.n39 GNDA 0.16531f
C1754 two_stage_opamp_dummy_magic_23_0.X.n40 GNDA 0.096905f
C1755 two_stage_opamp_dummy_magic_23_0.X.t2 GNDA 0.08934f
C1756 two_stage_opamp_dummy_magic_23_0.X.t6 GNDA 0.08934f
C1757 two_stage_opamp_dummy_magic_23_0.X.n41 GNDA 0.182755f
C1758 two_stage_opamp_dummy_magic_23_0.X.n42 GNDA 0.575548f
C1759 two_stage_opamp_dummy_magic_23_0.X.n43 GNDA 0.096905f
C1760 two_stage_opamp_dummy_magic_23_0.X.t12 GNDA 0.08934f
C1761 two_stage_opamp_dummy_magic_23_0.X.t10 GNDA 0.08934f
C1762 two_stage_opamp_dummy_magic_23_0.X.n44 GNDA 0.182755f
C1763 two_stage_opamp_dummy_magic_23_0.X.n45 GNDA 0.575548f
C1764 two_stage_opamp_dummy_magic_23_0.X.n46 GNDA 0.096905f
C1765 two_stage_opamp_dummy_magic_23_0.X.n47 GNDA 0.16531f
C1766 two_stage_opamp_dummy_magic_23_0.X.t0 GNDA 0.08934f
C1767 two_stage_opamp_dummy_magic_23_0.X.t9 GNDA 0.08934f
C1768 two_stage_opamp_dummy_magic_23_0.X.n48 GNDA 0.182755f
C1769 two_stage_opamp_dummy_magic_23_0.X.n49 GNDA 0.575548f
C1770 two_stage_opamp_dummy_magic_23_0.X.n50 GNDA 0.150696f
C1771 two_stage_opamp_dummy_magic_23_0.X.n51 GNDA 0.491162f
C1772 two_stage_opamp_dummy_magic_23_0.X.t44 GNDA 0.053604f
C1773 two_stage_opamp_dummy_magic_23_0.X.t30 GNDA 0.065091f
C1774 two_stage_opamp_dummy_magic_23_0.X.n52 GNDA 0.056954f
C1775 two_stage_opamp_dummy_magic_23_0.X.t27 GNDA 0.053604f
C1776 two_stage_opamp_dummy_magic_23_0.X.t45 GNDA 0.053604f
C1777 two_stage_opamp_dummy_magic_23_0.X.t28 GNDA 0.053604f
C1778 two_stage_opamp_dummy_magic_23_0.X.t42 GNDA 0.053604f
C1779 two_stage_opamp_dummy_magic_23_0.X.t25 GNDA 0.053604f
C1780 two_stage_opamp_dummy_magic_23_0.X.t40 GNDA 0.053604f
C1781 two_stage_opamp_dummy_magic_23_0.X.t54 GNDA 0.053604f
C1782 two_stage_opamp_dummy_magic_23_0.X.t38 GNDA 0.065091f
C1783 two_stage_opamp_dummy_magic_23_0.X.n53 GNDA 0.065091f
C1784 two_stage_opamp_dummy_magic_23_0.X.n54 GNDA 0.042118f
C1785 two_stage_opamp_dummy_magic_23_0.X.n55 GNDA 0.042118f
C1786 two_stage_opamp_dummy_magic_23_0.X.n56 GNDA 0.042118f
C1787 two_stage_opamp_dummy_magic_23_0.X.n57 GNDA 0.042118f
C1788 two_stage_opamp_dummy_magic_23_0.X.n58 GNDA 0.042118f
C1789 two_stage_opamp_dummy_magic_23_0.X.n59 GNDA 0.033981f
C1790 two_stage_opamp_dummy_magic_23_0.X.n60 GNDA 0.021431f
C1791 two_stage_opamp_dummy_magic_23_0.X.t49 GNDA 0.082321f
C1792 two_stage_opamp_dummy_magic_23_0.X.t35 GNDA 0.093585f
C1793 two_stage_opamp_dummy_magic_23_0.X.n61 GNDA 0.076321f
C1794 two_stage_opamp_dummy_magic_23_0.X.t32 GNDA 0.082321f
C1795 two_stage_opamp_dummy_magic_23_0.X.t50 GNDA 0.082321f
C1796 two_stage_opamp_dummy_magic_23_0.X.t33 GNDA 0.082321f
C1797 two_stage_opamp_dummy_magic_23_0.X.t47 GNDA 0.082321f
C1798 two_stage_opamp_dummy_magic_23_0.X.t29 GNDA 0.082321f
C1799 two_stage_opamp_dummy_magic_23_0.X.t43 GNDA 0.082321f
C1800 two_stage_opamp_dummy_magic_23_0.X.t26 GNDA 0.082321f
C1801 two_stage_opamp_dummy_magic_23_0.X.t41 GNDA 0.093585f
C1802 two_stage_opamp_dummy_magic_23_0.X.n62 GNDA 0.084458f
C1803 two_stage_opamp_dummy_magic_23_0.X.n63 GNDA 0.05169f
C1804 two_stage_opamp_dummy_magic_23_0.X.n64 GNDA 0.05169f
C1805 two_stage_opamp_dummy_magic_23_0.X.n65 GNDA 0.05169f
C1806 two_stage_opamp_dummy_magic_23_0.X.n66 GNDA 0.05169f
C1807 two_stage_opamp_dummy_magic_23_0.X.n67 GNDA 0.05169f
C1808 two_stage_opamp_dummy_magic_23_0.X.n68 GNDA 0.043554f
C1809 two_stage_opamp_dummy_magic_23_0.X.n69 GNDA 0.021431f
C1810 two_stage_opamp_dummy_magic_23_0.X.n70 GNDA 0.092553f
C1811 two_stage_opamp_dummy_magic_23_0.X.n71 GNDA 1.05185f
C1812 two_stage_opamp_dummy_magic_23_0.X.n72 GNDA 0.412424f
C1813 two_stage_opamp_dummy_magic_23_0.X.n73 GNDA 0.199954f
C1814 two_stage_opamp_dummy_magic_23_0.Vb1.n0 GNDA 0.03852f
C1815 two_stage_opamp_dummy_magic_23_0.Vb1.n1 GNDA 0.187378f
C1816 two_stage_opamp_dummy_magic_23_0.Vb1.t3 GNDA 0.01284f
C1817 two_stage_opamp_dummy_magic_23_0.Vb1.t0 GNDA 0.01284f
C1818 two_stage_opamp_dummy_magic_23_0.Vb1.n2 GNDA 0.032186f
C1819 two_stage_opamp_dummy_magic_23_0.Vb1.t1 GNDA 0.01284f
C1820 two_stage_opamp_dummy_magic_23_0.Vb1.t2 GNDA 0.01284f
C1821 two_stage_opamp_dummy_magic_23_0.Vb1.n3 GNDA 0.03197f
C1822 two_stage_opamp_dummy_magic_23_0.Vb1.n4 GNDA 0.351059f
C1823 two_stage_opamp_dummy_magic_23_0.Vb1.t28 GNDA 0.601753f
C1824 two_stage_opamp_dummy_magic_23_0.Vb1.n5 GNDA 0.166583f
C1825 two_stage_opamp_dummy_magic_23_0.Vb1.t5 GNDA 0.01926f
C1826 two_stage_opamp_dummy_magic_23_0.Vb1.t9 GNDA 0.01926f
C1827 two_stage_opamp_dummy_magic_23_0.Vb1.n6 GNDA 0.041908f
C1828 two_stage_opamp_dummy_magic_23_0.Vb1.n7 GNDA 0.16835f
C1829 two_stage_opamp_dummy_magic_23_0.Vb1.t10 GNDA 0.019742f
C1830 two_stage_opamp_dummy_magic_23_0.Vb1.t8 GNDA 0.025605f
C1831 two_stage_opamp_dummy_magic_23_0.Vb1.n8 GNDA 0.026326f
C1832 two_stage_opamp_dummy_magic_23_0.Vb1.t6 GNDA 0.019742f
C1833 two_stage_opamp_dummy_magic_23_0.Vb1.t12 GNDA 0.025605f
C1834 two_stage_opamp_dummy_magic_23_0.Vb1.n9 GNDA 0.026326f
C1835 two_stage_opamp_dummy_magic_23_0.Vb1.n10 GNDA 0.019623f
C1836 two_stage_opamp_dummy_magic_23_0.Vb1.t11 GNDA 0.01926f
C1837 two_stage_opamp_dummy_magic_23_0.Vb1.t7 GNDA 0.01926f
C1838 two_stage_opamp_dummy_magic_23_0.Vb1.n11 GNDA 0.041908f
C1839 two_stage_opamp_dummy_magic_23_0.Vb1.n12 GNDA 0.104283f
C1840 two_stage_opamp_dummy_magic_23_0.Vb1.t13 GNDA 0.01926f
C1841 two_stage_opamp_dummy_magic_23_0.Vb1.t4 GNDA 0.01926f
C1842 two_stage_opamp_dummy_magic_23_0.Vb1.n13 GNDA 0.041908f
C1843 two_stage_opamp_dummy_magic_23_0.Vb1.n14 GNDA 0.16835f
C1844 two_stage_opamp_dummy_magic_23_0.Vb1.n15 GNDA 0.299769f
C1845 two_stage_opamp_dummy_magic_23_0.Vb1.t33 GNDA 0.019742f
C1846 two_stage_opamp_dummy_magic_23_0.Vb1.t23 GNDA 0.019742f
C1847 two_stage_opamp_dummy_magic_23_0.Vb1.t31 GNDA 0.019742f
C1848 two_stage_opamp_dummy_magic_23_0.Vb1.t22 GNDA 0.019742f
C1849 two_stage_opamp_dummy_magic_23_0.Vb1.t30 GNDA 0.019742f
C1850 two_stage_opamp_dummy_magic_23_0.Vb1.t20 GNDA 0.019742f
C1851 two_stage_opamp_dummy_magic_23_0.Vb1.t15 GNDA 0.019742f
C1852 two_stage_opamp_dummy_magic_23_0.Vb1.t21 GNDA 0.019742f
C1853 two_stage_opamp_dummy_magic_23_0.Vb1.t29 GNDA 0.019742f
C1854 two_stage_opamp_dummy_magic_23_0.Vb1.t17 GNDA 0.019742f
C1855 two_stage_opamp_dummy_magic_23_0.Vb1.t27 GNDA 0.019742f
C1856 two_stage_opamp_dummy_magic_23_0.Vb1.t16 GNDA 0.019742f
C1857 two_stage_opamp_dummy_magic_23_0.Vb1.t25 GNDA 0.019742f
C1858 two_stage_opamp_dummy_magic_23_0.Vb1.t34 GNDA 0.019742f
C1859 two_stage_opamp_dummy_magic_23_0.Vb1.t26 GNDA 0.019742f
C1860 two_stage_opamp_dummy_magic_23_0.Vb1.t14 GNDA 0.019742f
C1861 two_stage_opamp_dummy_magic_23_0.Vb1.t24 GNDA 0.019742f
C1862 two_stage_opamp_dummy_magic_23_0.Vb1.t32 GNDA 0.019742f
C1863 two_stage_opamp_dummy_magic_23_0.Vb1.t18 GNDA 0.025605f
C1864 two_stage_opamp_dummy_magic_23_0.Vb1.n16 GNDA 0.027841f
C1865 two_stage_opamp_dummy_magic_23_0.Vb1.n17 GNDA 0.018779f
C1866 two_stage_opamp_dummy_magic_23_0.Vb1.n18 GNDA 0.018779f
C1867 two_stage_opamp_dummy_magic_23_0.Vb1.n19 GNDA 0.018779f
C1868 two_stage_opamp_dummy_magic_23_0.Vb1.n20 GNDA 0.018779f
C1869 two_stage_opamp_dummy_magic_23_0.Vb1.n21 GNDA 0.018779f
C1870 two_stage_opamp_dummy_magic_23_0.Vb1.n22 GNDA 0.018779f
C1871 two_stage_opamp_dummy_magic_23_0.Vb1.n23 GNDA 0.018779f
C1872 two_stage_opamp_dummy_magic_23_0.Vb1.n24 GNDA 0.145574f
C1873 two_stage_opamp_dummy_magic_23_0.Vb1.t19 GNDA 0.019742f
C1874 two_stage_opamp_dummy_magic_23_0.Vb1.n25 GNDA 0.145574f
C1875 two_stage_opamp_dummy_magic_23_0.Vb1.n26 GNDA 0.018779f
C1876 two_stage_opamp_dummy_magic_23_0.Vb1.n27 GNDA 0.018779f
C1877 two_stage_opamp_dummy_magic_23_0.Vb1.n28 GNDA 0.018779f
C1878 two_stage_opamp_dummy_magic_23_0.Vb1.n29 GNDA 0.018779f
C1879 two_stage_opamp_dummy_magic_23_0.Vb1.n30 GNDA 0.018779f
C1880 two_stage_opamp_dummy_magic_23_0.Vb1.n31 GNDA 0.018779f
C1881 two_stage_opamp_dummy_magic_23_0.Vb1.n32 GNDA 0.018779f
C1882 two_stage_opamp_dummy_magic_23_0.Vb1.n33 GNDA 0.018779f
C1883 two_stage_opamp_dummy_magic_23_0.Vb1.n34 GNDA 0.033467f
C1884 two_stage_opamp_dummy_magic_23_0.Vb1.n35 GNDA 1.22095f
C1885 bgr_11_0.VB1_CUR_BIAS GNDA 0.83841f
C1886 two_stage_opamp_dummy_magic_23_0.cap_res_X.t70 GNDA 0.344881f
C1887 two_stage_opamp_dummy_magic_23_0.cap_res_X.t103 GNDA 0.346131f
C1888 two_stage_opamp_dummy_magic_23_0.cap_res_X.t101 GNDA 0.344881f
C1889 two_stage_opamp_dummy_magic_23_0.cap_res_X.t4 GNDA 0.347585f
C1890 two_stage_opamp_dummy_magic_23_0.cap_res_X.t118 GNDA 0.378048f
C1891 two_stage_opamp_dummy_magic_23_0.cap_res_X.t107 GNDA 0.344881f
C1892 two_stage_opamp_dummy_magic_23_0.cap_res_X.t9 GNDA 0.346131f
C1893 two_stage_opamp_dummy_magic_23_0.cap_res_X.t62 GNDA 0.344881f
C1894 two_stage_opamp_dummy_magic_23_0.cap_res_X.t26 GNDA 0.346131f
C1895 two_stage_opamp_dummy_magic_23_0.cap_res_X.t138 GNDA 0.344881f
C1896 two_stage_opamp_dummy_magic_23_0.cap_res_X.t38 GNDA 0.346131f
C1897 two_stage_opamp_dummy_magic_23_0.cap_res_X.t13 GNDA 0.344881f
C1898 two_stage_opamp_dummy_magic_23_0.cap_res_X.t117 GNDA 0.346131f
C1899 two_stage_opamp_dummy_magic_23_0.cap_res_X.t43 GNDA 0.344881f
C1900 two_stage_opamp_dummy_magic_23_0.cap_res_X.t73 GNDA 0.346131f
C1901 two_stage_opamp_dummy_magic_23_0.cap_res_X.t57 GNDA 0.344881f
C1902 two_stage_opamp_dummy_magic_23_0.cap_res_X.t17 GNDA 0.346131f
C1903 two_stage_opamp_dummy_magic_23_0.cap_res_X.t3 GNDA 0.344881f
C1904 two_stage_opamp_dummy_magic_23_0.cap_res_X.t45 GNDA 0.346131f
C1905 two_stage_opamp_dummy_magic_23_0.cap_res_X.t19 GNDA 0.344881f
C1906 two_stage_opamp_dummy_magic_23_0.cap_res_X.t122 GNDA 0.346131f
C1907 two_stage_opamp_dummy_magic_23_0.cap_res_X.t49 GNDA 0.344881f
C1908 two_stage_opamp_dummy_magic_23_0.cap_res_X.t81 GNDA 0.346131f
C1909 two_stage_opamp_dummy_magic_23_0.cap_res_X.t61 GNDA 0.344881f
C1910 two_stage_opamp_dummy_magic_23_0.cap_res_X.t25 GNDA 0.346131f
C1911 two_stage_opamp_dummy_magic_23_0.cap_res_X.t85 GNDA 0.344881f
C1912 two_stage_opamp_dummy_magic_23_0.cap_res_X.t114 GNDA 0.346131f
C1913 two_stage_opamp_dummy_magic_23_0.cap_res_X.t97 GNDA 0.344881f
C1914 two_stage_opamp_dummy_magic_23_0.cap_res_X.t63 GNDA 0.346131f
C1915 two_stage_opamp_dummy_magic_23_0.cap_res_X.t52 GNDA 0.344881f
C1916 two_stage_opamp_dummy_magic_23_0.cap_res_X.t86 GNDA 0.346131f
C1917 two_stage_opamp_dummy_magic_23_0.cap_res_X.t64 GNDA 0.344881f
C1918 two_stage_opamp_dummy_magic_23_0.cap_res_X.t33 GNDA 0.346131f
C1919 two_stage_opamp_dummy_magic_23_0.cap_res_X.t89 GNDA 0.344881f
C1920 two_stage_opamp_dummy_magic_23_0.cap_res_X.t119 GNDA 0.346131f
C1921 two_stage_opamp_dummy_magic_23_0.cap_res_X.t99 GNDA 0.344881f
C1922 two_stage_opamp_dummy_magic_23_0.cap_res_X.t68 GNDA 0.346131f
C1923 two_stage_opamp_dummy_magic_23_0.cap_res_X.t129 GNDA 0.344881f
C1924 two_stage_opamp_dummy_magic_23_0.cap_res_X.t24 GNDA 0.346131f
C1925 two_stage_opamp_dummy_magic_23_0.cap_res_X.t5 GNDA 0.344881f
C1926 two_stage_opamp_dummy_magic_23_0.cap_res_X.t104 GNDA 0.346131f
C1927 two_stage_opamp_dummy_magic_23_0.cap_res_X.t95 GNDA 0.344881f
C1928 two_stage_opamp_dummy_magic_23_0.cap_res_X.t130 GNDA 0.346131f
C1929 two_stage_opamp_dummy_magic_23_0.cap_res_X.t106 GNDA 0.344881f
C1930 two_stage_opamp_dummy_magic_23_0.cap_res_X.t78 GNDA 0.346131f
C1931 two_stage_opamp_dummy_magic_23_0.cap_res_X.t135 GNDA 0.344881f
C1932 two_stage_opamp_dummy_magic_23_0.cap_res_X.t30 GNDA 0.346131f
C1933 two_stage_opamp_dummy_magic_23_0.cap_res_X.t10 GNDA 0.344881f
C1934 two_stage_opamp_dummy_magic_23_0.cap_res_X.t111 GNDA 0.346131f
C1935 two_stage_opamp_dummy_magic_23_0.cap_res_X.t37 GNDA 0.344881f
C1936 two_stage_opamp_dummy_magic_23_0.cap_res_X.t67 GNDA 0.346131f
C1937 two_stage_opamp_dummy_magic_23_0.cap_res_X.t54 GNDA 0.344881f
C1938 two_stage_opamp_dummy_magic_23_0.cap_res_X.t12 GNDA 0.346131f
C1939 two_stage_opamp_dummy_magic_23_0.cap_res_X.t72 GNDA 0.344881f
C1940 two_stage_opamp_dummy_magic_23_0.cap_res_X.t102 GNDA 0.346131f
C1941 two_stage_opamp_dummy_magic_23_0.cap_res_X.t91 GNDA 0.344881f
C1942 two_stage_opamp_dummy_magic_23_0.cap_res_X.t56 GNDA 0.346131f
C1943 two_stage_opamp_dummy_magic_23_0.cap_res_X.t44 GNDA 0.344881f
C1944 two_stage_opamp_dummy_magic_23_0.cap_res_X.t74 GNDA 0.346131f
C1945 two_stage_opamp_dummy_magic_23_0.cap_res_X.t55 GNDA 0.344881f
C1946 two_stage_opamp_dummy_magic_23_0.cap_res_X.t18 GNDA 0.346131f
C1947 two_stage_opamp_dummy_magic_23_0.cap_res_X.t96 GNDA 0.344881f
C1948 two_stage_opamp_dummy_magic_23_0.cap_res_X.t51 GNDA 0.346131f
C1949 two_stage_opamp_dummy_magic_23_0.cap_res_X.t84 GNDA 0.344881f
C1950 two_stage_opamp_dummy_magic_23_0.cap_res_X.t110 GNDA 0.361791f
C1951 two_stage_opamp_dummy_magic_23_0.cap_res_X.t36 GNDA 0.344881f
C1952 two_stage_opamp_dummy_magic_23_0.cap_res_X.t71 GNDA 0.185242f
C1953 two_stage_opamp_dummy_magic_23_0.cap_res_X.n0 GNDA 0.198255f
C1954 two_stage_opamp_dummy_magic_23_0.cap_res_X.t105 GNDA 0.344881f
C1955 two_stage_opamp_dummy_magic_23_0.cap_res_X.t7 GNDA 0.185242f
C1956 two_stage_opamp_dummy_magic_23_0.cap_res_X.n1 GNDA 0.196656f
C1957 two_stage_opamp_dummy_magic_23_0.cap_res_X.t76 GNDA 0.344881f
C1958 two_stage_opamp_dummy_magic_23_0.cap_res_X.t60 GNDA 0.185242f
C1959 two_stage_opamp_dummy_magic_23_0.cap_res_X.n2 GNDA 0.196656f
C1960 two_stage_opamp_dummy_magic_23_0.cap_res_X.t23 GNDA 0.344881f
C1961 two_stage_opamp_dummy_magic_23_0.cap_res_X.t15 GNDA 0.185242f
C1962 two_stage_opamp_dummy_magic_23_0.cap_res_X.n3 GNDA 0.196656f
C1963 two_stage_opamp_dummy_magic_23_0.cap_res_X.t128 GNDA 0.344881f
C1964 two_stage_opamp_dummy_magic_23_0.cap_res_X.t66 GNDA 0.185242f
C1965 two_stage_opamp_dummy_magic_23_0.cap_res_X.n4 GNDA 0.196656f
C1966 two_stage_opamp_dummy_magic_23_0.cap_res_X.t94 GNDA 0.344881f
C1967 two_stage_opamp_dummy_magic_23_0.cap_res_X.t115 GNDA 0.185242f
C1968 two_stage_opamp_dummy_magic_23_0.cap_res_X.n5 GNDA 0.196656f
C1969 two_stage_opamp_dummy_magic_23_0.cap_res_X.t59 GNDA 0.344881f
C1970 two_stage_opamp_dummy_magic_23_0.cap_res_X.t31 GNDA 0.185242f
C1971 two_stage_opamp_dummy_magic_23_0.cap_res_X.n6 GNDA 0.196656f
C1972 two_stage_opamp_dummy_magic_23_0.cap_res_X.t6 GNDA 0.344881f
C1973 two_stage_opamp_dummy_magic_23_0.cap_res_X.t126 GNDA 0.185242f
C1974 two_stage_opamp_dummy_magic_23_0.cap_res_X.n7 GNDA 0.196656f
C1975 two_stage_opamp_dummy_magic_23_0.cap_res_X.t109 GNDA 0.344881f
C1976 two_stage_opamp_dummy_magic_23_0.cap_res_X.t42 GNDA 0.185242f
C1977 two_stage_opamp_dummy_magic_23_0.cap_res_X.n8 GNDA 0.196656f
C1978 two_stage_opamp_dummy_magic_23_0.cap_res_X.t133 GNDA 0.344881f
C1979 two_stage_opamp_dummy_magic_23_0.cap_res_X.t28 GNDA 0.346131f
C1980 two_stage_opamp_dummy_magic_23_0.cap_res_X.t80 GNDA 0.166734f
C1981 two_stage_opamp_dummy_magic_23_0.cap_res_X.n9 GNDA 0.215061f
C1982 two_stage_opamp_dummy_magic_23_0.cap_res_X.t90 GNDA 0.184096f
C1983 two_stage_opamp_dummy_magic_23_0.cap_res_X.n10 GNDA 0.23357f
C1984 two_stage_opamp_dummy_magic_23_0.cap_res_X.t121 GNDA 0.184096f
C1985 two_stage_opamp_dummy_magic_23_0.cap_res_X.n11 GNDA 0.250829f
C1986 two_stage_opamp_dummy_magic_23_0.cap_res_X.t16 GNDA 0.184096f
C1987 two_stage_opamp_dummy_magic_23_0.cap_res_X.n12 GNDA 0.250829f
C1988 two_stage_opamp_dummy_magic_23_0.cap_res_X.t116 GNDA 0.184096f
C1989 two_stage_opamp_dummy_magic_23_0.cap_res_X.n13 GNDA 0.250829f
C1990 two_stage_opamp_dummy_magic_23_0.cap_res_X.t83 GNDA 0.184096f
C1991 two_stage_opamp_dummy_magic_23_0.cap_res_X.n14 GNDA 0.250829f
C1992 two_stage_opamp_dummy_magic_23_0.cap_res_X.t47 GNDA 0.184096f
C1993 two_stage_opamp_dummy_magic_23_0.cap_res_X.n15 GNDA 0.250829f
C1994 two_stage_opamp_dummy_magic_23_0.cap_res_X.t77 GNDA 0.184096f
C1995 two_stage_opamp_dummy_magic_23_0.cap_res_X.n16 GNDA 0.250829f
C1996 two_stage_opamp_dummy_magic_23_0.cap_res_X.t39 GNDA 0.184096f
C1997 two_stage_opamp_dummy_magic_23_0.cap_res_X.n17 GNDA 0.250829f
C1998 two_stage_opamp_dummy_magic_23_0.cap_res_X.t136 GNDA 0.184096f
C1999 two_stage_opamp_dummy_magic_23_0.cap_res_X.n18 GNDA 0.250829f
C2000 two_stage_opamp_dummy_magic_23_0.cap_res_X.t32 GNDA 0.184096f
C2001 two_stage_opamp_dummy_magic_23_0.cap_res_X.n19 GNDA 0.250829f
C2002 two_stage_opamp_dummy_magic_23_0.cap_res_X.t131 GNDA 0.184096f
C2003 two_stage_opamp_dummy_magic_23_0.cap_res_X.n20 GNDA 0.250829f
C2004 two_stage_opamp_dummy_magic_23_0.cap_res_X.t92 GNDA 0.184096f
C2005 two_stage_opamp_dummy_magic_23_0.cap_res_X.n21 GNDA 0.250829f
C2006 two_stage_opamp_dummy_magic_23_0.cap_res_X.t120 GNDA 0.184096f
C2007 two_stage_opamp_dummy_magic_23_0.cap_res_X.n22 GNDA 0.250829f
C2008 two_stage_opamp_dummy_magic_23_0.cap_res_X.t87 GNDA 0.184096f
C2009 two_stage_opamp_dummy_magic_23_0.cap_res_X.n23 GNDA 0.250829f
C2010 two_stage_opamp_dummy_magic_23_0.cap_res_X.t125 GNDA 0.184096f
C2011 two_stage_opamp_dummy_magic_23_0.cap_res_X.n24 GNDA 0.250829f
C2012 two_stage_opamp_dummy_magic_23_0.cap_res_X.t88 GNDA 0.184096f
C2013 two_stage_opamp_dummy_magic_23_0.cap_res_X.n25 GNDA 0.23357f
C2014 two_stage_opamp_dummy_magic_23_0.cap_res_X.t20 GNDA 0.343735f
C2015 two_stage_opamp_dummy_magic_23_0.cap_res_X.t123 GNDA 0.166734f
C2016 two_stage_opamp_dummy_magic_23_0.cap_res_X.n26 GNDA 0.216311f
C2017 two_stage_opamp_dummy_magic_23_0.cap_res_X.t58 GNDA 0.343735f
C2018 two_stage_opamp_dummy_magic_23_0.cap_res_X.t22 GNDA 0.166734f
C2019 two_stage_opamp_dummy_magic_23_0.cap_res_X.n27 GNDA 0.216311f
C2020 two_stage_opamp_dummy_magic_23_0.cap_res_X.t41 GNDA 0.343735f
C2021 two_stage_opamp_dummy_magic_23_0.cap_res_X.t100 GNDA 0.344881f
C2022 two_stage_opamp_dummy_magic_23_0.cap_res_X.t65 GNDA 0.36339f
C2023 two_stage_opamp_dummy_magic_23_0.cap_res_X.t48 GNDA 0.36339f
C2024 two_stage_opamp_dummy_magic_23_0.cap_res_X.t2 GNDA 0.185242f
C2025 two_stage_opamp_dummy_magic_23_0.cap_res_X.n28 GNDA 0.216311f
C2026 two_stage_opamp_dummy_magic_23_0.cap_res_X.t21 GNDA 0.343735f
C2027 two_stage_opamp_dummy_magic_23_0.cap_res_X.t29 GNDA 0.344881f
C2028 two_stage_opamp_dummy_magic_23_0.cap_res_X.t124 GNDA 0.185242f
C2029 two_stage_opamp_dummy_magic_23_0.cap_res_X.n29 GNDA 0.197803f
C2030 two_stage_opamp_dummy_magic_23_0.cap_res_X.t50 GNDA 0.343735f
C2031 two_stage_opamp_dummy_magic_23_0.cap_res_X.t53 GNDA 0.344881f
C2032 two_stage_opamp_dummy_magic_23_0.cap_res_X.t8 GNDA 0.185242f
C2033 two_stage_opamp_dummy_magic_23_0.cap_res_X.n30 GNDA 0.216311f
C2034 two_stage_opamp_dummy_magic_23_0.cap_res_X.t27 GNDA 0.343735f
C2035 two_stage_opamp_dummy_magic_23_0.cap_res_X.t35 GNDA 0.344881f
C2036 two_stage_opamp_dummy_magic_23_0.cap_res_X.t132 GNDA 0.185242f
C2037 two_stage_opamp_dummy_magic_23_0.cap_res_X.n31 GNDA 0.216311f
C2038 two_stage_opamp_dummy_magic_23_0.cap_res_X.t127 GNDA 0.343735f
C2039 two_stage_opamp_dummy_magic_23_0.cap_res_X.t134 GNDA 0.344881f
C2040 two_stage_opamp_dummy_magic_23_0.cap_res_X.t93 GNDA 0.185242f
C2041 two_stage_opamp_dummy_magic_23_0.cap_res_X.n32 GNDA 0.216311f
C2042 two_stage_opamp_dummy_magic_23_0.cap_res_X.t11 GNDA 0.343735f
C2043 two_stage_opamp_dummy_magic_23_0.cap_res_X.t69 GNDA 0.344881f
C2044 two_stage_opamp_dummy_magic_23_0.cap_res_X.t34 GNDA 0.36339f
C2045 two_stage_opamp_dummy_magic_23_0.cap_res_X.t14 GNDA 0.36339f
C2046 two_stage_opamp_dummy_magic_23_0.cap_res_X.t112 GNDA 0.185242f
C2047 two_stage_opamp_dummy_magic_23_0.cap_res_X.n33 GNDA 0.216311f
C2048 two_stage_opamp_dummy_magic_23_0.cap_res_X.t108 GNDA 0.343735f
C2049 two_stage_opamp_dummy_magic_23_0.cap_res_X.t40 GNDA 0.344881f
C2050 two_stage_opamp_dummy_magic_23_0.cap_res_X.t137 GNDA 0.36339f
C2051 two_stage_opamp_dummy_magic_23_0.cap_res_X.t113 GNDA 0.36339f
C2052 two_stage_opamp_dummy_magic_23_0.cap_res_X.t79 GNDA 0.185242f
C2053 two_stage_opamp_dummy_magic_23_0.cap_res_X.n34 GNDA 0.216311f
C2054 two_stage_opamp_dummy_magic_23_0.cap_res_X.t75 GNDA 0.343735f
C2055 two_stage_opamp_dummy_magic_23_0.cap_res_X.n35 GNDA 0.216311f
C2056 two_stage_opamp_dummy_magic_23_0.cap_res_X.t46 GNDA 0.185242f
C2057 two_stage_opamp_dummy_magic_23_0.cap_res_X.t82 GNDA 0.36339f
C2058 two_stage_opamp_dummy_magic_23_0.cap_res_X.t98 GNDA 0.36339f
C2059 two_stage_opamp_dummy_magic_23_0.cap_res_X.t1 GNDA 0.736617f
C2060 two_stage_opamp_dummy_magic_23_0.cap_res_X.t0 GNDA 0.297532f
C2061 VOUT-.t7 GNDA 0.047629f
C2062 VOUT-.t1 GNDA 0.047629f
C2063 VOUT-.n0 GNDA 0.097592f
C2064 VOUT-.n1 GNDA 0.249374f
C2065 VOUT-.n2 GNDA 0.03433f
C2066 VOUT-.n3 GNDA 0.060565f
C2067 VOUT-.t14 GNDA 0.047629f
C2068 VOUT-.t4 GNDA 0.047629f
C2069 VOUT-.n4 GNDA 0.097592f
C2070 VOUT-.n5 GNDA 0.290507f
C2071 VOUT-.t13 GNDA 0.047629f
C2072 VOUT-.t3 GNDA 0.047629f
C2073 VOUT-.n6 GNDA 0.097592f
C2074 VOUT-.n7 GNDA 0.285429f
C2075 VOUT-.n8 GNDA 0.060565f
C2076 VOUT-.n9 GNDA 0.03433f
C2077 VOUT-.t6 GNDA 0.047629f
C2078 VOUT-.t12 GNDA 0.047629f
C2079 VOUT-.n10 GNDA 0.097592f
C2080 VOUT-.n11 GNDA 0.285429f
C2081 VOUT-.n12 GNDA 0.03433f
C2082 VOUT-.t8 GNDA 0.047629f
C2083 VOUT-.t2 GNDA 0.047629f
C2084 VOUT-.n13 GNDA 0.097592f
C2085 VOUT-.n14 GNDA 0.285429f
C2086 VOUT-.n15 GNDA 0.03433f
C2087 VOUT-.n16 GNDA 0.060565f
C2088 VOUT-.t5 GNDA 0.047629f
C2089 VOUT-.t15 GNDA 0.047629f
C2090 VOUT-.n17 GNDA 0.097592f
C2091 VOUT-.n18 GNDA 0.290507f
C2092 VOUT-.n19 GNDA 0.050049f
C2093 VOUT-.n20 GNDA 0.198401f
C2094 VOUT-.t24 GNDA 0.322935f
C2095 VOUT-.t129 GNDA 0.317527f
C2096 VOUT-.n21 GNDA 0.212891f
C2097 VOUT-.t77 GNDA 0.317527f
C2098 VOUT-.n22 GNDA 0.138918f
C2099 VOUT-.t61 GNDA 0.322935f
C2100 VOUT-.t106 GNDA 0.317527f
C2101 VOUT-.n23 GNDA 0.212891f
C2102 VOUT-.t67 GNDA 0.317527f
C2103 VOUT-.t48 GNDA 0.322258f
C2104 VOUT-.t151 GNDA 0.322258f
C2105 VOUT-.t98 GNDA 0.322258f
C2106 VOUT-.t63 GNDA 0.322258f
C2107 VOUT-.t29 GNDA 0.322258f
C2108 VOUT-.t134 GNDA 0.322258f
C2109 VOUT-.t81 GNDA 0.322258f
C2110 VOUT-.t52 GNDA 0.322258f
C2111 VOUT-.t121 GNDA 0.322258f
C2112 VOUT-.t73 GNDA 0.322258f
C2113 VOUT-.t47 GNDA 0.317527f
C2114 VOUT-.n24 GNDA 0.213569f
C2115 VOUT-.t86 GNDA 0.317527f
C2116 VOUT-.n25 GNDA 0.273105f
C2117 VOUT-.t150 GNDA 0.317527f
C2118 VOUT-.n26 GNDA 0.273105f
C2119 VOUT-.t97 GNDA 0.317527f
C2120 VOUT-.n27 GNDA 0.273105f
C2121 VOUT-.t142 GNDA 0.317527f
C2122 VOUT-.n28 GNDA 0.273105f
C2123 VOUT-.t91 GNDA 0.317527f
C2124 VOUT-.n29 GNDA 0.273105f
C2125 VOUT-.t42 GNDA 0.317527f
C2126 VOUT-.n30 GNDA 0.273105f
C2127 VOUT-.t126 GNDA 0.317527f
C2128 VOUT-.n31 GNDA 0.273105f
C2129 VOUT-.t31 GNDA 0.317527f
C2130 VOUT-.n32 GNDA 0.273105f
C2131 VOUT-.t115 GNDA 0.317527f
C2132 VOUT-.n33 GNDA 0.273105f
C2133 VOUT-.n34 GNDA 0.257991f
C2134 VOUT-.t113 GNDA 0.322935f
C2135 VOUT-.t83 GNDA 0.317527f
C2136 VOUT-.n35 GNDA 0.212891f
C2137 VOUT-.t36 GNDA 0.317527f
C2138 VOUT-.t102 GNDA 0.322935f
C2139 VOUT-.t139 GNDA 0.317527f
C2140 VOUT-.n36 GNDA 0.212891f
C2141 VOUT-.n37 GNDA 0.257991f
C2142 VOUT-.t85 GNDA 0.322935f
C2143 VOUT-.t55 GNDA 0.317527f
C2144 VOUT-.n38 GNDA 0.212891f
C2145 VOUT-.t141 GNDA 0.317527f
C2146 VOUT-.t66 GNDA 0.322935f
C2147 VOUT-.t101 GNDA 0.317527f
C2148 VOUT-.n39 GNDA 0.212891f
C2149 VOUT-.n40 GNDA 0.257991f
C2150 VOUT-.t120 GNDA 0.322935f
C2151 VOUT-.t90 GNDA 0.317527f
C2152 VOUT-.n41 GNDA 0.212891f
C2153 VOUT-.t41 GNDA 0.317527f
C2154 VOUT-.t103 GNDA 0.322935f
C2155 VOUT-.t145 GNDA 0.317527f
C2156 VOUT-.n42 GNDA 0.212891f
C2157 VOUT-.n43 GNDA 0.257991f
C2158 VOUT-.t22 GNDA 0.322935f
C2159 VOUT-.t127 GNDA 0.317527f
C2160 VOUT-.n44 GNDA 0.212891f
C2161 VOUT-.t74 GNDA 0.317527f
C2162 VOUT-.t147 GNDA 0.322935f
C2163 VOUT-.t46 GNDA 0.317527f
C2164 VOUT-.n45 GNDA 0.212891f
C2165 VOUT-.n46 GNDA 0.257991f
C2166 VOUT-.t56 GNDA 0.322935f
C2167 VOUT-.t153 GNDA 0.317527f
C2168 VOUT-.n47 GNDA 0.212891f
C2169 VOUT-.t39 GNDA 0.317527f
C2170 VOUT-.n48 GNDA 0.138918f
C2171 VOUT-.t87 GNDA 0.322935f
C2172 VOUT-.t54 GNDA 0.317527f
C2173 VOUT-.n49 GNDA 0.212891f
C2174 VOUT-.t69 GNDA 0.317527f
C2175 VOUT-.t137 GNDA 0.322258f
C2176 VOUT-.t99 GNDA 0.322258f
C2177 VOUT-.t57 GNDA 0.322935f
C2178 VOUT-.t92 GNDA 0.317527f
C2179 VOUT-.n50 GNDA 0.212891f
C2180 VOUT-.t109 GNDA 0.317527f
C2181 VOUT-.n51 GNDA 0.133957f
C2182 VOUT-.t116 GNDA 0.322258f
C2183 VOUT-.t156 GNDA 0.322935f
C2184 VOUT-.t59 GNDA 0.317527f
C2185 VOUT-.n52 GNDA 0.212891f
C2186 VOUT-.t75 GNDA 0.317527f
C2187 VOUT-.n53 GNDA 0.133957f
C2188 VOUT-.t82 GNDA 0.322258f
C2189 VOUT-.t117 GNDA 0.322935f
C2190 VOUT-.t20 GNDA 0.317527f
C2191 VOUT-.n54 GNDA 0.212891f
C2192 VOUT-.t44 GNDA 0.317527f
C2193 VOUT-.n55 GNDA 0.133957f
C2194 VOUT-.t49 GNDA 0.322258f
C2195 VOUT-.t88 GNDA 0.322935f
C2196 VOUT-.t123 GNDA 0.317527f
C2197 VOUT-.n56 GNDA 0.212891f
C2198 VOUT-.t143 GNDA 0.317527f
C2199 VOUT-.n57 GNDA 0.133957f
C2200 VOUT-.t146 GNDA 0.322258f
C2201 VOUT-.t23 GNDA 0.322524f
C2202 VOUT-.t30 GNDA 0.322258f
C2203 VOUT-.t122 GNDA 0.322524f
C2204 VOUT-.t130 GNDA 0.322258f
C2205 VOUT-.t104 GNDA 0.322524f
C2206 VOUT-.t107 GNDA 0.322258f
C2207 VOUT-.t128 GNDA 0.322524f
C2208 VOUT-.t136 GNDA 0.322258f
C2209 VOUT-.t33 GNDA 0.317527f
C2210 VOUT-.n58 GNDA 0.351459f
C2211 VOUT-.t149 GNDA 0.317527f
C2212 VOUT-.n59 GNDA 0.410995f
C2213 VOUT-.t25 GNDA 0.317527f
C2214 VOUT-.n60 GNDA 0.410995f
C2215 VOUT-.t64 GNDA 0.317527f
C2216 VOUT-.n61 GNDA 0.410995f
C2217 VOUT-.t45 GNDA 0.317527f
C2218 VOUT-.n62 GNDA 0.337603f
C2219 VOUT-.t78 GNDA 0.317527f
C2220 VOUT-.n63 GNDA 0.337603f
C2221 VOUT-.t111 GNDA 0.317527f
C2222 VOUT-.n64 GNDA 0.337603f
C2223 VOUT-.t155 GNDA 0.317527f
C2224 VOUT-.n65 GNDA 0.337603f
C2225 VOUT-.t135 GNDA 0.317527f
C2226 VOUT-.n66 GNDA 0.273105f
C2227 VOUT-.t34 GNDA 0.317527f
C2228 VOUT-.n67 GNDA 0.273105f
C2229 VOUT-.n68 GNDA 0.257991f
C2230 VOUT-.t50 GNDA 0.322935f
C2231 VOUT-.t148 GNDA 0.317527f
C2232 VOUT-.n69 GNDA 0.212891f
C2233 VOUT-.t32 GNDA 0.317527f
C2234 VOUT-.t95 GNDA 0.322935f
C2235 VOUT-.t131 GNDA 0.317527f
C2236 VOUT-.n70 GNDA 0.212891f
C2237 VOUT-.n71 GNDA 0.257991f
C2238 VOUT-.t19 GNDA 0.322935f
C2239 VOUT-.t119 GNDA 0.317527f
C2240 VOUT-.n72 GNDA 0.212891f
C2241 VOUT-.t70 GNDA 0.317527f
C2242 VOUT-.t144 GNDA 0.322935f
C2243 VOUT-.t40 GNDA 0.317527f
C2244 VOUT-.n73 GNDA 0.212891f
C2245 VOUT-.n74 GNDA 0.257991f
C2246 VOUT-.t114 GNDA 0.322935f
C2247 VOUT-.t84 GNDA 0.317527f
C2248 VOUT-.n75 GNDA 0.212891f
C2249 VOUT-.t37 GNDA 0.317527f
C2250 VOUT-.t100 GNDA 0.322935f
C2251 VOUT-.t140 GNDA 0.317527f
C2252 VOUT-.n76 GNDA 0.212891f
C2253 VOUT-.n77 GNDA 0.257991f
C2254 VOUT-.t154 GNDA 0.322935f
C2255 VOUT-.t112 GNDA 0.317527f
C2256 VOUT-.n78 GNDA 0.212891f
C2257 VOUT-.t65 GNDA 0.317527f
C2258 VOUT-.t138 GNDA 0.322935f
C2259 VOUT-.t35 GNDA 0.317527f
C2260 VOUT-.n79 GNDA 0.212891f
C2261 VOUT-.n80 GNDA 0.257991f
C2262 VOUT-.t108 GNDA 0.322935f
C2263 VOUT-.t76 GNDA 0.317527f
C2264 VOUT-.n81 GNDA 0.212891f
C2265 VOUT-.t26 GNDA 0.317527f
C2266 VOUT-.t96 GNDA 0.322935f
C2267 VOUT-.t132 GNDA 0.317527f
C2268 VOUT-.n82 GNDA 0.212891f
C2269 VOUT-.n83 GNDA 0.257991f
C2270 VOUT-.t72 GNDA 0.322935f
C2271 VOUT-.t43 GNDA 0.317527f
C2272 VOUT-.n84 GNDA 0.212891f
C2273 VOUT-.t125 GNDA 0.317527f
C2274 VOUT-.t60 GNDA 0.322935f
C2275 VOUT-.t94 GNDA 0.317527f
C2276 VOUT-.n85 GNDA 0.212891f
C2277 VOUT-.n86 GNDA 0.257991f
C2278 VOUT-.t105 GNDA 0.322935f
C2279 VOUT-.t71 GNDA 0.317527f
C2280 VOUT-.n87 GNDA 0.212891f
C2281 VOUT-.t21 GNDA 0.317527f
C2282 VOUT-.t93 GNDA 0.322935f
C2283 VOUT-.t124 GNDA 0.317527f
C2284 VOUT-.n88 GNDA 0.212891f
C2285 VOUT-.n89 GNDA 0.257991f
C2286 VOUT-.t68 GNDA 0.322935f
C2287 VOUT-.t38 GNDA 0.317527f
C2288 VOUT-.n90 GNDA 0.212891f
C2289 VOUT-.t118 GNDA 0.317527f
C2290 VOUT-.t58 GNDA 0.322935f
C2291 VOUT-.t89 GNDA 0.317527f
C2292 VOUT-.n91 GNDA 0.212891f
C2293 VOUT-.n92 GNDA 0.257991f
C2294 VOUT-.t28 GNDA 0.322935f
C2295 VOUT-.t133 GNDA 0.317527f
C2296 VOUT-.n93 GNDA 0.212891f
C2297 VOUT-.t80 GNDA 0.317527f
C2298 VOUT-.t152 GNDA 0.322935f
C2299 VOUT-.t53 GNDA 0.317527f
C2300 VOUT-.n94 GNDA 0.212891f
C2301 VOUT-.n95 GNDA 0.257991f
C2302 VOUT-.t62 GNDA 0.322935f
C2303 VOUT-.t27 GNDA 0.317527f
C2304 VOUT-.n96 GNDA 0.212891f
C2305 VOUT-.t110 GNDA 0.317527f
C2306 VOUT-.n97 GNDA 0.257991f
C2307 VOUT-.t79 GNDA 0.317527f
C2308 VOUT-.n98 GNDA 0.138918f
C2309 VOUT-.t51 GNDA 0.317527f
C2310 VOUT-.n99 GNDA 0.252511f
C2311 VOUT-.n100 GNDA 0.309727f
C2312 VOUT-.n101 GNDA 0.084056f
C2313 VOUT-.t11 GNDA 0.055567f
C2314 VOUT-.t16 GNDA 0.055567f
C2315 VOUT-.n102 GNDA 0.119393f
C2316 VOUT-.n103 GNDA 0.333803f
C2317 VOUT-.t18 GNDA 0.055567f
C2318 VOUT-.t10 GNDA 0.055567f
C2319 VOUT-.n104 GNDA 0.119393f
C2320 VOUT-.n105 GNDA 0.321626f
C2321 VOUT-.n106 GNDA 0.11654f
C2322 VOUT-.t17 GNDA 0.055567f
C2323 VOUT-.t0 GNDA 0.055567f
C2324 VOUT-.n107 GNDA 0.119393f
C2325 VOUT-.n108 GNDA 0.326528f
C2326 VOUT-.n109 GNDA 0.056324f
C2327 VOUT-.t9 GNDA 0.091827f
C2328 VOUT-.n110 GNDA 0.111609f
C2329 bgr_11_0.cap_res2.t8 GNDA 0.358376f
C2330 bgr_11_0.cap_res2.t13 GNDA 0.359675f
C2331 bgr_11_0.cap_res2.t3 GNDA 0.340442f
C2332 bgr_11_0.cap_res2.t2 GNDA 0.358376f
C2333 bgr_11_0.cap_res2.t7 GNDA 0.359675f
C2334 bgr_11_0.cap_res2.t17 GNDA 0.340442f
C2335 bgr_11_0.cap_res2.t15 GNDA 0.358376f
C2336 bgr_11_0.cap_res2.t1 GNDA 0.359675f
C2337 bgr_11_0.cap_res2.t11 GNDA 0.340442f
C2338 bgr_11_0.cap_res2.t0 GNDA 0.358376f
C2339 bgr_11_0.cap_res2.t5 GNDA 0.359675f
C2340 bgr_11_0.cap_res2.t16 GNDA 0.340442f
C2341 bgr_11_0.cap_res2.t14 GNDA 0.358376f
C2342 bgr_11_0.cap_res2.t19 GNDA 0.359675f
C2343 bgr_11_0.cap_res2.t9 GNDA 0.340442f
C2344 bgr_11_0.cap_res2.n0 GNDA 0.24022f
C2345 bgr_11_0.cap_res2.t4 GNDA 0.1913f
C2346 bgr_11_0.cap_res2.n1 GNDA 0.260644f
C2347 bgr_11_0.cap_res2.t10 GNDA 0.1913f
C2348 bgr_11_0.cap_res2.n2 GNDA 0.260644f
C2349 bgr_11_0.cap_res2.t6 GNDA 0.1913f
C2350 bgr_11_0.cap_res2.n3 GNDA 0.260644f
C2351 bgr_11_0.cap_res2.t12 GNDA 0.1913f
C2352 bgr_11_0.cap_res2.n4 GNDA 0.260644f
C2353 bgr_11_0.cap_res2.t18 GNDA 0.373116f
C2354 bgr_11_0.cap_res2.t20 GNDA 0.086426f
C2355 bgr_11_0.1st_Vout_2.n0 GNDA 0.878946f
C2356 bgr_11_0.1st_Vout_2.n1 GNDA 0.288815f
C2357 bgr_11_0.1st_Vout_2.n2 GNDA 1.73947f
C2358 bgr_11_0.1st_Vout_2.n3 GNDA 0.126917f
C2359 bgr_11_0.1st_Vout_2.n4 GNDA 1.77207f
C2360 bgr_11_0.1st_Vout_2.n5 GNDA 0.012664f
C2361 bgr_11_0.1st_Vout_2.t6 GNDA 0.018465f
C2362 bgr_11_0.1st_Vout_2.n6 GNDA 0.191552f
C2363 bgr_11_0.1st_Vout_2.n7 GNDA 0.011458f
C2364 bgr_11_0.1st_Vout_2.t31 GNDA 0.021041f
C2365 bgr_11_0.1st_Vout_2.n8 GNDA 0.0221f
C2366 bgr_11_0.1st_Vout_2.t24 GNDA 0.013355f
C2367 bgr_11_0.1st_Vout_2.t12 GNDA 0.013355f
C2368 bgr_11_0.1st_Vout_2.n9 GNDA 0.029711f
C2369 bgr_11_0.1st_Vout_2.t26 GNDA 0.350679f
C2370 bgr_11_0.1st_Vout_2.t18 GNDA 0.356652f
C2371 bgr_11_0.1st_Vout_2.t11 GNDA 0.350679f
C2372 bgr_11_0.1st_Vout_2.t30 GNDA 0.350679f
C2373 bgr_11_0.1st_Vout_2.t23 GNDA 0.356652f
C2374 bgr_11_0.1st_Vout_2.t36 GNDA 0.356652f
C2375 bgr_11_0.1st_Vout_2.t29 GNDA 0.350679f
C2376 bgr_11_0.1st_Vout_2.t22 GNDA 0.350679f
C2377 bgr_11_0.1st_Vout_2.t15 GNDA 0.356652f
C2378 bgr_11_0.1st_Vout_2.t17 GNDA 0.356652f
C2379 bgr_11_0.1st_Vout_2.t35 GNDA 0.350679f
C2380 bgr_11_0.1st_Vout_2.t28 GNDA 0.350679f
C2381 bgr_11_0.1st_Vout_2.t21 GNDA 0.356652f
C2382 bgr_11_0.1st_Vout_2.t34 GNDA 0.356652f
C2383 bgr_11_0.1st_Vout_2.t27 GNDA 0.350679f
C2384 bgr_11_0.1st_Vout_2.t20 GNDA 0.350679f
C2385 bgr_11_0.1st_Vout_2.t14 GNDA 0.356652f
C2386 bgr_11_0.1st_Vout_2.t33 GNDA 0.356652f
C2387 bgr_11_0.1st_Vout_2.t13 GNDA 0.350679f
C2388 bgr_11_0.1st_Vout_2.t19 GNDA 0.350679f
C2389 bgr_11_0.1st_Vout_2.t32 GNDA 0.022909f
C2390 bgr_11_0.1st_Vout_2.n10 GNDA 0.0221f
C2391 bgr_11_0.1st_Vout_2.t25 GNDA 0.013355f
C2392 bgr_11_0.1st_Vout_2.t16 GNDA 0.013355f
C2393 bgr_11_0.1st_Vout_2.n11 GNDA 0.029711f
C2394 bgr_11_0.1st_Vout_2.n12 GNDA 0.021184f
C2395 VOUT+.n0 GNDA 0.08395f
C2396 VOUT+.t16 GNDA 0.055563f
C2397 VOUT+.t2 GNDA 0.055563f
C2398 VOUT+.n1 GNDA 0.119383f
C2399 VOUT+.n2 GNDA 0.333776f
C2400 VOUT+.t1 GNDA 0.055563f
C2401 VOUT+.t15 GNDA 0.055563f
C2402 VOUT+.n3 GNDA 0.119383f
C2403 VOUT+.n4 GNDA 0.321601f
C2404 VOUT+.n5 GNDA 0.116531f
C2405 VOUT+.t18 GNDA 0.055563f
C2406 VOUT+.t0 GNDA 0.055563f
C2407 VOUT+.n6 GNDA 0.119383f
C2408 VOUT+.n7 GNDA 0.327689f
C2409 VOUT+.n8 GNDA 0.060497f
C2410 VOUT+.t17 GNDA 0.091865f
C2411 VOUT+.n9 GNDA 0.11622f
C2412 VOUT+.t5 GNDA 0.047625f
C2413 VOUT+.t10 GNDA 0.047625f
C2414 VOUT+.n10 GNDA 0.097584f
C2415 VOUT+.n11 GNDA 0.249355f
C2416 VOUT+.t13 GNDA 0.047625f
C2417 VOUT+.t11 GNDA 0.047625f
C2418 VOUT+.n12 GNDA 0.097584f
C2419 VOUT+.n13 GNDA 0.290484f
C2420 VOUT+.n14 GNDA 0.034328f
C2421 VOUT+.n15 GNDA 0.06056f
C2422 VOUT+.t4 GNDA 0.047625f
C2423 VOUT+.t14 GNDA 0.047625f
C2424 VOUT+.n16 GNDA 0.097584f
C2425 VOUT+.n17 GNDA 0.290484f
C2426 VOUT+.n18 GNDA 0.06056f
C2427 VOUT+.t6 GNDA 0.047625f
C2428 VOUT+.t9 GNDA 0.047625f
C2429 VOUT+.n19 GNDA 0.097584f
C2430 VOUT+.n20 GNDA 0.285406f
C2431 VOUT+.n21 GNDA 0.06056f
C2432 VOUT+.t7 GNDA 0.047625f
C2433 VOUT+.t12 GNDA 0.047625f
C2434 VOUT+.n22 GNDA 0.097584f
C2435 VOUT+.n23 GNDA 0.285406f
C2436 VOUT+.n24 GNDA 0.034328f
C2437 VOUT+.n25 GNDA 0.034328f
C2438 VOUT+.t8 GNDA 0.047625f
C2439 VOUT+.t3 GNDA 0.047625f
C2440 VOUT+.n26 GNDA 0.097584f
C2441 VOUT+.n27 GNDA 0.285406f
C2442 VOUT+.n28 GNDA 0.034328f
C2443 VOUT+.n29 GNDA 0.050045f
C2444 VOUT+.n30 GNDA 0.198804f
C2445 VOUT+.t63 GNDA 0.317501f
C2446 VOUT+.t35 GNDA 0.322909f
C2447 VOUT+.t34 GNDA 0.317501f
C2448 VOUT+.n31 GNDA 0.212874f
C2449 VOUT+.n32 GNDA 0.138907f
C2450 VOUT+.t99 GNDA 0.322232f
C2451 VOUT+.t149 GNDA 0.322232f
C2452 VOUT+.t43 GNDA 0.322232f
C2453 VOUT+.t77 GNDA 0.322232f
C2454 VOUT+.t125 GNDA 0.322232f
C2455 VOUT+.t20 GNDA 0.322232f
C2456 VOUT+.t59 GNDA 0.322232f
C2457 VOUT+.t92 GNDA 0.322232f
C2458 VOUT+.t143 GNDA 0.322232f
C2459 VOUT+.t39 GNDA 0.322232f
C2460 VOUT+.t95 GNDA 0.317501f
C2461 VOUT+.n33 GNDA 0.213552f
C2462 VOUT+.t146 GNDA 0.317501f
C2463 VOUT+.n34 GNDA 0.273083f
C2464 VOUT+.t107 GNDA 0.317501f
C2465 VOUT+.n35 GNDA 0.273083f
C2466 VOUT+.t153 GNDA 0.317501f
C2467 VOUT+.n36 GNDA 0.273083f
C2468 VOUT+.t65 GNDA 0.317501f
C2469 VOUT+.n37 GNDA 0.273083f
C2470 VOUT+.t113 GNDA 0.317501f
C2471 VOUT+.n38 GNDA 0.273083f
C2472 VOUT+.t72 GNDA 0.317501f
C2473 VOUT+.n39 GNDA 0.273083f
C2474 VOUT+.t120 GNDA 0.317501f
C2475 VOUT+.n40 GNDA 0.273083f
C2476 VOUT+.t31 GNDA 0.317501f
C2477 VOUT+.n41 GNDA 0.273083f
C2478 VOUT+.t132 GNDA 0.317501f
C2479 VOUT+.n42 GNDA 0.273083f
C2480 VOUT+.t45 GNDA 0.317501f
C2481 VOUT+.t58 GNDA 0.322909f
C2482 VOUT+.t147 GNDA 0.317501f
C2483 VOUT+.n43 GNDA 0.212874f
C2484 VOUT+.n44 GNDA 0.25797f
C2485 VOUT+.t103 GNDA 0.322909f
C2486 VOUT+.t49 GNDA 0.317501f
C2487 VOUT+.n45 GNDA 0.212874f
C2488 VOUT+.t152 GNDA 0.317501f
C2489 VOUT+.t130 GNDA 0.322909f
C2490 VOUT+.t127 GNDA 0.317501f
C2491 VOUT+.n46 GNDA 0.212874f
C2492 VOUT+.n47 GNDA 0.25797f
C2493 VOUT+.t67 GNDA 0.322909f
C2494 VOUT+.t155 GNDA 0.317501f
C2495 VOUT+.n48 GNDA 0.212874f
C2496 VOUT+.t116 GNDA 0.317501f
C2497 VOUT+.t98 GNDA 0.322909f
C2498 VOUT+.t96 GNDA 0.317501f
C2499 VOUT+.n49 GNDA 0.212874f
C2500 VOUT+.n50 GNDA 0.25797f
C2501 VOUT+.t109 GNDA 0.322909f
C2502 VOUT+.t55 GNDA 0.317501f
C2503 VOUT+.n51 GNDA 0.212874f
C2504 VOUT+.t19 GNDA 0.317501f
C2505 VOUT+.t136 GNDA 0.322909f
C2506 VOUT+.t134 GNDA 0.317501f
C2507 VOUT+.n52 GNDA 0.212874f
C2508 VOUT+.n53 GNDA 0.25797f
C2509 VOUT+.t145 GNDA 0.322909f
C2510 VOUT+.t93 GNDA 0.317501f
C2511 VOUT+.n54 GNDA 0.212874f
C2512 VOUT+.t60 GNDA 0.317501f
C2513 VOUT+.t32 GNDA 0.322909f
C2514 VOUT+.t30 GNDA 0.317501f
C2515 VOUT+.n55 GNDA 0.212874f
C2516 VOUT+.n56 GNDA 0.25797f
C2517 VOUT+.t36 GNDA 0.317501f
C2518 VOUT+.t66 GNDA 0.322909f
C2519 VOUT+.t28 GNDA 0.317501f
C2520 VOUT+.n57 GNDA 0.212874f
C2521 VOUT+.n58 GNDA 0.138907f
C2522 VOUT+.t75 GNDA 0.322232f
C2523 VOUT+.t53 GNDA 0.322232f
C2524 VOUT+.t137 GNDA 0.322909f
C2525 VOUT+.t33 GNDA 0.317501f
C2526 VOUT+.n59 GNDA 0.212874f
C2527 VOUT+.t86 GNDA 0.317501f
C2528 VOUT+.n60 GNDA 0.133946f
C2529 VOUT+.t90 GNDA 0.322232f
C2530 VOUT+.t27 GNDA 0.322909f
C2531 VOUT+.t69 GNDA 0.317501f
C2532 VOUT+.n61 GNDA 0.212874f
C2533 VOUT+.t122 GNDA 0.317501f
C2534 VOUT+.n62 GNDA 0.133946f
C2535 VOUT+.t126 GNDA 0.322232f
C2536 VOUT+.t81 GNDA 0.322909f
C2537 VOUT+.t119 GNDA 0.317501f
C2538 VOUT+.n63 GNDA 0.212874f
C2539 VOUT+.t106 GNDA 0.317501f
C2540 VOUT+.n64 GNDA 0.133946f
C2541 VOUT+.t110 GNDA 0.322232f
C2542 VOUT+.t114 GNDA 0.322909f
C2543 VOUT+.t156 GNDA 0.317501f
C2544 VOUT+.n65 GNDA 0.212874f
C2545 VOUT+.t140 GNDA 0.317501f
C2546 VOUT+.n66 GNDA 0.133946f
C2547 VOUT+.t148 GNDA 0.322232f
C2548 VOUT+.t37 GNDA 0.322498f
C2549 VOUT+.t44 GNDA 0.322232f
C2550 VOUT+.t76 GNDA 0.322498f
C2551 VOUT+.t82 GNDA 0.322232f
C2552 VOUT+.t56 GNDA 0.322498f
C2553 VOUT+.t61 GNDA 0.322232f
C2554 VOUT+.t91 GNDA 0.322498f
C2555 VOUT+.t100 GNDA 0.322232f
C2556 VOUT+.t131 GNDA 0.317501f
C2557 VOUT+.n67 GNDA 0.351431f
C2558 VOUT+.t94 GNDA 0.317501f
C2559 VOUT+.n68 GNDA 0.410962f
C2560 VOUT+.t115 GNDA 0.317501f
C2561 VOUT+.n69 GNDA 0.410962f
C2562 VOUT+.t78 GNDA 0.317501f
C2563 VOUT+.n70 GNDA 0.410962f
C2564 VOUT+.t42 GNDA 0.317501f
C2565 VOUT+.n71 GNDA 0.337576f
C2566 VOUT+.t141 GNDA 0.317501f
C2567 VOUT+.n72 GNDA 0.337576f
C2568 VOUT+.t22 GNDA 0.317501f
C2569 VOUT+.n73 GNDA 0.337576f
C2570 VOUT+.t124 GNDA 0.317501f
C2571 VOUT+.n74 GNDA 0.337576f
C2572 VOUT+.t87 GNDA 0.317501f
C2573 VOUT+.n75 GNDA 0.273083f
C2574 VOUT+.t112 GNDA 0.317501f
C2575 VOUT+.n76 GNDA 0.273083f
C2576 VOUT+.t71 GNDA 0.317501f
C2577 VOUT+.t105 GNDA 0.322909f
C2578 VOUT+.t68 GNDA 0.317501f
C2579 VOUT+.n77 GNDA 0.212874f
C2580 VOUT+.n78 GNDA 0.25797f
C2581 VOUT+.t48 GNDA 0.322909f
C2582 VOUT+.t70 GNDA 0.317501f
C2583 VOUT+.n79 GNDA 0.212874f
C2584 VOUT+.t29 GNDA 0.317501f
C2585 VOUT+.t62 GNDA 0.322909f
C2586 VOUT+.t24 GNDA 0.317501f
C2587 VOUT+.n80 GNDA 0.212874f
C2588 VOUT+.n81 GNDA 0.25797f
C2589 VOUT+.t139 GNDA 0.322909f
C2590 VOUT+.t88 GNDA 0.317501f
C2591 VOUT+.n82 GNDA 0.212874f
C2592 VOUT+.t54 GNDA 0.317501f
C2593 VOUT+.t26 GNDA 0.322909f
C2594 VOUT+.t25 GNDA 0.317501f
C2595 VOUT+.n83 GNDA 0.212874f
C2596 VOUT+.n84 GNDA 0.25797f
C2597 VOUT+.t104 GNDA 0.322909f
C2598 VOUT+.t51 GNDA 0.317501f
C2599 VOUT+.n85 GNDA 0.212874f
C2600 VOUT+.t154 GNDA 0.317501f
C2601 VOUT+.t129 GNDA 0.322909f
C2602 VOUT+.t128 GNDA 0.317501f
C2603 VOUT+.n86 GNDA 0.212874f
C2604 VOUT+.n87 GNDA 0.25797f
C2605 VOUT+.t135 GNDA 0.322909f
C2606 VOUT+.t83 GNDA 0.317501f
C2607 VOUT+.n88 GNDA 0.212874f
C2608 VOUT+.t50 GNDA 0.317501f
C2609 VOUT+.t23 GNDA 0.322909f
C2610 VOUT+.t21 GNDA 0.317501f
C2611 VOUT+.n89 GNDA 0.212874f
C2612 VOUT+.n90 GNDA 0.25797f
C2613 VOUT+.t97 GNDA 0.322909f
C2614 VOUT+.t46 GNDA 0.317501f
C2615 VOUT+.n91 GNDA 0.212874f
C2616 VOUT+.t150 GNDA 0.317501f
C2617 VOUT+.t123 GNDA 0.322909f
C2618 VOUT+.t121 GNDA 0.317501f
C2619 VOUT+.n92 GNDA 0.212874f
C2620 VOUT+.n93 GNDA 0.25797f
C2621 VOUT+.t57 GNDA 0.322909f
C2622 VOUT+.t144 GNDA 0.317501f
C2623 VOUT+.n94 GNDA 0.212874f
C2624 VOUT+.t111 GNDA 0.317501f
C2625 VOUT+.t85 GNDA 0.322909f
C2626 VOUT+.t84 GNDA 0.317501f
C2627 VOUT+.n95 GNDA 0.212874f
C2628 VOUT+.n96 GNDA 0.25797f
C2629 VOUT+.t89 GNDA 0.322909f
C2630 VOUT+.t38 GNDA 0.317501f
C2631 VOUT+.n97 GNDA 0.212874f
C2632 VOUT+.t142 GNDA 0.317501f
C2633 VOUT+.t118 GNDA 0.322909f
C2634 VOUT+.t117 GNDA 0.317501f
C2635 VOUT+.n98 GNDA 0.212874f
C2636 VOUT+.n99 GNDA 0.25797f
C2637 VOUT+.t52 GNDA 0.322909f
C2638 VOUT+.t138 GNDA 0.317501f
C2639 VOUT+.n100 GNDA 0.212874f
C2640 VOUT+.t108 GNDA 0.317501f
C2641 VOUT+.t80 GNDA 0.322909f
C2642 VOUT+.t79 GNDA 0.317501f
C2643 VOUT+.n101 GNDA 0.212874f
C2644 VOUT+.n102 GNDA 0.25797f
C2645 VOUT+.t151 GNDA 0.322909f
C2646 VOUT+.t102 GNDA 0.317501f
C2647 VOUT+.n103 GNDA 0.212874f
C2648 VOUT+.t64 GNDA 0.317501f
C2649 VOUT+.t41 GNDA 0.322909f
C2650 VOUT+.t40 GNDA 0.317501f
C2651 VOUT+.n104 GNDA 0.212874f
C2652 VOUT+.n105 GNDA 0.25797f
C2653 VOUT+.t74 GNDA 0.322909f
C2654 VOUT+.t73 GNDA 0.317501f
C2655 VOUT+.n106 GNDA 0.212874f
C2656 VOUT+.t101 GNDA 0.317501f
C2657 VOUT+.n107 GNDA 0.25797f
C2658 VOUT+.t133 GNDA 0.317501f
C2659 VOUT+.n108 GNDA 0.138907f
C2660 VOUT+.t47 GNDA 0.317501f
C2661 VOUT+.n109 GNDA 0.252491f
C2662 VOUT+.n110 GNDA 0.308286f
C2663 VDDA.n3 GNDA 0.162507f
C2664 VDDA.n4 GNDA 0.14739f
C2665 VDDA.t480 GNDA 0.153744f
C2666 VDDA.t526 GNDA 0.151169f
C2667 VDDA.n5 GNDA 0.101354f
C2668 VDDA.t559 GNDA 0.151169f
C2669 VDDA.n6 GNDA 0.066136f
C2670 VDDA.t487 GNDA 0.151169f
C2671 VDDA.n7 GNDA 0.066136f
C2672 VDDA.t682 GNDA 0.151169f
C2673 VDDA.n8 GNDA 0.066136f
C2674 VDDA.t724 GNDA 0.151169f
C2675 VDDA.t474 GNDA 0.153744f
C2676 VDDA.t549 GNDA 0.151169f
C2677 VDDA.n9 GNDA 0.101354f
C2678 VDDA.t621 GNDA 0.151169f
C2679 VDDA.n10 GNDA 0.066136f
C2680 VDDA.t577 GNDA 0.151169f
C2681 VDDA.n11 GNDA 0.066136f
C2682 VDDA.t649 GNDA 0.151169f
C2683 VDDA.n12 GNDA 0.066136f
C2684 VDDA.n13 GNDA 0.094481f
C2685 VDDA.t670 GNDA 0.153744f
C2686 VDDA.t716 GNDA 0.151169f
C2687 VDDA.n14 GNDA 0.101354f
C2688 VDDA.t482 GNDA 0.151169f
C2689 VDDA.n15 GNDA 0.066136f
C2690 VDDA.t677 GNDA 0.151169f
C2691 VDDA.n16 GNDA 0.066136f
C2692 VDDA.t603 GNDA 0.151169f
C2693 VDDA.n17 GNDA 0.066136f
C2694 VDDA.t643 GNDA 0.151169f
C2695 VDDA.t662 GNDA 0.153744f
C2696 VDDA.t470 GNDA 0.151169f
C2697 VDDA.n18 GNDA 0.101354f
C2698 VDDA.t545 GNDA 0.151169f
C2699 VDDA.n19 GNDA 0.066136f
C2700 VDDA.t502 GNDA 0.151169f
C2701 VDDA.n20 GNDA 0.066136f
C2702 VDDA.t573 GNDA 0.151169f
C2703 VDDA.n21 GNDA 0.066136f
C2704 VDDA.n22 GNDA 0.122825f
C2705 VDDA.t469 GNDA 0.153744f
C2706 VDDA.t516 GNDA 0.151169f
C2707 VDDA.n23 GNDA 0.101354f
C2708 VDDA.t550 GNDA 0.151169f
C2709 VDDA.n24 GNDA 0.066136f
C2710 VDDA.t476 GNDA 0.151169f
C2711 VDDA.n25 GNDA 0.066136f
C2712 VDDA.t669 GNDA 0.151169f
C2713 VDDA.n26 GNDA 0.066136f
C2714 VDDA.t713 GNDA 0.151169f
C2715 VDDA.t734 GNDA 0.153744f
C2716 VDDA.t540 GNDA 0.151169f
C2717 VDDA.n27 GNDA 0.101354f
C2718 VDDA.t610 GNDA 0.151169f
C2719 VDDA.n28 GNDA 0.066136f
C2720 VDDA.t568 GNDA 0.151169f
C2721 VDDA.n29 GNDA 0.066136f
C2722 VDDA.t639 GNDA 0.151169f
C2723 VDDA.n30 GNDA 0.066136f
C2724 VDDA.n31 GNDA 0.122825f
C2725 VDDA.t659 GNDA 0.153744f
C2726 VDDA.t707 GNDA 0.151169f
C2727 VDDA.n32 GNDA 0.101354f
C2728 VDDA.t472 GNDA 0.151169f
C2729 VDDA.n33 GNDA 0.066136f
C2730 VDDA.t665 GNDA 0.151169f
C2731 VDDA.n34 GNDA 0.066136f
C2732 VDDA.t595 GNDA 0.151169f
C2733 VDDA.n35 GNDA 0.066136f
C2734 VDDA.t635 GNDA 0.151169f
C2735 VDDA.t655 GNDA 0.153744f
C2736 VDDA.t729 GNDA 0.151169f
C2737 VDDA.n36 GNDA 0.101354f
C2738 VDDA.t536 GNDA 0.151169f
C2739 VDDA.n37 GNDA 0.066136f
C2740 VDDA.t494 GNDA 0.151169f
C2741 VDDA.n38 GNDA 0.066136f
C2742 VDDA.t564 GNDA 0.151169f
C2743 VDDA.n39 GNDA 0.066136f
C2744 VDDA.n40 GNDA 0.122825f
C2745 VDDA.t585 GNDA 0.153744f
C2746 VDDA.t628 GNDA 0.151169f
C2747 VDDA.n41 GNDA 0.101354f
C2748 VDDA.t661 GNDA 0.151169f
C2749 VDDA.n42 GNDA 0.066136f
C2750 VDDA.t590 GNDA 0.151169f
C2751 VDDA.n43 GNDA 0.066136f
C2752 VDDA.t521 GNDA 0.151169f
C2753 VDDA.n44 GNDA 0.066136f
C2754 VDDA.t561 GNDA 0.151169f
C2755 VDDA.t580 GNDA 0.153744f
C2756 VDDA.t650 GNDA 0.151169f
C2757 VDDA.n45 GNDA 0.101354f
C2758 VDDA.t727 GNDA 0.151169f
C2759 VDDA.n46 GNDA 0.066136f
C2760 VDDA.t686 GNDA 0.151169f
C2761 VDDA.n47 GNDA 0.066136f
C2762 VDDA.t489 GNDA 0.151169f
C2763 VDDA.n48 GNDA 0.066136f
C2764 VDDA.n49 GNDA 0.122825f
C2765 VDDA.t512 GNDA 0.153744f
C2766 VDDA.t553 GNDA 0.151169f
C2767 VDDA.n50 GNDA 0.101354f
C2768 VDDA.t586 GNDA 0.151169f
C2769 VDDA.n51 GNDA 0.066136f
C2770 VDDA.t517 GNDA 0.151169f
C2771 VDDA.n52 GNDA 0.066136f
C2772 VDDA.t711 GNDA 0.151169f
C2773 VDDA.n53 GNDA 0.066136f
C2774 VDDA.t485 GNDA 0.151169f
C2775 VDDA.t506 GNDA 0.153744f
C2776 VDDA.t576 GNDA 0.151169f
C2777 VDDA.n54 GNDA 0.101354f
C2778 VDDA.t647 GNDA 0.151169f
C2779 VDDA.n55 GNDA 0.066136f
C2780 VDDA.t608 GNDA 0.151169f
C2781 VDDA.n56 GNDA 0.066136f
C2782 VDDA.t680 GNDA 0.151169f
C2783 VDDA.n57 GNDA 0.066136f
C2784 VDDA.n58 GNDA 0.122825f
C2785 VDDA.t575 GNDA 0.153744f
C2786 VDDA.t620 GNDA 0.151169f
C2787 VDDA.n59 GNDA 0.101354f
C2788 VDDA.t651 GNDA 0.151169f
C2789 VDDA.n60 GNDA 0.066136f
C2790 VDDA.t581 GNDA 0.151169f
C2791 VDDA.n61 GNDA 0.066136f
C2792 VDDA.t511 GNDA 0.151169f
C2793 VDDA.n62 GNDA 0.066136f
C2794 VDDA.t554 GNDA 0.151169f
C2795 VDDA.t569 GNDA 0.153744f
C2796 VDDA.t641 GNDA 0.151169f
C2797 VDDA.n63 GNDA 0.101354f
C2798 VDDA.t718 GNDA 0.151169f
C2799 VDDA.n64 GNDA 0.066136f
C2800 VDDA.t673 GNDA 0.151169f
C2801 VDDA.n65 GNDA 0.066136f
C2802 VDDA.t479 GNDA 0.151169f
C2803 VDDA.n66 GNDA 0.066136f
C2804 VDDA.n67 GNDA 0.122825f
C2805 VDDA.t501 GNDA 0.153744f
C2806 VDDA.t544 GNDA 0.151169f
C2807 VDDA.n68 GNDA 0.101354f
C2808 VDDA.t578 GNDA 0.151169f
C2809 VDDA.n69 GNDA 0.066136f
C2810 VDDA.t508 GNDA 0.151169f
C2811 VDDA.n70 GNDA 0.066136f
C2812 VDDA.t702 GNDA 0.151169f
C2813 VDDA.n71 GNDA 0.066136f
C2814 VDDA.t475 GNDA 0.151169f
C2815 VDDA.t495 GNDA 0.153744f
C2816 VDDA.t565 GNDA 0.151169f
C2817 VDDA.n72 GNDA 0.101354f
C2818 VDDA.t638 GNDA 0.151169f
C2819 VDDA.n73 GNDA 0.066136f
C2820 VDDA.t597 GNDA 0.151169f
C2821 VDDA.n74 GNDA 0.066136f
C2822 VDDA.t668 GNDA 0.151169f
C2823 VDDA.n75 GNDA 0.066136f
C2824 VDDA.n76 GNDA 0.122825f
C2825 VDDA.t694 GNDA 0.153744f
C2826 VDDA.t735 GNDA 0.151169f
C2827 VDDA.n77 GNDA 0.101354f
C2828 VDDA.t503 GNDA 0.151169f
C2829 VDDA.n78 GNDA 0.066136f
C2830 VDDA.t699 GNDA 0.151169f
C2831 VDDA.n79 GNDA 0.066136f
C2832 VDDA.t625 GNDA 0.151169f
C2833 VDDA.n80 GNDA 0.066136f
C2834 VDDA.t663 GNDA 0.151169f
C2835 VDDA.t688 GNDA 0.153744f
C2836 VDDA.t492 GNDA 0.151169f
C2837 VDDA.n81 GNDA 0.101354f
C2838 VDDA.t563 GNDA 0.151169f
C2839 VDDA.n82 GNDA 0.066136f
C2840 VDDA.t523 GNDA 0.151169f
C2841 VDDA.n83 GNDA 0.066136f
C2842 VDDA.t594 GNDA 0.151169f
C2843 VDDA.n84 GNDA 0.066136f
C2844 VDDA.n85 GNDA 0.122825f
C2845 VDDA.t491 GNDA 0.153744f
C2846 VDDA.t535 GNDA 0.151169f
C2847 VDDA.n86 GNDA 0.101354f
C2848 VDDA.t566 GNDA 0.151169f
C2849 VDDA.n87 GNDA 0.066136f
C2850 VDDA.t496 GNDA 0.151169f
C2851 VDDA.n88 GNDA 0.066136f
C2852 VDDA.t693 GNDA 0.151169f
C2853 VDDA.n89 GNDA 0.066136f
C2854 VDDA.t731 GNDA 0.151169f
C2855 VDDA.t486 GNDA 0.153744f
C2856 VDDA.t558 GNDA 0.151169f
C2857 VDDA.n90 GNDA 0.101354f
C2858 VDDA.t630 GNDA 0.151169f
C2859 VDDA.n91 GNDA 0.066136f
C2860 VDDA.t588 GNDA 0.151169f
C2861 VDDA.n92 GNDA 0.066136f
C2862 VDDA.t658 GNDA 0.151169f
C2863 VDDA.n93 GNDA 0.066136f
C2864 VDDA.n94 GNDA 0.122825f
C2865 VDDA.t683 GNDA 0.153744f
C2866 VDDA.t726 GNDA 0.151169f
C2867 VDDA.n95 GNDA 0.101354f
C2868 VDDA.t493 GNDA 0.151169f
C2869 VDDA.n96 GNDA 0.066136f
C2870 VDDA.t689 GNDA 0.151169f
C2871 VDDA.n97 GNDA 0.066136f
C2872 VDDA.t615 GNDA 0.151169f
C2873 VDDA.n98 GNDA 0.066136f
C2874 VDDA.t654 GNDA 0.151169f
C2875 VDDA.t675 GNDA 0.153744f
C2876 VDDA.t481 GNDA 0.151169f
C2877 VDDA.n99 GNDA 0.101354f
C2878 VDDA.t556 GNDA 0.151169f
C2879 VDDA.n100 GNDA 0.066136f
C2880 VDDA.t514 GNDA 0.151169f
C2881 VDDA.n101 GNDA 0.066136f
C2882 VDDA.t584 GNDA 0.151169f
C2883 VDDA.n102 GNDA 0.066136f
C2884 VDDA.n103 GNDA 0.122825f
C2885 VDDA.t606 GNDA 0.153744f
C2886 VDDA.t646 GNDA 0.151169f
C2887 VDDA.n104 GNDA 0.101354f
C2888 VDDA.t684 GNDA 0.151169f
C2889 VDDA.n105 GNDA 0.066136f
C2890 VDDA.t611 GNDA 0.151169f
C2891 VDDA.n106 GNDA 0.066136f
C2892 VDDA.t541 GNDA 0.151169f
C2893 VDDA.n107 GNDA 0.066136f
C2894 VDDA.t579 GNDA 0.151169f
C2895 VDDA.t600 GNDA 0.153744f
C2896 VDDA.t672 GNDA 0.151169f
C2897 VDDA.n108 GNDA 0.101354f
C2898 VDDA.t478 GNDA 0.151169f
C2899 VDDA.n109 GNDA 0.066136f
C2900 VDDA.t705 GNDA 0.151169f
C2901 VDDA.n110 GNDA 0.066136f
C2902 VDDA.t510 GNDA 0.151169f
C2903 VDDA.n111 GNDA 0.066136f
C2904 VDDA.n112 GNDA 0.122825f
C2905 VDDA.t671 GNDA 0.153744f
C2906 VDDA.t717 GNDA 0.151169f
C2907 VDDA.n113 GNDA 0.101354f
C2908 VDDA.t483 GNDA 0.151169f
C2909 VDDA.n114 GNDA 0.066136f
C2910 VDDA.t678 GNDA 0.151169f
C2911 VDDA.n115 GNDA 0.066136f
C2912 VDDA.t604 GNDA 0.151169f
C2913 VDDA.n116 GNDA 0.066136f
C2914 VDDA.t644 GNDA 0.151169f
C2915 VDDA.t664 GNDA 0.153744f
C2916 VDDA.t471 GNDA 0.151169f
C2917 VDDA.n117 GNDA 0.101354f
C2918 VDDA.t546 GNDA 0.151169f
C2919 VDDA.n118 GNDA 0.066136f
C2920 VDDA.t504 GNDA 0.151169f
C2921 VDDA.n119 GNDA 0.066136f
C2922 VDDA.t574 GNDA 0.151169f
C2923 VDDA.n120 GNDA 0.066136f
C2924 VDDA.n121 GNDA 0.122825f
C2925 VDDA.t596 GNDA 0.153744f
C2926 VDDA.t637 GNDA 0.151169f
C2927 VDDA.n122 GNDA 0.101354f
C2928 VDDA.t674 GNDA 0.151169f
C2929 VDDA.n123 GNDA 0.066136f
C2930 VDDA.t602 GNDA 0.151169f
C2931 VDDA.n124 GNDA 0.066136f
C2932 VDDA.t530 GNDA 0.151169f
C2933 VDDA.n125 GNDA 0.066136f
C2934 VDDA.t570 GNDA 0.151169f
C2935 VDDA.t589 GNDA 0.153744f
C2936 VDDA.t660 GNDA 0.151169f
C2937 VDDA.n126 GNDA 0.101354f
C2938 VDDA.t736 GNDA 0.151169f
C2939 VDDA.n127 GNDA 0.066136f
C2940 VDDA.t695 GNDA 0.151169f
C2941 VDDA.n128 GNDA 0.066136f
C2942 VDDA.t500 GNDA 0.151169f
C2943 VDDA.n129 GNDA 0.066136f
C2944 VDDA.n130 GNDA 0.122825f
C2945 VDDA.t532 GNDA 0.153744f
C2946 VDDA.t571 GNDA 0.151169f
C2947 VDDA.n131 GNDA 0.101354f
C2948 VDDA.t609 GNDA 0.151169f
C2949 VDDA.n132 GNDA 0.066136f
C2950 VDDA.t538 GNDA 0.151169f
C2951 VDDA.n133 GNDA 0.066136f
C2952 VDDA.t730 GNDA 0.151169f
C2953 VDDA.n134 GNDA 0.066136f
C2954 VDDA.t507 GNDA 0.151169f
C2955 VDDA.t528 GNDA 0.153744f
C2956 VDDA.t598 GNDA 0.151169f
C2957 VDDA.n135 GNDA 0.101354f
C2958 VDDA.t667 GNDA 0.151169f
C2959 VDDA.n136 GNDA 0.066136f
C2960 VDDA.t629 GNDA 0.151169f
C2961 VDDA.n137 GNDA 0.066136f
C2962 VDDA.t701 GNDA 0.151169f
C2963 VDDA.n138 GNDA 0.066136f
C2964 VDDA.n139 GNDA 0.122825f
C2965 VDDA.t723 GNDA 0.153744f
C2966 VDDA.t498 GNDA 0.151169f
C2967 VDDA.n140 GNDA 0.101354f
C2968 VDDA.t533 GNDA 0.151169f
C2969 VDDA.n141 GNDA 0.066136f
C2970 VDDA.t728 GNDA 0.151169f
C2971 VDDA.n142 GNDA 0.066136f
C2972 VDDA.t652 GNDA 0.151169f
C2973 VDDA.n143 GNDA 0.066136f
C2974 VDDA.t698 GNDA 0.151169f
C2975 VDDA.t719 GNDA 0.153744f
C2976 VDDA.t524 GNDA 0.151169f
C2977 VDDA.n144 GNDA 0.101354f
C2978 VDDA.t593 GNDA 0.151169f
C2979 VDDA.n145 GNDA 0.066136f
C2980 VDDA.t555 GNDA 0.151169f
C2981 VDDA.n146 GNDA 0.066136f
C2982 VDDA.t624 GNDA 0.151169f
C2983 VDDA.n147 GNDA 0.066136f
C2984 VDDA.n148 GNDA 0.122825f
C2985 VDDA.t522 GNDA 0.153744f
C2986 VDDA.t562 GNDA 0.151169f
C2987 VDDA.n149 GNDA 0.101354f
C2988 VDDA.t599 GNDA 0.151169f
C2989 VDDA.n150 GNDA 0.066136f
C2990 VDDA.t529 GNDA 0.151169f
C2991 VDDA.n151 GNDA 0.066136f
C2992 VDDA.t722 GNDA 0.151169f
C2993 VDDA.n152 GNDA 0.066136f
C2994 VDDA.t497 GNDA 0.151169f
C2995 VDDA.t519 GNDA 0.153744f
C2996 VDDA.t587 GNDA 0.151169f
C2997 VDDA.n153 GNDA 0.101354f
C2998 VDDA.t657 GNDA 0.151169f
C2999 VDDA.n154 GNDA 0.066136f
C3000 VDDA.t619 GNDA 0.151169f
C3001 VDDA.n155 GNDA 0.066136f
C3002 VDDA.t692 GNDA 0.151169f
C3003 VDDA.n156 GNDA 0.066136f
C3004 VDDA.n157 GNDA 0.122825f
C3005 VDDA.t712 GNDA 0.153744f
C3006 VDDA.t488 GNDA 0.151169f
C3007 VDDA.n158 GNDA 0.101354f
C3008 VDDA.t525 GNDA 0.151169f
C3009 VDDA.n159 GNDA 0.066136f
C3010 VDDA.t720 GNDA 0.151169f
C3011 VDDA.n160 GNDA 0.066136f
C3012 VDDA.t642 GNDA 0.151169f
C3013 VDDA.n161 GNDA 0.066136f
C3014 VDDA.t690 GNDA 0.151169f
C3015 VDDA.t708 GNDA 0.153744f
C3016 VDDA.t513 GNDA 0.151169f
C3017 VDDA.n162 GNDA 0.101354f
C3018 VDDA.t583 GNDA 0.151169f
C3019 VDDA.n163 GNDA 0.066136f
C3020 VDDA.t543 GNDA 0.151169f
C3021 VDDA.n164 GNDA 0.066136f
C3022 VDDA.t614 GNDA 0.151169f
C3023 VDDA.n165 GNDA 0.066136f
C3024 VDDA.n166 GNDA 0.122825f
C3025 VDDA.t634 GNDA 0.153744f
C3026 VDDA.t679 GNDA 0.151169f
C3027 VDDA.n167 GNDA 0.101354f
C3028 VDDA.t715 GNDA 0.151169f
C3029 VDDA.n168 GNDA 0.066136f
C3030 VDDA.t640 GNDA 0.151169f
C3031 VDDA.n169 GNDA 0.066136f
C3032 VDDA.t567 GNDA 0.151169f
C3033 VDDA.n170 GNDA 0.066136f
C3034 VDDA.t612 GNDA 0.151169f
C3035 VDDA.t631 GNDA 0.153744f
C3036 VDDA.t704 GNDA 0.151169f
C3037 VDDA.n171 GNDA 0.101354f
C3038 VDDA.t509 GNDA 0.151169f
C3039 VDDA.n172 GNDA 0.066136f
C3040 VDDA.t732 GNDA 0.151169f
C3041 VDDA.n173 GNDA 0.066136f
C3042 VDDA.t539 GNDA 0.151169f
C3043 VDDA.n174 GNDA 0.066136f
C3044 VDDA.n175 GNDA 0.122825f
C3045 VDDA.t703 GNDA 0.153744f
C3046 VDDA.t477 GNDA 0.151169f
C3047 VDDA.n176 GNDA 0.101354f
C3048 VDDA.t515 GNDA 0.151169f
C3049 VDDA.n177 GNDA 0.066136f
C3050 VDDA.t709 GNDA 0.151169f
C3051 VDDA.n178 GNDA 0.066136f
C3052 VDDA.t633 GNDA 0.151169f
C3053 VDDA.n179 GNDA 0.066136f
C3054 VDDA.t676 GNDA 0.151169f
C3055 VDDA.t700 GNDA 0.153744f
C3056 VDDA.t505 GNDA 0.151169f
C3057 VDDA.n180 GNDA 0.101354f
C3058 VDDA.t572 GNDA 0.151169f
C3059 VDDA.n181 GNDA 0.066136f
C3060 VDDA.t534 GNDA 0.151169f
C3061 VDDA.n182 GNDA 0.066136f
C3062 VDDA.t605 GNDA 0.151169f
C3063 VDDA.n183 GNDA 0.066136f
C3064 VDDA.n184 GNDA 0.122825f
C3065 VDDA.t626 GNDA 0.153744f
C3066 VDDA.t666 GNDA 0.151169f
C3067 VDDA.n185 GNDA 0.101354f
C3068 VDDA.t706 GNDA 0.151169f
C3069 VDDA.n186 GNDA 0.066136f
C3070 VDDA.t632 GNDA 0.151169f
C3071 VDDA.n187 GNDA 0.066136f
C3072 VDDA.t560 GNDA 0.151169f
C3073 VDDA.n188 GNDA 0.066136f
C3074 VDDA.t601 GNDA 0.151169f
C3075 VDDA.t622 GNDA 0.153744f
C3076 VDDA.t696 GNDA 0.151169f
C3077 VDDA.n189 GNDA 0.101354f
C3078 VDDA.t499 GNDA 0.151169f
C3079 VDDA.n190 GNDA 0.066136f
C3080 VDDA.t725 GNDA 0.151169f
C3081 VDDA.n191 GNDA 0.066136f
C3082 VDDA.t531 GNDA 0.151169f
C3083 VDDA.n192 GNDA 0.066136f
C3084 VDDA.n193 GNDA 0.122825f
C3085 VDDA.t552 GNDA 0.153744f
C3086 VDDA.t592 GNDA 0.151169f
C3087 VDDA.n194 GNDA 0.101354f
C3088 VDDA.t627 GNDA 0.151169f
C3089 VDDA.n195 GNDA 0.066136f
C3090 VDDA.t557 GNDA 0.151169f
C3091 VDDA.n196 GNDA 0.066136f
C3092 VDDA.t484 GNDA 0.151169f
C3093 VDDA.n197 GNDA 0.066136f
C3094 VDDA.t527 GNDA 0.151169f
C3095 VDDA.t547 GNDA 0.153744f
C3096 VDDA.t617 GNDA 0.151169f
C3097 VDDA.n198 GNDA 0.101354f
C3098 VDDA.t691 GNDA 0.151169f
C3099 VDDA.n199 GNDA 0.066136f
C3100 VDDA.t645 GNDA 0.151169f
C3101 VDDA.n200 GNDA 0.066136f
C3102 VDDA.t721 GNDA 0.151169f
C3103 VDDA.n201 GNDA 0.066136f
C3104 VDDA.n202 GNDA 0.122825f
C3105 VDDA.t616 GNDA 0.153744f
C3106 VDDA.t656 GNDA 0.151169f
C3107 VDDA.n203 GNDA 0.101354f
C3108 VDDA.t697 GNDA 0.151169f
C3109 VDDA.n204 GNDA 0.066136f
C3110 VDDA.t623 GNDA 0.151169f
C3111 VDDA.n205 GNDA 0.066136f
C3112 VDDA.t551 GNDA 0.151169f
C3113 VDDA.n206 GNDA 0.066136f
C3114 VDDA.t591 GNDA 0.151169f
C3115 VDDA.t613 GNDA 0.153744f
C3116 VDDA.t685 GNDA 0.151169f
C3117 VDDA.n207 GNDA 0.101354f
C3118 VDDA.t490 GNDA 0.151169f
C3119 VDDA.n208 GNDA 0.066136f
C3120 VDDA.t714 GNDA 0.151169f
C3121 VDDA.n209 GNDA 0.066136f
C3122 VDDA.t520 GNDA 0.151169f
C3123 VDDA.n210 GNDA 0.066136f
C3124 VDDA.n211 GNDA 0.122825f
C3125 VDDA.t542 GNDA 0.153744f
C3126 VDDA.t582 GNDA 0.151169f
C3127 VDDA.n212 GNDA 0.101354f
C3128 VDDA.t618 GNDA 0.151169f
C3129 VDDA.n213 GNDA 0.066136f
C3130 VDDA.t548 GNDA 0.151169f
C3131 VDDA.n214 GNDA 0.066136f
C3132 VDDA.t473 GNDA 0.151169f
C3133 VDDA.n215 GNDA 0.066136f
C3134 VDDA.t518 GNDA 0.151169f
C3135 VDDA.n216 GNDA 0.094481f
C3136 VDDA.t710 GNDA 0.151169f
C3137 VDDA.n217 GNDA 0.066136f
C3138 VDDA.t636 GNDA 0.151169f
C3139 VDDA.n218 GNDA 0.066136f
C3140 VDDA.t681 GNDA 0.151169f
C3141 VDDA.n219 GNDA 0.066136f
C3142 VDDA.t607 GNDA 0.151169f
C3143 VDDA.n220 GNDA 0.066136f
C3144 VDDA.t537 GNDA 0.151169f
C3145 VDDA.n221 GNDA 0.065321f
C3146 VDDA.n222 GNDA 0.014172f
C3147 VDDA.n225 GNDA 0.015306f
C3148 VDDA.n226 GNDA 0.015306f
C3149 VDDA.n227 GNDA 0.015873f
C3150 VDDA.n228 GNDA 0.014172f
C3151 VDDA.t733 GNDA 0.428762f
C3152 VDDA.t687 GNDA 0.445304f
C3153 VDDA.n229 GNDA 0.302641f
C3154 VDDA.t648 GNDA 0.44513f
C3155 VDDA.n230 GNDA 0.144475f
C3156 VDDA.t653 GNDA 0.417598f
C3157 VDDA.n231 GNDA 0.293881f
C3158 VDDA.n232 GNDA 0.323182f
C3159 VDDA.n233 GNDA 0.015306f
C3160 VDDA.n234 GNDA 0.015306f
C3161 VDDA.n235 GNDA 0.015306f
C3162 VDDA.n236 GNDA 0.015873f
C3163 VDDA.n237 GNDA 0.015873f
C3164 VDDA.n238 GNDA 0.015873f
C3165 VDDA.n239 GNDA 0.015873f
C3166 VDDA.n240 GNDA 0.043168f
C3167 VDDA.n241 GNDA 0.016069f
C3168 VDDA.n242 GNDA 0.014458f
C3169 VDDA.n243 GNDA 0.295595f
C3170 VDDA.n244 GNDA 0.014172f
C3171 VDDA.n247 GNDA 0.015306f
C3172 VDDA.n248 GNDA 0.015306f
C3173 VDDA.n249 GNDA 0.015873f
C3174 VDDA.n250 GNDA 0.014172f
C3175 VDDA.n252 GNDA 0.038491f
C3176 VDDA.n253 GNDA 0.015983f
C3177 VDDA.t335 GNDA 0.013146f
C3178 VDDA.n256 GNDA 0.038491f
C3179 VDDA.n258 GNDA 0.038491f
C3180 VDDA.n260 GNDA 0.038491f
C3181 VDDA.n262 GNDA 0.038491f
C3182 VDDA.n264 GNDA 0.038491f
C3183 VDDA.n266 GNDA 0.038491f
C3184 VDDA.n268 GNDA 0.038491f
C3185 VDDA.n270 GNDA 0.038491f
C3186 VDDA.n272 GNDA 0.038491f
C3187 VDDA.n273 GNDA 0.015983f
C3188 VDDA.t390 GNDA 0.013146f
C3189 VDDA.n275 GNDA 0.015983f
C3190 VDDA.n277 GNDA 0.038491f
C3191 VDDA.n279 GNDA 0.038491f
C3192 VDDA.n281 GNDA 0.038491f
C3193 VDDA.n283 GNDA 0.038491f
C3194 VDDA.n285 GNDA 0.038491f
C3195 VDDA.n287 GNDA 0.038491f
C3196 VDDA.n289 GNDA 0.038491f
C3197 VDDA.n291 GNDA 0.055313f
C3198 VDDA.n292 GNDA 0.014655f
C3199 VDDA.t373 GNDA 0.013944f
C3200 VDDA.t375 GNDA 0.013146f
C3201 VDDA.n294 GNDA 0.025299f
C3202 VDDA.n295 GNDA 0.046585f
C3203 VDDA.t374 GNDA 0.03922f
C3204 VDDA.t81 GNDA 0.031746f
C3205 VDDA.t126 GNDA 0.031746f
C3206 VDDA.t98 GNDA 0.031746f
C3207 VDDA.t219 GNDA 0.031746f
C3208 VDDA.t438 GNDA 0.031746f
C3209 VDDA.t65 GNDA 0.031746f
C3210 VDDA.t41 GNDA 0.031746f
C3211 VDDA.t83 GNDA 0.031746f
C3212 VDDA.t0 GNDA 0.031746f
C3213 VDDA.t460 GNDA 0.031746f
C3214 VDDA.t7 GNDA 0.031746f
C3215 VDDA.t70 GNDA 0.031746f
C3216 VDDA.t63 GNDA 0.031746f
C3217 VDDA.t116 GNDA 0.031746f
C3218 VDDA.t227 GNDA 0.031746f
C3219 VDDA.t51 GNDA 0.031746f
C3220 VDDA.t443 GNDA 0.031746f
C3221 VDDA.t79 GNDA 0.031746f
C3222 VDDA.t389 GNDA 0.03922f
C3223 VDDA.n296 GNDA 0.046585f
C3224 VDDA.n297 GNDA 0.025198f
C3225 VDDA.t388 GNDA 0.013951f
C3226 VDDA.n298 GNDA 0.013907f
C3227 VDDA.n299 GNDA 0.028152f
C3228 VDDA.n300 GNDA 0.028152f
C3229 VDDA.n301 GNDA 0.01546f
C3230 VDDA.t381 GNDA 0.013237f
C3231 VDDA.n302 GNDA 0.068949f
C3232 VDDA.t380 GNDA 0.048423f
C3233 VDDA.t107 GNDA 0.031746f
C3234 VDDA.t134 GNDA 0.031746f
C3235 VDDA.t20 GNDA 0.031746f
C3236 VDDA.t25 GNDA 0.031746f
C3237 VDDA.t235 GNDA 0.031746f
C3238 VDDA.t5 GNDA 0.031746f
C3239 VDDA.t114 GNDA 0.031746f
C3240 VDDA.t243 GNDA 0.031746f
C3241 VDDA.t432 GNDA 0.031746f
C3242 VDDA.t112 GNDA 0.031746f
C3243 VDDA.t267 GNDA 0.031746f
C3244 VDDA.t61 GNDA 0.031746f
C3245 VDDA.t105 GNDA 0.031746f
C3246 VDDA.t38 GNDA 0.031746f
C3247 VDDA.t249 GNDA 0.031746f
C3248 VDDA.t245 GNDA 0.031746f
C3249 VDDA.t424 GNDA 0.031746f
C3250 VDDA.t30 GNDA 0.031746f
C3251 VDDA.t334 GNDA 0.03922f
C3252 VDDA.n303 GNDA 0.046585f
C3253 VDDA.n304 GNDA 0.025198f
C3254 VDDA.t333 GNDA 0.013951f
C3255 VDDA.n305 GNDA 0.013907f
C3256 VDDA.n306 GNDA 0.105725f
C3257 VDDA.n307 GNDA 0.219285f
C3258 VDDA.n308 GNDA 0.015306f
C3259 VDDA.n309 GNDA 0.015306f
C3260 VDDA.n310 GNDA 0.015306f
C3261 VDDA.n311 GNDA 0.015873f
C3262 VDDA.n312 GNDA 0.015873f
C3263 VDDA.n313 GNDA 0.015873f
C3264 VDDA.n314 GNDA 0.015873f
C3265 VDDA.n315 GNDA 0.043168f
C3266 VDDA.n316 GNDA 0.016069f
C3267 VDDA.n317 GNDA 0.014458f
C3268 VDDA.n318 GNDA 1.60239f
C3269 VDDA.n319 GNDA 0.01181f
C3270 VDDA.n322 GNDA 0.012755f
C3271 VDDA.n323 GNDA 0.012755f
C3272 VDDA.n324 GNDA 0.013227f
C3273 VDDA.n325 GNDA 0.01181f
C3274 VDDA.n327 GNDA 0.033295f
C3275 VDDA.n329 GNDA 0.033278f
C3276 VDDA.t344 GNDA 0.013778f
C3277 VDDA.t420 GNDA 0.013778f
C3278 VDDA.n331 GNDA 0.045545f
C3279 VDDA.n332 GNDA 0.015807f
C3280 VDDA.n333 GNDA 0.039346f
C3281 VDDA.t419 GNDA 0.041458f
C3282 VDDA.t118 GNDA 0.0291f
C3283 VDDA.t225 GNDA 0.0291f
C3284 VDDA.t456 GNDA 0.0291f
C3285 VDDA.t449 GNDA 0.0291f
C3286 VDDA.t343 GNDA 0.041458f
C3287 VDDA.n334 GNDA 0.039346f
C3288 VDDA.n335 GNDA 0.015307f
C3289 VDDA.n336 GNDA 0.022971f
C3290 VDDA.n338 GNDA 0.033274f
C3291 VDDA.t323 GNDA 0.013786f
C3292 VDDA.t402 GNDA 0.013786f
C3293 VDDA.n340 GNDA 0.045541f
C3294 VDDA.n341 GNDA 0.015807f
C3295 VDDA.n342 GNDA 0.039339f
C3296 VDDA.t401 GNDA 0.041458f
C3297 VDDA.t11 GNDA 0.0291f
C3298 VDDA.t147 GNDA 0.0291f
C3299 VDDA.t47 GNDA 0.0291f
C3300 VDDA.t45 GNDA 0.0291f
C3301 VDDA.t322 GNDA 0.041458f
C3302 VDDA.n343 GNDA 0.039339f
C3303 VDDA.n344 GNDA 0.015543f
C3304 VDDA.n345 GNDA 0.022971f
C3305 VDDA.n347 GNDA 0.033295f
C3306 VDDA.n348 GNDA 0.022971f
C3307 VDDA.n349 GNDA 0.014704f
C3308 VDDA.t329 GNDA 0.01321f
C3309 VDDA.n350 GNDA 0.040411f
C3310 VDDA.t328 GNDA 0.041564f
C3311 VDDA.t464 GNDA 0.0291f
C3312 VDDA.t100 GNDA 0.0291f
C3313 VDDA.t149 GNDA 0.0291f
C3314 VDDA.t120 GNDA 0.0291f
C3315 VDDA.t436 GNDA 0.0291f
C3316 VDDA.t462 GNDA 0.0291f
C3317 VDDA.t447 GNDA 0.0291f
C3318 VDDA.t109 GNDA 0.0291f
C3319 VDDA.t128 GNDA 0.0291f
C3320 VDDA.t445 GNDA 0.0291f
C3321 VDDA.t392 GNDA 0.041564f
C3322 VDDA.t393 GNDA 0.01321f
C3323 VDDA.n351 GNDA 0.040411f
C3324 VDDA.n352 GNDA 0.014704f
C3325 VDDA.n353 GNDA 0.022971f
C3326 VDDA.n355 GNDA 0.033295f
C3327 VDDA.n357 GNDA 0.033295f
C3328 VDDA.n358 GNDA 0.011338f
C3329 VDDA.n360 GNDA 0.064168f
C3330 VDDA.n361 GNDA 0.053038f
C3331 VDDA.n362 GNDA 0.012755f
C3332 VDDA.n363 GNDA 0.012755f
C3333 VDDA.n364 GNDA 0.012755f
C3334 VDDA.n365 GNDA 0.013227f
C3335 VDDA.n366 GNDA 0.013227f
C3336 VDDA.n367 GNDA 0.013227f
C3337 VDDA.n368 GNDA 0.013227f
C3338 VDDA.n369 GNDA 0.013227f
C3339 VDDA.n370 GNDA 0.012755f
C3340 VDDA.t97 GNDA 0.013227f
C3341 VDDA.t16 GNDA 0.013227f
C3342 VDDA.n371 GNDA 0.028089f
C3343 VDDA.t454 GNDA 0.013227f
C3344 VDDA.t154 GNDA 0.013227f
C3345 VDDA.n372 GNDA 0.033575f
C3346 VDDA.n373 GNDA 0.093785f
C3347 VDDA.t394 GNDA 0.023194f
C3348 VDDA.t326 GNDA 0.047051f
C3349 VDDA.t467 GNDA 0.013227f
C3350 VDDA.t86 GNDA 0.013227f
C3351 VDDA.n374 GNDA 0.033575f
C3352 VDDA.n375 GNDA 0.104754f
C3353 VDDA.t324 GNDA 0.023194f
C3354 VDDA.n376 GNDA 0.068916f
C3355 VDDA.n377 GNDA 0.136492f
C3356 VDDA.t325 GNDA 0.112748f
C3357 VDDA.t466 GNDA 0.088434f
C3358 VDDA.t85 GNDA 0.088434f
C3359 VDDA.t453 GNDA 0.088434f
C3360 VDDA.t153 GNDA 0.088434f
C3361 VDDA.t96 GNDA 0.088434f
C3362 VDDA.t15 GNDA 0.088434f
C3363 VDDA.t451 GNDA 0.088434f
C3364 VDDA.t124 GNDA 0.088434f
C3365 VDDA.t130 GNDA 0.088434f
C3366 VDDA.t67 GNDA 0.088434f
C3367 VDDA.t395 GNDA 0.114222f
C3368 VDDA.t396 GNDA 0.047051f
C3369 VDDA.n378 GNDA 0.142388f
C3370 VDDA.n379 GNDA 0.068916f
C3371 VDDA.t131 GNDA 0.013227f
C3372 VDDA.t68 GNDA 0.013227f
C3373 VDDA.n380 GNDA 0.033575f
C3374 VDDA.n381 GNDA 0.104754f
C3375 VDDA.t452 GNDA 0.013227f
C3376 VDDA.t125 GNDA 0.013227f
C3377 VDDA.n382 GNDA 0.033575f
C3378 VDDA.n383 GNDA 0.093785f
C3379 VDDA.n384 GNDA 0.012094f
C3380 VDDA.n385 GNDA 0.104165f
C3381 VDDA.t440 GNDA 0.011338f
C3382 VDDA.t259 GNDA 0.011338f
C3383 VDDA.n386 GNDA 0.038852f
C3384 VDDA.t189 GNDA 0.011338f
C3385 VDDA.t176 GNDA 0.011338f
C3386 VDDA.n387 GNDA 0.037525f
C3387 VDDA.n388 GNDA 0.143952f
C3388 VDDA.t181 GNDA 0.011338f
C3389 VDDA.t172 GNDA 0.011338f
C3390 VDDA.n389 GNDA 0.037525f
C3391 VDDA.n390 GNDA 0.073963f
C3392 VDDA.t242 GNDA 0.011338f
C3393 VDDA.t255 GNDA 0.011338f
C3394 VDDA.n391 GNDA 0.037525f
C3395 VDDA.n392 GNDA 0.073963f
C3396 VDDA.t241 GNDA 0.011338f
C3397 VDDA.t165 GNDA 0.011338f
C3398 VDDA.n393 GNDA 0.037525f
C3399 VDDA.n394 GNDA 0.073963f
C3400 VDDA.t188 GNDA 0.011338f
C3401 VDDA.t44 GNDA 0.011338f
C3402 VDDA.n395 GNDA 0.037525f
C3403 VDDA.n396 GNDA 0.108358f
C3404 VDDA.t318 GNDA 0.01104f
C3405 VDDA.n397 GNDA 0.057724f
C3406 VDDA.t320 GNDA 0.026966f
C3407 VDDA.n398 GNDA 0.082842f
C3408 VDDA.t319 GNDA 0.06718f
C3409 VDDA.t177 GNDA 0.049886f
C3410 VDDA.t158 GNDA 0.049886f
C3411 VDDA.t258 GNDA 0.049886f
C3412 VDDA.t215 GNDA 0.049886f
C3413 VDDA.t175 GNDA 0.049886f
C3414 VDDA.t180 GNDA 0.049886f
C3415 VDDA.t174 GNDA 0.049886f
C3416 VDDA.t190 GNDA 0.049886f
C3417 VDDA.t173 GNDA 0.049886f
C3418 VDDA.t260 GNDA 0.049886f
C3419 VDDA.t337 GNDA 0.06718f
C3420 VDDA.t338 GNDA 0.026966f
C3421 VDDA.n399 GNDA 0.082842f
C3422 VDDA.t336 GNDA 0.01104f
C3423 VDDA.n400 GNDA 0.044086f
C3424 VDDA.n401 GNDA 0.058814f
C3425 VDDA.n402 GNDA 0.070259f
C3426 VDDA.n403 GNDA 0.047522f
C3427 VDDA.n404 GNDA 0.021466f
C3428 VDDA.t407 GNDA 0.028297f
C3429 VDDA.t426 GNDA 0.018707f
C3430 VDDA.t43 GNDA 0.018707f
C3431 VDDA.t455 GNDA 0.018707f
C3432 VDDA.t19 GNDA 0.018707f
C3433 VDDA.t431 GNDA 0.018707f
C3434 VDDA.t92 GNDA 0.018707f
C3435 VDDA.t91 GNDA 0.018707f
C3436 VDDA.t24 GNDA 0.018707f
C3437 VDDA.t18 GNDA 0.018707f
C3438 VDDA.t104 GNDA 0.018707f
C3439 VDDA.t416 GNDA 0.028297f
C3440 VDDA.n405 GNDA 0.021466f
C3441 VDDA.n406 GNDA 0.033929f
C3442 VDDA.n407 GNDA 0.067623f
C3443 VDDA.n408 GNDA 0.040374f
C3444 VDDA.t160 GNDA 0.022675f
C3445 VDDA.t179 GNDA 0.022675f
C3446 VDDA.n409 GNDA 0.067557f
C3447 VDDA.n410 GNDA 0.1386f
C3448 VDDA.t411 GNDA 0.0798f
C3449 VDDA.t162 GNDA 0.022675f
C3450 VDDA.t208 GNDA 0.022675f
C3451 VDDA.n411 GNDA 0.067557f
C3452 VDDA.n412 GNDA 0.1386f
C3453 VDDA.t257 GNDA 0.022675f
C3454 VDDA.t210 GNDA 0.022675f
C3455 VDDA.n413 GNDA 0.067557f
C3456 VDDA.n414 GNDA 0.1386f
C3457 VDDA.t164 GNDA 0.022675f
C3458 VDDA.t187 GNDA 0.022675f
C3459 VDDA.n415 GNDA 0.067557f
C3460 VDDA.n416 GNDA 0.1386f
C3461 VDDA.t171 GNDA 0.022675f
C3462 VDDA.t262 GNDA 0.022675f
C3463 VDDA.n417 GNDA 0.067557f
C3464 VDDA.n418 GNDA 0.146729f
C3465 VDDA.t409 GNDA 0.027511f
C3466 VDDA.n419 GNDA 0.062825f
C3467 VDDA.n420 GNDA 0.266939f
C3468 VDDA.t410 GNDA 0.172889f
C3469 VDDA.t170 GNDA 0.133029f
C3470 VDDA.t261 GNDA 0.133029f
C3471 VDDA.t163 GNDA 0.133029f
C3472 VDDA.t186 GNDA 0.133029f
C3473 VDDA.t256 GNDA 0.133029f
C3474 VDDA.t209 GNDA 0.133029f
C3475 VDDA.t161 GNDA 0.133029f
C3476 VDDA.t207 GNDA 0.133029f
C3477 VDDA.t159 GNDA 0.133029f
C3478 VDDA.t178 GNDA 0.133029f
C3479 VDDA.t422 GNDA 0.172889f
C3480 VDDA.t423 GNDA 0.0798f
C3481 VDDA.n421 GNDA 0.266939f
C3482 VDDA.t421 GNDA 0.027511f
C3483 VDDA.n422 GNDA 0.061862f
C3484 VDDA.n423 GNDA 0.013059f
C3485 VDDA.n425 GNDA 0.036948f
C3486 VDDA.n427 GNDA 0.036948f
C3487 VDDA.n429 GNDA 0.036948f
C3488 VDDA.n431 GNDA 0.036948f
C3489 VDDA.n433 GNDA 0.036948f
C3490 VDDA.n435 GNDA 0.036948f
C3491 VDDA.n437 GNDA 0.036948f
C3492 VDDA.n439 GNDA 0.036948f
C3493 VDDA.n441 GNDA 0.036948f
C3494 VDDA.n443 GNDA 0.045893f
C3495 VDDA.n444 GNDA 0.03556f
C3496 VDDA.n445 GNDA 0.021317f
C3497 VDDA.t356 GNDA 0.028297f
C3498 VDDA.t211 GNDA 0.018707f
C3499 VDDA.t197 GNDA 0.018707f
C3500 VDDA.t184 GNDA 0.018707f
C3501 VDDA.t199 GNDA 0.018707f
C3502 VDDA.t203 GNDA 0.018707f
C3503 VDDA.t265 GNDA 0.018707f
C3504 VDDA.t77 GNDA 0.018707f
C3505 VDDA.t263 GNDA 0.018707f
C3506 VDDA.t201 GNDA 0.018707f
C3507 VDDA.t205 GNDA 0.018707f
C3508 VDDA.t213 GNDA 0.018707f
C3509 VDDA.t253 GNDA 0.018707f
C3510 VDDA.t193 GNDA 0.018707f
C3511 VDDA.t168 GNDA 0.018707f
C3512 VDDA.t191 GNDA 0.018707f
C3513 VDDA.t166 GNDA 0.018707f
C3514 VDDA.t195 GNDA 0.018707f
C3515 VDDA.t182 GNDA 0.018707f
C3516 VDDA.t251 GNDA 0.018707f
C3517 VDDA.t75 GNDA 0.018707f
C3518 VDDA.t362 GNDA 0.028297f
C3519 VDDA.n446 GNDA 0.021317f
C3520 VDDA.n447 GNDA 0.034562f
C3521 VDDA.n448 GNDA 0.028083f
C3522 VDDA.n449 GNDA 0.028155f
C3523 VDDA.n450 GNDA 0.074839f
C3524 VDDA.n451 GNDA 0.096757f
C3525 VDDA.t73 GNDA 0.013227f
C3526 VDDA.t88 GNDA 0.013227f
C3527 VDDA.n452 GNDA 0.028089f
C3528 VDDA.t123 GNDA 0.013227f
C3529 VDDA.t50 GNDA 0.013227f
C3530 VDDA.n453 GNDA 0.033575f
C3531 VDDA.n454 GNDA 0.093785f
C3532 VDDA.t352 GNDA 0.023194f
C3533 VDDA.t399 GNDA 0.047051f
C3534 VDDA.t23 GNDA 0.013227f
C3535 VDDA.t459 GNDA 0.013227f
C3536 VDDA.n455 GNDA 0.033575f
C3537 VDDA.n456 GNDA 0.104754f
C3538 VDDA.t397 GNDA 0.023194f
C3539 VDDA.n457 GNDA 0.068916f
C3540 VDDA.n458 GNDA 0.136492f
C3541 VDDA.t398 GNDA 0.112748f
C3542 VDDA.t22 GNDA 0.088434f
C3543 VDDA.t458 GNDA 0.088434f
C3544 VDDA.t122 GNDA 0.088434f
C3545 VDDA.t49 GNDA 0.088434f
C3546 VDDA.t72 GNDA 0.088434f
C3547 VDDA.t87 GNDA 0.088434f
C3548 VDDA.t102 GNDA 0.088434f
C3549 VDDA.t155 GNDA 0.088434f
C3550 VDDA.t13 GNDA 0.088434f
C3551 VDDA.t89 GNDA 0.088434f
C3552 VDDA.t353 GNDA 0.112748f
C3553 VDDA.t354 GNDA 0.047051f
C3554 VDDA.n459 GNDA 0.136492f
C3555 VDDA.n460 GNDA 0.068916f
C3556 VDDA.t14 GNDA 0.013227f
C3557 VDDA.t90 GNDA 0.013227f
C3558 VDDA.n461 GNDA 0.033575f
C3559 VDDA.n462 GNDA 0.104754f
C3560 VDDA.t103 GNDA 0.013227f
C3561 VDDA.t156 GNDA 0.013227f
C3562 VDDA.n463 GNDA 0.033575f
C3563 VDDA.n464 GNDA 0.093785f
C3564 VDDA.n465 GNDA 0.012094f
C3565 VDDA.n466 GNDA 0.104165f
C3566 VDDA.t277 GNDA 0.011338f
C3567 VDDA.t441 GNDA 0.011338f
C3568 VDDA.n467 GNDA 0.038852f
C3569 VDDA.t290 GNDA 0.011338f
C3570 VDDA.t289 GNDA 0.011338f
C3571 VDDA.n468 GNDA 0.037525f
C3572 VDDA.n469 GNDA 0.143952f
C3573 VDDA.t294 GNDA 0.011338f
C3574 VDDA.t273 GNDA 0.011338f
C3575 VDDA.n470 GNDA 0.037525f
C3576 VDDA.n471 GNDA 0.073963f
C3577 VDDA.t298 GNDA 0.011338f
C3578 VDDA.t278 GNDA 0.011338f
C3579 VDDA.n472 GNDA 0.037525f
C3580 VDDA.n473 GNDA 0.073963f
C3581 VDDA.t286 GNDA 0.011338f
C3582 VDDA.t305 GNDA 0.011338f
C3583 VDDA.n474 GNDA 0.037525f
C3584 VDDA.n475 GNDA 0.073963f
C3585 VDDA.t40 GNDA 0.011338f
C3586 VDDA.t269 GNDA 0.011338f
C3587 VDDA.n476 GNDA 0.037525f
C3588 VDDA.n477 GNDA 0.108358f
C3589 VDDA.t403 GNDA 0.01104f
C3590 VDDA.n478 GNDA 0.057724f
C3591 VDDA.t405 GNDA 0.026966f
C3592 VDDA.n479 GNDA 0.082842f
C3593 VDDA.t404 GNDA 0.06718f
C3594 VDDA.t283 GNDA 0.049886f
C3595 VDDA.t306 GNDA 0.049886f
C3596 VDDA.t297 GNDA 0.049886f
C3597 VDDA.t279 GNDA 0.049886f
C3598 VDDA.t299 GNDA 0.049886f
C3599 VDDA.t280 GNDA 0.049886f
C3600 VDDA.t302 GNDA 0.049886f
C3601 VDDA.t272 GNDA 0.049886f
C3602 VDDA.t293 GNDA 0.049886f
C3603 VDDA.t276 GNDA 0.049886f
C3604 VDDA.t383 GNDA 0.06718f
C3605 VDDA.t384 GNDA 0.026966f
C3606 VDDA.n480 GNDA 0.082842f
C3607 VDDA.t382 GNDA 0.01104f
C3608 VDDA.n481 GNDA 0.044086f
C3609 VDDA.n482 GNDA 0.058814f
C3610 VDDA.n483 GNDA 0.070259f
C3611 VDDA.n484 GNDA 0.047522f
C3612 VDDA.n485 GNDA 0.021466f
C3613 VDDA.t413 GNDA 0.028297f
C3614 VDDA.t468 GNDA 0.018707f
C3615 VDDA.t74 GNDA 0.018707f
C3616 VDDA.t442 GNDA 0.018707f
C3617 VDDA.t140 GNDA 0.018707f
C3618 VDDA.t240 GNDA 0.018707f
C3619 VDDA.t69 GNDA 0.018707f
C3620 VDDA.t17 GNDA 0.018707f
C3621 VDDA.t4 GNDA 0.018707f
C3622 VDDA.t248 GNDA 0.018707f
C3623 VDDA.t111 GNDA 0.018707f
C3624 VDDA.t310 GNDA 0.028297f
C3625 VDDA.n486 GNDA 0.021466f
C3626 VDDA.n487 GNDA 0.033929f
C3627 VDDA.n488 GNDA 0.06735f
C3628 VDDA.n489 GNDA 0.040268f
C3629 VDDA.t304 GNDA 0.022675f
C3630 VDDA.t282 GNDA 0.022675f
C3631 VDDA.n490 GNDA 0.067557f
C3632 VDDA.n491 GNDA 0.1386f
C3633 VDDA.t372 GNDA 0.0798f
C3634 VDDA.t301 GNDA 0.022675f
C3635 VDDA.t292 GNDA 0.022675f
C3636 VDDA.n492 GNDA 0.067557f
C3637 VDDA.n493 GNDA 0.1386f
C3638 VDDA.t271 GNDA 0.022675f
C3639 VDDA.t288 GNDA 0.022675f
C3640 VDDA.n494 GNDA 0.067557f
C3641 VDDA.n495 GNDA 0.1386f
C3642 VDDA.t308 GNDA 0.022675f
C3643 VDDA.t285 GNDA 0.022675f
C3644 VDDA.n496 GNDA 0.067557f
C3645 VDDA.n497 GNDA 0.1386f
C3646 VDDA.t296 GNDA 0.022675f
C3647 VDDA.t275 GNDA 0.022675f
C3648 VDDA.n498 GNDA 0.067557f
C3649 VDDA.n499 GNDA 0.146729f
C3650 VDDA.t370 GNDA 0.027511f
C3651 VDDA.n500 GNDA 0.062825f
C3652 VDDA.n501 GNDA 0.266939f
C3653 VDDA.t371 GNDA 0.172889f
C3654 VDDA.t274 GNDA 0.133029f
C3655 VDDA.t295 GNDA 0.133029f
C3656 VDDA.t284 GNDA 0.133029f
C3657 VDDA.t307 GNDA 0.133029f
C3658 VDDA.t287 GNDA 0.133029f
C3659 VDDA.t270 GNDA 0.133029f
C3660 VDDA.t291 GNDA 0.133029f
C3661 VDDA.t300 GNDA 0.133029f
C3662 VDDA.t281 GNDA 0.133029f
C3663 VDDA.t303 GNDA 0.133029f
C3664 VDDA.t359 GNDA 0.172889f
C3665 VDDA.t360 GNDA 0.0798f
C3666 VDDA.n502 GNDA 0.266939f
C3667 VDDA.t358 GNDA 0.027511f
C3668 VDDA.n503 GNDA 0.061862f
C3669 VDDA.n504 GNDA 0.021593f
C3670 VDDA.n505 GNDA 0.07632f
C3671 VDDA.n506 GNDA 0.096568f
C3672 VDDA.n507 GNDA 0.094409f
C3673 VDDA.n508 GNDA 0.015387f
C3674 VDDA.n509 GNDA 0.061352f
C3675 VDDA.t330 GNDA 0.014217f
C3676 VDDA.t348 GNDA 0.024554f
C3677 VDDA.t345 GNDA 0.014217f
C3678 VDDA.n510 GNDA 0.037638f
C3679 VDDA.n511 GNDA 0.073928f
C3680 VDDA.t346 GNDA 0.065816f
C3681 VDDA.t2 GNDA 0.049886f
C3682 VDDA.t331 GNDA 0.065816f
C3683 VDDA.t332 GNDA 0.024554f
C3684 VDDA.n512 GNDA 0.073928f
C3685 VDDA.n513 GNDA 0.03728f
C3686 VDDA.n514 GNDA 0.021572f
C3687 VDDA.n515 GNDA 0.0384f
C3688 VDDA.n516 GNDA 0.094908f
C3689 VDDA.t376 GNDA 0.023424f
C3690 VDDA.t230 GNDA 0.013227f
C3691 VDDA.n517 GNDA 0.033228f
C3692 VDDA.t341 GNDA 0.060279f
C3693 VDDA.t339 GNDA 0.023424f
C3694 VDDA.n518 GNDA 0.049476f
C3695 VDDA.n519 GNDA 0.150495f
C3696 VDDA.t340 GNDA 0.112748f
C3697 VDDA.t229 GNDA 0.088434f
C3698 VDDA.t377 GNDA 0.112748f
C3699 VDDA.t378 GNDA 0.047051f
C3700 VDDA.n520 GNDA 0.150495f
C3701 VDDA.n521 GNDA 0.049118f
C3702 VDDA.n522 GNDA 0.021572f
C3703 VDDA.n523 GNDA 0.07035f
C3704 VDDA.n524 GNDA 0.069545f
C3705 VDDA.n525 GNDA 0.01181f
C3706 VDDA.n526 GNDA 0.01181f
C3707 VDDA.n527 GNDA 2.31289f
C3708 VDDA.n528 GNDA 0.014172f
C3709 VDDA.n531 GNDA 0.015306f
C3710 VDDA.n532 GNDA 0.015306f
C3711 VDDA.n533 GNDA 0.015873f
C3712 VDDA.n534 GNDA 0.014172f
C3713 VDDA.n535 GNDA 0.014913f
C3714 VDDA.t366 GNDA 0.013237f
C3715 VDDA.t369 GNDA 0.013237f
C3716 VDDA.n536 GNDA 0.06585f
C3717 VDDA.t368 GNDA 0.045858f
C3718 VDDA.t9 GNDA 0.0291f
C3719 VDDA.t151 GNDA 0.0291f
C3720 VDDA.t365 GNDA 0.045858f
C3721 VDDA.n537 GNDA 0.06585f
C3722 VDDA.n538 GNDA 0.014913f
C3723 VDDA.n539 GNDA 0.035872f
C3724 VDDA.n541 GNDA 0.02452f
C3725 VDDA.t33 GNDA 0.011338f
C3726 VDDA.t55 GNDA 0.011338f
C3727 VDDA.n542 GNDA 0.037456f
C3728 VDDA.n543 GNDA 0.048332f
C3729 VDDA.n550 GNDA 0.013148f
C3730 VDDA.n554 GNDA 0.013227f
C3731 VDDA.t349 GNDA 0.054063f
C3732 VDDA.n555 GNDA 0.018565f
C3733 VDDA.t317 GNDA 0.015089f
C3734 VDDA.t387 GNDA 0.013237f
C3735 VDDA.n556 GNDA 0.066223f
C3736 VDDA.t386 GNDA 0.045858f
C3737 VDDA.t247 GNDA 0.0291f
C3738 VDDA.t157 GNDA 0.0291f
C3739 VDDA.t316 GNDA 0.046868f
C3740 VDDA.n557 GNDA 0.069357f
C3741 VDDA.n558 GNDA 0.018424f
C3742 VDDA.n559 GNDA 0.055422f
C3743 VDDA.t224 GNDA 0.011338f
C3744 VDDA.t232 GNDA 0.011338f
C3745 VDDA.n560 GNDA 0.037456f
C3746 VDDA.n561 GNDA 0.048332f
C3747 VDDA.t139 GNDA 0.011338f
C3748 VDDA.t145 GNDA 0.011338f
C3749 VDDA.n562 GNDA 0.037456f
C3750 VDDA.n563 GNDA 0.048332f
C3751 VDDA.t234 GNDA 0.011338f
C3752 VDDA.t35 GNDA 0.011338f
C3753 VDDA.n564 GNDA 0.037456f
C3754 VDDA.n565 GNDA 0.048332f
C3755 VDDA.t143 GNDA 0.011338f
C3756 VDDA.t239 GNDA 0.011338f
C3757 VDDA.n566 GNDA 0.037456f
C3758 VDDA.n567 GNDA 0.048332f
C3759 VDDA.t94 GNDA 0.011338f
C3760 VDDA.t217 GNDA 0.011338f
C3761 VDDA.n568 GNDA 0.037456f
C3762 VDDA.n569 GNDA 0.048332f
C3763 VDDA.t137 GNDA 0.011338f
C3764 VDDA.t222 GNDA 0.011338f
C3765 VDDA.n570 GNDA 0.037456f
C3766 VDDA.n571 GNDA 0.048332f
C3767 VDDA.t28 GNDA 0.011338f
C3768 VDDA.t60 GNDA 0.011338f
C3769 VDDA.n572 GNDA 0.037456f
C3770 VDDA.n573 GNDA 0.048332f
C3771 VDDA.n574 GNDA 0.025806f
C3772 VDDA.n575 GNDA 0.020191f
C3773 VDDA.n576 GNDA 0.01499f
C3774 VDDA.n578 GNDA 0.013148f
C3775 VDDA.n579 GNDA 0.013227f
C3776 VDDA.n580 GNDA 0.013227f
C3777 VDDA.n581 GNDA 0.013227f
C3778 VDDA.n582 GNDA 0.019146f
C3779 VDDA.n584 GNDA 0.106007f
C3780 VDDA.t350 GNDA 0.112432f
C3781 VDDA.t27 GNDA 0.115644f
C3782 VDDA.t59 GNDA 0.115644f
C3783 VDDA.t136 GNDA 0.115644f
C3784 VDDA.t221 GNDA 0.115644f
C3785 VDDA.t93 GNDA 0.115644f
C3786 VDDA.t216 GNDA 0.115644f
C3787 VDDA.t142 GNDA 0.115644f
C3788 VDDA.t238 GNDA 0.115644f
C3789 VDDA.t233 GNDA 0.115644f
C3790 VDDA.t34 GNDA 0.115644f
C3791 VDDA.t138 GNDA 0.115644f
C3792 VDDA.t144 GNDA 0.115644f
C3793 VDDA.t223 GNDA 0.115644f
C3794 VDDA.t231 GNDA 0.115644f
C3795 VDDA.t32 GNDA 0.115644f
C3796 VDDA.t54 GNDA 0.115644f
C3797 VDDA.t313 GNDA 0.112432f
C3798 VDDA.n588 GNDA 0.013227f
C3799 VDDA.n589 GNDA 0.013148f
C3800 VDDA.n590 GNDA 0.013227f
C3801 VDDA.n592 GNDA 0.013227f
C3802 VDDA.n593 GNDA 0.013227f
C3803 VDDA.n594 GNDA 0.013148f
C3804 VDDA.n595 GNDA 0.020888f
C3805 VDDA.n597 GNDA 0.106007f
C3806 VDDA.n599 GNDA 0.01499f
C3807 VDDA.t312 GNDA 0.054063f
C3808 VDDA.n600 GNDA 0.020191f
C3809 VDDA.n601 GNDA 0.042893f
C3810 VDDA.n602 GNDA 0.092357f
C3811 VDDA.n603 GNDA 0.090855f
C3812 VDDA.n604 GNDA 0.015306f
C3813 VDDA.n605 GNDA 0.015306f
C3814 VDDA.n606 GNDA 0.015306f
C3815 VDDA.n607 GNDA 0.015873f
C3816 VDDA.n608 GNDA 0.015873f
C3817 VDDA.n609 GNDA 0.015873f
C3818 VDDA.n610 GNDA 0.015873f
C3819 VDDA.n611 GNDA 0.043168f
C3820 VDDA.n612 GNDA 0.016069f
C3821 VDDA.n613 GNDA 0.014458f
C3822 VDDA.n614 GNDA 1.57594f
C3823 VDDA.n615 GNDA 0.014172f
C3824 VDDA.n618 GNDA 0.015306f
C3825 VDDA.n619 GNDA 0.015306f
C3826 VDDA.n620 GNDA 0.015873f
C3827 VDDA.n621 GNDA 0.014172f
C3828 VDDA.t53 GNDA 0.211259f
C3829 VDDA.t146 GNDA 0.212024f
C3830 VDDA.t57 GNDA 0.200687f
C3831 VDDA.t427 GNDA 0.211259f
C3832 VDDA.t29 GNDA 0.212024f
C3833 VDDA.t36 GNDA 0.200687f
C3834 VDDA.t133 GNDA 0.211259f
C3835 VDDA.t434 GNDA 0.212024f
C3836 VDDA.t141 GNDA 0.200687f
C3837 VDDA.t428 GNDA 0.211259f
C3838 VDDA.t95 GNDA 0.212024f
C3839 VDDA.t37 GNDA 0.200687f
C3840 VDDA.t56 GNDA 0.211259f
C3841 VDDA.t435 GNDA 0.212024f
C3842 VDDA.t430 GNDA 0.200687f
C3843 VDDA.n622 GNDA 0.141607f
C3844 VDDA.t132 GNDA 0.112769f
C3845 VDDA.n623 GNDA 0.153647f
C3846 VDDA.t429 GNDA 0.112769f
C3847 VDDA.n624 GNDA 0.153647f
C3848 VDDA.t58 GNDA 0.112769f
C3849 VDDA.n625 GNDA 0.153647f
C3850 VDDA.t218 GNDA 0.112769f
C3851 VDDA.n626 GNDA 0.153647f
C3852 VDDA.t237 GNDA 0.468095f
C3853 VDDA.n627 GNDA 0.762326f
C3854 VDDA.n628 GNDA 0.015306f
C3855 VDDA.n629 GNDA 0.015306f
C3856 VDDA.n630 GNDA 0.015306f
C3857 VDDA.n631 GNDA 0.015873f
C3858 VDDA.n632 GNDA 0.015873f
C3859 VDDA.n633 GNDA 0.015873f
C3860 VDDA.n634 GNDA 0.015873f
C3861 VDDA.n635 GNDA 0.043168f
C3862 VDDA.n636 GNDA 0.016069f
C3863 VDDA.n637 GNDA 0.014458f
C3864 VDDA.n638 GNDA 3.74899f
C3865 VDDA.n639 GNDA 0.287221f
C3866 VDDA.n640 GNDA 0.143611f
C3867 VDDA.n642 GNDA 0.287221f
C3868 VDDA.n645 GNDA 0.151169f
C3869 VDDA.n646 GNDA 0.14739f
C3870 VDDA.n647 GNDA 0.143611f
C3871 VDDA.n650 GNDA 0.151169f
C3872 VDDA.n651 GNDA 0.317455f
C3873 VDDA.n652 GNDA 3.17455f
C3874 VDDA.n653 GNDA 2.19951f
C3875 two_stage_opamp_dummy_magic_23_0.Y.t11 GNDA 0.037911f
C3876 two_stage_opamp_dummy_magic_23_0.Y.t5 GNDA 0.037911f
C3877 two_stage_opamp_dummy_magic_23_0.Y.n0 GNDA 0.082489f
C3878 two_stage_opamp_dummy_magic_23_0.Y.n1 GNDA 0.256901f
C3879 two_stage_opamp_dummy_magic_23_0.Y.n2 GNDA 0.080625f
C3880 two_stage_opamp_dummy_magic_23_0.Y.t4 GNDA 0.037911f
C3881 two_stage_opamp_dummy_magic_23_0.Y.t15 GNDA 0.037911f
C3882 two_stage_opamp_dummy_magic_23_0.Y.n3 GNDA 0.082489f
C3883 two_stage_opamp_dummy_magic_23_0.Y.n4 GNDA 0.327754f
C3884 two_stage_opamp_dummy_magic_23_0.Y.t24 GNDA 0.037911f
C3885 two_stage_opamp_dummy_magic_23_0.Y.t19 GNDA 0.037911f
C3886 two_stage_opamp_dummy_magic_23_0.Y.n5 GNDA 0.082489f
C3887 two_stage_opamp_dummy_magic_23_0.Y.n6 GNDA 0.327754f
C3888 two_stage_opamp_dummy_magic_23_0.Y.n7 GNDA 0.137048f
C3889 two_stage_opamp_dummy_magic_23_0.Y.t10 GNDA 0.037911f
C3890 two_stage_opamp_dummy_magic_23_0.Y.t8 GNDA 0.037911f
C3891 two_stage_opamp_dummy_magic_23_0.Y.n8 GNDA 0.082489f
C3892 two_stage_opamp_dummy_magic_23_0.Y.n9 GNDA 0.314545f
C3893 two_stage_opamp_dummy_magic_23_0.Y.n10 GNDA 0.144975f
C3894 two_stage_opamp_dummy_magic_23_0.Y.t9 GNDA 0.037911f
C3895 two_stage_opamp_dummy_magic_23_0.Y.t7 GNDA 0.037911f
C3896 two_stage_opamp_dummy_magic_23_0.Y.n11 GNDA 0.082489f
C3897 two_stage_opamp_dummy_magic_23_0.Y.n12 GNDA 0.314545f
C3898 two_stage_opamp_dummy_magic_23_0.Y.n13 GNDA 0.084683f
C3899 two_stage_opamp_dummy_magic_23_0.Y.n14 GNDA 0.084683f
C3900 two_stage_opamp_dummy_magic_23_0.Y.n15 GNDA 0.144975f
C3901 two_stage_opamp_dummy_magic_23_0.Y.t12 GNDA 0.037911f
C3902 two_stage_opamp_dummy_magic_23_0.Y.t6 GNDA 0.037911f
C3903 two_stage_opamp_dummy_magic_23_0.Y.n16 GNDA 0.082489f
C3904 two_stage_opamp_dummy_magic_23_0.Y.n17 GNDA 0.314545f
C3905 two_stage_opamp_dummy_magic_23_0.Y.n18 GNDA 0.137048f
C3906 two_stage_opamp_dummy_magic_23_0.Y.n19 GNDA 0.075821f
C3907 two_stage_opamp_dummy_magic_23_0.Y.n20 GNDA 0.3074f
C3908 two_stage_opamp_dummy_magic_23_0.Y.t1 GNDA 0.088458f
C3909 two_stage_opamp_dummy_magic_23_0.Y.t17 GNDA 0.088458f
C3910 two_stage_opamp_dummy_magic_23_0.Y.n21 GNDA 0.180951f
C3911 two_stage_opamp_dummy_magic_23_0.Y.n22 GNDA 0.492191f
C3912 two_stage_opamp_dummy_magic_23_0.Y.n23 GNDA 0.095948f
C3913 two_stage_opamp_dummy_magic_23_0.Y.n24 GNDA 0.163678f
C3914 two_stage_opamp_dummy_magic_23_0.Y.t3 GNDA 0.088458f
C3915 two_stage_opamp_dummy_magic_23_0.Y.t0 GNDA 0.088458f
C3916 two_stage_opamp_dummy_magic_23_0.Y.n25 GNDA 0.180951f
C3917 two_stage_opamp_dummy_magic_23_0.Y.n26 GNDA 0.585864f
C3918 two_stage_opamp_dummy_magic_23_0.Y.t13 GNDA 0.088458f
C3919 two_stage_opamp_dummy_magic_23_0.Y.t20 GNDA 0.088458f
C3920 two_stage_opamp_dummy_magic_23_0.Y.n27 GNDA 0.180951f
C3921 two_stage_opamp_dummy_magic_23_0.Y.n28 GNDA 0.569865f
C3922 two_stage_opamp_dummy_magic_23_0.Y.n29 GNDA 0.163678f
C3923 two_stage_opamp_dummy_magic_23_0.Y.n30 GNDA 0.095948f
C3924 two_stage_opamp_dummy_magic_23_0.Y.t22 GNDA 0.088458f
C3925 two_stage_opamp_dummy_magic_23_0.Y.t23 GNDA 0.088458f
C3926 two_stage_opamp_dummy_magic_23_0.Y.n31 GNDA 0.180951f
C3927 two_stage_opamp_dummy_magic_23_0.Y.n32 GNDA 0.569865f
C3928 two_stage_opamp_dummy_magic_23_0.Y.n33 GNDA 0.095948f
C3929 two_stage_opamp_dummy_magic_23_0.Y.t21 GNDA 0.088458f
C3930 two_stage_opamp_dummy_magic_23_0.Y.t14 GNDA 0.088458f
C3931 two_stage_opamp_dummy_magic_23_0.Y.n34 GNDA 0.180951f
C3932 two_stage_opamp_dummy_magic_23_0.Y.n35 GNDA 0.569865f
C3933 two_stage_opamp_dummy_magic_23_0.Y.n36 GNDA 0.095948f
C3934 two_stage_opamp_dummy_magic_23_0.Y.n37 GNDA 0.163678f
C3935 two_stage_opamp_dummy_magic_23_0.Y.t2 GNDA 0.088458f
C3936 two_stage_opamp_dummy_magic_23_0.Y.t18 GNDA 0.088458f
C3937 two_stage_opamp_dummy_magic_23_0.Y.n38 GNDA 0.180951f
C3938 two_stage_opamp_dummy_magic_23_0.Y.n39 GNDA 0.569865f
C3939 two_stage_opamp_dummy_magic_23_0.Y.n40 GNDA 0.149208f
C3940 two_stage_opamp_dummy_magic_23_0.Y.n41 GNDA 0.48498f
C3941 two_stage_opamp_dummy_magic_23_0.Y.t52 GNDA 0.053075f
C3942 two_stage_opamp_dummy_magic_23_0.Y.t29 GNDA 0.053075f
C3943 two_stage_opamp_dummy_magic_23_0.Y.t45 GNDA 0.053075f
C3944 two_stage_opamp_dummy_magic_23_0.Y.t31 GNDA 0.053075f
C3945 two_stage_opamp_dummy_magic_23_0.Y.t46 GNDA 0.053075f
C3946 two_stage_opamp_dummy_magic_23_0.Y.t34 GNDA 0.053075f
C3947 two_stage_opamp_dummy_magic_23_0.Y.t27 GNDA 0.053075f
C3948 two_stage_opamp_dummy_magic_23_0.Y.t43 GNDA 0.064448f
C3949 two_stage_opamp_dummy_magic_23_0.Y.n42 GNDA 0.064448f
C3950 two_stage_opamp_dummy_magic_23_0.Y.n43 GNDA 0.041702f
C3951 two_stage_opamp_dummy_magic_23_0.Y.n44 GNDA 0.041702f
C3952 two_stage_opamp_dummy_magic_23_0.Y.n45 GNDA 0.041702f
C3953 two_stage_opamp_dummy_magic_23_0.Y.n46 GNDA 0.041702f
C3954 two_stage_opamp_dummy_magic_23_0.Y.n47 GNDA 0.041702f
C3955 two_stage_opamp_dummy_magic_23_0.Y.n48 GNDA 0.033646f
C3956 two_stage_opamp_dummy_magic_23_0.Y.t37 GNDA 0.053075f
C3957 two_stage_opamp_dummy_magic_23_0.Y.t49 GNDA 0.064448f
C3958 two_stage_opamp_dummy_magic_23_0.Y.n49 GNDA 0.056392f
C3959 two_stage_opamp_dummy_magic_23_0.Y.n50 GNDA 0.021219f
C3960 two_stage_opamp_dummy_magic_23_0.Y.t26 GNDA 0.081508f
C3961 two_stage_opamp_dummy_magic_23_0.Y.t33 GNDA 0.081508f
C3962 two_stage_opamp_dummy_magic_23_0.Y.t48 GNDA 0.081508f
C3963 two_stage_opamp_dummy_magic_23_0.Y.t36 GNDA 0.081508f
C3964 two_stage_opamp_dummy_magic_23_0.Y.t51 GNDA 0.081508f
C3965 two_stage_opamp_dummy_magic_23_0.Y.t39 GNDA 0.081508f
C3966 two_stage_opamp_dummy_magic_23_0.Y.t32 GNDA 0.081508f
C3967 two_stage_opamp_dummy_magic_23_0.Y.t47 GNDA 0.092661f
C3968 two_stage_opamp_dummy_magic_23_0.Y.n51 GNDA 0.083624f
C3969 two_stage_opamp_dummy_magic_23_0.Y.n52 GNDA 0.05118f
C3970 two_stage_opamp_dummy_magic_23_0.Y.n53 GNDA 0.05118f
C3971 two_stage_opamp_dummy_magic_23_0.Y.n54 GNDA 0.05118f
C3972 two_stage_opamp_dummy_magic_23_0.Y.n55 GNDA 0.05118f
C3973 two_stage_opamp_dummy_magic_23_0.Y.n56 GNDA 0.05118f
C3974 two_stage_opamp_dummy_magic_23_0.Y.n57 GNDA 0.043123f
C3975 two_stage_opamp_dummy_magic_23_0.Y.t41 GNDA 0.081508f
C3976 two_stage_opamp_dummy_magic_23_0.Y.t54 GNDA 0.092661f
C3977 two_stage_opamp_dummy_magic_23_0.Y.n58 GNDA 0.075568f
C3978 two_stage_opamp_dummy_magic_23_0.Y.n59 GNDA 0.021219f
C3979 two_stage_opamp_dummy_magic_23_0.Y.n60 GNDA 0.091639f
C3980 two_stage_opamp_dummy_magic_23_0.Y.n61 GNDA 1.04027f
C3981 two_stage_opamp_dummy_magic_23_0.Y.n62 GNDA 0.450882f
C3982 two_stage_opamp_dummy_magic_23_0.Y.t42 GNDA 0.166807f
C3983 two_stage_opamp_dummy_magic_23_0.Y.t35 GNDA 0.166807f
C3984 two_stage_opamp_dummy_magic_23_0.Y.t50 GNDA 0.177661f
C3985 two_stage_opamp_dummy_magic_23_0.Y.n63 GNDA 0.140789f
C3986 two_stage_opamp_dummy_magic_23_0.Y.n64 GNDA 0.071557f
C3987 two_stage_opamp_dummy_magic_23_0.Y.t25 GNDA 0.166807f
C3988 two_stage_opamp_dummy_magic_23_0.Y.t40 GNDA 0.166807f
C3989 two_stage_opamp_dummy_magic_23_0.Y.t53 GNDA 0.166807f
C3990 two_stage_opamp_dummy_magic_23_0.Y.t38 GNDA 0.166807f
C3991 two_stage_opamp_dummy_magic_23_0.Y.t30 GNDA 0.166807f
C3992 two_stage_opamp_dummy_magic_23_0.Y.t44 GNDA 0.166807f
C3993 two_stage_opamp_dummy_magic_23_0.Y.t28 GNDA 0.177661f
C3994 two_stage_opamp_dummy_magic_23_0.Y.n65 GNDA 0.140789f
C3995 two_stage_opamp_dummy_magic_23_0.Y.n66 GNDA 0.079613f
C3996 two_stage_opamp_dummy_magic_23_0.Y.n67 GNDA 0.079613f
C3997 two_stage_opamp_dummy_magic_23_0.Y.n68 GNDA 0.079613f
C3998 two_stage_opamp_dummy_magic_23_0.Y.n69 GNDA 0.079613f
C3999 two_stage_opamp_dummy_magic_23_0.Y.n70 GNDA 0.071557f
C4000 two_stage_opamp_dummy_magic_23_0.Y.n71 GNDA 0.036197f
C4001 two_stage_opamp_dummy_magic_23_0.Y.n72 GNDA 1.26467f
C4002 two_stage_opamp_dummy_magic_23_0.Y.t16 GNDA 1.21199f
.ends

