** sch_path: /foss/designs/projects/bandgapref/xschem_ngspice/new_files/tb_low_voltage_BGR_7.sch
**.subckt tb_low_voltage_BGR_7
V1 VDD GND 1.8
XM1 V1 Vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 V2 Vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vmeas V1 Vbiasn 0
.save i(vmeas)
Vmeas1 V2 Vreg 0
.save i(vmeas1)
XM5 net2 net2 GND GND sky130_fd_pr__nfet_01v8 L=5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 start_up Vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 start_up Vbiasp VDD sky130_fd_pr__pfet_01v8 L=0.6 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 Vbiasn Vbiasn GND GND sky130_fd_pr__nfet_01v8 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 Vreg Vreg net3 GND sky130_fd_pr__nfet_01v8 L=0.6 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vmeas2 net1 V1 0
.save i(vmeas2)
Vmeas3 start_up net2 0
.save i(vmeas3)
XM9 net4 Vreg GND GND sky130_fd_pr__nfet_01v8 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 Vbiasp Vbiasn GND GND sky130_fd_pr__nfet_01v8 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 net4 net4 VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 Vbiasp net4 VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR7 GND net3 GND sky130_fd_pr__res_xhigh_po_0p35 L=0.90 mult=1 m=1
**** begin user architecture code
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt



.option method=gear
.option wnflag=1
.option savecurrents
* .temp =140

.save
+@m.xm1.msky130_fd_pr__pfet_01v8[gm]
+@m.xm1.msky130_fd_pr__pfet_01v8[vth]
+@m.xm1.msky130_fd_pr__pfet_01v8[vgs]
+@m.xm1.msky130_fd_pr__pfet_01v8[vds]
+@m.xm2.msky130_fd_pr__pfet_01v8[gm]
+@m.xm2.msky130_fd_pr__pfet_01v8[vth]
+@m.xm2.msky130_fd_pr__pfet_01v8[vgs]
+@m.xm2.msky130_fd_pr__pfet_01v8[vds]
+@m.xm3.msky130_fd_pr__pfet_01v8[gm]
+@m.xm4.msky130_fd_pr__pfet_01v8[gm]
+@m.xm4.msky130_fd_pr__nfet_01v8[gm]
+@m.x1.xm1.msky130_fd_pr__nfet_01v8[gm]
+@m.x1.xm2.msky130_fd_pr__nfet_01v8[gm]
+@m.x1.xm3.msky130_fd_pr__nfet_01v8[gm]
+@m.x1.xm4.msky130_fd_pr__pfet_01v8[gm]
+@m.x1.xm5.msky130_fd_pr__pfet_01v8[gm]
+@m.x1.xm6.msky130_fd_pr__nfet_01v8[gm]
+@m.x1.xm7.msky130_fd_pr__pfet_01v8[gm]
+@m.x2.xm1.msky130_fd_pr__nfet_01v8[gm]
+@m.x2.xm2.msky130_fd_pr__nfet_01v8[gm]
+@m.x2.xm3.msky130_fd_pr__nfet_01v8[gm]
+@m.x2.xm4.msky130_fd_pr__pfet_01v8[gm]
+@m.x2.xm5.msky130_fd_pr__pfet_01v8[gm]
+@m.x2.xm6.msky130_fd_pr__pfet_01v8[gm]
+@m.x2.xm7.msky130_fd_pr__pfet_01v8[gm]

* .ic v(vin-) = 0.8
* .ic v(vin+) = 0.8
* .ic v(v_top) = 1.8

.control

  * let start_vdd = 0.3
  * let stop_vdd = 1.8
  * let delta_vdd = 0.3
  * let w_act = start_vdd
  * while w_act le stop_vdd
    * echo $&w_act
    * alter V1 = w_act
    * echo v[vdd]
    * alter @V1[pwl] = [ 0 0 1us 0 2us $&w_act ]
    * reset
    save all
    * run
    * dc temp -40 120 5 V1 1.6 2.0 0.05
    * dc V1 1.7 1.9 0.001 temp -40 120 40
    * dc V1 0 2.0 0.01 temp -40 120 40
    dc V1 0 2.0 0.01
    * tran 1ns 8us
    remzerovec
    write tb_low_voltage_BGR_7.raw
    * let w_act = w_act + delta_vdd
    set appendwrite
  * end

.endc



**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
