magic
tech sky130A
timestamp 1739026514
<< nwell >>
rect 9230 2165 10840 2455
<< nmos >>
rect 9250 1805 9310 2005
rect 9360 1805 9420 2005
rect 9470 1805 9530 2005
rect 9580 1805 9640 2005
rect 9790 1805 9850 2005
rect 9900 1805 9960 2005
rect 10010 1805 10070 2005
rect 10120 1805 10180 2005
rect 10330 1805 10390 2005
rect 10440 1805 10500 2005
rect 10550 1805 10610 2005
rect 10660 1805 10720 2005
<< pmos >>
rect 9350 2235 9410 2435
rect 9460 2235 9520 2435
rect 9570 2235 9630 2435
rect 9680 2235 9740 2435
rect 9790 2235 9850 2435
rect 9900 2235 9960 2435
rect 10110 2235 10170 2435
rect 10220 2235 10280 2435
rect 10330 2235 10390 2435
rect 10440 2235 10500 2435
rect 10550 2235 10610 2435
rect 10660 2235 10720 2435
<< ndiff >>
rect 9200 1990 9250 2005
rect 9200 1820 9215 1990
rect 9235 1820 9250 1990
rect 9200 1805 9250 1820
rect 9310 1990 9360 2005
rect 9310 1820 9325 1990
rect 9345 1820 9360 1990
rect 9310 1805 9360 1820
rect 9420 1990 9470 2005
rect 9420 1820 9435 1990
rect 9455 1820 9470 1990
rect 9420 1805 9470 1820
rect 9530 1990 9580 2005
rect 9530 1820 9545 1990
rect 9565 1820 9580 1990
rect 9530 1805 9580 1820
rect 9640 1990 9690 2005
rect 9740 1990 9790 2005
rect 9640 1820 9655 1990
rect 9675 1820 9690 1990
rect 9740 1820 9755 1990
rect 9775 1820 9790 1990
rect 9640 1805 9690 1820
rect 9740 1805 9790 1820
rect 9850 1990 9900 2005
rect 9850 1820 9865 1990
rect 9885 1820 9900 1990
rect 9850 1805 9900 1820
rect 9960 1990 10010 2005
rect 9960 1820 9975 1990
rect 9995 1820 10010 1990
rect 9960 1805 10010 1820
rect 10070 1990 10120 2005
rect 10070 1820 10085 1990
rect 10105 1820 10120 1990
rect 10070 1805 10120 1820
rect 10180 1990 10230 2005
rect 10280 1990 10330 2005
rect 10180 1820 10195 1990
rect 10215 1820 10230 1990
rect 10280 1820 10295 1990
rect 10315 1820 10330 1990
rect 10180 1805 10230 1820
rect 10280 1805 10330 1820
rect 10390 1990 10440 2005
rect 10390 1820 10405 1990
rect 10425 1820 10440 1990
rect 10390 1805 10440 1820
rect 10500 1990 10550 2005
rect 10500 1820 10515 1990
rect 10535 1820 10550 1990
rect 10500 1805 10550 1820
rect 10610 1990 10660 2005
rect 10610 1820 10625 1990
rect 10645 1820 10660 1990
rect 10610 1805 10660 1820
rect 10720 1990 10770 2005
rect 10720 1820 10735 1990
rect 10755 1820 10770 1990
rect 10720 1805 10770 1820
<< pdiff >>
rect 9300 2420 9350 2435
rect 9300 2250 9315 2420
rect 9335 2250 9350 2420
rect 9300 2235 9350 2250
rect 9410 2420 9460 2435
rect 9410 2250 9425 2420
rect 9445 2250 9460 2420
rect 9410 2235 9460 2250
rect 9520 2420 9570 2435
rect 9520 2250 9535 2420
rect 9555 2250 9570 2420
rect 9520 2235 9570 2250
rect 9630 2420 9680 2435
rect 9630 2250 9645 2420
rect 9665 2250 9680 2420
rect 9630 2235 9680 2250
rect 9740 2420 9790 2435
rect 9740 2250 9755 2420
rect 9775 2250 9790 2420
rect 9740 2235 9790 2250
rect 9850 2420 9900 2435
rect 9850 2250 9865 2420
rect 9885 2250 9900 2420
rect 9850 2235 9900 2250
rect 9960 2420 10010 2435
rect 10060 2420 10110 2435
rect 9960 2250 9975 2420
rect 9995 2250 10010 2420
rect 10060 2250 10075 2420
rect 10095 2250 10110 2420
rect 9960 2235 10010 2250
rect 10060 2235 10110 2250
rect 10170 2420 10220 2435
rect 10170 2250 10185 2420
rect 10205 2250 10220 2420
rect 10170 2235 10220 2250
rect 10280 2420 10330 2435
rect 10280 2250 10295 2420
rect 10315 2250 10330 2420
rect 10280 2235 10330 2250
rect 10390 2420 10440 2435
rect 10390 2250 10405 2420
rect 10425 2250 10440 2420
rect 10390 2235 10440 2250
rect 10500 2420 10550 2435
rect 10500 2250 10515 2420
rect 10535 2250 10550 2420
rect 10500 2235 10550 2250
rect 10610 2420 10660 2435
rect 10610 2250 10625 2420
rect 10645 2250 10660 2420
rect 10610 2235 10660 2250
rect 10720 2420 10770 2435
rect 10720 2250 10735 2420
rect 10755 2250 10770 2420
rect 10720 2235 10770 2250
<< ndiffc >>
rect 9215 1820 9235 1990
rect 9325 1820 9345 1990
rect 9435 1820 9455 1990
rect 9545 1820 9565 1990
rect 9655 1820 9675 1990
rect 9755 1820 9775 1990
rect 9865 1820 9885 1990
rect 9975 1820 9995 1990
rect 10085 1820 10105 1990
rect 10195 1820 10215 1990
rect 10295 1820 10315 1990
rect 10405 1820 10425 1990
rect 10515 1820 10535 1990
rect 10625 1820 10645 1990
rect 10735 1820 10755 1990
<< pdiffc >>
rect 9315 2250 9335 2420
rect 9425 2250 9445 2420
rect 9535 2250 9555 2420
rect 9645 2250 9665 2420
rect 9755 2250 9775 2420
rect 9865 2250 9885 2420
rect 9975 2250 9995 2420
rect 10075 2250 10095 2420
rect 10185 2250 10205 2420
rect 10295 2250 10315 2420
rect 10405 2250 10425 2420
rect 10515 2250 10535 2420
rect 10625 2250 10645 2420
rect 10735 2250 10755 2420
<< psubdiff >>
rect 9150 1990 9200 2005
rect 9150 1820 9165 1990
rect 9185 1820 9200 1990
rect 9150 1805 9200 1820
rect 9690 1990 9740 2005
rect 9690 1820 9705 1990
rect 9725 1820 9740 1990
rect 9690 1805 9740 1820
rect 10230 1990 10280 2005
rect 10230 1820 10245 1990
rect 10265 1820 10280 1990
rect 10230 1805 10280 1820
rect 10770 1990 10820 2005
rect 10770 1820 10785 1990
rect 10805 1820 10820 1990
rect 10770 1805 10820 1820
<< nsubdiff >>
rect 9250 2420 9300 2435
rect 9250 2250 9265 2420
rect 9285 2250 9300 2420
rect 9250 2235 9300 2250
rect 10010 2420 10060 2435
rect 10010 2250 10025 2420
rect 10045 2250 10060 2420
rect 10010 2235 10060 2250
rect 10770 2420 10820 2435
rect 10770 2250 10785 2420
rect 10805 2250 10820 2420
rect 10770 2235 10820 2250
<< psubdiffcont >>
rect 9165 1820 9185 1990
rect 9705 1820 9725 1990
rect 10245 1820 10265 1990
rect 10785 1820 10805 1990
<< nsubdiffcont >>
rect 9265 2250 9285 2420
rect 10025 2250 10045 2420
rect 10785 2250 10805 2420
<< poly >>
rect 10555 2505 10610 2515
rect 10555 2470 10565 2505
rect 10600 2470 10610 2505
rect 10555 2460 10610 2470
rect 9350 2435 9410 2450
rect 9460 2435 9520 2450
rect 9570 2435 9630 2450
rect 9680 2435 9740 2450
rect 9790 2435 9850 2450
rect 9900 2435 9960 2450
rect 10110 2435 10170 2450
rect 10220 2445 10610 2460
rect 10220 2435 10280 2445
rect 10330 2435 10390 2445
rect 10440 2435 10500 2445
rect 10550 2435 10610 2445
rect 10660 2435 10720 2450
rect 9350 2225 9410 2235
rect 9305 2210 9410 2225
rect 9305 2190 9315 2210
rect 9335 2205 9410 2210
rect 9460 2225 9520 2235
rect 9570 2225 9630 2235
rect 9680 2225 9740 2235
rect 9790 2225 9850 2235
rect 9460 2205 9850 2225
rect 9900 2225 9960 2235
rect 10110 2225 10170 2235
rect 9900 2210 10170 2225
rect 10220 2220 10280 2235
rect 10330 2220 10390 2235
rect 10440 2220 10500 2235
rect 10550 2220 10610 2235
rect 10660 2225 10720 2235
rect 10660 2210 10765 2225
rect 9335 2190 9345 2205
rect 9305 2180 9345 2190
rect 10015 2190 10025 2210
rect 10045 2190 10055 2210
rect 10015 2180 10055 2190
rect 10725 2190 10735 2210
rect 10755 2190 10765 2210
rect 10725 2180 10765 2190
rect 9205 2050 9245 2060
rect 9205 2030 9215 2050
rect 9235 2030 9245 2050
rect 9370 2050 9410 2060
rect 9370 2030 9380 2050
rect 9400 2030 9410 2050
rect 9480 2050 9520 2060
rect 9480 2030 9490 2050
rect 9510 2030 9520 2050
rect 9695 2050 9735 2060
rect 9695 2030 9705 2050
rect 9725 2030 9735 2050
rect 10235 2050 10275 2060
rect 10235 2030 10245 2050
rect 10265 2030 10275 2050
rect 10725 2050 10765 2060
rect 10725 2030 10735 2050
rect 10755 2030 10765 2050
rect 9205 2015 9310 2030
rect 9250 2005 9310 2015
rect 9360 2015 9530 2030
rect 9360 2005 9420 2015
rect 9470 2005 9530 2015
rect 9580 2015 9850 2030
rect 9580 2005 9640 2015
rect 9790 2005 9850 2015
rect 9900 2015 10070 2030
rect 9900 2005 9960 2015
rect 10010 2005 10070 2015
rect 10120 2015 10390 2030
rect 10120 2005 10180 2015
rect 10330 2005 10390 2015
rect 10440 2005 10500 2020
rect 10550 2005 10610 2020
rect 10660 2015 10765 2030
rect 10660 2005 10720 2015
rect 9250 1790 9310 1805
rect 9360 1790 9420 1805
rect 9470 1765 9530 1805
rect 9580 1790 9640 1805
rect 9790 1790 9850 1805
rect 9900 1765 9960 1805
rect 10010 1790 10070 1805
rect 10120 1790 10180 1805
rect 10330 1790 10390 1805
rect 10440 1795 10500 1805
rect 10550 1795 10610 1805
rect 10440 1780 10610 1795
rect 10660 1790 10720 1805
rect 9470 1750 9960 1765
rect 10555 1770 10610 1780
rect 10555 1735 10565 1770
rect 10600 1735 10610 1770
rect 10555 1725 10610 1735
<< polycont >>
rect 10565 2470 10600 2505
rect 9315 2190 9335 2210
rect 10025 2190 10045 2210
rect 10735 2190 10755 2210
rect 9215 2030 9235 2050
rect 9380 2030 9400 2050
rect 9490 2030 9510 2050
rect 9705 2030 9725 2050
rect 10245 2030 10265 2050
rect 10735 2030 10755 2050
rect 10565 1735 10600 1770
<< locali >>
rect 8205 2885 10905 2895
rect 8205 2850 10860 2885
rect 10895 2850 10905 2885
rect 8205 2840 10905 2850
rect 10555 2505 10905 2515
rect 10555 2470 10565 2505
rect 10600 2470 10860 2505
rect 10895 2470 10905 2505
rect 10555 2460 10905 2470
rect 9255 2420 9345 2430
rect 9255 2250 9265 2420
rect 9285 2250 9315 2420
rect 9335 2250 9345 2420
rect 9255 2240 9345 2250
rect 9415 2420 9455 2430
rect 9415 2250 9425 2420
rect 9445 2250 9455 2420
rect 9415 2240 9455 2250
rect 9525 2420 9565 2430
rect 9525 2250 9535 2420
rect 9555 2250 9565 2420
rect 9305 2210 9345 2240
rect 9305 2190 9315 2210
rect 9335 2190 9345 2210
rect 9305 2180 9345 2190
rect 9525 2220 9565 2250
rect 9635 2420 9675 2430
rect 9635 2250 9645 2420
rect 9665 2250 9675 2420
rect 9635 2240 9675 2250
rect 9745 2420 9785 2430
rect 9745 2250 9755 2420
rect 9775 2250 9785 2420
rect 9745 2220 9785 2250
rect 9855 2420 9895 2430
rect 9855 2250 9865 2420
rect 9885 2250 9895 2420
rect 9855 2240 9895 2250
rect 9965 2420 10105 2430
rect 9965 2250 9975 2420
rect 9995 2250 10025 2420
rect 10045 2250 10075 2420
rect 10095 2250 10105 2420
rect 9965 2240 10105 2250
rect 10175 2420 10215 2430
rect 10175 2250 10185 2420
rect 10205 2250 10215 2420
rect 10175 2240 10215 2250
rect 10285 2420 10325 2430
rect 10285 2250 10295 2420
rect 10315 2250 10325 2420
rect 9525 2180 9785 2220
rect 10015 2210 10055 2240
rect 10015 2190 10025 2210
rect 10045 2190 10055 2210
rect 10015 2180 10055 2190
rect 10285 2220 10325 2250
rect 10395 2420 10435 2430
rect 10395 2250 10405 2420
rect 10425 2250 10435 2420
rect 10395 2240 10435 2250
rect 10505 2420 10545 2430
rect 10505 2250 10515 2420
rect 10535 2250 10545 2420
rect 10505 2220 10545 2250
rect 10615 2420 10655 2430
rect 10615 2250 10625 2420
rect 10645 2250 10655 2420
rect 10615 2240 10655 2250
rect 10725 2420 10815 2430
rect 10725 2250 10735 2420
rect 10755 2250 10785 2420
rect 10805 2250 10815 2420
rect 10725 2240 10815 2250
rect 10285 2180 10545 2220
rect 10725 2210 10765 2240
rect 10725 2190 10735 2210
rect 10755 2190 10765 2210
rect 10725 2180 10765 2190
rect 9745 2135 9785 2180
rect 8815 2080 9410 2100
rect 9745 2095 10005 2135
rect 9370 2060 9410 2080
rect 9205 2050 9245 2060
rect 9205 2030 9215 2050
rect 9235 2030 9245 2050
rect 9205 2000 9245 2030
rect 9370 2050 9520 2060
rect 9370 2030 9380 2050
rect 9400 2030 9490 2050
rect 9510 2030 9520 2050
rect 9370 2020 9520 2030
rect 9695 2050 9735 2060
rect 9695 2030 9705 2050
rect 9725 2030 9735 2050
rect 9155 1990 9245 2000
rect 9155 1820 9165 1990
rect 9185 1820 9215 1990
rect 9235 1820 9245 1990
rect 9155 1810 9245 1820
rect 9315 1990 9355 2000
rect 9315 1820 9325 1990
rect 9345 1820 9355 1990
rect 9315 1810 9355 1820
rect 9425 1990 9465 2020
rect 9695 2000 9735 2030
rect 9425 1820 9435 1990
rect 9455 1820 9465 1990
rect 9425 1810 9465 1820
rect 9535 1990 9575 2000
rect 9535 1820 9545 1990
rect 9565 1820 9575 1990
rect 9535 1810 9575 1820
rect 9645 1990 9785 2000
rect 9645 1820 9655 1990
rect 9675 1820 9705 1990
rect 9725 1820 9755 1990
rect 9775 1820 9785 1990
rect 9645 1810 9785 1820
rect 9855 1990 9895 2000
rect 9855 1820 9865 1990
rect 9885 1820 9895 1990
rect 9855 1810 9895 1820
rect 9965 1990 10005 2095
rect 10235 2050 10275 2060
rect 10235 2030 10245 2050
rect 10265 2030 10275 2050
rect 10235 2000 10275 2030
rect 9965 1820 9975 1990
rect 9995 1820 10005 1990
rect 9965 1810 10005 1820
rect 10075 1990 10115 2000
rect 10075 1820 10085 1990
rect 10105 1820 10115 1990
rect 10075 1810 10115 1820
rect 10185 1990 10325 2000
rect 10185 1820 10195 1990
rect 10215 1820 10245 1990
rect 10265 1820 10295 1990
rect 10315 1820 10325 1990
rect 10185 1810 10325 1820
rect 10395 1990 10435 2000
rect 10395 1820 10405 1990
rect 10425 1820 10435 1990
rect 10395 1810 10435 1820
rect 10505 1990 10545 2180
rect 10725 2050 10765 2060
rect 10725 2030 10735 2050
rect 10755 2030 10765 2050
rect 10725 2000 10765 2030
rect 10505 1820 10515 1990
rect 10535 1820 10545 1990
rect 10505 1810 10545 1820
rect 10615 1990 10655 2000
rect 10615 1820 10625 1990
rect 10645 1820 10655 1990
rect 10615 1810 10655 1820
rect 10725 1990 10815 2000
rect 10725 1820 10735 1990
rect 10755 1820 10785 1990
rect 10805 1820 10815 1990
rect 10725 1810 10815 1820
rect 10555 1770 10945 1780
rect 10555 1735 10565 1770
rect 10600 1735 10900 1770
rect 10935 1735 10945 1770
rect 10555 1725 10945 1735
rect 8250 1550 10945 1560
rect 8250 1515 10900 1550
rect 10935 1515 10945 1550
rect 8250 1505 10945 1515
<< viali >>
rect 10860 2850 10895 2885
rect 10860 2470 10895 2505
rect 9265 2250 9285 2420
rect 9315 2250 9335 2420
rect 9425 2250 9445 2420
rect 9645 2250 9665 2420
rect 9865 2250 9885 2420
rect 9975 2250 9995 2420
rect 10025 2250 10045 2420
rect 10075 2250 10095 2420
rect 10185 2250 10205 2420
rect 10405 2250 10425 2420
rect 10625 2250 10645 2420
rect 10735 2250 10755 2420
rect 10785 2250 10805 2420
rect 9165 1820 9185 1990
rect 9215 1820 9235 1990
rect 9325 1820 9345 1990
rect 9545 1820 9565 1990
rect 9655 1820 9675 1990
rect 9705 1820 9725 1990
rect 9755 1820 9775 1990
rect 9865 1820 9885 1990
rect 10085 1820 10105 1990
rect 10195 1820 10215 1990
rect 10245 1820 10265 1990
rect 10295 1820 10315 1990
rect 10405 1820 10425 1990
rect 10625 1820 10645 1990
rect 10735 1820 10755 1990
rect 10785 1820 10805 1990
rect 10900 1735 10935 1770
rect 10900 1515 10935 1550
<< metal1 >>
rect 10850 2885 10905 2895
rect 10850 2850 10860 2885
rect 10895 2850 10905 2885
rect 10850 2840 10905 2850
rect 10850 2505 10905 2515
rect 10850 2470 10860 2505
rect 10895 2470 10905 2505
rect 10850 2460 10905 2470
rect 9250 2430 10820 2435
rect 9220 2420 10820 2430
rect 9220 2250 9265 2420
rect 9285 2250 9315 2420
rect 9335 2250 9425 2420
rect 9445 2250 9645 2420
rect 9665 2250 9865 2420
rect 9885 2250 9975 2420
rect 9995 2250 10025 2420
rect 10045 2250 10075 2420
rect 10095 2250 10185 2420
rect 10205 2250 10405 2420
rect 10425 2250 10625 2420
rect 10645 2250 10735 2420
rect 10755 2250 10785 2420
rect 10805 2250 10820 2420
rect 9220 2240 10820 2250
rect 9250 2235 10820 2240
rect 9060 1990 10820 2005
rect 9060 1820 9165 1990
rect 9185 1820 9215 1990
rect 9235 1820 9325 1990
rect 9345 1820 9545 1990
rect 9565 1820 9655 1990
rect 9675 1820 9705 1990
rect 9725 1820 9755 1990
rect 9775 1820 9865 1990
rect 9885 1820 10085 1990
rect 10105 1820 10195 1990
rect 10215 1820 10245 1990
rect 10265 1820 10295 1990
rect 10315 1820 10405 1990
rect 10425 1820 10625 1990
rect 10645 1820 10735 1990
rect 10755 1820 10785 1990
rect 10805 1820 10820 1990
rect 9060 1805 10820 1820
rect 10890 1770 10945 1780
rect 10890 1735 10900 1770
rect 10935 1735 10945 1770
rect 10890 1725 10945 1735
rect 10890 1550 10945 1560
rect 10890 1515 10900 1550
rect 10935 1515 10945 1550
rect 10890 1505 10945 1515
<< via1 >>
rect 10860 2850 10895 2885
rect 10860 2470 10895 2505
rect 10900 1735 10935 1770
rect 10900 1515 10935 1550
<< metal2 >>
rect 10850 2885 10905 2895
rect 10850 2850 10860 2885
rect 10895 2850 10905 2885
rect 10850 2840 10905 2850
rect 10850 2505 10905 2515
rect 10850 2470 10860 2505
rect 10895 2470 10905 2505
rect 10850 2460 10905 2470
rect 10890 1770 10945 1780
rect 10890 1735 10900 1770
rect 10935 1735 10945 1770
rect 10890 1725 10945 1735
rect 10890 1550 10945 1560
rect 10890 1515 10900 1550
rect 10935 1515 10945 1550
rect 10890 1505 10945 1515
<< via2 >>
rect 10860 2850 10895 2885
rect 10860 2470 10895 2505
rect 10900 1735 10935 1770
rect 10900 1515 10935 1550
<< metal3 >>
rect 10850 2885 11655 2895
rect 10850 2850 10860 2885
rect 10895 2850 11655 2885
rect 10850 2840 11655 2850
rect 10850 2505 10905 2515
rect 10850 2470 10860 2505
rect 10895 2470 10905 2505
rect 10850 2460 10905 2470
rect 11025 2445 11655 2840
rect 10890 1770 10945 1780
rect 10890 1735 10900 1770
rect 10935 1735 10945 1770
rect 10890 1725 10945 1735
rect 11065 1560 11355 1795
rect 10890 1550 11355 1560
rect 10890 1515 10900 1550
rect 10935 1515 11355 1550
rect 10890 1505 11355 1515
<< via3 >>
rect 10860 2470 10895 2505
rect 10900 1735 10935 1770
<< mimcap >>
rect 11040 2505 11640 2880
rect 11040 2470 11050 2505
rect 11085 2470 11640 2505
rect 11040 2460 11640 2470
rect 11080 1770 11340 1780
rect 11080 1735 11090 1770
rect 11125 1735 11340 1770
rect 11080 1520 11340 1735
<< mimcapcontact >>
rect 11050 2470 11085 2505
rect 11090 1735 11125 1770
<< metal4 >>
rect 10850 2505 11095 2515
rect 10850 2470 10860 2505
rect 10895 2470 11050 2505
rect 11085 2470 11095 2505
rect 10850 2460 11095 2470
rect 10890 1770 11135 1780
rect 10890 1735 10900 1770
rect 10935 1735 11090 1770
rect 11125 1735 11135 1770
rect 10890 1725 11135 1735
<< labels >>
flabel locali 8815 2090 8815 2090 7 FreeSans 400 0 -200 0 I_IN
flabel locali 10545 2105 10545 2105 3 FreeSans 400 0 160 0 vout
flabel metal1 9220 2285 9220 2285 7 FreeSans 400 0 -200 0 VDDA
flabel metal1 9060 1950 9060 1950 7 FreeSans 400 0 -200 0 GNDA
flabel locali 8250 1530 8250 1530 7 FreeSans 400 0 -200 0 DOWN
flabel locali 10005 2120 10005 2120 3 FreeSans 400 0 200 0 x
flabel locali 8205 2870 8205 2870 7 FreeSans 400 0 -200 0 UP_b
<< end >>
