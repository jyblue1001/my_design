* PEX produced on Thu Jul  3 03:10:36 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic_5.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic_5 VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 VDDA.t300 bgr_0.V_TOP.t14 bgr_0.Vin-.t7 VDDA.t299 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X1 bgr_0.1st_Vout_1.t11 bgr_0.cap_res1.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2 a_14640_5738.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 GNDA.t176 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X3 bgr_0.V_TOP.t15 VDDA.t298 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4 two_stage_opamp_dummy_magic_0.VD2.t19 GNDA.t334 GNDA.t336 GNDA.t335 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X5 VOUT-.t19 two_stage_opamp_dummy_magic_0.cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 GNDA.t243 GNDA.t333 bgr_0.Vbe2.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X7 VOUT-.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8 VOUT-.t21 two_stage_opamp_dummy_magic_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 bgr_0.NFET_GATE_10uA.t1 bgr_0.NFET_GATE_10uA.t0 GNDA.t118 GNDA.t117 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X10 bgr_0.1st_Vout_1.t12 bgr_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X11 bgr_0.V_TOP.t16 VDDA.t297 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 VDDA.t457 bgr_0.V_mir2.t15 bgr_0.V_mir2.t16 VDDA.t456 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X13 VOUT-.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X14 two_stage_opamp_dummy_magic_0.V_err_gate.t4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X15 VOUT-.t23 two_stage_opamp_dummy_magic_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 GNDA.t63 two_stage_opamp_dummy_magic_0.X.t25 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X17 two_stage_opamp_dummy_magic_0.X.t22 GNDA.t330 GNDA.t332 GNDA.t331 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X18 VOUT-.t24 two_stage_opamp_dummy_magic_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X19 VOUT-.t25 two_stage_opamp_dummy_magic_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 VOUT-.t26 two_stage_opamp_dummy_magic_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 VDDA.t17 two_stage_opamp_dummy_magic_0.X.t26 VOUT-.t2 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X22 VDDA.t104 bgr_0.PFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X23 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 two_stage_opamp_dummy_magic_0.Y.t25 VDDA.t145 GNDA.t126 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X24 bgr_0.V_TOP.t17 VDDA.t296 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 VDDA.t438 bgr_0.V_mir1.t17 bgr_0.1st_Vout_1.t8 VDDA.t437 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X26 VOUT+.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 bgr_0.START_UP_NFET1.t0 bgr_0.START_UP_NFET1 GNDA.t100 GNDA.t99 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X28 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 a_5750_2946.t0 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X29 VOUT+.t20 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 VOUT+.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 VOUT-.t27 two_stage_opamp_dummy_magic_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 VDDA.t190 two_stage_opamp_dummy_magic_0.V_err_gate.t14 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 VDDA.t189 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X33 two_stage_opamp_dummy_magic_0.VD3.t15 two_stage_opamp_dummy_magic_0.VD3.t13 two_stage_opamp_dummy_magic_0.X.t13 two_stage_opamp_dummy_magic_0.VD3.t14 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X34 VOUT-.t28 two_stage_opamp_dummy_magic_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 VOUT-.t29 two_stage_opamp_dummy_magic_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 VOUT+.t22 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 bgr_0.1st_Vout_1.t13 bgr_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 GNDA.t48 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X39 VOUT-.t30 two_stage_opamp_dummy_magic_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 bgr_0.V_mir2.t1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 bgr_0.V_p_2.t5 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X41 bgr_0.Vin-.t5 bgr_0.V_TOP.t18 VDDA.t295 VDDA.t294 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X42 GNDA.t167 bgr_0.NFET_GATE_10uA.t5 two_stage_opamp_dummy_magic_0.Vb2.t5 GNDA.t166 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X43 VDDA.t166 two_stage_opamp_dummy_magic_0.Vb3.t8 two_stage_opamp_dummy_magic_0.VD3.t19 VDDA.t165 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X44 GNDA.t169 bgr_0.NFET_GATE_10uA.t6 two_stage_opamp_dummy_magic_0.Vb2.t4 GNDA.t168 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X45 VDDA.t415 VDDA.t413 two_stage_opamp_dummy_magic_0.V_err_gate.t12 VDDA.t414 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X46 VOUT-.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 VOUT+.t23 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X48 two_stage_opamp_dummy_magic_0.Y.t22 GNDA.t327 GNDA.t329 GNDA.t328 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X49 two_stage_opamp_dummy_magic_0.Y.t1 two_stage_opamp_dummy_magic_0.Vb1.t6 two_stage_opamp_dummy_magic_0.VD1.t15 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X50 VOUT+.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 VOUT+.t25 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 two_stage_opamp_dummy_magic_0.V_err_p.t15 two_stage_opamp_dummy_magic_0.V_err_gate.t15 VDDA.t443 VDDA.t442 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X53 VOUT-.t3 two_stage_opamp_dummy_magic_0.X.t27 VDDA.t19 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X54 bgr_0.1st_Vout_1.t1 bgr_0.Vin+.t6 bgr_0.V_p_1.t4 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X55 two_stage_opamp_dummy_magic_0.V_err_p.t16 two_stage_opamp_dummy_magic_0.V_tot.t4 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 VDDA.t228 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X56 VOUT+.t26 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X57 bgr_0.1st_Vout_2.t11 bgr_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X58 VDDA.t412 VDDA.t410 bgr_0.V_TOP.t1 VDDA.t411 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X59 two_stage_opamp_dummy_magic_0.VD1.t16 VIN-.t0 two_stage_opamp_dummy_magic_0.V_p.t25 GNDA.t185 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X60 VOUT+.t27 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 GNDA.t171 bgr_0.NFET_GATE_10uA.t7 two_stage_opamp_dummy_magic_0.Vb2.t3 GNDA.t170 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X62 GNDA.t326 GNDA.t324 two_stage_opamp_dummy_magic_0.Vb2.t8 GNDA.t325 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X63 VDDA.t129 bgr_0.V_mir1.t18 bgr_0.1st_Vout_1.t3 VDDA.t128 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X64 VOUT-.t32 two_stage_opamp_dummy_magic_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X65 VOUT+.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 two_stage_opamp_dummy_magic_0.V_err_p.t14 two_stage_opamp_dummy_magic_0.V_err_gate.t16 VDDA.t40 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X67 VOUT+.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 VOUT+.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X69 GNDA.t194 two_stage_opamp_dummy_magic_0.Y.t26 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 VDDA.t226 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X70 VOUT-.t33 two_stage_opamp_dummy_magic_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X71 two_stage_opamp_dummy_magic_0.VD1.t0 VIN-.t1 two_stage_opamp_dummy_magic_0.V_p.t24 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X72 VDDA.t195 two_stage_opamp_dummy_magic_0.Vb3.t9 two_stage_opamp_dummy_magic_0.VD3.t20 VDDA.t194 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X73 VOUT+.t31 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 two_stage_opamp_dummy_magic_0.X.t1 two_stage_opamp_dummy_magic_0.Vb2.t11 two_stage_opamp_dummy_magic_0.VD3.t3 two_stage_opamp_dummy_magic_0.VD3.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X75 bgr_0.NFET_GATE_10uA.t2 bgr_0.PFET_GATE_10uA.t11 VDDA.t110 VDDA.t109 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X76 bgr_0.1st_Vout_2.t12 bgr_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X77 VDDA.t455 bgr_0.PFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 VDDA.t454 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X78 VOUT-.t34 two_stage_opamp_dummy_magic_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 GNDA.t137 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 VOUT+.t3 GNDA.t136 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X80 VDDA.t409 VDDA.t407 bgr_0.NFET_GATE_10uA.t3 VDDA.t408 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X81 GNDA.t82 two_stage_opamp_dummy_magic_0.X.t28 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X82 GNDA.t152 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 two_stage_opamp_dummy_magic_0.V_p.t28 GNDA.t151 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X83 VDDA.t206 bgr_0.1st_Vout_1.t14 bgr_0.V_TOP.t5 VDDA.t205 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X84 VOUT+.t32 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 GNDA.t323 GNDA.t321 two_stage_opamp_dummy_magic_0.VD1.t19 GNDA.t322 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X86 VOUT+.t33 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X87 VOUT-.t35 two_stage_opamp_dummy_magic_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 VOUT+.t34 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 VDDA.t204 bgr_0.V_mir2.t13 bgr_0.V_mir2.t14 VDDA.t203 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X90 GNDA.t163 bgr_0.NFET_GATE_10uA.t8 two_stage_opamp_dummy_magic_0.Vb3.t5 GNDA.t162 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X91 VOUT-.t36 two_stage_opamp_dummy_magic_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X92 two_stage_opamp_dummy_magic_0.Vb3.t4 bgr_0.NFET_GATE_10uA.t9 GNDA.t165 GNDA.t164 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X93 VOUT+.t18 two_stage_opamp_dummy_magic_0.Y.t27 VDDA.t121 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X94 GNDA.t320 GNDA.t318 GNDA.t320 GNDA.t319 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0 ps=0 w=2.5 l=0.15
X95 GNDA.t317 GNDA.t315 two_stage_opamp_dummy_magic_0.VD1.t18 GNDA.t316 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X96 VDDA.t208 bgr_0.1st_Vout_1.t15 bgr_0.V_TOP.t6 VDDA.t207 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X97 VDDA.t67 two_stage_opamp_dummy_magic_0.V_err_gate.t17 two_stage_opamp_dummy_magic_0.V_err_p.t13 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X98 VOUT+.t35 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X99 bgr_0.V_TOP.t4 bgr_0.cap_res1.t0 GNDA.t112 sky130_fd_pr__res_high_po_0p35 l=2.05
X100 GNDA.t314 GNDA.t312 VOUT+.t8 GNDA.t313 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X101 a_11220_17410.t0 GNDA.t71 GNDA.t53 sky130_fd_pr__res_xhigh_po_0p35 l=6
X102 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 two_stage_opamp_dummy_magic_0.X.t29 VDDA.t87 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X103 two_stage_opamp_dummy_magic_0.X.t17 two_stage_opamp_dummy_magic_0.Vb2.t12 two_stage_opamp_dummy_magic_0.VD3.t27 two_stage_opamp_dummy_magic_0.VD3.t26 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X104 two_stage_opamp_dummy_magic_0.Vb1.t1 bgr_0.PFET_GATE_10uA.t13 VDDA.t27 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X105 GNDA.t311 GNDA.t309 two_stage_opamp_dummy_magic_0.X.t21 GNDA.t310 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X106 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 two_stage_opamp_dummy_magic_0.V_err_gate.t18 VDDA.t192 VDDA.t191 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X107 VOUT-.t7 two_stage_opamp_dummy_magic_0.X.t30 VDDA.t94 VDDA.t93 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X108 VOUT+.t36 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X109 bgr_0.PFET_GATE_10uA.t5 bgr_0.1st_Vout_2.t13 VDDA.t246 VDDA.t245 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X110 VOUT+.t37 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 VOUT+.t38 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X112 VOUT+.t39 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 VOUT+.t40 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 a_14640_5738.t0 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA.t69 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X115 VOUT-.t37 two_stage_opamp_dummy_magic_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X116 VOUT-.t38 two_stage_opamp_dummy_magic_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X117 VDDA.t23 bgr_0.V_mir1.t10 bgr_0.V_mir1.t11 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X118 VOUT-.t39 two_stage_opamp_dummy_magic_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 VDDA.t406 VDDA.t404 two_stage_opamp_dummy_magic_0.VD3.t32 VDDA.t405 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X120 VOUT-.t40 two_stage_opamp_dummy_magic_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 GNDA.t186 two_stage_opamp_dummy_magic_0.Y.t28 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 VDDA.t216 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X122 VOUT-.t41 two_stage_opamp_dummy_magic_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 bgr_0.1st_Vout_1.t16 bgr_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 VDDA.t29 bgr_0.1st_Vout_2.t14 bgr_0.PFET_GATE_10uA.t1 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X125 bgr_0.V_TOP.t19 VDDA.t293 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 VDDA.t95 two_stage_opamp_dummy_magic_0.X.t31 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X127 two_stage_opamp_dummy_magic_0.VD4.t21 two_stage_opamp_dummy_magic_0.Vb2.t13 two_stage_opamp_dummy_magic_0.Y.t8 two_stage_opamp_dummy_magic_0.VD4.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X128 VOUT+.t41 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 bgr_0.1st_Vout_1.t17 bgr_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 GNDA.t308 GNDA.t306 two_stage_opamp_dummy_magic_0.Y.t21 GNDA.t307 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X131 GNDA.t129 two_stage_opamp_dummy_magic_0.X.t32 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 VDDA.t152 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X132 VOUT+.t42 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 GNDA.t144 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 two_stage_opamp_dummy_magic_0.V_p.t27 GNDA.t143 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X134 GNDA.t130 two_stage_opamp_dummy_magic_0.X.t33 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X135 two_stage_opamp_dummy_magic_0.X.t23 two_stage_opamp_dummy_magic_0.Vb1.t7 two_stage_opamp_dummy_magic_0.VD2.t20 GNDA.t349 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X136 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 GNDA.t303 GNDA.t305 GNDA.t304 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X137 VOUT+.t43 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 VOUT-.t42 two_stage_opamp_dummy_magic_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 two_stage_opamp_dummy_magic_0.V_p.t3 VIN+.t0 two_stage_opamp_dummy_magic_0.VD2.t1 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X140 VOUT+.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X141 VDDA.t97 bgr_0.V_mir2.t17 bgr_0.1st_Vout_2.t7 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X142 VOUT-.t12 a_5750_2946.t1 GNDA.t142 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X143 VOUT-.t43 two_stage_opamp_dummy_magic_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 VOUT-.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 bgr_0.1st_Vout_1.t18 bgr_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X146 a_13730_17020.t0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 GNDA.t33 sky130_fd_pr__res_xhigh_po_0p35 l=6.3
X147 VOUT+.t17 two_stage_opamp_dummy_magic_0.Y.t29 VDDA.t157 VDDA.t156 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X148 two_stage_opamp_dummy_magic_0.V_p.t0 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 GNDA.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X149 two_stage_opamp_dummy_magic_0.V_p.t4 VIN+.t1 two_stage_opamp_dummy_magic_0.VD2.t2 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X150 VOUT+.t45 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 bgr_0.V_CUR_REF_REG.t2 VDDA.t401 VDDA.t403 VDDA.t402 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X152 a_11220_17410.t1 a_12828_17530.t0 GNDA.t53 sky130_fd_pr__res_xhigh_po_0p35 l=6
X153 VOUT+.t46 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 two_stage_opamp_dummy_magic_0.VD3.t35 two_stage_opamp_dummy_magic_0.Vb3.t10 VDDA.t421 VDDA.t420 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X155 VOUT-.t45 two_stage_opamp_dummy_magic_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X156 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 bgr_0.PFET_GATE_10uA.t14 VDDA.t178 VDDA.t177 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X157 VOUT+.t47 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 VOUT+.t48 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 VDDA.t213 bgr_0.PFET_GATE_10uA.t15 bgr_0.V_CUR_REF_REG.t1 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X160 VOUT+.t49 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X161 bgr_0.PFET_GATE_10uA.t3 bgr_0.cap_res2.t20 GNDA.t112 sky130_fd_pr__res_high_po_0p35 l=2.05
X162 VOUT+.t7 GNDA.t300 GNDA.t302 GNDA.t301 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X163 bgr_0.V_p_1.t9 bgr_0.Vin-.t8 bgr_0.V_mir1.t16 GNDA.t225 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X164 VDDA.t1 bgr_0.V_mir1.t8 bgr_0.V_mir1.t9 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X165 VOUT+.t50 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 VOUT+.t51 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X167 two_stage_opamp_dummy_magic_0.VD2.t16 two_stage_opamp_dummy_magic_0.Vb1.t8 two_stage_opamp_dummy_magic_0.X.t19 GNDA.t212 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X168 bgr_0.1st_Vout_2.t15 bgr_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X169 VOUT-.t46 two_stage_opamp_dummy_magic_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X170 VOUT-.t47 two_stage_opamp_dummy_magic_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 VDDA.t417 bgr_0.1st_Vout_1.t19 bgr_0.V_TOP.t11 VDDA.t416 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X172 VOUT-.t10 two_stage_opamp_dummy_magic_0.X.t34 VDDA.t168 VDDA.t167 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X173 VDDA.t292 bgr_0.V_TOP.t20 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 VDDA.t291 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X174 VOUT-.t11 two_stage_opamp_dummy_magic_0.X.t35 VDDA.t170 VDDA.t169 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X175 VDDA.t227 two_stage_opamp_dummy_magic_0.Y.t30 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 GNDA.t195 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X176 VOUT-.t48 two_stage_opamp_dummy_magic_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 VOUT-.t49 two_stage_opamp_dummy_magic_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X178 bgr_0.V_p_2.t8 bgr_0.V_CUR_REF_REG.t3 bgr_0.1st_Vout_2.t9 GNDA.t216 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X179 VOUT-.t9 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 GNDA.t132 GNDA.t131 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X180 two_stage_opamp_dummy_magic_0.cap_res_X.t0 two_stage_opamp_dummy_magic_0.X.t11 GNDA.t111 sky130_fd_pr__res_high_po_1p41 l=1.41
X181 VOUT-.t50 two_stage_opamp_dummy_magic_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 GNDA.t191 two_stage_opamp_dummy_magic_0.Y.t31 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 VDDA.t225 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X183 VOUT+.t52 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X184 two_stage_opamp_dummy_magic_0.VD3.t30 two_stage_opamp_dummy_magic_0.Vb3.t11 VDDA.t243 VDDA.t242 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X185 VOUT+.t53 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 bgr_0.V_p_1.t8 bgr_0.Vin-.t9 bgr_0.V_mir1.t13 GNDA.t224 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X187 two_stage_opamp_dummy_magic_0.VD3.t29 two_stage_opamp_dummy_magic_0.Vb2.t14 two_stage_opamp_dummy_magic_0.X.t18 two_stage_opamp_dummy_magic_0.VD3.t28 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X188 bgr_0.1st_Vout_2.t16 bgr_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 two_stage_opamp_dummy_magic_0.err_amp_out.t9 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 GNDA.t59 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X190 bgr_0.V_TOP.t13 VDDA.t398 VDDA.t400 VDDA.t399 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X191 VDDA.t79 two_stage_opamp_dummy_magic_0.X.t36 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X192 VOUT-.t51 two_stage_opamp_dummy_magic_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X193 bgr_0.Vin-.t1 bgr_0.START_UP.t6 bgr_0.V_TOP.t3 VDDA.t193 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X194 two_stage_opamp_dummy_magic_0.VD1.t14 two_stage_opamp_dummy_magic_0.Vb1.t9 two_stage_opamp_dummy_magic_0.Y.t20 GNDA.t235 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X195 VOUT-.t52 two_stage_opamp_dummy_magic_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 VOUT+.t54 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 bgr_0.1st_Vout_1.t20 bgr_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 bgr_0.V_TOP.t21 VDDA.t282 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 VDDA.t397 VDDA.t395 two_stage_opamp_dummy_magic_0.V_err_p.t18 VDDA.t396 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X200 VOUT-.t53 two_stage_opamp_dummy_magic_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X201 VOUT-.t54 two_stage_opamp_dummy_magic_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 VOUT-.t55 two_stage_opamp_dummy_magic_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X203 GNDA.t351 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 two_stage_opamp_dummy_magic_0.V_p.t40 GNDA.t350 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X204 two_stage_opamp_dummy_magic_0.err_amp_out.t4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 two_stage_opamp_dummy_magic_0.V_err_p.t2 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X205 GNDA.t78 two_stage_opamp_dummy_magic_0.X.t37 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 VDDA.t80 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X206 a_5230_5738.t1 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA.t32 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X207 a_13730_17020.t1 GNDA.t98 GNDA.t33 sky130_fd_pr__res_xhigh_po_0p35 l=6.3
X208 bgr_0.1st_Vout_1.t21 bgr_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 bgr_0.V_TOP.t22 VDDA.t281 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 VDDA.t392 VDDA.t394 VDDA.t393 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X211 a_11220_17290.t1 a_12828_17650.t1 GNDA.t53 sky130_fd_pr__res_xhigh_po_0p35 l=6
X212 VOUT+.t55 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 VOUT+.t56 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X214 VOUT+.t57 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X215 VOUT-.t56 two_stage_opamp_dummy_magic_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 bgr_0.V_p_2.t6 bgr_0.V_CUR_REF_REG.t4 bgr_0.1st_Vout_2.t1 GNDA.t138 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X217 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 bgr_0.PFET_GATE_10uA.t16 VDDA.t202 VDDA.t201 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X218 VOUT+.t58 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X219 VDDA.t453 bgr_0.PFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 VDDA.t452 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X220 two_stage_opamp_dummy_magic_0.V_p.t15 VIN+.t2 two_stage_opamp_dummy_magic_0.VD2.t11 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X221 VOUT-.t57 two_stage_opamp_dummy_magic_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 two_stage_opamp_dummy_magic_0.V_p.t39 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 GNDA.t343 GNDA.t342 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X223 VDDA.t182 two_stage_opamp_dummy_magic_0.Vb3.t12 two_stage_opamp_dummy_magic_0.VD4.t37 VDDA.t181 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X224 VOUT+.t16 two_stage_opamp_dummy_magic_0.Y.t32 VDDA.t133 VDDA.t132 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X225 a_11220_17290.t0 GNDA.t119 GNDA.t53 sky130_fd_pr__res_xhigh_po_0p35 l=6
X226 two_stage_opamp_dummy_magic_0.Y.t3 two_stage_opamp_dummy_magic_0.VD4.t25 two_stage_opamp_dummy_magic_0.VD4.t27 two_stage_opamp_dummy_magic_0.VD4.t26 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X227 two_stage_opamp_dummy_magic_0.V_p.t23 VIN-.t2 two_stage_opamp_dummy_magic_0.VD1.t20 GNDA.t344 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X228 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 GNDA.t297 GNDA.t299 GNDA.t298 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X229 bgr_0.1st_Vout_1.t22 bgr_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 VOUT-.t58 two_stage_opamp_dummy_magic_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X231 bgr_0.START_UP.t3 bgr_0.V_TOP.t23 VDDA.t290 VDDA.t289 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X232 bgr_0.1st_Vout_2.t6 bgr_0.V_mir2.t18 VDDA.t112 VDDA.t111 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X233 bgr_0.V_TOP.t24 VDDA.t288 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X234 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t3 VDDA.t198 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X235 VOUT-.t59 two_stage_opamp_dummy_magic_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 VOUT-.t60 two_stage_opamp_dummy_magic_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X237 VOUT+.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X238 VOUT+.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 VDDA.t125 bgr_0.V_mir1.t19 bgr_0.1st_Vout_1.t2 VDDA.t124 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X240 two_stage_opamp_dummy_magic_0.VD2.t10 two_stage_opamp_dummy_magic_0.Vb1.t10 two_stage_opamp_dummy_magic_0.X.t9 GNDA.t92 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X241 VOUT-.t61 two_stage_opamp_dummy_magic_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X242 a_14520_5738.t0 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA.t110 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X243 VOUT-.t4 two_stage_opamp_dummy_magic_0.X.t38 VDDA.t77 VDDA.t76 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X244 VOUT-.t62 two_stage_opamp_dummy_magic_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 bgr_0.1st_Vout_1.t23 bgr_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 VDDA.t459 two_stage_opamp_dummy_magic_0.Y.t33 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 GNDA.t346 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X247 bgr_0.V_p_2.t10 bgr_0.V_CUR_REF_REG.t5 bgr_0.1st_Vout_2.t10 GNDA.t354 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X248 VOUT+.t61 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X249 VOUT+.t62 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 VOUT-.t63 two_stage_opamp_dummy_magic_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X251 VOUT-.t64 two_stage_opamp_dummy_magic_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X252 VOUT+.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 bgr_0.V_TOP.t25 VDDA.t287 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 GNDA.t250 GNDA.t293 bgr_0.Vbe2.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X255 two_stage_opamp_dummy_magic_0.V_err_p.t17 VDDA.t389 VDDA.t391 VDDA.t390 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X256 GNDA.t139 two_stage_opamp_dummy_magic_0.Y.t34 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 VDDA.t183 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X257 VOUT+.t64 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 two_stage_opamp_dummy_magic_0.Y.t18 two_stage_opamp_dummy_magic_0.Vb2.t15 two_stage_opamp_dummy_magic_0.VD4.t19 two_stage_opamp_dummy_magic_0.VD4.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X259 GNDA.t75 two_stage_opamp_dummy_magic_0.Y.t35 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X260 VOUT-.t65 two_stage_opamp_dummy_magic_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X261 VOUT-.t66 two_stage_opamp_dummy_magic_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 two_stage_opamp_dummy_magic_0.err_amp_out.t8 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 GNDA.t107 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X263 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 GNDA.t348 GNDA.t347 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X264 VDDA.t78 two_stage_opamp_dummy_magic_0.X.t39 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X265 VOUT+.t65 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 bgr_0.1st_Vout_2.t17 bgr_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X267 GNDA.t159 bgr_0.NFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t6 GNDA.t158 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X268 two_stage_opamp_dummy_magic_0.Vb3.t7 two_stage_opamp_dummy_magic_0.Vb2.t16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4 as=0.72 ps=4 w=3.6 l=0.2
X269 VDDA.t43 two_stage_opamp_dummy_magic_0.X.t40 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X270 VOUT-.t67 two_stage_opamp_dummy_magic_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 VOUT+.t66 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X272 two_stage_opamp_dummy_magic_0.VD1.t13 two_stage_opamp_dummy_magic_0.Vb1.t11 two_stage_opamp_dummy_magic_0.Y.t17 GNDA.t204 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X273 VOUT-.t68 two_stage_opamp_dummy_magic_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X274 VDDA.t50 two_stage_opamp_dummy_magic_0.V_err_gate.t19 two_stage_opamp_dummy_magic_0.V_err_p.t12 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X275 VDDA.t116 two_stage_opamp_dummy_magic_0.V_err_gate.t20 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 VDDA.t115 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X276 bgr_0.V_mir2.t12 bgr_0.V_mir2.t11 VDDA.t465 VDDA.t464 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X277 VDDA.t286 bgr_0.V_TOP.t26 bgr_0.Vin-.t4 VDDA.t285 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X278 GNDA.t219 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 two_stage_opamp_dummy_magic_0.V_p.t35 GNDA.t218 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X279 VDDA.t388 VDDA.t386 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 VDDA.t387 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X280 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 two_stage_opamp_dummy_magic_0.V_tot.t5 two_stage_opamp_dummy_magic_0.V_err_p.t19 VDDA.t426 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X281 GNDA.t18 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 VOUT-.t0 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X282 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 bgr_0.PFET_GATE_10uA.t18 VDDA.t467 VDDA.t466 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X283 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 VIN+.t3 two_stage_opamp_dummy_magic_0.V_p_mir.t0 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X284 two_stage_opamp_dummy_magic_0.V_p.t22 VIN-.t3 two_stage_opamp_dummy_magic_0.VD1.t17 GNDA.t200 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X285 VOUT+.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 GNDA.t339 two_stage_opamp_dummy_magic_0.err_amp_out.t12 two_stage_opamp_dummy_magic_0.V_p.t38 GNDA.t338 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X287 VOUT-.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X288 VOUT+.t68 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X289 bgr_0.Vin-.t0 a_12828_17650.t0 GNDA.t53 sky130_fd_pr__res_xhigh_po_0p35 l=6
X290 VOUT+.t69 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X291 VOUT-.t70 two_stage_opamp_dummy_magic_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 VDDA.t430 two_stage_opamp_dummy_magic_0.Vb3.t13 two_stage_opamp_dummy_magic_0.VD3.t36 VDDA.t429 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X293 VOUT-.t71 two_stage_opamp_dummy_magic_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X294 GNDA.t252 GNDA.t292 bgr_0.Vbe2.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X295 VOUT+.t15 two_stage_opamp_dummy_magic_0.Y.t36 VDDA.t143 VDDA.t142 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X296 two_stage_opamp_dummy_magic_0.V_p.t21 VIN-.t4 two_stage_opamp_dummy_magic_0.VD1.t1 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X297 two_stage_opamp_dummy_magic_0.V_p.t9 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 GNDA.t52 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X298 VOUT+.t14 two_stage_opamp_dummy_magic_0.Y.t37 VDDA.t219 VDDA.t218 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X299 VOUT-.t72 two_stage_opamp_dummy_magic_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 VOUT+.t70 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 bgr_0.1st_Vout_2.t18 bgr_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 GNDA.t161 bgr_0.NFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 GNDA.t160 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X303 bgr_0.PFET_GATE_10uA.t9 bgr_0.1st_Vout_2.t19 VDDA.t425 VDDA.t424 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X304 VOUT-.t73 two_stage_opamp_dummy_magic_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X305 VOUT-.t74 two_stage_opamp_dummy_magic_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X306 VOUT-.t75 two_stage_opamp_dummy_magic_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X307 two_stage_opamp_dummy_magic_0.Vb2.t7 GNDA.t294 GNDA.t296 GNDA.t295 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X308 GNDA.t291 GNDA.t289 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 GNDA.t290 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X309 two_stage_opamp_dummy_magic_0.Vb2.t2 bgr_0.NFET_GATE_10uA.t12 GNDA.t173 GNDA.t172 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X310 bgr_0.START_UP.t5 bgr_0.START_UP.t4 bgr_0.START_UP_NFET1.t0 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X311 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 two_stage_opamp_dummy_magic_0.V_tot.t6 two_stage_opamp_dummy_magic_0.V_err_gate.t10 VDDA.t229 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X312 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 two_stage_opamp_dummy_magic_0.V_tot.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t9 VDDA.t209 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X313 two_stage_opamp_dummy_magic_0.Y.t7 two_stage_opamp_dummy_magic_0.Vb2.t17 two_stage_opamp_dummy_magic_0.VD4.t17 two_stage_opamp_dummy_magic_0.VD4.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X314 VOUT-.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 VOUT+.t71 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 VDDA.t184 two_stage_opamp_dummy_magic_0.Y.t38 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 GNDA.t140 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X317 VOUT+.t72 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 VOUT+.t73 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 VOUT+.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 VOUT-.t77 two_stage_opamp_dummy_magic_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X321 VOUT-.t78 two_stage_opamp_dummy_magic_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X322 VOUT-.t79 two_stage_opamp_dummy_magic_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 GNDA.t175 bgr_0.NFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 GNDA.t174 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X324 bgr_0.V_p_1.t3 bgr_0.Vin+.t7 bgr_0.1st_Vout_1.t4 GNDA.t113 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X325 two_stage_opamp_dummy_magic_0.Vb2.t1 bgr_0.NFET_GATE_10uA.t14 GNDA.t182 GNDA.t181 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X326 two_stage_opamp_dummy_magic_0.Vb2.t0 bgr_0.NFET_GATE_10uA.t15 GNDA.t184 GNDA.t183 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X327 two_stage_opamp_dummy_magic_0.VD4.t1 VDDA.t383 VDDA.t385 VDDA.t384 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X328 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 two_stage_opamp_dummy_magic_0.V_err_gate.t21 VDDA.t440 VDDA.t439 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X329 GNDA.t228 VDDA.t380 VDDA.t382 VDDA.t381 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X330 bgr_0.1st_Vout_2.t20 bgr_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X331 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 GNDA.t215 GNDA.t214 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X332 bgr_0.Vin+.t5 bgr_0.V_TOP.t27 VDDA.t284 VDDA.t283 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X333 VOUT+.t75 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X334 VOUT+.t76 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X335 VOUT+.t77 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X336 VDDA.t44 two_stage_opamp_dummy_magic_0.X.t41 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X337 VOUT-.t80 two_stage_opamp_dummy_magic_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X338 VDDA.t176 bgr_0.PFET_GATE_10uA.t19 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 VDDA.t175 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X339 VOUT+.t78 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X340 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 bgr_0.PFET_GATE_10uA.t20 VDDA.t102 VDDA.t101 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X341 two_stage_opamp_dummy_magic_0.VD1.t12 two_stage_opamp_dummy_magic_0.Vb1.t12 two_stage_opamp_dummy_magic_0.Y.t4 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X342 VDDA.t65 two_stage_opamp_dummy_magic_0.V_err_gate.t22 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X343 a_5350_5738.t0 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA.t31 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X344 VOUT+.t79 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 GNDA.t208 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 two_stage_opamp_dummy_magic_0.V_p_mir.t3 GNDA.t207 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X346 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 two_stage_opamp_dummy_magic_0.V_tot.t8 two_stage_opamp_dummy_magic_0.V_err_p.t21 VDDA.t441 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X347 VOUT+.t80 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X348 VOUT-.t81 two_stage_opamp_dummy_magic_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X349 VOUT-.t82 two_stage_opamp_dummy_magic_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 bgr_0.V_TOP.t28 VDDA.t280 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 GNDA.t13 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 two_stage_opamp_dummy_magic_0.V_p.t2 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X352 bgr_0.Vin+.t1 a_12828_17530.t1 GNDA.t53 sky130_fd_pr__res_xhigh_po_0p35 l=6
X353 two_stage_opamp_dummy_magic_0.err_amp_out.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 two_stage_opamp_dummy_magic_0.V_err_p.t4 VDDA.t199 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X354 two_stage_opamp_dummy_magic_0.V_p.t5 VIN+.t4 two_stage_opamp_dummy_magic_0.VD2.t3 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X355 VOUT-.t83 two_stage_opamp_dummy_magic_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X356 VOUT+.t81 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X357 two_stage_opamp_dummy_magic_0.VD4.t36 two_stage_opamp_dummy_magic_0.Vb3.t14 VDDA.t70 VDDA.t69 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X358 bgr_0.1st_Vout_1.t24 bgr_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 two_stage_opamp_dummy_magic_0.Vb3.t6 GNDA.t286 GNDA.t288 GNDA.t287 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X360 two_stage_opamp_dummy_magic_0.VD4.t15 two_stage_opamp_dummy_magic_0.Vb2.t18 two_stage_opamp_dummy_magic_0.Y.t5 two_stage_opamp_dummy_magic_0.VD4.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X361 two_stage_opamp_dummy_magic_0.Vb3.t3 bgr_0.NFET_GATE_10uA.t16 GNDA.t95 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X362 VDDA.t379 VDDA.t376 VDDA.t378 VDDA.t377 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.06 as=0 ps=0 w=0.63 l=0.2
X363 GNDA.t97 bgr_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_0.Vb3.t2 GNDA.t96 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X364 VOUT+.t6 VDDA.t373 VDDA.t375 VDDA.t374 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X365 two_stage_opamp_dummy_magic_0.V_p.t34 VIN+.t5 two_stage_opamp_dummy_magic_0.VD2.t15 GNDA.t211 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X366 two_stage_opamp_dummy_magic_0.V_p.t7 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 GNDA.t43 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X367 bgr_0.V_mir1.t7 bgr_0.V_mir1.t6 VDDA.t436 VDDA.t435 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X368 VOUT+.t82 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X369 VOUT+.t83 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X370 VOUT+.t84 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X371 bgr_0.V_p_2.t4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 bgr_0.V_mir2.t2 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X372 VOUT+.t85 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 VDDA.t108 bgr_0.PFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_0.Vb1.t0 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X374 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 two_stage_opamp_dummy_magic_0.V_err_gate.t2 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X375 two_stage_opamp_dummy_magic_0.VD2.t9 two_stage_opamp_dummy_magic_0.Vb1.t13 two_stage_opamp_dummy_magic_0.X.t8 GNDA.t88 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X376 VOUT-.t84 two_stage_opamp_dummy_magic_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X377 VOUT+.t86 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X378 VDDA.t164 two_stage_opamp_dummy_magic_0.Y.t39 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 GNDA.t135 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X379 VOUT-.t85 two_stage_opamp_dummy_magic_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X380 VDDA.t98 two_stage_opamp_dummy_magic_0.Y.t40 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X381 bgr_0.V_p_1.t2 bgr_0.Vin+.t8 bgr_0.1st_Vout_1.t6 GNDA.t141 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X382 VOUT+.t87 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 VDDA.t279 bgr_0.V_TOP.t29 bgr_0.START_UP.t2 VDDA.t278 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X384 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_0.Y.t11 GNDA.t124 sky130_fd_pr__res_high_po_1p41 l=1.41
X385 two_stage_opamp_dummy_magic_0.VD4.t13 two_stage_opamp_dummy_magic_0.Vb2.t19 two_stage_opamp_dummy_magic_0.Y.t13 two_stage_opamp_dummy_magic_0.VD4.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X386 VOUT+.t88 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X387 bgr_0.1st_Vout_2.t21 bgr_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 bgr_0.V_mir1.t5 bgr_0.V_mir1.t4 VDDA.t74 VDDA.t73 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X389 two_stage_opamp_dummy_magic_0.V_err_p.t11 two_stage_opamp_dummy_magic_0.V_err_gate.t23 VDDA.t5 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X390 VOUT-.t86 two_stage_opamp_dummy_magic_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X391 two_stage_opamp_dummy_magic_0.X.t12 two_stage_opamp_dummy_magic_0.Vb2.t20 two_stage_opamp_dummy_magic_0.VD3.t18 two_stage_opamp_dummy_magic_0.VD3.t17 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X392 VOUT+.t89 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X393 two_stage_opamp_dummy_magic_0.err_amp_out.t7 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 GNDA.t74 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X394 bgr_0.V_p_2.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 bgr_0.V_mir2.t3 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X395 VOUT-.t87 two_stage_opamp_dummy_magic_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X396 VOUT+.t90 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X397 bgr_0.1st_Vout_2.t22 bgr_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X398 two_stage_opamp_dummy_magic_0.VD4.t35 two_stage_opamp_dummy_magic_0.Vb3.t15 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X399 two_stage_opamp_dummy_magic_0.VD1.t11 two_stage_opamp_dummy_magic_0.Vb1.t14 two_stage_opamp_dummy_magic_0.Y.t16 GNDA.t203 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X400 VDDA.t34 two_stage_opamp_dummy_magic_0.V_err_gate.t24 two_stage_opamp_dummy_magic_0.V_err_p.t10 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X401 two_stage_opamp_dummy_magic_0.VD4.t11 two_stage_opamp_dummy_magic_0.Vb2.t21 two_stage_opamp_dummy_magic_0.Y.t23 two_stage_opamp_dummy_magic_0.VD4.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X402 two_stage_opamp_dummy_magic_0.VD1.t10 two_stage_opamp_dummy_magic_0.Vb1.t15 two_stage_opamp_dummy_magic_0.Y.t0 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X403 VOUT-.t88 two_stage_opamp_dummy_magic_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 VOUT-.t89 two_stage_opamp_dummy_magic_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X405 VOUT-.t90 two_stage_opamp_dummy_magic_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 GNDA.t285 GNDA.t282 GNDA.t284 GNDA.t283 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X407 two_stage_opamp_dummy_magic_0.err_amp_out.t2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 two_stage_opamp_dummy_magic_0.V_err_p.t3 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X408 GNDA.t234 VDDA.t370 VDDA.t372 VDDA.t371 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X409 VDDA.t100 two_stage_opamp_dummy_magic_0.Vb3.t16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=0.64 pd=3.6 as=0.64 ps=3.6 w=3.2 l=0.2
X410 VOUT-.t91 two_stage_opamp_dummy_magic_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 two_stage_opamp_dummy_magic_0.V_p.t20 VIN-.t5 two_stage_opamp_dummy_magic_0.VD1.t5 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X412 bgr_0.1st_Vout_1.t10 bgr_0.V_mir1.t20 VDDA.t461 VDDA.t460 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X413 GNDA.t232 VDDA.t469 bgr_0.V_TOP.t2 GNDA.t223 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X414 VOUT+.t91 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X415 VOUT+.t92 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 VOUT+.t93 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 bgr_0.1st_Vout_2.t5 bgr_0.V_mir2.t19 VDDA.t114 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X418 VDDA.t240 two_stage_opamp_dummy_magic_0.V_err_gate.t25 two_stage_opamp_dummy_magic_0.V_err_p.t9 VDDA.t239 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X419 VDDA.t369 VDDA.t367 GNDA.t233 VDDA.t368 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X420 VOUT+.t94 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 VOUT+.t95 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X422 bgr_0.1st_Vout_2.t23 bgr_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 GNDA.t20 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 two_stage_opamp_dummy_magic_0.err_amp_out.t6 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X424 VOUT-.t92 two_stage_opamp_dummy_magic_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X425 VOUT+.t1 a_14240_2946.t0 GNDA.t86 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X426 bgr_0.1st_Vout_2.t24 bgr_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 VDDA.t451 bgr_0.PFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 VDDA.t450 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X428 VOUT-.t93 two_stage_opamp_dummy_magic_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X429 bgr_0.1st_Vout_1.t25 bgr_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X430 VOUT+.t96 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 bgr_0.V_TOP.t30 VDDA.t277 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 VOUT-.t94 two_stage_opamp_dummy_magic_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 bgr_0.START_UP.t1 bgr_0.V_TOP.t31 VDDA.t276 VDDA.t275 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X434 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 two_stage_opamp_dummy_magic_0.V_err_gate.t26 VDDA.t238 VDDA.t237 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X435 VOUT-.t95 two_stage_opamp_dummy_magic_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 VOUT+.t97 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 VOUT+.t98 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 two_stage_opamp_dummy_magic_0.V_tot.t9 two_stage_opamp_dummy_magic_0.V_err_gate.t7 VDDA.t117 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X439 two_stage_opamp_dummy_magic_0.VD4.t9 two_stage_opamp_dummy_magic_0.Vb2.t22 two_stage_opamp_dummy_magic_0.Y.t12 two_stage_opamp_dummy_magic_0.VD4.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X440 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 two_stage_opamp_dummy_magic_0.X.t42 GNDA.t23 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X441 VOUT-.t15 VDDA.t364 VDDA.t366 VDDA.t365 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X442 VDDA.t30 GNDA.t279 GNDA.t281 GNDA.t280 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X443 bgr_0.1st_Vout_1.t26 bgr_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X444 bgr_0.V_mir2.t10 bgr_0.V_mir2.t9 VDDA.t106 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X445 VDDA.t54 two_stage_opamp_dummy_magic_0.Vb3.t17 two_stage_opamp_dummy_magic_0.VD4.t34 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X446 VOUT+.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X447 VOUT+.t100 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X448 bgr_0.1st_Vout_2.t25 bgr_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X449 VOUT+.t101 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X450 bgr_0.V_TOP.t8 bgr_0.1st_Vout_1.t27 VDDA.t234 VDDA.t233 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X451 VDDA.t363 VDDA.t361 VOUT+.t5 VDDA.t362 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X452 VOUT-.t96 two_stage_opamp_dummy_magic_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X453 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_0.V_err_gate.t27 VDDA.t38 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X454 VOUT-.t97 two_stage_opamp_dummy_magic_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X455 VOUT-.t98 two_stage_opamp_dummy_magic_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 bgr_0.1st_Vout_1.t28 bgr_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X457 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 GNDA.t277 GNDA.t278 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X458 VOUT+.t2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 GNDA.t109 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X459 GNDA.t243 GNDA.t267 bgr_0.Vbe2.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X460 bgr_0.V_mir2.t8 bgr_0.V_mir2.t7 VDDA.t58 VDDA.t57 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X461 VDDA.t274 bgr_0.V_TOP.t32 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 VDDA.t273 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X462 VOUT-.t99 two_stage_opamp_dummy_magic_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 VOUT-.t100 two_stage_opamp_dummy_magic_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X464 VDDA.t360 VDDA.t358 bgr_0.V_TOP.t9 VDDA.t359 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X465 a_5350_5738.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 GNDA.t210 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X466 VOUT+.t102 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X467 two_stage_opamp_dummy_magic_0.V_err_gate.t1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X468 VOUT-.t101 two_stage_opamp_dummy_magic_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X469 bgr_0.V_TOP.t33 VDDA.t272 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 VDDA.t63 two_stage_opamp_dummy_magic_0.V_err_gate.t28 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X471 VDDA.t15 two_stage_opamp_dummy_magic_0.X.t43 VOUT-.t1 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X472 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 VDDA.t355 VDDA.t357 VDDA.t356 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X473 VDDA.t42 two_stage_opamp_dummy_magic_0.Vb3.t18 two_stage_opamp_dummy_magic_0.VD4.t33 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X474 VOUT+.t103 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X475 VOUT+.t104 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X476 VOUT+.t105 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X477 GNDA.t250 GNDA.t266 bgr_0.Vbe2.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X478 bgr_0.1st_Vout_1.t29 bgr_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X479 two_stage_opamp_dummy_magic_0.Y.t10 two_stage_opamp_dummy_magic_0.Vb2.t23 two_stage_opamp_dummy_magic_0.VD4.t7 two_stage_opamp_dummy_magic_0.VD4.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X480 two_stage_opamp_dummy_magic_0.V_p.t36 VIN+.t6 two_stage_opamp_dummy_magic_0.VD2.t17 GNDA.t220 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X481 bgr_0.V_TOP.t34 VDDA.t271 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 two_stage_opamp_dummy_magic_0.VD3.t9 two_stage_opamp_dummy_magic_0.Vb3.t19 VDDA.t56 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X483 VOUT+.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X484 VOUT+.t4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 GNDA.t193 GNDA.t192 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X485 two_stage_opamp_dummy_magic_0.VD3.t23 two_stage_opamp_dummy_magic_0.Vb2.t24 two_stage_opamp_dummy_magic_0.X.t14 two_stage_opamp_dummy_magic_0.VD3.t22 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X486 VOUT-.t102 two_stage_opamp_dummy_magic_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X487 bgr_0.PFET_GATE_10uA.t4 bgr_0.1st_Vout_2.t26 VDDA.t155 VDDA.t154 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X488 a_13790_17550.t1 bgr_0.V_CUR_REF_REG.t0 GNDA.t29 sky130_fd_pr__res_xhigh_po_0p35 l=6
X489 VOUT-.t103 two_stage_opamp_dummy_magic_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 VDDA.t25 bgr_0.PFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X491 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 two_stage_opamp_dummy_magic_0.Y.t41 GNDA.t128 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X492 VDDA.t270 bgr_0.V_TOP.t35 bgr_0.Vin+.t4 VDDA.t269 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X493 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 VDDA.t352 VDDA.t354 VDDA.t353 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X494 bgr_0.1st_Vout_2.t27 bgr_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X495 VOUT-.t104 two_stage_opamp_dummy_magic_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X496 GNDA.t231 VDDA.t470 bgr_0.V_p_2.t9 GNDA.t138 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X497 VOUT-.t105 two_stage_opamp_dummy_magic_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 VDDA.t248 two_stage_opamp_dummy_magic_0.Vb3.t20 two_stage_opamp_dummy_magic_0.VD4.t32 VDDA.t247 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X499 VDDA.t351 VDDA.t349 two_stage_opamp_dummy_magic_0.Vb2.t6 VDDA.t350 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.06 as=0.126 ps=1.03 w=0.63 l=0.2
X500 bgr_0.V_p_1.t7 bgr_0.Vin-.t10 bgr_0.V_mir1.t15 GNDA.t223 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X501 VOUT-.t106 two_stage_opamp_dummy_magic_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X502 VOUT+.t107 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X503 two_stage_opamp_dummy_magic_0.V_p.t32 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 GNDA.t202 GNDA.t201 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X504 two_stage_opamp_dummy_magic_0.V_p.t1 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 GNDA.t7 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X505 bgr_0.V_TOP.t0 bgr_0.1st_Vout_1.t30 VDDA.t48 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X506 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 two_stage_opamp_dummy_magic_0.X.t44 GNDA.t81 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X507 two_stage_opamp_dummy_magic_0.VD2.t4 two_stage_opamp_dummy_magic_0.Vb1.t16 two_stage_opamp_dummy_magic_0.X.t4 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X508 VDDA.t348 VDDA.t346 GNDA.t230 VDDA.t347 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X509 VOUT+.t108 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 bgr_0.V_TOP.t36 VDDA.t268 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 VOUT+.t109 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X512 GNDA.t252 GNDA.t265 bgr_0.Vbe2.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X513 two_stage_opamp_dummy_magic_0.VD1.t21 VIN-.t6 two_stage_opamp_dummy_magic_0.V_p.t19 GNDA.t352 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X514 bgr_0.1st_Vout_1.t9 bgr_0.V_mir1.t21 VDDA.t445 VDDA.t444 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X515 VOUT-.t107 two_stage_opamp_dummy_magic_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X516 VOUT-.t108 two_stage_opamp_dummy_magic_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X517 VOUT-.t109 two_stage_opamp_dummy_magic_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X518 VOUT-.t110 two_stage_opamp_dummy_magic_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X519 VOUT-.t111 two_stage_opamp_dummy_magic_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X520 VOUT-.t112 two_stage_opamp_dummy_magic_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X521 bgr_0.Vin+.t3 bgr_0.V_TOP.t37 VDDA.t267 VDDA.t266 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X522 two_stage_opamp_dummy_magic_0.VD3.t25 two_stage_opamp_dummy_magic_0.Vb2.t25 two_stage_opamp_dummy_magic_0.X.t16 two_stage_opamp_dummy_magic_0.VD3.t24 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X523 bgr_0.V_mir2.t0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 bgr_0.V_p_2.t2 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X524 bgr_0.1st_Vout_2.t28 bgr_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 GNDA.t91 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 two_stage_opamp_dummy_magic_0.V_p.t14 GNDA.t90 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X526 bgr_0.PFET_GATE_10uA.t8 VDDA.t471 GNDA.t229 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X527 VDDA.t236 two_stage_opamp_dummy_magic_0.Y.t42 VOUT+.t13 VDDA.t235 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X528 two_stage_opamp_dummy_magic_0.VD1.t2 VIN-.t7 two_stage_opamp_dummy_magic_0.V_p.t18 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X529 VOUT+.t110 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X530 bgr_0.1st_Vout_2.t29 bgr_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X531 VOUT-.t113 two_stage_opamp_dummy_magic_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 VOUT-.t114 two_stage_opamp_dummy_magic_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X533 VOUT+.t111 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X534 GNDA.t270 GNDA.t268 bgr_0.NFET_GATE_10uA.t4 GNDA.t269 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X535 VOUT+.t112 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X536 VOUT+.t113 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X537 two_stage_opamp_dummy_magic_0.V_err_gate.t5 bgr_0.NFET_GATE_10uA.t18 GNDA.t178 GNDA.t177 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X538 bgr_0.1st_Vout_1.t7 bgr_0.Vin+.t9 bgr_0.V_p_1.t1 GNDA.t226 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X539 VDDA.t119 two_stage_opamp_dummy_magic_0.Vb3.t21 two_stage_opamp_dummy_magic_0.VD4.t31 VDDA.t118 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X540 VDDA.t232 GNDA.t271 GNDA.t273 GNDA.t272 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X541 two_stage_opamp_dummy_magic_0.Y.t9 two_stage_opamp_dummy_magic_0.Vb2.t26 two_stage_opamp_dummy_magic_0.VD4.t5 two_stage_opamp_dummy_magic_0.VD4.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X542 bgr_0.V_TOP.t12 bgr_0.1st_Vout_1.t31 VDDA.t434 VDDA.t433 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X543 two_stage_opamp_dummy_magic_0.X.t5 two_stage_opamp_dummy_magic_0.Vb1.t17 two_stage_opamp_dummy_magic_0.VD2.t5 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X544 VOUT-.t115 two_stage_opamp_dummy_magic_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X545 VDDA.t85 two_stage_opamp_dummy_magic_0.X.t45 VOUT-.t5 VDDA.t84 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X546 VOUT+.t114 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 VDDA.t345 VDDA.t343 VOUT-.t14 VDDA.t344 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X548 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 bgr_0.PFET_GATE_10uA.t24 VDDA.t174 VDDA.t173 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X549 GNDA.t276 GNDA.t274 VDDA.t222 GNDA.t275 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X550 VOUT-.t116 two_stage_opamp_dummy_magic_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X551 VOUT-.t117 two_stage_opamp_dummy_magic_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X552 bgr_0.Vin-.t6 bgr_0.V_TOP.t38 VDDA.t265 VDDA.t264 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X553 VDDA.t211 bgr_0.PFET_GATE_10uA.t25 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X554 VOUT+.t115 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X555 VOUT-.t118 two_stage_opamp_dummy_magic_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X556 a_13790_17550.t0 GNDA.t30 GNDA.t29 sky130_fd_pr__res_xhigh_po_0p35 l=6
X557 VOUT+.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X558 VOUT+.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X559 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 a_14240_2946.t1 GNDA.t103 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X560 bgr_0.V_TOP.t7 VDDA.t340 VDDA.t342 VDDA.t341 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X561 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 two_stage_opamp_dummy_magic_0.Y.t43 GNDA.t64 VDDA.t46 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X562 VOUT+.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X563 VOUT+.t119 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X564 VOUT-.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X565 GNDA.t264 GNDA.t262 two_stage_opamp_dummy_magic_0.err_amp_out.t11 GNDA.t263 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X566 two_stage_opamp_dummy_magic_0.X.t7 two_stage_opamp_dummy_magic_0.VD3.t10 two_stage_opamp_dummy_magic_0.VD3.t12 two_stage_opamp_dummy_magic_0.VD3.t11 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X567 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 two_stage_opamp_dummy_magic_0.X.t46 VDDA.t140 GNDA.t122 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X568 bgr_0.V_TOP.t39 VDDA.t263 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X569 VOUT+.t120 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 VOUT-.t120 two_stage_opamp_dummy_magic_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X571 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 bgr_0.NFET_GATE_10uA.t19 GNDA.t180 GNDA.t179 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X572 two_stage_opamp_dummy_magic_0.Y.t24 two_stage_opamp_dummy_magic_0.Vb2.t27 two_stage_opamp_dummy_magic_0.VD4.t3 two_stage_opamp_dummy_magic_0.VD4.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X573 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 bgr_0.NFET_GATE_10uA.t20 GNDA.t155 GNDA.t154 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X574 VOUT-.t121 two_stage_opamp_dummy_magic_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X575 GNDA.t190 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 VOUT-.t13 GNDA.t189 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X576 VOUT+.t121 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X577 bgr_0.1st_Vout_1.t32 bgr_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X578 VDDA.t149 bgr_0.V_mir2.t20 bgr_0.1st_Vout_2.t4 VDDA.t148 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X579 two_stage_opamp_dummy_magic_0.Y.t19 two_stage_opamp_dummy_magic_0.Vb1.t18 two_stage_opamp_dummy_magic_0.VD1.t9 GNDA.t217 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X580 VOUT-.t122 two_stage_opamp_dummy_magic_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X581 bgr_0.V_TOP.t40 VDDA.t262 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X582 VDDA.t261 bgr_0.V_TOP.t41 bgr_0.Vin+.t2 VDDA.t260 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X583 two_stage_opamp_dummy_magic_0.VD4.t30 two_stage_opamp_dummy_magic_0.Vb3.t22 VDDA.t60 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X584 VOUT-.t123 two_stage_opamp_dummy_magic_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X585 two_stage_opamp_dummy_magic_0.VD2.t14 two_stage_opamp_dummy_magic_0.Vb1.t19 two_stage_opamp_dummy_magic_0.X.t15 GNDA.t187 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X586 two_stage_opamp_dummy_magic_0.V_p.t10 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 GNDA.t55 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X587 VDDA.t339 VDDA.t337 two_stage_opamp_dummy_magic_0.err_amp_out.t10 VDDA.t338 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X588 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 two_stage_opamp_dummy_magic_0.X.t47 GNDA.t123 VDDA.t141 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X589 bgr_0.V_mir1.t3 bgr_0.V_mir1.t2 VDDA.t186 VDDA.t185 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X590 VDDA.t9 two_stage_opamp_dummy_magic_0.Vb3.t23 two_stage_opamp_dummy_magic_0.VD3.t6 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X591 GNDA.t28 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 VOUT+.t0 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X592 VOUT-.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X593 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 bgr_0.NFET_GATE_10uA.t21 GNDA.t157 GNDA.t156 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X594 GNDA.t250 GNDA.t249 bgr_0.Vbe2.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X595 bgr_0.V_mir2.t4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 bgr_0.V_p_2.t1 GNDA.t72 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X596 bgr_0.PFET_GATE_10uA.t7 VDDA.t334 VDDA.t336 VDDA.t335 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X597 GNDA.t206 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 two_stage_opamp_dummy_magic_0.V_p.t33 GNDA.t205 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X598 VDDA.t52 two_stage_opamp_dummy_magic_0.Y.t44 VOUT+.t12 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X599 a_5230_5738.t0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 GNDA.t2 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X600 GNDA.t261 GNDA.t259 VOUT-.t17 GNDA.t260 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X601 two_stage_opamp_dummy_magic_0.VD2.t12 VIN+.t7 two_stage_opamp_dummy_magic_0.V_p.t26 GNDA.t104 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X602 VOUT+.t122 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X603 VOUT-.t125 two_stage_opamp_dummy_magic_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X604 VOUT+.t123 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X605 VDDA.t333 VDDA.t331 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 VDDA.t332 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X606 two_stage_opamp_dummy_magic_0.V_err_gate.t8 two_stage_opamp_dummy_magic_0.V_tot.t10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 VDDA.t200 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X607 VOUT-.t126 two_stage_opamp_dummy_magic_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X608 bgr_0.V_TOP.t42 VDDA.t259 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X609 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 bgr_0.PFET_GATE_10uA.t26 VDDA.t449 VDDA.t448 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X610 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 VDDA.t328 VDDA.t330 VDDA.t329 sky130_fd_pr__pfet_01v8 ad=0.64 pd=3.6 as=1.28 ps=7.2 w=3.2 l=0.2
X611 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_0.Vb3.t0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 sky130_fd_pr__pfet_01v8 ad=1.44 pd=8 as=0.72 ps=4 w=3.6 l=0.2
X612 VOUT+.t124 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X613 VOUT+.t125 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X614 two_stage_opamp_dummy_magic_0.X.t10 two_stage_opamp_dummy_magic_0.Vb1.t20 two_stage_opamp_dummy_magic_0.VD2.t13 GNDA.t105 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X615 VOUT-.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X616 VOUT-.t128 two_stage_opamp_dummy_magic_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X617 VDDA.t136 two_stage_opamp_dummy_magic_0.X.t48 VOUT-.t8 VDDA.t135 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X618 bgr_0.1st_Vout_2.t3 bgr_0.V_mir2.t21 VDDA.t151 VDDA.t150 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X619 VDDA.t432 two_stage_opamp_dummy_magic_0.Vb3.t24 two_stage_opamp_dummy_magic_0.VD3.t37 VDDA.t431 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X620 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 two_stage_opamp_dummy_magic_0.Y.t45 VDDA.t458 GNDA.t345 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X621 two_stage_opamp_dummy_magic_0.X.t20 two_stage_opamp_dummy_magic_0.Vb2.t28 two_stage_opamp_dummy_magic_0.VD3.t34 two_stage_opamp_dummy_magic_0.VD3.t33 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X622 bgr_0.1st_Vout_2.t30 bgr_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X623 GNDA.t252 GNDA.t251 bgr_0.Vin-.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X624 VOUT+.t126 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X625 GNDA.t148 bgr_0.NFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_0.Vb3.t1 GNDA.t147 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X626 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 two_stage_opamp_dummy_magic_0.Y.t46 GNDA.t188 VDDA.t217 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X627 VOUT+.t127 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X628 VOUT+.t128 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X629 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 two_stage_opamp_dummy_magic_0.Y.t47 GNDA.t134 VDDA.t161 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X630 VOUT-.t129 two_stage_opamp_dummy_magic_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X631 two_stage_opamp_dummy_magic_0.VD4.t29 two_stage_opamp_dummy_magic_0.Vb3.t25 VDDA.t224 VDDA.t223 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X632 VOUT+.t129 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X633 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 bgr_0.V_TOP.t43 VDDA.t258 VDDA.t257 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X634 bgr_0.1st_Vout_2.t31 bgr_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X635 GNDA.t10 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X636 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 two_stage_opamp_dummy_magic_0.X.t49 VDDA.t137 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X637 GNDA.t258 GNDA.t256 VDDA.t241 GNDA.t257 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X638 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 VDDA.t325 VDDA.t327 VDDA.t326 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X639 VOUT-.t130 two_stage_opamp_dummy_magic_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X640 VOUT-.t131 two_stage_opamp_dummy_magic_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X641 two_stage_opamp_dummy_magic_0.Y.t15 two_stage_opamp_dummy_magic_0.Vb1.t21 two_stage_opamp_dummy_magic_0.VD1.t8 GNDA.t153 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X642 VDDA.t72 bgr_0.1st_Vout_2.t32 bgr_0.PFET_GATE_10uA.t2 VDDA.t71 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X643 VDDA.t324 VDDA.t322 two_stage_opamp_dummy_magic_0.Vb1.t5 VDDA.t323 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X644 VOUT+.t130 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X645 two_stage_opamp_dummy_magic_0.Vb1.t4 VDDA.t319 VDDA.t321 VDDA.t320 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X646 VOUT+.t131 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X647 two_stage_opamp_dummy_magic_0.V_err_p.t8 two_stage_opamp_dummy_magic_0.V_err_gate.t29 VDDA.t180 VDDA.t179 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X648 two_stage_opamp_dummy_magic_0.V_p.t31 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 GNDA.t199 GNDA.t198 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X649 two_stage_opamp_dummy_magic_0.V_err_p.t0 two_stage_opamp_dummy_magic_0.V_tot.t11 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 VDDA.t61 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X650 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 two_stage_opamp_dummy_magic_0.X.t50 GNDA.t84 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X651 two_stage_opamp_dummy_magic_0.VD2.t8 VIN+.t8 two_stage_opamp_dummy_magic_0.V_p.t13 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X652 GNDA.t255 GNDA.t253 GNDA.t255 GNDA.t254 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0 ps=0 w=2.5 l=0.15
X653 two_stage_opamp_dummy_magic_0.X.t0 two_stage_opamp_dummy_magic_0.Vb2.t29 two_stage_opamp_dummy_magic_0.VD3.t1 two_stage_opamp_dummy_magic_0.VD3.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X654 GNDA.t248 GNDA.t247 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X655 bgr_0.1st_Vout_2.t33 bgr_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X656 VOUT+.t132 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X657 VOUT+.t133 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X658 bgr_0.1st_Vout_2.t34 bgr_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X659 VOUT+.t134 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X660 two_stage_opamp_dummy_magic_0.VD3.t31 VDDA.t316 VDDA.t318 VDDA.t317 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X661 VOUT-.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X662 bgr_0.V_mir1.t14 bgr_0.Vin-.t11 bgr_0.V_p_1.t6 GNDA.t222 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X663 VDDA.t215 two_stage_opamp_dummy_magic_0.Y.t48 VOUT+.t11 VDDA.t214 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X664 VOUT+.t135 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X665 VOUT+.t136 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X666 two_stage_opamp_dummy_magic_0.VD2.t6 VIN+.t9 two_stage_opamp_dummy_magic_0.V_p.t8 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X667 two_stage_opamp_dummy_magic_0.VD4.t28 two_stage_opamp_dummy_magic_0.Vb3.t26 VDDA.t419 VDDA.t418 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X668 VDDA.t160 two_stage_opamp_dummy_magic_0.Y.t49 VOUT+.t10 VDDA.t159 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X669 VOUT-.t133 two_stage_opamp_dummy_magic_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X670 GNDA.t197 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 two_stage_opamp_dummy_magic_0.V_p.t30 GNDA.t196 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X671 bgr_0.1st_Vout_1.t33 bgr_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X672 a_14520_5738.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 GNDA.t116 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X673 VOUT-.t16 GNDA.t244 GNDA.t246 GNDA.t245 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X674 two_stage_opamp_dummy_magic_0.V_err_gate.t0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X675 two_stage_opamp_dummy_magic_0.X.t24 two_stage_opamp_dummy_magic_0.Vb1.t22 two_stage_opamp_dummy_magic_0.VD2.t21 GNDA.t353 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X676 GNDA.t150 bgr_0.NFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 GNDA.t149 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X677 two_stage_opamp_dummy_magic_0.V_p.t29 two_stage_opamp_dummy_magic_0.Vb1.t2 two_stage_opamp_dummy_magic_0.Vb1.t3 GNDA.t337 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=2.9
X678 VDDA.t256 bgr_0.V_TOP.t44 bgr_0.START_UP.t0 VDDA.t255 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X679 VDDA.t92 two_stage_opamp_dummy_magic_0.X.t51 VOUT-.t6 VDDA.t91 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X680 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 two_stage_opamp_dummy_magic_0.Y.t50 VDDA.t158 GNDA.t133 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X681 VOUT+.t137 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X682 VOUT+.t138 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X683 VOUT+.t139 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X684 VOUT-.t134 two_stage_opamp_dummy_magic_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X685 GNDA.t243 GNDA.t242 bgr_0.Vbe2.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X686 VOUT-.t18 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 GNDA.t341 GNDA.t340 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X687 VOUT-.t135 two_stage_opamp_dummy_magic_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X688 VDDA.t188 two_stage_opamp_dummy_magic_0.V_err_gate.t30 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 VDDA.t187 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X689 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 two_stage_opamp_dummy_magic_0.Y.t51 GNDA.t125 VDDA.t144 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X690 VOUT-.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X691 two_stage_opamp_dummy_magic_0.VD4.t24 two_stage_opamp_dummy_magic_0.VD4.t22 two_stage_opamp_dummy_magic_0.Y.t14 two_stage_opamp_dummy_magic_0.VD4.t23 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X692 GNDA.t102 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 GNDA.t101 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X693 two_stage_opamp_dummy_magic_0.Vb2.t10 two_stage_opamp_dummy_magic_0.Vb2.t9 VDDA.t423 VDDA.t422 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.03 as=0.126 ps=1.03 w=0.63 l=0.2
X694 VDDA.t123 bgr_0.V_mir2.t5 bgr_0.V_mir2.t6 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X695 VDDA.t447 bgr_0.PFET_GATE_10uA.t27 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 VDDA.t446 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X696 VOUT+.t140 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X697 bgr_0.1st_Vout_1.t34 bgr_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X698 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 bgr_0.PFET_GATE_10uA.t28 VDDA.t463 VDDA.t462 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X699 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 two_stage_opamp_dummy_magic_0.X.t52 VDDA.t138 GNDA.t120 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X700 VOUT-.t137 two_stage_opamp_dummy_magic_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X701 bgr_0.V_TOP.t45 VDDA.t254 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X702 bgr_0.1st_Vout_1.t5 bgr_0.V_mir1.t22 VDDA.t172 VDDA.t171 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X703 two_stage_opamp_dummy_magic_0.Y.t2 two_stage_opamp_dummy_magic_0.Vb1.t23 two_stage_opamp_dummy_magic_0.VD1.t7 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X704 VOUT-.t138 two_stage_opamp_dummy_magic_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X705 two_stage_opamp_dummy_magic_0.V_err_p.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t31 VDDA.t21 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X706 two_stage_opamp_dummy_magic_0.VD3.t21 two_stage_opamp_dummy_magic_0.Vb3.t27 VDDA.t197 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X707 VOUT+.t141 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X708 two_stage_opamp_dummy_magic_0.V_err_p.t20 two_stage_opamp_dummy_magic_0.V_tot.t12 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 VDDA.t427 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X709 bgr_0.1st_Vout_1.t35 bgr_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X710 bgr_0.1st_Vout_2.t0 bgr_0.V_CUR_REF_REG.t6 bgr_0.V_p_2.t0 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X711 bgr_0.V_TOP.t46 VDDA.t253 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X712 two_stage_opamp_dummy_magic_0.V_p.t6 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 GNDA.t41 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X713 two_stage_opamp_dummy_magic_0.V_err_p.t1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 two_stage_opamp_dummy_magic_0.err_amp_out.t1 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X714 two_stage_opamp_dummy_magic_0.V_p.t37 GNDA.t239 GNDA.t241 GNDA.t240 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X715 two_stage_opamp_dummy_magic_0.V_p_mir.t1 VIN-.t8 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 GNDA.t213 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X716 two_stage_opamp_dummy_magic_0.VD1.t3 VIN-.t9 two_stage_opamp_dummy_magic_0.V_p.t17 GNDA.t50 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X717 VOUT+.t142 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X718 VOUT-.t139 two_stage_opamp_dummy_magic_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X719 VOUT-.t140 two_stage_opamp_dummy_magic_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X720 VOUT-.t141 two_stage_opamp_dummy_magic_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X721 bgr_0.V_p_1.t10 VDDA.t472 GNDA.t227 GNDA.t226 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X722 bgr_0.1st_Vout_2.t35 bgr_0.cap_res2.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X723 bgr_0.V_mir1.t12 bgr_0.Vin-.t12 bgr_0.V_p_1.t5 GNDA.t221 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X724 VDDA.t315 VDDA.t313 bgr_0.PFET_GATE_10uA.t6 VDDA.t314 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X725 VOUT-.t142 two_stage_opamp_dummy_magic_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X726 VOUT-.t143 two_stage_opamp_dummy_magic_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X727 VDDA.t82 two_stage_opamp_dummy_magic_0.Y.t52 VOUT+.t9 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X728 VOUT+.t143 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X729 two_stage_opamp_dummy_magic_0.VD1.t4 VIN-.t10 two_stage_opamp_dummy_magic_0.V_p.t16 GNDA.t145 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X730 GNDA.t67 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 two_stage_opamp_dummy_magic_0.V_p.t11 GNDA.t66 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X731 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 sky130_fd_pr__pfet_01v8 ad=1.44 pd=8 as=0 ps=0 w=3.6 l=0.2
X732 bgr_0.V_TOP.t47 VDDA.t252 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X733 VDDA.t221 bgr_0.V_mir1.t0 bgr_0.V_mir1.t1 VDDA.t220 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X734 VOUT+.t144 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X735 VOUT+.t145 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X736 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 bgr_0.V_TOP.t48 VDDA.t251 VDDA.t250 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X737 bgr_0.V_TOP.t10 bgr_0.START_UP.t7 bgr_0.Vin-.t3 VDDA.t244 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X738 VOUT-.t144 two_stage_opamp_dummy_magic_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X739 bgr_0.1st_Vout_2.t8 bgr_0.V_CUR_REF_REG.t7 bgr_0.V_p_2.t7 GNDA.t209 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X740 VOUT+.t146 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X741 VDDA.t11 bgr_0.1st_Vout_2.t36 bgr_0.PFET_GATE_10uA.t0 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X742 two_stage_opamp_dummy_magic_0.V_err_gate.t11 VDDA.t310 VDDA.t312 VDDA.t311 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X743 bgr_0.1st_Vout_1.t36 bgr_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X744 two_stage_opamp_dummy_magic_0.V_err_gate.t13 two_stage_opamp_dummy_magic_0.V_tot.t13 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 VDDA.t428 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X745 two_stage_opamp_dummy_magic_0.VD3.t16 two_stage_opamp_dummy_magic_0.Vb3.t28 VDDA.t127 VDDA.t126 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X746 two_stage_opamp_dummy_magic_0.X.t3 two_stage_opamp_dummy_magic_0.Vb1.t24 two_stage_opamp_dummy_magic_0.VD2.t0 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X747 two_stage_opamp_dummy_magic_0.VD3.t5 two_stage_opamp_dummy_magic_0.Vb2.t30 two_stage_opamp_dummy_magic_0.X.t2 two_stage_opamp_dummy_magic_0.VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X748 VOUT+.t147 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X749 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 two_stage_opamp_dummy_magic_0.Y.t53 VDDA.t146 GNDA.t127 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X750 VOUT-.t145 two_stage_opamp_dummy_magic_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X751 VOUT-.t146 two_stage_opamp_dummy_magic_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X752 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 two_stage_opamp_dummy_magic_0.Y.t54 VDDA.t468 GNDA.t355 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X753 VOUT-.t147 two_stage_opamp_dummy_magic_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X754 VOUT+.t148 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X755 VOUT+.t149 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X756 VDDA.t309 VDDA.t307 VDDA.t309 VDDA.t308 sky130_fd_pr__pfet_01v8 ad=0.64 pd=3.6 as=0 ps=0 w=3.2 l=0.2
X757 VOUT-.t148 two_stage_opamp_dummy_magic_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X758 VOUT-.t149 two_stage_opamp_dummy_magic_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X759 VOUT+.t150 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X760 VDDA.t306 VDDA.t304 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 VDDA.t305 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X761 VOUT-.t150 two_stage_opamp_dummy_magic_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X762 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 bgr_0.PFET_GATE_10uA.t29 VDDA.t131 VDDA.t130 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X763 VDDA.t231 two_stage_opamp_dummy_magic_0.V_err_gate.t32 two_stage_opamp_dummy_magic_0.V_err_p.t6 VDDA.t230 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X764 VOUT+.t151 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X765 GNDA.t57 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 two_stage_opamp_dummy_magic_0.err_amp_out.t5 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X766 VDDA.t163 bgr_0.V_mir2.t22 bgr_0.1st_Vout_2.t2 VDDA.t162 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X767 VOUT-.t151 two_stage_opamp_dummy_magic_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X768 VOUT+.t152 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X769 VOUT+.t153 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X770 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 two_stage_opamp_dummy_magic_0.X.t53 VDDA.t139 GNDA.t121 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X771 VOUT-.t152 two_stage_opamp_dummy_magic_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X772 two_stage_opamp_dummy_magic_0.Y.t6 two_stage_opamp_dummy_magic_0.Vb1.t25 two_stage_opamp_dummy_magic_0.VD1.t6 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X773 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 two_stage_opamp_dummy_magic_0.V_err_gate.t33 VDDA.t89 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X774 two_stage_opamp_dummy_magic_0.VD3.t8 two_stage_opamp_dummy_magic_0.Vb2.t31 two_stage_opamp_dummy_magic_0.X.t6 two_stage_opamp_dummy_magic_0.VD3.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X775 VOUT-.t153 two_stage_opamp_dummy_magic_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X776 VOUT-.t154 two_stage_opamp_dummy_magic_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X777 VOUT+.t154 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X778 VOUT+.t155 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X779 two_stage_opamp_dummy_magic_0.V_p_mir.t2 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 GNDA.t37 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X780 two_stage_opamp_dummy_magic_0.V_err_p.t5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 two_stage_opamp_dummy_magic_0.err_amp_out.t0 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X781 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 two_stage_opamp_dummy_magic_0.X.t54 GNDA.t114 VDDA.t134 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X782 VOUT-.t155 two_stage_opamp_dummy_magic_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X783 bgr_0.V_TOP.t49 VDDA.t249 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X784 bgr_0.1st_Vout_1.t0 bgr_0.Vin+.t10 bgr_0.V_p_1.t0 GNDA.t65 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X785 two_stage_opamp_dummy_magic_0.VD2.t18 GNDA.t236 GNDA.t238 GNDA.t237 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X786 VOUT-.t156 two_stage_opamp_dummy_magic_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X787 two_stage_opamp_dummy_magic_0.VD2.t7 VIN+.t10 two_stage_opamp_dummy_magic_0.V_p.t12 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X788 bgr_0.Vin+.t0 bgr_0.Vbe2.t0 GNDA.t70 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X789 VDDA.t303 VDDA.t301 two_stage_opamp_dummy_magic_0.VD4.t0 VDDA.t302 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X790 VOUT+.t156 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 bgr_0.V_TOP.n0 bgr_0.V_TOP.t43 369.534
R1 bgr_0.V_TOP.n11 bgr_0.V_TOP.n9 339.961
R2 bgr_0.V_TOP.n11 bgr_0.V_TOP.n10 339.272
R3 bgr_0.V_TOP.n7 bgr_0.V_TOP.n6 339.272
R4 bgr_0.V_TOP.n15 bgr_0.V_TOP.n14 339.272
R5 bgr_0.V_TOP.n17 bgr_0.V_TOP.n16 339.272
R6 bgr_0.V_TOP.n12 bgr_0.V_TOP.n8 334.772
R7 bgr_0.V_TOP.n27 bgr_0.V_TOP.n26 224.934
R8 bgr_0.V_TOP.n26 bgr_0.V_TOP.n25 224.934
R9 bgr_0.V_TOP.n25 bgr_0.V_TOP.n24 224.934
R10 bgr_0.V_TOP.n24 bgr_0.V_TOP.n23 224.934
R11 bgr_0.V_TOP.n23 bgr_0.V_TOP.n22 224.934
R12 bgr_0.V_TOP.n22 bgr_0.V_TOP.n21 224.934
R13 bgr_0.V_TOP.n21 bgr_0.V_TOP.n20 224.934
R14 bgr_0.V_TOP.n1 bgr_0.V_TOP.n0 224.934
R15 bgr_0.V_TOP.n2 bgr_0.V_TOP.n1 224.934
R16 bgr_0.V_TOP.n3 bgr_0.V_TOP.n2 224.934
R17 bgr_0.V_TOP.n4 bgr_0.V_TOP.n3 224.934
R18 bgr_0.V_TOP.n5 bgr_0.V_TOP.n4 224.934
R19 bgr_0.V_TOP bgr_0.V_TOP.t32 214.222
R20 bgr_0.V_TOP bgr_0.V_TOP.n40 205.502
R21 bgr_0.V_TOP.n7 bgr_0.V_TOP.t4 176.114
R22 bgr_0.V_TOP.n19 bgr_0.V_TOP.n18 163.175
R23 bgr_0.V_TOP.n27 bgr_0.V_TOP.t31 144.601
R24 bgr_0.V_TOP.n26 bgr_0.V_TOP.t44 144.601
R25 bgr_0.V_TOP.n25 bgr_0.V_TOP.t18 144.601
R26 bgr_0.V_TOP.n24 bgr_0.V_TOP.t26 144.601
R27 bgr_0.V_TOP.n23 bgr_0.V_TOP.t37 144.601
R28 bgr_0.V_TOP.n22 bgr_0.V_TOP.t35 144.601
R29 bgr_0.V_TOP.n21 bgr_0.V_TOP.t48 144.601
R30 bgr_0.V_TOP.n20 bgr_0.V_TOP.t20 144.601
R31 bgr_0.V_TOP.n0 bgr_0.V_TOP.t29 144.601
R32 bgr_0.V_TOP.n1 bgr_0.V_TOP.t23 144.601
R33 bgr_0.V_TOP.n2 bgr_0.V_TOP.t14 144.601
R34 bgr_0.V_TOP.n3 bgr_0.V_TOP.t38 144.601
R35 bgr_0.V_TOP.n4 bgr_0.V_TOP.t41 144.601
R36 bgr_0.V_TOP.n5 bgr_0.V_TOP.t27 144.601
R37 bgr_0.V_TOP.n18 bgr_0.V_TOP.t2 95.4466
R38 bgr_0.V_TOP bgr_0.V_TOP.n27 69.6227
R39 bgr_0.V_TOP.n20 bgr_0.V_TOP.n19 69.6227
R40 bgr_0.V_TOP.n19 bgr_0.V_TOP.n5 69.6227
R41 bgr_0.V_TOP.n6 bgr_0.V_TOP.t1 39.4005
R42 bgr_0.V_TOP.n6 bgr_0.V_TOP.t0 39.4005
R43 bgr_0.V_TOP.n8 bgr_0.V_TOP.t5 39.4005
R44 bgr_0.V_TOP.n8 bgr_0.V_TOP.t12 39.4005
R45 bgr_0.V_TOP.n10 bgr_0.V_TOP.t3 39.4005
R46 bgr_0.V_TOP.n10 bgr_0.V_TOP.t13 39.4005
R47 bgr_0.V_TOP.n9 bgr_0.V_TOP.t9 39.4005
R48 bgr_0.V_TOP.n9 bgr_0.V_TOP.t10 39.4005
R49 bgr_0.V_TOP.n14 bgr_0.V_TOP.t11 39.4005
R50 bgr_0.V_TOP.n14 bgr_0.V_TOP.t8 39.4005
R51 bgr_0.V_TOP.n16 bgr_0.V_TOP.t6 39.4005
R52 bgr_0.V_TOP.n16 bgr_0.V_TOP.t7 39.4005
R53 bgr_0.V_TOP.n12 bgr_0.V_TOP.n11 8.313
R54 bgr_0.V_TOP.n18 bgr_0.V_TOP.n17 5.188
R55 bgr_0.V_TOP.n28 bgr_0.V_TOP.t49 4.8295
R56 bgr_0.V_TOP.n29 bgr_0.V_TOP.t25 4.8295
R57 bgr_0.V_TOP.n31 bgr_0.V_TOP.t21 4.8295
R58 bgr_0.V_TOP.n32 bgr_0.V_TOP.t34 4.8295
R59 bgr_0.V_TOP.n34 bgr_0.V_TOP.t30 4.8295
R60 bgr_0.V_TOP.n35 bgr_0.V_TOP.t46 4.8295
R61 bgr_0.V_TOP.n37 bgr_0.V_TOP.t24 4.8295
R62 bgr_0.V_TOP.n28 bgr_0.V_TOP.t39 4.5005
R63 bgr_0.V_TOP.n30 bgr_0.V_TOP.t28 4.5005
R64 bgr_0.V_TOP.n29 bgr_0.V_TOP.t33 4.5005
R65 bgr_0.V_TOP.n31 bgr_0.V_TOP.t15 4.5005
R66 bgr_0.V_TOP.n33 bgr_0.V_TOP.t40 4.5005
R67 bgr_0.V_TOP.n32 bgr_0.V_TOP.t45 4.5005
R68 bgr_0.V_TOP.n34 bgr_0.V_TOP.t22 4.5005
R69 bgr_0.V_TOP.n36 bgr_0.V_TOP.t16 4.5005
R70 bgr_0.V_TOP.n35 bgr_0.V_TOP.t19 4.5005
R71 bgr_0.V_TOP.n37 bgr_0.V_TOP.t17 4.5005
R72 bgr_0.V_TOP.n38 bgr_0.V_TOP.t42 4.5005
R73 bgr_0.V_TOP.n39 bgr_0.V_TOP.t47 4.5005
R74 bgr_0.V_TOP.n40 bgr_0.V_TOP.t36 4.5005
R75 bgr_0.V_TOP.n13 bgr_0.V_TOP.n12 4.5005
R76 bgr_0.V_TOP.n17 bgr_0.V_TOP.n15 2.1255
R77 bgr_0.V_TOP.n15 bgr_0.V_TOP.n13 2.1255
R78 bgr_0.V_TOP.n13 bgr_0.V_TOP.n7 2.1255
R79 bgr_0.V_TOP.n30 bgr_0.V_TOP.n28 0.3295
R80 bgr_0.V_TOP.n30 bgr_0.V_TOP.n29 0.3295
R81 bgr_0.V_TOP.n33 bgr_0.V_TOP.n31 0.3295
R82 bgr_0.V_TOP.n33 bgr_0.V_TOP.n32 0.3295
R83 bgr_0.V_TOP.n36 bgr_0.V_TOP.n34 0.3295
R84 bgr_0.V_TOP.n36 bgr_0.V_TOP.n35 0.3295
R85 bgr_0.V_TOP.n38 bgr_0.V_TOP.n37 0.3295
R86 bgr_0.V_TOP.n39 bgr_0.V_TOP.n38 0.3295
R87 bgr_0.V_TOP.n40 bgr_0.V_TOP.n39 0.3295
R88 bgr_0.V_TOP.n33 bgr_0.V_TOP.n30 0.2825
R89 bgr_0.V_TOP.n36 bgr_0.V_TOP.n33 0.2825
R90 bgr_0.V_TOP.n38 bgr_0.V_TOP.n36 0.2825
R91 bgr_0.Vin-.n14 bgr_0.Vin-.t10 688.859
R92 bgr_0.Vin-.n16 bgr_0.Vin-.n15 514.134
R93 bgr_0.Vin-.n12 bgr_0.Vin-.n11 345.115
R94 bgr_0.Vin-.n18 bgr_0.Vin-.n17 214.713
R95 bgr_0.Vin-.n14 bgr_0.Vin-.t12 174.726
R96 bgr_0.Vin-.n15 bgr_0.Vin-.t8 174.726
R97 bgr_0.Vin-.n16 bgr_0.Vin-.t11 174.726
R98 bgr_0.Vin-.n17 bgr_0.Vin-.t9 174.726
R99 bgr_0.Vin-.n10 bgr_0.Vin-.n8 173.029
R100 bgr_0.Vin-.n10 bgr_0.Vin-.n9 168.654
R101 bgr_0.Vin-.n12 bgr_0.Vin-.t0 162.921
R102 bgr_0.Vin-.n15 bgr_0.Vin-.n14 128.534
R103 bgr_0.Vin-.n17 bgr_0.Vin-.n16 128.534
R104 bgr_0.Vin-.n5 bgr_0.Vin-.n4 83.5719
R105 bgr_0.Vin-.n3 bgr_0.Vin-.n0 83.5719
R106 bgr_0.Vin-.n3 bgr_0.Vin-.n1 73.3165
R107 bgr_0.Vin-.t2 bgr_0.Vin-.n2 65.0341
R108 bgr_0.Vin-.n11 bgr_0.Vin-.t3 39.4005
R109 bgr_0.Vin-.n11 bgr_0.Vin-.t1 39.4005
R110 bgr_0.Vin-.n4 bgr_0.Vin-.n3 26.074
R111 bgr_0.Vin-.n19 bgr_0.Vin-.n18 17.526
R112 bgr_0.Vin-.n9 bgr_0.Vin-.t7 13.1338
R113 bgr_0.Vin-.n9 bgr_0.Vin-.t6 13.1338
R114 bgr_0.Vin-.n8 bgr_0.Vin-.t4 13.1338
R115 bgr_0.Vin-.n8 bgr_0.Vin-.t5 13.1338
R116 bgr_0.Vin-.n18 bgr_0.Vin-.n13 12.5317
R117 bgr_0.Vin-.n13 bgr_0.Vin-.n12 6.40675
R118 bgr_0.Vin-.n13 bgr_0.Vin-.n10 3.8755
R119 bgr_0.Vin-.n19 bgr_0.Vin-.n1 2.19742
R120 bgr_0.Vin-.n5 bgr_0.Vin-.n2 1.56483
R121 bgr_0.Vin-.n21 bgr_0.Vin-.n20 1.5505
R122 bgr_0.Vin-.n7 bgr_0.Vin-.n6 1.5505
R123 bgr_0.Vin-.n21 bgr_0.Vin-.n1 1.19225
R124 bgr_0.Vin-.n6 bgr_0.Vin-.n0 0.885803
R125 bgr_0.Vin-.n6 bgr_0.Vin-.n5 0.77514
R126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter bgr_0.Vin-.n0 0.756696
R127 bgr_0.Vin-.n7 bgr_0.Vin-.n2 0.539177
R128 bgr_0.Vin-.n4 bgr_0.Vin-.t2 0.290206
R129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter bgr_0.Vin-.n21 0.203382
R130 bgr_0.Vin-.n20 bgr_0.Vin-.n7 0.0183571
R131 bgr_0.Vin-.n20 bgr_0.Vin-.n19 0.0183571
R132 VDDA.n376 VDDA.n343 6600
R133 VDDA.n378 VDDA.n343 6600
R134 VDDA.n378 VDDA.n344 6570
R135 VDDA.n376 VDDA.n344 6570
R136 VDDA.n331 VDDA.n266 4710
R137 VDDA.n331 VDDA.n267 4710
R138 VDDA.n333 VDDA.n266 4710
R139 VDDA.n333 VDDA.n267 4710
R140 VDDA.n289 VDDA.n288 4710
R141 VDDA.n291 VDDA.n288 4710
R142 VDDA.n289 VDDA.n282 4710
R143 VDDA.n291 VDDA.n282 4710
R144 VDDA.n141 VDDA.n137 4605
R145 VDDA.n141 VDDA.n138 4605
R146 VDDA.n42 VDDA.n28 4605
R147 VDDA.n44 VDDA.n28 4605
R148 VDDA.n206 VDDA.n182 4590
R149 VDDA.n208 VDDA.n182 4590
R150 VDDA.n208 VDDA.n183 4590
R151 VDDA.n206 VDDA.n183 4590
R152 VDDA.n143 VDDA.n137 4575
R153 VDDA.n143 VDDA.n138 4575
R154 VDDA.n42 VDDA.n29 4575
R155 VDDA.n44 VDDA.n29 4575
R156 VDDA.n101 VDDA.n94 4020
R157 VDDA.n103 VDDA.n94 4020
R158 VDDA.n101 VDDA.n100 4020
R159 VDDA.n103 VDDA.n100 4020
R160 VDDA.n77 VDDA.n70 4020
R161 VDDA.n79 VDDA.n70 4020
R162 VDDA.n77 VDDA.n76 4020
R163 VDDA.n79 VDDA.n76 4020
R164 VDDA.n442 VDDA.n410 3420
R165 VDDA.n442 VDDA.n411 3420
R166 VDDA.n121 VDDA.n114 3390
R167 VDDA.n123 VDDA.n114 3390
R168 VDDA.n121 VDDA.n120 3390
R169 VDDA.n123 VDDA.n120 3390
R170 VDDA.n21 VDDA.n14 3390
R171 VDDA.n23 VDDA.n14 3390
R172 VDDA.n21 VDDA.n20 3390
R173 VDDA.n23 VDDA.n20 3390
R174 VDDA.n163 VDDA.n157 2940
R175 VDDA.n165 VDDA.n157 2940
R176 VDDA.n165 VDDA.n162 2940
R177 VDDA.n163 VDDA.n162 2940
R178 VDDA.n171 VDDA.n152 2940
R179 VDDA.n173 VDDA.n152 2940
R180 VDDA.n173 VDDA.n170 2940
R181 VDDA.n171 VDDA.n170 2940
R182 VDDA.n444 VDDA.n410 2760
R183 VDDA.n444 VDDA.n411 2760
R184 VDDA.n235 VDDA.n224 2415
R185 VDDA.n235 VDDA.n225 2370
R186 VDDA.n232 VDDA.n225 2280
R187 VDDA.n232 VDDA.n224 2235
R188 VDDA.n458 VDDA.n404 2145
R189 VDDA.n458 VDDA.n405 2100
R190 VDDA.n455 VDDA.n405 2100
R191 VDDA.n423 VDDA.n416 2100
R192 VDDA.n425 VDDA.n416 2100
R193 VDDA.n425 VDDA.n417 2100
R194 VDDA.n423 VDDA.n417 2100
R195 VDDA.n455 VDDA.n404 2055
R196 VDDA.n391 VDDA.n389 1770
R197 VDDA.n393 VDDA.n389 1770
R198 VDDA.n391 VDDA.n386 1770
R199 VDDA.n393 VDDA.n386 1770
R200 VDDA.n352 VDDA.n350 1770
R201 VDDA.n354 VDDA.n350 1770
R202 VDDA.n352 VDDA.n347 1770
R203 VDDA.n354 VDDA.n347 1770
R204 VDDA.n247 VDDA.n220 1575
R205 VDDA.n246 VDDA.n220 1575
R206 VDDA.n246 VDDA.n219 1545
R207 VDDA.n247 VDDA.n219 1545
R208 VDDA.n135 VDDA.t364 1216.42
R209 VDDA.n146 VDDA.t343 1216.42
R210 VDDA.n39 VDDA.t361 1216.42
R211 VDDA.n47 VDDA.t373 1216.42
R212 VDDA.n375 VDDA.n342 704
R213 VDDA.n379 VDDA.n342 704
R214 VDDA.n159 VDDA.t339 689.4
R215 VDDA.n158 VDDA.t357 689.4
R216 VDDA.n154 VDDA.t415 689.4
R217 VDDA.n153 VDDA.t312 689.4
R218 VDDA.n202 VDDA.t397 663.801
R219 VDDA.n212 VDDA.t391 663.801
R220 VDDA.n97 VDDA.t404 660.109
R221 VDDA.n95 VDDA.t316 660.109
R222 VDDA.n73 VDDA.t301 660.109
R223 VDDA.n71 VDDA.t383 660.109
R224 VDDA.n242 VDDA.t351 647.54
R225 VDDA.n251 VDDA.t379 647.54
R226 VDDA.n216 VDDA.n215 633.361
R227 VDDA.n179 VDDA.n178 626.534
R228 VDDA.n185 VDDA.n184 626.534
R229 VDDA.n187 VDDA.n186 626.534
R230 VDDA.n189 VDDA.n188 626.534
R231 VDDA.n191 VDDA.n190 626.534
R232 VDDA.n193 VDDA.n192 626.534
R233 VDDA.n195 VDDA.n194 626.534
R234 VDDA.n197 VDDA.n196 626.534
R235 VDDA.n199 VDDA.n198 626.534
R236 VDDA.n201 VDDA.n200 626.534
R237 VDDA.n229 VDDA.t307 623.958
R238 VDDA.n238 VDDA.t328 623.958
R239 VDDA.t307 VDDA.n228 615.926
R240 VDDA.n117 VDDA.t346 573.75
R241 VDDA.n115 VDDA.t370 573.75
R242 VDDA.n17 VDDA.t367 573.75
R243 VDDA.n15 VDDA.t380 573.75
R244 VDDA.n374 VDDA.n341 518.4
R245 VDDA.n380 VDDA.n341 518.4
R246 VDDA.n293 VDDA.n292 496
R247 VDDA.n293 VDDA.n281 496
R248 VDDA.n140 VDDA.n112 491.2
R249 VDDA.n140 VDDA.n139 491.2
R250 VDDA.n45 VDDA.n27 491.2
R251 VDDA.n41 VDDA.n27 491.2
R252 VDDA.n205 VDDA.n181 489.601
R253 VDDA.n209 VDDA.n181 489.601
R254 VDDA.n105 VDDA.n104 428.8
R255 VDDA.n105 VDDA.n93 428.8
R256 VDDA.n81 VDDA.n80 428.8
R257 VDDA.n81 VDDA.n69 428.8
R258 VDDA.n387 VDDA.t319 419.108
R259 VDDA.n384 VDDA.t322 419.108
R260 VDDA.n348 VDDA.t398 413.084
R261 VDDA.n345 VDDA.t358 413.084
R262 VDDA.n452 VDDA.t386 409.067
R263 VDDA.n461 VDDA.t325 409.067
R264 VDDA.n439 VDDA.t407 409.067
R265 VDDA.n447 VDDA.t401 409.067
R266 VDDA.n420 VDDA.t304 409.067
R267 VDDA.n428 VDDA.t352 390.322
R268 VDDA.t396 VDDA.n206 389.375
R269 VDDA.n208 VDDA.t390 389.375
R270 VDDA.t414 VDDA.n170 389.375
R271 VDDA.t311 VDDA.n152 389.375
R272 VDDA.n387 VDDA.t321 389.185
R273 VDDA.n384 VDDA.t324 389.185
R274 VDDA.n204 VDDA.n180 387.2
R275 VDDA.n210 VDDA.n180 387.2
R276 VDDA.n439 VDDA.t409 387.051
R277 VDDA.n447 VDDA.t403 387.051
R278 VDDA.n264 VDDA.t336 384.918
R279 VDDA.n268 VDDA.t315 384.918
R280 VDDA.n283 VDDA.t342 384.918
R281 VDDA.n285 VDDA.t412 384.918
R282 VDDA.n348 VDDA.t400 384.918
R283 VDDA.n345 VDDA.t360 384.918
R284 VDDA.t338 VDDA.n162 384.168
R285 VDDA.t356 VDDA.n157 384.168
R286 VDDA.n270 VDDA.n269 384
R287 VDDA.n269 VDDA.n265 384
R288 VDDA.n287 VDDA.n286 384
R289 VDDA.n287 VDDA.n284 384
R290 VDDA.n420 VDDA.t306 370.728
R291 VDDA.n428 VDDA.t354 370.728
R292 VDDA.n452 VDDA.t388 370.3
R293 VDDA.n461 VDDA.t327 370.3
R294 VDDA.n441 VDDA.n409 364.8
R295 VDDA.n373 VDDA.t331 360.868
R296 VDDA.n381 VDDA.t392 360.868
R297 VDDA.n264 VDDA.t334 358.858
R298 VDDA.n268 VDDA.t313 358.858
R299 VDDA.n283 VDDA.t340 358.858
R300 VDDA.n285 VDDA.t410 358.858
R301 VDDA.n125 VDDA.n124 355.2
R302 VDDA.n125 VDDA.n113 355.2
R303 VDDA.n25 VDDA.n24 355.2
R304 VDDA.n25 VDDA.n13 355.2
R305 VDDA.t314 VDDA.n331 351.591
R306 VDDA.n333 VDDA.t335 351.591
R307 VDDA.t411 VDDA.n289 351.591
R308 VDDA.n291 VDDA.t341 351.591
R309 VDDA.t350 VDDA.n246 346.668
R310 VDDA.n247 VDDA.t377 346.668
R311 VDDA.n413 VDDA.n412 345.127
R312 VDDA.n419 VDDA.n418 345.127
R313 VDDA.n401 VDDA.n400 344.7
R314 VDDA.n450 VDDA.n449 344.7
R315 VDDA.t323 VDDA.n391 344.394
R316 VDDA.n393 VDDA.t320 344.394
R317 VDDA.t359 VDDA.n352 344.394
R318 VDDA.n354 VDDA.t399 344.394
R319 VDDA.t387 VDDA.n455 344.394
R320 VDDA.n458 VDDA.t326 344.394
R321 VDDA.n275 VDDA.n273 342.3
R322 VDDA.n303 VDDA.n302 341.675
R323 VDDA.n301 VDDA.n300 341.675
R324 VDDA.n299 VDDA.n298 341.675
R325 VDDA.n297 VDDA.n296 341.675
R326 VDDA.n279 VDDA.n278 341.675
R327 VDDA.n277 VDDA.n276 341.675
R328 VDDA.n275 VDDA.n274 341.675
R329 VDDA.t408 VDDA.n442 340.635
R330 VDDA.n444 VDDA.t402 340.635
R331 VDDA.t305 VDDA.n423 340.635
R332 VDDA.n425 VDDA.t353 340.635
R333 VDDA.n407 VDDA.n406 339.272
R334 VDDA.n431 VDDA.n430 339.272
R335 VDDA.n433 VDDA.n432 339.272
R336 VDDA.n435 VDDA.n434 339.272
R337 VDDA.n437 VDDA.n436 339.272
R338 VDDA.n336 VDDA.n260 337.175
R339 VDDA.n262 VDDA.n261 337.175
R340 VDDA.n312 VDDA.n311 337.175
R341 VDDA.n315 VDDA.n309 337.175
R342 VDDA.n307 VDDA.n306 337.175
R343 VDDA.n319 VDDA.n318 337.175
R344 VDDA.n322 VDDA.n305 337.175
R345 VDDA.n325 VDDA.n324 337.175
R346 VDDA.n328 VDDA.n272 337.175
R347 VDDA.n294 VDDA.n280 337.175
R348 VDDA.n397 VDDA.n383 335.022
R349 VDDA.n203 VDDA.t395 332.75
R350 VDDA.n211 VDDA.t389 332.75
R351 VDDA.n159 VDDA.t337 332.75
R352 VDDA.n158 VDDA.t355 332.75
R353 VDDA.n154 VDDA.t413 332.75
R354 VDDA.n153 VDDA.t310 332.75
R355 VDDA.n243 VDDA.t349 314.274
R356 VDDA.n250 VDDA.t376 314.274
R357 VDDA.n161 VDDA.n156 313.601
R358 VDDA.n168 VDDA.n156 307.2
R359 VDDA.n176 VDDA.n151 307.2
R360 VDDA.n169 VDDA.n151 307.2
R361 VDDA.n445 VDDA.n409 294.401
R362 VDDA.t347 VDDA.n121 285.815
R363 VDDA.n123 VDDA.t371 285.815
R364 VDDA.t368 VDDA.n21 285.815
R365 VDDA.n23 VDDA.t381 285.815
R366 VDDA.t332 VDDA.n376 278.95
R367 VDDA.n378 VDDA.t393 278.95
R368 VDDA.n117 VDDA.t348 277.916
R369 VDDA.n115 VDDA.t372 277.916
R370 VDDA.n17 VDDA.t369 277.916
R371 VDDA.n15 VDDA.t382 277.916
R372 VDDA.n145 VDDA.n112 276.8
R373 VDDA.n139 VDDA.n136 276.8
R374 VDDA.n46 VDDA.n45 276.8
R375 VDDA.n41 VDDA.n40 276.8
R376 VDDA.n373 VDDA.t333 270.705
R377 VDDA.n381 VDDA.t394 270.705
R378 VDDA.n236 VDDA.n223 257.601
R379 VDDA.n440 VDDA.n408 246.4
R380 VDDA.t405 VDDA.n101 239.915
R381 VDDA.n103 VDDA.t317 239.915
R382 VDDA.t302 VDDA.n77 239.915
R383 VDDA.n79 VDDA.t384 239.915
R384 VDDA.n231 VDDA.n223 238.4
R385 VDDA.n99 VDDA.n98 230.4
R386 VDDA.n99 VDDA.n96 230.4
R387 VDDA.n75 VDDA.n74 230.4
R388 VDDA.n75 VDDA.n72 230.4
R389 VDDA.n459 VDDA.n403 228.8
R390 VDDA.n422 VDDA.n415 224
R391 VDDA.n426 VDDA.n415 224
R392 VDDA.n454 VDDA.n403 219.201
R393 VDDA.n166 VDDA.n160 211.201
R394 VDDA.n167 VDDA.n166 211.201
R395 VDDA.n175 VDDA.n174 211.201
R396 VDDA.n119 VDDA.n118 211.201
R397 VDDA.n119 VDDA.n116 211.201
R398 VDDA.n19 VDDA.n18 211.201
R399 VDDA.n19 VDDA.n16 211.201
R400 VDDA.n145 VDDA.n144 204.8
R401 VDDA.n144 VDDA.n136 204.8
R402 VDDA.n40 VDDA.n26 204.8
R403 VDDA.n46 VDDA.n26 204.8
R404 VDDA.n174 VDDA.n155 202.971
R405 VDDA.n104 VDDA.n96 198.4
R406 VDDA.n98 VDDA.n93 198.4
R407 VDDA.n80 VDDA.n72 198.4
R408 VDDA.n74 VDDA.n69 198.4
R409 VDDA.n231 VDDA.n230 192
R410 VDDA.t422 VDDA.t350 190
R411 VDDA.t377 VDDA.t422 190
R412 VDDA.n237 VDDA.n236 188.8
R413 VDDA.n335 VDDA.n334 188.8
R414 VDDA.n330 VDDA.n329 188.8
R415 VDDA.n394 VDDA.n388 188.8
R416 VDDA.n390 VDDA.n388 188.8
R417 VDDA.n355 VDDA.n349 188.8
R418 VDDA.n351 VDDA.n349 188.8
R419 VDDA.t179 VDDA.t396 186.607
R420 VDDA.t115 VDDA.t179 186.607
R421 VDDA.t237 VDDA.t115 186.607
R422 VDDA.t49 VDDA.t237 186.607
R423 VDDA.t20 VDDA.t49 186.607
R424 VDDA.t64 VDDA.t20 186.607
R425 VDDA.t88 VDDA.t64 186.607
R426 VDDA.t33 VDDA.t88 186.607
R427 VDDA.t442 VDDA.t33 186.607
R428 VDDA.t62 VDDA.t442 186.607
R429 VDDA.t239 VDDA.t191 186.607
R430 VDDA.t39 VDDA.t239 186.607
R431 VDDA.t187 VDDA.t39 186.607
R432 VDDA.t439 VDDA.t187 186.607
R433 VDDA.t230 VDDA.t439 186.607
R434 VDDA.t4 VDDA.t230 186.607
R435 VDDA.t189 VDDA.t4 186.607
R436 VDDA.t37 VDDA.t189 186.607
R437 VDDA.t66 VDDA.t37 186.607
R438 VDDA.t390 VDDA.t66 186.607
R439 VDDA.t6 VDDA.t414 186.607
R440 VDDA.t209 VDDA.t6 186.607
R441 VDDA.t428 VDDA.t209 186.607
R442 VDDA.t12 VDDA.t428 186.607
R443 VDDA.t36 VDDA.t12 186.607
R444 VDDA.t117 VDDA.t200 186.607
R445 VDDA.t200 VDDA.t198 186.607
R446 VDDA.t198 VDDA.t68 186.607
R447 VDDA.t68 VDDA.t229 186.607
R448 VDDA.t229 VDDA.t311 186.607
R449 VDDA.t7 VDDA.t338 183.333
R450 VDDA.t61 VDDA.t7 183.333
R451 VDDA.t426 VDDA.t61 183.333
R452 VDDA.t31 VDDA.t426 183.333
R453 VDDA.t199 VDDA.t31 183.333
R454 VDDA.t427 VDDA.t441 183.333
R455 VDDA.t441 VDDA.t32 183.333
R456 VDDA.t32 VDDA.t35 183.333
R457 VDDA.t35 VDDA.t228 183.333
R458 VDDA.t228 VDDA.t356 183.333
R459 VDDA.n375 VDDA.n374 182.4
R460 VDDA.n380 VDDA.n379 182.4
R461 VDDA.n134 VDDA.t366 178.124
R462 VDDA.n147 VDDA.t345 178.124
R463 VDDA.n38 VDDA.t363 178.124
R464 VDDA.n48 VDDA.t375 178.124
R465 VDDA.n446 VDDA.n408 176
R466 VDDA.n226 VDDA.n221 174.393
R467 VDDA.t245 VDDA.t314 172.727
R468 VDDA.t148 VDDA.t245 172.727
R469 VDDA.t111 VDDA.t148 172.727
R470 VDDA.t122 VDDA.t111 172.727
R471 VDDA.t105 VDDA.t122 172.727
R472 VDDA.t71 VDDA.t105 172.727
R473 VDDA.t424 VDDA.t71 172.727
R474 VDDA.t162 VDDA.t424 172.727
R475 VDDA.t113 VDDA.t162 172.727
R476 VDDA.t464 VDDA.t203 172.727
R477 VDDA.t10 VDDA.t464 172.727
R478 VDDA.t154 VDDA.t10 172.727
R479 VDDA.t96 VDDA.t154 172.727
R480 VDDA.t150 VDDA.t96 172.727
R481 VDDA.t456 VDDA.t150 172.727
R482 VDDA.t57 VDDA.t456 172.727
R483 VDDA.t28 VDDA.t57 172.727
R484 VDDA.t335 VDDA.t28 172.727
R485 VDDA.t47 VDDA.t411 172.727
R486 VDDA.t0 VDDA.t47 172.727
R487 VDDA.t435 VDDA.t0 172.727
R488 VDDA.t437 VDDA.t435 172.727
R489 VDDA.t460 VDDA.t437 172.727
R490 VDDA.t205 VDDA.t460 172.727
R491 VDDA.t433 VDDA.t205 172.727
R492 VDDA.t220 VDDA.t433 172.727
R493 VDDA.t73 VDDA.t220 172.727
R494 VDDA.t444 VDDA.t128 172.727
R495 VDDA.t416 VDDA.t444 172.727
R496 VDDA.t233 VDDA.t416 172.727
R497 VDDA.t22 VDDA.t233 172.727
R498 VDDA.t185 VDDA.t22 172.727
R499 VDDA.t124 VDDA.t185 172.727
R500 VDDA.t171 VDDA.t124 172.727
R501 VDDA.t207 VDDA.t171 172.727
R502 VDDA.t341 VDDA.t207 172.727
R503 VDDA.t308 VDDA.n232 172.554
R504 VDDA.n235 VDDA.t329 172.554
R505 VDDA.n340 VDDA.n339 168.435
R506 VDDA.n359 VDDA.n358 168.435
R507 VDDA.n361 VDDA.n360 168.435
R508 VDDA.n363 VDDA.n362 168.435
R509 VDDA.n365 VDDA.n364 168.435
R510 VDDA.n367 VDDA.n366 168.435
R511 VDDA.n369 VDDA.n368 168.435
R512 VDDA.n371 VDDA.n370 168.435
R513 VDDA.n245 VDDA.n218 164.8
R514 VDDA.n248 VDDA.n218 164.8
R515 VDDA.t344 VDDA.n137 161.817
R516 VDDA.t365 VDDA.n138 161.817
R517 VDDA.t362 VDDA.n42 161.817
R518 VDDA.n44 VDDA.t374 161.817
R519 VDDA.n91 VDDA.n89 160.428
R520 VDDA.n88 VDDA.n86 160.428
R521 VDDA.n67 VDDA.n65 160.428
R522 VDDA.n64 VDDA.n62 160.428
R523 VDDA.t257 VDDA.t332 159.814
R524 VDDA.t278 VDDA.t257 159.814
R525 VDDA.t289 VDDA.t278 159.814
R526 VDDA.t299 VDDA.t289 159.814
R527 VDDA.t264 VDDA.t299 159.814
R528 VDDA.t260 VDDA.t264 159.814
R529 VDDA.t283 VDDA.t260 159.814
R530 VDDA.t291 VDDA.t283 159.814
R531 VDDA.t269 VDDA.t250 159.814
R532 VDDA.t266 VDDA.t269 159.814
R533 VDDA.t285 VDDA.t266 159.814
R534 VDDA.t294 VDDA.t285 159.814
R535 VDDA.t255 VDDA.t294 159.814
R536 VDDA.t275 VDDA.t255 159.814
R537 VDDA.t273 VDDA.t275 159.814
R538 VDDA.t393 VDDA.t273 159.814
R539 VDDA.n91 VDDA.n90 159.803
R540 VDDA.n88 VDDA.n87 159.803
R541 VDDA.n67 VDDA.n66 159.803
R542 VDDA.n64 VDDA.n63 159.803
R543 VDDA.t26 VDDA.t323 158.333
R544 VDDA.t320 VDDA.t107 158.333
R545 VDDA.t244 VDDA.t359 158.333
R546 VDDA.t399 VDDA.t193 158.333
R547 VDDA.t173 VDDA.t387 158.333
R548 VDDA.t103 VDDA.t173 158.333
R549 VDDA.t210 VDDA.t466 158.333
R550 VDDA.t326 VDDA.t210 158.333
R551 VDDA.t109 VDDA.t408 155.97
R552 VDDA.t175 VDDA.t109 155.97
R553 VDDA.t448 VDDA.t175 155.97
R554 VDDA.t454 VDDA.t448 155.97
R555 VDDA.t101 VDDA.t454 155.97
R556 VDDA.t446 VDDA.t101 155.97
R557 VDDA.t450 VDDA.t177 155.97
R558 VDDA.t462 VDDA.t450 155.97
R559 VDDA.t212 VDDA.t462 155.97
R560 VDDA.t402 VDDA.t212 155.97
R561 VDDA.t201 VDDA.t305 155.97
R562 VDDA.t24 VDDA.t201 155.97
R563 VDDA.t452 VDDA.t130 155.97
R564 VDDA.t353 VDDA.t452 155.97
R565 VDDA.n97 VDDA.t406 155.125
R566 VDDA.n95 VDDA.t318 155.125
R567 VDDA.n73 VDDA.t303 155.125
R568 VDDA.n71 VDDA.t385 155.125
R569 VDDA.n134 VDDA.n133 151.882
R570 VDDA.n38 VDDA.n37 151.882
R571 VDDA.n148 VDDA.n147 151.321
R572 VDDA.n49 VDDA.n48 151.321
R573 VDDA.n124 VDDA.n116 150.4
R574 VDDA.n118 VDDA.n113 150.4
R575 VDDA.n24 VDDA.n16 150.4
R576 VDDA.n18 VDDA.n13 150.4
R577 VDDA.n107 VDDA.n106 146.002
R578 VDDA.n83 VDDA.n82 146.002
R579 VDDA.n111 VDDA.n110 145.429
R580 VDDA.n127 VDDA.n126 145.429
R581 VDDA.n129 VDDA.n128 145.429
R582 VDDA.n131 VDDA.n130 145.429
R583 VDDA.n133 VDDA.n132 145.429
R584 VDDA.n12 VDDA.n11 145.429
R585 VDDA.n31 VDDA.n30 145.429
R586 VDDA.n33 VDDA.n32 145.429
R587 VDDA.n35 VDDA.n34 145.429
R588 VDDA.n37 VDDA.n36 145.429
R589 VDDA.n147 VDDA.n146 135.387
R590 VDDA.n135 VDDA.n134 135.387
R591 VDDA.n48 VDDA.n47 135.387
R592 VDDA.n39 VDDA.n38 135.387
R593 VDDA.t153 VDDA.t347 121.513
R594 VDDA.t141 VDDA.t153 121.513
R595 VDDA.t80 VDDA.t141 121.513
R596 VDDA.t90 VDDA.t80 121.513
R597 VDDA.t45 VDDA.t90 121.513
R598 VDDA.t86 VDDA.t13 121.513
R599 VDDA.t83 VDDA.t86 121.513
R600 VDDA.t152 VDDA.t83 121.513
R601 VDDA.t134 VDDA.t152 121.513
R602 VDDA.t371 VDDA.t134 121.513
R603 VDDA.t226 VDDA.t368 121.513
R604 VDDA.t147 VDDA.t226 121.513
R605 VDDA.t216 VDDA.t147 121.513
R606 VDDA.t46 VDDA.t216 121.513
R607 VDDA.t225 VDDA.t46 121.513
R608 VDDA.t75 VDDA.t161 121.513
R609 VDDA.t217 VDDA.t75 121.513
R610 VDDA.t183 VDDA.t217 121.513
R611 VDDA.t144 VDDA.t183 121.513
R612 VDDA.t381 VDDA.t144 121.513
R613 VDDA.n334 VDDA.n265 118.4
R614 VDDA.n330 VDDA.n270 118.4
R615 VDDA.n292 VDDA.n284 118.4
R616 VDDA.n286 VDDA.n281 118.4
R617 VDDA.n395 VDDA.n394 118.4
R618 VDDA.n390 VDDA.n385 118.4
R619 VDDA.n356 VDDA.n355 118.4
R620 VDDA.n351 VDDA.n346 118.4
R621 VDDA.n454 VDDA.n453 118.4
R622 VDDA.n460 VDDA.n459 118.4
R623 VDDA.n441 VDDA.n440 118.4
R624 VDDA.n446 VDDA.n445 118.4
R625 VDDA.n422 VDDA.n421 118.4
R626 VDDA.n427 VDDA.n426 118.4
R627 VDDA.n245 VDDA.n244 110.4
R628 VDDA.n249 VDDA.n248 110.4
R629 VDDA.n453 VDDA.n402 105.6
R630 VDDA.n460 VDDA.n402 105.6
R631 VDDA.n421 VDDA.n414 105.6
R632 VDDA.n427 VDDA.n414 105.6
R633 VDDA.t329 VDDA.t99 102.704
R634 VDDA.n205 VDDA.n204 102.4
R635 VDDA.n210 VDDA.n209 102.4
R636 VDDA.n161 VDDA.n160 102.4
R637 VDDA.n240 VDDA.n239 101.267
R638 VDDA.t242 VDDA.t405 98.2764
R639 VDDA.t194 VDDA.t242 98.2764
R640 VDDA.t126 VDDA.t194 98.2764
R641 VDDA.t431 VDDA.t126 98.2764
R642 VDDA.t55 VDDA.t431 98.2764
R643 VDDA.t420 VDDA.t429 98.2764
R644 VDDA.t165 VDDA.t420 98.2764
R645 VDDA.t196 VDDA.t165 98.2764
R646 VDDA.t8 VDDA.t196 98.2764
R647 VDDA.t317 VDDA.t8 98.2764
R648 VDDA.t418 VDDA.t302 98.2764
R649 VDDA.t118 VDDA.t418 98.2764
R650 VDDA.t2 VDDA.t118 98.2764
R651 VDDA.t41 VDDA.t2 98.2764
R652 VDDA.t69 VDDA.t41 98.2764
R653 VDDA.t223 VDDA.t181 98.2764
R654 VDDA.t247 VDDA.t223 98.2764
R655 VDDA.t59 VDDA.t247 98.2764
R656 VDDA.t53 VDDA.t59 98.2764
R657 VDDA.t384 VDDA.t53 98.2764
R658 VDDA.n52 VDDA.n50 97.4034
R659 VDDA.n2 VDDA.n0 97.4034
R660 VDDA.n60 VDDA.n59 96.8409
R661 VDDA.n58 VDDA.n57 96.8409
R662 VDDA.n56 VDDA.n55 96.8409
R663 VDDA.n54 VDDA.n53 96.8409
R664 VDDA.n52 VDDA.n51 96.8409
R665 VDDA.n10 VDDA.n9 96.8409
R666 VDDA.n8 VDDA.n7 96.8409
R667 VDDA.n6 VDDA.n5 96.8409
R668 VDDA.n4 VDDA.n3 96.8409
R669 VDDA.n2 VDDA.n1 96.8409
R670 VDDA.n168 VDDA.n167 96.0005
R671 VDDA.n169 VDDA.n155 96.0005
R672 VDDA.n176 VDDA.n175 96.0005
R673 VDDA.n207 VDDA.t62 93.3041
R674 VDDA.t191 VDDA.n207 93.3041
R675 VDDA.n172 VDDA.t36 93.3041
R676 VDDA.n172 VDDA.t117 93.3041
R677 VDDA.n219 VDDA.n218 92.5005
R678 VDDA.t422 VDDA.n219 92.5005
R679 VDDA.n220 VDDA.n217 92.5005
R680 VDDA.t422 VDDA.n220 92.5005
R681 VDDA.n224 VDDA.n223 92.5005
R682 VDDA.n233 VDDA.n224 92.5005
R683 VDDA.n225 VDDA.n222 92.5005
R684 VDDA.n234 VDDA.n225 92.5005
R685 VDDA.n206 VDDA.n205 92.5005
R686 VDDA.n182 VDDA.n181 92.5005
R687 VDDA.n207 VDDA.n182 92.5005
R688 VDDA.n209 VDDA.n208 92.5005
R689 VDDA.n183 VDDA.n180 92.5005
R690 VDDA.n207 VDDA.n183 92.5005
R691 VDDA.n163 VDDA.n156 92.5005
R692 VDDA.n164 VDDA.n163 92.5005
R693 VDDA.n162 VDDA.n161 92.5005
R694 VDDA.n166 VDDA.n165 92.5005
R695 VDDA.n165 VDDA.n164 92.5005
R696 VDDA.n168 VDDA.n157 92.5005
R697 VDDA.n171 VDDA.n151 92.5005
R698 VDDA.n172 VDDA.n171 92.5005
R699 VDDA.n170 VDDA.n169 92.5005
R700 VDDA.n174 VDDA.n173 92.5005
R701 VDDA.n173 VDDA.n172 92.5005
R702 VDDA.n176 VDDA.n152 92.5005
R703 VDDA.n124 VDDA.n123 92.5005
R704 VDDA.n120 VDDA.n119 92.5005
R705 VDDA.n122 VDDA.n120 92.5005
R706 VDDA.n121 VDDA.n113 92.5005
R707 VDDA.n125 VDDA.n114 92.5005
R708 VDDA.n122 VDDA.n114 92.5005
R709 VDDA.n144 VDDA.n143 92.5005
R710 VDDA.n143 VDDA.n142 92.5005
R711 VDDA.n141 VDDA.n140 92.5005
R712 VDDA.n142 VDDA.n141 92.5005
R713 VDDA.n104 VDDA.n103 92.5005
R714 VDDA.n100 VDDA.n99 92.5005
R715 VDDA.n102 VDDA.n100 92.5005
R716 VDDA.n101 VDDA.n93 92.5005
R717 VDDA.n105 VDDA.n94 92.5005
R718 VDDA.n102 VDDA.n94 92.5005
R719 VDDA.n80 VDDA.n79 92.5005
R720 VDDA.n76 VDDA.n75 92.5005
R721 VDDA.n78 VDDA.n76 92.5005
R722 VDDA.n77 VDDA.n69 92.5005
R723 VDDA.n81 VDDA.n70 92.5005
R724 VDDA.n78 VDDA.n70 92.5005
R725 VDDA.n24 VDDA.n23 92.5005
R726 VDDA.n20 VDDA.n19 92.5005
R727 VDDA.n22 VDDA.n20 92.5005
R728 VDDA.n21 VDDA.n13 92.5005
R729 VDDA.n25 VDDA.n14 92.5005
R730 VDDA.n22 VDDA.n14 92.5005
R731 VDDA.n29 VDDA.n26 92.5005
R732 VDDA.n43 VDDA.n29 92.5005
R733 VDDA.n28 VDDA.n27 92.5005
R734 VDDA.n43 VDDA.n28 92.5005
R735 VDDA.n317 VDDA.n267 92.5005
R736 VDDA.n332 VDDA.n267 92.5005
R737 VDDA.n334 VDDA.n333 92.5005
R738 VDDA.n269 VDDA.n266 92.5005
R739 VDDA.n332 VDDA.n266 92.5005
R740 VDDA.n331 VDDA.n330 92.5005
R741 VDDA.n292 VDDA.n291 92.5005
R742 VDDA.n288 VDDA.n287 92.5005
R743 VDDA.n290 VDDA.n288 92.5005
R744 VDDA.n289 VDDA.n281 92.5005
R745 VDDA.n293 VDDA.n282 92.5005
R746 VDDA.n290 VDDA.n282 92.5005
R747 VDDA.n394 VDDA.n393 92.5005
R748 VDDA.n389 VDDA.n388 92.5005
R749 VDDA.n392 VDDA.n389 92.5005
R750 VDDA.n391 VDDA.n390 92.5005
R751 VDDA.n396 VDDA.n386 92.5005
R752 VDDA.n392 VDDA.n386 92.5005
R753 VDDA.n376 VDDA.n375 92.5005
R754 VDDA.n343 VDDA.n342 92.5005
R755 VDDA.n377 VDDA.n343 92.5005
R756 VDDA.n379 VDDA.n378 92.5005
R757 VDDA.n344 VDDA.n341 92.5005
R758 VDDA.n377 VDDA.n344 92.5005
R759 VDDA.n355 VDDA.n354 92.5005
R760 VDDA.n350 VDDA.n349 92.5005
R761 VDDA.n353 VDDA.n350 92.5005
R762 VDDA.n352 VDDA.n351 92.5005
R763 VDDA.n357 VDDA.n347 92.5005
R764 VDDA.n353 VDDA.n347 92.5005
R765 VDDA.n455 VDDA.n454 92.5005
R766 VDDA.n404 VDDA.n403 92.5005
R767 VDDA.n456 VDDA.n404 92.5005
R768 VDDA.n459 VDDA.n458 92.5005
R769 VDDA.n405 VDDA.n402 92.5005
R770 VDDA.n457 VDDA.n405 92.5005
R771 VDDA.n442 VDDA.n441 92.5005
R772 VDDA.n410 VDDA.n409 92.5005
R773 VDDA.n443 VDDA.n410 92.5005
R774 VDDA.n445 VDDA.n444 92.5005
R775 VDDA.n411 VDDA.n408 92.5005
R776 VDDA.n443 VDDA.n411 92.5005
R777 VDDA.n423 VDDA.n422 92.5005
R778 VDDA.n416 VDDA.n415 92.5005
R779 VDDA.n424 VDDA.n416 92.5005
R780 VDDA.n426 VDDA.n425 92.5005
R781 VDDA.n417 VDDA.n414 92.5005
R782 VDDA.n424 VDDA.n417 92.5005
R783 VDDA.n164 VDDA.t199 91.6672
R784 VDDA.n164 VDDA.t427 91.6672
R785 VDDA.n228 VDDA.n227 87.4672
R786 VDDA.n332 VDDA.t113 86.3641
R787 VDDA.t203 VDDA.n332 86.3641
R788 VDDA.n290 VDDA.t73 86.3641
R789 VDDA.t128 VDDA.n290 86.3641
R790 VDDA.n227 VDDA.t309 85.438
R791 VDDA.n239 VDDA.t330 85.438
R792 VDDA.n233 VDDA.t308 81.3068
R793 VDDA.n239 VDDA.n238 81.0672
R794 VDDA.n229 VDDA.n227 81.0672
R795 VDDA.n377 VDDA.t291 79.907
R796 VDDA.t250 VDDA.n377 79.907
R797 VDDA.n392 VDDA.t26 79.1672
R798 VDDA.t107 VDDA.n392 79.1672
R799 VDDA.n353 VDDA.t244 79.1672
R800 VDDA.t193 VDDA.n353 79.1672
R801 VDDA.t466 VDDA.n457 79.1672
R802 VDDA.n178 VDDA.t38 78.8005
R803 VDDA.n178 VDDA.t67 78.8005
R804 VDDA.n184 VDDA.t5 78.8005
R805 VDDA.n184 VDDA.t190 78.8005
R806 VDDA.n186 VDDA.t440 78.8005
R807 VDDA.n186 VDDA.t231 78.8005
R808 VDDA.n188 VDDA.t40 78.8005
R809 VDDA.n188 VDDA.t188 78.8005
R810 VDDA.n190 VDDA.t192 78.8005
R811 VDDA.n190 VDDA.t240 78.8005
R812 VDDA.n192 VDDA.t443 78.8005
R813 VDDA.n192 VDDA.t63 78.8005
R814 VDDA.n194 VDDA.t89 78.8005
R815 VDDA.n194 VDDA.t34 78.8005
R816 VDDA.n196 VDDA.t21 78.8005
R817 VDDA.n196 VDDA.t65 78.8005
R818 VDDA.n198 VDDA.t238 78.8005
R819 VDDA.n198 VDDA.t50 78.8005
R820 VDDA.n200 VDDA.t180 78.8005
R821 VDDA.n200 VDDA.t116 78.8005
R822 VDDA.n443 VDDA.t446 77.9856
R823 VDDA.t177 VDDA.n443 77.9856
R824 VDDA.n424 VDDA.t24 77.9856
R825 VDDA.t130 VDDA.n424 77.9856
R826 VDDA.n237 VDDA.n222 64.0005
R827 VDDA.n329 VDDA.n271 64.0005
R828 VDDA.n321 VDDA.n271 64.0005
R829 VDDA.n321 VDDA.n320 64.0005
R830 VDDA.n320 VDDA.n317 64.0005
R831 VDDA.n317 VDDA.n316 64.0005
R832 VDDA.n316 VDDA.n308 64.0005
R833 VDDA.n308 VDDA.n263 64.0005
R834 VDDA.n335 VDDA.n263 64.0005
R835 VDDA.n357 VDDA.n356 64.0005
R836 VDDA.n357 VDDA.n346 64.0005
R837 VDDA.t169 VDDA.t344 62.9523
R838 VDDA.t135 VDDA.t169 62.9523
R839 VDDA.t76 VDDA.t135 62.9523
R840 VDDA.t91 VDDA.t76 62.9523
R841 VDDA.t18 VDDA.t91 62.9523
R842 VDDA.t14 VDDA.t93 62.9523
R843 VDDA.t93 VDDA.t84 62.9523
R844 VDDA.t84 VDDA.t167 62.9523
R845 VDDA.t167 VDDA.t16 62.9523
R846 VDDA.t16 VDDA.t365 62.9523
R847 VDDA.t120 VDDA.t362 62.9523
R848 VDDA.t235 VDDA.t120 62.9523
R849 VDDA.t156 VDDA.t235 62.9523
R850 VDDA.t51 VDDA.t156 62.9523
R851 VDDA.t132 VDDA.t51 62.9523
R852 VDDA.t218 VDDA.t159 62.9523
R853 VDDA.t214 VDDA.t218 62.9523
R854 VDDA.t142 VDDA.t214 62.9523
R855 VDDA.t81 VDDA.t142 62.9523
R856 VDDA.t374 VDDA.t81 62.9523
R857 VDDA.n396 VDDA.n395 62.7205
R858 VDDA.n396 VDDA.n385 62.7205
R859 VDDA.n215 VDDA.t423 62.5402
R860 VDDA.n215 VDDA.t378 62.5402
R861 VDDA.n246 VDDA.n245 61.6672
R862 VDDA.n248 VDDA.n247 61.6672
R863 VDDA.n137 VDDA.n112 61.6672
R864 VDDA.n139 VDDA.n138 61.6672
R865 VDDA.n45 VDDA.n44 61.6672
R866 VDDA.n42 VDDA.n41 61.6672
R867 VDDA.n122 VDDA.t45 60.7563
R868 VDDA.t13 VDDA.n122 60.7563
R869 VDDA.n22 VDDA.t225 60.7563
R870 VDDA.t161 VDDA.n22 60.7563
R871 VDDA.n256 VDDA.t471 59.5681
R872 VDDA.n255 VDDA.t469 59.5681
R873 VDDA.n244 VDDA.n217 57.6005
R874 VDDA.n249 VDDA.n217 57.6005
R875 VDDA.n456 VDDA.t103 57.5763
R876 VDDA.n255 VDDA.t472 51.8888
R877 VDDA.n230 VDDA.n222 51.2005
R878 VDDA.n102 VDDA.t55 49.1384
R879 VDDA.t429 VDDA.n102 49.1384
R880 VDDA.n78 VDDA.t69 49.1384
R881 VDDA.t181 VDDA.n78 49.1384
R882 VDDA.n257 VDDA.t470 48.9557
R883 VDDA.n252 VDDA.n251 48.3605
R884 VDDA.n242 VDDA.n241 43.8605
R885 VDDA.n202 VDDA.n201 42.0963
R886 VDDA.n213 VDDA.n212 41.5338
R887 VDDA.n260 VDDA.t58 39.4005
R888 VDDA.n260 VDDA.t29 39.4005
R889 VDDA.n261 VDDA.t151 39.4005
R890 VDDA.n261 VDDA.t457 39.4005
R891 VDDA.n311 VDDA.t155 39.4005
R892 VDDA.n311 VDDA.t97 39.4005
R893 VDDA.n309 VDDA.t465 39.4005
R894 VDDA.n309 VDDA.t11 39.4005
R895 VDDA.n306 VDDA.t114 39.4005
R896 VDDA.n306 VDDA.t204 39.4005
R897 VDDA.n318 VDDA.t425 39.4005
R898 VDDA.n318 VDDA.t163 39.4005
R899 VDDA.n305 VDDA.t106 39.4005
R900 VDDA.n305 VDDA.t72 39.4005
R901 VDDA.n324 VDDA.t112 39.4005
R902 VDDA.n324 VDDA.t123 39.4005
R903 VDDA.n272 VDDA.t246 39.4005
R904 VDDA.n272 VDDA.t149 39.4005
R905 VDDA.n302 VDDA.t172 39.4005
R906 VDDA.n302 VDDA.t208 39.4005
R907 VDDA.n300 VDDA.t186 39.4005
R908 VDDA.n300 VDDA.t125 39.4005
R909 VDDA.n298 VDDA.t234 39.4005
R910 VDDA.n298 VDDA.t23 39.4005
R911 VDDA.n296 VDDA.t445 39.4005
R912 VDDA.n296 VDDA.t417 39.4005
R913 VDDA.n280 VDDA.t74 39.4005
R914 VDDA.n280 VDDA.t129 39.4005
R915 VDDA.n278 VDDA.t434 39.4005
R916 VDDA.n278 VDDA.t221 39.4005
R917 VDDA.n276 VDDA.t461 39.4005
R918 VDDA.n276 VDDA.t206 39.4005
R919 VDDA.n274 VDDA.t436 39.4005
R920 VDDA.n274 VDDA.t438 39.4005
R921 VDDA.n273 VDDA.t48 39.4005
R922 VDDA.n273 VDDA.t1 39.4005
R923 VDDA.n383 VDDA.t27 39.4005
R924 VDDA.n383 VDDA.t108 39.4005
R925 VDDA.n400 VDDA.t467 39.4005
R926 VDDA.n400 VDDA.t211 39.4005
R927 VDDA.n449 VDDA.t174 39.4005
R928 VDDA.n449 VDDA.t104 39.4005
R929 VDDA.n406 VDDA.t463 39.4005
R930 VDDA.n406 VDDA.t213 39.4005
R931 VDDA.n430 VDDA.t178 39.4005
R932 VDDA.n430 VDDA.t451 39.4005
R933 VDDA.n432 VDDA.t102 39.4005
R934 VDDA.n432 VDDA.t447 39.4005
R935 VDDA.n434 VDDA.t449 39.4005
R936 VDDA.n434 VDDA.t455 39.4005
R937 VDDA.n436 VDDA.t110 39.4005
R938 VDDA.n436 VDDA.t176 39.4005
R939 VDDA.n412 VDDA.t131 39.4005
R940 VDDA.n412 VDDA.t453 39.4005
R941 VDDA.n418 VDDA.t202 39.4005
R942 VDDA.n418 VDDA.t25 39.4005
R943 VDDA.n142 VDDA.t18 31.4764
R944 VDDA.n142 VDDA.t14 31.4764
R945 VDDA.n43 VDDA.t132 31.4764
R946 VDDA.t159 VDDA.n43 31.4764
R947 VDDA.n169 VDDA.n168 28.663
R948 VDDA.n251 VDDA.n250 25.6005
R949 VDDA.n243 VDDA.n242 25.6005
R950 VDDA.n212 VDDA.n211 25.6005
R951 VDDA.n203 VDDA.n202 25.6005
R952 VDDA.n258 VDDA.n254 24.7453
R953 VDDA.n250 VDDA.n249 24.5338
R954 VDDA.n244 VDDA.n243 24.5338
R955 VDDA.n238 VDDA.n237 24.5338
R956 VDDA.n230 VDDA.n229 24.5338
R957 VDDA.n457 VDDA.n456 21.5914
R958 VDDA.n211 VDDA.n210 21.3338
R959 VDDA.n204 VDDA.n203 21.3338
R960 VDDA.n160 VDDA.n159 21.3338
R961 VDDA.n167 VDDA.n158 21.3338
R962 VDDA.n155 VDDA.n154 21.3338
R963 VDDA.n175 VDDA.n153 21.3338
R964 VDDA.n118 VDDA.n117 21.3338
R965 VDDA.n116 VDDA.n115 21.3338
R966 VDDA.n146 VDDA.n145 21.3338
R967 VDDA.n136 VDDA.n135 21.3338
R968 VDDA.n98 VDDA.n97 21.3338
R969 VDDA.n96 VDDA.n95 21.3338
R970 VDDA.n74 VDDA.n73 21.3338
R971 VDDA.n72 VDDA.n71 21.3338
R972 VDDA.n18 VDDA.n17 21.3338
R973 VDDA.n16 VDDA.n15 21.3338
R974 VDDA.n47 VDDA.n46 21.3338
R975 VDDA.n40 VDDA.n39 21.3338
R976 VDDA.n265 VDDA.n264 21.3338
R977 VDDA.n270 VDDA.n268 21.3338
R978 VDDA.n284 VDDA.n283 21.3338
R979 VDDA.n286 VDDA.n285 21.3338
R980 VDDA.n395 VDDA.n387 21.3338
R981 VDDA.n385 VDDA.n384 21.3338
R982 VDDA.n356 VDDA.n348 21.3338
R983 VDDA.n346 VDDA.n345 21.3338
R984 VDDA.n61 VDDA.n60 21.1567
R985 VDDA.n177 VDDA.n176 19.5505
R986 VDDA.n144 VDDA.n125 19.538
R987 VDDA.n26 VDDA.n25 19.538
R988 VDDA.n254 VDDA.n253 19.4142
R989 VDDA.n107 VDDA.n105 19.2005
R990 VDDA.n83 VDDA.n81 19.2005
R991 VDDA.n381 VDDA.n380 19.2005
R992 VDDA.n374 VDDA.n373 19.2005
R993 VDDA.n461 VDDA.n460 19.2005
R994 VDDA.n453 VDDA.n452 19.2005
R995 VDDA.n447 VDDA.n446 19.2005
R996 VDDA.n440 VDDA.n439 19.2005
R997 VDDA.n428 VDDA.n427 19.2005
R998 VDDA.n421 VDDA.n420 19.2005
R999 VDDA.n232 VDDA.n231 18.5005
R1000 VDDA.n236 VDDA.n235 18.5005
R1001 VDDA.t99 VDDA.n234 17.1176
R1002 VDDA.n150 VDDA.n10 16.8443
R1003 VDDA.n372 VDDA.n357 16.363
R1004 VDDA.n468 VDDA.t259 15.0181
R1005 VDDA.n420 VDDA.n419 14.363
R1006 VDDA.n228 VDDA.n221 14.0505
R1007 VDDA.n373 VDDA.n372 13.8005
R1008 VDDA.n382 VDDA.n381 13.8005
R1009 VDDA.n452 VDDA.n451 13.8005
R1010 VDDA.n439 VDDA.n438 13.8005
R1011 VDDA.n429 VDDA.n428 13.8005
R1012 VDDA.n448 VDDA.n447 13.8005
R1013 VDDA.n462 VDDA.n461 13.8005
R1014 VDDA.n339 VDDA.t276 13.1338
R1015 VDDA.n339 VDDA.t274 13.1338
R1016 VDDA.n358 VDDA.t295 13.1338
R1017 VDDA.n358 VDDA.t256 13.1338
R1018 VDDA.n360 VDDA.t267 13.1338
R1019 VDDA.n360 VDDA.t286 13.1338
R1020 VDDA.n362 VDDA.t251 13.1338
R1021 VDDA.n362 VDDA.t270 13.1338
R1022 VDDA.n364 VDDA.t284 13.1338
R1023 VDDA.n364 VDDA.t292 13.1338
R1024 VDDA.n366 VDDA.t265 13.1338
R1025 VDDA.n366 VDDA.t261 13.1338
R1026 VDDA.n368 VDDA.t290 13.1338
R1027 VDDA.n368 VDDA.t300 13.1338
R1028 VDDA.n370 VDDA.t258 13.1338
R1029 VDDA.n370 VDDA.t279 13.1338
R1030 VDDA.t309 VDDA.n226 12.313
R1031 VDDA.n226 VDDA.t100 12.313
R1032 VDDA.n106 VDDA.t56 11.2576
R1033 VDDA.n106 VDDA.t430 11.2576
R1034 VDDA.n90 VDDA.t421 11.2576
R1035 VDDA.n90 VDDA.t166 11.2576
R1036 VDDA.n89 VDDA.t197 11.2576
R1037 VDDA.n89 VDDA.t9 11.2576
R1038 VDDA.n87 VDDA.t127 11.2576
R1039 VDDA.n87 VDDA.t432 11.2576
R1040 VDDA.n86 VDDA.t243 11.2576
R1041 VDDA.n86 VDDA.t195 11.2576
R1042 VDDA.n82 VDDA.t70 11.2576
R1043 VDDA.n82 VDDA.t182 11.2576
R1044 VDDA.n66 VDDA.t224 11.2576
R1045 VDDA.n66 VDDA.t248 11.2576
R1046 VDDA.n65 VDDA.t60 11.2576
R1047 VDDA.n65 VDDA.t54 11.2576
R1048 VDDA.n63 VDDA.t3 11.2576
R1049 VDDA.n63 VDDA.t42 11.2576
R1050 VDDA.n62 VDDA.t419 11.2576
R1051 VDDA.n62 VDDA.t119 11.2576
R1052 VDDA.n108 VDDA.n107 9.3005
R1053 VDDA.n84 VDDA.n83 9.3005
R1054 VDDA.n325 VDDA.n271 9.3005
R1055 VDDA.n322 VDDA.n321 9.3005
R1056 VDDA.n320 VDDA.n319 9.3005
R1057 VDDA.n317 VDDA.n307 9.3005
R1058 VDDA.n316 VDDA.n315 9.3005
R1059 VDDA.n312 VDDA.n308 9.3005
R1060 VDDA.n263 VDDA.n262 9.3005
R1061 VDDA.n336 VDDA.n335 9.3005
R1062 VDDA.n329 VDDA.n328 9.3005
R1063 VDDA.n294 VDDA.n293 9.3005
R1064 VDDA.n397 VDDA.n396 9.3005
R1065 VDDA.n241 VDDA.n240 8.53175
R1066 VDDA.n258 VDDA.n257 8.03219
R1067 VDDA.n59 VDDA.t145 8.0005
R1068 VDDA.n59 VDDA.t30 8.0005
R1069 VDDA.n57 VDDA.t146 8.0005
R1070 VDDA.n57 VDDA.t164 8.0005
R1071 VDDA.n55 VDDA.t468 8.0005
R1072 VDDA.n55 VDDA.t98 8.0005
R1073 VDDA.n53 VDDA.t158 8.0005
R1074 VDDA.n53 VDDA.t184 8.0005
R1075 VDDA.n51 VDDA.t458 8.0005
R1076 VDDA.n51 VDDA.t459 8.0005
R1077 VDDA.n50 VDDA.t222 8.0005
R1078 VDDA.n50 VDDA.t227 8.0005
R1079 VDDA.n9 VDDA.t241 8.0005
R1080 VDDA.n9 VDDA.t43 8.0005
R1081 VDDA.n7 VDDA.t138 8.0005
R1082 VDDA.n7 VDDA.t44 8.0005
R1083 VDDA.n5 VDDA.t139 8.0005
R1084 VDDA.n5 VDDA.t95 8.0005
R1085 VDDA.n3 VDDA.t140 8.0005
R1086 VDDA.n3 VDDA.t79 8.0005
R1087 VDDA.n1 VDDA.t137 8.0005
R1088 VDDA.n1 VDDA.t78 8.0005
R1089 VDDA.n0 VDDA.t87 8.0005
R1090 VDDA.n0 VDDA.t232 8.0005
R1091 VDDA.n463 VDDA.n462 7.44175
R1092 VDDA.n214 VDDA.n213 7.438
R1093 VDDA.n110 VDDA.t170 6.56717
R1094 VDDA.n110 VDDA.t136 6.56717
R1095 VDDA.n126 VDDA.t77 6.56717
R1096 VDDA.n126 VDDA.t92 6.56717
R1097 VDDA.n128 VDDA.t19 6.56717
R1098 VDDA.n128 VDDA.t15 6.56717
R1099 VDDA.n130 VDDA.t94 6.56717
R1100 VDDA.n130 VDDA.t85 6.56717
R1101 VDDA.n132 VDDA.t168 6.56717
R1102 VDDA.n132 VDDA.t17 6.56717
R1103 VDDA.n11 VDDA.t143 6.56717
R1104 VDDA.n11 VDDA.t82 6.56717
R1105 VDDA.n30 VDDA.t219 6.56717
R1106 VDDA.n30 VDDA.t215 6.56717
R1107 VDDA.n32 VDDA.t133 6.56717
R1108 VDDA.n32 VDDA.t160 6.56717
R1109 VDDA.n34 VDDA.t157 6.56717
R1110 VDDA.n34 VDDA.t52 6.56717
R1111 VDDA.n36 VDDA.t121 6.56717
R1112 VDDA.n36 VDDA.t236 6.56717
R1113 VDDA.n109 VDDA.n85 6.313
R1114 VDDA.n399 VDDA.n398 6.13371
R1115 VDDA.n338 VDDA.n337 6.098
R1116 VDDA.n253 VDDA.n252 6.0005
R1117 VDDA.n241 VDDA.n216 5.1255
R1118 VDDA.n109 VDDA.n108 5.063
R1119 VDDA.n85 VDDA.n84 5.063
R1120 VDDA.n108 VDDA.n92 4.5005
R1121 VDDA.n84 VDDA.n68 4.5005
R1122 VDDA.n150 VDDA.n149 4.5005
R1123 VDDA.n295 VDDA.n294 4.5005
R1124 VDDA.n328 VDDA.n327 4.5005
R1125 VDDA.n326 VDDA.n325 4.5005
R1126 VDDA.n323 VDDA.n322 4.5005
R1127 VDDA.n319 VDDA.n304 4.5005
R1128 VDDA.n310 VDDA.n307 4.5005
R1129 VDDA.n315 VDDA.n314 4.5005
R1130 VDDA.n313 VDDA.n312 4.5005
R1131 VDDA.n262 VDDA.n259 4.5005
R1132 VDDA.n337 VDDA.n336 4.5005
R1133 VDDA.n398 VDDA.n397 4.5005
R1134 VDDA.n234 VDDA.n233 4.27978
R1135 VDDA.n256 VDDA.n255 4.12334
R1136 VDDA.n469 VDDA 4.08025
R1137 VDDA.n85 VDDA.n61 3.688
R1138 VDDA.n149 VDDA.n109 3.5005
R1139 VDDA.n327 VDDA.n303 3.3755
R1140 VDDA.n257 VDDA.n256 2.93377
R1141 VDDA.n214 VDDA.n177 2.813
R1142 VDDA.n253 VDDA.n214 2.563
R1143 VDDA.n451 VDDA.n448 2.5005
R1144 VDDA.n398 VDDA.n382 2.47371
R1145 VDDA.n438 VDDA.n429 1.813
R1146 VDDA.n177 VDDA.n150 1.46925
R1147 VDDA VDDA.n469 1.20605
R1148 VDDA VDDA.n468 1.0815
R1149 VDDA.n372 VDDA.n371 1.0005
R1150 VDDA.n371 VDDA.n369 1.0005
R1151 VDDA.n369 VDDA.n367 1.0005
R1152 VDDA.n367 VDDA.n365 1.0005
R1153 VDDA.n365 VDDA.n363 1.0005
R1154 VDDA.n363 VDDA.n361 1.0005
R1155 VDDA.n361 VDDA.n359 1.0005
R1156 VDDA.n359 VDDA.n340 1.0005
R1157 VDDA.n382 VDDA.n340 1.0005
R1158 VDDA.n149 VDDA.n148 0.938
R1159 VDDA.n338 VDDA.n258 0.840625
R1160 VDDA.n469 VDDA.n254 0.7948
R1161 VDDA.n61 VDDA.n49 0.7505
R1162 VDDA.n399 VDDA.n338 0.74075
R1163 VDDA.n240 VDDA.n221 0.6255
R1164 VDDA.n92 VDDA.n91 0.6255
R1165 VDDA.n92 VDDA.n88 0.6255
R1166 VDDA.n68 VDDA.n67 0.6255
R1167 VDDA.n68 VDDA.n64 0.6255
R1168 VDDA.n277 VDDA.n275 0.6255
R1169 VDDA.n279 VDDA.n277 0.6255
R1170 VDDA.n295 VDDA.n279 0.6255
R1171 VDDA.n297 VDDA.n295 0.6255
R1172 VDDA.n299 VDDA.n297 0.6255
R1173 VDDA.n301 VDDA.n299 0.6255
R1174 VDDA.n303 VDDA.n301 0.6255
R1175 VDDA.n327 VDDA.n326 0.6255
R1176 VDDA.n326 VDDA.n323 0.6255
R1177 VDDA.n323 VDDA.n304 0.6255
R1178 VDDA.n310 VDDA.n304 0.6255
R1179 VDDA.n314 VDDA.n310 0.6255
R1180 VDDA.n314 VDDA.n313 0.6255
R1181 VDDA.n313 VDDA.n259 0.6255
R1182 VDDA.n337 VDDA.n259 0.6255
R1183 VDDA.n201 VDDA.n199 0.563
R1184 VDDA.n199 VDDA.n197 0.563
R1185 VDDA.n197 VDDA.n195 0.563
R1186 VDDA.n195 VDDA.n193 0.563
R1187 VDDA.n193 VDDA.n191 0.563
R1188 VDDA.n191 VDDA.n189 0.563
R1189 VDDA.n189 VDDA.n187 0.563
R1190 VDDA.n187 VDDA.n185 0.563
R1191 VDDA.n185 VDDA.n179 0.563
R1192 VDDA.n213 VDDA.n179 0.563
R1193 VDDA.n133 VDDA.n131 0.563
R1194 VDDA.n131 VDDA.n129 0.563
R1195 VDDA.n129 VDDA.n127 0.563
R1196 VDDA.n127 VDDA.n111 0.563
R1197 VDDA.n148 VDDA.n111 0.563
R1198 VDDA.n54 VDDA.n52 0.563
R1199 VDDA.n56 VDDA.n54 0.563
R1200 VDDA.n58 VDDA.n56 0.563
R1201 VDDA.n60 VDDA.n58 0.563
R1202 VDDA.n37 VDDA.n35 0.563
R1203 VDDA.n35 VDDA.n33 0.563
R1204 VDDA.n33 VDDA.n31 0.563
R1205 VDDA.n31 VDDA.n12 0.563
R1206 VDDA.n49 VDDA.n12 0.563
R1207 VDDA.n4 VDDA.n2 0.563
R1208 VDDA.n6 VDDA.n4 0.563
R1209 VDDA.n8 VDDA.n6 0.563
R1210 VDDA.n10 VDDA.n8 0.563
R1211 VDDA.n419 VDDA.n413 0.563
R1212 VDDA.n429 VDDA.n413 0.563
R1213 VDDA.n438 VDDA.n437 0.563
R1214 VDDA.n437 VDDA.n435 0.563
R1215 VDDA.n435 VDDA.n433 0.563
R1216 VDDA.n433 VDDA.n431 0.563
R1217 VDDA.n431 VDDA.n407 0.563
R1218 VDDA.n448 VDDA.n407 0.563
R1219 VDDA.n451 VDDA.n450 0.563
R1220 VDDA.n450 VDDA.n401 0.563
R1221 VDDA.n462 VDDA.n401 0.563
R1222 VDDA.n463 VDDA.n399 0.546875
R1223 VDDA.n468 VDDA.n463 0.370625
R1224 VDDA.n252 VDDA.n216 0.2505
R1225 VDDA.t252 VDDA.t268 0.1603
R1226 VDDA.t296 VDDA.t288 0.1603
R1227 VDDA.t293 VDDA.t253 0.1603
R1228 VDDA.t281 VDDA.t277 0.1603
R1229 VDDA.t254 VDDA.t271 0.1603
R1230 VDDA.t298 VDDA.t282 0.1603
R1231 VDDA.t272 VDDA.t287 0.1603
R1232 VDDA.t263 VDDA.t249 0.1603
R1233 VDDA.n465 VDDA.t280 0.159278
R1234 VDDA.n466 VDDA.t262 0.159278
R1235 VDDA.n467 VDDA.t297 0.159278
R1236 VDDA.n467 VDDA.t252 0.1368
R1237 VDDA.n467 VDDA.t296 0.1368
R1238 VDDA.n466 VDDA.t293 0.1368
R1239 VDDA.n466 VDDA.t281 0.1368
R1240 VDDA.n465 VDDA.t254 0.1368
R1241 VDDA.n465 VDDA.t298 0.1368
R1242 VDDA.n464 VDDA.t272 0.1368
R1243 VDDA.n464 VDDA.t263 0.1368
R1244 VDDA.t280 VDDA.n464 0.00152174
R1245 VDDA.t262 VDDA.n465 0.00152174
R1246 VDDA.t297 VDDA.n466 0.00152174
R1247 VDDA.t259 VDDA.n467 0.00152174
R1248 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.t15 354.854
R1249 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t30 346.8
R1250 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n11 339.522
R1251 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n4 339.522
R1252 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n9 335.022
R1253 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.t7 275.909
R1254 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.n6 227.909
R1255 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n8 222.034
R1256 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t27 184.097
R1257 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t19 184.097
R1258 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t31 184.097
R1259 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t14 184.097
R1260 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n10 166.05
R1261 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n5 166.05
R1262 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t4 48.0005
R1263 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t0 48.0005
R1264 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t6 48.0005
R1265 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t1 48.0005
R1266 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.t3 39.4005
R1267 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.t9 39.4005
R1268 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t8 39.4005
R1269 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t10 39.4005
R1270 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t2 39.4005
R1271 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t5 39.4005
R1272 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n2 33.1711
R1273 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n0 5.6255
R1274 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n3 5.28175
R1275 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t20 4.8295
R1276 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t29 4.8295
R1277 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t25 4.8295
R1278 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t35 4.8295
R1279 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t33 4.8295
R1280 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t17 4.8295
R1281 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t28 4.8295
R1282 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n7 4.5005
R1283 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t11 4.5005
R1284 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t32 4.5005
R1285 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t34 4.5005
R1286 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t21 4.5005
R1287 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t12 4.5005
R1288 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t16 4.5005
R1289 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t26 4.5005
R1290 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t22 4.5005
R1291 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t24 4.5005
R1292 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t23 4.5005
R1293 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t13 4.5005
R1294 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t18 4.5005
R1295 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t36 4.5005
R1296 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.n1 3.8075
R1297 bgr_0.cap_res1.t0 bgr_0.cap_res1.t18 178.633
R1298 bgr_0.cap_res1.t15 bgr_0.cap_res1.t1 0.1603
R1299 bgr_0.cap_res1.t11 bgr_0.cap_res1.t7 0.1603
R1300 bgr_0.cap_res1.t10 bgr_0.cap_res1.t16 0.1603
R1301 bgr_0.cap_res1.t8 bgr_0.cap_res1.t4 0.1603
R1302 bgr_0.cap_res1.t17 bgr_0.cap_res1.t2 0.1603
R1303 bgr_0.cap_res1.t13 bgr_0.cap_res1.t9 0.1603
R1304 bgr_0.cap_res1.t3 bgr_0.cap_res1.t6 0.1603
R1305 bgr_0.cap_res1.t20 bgr_0.cap_res1.t14 0.1603
R1306 bgr_0.cap_res1.n1 bgr_0.cap_res1.t5 0.159278
R1307 bgr_0.cap_res1.n2 bgr_0.cap_res1.t19 0.159278
R1308 bgr_0.cap_res1.n3 bgr_0.cap_res1.t12 0.159278
R1309 bgr_0.cap_res1.n3 bgr_0.cap_res1.t15 0.1368
R1310 bgr_0.cap_res1.n3 bgr_0.cap_res1.t11 0.1368
R1311 bgr_0.cap_res1.n2 bgr_0.cap_res1.t10 0.1368
R1312 bgr_0.cap_res1.n2 bgr_0.cap_res1.t8 0.1368
R1313 bgr_0.cap_res1.n1 bgr_0.cap_res1.t17 0.1368
R1314 bgr_0.cap_res1.n1 bgr_0.cap_res1.t13 0.1368
R1315 bgr_0.cap_res1.n0 bgr_0.cap_res1.t3 0.1368
R1316 bgr_0.cap_res1.n0 bgr_0.cap_res1.t20 0.1368
R1317 bgr_0.cap_res1.t5 bgr_0.cap_res1.n0 0.00152174
R1318 bgr_0.cap_res1.t19 bgr_0.cap_res1.n1 0.00152174
R1319 bgr_0.cap_res1.t12 bgr_0.cap_res1.n2 0.00152174
R1320 bgr_0.cap_res1.t18 bgr_0.cap_res1.n3 0.00152174
R1321 a_14640_5738.t0 a_14640_5738.t1 169.905
R1322 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 345.264
R1323 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 344.7
R1324 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 344.7
R1325 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 206.052
R1326 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 205.488
R1327 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 205.488
R1328 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 205.488
R1329 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 205.488
R1330 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 122.474
R1331 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 81.2505
R1332 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 39.4005
R1333 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 39.4005
R1334 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 39.4005
R1335 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 39.4005
R1336 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 39.4005
R1337 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 39.4005
R1338 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 19.7005
R1339 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 19.7005
R1340 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 19.7005
R1341 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 19.7005
R1342 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 19.7005
R1343 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 19.7005
R1344 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 19.7005
R1345 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 19.7005
R1346 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 19.7005
R1347 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 19.7005
R1348 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 6.15675
R1349 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 6.1255
R1350 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 0.563
R1351 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 0.563
R1352 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 0.563
R1353 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 0.563
R1354 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 0.21925
R1355 GNDA.n2297 GNDA.n85 558653
R1356 GNDA.n2294 GNDA.n2293 138008
R1357 GNDA.n2293 GNDA.n2292 68623.1
R1358 GNDA.n2297 GNDA.n2296 63946.7
R1359 GNDA.n2287 GNDA.n2286 41223.8
R1360 GNDA.n2342 GNDA.n46 35574.1
R1361 GNDA.n2341 GNDA.n47 34650
R1362 GNDA.n86 GNDA.n50 33145.9
R1363 GNDA.n2288 GNDA.n24 32661.5
R1364 GNDA.n2435 GNDA.n24 32661.5
R1365 GNDA.n2289 GNDA.n46 29770.1
R1366 GNDA.n2287 GNDA.n2191 28842.3
R1367 GNDA.n2436 GNDA.n45 28430.8
R1368 GNDA.n2292 GNDA.n47 27818.3
R1369 GNDA.n867 GNDA.n866 26648.4
R1370 GNDA.n867 GNDA.n51 26648.4
R1371 GNDA.n2290 GNDA.n2289 24234.9
R1372 GNDA.n2296 GNDA.n87 24147.7
R1373 GNDA.n2295 GNDA.n2294 22990.2
R1374 GNDA.n86 GNDA.n48 21292.6
R1375 GNDA.n46 GNDA.n24 19630.8
R1376 GNDA.n2489 GNDA.n24 19630.8
R1377 GNDA.n2340 GNDA.n49 17297.8
R1378 GNDA.n2338 GNDA.n51 17265.8
R1379 GNDA.n2294 GNDA.n49 16323.6
R1380 GNDA.n51 GNDA.n50 15861.4
R1381 GNDA.n2289 GNDA.n2288 14714.3
R1382 GNDA.n2435 GNDA.n2434 14314.3
R1383 GNDA.n87 GNDA.n86 13428.1
R1384 GNDA.n870 GNDA.n869 12361.8
R1385 GNDA.n871 GNDA.n869 12312.5
R1386 GNDA.n875 GNDA.n870 11918.5
R1387 GNDA.n875 GNDA.n871 11869.2
R1388 GNDA.n866 GNDA.n87 11169.2
R1389 GNDA.n2490 GNDA.n23 10835
R1390 GNDA.n2488 GNDA.n23 10835
R1391 GNDA.n2488 GNDA.n22 10835
R1392 GNDA.n2490 GNDA.n22 10835
R1393 GNDA.n949 GNDA.n867 10371.4
R1394 GNDA.n2437 GNDA.n2436 10371.4
R1395 GNDA.n2102 GNDA.n85 9680
R1396 GNDA.n2292 GNDA.n46 9476.92
R1397 GNDA.n2194 GNDA.n6 9308.25
R1398 GNDA.n2494 GNDA.n6 9308.25
R1399 GNDA.n2194 GNDA.n7 9308.25
R1400 GNDA.n2494 GNDA.n7 9308.25
R1401 GNDA.n2447 GNDA.n2440 9259
R1402 GNDA.n2329 GNDA.n57 9062
R1403 GNDA.n2449 GNDA.n2440 8914.25
R1404 GNDA.n49 GNDA.n47 8695.24
R1405 GNDA.n2447 GNDA.n43 8175.5
R1406 GNDA.n2299 GNDA.n82 8175.5
R1407 GNDA.n2299 GNDA.n81 8126.25
R1408 GNDA.n866 GNDA.n85 7953.85
R1409 GNDA.n2332 GNDA.n53 7880
R1410 GNDA.n2336 GNDA.n53 7880
R1411 GNDA.n955 GNDA.n863 7880
R1412 GNDA.n951 GNDA.n863 7880
R1413 GNDA.n2449 GNDA.n43 7830.75
R1414 GNDA.n2332 GNDA.n54 7830.75
R1415 GNDA.n2336 GNDA.n54 7830.75
R1416 GNDA.n955 GNDA.n864 7830.75
R1417 GNDA.n951 GNDA.n864 7830.75
R1418 GNDA.n2290 GNDA.n2190 7752.38
R1419 GNDA.n2259 GNDA.n2200 7732.25
R1420 GNDA.n2259 GNDA.n2201 7732.25
R1421 GNDA.n2261 GNDA.n2200 7732.25
R1422 GNDA.n2261 GNDA.n2201 7732.25
R1423 GNDA.n2393 GNDA.n2353 7732.25
R1424 GNDA.n2424 GNDA.n2353 7732.25
R1425 GNDA.n2393 GNDA.n2361 7732.25
R1426 GNDA.n2424 GNDA.n2361 7732.25
R1427 GNDA.n2303 GNDA.n82 7732.25
R1428 GNDA.n2303 GNDA.n81 7683
R1429 GNDA.n2293 GNDA.n2291 7617.62
R1430 GNDA.n2372 GNDA.n2343 7338.25
R1431 GNDA.n2239 GNDA.n2217 7338.25
R1432 GNDA.n2432 GNDA.n2343 7289
R1433 GNDA.n2234 GNDA.n2217 7092
R1434 GNDA.n1648 GNDA.n515 6845.75
R1435 GNDA.n1649 GNDA.n515 6845.75
R1436 GNDA.n1655 GNDA.n1648 6796.5
R1437 GNDA.n1655 GNDA.n1649 6796.5
R1438 GNDA.n1646 GNDA.n72 6698
R1439 GNDA.n2313 GNDA.n72 6698
R1440 GNDA.n1646 GNDA.n68 6648.75
R1441 GNDA.n2313 GNDA.n68 6648.75
R1442 GNDA.n2250 GNDA.n2208 6057.75
R1443 GNDA.n2252 GNDA.n2250 6057.75
R1444 GNDA.n2208 GNDA.n2205 6057.75
R1445 GNDA.n2252 GNDA.n2205 6057.75
R1446 GNDA.n2358 GNDA.n2351 6057.75
R1447 GNDA.n2427 GNDA.n2351 6057.75
R1448 GNDA.n2358 GNDA.n2352 6057.75
R1449 GNDA.n2427 GNDA.n2352 6057.75
R1450 GNDA.n2372 GNDA.n2344 5319
R1451 GNDA.n2239 GNDA.n2218 5319
R1452 GNDA.n2432 GNDA.n2344 5269.75
R1453 GNDA.n2234 GNDA.n2218 5269.75
R1454 GNDA.n2246 GNDA.n2212 5171.25
R1455 GNDA.n2386 GNDA.n2366 5171.25
R1456 GNDA.n2242 GNDA.n2212 5122
R1457 GNDA.n2368 GNDA.n2366 5122
R1458 GNDA.n2329 GNDA.n58 4974.25
R1459 GNDA.n936 GNDA.n923 4974.25
R1460 GNDA.n937 GNDA.n936 4974.25
R1461 GNDA.n2246 GNDA.n2213 4944.7
R1462 GNDA.n2386 GNDA.n2385 4944.7
R1463 GNDA.n2461 GNDA.n25 4925
R1464 GNDA.n2475 GNDA.n25 4925
R1465 GNDA.n2242 GNDA.n2213 4895.45
R1466 GNDA.n2385 GNDA.n2368 4895.45
R1467 GNDA.n2461 GNDA.n26 4728
R1468 GNDA.n2475 GNDA.n26 4728
R1469 GNDA.n2114 GNDA.n2108 4678.75
R1470 GNDA.n2114 GNDA.n2106 4629.5
R1471 GNDA.n2110 GNDA.n2108 4629.5
R1472 GNDA.n2173 GNDA.n106 4580.25
R1473 GNDA.n106 GNDA.n102 4580.25
R1474 GNDA.n2110 GNDA.n2106 4580.25
R1475 GNDA.n2167 GNDA.n104 4580.25
R1476 GNDA.n2167 GNDA.n103 4580.25
R1477 GNDA.n948 GNDA.n876 4531
R1478 GNDA.n948 GNDA.n877 4531
R1479 GNDA.n876 GNDA.n868 4531
R1480 GNDA.n877 GNDA.n868 4531
R1481 GNDA.n923 GNDA.n922 4531
R1482 GNDA.n937 GNDA.n922 4531
R1483 GNDA.n2173 GNDA.n105 4481.75
R1484 GNDA.n105 GNDA.n102 4481.75
R1485 GNDA.n519 GNDA.n104 4481.75
R1486 GNDA.n519 GNDA.n103 4481.75
R1487 GNDA.n2296 GNDA.n2295 3708.05
R1488 GNDA.n2283 GNDA.n32 3595.25
R1489 GNDA.n2458 GNDA.n32 3595.25
R1490 GNDA.n2497 GNDA.n4 3349
R1491 GNDA.n2443 GNDA.n4 3299.75
R1492 GNDA.n2338 GNDA.n2337 3287.9
R1493 GNDA.n2283 GNDA.n33 3250.5
R1494 GNDA.n2458 GNDA.n33 3250.5
R1495 GNDA.n2497 GNDA.n5 3250.5
R1496 GNDA.n2443 GNDA.n5 3201.25
R1497 GNDA.n2339 GNDA.n50 3156.82
R1498 GNDA.n2436 GNDA.n2435 2933.33
R1499 GNDA.n2288 GNDA.n2287 2933.33
R1500 GNDA.n2225 GNDA.n2190 2928.06
R1501 GNDA.n2341 GNDA.n2340 2386.89
R1502 GNDA.n2224 GNDA.n2223 2326.02
R1503 GNDA.n2223 GNDA.n2222 2326.02
R1504 GNDA.n2382 GNDA.n2369 2326.02
R1505 GNDA.n2375 GNDA.n2369 2326.02
R1506 GNDA.n912 GNDA.n908 2142.38
R1507 GNDA.n931 GNDA.n921 2142.38
R1508 GNDA.n908 GNDA.n883 1846.88
R1509 GNDA.n941 GNDA.n921 1846.88
R1510 GNDA.n1070 GNDA.n842 1672.5
R1511 GNDA.n2340 GNDA.n2339 1609.95
R1512 GNDA.n2233 GNDA.n2190 1255.01
R1513 GNDA.n2339 GNDA.n2338 1226.55
R1514 GNDA.n1536 GNDA.n828 1214.72
R1515 GNDA.n1530 GNDA.n828 1214.72
R1516 GNDA.n1530 GNDA.n1094 1214.72
R1517 GNDA.n1520 GNDA.n1094 1214.72
R1518 GNDA.n1520 GNDA.n619 1214.72
R1519 GNDA.n1513 GNDA.n620 1214.72
R1520 GNDA.n1513 GNDA.n1106 1214.72
R1521 GNDA.n1190 GNDA.n1106 1214.72
R1522 GNDA.n1502 GNDA.n1190 1214.72
R1523 GNDA.n1502 GNDA.n621 1214.72
R1524 GNDA.n2228 GNDA.n2223 1114.8
R1525 GNDA.n2379 GNDA.n2369 1114.8
R1526 GNDA.t250 GNDA.n807 1064.42
R1527 GNDA.n827 GNDA.n826 1064.42
R1528 GNDA.n2434 GNDA.n2433 1055.59
R1529 GNDA.t250 GNDA.n1559 1041.66
R1530 GNDA.n833 GNDA.n827 1041.66
R1531 GNDA.n915 GNDA.n908 991.841
R1532 GNDA.n933 GNDA.n921 991.841
R1533 GNDA.n1647 GNDA.n516 964.235
R1534 GNDA.n2340 GNDA.n48 919.673
R1535 GNDA.t250 GNDA.n619 823.313
R1536 GNDA.n872 GNDA.n61 803.201
R1537 GNDA.n873 GNDA.n61 800
R1538 GNDA.n874 GNDA.n872 774.4
R1539 GNDA.n874 GNDA.n873 771.201
R1540 GNDA.n2348 GNDA.t271 734.418
R1541 GNDA.n2354 GNDA.t256 734.418
R1542 GNDA.n2206 GNDA.t279 734.418
R1543 GNDA.n2209 GNDA.t274 734.418
R1544 GNDA.n2487 GNDA.n2481 704
R1545 GNDA.n2487 GNDA.n2486 697.601
R1546 GNDA.n2295 GNDA.n48 685.899
R1547 GNDA.n2455 GNDA.t239 682.201
R1548 GNDA.n2415 GNDA.t282 682.201
R1549 GNDA.n573 GNDA.n572 669.307
R1550 GNDA.n2280 GNDA.t253 666.134
R1551 GNDA.n2452 GNDA.t318 666.134
R1552 GNDA.n1872 GNDA.n401 662.155
R1553 GNDA.n2144 GNDA.n127 662.155
R1554 GNDA.n2381 GNDA.n2370 617.601
R1555 GNDA.n2221 GNDA.n2220 617.601
R1556 GNDA.n2446 GNDA.n2445 601.601
R1557 GNDA.n2493 GNDA.n2492 598.4
R1558 GNDA.n2492 GNDA.n17 598.4
R1559 GNDA.n571 GNDA.n568 585
R1560 GNDA.n570 GNDA.n569 585
R1561 GNDA.n570 GNDA.n360 585
R1562 GNDA.n1214 GNDA.n1213 585
R1563 GNDA.n1212 GNDA.n1211 585
R1564 GNDA.n1210 GNDA.n1209 585
R1565 GNDA.n1208 GNDA.n1207 585
R1566 GNDA.n1206 GNDA.n1205 585
R1567 GNDA.n1204 GNDA.n1203 585
R1568 GNDA.n1202 GNDA.n1201 585
R1569 GNDA.n1200 GNDA.n1199 585
R1570 GNDA.n1198 GNDA.n1197 585
R1571 GNDA.n1196 GNDA.n1195 585
R1572 GNDA.n353 GNDA.n352 585
R1573 GNDA.n1964 GNDA.n1963 585
R1574 GNDA.n1535 GNDA.n1534 585
R1575 GNDA.n1536 GNDA.n1535 585
R1576 GNDA.n1533 GNDA.n830 585
R1577 GNDA.n830 GNDA.n828 585
R1578 GNDA.n1532 GNDA.n1531 585
R1579 GNDA.n1531 GNDA.n1530 585
R1580 GNDA.n1093 GNDA.n1092 585
R1581 GNDA.n1094 GNDA.n1093 585
R1582 GNDA.n1519 GNDA.n1518 585
R1583 GNDA.n1520 GNDA.n1519 585
R1584 GNDA.n1517 GNDA.n1103 585
R1585 GNDA.n1103 GNDA.n619 585
R1586 GNDA.n1516 GNDA.n1515 585
R1587 GNDA.n1515 GNDA.n620 585
R1588 GNDA.n1514 GNDA.n1104 585
R1589 GNDA.n1514 GNDA.n1513 585
R1590 GNDA.n1193 GNDA.n1105 585
R1591 GNDA.n1106 GNDA.n1105 585
R1592 GNDA.n1194 GNDA.n1191 585
R1593 GNDA.n1191 GNDA.n1190 585
R1594 GNDA.n1501 GNDA.n1500 585
R1595 GNDA.n1502 GNDA.n1501 585
R1596 GNDA.n1499 GNDA.n1192 585
R1597 GNDA.n1192 GNDA.n621 585
R1598 GNDA.n1866 GNDA.n402 585
R1599 GNDA.n1477 GNDA.n404 585
R1600 GNDA.n1478 GNDA.n1475 585
R1601 GNDA.n1481 GNDA.n1474 585
R1602 GNDA.n1482 GNDA.n1473 585
R1603 GNDA.n1485 GNDA.n1472 585
R1604 GNDA.n1486 GNDA.n1471 585
R1605 GNDA.n1489 GNDA.n1470 585
R1606 GNDA.n1490 GNDA.n1469 585
R1607 GNDA.n1493 GNDA.n1468 585
R1608 GNDA.n1494 GNDA.n416 585
R1609 GNDA.n1866 GNDA.n416 585
R1610 GNDA.n1497 GNDA.n1496 585
R1611 GNDA.n1496 GNDA.n590 585
R1612 GNDA.n1495 GNDA.n1494 585
R1613 GNDA.n1493 GNDA.n1492 585
R1614 GNDA.n1491 GNDA.n1490 585
R1615 GNDA.n1489 GNDA.n1488 585
R1616 GNDA.n1487 GNDA.n1486 585
R1617 GNDA.n1485 GNDA.n1484 585
R1618 GNDA.n1483 GNDA.n1482 585
R1619 GNDA.n1481 GNDA.n1480 585
R1620 GNDA.n1479 GNDA.n1478 585
R1621 GNDA.n1477 GNDA.n1476 585
R1622 GNDA.n1568 GNDA.n601 585
R1623 GNDA.n1568 GNDA.n607 585
R1624 GNDA.n1408 GNDA.n1407 585
R1625 GNDA.n1405 GNDA.n1348 585
R1626 GNDA.n1404 GNDA.n1349 585
R1627 GNDA.n1402 GNDA.n1401 585
R1628 GNDA.n1400 GNDA.n1350 585
R1629 GNDA.n1399 GNDA.n1398 585
R1630 GNDA.n1397 GNDA.n1351 585
R1631 GNDA.n1395 GNDA.n1394 585
R1632 GNDA.n1393 GNDA.n1353 585
R1633 GNDA.n1392 GNDA.n1391 585
R1634 GNDA.n1390 GNDA.n1354 585
R1635 GNDA.n1388 GNDA.n1387 585
R1636 GNDA.n1866 GNDA.n411 585
R1637 GNDA.n1249 GNDA.n1248 585
R1638 GNDA.n1241 GNDA.n1240 585
R1639 GNDA.n1320 GNDA.n1319 585
R1640 GNDA.n1323 GNDA.n1322 585
R1641 GNDA.n1239 GNDA.n1236 585
R1642 GNDA.n1232 GNDA.n1231 585
R1643 GNDA.n1331 GNDA.n1330 585
R1644 GNDA.n1334 GNDA.n1333 585
R1645 GNDA.n1230 GNDA.n1227 585
R1646 GNDA.n1223 GNDA.n1222 585
R1647 GNDA.n1342 GNDA.n1341 585
R1648 GNDA.n1345 GNDA.n1344 585
R1649 GNDA.n1215 GNDA.n1189 585
R1650 GNDA.n1189 GNDA.n621 585
R1651 GNDA.n1504 GNDA.n1503 585
R1652 GNDA.n1503 GNDA.n1502 585
R1653 GNDA.n1188 GNDA.n1120 585
R1654 GNDA.n1190 GNDA.n1188 585
R1655 GNDA.n1110 GNDA.n1108 585
R1656 GNDA.n1108 GNDA.n1106 585
R1657 GNDA.n1512 GNDA.n1511 585
R1658 GNDA.n1513 GNDA.n1512 585
R1659 GNDA.n1113 GNDA.n1107 585
R1660 GNDA.n1107 GNDA.n620 585
R1661 GNDA.n1112 GNDA.n1102 585
R1662 GNDA.n1102 GNDA.n619 585
R1663 GNDA.n1522 GNDA.n1521 585
R1664 GNDA.n1521 GNDA.n1520 585
R1665 GNDA.n1098 GNDA.n1095 585
R1666 GNDA.n1095 GNDA.n1094 585
R1667 GNDA.n1529 GNDA.n1528 585
R1668 GNDA.n1530 GNDA.n1529 585
R1669 GNDA.n1096 GNDA.n823 585
R1670 GNDA.n828 GNDA.n823 585
R1671 GNDA.n1538 GNDA.n1537 585
R1672 GNDA.n1537 GNDA.n1536 585
R1673 GNDA.n1217 GNDA.n1216 585
R1674 GNDA.n1216 GNDA.n590 585
R1675 GNDA.n1568 GNDA.n608 585
R1676 GNDA.n1466 GNDA.n1464 585
R1677 GNDA.n1463 GNDA.n1462 585
R1678 GNDA.n1461 GNDA.n1459 585
R1679 GNDA.n1458 GNDA.n1457 585
R1680 GNDA.n1454 GNDA.n1453 585
R1681 GNDA.n1452 GNDA.n1451 585
R1682 GNDA.n1448 GNDA.n1447 585
R1683 GNDA.n1446 GNDA.n1445 585
R1684 GNDA.n1442 GNDA.n1441 585
R1685 GNDA.n1440 GNDA.n422 585
R1686 GNDA.n1866 GNDA.n422 585
R1687 GNDA.n1438 GNDA.n1347 585
R1688 GNDA.n1438 GNDA.n590 585
R1689 GNDA.n1440 GNDA.n1439 585
R1690 GNDA.n1443 GNDA.n1442 585
R1691 GNDA.n1445 GNDA.n1444 585
R1692 GNDA.n1449 GNDA.n1448 585
R1693 GNDA.n1451 GNDA.n1450 585
R1694 GNDA.n1455 GNDA.n1454 585
R1695 GNDA.n1457 GNDA.n1456 585
R1696 GNDA.n1461 GNDA.n1460 585
R1697 GNDA.n1462 GNDA.n595 585
R1698 GNDA.n1568 GNDA.n595 585
R1699 GNDA.n1466 GNDA.n1465 585
R1700 GNDA.n811 GNDA.n809 585
R1701 GNDA.n1417 GNDA.n1416 585
R1702 GNDA.n1419 GNDA.n1418 585
R1703 GNDA.n1421 GNDA.n1414 585
R1704 GNDA.n1424 GNDA.n1423 585
R1705 GNDA.n1425 GNDA.n1413 585
R1706 GNDA.n1427 GNDA.n1426 585
R1707 GNDA.n1429 GNDA.n1412 585
R1708 GNDA.n1432 GNDA.n1431 585
R1709 GNDA.n1433 GNDA.n1411 585
R1710 GNDA.n1435 GNDA.n1434 585
R1711 GNDA.n1437 GNDA.n1410 585
R1712 GNDA.n826 GNDA.n822 585
R1713 GNDA.n825 GNDA.n824 585
R1714 GNDA.n1540 GNDA.n819 585
R1715 GNDA.n819 GNDA.n818 585
R1716 GNDA.n1542 GNDA.n1541 585
R1717 GNDA.n1543 GNDA.n1542 585
R1718 GNDA.n817 GNDA.n816 585
R1719 GNDA.n1544 GNDA.n817 585
R1720 GNDA.n1547 GNDA.n1546 585
R1721 GNDA.n1546 GNDA.n1545 585
R1722 GNDA.n1548 GNDA.n815 585
R1723 GNDA.n815 GNDA.n814 585
R1724 GNDA.n1550 GNDA.n1549 585
R1725 GNDA.n1551 GNDA.n1550 585
R1726 GNDA.n813 GNDA.n812 585
R1727 GNDA.n1552 GNDA.n813 585
R1728 GNDA.n1555 GNDA.n1554 585
R1729 GNDA.n1554 GNDA.n1553 585
R1730 GNDA.n1556 GNDA.n810 585
R1731 GNDA.n810 GNDA.n808 585
R1732 GNDA.n1558 GNDA.n1557 585
R1733 GNDA.n1559 GNDA.n1558 585
R1734 GNDA.n1091 GNDA.n829 585
R1735 GNDA.n833 GNDA.n829 585
R1736 GNDA.n1090 GNDA.n1089 585
R1737 GNDA.n1089 GNDA.n1088 585
R1738 GNDA.n832 GNDA.n831 585
R1739 GNDA.n1087 GNDA.n832 585
R1740 GNDA.n1085 GNDA.n1084 585
R1741 GNDA.n1086 GNDA.n1085 585
R1742 GNDA.n1083 GNDA.n835 585
R1743 GNDA.n835 GNDA.n834 585
R1744 GNDA.n1082 GNDA.n1081 585
R1745 GNDA.n1081 GNDA.n1080 585
R1746 GNDA.n837 GNDA.n836 585
R1747 GNDA.n1079 GNDA.n837 585
R1748 GNDA.n1077 GNDA.n1076 585
R1749 GNDA.n1078 GNDA.n1077 585
R1750 GNDA.n1075 GNDA.n839 585
R1751 GNDA.n839 GNDA.n838 585
R1752 GNDA.n1074 GNDA.n1073 585
R1753 GNDA.n1073 GNDA.n1072 585
R1754 GNDA.n1071 GNDA.n841 585
R1755 GNDA.n1070 GNDA.n1069 585
R1756 GNDA.n693 GNDA.n692 585
R1757 GNDA.n692 GNDA.n691 585
R1758 GNDA.n628 GNDA.n627 585
R1759 GNDA.n690 GNDA.n628 585
R1760 GNDA.n688 GNDA.n687 585
R1761 GNDA.n689 GNDA.n688 585
R1762 GNDA.n686 GNDA.n631 585
R1763 GNDA.n631 GNDA.n630 585
R1764 GNDA.n685 GNDA.n684 585
R1765 GNDA.n684 GNDA.n683 585
R1766 GNDA.n633 GNDA.n632 585
R1767 GNDA.n682 GNDA.n633 585
R1768 GNDA.n680 GNDA.n679 585
R1769 GNDA.n681 GNDA.n680 585
R1770 GNDA.n678 GNDA.n635 585
R1771 GNDA.n635 GNDA.n634 585
R1772 GNDA.n677 GNDA.n676 585
R1773 GNDA.n676 GNDA.n675 585
R1774 GNDA.n637 GNDA.n636 585
R1775 GNDA.n674 GNDA.n637 585
R1776 GNDA.n672 GNDA.n671 585
R1777 GNDA.n673 GNDA.n672 585
R1778 GNDA.n670 GNDA.n639 585
R1779 GNDA.n639 GNDA.n638 585
R1780 GNDA.n669 GNDA.n668 585
R1781 GNDA.n668 GNDA.n667 585
R1782 GNDA.n641 GNDA.n640 585
R1783 GNDA.n666 GNDA.n641 585
R1784 GNDA.n664 GNDA.n663 585
R1785 GNDA.n665 GNDA.n664 585
R1786 GNDA.n662 GNDA.n642 585
R1787 GNDA.n642 GNDA.n617 585
R1788 GNDA.n661 GNDA.n660 585
R1789 GNDA.n660 GNDA.n618 585
R1790 GNDA.n659 GNDA.n643 585
R1791 GNDA.n659 GNDA.n658 585
R1792 GNDA.n647 GNDA.n644 585
R1793 GNDA.n657 GNDA.n644 585
R1794 GNDA.n655 GNDA.n654 585
R1795 GNDA.n656 GNDA.n655 585
R1796 GNDA.n653 GNDA.n646 585
R1797 GNDA.n646 GNDA.n645 585
R1798 GNDA.n652 GNDA.n651 585
R1799 GNDA.n651 GNDA.n650 585
R1800 GNDA.n648 GNDA.n579 585
R1801 GNDA.n649 GNDA.n648 585
R1802 GNDA.n1588 GNDA.n580 585
R1803 GNDA.n1587 GNDA.n581 585
R1804 GNDA.n1584 GNDA.n582 585
R1805 GNDA.n1583 GNDA.n583 585
R1806 GNDA.n1580 GNDA.n584 585
R1807 GNDA.n1579 GNDA.n585 585
R1808 GNDA.n1576 GNDA.n586 585
R1809 GNDA.n1575 GNDA.n587 585
R1810 GNDA.n1572 GNDA.n588 585
R1811 GNDA.n1571 GNDA.n1570 585
R1812 GNDA.n1571 GNDA.n423 585
R1813 GNDA.n1573 GNDA.n1572 585
R1814 GNDA.n1575 GNDA.n1574 585
R1815 GNDA.n1577 GNDA.n1576 585
R1816 GNDA.n1579 GNDA.n1578 585
R1817 GNDA.n1581 GNDA.n1580 585
R1818 GNDA.n1583 GNDA.n1582 585
R1819 GNDA.n1585 GNDA.n1584 585
R1820 GNDA.n1587 GNDA.n1586 585
R1821 GNDA.n1589 GNDA.n1588 585
R1822 GNDA.n1592 GNDA.n1591 585
R1823 GNDA.n1591 GNDA.n1590 585
R1824 GNDA.n1593 GNDA.n577 585
R1825 GNDA.n577 GNDA.n576 585
R1826 GNDA.n1595 GNDA.n1594 585
R1827 GNDA.n1596 GNDA.n1595 585
R1828 GNDA.n575 GNDA.n574 585
R1829 GNDA.n1597 GNDA.n575 585
R1830 GNDA.n1600 GNDA.n1599 585
R1831 GNDA.n1599 GNDA.n1598 585
R1832 GNDA.n1601 GNDA.n567 585
R1833 GNDA.n567 GNDA.n359 585
R1834 GNDA.n1604 GNDA.n1603 585
R1835 GNDA.n1605 GNDA.n1604 585
R1836 GNDA.n566 GNDA.n565 585
R1837 GNDA.n1606 GNDA.n566 585
R1838 GNDA.n1609 GNDA.n1608 585
R1839 GNDA.n1608 GNDA.n1607 585
R1840 GNDA.n1610 GNDA.n564 585
R1841 GNDA.n564 GNDA.n563 585
R1842 GNDA.n1612 GNDA.n1611 585
R1843 GNDA.n1613 GNDA.n1612 585
R1844 GNDA.n561 GNDA.n534 585
R1845 GNDA.n1614 GNDA.n561 585
R1846 GNDA.n1617 GNDA.n1616 585
R1847 GNDA.n1616 GNDA.n1615 585
R1848 GNDA.n1621 GNDA.n1620 585
R1849 GNDA.n1620 GNDA.n1619 585
R1850 GNDA.n1622 GNDA.n533 585
R1851 GNDA.n533 GNDA.n532 585
R1852 GNDA.n1625 GNDA.n1624 585
R1853 GNDA.n1626 GNDA.n1625 585
R1854 GNDA.n1623 GNDA.n531 585
R1855 GNDA.n1627 GNDA.n531 585
R1856 GNDA.n1629 GNDA.n530 585
R1857 GNDA.n1629 GNDA.n1628 585
R1858 GNDA.n1631 GNDA.n1630 585
R1859 GNDA.n1630 GNDA.n95 585
R1860 GNDA.n1632 GNDA.n529 585
R1861 GNDA.n529 GNDA.n96 585
R1862 GNDA.n1634 GNDA.n1633 585
R1863 GNDA.n1635 GNDA.n1634 585
R1864 GNDA.n528 GNDA.n527 585
R1865 GNDA.n1636 GNDA.n528 585
R1866 GNDA.n1640 GNDA.n1639 585
R1867 GNDA.n1639 GNDA.n1638 585
R1868 GNDA.n1641 GNDA.n526 585
R1869 GNDA.n1637 GNDA.n526 585
R1870 GNDA.n1643 GNDA.n1642 585
R1871 GNDA.n1643 GNDA.n516 585
R1872 GNDA.n1866 GNDA.n405 585
R1873 GNDA.n1866 GNDA.n1865 585
R1874 GNDA.n1766 GNDA.n1765 585
R1875 GNDA.n445 GNDA.n444 585
R1876 GNDA.n1837 GNDA.n1836 585
R1877 GNDA.n1840 GNDA.n1839 585
R1878 GNDA.n443 GNDA.n440 585
R1879 GNDA.n436 GNDA.n435 585
R1880 GNDA.n1848 GNDA.n1847 585
R1881 GNDA.n1851 GNDA.n1850 585
R1882 GNDA.n434 GNDA.n431 585
R1883 GNDA.n427 GNDA.n426 585
R1884 GNDA.n1859 GNDA.n1858 585
R1885 GNDA.n1862 GNDA.n1861 585
R1886 GNDA.n807 GNDA.n806 585
R1887 GNDA.n629 GNDA.n625 585
R1888 GNDA.n1563 GNDA.n1562 585
R1889 GNDA.n705 GNDA.n611 585
R1890 GNDA.n776 GNDA.n775 585
R1891 GNDA.n780 GNDA.n779 585
R1892 GNDA.n778 GNDA.n701 585
R1893 GNDA.n787 GNDA.n786 585
R1894 GNDA.n789 GNDA.n788 585
R1895 GNDA.n793 GNDA.n792 585
R1896 GNDA.n791 GNDA.n697 585
R1897 GNDA.n800 GNDA.n799 585
R1898 GNDA.n802 GNDA.n801 585
R1899 GNDA.n805 GNDA.n804 585
R1900 GNDA.n1564 GNDA.n609 585
R1901 GNDA.n609 GNDA.n590 585
R1902 GNDA.n1568 GNDA.n589 585
R1903 GNDA.n1568 GNDA.n1567 585
R1904 GNDA.n1662 GNDA.n1661 585
R1905 GNDA.n510 GNDA.n509 585
R1906 GNDA.n1733 GNDA.n1732 585
R1907 GNDA.n1736 GNDA.n1735 585
R1908 GNDA.n508 GNDA.n505 585
R1909 GNDA.n501 GNDA.n500 585
R1910 GNDA.n1744 GNDA.n1743 585
R1911 GNDA.n1747 GNDA.n1746 585
R1912 GNDA.n499 GNDA.n496 585
R1913 GNDA.n492 GNDA.n491 585
R1914 GNDA.n1755 GNDA.n1754 585
R1915 GNDA.n1758 GNDA.n1757 585
R1916 GNDA.n485 GNDA.n484 585
R1917 GNDA.n482 GNDA.n448 585
R1918 GNDA.n481 GNDA.n480 585
R1919 GNDA.n479 GNDA.n478 585
R1920 GNDA.n477 GNDA.n450 585
R1921 GNDA.n475 GNDA.n474 585
R1922 GNDA.n473 GNDA.n451 585
R1923 GNDA.n472 GNDA.n471 585
R1924 GNDA.n469 GNDA.n452 585
R1925 GNDA.n467 GNDA.n466 585
R1926 GNDA.n465 GNDA.n453 585
R1927 GNDA.n464 GNDA.n463 585
R1928 GNDA.n315 GNDA.n314 585
R1929 GNDA.n318 GNDA.n317 585
R1930 GNDA.n320 GNDA.n319 585
R1931 GNDA.n324 GNDA.n323 585
R1932 GNDA.n322 GNDA.n236 585
R1933 GNDA.n331 GNDA.n330 585
R1934 GNDA.n333 GNDA.n332 585
R1935 GNDA.n337 GNDA.n336 585
R1936 GNDA.n335 GNDA.n232 585
R1937 GNDA.n344 GNDA.n343 585
R1938 GNDA.n346 GNDA.n345 585
R1939 GNDA.n349 GNDA.n348 585
R1940 GNDA.n1966 GNDA.n148 585
R1941 GNDA.n1967 GNDA.n228 585
R1942 GNDA.n1969 GNDA.n1968 585
R1943 GNDA.n1971 GNDA.n226 585
R1944 GNDA.n1974 GNDA.n1973 585
R1945 GNDA.n1975 GNDA.n225 585
R1946 GNDA.n1977 GNDA.n1976 585
R1947 GNDA.n1979 GNDA.n224 585
R1948 GNDA.n1982 GNDA.n1981 585
R1949 GNDA.n1983 GNDA.n223 585
R1950 GNDA.n1985 GNDA.n1984 585
R1951 GNDA.n1987 GNDA.n222 585
R1952 GNDA.n2157 GNDA.n130 585
R1953 GNDA.n542 GNDA.n488 585
R1954 GNDA.n544 GNDA.n543 585
R1955 GNDA.n547 GNDA.n541 585
R1956 GNDA.n548 GNDA.n540 585
R1957 GNDA.n551 GNDA.n539 585
R1958 GNDA.n552 GNDA.n538 585
R1959 GNDA.n555 GNDA.n537 585
R1960 GNDA.n556 GNDA.n536 585
R1961 GNDA.n559 GNDA.n535 585
R1962 GNDA.n560 GNDA.n136 585
R1963 GNDA.n2157 GNDA.n136 585
R1964 GNDA.n2157 GNDA.n129 585
R1965 GNDA.n1367 GNDA.n1365 585
R1966 GNDA.n1368 GNDA.n1364 585
R1967 GNDA.n1371 GNDA.n1363 585
R1968 GNDA.n1372 GNDA.n1362 585
R1969 GNDA.n1375 GNDA.n1361 585
R1970 GNDA.n1376 GNDA.n1360 585
R1971 GNDA.n1379 GNDA.n1359 585
R1972 GNDA.n1380 GNDA.n1358 585
R1973 GNDA.n1383 GNDA.n1357 585
R1974 GNDA.n1384 GNDA.n142 585
R1975 GNDA.n2157 GNDA.n142 585
R1976 GNDA.n2157 GNDA.n128 585
R1977 GNDA.n199 GNDA.n197 585
R1978 GNDA.n196 GNDA.n195 585
R1979 GNDA.n192 GNDA.n191 585
R1980 GNDA.n190 GNDA.n189 585
R1981 GNDA.n186 GNDA.n185 585
R1982 GNDA.n184 GNDA.n183 585
R1983 GNDA.n180 GNDA.n179 585
R1984 GNDA.n178 GNDA.n177 585
R1985 GNDA.n151 GNDA.n149 585
R1986 GNDA.n2156 GNDA.n2155 585
R1987 GNDA.n2157 GNDA.n2156 585
R1988 GNDA.n1764 GNDA.n1762 585
R1989 GNDA.n1764 GNDA.n154 585
R1990 GNDA.n562 GNDA.n560 585
R1991 GNDA.n559 GNDA.n558 585
R1992 GNDA.n557 GNDA.n556 585
R1993 GNDA.n555 GNDA.n554 585
R1994 GNDA.n553 GNDA.n552 585
R1995 GNDA.n551 GNDA.n550 585
R1996 GNDA.n549 GNDA.n548 585
R1997 GNDA.n547 GNDA.n546 585
R1998 GNDA.n545 GNDA.n544 585
R1999 GNDA.n488 GNDA.n487 585
R2000 GNDA.n2152 GNDA.n166 585
R2001 GNDA.n2152 GNDA.n172 585
R2002 GNDA.n1247 GNDA.n1245 585
R2003 GNDA.n1247 GNDA.n154 585
R2004 GNDA.n1386 GNDA.n1356 585
R2005 GNDA.n1386 GNDA.n154 585
R2006 GNDA.n1385 GNDA.n1384 585
R2007 GNDA.n1383 GNDA.n1382 585
R2008 GNDA.n1381 GNDA.n1380 585
R2009 GNDA.n1379 GNDA.n1378 585
R2010 GNDA.n1377 GNDA.n1376 585
R2011 GNDA.n1375 GNDA.n1374 585
R2012 GNDA.n1373 GNDA.n1372 585
R2013 GNDA.n1371 GNDA.n1370 585
R2014 GNDA.n1369 GNDA.n1368 585
R2015 GNDA.n1367 GNDA.n1366 585
R2016 GNDA.n2152 GNDA.n160 585
R2017 GNDA.n2152 GNDA.n173 585
R2018 GNDA.n152 GNDA.n150 585
R2019 GNDA.n154 GNDA.n152 585
R2020 GNDA.n2155 GNDA.n2154 585
R2021 GNDA.n153 GNDA.n151 585
R2022 GNDA.n177 GNDA.n176 585
R2023 GNDA.n181 GNDA.n180 585
R2024 GNDA.n183 GNDA.n182 585
R2025 GNDA.n187 GNDA.n186 585
R2026 GNDA.n189 GNDA.n188 585
R2027 GNDA.n193 GNDA.n192 585
R2028 GNDA.n195 GNDA.n194 585
R2029 GNDA.n199 GNDA.n198 585
R2030 GNDA.n2152 GNDA.n155 585
R2031 GNDA.n2152 GNDA.n2151 585
R2032 GNDA.n2105 GNDA.n2006 585
R2033 GNDA.n2105 GNDA.n2104 585
R2034 GNDA.n2011 GNDA.n2007 585
R2035 GNDA.n2103 GNDA.n2007 585
R2036 GNDA.n2100 GNDA.n2099 585
R2037 GNDA.n2101 GNDA.n2100 585
R2038 GNDA.n2024 GNDA.n2009 585
R2039 GNDA.n2009 GNDA.n2008 585
R2040 GNDA.n2023 GNDA.n2022 585
R2041 GNDA.n2022 GNDA.n2021 585
R2042 GNDA.n2020 GNDA.n2019 585
R2043 GNDA.n2020 GNDA.n212 585
R2044 GNDA.n2014 GNDA.n211 585
R2045 GNDA.n2131 GNDA.n211 585
R2046 GNDA.n2134 GNDA.n2133 585
R2047 GNDA.n2133 GNDA.n2132 585
R2048 GNDA.n207 GNDA.n204 585
R2049 GNDA.n204 GNDA.n203 585
R2050 GNDA.n2141 GNDA.n2140 585
R2051 GNDA.n2142 GNDA.n2141 585
R2052 GNDA.n205 GNDA.n202 585
R2053 GNDA.n2143 GNDA.n202 585
R2054 GNDA.n2146 GNDA.n2145 585
R2055 GNDA.n2145 GNDA.n2144 585
R2056 GNDA.n1944 GNDA.n376 585
R2057 GNDA.n376 GNDA.n375 585
R2058 GNDA.n1947 GNDA.n1946 585
R2059 GNDA.n1948 GNDA.n1947 585
R2060 GNDA.n377 GNDA.n373 585
R2061 GNDA.n1949 GNDA.n373 585
R2062 GNDA.n1952 GNDA.n1951 585
R2063 GNDA.n1951 GNDA.n1950 585
R2064 GNDA.n369 GNDA.n367 585
R2065 GNDA.n367 GNDA.n365 585
R2066 GNDA.n1959 GNDA.n1958 585
R2067 GNDA.n1960 GNDA.n1959 585
R2068 GNDA.n1876 GNDA.n366 585
R2069 GNDA.n366 GNDA.n364 585
R2070 GNDA.n1883 GNDA.n1882 585
R2071 GNDA.n1884 GNDA.n1883 585
R2072 GNDA.n1874 GNDA.n400 585
R2073 GNDA.n1885 GNDA.n400 585
R2074 GNDA.n1888 GNDA.n1887 585
R2075 GNDA.n1887 GNDA.n1886 585
R2076 GNDA.n399 GNDA.n397 585
R2077 GNDA.n1873 GNDA.n399 585
R2078 GNDA.n1871 GNDA.n1870 585
R2079 GNDA.n1872 GNDA.n1871 585
R2080 GNDA.n175 GNDA.n174 585
R2081 GNDA.n374 GNDA.n174 585
R2082 GNDA.n1034 GNDA.n958 585
R2083 GNDA.n1030 GNDA.n958 585
R2084 GNDA.n1037 GNDA.n1036 585
R2085 GNDA.n1038 GNDA.n1037 585
R2086 GNDA.n959 GNDA.n860 585
R2087 GNDA.n1039 GNDA.n860 585
R2088 GNDA.n1042 GNDA.n1041 585
R2089 GNDA.n1041 GNDA.n1040 585
R2090 GNDA.n859 GNDA.n857 585
R2091 GNDA.n861 GNDA.n859 585
R2092 GNDA.n853 GNDA.n852 585
R2093 GNDA.n852 GNDA.n623 585
R2094 GNDA.n1050 GNDA.n1049 585
R2095 GNDA.n1050 GNDA.n622 585
R2096 GNDA.n1057 GNDA.n1056 585
R2097 GNDA.n1056 GNDA.n1055 585
R2098 GNDA.n851 GNDA.n849 585
R2099 GNDA.n1054 GNDA.n851 585
R2100 GNDA.n1052 GNDA.n845 585
R2101 GNDA.n1053 GNDA.n1052 585
R2102 GNDA.n1064 GNDA.n843 585
R2103 GNDA.n1051 GNDA.n843 585
R2104 GNDA.n1067 GNDA.n1066 585
R2105 GNDA.n1067 GNDA.n842 585
R2106 GNDA.n1033 GNDA.n1032 585
R2107 GNDA.n1032 GNDA.n1031 585
R2108 GNDA.n1660 GNDA.n512 585
R2109 GNDA.n1660 GNDA.n123 585
R2110 GNDA.n1644 GNDA.n518 585
R2111 GNDA.n1645 GNDA.n1644 585
R2112 GNDA.n525 GNDA.n524 585
R2113 GNDA.n525 GNDA.n517 585
R2114 GNDA.n523 GNDA.n522 585
R2115 GNDA.n522 GNDA.n521 585
R2116 GNDA.n92 GNDA.n90 585
R2117 GNDA.n90 GNDA.n88 585
R2118 GNDA.n2188 GNDA.n2187 585
R2119 GNDA.n2189 GNDA.n2188 585
R2120 GNDA.n2186 GNDA.n91 585
R2121 GNDA.n91 GNDA.n89 585
R2122 GNDA.n2185 GNDA.n2184 585
R2123 GNDA.n2184 GNDA.n2183 585
R2124 GNDA.n94 GNDA.n93 585
R2125 GNDA.n2182 GNDA.n94 585
R2126 GNDA.n2180 GNDA.n2179 585
R2127 GNDA.n2181 GNDA.n2180 585
R2128 GNDA.n2178 GNDA.n99 585
R2129 GNDA.n99 GNDA.n98 585
R2130 GNDA.n2177 GNDA.n2176 585
R2131 GNDA.n2176 GNDA.n2175 585
R2132 GNDA.n1657 GNDA.n101 585
R2133 GNDA.n1659 GNDA.n1658 585
R2134 GNDA.n313 GNDA.n309 585
R2135 GNDA.n313 GNDA.n125 585
R2136 GNDA.n461 GNDA.n454 585
R2137 GNDA.n461 GNDA.n122 585
R2138 GNDA.n460 GNDA.n457 585
R2139 GNDA.n460 GNDA.n459 585
R2140 GNDA.n456 GNDA.n455 585
R2141 GNDA.n458 GNDA.n455 585
R2142 GNDA.n113 GNDA.n111 585
R2143 GNDA.n111 GNDA.n109 585
R2144 GNDA.n2164 GNDA.n2163 585
R2145 GNDA.n2165 GNDA.n2164 585
R2146 GNDA.n2162 GNDA.n112 585
R2147 GNDA.n112 GNDA.n110 585
R2148 GNDA.n2161 GNDA.n2160 585
R2149 GNDA.n2160 GNDA.n2159 585
R2150 GNDA.n114 GNDA.n75 585
R2151 GNDA.n75 GNDA.n73 585
R2152 GNDA.n2310 GNDA.n2309 585
R2153 GNDA.n2311 GNDA.n2310 585
R2154 GNDA.n2308 GNDA.n76 585
R2155 GNDA.n79 GNDA.n76 585
R2156 GNDA.n2307 GNDA.n2306 585
R2157 GNDA.n2306 GNDA.n2305 585
R2158 GNDA.n80 GNDA.n78 585
R2159 GNDA.n312 GNDA.n311 585
R2160 GNDA.n2118 GNDA.n2117 585
R2161 GNDA.n2117 GNDA.n2116 585
R2162 GNDA.n1988 GNDA.n221 585
R2163 GNDA.n1989 GNDA.n1988 585
R2164 GNDA.n1992 GNDA.n1991 585
R2165 GNDA.n1991 GNDA.n1990 585
R2166 GNDA.n1993 GNDA.n220 585
R2167 GNDA.n220 GNDA.n219 585
R2168 GNDA.n1995 GNDA.n1994 585
R2169 GNDA.n1996 GNDA.n1995 585
R2170 GNDA.n218 GNDA.n217 585
R2171 GNDA.n1997 GNDA.n218 585
R2172 GNDA.n2000 GNDA.n1999 585
R2173 GNDA.n1999 GNDA.n1998 585
R2174 GNDA.n2001 GNDA.n215 585
R2175 GNDA.n215 GNDA.n213 585
R2176 GNDA.n2129 GNDA.n2128 585
R2177 GNDA.n2130 GNDA.n2129 585
R2178 GNDA.n2127 GNDA.n216 585
R2179 GNDA.n216 GNDA.n214 585
R2180 GNDA.n2126 GNDA.n2125 585
R2181 GNDA.n2125 GNDA.n2124 585
R2182 GNDA.n2003 GNDA.n2002 585
R2183 GNDA.n2123 GNDA.n2003 585
R2184 GNDA.n2122 GNDA.n2121 585
R2185 GNDA.n2005 GNDA.n2004 585
R2186 GNDA.n674 GNDA.n673 579.628
R2187 GNDA.n957 GNDA.n956 556.322
R2188 GNDA.n2362 GNDA.t244 535.191
R2189 GNDA.n2389 GNDA.t259 535.191
R2190 GNDA.n2202 GNDA.t312 535.191
R2191 GNDA.n2256 GNDA.t300 535.191
R2192 GNDA.n2446 GNDA.n39 531.201
R2193 GNDA.n2301 GNDA.n2300 531.201
R2194 GNDA.n2300 GNDA.n83 528
R2195 GNDA.t250 GNDA.n621 512.884
R2196 GNDA.n675 GNDA.n674 512.29
R2197 GNDA.n675 GNDA.n634 512.29
R2198 GNDA.n681 GNDA.n634 512.29
R2199 GNDA.n682 GNDA.n681 512.29
R2200 GNDA.n683 GNDA.n682 512.29
R2201 GNDA.n689 GNDA.n630 512.29
R2202 GNDA.n690 GNDA.n689 512.29
R2203 GNDA.n691 GNDA.n690 512.29
R2204 GNDA.n691 GNDA.n625 512.29
R2205 GNDA.n807 GNDA.n625 512.29
R2206 GNDA.n1559 GNDA.n808 512.29
R2207 GNDA.n1553 GNDA.n808 512.29
R2208 GNDA.n1553 GNDA.n1552 512.29
R2209 GNDA.n1552 GNDA.n1551 512.29
R2210 GNDA.n1551 GNDA.n814 512.29
R2211 GNDA.n1545 GNDA.n1544 512.29
R2212 GNDA.n1544 GNDA.n1543 512.29
R2213 GNDA.n1543 GNDA.n818 512.29
R2214 GNDA.n825 GNDA.n818 512.29
R2215 GNDA.n826 GNDA.n825 512.29
R2216 GNDA.n1088 GNDA.n833 512.29
R2217 GNDA.n1088 GNDA.n1087 512.29
R2218 GNDA.n1087 GNDA.n1086 512.29
R2219 GNDA.n1086 GNDA.n834 512.29
R2220 GNDA.n1080 GNDA.n834 512.29
R2221 GNDA.n1079 GNDA.n1078 512.29
R2222 GNDA.n1078 GNDA.n838 512.29
R2223 GNDA.n1072 GNDA.n838 512.29
R2224 GNDA.n1072 GNDA.n1071 512.29
R2225 GNDA.n1071 GNDA.n1070 512.29
R2226 GNDA.n2333 GNDA.n55 512
R2227 GNDA.n2335 GNDA.n55 512
R2228 GNDA.n952 GNDA.n865 512
R2229 GNDA.n954 GNDA.n865 512
R2230 GNDA.n2334 GNDA.n2333 508.8
R2231 GNDA.n2335 GNDA.n2334 508.8
R2232 GNDA.n953 GNDA.n952 508.8
R2233 GNDA.n954 GNDA.n953 508.8
R2234 GNDA.n2302 GNDA.n2301 499.2
R2235 GNDA.n2422 GNDA.n2394 496
R2236 GNDA.n2262 GNDA.n2199 496
R2237 GNDA.n8 GNDA.t330 493.418
R2238 GNDA.n12 GNDA.t309 493.418
R2239 GNDA.n11 GNDA.t327 493.418
R2240 GNDA.n10 GNDA.t306 493.418
R2241 GNDA.n2482 GNDA.t334 493.418
R2242 GNDA.n2483 GNDA.t315 493.418
R2243 GNDA.n20 GNDA.t297 493.418
R2244 GNDA.n18 GNDA.t247 493.418
R2245 GNDA.n2478 GNDA.t236 493.418
R2246 GNDA.n2477 GNDA.t321 493.418
R2247 GNDA.n2423 GNDA.n2422 489.601
R2248 GNDA.n2262 GNDA.n2198 489.601
R2249 GNDA.n83 GNDA.n69 486.401
R2250 GNDA.n2347 GNDA.n2346 476.8
R2251 GNDA.n2238 GNDA.n2219 476.8
R2252 GNDA.n2431 GNDA.n2345 448
R2253 GNDA.n2235 GNDA.n2231 448
R2254 GNDA.n1653 GNDA.n1652 444.8
R2255 GNDA.n1652 GNDA.n1651 444.8
R2256 GNDA.n1654 GNDA.n1653 441.601
R2257 GNDA.n1651 GNDA.n1650 438.401
R2258 GNDA.n71 GNDA.n67 435.2
R2259 GNDA.n1031 GNDA.n401 434.906
R2260 GNDA.n374 GNDA.n127 434.906
R2261 GNDA.n2450 GNDA.n40 428.8
R2262 GNDA.n2315 GNDA.n67 425.601
R2263 GNDA.n2314 GNDA.n70 422.401
R2264 GNDA.n16 GNDA.n15 422.401
R2265 GNDA.n13 GNDA.n9 422.401
R2266 GNDA.n2485 GNDA.n2484 422.401
R2267 GNDA.n2480 GNDA.n2479 422.401
R2268 GNDA.n2315 GNDA.n2314 419.2
R2269 GNDA.n2342 GNDA.n2341 418.483
R2270 GNDA.n884 GNDA.t294 413.084
R2271 GNDA.n881 GNDA.t289 413.084
R2272 GNDA.n880 GNDA.t286 413.084
R2273 GNDA.n878 GNDA.t268 413.084
R2274 GNDA.n918 GNDA.t303 413.084
R2275 GNDA.n928 GNDA.t324 413.084
R2276 GNDA.n2227 GNDA.n2191 411.512
R2277 GNDA.t250 GNDA.n620 391.411
R2278 GNDA.n2357 GNDA.n2350 387.2
R2279 GNDA.n2254 GNDA.n2253 387.2
R2280 GNDA.n59 GNDA.n57 383.118
R2281 GNDA.n2428 GNDA.n2350 380.8
R2282 GNDA.n2254 GNDA.n2204 380.8
R2283 GNDA.n2291 GNDA.n2290 368.283
R2284 GNDA.n2451 GNDA.n2450 355.2
R2285 GNDA.n927 GNDA.n862 354.024
R2286 GNDA.n1051 GNDA.n842 352.627
R2287 GNDA.n1053 GNDA.n1051 352.627
R2288 GNDA.n1054 GNDA.n1053 352.627
R2289 GNDA.n1055 GNDA.n1054 352.627
R2290 GNDA.n1055 GNDA.n622 352.627
R2291 GNDA.n861 GNDA.n623 352.627
R2292 GNDA.n1040 GNDA.n861 352.627
R2293 GNDA.n1040 GNDA.n1039 352.627
R2294 GNDA.n1039 GNDA.n1038 352.627
R2295 GNDA.n1031 GNDA.n1030 352.627
R2296 GNDA.n1873 GNDA.n1872 352.627
R2297 GNDA.n1886 GNDA.n1873 352.627
R2298 GNDA.n1886 GNDA.n1885 352.627
R2299 GNDA.n1885 GNDA.n1884 352.627
R2300 GNDA.n1884 GNDA.n364 352.627
R2301 GNDA.n1960 GNDA.n365 352.627
R2302 GNDA.n1950 GNDA.n365 352.627
R2303 GNDA.n1950 GNDA.n1949 352.627
R2304 GNDA.n1949 GNDA.n1948 352.627
R2305 GNDA.n1948 GNDA.n375 352.627
R2306 GNDA.n375 GNDA.n374 352.627
R2307 GNDA.n2144 GNDA.n2143 352.627
R2308 GNDA.n2143 GNDA.n2142 352.627
R2309 GNDA.n2142 GNDA.n203 352.627
R2310 GNDA.n2132 GNDA.n203 352.627
R2311 GNDA.n2132 GNDA.n2131 352.627
R2312 GNDA.n2021 GNDA.n212 352.627
R2313 GNDA.n2021 GNDA.n2008 352.627
R2314 GNDA.n2101 GNDA.n2008 352.627
R2315 GNDA.n2104 GNDA.n2103 352.627
R2316 GNDA.n2431 GNDA.n2430 342.401
R2317 GNDA.n2236 GNDA.n2235 342.401
R2318 GNDA.n911 GNDA.n52 341.38
R2319 GNDA.n2367 GNDA.n2364 332.8
R2320 GNDA.n2243 GNDA.n2215 332.8
R2321 GNDA.n27 GNDA.t277 332.75
R2322 GNDA.n29 GNDA.t262 332.75
R2323 GNDA.t252 GNDA.n361 172.876
R2324 GNDA.t252 GNDA.n362 172.876
R2325 GNDA.t243 GNDA.n97 172.876
R2326 GNDA.t243 GNDA.n2158 172.876
R2327 GNDA.n1961 GNDA.t252 172.615
R2328 GNDA.t252 GNDA.n363 172.615
R2329 GNDA.t243 GNDA.n115 172.615
R2330 GNDA.t243 GNDA.n126 172.615
R2331 GNDA.n926 GNDA.n925 323.2
R2332 GNDA.n59 GNDA.n58 322.861
R2333 GNDA.n2387 GNDA.n2365 321.281
R2334 GNDA.n2245 GNDA.n2244 321.281
R2335 GNDA.n2367 GNDA.n2365 318.08
R2336 GNDA.n2244 GNDA.n2243 318.08
R2337 GNDA.n926 GNDA.n60 316.8
R2338 GNDA.n2394 GNDA.n2392 310.401
R2339 GNDA.n2257 GNDA.n2199 310.401
R2340 GNDA.n2113 GNDA.n2112 304
R2341 GNDA.n2423 GNDA.n2363 304
R2342 GNDA.n2203 GNDA.n2198 304
R2343 GNDA.n2474 GNDA.n2473 300.8
R2344 GNDA.n2473 GNDA.n2462 300.8
R2345 GNDA.n2112 GNDA.n2111 300.8
R2346 GNDA.n2113 GNDA.n2109 300.8
R2347 GNDA.n2388 GNDA.n2364 300.8
R2348 GNDA.n2215 GNDA.n2214 300.8
R2349 GNDA.n2172 GNDA.n2171 297.601
R2350 GNDA.n2171 GNDA.n2170 297.601
R2351 GNDA.n2111 GNDA.n2109 297.601
R2352 GNDA.n2169 GNDA.n2168 297.601
R2353 GNDA.n2168 GNDA.n66 297.601
R2354 GNDA.n2381 GNDA.n2380 296
R2355 GNDA.n2229 GNDA.n2221 296
R2356 GNDA.n945 GNDA.n944 294.401
R2357 GNDA.n944 GNDA.n943 294.401
R2358 GNDA.n925 GNDA.n924 294.401
R2359 GNDA.n937 GNDA.n60 292.5
R2360 GNDA.n938 GNDA.n937 292.5
R2361 GNDA.n936 GNDA.n926 292.5
R2362 GNDA.n936 GNDA.n935 292.5
R2363 GNDA.n925 GNDA.n923 292.5
R2364 GNDA.n927 GNDA.n923 292.5
R2365 GNDA.n924 GNDA.n922 292.5
R2366 GNDA.n935 GNDA.n922 292.5
R2367 GNDA.n911 GNDA.n57 292.5
R2368 GNDA.n910 GNDA.n58 292.5
R2369 GNDA.n2329 GNDA.n2328 292.5
R2370 GNDA.n2330 GNDA.n2329 292.5
R2371 GNDA.n2336 GNDA.n2335 292.5
R2372 GNDA.n2337 GNDA.n2336 292.5
R2373 GNDA.n2334 GNDA.n54 292.5
R2374 GNDA.n910 GNDA.n54 292.5
R2375 GNDA.n2333 GNDA.n2332 292.5
R2376 GNDA.n2332 GNDA.n2331 292.5
R2377 GNDA.n55 GNDA.n53 292.5
R2378 GNDA.n910 GNDA.n53 292.5
R2379 GNDA.n873 GNDA.n871 292.5
R2380 GNDA.n871 GNDA.n52 292.5
R2381 GNDA.n869 GNDA.n61 292.5
R2382 GNDA.n949 GNDA.n869 292.5
R2383 GNDA.n872 GNDA.n870 292.5
R2384 GNDA.n870 GNDA.n862 292.5
R2385 GNDA.n875 GNDA.n874 292.5
R2386 GNDA.n949 GNDA.n875 292.5
R2387 GNDA.n942 GNDA.n941 292.5
R2388 GNDA.n941 GNDA.n940 292.5
R2389 GNDA.n933 GNDA.n920 292.5
R2390 GNDA.n934 GNDA.n933 292.5
R2391 GNDA.n931 GNDA.n930 292.5
R2392 GNDA.n932 GNDA.n931 292.5
R2393 GNDA.n945 GNDA.n877 292.5
R2394 GNDA.n877 GNDA.n56 292.5
R2395 GNDA.n944 GNDA.n868 292.5
R2396 GNDA.n949 GNDA.n868 292.5
R2397 GNDA.n943 GNDA.n876 292.5
R2398 GNDA.n939 GNDA.n876 292.5
R2399 GNDA.n948 GNDA.n947 292.5
R2400 GNDA.n949 GNDA.n948 292.5
R2401 GNDA.n912 GNDA.n907 292.5
R2402 GNDA.n913 GNDA.n912 292.5
R2403 GNDA.n916 GNDA.n915 292.5
R2404 GNDA.n915 GNDA.n914 292.5
R2405 GNDA.n917 GNDA.n883 292.5
R2406 GNDA.n909 GNDA.n883 292.5
R2407 GNDA.n952 GNDA.n951 292.5
R2408 GNDA.n951 GNDA.n950 292.5
R2409 GNDA.n953 GNDA.n864 292.5
R2410 GNDA.n935 GNDA.n864 292.5
R2411 GNDA.n955 GNDA.n954 292.5
R2412 GNDA.n956 GNDA.n955 292.5
R2413 GNDA.n865 GNDA.n863 292.5
R2414 GNDA.n935 GNDA.n863 292.5
R2415 GNDA.n1653 GNDA.n1649 292.5
R2416 GNDA.n1649 GNDA.n74 292.5
R2417 GNDA.n1652 GNDA.n515 292.5
R2418 GNDA.n1656 GNDA.n515 292.5
R2419 GNDA.n1651 GNDA.n1648 292.5
R2420 GNDA.n1648 GNDA.n1647 292.5
R2421 GNDA.n1655 GNDA.n1654 292.5
R2422 GNDA.n1656 GNDA.n1655 292.5
R2423 GNDA.n2314 GNDA.n2313 292.5
R2424 GNDA.n2313 GNDA.n2312 292.5
R2425 GNDA.n72 GNDA.n71 292.5
R2426 GNDA.n2174 GNDA.n72 292.5
R2427 GNDA.n1646 GNDA.n67 292.5
R2428 GNDA.n1647 GNDA.n1646 292.5
R2429 GNDA.n2315 GNDA.n68 292.5
R2430 GNDA.n2174 GNDA.n68 292.5
R2431 GNDA.n2300 GNDA.n2299 292.5
R2432 GNDA.n2299 GNDA.n2298 292.5
R2433 GNDA.n2301 GNDA.n82 292.5
R2434 GNDA.n2107 GNDA.n82 292.5
R2435 GNDA.n2303 GNDA.n2302 292.5
R2436 GNDA.n2304 GNDA.n2303 292.5
R2437 GNDA.n83 GNDA.n81 292.5
R2438 GNDA.n2107 GNDA.n81 292.5
R2439 GNDA.n2168 GNDA.n2167 292.5
R2440 GNDA.n2167 GNDA.n2166 292.5
R2441 GNDA.n103 GNDA.n66 292.5
R2442 GNDA.n2174 GNDA.n103 292.5
R2443 GNDA.n519 GNDA.n108 292.5
R2444 GNDA.n520 GNDA.n519 292.5
R2445 GNDA.n2169 GNDA.n104 292.5
R2446 GNDA.n2174 GNDA.n104 292.5
R2447 GNDA.n2114 GNDA.n2113 292.5
R2448 GNDA.n2115 GNDA.n2114 292.5
R2449 GNDA.n2112 GNDA.n2108 292.5
R2450 GNDA.n2108 GNDA.n2107 292.5
R2451 GNDA.n2111 GNDA.n2110 292.5
R2452 GNDA.n2110 GNDA.n124 292.5
R2453 GNDA.n2109 GNDA.n2106 292.5
R2454 GNDA.n2107 GNDA.n2106 292.5
R2455 GNDA.n2171 GNDA.n106 292.5
R2456 GNDA.n2166 GNDA.n106 292.5
R2457 GNDA.n2170 GNDA.n102 292.5
R2458 GNDA.n2174 GNDA.n102 292.5
R2459 GNDA.n107 GNDA.n105 292.5
R2460 GNDA.n520 GNDA.n105 292.5
R2461 GNDA.n2173 GNDA.n2172 292.5
R2462 GNDA.n2174 GNDA.n2173 292.5
R2463 GNDA.n2428 GNDA.n2427 292.5
R2464 GNDA.n2427 GNDA.n2426 292.5
R2465 GNDA.n2352 GNDA.n2350 292.5
R2466 GNDA.t340 GNDA.n2352 292.5
R2467 GNDA.n2358 GNDA.n2357 292.5
R2468 GNDA.n2359 GNDA.n2358 292.5
R2469 GNDA.n2355 GNDA.n2351 292.5
R2470 GNDA.t340 GNDA.n2351 292.5
R2471 GNDA.n2432 GNDA.n2431 292.5
R2472 GNDA.n2433 GNDA.n2432 292.5
R2473 GNDA.n2430 GNDA.n2344 292.5
R2474 GNDA.n2377 GNDA.n2344 292.5
R2475 GNDA.n2372 GNDA.n2347 292.5
R2476 GNDA.n2373 GNDA.n2372 292.5
R2477 GNDA.n2346 GNDA.n2343 292.5
R2478 GNDA.n2377 GNDA.n2343 292.5
R2479 GNDA.n2380 GNDA.n2379 292.5
R2480 GNDA.n2379 GNDA.n2378 292.5
R2481 GNDA.n2366 GNDA.n2364 292.5
R2482 GNDA.n2384 GNDA.n2366 292.5
R2483 GNDA.n2368 GNDA.n2367 292.5
R2484 GNDA.n2374 GNDA.n2368 292.5
R2485 GNDA.n2385 GNDA.n2365 292.5
R2486 GNDA.n2385 GNDA.n2384 292.5
R2487 GNDA.n2387 GNDA.n2386 292.5
R2488 GNDA.n2386 GNDA.n45 292.5
R2489 GNDA.n2424 GNDA.n2423 292.5
R2490 GNDA.n2425 GNDA.n2424 292.5
R2491 GNDA.n2391 GNDA.n2353 292.5
R2492 GNDA.n2360 GNDA.n2353 292.5
R2493 GNDA.n2394 GNDA.n2393 292.5
R2494 GNDA.n2393 GNDA.n44 292.5
R2495 GNDA.n2422 GNDA.n2361 292.5
R2496 GNDA.n2361 GNDA.n2360 292.5
R2497 GNDA.n2246 GNDA.n2245 292.5
R2498 GNDA.n2247 GNDA.n2246 292.5
R2499 GNDA.n2244 GNDA.n2213 292.5
R2500 GNDA.n2216 GNDA.n2213 292.5
R2501 GNDA.n2243 GNDA.n2242 292.5
R2502 GNDA.n2242 GNDA.n2241 292.5
R2503 GNDA.n2215 GNDA.n2212 292.5
R2504 GNDA.n2216 GNDA.n2212 292.5
R2505 GNDA.n2201 GNDA.n2199 292.5
R2506 GNDA.n2201 GNDA.n2192 292.5
R2507 GNDA.n2262 GNDA.n2261 292.5
R2508 GNDA.n2261 GNDA.n2260 292.5
R2509 GNDA.n2200 GNDA.n2198 292.5
R2510 GNDA.n2249 GNDA.n2200 292.5
R2511 GNDA.n2259 GNDA.n2258 292.5
R2512 GNDA.n2260 GNDA.n2259 292.5
R2513 GNDA.n2253 GNDA.n2252 292.5
R2514 GNDA.n2252 GNDA.n2251 292.5
R2515 GNDA.n2254 GNDA.n2205 292.5
R2516 GNDA.t136 GNDA.n2205 292.5
R2517 GNDA.n2208 GNDA.n2204 292.5
R2518 GNDA.n2248 GNDA.n2208 292.5
R2519 GNDA.n2250 GNDA.n2211 292.5
R2520 GNDA.n2250 GNDA.t136 292.5
R2521 GNDA.n2235 GNDA.n2234 292.5
R2522 GNDA.n2234 GNDA.n2233 292.5
R2523 GNDA.n2236 GNDA.n2218 292.5
R2524 GNDA.n2232 GNDA.n2218 292.5
R2525 GNDA.n2239 GNDA.n2238 292.5
R2526 GNDA.n2240 GNDA.n2239 292.5
R2527 GNDA.n2219 GNDA.n2217 292.5
R2528 GNDA.n2226 GNDA.n2217 292.5
R2529 GNDA.n2229 GNDA.n2228 292.5
R2530 GNDA.n2228 GNDA.n2227 292.5
R2531 GNDA.n2475 GNDA.n2474 292.5
R2532 GNDA.n2476 GNDA.n2475 292.5
R2533 GNDA.n2473 GNDA.n26 292.5
R2534 GNDA.n41 GNDA.n26 292.5
R2535 GNDA.n2462 GNDA.n2461 292.5
R2536 GNDA.n2461 GNDA.n2460 292.5
R2537 GNDA.n30 GNDA.n25 292.5
R2538 GNDA.n41 GNDA.n25 292.5
R2539 GNDA.n2498 GNDA.n2497 292.5
R2540 GNDA.n2497 GNDA.n2496 292.5
R2541 GNDA.n5 GNDA.n2 292.5
R2542 GNDA.n2441 GNDA.n5 292.5
R2543 GNDA.n2443 GNDA.n2442 292.5
R2544 GNDA.n2444 GNDA.n2443 292.5
R2545 GNDA.n4 GNDA.n3 292.5
R2546 GNDA.n2441 GNDA.n4 292.5
R2547 GNDA.n2458 GNDA.n2457 292.5
R2548 GNDA.n2459 GNDA.n2458 292.5
R2549 GNDA.n35 GNDA.n33 292.5
R2550 GNDA.n2193 GNDA.n33 292.5
R2551 GNDA.n2283 GNDA.n2282 292.5
R2552 GNDA.n2284 GNDA.n2283 292.5
R2553 GNDA.n34 GNDA.n32 292.5
R2554 GNDA.n2193 GNDA.n32 292.5
R2555 GNDA.n2445 GNDA.n2440 292.5
R2556 GNDA.n2440 GNDA.n2439 292.5
R2557 GNDA.n2450 GNDA.n2449 292.5
R2558 GNDA.n2449 GNDA.n2448 292.5
R2559 GNDA.n43 GNDA.n39 292.5
R2560 GNDA.n43 GNDA.n42 292.5
R2561 GNDA.n2447 GNDA.n2446 292.5
R2562 GNDA.n2448 GNDA.n2447 292.5
R2563 GNDA.n2494 GNDA.n2493 292.5
R2564 GNDA.n2495 GNDA.n2494 292.5
R2565 GNDA.n14 GNDA.n6 292.5
R2566 GNDA.n2489 GNDA.n6 292.5
R2567 GNDA.n2194 GNDA.n17 292.5
R2568 GNDA.n2195 GNDA.n2194 292.5
R2569 GNDA.n2492 GNDA.n7 292.5
R2570 GNDA.n2489 GNDA.n7 292.5
R2571 GNDA.n2491 GNDA.n2490 292.5
R2572 GNDA.n2490 GNDA.n2489 292.5
R2573 GNDA.n2481 GNDA.n22 292.5
R2574 GNDA.n2285 GNDA.n22 292.5
R2575 GNDA.n2488 GNDA.n2487 292.5
R2576 GNDA.n2489 GNDA.n2488 292.5
R2577 GNDA.n2486 GNDA.n23 292.5
R2578 GNDA.n2438 GNDA.n23 292.5
R2579 GNDA.n2172 GNDA.n107 291.2
R2580 GNDA.n2170 GNDA.n107 291.2
R2581 GNDA.n2169 GNDA.n108 291.2
R2582 GNDA.n108 GNDA.n66 291.2
R2583 GNDA.n924 GNDA.n60 288
R2584 GNDA.n885 GNDA.n882 281.601
R2585 GNDA.n929 GNDA.n919 281.601
R2586 GNDA.n916 GNDA.n907 278.401
R2587 GNDA.n930 GNDA.n920 278.401
R2588 GNDA.n683 GNDA.t250 267.529
R2589 GNDA.t250 GNDA.n814 267.529
R2590 GNDA.n1080 GNDA.t250 267.529
R2591 GNDA.n2337 GNDA.n52 265.517
R2592 GNDA.n2145 GNDA.n128 259.416
R2593 GNDA.n348 GNDA.n129 259.416
R2594 GNDA.n1757 GNDA.n130 259.416
R2595 GNDA.n1537 GNDA.n822 259.416
R2596 GNDA.n1069 GNDA.n1067 259.416
R2597 GNDA.n1871 GNDA.n402 259.416
R2598 GNDA.n1344 GNDA.n411 259.416
R2599 GNDA.n806 GNDA.n805 259.416
R2600 GNDA.n1861 GNDA.n405 259.416
R2601 GNDA.n27 GNDA.t278 258.601
R2602 GNDA.n29 GNDA.t264 258.601
R2603 GNDA.n2103 GNDA.n2102 254.675
R2604 GNDA.n1068 GNDA.n840 254.494
R2605 GNDA.n1539 GNDA.n820 254.392
R2606 GNDA.n694 GNDA.n626 254.392
R2607 GNDA.n1961 GNDA.n358 254.34
R2608 GNDA.n1961 GNDA.n357 254.34
R2609 GNDA.n1961 GNDA.n356 254.34
R2610 GNDA.n1961 GNDA.n355 254.34
R2611 GNDA.n1961 GNDA.n354 254.34
R2612 GNDA.n1962 GNDA.n1961 254.34
R2613 GNDA.n1869 GNDA.n1868 254.34
R2614 GNDA.n1867 GNDA.n1866 254.34
R2615 GNDA.n1866 GNDA.n412 254.34
R2616 GNDA.n1866 GNDA.n413 254.34
R2617 GNDA.n1866 GNDA.n414 254.34
R2618 GNDA.n1866 GNDA.n415 254.34
R2619 GNDA.n1568 GNDA.n606 254.34
R2620 GNDA.n1568 GNDA.n605 254.34
R2621 GNDA.n1568 GNDA.n604 254.34
R2622 GNDA.n1568 GNDA.n603 254.34
R2623 GNDA.n1568 GNDA.n602 254.34
R2624 GNDA.n1029 GNDA.n1028 254.34
R2625 GNDA.n1406 GNDA.n363 254.34
R2626 GNDA.n1403 GNDA.n363 254.34
R2627 GNDA.n1352 GNDA.n363 254.34
R2628 GNDA.n1396 GNDA.n363 254.34
R2629 GNDA.n1355 GNDA.n363 254.34
R2630 GNDA.n1389 GNDA.n363 254.34
R2631 GNDA.n1346 GNDA.n1220 254.34
R2632 GNDA.n1866 GNDA.n417 254.34
R2633 GNDA.n1246 GNDA.n361 254.34
R2634 GNDA.n1321 GNDA.n361 254.34
R2635 GNDA.n1238 GNDA.n361 254.34
R2636 GNDA.n1332 GNDA.n361 254.34
R2637 GNDA.n1229 GNDA.n361 254.34
R2638 GNDA.n1343 GNDA.n361 254.34
R2639 GNDA.n1219 GNDA.n1218 254.34
R2640 GNDA.n1568 GNDA.n600 254.34
R2641 GNDA.n1866 GNDA.n418 254.34
R2642 GNDA.n1866 GNDA.n419 254.34
R2643 GNDA.n1866 GNDA.n420 254.34
R2644 GNDA.n1866 GNDA.n421 254.34
R2645 GNDA.n1568 GNDA.n599 254.34
R2646 GNDA.n1568 GNDA.n598 254.34
R2647 GNDA.n1568 GNDA.n597 254.34
R2648 GNDA.n1568 GNDA.n596 254.34
R2649 GNDA.n1415 GNDA.n624 254.34
R2650 GNDA.n1420 GNDA.n624 254.34
R2651 GNDA.n1422 GNDA.n624 254.34
R2652 GNDA.n1428 GNDA.n624 254.34
R2653 GNDA.n1430 GNDA.n624 254.34
R2654 GNDA.n1436 GNDA.n624 254.34
R2655 GNDA.n1568 GNDA.n594 254.34
R2656 GNDA.n1568 GNDA.n593 254.34
R2657 GNDA.n1568 GNDA.n592 254.34
R2658 GNDA.n1568 GNDA.n591 254.34
R2659 GNDA.n1569 GNDA.n1568 254.34
R2660 GNDA.n1866 GNDA.n410 254.34
R2661 GNDA.n1866 GNDA.n409 254.34
R2662 GNDA.n1866 GNDA.n408 254.34
R2663 GNDA.n1866 GNDA.n407 254.34
R2664 GNDA.n1866 GNDA.n406 254.34
R2665 GNDA.n1864 GNDA.n1863 254.34
R2666 GNDA.n1763 GNDA.n362 254.34
R2667 GNDA.n1838 GNDA.n362 254.34
R2668 GNDA.n442 GNDA.n362 254.34
R2669 GNDA.n1849 GNDA.n362 254.34
R2670 GNDA.n433 GNDA.n362 254.34
R2671 GNDA.n1860 GNDA.n362 254.34
R2672 GNDA.n1561 GNDA.n1560 254.34
R2673 GNDA.n1560 GNDA.n616 254.34
R2674 GNDA.n1560 GNDA.n615 254.34
R2675 GNDA.n1560 GNDA.n614 254.34
R2676 GNDA.n1560 GNDA.n613 254.34
R2677 GNDA.n1560 GNDA.n612 254.34
R2678 GNDA.n1566 GNDA.n1565 254.34
R2679 GNDA.n513 GNDA.n97 254.34
R2680 GNDA.n1734 GNDA.n97 254.34
R2681 GNDA.n507 GNDA.n97 254.34
R2682 GNDA.n1745 GNDA.n97 254.34
R2683 GNDA.n498 GNDA.n97 254.34
R2684 GNDA.n1756 GNDA.n97 254.34
R2685 GNDA.n483 GNDA.n115 254.34
R2686 GNDA.n449 GNDA.n115 254.34
R2687 GNDA.n476 GNDA.n115 254.34
R2688 GNDA.n470 GNDA.n115 254.34
R2689 GNDA.n468 GNDA.n115 254.34
R2690 GNDA.n462 GNDA.n115 254.34
R2691 GNDA.n2158 GNDA.n121 254.34
R2692 GNDA.n2158 GNDA.n120 254.34
R2693 GNDA.n2158 GNDA.n119 254.34
R2694 GNDA.n2158 GNDA.n118 254.34
R2695 GNDA.n2158 GNDA.n117 254.34
R2696 GNDA.n2158 GNDA.n116 254.34
R2697 GNDA.n227 GNDA.n126 254.34
R2698 GNDA.n1970 GNDA.n126 254.34
R2699 GNDA.n1972 GNDA.n126 254.34
R2700 GNDA.n1978 GNDA.n126 254.34
R2701 GNDA.n1980 GNDA.n126 254.34
R2702 GNDA.n1986 GNDA.n126 254.34
R2703 GNDA.n1759 GNDA.n489 254.34
R2704 GNDA.n2157 GNDA.n131 254.34
R2705 GNDA.n2157 GNDA.n132 254.34
R2706 GNDA.n2157 GNDA.n133 254.34
R2707 GNDA.n2157 GNDA.n134 254.34
R2708 GNDA.n2157 GNDA.n135 254.34
R2709 GNDA.n350 GNDA.n229 254.34
R2710 GNDA.n2157 GNDA.n137 254.34
R2711 GNDA.n2157 GNDA.n138 254.34
R2712 GNDA.n2157 GNDA.n139 254.34
R2713 GNDA.n2157 GNDA.n140 254.34
R2714 GNDA.n2157 GNDA.n141 254.34
R2715 GNDA.n2147 GNDA.n200 254.34
R2716 GNDA.n2157 GNDA.n143 254.34
R2717 GNDA.n2157 GNDA.n144 254.34
R2718 GNDA.n2157 GNDA.n145 254.34
R2719 GNDA.n2157 GNDA.n146 254.34
R2720 GNDA.n2157 GNDA.n147 254.34
R2721 GNDA.n2152 GNDA.n171 254.34
R2722 GNDA.n2152 GNDA.n170 254.34
R2723 GNDA.n2152 GNDA.n169 254.34
R2724 GNDA.n2152 GNDA.n168 254.34
R2725 GNDA.n2152 GNDA.n167 254.34
R2726 GNDA.n1761 GNDA.n447 254.34
R2727 GNDA.n2152 GNDA.n165 254.34
R2728 GNDA.n2152 GNDA.n164 254.34
R2729 GNDA.n2152 GNDA.n163 254.34
R2730 GNDA.n2152 GNDA.n162 254.34
R2731 GNDA.n2152 GNDA.n161 254.34
R2732 GNDA.n1244 GNDA.n1243 254.34
R2733 GNDA.n2153 GNDA.n2152 254.34
R2734 GNDA.n2152 GNDA.n159 254.34
R2735 GNDA.n2152 GNDA.n158 254.34
R2736 GNDA.n2152 GNDA.n157 254.34
R2737 GNDA.n2152 GNDA.n156 254.34
R2738 GNDA.n2150 GNDA.n2149 254.34
R2739 GNDA.n514 GNDA.n100 254.34
R2740 GNDA.n310 GNDA.n77 254.34
R2741 GNDA.n2120 GNDA.n2119 254.34
R2742 GNDA.n2226 GNDA.n2225 253.238
R2743 GNDA.n956 GNDA.n862 252.875
R2744 GNDA.n572 GNDA.n360 250.349
R2745 GNDA.n2156 GNDA.n148 249.663
R2746 GNDA.n484 GNDA.n142 249.663
R2747 GNDA.n1620 GNDA.n136 249.663
R2748 GNDA.n1558 GNDA.n809 249.663
R2749 GNDA.n1535 GNDA.n829 249.663
R2750 GNDA.n1213 GNDA.n416 249.663
R2751 GNDA.n1407 GNDA.n422 249.663
R2752 GNDA.n672 GNDA.n637 249.663
R2753 GNDA.n1591 GNDA.n1589 249.663
R2754 GNDA.n2430 GNDA.n2429 246.4
R2755 GNDA.n2237 GNDA.n2236 246.4
R2756 GNDA.t250 GNDA.n630 244.762
R2757 GNDA.n1545 GNDA.t250 244.762
R2758 GNDA.t250 GNDA.n1079 244.762
R2759 GNDA.n917 GNDA.n916 240
R2760 GNDA.n942 GNDA.n920 240
R2761 GNDA.t250 GNDA.n622 239.004
R2762 GNDA.n1038 GNDA.n957 239.004
R2763 GNDA.t252 GNDA.n364 239.004
R2764 GNDA.n2131 GNDA.t243 239.004
R2765 GNDA.n2371 GNDA.n2370 238.4
R2766 GNDA.n2230 GNDA.n2220 238.4
R2767 GNDA.n2282 GNDA.n34 233.601
R2768 GNDA.n2457 GNDA.n34 233.601
R2769 GNDA.n2468 GNDA.n2466 227.096
R2770 GNDA.n2465 GNDA.n2463 227.096
R2771 GNDA.n2468 GNDA.n2467 226.534
R2772 GNDA.n2465 GNDA.n2464 226.534
R2773 GNDA.n2362 GNDA.t246 224.525
R2774 GNDA.n2389 GNDA.t261 224.525
R2775 GNDA.n2202 GNDA.t314 224.525
R2776 GNDA.n2256 GNDA.t302 224.525
R2777 GNDA.n2471 GNDA.n2470 222.034
R2778 GNDA.n756 GNDA.n755 221.667
R2779 GNDA.n1817 GNDA.n1816 221.667
R2780 GNDA.n1713 GNDA.n1712 221.667
R2781 GNDA.n1171 GNDA.n1125 221.667
R2782 GNDA.n1300 GNDA.n1299 221.667
R2783 GNDA.n293 GNDA.n248 221.667
R2784 GNDA.n1012 GNDA.n968 221.667
R2785 GNDA.n1928 GNDA.n386 221.667
R2786 GNDA.n2080 GNDA.n2079 221.667
R2787 GNDA.n2116 GNDA.n2115 218.715
R2788 GNDA.n2498 GNDA.n3 217.601
R2789 GNDA.n2442 GNDA.n3 214.4
R2790 GNDA.n31 GNDA.n30 211.201
R2791 GNDA.n30 GNDA.n28 211.201
R2792 GNDA.n2356 GNDA.n2355 211.201
R2793 GNDA.n2355 GNDA.n2349 211.201
R2794 GNDA.n2211 GNDA.n2210 211.201
R2795 GNDA.n2211 GNDA.n2207 211.201
R2796 GNDA.n2503 GNDA.n2501 206.052
R2797 GNDA.n2268 GNDA.n2266 206.052
R2798 GNDA.n2511 GNDA.n2510 205.488
R2799 GNDA.n2509 GNDA.n2508 205.488
R2800 GNDA.n2507 GNDA.n2506 205.488
R2801 GNDA.n2505 GNDA.n2504 205.488
R2802 GNDA.n2503 GNDA.n2502 205.488
R2803 GNDA.n2276 GNDA.n2275 205.488
R2804 GNDA.n2274 GNDA.n2273 205.488
R2805 GNDA.n2272 GNDA.n2271 205.488
R2806 GNDA.n2270 GNDA.n2269 205.488
R2807 GNDA.n2268 GNDA.n2267 205.488
R2808 GNDA.n2442 GNDA.n2 203.201
R2809 GNDA.n2499 GNDA.n2498 201.601
R2810 GNDA.n1590 GNDA.n401 200.81
R2811 GNDA.n1619 GNDA.n127 200.81
R2812 GNDA.n2117 GNDA.n2005 197
R2813 GNDA.n313 GNDA.n312 197
R2814 GNDA.n1660 GNDA.n1659 197
R2815 GNDA.n571 GNDA.n570 197
R2816 GNDA.n1216 GNDA.n608 197
R2817 GNDA.n1032 GNDA.n607 197
R2818 GNDA.n2151 GNDA.n174 197
R2819 GNDA.n1247 GNDA.n173 197
R2820 GNDA.n1567 GNDA.n609 197
R2821 GNDA.n1764 GNDA.n172 197
R2822 GNDA.n2375 GNDA.n2370 195
R2823 GNDA.n2376 GNDA.n2375 195
R2824 GNDA.n2382 GNDA.n2381 195
R2825 GNDA.n2383 GNDA.n2382 195
R2826 GNDA.n2222 GNDA.n2221 195
R2827 GNDA.n2222 GNDA.n2191 195
R2828 GNDA.n2224 GNDA.n2220 195
R2829 GNDA.n2225 GNDA.n2224 195
R2830 GNDA.n2392 GNDA.n2391 192
R2831 GNDA.n2258 GNDA.n2257 192
R2832 GNDA.n1991 GNDA.n1988 187.249
R2833 GNDA.n461 GNDA.n460 187.249
R2834 GNDA.n1644 GNDA.n525 187.249
R2835 GNDA.n1439 GNDA.n1438 187.249
R2836 GNDA.n1496 GNDA.n1495 187.249
R2837 GNDA.n2154 GNDA.n152 187.249
R2838 GNDA.n1386 GNDA.n1385 187.249
R2839 GNDA.n648 GNDA.n580 187.249
R2840 GNDA.n1616 GNDA.n562 187.249
R2841 GNDA.n722 GNDA.n695 185
R2842 GNDA.n723 GNDA.n720 185
R2843 GNDA.n723 GNDA.t293 185
R2844 GNDA.n726 GNDA.n725 185
R2845 GNDA.n727 GNDA.n719 185
R2846 GNDA.n729 GNDA.n728 185
R2847 GNDA.n731 GNDA.n718 185
R2848 GNDA.n734 GNDA.n733 185
R2849 GNDA.n735 GNDA.n717 185
R2850 GNDA.n737 GNDA.n736 185
R2851 GNDA.n739 GNDA.n716 185
R2852 GNDA.n742 GNDA.n741 185
R2853 GNDA.n743 GNDA.n715 185
R2854 GNDA.n745 GNDA.n744 185
R2855 GNDA.n747 GNDA.n714 185
R2856 GNDA.n750 GNDA.n749 185
R2857 GNDA.n751 GNDA.n713 185
R2858 GNDA.n753 GNDA.n752 185
R2859 GNDA.n755 GNDA.n712 185
R2860 GNDA.n772 GNDA.n707 185
R2861 GNDA.n770 GNDA.n769 185
R2862 GNDA.n768 GNDA.n708 185
R2863 GNDA.n767 GNDA.n766 185
R2864 GNDA.n764 GNDA.n709 185
R2865 GNDA.n762 GNDA.n761 185
R2866 GNDA.n760 GNDA.n710 185
R2867 GNDA.n710 GNDA.t293 185
R2868 GNDA.n759 GNDA.n758 185
R2869 GNDA.n756 GNDA.n711 185
R2870 GNDA.n1783 GNDA.n1782 185
R2871 GNDA.n1784 GNDA.n1781 185
R2872 GNDA.n1784 GNDA.t292 185
R2873 GNDA.n1787 GNDA.n1786 185
R2874 GNDA.n1788 GNDA.n1780 185
R2875 GNDA.n1790 GNDA.n1789 185
R2876 GNDA.n1792 GNDA.n1779 185
R2877 GNDA.n1795 GNDA.n1794 185
R2878 GNDA.n1796 GNDA.n1778 185
R2879 GNDA.n1798 GNDA.n1797 185
R2880 GNDA.n1800 GNDA.n1777 185
R2881 GNDA.n1803 GNDA.n1802 185
R2882 GNDA.n1804 GNDA.n1776 185
R2883 GNDA.n1806 GNDA.n1805 185
R2884 GNDA.n1808 GNDA.n1775 185
R2885 GNDA.n1811 GNDA.n1810 185
R2886 GNDA.n1812 GNDA.n1774 185
R2887 GNDA.n1814 GNDA.n1813 185
R2888 GNDA.n1816 GNDA.n1773 185
R2889 GNDA.n1833 GNDA.n1768 185
R2890 GNDA.n1831 GNDA.n1830 185
R2891 GNDA.n1829 GNDA.n1769 185
R2892 GNDA.n1828 GNDA.n1827 185
R2893 GNDA.n1825 GNDA.n1770 185
R2894 GNDA.n1823 GNDA.n1822 185
R2895 GNDA.n1821 GNDA.n1771 185
R2896 GNDA.n1771 GNDA.t292 185
R2897 GNDA.n1820 GNDA.n1819 185
R2898 GNDA.n1817 GNDA.n1772 185
R2899 GNDA.n1679 GNDA.n1678 185
R2900 GNDA.n1680 GNDA.n1677 185
R2901 GNDA.n1680 GNDA.t267 185
R2902 GNDA.n1683 GNDA.n1682 185
R2903 GNDA.n1684 GNDA.n1676 185
R2904 GNDA.n1686 GNDA.n1685 185
R2905 GNDA.n1688 GNDA.n1675 185
R2906 GNDA.n1691 GNDA.n1690 185
R2907 GNDA.n1692 GNDA.n1674 185
R2908 GNDA.n1694 GNDA.n1693 185
R2909 GNDA.n1696 GNDA.n1673 185
R2910 GNDA.n1699 GNDA.n1698 185
R2911 GNDA.n1700 GNDA.n1672 185
R2912 GNDA.n1702 GNDA.n1701 185
R2913 GNDA.n1704 GNDA.n1671 185
R2914 GNDA.n1707 GNDA.n1706 185
R2915 GNDA.n1708 GNDA.n1670 185
R2916 GNDA.n1710 GNDA.n1709 185
R2917 GNDA.n1712 GNDA.n1669 185
R2918 GNDA.n1729 GNDA.n1664 185
R2919 GNDA.n1727 GNDA.n1726 185
R2920 GNDA.n1725 GNDA.n1665 185
R2921 GNDA.n1724 GNDA.n1723 185
R2922 GNDA.n1721 GNDA.n1666 185
R2923 GNDA.n1719 GNDA.n1718 185
R2924 GNDA.n1717 GNDA.n1667 185
R2925 GNDA.n1667 GNDA.t267 185
R2926 GNDA.n1716 GNDA.n1715 185
R2927 GNDA.n1713 GNDA.n1668 185
R2928 GNDA.n1136 GNDA.n1135 185
R2929 GNDA.n1137 GNDA.n1133 185
R2930 GNDA.n1133 GNDA.t249 185
R2931 GNDA.n1139 GNDA.n1138 185
R2932 GNDA.n1141 GNDA.n1132 185
R2933 GNDA.n1144 GNDA.n1143 185
R2934 GNDA.n1145 GNDA.n1131 185
R2935 GNDA.n1147 GNDA.n1146 185
R2936 GNDA.n1149 GNDA.n1130 185
R2937 GNDA.n1152 GNDA.n1151 185
R2938 GNDA.n1153 GNDA.n1129 185
R2939 GNDA.n1155 GNDA.n1154 185
R2940 GNDA.n1157 GNDA.n1128 185
R2941 GNDA.n1160 GNDA.n1159 185
R2942 GNDA.n1161 GNDA.n1127 185
R2943 GNDA.n1163 GNDA.n1162 185
R2944 GNDA.n1165 GNDA.n1126 185
R2945 GNDA.n1168 GNDA.n1167 185
R2946 GNDA.n1169 GNDA.n1125 185
R2947 GNDA.n1186 GNDA.n1119 185
R2948 GNDA.n1185 GNDA.n1184 185
R2949 GNDA.n1182 GNDA.n1121 185
R2950 GNDA.n1180 GNDA.n1179 185
R2951 GNDA.n1178 GNDA.n1122 185
R2952 GNDA.n1177 GNDA.n1176 185
R2953 GNDA.n1174 GNDA.n1123 185
R2954 GNDA.n1174 GNDA.t249 185
R2955 GNDA.n1173 GNDA.n1124 185
R2956 GNDA.n1171 GNDA.n1170 185
R2957 GNDA.n1266 GNDA.n1265 185
R2958 GNDA.n1267 GNDA.n1264 185
R2959 GNDA.n1267 GNDA.t251 185
R2960 GNDA.n1270 GNDA.n1269 185
R2961 GNDA.n1271 GNDA.n1263 185
R2962 GNDA.n1273 GNDA.n1272 185
R2963 GNDA.n1275 GNDA.n1262 185
R2964 GNDA.n1278 GNDA.n1277 185
R2965 GNDA.n1279 GNDA.n1261 185
R2966 GNDA.n1281 GNDA.n1280 185
R2967 GNDA.n1283 GNDA.n1260 185
R2968 GNDA.n1286 GNDA.n1285 185
R2969 GNDA.n1287 GNDA.n1259 185
R2970 GNDA.n1289 GNDA.n1288 185
R2971 GNDA.n1291 GNDA.n1258 185
R2972 GNDA.n1294 GNDA.n1293 185
R2973 GNDA.n1295 GNDA.n1257 185
R2974 GNDA.n1297 GNDA.n1296 185
R2975 GNDA.n1299 GNDA.n1256 185
R2976 GNDA.n1316 GNDA.n1251 185
R2977 GNDA.n1314 GNDA.n1313 185
R2978 GNDA.n1312 GNDA.n1252 185
R2979 GNDA.n1311 GNDA.n1310 185
R2980 GNDA.n1308 GNDA.n1253 185
R2981 GNDA.n1306 GNDA.n1305 185
R2982 GNDA.n1304 GNDA.n1254 185
R2983 GNDA.n1254 GNDA.t251 185
R2984 GNDA.n1303 GNDA.n1302 185
R2985 GNDA.n1300 GNDA.n1255 185
R2986 GNDA.n257 GNDA.n230 185
R2987 GNDA.n259 GNDA.n258 185
R2988 GNDA.n258 GNDA.t333 185
R2989 GNDA.n261 GNDA.n260 185
R2990 GNDA.n263 GNDA.n255 185
R2991 GNDA.n266 GNDA.n265 185
R2992 GNDA.n267 GNDA.n254 185
R2993 GNDA.n269 GNDA.n268 185
R2994 GNDA.n271 GNDA.n253 185
R2995 GNDA.n274 GNDA.n273 185
R2996 GNDA.n275 GNDA.n252 185
R2997 GNDA.n277 GNDA.n276 185
R2998 GNDA.n279 GNDA.n251 185
R2999 GNDA.n282 GNDA.n281 185
R3000 GNDA.n283 GNDA.n250 185
R3001 GNDA.n285 GNDA.n284 185
R3002 GNDA.n287 GNDA.n249 185
R3003 GNDA.n290 GNDA.n289 185
R3004 GNDA.n291 GNDA.n248 185
R3005 GNDA.n308 GNDA.n307 185
R3006 GNDA.n305 GNDA.n241 185
R3007 GNDA.n304 GNDA.n244 185
R3008 GNDA.n302 GNDA.n301 185
R3009 GNDA.n300 GNDA.n245 185
R3010 GNDA.n299 GNDA.n298 185
R3011 GNDA.n296 GNDA.n246 185
R3012 GNDA.n296 GNDA.t333 185
R3013 GNDA.n295 GNDA.n247 185
R3014 GNDA.n293 GNDA.n292 185
R3015 GNDA.n976 GNDA.n844 185
R3016 GNDA.n978 GNDA.n977 185
R3017 GNDA.n977 GNDA.t266 185
R3018 GNDA.n980 GNDA.n979 185
R3019 GNDA.n982 GNDA.n975 185
R3020 GNDA.n985 GNDA.n984 185
R3021 GNDA.n986 GNDA.n974 185
R3022 GNDA.n988 GNDA.n987 185
R3023 GNDA.n990 GNDA.n973 185
R3024 GNDA.n993 GNDA.n992 185
R3025 GNDA.n994 GNDA.n972 185
R3026 GNDA.n996 GNDA.n995 185
R3027 GNDA.n998 GNDA.n971 185
R3028 GNDA.n1001 GNDA.n1000 185
R3029 GNDA.n1002 GNDA.n970 185
R3030 GNDA.n1004 GNDA.n1003 185
R3031 GNDA.n1006 GNDA.n969 185
R3032 GNDA.n1009 GNDA.n1008 185
R3033 GNDA.n1010 GNDA.n968 185
R3034 GNDA.n1027 GNDA.n1026 185
R3035 GNDA.n1024 GNDA.n961 185
R3036 GNDA.n1023 GNDA.n964 185
R3037 GNDA.n1021 GNDA.n1020 185
R3038 GNDA.n1019 GNDA.n965 185
R3039 GNDA.n1018 GNDA.n1017 185
R3040 GNDA.n1015 GNDA.n966 185
R3041 GNDA.n1015 GNDA.t266 185
R3042 GNDA.n1014 GNDA.n967 185
R3043 GNDA.n1012 GNDA.n1011 185
R3044 GNDA.n1893 GNDA.n1892 185
R3045 GNDA.n1894 GNDA.n394 185
R3046 GNDA.n394 GNDA.t265 185
R3047 GNDA.n1896 GNDA.n1895 185
R3048 GNDA.n1898 GNDA.n393 185
R3049 GNDA.n1901 GNDA.n1900 185
R3050 GNDA.n1902 GNDA.n392 185
R3051 GNDA.n1904 GNDA.n1903 185
R3052 GNDA.n1906 GNDA.n391 185
R3053 GNDA.n1909 GNDA.n1908 185
R3054 GNDA.n1910 GNDA.n390 185
R3055 GNDA.n1912 GNDA.n1911 185
R3056 GNDA.n1914 GNDA.n389 185
R3057 GNDA.n1917 GNDA.n1916 185
R3058 GNDA.n1918 GNDA.n388 185
R3059 GNDA.n1920 GNDA.n1919 185
R3060 GNDA.n1922 GNDA.n387 185
R3061 GNDA.n1925 GNDA.n1924 185
R3062 GNDA.n1926 GNDA.n386 185
R3063 GNDA.n1943 GNDA.n1942 185
R3064 GNDA.n1940 GNDA.n379 185
R3065 GNDA.n1939 GNDA.n382 185
R3066 GNDA.n1937 GNDA.n1936 185
R3067 GNDA.n1935 GNDA.n383 185
R3068 GNDA.n1934 GNDA.n1933 185
R3069 GNDA.n1931 GNDA.n384 185
R3070 GNDA.n1931 GNDA.t265 185
R3071 GNDA.n1930 GNDA.n385 185
R3072 GNDA.n1928 GNDA.n1927 185
R3073 GNDA.n2046 GNDA.n2044 185
R3074 GNDA.n2047 GNDA.n2043 185
R3075 GNDA.n2047 GNDA.t242 185
R3076 GNDA.n2050 GNDA.n2049 185
R3077 GNDA.n2051 GNDA.n2042 185
R3078 GNDA.n2053 GNDA.n2052 185
R3079 GNDA.n2055 GNDA.n2041 185
R3080 GNDA.n2058 GNDA.n2057 185
R3081 GNDA.n2059 GNDA.n2040 185
R3082 GNDA.n2061 GNDA.n2060 185
R3083 GNDA.n2063 GNDA.n2039 185
R3084 GNDA.n2066 GNDA.n2065 185
R3085 GNDA.n2067 GNDA.n2038 185
R3086 GNDA.n2069 GNDA.n2068 185
R3087 GNDA.n2071 GNDA.n2037 185
R3088 GNDA.n2074 GNDA.n2073 185
R3089 GNDA.n2075 GNDA.n2036 185
R3090 GNDA.n2077 GNDA.n2076 185
R3091 GNDA.n2079 GNDA.n2035 185
R3092 GNDA.n2096 GNDA.n2030 185
R3093 GNDA.n2094 GNDA.n2093 185
R3094 GNDA.n2092 GNDA.n2031 185
R3095 GNDA.n2091 GNDA.n2090 185
R3096 GNDA.n2088 GNDA.n2032 185
R3097 GNDA.n2086 GNDA.n2085 185
R3098 GNDA.n2084 GNDA.n2033 185
R3099 GNDA.n2033 GNDA.t242 185
R3100 GNDA.n2083 GNDA.n2082 185
R3101 GNDA.n2080 GNDA.n2034 185
R3102 GNDA.n2098 GNDA.n2097 185
R3103 GNDA.n2027 GNDA.n2010 185
R3104 GNDA.n2026 GNDA.n2025 185
R3105 GNDA.n2016 GNDA.n2013 185
R3106 GNDA.n2018 GNDA.n2017 185
R3107 GNDA.n210 GNDA.n209 185
R3108 GNDA.n2136 GNDA.n2135 185
R3109 GNDA.n2139 GNDA.n2138 185
R3110 GNDA.n208 GNDA.n206 185
R3111 GNDA.n381 GNDA.n378 185
R3112 GNDA.n372 GNDA.n371 185
R3113 GNDA.n1954 GNDA.n1953 185
R3114 GNDA.n1957 GNDA.n1956 185
R3115 GNDA.n370 GNDA.n368 185
R3116 GNDA.n1881 GNDA.n1880 185
R3117 GNDA.n1878 GNDA.n1875 185
R3118 GNDA.n398 GNDA.n396 185
R3119 GNDA.n1890 GNDA.n1889 185
R3120 GNDA.n963 GNDA.n960 185
R3121 GNDA.n858 GNDA.n856 185
R3122 GNDA.n1044 GNDA.n1043 185
R3123 GNDA.n1046 GNDA.n855 185
R3124 GNDA.n1048 GNDA.n1047 185
R3125 GNDA.n850 GNDA.n848 185
R3126 GNDA.n1059 GNDA.n1058 185
R3127 GNDA.n1061 GNDA.n847 185
R3128 GNDA.n1063 GNDA.n1062 185
R3129 GNDA.n243 GNDA.n240 185
R3130 GNDA.n321 GNDA.n239 185
R3131 GNDA.n326 GNDA.n325 185
R3132 GNDA.n329 GNDA.n328 185
R3133 GNDA.n238 GNDA.n235 185
R3134 GNDA.n334 GNDA.n234 185
R3135 GNDA.n339 GNDA.n338 185
R3136 GNDA.n342 GNDA.n341 185
R3137 GNDA.n233 GNDA.n231 185
R3138 GNDA.n1318 GNDA.n1317 185
R3139 GNDA.n1237 GNDA.n1235 185
R3140 GNDA.n1325 GNDA.n1324 185
R3141 GNDA.n1327 GNDA.n1234 185
R3142 GNDA.n1329 GNDA.n1328 185
R3143 GNDA.n1228 GNDA.n1226 185
R3144 GNDA.n1336 GNDA.n1335 185
R3145 GNDA.n1338 GNDA.n1225 185
R3146 GNDA.n1340 GNDA.n1339 185
R3147 GNDA.n1506 GNDA.n1505 185
R3148 GNDA.n1508 GNDA.n1118 185
R3149 GNDA.n1510 GNDA.n1509 185
R3150 GNDA.n1116 GNDA.n1109 185
R3151 GNDA.n1115 GNDA.n1114 185
R3152 GNDA.n1101 GNDA.n1100 185
R3153 GNDA.n1524 GNDA.n1523 185
R3154 GNDA.n1527 GNDA.n1526 185
R3155 GNDA.n1099 GNDA.n1097 185
R3156 GNDA.n1731 GNDA.n1730 185
R3157 GNDA.n506 GNDA.n504 185
R3158 GNDA.n1738 GNDA.n1737 185
R3159 GNDA.n1740 GNDA.n503 185
R3160 GNDA.n1742 GNDA.n1741 185
R3161 GNDA.n497 GNDA.n495 185
R3162 GNDA.n1749 GNDA.n1748 185
R3163 GNDA.n1751 GNDA.n494 185
R3164 GNDA.n1753 GNDA.n1752 185
R3165 GNDA.n1835 GNDA.n1834 185
R3166 GNDA.n441 GNDA.n439 185
R3167 GNDA.n1842 GNDA.n1841 185
R3168 GNDA.n1844 GNDA.n438 185
R3169 GNDA.n1846 GNDA.n1845 185
R3170 GNDA.n432 GNDA.n430 185
R3171 GNDA.n1853 GNDA.n1852 185
R3172 GNDA.n1855 GNDA.n429 185
R3173 GNDA.n1857 GNDA.n1856 185
R3174 GNDA.n774 GNDA.n773 185
R3175 GNDA.n777 GNDA.n704 185
R3176 GNDA.n782 GNDA.n781 185
R3177 GNDA.n785 GNDA.n784 185
R3178 GNDA.n703 GNDA.n700 185
R3179 GNDA.n790 GNDA.n699 185
R3180 GNDA.n795 GNDA.n794 185
R3181 GNDA.n798 GNDA.n797 185
R3182 GNDA.n698 GNDA.n696 185
R3183 GNDA.n2357 GNDA.n2356 182.4
R3184 GNDA.n2253 GNDA.n2207 182.4
R3185 GNDA.n2328 GNDA.n59 179.917
R3186 GNDA.n2438 GNDA.n2437 179.363
R3187 GNDA.n947 GNDA.n879 176
R3188 GNDA.n947 GNDA.n946 176
R3189 GNDA.n2428 GNDA.n2349 176
R3190 GNDA.n2210 GNDA.n2204 176
R3191 GNDA.n2145 GNDA.n202 175.546
R3192 GNDA.n2141 GNDA.n202 175.546
R3193 GNDA.n2141 GNDA.n204 175.546
R3194 GNDA.n2133 GNDA.n204 175.546
R3195 GNDA.n2133 GNDA.n211 175.546
R3196 GNDA.n2020 GNDA.n211 175.546
R3197 GNDA.n2022 GNDA.n2020 175.546
R3198 GNDA.n2022 GNDA.n2009 175.546
R3199 GNDA.n2100 GNDA.n2009 175.546
R3200 GNDA.n2100 GNDA.n2007 175.546
R3201 GNDA.n2105 GNDA.n2007 175.546
R3202 GNDA.n2156 GNDA.n149 175.546
R3203 GNDA.n179 GNDA.n178 175.546
R3204 GNDA.n185 GNDA.n184 175.546
R3205 GNDA.n191 GNDA.n190 175.546
R3206 GNDA.n197 GNDA.n196 175.546
R3207 GNDA.n1991 GNDA.n220 175.546
R3208 GNDA.n1995 GNDA.n220 175.546
R3209 GNDA.n1995 GNDA.n218 175.546
R3210 GNDA.n1999 GNDA.n218 175.546
R3211 GNDA.n1999 GNDA.n215 175.546
R3212 GNDA.n2129 GNDA.n215 175.546
R3213 GNDA.n2129 GNDA.n216 175.546
R3214 GNDA.n2125 GNDA.n216 175.546
R3215 GNDA.n2125 GNDA.n2003 175.546
R3216 GNDA.n2121 GNDA.n2003 175.546
R3217 GNDA.n1969 GNDA.n228 175.546
R3218 GNDA.n1973 GNDA.n1971 175.546
R3219 GNDA.n1977 GNDA.n225 175.546
R3220 GNDA.n1981 GNDA.n1979 175.546
R3221 GNDA.n1985 GNDA.n223 175.546
R3222 GNDA.n345 GNDA.n344 175.546
R3223 GNDA.n336 GNDA.n335 175.546
R3224 GNDA.n332 GNDA.n331 175.546
R3225 GNDA.n323 GNDA.n322 175.546
R3226 GNDA.n319 GNDA.n318 175.546
R3227 GNDA.n1357 GNDA.n142 175.546
R3228 GNDA.n1359 GNDA.n1358 175.546
R3229 GNDA.n1361 GNDA.n1360 175.546
R3230 GNDA.n1363 GNDA.n1362 175.546
R3231 GNDA.n1365 GNDA.n1364 175.546
R3232 GNDA.n460 GNDA.n455 175.546
R3233 GNDA.n455 GNDA.n111 175.546
R3234 GNDA.n2164 GNDA.n111 175.546
R3235 GNDA.n2164 GNDA.n112 175.546
R3236 GNDA.n2160 GNDA.n112 175.546
R3237 GNDA.n2160 GNDA.n75 175.546
R3238 GNDA.n2310 GNDA.n75 175.546
R3239 GNDA.n2310 GNDA.n76 175.546
R3240 GNDA.n2306 GNDA.n76 175.546
R3241 GNDA.n2306 GNDA.n78 175.546
R3242 GNDA.n482 GNDA.n481 175.546
R3243 GNDA.n478 GNDA.n477 175.546
R3244 GNDA.n475 GNDA.n451 175.546
R3245 GNDA.n471 GNDA.n469 175.546
R3246 GNDA.n467 GNDA.n453 175.546
R3247 GNDA.n1755 GNDA.n491 175.546
R3248 GNDA.n1746 GNDA.n499 175.546
R3249 GNDA.n1744 GNDA.n500 175.546
R3250 GNDA.n1735 GNDA.n508 175.546
R3251 GNDA.n1733 GNDA.n509 175.546
R3252 GNDA.n535 GNDA.n136 175.546
R3253 GNDA.n537 GNDA.n536 175.546
R3254 GNDA.n539 GNDA.n538 175.546
R3255 GNDA.n541 GNDA.n540 175.546
R3256 GNDA.n543 GNDA.n542 175.546
R3257 GNDA.n525 GNDA.n522 175.546
R3258 GNDA.n522 GNDA.n90 175.546
R3259 GNDA.n2188 GNDA.n90 175.546
R3260 GNDA.n2188 GNDA.n91 175.546
R3261 GNDA.n2184 GNDA.n91 175.546
R3262 GNDA.n2184 GNDA.n94 175.546
R3263 GNDA.n2180 GNDA.n94 175.546
R3264 GNDA.n2180 GNDA.n99 175.546
R3265 GNDA.n2176 GNDA.n99 175.546
R3266 GNDA.n2176 GNDA.n101 175.546
R3267 GNDA.n1620 GNDA.n533 175.546
R3268 GNDA.n1625 GNDA.n533 175.546
R3269 GNDA.n1625 GNDA.n531 175.546
R3270 GNDA.n1629 GNDA.n531 175.546
R3271 GNDA.n1630 GNDA.n1629 175.546
R3272 GNDA.n1630 GNDA.n529 175.546
R3273 GNDA.n1634 GNDA.n529 175.546
R3274 GNDA.n1634 GNDA.n528 175.546
R3275 GNDA.n1639 GNDA.n528 175.546
R3276 GNDA.n1639 GNDA.n526 175.546
R3277 GNDA.n1643 GNDA.n526 175.546
R3278 GNDA.n1419 GNDA.n1416 175.546
R3279 GNDA.n1423 GNDA.n1421 175.546
R3280 GNDA.n1427 GNDA.n1413 175.546
R3281 GNDA.n1431 GNDA.n1429 175.546
R3282 GNDA.n1435 GNDA.n1411 175.546
R3283 GNDA.n1558 GNDA.n810 175.546
R3284 GNDA.n1554 GNDA.n810 175.546
R3285 GNDA.n1554 GNDA.n813 175.546
R3286 GNDA.n1550 GNDA.n813 175.546
R3287 GNDA.n1550 GNDA.n815 175.546
R3288 GNDA.n1546 GNDA.n815 175.546
R3289 GNDA.n1546 GNDA.n817 175.546
R3290 GNDA.n1542 GNDA.n817 175.546
R3291 GNDA.n1542 GNDA.n819 175.546
R3292 GNDA.n824 GNDA.n819 175.546
R3293 GNDA.n1444 GNDA.n1443 175.546
R3294 GNDA.n1450 GNDA.n1449 175.546
R3295 GNDA.n1456 GNDA.n1455 175.546
R3296 GNDA.n1460 GNDA.n595 175.546
R3297 GNDA.n1465 GNDA.n595 175.546
R3298 GNDA.n1537 GNDA.n823 175.546
R3299 GNDA.n1529 GNDA.n823 175.546
R3300 GNDA.n1529 GNDA.n1095 175.546
R3301 GNDA.n1521 GNDA.n1095 175.546
R3302 GNDA.n1521 GNDA.n1102 175.546
R3303 GNDA.n1107 GNDA.n1102 175.546
R3304 GNDA.n1512 GNDA.n1107 175.546
R3305 GNDA.n1512 GNDA.n1108 175.546
R3306 GNDA.n1188 GNDA.n1108 175.546
R3307 GNDA.n1503 GNDA.n1188 175.546
R3308 GNDA.n1503 GNDA.n1189 175.546
R3309 GNDA.n1067 GNDA.n843 175.546
R3310 GNDA.n1052 GNDA.n843 175.546
R3311 GNDA.n1052 GNDA.n851 175.546
R3312 GNDA.n1056 GNDA.n851 175.546
R3313 GNDA.n1056 GNDA.n1050 175.546
R3314 GNDA.n1050 GNDA.n852 175.546
R3315 GNDA.n859 GNDA.n852 175.546
R3316 GNDA.n1041 GNDA.n859 175.546
R3317 GNDA.n1041 GNDA.n860 175.546
R3318 GNDA.n1037 GNDA.n860 175.546
R3319 GNDA.n1037 GNDA.n958 175.546
R3320 GNDA.n1089 GNDA.n829 175.546
R3321 GNDA.n1089 GNDA.n832 175.546
R3322 GNDA.n1085 GNDA.n832 175.546
R3323 GNDA.n1085 GNDA.n835 175.546
R3324 GNDA.n1081 GNDA.n835 175.546
R3325 GNDA.n1081 GNDA.n837 175.546
R3326 GNDA.n1077 GNDA.n837 175.546
R3327 GNDA.n1077 GNDA.n839 175.546
R3328 GNDA.n1073 GNDA.n839 175.546
R3329 GNDA.n1073 GNDA.n841 175.546
R3330 GNDA.n1492 GNDA.n1491 175.546
R3331 GNDA.n1488 GNDA.n1487 175.546
R3332 GNDA.n1484 GNDA.n1483 175.546
R3333 GNDA.n1480 GNDA.n1479 175.546
R3334 GNDA.n1476 GNDA.n601 175.546
R3335 GNDA.n1535 GNDA.n830 175.546
R3336 GNDA.n1531 GNDA.n830 175.546
R3337 GNDA.n1531 GNDA.n1093 175.546
R3338 GNDA.n1519 GNDA.n1093 175.546
R3339 GNDA.n1519 GNDA.n1103 175.546
R3340 GNDA.n1515 GNDA.n1103 175.546
R3341 GNDA.n1515 GNDA.n1514 175.546
R3342 GNDA.n1514 GNDA.n1105 175.546
R3343 GNDA.n1191 GNDA.n1105 175.546
R3344 GNDA.n1501 GNDA.n1191 175.546
R3345 GNDA.n1501 GNDA.n1192 175.546
R3346 GNDA.n1871 GNDA.n399 175.546
R3347 GNDA.n1887 GNDA.n399 175.546
R3348 GNDA.n1887 GNDA.n400 175.546
R3349 GNDA.n1883 GNDA.n400 175.546
R3350 GNDA.n1883 GNDA.n366 175.546
R3351 GNDA.n1959 GNDA.n366 175.546
R3352 GNDA.n1959 GNDA.n367 175.546
R3353 GNDA.n1951 GNDA.n367 175.546
R3354 GNDA.n1951 GNDA.n373 175.546
R3355 GNDA.n1947 GNDA.n373 175.546
R3356 GNDA.n1947 GNDA.n376 175.546
R3357 GNDA.n1468 GNDA.n416 175.546
R3358 GNDA.n1470 GNDA.n1469 175.546
R3359 GNDA.n1472 GNDA.n1471 175.546
R3360 GNDA.n1474 GNDA.n1473 175.546
R3361 GNDA.n1475 GNDA.n404 175.546
R3362 GNDA.n176 GNDA.n153 175.546
R3363 GNDA.n182 GNDA.n181 175.546
R3364 GNDA.n188 GNDA.n187 175.546
R3365 GNDA.n194 GNDA.n193 175.546
R3366 GNDA.n198 GNDA.n155 175.546
R3367 GNDA.n1211 GNDA.n1210 175.546
R3368 GNDA.n1207 GNDA.n1206 175.546
R3369 GNDA.n1203 GNDA.n1202 175.546
R3370 GNDA.n1199 GNDA.n1198 175.546
R3371 GNDA.n1195 GNDA.n353 175.546
R3372 GNDA.n1342 GNDA.n1222 175.546
R3373 GNDA.n1333 GNDA.n1230 175.546
R3374 GNDA.n1331 GNDA.n1231 175.546
R3375 GNDA.n1322 GNDA.n1239 175.546
R3376 GNDA.n1320 GNDA.n1240 175.546
R3377 GNDA.n1441 GNDA.n422 175.546
R3378 GNDA.n1447 GNDA.n1446 175.546
R3379 GNDA.n1453 GNDA.n1452 175.546
R3380 GNDA.n1459 GNDA.n1458 175.546
R3381 GNDA.n1464 GNDA.n1463 175.546
R3382 GNDA.n1382 GNDA.n1381 175.546
R3383 GNDA.n1378 GNDA.n1377 175.546
R3384 GNDA.n1374 GNDA.n1373 175.546
R3385 GNDA.n1370 GNDA.n1369 175.546
R3386 GNDA.n1366 GNDA.n160 175.546
R3387 GNDA.n1405 GNDA.n1404 175.546
R3388 GNDA.n1402 GNDA.n1350 175.546
R3389 GNDA.n1398 GNDA.n1397 175.546
R3390 GNDA.n1395 GNDA.n1353 175.546
R3391 GNDA.n1391 GNDA.n1390 175.546
R3392 GNDA.n801 GNDA.n800 175.546
R3393 GNDA.n792 GNDA.n791 175.546
R3394 GNDA.n788 GNDA.n787 175.546
R3395 GNDA.n779 GNDA.n778 175.546
R3396 GNDA.n775 GNDA.n611 175.546
R3397 GNDA.n582 GNDA.n581 175.546
R3398 GNDA.n584 GNDA.n583 175.546
R3399 GNDA.n586 GNDA.n585 175.546
R3400 GNDA.n588 GNDA.n587 175.546
R3401 GNDA.n1570 GNDA.n589 175.546
R3402 GNDA.n672 GNDA.n639 175.546
R3403 GNDA.n668 GNDA.n639 175.546
R3404 GNDA.n668 GNDA.n641 175.546
R3405 GNDA.n664 GNDA.n641 175.546
R3406 GNDA.n664 GNDA.n642 175.546
R3407 GNDA.n660 GNDA.n642 175.546
R3408 GNDA.n660 GNDA.n659 175.546
R3409 GNDA.n659 GNDA.n644 175.546
R3410 GNDA.n655 GNDA.n644 175.546
R3411 GNDA.n655 GNDA.n646 175.546
R3412 GNDA.n651 GNDA.n646 175.546
R3413 GNDA.n676 GNDA.n637 175.546
R3414 GNDA.n676 GNDA.n635 175.546
R3415 GNDA.n680 GNDA.n635 175.546
R3416 GNDA.n680 GNDA.n633 175.546
R3417 GNDA.n684 GNDA.n633 175.546
R3418 GNDA.n684 GNDA.n631 175.546
R3419 GNDA.n688 GNDA.n631 175.546
R3420 GNDA.n688 GNDA.n628 175.546
R3421 GNDA.n692 GNDA.n628 175.546
R3422 GNDA.n692 GNDA.n629 175.546
R3423 GNDA.n1859 GNDA.n426 175.546
R3424 GNDA.n1850 GNDA.n434 175.546
R3425 GNDA.n1848 GNDA.n435 175.546
R3426 GNDA.n1839 GNDA.n443 175.546
R3427 GNDA.n1837 GNDA.n444 175.546
R3428 GNDA.n1586 GNDA.n1585 175.546
R3429 GNDA.n1582 GNDA.n1581 175.546
R3430 GNDA.n1578 GNDA.n1577 175.546
R3431 GNDA.n1574 GNDA.n1573 175.546
R3432 GNDA.n1865 GNDA.n423 175.546
R3433 GNDA.n1591 GNDA.n577 175.546
R3434 GNDA.n1595 GNDA.n577 175.546
R3435 GNDA.n1595 GNDA.n575 175.546
R3436 GNDA.n1599 GNDA.n575 175.546
R3437 GNDA.n1599 GNDA.n567 175.546
R3438 GNDA.n1604 GNDA.n567 175.546
R3439 GNDA.n1604 GNDA.n566 175.546
R3440 GNDA.n1608 GNDA.n566 175.546
R3441 GNDA.n1608 GNDA.n564 175.546
R3442 GNDA.n1612 GNDA.n564 175.546
R3443 GNDA.n1612 GNDA.n561 175.546
R3444 GNDA.n558 GNDA.n557 175.546
R3445 GNDA.n554 GNDA.n553 175.546
R3446 GNDA.n550 GNDA.n549 175.546
R3447 GNDA.n546 GNDA.n545 175.546
R3448 GNDA.n487 GNDA.n166 175.546
R3449 GNDA.n2298 GNDA.n84 173.898
R3450 GNDA.n1560 GNDA.t250 172.876
R3451 GNDA.t250 GNDA.n624 172.615
R3452 GNDA.n2437 GNDA.n44 171.817
R3453 GNDA.n2439 GNDA.n2438 164.906
R3454 GNDA.n939 GNDA.n938 164.369
R3455 GNDA.n2330 GNDA.n56 164.369
R3456 GNDA.n773 GNDA.n772 163.333
R3457 GNDA.n1834 GNDA.n1833 163.333
R3458 GNDA.n1730 GNDA.n1729 163.333
R3459 GNDA.n1506 GNDA.n1119 163.333
R3460 GNDA.n1317 GNDA.n1316 163.333
R3461 GNDA.n307 GNDA.n243 163.333
R3462 GNDA.n1026 GNDA.n963 163.333
R3463 GNDA.n1942 GNDA.n381 163.333
R3464 GNDA.n2097 GNDA.n2096 163.333
R3465 GNDA.n2298 GNDA.n2297 161.347
R3466 GNDA.n884 GNDA.t296 160.725
R3467 GNDA.n881 GNDA.t291 160.725
R3468 GNDA.n880 GNDA.t288 160.725
R3469 GNDA.n878 GNDA.t270 160.725
R3470 GNDA.n918 GNDA.t305 160.725
R3471 GNDA.n928 GNDA.t326 160.725
R3472 GNDA.n2493 GNDA.n9 160
R3473 GNDA.n17 GNDA.n16 160
R3474 GNDA.n2481 GNDA.n2480 160
R3475 GNDA.n2317 GNDA.t30 157.555
R3476 GNDA.n2318 GNDA.t98 157.555
R3477 GNDA.n2282 GNDA.n2281 156.8
R3478 GNDA.t124 GNDA.n2226 156.691
R3479 GNDA.n2451 GNDA.n39 153.601
R3480 GNDA.n2390 GNDA.n2363 153.601
R3481 GNDA.n2255 GNDA.n2203 153.601
R3482 GNDA.n2486 GNDA.n2485 153.601
R3483 GNDA.n64 GNDA.t100 153.294
R3484 GNDA.n2348 GNDA.t273 152.994
R3485 GNDA.n2354 GNDA.t258 152.994
R3486 GNDA.n2206 GNDA.t281 152.994
R3487 GNDA.n2209 GNDA.t276 152.994
R3488 GNDA.n200 GNDA.n143 152.643
R3489 GNDA.n229 GNDA.n137 152.643
R3490 GNDA.n489 GNDA.n131 152.643
R3491 GNDA.n1218 GNDA.n600 152.643
R3492 GNDA.n1868 GNDA.n1867 152.643
R3493 GNDA.n1220 GNDA.n417 152.643
R3494 GNDA.n2457 GNDA.n2456 150.4
R3495 GNDA.n2445 GNDA.n40 150.4
R3496 GNDA.n797 GNDA.n698 150
R3497 GNDA.n795 GNDA.n699 150
R3498 GNDA.n784 GNDA.n703 150
R3499 GNDA.n782 GNDA.n704 150
R3500 GNDA.n758 GNDA.n710 150
R3501 GNDA.n762 GNDA.n710 150
R3502 GNDA.n766 GNDA.n764 150
R3503 GNDA.n770 GNDA.n708 150
R3504 GNDA.n741 GNDA.n739 150
R3505 GNDA.n745 GNDA.n715 150
R3506 GNDA.n749 GNDA.n747 150
R3507 GNDA.n753 GNDA.n713 150
R3508 GNDA.n737 GNDA.n717 150
R3509 GNDA.n733 GNDA.n731 150
R3510 GNDA.n729 GNDA.n719 150
R3511 GNDA.n725 GNDA.n723 150
R3512 GNDA.n723 GNDA.n722 150
R3513 GNDA.n1856 GNDA.n1855 150
R3514 GNDA.n1853 GNDA.n430 150
R3515 GNDA.n1845 GNDA.n1844 150
R3516 GNDA.n1842 GNDA.n439 150
R3517 GNDA.n1819 GNDA.n1771 150
R3518 GNDA.n1823 GNDA.n1771 150
R3519 GNDA.n1827 GNDA.n1825 150
R3520 GNDA.n1831 GNDA.n1769 150
R3521 GNDA.n1802 GNDA.n1800 150
R3522 GNDA.n1806 GNDA.n1776 150
R3523 GNDA.n1810 GNDA.n1808 150
R3524 GNDA.n1814 GNDA.n1774 150
R3525 GNDA.n1798 GNDA.n1778 150
R3526 GNDA.n1794 GNDA.n1792 150
R3527 GNDA.n1790 GNDA.n1780 150
R3528 GNDA.n1786 GNDA.n1784 150
R3529 GNDA.n1784 GNDA.n1783 150
R3530 GNDA.n1752 GNDA.n1751 150
R3531 GNDA.n1749 GNDA.n495 150
R3532 GNDA.n1741 GNDA.n1740 150
R3533 GNDA.n1738 GNDA.n504 150
R3534 GNDA.n1715 GNDA.n1667 150
R3535 GNDA.n1719 GNDA.n1667 150
R3536 GNDA.n1723 GNDA.n1721 150
R3537 GNDA.n1727 GNDA.n1665 150
R3538 GNDA.n1698 GNDA.n1696 150
R3539 GNDA.n1702 GNDA.n1672 150
R3540 GNDA.n1706 GNDA.n1704 150
R3541 GNDA.n1710 GNDA.n1670 150
R3542 GNDA.n1694 GNDA.n1674 150
R3543 GNDA.n1690 GNDA.n1688 150
R3544 GNDA.n1686 GNDA.n1676 150
R3545 GNDA.n1682 GNDA.n1680 150
R3546 GNDA.n1680 GNDA.n1679 150
R3547 GNDA.n1526 GNDA.n1099 150
R3548 GNDA.n1524 GNDA.n1100 150
R3549 GNDA.n1116 GNDA.n1115 150
R3550 GNDA.n1509 GNDA.n1508 150
R3551 GNDA.n1174 GNDA.n1173 150
R3552 GNDA.n1176 GNDA.n1174 150
R3553 GNDA.n1180 GNDA.n1122 150
R3554 GNDA.n1184 GNDA.n1182 150
R3555 GNDA.n1155 GNDA.n1129 150
R3556 GNDA.n1159 GNDA.n1157 150
R3557 GNDA.n1163 GNDA.n1127 150
R3558 GNDA.n1167 GNDA.n1165 150
R3559 GNDA.n1151 GNDA.n1149 150
R3560 GNDA.n1147 GNDA.n1131 150
R3561 GNDA.n1143 GNDA.n1141 150
R3562 GNDA.n1139 GNDA.n1133 150
R3563 GNDA.n1135 GNDA.n1133 150
R3564 GNDA.n1339 GNDA.n1338 150
R3565 GNDA.n1336 GNDA.n1226 150
R3566 GNDA.n1328 GNDA.n1327 150
R3567 GNDA.n1325 GNDA.n1235 150
R3568 GNDA.n1302 GNDA.n1254 150
R3569 GNDA.n1306 GNDA.n1254 150
R3570 GNDA.n1310 GNDA.n1308 150
R3571 GNDA.n1314 GNDA.n1252 150
R3572 GNDA.n1285 GNDA.n1283 150
R3573 GNDA.n1289 GNDA.n1259 150
R3574 GNDA.n1293 GNDA.n1291 150
R3575 GNDA.n1297 GNDA.n1257 150
R3576 GNDA.n1281 GNDA.n1261 150
R3577 GNDA.n1277 GNDA.n1275 150
R3578 GNDA.n1273 GNDA.n1263 150
R3579 GNDA.n1269 GNDA.n1267 150
R3580 GNDA.n1267 GNDA.n1266 150
R3581 GNDA.n341 GNDA.n233 150
R3582 GNDA.n339 GNDA.n234 150
R3583 GNDA.n328 GNDA.n238 150
R3584 GNDA.n326 GNDA.n239 150
R3585 GNDA.n296 GNDA.n295 150
R3586 GNDA.n298 GNDA.n296 150
R3587 GNDA.n302 GNDA.n245 150
R3588 GNDA.n305 GNDA.n304 150
R3589 GNDA.n277 GNDA.n252 150
R3590 GNDA.n281 GNDA.n279 150
R3591 GNDA.n285 GNDA.n250 150
R3592 GNDA.n289 GNDA.n287 150
R3593 GNDA.n273 GNDA.n271 150
R3594 GNDA.n269 GNDA.n254 150
R3595 GNDA.n265 GNDA.n263 150
R3596 GNDA.n261 GNDA.n258 150
R3597 GNDA.n258 GNDA.n257 150
R3598 GNDA.n1062 GNDA.n1061 150
R3599 GNDA.n1059 GNDA.n848 150
R3600 GNDA.n1047 GNDA.n1046 150
R3601 GNDA.n1044 GNDA.n856 150
R3602 GNDA.n1015 GNDA.n1014 150
R3603 GNDA.n1017 GNDA.n1015 150
R3604 GNDA.n1021 GNDA.n965 150
R3605 GNDA.n1024 GNDA.n1023 150
R3606 GNDA.n996 GNDA.n972 150
R3607 GNDA.n1000 GNDA.n998 150
R3608 GNDA.n1004 GNDA.n970 150
R3609 GNDA.n1008 GNDA.n1006 150
R3610 GNDA.n992 GNDA.n990 150
R3611 GNDA.n988 GNDA.n974 150
R3612 GNDA.n984 GNDA.n982 150
R3613 GNDA.n980 GNDA.n977 150
R3614 GNDA.n977 GNDA.n976 150
R3615 GNDA.n1890 GNDA.n396 150
R3616 GNDA.n1880 GNDA.n1878 150
R3617 GNDA.n1956 GNDA.n370 150
R3618 GNDA.n1954 GNDA.n371 150
R3619 GNDA.n1931 GNDA.n1930 150
R3620 GNDA.n1933 GNDA.n1931 150
R3621 GNDA.n1937 GNDA.n383 150
R3622 GNDA.n1940 GNDA.n1939 150
R3623 GNDA.n1912 GNDA.n390 150
R3624 GNDA.n1916 GNDA.n1914 150
R3625 GNDA.n1920 GNDA.n388 150
R3626 GNDA.n1924 GNDA.n1922 150
R3627 GNDA.n1908 GNDA.n1906 150
R3628 GNDA.n1904 GNDA.n392 150
R3629 GNDA.n1900 GNDA.n1898 150
R3630 GNDA.n1896 GNDA.n394 150
R3631 GNDA.n1892 GNDA.n394 150
R3632 GNDA.n2138 GNDA.n208 150
R3633 GNDA.n2136 GNDA.n209 150
R3634 GNDA.n2017 GNDA.n2016 150
R3635 GNDA.n2027 GNDA.n2026 150
R3636 GNDA.n2082 GNDA.n2033 150
R3637 GNDA.n2086 GNDA.n2033 150
R3638 GNDA.n2090 GNDA.n2088 150
R3639 GNDA.n2094 GNDA.n2031 150
R3640 GNDA.n2065 GNDA.n2063 150
R3641 GNDA.n2069 GNDA.n2038 150
R3642 GNDA.n2073 GNDA.n2071 150
R3643 GNDA.n2077 GNDA.n2036 150
R3644 GNDA.n2061 GNDA.n2040 150
R3645 GNDA.n2057 GNDA.n2055 150
R3646 GNDA.n2053 GNDA.n2042 150
R3647 GNDA.n2049 GNDA.n2047 150
R3648 GNDA.n2047 GNDA.n2046 150
R3649 GNDA.n2319 GNDA.t71 148.906
R3650 GNDA.n2104 GNDA.n84 148.887
R3651 GNDA.n2319 GNDA.t119 148.653
R3652 GNDA.t304 GNDA.t79 145.403
R3653 GNDA.t290 GNDA.t216 145.403
R3654 GNDA.n1647 GNDA.n1645 141.627
R3655 GNDA.n888 GNDA.n886 139.638
R3656 GNDA.t269 GNDA.t117 139.081
R3657 GNDA.t117 GNDA.t158 139.081
R3658 GNDA.t158 GNDA.t177 139.081
R3659 GNDA.t147 GNDA.t164 139.081
R3660 GNDA.t164 GNDA.t96 139.081
R3661 GNDA.t96 GNDA.t287 139.081
R3662 GNDA.n904 GNDA.n903 139.077
R3663 GNDA.n902 GNDA.n901 139.077
R3664 GNDA.n900 GNDA.n899 139.077
R3665 GNDA.n898 GNDA.n897 139.077
R3666 GNDA.n896 GNDA.n895 139.077
R3667 GNDA.n894 GNDA.n893 139.077
R3668 GNDA.n892 GNDA.n891 139.077
R3669 GNDA.n890 GNDA.n889 139.077
R3670 GNDA.n888 GNDA.n887 139.077
R3671 GNDA.n950 GNDA.t177 132.76
R3672 GNDA.n2331 GNDA.t147 132.76
R3673 GNDA.n649 GNDA.n401 131.893
R3674 GNDA.n1615 GNDA.n127 131.893
R3675 GNDA.t257 GNDA.n2359 130.731
R3676 GNDA.n2251 GNDA.t280 130.731
R3677 GNDA.n2286 GNDA.n2285 127.249
R3678 GNDA.t226 GNDA.n932 126.438
R3679 GNDA.t138 GNDA.n913 126.438
R3680 GNDA.n2117 GNDA.n2105 124.832
R3681 GNDA.n1988 GNDA.n1987 124.832
R3682 GNDA.n314 GNDA.n313 124.832
R3683 GNDA.n463 GNDA.n461 124.832
R3684 GNDA.n1661 GNDA.n1660 124.832
R3685 GNDA.n1644 GNDA.n1643 124.832
R3686 GNDA.n1438 GNDA.n1437 124.832
R3687 GNDA.n1216 GNDA.n1189 124.832
R3688 GNDA.n1032 GNDA.n958 124.832
R3689 GNDA.n1496 GNDA.n1192 124.832
R3690 GNDA.n376 GNDA.n174 124.832
R3691 GNDA.n1963 GNDA.n152 124.832
R3692 GNDA.n1248 GNDA.n1247 124.832
R3693 GNDA.n1388 GNDA.n1386 124.832
R3694 GNDA.n1562 GNDA.n609 124.832
R3695 GNDA.n651 GNDA.n648 124.832
R3696 GNDA.n1765 GNDA.n1764 124.832
R3697 GNDA.n1616 GNDA.n561 124.832
R3698 GNDA.t181 GNDA.t221 120.115
R3699 GNDA.t168 GNDA.t49 120.115
R3700 GNDA.n2426 GNDA.n2425 119.525
R3701 GNDA.n2249 GNDA.n2248 119.525
R3702 GNDA.n917 GNDA.n882 118.4
R3703 GNDA.n907 GNDA.n885 118.4
R3704 GNDA.n943 GNDA.n879 118.4
R3705 GNDA.n946 GNDA.n945 118.4
R3706 GNDA.n930 GNDA.n929 118.4
R3707 GNDA.n942 GNDA.n919 118.4
R3708 GNDA.n2233 GNDA.t110 115.79
R3709 GNDA.n2247 GNDA.t86 115.79
R3710 GNDA.n8 GNDA.t332 113.974
R3711 GNDA.n12 GNDA.t311 113.974
R3712 GNDA.n11 GNDA.t329 113.974
R3713 GNDA.n10 GNDA.t308 113.974
R3714 GNDA.n2482 GNDA.t336 113.974
R3715 GNDA.n2483 GNDA.t317 113.974
R3716 GNDA.n20 GNDA.t299 113.974
R3717 GNDA.n18 GNDA.t248 113.974
R3718 GNDA.n2478 GNDA.t238 113.974
R3719 GNDA.n2477 GNDA.t323 113.974
R3720 GNDA.t250 GNDA.n623 113.624
R3721 GNDA.n1030 GNDA.n957 113.624
R3722 GNDA.t252 GNDA.n1960 113.624
R3723 GNDA.t243 GNDA.n212 113.624
R3724 GNDA.n2241 GNDA.n2240 112.055
R3725 GNDA.n2474 GNDA.n28 108.8
R3726 GNDA.n2462 GNDA.n31 108.8
R3727 GNDA.n673 GNDA.n638 106.941
R3728 GNDA.n667 GNDA.n638 106.941
R3729 GNDA.n667 GNDA.n666 106.941
R3730 GNDA.n666 GNDA.n665 106.941
R3731 GNDA.n665 GNDA.n617 106.941
R3732 GNDA.n658 GNDA.n618 106.941
R3733 GNDA.n658 GNDA.n657 106.941
R3734 GNDA.n657 GNDA.n656 106.941
R3735 GNDA.n656 GNDA.n645 106.941
R3736 GNDA.n650 GNDA.n645 106.941
R3737 GNDA.n650 GNDA.n649 106.941
R3738 GNDA.n1590 GNDA.n576 106.941
R3739 GNDA.n1596 GNDA.n576 106.941
R3740 GNDA.n1597 GNDA.n1596 106.941
R3741 GNDA.n1598 GNDA.n1597 106.941
R3742 GNDA.n1598 GNDA.n359 106.941
R3743 GNDA.n1606 GNDA.n1605 106.941
R3744 GNDA.n1607 GNDA.n1606 106.941
R3745 GNDA.n1607 GNDA.n563 106.941
R3746 GNDA.n1613 GNDA.n563 106.941
R3747 GNDA.n1614 GNDA.n1613 106.941
R3748 GNDA.n1615 GNDA.n1614 106.941
R3749 GNDA.n1619 GNDA.n532 106.941
R3750 GNDA.n1626 GNDA.n532 106.941
R3751 GNDA.n1627 GNDA.n1626 106.941
R3752 GNDA.n1628 GNDA.n1627 106.941
R3753 GNDA.n1628 GNDA.n95 106.941
R3754 GNDA.n1635 GNDA.n96 106.941
R3755 GNDA.n1636 GNDA.n1635 106.941
R3756 GNDA.n1638 GNDA.n1636 106.941
R3757 GNDA.n1638 GNDA.n1637 106.941
R3758 GNDA.n1637 GNDA.n516 106.941
R3759 GNDA.n1568 GNDA.n401 103.144
R3760 GNDA.n2152 GNDA.n127 103.144
R3761 GNDA.n2284 GNDA.t322 101.194
R3762 GNDA.n932 GNDA.n927 101.15
R3763 GNDA.t34 GNDA.t141 101.15
R3764 GNDA.t99 GNDA.t209 101.15
R3765 GNDA.n913 GNDA.n911 101.15
R3766 GNDA.n1866 GNDA.n401 99.6276
R3767 GNDA.n2157 GNDA.n127 99.6276
R3768 GNDA.n2196 GNDA.n36 99.0842
R3769 GNDA.n38 GNDA.n37 99.0842
R3770 GNDA.n2396 GNDA.n2395 99.0842
R3771 GNDA.n2398 GNDA.n2397 99.0842
R3772 GNDA.n2400 GNDA.n2399 99.0842
R3773 GNDA.n2402 GNDA.n2401 99.0842
R3774 GNDA.n2404 GNDA.n2403 99.0842
R3775 GNDA.n2406 GNDA.n2405 99.0842
R3776 GNDA.n2408 GNDA.n2407 99.0842
R3777 GNDA.n2410 GNDA.n2409 99.0842
R3778 GNDA.n2412 GNDA.n2411 99.0842
R3779 GNDA.n2414 GNDA.n2413 99.0842
R3780 GNDA.n2102 GNDA.n2101 97.9524
R3781 GNDA.n2421 GNDA.n2420 95.101
R3782 GNDA.n2263 GNDA.n2197 95.101
R3783 GNDA.n2455 GNDA.t241 94.8842
R3784 GNDA.n2280 GNDA.t255 94.8842
R3785 GNDA.n2415 GNDA.t285 94.8842
R3786 GNDA.n2452 GNDA.t320 94.8842
R3787 GNDA.t325 GNDA.t226 94.8281
R3788 GNDA.t65 GNDA.t156 94.8281
R3789 GNDA.t354 GNDA.t160 94.8281
R3790 GNDA.t295 GNDA.t138 94.8281
R3791 GNDA.n2265 GNDA.n2264 94.601
R3792 GNDA.n2419 GNDA.n2418 94.601
R3793 GNDA.n1866 GNDA.t252 91.423
R3794 GNDA.t243 GNDA.n2157 91.423
R3795 GNDA.n2285 GNDA.n2284 89.9494
R3796 GNDA.t110 GNDA.t69 89.644
R3797 GNDA.t176 GNDA.t116 89.644
R3798 GNDA.n2429 GNDA.n2347 86.4005
R3799 GNDA.n2238 GNDA.n2237 86.4005
R3800 GNDA.n2323 GNDA.n2322 85.2845
R3801 GNDA.n63 GNDA.n62 85.2845
R3802 GNDA.n572 GNDA.n571 84.306
R3803 GNDA.t183 GNDA.t224 82.1844
R3804 GNDA.t113 GNDA.t174 82.1844
R3805 GNDA.t25 GNDA.t179 82.1844
R3806 GNDA.t166 GNDA.t15 82.1844
R3807 GNDA.t62 GNDA.t120 82.1737
R3808 GNDA.t122 GNDA.t77 82.1737
R3809 GNDA.t115 GNDA.t76 82.1737
R3810 GNDA.t83 GNDA.t272 82.1737
R3811 GNDA.t195 GNDA.t275 82.1737
R3812 GNDA.t346 GNDA.t345 82.1737
R3813 GNDA.t140 GNDA.t133 82.1737
R3814 GNDA.t135 GNDA.t127 82.1737
R3815 GNDA.n1536 GNDA.n827 80.9821
R3816 GNDA.t142 GNDA.n45 78.6626
R3817 GNDA.n2433 GNDA.t32 78.6626
R3818 GNDA.t61 GNDA.t260 78.4385
R3819 GNDA.t301 GNDA.t126 78.4385
R3820 GNDA.n178 GNDA.n147 76.3222
R3821 GNDA.n184 GNDA.n146 76.3222
R3822 GNDA.n190 GNDA.n145 76.3222
R3823 GNDA.n196 GNDA.n144 76.3222
R3824 GNDA.n200 GNDA.n128 76.3222
R3825 GNDA.n2121 GNDA.n2120 76.3222
R3826 GNDA.n227 GNDA.n148 76.3222
R3827 GNDA.n1970 GNDA.n1969 76.3222
R3828 GNDA.n1973 GNDA.n1972 76.3222
R3829 GNDA.n1978 GNDA.n1977 76.3222
R3830 GNDA.n1981 GNDA.n1980 76.3222
R3831 GNDA.n1986 GNDA.n1985 76.3222
R3832 GNDA.n345 GNDA.n116 76.3222
R3833 GNDA.n335 GNDA.n117 76.3222
R3834 GNDA.n332 GNDA.n118 76.3222
R3835 GNDA.n322 GNDA.n119 76.3222
R3836 GNDA.n319 GNDA.n120 76.3222
R3837 GNDA.n314 GNDA.n121 76.3222
R3838 GNDA.n1358 GNDA.n141 76.3222
R3839 GNDA.n1360 GNDA.n140 76.3222
R3840 GNDA.n1362 GNDA.n139 76.3222
R3841 GNDA.n1364 GNDA.n138 76.3222
R3842 GNDA.n229 GNDA.n129 76.3222
R3843 GNDA.n310 GNDA.n78 76.3222
R3844 GNDA.n484 GNDA.n483 76.3222
R3845 GNDA.n481 GNDA.n449 76.3222
R3846 GNDA.n477 GNDA.n476 76.3222
R3847 GNDA.n470 GNDA.n451 76.3222
R3848 GNDA.n469 GNDA.n468 76.3222
R3849 GNDA.n462 GNDA.n453 76.3222
R3850 GNDA.n1756 GNDA.n1755 76.3222
R3851 GNDA.n499 GNDA.n498 76.3222
R3852 GNDA.n1745 GNDA.n1744 76.3222
R3853 GNDA.n508 GNDA.n507 76.3222
R3854 GNDA.n1734 GNDA.n1733 76.3222
R3855 GNDA.n1661 GNDA.n513 76.3222
R3856 GNDA.n536 GNDA.n135 76.3222
R3857 GNDA.n538 GNDA.n134 76.3222
R3858 GNDA.n540 GNDA.n133 76.3222
R3859 GNDA.n543 GNDA.n132 76.3222
R3860 GNDA.n489 GNDA.n130 76.3222
R3861 GNDA.n514 GNDA.n101 76.3222
R3862 GNDA.n1415 GNDA.n809 76.3222
R3863 GNDA.n1420 GNDA.n1419 76.3222
R3864 GNDA.n1423 GNDA.n1422 76.3222
R3865 GNDA.n1428 GNDA.n1427 76.3222
R3866 GNDA.n1431 GNDA.n1430 76.3222
R3867 GNDA.n1436 GNDA.n1435 76.3222
R3868 GNDA.n822 GNDA.n820 76.3222
R3869 GNDA.n1439 GNDA.n599 76.3222
R3870 GNDA.n1444 GNDA.n598 76.3222
R3871 GNDA.n1450 GNDA.n597 76.3222
R3872 GNDA.n1456 GNDA.n596 76.3222
R3873 GNDA.n1068 GNDA.n841 76.3222
R3874 GNDA.n1495 GNDA.n606 76.3222
R3875 GNDA.n1491 GNDA.n605 76.3222
R3876 GNDA.n1487 GNDA.n604 76.3222
R3877 GNDA.n1483 GNDA.n603 76.3222
R3878 GNDA.n1479 GNDA.n602 76.3222
R3879 GNDA.n1028 GNDA.n601 76.3222
R3880 GNDA.n1469 GNDA.n415 76.3222
R3881 GNDA.n1471 GNDA.n414 76.3222
R3882 GNDA.n1473 GNDA.n413 76.3222
R3883 GNDA.n1475 GNDA.n412 76.3222
R3884 GNDA.n2154 GNDA.n2153 76.3222
R3885 GNDA.n176 GNDA.n159 76.3222
R3886 GNDA.n182 GNDA.n158 76.3222
R3887 GNDA.n188 GNDA.n157 76.3222
R3888 GNDA.n194 GNDA.n156 76.3222
R3889 GNDA.n2150 GNDA.n155 76.3222
R3890 GNDA.n1211 GNDA.n358 76.3222
R3891 GNDA.n1207 GNDA.n357 76.3222
R3892 GNDA.n1203 GNDA.n356 76.3222
R3893 GNDA.n1199 GNDA.n355 76.3222
R3894 GNDA.n1195 GNDA.n354 76.3222
R3895 GNDA.n1963 GNDA.n1962 76.3222
R3896 GNDA.n1213 GNDA.n358 76.3222
R3897 GNDA.n1210 GNDA.n357 76.3222
R3898 GNDA.n1206 GNDA.n356 76.3222
R3899 GNDA.n1202 GNDA.n355 76.3222
R3900 GNDA.n1198 GNDA.n354 76.3222
R3901 GNDA.n1962 GNDA.n353 76.3222
R3902 GNDA.n1868 GNDA.n402 76.3222
R3903 GNDA.n1867 GNDA.n404 76.3222
R3904 GNDA.n1474 GNDA.n412 76.3222
R3905 GNDA.n1472 GNDA.n413 76.3222
R3906 GNDA.n1470 GNDA.n414 76.3222
R3907 GNDA.n1468 GNDA.n415 76.3222
R3908 GNDA.n1492 GNDA.n606 76.3222
R3909 GNDA.n1488 GNDA.n605 76.3222
R3910 GNDA.n1484 GNDA.n604 76.3222
R3911 GNDA.n1480 GNDA.n603 76.3222
R3912 GNDA.n1476 GNDA.n602 76.3222
R3913 GNDA.n1028 GNDA.n607 76.3222
R3914 GNDA.n1343 GNDA.n1342 76.3222
R3915 GNDA.n1230 GNDA.n1229 76.3222
R3916 GNDA.n1332 GNDA.n1331 76.3222
R3917 GNDA.n1239 GNDA.n1238 76.3222
R3918 GNDA.n1321 GNDA.n1320 76.3222
R3919 GNDA.n1248 GNDA.n1246 76.3222
R3920 GNDA.n1446 GNDA.n421 76.3222
R3921 GNDA.n1452 GNDA.n420 76.3222
R3922 GNDA.n1458 GNDA.n419 76.3222
R3923 GNDA.n1463 GNDA.n418 76.3222
R3924 GNDA.n1220 GNDA.n411 76.3222
R3925 GNDA.n1385 GNDA.n165 76.3222
R3926 GNDA.n1381 GNDA.n164 76.3222
R3927 GNDA.n1377 GNDA.n163 76.3222
R3928 GNDA.n1373 GNDA.n162 76.3222
R3929 GNDA.n1369 GNDA.n161 76.3222
R3930 GNDA.n1243 GNDA.n160 76.3222
R3931 GNDA.n1406 GNDA.n1405 76.3222
R3932 GNDA.n1403 GNDA.n1402 76.3222
R3933 GNDA.n1398 GNDA.n1352 76.3222
R3934 GNDA.n1396 GNDA.n1395 76.3222
R3935 GNDA.n1391 GNDA.n1355 76.3222
R3936 GNDA.n1389 GNDA.n1388 76.3222
R3937 GNDA.n1407 GNDA.n1406 76.3222
R3938 GNDA.n1404 GNDA.n1403 76.3222
R3939 GNDA.n1352 GNDA.n1350 76.3222
R3940 GNDA.n1397 GNDA.n1396 76.3222
R3941 GNDA.n1355 GNDA.n1353 76.3222
R3942 GNDA.n1390 GNDA.n1389 76.3222
R3943 GNDA.n1246 GNDA.n1240 76.3222
R3944 GNDA.n1322 GNDA.n1321 76.3222
R3945 GNDA.n1238 GNDA.n1231 76.3222
R3946 GNDA.n1333 GNDA.n1332 76.3222
R3947 GNDA.n1229 GNDA.n1222 76.3222
R3948 GNDA.n1344 GNDA.n1343 76.3222
R3949 GNDA.n1218 GNDA.n608 76.3222
R3950 GNDA.n1464 GNDA.n417 76.3222
R3951 GNDA.n1459 GNDA.n418 76.3222
R3952 GNDA.n1453 GNDA.n419 76.3222
R3953 GNDA.n1447 GNDA.n420 76.3222
R3954 GNDA.n1441 GNDA.n421 76.3222
R3955 GNDA.n1443 GNDA.n599 76.3222
R3956 GNDA.n1449 GNDA.n598 76.3222
R3957 GNDA.n1455 GNDA.n597 76.3222
R3958 GNDA.n1460 GNDA.n596 76.3222
R3959 GNDA.n1465 GNDA.n600 76.3222
R3960 GNDA.n1416 GNDA.n1415 76.3222
R3961 GNDA.n1421 GNDA.n1420 76.3222
R3962 GNDA.n1422 GNDA.n1413 76.3222
R3963 GNDA.n1429 GNDA.n1428 76.3222
R3964 GNDA.n1430 GNDA.n1411 76.3222
R3965 GNDA.n1437 GNDA.n1436 76.3222
R3966 GNDA.n824 GNDA.n820 76.3222
R3967 GNDA.n1069 GNDA.n1068 76.3222
R3968 GNDA.n801 GNDA.n612 76.3222
R3969 GNDA.n791 GNDA.n613 76.3222
R3970 GNDA.n788 GNDA.n614 76.3222
R3971 GNDA.n778 GNDA.n615 76.3222
R3972 GNDA.n775 GNDA.n616 76.3222
R3973 GNDA.n1562 GNDA.n1561 76.3222
R3974 GNDA.n594 GNDA.n580 76.3222
R3975 GNDA.n593 GNDA.n582 76.3222
R3976 GNDA.n592 GNDA.n584 76.3222
R3977 GNDA.n591 GNDA.n586 76.3222
R3978 GNDA.n1569 GNDA.n588 76.3222
R3979 GNDA.n1566 GNDA.n589 76.3222
R3980 GNDA.n806 GNDA.n626 76.3222
R3981 GNDA.n594 GNDA.n581 76.3222
R3982 GNDA.n593 GNDA.n583 76.3222
R3983 GNDA.n592 GNDA.n585 76.3222
R3984 GNDA.n591 GNDA.n587 76.3222
R3985 GNDA.n1570 GNDA.n1569 76.3222
R3986 GNDA.n1860 GNDA.n1859 76.3222
R3987 GNDA.n434 GNDA.n433 76.3222
R3988 GNDA.n1849 GNDA.n1848 76.3222
R3989 GNDA.n443 GNDA.n442 76.3222
R3990 GNDA.n1838 GNDA.n1837 76.3222
R3991 GNDA.n1765 GNDA.n1763 76.3222
R3992 GNDA.n1586 GNDA.n406 76.3222
R3993 GNDA.n1582 GNDA.n407 76.3222
R3994 GNDA.n1578 GNDA.n408 76.3222
R3995 GNDA.n1574 GNDA.n409 76.3222
R3996 GNDA.n423 GNDA.n410 76.3222
R3997 GNDA.n1864 GNDA.n405 76.3222
R3998 GNDA.n1573 GNDA.n410 76.3222
R3999 GNDA.n1577 GNDA.n409 76.3222
R4000 GNDA.n1581 GNDA.n408 76.3222
R4001 GNDA.n1585 GNDA.n407 76.3222
R4002 GNDA.n1589 GNDA.n406 76.3222
R4003 GNDA.n562 GNDA.n171 76.3222
R4004 GNDA.n557 GNDA.n170 76.3222
R4005 GNDA.n553 GNDA.n169 76.3222
R4006 GNDA.n549 GNDA.n168 76.3222
R4007 GNDA.n545 GNDA.n167 76.3222
R4008 GNDA.n447 GNDA.n166 76.3222
R4009 GNDA.n1865 GNDA.n1864 76.3222
R4010 GNDA.n1763 GNDA.n444 76.3222
R4011 GNDA.n1839 GNDA.n1838 76.3222
R4012 GNDA.n442 GNDA.n435 76.3222
R4013 GNDA.n1850 GNDA.n1849 76.3222
R4014 GNDA.n433 GNDA.n426 76.3222
R4015 GNDA.n1861 GNDA.n1860 76.3222
R4016 GNDA.n629 GNDA.n626 76.3222
R4017 GNDA.n1561 GNDA.n611 76.3222
R4018 GNDA.n779 GNDA.n616 76.3222
R4019 GNDA.n787 GNDA.n615 76.3222
R4020 GNDA.n792 GNDA.n614 76.3222
R4021 GNDA.n800 GNDA.n613 76.3222
R4022 GNDA.n805 GNDA.n612 76.3222
R4023 GNDA.n1567 GNDA.n1566 76.3222
R4024 GNDA.n513 GNDA.n509 76.3222
R4025 GNDA.n1735 GNDA.n1734 76.3222
R4026 GNDA.n507 GNDA.n500 76.3222
R4027 GNDA.n1746 GNDA.n1745 76.3222
R4028 GNDA.n498 GNDA.n491 76.3222
R4029 GNDA.n1757 GNDA.n1756 76.3222
R4030 GNDA.n483 GNDA.n482 76.3222
R4031 GNDA.n478 GNDA.n449 76.3222
R4032 GNDA.n476 GNDA.n475 76.3222
R4033 GNDA.n471 GNDA.n470 76.3222
R4034 GNDA.n468 GNDA.n467 76.3222
R4035 GNDA.n463 GNDA.n462 76.3222
R4036 GNDA.n318 GNDA.n121 76.3222
R4037 GNDA.n323 GNDA.n120 76.3222
R4038 GNDA.n331 GNDA.n119 76.3222
R4039 GNDA.n336 GNDA.n118 76.3222
R4040 GNDA.n344 GNDA.n117 76.3222
R4041 GNDA.n348 GNDA.n116 76.3222
R4042 GNDA.n228 GNDA.n227 76.3222
R4043 GNDA.n1971 GNDA.n1970 76.3222
R4044 GNDA.n1972 GNDA.n225 76.3222
R4045 GNDA.n1979 GNDA.n1978 76.3222
R4046 GNDA.n1980 GNDA.n223 76.3222
R4047 GNDA.n1987 GNDA.n1986 76.3222
R4048 GNDA.n542 GNDA.n131 76.3222
R4049 GNDA.n541 GNDA.n132 76.3222
R4050 GNDA.n539 GNDA.n133 76.3222
R4051 GNDA.n537 GNDA.n134 76.3222
R4052 GNDA.n535 GNDA.n135 76.3222
R4053 GNDA.n1365 GNDA.n137 76.3222
R4054 GNDA.n1363 GNDA.n138 76.3222
R4055 GNDA.n1361 GNDA.n139 76.3222
R4056 GNDA.n1359 GNDA.n140 76.3222
R4057 GNDA.n1357 GNDA.n141 76.3222
R4058 GNDA.n197 GNDA.n143 76.3222
R4059 GNDA.n191 GNDA.n144 76.3222
R4060 GNDA.n185 GNDA.n145 76.3222
R4061 GNDA.n179 GNDA.n146 76.3222
R4062 GNDA.n149 GNDA.n147 76.3222
R4063 GNDA.n558 GNDA.n171 76.3222
R4064 GNDA.n554 GNDA.n170 76.3222
R4065 GNDA.n550 GNDA.n169 76.3222
R4066 GNDA.n546 GNDA.n168 76.3222
R4067 GNDA.n487 GNDA.n167 76.3222
R4068 GNDA.n447 GNDA.n172 76.3222
R4069 GNDA.n1382 GNDA.n165 76.3222
R4070 GNDA.n1378 GNDA.n164 76.3222
R4071 GNDA.n1374 GNDA.n163 76.3222
R4072 GNDA.n1370 GNDA.n162 76.3222
R4073 GNDA.n1366 GNDA.n161 76.3222
R4074 GNDA.n1243 GNDA.n173 76.3222
R4075 GNDA.n2153 GNDA.n153 76.3222
R4076 GNDA.n181 GNDA.n159 76.3222
R4077 GNDA.n187 GNDA.n158 76.3222
R4078 GNDA.n193 GNDA.n157 76.3222
R4079 GNDA.n198 GNDA.n156 76.3222
R4080 GNDA.n2151 GNDA.n2150 76.3222
R4081 GNDA.n1659 GNDA.n514 76.3222
R4082 GNDA.n312 GNDA.n310 76.3222
R4083 GNDA.n2120 GNDA.n2005 76.3222
R4084 GNDA.n2374 GNDA.n2373 76.1251
R4085 GNDA.n739 GNDA.n738 76.062
R4086 GNDA.n738 GNDA.n737 76.062
R4087 GNDA.n1800 GNDA.n1799 76.062
R4088 GNDA.n1799 GNDA.n1798 76.062
R4089 GNDA.n1696 GNDA.n1695 76.062
R4090 GNDA.n1695 GNDA.n1694 76.062
R4091 GNDA.n1150 GNDA.n1129 76.062
R4092 GNDA.n1151 GNDA.n1150 76.062
R4093 GNDA.n1283 GNDA.n1282 76.062
R4094 GNDA.n1282 GNDA.n1281 76.062
R4095 GNDA.n272 GNDA.n252 76.062
R4096 GNDA.n273 GNDA.n272 76.062
R4097 GNDA.n991 GNDA.n972 76.062
R4098 GNDA.n992 GNDA.n991 76.062
R4099 GNDA.n1907 GNDA.n390 76.062
R4100 GNDA.n1908 GNDA.n1907 76.062
R4101 GNDA.n2063 GNDA.n2062 76.062
R4102 GNDA.n2062 GNDA.n2061 76.062
R4103 GNDA.n935 GNDA.t225 75.8626
R4104 GNDA.n940 GNDA.t79 75.8626
R4105 GNDA.n940 GNDA.t223 75.8626
R4106 GNDA.n909 GNDA.t14 75.8626
R4107 GNDA.t216 GNDA.n909 75.8626
R4108 GNDA.n910 GNDA.t72 75.8626
R4109 GNDA.n721 GNDA.n698 74.5978
R4110 GNDA.n722 GNDA.n721 74.5978
R4111 GNDA.n1856 GNDA.n428 74.5978
R4112 GNDA.n1783 GNDA.n428 74.5978
R4113 GNDA.n1752 GNDA.n493 74.5978
R4114 GNDA.n1679 GNDA.n493 74.5978
R4115 GNDA.n1134 GNDA.n1099 74.5978
R4116 GNDA.n1135 GNDA.n1134 74.5978
R4117 GNDA.n1339 GNDA.n1224 74.5978
R4118 GNDA.n1266 GNDA.n1224 74.5978
R4119 GNDA.n256 GNDA.n233 74.5978
R4120 GNDA.n257 GNDA.n256 74.5978
R4121 GNDA.n1062 GNDA.n846 74.5978
R4122 GNDA.n976 GNDA.n846 74.5978
R4123 GNDA.n1891 GNDA.n1890 74.5978
R4124 GNDA.n1892 GNDA.n1891 74.5978
R4125 GNDA.n2045 GNDA.n208 74.5978
R4126 GNDA.n2046 GNDA.n2045 74.5978
R4127 GNDA.t250 GNDA.n617 72.4823
R4128 GNDA.t252 GNDA.n359 72.4823
R4129 GNDA.t243 GNDA.n95 72.4823
R4130 GNDA.n2115 GNDA.n84 71.1128
R4131 GNDA.t131 GNDA.t61 70.9682
R4132 GNDA.t245 GNDA.t83 70.9682
R4133 GNDA.t313 GNDA.t195 70.9682
R4134 GNDA.t126 GNDA.t27 70.9682
R4135 GNDA.t222 GNDA.t183 69.5407
R4136 GNDA.t174 GNDA.t222 69.5407
R4137 GNDA.t162 GNDA.n949 69.5407
R4138 GNDA.n949 GNDA.t94 69.5407
R4139 GNDA.t179 GNDA.t22 69.5407
R4140 GNDA.t22 GNDA.t166 69.5407
R4141 GNDA.n724 GNDA.t293 65.8183
R4142 GNDA.n730 GNDA.t293 65.8183
R4143 GNDA.n732 GNDA.t293 65.8183
R4144 GNDA.n740 GNDA.t293 65.8183
R4145 GNDA.n746 GNDA.t293 65.8183
R4146 GNDA.n748 GNDA.t293 65.8183
R4147 GNDA.n754 GNDA.t293 65.8183
R4148 GNDA.n771 GNDA.t293 65.8183
R4149 GNDA.n765 GNDA.t293 65.8183
R4150 GNDA.n763 GNDA.t293 65.8183
R4151 GNDA.n757 GNDA.t293 65.8183
R4152 GNDA.n1785 GNDA.t292 65.8183
R4153 GNDA.n1791 GNDA.t292 65.8183
R4154 GNDA.n1793 GNDA.t292 65.8183
R4155 GNDA.n1801 GNDA.t292 65.8183
R4156 GNDA.n1807 GNDA.t292 65.8183
R4157 GNDA.n1809 GNDA.t292 65.8183
R4158 GNDA.n1815 GNDA.t292 65.8183
R4159 GNDA.n1832 GNDA.t292 65.8183
R4160 GNDA.n1826 GNDA.t292 65.8183
R4161 GNDA.n1824 GNDA.t292 65.8183
R4162 GNDA.n1818 GNDA.t292 65.8183
R4163 GNDA.n1681 GNDA.t267 65.8183
R4164 GNDA.n1687 GNDA.t267 65.8183
R4165 GNDA.n1689 GNDA.t267 65.8183
R4166 GNDA.n1697 GNDA.t267 65.8183
R4167 GNDA.n1703 GNDA.t267 65.8183
R4168 GNDA.n1705 GNDA.t267 65.8183
R4169 GNDA.n1711 GNDA.t267 65.8183
R4170 GNDA.n1728 GNDA.t267 65.8183
R4171 GNDA.n1722 GNDA.t267 65.8183
R4172 GNDA.n1720 GNDA.t267 65.8183
R4173 GNDA.n1714 GNDA.t267 65.8183
R4174 GNDA.n1140 GNDA.t249 65.8183
R4175 GNDA.n1142 GNDA.t249 65.8183
R4176 GNDA.n1148 GNDA.t249 65.8183
R4177 GNDA.n1156 GNDA.t249 65.8183
R4178 GNDA.n1158 GNDA.t249 65.8183
R4179 GNDA.n1164 GNDA.t249 65.8183
R4180 GNDA.n1166 GNDA.t249 65.8183
R4181 GNDA.n1183 GNDA.t249 65.8183
R4182 GNDA.n1181 GNDA.t249 65.8183
R4183 GNDA.n1175 GNDA.t249 65.8183
R4184 GNDA.n1172 GNDA.t249 65.8183
R4185 GNDA.n1268 GNDA.t251 65.8183
R4186 GNDA.n1274 GNDA.t251 65.8183
R4187 GNDA.n1276 GNDA.t251 65.8183
R4188 GNDA.n1284 GNDA.t251 65.8183
R4189 GNDA.n1290 GNDA.t251 65.8183
R4190 GNDA.n1292 GNDA.t251 65.8183
R4191 GNDA.n1298 GNDA.t251 65.8183
R4192 GNDA.n1315 GNDA.t251 65.8183
R4193 GNDA.n1309 GNDA.t251 65.8183
R4194 GNDA.n1307 GNDA.t251 65.8183
R4195 GNDA.n1301 GNDA.t251 65.8183
R4196 GNDA.n262 GNDA.t333 65.8183
R4197 GNDA.n264 GNDA.t333 65.8183
R4198 GNDA.n270 GNDA.t333 65.8183
R4199 GNDA.n278 GNDA.t333 65.8183
R4200 GNDA.n280 GNDA.t333 65.8183
R4201 GNDA.n286 GNDA.t333 65.8183
R4202 GNDA.n288 GNDA.t333 65.8183
R4203 GNDA.n306 GNDA.t333 65.8183
R4204 GNDA.n303 GNDA.t333 65.8183
R4205 GNDA.n297 GNDA.t333 65.8183
R4206 GNDA.n294 GNDA.t333 65.8183
R4207 GNDA.n981 GNDA.t266 65.8183
R4208 GNDA.n983 GNDA.t266 65.8183
R4209 GNDA.n989 GNDA.t266 65.8183
R4210 GNDA.n997 GNDA.t266 65.8183
R4211 GNDA.n999 GNDA.t266 65.8183
R4212 GNDA.n1005 GNDA.t266 65.8183
R4213 GNDA.n1007 GNDA.t266 65.8183
R4214 GNDA.n1025 GNDA.t266 65.8183
R4215 GNDA.n1022 GNDA.t266 65.8183
R4216 GNDA.n1016 GNDA.t266 65.8183
R4217 GNDA.n1013 GNDA.t266 65.8183
R4218 GNDA.n1897 GNDA.t265 65.8183
R4219 GNDA.n1899 GNDA.t265 65.8183
R4220 GNDA.n1905 GNDA.t265 65.8183
R4221 GNDA.n1913 GNDA.t265 65.8183
R4222 GNDA.n1915 GNDA.t265 65.8183
R4223 GNDA.n1921 GNDA.t265 65.8183
R4224 GNDA.n1923 GNDA.t265 65.8183
R4225 GNDA.n1941 GNDA.t265 65.8183
R4226 GNDA.n1938 GNDA.t265 65.8183
R4227 GNDA.n1932 GNDA.t265 65.8183
R4228 GNDA.n1929 GNDA.t265 65.8183
R4229 GNDA.n2048 GNDA.t242 65.8183
R4230 GNDA.n2054 GNDA.t242 65.8183
R4231 GNDA.n2056 GNDA.t242 65.8183
R4232 GNDA.n2064 GNDA.t242 65.8183
R4233 GNDA.n2070 GNDA.t242 65.8183
R4234 GNDA.n2072 GNDA.t242 65.8183
R4235 GNDA.n2078 GNDA.t242 65.8183
R4236 GNDA.n2095 GNDA.t242 65.8183
R4237 GNDA.n2089 GNDA.t242 65.8183
R4238 GNDA.n2087 GNDA.t242 65.8183
R4239 GNDA.n2081 GNDA.t242 65.8183
R4240 GNDA.n2028 GNDA.t242 65.8183
R4241 GNDA.n2012 GNDA.t242 65.8183
R4242 GNDA.n2015 GNDA.t242 65.8183
R4243 GNDA.n2137 GNDA.t242 65.8183
R4244 GNDA.n380 GNDA.t265 65.8183
R4245 GNDA.n1955 GNDA.t265 65.8183
R4246 GNDA.n1879 GNDA.t265 65.8183
R4247 GNDA.n1877 GNDA.t265 65.8183
R4248 GNDA.n962 GNDA.t266 65.8183
R4249 GNDA.n1045 GNDA.t266 65.8183
R4250 GNDA.n854 GNDA.t266 65.8183
R4251 GNDA.n1060 GNDA.t266 65.8183
R4252 GNDA.n242 GNDA.t333 65.8183
R4253 GNDA.n327 GNDA.t333 65.8183
R4254 GNDA.n237 GNDA.t333 65.8183
R4255 GNDA.n340 GNDA.t333 65.8183
R4256 GNDA.n1242 GNDA.t251 65.8183
R4257 GNDA.n1326 GNDA.t251 65.8183
R4258 GNDA.n1233 GNDA.t251 65.8183
R4259 GNDA.n1337 GNDA.t251 65.8183
R4260 GNDA.n1507 GNDA.t249 65.8183
R4261 GNDA.n1117 GNDA.t249 65.8183
R4262 GNDA.n1111 GNDA.t249 65.8183
R4263 GNDA.n1525 GNDA.t249 65.8183
R4264 GNDA.n511 GNDA.t267 65.8183
R4265 GNDA.n1739 GNDA.t267 65.8183
R4266 GNDA.n502 GNDA.t267 65.8183
R4267 GNDA.n1750 GNDA.t267 65.8183
R4268 GNDA.n446 GNDA.t292 65.8183
R4269 GNDA.n1843 GNDA.t292 65.8183
R4270 GNDA.n437 GNDA.t292 65.8183
R4271 GNDA.n1854 GNDA.t292 65.8183
R4272 GNDA.n706 GNDA.t293 65.8183
R4273 GNDA.n783 GNDA.t293 65.8183
R4274 GNDA.n702 GNDA.t293 65.8183
R4275 GNDA.n796 GNDA.t293 65.8183
R4276 GNDA.n2491 GNDA.n21 64.0005
R4277 GNDA.n2491 GNDA.n19 64.0005
R4278 GNDA.t223 GNDA.n939 63.2189
R4279 GNDA.t14 GNDA.n56 63.2189
R4280 GNDA.t250 GNDA.n590 60.9488
R4281 GNDA.t252 GNDA.n154 60.9488
R4282 GNDA.n2456 GNDA.n35 60.8005
R4283 GNDA.n1658 GNDA.n123 60.3563
R4284 GNDA.n311 GNDA.n125 60.3563
R4285 GNDA.n2116 GNDA.n2004 60.3563
R4286 GNDA.n1645 GNDA.n517 57.3684
R4287 GNDA.n459 GNDA.n122 57.3684
R4288 GNDA.n1990 GNDA.n1989 57.3684
R4289 GNDA.t224 GNDA.t325 56.897
R4290 GNDA.t156 GNDA.t113 56.897
R4291 GNDA.n938 GNDA.t269 56.897
R4292 GNDA.t287 GNDA.n2330 56.897
R4293 GNDA.t160 GNDA.t25 56.897
R4294 GNDA.t15 GNDA.t295 56.897
R4295 GNDA.t189 GNDA.t62 56.0277
R4296 GNDA.t17 GNDA.t115 56.0277
R4297 GNDA.t192 GNDA.t346 56.0277
R4298 GNDA.t127 GNDA.t108 56.0277
R4299 GNDA.n2045 GNDA.t242 55.2026
R4300 GNDA.n1891 GNDA.t265 55.2026
R4301 GNDA.t266 GNDA.n846 55.2026
R4302 GNDA.n256 GNDA.t333 55.2026
R4303 GNDA.t251 GNDA.n1224 55.2026
R4304 GNDA.n1134 GNDA.t249 55.2026
R4305 GNDA.t267 GNDA.n493 55.2026
R4306 GNDA.t292 GNDA.n428 55.2026
R4307 GNDA.n721 GNDA.t293 55.2026
R4308 GNDA.n738 GNDA.t293 54.4705
R4309 GNDA.n1799 GNDA.t292 54.4705
R4310 GNDA.n1695 GNDA.t267 54.4705
R4311 GNDA.n1150 GNDA.t249 54.4705
R4312 GNDA.n1282 GNDA.t251 54.4705
R4313 GNDA.n272 GNDA.t333 54.4705
R4314 GNDA.n991 GNDA.t266 54.4705
R4315 GNDA.n1907 GNDA.t265 54.4705
R4316 GNDA.n2062 GNDA.t242 54.4705
R4317 GNDA.n2281 GNDA.n35 54.4005
R4318 GNDA.n521 GNDA.n88 53.7829
R4319 GNDA.n2189 GNDA.n89 53.7829
R4320 GNDA.n2183 GNDA.n89 53.7829
R4321 GNDA.n2182 GNDA.n2181 53.7829
R4322 GNDA.n2181 GNDA.n98 53.7829
R4323 GNDA.n2175 GNDA.n98 53.7829
R4324 GNDA.n1658 GNDA.n1657 53.7829
R4325 GNDA.n459 GNDA.n458 53.7829
R4326 GNDA.n458 GNDA.n109 53.7829
R4327 GNDA.n2165 GNDA.n110 53.7829
R4328 GNDA.n2159 GNDA.n110 53.7829
R4329 GNDA.n2305 GNDA.n79 53.7829
R4330 GNDA.n311 GNDA.n80 53.7829
R4331 GNDA.n1990 GNDA.n219 53.7829
R4332 GNDA.n1996 GNDA.n219 53.7829
R4333 GNDA.n1997 GNDA.n1996 53.7829
R4334 GNDA.n1998 GNDA.n1997 53.7829
R4335 GNDA.n1998 GNDA.n213 53.7829
R4336 GNDA.n2130 GNDA.n214 53.7829
R4337 GNDA.n2124 GNDA.n2123 53.7829
R4338 GNDA.n2123 GNDA.n2122 53.7829
R4339 GNDA.n2122 GNDA.n2004 53.7829
R4340 GNDA.n796 GNDA.n795 53.3664
R4341 GNDA.n703 GNDA.n702 53.3664
R4342 GNDA.n783 GNDA.n782 53.3664
R4343 GNDA.n773 GNDA.n706 53.3664
R4344 GNDA.n757 GNDA.n756 53.3664
R4345 GNDA.n763 GNDA.n762 53.3664
R4346 GNDA.n766 GNDA.n765 53.3664
R4347 GNDA.n771 GNDA.n770 53.3664
R4348 GNDA.n741 GNDA.n740 53.3664
R4349 GNDA.n746 GNDA.n745 53.3664
R4350 GNDA.n749 GNDA.n748 53.3664
R4351 GNDA.n754 GNDA.n753 53.3664
R4352 GNDA.n732 GNDA.n717 53.3664
R4353 GNDA.n731 GNDA.n730 53.3664
R4354 GNDA.n724 GNDA.n719 53.3664
R4355 GNDA.n725 GNDA.n724 53.3664
R4356 GNDA.n730 GNDA.n729 53.3664
R4357 GNDA.n733 GNDA.n732 53.3664
R4358 GNDA.n740 GNDA.n715 53.3664
R4359 GNDA.n747 GNDA.n746 53.3664
R4360 GNDA.n748 GNDA.n713 53.3664
R4361 GNDA.n755 GNDA.n754 53.3664
R4362 GNDA.n772 GNDA.n771 53.3664
R4363 GNDA.n765 GNDA.n708 53.3664
R4364 GNDA.n764 GNDA.n763 53.3664
R4365 GNDA.n758 GNDA.n757 53.3664
R4366 GNDA.n1854 GNDA.n1853 53.3664
R4367 GNDA.n1845 GNDA.n437 53.3664
R4368 GNDA.n1843 GNDA.n1842 53.3664
R4369 GNDA.n1834 GNDA.n446 53.3664
R4370 GNDA.n1818 GNDA.n1817 53.3664
R4371 GNDA.n1824 GNDA.n1823 53.3664
R4372 GNDA.n1827 GNDA.n1826 53.3664
R4373 GNDA.n1832 GNDA.n1831 53.3664
R4374 GNDA.n1802 GNDA.n1801 53.3664
R4375 GNDA.n1807 GNDA.n1806 53.3664
R4376 GNDA.n1810 GNDA.n1809 53.3664
R4377 GNDA.n1815 GNDA.n1814 53.3664
R4378 GNDA.n1793 GNDA.n1778 53.3664
R4379 GNDA.n1792 GNDA.n1791 53.3664
R4380 GNDA.n1785 GNDA.n1780 53.3664
R4381 GNDA.n1786 GNDA.n1785 53.3664
R4382 GNDA.n1791 GNDA.n1790 53.3664
R4383 GNDA.n1794 GNDA.n1793 53.3664
R4384 GNDA.n1801 GNDA.n1776 53.3664
R4385 GNDA.n1808 GNDA.n1807 53.3664
R4386 GNDA.n1809 GNDA.n1774 53.3664
R4387 GNDA.n1816 GNDA.n1815 53.3664
R4388 GNDA.n1833 GNDA.n1832 53.3664
R4389 GNDA.n1826 GNDA.n1769 53.3664
R4390 GNDA.n1825 GNDA.n1824 53.3664
R4391 GNDA.n1819 GNDA.n1818 53.3664
R4392 GNDA.n1750 GNDA.n1749 53.3664
R4393 GNDA.n1741 GNDA.n502 53.3664
R4394 GNDA.n1739 GNDA.n1738 53.3664
R4395 GNDA.n1730 GNDA.n511 53.3664
R4396 GNDA.n1714 GNDA.n1713 53.3664
R4397 GNDA.n1720 GNDA.n1719 53.3664
R4398 GNDA.n1723 GNDA.n1722 53.3664
R4399 GNDA.n1728 GNDA.n1727 53.3664
R4400 GNDA.n1698 GNDA.n1697 53.3664
R4401 GNDA.n1703 GNDA.n1702 53.3664
R4402 GNDA.n1706 GNDA.n1705 53.3664
R4403 GNDA.n1711 GNDA.n1710 53.3664
R4404 GNDA.n1689 GNDA.n1674 53.3664
R4405 GNDA.n1688 GNDA.n1687 53.3664
R4406 GNDA.n1681 GNDA.n1676 53.3664
R4407 GNDA.n1682 GNDA.n1681 53.3664
R4408 GNDA.n1687 GNDA.n1686 53.3664
R4409 GNDA.n1690 GNDA.n1689 53.3664
R4410 GNDA.n1697 GNDA.n1672 53.3664
R4411 GNDA.n1704 GNDA.n1703 53.3664
R4412 GNDA.n1705 GNDA.n1670 53.3664
R4413 GNDA.n1712 GNDA.n1711 53.3664
R4414 GNDA.n1729 GNDA.n1728 53.3664
R4415 GNDA.n1722 GNDA.n1665 53.3664
R4416 GNDA.n1721 GNDA.n1720 53.3664
R4417 GNDA.n1715 GNDA.n1714 53.3664
R4418 GNDA.n1525 GNDA.n1524 53.3664
R4419 GNDA.n1115 GNDA.n1111 53.3664
R4420 GNDA.n1509 GNDA.n1117 53.3664
R4421 GNDA.n1507 GNDA.n1506 53.3664
R4422 GNDA.n1172 GNDA.n1171 53.3664
R4423 GNDA.n1176 GNDA.n1175 53.3664
R4424 GNDA.n1181 GNDA.n1180 53.3664
R4425 GNDA.n1184 GNDA.n1183 53.3664
R4426 GNDA.n1156 GNDA.n1155 53.3664
R4427 GNDA.n1159 GNDA.n1158 53.3664
R4428 GNDA.n1164 GNDA.n1163 53.3664
R4429 GNDA.n1167 GNDA.n1166 53.3664
R4430 GNDA.n1149 GNDA.n1148 53.3664
R4431 GNDA.n1142 GNDA.n1131 53.3664
R4432 GNDA.n1141 GNDA.n1140 53.3664
R4433 GNDA.n1140 GNDA.n1139 53.3664
R4434 GNDA.n1143 GNDA.n1142 53.3664
R4435 GNDA.n1148 GNDA.n1147 53.3664
R4436 GNDA.n1157 GNDA.n1156 53.3664
R4437 GNDA.n1158 GNDA.n1127 53.3664
R4438 GNDA.n1165 GNDA.n1164 53.3664
R4439 GNDA.n1166 GNDA.n1125 53.3664
R4440 GNDA.n1183 GNDA.n1119 53.3664
R4441 GNDA.n1182 GNDA.n1181 53.3664
R4442 GNDA.n1175 GNDA.n1122 53.3664
R4443 GNDA.n1173 GNDA.n1172 53.3664
R4444 GNDA.n1337 GNDA.n1336 53.3664
R4445 GNDA.n1328 GNDA.n1233 53.3664
R4446 GNDA.n1326 GNDA.n1325 53.3664
R4447 GNDA.n1317 GNDA.n1242 53.3664
R4448 GNDA.n1301 GNDA.n1300 53.3664
R4449 GNDA.n1307 GNDA.n1306 53.3664
R4450 GNDA.n1310 GNDA.n1309 53.3664
R4451 GNDA.n1315 GNDA.n1314 53.3664
R4452 GNDA.n1285 GNDA.n1284 53.3664
R4453 GNDA.n1290 GNDA.n1289 53.3664
R4454 GNDA.n1293 GNDA.n1292 53.3664
R4455 GNDA.n1298 GNDA.n1297 53.3664
R4456 GNDA.n1276 GNDA.n1261 53.3664
R4457 GNDA.n1275 GNDA.n1274 53.3664
R4458 GNDA.n1268 GNDA.n1263 53.3664
R4459 GNDA.n1269 GNDA.n1268 53.3664
R4460 GNDA.n1274 GNDA.n1273 53.3664
R4461 GNDA.n1277 GNDA.n1276 53.3664
R4462 GNDA.n1284 GNDA.n1259 53.3664
R4463 GNDA.n1291 GNDA.n1290 53.3664
R4464 GNDA.n1292 GNDA.n1257 53.3664
R4465 GNDA.n1299 GNDA.n1298 53.3664
R4466 GNDA.n1316 GNDA.n1315 53.3664
R4467 GNDA.n1309 GNDA.n1252 53.3664
R4468 GNDA.n1308 GNDA.n1307 53.3664
R4469 GNDA.n1302 GNDA.n1301 53.3664
R4470 GNDA.n340 GNDA.n339 53.3664
R4471 GNDA.n238 GNDA.n237 53.3664
R4472 GNDA.n327 GNDA.n326 53.3664
R4473 GNDA.n243 GNDA.n242 53.3664
R4474 GNDA.n294 GNDA.n293 53.3664
R4475 GNDA.n298 GNDA.n297 53.3664
R4476 GNDA.n303 GNDA.n302 53.3664
R4477 GNDA.n306 GNDA.n305 53.3664
R4478 GNDA.n278 GNDA.n277 53.3664
R4479 GNDA.n281 GNDA.n280 53.3664
R4480 GNDA.n286 GNDA.n285 53.3664
R4481 GNDA.n289 GNDA.n288 53.3664
R4482 GNDA.n271 GNDA.n270 53.3664
R4483 GNDA.n264 GNDA.n254 53.3664
R4484 GNDA.n263 GNDA.n262 53.3664
R4485 GNDA.n262 GNDA.n261 53.3664
R4486 GNDA.n265 GNDA.n264 53.3664
R4487 GNDA.n270 GNDA.n269 53.3664
R4488 GNDA.n279 GNDA.n278 53.3664
R4489 GNDA.n280 GNDA.n250 53.3664
R4490 GNDA.n287 GNDA.n286 53.3664
R4491 GNDA.n288 GNDA.n248 53.3664
R4492 GNDA.n307 GNDA.n306 53.3664
R4493 GNDA.n304 GNDA.n303 53.3664
R4494 GNDA.n297 GNDA.n245 53.3664
R4495 GNDA.n295 GNDA.n294 53.3664
R4496 GNDA.n1060 GNDA.n1059 53.3664
R4497 GNDA.n1047 GNDA.n854 53.3664
R4498 GNDA.n1045 GNDA.n1044 53.3664
R4499 GNDA.n963 GNDA.n962 53.3664
R4500 GNDA.n1013 GNDA.n1012 53.3664
R4501 GNDA.n1017 GNDA.n1016 53.3664
R4502 GNDA.n1022 GNDA.n1021 53.3664
R4503 GNDA.n1025 GNDA.n1024 53.3664
R4504 GNDA.n997 GNDA.n996 53.3664
R4505 GNDA.n1000 GNDA.n999 53.3664
R4506 GNDA.n1005 GNDA.n1004 53.3664
R4507 GNDA.n1008 GNDA.n1007 53.3664
R4508 GNDA.n990 GNDA.n989 53.3664
R4509 GNDA.n983 GNDA.n974 53.3664
R4510 GNDA.n982 GNDA.n981 53.3664
R4511 GNDA.n981 GNDA.n980 53.3664
R4512 GNDA.n984 GNDA.n983 53.3664
R4513 GNDA.n989 GNDA.n988 53.3664
R4514 GNDA.n998 GNDA.n997 53.3664
R4515 GNDA.n999 GNDA.n970 53.3664
R4516 GNDA.n1006 GNDA.n1005 53.3664
R4517 GNDA.n1007 GNDA.n968 53.3664
R4518 GNDA.n1026 GNDA.n1025 53.3664
R4519 GNDA.n1023 GNDA.n1022 53.3664
R4520 GNDA.n1016 GNDA.n965 53.3664
R4521 GNDA.n1014 GNDA.n1013 53.3664
R4522 GNDA.n1878 GNDA.n1877 53.3664
R4523 GNDA.n1879 GNDA.n370 53.3664
R4524 GNDA.n1955 GNDA.n1954 53.3664
R4525 GNDA.n381 GNDA.n380 53.3664
R4526 GNDA.n1929 GNDA.n1928 53.3664
R4527 GNDA.n1933 GNDA.n1932 53.3664
R4528 GNDA.n1938 GNDA.n1937 53.3664
R4529 GNDA.n1941 GNDA.n1940 53.3664
R4530 GNDA.n1913 GNDA.n1912 53.3664
R4531 GNDA.n1916 GNDA.n1915 53.3664
R4532 GNDA.n1921 GNDA.n1920 53.3664
R4533 GNDA.n1924 GNDA.n1923 53.3664
R4534 GNDA.n1906 GNDA.n1905 53.3664
R4535 GNDA.n1899 GNDA.n392 53.3664
R4536 GNDA.n1898 GNDA.n1897 53.3664
R4537 GNDA.n1897 GNDA.n1896 53.3664
R4538 GNDA.n1900 GNDA.n1899 53.3664
R4539 GNDA.n1905 GNDA.n1904 53.3664
R4540 GNDA.n1914 GNDA.n1913 53.3664
R4541 GNDA.n1915 GNDA.n388 53.3664
R4542 GNDA.n1922 GNDA.n1921 53.3664
R4543 GNDA.n1923 GNDA.n386 53.3664
R4544 GNDA.n1942 GNDA.n1941 53.3664
R4545 GNDA.n1939 GNDA.n1938 53.3664
R4546 GNDA.n1932 GNDA.n383 53.3664
R4547 GNDA.n1930 GNDA.n1929 53.3664
R4548 GNDA.n2137 GNDA.n2136 53.3664
R4549 GNDA.n2017 GNDA.n2015 53.3664
R4550 GNDA.n2026 GNDA.n2012 53.3664
R4551 GNDA.n2097 GNDA.n2028 53.3664
R4552 GNDA.n2081 GNDA.n2080 53.3664
R4553 GNDA.n2087 GNDA.n2086 53.3664
R4554 GNDA.n2090 GNDA.n2089 53.3664
R4555 GNDA.n2095 GNDA.n2094 53.3664
R4556 GNDA.n2065 GNDA.n2064 53.3664
R4557 GNDA.n2070 GNDA.n2069 53.3664
R4558 GNDA.n2073 GNDA.n2072 53.3664
R4559 GNDA.n2078 GNDA.n2077 53.3664
R4560 GNDA.n2056 GNDA.n2040 53.3664
R4561 GNDA.n2055 GNDA.n2054 53.3664
R4562 GNDA.n2048 GNDA.n2042 53.3664
R4563 GNDA.n2049 GNDA.n2048 53.3664
R4564 GNDA.n2054 GNDA.n2053 53.3664
R4565 GNDA.n2057 GNDA.n2056 53.3664
R4566 GNDA.n2064 GNDA.n2038 53.3664
R4567 GNDA.n2071 GNDA.n2070 53.3664
R4568 GNDA.n2072 GNDA.n2036 53.3664
R4569 GNDA.n2079 GNDA.n2078 53.3664
R4570 GNDA.n2096 GNDA.n2095 53.3664
R4571 GNDA.n2089 GNDA.n2031 53.3664
R4572 GNDA.n2088 GNDA.n2087 53.3664
R4573 GNDA.n2082 GNDA.n2081 53.3664
R4574 GNDA.n2028 GNDA.n2027 53.3664
R4575 GNDA.n2016 GNDA.n2012 53.3664
R4576 GNDA.n2015 GNDA.n209 53.3664
R4577 GNDA.n2138 GNDA.n2137 53.3664
R4578 GNDA.n380 GNDA.n371 53.3664
R4579 GNDA.n1956 GNDA.n1955 53.3664
R4580 GNDA.n1880 GNDA.n1879 53.3664
R4581 GNDA.n1877 GNDA.n396 53.3664
R4582 GNDA.n962 GNDA.n856 53.3664
R4583 GNDA.n1046 GNDA.n1045 53.3664
R4584 GNDA.n854 GNDA.n848 53.3664
R4585 GNDA.n1061 GNDA.n1060 53.3664
R4586 GNDA.n242 GNDA.n239 53.3664
R4587 GNDA.n328 GNDA.n327 53.3664
R4588 GNDA.n237 GNDA.n234 53.3664
R4589 GNDA.n341 GNDA.n340 53.3664
R4590 GNDA.n1242 GNDA.n1235 53.3664
R4591 GNDA.n1327 GNDA.n1326 53.3664
R4592 GNDA.n1233 GNDA.n1226 53.3664
R4593 GNDA.n1338 GNDA.n1337 53.3664
R4594 GNDA.n1508 GNDA.n1507 53.3664
R4595 GNDA.n1117 GNDA.n1116 53.3664
R4596 GNDA.n1111 GNDA.n1100 53.3664
R4597 GNDA.n1526 GNDA.n1525 53.3664
R4598 GNDA.n511 GNDA.n504 53.3664
R4599 GNDA.n1740 GNDA.n1739 53.3664
R4600 GNDA.n502 GNDA.n495 53.3664
R4601 GNDA.n1751 GNDA.n1750 53.3664
R4602 GNDA.n446 GNDA.n439 53.3664
R4603 GNDA.n1844 GNDA.n1843 53.3664
R4604 GNDA.n437 GNDA.n430 53.3664
R4605 GNDA.n1855 GNDA.n1854 53.3664
R4606 GNDA.n706 GNDA.n704 53.3664
R4607 GNDA.n784 GNDA.n783 53.3664
R4608 GNDA.n702 GNDA.n699 53.3664
R4609 GNDA.n797 GNDA.n796 53.3664
R4610 GNDA.t31 GNDA.n2376 53.2877
R4611 GNDA.t68 GNDA.t73 52.4707
R4612 GNDA.t203 GNDA.t47 52.4707
R4613 GNDA.t328 GNDA.t1 52.4707
R4614 GNDA.t243 GNDA.n122 51.9902
R4615 GNDA.n2312 GNDA.n73 51.9902
R4616 GNDA.t243 GNDA.n123 51.3926
R4617 GNDA.t243 GNDA.n125 51.3926
R4618 GNDA.n2484 GNDA.n21 51.2005
R4619 GNDA.n2479 GNDA.n19 51.2005
R4620 GNDA.n2496 GNDA.t283 48.7228
R4621 GNDA.n2360 GNDA.t121 48.5574
R4622 GNDA.n2232 GNDA.t176 48.5574
R4623 GNDA.n2216 GNDA.t86 48.5574
R4624 GNDA.n2260 GNDA.t89 48.5574
R4625 GNDA.n2470 GNDA.t107 48.0005
R4626 GNDA.n2470 GNDA.t102 48.0005
R4627 GNDA.n2467 GNDA.t215 48.0005
R4628 GNDA.n2467 GNDA.t57 48.0005
R4629 GNDA.n2466 GNDA.t74 48.0005
R4630 GNDA.n2466 GNDA.t48 48.0005
R4631 GNDA.n2464 GNDA.t348 48.0005
R4632 GNDA.n2464 GNDA.t20 48.0005
R4633 GNDA.n2463 GNDA.t59 48.0005
R4634 GNDA.n2463 GNDA.t10 48.0005
R4635 GNDA.n2166 GNDA.n109 46.0144
R4636 GNDA.t212 GNDA.t143 44.9749
R4637 GNDA.t105 GNDA.t54 44.9749
R4638 GNDA.t92 GNDA.t350 44.9749
R4639 GNDA.t353 GNDA.t198 44.9749
R4640 GNDA.t44 GNDA.t218 44.9749
R4641 GNDA.t349 GNDA.t40 44.9749
R4642 GNDA.t187 GNDA.t12 44.9749
R4643 GNDA.t16 GNDA.t6 44.9749
R4644 GNDA.t88 GNDA.t207 44.9749
R4645 GNDA.t331 GNDA.t36 44.9749
R4646 GNDA.n2426 GNDA.n45 44.8222
R4647 GNDA.n2248 GNDA.n2247 44.8222
R4648 GNDA.n2380 GNDA.n2371 44.8005
R4649 GNDA.n2230 GNDA.n2229 44.8005
R4650 GNDA.t170 GNDA.t65 44.2534
R4651 GNDA.t172 GNDA.t354 44.2534
R4652 GNDA.n2378 GNDA.t2 43.1378
R4653 GNDA.n2195 GNDA.t352 41.2271
R4654 GNDA.n2489 GNDA.t213 41.2271
R4655 GNDA.n2448 GNDA.t201 41.2271
R4656 GNDA.t211 GNDA.n2495 41.2271
R4657 GNDA.n2495 GNDA.t335 41.2271
R4658 GNDA.t85 GNDA.t340 41.0871
R4659 GNDA.t340 GNDA.t122 41.0871
R4660 GNDA.t69 GNDA.n2232 41.0871
R4661 GNDA.t103 GNDA.n2216 41.0871
R4662 GNDA.t136 GNDA.t140 41.0871
R4663 GNDA.t136 GNDA.t355 41.0871
R4664 GNDA.n2305 GNDA.n2304 40.0385
R4665 GNDA.n2291 GNDA.n2189 37.6482
R4666 GNDA.t322 GNDA.t254 37.4792
R4667 GNDA.t21 GNDA.t240 37.4792
R4668 GNDA.t80 GNDA.t263 37.4792
R4669 GNDA.t9 GNDA.t185 37.4792
R4670 GNDA.t87 GNDA.t19 37.4792
R4671 GNDA.t200 GNDA.t106 37.4792
R4672 GNDA.t50 GNDA.t101 37.4792
R4673 GNDA.t39 GNDA.t214 37.4792
R4674 GNDA.t237 GNDA.t56 37.4792
R4675 GNDA.t45 GNDA.t151 37.4792
R4676 GNDA.t201 GNDA.t212 37.4792
R4677 GNDA.n2512 GNDA.n2511 36.9067
R4678 GNDA.n2277 GNDA.n2276 36.6567
R4679 GNDA.n2434 GNDA.n2342 36.2041
R4680 GNDA.t250 GNDA.n618 34.459
R4681 GNDA.t243 GNDA.n96 34.459
R4682 GNDA.n520 GNDA.n517 34.0627
R4683 GNDA.n2311 GNDA.n74 34.0627
R4684 GNDA.n1989 GNDA.n124 34.0627
R4685 GNDA.t352 GNDA.n2193 33.7313
R4686 GNDA.n2460 GNDA.t338 33.7313
R4687 GNDA.n2459 GNDA.t58 33.7313
R4688 GNDA.n42 GNDA.t347 33.7313
R4689 GNDA.t42 GNDA.n2476 33.7313
R4690 GNDA.n2360 GNDA.t85 33.6168
R4691 GNDA.n2260 GNDA.t355 33.6168
R4692 GNDA.n2384 GNDA.t142 32.9878
R4693 GNDA.t210 GNDA.n2377 32.9878
R4694 GNDA.t225 GNDA.t181 31.6097
R4695 GNDA.t149 GNDA.t34 31.6097
R4696 GNDA.t154 GNDA.t99 31.6097
R4697 GNDA.t72 GNDA.t168 31.6097
R4698 GNDA.t240 GNDA.t307 29.9835
R4699 GNDA.t263 GNDA.t217 29.9835
R4700 GNDA.t8 GNDA.t58 29.9835
R4701 GNDA.t11 GNDA.t9 29.9835
R4702 GNDA.t347 GNDA.t235 29.9835
R4703 GNDA.t298 GNDA.t310 29.9835
R4704 GNDA.n2359 GNDA.n44 29.8817
R4705 GNDA.n2251 GNDA.n2192 29.8817
R4706 GNDA.n2429 GNDA.n2428 28.413
R4707 GNDA.n2237 GNDA.n2204 28.413
R4708 GNDA.n2314 GNDA.n69 28.1318
R4709 GNDA.n2183 GNDA.t243 28.0869
R4710 GNDA.n2159 GNDA.t243 28.0869
R4711 GNDA.t243 GNDA.n213 28.0869
R4712 GNDA.n2423 GNDA.n2388 28.038
R4713 GNDA.n2214 GNDA.n2198 28.038
R4714 GNDA.n2377 GNDA.t31 27.9128
R4715 GNDA.n945 GNDA.n917 27.8193
R4716 GNDA.n943 GNDA.n942 27.8193
R4717 GNDA.n736 GNDA.n716 27.5561
R4718 GNDA.n1797 GNDA.n1777 27.5561
R4719 GNDA.n1693 GNDA.n1673 27.5561
R4720 GNDA.n1153 GNDA.n1152 27.5561
R4721 GNDA.n1280 GNDA.n1260 27.5561
R4722 GNDA.n275 GNDA.n274 27.5561
R4723 GNDA.n994 GNDA.n993 27.5561
R4724 GNDA.n1910 GNDA.n1909 27.5561
R4725 GNDA.n2060 GNDA.n2039 27.5561
R4726 GNDA.n1568 GNDA.n590 26.9584
R4727 GNDA.n2152 GNDA.n154 26.9584
R4728 GNDA.n2489 GNDA.t66 26.2356
R4729 GNDA.n2439 GNDA.t335 26.2356
R4730 GNDA.t121 GNDA.t189 26.1465
R4731 GNDA.t77 GNDA.t17 26.1465
R4732 GNDA.t133 GNDA.t192 26.1465
R4733 GNDA.t108 GNDA.t89 26.1465
R4734 GNDA.t243 GNDA.n2182 25.6965
R4735 GNDA.t243 GNDA.n73 25.6965
R4736 GNDA.t243 GNDA.n2130 25.6965
R4737 GNDA.n2391 GNDA.n2390 25.6005
R4738 GNDA.n2258 GNDA.n2255 25.6005
R4739 GNDA.n935 GNDA.n934 25.2879
R4740 GNDA.n914 GNDA.n910 25.2879
R4741 GNDA.n903 GNDA.t180 24.0005
R4742 GNDA.n903 GNDA.t167 24.0005
R4743 GNDA.n901 GNDA.t173 24.0005
R4744 GNDA.n901 GNDA.t161 24.0005
R4745 GNDA.n899 GNDA.t155 24.0005
R4746 GNDA.n899 GNDA.t169 24.0005
R4747 GNDA.n897 GNDA.t165 24.0005
R4748 GNDA.n897 GNDA.t97 24.0005
R4749 GNDA.n895 GNDA.t95 24.0005
R4750 GNDA.n895 GNDA.t148 24.0005
R4751 GNDA.n893 GNDA.t178 24.0005
R4752 GNDA.n893 GNDA.t163 24.0005
R4753 GNDA.n891 GNDA.t118 24.0005
R4754 GNDA.n891 GNDA.t159 24.0005
R4755 GNDA.n889 GNDA.t182 24.0005
R4756 GNDA.n889 GNDA.t150 24.0005
R4757 GNDA.n887 GNDA.t157 24.0005
R4758 GNDA.n887 GNDA.t171 24.0005
R4759 GNDA.n886 GNDA.t184 24.0005
R4760 GNDA.n886 GNDA.t175 24.0005
R4761 GNDA.t70 GNDA.t53 23.9038
R4762 GNDA.t252 GNDA.n360 23.765
R4763 GNDA.n712 GNDA.n711 23.6449
R4764 GNDA.n1773 GNDA.n1772 23.6449
R4765 GNDA.n1669 GNDA.n1668 23.6449
R4766 GNDA.n1170 GNDA.n1169 23.6449
R4767 GNDA.n1256 GNDA.n1255 23.6449
R4768 GNDA.n292 GNDA.n291 23.6449
R4769 GNDA.n1011 GNDA.n1010 23.6449
R4770 GNDA.n1927 GNDA.n1926 23.6449
R4771 GNDA.n2035 GNDA.n2034 23.6449
R4772 GNDA.n2486 GNDA.n0 23.488
R4773 GNDA.t143 GNDA.t316 22.4877
R4774 GNDA.t350 GNDA.t35 22.4877
R4775 GNDA.t198 GNDA.t104 22.4877
R4776 GNDA.t218 GNDA.t344 22.4877
R4777 GNDA.t12 GNDA.t93 22.4877
R4778 GNDA.t6 GNDA.t46 22.4877
R4779 GNDA.t207 GNDA.t26 22.4877
R4780 GNDA.t36 GNDA.t145 22.4877
R4781 GNDA.t283 GNDA.t211 22.4877
R4782 GNDA.n2281 GNDA.n2280 22.4005
R4783 GNDA.n2456 GNDA.n2455 22.4005
R4784 GNDA.n2452 GNDA.n2451 22.4005
R4785 GNDA.n2415 GNDA.n40 22.4005
R4786 GNDA.n2388 GNDA.n2387 22.4005
R4787 GNDA.n2245 GNDA.n2214 22.4005
R4788 GNDA.n15 GNDA.n14 22.4005
R4789 GNDA.n14 GNDA.n13 22.4005
R4790 GNDA.n2316 GNDA.n2315 21.4917
R4791 GNDA.n28 GNDA.n27 21.3338
R4792 GNDA.n31 GNDA.n29 21.3338
R4793 GNDA.n885 GNDA.n884 21.3338
R4794 GNDA.n882 GNDA.n881 21.3338
R4795 GNDA.n946 GNDA.n880 21.3338
R4796 GNDA.n879 GNDA.n878 21.3338
R4797 GNDA.n919 GNDA.n918 21.3338
R4798 GNDA.n929 GNDA.n928 21.3338
R4799 GNDA.n2349 GNDA.n2348 21.3338
R4800 GNDA.n2356 GNDA.n2354 21.3338
R4801 GNDA.n2363 GNDA.n2362 21.3338
R4802 GNDA.n2392 GNDA.n2389 21.3338
R4803 GNDA.n2207 GNDA.n2206 21.3338
R4804 GNDA.n2210 GNDA.n2209 21.3338
R4805 GNDA.n2203 GNDA.n2202 21.3338
R4806 GNDA.n2257 GNDA.n2256 21.3338
R4807 GNDA.n9 GNDA.n8 21.3338
R4808 GNDA.n13 GNDA.n12 21.3338
R4809 GNDA.n15 GNDA.n11 21.3338
R4810 GNDA.n16 GNDA.n10 21.3338
R4811 GNDA.n2485 GNDA.n2482 21.3338
R4812 GNDA.n2484 GNDA.n2483 21.3338
R4813 GNDA.n21 GNDA.n20 21.3338
R4814 GNDA.n19 GNDA.n18 21.3338
R4815 GNDA.n2479 GNDA.n2478 21.3338
R4816 GNDA.n2480 GNDA.n2477 21.3338
R4817 GNDA.n907 GNDA.n906 21.1792
R4818 GNDA.n2384 GNDA.n2383 20.3004
R4819 GNDA GNDA.n2513 20.281
R4820 GNDA.n521 GNDA.n520 19.7207
R4821 GNDA.n79 GNDA.n74 19.7207
R4822 GNDA.n2510 GNDA.t114 19.7005
R4823 GNDA.n2510 GNDA.t234 19.7005
R4824 GNDA.n2508 GNDA.t81 19.7005
R4825 GNDA.n2508 GNDA.t129 19.7005
R4826 GNDA.n2506 GNDA.t23 19.7005
R4827 GNDA.n2506 GNDA.t82 19.7005
R4828 GNDA.n2504 GNDA.t84 19.7005
R4829 GNDA.n2504 GNDA.t63 19.7005
R4830 GNDA.n2502 GNDA.t123 19.7005
R4831 GNDA.n2502 GNDA.t78 19.7005
R4832 GNDA.n2501 GNDA.t230 19.7005
R4833 GNDA.n2501 GNDA.t130 19.7005
R4834 GNDA.n2275 GNDA.t233 19.7005
R4835 GNDA.n2275 GNDA.t194 19.7005
R4836 GNDA.n2273 GNDA.t128 19.7005
R4837 GNDA.n2273 GNDA.t186 19.7005
R4838 GNDA.n2271 GNDA.t64 19.7005
R4839 GNDA.n2271 GNDA.t191 19.7005
R4840 GNDA.n2269 GNDA.t134 19.7005
R4841 GNDA.n2269 GNDA.t75 19.7005
R4842 GNDA.n2267 GNDA.t188 19.7005
R4843 GNDA.n2267 GNDA.t139 19.7005
R4844 GNDA.n2266 GNDA.t125 19.7005
R4845 GNDA.n2266 GNDA.t228 19.7005
R4846 GNDA.n2320 GNDA.n2319 19.4279
R4847 GNDA.n2371 GNDA.n2345 19.3505
R4848 GNDA.n2231 GNDA.n2230 19.3505
R4849 GNDA.n2492 GNDA.n2491 19.288
R4850 GNDA.n2170 GNDA.n2169 19.2005
R4851 GNDA.n2112 GNDA.n83 19.2005
R4852 GNDA.n2315 GNDA.n66 19.2005
R4853 GNDA.n1650 GNDA.n70 19.2005
R4854 GNDA.n2323 GNDA.n55 19.2005
R4855 GNDA.n865 GNDA.n63 19.2005
R4856 GNDA.n2390 GNDA.n2350 19.1005
R4857 GNDA.n2255 GNDA.n2254 19.1005
R4858 GNDA.t221 GNDA.t149 18.966
R4859 GNDA.t49 GNDA.t154 18.966
R4860 GNDA.t40 GNDA.n2441 18.7399
R4861 GNDA.t243 GNDA.n124 17.928
R4862 GNDA.n2325 GNDA.n63 17.613
R4863 GNDA.n569 GNDA.n65 17.4917
R4864 GNDA.t111 GNDA.t210 17.2554
R4865 GNDA.n1602 GNDA.n573 16.9605
R4866 GNDA.n1557 GNDA.n811 16.9379
R4867 GNDA.n1534 GNDA.n1091 16.9379
R4868 GNDA.n671 GNDA.n636 16.9379
R4869 GNDA.n2291 GNDA.n88 16.1352
R4870 GNDA.n1657 GNDA.t33 16.1352
R4871 GNDA.n2124 GNDA.t53 16.1352
R4872 GNDA.n736 GNDA.n735 16.0005
R4873 GNDA.n735 GNDA.n734 16.0005
R4874 GNDA.n734 GNDA.n718 16.0005
R4875 GNDA.n728 GNDA.n718 16.0005
R4876 GNDA.n728 GNDA.n727 16.0005
R4877 GNDA.n727 GNDA.n726 16.0005
R4878 GNDA.n726 GNDA.n720 16.0005
R4879 GNDA.n720 GNDA.n695 16.0005
R4880 GNDA.n742 GNDA.n716 16.0005
R4881 GNDA.n743 GNDA.n742 16.0005
R4882 GNDA.n744 GNDA.n743 16.0005
R4883 GNDA.n744 GNDA.n714 16.0005
R4884 GNDA.n750 GNDA.n714 16.0005
R4885 GNDA.n751 GNDA.n750 16.0005
R4886 GNDA.n752 GNDA.n751 16.0005
R4887 GNDA.n752 GNDA.n712 16.0005
R4888 GNDA.n759 GNDA.n711 16.0005
R4889 GNDA.n760 GNDA.n759 16.0005
R4890 GNDA.n761 GNDA.n760 16.0005
R4891 GNDA.n761 GNDA.n709 16.0005
R4892 GNDA.n768 GNDA.n767 16.0005
R4893 GNDA.n769 GNDA.n768 16.0005
R4894 GNDA.n769 GNDA.n707 16.0005
R4895 GNDA.n1797 GNDA.n1796 16.0005
R4896 GNDA.n1796 GNDA.n1795 16.0005
R4897 GNDA.n1795 GNDA.n1779 16.0005
R4898 GNDA.n1789 GNDA.n1779 16.0005
R4899 GNDA.n1789 GNDA.n1788 16.0005
R4900 GNDA.n1788 GNDA.n1787 16.0005
R4901 GNDA.n1787 GNDA.n1781 16.0005
R4902 GNDA.n1782 GNDA.n1781 16.0005
R4903 GNDA.n1803 GNDA.n1777 16.0005
R4904 GNDA.n1804 GNDA.n1803 16.0005
R4905 GNDA.n1805 GNDA.n1804 16.0005
R4906 GNDA.n1805 GNDA.n1775 16.0005
R4907 GNDA.n1811 GNDA.n1775 16.0005
R4908 GNDA.n1812 GNDA.n1811 16.0005
R4909 GNDA.n1813 GNDA.n1812 16.0005
R4910 GNDA.n1813 GNDA.n1773 16.0005
R4911 GNDA.n1820 GNDA.n1772 16.0005
R4912 GNDA.n1821 GNDA.n1820 16.0005
R4913 GNDA.n1822 GNDA.n1821 16.0005
R4914 GNDA.n1822 GNDA.n1770 16.0005
R4915 GNDA.n1829 GNDA.n1828 16.0005
R4916 GNDA.n1830 GNDA.n1829 16.0005
R4917 GNDA.n1830 GNDA.n1768 16.0005
R4918 GNDA.n1693 GNDA.n1692 16.0005
R4919 GNDA.n1692 GNDA.n1691 16.0005
R4920 GNDA.n1691 GNDA.n1675 16.0005
R4921 GNDA.n1685 GNDA.n1675 16.0005
R4922 GNDA.n1685 GNDA.n1684 16.0005
R4923 GNDA.n1684 GNDA.n1683 16.0005
R4924 GNDA.n1683 GNDA.n1677 16.0005
R4925 GNDA.n1678 GNDA.n1677 16.0005
R4926 GNDA.n1699 GNDA.n1673 16.0005
R4927 GNDA.n1700 GNDA.n1699 16.0005
R4928 GNDA.n1701 GNDA.n1700 16.0005
R4929 GNDA.n1701 GNDA.n1671 16.0005
R4930 GNDA.n1707 GNDA.n1671 16.0005
R4931 GNDA.n1708 GNDA.n1707 16.0005
R4932 GNDA.n1709 GNDA.n1708 16.0005
R4933 GNDA.n1709 GNDA.n1669 16.0005
R4934 GNDA.n1716 GNDA.n1668 16.0005
R4935 GNDA.n1717 GNDA.n1716 16.0005
R4936 GNDA.n1718 GNDA.n1717 16.0005
R4937 GNDA.n1718 GNDA.n1666 16.0005
R4938 GNDA.n1725 GNDA.n1724 16.0005
R4939 GNDA.n1726 GNDA.n1725 16.0005
R4940 GNDA.n1726 GNDA.n1664 16.0005
R4941 GNDA.n569 GNDA.n568 16.0005
R4942 GNDA.n573 GNDA.n568 16.0005
R4943 GNDA.n1152 GNDA.n1130 16.0005
R4944 GNDA.n1146 GNDA.n1130 16.0005
R4945 GNDA.n1146 GNDA.n1145 16.0005
R4946 GNDA.n1145 GNDA.n1144 16.0005
R4947 GNDA.n1144 GNDA.n1132 16.0005
R4948 GNDA.n1138 GNDA.n1132 16.0005
R4949 GNDA.n1138 GNDA.n1137 16.0005
R4950 GNDA.n1137 GNDA.n1136 16.0005
R4951 GNDA.n1154 GNDA.n1153 16.0005
R4952 GNDA.n1154 GNDA.n1128 16.0005
R4953 GNDA.n1160 GNDA.n1128 16.0005
R4954 GNDA.n1161 GNDA.n1160 16.0005
R4955 GNDA.n1162 GNDA.n1161 16.0005
R4956 GNDA.n1162 GNDA.n1126 16.0005
R4957 GNDA.n1168 GNDA.n1126 16.0005
R4958 GNDA.n1169 GNDA.n1168 16.0005
R4959 GNDA.n1170 GNDA.n1124 16.0005
R4960 GNDA.n1124 GNDA.n1123 16.0005
R4961 GNDA.n1177 GNDA.n1123 16.0005
R4962 GNDA.n1178 GNDA.n1177 16.0005
R4963 GNDA.n1179 GNDA.n1121 16.0005
R4964 GNDA.n1185 GNDA.n1121 16.0005
R4965 GNDA.n1186 GNDA.n1185 16.0005
R4966 GNDA.n1280 GNDA.n1279 16.0005
R4967 GNDA.n1279 GNDA.n1278 16.0005
R4968 GNDA.n1278 GNDA.n1262 16.0005
R4969 GNDA.n1272 GNDA.n1262 16.0005
R4970 GNDA.n1272 GNDA.n1271 16.0005
R4971 GNDA.n1271 GNDA.n1270 16.0005
R4972 GNDA.n1270 GNDA.n1264 16.0005
R4973 GNDA.n1265 GNDA.n1264 16.0005
R4974 GNDA.n1286 GNDA.n1260 16.0005
R4975 GNDA.n1287 GNDA.n1286 16.0005
R4976 GNDA.n1288 GNDA.n1287 16.0005
R4977 GNDA.n1288 GNDA.n1258 16.0005
R4978 GNDA.n1294 GNDA.n1258 16.0005
R4979 GNDA.n1295 GNDA.n1294 16.0005
R4980 GNDA.n1296 GNDA.n1295 16.0005
R4981 GNDA.n1296 GNDA.n1256 16.0005
R4982 GNDA.n1303 GNDA.n1255 16.0005
R4983 GNDA.n1304 GNDA.n1303 16.0005
R4984 GNDA.n1305 GNDA.n1304 16.0005
R4985 GNDA.n1305 GNDA.n1253 16.0005
R4986 GNDA.n1312 GNDA.n1311 16.0005
R4987 GNDA.n1313 GNDA.n1312 16.0005
R4988 GNDA.n1313 GNDA.n1251 16.0005
R4989 GNDA.n274 GNDA.n253 16.0005
R4990 GNDA.n268 GNDA.n253 16.0005
R4991 GNDA.n268 GNDA.n267 16.0005
R4992 GNDA.n267 GNDA.n266 16.0005
R4993 GNDA.n266 GNDA.n255 16.0005
R4994 GNDA.n260 GNDA.n255 16.0005
R4995 GNDA.n260 GNDA.n259 16.0005
R4996 GNDA.n259 GNDA.n230 16.0005
R4997 GNDA.n276 GNDA.n275 16.0005
R4998 GNDA.n276 GNDA.n251 16.0005
R4999 GNDA.n282 GNDA.n251 16.0005
R5000 GNDA.n283 GNDA.n282 16.0005
R5001 GNDA.n284 GNDA.n283 16.0005
R5002 GNDA.n284 GNDA.n249 16.0005
R5003 GNDA.n290 GNDA.n249 16.0005
R5004 GNDA.n291 GNDA.n290 16.0005
R5005 GNDA.n292 GNDA.n247 16.0005
R5006 GNDA.n247 GNDA.n246 16.0005
R5007 GNDA.n299 GNDA.n246 16.0005
R5008 GNDA.n300 GNDA.n299 16.0005
R5009 GNDA.n301 GNDA.n244 16.0005
R5010 GNDA.n244 GNDA.n241 16.0005
R5011 GNDA.n308 GNDA.n241 16.0005
R5012 GNDA.n993 GNDA.n973 16.0005
R5013 GNDA.n987 GNDA.n973 16.0005
R5014 GNDA.n987 GNDA.n986 16.0005
R5015 GNDA.n986 GNDA.n985 16.0005
R5016 GNDA.n985 GNDA.n975 16.0005
R5017 GNDA.n979 GNDA.n975 16.0005
R5018 GNDA.n979 GNDA.n978 16.0005
R5019 GNDA.n978 GNDA.n844 16.0005
R5020 GNDA.n995 GNDA.n994 16.0005
R5021 GNDA.n995 GNDA.n971 16.0005
R5022 GNDA.n1001 GNDA.n971 16.0005
R5023 GNDA.n1002 GNDA.n1001 16.0005
R5024 GNDA.n1003 GNDA.n1002 16.0005
R5025 GNDA.n1003 GNDA.n969 16.0005
R5026 GNDA.n1009 GNDA.n969 16.0005
R5027 GNDA.n1010 GNDA.n1009 16.0005
R5028 GNDA.n1011 GNDA.n967 16.0005
R5029 GNDA.n967 GNDA.n966 16.0005
R5030 GNDA.n1018 GNDA.n966 16.0005
R5031 GNDA.n1019 GNDA.n1018 16.0005
R5032 GNDA.n1020 GNDA.n964 16.0005
R5033 GNDA.n964 GNDA.n961 16.0005
R5034 GNDA.n1027 GNDA.n961 16.0005
R5035 GNDA.n1909 GNDA.n391 16.0005
R5036 GNDA.n1903 GNDA.n391 16.0005
R5037 GNDA.n1903 GNDA.n1902 16.0005
R5038 GNDA.n1902 GNDA.n1901 16.0005
R5039 GNDA.n1901 GNDA.n393 16.0005
R5040 GNDA.n1895 GNDA.n393 16.0005
R5041 GNDA.n1895 GNDA.n1894 16.0005
R5042 GNDA.n1894 GNDA.n1893 16.0005
R5043 GNDA.n1911 GNDA.n1910 16.0005
R5044 GNDA.n1911 GNDA.n389 16.0005
R5045 GNDA.n1917 GNDA.n389 16.0005
R5046 GNDA.n1918 GNDA.n1917 16.0005
R5047 GNDA.n1919 GNDA.n1918 16.0005
R5048 GNDA.n1919 GNDA.n387 16.0005
R5049 GNDA.n1925 GNDA.n387 16.0005
R5050 GNDA.n1926 GNDA.n1925 16.0005
R5051 GNDA.n1927 GNDA.n385 16.0005
R5052 GNDA.n385 GNDA.n384 16.0005
R5053 GNDA.n1934 GNDA.n384 16.0005
R5054 GNDA.n1935 GNDA.n1934 16.0005
R5055 GNDA.n1936 GNDA.n382 16.0005
R5056 GNDA.n382 GNDA.n379 16.0005
R5057 GNDA.n1943 GNDA.n379 16.0005
R5058 GNDA.n2060 GNDA.n2059 16.0005
R5059 GNDA.n2059 GNDA.n2058 16.0005
R5060 GNDA.n2058 GNDA.n2041 16.0005
R5061 GNDA.n2052 GNDA.n2041 16.0005
R5062 GNDA.n2052 GNDA.n2051 16.0005
R5063 GNDA.n2051 GNDA.n2050 16.0005
R5064 GNDA.n2050 GNDA.n2043 16.0005
R5065 GNDA.n2044 GNDA.n2043 16.0005
R5066 GNDA.n2066 GNDA.n2039 16.0005
R5067 GNDA.n2067 GNDA.n2066 16.0005
R5068 GNDA.n2068 GNDA.n2067 16.0005
R5069 GNDA.n2068 GNDA.n2037 16.0005
R5070 GNDA.n2074 GNDA.n2037 16.0005
R5071 GNDA.n2075 GNDA.n2074 16.0005
R5072 GNDA.n2076 GNDA.n2075 16.0005
R5073 GNDA.n2076 GNDA.n2035 16.0005
R5074 GNDA.n2083 GNDA.n2034 16.0005
R5075 GNDA.n2084 GNDA.n2083 16.0005
R5076 GNDA.n2085 GNDA.n2084 16.0005
R5077 GNDA.n2085 GNDA.n2032 16.0005
R5078 GNDA.n2092 GNDA.n2091 16.0005
R5079 GNDA.n2093 GNDA.n2092 16.0005
R5080 GNDA.n2093 GNDA.n2030 16.0005
R5081 GNDA.n2328 GNDA.n2327 15.363
R5082 GNDA.n2327 GNDA.n60 15.363
R5083 GNDA.t307 GNDA.t80 14.992
R5084 GNDA.t217 GNDA.t146 14.992
R5085 GNDA.t185 GNDA.t8 14.992
R5086 GNDA.t220 GNDA.t11 14.992
R5087 GNDA.t235 GNDA.t87 14.992
R5088 GNDA.t19 GNDA.t319 14.992
R5089 GNDA.t319 GNDA.t153 14.992
R5090 GNDA.t153 GNDA.t200 14.992
R5091 GNDA.t106 GNDA.t90 14.992
R5092 GNDA.t90 GNDA.t204 14.992
R5093 GNDA.t101 GNDA.t4 14.992
R5094 GNDA.t4 GNDA.t24 14.992
R5095 GNDA.t24 GNDA.t39 14.992
R5096 GNDA.t214 GNDA.t205 14.992
R5097 GNDA.t205 GNDA.t60 14.992
R5098 GNDA.t60 GNDA.t237 14.992
R5099 GNDA.t56 GNDA.t342 14.992
R5100 GNDA.t342 GNDA.t68 14.992
R5101 GNDA.t73 GNDA.t196 14.992
R5102 GNDA.t196 GNDA.t203 14.992
R5103 GNDA.t47 GNDA.t51 14.992
R5104 GNDA.t51 GNDA.t328 14.992
R5105 GNDA.t1 GNDA.t66 14.992
R5106 GNDA.t213 GNDA.t42 14.992
R5107 GNDA.t151 GNDA.t298 14.992
R5108 GNDA.t316 GNDA.t105 14.992
R5109 GNDA.t38 GNDA.t92 14.992
R5110 GNDA.t35 GNDA.t353 14.992
R5111 GNDA.t104 GNDA.t44 14.992
R5112 GNDA.t344 GNDA.t349 14.992
R5113 GNDA.t93 GNDA.t16 14.992
R5114 GNDA.t46 GNDA.t88 14.992
R5115 GNDA.t26 GNDA.t331 14.992
R5116 GNDA.n2286 GNDA.n2192 14.9411
R5117 GNDA GNDA.n2320 14.6989
R5118 GNDA.n2422 GNDA.n2421 14.0505
R5119 GNDA.n2263 GNDA.n2262 14.0505
R5120 GNDA.n767 GNDA 14.0449
R5121 GNDA.n1828 GNDA 14.0449
R5122 GNDA.n1724 GNDA 14.0449
R5123 GNDA.n1179 GNDA 14.0449
R5124 GNDA.n1311 GNDA 14.0449
R5125 GNDA.n301 GNDA 14.0449
R5126 GNDA.n1020 GNDA 14.0449
R5127 GNDA.n1936 GNDA 14.0449
R5128 GNDA.n2091 GNDA 14.0449
R5129 GNDA.n2500 GNDA.n2499 14.0193
R5130 GNDA.n2455 GNDA.n2454 13.8005
R5131 GNDA.n2416 GNDA.n2415 13.8005
R5132 GNDA.n2324 GNDA.n2323 13.8005
R5133 GNDA.n2453 GNDA.n2452 13.8005
R5134 GNDA.n2280 GNDA.n2279 13.8005
R5135 GNDA.n906 GNDA.n65 13.7706
R5136 GNDA.n2304 GNDA.n80 13.7449
R5137 GNDA.n1965 GNDA.n351 12.9309
R5138 GNDA.n1498 GNDA.n1467 12.9309
R5139 GNDA.n1760 GNDA.n486 12.9309
R5140 GNDA.n1409 GNDA.n424 12.9309
R5141 GNDA.n2346 GNDA.n2345 12.8005
R5142 GNDA.n2231 GNDA.n2219 12.8005
R5143 GNDA.n1992 GNDA.n221 12.4126
R5144 GNDA.n457 GNDA.n454 12.4126
R5145 GNDA.n524 GNDA.n518 12.4126
R5146 GNDA.n1557 GNDA.n1556 11.6369
R5147 GNDA.n1556 GNDA.n1555 11.6369
R5148 GNDA.n1555 GNDA.n812 11.6369
R5149 GNDA.n1549 GNDA.n812 11.6369
R5150 GNDA.n1549 GNDA.n1548 11.6369
R5151 GNDA.n1548 GNDA.n1547 11.6369
R5152 GNDA.n1547 GNDA.n816 11.6369
R5153 GNDA.n1541 GNDA.n816 11.6369
R5154 GNDA.n1541 GNDA.n1540 11.6369
R5155 GNDA.n1993 GNDA.n1992 11.6369
R5156 GNDA.n1994 GNDA.n1993 11.6369
R5157 GNDA.n1994 GNDA.n217 11.6369
R5158 GNDA.n2000 GNDA.n217 11.6369
R5159 GNDA.n2001 GNDA.n2000 11.6369
R5160 GNDA.n2128 GNDA.n2001 11.6369
R5161 GNDA.n2127 GNDA.n2126 11.6369
R5162 GNDA.n2126 GNDA.n2002 11.6369
R5163 GNDA.n1967 GNDA.n1966 11.6369
R5164 GNDA.n1968 GNDA.n1967 11.6369
R5165 GNDA.n1968 GNDA.n226 11.6369
R5166 GNDA.n1974 GNDA.n226 11.6369
R5167 GNDA.n1975 GNDA.n1974 11.6369
R5168 GNDA.n1976 GNDA.n1975 11.6369
R5169 GNDA.n1976 GNDA.n224 11.6369
R5170 GNDA.n1982 GNDA.n224 11.6369
R5171 GNDA.n1983 GNDA.n1982 11.6369
R5172 GNDA.n1984 GNDA.n1983 11.6369
R5173 GNDA.n1984 GNDA.n222 11.6369
R5174 GNDA.n1214 GNDA.n1212 11.6369
R5175 GNDA.n1212 GNDA.n1209 11.6369
R5176 GNDA.n1209 GNDA.n1208 11.6369
R5177 GNDA.n1208 GNDA.n1205 11.6369
R5178 GNDA.n1205 GNDA.n1204 11.6369
R5179 GNDA.n1204 GNDA.n1201 11.6369
R5180 GNDA.n1201 GNDA.n1200 11.6369
R5181 GNDA.n1200 GNDA.n1197 11.6369
R5182 GNDA.n1197 GNDA.n1196 11.6369
R5183 GNDA.n1196 GNDA.n352 11.6369
R5184 GNDA.n1964 GNDA.n352 11.6369
R5185 GNDA.n1534 GNDA.n1533 11.6369
R5186 GNDA.n1533 GNDA.n1532 11.6369
R5187 GNDA.n1532 GNDA.n1092 11.6369
R5188 GNDA.n1518 GNDA.n1092 11.6369
R5189 GNDA.n1518 GNDA.n1517 11.6369
R5190 GNDA.n1517 GNDA.n1516 11.6369
R5191 GNDA.n1516 GNDA.n1104 11.6369
R5192 GNDA.n1193 GNDA.n1104 11.6369
R5193 GNDA.n1194 GNDA.n1193 11.6369
R5194 GNDA.n1500 GNDA.n1194 11.6369
R5195 GNDA.n1500 GNDA.n1499 11.6369
R5196 GNDA.n1091 GNDA.n1090 11.6369
R5197 GNDA.n1090 GNDA.n831 11.6369
R5198 GNDA.n1084 GNDA.n831 11.6369
R5199 GNDA.n1084 GNDA.n1083 11.6369
R5200 GNDA.n1083 GNDA.n1082 11.6369
R5201 GNDA.n1082 GNDA.n836 11.6369
R5202 GNDA.n1076 GNDA.n836 11.6369
R5203 GNDA.n1076 GNDA.n1075 11.6369
R5204 GNDA.n1075 GNDA.n1074 11.6369
R5205 GNDA.n1408 GNDA.n1348 11.6369
R5206 GNDA.n1349 GNDA.n1348 11.6369
R5207 GNDA.n1401 GNDA.n1349 11.6369
R5208 GNDA.n1401 GNDA.n1400 11.6369
R5209 GNDA.n1400 GNDA.n1399 11.6369
R5210 GNDA.n1399 GNDA.n1351 11.6369
R5211 GNDA.n1394 GNDA.n1351 11.6369
R5212 GNDA.n1394 GNDA.n1393 11.6369
R5213 GNDA.n1393 GNDA.n1392 11.6369
R5214 GNDA.n1392 GNDA.n1354 11.6369
R5215 GNDA.n1387 GNDA.n1354 11.6369
R5216 GNDA.n485 GNDA.n448 11.6369
R5217 GNDA.n480 GNDA.n448 11.6369
R5218 GNDA.n480 GNDA.n479 11.6369
R5219 GNDA.n479 GNDA.n450 11.6369
R5220 GNDA.n474 GNDA.n450 11.6369
R5221 GNDA.n474 GNDA.n473 11.6369
R5222 GNDA.n473 GNDA.n472 11.6369
R5223 GNDA.n472 GNDA.n452 11.6369
R5224 GNDA.n466 GNDA.n452 11.6369
R5225 GNDA.n466 GNDA.n465 11.6369
R5226 GNDA.n465 GNDA.n464 11.6369
R5227 GNDA.n457 GNDA.n456 11.6369
R5228 GNDA.n456 GNDA.n113 11.6369
R5229 GNDA.n2163 GNDA.n113 11.6369
R5230 GNDA.n2163 GNDA.n2162 11.6369
R5231 GNDA.n2162 GNDA.n2161 11.6369
R5232 GNDA.n2161 GNDA.n114 11.6369
R5233 GNDA.n2309 GNDA.n2308 11.6369
R5234 GNDA.n2308 GNDA.n2307 11.6369
R5235 GNDA.n1417 GNDA.n811 11.6369
R5236 GNDA.n1418 GNDA.n1417 11.6369
R5237 GNDA.n1418 GNDA.n1414 11.6369
R5238 GNDA.n1424 GNDA.n1414 11.6369
R5239 GNDA.n1425 GNDA.n1424 11.6369
R5240 GNDA.n1426 GNDA.n1425 11.6369
R5241 GNDA.n1426 GNDA.n1412 11.6369
R5242 GNDA.n1432 GNDA.n1412 11.6369
R5243 GNDA.n1433 GNDA.n1432 11.6369
R5244 GNDA.n1434 GNDA.n1433 11.6369
R5245 GNDA.n1434 GNDA.n1410 11.6369
R5246 GNDA.n677 GNDA.n636 11.6369
R5247 GNDA.n678 GNDA.n677 11.6369
R5248 GNDA.n679 GNDA.n678 11.6369
R5249 GNDA.n679 GNDA.n632 11.6369
R5250 GNDA.n685 GNDA.n632 11.6369
R5251 GNDA.n686 GNDA.n685 11.6369
R5252 GNDA.n687 GNDA.n686 11.6369
R5253 GNDA.n687 GNDA.n627 11.6369
R5254 GNDA.n693 GNDA.n627 11.6369
R5255 GNDA.n671 GNDA.n670 11.6369
R5256 GNDA.n670 GNDA.n669 11.6369
R5257 GNDA.n669 GNDA.n640 11.6369
R5258 GNDA.n663 GNDA.n640 11.6369
R5259 GNDA.n663 GNDA.n662 11.6369
R5260 GNDA.n662 GNDA.n661 11.6369
R5261 GNDA.n661 GNDA.n643 11.6369
R5262 GNDA.n647 GNDA.n643 11.6369
R5263 GNDA.n654 GNDA.n647 11.6369
R5264 GNDA.n654 GNDA.n653 11.6369
R5265 GNDA.n653 GNDA.n652 11.6369
R5266 GNDA.n1593 GNDA.n1592 11.6369
R5267 GNDA.n1594 GNDA.n1593 11.6369
R5268 GNDA.n1594 GNDA.n574 11.6369
R5269 GNDA.n1600 GNDA.n574 11.6369
R5270 GNDA.n1601 GNDA.n1600 11.6369
R5271 GNDA.n1603 GNDA.n565 11.6369
R5272 GNDA.n1609 GNDA.n565 11.6369
R5273 GNDA.n1610 GNDA.n1609 11.6369
R5274 GNDA.n1611 GNDA.n1610 11.6369
R5275 GNDA.n1611 GNDA.n534 11.6369
R5276 GNDA.n1622 GNDA.n1621 11.6369
R5277 GNDA.n1624 GNDA.n1622 11.6369
R5278 GNDA.n1624 GNDA.n1623 11.6369
R5279 GNDA.n1623 GNDA.n530 11.6369
R5280 GNDA.n1631 GNDA.n530 11.6369
R5281 GNDA.n1632 GNDA.n1631 11.6369
R5282 GNDA.n1633 GNDA.n1632 11.6369
R5283 GNDA.n1633 GNDA.n527 11.6369
R5284 GNDA.n1640 GNDA.n527 11.6369
R5285 GNDA.n1641 GNDA.n1640 11.6369
R5286 GNDA.n1642 GNDA.n1641 11.6369
R5287 GNDA.n524 GNDA.n523 11.6369
R5288 GNDA.n523 GNDA.n92 11.6369
R5289 GNDA.n2187 GNDA.n92 11.6369
R5290 GNDA.n2187 GNDA.n2186 11.6369
R5291 GNDA.n2186 GNDA.n2185 11.6369
R5292 GNDA.n2185 GNDA.n93 11.6369
R5293 GNDA.n2179 GNDA.n2178 11.6369
R5294 GNDA.n2178 GNDA.n2177 11.6369
R5295 GNDA.n2278 GNDA.n2277 11.6255
R5296 GNDA GNDA.n2127 11.5076
R5297 GNDA.n2309 GNDA 11.5076
R5298 GNDA.n2179 GNDA 11.5076
R5299 GNDA.n2119 GNDA.n2002 11.4026
R5300 GNDA.n2307 GNDA.n77 11.4026
R5301 GNDA.n2177 GNDA.n100 11.4026
R5302 GNDA.n1540 GNDA.n1539 11.249
R5303 GNDA.n1074 GNDA.n840 11.249
R5304 GNDA.n694 GNDA.n693 11.249
R5305 GNDA.n2460 GNDA.t21 11.2441
R5306 GNDA.t204 GNDA.n41 11.2441
R5307 GNDA.t54 GNDA.n2444 11.2441
R5308 GNDA.n2444 GNDA.t38 11.2441
R5309 GNDA.t337 GNDA.t187 11.2441
R5310 GNDA.n2496 GNDA.t145 11.2441
R5311 GNDA.t120 GNDA.t131 11.2059
R5312 GNDA.t76 GNDA.t245 11.2059
R5313 GNDA.n2425 GNDA.t272 11.2059
R5314 GNDA.t275 GNDA.n2249 11.2059
R5315 GNDA.t345 GNDA.t313 11.2059
R5316 GNDA.t27 GNDA.t135 11.2059
R5317 GNDA.n1605 GNDA.n360 10.6945
R5318 GNDA.n1602 GNDA.n1601 10.4732
R5319 GNDA.n2175 GNDA.n2174 10.1594
R5320 GNDA.n2107 GNDA.n214 10.1594
R5321 GNDA.n2326 GNDA.n61 9.78488
R5322 GNDA.t255 GNDA.n2196 9.6005
R5323 GNDA.n2196 GNDA.t339 9.6005
R5324 GNDA.t320 GNDA.n38 9.6005
R5325 GNDA.n38 GNDA.t91 9.6005
R5326 GNDA.n2395 GNDA.t5 9.6005
R5327 GNDA.n2395 GNDA.t206 9.6005
R5328 GNDA.n2397 GNDA.t343 9.6005
R5329 GNDA.n2397 GNDA.t197 9.6005
R5330 GNDA.n2399 GNDA.t52 9.6005
R5331 GNDA.n2399 GNDA.t67 9.6005
R5332 GNDA.n2401 GNDA.t43 9.6005
R5333 GNDA.n2401 GNDA.t152 9.6005
R5334 GNDA.n2403 GNDA.t202 9.6005
R5335 GNDA.n2403 GNDA.t144 9.6005
R5336 GNDA.n2405 GNDA.t55 9.6005
R5337 GNDA.n2405 GNDA.t351 9.6005
R5338 GNDA.n2407 GNDA.t199 9.6005
R5339 GNDA.n2407 GNDA.t219 9.6005
R5340 GNDA.n2409 GNDA.t41 9.6005
R5341 GNDA.n2409 GNDA.t13 9.6005
R5342 GNDA.n2411 GNDA.t7 9.6005
R5343 GNDA.n2411 GNDA.t208 9.6005
R5344 GNDA.n2413 GNDA.t37 9.6005
R5345 GNDA.n2413 GNDA.t284 9.6005
R5346 GNDA.n2322 GNDA.t229 9.6005
R5347 GNDA.n2322 GNDA.t231 9.6005
R5348 GNDA.n62 GNDA.t227 9.6005
R5349 GNDA.n62 GNDA.t232 9.6005
R5350 GNDA.t33 GNDA.n1656 9.56182
R5351 GNDA.n2324 GNDA.n2321 9.37925
R5352 GNDA.n2473 GNDA.n2472 9.3005
R5353 GNDA.n222 GNDA.n221 8.66313
R5354 GNDA.n464 GNDA.n454 8.66313
R5355 GNDA.n1642 GNDA.n518 8.66313
R5356 GNDA.n1965 GNDA.n1964 8.53383
R5357 GNDA.n1499 GNDA.n1498 8.53383
R5358 GNDA.n1387 GNDA.n486 8.53383
R5359 GNDA.n1410 GNDA.n1409 8.53383
R5360 GNDA.n652 GNDA.n578 8.53383
R5361 GNDA.n1618 GNDA.n534 8.53383
R5362 GNDA.n905 GNDA.n904 8.44175
R5363 GNDA.n1656 GNDA.t29 8.36666
R5364 GNDA.n803 GNDA.n695 8.35606
R5365 GNDA.n1782 GNDA.n425 8.35606
R5366 GNDA.n1678 GNDA.n490 8.35606
R5367 GNDA.n1136 GNDA.n821 8.35606
R5368 GNDA.n1265 GNDA.n1221 8.35606
R5369 GNDA.n347 GNDA.n230 8.35606
R5370 GNDA.n1065 GNDA.n844 8.35606
R5371 GNDA.n1893 GNDA.n395 8.35606
R5372 GNDA.n2044 GNDA.n201 8.35606
R5373 GNDA.n2166 GNDA.n2165 7.76907
R5374 GNDA.n2327 GNDA.n2326 7.71925
R5375 GNDA.n2383 GNDA.t3 7.61296
R5376 GNDA.n2376 GNDA.t32 7.61296
R5377 GNDA.n71 GNDA.n70 6.4005
R5378 GNDA.n934 GNDA.t170 6.32234
R5379 GNDA.t141 GNDA.t304 6.32234
R5380 GNDA.n950 GNDA.t162 6.32234
R5381 GNDA.n2331 GNDA.t94 6.32234
R5382 GNDA.t209 GNDA.t290 6.32234
R5383 GNDA.n914 GNDA.t172 6.32234
R5384 GNDA.n2174 GNDA.t112 5.37874
R5385 GNDA.n2500 GNDA.n1 5.03175
R5386 GNDA.n2277 GNDA.n1 4.90675
R5387 GNDA.n2472 GNDA.n1 4.7505
R5388 GNDA.n1034 GNDA.n1033 4.6085
R5389 GNDA.n1944 GNDA.n175 4.6085
R5390 GNDA.n2118 GNDA.n2006 4.6085
R5391 GNDA.n1217 GNDA.n1215 4.6085
R5392 GNDA.n1249 GNDA.n1245 4.6085
R5393 GNDA.n315 GNDA.n309 4.6085
R5394 GNDA.n1564 GNDA.n1563 4.6085
R5395 GNDA.n1766 GNDA.n1762 4.6085
R5396 GNDA.n1662 GNDA.n512 4.6085
R5397 GNDA.n2155 GNDA.n150 4.55161
R5398 GNDA.n1497 GNDA.n1494 4.55161
R5399 GNDA.n1384 GNDA.n1356 4.55161
R5400 GNDA.n1440 GNDA.n1347 4.55161
R5401 GNDA.n1588 GNDA.n579 4.55161
R5402 GNDA.n1617 GNDA.n560 4.55161
R5403 GNDA.n1029 GNDA.n403 4.5061
R5404 GNDA.n2149 GNDA.n2148 4.5061
R5405 GNDA.n1467 GNDA.n1219 4.5061
R5406 GNDA.n1244 GNDA.n351 4.5061
R5407 GNDA.n1565 GNDA.n424 4.5061
R5408 GNDA.n1761 GNDA.n1760 4.5061
R5409 GNDA.n2471 GNDA.n2469 4.5005
R5410 GNDA.n2326 GNDA.n2325 4.5005
R5411 GNDA.n2417 GNDA.n0 4.5005
R5412 GNDA.n2513 GNDA.n2512 4.5005
R5413 GNDA.n1966 GNDA.n1965 4.39646
R5414 GNDA.n1498 GNDA.n1214 4.39646
R5415 GNDA.n1409 GNDA.n1408 4.39646
R5416 GNDA.n486 GNDA.n485 4.39646
R5417 GNDA.n1592 GNDA.n578 4.39646
R5418 GNDA.n1621 GNDA.n1618 4.39646
R5419 GNDA.n1869 GNDA.n403 4.3525
R5420 GNDA.n2148 GNDA.n2147 4.3525
R5421 GNDA.n1467 GNDA.n1346 4.3525
R5422 GNDA.n351 GNDA.n350 4.3525
R5423 GNDA.n1863 GNDA.n424 4.3525
R5424 GNDA.n1760 GNDA.n1759 4.3525
R5425 GNDA.n1870 GNDA.n1869 4.3013
R5426 GNDA.n2147 GNDA.n2146 4.3013
R5427 GNDA.n1346 GNDA.n1345 4.3013
R5428 GNDA.n350 GNDA.n349 4.3013
R5429 GNDA.n1863 GNDA.n1862 4.3013
R5430 GNDA.n1759 GNDA.n1758 4.3013
R5431 GNDA.n2155 GNDA.n151 4.26717
R5432 GNDA.n177 GNDA.n151 4.26717
R5433 GNDA.n180 GNDA.n177 4.26717
R5434 GNDA.n183 GNDA.n180 4.26717
R5435 GNDA.n186 GNDA.n183 4.26717
R5436 GNDA.n189 GNDA.n186 4.26717
R5437 GNDA.n195 GNDA.n192 4.26717
R5438 GNDA.n199 GNDA.n195 4.26717
R5439 GNDA.n1494 GNDA.n1493 4.26717
R5440 GNDA.n1493 GNDA.n1490 4.26717
R5441 GNDA.n1490 GNDA.n1489 4.26717
R5442 GNDA.n1489 GNDA.n1486 4.26717
R5443 GNDA.n1486 GNDA.n1485 4.26717
R5444 GNDA.n1485 GNDA.n1482 4.26717
R5445 GNDA.n1481 GNDA.n1478 4.26717
R5446 GNDA.n1478 GNDA.n1477 4.26717
R5447 GNDA.n1384 GNDA.n1383 4.26717
R5448 GNDA.n1383 GNDA.n1380 4.26717
R5449 GNDA.n1380 GNDA.n1379 4.26717
R5450 GNDA.n1379 GNDA.n1376 4.26717
R5451 GNDA.n1376 GNDA.n1375 4.26717
R5452 GNDA.n1375 GNDA.n1372 4.26717
R5453 GNDA.n1371 GNDA.n1368 4.26717
R5454 GNDA.n1368 GNDA.n1367 4.26717
R5455 GNDA.n1442 GNDA.n1440 4.26717
R5456 GNDA.n1445 GNDA.n1442 4.26717
R5457 GNDA.n1448 GNDA.n1445 4.26717
R5458 GNDA.n1451 GNDA.n1448 4.26717
R5459 GNDA.n1454 GNDA.n1451 4.26717
R5460 GNDA.n1457 GNDA.n1454 4.26717
R5461 GNDA.n1462 GNDA.n1461 4.26717
R5462 GNDA.n1466 GNDA.n1462 4.26717
R5463 GNDA.n1588 GNDA.n1587 4.26717
R5464 GNDA.n1587 GNDA.n1584 4.26717
R5465 GNDA.n1584 GNDA.n1583 4.26717
R5466 GNDA.n1583 GNDA.n1580 4.26717
R5467 GNDA.n1580 GNDA.n1579 4.26717
R5468 GNDA.n1579 GNDA.n1576 4.26717
R5469 GNDA.n1575 GNDA.n1572 4.26717
R5470 GNDA.n1572 GNDA.n1571 4.26717
R5471 GNDA.n560 GNDA.n559 4.26717
R5472 GNDA.n559 GNDA.n556 4.26717
R5473 GNDA.n556 GNDA.n555 4.26717
R5474 GNDA.n555 GNDA.n552 4.26717
R5475 GNDA.n552 GNDA.n551 4.26717
R5476 GNDA.n551 GNDA.n548 4.26717
R5477 GNDA.n547 GNDA.n544 4.26717
R5478 GNDA.n544 GNDA.n488 4.26717
R5479 GNDA.n1539 GNDA.n1538 4.2501
R5480 GNDA.n804 GNDA.n694 4.2501
R5481 GNDA.n192 GNDA 4.21976
R5482 GNDA GNDA.n1481 4.21976
R5483 GNDA GNDA.n1371 4.21976
R5484 GNDA.n1461 GNDA 4.21976
R5485 GNDA GNDA.n1575 4.21976
R5486 GNDA GNDA.n547 4.21976
R5487 GNDA.t29 GNDA.t112 4.18358
R5488 GNDA.n1066 GNDA.n840 4.1477
R5489 GNDA.n2148 GNDA.n199 4.12494
R5490 GNDA.n1477 GNDA.n403 4.12494
R5491 GNDA.n1367 GNDA.n351 4.12494
R5492 GNDA.n1467 GNDA.n1466 4.12494
R5493 GNDA.n1571 GNDA.n424 4.12494
R5494 GNDA.n1760 GNDA.n488 4.12494
R5495 GNDA.n2325 GNDA.n2324 3.813
R5496 GNDA.t254 GNDA.n2195 3.74837
R5497 GNDA.n2193 GNDA.t338 3.74837
R5498 GNDA.t146 GNDA.n2459 3.74837
R5499 GNDA.n42 GNDA.t220 3.74837
R5500 GNDA.n41 GNDA.t50 3.74837
R5501 GNDA.n2476 GNDA.t310 3.74837
R5502 GNDA.n2448 GNDA.t45 3.74837
R5503 GNDA.n2441 GNDA.t0 3.74837
R5504 GNDA.t0 GNDA.t337 3.74837
R5505 GNDA.t260 GNDA.t257 3.73564
R5506 GNDA.n2241 GNDA.t116 3.73564
R5507 GNDA.n2240 GNDA.t103 3.73564
R5508 GNDA.t280 GNDA.t301 3.73564
R5509 GNDA.n2321 GNDA 3.68412
R5510 GNDA.n2512 GNDA.n2500 3.6255
R5511 GNDA.n2107 GNDA.t70 3.586
R5512 GNDA.n1064 GNDA.n1063 3.5845
R5513 GNDA.n847 GNDA.n845 3.5845
R5514 GNDA.n1058 GNDA.n849 3.5845
R5515 GNDA.n1057 GNDA.n850 3.5845
R5516 GNDA.n1049 GNDA.n1048 3.5845
R5517 GNDA.n855 GNDA.n853 3.5845
R5518 GNDA.n1043 GNDA.n857 3.5845
R5519 GNDA.n1042 GNDA.n858 3.5845
R5520 GNDA.n960 GNDA.n959 3.5845
R5521 GNDA.n1889 GNDA.n397 3.5845
R5522 GNDA.n1888 GNDA.n398 3.5845
R5523 GNDA.n1875 GNDA.n1874 3.5845
R5524 GNDA.n1882 GNDA.n1881 3.5845
R5525 GNDA.n1876 GNDA.n368 3.5845
R5526 GNDA.n1958 GNDA.n1957 3.5845
R5527 GNDA.n1953 GNDA.n369 3.5845
R5528 GNDA.n1952 GNDA.n372 3.5845
R5529 GNDA.n378 GNDA.n377 3.5845
R5530 GNDA.n206 GNDA.n205 3.5845
R5531 GNDA.n2140 GNDA.n2139 3.5845
R5532 GNDA.n2135 GNDA.n207 3.5845
R5533 GNDA.n2134 GNDA.n210 3.5845
R5534 GNDA.n2018 GNDA.n2014 3.5845
R5535 GNDA.n2019 GNDA.n2013 3.5845
R5536 GNDA.n2025 GNDA.n2023 3.5845
R5537 GNDA.n2024 GNDA.n2010 3.5845
R5538 GNDA.n2099 GNDA.n2098 3.5845
R5539 GNDA.n1097 GNDA.n1096 3.5845
R5540 GNDA.n1528 GNDA.n1527 3.5845
R5541 GNDA.n1523 GNDA.n1098 3.5845
R5542 GNDA.n1522 GNDA.n1101 3.5845
R5543 GNDA.n1114 GNDA.n1112 3.5845
R5544 GNDA.n1113 GNDA.n1109 3.5845
R5545 GNDA.n1511 GNDA.n1510 3.5845
R5546 GNDA.n1118 GNDA.n1110 3.5845
R5547 GNDA.n1505 GNDA.n1120 3.5845
R5548 GNDA.n1341 GNDA.n1340 3.5845
R5549 GNDA.n1225 GNDA.n1223 3.5845
R5550 GNDA.n1335 GNDA.n1227 3.5845
R5551 GNDA.n1334 GNDA.n1228 3.5845
R5552 GNDA.n1330 GNDA.n1329 3.5845
R5553 GNDA.n1234 GNDA.n1232 3.5845
R5554 GNDA.n1324 GNDA.n1236 3.5845
R5555 GNDA.n1323 GNDA.n1237 3.5845
R5556 GNDA.n1319 GNDA.n1318 3.5845
R5557 GNDA.n346 GNDA.n231 3.5845
R5558 GNDA.n343 GNDA.n342 3.5845
R5559 GNDA.n338 GNDA.n232 3.5845
R5560 GNDA.n337 GNDA.n334 3.5845
R5561 GNDA.n333 GNDA.n235 3.5845
R5562 GNDA.n330 GNDA.n329 3.5845
R5563 GNDA.n325 GNDA.n236 3.5845
R5564 GNDA.n324 GNDA.n321 3.5845
R5565 GNDA.n320 GNDA.n240 3.5845
R5566 GNDA.n802 GNDA.n696 3.5845
R5567 GNDA.n799 GNDA.n798 3.5845
R5568 GNDA.n794 GNDA.n697 3.5845
R5569 GNDA.n793 GNDA.n790 3.5845
R5570 GNDA.n789 GNDA.n700 3.5845
R5571 GNDA.n786 GNDA.n785 3.5845
R5572 GNDA.n781 GNDA.n701 3.5845
R5573 GNDA.n780 GNDA.n777 3.5845
R5574 GNDA.n776 GNDA.n774 3.5845
R5575 GNDA.n1858 GNDA.n1857 3.5845
R5576 GNDA.n429 GNDA.n427 3.5845
R5577 GNDA.n1852 GNDA.n431 3.5845
R5578 GNDA.n1851 GNDA.n432 3.5845
R5579 GNDA.n1847 GNDA.n1846 3.5845
R5580 GNDA.n438 GNDA.n436 3.5845
R5581 GNDA.n1841 GNDA.n440 3.5845
R5582 GNDA.n1840 GNDA.n441 3.5845
R5583 GNDA.n1836 GNDA.n1835 3.5845
R5584 GNDA.n1754 GNDA.n1753 3.5845
R5585 GNDA.n494 GNDA.n492 3.5845
R5586 GNDA.n1748 GNDA.n496 3.5845
R5587 GNDA.n1747 GNDA.n497 3.5845
R5588 GNDA.n1743 GNDA.n1742 3.5845
R5589 GNDA.n503 GNDA.n501 3.5845
R5590 GNDA.n1737 GNDA.n505 3.5845
R5591 GNDA.n1736 GNDA.n506 3.5845
R5592 GNDA.n1732 GNDA.n1731 3.5845
R5593 GNDA.n2264 GNDA.t109 3.42907
R5594 GNDA.n2264 GNDA.t28 3.42907
R5595 GNDA.n2418 GNDA.t132 3.42907
R5596 GNDA.n2418 GNDA.t190 3.42907
R5597 GNDA.n2420 GNDA.t341 3.42907
R5598 GNDA.n2420 GNDA.t18 3.42907
R5599 GNDA.n2197 GNDA.t193 3.42907
R5600 GNDA.n2197 GNDA.t137 3.42907
R5601 GNDA.n1066 GNDA.n1065 3.3797
R5602 GNDA.n1870 GNDA.n395 3.3797
R5603 GNDA.n2146 GNDA.n201 3.3797
R5604 GNDA.n1538 GNDA.n821 3.3797
R5605 GNDA.n1345 GNDA.n1221 3.3797
R5606 GNDA.n349 GNDA.n347 3.3797
R5607 GNDA.n804 GNDA.n803 3.3797
R5608 GNDA.n1862 GNDA.n425 3.3797
R5609 GNDA.n1758 GNDA.n490 3.3797
R5610 GNDA.n2302 GNDA.n69 3.2005
R5611 GNDA.n1654 GNDA.n1650 3.2005
R5612 GNDA.n1036 GNDA.n1035 2.8677
R5613 GNDA.n1946 GNDA.n1945 2.8677
R5614 GNDA.n2029 GNDA.n2011 2.8677
R5615 GNDA.n1504 GNDA.n1187 2.8677
R5616 GNDA.n1250 GNDA.n1241 2.8677
R5617 GNDA.n317 GNDA.n316 2.8677
R5618 GNDA.n705 GNDA.n610 2.8677
R5619 GNDA.n1767 GNDA.n445 2.8677
R5620 GNDA.n1663 GNDA.n510 2.8677
R5621 GNDA.n2373 GNDA.t3 2.53799
R5622 GNDA.t2 GNDA.n2374 2.53799
R5623 GNDA.n2513 GNDA.n0 2.5005
R5624 GNDA.n892 GNDA.n890 2.34425
R5625 GNDA.n900 GNDA.n898 2.34425
R5626 GNDA.n707 GNDA.n610 2.31161
R5627 GNDA.n1768 GNDA.n1767 2.31161
R5628 GNDA.n1664 GNDA.n1663 2.31161
R5629 GNDA.n1187 GNDA.n1186 2.31161
R5630 GNDA.n1251 GNDA.n1250 2.31161
R5631 GNDA.n316 GNDA.n308 2.31161
R5632 GNDA.n1035 GNDA.n1027 2.31161
R5633 GNDA.n1945 GNDA.n1943 2.31161
R5634 GNDA.n2030 GNDA.n2029 2.31161
R5635 GNDA.n2419 GNDA.n2417 2.063
R5636 GNDA.n709 GNDA 1.95606
R5637 GNDA.n1770 GNDA 1.95606
R5638 GNDA.n1666 GNDA 1.95606
R5639 GNDA GNDA.n1178 1.95606
R5640 GNDA.n1253 GNDA 1.95606
R5641 GNDA GNDA.n300 1.95606
R5642 GNDA GNDA.n1019 1.95606
R5643 GNDA GNDA.n1935 1.95606
R5644 GNDA.n2032 GNDA 1.95606
R5645 GNDA.n2278 GNDA.n2265 1.813
R5646 GNDA.n2312 GNDA.n2311 1.79325
R5647 GNDA.n2417 GNDA.n2416 1.78175
R5648 GNDA.n2279 GNDA.n2278 1.78175
R5649 GNDA.n1035 GNDA.n1034 1.7413
R5650 GNDA.n1945 GNDA.n1944 1.7413
R5651 GNDA.n2029 GNDA.n2006 1.7413
R5652 GNDA.n1215 GNDA.n1187 1.7413
R5653 GNDA.n1250 GNDA.n1249 1.7413
R5654 GNDA.n316 GNDA.n315 1.7413
R5655 GNDA.n1563 GNDA.n610 1.7413
R5656 GNDA.n1767 GNDA.n1766 1.7413
R5657 GNDA.n1663 GNDA.n1662 1.7413
R5658 GNDA.n2316 GNDA.n65 1.73362
R5659 GNDA.n2499 GNDA.n2 1.6005
R5660 GNDA.n2227 GNDA.t124 1.58323
R5661 GNDA.n1065 GNDA.n1064 1.2293
R5662 GNDA.n397 GNDA.n395 1.2293
R5663 GNDA.n205 GNDA.n201 1.2293
R5664 GNDA.n1096 GNDA.n821 1.2293
R5665 GNDA.n1341 GNDA.n1221 1.2293
R5666 GNDA.n347 GNDA.n346 1.2293
R5667 GNDA.n803 GNDA.n802 1.2293
R5668 GNDA.n1858 GNDA.n425 1.2293
R5669 GNDA.n1754 GNDA.n490 1.2293
R5670 GNDA.n2454 GNDA.n2453 1.21925
R5671 GNDA.n1033 GNDA.n1029 1.1781
R5672 GNDA.n2149 GNDA.n175 1.1781
R5673 GNDA.n2119 GNDA.n2118 1.1781
R5674 GNDA.n1219 GNDA.n1217 1.1781
R5675 GNDA.n1245 GNDA.n1244 1.1781
R5676 GNDA.n309 GNDA.n77 1.1781
R5677 GNDA.n1565 GNDA.n1564 1.1781
R5678 GNDA.n1762 GNDA.n1761 1.1781
R5679 GNDA.n512 GNDA.n100 1.1781
R5680 GNDA.n1603 GNDA.n1602 1.16414
R5681 GNDA.n1063 GNDA.n845 1.0245
R5682 GNDA.n849 GNDA.n847 1.0245
R5683 GNDA.n1058 GNDA.n1057 1.0245
R5684 GNDA.n1049 GNDA.n850 1.0245
R5685 GNDA.n1048 GNDA.n853 1.0245
R5686 GNDA.n857 GNDA.n855 1.0245
R5687 GNDA.n1043 GNDA.n1042 1.0245
R5688 GNDA.n959 GNDA.n858 1.0245
R5689 GNDA.n1036 GNDA.n960 1.0245
R5690 GNDA.n1889 GNDA.n1888 1.0245
R5691 GNDA.n1874 GNDA.n398 1.0245
R5692 GNDA.n1882 GNDA.n1875 1.0245
R5693 GNDA.n1881 GNDA.n1876 1.0245
R5694 GNDA.n1958 GNDA.n368 1.0245
R5695 GNDA.n1957 GNDA.n369 1.0245
R5696 GNDA.n1953 GNDA.n1952 1.0245
R5697 GNDA.n377 GNDA.n372 1.0245
R5698 GNDA.n1946 GNDA.n378 1.0245
R5699 GNDA.n2140 GNDA.n206 1.0245
R5700 GNDA.n2139 GNDA.n207 1.0245
R5701 GNDA.n2135 GNDA.n2134 1.0245
R5702 GNDA.n2014 GNDA.n210 1.0245
R5703 GNDA.n2019 GNDA.n2018 1.0245
R5704 GNDA.n2023 GNDA.n2013 1.0245
R5705 GNDA.n2025 GNDA.n2024 1.0245
R5706 GNDA.n2099 GNDA.n2010 1.0245
R5707 GNDA.n2098 GNDA.n2011 1.0245
R5708 GNDA.n1528 GNDA.n1097 1.0245
R5709 GNDA.n1527 GNDA.n1098 1.0245
R5710 GNDA.n1523 GNDA.n1522 1.0245
R5711 GNDA.n1112 GNDA.n1101 1.0245
R5712 GNDA.n1114 GNDA.n1113 1.0245
R5713 GNDA.n1511 GNDA.n1109 1.0245
R5714 GNDA.n1510 GNDA.n1110 1.0245
R5715 GNDA.n1120 GNDA.n1118 1.0245
R5716 GNDA.n1505 GNDA.n1504 1.0245
R5717 GNDA.n1340 GNDA.n1223 1.0245
R5718 GNDA.n1227 GNDA.n1225 1.0245
R5719 GNDA.n1335 GNDA.n1334 1.0245
R5720 GNDA.n1330 GNDA.n1228 1.0245
R5721 GNDA.n1329 GNDA.n1232 1.0245
R5722 GNDA.n1236 GNDA.n1234 1.0245
R5723 GNDA.n1324 GNDA.n1323 1.0245
R5724 GNDA.n1319 GNDA.n1237 1.0245
R5725 GNDA.n1318 GNDA.n1241 1.0245
R5726 GNDA.n343 GNDA.n231 1.0245
R5727 GNDA.n342 GNDA.n232 1.0245
R5728 GNDA.n338 GNDA.n337 1.0245
R5729 GNDA.n334 GNDA.n333 1.0245
R5730 GNDA.n330 GNDA.n235 1.0245
R5731 GNDA.n329 GNDA.n236 1.0245
R5732 GNDA.n325 GNDA.n324 1.0245
R5733 GNDA.n321 GNDA.n320 1.0245
R5734 GNDA.n317 GNDA.n240 1.0245
R5735 GNDA.n799 GNDA.n696 1.0245
R5736 GNDA.n798 GNDA.n697 1.0245
R5737 GNDA.n794 GNDA.n793 1.0245
R5738 GNDA.n790 GNDA.n789 1.0245
R5739 GNDA.n786 GNDA.n700 1.0245
R5740 GNDA.n785 GNDA.n701 1.0245
R5741 GNDA.n781 GNDA.n780 1.0245
R5742 GNDA.n777 GNDA.n776 1.0245
R5743 GNDA.n774 GNDA.n705 1.0245
R5744 GNDA.n1857 GNDA.n427 1.0245
R5745 GNDA.n431 GNDA.n429 1.0245
R5746 GNDA.n1852 GNDA.n1851 1.0245
R5747 GNDA.n1847 GNDA.n432 1.0245
R5748 GNDA.n1846 GNDA.n436 1.0245
R5749 GNDA.n440 GNDA.n438 1.0245
R5750 GNDA.n1841 GNDA.n1840 1.0245
R5751 GNDA.n1836 GNDA.n441 1.0245
R5752 GNDA.n1835 GNDA.n445 1.0245
R5753 GNDA.n1753 GNDA.n492 1.0245
R5754 GNDA.n496 GNDA.n494 1.0245
R5755 GNDA.n1748 GNDA.n1747 1.0245
R5756 GNDA.n1743 GNDA.n497 1.0245
R5757 GNDA.n1742 GNDA.n501 1.0245
R5758 GNDA.n505 GNDA.n503 1.0245
R5759 GNDA.n1737 GNDA.n1736 1.0245
R5760 GNDA.n1732 GNDA.n506 1.0245
R5761 GNDA.n1731 GNDA.n510 1.0245
R5762 GNDA.n2454 GNDA.n36 0.6255
R5763 GNDA.n2469 GNDA.n2468 0.563
R5764 GNDA.n2469 GNDA.n2465 0.563
R5765 GNDA.n2505 GNDA.n2503 0.563
R5766 GNDA.n2507 GNDA.n2505 0.563
R5767 GNDA.n2509 GNDA.n2507 0.563
R5768 GNDA.n2511 GNDA.n2509 0.563
R5769 GNDA.n2270 GNDA.n2268 0.563
R5770 GNDA.n2272 GNDA.n2270 0.563
R5771 GNDA.n2274 GNDA.n2272 0.563
R5772 GNDA.n2276 GNDA.n2274 0.563
R5773 GNDA.n890 GNDA.n888 0.563
R5774 GNDA.n894 GNDA.n892 0.563
R5775 GNDA.n896 GNDA.n894 0.563
R5776 GNDA.n898 GNDA.n896 0.563
R5777 GNDA.n902 GNDA.n900 0.563
R5778 GNDA.n904 GNDA.n902 0.563
R5779 GNDA.n2414 GNDA.n2412 0.563
R5780 GNDA.n2412 GNDA.n2410 0.563
R5781 GNDA.n2410 GNDA.n2408 0.563
R5782 GNDA.n2408 GNDA.n2406 0.563
R5783 GNDA.n2406 GNDA.n2404 0.563
R5784 GNDA.n2404 GNDA.n2402 0.563
R5785 GNDA.n2402 GNDA.n2400 0.563
R5786 GNDA.n2400 GNDA.n2398 0.563
R5787 GNDA.n2398 GNDA.n2396 0.563
R5788 GNDA.n2396 GNDA.n37 0.563
R5789 GNDA.n2378 GNDA.t111 0.507997
R5790 GNDA.n2421 GNDA.n2419 0.5005
R5791 GNDA.n2265 GNDA.n2263 0.5005
R5792 GNDA.n2320 GNDA.n2318 0.41175
R5793 GNDA.n2318 GNDA.n2317 0.311875
R5794 GNDA.n2416 GNDA.n2414 0.28175
R5795 GNDA.n2321 GNDA.n64 0.276625
R5796 GNDA.n2472 GNDA.n2471 0.2505
R5797 GNDA.n2453 GNDA.n37 0.2505
R5798 GNDA.n2279 GNDA.n36 0.2505
R5799 GNDA.n905 GNDA.n64 0.22375
R5800 GNDA.n2128 GNDA 0.129793
R5801 GNDA.n114 GNDA 0.129793
R5802 GNDA GNDA.n93 0.129793
R5803 GNDA.n906 GNDA.n905 0.100375
R5804 GNDA.n2317 GNDA.n2316 0.076875
R5805 GNDA.n1965 GNDA.n150 0.0479074
R5806 GNDA.n189 GNDA 0.0479074
R5807 GNDA.n1498 GNDA.n1497 0.0479074
R5808 GNDA.n1482 GNDA 0.0479074
R5809 GNDA.n1356 GNDA.n486 0.0479074
R5810 GNDA.n1372 GNDA 0.0479074
R5811 GNDA.n1409 GNDA.n1347 0.0479074
R5812 GNDA.n1457 GNDA 0.0479074
R5813 GNDA.n579 GNDA.n578 0.0479074
R5814 GNDA.n1576 GNDA 0.0479074
R5815 GNDA.n1618 GNDA.n1617 0.0479074
R5816 GNDA.n548 GNDA 0.0479074
R5817 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n9 114.719
R5818 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.n6 114.719
R5819 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n10 114.156
R5820 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.n7 114.156
R5821 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.n0 112.456
R5822 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.n18 112.454
R5823 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n17 111.206
R5824 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.n3 111.206
R5825 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.n1 111.206
R5826 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n5 109.656
R5827 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.n14 106.706
R5828 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.t11 16.0005
R5829 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.t6 16.0005
R5830 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t20 16.0005
R5831 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t14 16.0005
R5832 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.t0 16.0005
R5833 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.t9 16.0005
R5834 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.t13 16.0005
R5835 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.t10 16.0005
R5836 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.t5 16.0005
R5837 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.t16 16.0005
R5838 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t21 16.0005
R5839 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t4 16.0005
R5840 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t2 16.0005
R5841 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t12 16.0005
R5842 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t3 16.0005
R5843 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t18 16.0005
R5844 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t17 16.0005
R5845 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t8 16.0005
R5846 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.t1 16.0005
R5847 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.t7 16.0005
R5848 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.t15 16.0005
R5849 two_stage_opamp_dummy_magic_0.VD2.t19 two_stage_opamp_dummy_magic_0.VD2.n19 16.0005
R5850 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n12 4.5005
R5851 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n15 4.5005
R5852 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n4 3.6255
R5853 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.n2 1.2505
R5854 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n16 1.2505
R5855 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.n13 0.78175
R5856 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.n11 0.563
R5857 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.n8 0.563
R5858 VOUT-.n14 VOUT-.n6 145.989
R5859 VOUT-.n9 VOUT-.n7 145.989
R5860 VOUT-.n13 VOUT-.n12 145.427
R5861 VOUT-.n11 VOUT-.n10 145.427
R5862 VOUT-.n9 VOUT-.n8 145.427
R5863 VOUT-.n16 VOUT-.n15 140.927
R5864 VOUT-.n5 VOUT-.t12 113.192
R5865 VOUT-.n2 VOUT-.n0 95.7303
R5866 VOUT-.n4 VOUT-.n3 94.6053
R5867 VOUT-.n2 VOUT-.n1 94.6053
R5868 VOUT-.n100 VOUT-.n16 20.5943
R5869 VOUT-.n100 VOUT-.n99 11.7059
R5870 VOUT- VOUT-.n100 7.813
R5871 VOUT-.n15 VOUT-.t8 6.56717
R5872 VOUT-.n15 VOUT-.t4 6.56717
R5873 VOUT-.n12 VOUT-.t6 6.56717
R5874 VOUT-.n12 VOUT-.t3 6.56717
R5875 VOUT-.n10 VOUT-.t1 6.56717
R5876 VOUT-.n10 VOUT-.t7 6.56717
R5877 VOUT-.n8 VOUT-.t5 6.56717
R5878 VOUT-.n8 VOUT-.t10 6.56717
R5879 VOUT-.n7 VOUT-.t2 6.56717
R5880 VOUT-.n7 VOUT-.t15 6.56717
R5881 VOUT-.n6 VOUT-.t14 6.56717
R5882 VOUT-.n6 VOUT-.t11 6.56717
R5883 VOUT-.n46 VOUT-.t83 4.8295
R5884 VOUT-.n48 VOUT-.t90 4.8295
R5885 VOUT-.n51 VOUT-.t128 4.8295
R5886 VOUT-.n54 VOUT-.t26 4.8295
R5887 VOUT-.n57 VOUT-.t74 4.8295
R5888 VOUT-.n70 VOUT-.t39 4.8295
R5889 VOUT-.n72 VOUT-.t34 4.8295
R5890 VOUT-.n73 VOUT-.t136 4.8295
R5891 VOUT-.n75 VOUT-.t68 4.8295
R5892 VOUT-.n76 VOUT-.t36 4.8295
R5893 VOUT-.n78 VOUT-.t94 4.8295
R5894 VOUT-.n79 VOUT-.t64 4.8295
R5895 VOUT-.n81 VOUT-.t54 4.8295
R5896 VOUT-.n82 VOUT-.t29 4.8295
R5897 VOUT-.n84 VOUT-.t89 4.8295
R5898 VOUT-.n85 VOUT-.t57 4.8295
R5899 VOUT-.n87 VOUT-.t48 4.8295
R5900 VOUT-.n88 VOUT-.t20 4.8295
R5901 VOUT-.n90 VOUT-.t148 4.8295
R5902 VOUT-.n91 VOUT-.t121 4.8295
R5903 VOUT-.n93 VOUT-.t43 4.8295
R5904 VOUT-.n94 VOUT-.t152 4.8295
R5905 VOUT-.n17 VOUT-.t107 4.8295
R5906 VOUT-.n29 VOUT-.t28 4.8295
R5907 VOUT-.n31 VOUT-.t24 4.8295
R5908 VOUT-.n32 VOUT-.t129 4.8295
R5909 VOUT-.n34 VOUT-.t59 4.8295
R5910 VOUT-.n35 VOUT-.t32 4.8295
R5911 VOUT-.n37 VOUT-.t99 4.8295
R5912 VOUT-.n38 VOUT-.t69 4.8295
R5913 VOUT-.n40 VOUT-.t67 4.8295
R5914 VOUT-.n41 VOUT-.t35 4.8295
R5915 VOUT-.n43 VOUT-.t104 4.8295
R5916 VOUT-.n44 VOUT-.t76 4.8295
R5917 VOUT-.n96 VOUT-.t115 4.8295
R5918 VOUT-.n69 VOUT-.t132 4.806
R5919 VOUT-.n68 VOUT-.t114 4.806
R5920 VOUT-.n67 VOUT-.t146 4.806
R5921 VOUT-.n66 VOUT-.t45 4.806
R5922 VOUT-.n65 VOUT-.t85 4.806
R5923 VOUT-.n64 VOUT-.t63 4.806
R5924 VOUT-.n63 VOUT-.t101 4.806
R5925 VOUT-.n62 VOUT-.t134 4.806
R5926 VOUT-.n61 VOUT-.t119 4.806
R5927 VOUT-.n60 VOUT-.t155 4.806
R5928 VOUT-.n28 VOUT-.t47 4.806
R5929 VOUT-.n27 VOUT-.t91 4.806
R5930 VOUT-.n26 VOUT-.t41 4.806
R5931 VOUT-.n25 VOUT-.t130 4.806
R5932 VOUT-.n24 VOUT-.t82 4.806
R5933 VOUT-.n23 VOUT-.t124 4.806
R5934 VOUT-.n22 VOUT-.t72 4.806
R5935 VOUT-.n21 VOUT-.t23 4.806
R5936 VOUT-.n20 VOUT-.t62 4.806
R5937 VOUT-.n19 VOUT-.t150 4.806
R5938 VOUT-.n47 VOUT-.t95 4.5005
R5939 VOUT-.n46 VOUT-.t56 4.5005
R5940 VOUT-.n48 VOUT-.t131 4.5005
R5941 VOUT-.n49 VOUT-.t103 4.5005
R5942 VOUT-.n50 VOUT-.t71 4.5005
R5943 VOUT-.n51 VOUT-.t31 4.5005
R5944 VOUT-.n52 VOUT-.t138 4.5005
R5945 VOUT-.n53 VOUT-.t106 4.5005
R5946 VOUT-.n54 VOUT-.t60 4.5005
R5947 VOUT-.n55 VOUT-.t40 4.5005
R5948 VOUT-.n56 VOUT-.t143 4.5005
R5949 VOUT-.n57 VOUT-.t113 4.5005
R5950 VOUT-.n58 VOUT-.t21 4.5005
R5951 VOUT-.n59 VOUT-.t125 4.5005
R5952 VOUT-.n60 VOUT-.t118 4.5005
R5953 VOUT-.n61 VOUT-.t80 4.5005
R5954 VOUT-.n62 VOUT-.t96 4.5005
R5955 VOUT-.n63 VOUT-.t61 4.5005
R5956 VOUT-.n64 VOUT-.t27 4.5005
R5957 VOUT-.n65 VOUT-.t44 4.5005
R5958 VOUT-.n66 VOUT-.t144 4.5005
R5959 VOUT-.n67 VOUT-.t111 4.5005
R5960 VOUT-.n68 VOUT-.t75 4.5005
R5961 VOUT-.n69 VOUT-.t92 4.5005
R5962 VOUT-.n71 VOUT-.t55 4.5005
R5963 VOUT-.n70 VOUT-.t19 4.5005
R5964 VOUT-.n72 VOUT-.t51 4.5005
R5965 VOUT-.n74 VOUT-.t156 4.5005
R5966 VOUT-.n73 VOUT-.t120 4.5005
R5967 VOUT-.n75 VOUT-.t87 4.5005
R5968 VOUT-.n77 VOUT-.t49 4.5005
R5969 VOUT-.n76 VOUT-.t151 4.5005
R5970 VOUT-.n78 VOUT-.t42 4.5005
R5971 VOUT-.n80 VOUT-.t145 4.5005
R5972 VOUT-.n79 VOUT-.t117 4.5005
R5973 VOUT-.n81 VOUT-.t141 4.5005
R5974 VOUT-.n83 VOUT-.t110 4.5005
R5975 VOUT-.n82 VOUT-.t79 4.5005
R5976 VOUT-.n84 VOUT-.t38 4.5005
R5977 VOUT-.n86 VOUT-.t139 4.5005
R5978 VOUT-.n85 VOUT-.t108 4.5005
R5979 VOUT-.n87 VOUT-.t135 4.5005
R5980 VOUT-.n89 VOUT-.t102 4.5005
R5981 VOUT-.n88 VOUT-.t70 4.5005
R5982 VOUT-.n90 VOUT-.t98 4.5005
R5983 VOUT-.n92 VOUT-.t66 4.5005
R5984 VOUT-.n91 VOUT-.t33 4.5005
R5985 VOUT-.n93 VOUT-.t133 4.5005
R5986 VOUT-.n95 VOUT-.t97 4.5005
R5987 VOUT-.n94 VOUT-.t65 4.5005
R5988 VOUT-.n18 VOUT-.t100 4.5005
R5989 VOUT-.n17 VOUT-.t149 4.5005
R5990 VOUT-.n19 VOUT-.t86 4.5005
R5991 VOUT-.n20 VOUT-.t50 4.5005
R5992 VOUT-.n21 VOUT-.t137 4.5005
R5993 VOUT-.n22 VOUT-.t105 4.5005
R5994 VOUT-.n23 VOUT-.t73 4.5005
R5995 VOUT-.n24 VOUT-.t25 4.5005
R5996 VOUT-.n25 VOUT-.t127 4.5005
R5997 VOUT-.n26 VOUT-.t88 4.5005
R5998 VOUT-.n27 VOUT-.t53 4.5005
R5999 VOUT-.n28 VOUT-.t140 4.5005
R6000 VOUT-.n30 VOUT-.t109 4.5005
R6001 VOUT-.n29 VOUT-.t78 4.5005
R6002 VOUT-.n31 VOUT-.t112 4.5005
R6003 VOUT-.n33 VOUT-.t77 4.5005
R6004 VOUT-.n32 VOUT-.t37 4.5005
R6005 VOUT-.n34 VOUT-.t147 4.5005
R6006 VOUT-.n36 VOUT-.t116 4.5005
R6007 VOUT-.n35 VOUT-.t81 4.5005
R6008 VOUT-.n37 VOUT-.t46 4.5005
R6009 VOUT-.n39 VOUT-.t153 4.5005
R6010 VOUT-.n38 VOUT-.t122 4.5005
R6011 VOUT-.n40 VOUT-.t154 4.5005
R6012 VOUT-.n42 VOUT-.t123 4.5005
R6013 VOUT-.n41 VOUT-.t84 4.5005
R6014 VOUT-.n43 VOUT-.t52 4.5005
R6015 VOUT-.n45 VOUT-.t22 4.5005
R6016 VOUT-.n44 VOUT-.t126 4.5005
R6017 VOUT-.n99 VOUT-.t142 4.5005
R6018 VOUT-.n98 VOUT-.t93 4.5005
R6019 VOUT-.n97 VOUT-.t58 4.5005
R6020 VOUT-.n96 VOUT-.t30 4.5005
R6021 VOUT-.n16 VOUT-.n14 4.5005
R6022 VOUT-.n3 VOUT-.t0 3.42907
R6023 VOUT-.n3 VOUT-.t16 3.42907
R6024 VOUT-.n1 VOUT-.t13 3.42907
R6025 VOUT-.n1 VOUT-.t18 3.42907
R6026 VOUT-.n0 VOUT-.t17 3.42907
R6027 VOUT-.n0 VOUT-.t9 3.42907
R6028 VOUT- VOUT-.n5 2.84425
R6029 VOUT-.n5 VOUT-.n4 2.03175
R6030 VOUT-.n4 VOUT-.n2 1.1255
R6031 VOUT-.n11 VOUT-.n9 0.563
R6032 VOUT-.n13 VOUT-.n11 0.563
R6033 VOUT-.n14 VOUT-.n13 0.563
R6034 VOUT-.n47 VOUT-.n46 0.3295
R6035 VOUT-.n50 VOUT-.n49 0.3295
R6036 VOUT-.n49 VOUT-.n48 0.3295
R6037 VOUT-.n53 VOUT-.n52 0.3295
R6038 VOUT-.n52 VOUT-.n51 0.3295
R6039 VOUT-.n56 VOUT-.n55 0.3295
R6040 VOUT-.n55 VOUT-.n54 0.3295
R6041 VOUT-.n59 VOUT-.n58 0.3295
R6042 VOUT-.n58 VOUT-.n57 0.3295
R6043 VOUT-.n61 VOUT-.n60 0.3295
R6044 VOUT-.n62 VOUT-.n61 0.3295
R6045 VOUT-.n63 VOUT-.n62 0.3295
R6046 VOUT-.n64 VOUT-.n63 0.3295
R6047 VOUT-.n65 VOUT-.n64 0.3295
R6048 VOUT-.n66 VOUT-.n65 0.3295
R6049 VOUT-.n67 VOUT-.n66 0.3295
R6050 VOUT-.n68 VOUT-.n67 0.3295
R6051 VOUT-.n69 VOUT-.n68 0.3295
R6052 VOUT-.n71 VOUT-.n69 0.3295
R6053 VOUT-.n71 VOUT-.n70 0.3295
R6054 VOUT-.n74 VOUT-.n72 0.3295
R6055 VOUT-.n74 VOUT-.n73 0.3295
R6056 VOUT-.n77 VOUT-.n75 0.3295
R6057 VOUT-.n77 VOUT-.n76 0.3295
R6058 VOUT-.n80 VOUT-.n78 0.3295
R6059 VOUT-.n80 VOUT-.n79 0.3295
R6060 VOUT-.n83 VOUT-.n81 0.3295
R6061 VOUT-.n83 VOUT-.n82 0.3295
R6062 VOUT-.n86 VOUT-.n84 0.3295
R6063 VOUT-.n86 VOUT-.n85 0.3295
R6064 VOUT-.n89 VOUT-.n87 0.3295
R6065 VOUT-.n89 VOUT-.n88 0.3295
R6066 VOUT-.n92 VOUT-.n90 0.3295
R6067 VOUT-.n92 VOUT-.n91 0.3295
R6068 VOUT-.n95 VOUT-.n93 0.3295
R6069 VOUT-.n95 VOUT-.n94 0.3295
R6070 VOUT-.n18 VOUT-.n17 0.3295
R6071 VOUT-.n20 VOUT-.n19 0.3295
R6072 VOUT-.n21 VOUT-.n20 0.3295
R6073 VOUT-.n22 VOUT-.n21 0.3295
R6074 VOUT-.n23 VOUT-.n22 0.3295
R6075 VOUT-.n24 VOUT-.n23 0.3295
R6076 VOUT-.n25 VOUT-.n24 0.3295
R6077 VOUT-.n26 VOUT-.n25 0.3295
R6078 VOUT-.n27 VOUT-.n26 0.3295
R6079 VOUT-.n28 VOUT-.n27 0.3295
R6080 VOUT-.n30 VOUT-.n28 0.3295
R6081 VOUT-.n30 VOUT-.n29 0.3295
R6082 VOUT-.n33 VOUT-.n31 0.3295
R6083 VOUT-.n33 VOUT-.n32 0.3295
R6084 VOUT-.n36 VOUT-.n34 0.3295
R6085 VOUT-.n36 VOUT-.n35 0.3295
R6086 VOUT-.n39 VOUT-.n37 0.3295
R6087 VOUT-.n39 VOUT-.n38 0.3295
R6088 VOUT-.n42 VOUT-.n40 0.3295
R6089 VOUT-.n42 VOUT-.n41 0.3295
R6090 VOUT-.n45 VOUT-.n43 0.3295
R6091 VOUT-.n45 VOUT-.n44 0.3295
R6092 VOUT-.n99 VOUT-.n98 0.3295
R6093 VOUT-.n98 VOUT-.n97 0.3295
R6094 VOUT-.n97 VOUT-.n96 0.3295
R6095 VOUT-.n67 VOUT-.n50 0.306
R6096 VOUT-.n66 VOUT-.n53 0.306
R6097 VOUT-.n65 VOUT-.n56 0.306
R6098 VOUT-.n64 VOUT-.n59 0.306
R6099 VOUT-.n71 VOUT-.n47 0.2825
R6100 VOUT-.n74 VOUT-.n71 0.2825
R6101 VOUT-.n77 VOUT-.n74 0.2825
R6102 VOUT-.n80 VOUT-.n77 0.2825
R6103 VOUT-.n83 VOUT-.n80 0.2825
R6104 VOUT-.n86 VOUT-.n83 0.2825
R6105 VOUT-.n89 VOUT-.n86 0.2825
R6106 VOUT-.n92 VOUT-.n89 0.2825
R6107 VOUT-.n95 VOUT-.n92 0.2825
R6108 VOUT-.n30 VOUT-.n18 0.2825
R6109 VOUT-.n33 VOUT-.n30 0.2825
R6110 VOUT-.n36 VOUT-.n33 0.2825
R6111 VOUT-.n39 VOUT-.n36 0.2825
R6112 VOUT-.n42 VOUT-.n39 0.2825
R6113 VOUT-.n45 VOUT-.n42 0.2825
R6114 VOUT-.n97 VOUT-.n45 0.2825
R6115 VOUT-.n97 VOUT-.n95 0.2825
R6116 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.cap_res_X.t0 49.083
R6117 two_stage_opamp_dummy_magic_0.cap_res_X.t138 two_stage_opamp_dummy_magic_0.cap_res_X.t118 0.1603
R6118 two_stage_opamp_dummy_magic_0.cap_res_X.t101 two_stage_opamp_dummy_magic_0.cap_res_X.t74 0.1603
R6119 two_stage_opamp_dummy_magic_0.cap_res_X.t37 two_stage_opamp_dummy_magic_0.cap_res_X.t21 0.1603
R6120 two_stage_opamp_dummy_magic_0.cap_res_X.t106 two_stage_opamp_dummy_magic_0.cap_res_X.t123 0.1603
R6121 two_stage_opamp_dummy_magic_0.cap_res_X.t6 two_stage_opamp_dummy_magic_0.cap_res_X.t121 0.1603
R6122 two_stage_opamp_dummy_magic_0.cap_res_X.t70 two_stage_opamp_dummy_magic_0.cap_res_X.t89 0.1603
R6123 two_stage_opamp_dummy_magic_0.cap_res_X.t40 two_stage_opamp_dummy_magic_0.cap_res_X.t93 0.1603
R6124 two_stage_opamp_dummy_magic_0.cap_res_X.t115 two_stage_opamp_dummy_magic_0.cap_res_X.t63 0.1603
R6125 two_stage_opamp_dummy_magic_0.cap_res_X.t78 two_stage_opamp_dummy_magic_0.cap_res_X.t128 0.1603
R6126 two_stage_opamp_dummy_magic_0.cap_res_X.t16 two_stage_opamp_dummy_magic_0.cap_res_X.t103 0.1603
R6127 two_stage_opamp_dummy_magic_0.cap_res_X.t49 two_stage_opamp_dummy_magic_0.cap_res_X.t100 0.1603
R6128 two_stage_opamp_dummy_magic_0.cap_res_X.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t68 0.1603
R6129 two_stage_opamp_dummy_magic_0.cap_res_X.t87 two_stage_opamp_dummy_magic_0.cap_res_X.t137 0.1603
R6130 two_stage_opamp_dummy_magic_0.cap_res_X.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t109 0.1603
R6131 two_stage_opamp_dummy_magic_0.cap_res_X.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t36 0.1603
R6132 two_stage_opamp_dummy_magic_0.cap_res_X.t59 two_stage_opamp_dummy_magic_0.cap_res_X.t9 0.1603
R6133 two_stage_opamp_dummy_magic_0.cap_res_X.t92 two_stage_opamp_dummy_magic_0.cap_res_X.t5 0.1603
R6134 two_stage_opamp_dummy_magic_0.cap_res_X.t24 two_stage_opamp_dummy_magic_0.cap_res_X.t114 0.1603
R6135 two_stage_opamp_dummy_magic_0.cap_res_X.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t42 0.1603
R6136 two_stage_opamp_dummy_magic_0.cap_res_X.t64 two_stage_opamp_dummy_magic_0.cap_res_X.t15 0.1603
R6137 two_stage_opamp_dummy_magic_0.cap_res_X.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t81 0.1603
R6138 two_stage_opamp_dummy_magic_0.cap_res_X.t105 two_stage_opamp_dummy_magic_0.cap_res_X.t53 0.1603
R6139 two_stage_opamp_dummy_magic_0.cap_res_X.t73 two_stage_opamp_dummy_magic_0.cap_res_X.t122 0.1603
R6140 two_stage_opamp_dummy_magic_0.cap_res_X.t3 two_stage_opamp_dummy_magic_0.cap_res_X.t90 0.1603
R6141 two_stage_opamp_dummy_magic_0.cap_res_X.t35 two_stage_opamp_dummy_magic_0.cap_res_X.t88 0.1603
R6142 two_stage_opamp_dummy_magic_0.cap_res_X.t111 two_stage_opamp_dummy_magic_0.cap_res_X.t58 0.1603
R6143 two_stage_opamp_dummy_magic_0.cap_res_X.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t125 0.1603
R6144 two_stage_opamp_dummy_magic_0.cap_res_X.t10 two_stage_opamp_dummy_magic_0.cap_res_X.t98 0.1603
R6145 two_stage_opamp_dummy_magic_0.cap_res_X.t120 two_stage_opamp_dummy_magic_0.cap_res_X.t28 0.1603
R6146 two_stage_opamp_dummy_magic_0.cap_res_X.t45 two_stage_opamp_dummy_magic_0.cap_res_X.t133 0.1603
R6147 two_stage_opamp_dummy_magic_0.cap_res_X.t79 two_stage_opamp_dummy_magic_0.cap_res_X.t129 0.1603
R6148 two_stage_opamp_dummy_magic_0.cap_res_X.t71 two_stage_opamp_dummy_magic_0.cap_res_X.t7 0.1603
R6149 two_stage_opamp_dummy_magic_0.cap_res_X.t107 two_stage_opamp_dummy_magic_0.cap_res_X.t95 0.1603
R6150 two_stage_opamp_dummy_magic_0.cap_res_X.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t134 0.1603
R6151 two_stage_opamp_dummy_magic_0.cap_res_X.t52 two_stage_opamp_dummy_magic_0.cap_res_X.t85 0.1603
R6152 two_stage_opamp_dummy_magic_0.cap_res_X.t84 two_stage_opamp_dummy_magic_0.cap_res_X.t33 0.1603
R6153 two_stage_opamp_dummy_magic_0.cap_res_X.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t75 0.1603
R6154 two_stage_opamp_dummy_magic_0.cap_res_X.t30 two_stage_opamp_dummy_magic_0.cap_res_X.t27 0.1603
R6155 two_stage_opamp_dummy_magic_0.cap_res_X.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t116 0.1603
R6156 two_stage_opamp_dummy_magic_0.cap_res_X.t104 two_stage_opamp_dummy_magic_0.cap_res_X.t66 0.1603
R6157 two_stage_opamp_dummy_magic_0.cap_res_X.t17 two_stage_opamp_dummy_magic_0.cap_res_X.t110 0.1603
R6158 two_stage_opamp_dummy_magic_0.cap_res_X.t8 two_stage_opamp_dummy_magic_0.cap_res_X.t50 0.1603
R6159 two_stage_opamp_dummy_magic_0.cap_res_X.t26 two_stage_opamp_dummy_magic_0.cap_res_X.t67 0.1603
R6160 two_stage_opamp_dummy_magic_0.cap_res_X.t54 two_stage_opamp_dummy_magic_0.cap_res_X.t26 0.1603
R6161 two_stage_opamp_dummy_magic_0.cap_res_X.t86 two_stage_opamp_dummy_magic_0.cap_res_X.t54 0.1603
R6162 two_stage_opamp_dummy_magic_0.cap_res_X.t46 two_stage_opamp_dummy_magic_0.cap_res_X.t86 0.1603
R6163 two_stage_opamp_dummy_magic_0.cap_res_X.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t83 0.1603
R6164 two_stage_opamp_dummy_magic_0.cap_res_X.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t44 0.1603
R6165 two_stage_opamp_dummy_magic_0.cap_res_X.t32 two_stage_opamp_dummy_magic_0.cap_res_X.t136 0.1603
R6166 two_stage_opamp_dummy_magic_0.cap_res_X.t130 two_stage_opamp_dummy_magic_0.cap_res_X.t32 0.1603
R6167 two_stage_opamp_dummy_magic_0.cap_res_X.t97 two_stage_opamp_dummy_magic_0.cap_res_X.t131 0.1603
R6168 two_stage_opamp_dummy_magic_0.cap_res_X.t117 two_stage_opamp_dummy_magic_0.cap_res_X.t97 0.1603
R6169 two_stage_opamp_dummy_magic_0.cap_res_X.t14 two_stage_opamp_dummy_magic_0.cap_res_X.t117 0.1603
R6170 two_stage_opamp_dummy_magic_0.cap_res_X.t113 two_stage_opamp_dummy_magic_0.cap_res_X.t14 0.1603
R6171 two_stage_opamp_dummy_magic_0.cap_res_X.t51 two_stage_opamp_dummy_magic_0.cap_res_X.t13 0.1603
R6172 two_stage_opamp_dummy_magic_0.cap_res_X.t19 two_stage_opamp_dummy_magic_0.cap_res_X.t51 0.1603
R6173 two_stage_opamp_dummy_magic_0.cap_res_X.t126 two_stage_opamp_dummy_magic_0.cap_res_X.t19 0.1603
R6174 two_stage_opamp_dummy_magic_0.cap_res_X.t29 two_stage_opamp_dummy_magic_0.cap_res_X.t126 0.1603
R6175 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t62 0.159278
R6176 two_stage_opamp_dummy_magic_0.cap_res_X.t48 two_stage_opamp_dummy_magic_0.cap_res_X.n15 0.159278
R6177 two_stage_opamp_dummy_magic_0.cap_res_X.t80 two_stage_opamp_dummy_magic_0.cap_res_X.n16 0.159278
R6178 two_stage_opamp_dummy_magic_0.cap_res_X.t41 two_stage_opamp_dummy_magic_0.cap_res_X.n17 0.159278
R6179 two_stage_opamp_dummy_magic_0.cap_res_X.t4 two_stage_opamp_dummy_magic_0.cap_res_X.n18 0.159278
R6180 two_stage_opamp_dummy_magic_0.cap_res_X.t34 two_stage_opamp_dummy_magic_0.cap_res_X.n19 0.159278
R6181 two_stage_opamp_dummy_magic_0.cap_res_X.t135 two_stage_opamp_dummy_magic_0.cap_res_X.n20 0.159278
R6182 two_stage_opamp_dummy_magic_0.cap_res_X.t99 two_stage_opamp_dummy_magic_0.cap_res_X.n21 0.159278
R6183 two_stage_opamp_dummy_magic_0.cap_res_X.t60 two_stage_opamp_dummy_magic_0.cap_res_X.n22 0.159278
R6184 two_stage_opamp_dummy_magic_0.cap_res_X.t91 two_stage_opamp_dummy_magic_0.cap_res_X.n23 0.159278
R6185 two_stage_opamp_dummy_magic_0.cap_res_X.t55 two_stage_opamp_dummy_magic_0.cap_res_X.n24 0.159278
R6186 two_stage_opamp_dummy_magic_0.cap_res_X.t18 two_stage_opamp_dummy_magic_0.cap_res_X.n25 0.159278
R6187 two_stage_opamp_dummy_magic_0.cap_res_X.t47 two_stage_opamp_dummy_magic_0.cap_res_X.n26 0.159278
R6188 two_stage_opamp_dummy_magic_0.cap_res_X.t12 two_stage_opamp_dummy_magic_0.cap_res_X.n27 0.159278
R6189 two_stage_opamp_dummy_magic_0.cap_res_X.t108 two_stage_opamp_dummy_magic_0.cap_res_X.n28 0.159278
R6190 two_stage_opamp_dummy_magic_0.cap_res_X.t1 two_stage_opamp_dummy_magic_0.cap_res_X.n29 0.159278
R6191 two_stage_opamp_dummy_magic_0.cap_res_X.t102 two_stage_opamp_dummy_magic_0.cap_res_X.n30 0.159278
R6192 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t25 0.159278
R6193 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t43 0.159278
R6194 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t11 0.159278
R6195 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t2 0.159278
R6196 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.t38 0.159278
R6197 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.t23 0.159278
R6198 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.t56 0.159278
R6199 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.t94 0.159278
R6200 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.t72 0.159278
R6201 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.t112 0.159278
R6202 two_stage_opamp_dummy_magic_0.cap_res_X.t62 two_stage_opamp_dummy_magic_0.cap_res_X.t101 0.137822
R6203 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t138 0.1368
R6204 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t37 0.1368
R6205 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t106 0.1368
R6206 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t6 0.1368
R6207 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t70 0.1368
R6208 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t40 0.1368
R6209 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t115 0.1368
R6210 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t78 0.1368
R6211 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t16 0.1368
R6212 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t49 0.1368
R6213 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t119 0.1368
R6214 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t87 0.1368
R6215 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t22 0.1368
R6216 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t124 0.1368
R6217 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t59 0.1368
R6218 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t92 0.1368
R6219 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t24 0.1368
R6220 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t127 0.1368
R6221 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t64 0.1368
R6222 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t31 0.1368
R6223 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t105 0.1368
R6224 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t73 0.1368
R6225 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t3 0.1368
R6226 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t35 0.1368
R6227 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t111 0.1368
R6228 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t76 0.1368
R6229 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t10 0.1368
R6230 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t120 0.1368
R6231 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t45 0.1368
R6232 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t79 0.1368
R6233 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t8 0.1368
R6234 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.cap_res_X.t29 0.118
R6235 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.t71 0.114322
R6236 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.n6 0.1133
R6237 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.n7 0.1133
R6238 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.n8 0.1133
R6239 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.n9 0.1133
R6240 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.n10 0.1133
R6241 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.n11 0.1133
R6242 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.n12 0.1133
R6243 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.n13 0.1133
R6244 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.n14 0.1133
R6245 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.n31 0.1133
R6246 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.n32 0.1133
R6247 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.n33 0.1133
R6248 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.n0 0.1133
R6249 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.n1 0.1133
R6250 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.n2 0.1133
R6251 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.n3 0.1133
R6252 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.n4 0.1133
R6253 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n5 0.1133
R6254 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n34 0.1133
R6255 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.t107 0.00152174
R6256 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.t20 0.00152174
R6257 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.t52 0.00152174
R6258 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.t84 0.00152174
R6259 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.t132 0.00152174
R6260 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t30 0.00152174
R6261 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t69 0.00152174
R6262 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t104 0.00152174
R6263 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t17 0.00152174
R6264 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t57 0.00152174
R6265 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t48 0.00152174
R6266 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t80 0.00152174
R6267 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t41 0.00152174
R6268 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t4 0.00152174
R6269 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t34 0.00152174
R6270 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t135 0.00152174
R6271 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t99 0.00152174
R6272 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t60 0.00152174
R6273 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t91 0.00152174
R6274 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t55 0.00152174
R6275 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t18 0.00152174
R6276 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t47 0.00152174
R6277 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t12 0.00152174
R6278 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t108 0.00152174
R6279 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t1 0.00152174
R6280 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t102 0.00152174
R6281 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t65 0.00152174
R6282 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t82 0.00152174
R6283 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t46 0.00152174
R6284 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t39 0.00152174
R6285 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.t77 0.00152174
R6286 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.t61 0.00152174
R6287 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.t96 0.00152174
R6288 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.t130 0.00152174
R6289 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.t113 0.00152174
R6290 two_stage_opamp_dummy_magic_0.cap_res_X.t13 two_stage_opamp_dummy_magic_0.cap_res_X.n35 0.00152174
R6291 bgr_0.Vbe2.n125 bgr_0.Vbe2.t0 162.458
R6292 bgr_0.Vbe2.n142 bgr_0.Vbe2.n1 83.5719
R6293 bgr_0.Vbe2.n134 bgr_0.Vbe2.n2 83.5719
R6294 bgr_0.Vbe2.n136 bgr_0.Vbe2.n135 83.5719
R6295 bgr_0.Vbe2.n128 bgr_0.Vbe2.n7 83.5719
R6296 bgr_0.Vbe2.n120 bgr_0.Vbe2.n8 83.5719
R6297 bgr_0.Vbe2.n122 bgr_0.Vbe2.n121 83.5719
R6298 bgr_0.Vbe2.n114 bgr_0.Vbe2.n12 83.5719
R6299 bgr_0.Vbe2.n109 bgr_0.Vbe2.n13 83.5719
R6300 bgr_0.Vbe2.n51 bgr_0.Vbe2.n50 83.5719
R6301 bgr_0.Vbe2.n49 bgr_0.Vbe2.n48 83.5719
R6302 bgr_0.Vbe2.n47 bgr_0.Vbe2.n46 83.5719
R6303 bgr_0.Vbe2.n65 bgr_0.Vbe2.n64 83.5719
R6304 bgr_0.Vbe2.n63 bgr_0.Vbe2.n62 83.5719
R6305 bgr_0.Vbe2.n33 bgr_0.Vbe2.n32 83.5719
R6306 bgr_0.Vbe2.n73 bgr_0.Vbe2.n72 83.5719
R6307 bgr_0.Vbe2.n28 bgr_0.Vbe2.n26 83.5719
R6308 bgr_0.Vbe2.n78 bgr_0.Vbe2.n25 83.5719
R6309 bgr_0.Vbe2.n86 bgr_0.Vbe2.n85 83.5719
R6310 bgr_0.Vbe2.n23 bgr_0.Vbe2.n22 83.5719
R6311 bgr_0.Vbe2.n101 bgr_0.Vbe2.n100 83.5719
R6312 bgr_0.Vbe2.n99 bgr_0.Vbe2.n98 83.5719
R6313 bgr_0.Vbe2.n97 bgr_0.Vbe2.n96 83.5719
R6314 bgr_0.Vbe2.n59 bgr_0.Vbe2.n32 73.8495
R6315 bgr_0.Vbe2.n144 bgr_0.Vbe2.n1 73.3165
R6316 bgr_0.Vbe2.n130 bgr_0.Vbe2.n7 73.3165
R6317 bgr_0.Vbe2.n116 bgr_0.Vbe2.n12 73.3165
R6318 bgr_0.Vbe2.n50 bgr_0.Vbe2.n42 73.3165
R6319 bgr_0.Vbe2.n72 bgr_0.Vbe2.n71 73.3165
R6320 bgr_0.Vbe2.n85 bgr_0.Vbe2.n84 73.3165
R6321 bgr_0.Vbe2.n102 bgr_0.Vbe2.n101 73.3165
R6322 bgr_0.Vbe2.n135 bgr_0.Vbe2.n133 73.19
R6323 bgr_0.Vbe2.n121 bgr_0.Vbe2.n119 73.19
R6324 bgr_0.Vbe2.n47 bgr_0.Vbe2.n45 73.19
R6325 bgr_0.Vbe2.n64 bgr_0.Vbe2.n29 73.19
R6326 bgr_0.Vbe2.n80 bgr_0.Vbe2.n25 73.19
R6327 bgr_0.Vbe2.n97 bgr_0.Vbe2.n19 73.19
R6328 bgr_0.Vbe2.n110 bgr_0.Vbe2.t5 65.0299
R6329 bgr_0.Vbe2.t7 bgr_0.Vbe2.n20 65.0299
R6330 bgr_0.Vbe2.n134 bgr_0.Vbe2.n1 26.074
R6331 bgr_0.Vbe2.n120 bgr_0.Vbe2.n7 26.074
R6332 bgr_0.Vbe2.n109 bgr_0.Vbe2.n12 26.074
R6333 bgr_0.Vbe2.n50 bgr_0.Vbe2.n49 26.074
R6334 bgr_0.Vbe2.n63 bgr_0.Vbe2.n32 26.074
R6335 bgr_0.Vbe2.n72 bgr_0.Vbe2.n28 26.074
R6336 bgr_0.Vbe2.n85 bgr_0.Vbe2.n23 26.074
R6337 bgr_0.Vbe2.n101 bgr_0.Vbe2.n99 26.074
R6338 bgr_0.Vbe2.n135 bgr_0.Vbe2.t1 25.7843
R6339 bgr_0.Vbe2.n121 bgr_0.Vbe2.t8 25.7843
R6340 bgr_0.Vbe2.t3 bgr_0.Vbe2.n47 25.7843
R6341 bgr_0.Vbe2.n64 bgr_0.Vbe2.t4 25.7843
R6342 bgr_0.Vbe2.t2 bgr_0.Vbe2.n25 25.7843
R6343 bgr_0.Vbe2.t6 bgr_0.Vbe2.n97 25.7843
R6344 bgr_0.Vbe2.n103 bgr_0.Vbe2.n91 9.3005
R6345 bgr_0.Vbe2.n91 bgr_0.Vbe2.n17 9.3005
R6346 bgr_0.Vbe2.n91 bgr_0.Vbe2.n18 9.3005
R6347 bgr_0.Vbe2.n107 bgr_0.Vbe2.n91 9.3005
R6348 bgr_0.Vbe2.n93 bgr_0.Vbe2.n17 9.3005
R6349 bgr_0.Vbe2.n93 bgr_0.Vbe2.n18 9.3005
R6350 bgr_0.Vbe2.n93 bgr_0.Vbe2.n15 9.3005
R6351 bgr_0.Vbe2.n107 bgr_0.Vbe2.n93 9.3005
R6352 bgr_0.Vbe2.n108 bgr_0.Vbe2.n17 9.3005
R6353 bgr_0.Vbe2.n108 bgr_0.Vbe2.n16 9.3005
R6354 bgr_0.Vbe2.n108 bgr_0.Vbe2.n18 9.3005
R6355 bgr_0.Vbe2.n108 bgr_0.Vbe2.n15 9.3005
R6356 bgr_0.Vbe2.n108 bgr_0.Vbe2.n107 9.3005
R6357 bgr_0.Vbe2.n107 bgr_0.Vbe2.n95 9.3005
R6358 bgr_0.Vbe2.n95 bgr_0.Vbe2.n15 9.3005
R6359 bgr_0.Vbe2.n95 bgr_0.Vbe2.n18 9.3005
R6360 bgr_0.Vbe2.n95 bgr_0.Vbe2.n16 9.3005
R6361 bgr_0.Vbe2.n107 bgr_0.Vbe2.n90 9.3005
R6362 bgr_0.Vbe2.n90 bgr_0.Vbe2.n15 9.3005
R6363 bgr_0.Vbe2.n90 bgr_0.Vbe2.n18 9.3005
R6364 bgr_0.Vbe2.n90 bgr_0.Vbe2.n16 9.3005
R6365 bgr_0.Vbe2.n103 bgr_0.Vbe2.n90 9.3005
R6366 bgr_0.Vbe2.n106 bgr_0.Vbe2.n17 9.3005
R6367 bgr_0.Vbe2.n106 bgr_0.Vbe2.n16 9.3005
R6368 bgr_0.Vbe2.n106 bgr_0.Vbe2.n18 9.3005
R6369 bgr_0.Vbe2.n107 bgr_0.Vbe2.n106 9.3005
R6370 bgr_0.Vbe2.n56 bgr_0.Vbe2.n55 9.3005
R6371 bgr_0.Vbe2.n55 bgr_0.Vbe2.n54 9.3005
R6372 bgr_0.Vbe2.n55 bgr_0.Vbe2.n35 9.3005
R6373 bgr_0.Vbe2.n55 bgr_0.Vbe2.n36 9.3005
R6374 bgr_0.Vbe2.n54 bgr_0.Vbe2.n52 9.3005
R6375 bgr_0.Vbe2.n52 bgr_0.Vbe2.n35 9.3005
R6376 bgr_0.Vbe2.n52 bgr_0.Vbe2.n37 9.3005
R6377 bgr_0.Vbe2.n52 bgr_0.Vbe2.n36 9.3005
R6378 bgr_0.Vbe2.n54 bgr_0.Vbe2.n3 9.3005
R6379 bgr_0.Vbe2.n38 bgr_0.Vbe2.n3 9.3005
R6380 bgr_0.Vbe2.n35 bgr_0.Vbe2.n3 9.3005
R6381 bgr_0.Vbe2.n37 bgr_0.Vbe2.n3 9.3005
R6382 bgr_0.Vbe2.n36 bgr_0.Vbe2.n3 9.3005
R6383 bgr_0.Vbe2.n39 bgr_0.Vbe2.n36 9.3005
R6384 bgr_0.Vbe2.n39 bgr_0.Vbe2.n37 9.3005
R6385 bgr_0.Vbe2.n39 bgr_0.Vbe2.n35 9.3005
R6386 bgr_0.Vbe2.n39 bgr_0.Vbe2.n38 9.3005
R6387 bgr_0.Vbe2.n57 bgr_0.Vbe2.n36 9.3005
R6388 bgr_0.Vbe2.n57 bgr_0.Vbe2.n37 9.3005
R6389 bgr_0.Vbe2.n57 bgr_0.Vbe2.n35 9.3005
R6390 bgr_0.Vbe2.n57 bgr_0.Vbe2.n38 9.3005
R6391 bgr_0.Vbe2.n57 bgr_0.Vbe2.n56 9.3005
R6392 bgr_0.Vbe2.n54 bgr_0.Vbe2.n53 9.3005
R6393 bgr_0.Vbe2.n53 bgr_0.Vbe2.n38 9.3005
R6394 bgr_0.Vbe2.n53 bgr_0.Vbe2.n35 9.3005
R6395 bgr_0.Vbe2.n53 bgr_0.Vbe2.n36 9.3005
R6396 bgr_0.Vbe2.n105 bgr_0.Vbe2.n15 4.64654
R6397 bgr_0.Vbe2.n92 bgr_0.Vbe2.n16 4.64654
R6398 bgr_0.Vbe2.n103 bgr_0.Vbe2.n14 4.64654
R6399 bgr_0.Vbe2.n94 bgr_0.Vbe2.n17 4.64654
R6400 bgr_0.Vbe2.n104 bgr_0.Vbe2.n103 4.64654
R6401 bgr_0.Vbe2.n43 bgr_0.Vbe2.n37 4.64654
R6402 bgr_0.Vbe2.n44 bgr_0.Vbe2.n38 4.64654
R6403 bgr_0.Vbe2.n56 bgr_0.Vbe2.n41 4.64654
R6404 bgr_0.Vbe2.n54 bgr_0.Vbe2.n34 4.64654
R6405 bgr_0.Vbe2.n56 bgr_0.Vbe2.n40 4.64654
R6406 bgr_0.Vbe2.n133 bgr_0.Vbe2.n132 2.36206
R6407 bgr_0.Vbe2.n119 bgr_0.Vbe2.n118 2.36206
R6408 bgr_0.Vbe2.n68 bgr_0.Vbe2.n29 2.36206
R6409 bgr_0.Vbe2.n81 bgr_0.Vbe2.n80 2.36206
R6410 bgr_0.Vbe2.n145 bgr_0.Vbe2.n144 2.19742
R6411 bgr_0.Vbe2.n131 bgr_0.Vbe2.n130 2.19742
R6412 bgr_0.Vbe2.n117 bgr_0.Vbe2.n116 2.19742
R6413 bgr_0.Vbe2.n71 bgr_0.Vbe2.n69 2.19742
R6414 bgr_0.Vbe2.n84 bgr_0.Vbe2.n82 2.19742
R6415 bgr_0.Vbe2.n110 bgr_0.Vbe2.n13 1.56363
R6416 bgr_0.Vbe2.n22 bgr_0.Vbe2.n20 1.56363
R6417 bgr_0.Vbe2.n83 bgr_0.Vbe2.n21 1.5505
R6418 bgr_0.Vbe2.n88 bgr_0.Vbe2.n87 1.5505
R6419 bgr_0.Vbe2.n70 bgr_0.Vbe2.n27 1.5505
R6420 bgr_0.Vbe2.n75 bgr_0.Vbe2.n74 1.5505
R6421 bgr_0.Vbe2.n77 bgr_0.Vbe2.n76 1.5505
R6422 bgr_0.Vbe2.n79 bgr_0.Vbe2.n24 1.5505
R6423 bgr_0.Vbe2.n61 bgr_0.Vbe2.n60 1.5505
R6424 bgr_0.Vbe2.n67 bgr_0.Vbe2.n66 1.5505
R6425 bgr_0.Vbe2.n31 bgr_0.Vbe2.n30 1.5505
R6426 bgr_0.Vbe2.n115 bgr_0.Vbe2.n11 1.5505
R6427 bgr_0.Vbe2.n113 bgr_0.Vbe2.n112 1.5505
R6428 bgr_0.Vbe2.n129 bgr_0.Vbe2.n6 1.5505
R6429 bgr_0.Vbe2.n127 bgr_0.Vbe2.n126 1.5505
R6430 bgr_0.Vbe2.n124 bgr_0.Vbe2.n123 1.5505
R6431 bgr_0.Vbe2.n10 bgr_0.Vbe2.n9 1.5505
R6432 bgr_0.Vbe2.n143 bgr_0.Vbe2.n0 1.5505
R6433 bgr_0.Vbe2.n141 bgr_0.Vbe2.n140 1.5505
R6434 bgr_0.Vbe2.n138 bgr_0.Vbe2.n137 1.5505
R6435 bgr_0.Vbe2.n5 bgr_0.Vbe2.n4 1.5505
R6436 bgr_0.Vbe2.n136 bgr_0.Vbe2.n5 1.25468
R6437 bgr_0.Vbe2.n122 bgr_0.Vbe2.n10 1.25468
R6438 bgr_0.Vbe2.n46 bgr_0.Vbe2.n37 1.25468
R6439 bgr_0.Vbe2.n66 bgr_0.Vbe2.n65 1.25468
R6440 bgr_0.Vbe2.n79 bgr_0.Vbe2.n78 1.25468
R6441 bgr_0.Vbe2.n96 bgr_0.Vbe2.n15 1.25468
R6442 bgr_0.Vbe2.n144 bgr_0.Vbe2.n143 1.19225
R6443 bgr_0.Vbe2.n130 bgr_0.Vbe2.n129 1.19225
R6444 bgr_0.Vbe2.n116 bgr_0.Vbe2.n115 1.19225
R6445 bgr_0.Vbe2.n54 bgr_0.Vbe2.n42 1.19225
R6446 bgr_0.Vbe2.n71 bgr_0.Vbe2.n70 1.19225
R6447 bgr_0.Vbe2.n84 bgr_0.Vbe2.n83 1.19225
R6448 bgr_0.Vbe2.n102 bgr_0.Vbe2.n17 1.19225
R6449 bgr_0.Vbe2.n137 bgr_0.Vbe2.n2 1.07024
R6450 bgr_0.Vbe2.n123 bgr_0.Vbe2.n8 1.07024
R6451 bgr_0.Vbe2.n48 bgr_0.Vbe2.n35 1.07024
R6452 bgr_0.Vbe2.n62 bgr_0.Vbe2.n31 1.07024
R6453 bgr_0.Vbe2.n77 bgr_0.Vbe2.n26 1.07024
R6454 bgr_0.Vbe2.n98 bgr_0.Vbe2.n18 1.07024
R6455 bgr_0.Vbe2.n133 bgr_0.Vbe2.n5 1.0237
R6456 bgr_0.Vbe2.n119 bgr_0.Vbe2.n10 1.0237
R6457 bgr_0.Vbe2.n45 bgr_0.Vbe2.n37 1.0237
R6458 bgr_0.Vbe2.n66 bgr_0.Vbe2.n29 1.0237
R6459 bgr_0.Vbe2.n80 bgr_0.Vbe2.n79 1.0237
R6460 bgr_0.Vbe2.n19 bgr_0.Vbe2.n15 1.0237
R6461 bgr_0.Vbe2.n142 bgr_0.Vbe2.n141 0.885803
R6462 bgr_0.Vbe2.n128 bgr_0.Vbe2.n127 0.885803
R6463 bgr_0.Vbe2.n114 bgr_0.Vbe2.n113 0.885803
R6464 bgr_0.Vbe2.n51 bgr_0.Vbe2.n38 0.885803
R6465 bgr_0.Vbe2.n61 bgr_0.Vbe2.n33 0.885803
R6466 bgr_0.Vbe2.n74 bgr_0.Vbe2.n73 0.885803
R6467 bgr_0.Vbe2.n87 bgr_0.Vbe2.n86 0.885803
R6468 bgr_0.Vbe2.n100 bgr_0.Vbe2.n16 0.885803
R6469 bgr_0.Vbe2.n45 bgr_0.Vbe2.n36 0.812055
R6470 bgr_0.Vbe2.n107 bgr_0.Vbe2.n19 0.812055
R6471 bgr_0.Vbe2.n141 bgr_0.Vbe2.n2 0.77514
R6472 bgr_0.Vbe2.n127 bgr_0.Vbe2.n8 0.77514
R6473 bgr_0.Vbe2.n113 bgr_0.Vbe2.n13 0.77514
R6474 bgr_0.Vbe2.n48 bgr_0.Vbe2.n38 0.77514
R6475 bgr_0.Vbe2.n62 bgr_0.Vbe2.n61 0.77514
R6476 bgr_0.Vbe2.n74 bgr_0.Vbe2.n26 0.77514
R6477 bgr_0.Vbe2.n87 bgr_0.Vbe2.n22 0.77514
R6478 bgr_0.Vbe2.n98 bgr_0.Vbe2.n16 0.77514
R6479 bgr_0.Vbe2 bgr_0.Vbe2.n142 0.756696
R6480 bgr_0.Vbe2 bgr_0.Vbe2.n128 0.756696
R6481 bgr_0.Vbe2 bgr_0.Vbe2.n114 0.756696
R6482 bgr_0.Vbe2 bgr_0.Vbe2.n51 0.756696
R6483 bgr_0.Vbe2 bgr_0.Vbe2.n33 0.756696
R6484 bgr_0.Vbe2.n73 bgr_0.Vbe2 0.756696
R6485 bgr_0.Vbe2.n86 bgr_0.Vbe2 0.756696
R6486 bgr_0.Vbe2.n100 bgr_0.Vbe2 0.756696
R6487 bgr_0.Vbe2.n60 bgr_0.Vbe2.n59 0.711459
R6488 bgr_0.Vbe2.n56 bgr_0.Vbe2.n42 0.647417
R6489 bgr_0.Vbe2.n103 bgr_0.Vbe2.n102 0.647417
R6490 bgr_0.Vbe2.n137 bgr_0.Vbe2.n136 0.590702
R6491 bgr_0.Vbe2.n123 bgr_0.Vbe2.n122 0.590702
R6492 bgr_0.Vbe2.n46 bgr_0.Vbe2.n35 0.590702
R6493 bgr_0.Vbe2.n65 bgr_0.Vbe2.n31 0.590702
R6494 bgr_0.Vbe2.n78 bgr_0.Vbe2.n77 0.590702
R6495 bgr_0.Vbe2.n96 bgr_0.Vbe2.n18 0.590702
R6496 bgr_0.Vbe2.n59 bgr_0.Vbe2 0.576566
R6497 bgr_0.Vbe2.n89 bgr_0.Vbe2.n20 0.530034
R6498 bgr_0.Vbe2.n111 bgr_0.Vbe2.n110 0.530034
R6499 bgr_0.Vbe2.t1 bgr_0.Vbe2.n134 0.290206
R6500 bgr_0.Vbe2.t8 bgr_0.Vbe2.n120 0.290206
R6501 bgr_0.Vbe2.t5 bgr_0.Vbe2.n109 0.290206
R6502 bgr_0.Vbe2.n49 bgr_0.Vbe2.t3 0.290206
R6503 bgr_0.Vbe2.t4 bgr_0.Vbe2.n63 0.290206
R6504 bgr_0.Vbe2.n28 bgr_0.Vbe2.t2 0.290206
R6505 bgr_0.Vbe2.n23 bgr_0.Vbe2.t7 0.290206
R6506 bgr_0.Vbe2.n99 bgr_0.Vbe2.t6 0.290206
R6507 bgr_0.Vbe2.n143 bgr_0.Vbe2 0.203382
R6508 bgr_0.Vbe2.n129 bgr_0.Vbe2 0.203382
R6509 bgr_0.Vbe2.n115 bgr_0.Vbe2 0.203382
R6510 bgr_0.Vbe2.n54 bgr_0.Vbe2 0.203382
R6511 bgr_0.Vbe2.n70 bgr_0.Vbe2 0.203382
R6512 bgr_0.Vbe2.n83 bgr_0.Vbe2 0.203382
R6513 bgr_0.Vbe2 bgr_0.Vbe2.n17 0.203382
R6514 bgr_0.Vbe2.n82 bgr_0.Vbe2.n81 0.154071
R6515 bgr_0.Vbe2.n69 bgr_0.Vbe2.n68 0.154071
R6516 bgr_0.Vbe2.n118 bgr_0.Vbe2.n117 0.154071
R6517 bgr_0.Vbe2.n132 bgr_0.Vbe2.n131 0.154071
R6518 bgr_0.Vbe2.n111 bgr_0.Vbe2.n108 0.137464
R6519 bgr_0.Vbe2.n139 bgr_0.Vbe2.n3 0.137464
R6520 bgr_0.Vbe2.n90 bgr_0.Vbe2.n89 0.134964
R6521 bgr_0.Vbe2.n58 bgr_0.Vbe2.n57 0.134964
R6522 bgr_0.Vbe2 bgr_0.Vbe2.n145 0.0196071
R6523 bgr_0.Vbe2.n88 bgr_0.Vbe2.n21 0.0183571
R6524 bgr_0.Vbe2.n82 bgr_0.Vbe2.n21 0.0183571
R6525 bgr_0.Vbe2.n81 bgr_0.Vbe2.n24 0.0183571
R6526 bgr_0.Vbe2.n76 bgr_0.Vbe2.n24 0.0183571
R6527 bgr_0.Vbe2.n76 bgr_0.Vbe2.n75 0.0183571
R6528 bgr_0.Vbe2.n75 bgr_0.Vbe2.n27 0.0183571
R6529 bgr_0.Vbe2.n69 bgr_0.Vbe2.n27 0.0183571
R6530 bgr_0.Vbe2.n68 bgr_0.Vbe2.n67 0.0183571
R6531 bgr_0.Vbe2.n67 bgr_0.Vbe2.n30 0.0183571
R6532 bgr_0.Vbe2.n112 bgr_0.Vbe2.n11 0.0183571
R6533 bgr_0.Vbe2.n117 bgr_0.Vbe2.n11 0.0183571
R6534 bgr_0.Vbe2.n118 bgr_0.Vbe2.n9 0.0183571
R6535 bgr_0.Vbe2.n124 bgr_0.Vbe2.n9 0.0183571
R6536 bgr_0.Vbe2.n126 bgr_0.Vbe2.n6 0.0183571
R6537 bgr_0.Vbe2.n131 bgr_0.Vbe2.n6 0.0183571
R6538 bgr_0.Vbe2.n132 bgr_0.Vbe2.n4 0.0183571
R6539 bgr_0.Vbe2.n138 bgr_0.Vbe2.n4 0.0183571
R6540 bgr_0.Vbe2.n140 bgr_0.Vbe2.n0 0.0183571
R6541 bgr_0.Vbe2.n145 bgr_0.Vbe2.n0 0.0183571
R6542 bgr_0.Vbe2.n58 bgr_0.Vbe2.n30 0.0106786
R6543 bgr_0.Vbe2.n139 bgr_0.Vbe2.n138 0.0106786
R6544 bgr_0.Vbe2.n126 bgr_0.Vbe2.n125 0.00996429
R6545 bgr_0.Vbe2.n95 bgr_0.Vbe2.n94 0.00992001
R6546 bgr_0.Vbe2.n106 bgr_0.Vbe2.n104 0.00992001
R6547 bgr_0.Vbe2.n105 bgr_0.Vbe2.n91 0.00992001
R6548 bgr_0.Vbe2.n93 bgr_0.Vbe2.n92 0.00992001
R6549 bgr_0.Vbe2.n108 bgr_0.Vbe2.n14 0.00992001
R6550 bgr_0.Vbe2.n92 bgr_0.Vbe2.n91 0.00992001
R6551 bgr_0.Vbe2.n93 bgr_0.Vbe2.n14 0.00992001
R6552 bgr_0.Vbe2.n104 bgr_0.Vbe2.n95 0.00992001
R6553 bgr_0.Vbe2.n94 bgr_0.Vbe2.n90 0.00992001
R6554 bgr_0.Vbe2.n106 bgr_0.Vbe2.n105 0.00992001
R6555 bgr_0.Vbe2.n39 bgr_0.Vbe2.n34 0.00992001
R6556 bgr_0.Vbe2.n53 bgr_0.Vbe2.n40 0.00992001
R6557 bgr_0.Vbe2.n55 bgr_0.Vbe2.n43 0.00992001
R6558 bgr_0.Vbe2.n52 bgr_0.Vbe2.n44 0.00992001
R6559 bgr_0.Vbe2.n41 bgr_0.Vbe2.n3 0.00992001
R6560 bgr_0.Vbe2.n55 bgr_0.Vbe2.n44 0.00992001
R6561 bgr_0.Vbe2.n52 bgr_0.Vbe2.n41 0.00992001
R6562 bgr_0.Vbe2.n40 bgr_0.Vbe2.n39 0.00992001
R6563 bgr_0.Vbe2.n57 bgr_0.Vbe2.n34 0.00992001
R6564 bgr_0.Vbe2.n53 bgr_0.Vbe2.n43 0.00992001
R6565 bgr_0.Vbe2.n125 bgr_0.Vbe2.n124 0.00889286
R6566 bgr_0.Vbe2.n89 bgr_0.Vbe2.n88 0.00817857
R6567 bgr_0.Vbe2.n60 bgr_0.Vbe2.n58 0.00817857
R6568 bgr_0.Vbe2.n112 bgr_0.Vbe2.n111 0.00817857
R6569 bgr_0.Vbe2.n140 bgr_0.Vbe2.n139 0.00817857
R6570 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.t0 384.967
R6571 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t5 369.534
R6572 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t20 369.534
R6573 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t23 369.534
R6574 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t15 369.534
R6575 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t17 369.534
R6576 bgr_0.NFET_GATE_10uA.t0 bgr_0.NFET_GATE_10uA.n18 369.534
R6577 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n20 365.491
R6578 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.t12 192.8
R6579 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.t11 192.8
R6580 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t19 192.8
R6581 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t6 192.8
R6582 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t14 192.8
R6583 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t13 192.8
R6584 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.t21 192.8
R6585 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.t7 192.8
R6586 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.t16 192.8
R6587 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.t22 192.8
R6588 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t9 192.8
R6589 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.t10 192.8
R6590 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.t18 192.8
R6591 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.t8 192.8
R6592 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.n11 176.733
R6593 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.n10 176.733
R6594 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.n4 176.733
R6595 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.n5 176.733
R6596 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.n2 176.733
R6597 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.n1 176.733
R6598 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.n17 176.733
R6599 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.n16 176.733
R6600 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n13 169.852
R6601 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n8 169.852
R6602 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n14 166.133
R6603 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.n0 126.877
R6604 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n12 56.2338
R6605 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n9 56.2338
R6606 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n7 56.2338
R6607 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n6 56.2338
R6608 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n3 56.2338
R6609 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.n15 56.2338
R6610 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t3 39.4005
R6611 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t2 39.4005
R6612 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n19 28.6755
R6613 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t4 24.0005
R6614 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t1 24.0005
R6615 bgr_0.V_mir2.n20 bgr_0.V_mir2.n19 325.473
R6616 bgr_0.V_mir2.n13 bgr_0.V_mir2.n12 325.473
R6617 bgr_0.V_mir2.n8 bgr_0.V_mir2.n7 325.473
R6618 bgr_0.V_mir2.n16 bgr_0.V_mir2.t22 310.488
R6619 bgr_0.V_mir2.n9 bgr_0.V_mir2.t17 310.488
R6620 bgr_0.V_mir2.n4 bgr_0.V_mir2.t20 310.488
R6621 bgr_0.V_mir2.n2 bgr_0.V_mir2.t0 278.312
R6622 bgr_0.V_mir2.n2 bgr_0.V_mir2.n1 228.939
R6623 bgr_0.V_mir2.n3 bgr_0.V_mir2.n0 224.439
R6624 bgr_0.V_mir2.n18 bgr_0.V_mir2.t11 184.097
R6625 bgr_0.V_mir2.n11 bgr_0.V_mir2.t7 184.097
R6626 bgr_0.V_mir2.n6 bgr_0.V_mir2.t9 184.097
R6627 bgr_0.V_mir2.n17 bgr_0.V_mir2.n16 167.094
R6628 bgr_0.V_mir2.n10 bgr_0.V_mir2.n9 167.094
R6629 bgr_0.V_mir2.n5 bgr_0.V_mir2.n4 167.094
R6630 bgr_0.V_mir2.n13 bgr_0.V_mir2.n11 152
R6631 bgr_0.V_mir2.n8 bgr_0.V_mir2.n6 152
R6632 bgr_0.V_mir2.n19 bgr_0.V_mir2.n18 152
R6633 bgr_0.V_mir2.n16 bgr_0.V_mir2.t19 120.501
R6634 bgr_0.V_mir2.n17 bgr_0.V_mir2.t13 120.501
R6635 bgr_0.V_mir2.n9 bgr_0.V_mir2.t21 120.501
R6636 bgr_0.V_mir2.n10 bgr_0.V_mir2.t15 120.501
R6637 bgr_0.V_mir2.n4 bgr_0.V_mir2.t18 120.501
R6638 bgr_0.V_mir2.n5 bgr_0.V_mir2.t5 120.501
R6639 bgr_0.V_mir2.n1 bgr_0.V_mir2.t3 48.0005
R6640 bgr_0.V_mir2.n1 bgr_0.V_mir2.t4 48.0005
R6641 bgr_0.V_mir2.n0 bgr_0.V_mir2.t2 48.0005
R6642 bgr_0.V_mir2.n0 bgr_0.V_mir2.t1 48.0005
R6643 bgr_0.V_mir2.n18 bgr_0.V_mir2.n17 40.7027
R6644 bgr_0.V_mir2.n11 bgr_0.V_mir2.n10 40.7027
R6645 bgr_0.V_mir2.n6 bgr_0.V_mir2.n5 40.7027
R6646 bgr_0.V_mir2.n12 bgr_0.V_mir2.t16 39.4005
R6647 bgr_0.V_mir2.n12 bgr_0.V_mir2.t8 39.4005
R6648 bgr_0.V_mir2.n7 bgr_0.V_mir2.t6 39.4005
R6649 bgr_0.V_mir2.n7 bgr_0.V_mir2.t10 39.4005
R6650 bgr_0.V_mir2.t14 bgr_0.V_mir2.n20 39.4005
R6651 bgr_0.V_mir2.n20 bgr_0.V_mir2.t12 39.4005
R6652 bgr_0.V_mir2.n14 bgr_0.V_mir2.n13 15.8005
R6653 bgr_0.V_mir2.n14 bgr_0.V_mir2.n8 15.8005
R6654 bgr_0.V_mir2.n19 bgr_0.V_mir2.n15 9.3005
R6655 bgr_0.V_mir2.n3 bgr_0.V_mir2.n2 5.8755
R6656 bgr_0.V_mir2.n15 bgr_0.V_mir2.n14 4.5005
R6657 bgr_0.V_mir2.n15 bgr_0.V_mir2.n3 0.78175
R6658 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 688.859
R6659 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 514.134
R6660 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 323.491
R6661 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 322.692
R6662 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 270.591
R6663 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 270.591
R6664 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 270.591
R6665 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 270.591
R6666 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 233.374
R6667 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 233.374
R6668 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 233.374
R6669 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 233.374
R6670 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 208.838
R6671 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 197.964
R6672 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 174.726
R6673 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 174.726
R6674 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 174.726
R6675 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 174.726
R6676 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 169.216
R6677 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 169.216
R6678 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 169.216
R6679 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 129.24
R6680 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 129.24
R6681 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 129.24
R6682 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 129.24
R6683 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 128.534
R6684 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 128.534
R6685 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 16.8443
R6686 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 13.1338
R6687 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 13.1338
R6688 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 13.1338
R6689 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 13.1338
R6690 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 13.1338
R6691 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 13.1338
R6692 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 4.3755
R6693 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 4.3755
R6694 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 3.688
R6695 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 3.2505
R6696 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 3.1255
R6697 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 1.2755
R6698 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 1.2755
R6699 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 0.8005
R6700 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 632.186
R6701 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 630.264
R6702 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 630.264
R6703 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 630.264
R6704 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 628.003
R6705 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 628.003
R6706 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 626.753
R6707 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 626.753
R6708 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 625.756
R6709 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 622.231
R6710 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 78.8005
R6711 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 78.8005
R6712 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 78.8005
R6713 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 78.8005
R6714 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 78.8005
R6715 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 78.8005
R6716 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 78.8005
R6717 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 78.8005
R6718 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 78.8005
R6719 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 78.8005
R6720 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 78.8005
R6721 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 78.8005
R6722 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 78.8005
R6723 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 78.8005
R6724 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 78.8005
R6725 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 78.8005
R6726 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 78.8005
R6727 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 78.8005
R6728 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 78.8005
R6729 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 78.8005
R6730 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 7.94147
R6731 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 6.188
R6732 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n27 630.264
R6733 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n2 627.316
R6734 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n4 626.784
R6735 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n3 626.784
R6736 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n26 626.784
R6737 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate.n24 585
R6738 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.t17 289.2
R6739 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.t29 289.2
R6740 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.n21 176.733
R6741 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.n5 176.733
R6742 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.n6 176.733
R6743 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.n7 176.733
R6744 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.n8 176.733
R6745 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.n9 176.733
R6746 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.n10 176.733
R6747 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.n11 176.733
R6748 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.n12 176.733
R6749 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.n13 176.733
R6750 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.n14 176.733
R6751 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.n15 176.733
R6752 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.n16 176.733
R6753 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.n17 176.733
R6754 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.n18 176.733
R6755 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.n19 176.733
R6756 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n23 162.214
R6757 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n28 135.81
R6758 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n1 124.484
R6759 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.t14 112.468
R6760 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.t27 112.468
R6761 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.t20 112.468
R6762 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.t26 112.468
R6763 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.t19 112.468
R6764 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.t31 112.468
R6765 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.t22 112.468
R6766 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.t33 112.468
R6767 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.t24 112.468
R6768 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.t15 112.468
R6769 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.t28 112.468
R6770 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.t18 112.468
R6771 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.t25 112.468
R6772 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.t16 112.468
R6773 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.t30 112.468
R6774 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.t21 112.468
R6775 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.t32 112.468
R6776 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.t23 112.468
R6777 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.t7 78.8005
R6778 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.t8 78.8005
R6779 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.t3 78.8005
R6780 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.t0 78.8005
R6781 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.t10 78.8005
R6782 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.t11 78.8005
R6783 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate.t9 78.8005
R6784 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate.t13 78.8005
R6785 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t12 78.8005
R6786 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t1 78.8005
R6787 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.t2 78.8005
R6788 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.t4 78.8005
R6789 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.n22 49.8072
R6790 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.n20 49.8072
R6791 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n25 41.7838
R6792 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate 39.8442
R6793 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.t6 24.0005
R6794 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.t5 24.0005
R6795 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n0 2.313
R6796 two_stage_opamp_dummy_magic_0.X.n49 two_stage_opamp_dummy_magic_0.X.t26 1172.87
R6797 two_stage_opamp_dummy_magic_0.X.n43 two_stage_opamp_dummy_magic_0.X.t35 1172.87
R6798 two_stage_opamp_dummy_magic_0.X.n50 two_stage_opamp_dummy_magic_0.X.t45 996.134
R6799 two_stage_opamp_dummy_magic_0.X.n49 two_stage_opamp_dummy_magic_0.X.t34 996.134
R6800 two_stage_opamp_dummy_magic_0.X.n43 two_stage_opamp_dummy_magic_0.X.t48 996.134
R6801 two_stage_opamp_dummy_magic_0.X.n44 two_stage_opamp_dummy_magic_0.X.t38 996.134
R6802 two_stage_opamp_dummy_magic_0.X.n45 two_stage_opamp_dummy_magic_0.X.t51 996.134
R6803 two_stage_opamp_dummy_magic_0.X.n46 two_stage_opamp_dummy_magic_0.X.t27 996.134
R6804 two_stage_opamp_dummy_magic_0.X.n47 two_stage_opamp_dummy_magic_0.X.t43 996.134
R6805 two_stage_opamp_dummy_magic_0.X.n48 two_stage_opamp_dummy_magic_0.X.t30 996.134
R6806 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.t29 690.867
R6807 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.t40 690.867
R6808 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.t54 530.201
R6809 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.t33 530.201
R6810 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.t39 514.134
R6811 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.t49 514.134
R6812 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.t36 514.134
R6813 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.t46 514.134
R6814 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.t31 514.134
R6815 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.t53 514.134
R6816 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.t41 514.134
R6817 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.t52 514.134
R6818 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.t37 353.467
R6819 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.t50 353.467
R6820 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.t25 353.467
R6821 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.t42 353.467
R6822 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.t28 353.467
R6823 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.t44 353.467
R6824 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.t32 353.467
R6825 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.t47 353.467
R6826 two_stage_opamp_dummy_magic_0.X.n50 two_stage_opamp_dummy_magic_0.X.n49 176.733
R6827 two_stage_opamp_dummy_magic_0.X.n44 two_stage_opamp_dummy_magic_0.X.n43 176.733
R6828 two_stage_opamp_dummy_magic_0.X.n45 two_stage_opamp_dummy_magic_0.X.n44 176.733
R6829 two_stage_opamp_dummy_magic_0.X.n46 two_stage_opamp_dummy_magic_0.X.n45 176.733
R6830 two_stage_opamp_dummy_magic_0.X.n47 two_stage_opamp_dummy_magic_0.X.n46 176.733
R6831 two_stage_opamp_dummy_magic_0.X.n48 two_stage_opamp_dummy_magic_0.X.n47 176.733
R6832 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.n29 176.733
R6833 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.n28 176.733
R6834 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.n27 176.733
R6835 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.n26 176.733
R6836 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.n25 176.733
R6837 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.n24 176.733
R6838 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.n38 176.733
R6839 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.n37 176.733
R6840 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.n36 176.733
R6841 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.n35 176.733
R6842 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.n34 176.733
R6843 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.n33 176.733
R6844 two_stage_opamp_dummy_magic_0.X.n52 two_stage_opamp_dummy_magic_0.X.n51 166.436
R6845 two_stage_opamp_dummy_magic_0.X.n41 two_stage_opamp_dummy_magic_0.X.n31 161.875
R6846 two_stage_opamp_dummy_magic_0.X.n41 two_stage_opamp_dummy_magic_0.X.n40 161.686
R6847 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.n0 160.427
R6848 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.n7 159.802
R6849 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.n5 159.802
R6850 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.n3 159.802
R6851 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.n1 159.802
R6852 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n9 155.302
R6853 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.n13 114.689
R6854 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.n12 114.689
R6855 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n18 114.126
R6856 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.n16 114.126
R6857 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.n14 114.126
R6858 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.n11 109.626
R6859 two_stage_opamp_dummy_magic_0.X.n51 two_stage_opamp_dummy_magic_0.X.n50 51.9494
R6860 two_stage_opamp_dummy_magic_0.X.n51 two_stage_opamp_dummy_magic_0.X.n48 51.9494
R6861 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.n30 51.9494
R6862 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.n23 51.9494
R6863 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n39 51.9494
R6864 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n32 51.9494
R6865 two_stage_opamp_dummy_magic_0.X.t11 two_stage_opamp_dummy_magic_0.X.n52 49.3036
R6866 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.t9 16.0005
R6867 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.t24 16.0005
R6868 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.t4 16.0005
R6869 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.t23 16.0005
R6870 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.t15 16.0005
R6871 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.t3 16.0005
R6872 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.t8 16.0005
R6873 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.t22 16.0005
R6874 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.t21 16.0005
R6875 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.t5 16.0005
R6876 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t19 16.0005
R6877 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t10 16.0005
R6878 two_stage_opamp_dummy_magic_0.X.n52 two_stage_opamp_dummy_magic_0.X.n42 15.7193
R6879 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.t13 11.2576
R6880 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.t17 11.2576
R6881 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.t6 11.2576
R6882 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.t0 11.2576
R6883 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.t16 11.2576
R6884 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.t12 11.2576
R6885 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.t18 11.2576
R6886 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.t1 11.2576
R6887 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t2 11.2576
R6888 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t20 11.2576
R6889 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t14 11.2576
R6890 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t7 11.2576
R6891 two_stage_opamp_dummy_magic_0.X.n42 two_stage_opamp_dummy_magic_0.X.n22 10.188
R6892 two_stage_opamp_dummy_magic_0.X.n42 two_stage_opamp_dummy_magic_0.X.n41 6.188
R6893 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n8 5.1255
R6894 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.n20 4.5005
R6895 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.n2 0.6255
R6896 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.n4 0.6255
R6897 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.n6 0.6255
R6898 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.n15 0.563
R6899 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n17 0.563
R6900 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.n19 0.563
R6901 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.n10 0.5005
R6902 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.n21 0.438
R6903 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 344.837
R6904 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 344.274
R6905 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 292.5
R6906 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 206.052
R6907 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 205.488
R6908 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 205.488
R6909 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 205.488
R6910 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 205.488
R6911 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 122.504
R6912 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 71.2813
R6913 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 52.4067
R6914 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 52.3363
R6915 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 39.4005
R6916 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 39.4005
R6917 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 39.4005
R6918 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 39.4005
R6919 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 39.4005
R6920 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 39.4005
R6921 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 19.7005
R6922 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 19.7005
R6923 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 19.7005
R6924 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 19.7005
R6925 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 19.7005
R6926 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 19.7005
R6927 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 19.7005
R6928 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 19.7005
R6929 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 19.7005
R6930 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 19.7005
R6931 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 6.09425
R6932 bgr_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 1.15675
R6933 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 0.563
R6934 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 0.563
R6935 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 0.563
R6936 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t25 369.534
R6937 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t24 369.534
R6938 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t15 369.534
R6939 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t11 369.534
R6940 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t17 369.534
R6941 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t16 369.534
R6942 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n6 341.397
R6943 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n9 339.272
R6944 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n7 339.272
R6945 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n12 334.772
R6946 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.t21 238.322
R6947 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.t13 238.322
R6948 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.t3 194.895
R6949 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t18 192.8
R6950 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t10 192.8
R6951 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.t14 192.8
R6952 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.t22 192.8
R6953 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t28 192.8
R6954 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t19 192.8
R6955 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.t26 192.8
R6956 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.t12 192.8
R6957 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.t20 192.8
R6958 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.t27 192.8
R6959 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t29 192.8
R6960 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t23 192.8
R6961 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.n24 176.733
R6962 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.n23 176.733
R6963 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.n18 176.733
R6964 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.n19 176.733
R6965 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.n20 176.733
R6966 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.n21 176.733
R6967 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n2 171.321
R6968 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n15 169.394
R6969 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n5 168.166
R6970 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n26 166.071
R6971 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.t8 100.635
R6972 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n4 56.2338
R6973 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n3 56.2338
R6974 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n25 56.2338
R6975 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n22 56.2338
R6976 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n1 56.2338
R6977 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n0 56.2338
R6978 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t6 39.4005
R6979 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t5 39.4005
R6980 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t2 39.4005
R6981 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t9 39.4005
R6982 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t0 39.4005
R6983 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t4 39.4005
R6984 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t1 39.4005
R6985 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t7 39.4005
R6986 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n16 26.9067
R6987 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.n13 5.15675
R6988 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n11 4.5005
R6989 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n14 4.188
R6990 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n17 3.03175
R6991 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n8 2.1255
R6992 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.n10 2.1255
R6993 two_stage_opamp_dummy_magic_0.Y.n43 two_stage_opamp_dummy_magic_0.Y.t52 1172.87
R6994 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.t27 1172.87
R6995 two_stage_opamp_dummy_magic_0.Y.n48 two_stage_opamp_dummy_magic_0.Y.t44 996.134
R6996 two_stage_opamp_dummy_magic_0.Y.n47 two_stage_opamp_dummy_magic_0.Y.t32 996.134
R6997 two_stage_opamp_dummy_magic_0.Y.n46 two_stage_opamp_dummy_magic_0.Y.t49 996.134
R6998 two_stage_opamp_dummy_magic_0.Y.n45 two_stage_opamp_dummy_magic_0.Y.t37 996.134
R6999 two_stage_opamp_dummy_magic_0.Y.n44 two_stage_opamp_dummy_magic_0.Y.t48 996.134
R7000 two_stage_opamp_dummy_magic_0.Y.n43 two_stage_opamp_dummy_magic_0.Y.t36 996.134
R7001 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.t42 996.134
R7002 two_stage_opamp_dummy_magic_0.Y.n42 two_stage_opamp_dummy_magic_0.Y.t29 996.134
R7003 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.t25 690.867
R7004 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.t30 690.867
R7005 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.t51 530.201
R7006 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.t26 530.201
R7007 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.t39 514.134
R7008 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.t53 514.134
R7009 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.t40 514.134
R7010 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.t54 514.134
R7011 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.t38 514.134
R7012 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.t50 514.134
R7013 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.t33 514.134
R7014 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.t45 514.134
R7015 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.t34 353.467
R7016 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.t41 353.467
R7017 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.t28 353.467
R7018 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.t43 353.467
R7019 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.t31 353.467
R7020 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.t47 353.467
R7021 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.t35 353.467
R7022 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.t46 353.467
R7023 two_stage_opamp_dummy_magic_0.Y.n48 two_stage_opamp_dummy_magic_0.Y.n47 176.733
R7024 two_stage_opamp_dummy_magic_0.Y.n47 two_stage_opamp_dummy_magic_0.Y.n46 176.733
R7025 two_stage_opamp_dummy_magic_0.Y.n46 two_stage_opamp_dummy_magic_0.Y.n45 176.733
R7026 two_stage_opamp_dummy_magic_0.Y.n45 two_stage_opamp_dummy_magic_0.Y.n44 176.733
R7027 two_stage_opamp_dummy_magic_0.Y.n44 two_stage_opamp_dummy_magic_0.Y.n43 176.733
R7028 two_stage_opamp_dummy_magic_0.Y.n42 two_stage_opamp_dummy_magic_0.Y.n41 176.733
R7029 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.n22 176.733
R7030 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.n23 176.733
R7031 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.n24 176.733
R7032 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.n25 176.733
R7033 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.n26 176.733
R7034 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.n27 176.733
R7035 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.n31 176.733
R7036 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.n32 176.733
R7037 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.n33 176.733
R7038 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.n34 176.733
R7039 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.n35 176.733
R7040 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.n36 176.733
R7041 two_stage_opamp_dummy_magic_0.Y.n50 two_stage_opamp_dummy_magic_0.Y.n49 166.375
R7042 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n30 161.875
R7043 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n39 161.686
R7044 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.n0 160.427
R7045 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.n7 159.802
R7046 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.n5 159.802
R7047 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.n3 159.802
R7048 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.n1 159.802
R7049 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n9 155.302
R7050 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.n19 114.689
R7051 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.n12 114.689
R7052 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.n17 114.126
R7053 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.n15 114.126
R7054 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.n13 114.126
R7055 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.n11 109.626
R7056 two_stage_opamp_dummy_magic_0.Y.n49 two_stage_opamp_dummy_magic_0.Y.n48 51.9494
R7057 two_stage_opamp_dummy_magic_0.Y.n49 two_stage_opamp_dummy_magic_0.Y.n42 51.9494
R7058 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.n29 51.9494
R7059 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.n28 51.9494
R7060 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n38 51.9494
R7061 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n37 51.9494
R7062 two_stage_opamp_dummy_magic_0.Y.n50 two_stage_opamp_dummy_magic_0.Y.t11 49.2412
R7063 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.t16 16.0005
R7064 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.t22 16.0005
R7065 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.t17 16.0005
R7066 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.t2 16.0005
R7067 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.t20 16.0005
R7068 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.t15 16.0005
R7069 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.t0 16.0005
R7070 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.t1 16.0005
R7071 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.t21 16.0005
R7072 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.t19 16.0005
R7073 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t4 16.0005
R7074 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t6 16.0005
R7075 two_stage_opamp_dummy_magic_0.Y.n51 two_stage_opamp_dummy_magic_0.Y.n50 15.6567
R7076 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.t5 11.2576
R7077 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.t3 11.2576
R7078 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.t23 11.2576
R7079 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.t10 11.2576
R7080 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.t8 11.2576
R7081 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.t9 11.2576
R7082 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.t13 11.2576
R7083 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.t18 11.2576
R7084 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t12 11.2576
R7085 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t7 11.2576
R7086 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t14 11.2576
R7087 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t24 11.2576
R7088 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.Y.n51 10.313
R7089 two_stage_opamp_dummy_magic_0.Y.n51 two_stage_opamp_dummy_magic_0.Y.n40 6.063
R7090 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n8 5.1255
R7091 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.n20 4.5005
R7092 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.n2 0.6255
R7093 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.n4 0.6255
R7094 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.n6 0.6255
R7095 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.n14 0.563
R7096 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.n16 0.563
R7097 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.n18 0.563
R7098 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.Y.n10 0.5005
R7099 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.Y.n21 0.438
R7100 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 144.827
R7101 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 134.577
R7102 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 120.629
R7103 bgr_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 112.281
R7104 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 97.4009
R7105 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 96.8384
R7106 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 96.8384
R7107 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 96.8384
R7108 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 96.8384
R7109 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 24.0005
R7110 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 24.0005
R7111 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 24.0005
R7112 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 24.0005
R7113 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 8.0005
R7114 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 8.0005
R7115 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 8.0005
R7116 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 8.0005
R7117 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 8.0005
R7118 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 8.0005
R7119 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 8.0005
R7120 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 8.0005
R7121 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 8.0005
R7122 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 8.0005
R7123 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 5.84425
R7124 bgr_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 1.46925
R7125 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 0.563
R7126 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 0.563
R7127 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 0.563
R7128 bgr_0.V_mir1.n20 bgr_0.V_mir1.n19 325.473
R7129 bgr_0.V_mir1.n13 bgr_0.V_mir1.n12 325.473
R7130 bgr_0.V_mir1.n4 bgr_0.V_mir1.n3 325.473
R7131 bgr_0.V_mir1.n16 bgr_0.V_mir1.t22 310.488
R7132 bgr_0.V_mir1.n9 bgr_0.V_mir1.t21 310.488
R7133 bgr_0.V_mir1.n0 bgr_0.V_mir1.t20 310.488
R7134 bgr_0.V_mir1.n7 bgr_0.V_mir1.t15 278.312
R7135 bgr_0.V_mir1.n7 bgr_0.V_mir1.n6 228.939
R7136 bgr_0.V_mir1.n8 bgr_0.V_mir1.n5 224.439
R7137 bgr_0.V_mir1.n18 bgr_0.V_mir1.t10 184.097
R7138 bgr_0.V_mir1.n11 bgr_0.V_mir1.t0 184.097
R7139 bgr_0.V_mir1.n2 bgr_0.V_mir1.t8 184.097
R7140 bgr_0.V_mir1.n17 bgr_0.V_mir1.n16 167.094
R7141 bgr_0.V_mir1.n10 bgr_0.V_mir1.n9 167.094
R7142 bgr_0.V_mir1.n1 bgr_0.V_mir1.n0 167.094
R7143 bgr_0.V_mir1.n13 bgr_0.V_mir1.n11 152
R7144 bgr_0.V_mir1.n4 bgr_0.V_mir1.n2 152
R7145 bgr_0.V_mir1.n19 bgr_0.V_mir1.n18 152
R7146 bgr_0.V_mir1.n16 bgr_0.V_mir1.t19 120.501
R7147 bgr_0.V_mir1.n17 bgr_0.V_mir1.t2 120.501
R7148 bgr_0.V_mir1.n9 bgr_0.V_mir1.t18 120.501
R7149 bgr_0.V_mir1.n10 bgr_0.V_mir1.t4 120.501
R7150 bgr_0.V_mir1.n0 bgr_0.V_mir1.t17 120.501
R7151 bgr_0.V_mir1.n1 bgr_0.V_mir1.t6 120.501
R7152 bgr_0.V_mir1.n6 bgr_0.V_mir1.t16 48.0005
R7153 bgr_0.V_mir1.n6 bgr_0.V_mir1.t12 48.0005
R7154 bgr_0.V_mir1.n5 bgr_0.V_mir1.t13 48.0005
R7155 bgr_0.V_mir1.n5 bgr_0.V_mir1.t14 48.0005
R7156 bgr_0.V_mir1.n18 bgr_0.V_mir1.n17 40.7027
R7157 bgr_0.V_mir1.n11 bgr_0.V_mir1.n10 40.7027
R7158 bgr_0.V_mir1.n2 bgr_0.V_mir1.n1 40.7027
R7159 bgr_0.V_mir1.n12 bgr_0.V_mir1.t1 39.4005
R7160 bgr_0.V_mir1.n12 bgr_0.V_mir1.t5 39.4005
R7161 bgr_0.V_mir1.n3 bgr_0.V_mir1.t9 39.4005
R7162 bgr_0.V_mir1.n3 bgr_0.V_mir1.t7 39.4005
R7163 bgr_0.V_mir1.t11 bgr_0.V_mir1.n20 39.4005
R7164 bgr_0.V_mir1.n20 bgr_0.V_mir1.t3 39.4005
R7165 bgr_0.V_mir1.n15 bgr_0.V_mir1.n4 15.8005
R7166 bgr_0.V_mir1.n19 bgr_0.V_mir1.n15 15.8005
R7167 bgr_0.V_mir1.n14 bgr_0.V_mir1.n13 9.3005
R7168 bgr_0.V_mir1.n8 bgr_0.V_mir1.n7 5.8755
R7169 bgr_0.V_mir1.n15 bgr_0.V_mir1.n14 4.5005
R7170 bgr_0.V_mir1.n14 bgr_0.V_mir1.n8 0.78175
R7171 VOUT+.n2 VOUT+.n0 145.989
R7172 VOUT+.n8 VOUT+.n7 145.989
R7173 VOUT+.n6 VOUT+.n5 145.427
R7174 VOUT+.n4 VOUT+.n3 145.427
R7175 VOUT+.n2 VOUT+.n1 145.427
R7176 VOUT+.n10 VOUT+.n9 140.927
R7177 VOUT+.n100 VOUT+.t1 113.192
R7178 VOUT+.n97 VOUT+.n95 95.7303
R7179 VOUT+.n99 VOUT+.n98 94.6053
R7180 VOUT+.n97 VOUT+.n96 94.6053
R7181 VOUT+.n94 VOUT+.n10 20.5943
R7182 VOUT+.n94 VOUT+.n93 11.7059
R7183 VOUT+ VOUT+.n94 7.813
R7184 VOUT+.n9 VOUT+.t11 6.56717
R7185 VOUT+.n9 VOUT+.t15 6.56717
R7186 VOUT+.n7 VOUT+.t9 6.56717
R7187 VOUT+.n7 VOUT+.t6 6.56717
R7188 VOUT+.n5 VOUT+.t10 6.56717
R7189 VOUT+.n5 VOUT+.t14 6.56717
R7190 VOUT+.n3 VOUT+.t12 6.56717
R7191 VOUT+.n3 VOUT+.t16 6.56717
R7192 VOUT+.n1 VOUT+.t13 6.56717
R7193 VOUT+.n1 VOUT+.t17 6.56717
R7194 VOUT+.n0 VOUT+.t5 6.56717
R7195 VOUT+.n0 VOUT+.t18 6.56717
R7196 VOUT+.n40 VOUT+.t108 4.8295
R7197 VOUT+.n52 VOUT+.t25 4.8295
R7198 VOUT+.n49 VOUT+.t76 4.8295
R7199 VOUT+.n46 VOUT+.t113 4.8295
R7200 VOUT+.n43 VOUT+.t145 4.8295
R7201 VOUT+.n42 VOUT+.t68 4.8295
R7202 VOUT+.n66 VOUT+.t28 4.8295
R7203 VOUT+.n67 VOUT+.t77 4.8295
R7204 VOUT+.n69 VOUT+.t63 4.8295
R7205 VOUT+.n70 VOUT+.t111 4.8295
R7206 VOUT+.n72 VOUT+.t114 4.8295
R7207 VOUT+.n73 VOUT+.t99 4.8295
R7208 VOUT+.n75 VOUT+.t74 4.8295
R7209 VOUT+.n76 VOUT+.t56 4.8295
R7210 VOUT+.n78 VOUT+.t109 4.8295
R7211 VOUT+.n79 VOUT+.t92 4.8295
R7212 VOUT+.n81 VOUT+.t69 4.8295
R7213 VOUT+.n82 VOUT+.t53 4.8295
R7214 VOUT+.n84 VOUT+.t30 4.8295
R7215 VOUT+.n85 VOUT+.t153 4.8295
R7216 VOUT+.n87 VOUT+.t64 4.8295
R7217 VOUT+.n88 VOUT+.t47 4.8295
R7218 VOUT+.n11 VOUT+.t117 4.8295
R7219 VOUT+.n13 VOUT+.t72 4.8295
R7220 VOUT+.n25 VOUT+.t38 4.8295
R7221 VOUT+.n26 VOUT+.t20 4.8295
R7222 VOUT+.n28 VOUT+.t80 4.8295
R7223 VOUT+.n29 VOUT+.t61 4.8295
R7224 VOUT+.n31 VOUT+.t121 4.8295
R7225 VOUT+.n32 VOUT+.t104 4.8295
R7226 VOUT+.n34 VOUT+.t85 4.8295
R7227 VOUT+.n35 VOUT+.t67 4.8295
R7228 VOUT+.n37 VOUT+.t123 4.8295
R7229 VOUT+.n38 VOUT+.t107 4.8295
R7230 VOUT+.n90 VOUT+.t22 4.8295
R7231 VOUT+.n55 VOUT+.t33 4.806
R7232 VOUT+.n56 VOUT+.t150 4.806
R7233 VOUT+.n57 VOUT+.t51 4.806
R7234 VOUT+.n58 VOUT+.t88 4.806
R7235 VOUT+.n59 VOUT+.t125 4.806
R7236 VOUT+.n60 VOUT+.t105 4.806
R7237 VOUT+.n61 VOUT+.t140 4.806
R7238 VOUT+.n62 VOUT+.t37 4.806
R7239 VOUT+.n63 VOUT+.t156 4.806
R7240 VOUT+.n64 VOUT+.t54 4.806
R7241 VOUT+.n14 VOUT+.t73 4.806
R7242 VOUT+.n15 VOUT+.t116 4.806
R7243 VOUT+.n16 VOUT+.t65 4.806
R7244 VOUT+.n17 VOUT+.t154 4.806
R7245 VOUT+.n18 VOUT+.t106 4.806
R7246 VOUT+.n19 VOUT+.t143 4.806
R7247 VOUT+.n20 VOUT+.t96 4.806
R7248 VOUT+.n21 VOUT+.t43 4.806
R7249 VOUT+.n22 VOUT+.t87 4.806
R7250 VOUT+.n23 VOUT+.t35 4.806
R7251 VOUT+.n40 VOUT+.t70 4.5005
R7252 VOUT+.n41 VOUT+.t91 4.5005
R7253 VOUT+.n52 VOUT+.t66 4.5005
R7254 VOUT+.n53 VOUT+.t81 4.5005
R7255 VOUT+.n54 VOUT+.t44 4.5005
R7256 VOUT+.n49 VOUT+.t118 4.5005
R7257 VOUT+.n50 VOUT+.t57 4.5005
R7258 VOUT+.n51 VOUT+.t21 4.5005
R7259 VOUT+.n46 VOUT+.t151 4.5005
R7260 VOUT+.n47 VOUT+.t98 4.5005
R7261 VOUT+.n48 VOUT+.t60 4.5005
R7262 VOUT+.n43 VOUT+.t45 4.5005
R7263 VOUT+.n44 VOUT+.t136 4.5005
R7264 VOUT+.n45 VOUT+.t101 4.5005
R7265 VOUT+.n42 VOUT+.t31 4.5005
R7266 VOUT+.n65 VOUT+.t52 4.5005
R7267 VOUT+.n64 VOUT+.t155 4.5005
R7268 VOUT+.n63 VOUT+.t119 4.5005
R7269 VOUT+.n62 VOUT+.t139 4.5005
R7270 VOUT+.n61 VOUT+.t102 4.5005
R7271 VOUT+.n60 VOUT+.t62 4.5005
R7272 VOUT+.n59 VOUT+.t86 4.5005
R7273 VOUT+.n58 VOUT+.t46 4.5005
R7274 VOUT+.n57 VOUT+.t147 4.5005
R7275 VOUT+.n56 VOUT+.t110 4.5005
R7276 VOUT+.n55 VOUT+.t134 4.5005
R7277 VOUT+.n66 VOUT+.t130 4.5005
R7278 VOUT+.n68 VOUT+.t152 4.5005
R7279 VOUT+.n67 VOUT+.t115 4.5005
R7280 VOUT+.n69 VOUT+.t23 4.5005
R7281 VOUT+.n71 VOUT+.t48 4.5005
R7282 VOUT+.n70 VOUT+.t148 4.5005
R7283 VOUT+.n72 VOUT+.t79 4.5005
R7284 VOUT+.n74 VOUT+.t27 4.5005
R7285 VOUT+.n73 VOUT+.t132 4.5005
R7286 VOUT+.n75 VOUT+.t40 4.5005
R7287 VOUT+.n77 VOUT+.t128 4.5005
R7288 VOUT+.n76 VOUT+.t93 4.5005
R7289 VOUT+.n78 VOUT+.t71 4.5005
R7290 VOUT+.n80 VOUT+.t19 4.5005
R7291 VOUT+.n79 VOUT+.t126 4.5005
R7292 VOUT+.n81 VOUT+.t34 4.5005
R7293 VOUT+.n83 VOUT+.t122 4.5005
R7294 VOUT+.n82 VOUT+.t89 4.5005
R7295 VOUT+.n84 VOUT+.t135 4.5005
R7296 VOUT+.n86 VOUT+.t83 4.5005
R7297 VOUT+.n85 VOUT+.t49 4.5005
R7298 VOUT+.n87 VOUT+.t29 4.5005
R7299 VOUT+.n89 VOUT+.t120 4.5005
R7300 VOUT+.n88 VOUT+.t82 4.5005
R7301 VOUT+.n11 VOUT+.t26 4.5005
R7302 VOUT+.n12 VOUT+.t124 4.5005
R7303 VOUT+.n13 VOUT+.t39 4.5005
R7304 VOUT+.n24 VOUT+.t127 4.5005
R7305 VOUT+.n23 VOUT+.t95 4.5005
R7306 VOUT+.n22 VOUT+.t55 4.5005
R7307 VOUT+.n21 VOUT+.t144 4.5005
R7308 VOUT+.n20 VOUT+.t112 4.5005
R7309 VOUT+.n19 VOUT+.t75 4.5005
R7310 VOUT+.n18 VOUT+.t24 4.5005
R7311 VOUT+.n17 VOUT+.t131 4.5005
R7312 VOUT+.n16 VOUT+.t97 4.5005
R7313 VOUT+.n15 VOUT+.t59 4.5005
R7314 VOUT+.n14 VOUT+.t149 4.5005
R7315 VOUT+.n25 VOUT+.t142 4.5005
R7316 VOUT+.n27 VOUT+.t94 4.5005
R7317 VOUT+.n26 VOUT+.t58 4.5005
R7318 VOUT+.n28 VOUT+.t42 4.5005
R7319 VOUT+.n30 VOUT+.t133 4.5005
R7320 VOUT+.n29 VOUT+.t100 4.5005
R7321 VOUT+.n31 VOUT+.t84 4.5005
R7322 VOUT+.n33 VOUT+.t32 4.5005
R7323 VOUT+.n32 VOUT+.t137 4.5005
R7324 VOUT+.n34 VOUT+.t50 4.5005
R7325 VOUT+.n36 VOUT+.t138 4.5005
R7326 VOUT+.n35 VOUT+.t103 4.5005
R7327 VOUT+.n37 VOUT+.t90 4.5005
R7328 VOUT+.n39 VOUT+.t36 4.5005
R7329 VOUT+.n38 VOUT+.t141 4.5005
R7330 VOUT+.n90 VOUT+.t129 4.5005
R7331 VOUT+.n91 VOUT+.t78 4.5005
R7332 VOUT+.n92 VOUT+.t41 4.5005
R7333 VOUT+.n93 VOUT+.t146 4.5005
R7334 VOUT+.n10 VOUT+.n8 4.5005
R7335 VOUT+.n98 VOUT+.t8 3.42907
R7336 VOUT+.n98 VOUT+.t4 3.42907
R7337 VOUT+.n96 VOUT+.t3 3.42907
R7338 VOUT+.n96 VOUT+.t2 3.42907
R7339 VOUT+.n95 VOUT+.t0 3.42907
R7340 VOUT+.n95 VOUT+.t7 3.42907
R7341 VOUT+ VOUT+.n100 2.84425
R7342 VOUT+.n100 VOUT+.n99 2.03175
R7343 VOUT+.n99 VOUT+.n97 1.1255
R7344 VOUT+.n4 VOUT+.n2 0.563
R7345 VOUT+.n6 VOUT+.n4 0.563
R7346 VOUT+.n8 VOUT+.n6 0.563
R7347 VOUT+.n41 VOUT+.n40 0.3295
R7348 VOUT+.n54 VOUT+.n53 0.3295
R7349 VOUT+.n53 VOUT+.n52 0.3295
R7350 VOUT+.n51 VOUT+.n50 0.3295
R7351 VOUT+.n50 VOUT+.n49 0.3295
R7352 VOUT+.n48 VOUT+.n47 0.3295
R7353 VOUT+.n47 VOUT+.n46 0.3295
R7354 VOUT+.n45 VOUT+.n44 0.3295
R7355 VOUT+.n44 VOUT+.n43 0.3295
R7356 VOUT+.n65 VOUT+.n42 0.3295
R7357 VOUT+.n65 VOUT+.n64 0.3295
R7358 VOUT+.n64 VOUT+.n63 0.3295
R7359 VOUT+.n63 VOUT+.n62 0.3295
R7360 VOUT+.n62 VOUT+.n61 0.3295
R7361 VOUT+.n61 VOUT+.n60 0.3295
R7362 VOUT+.n60 VOUT+.n59 0.3295
R7363 VOUT+.n59 VOUT+.n58 0.3295
R7364 VOUT+.n58 VOUT+.n57 0.3295
R7365 VOUT+.n57 VOUT+.n56 0.3295
R7366 VOUT+.n56 VOUT+.n55 0.3295
R7367 VOUT+.n68 VOUT+.n66 0.3295
R7368 VOUT+.n68 VOUT+.n67 0.3295
R7369 VOUT+.n71 VOUT+.n69 0.3295
R7370 VOUT+.n71 VOUT+.n70 0.3295
R7371 VOUT+.n74 VOUT+.n72 0.3295
R7372 VOUT+.n74 VOUT+.n73 0.3295
R7373 VOUT+.n77 VOUT+.n75 0.3295
R7374 VOUT+.n77 VOUT+.n76 0.3295
R7375 VOUT+.n80 VOUT+.n78 0.3295
R7376 VOUT+.n80 VOUT+.n79 0.3295
R7377 VOUT+.n83 VOUT+.n81 0.3295
R7378 VOUT+.n83 VOUT+.n82 0.3295
R7379 VOUT+.n86 VOUT+.n84 0.3295
R7380 VOUT+.n86 VOUT+.n85 0.3295
R7381 VOUT+.n89 VOUT+.n87 0.3295
R7382 VOUT+.n89 VOUT+.n88 0.3295
R7383 VOUT+.n12 VOUT+.n11 0.3295
R7384 VOUT+.n24 VOUT+.n13 0.3295
R7385 VOUT+.n24 VOUT+.n23 0.3295
R7386 VOUT+.n23 VOUT+.n22 0.3295
R7387 VOUT+.n22 VOUT+.n21 0.3295
R7388 VOUT+.n21 VOUT+.n20 0.3295
R7389 VOUT+.n20 VOUT+.n19 0.3295
R7390 VOUT+.n19 VOUT+.n18 0.3295
R7391 VOUT+.n18 VOUT+.n17 0.3295
R7392 VOUT+.n17 VOUT+.n16 0.3295
R7393 VOUT+.n16 VOUT+.n15 0.3295
R7394 VOUT+.n15 VOUT+.n14 0.3295
R7395 VOUT+.n27 VOUT+.n25 0.3295
R7396 VOUT+.n27 VOUT+.n26 0.3295
R7397 VOUT+.n30 VOUT+.n28 0.3295
R7398 VOUT+.n30 VOUT+.n29 0.3295
R7399 VOUT+.n33 VOUT+.n31 0.3295
R7400 VOUT+.n33 VOUT+.n32 0.3295
R7401 VOUT+.n36 VOUT+.n34 0.3295
R7402 VOUT+.n36 VOUT+.n35 0.3295
R7403 VOUT+.n39 VOUT+.n37 0.3295
R7404 VOUT+.n39 VOUT+.n38 0.3295
R7405 VOUT+.n91 VOUT+.n90 0.3295
R7406 VOUT+.n92 VOUT+.n91 0.3295
R7407 VOUT+.n93 VOUT+.n92 0.3295
R7408 VOUT+.n59 VOUT+.n54 0.306
R7409 VOUT+.n60 VOUT+.n51 0.306
R7410 VOUT+.n61 VOUT+.n48 0.306
R7411 VOUT+.n62 VOUT+.n45 0.306
R7412 VOUT+.n65 VOUT+.n41 0.2825
R7413 VOUT+.n68 VOUT+.n65 0.2825
R7414 VOUT+.n71 VOUT+.n68 0.2825
R7415 VOUT+.n74 VOUT+.n71 0.2825
R7416 VOUT+.n77 VOUT+.n74 0.2825
R7417 VOUT+.n80 VOUT+.n77 0.2825
R7418 VOUT+.n83 VOUT+.n80 0.2825
R7419 VOUT+.n86 VOUT+.n83 0.2825
R7420 VOUT+.n89 VOUT+.n86 0.2825
R7421 VOUT+.n24 VOUT+.n12 0.2825
R7422 VOUT+.n27 VOUT+.n24 0.2825
R7423 VOUT+.n30 VOUT+.n27 0.2825
R7424 VOUT+.n33 VOUT+.n30 0.2825
R7425 VOUT+.n36 VOUT+.n33 0.2825
R7426 VOUT+.n39 VOUT+.n36 0.2825
R7427 VOUT+.n91 VOUT+.n39 0.2825
R7428 VOUT+.n91 VOUT+.n89 0.2825
R7429 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 49.2006
R7430 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 0.1603
R7431 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 0.1603
R7432 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 0.1603
R7433 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 0.1603
R7434 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 0.1603
R7435 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 0.1603
R7436 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 0.1603
R7437 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 0.1603
R7438 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 0.1603
R7439 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 0.1603
R7440 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 0.1603
R7441 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 0.1603
R7442 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 0.1603
R7443 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 0.1603
R7444 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 0.1603
R7445 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 0.1603
R7446 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 0.1603
R7447 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 0.1603
R7448 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 0.1603
R7449 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 0.1603
R7450 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 0.1603
R7451 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 0.1603
R7452 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 0.1603
R7453 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 0.1603
R7454 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 0.1603
R7455 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 0.1603
R7456 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 0.1603
R7457 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 0.1603
R7458 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 0.1603
R7459 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 0.1603
R7460 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 0.1603
R7461 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 0.1603
R7462 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 0.1603
R7463 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 0.1603
R7464 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 0.1603
R7465 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 0.1603
R7466 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 0.1603
R7467 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 0.1603
R7468 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 0.1603
R7469 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 0.1603
R7470 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 0.1603
R7471 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 0.1603
R7472 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 0.1603
R7473 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 0.1603
R7474 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 0.1603
R7475 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 0.1603
R7476 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 0.1603
R7477 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 0.1603
R7478 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 0.1603
R7479 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 0.1603
R7480 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 0.1603
R7481 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 0.1603
R7482 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 0.1603
R7483 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 0.1603
R7484 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 0.1603
R7485 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 0.1603
R7486 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 0.1603
R7487 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 0.1603
R7488 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 0.159278
R7489 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 0.159278
R7490 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 0.159278
R7491 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 0.159278
R7492 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 0.159278
R7493 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 0.159278
R7494 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 0.159278
R7495 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 0.159278
R7496 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 0.159278
R7497 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 0.159278
R7498 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 0.159278
R7499 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 0.159278
R7500 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 0.159278
R7501 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 0.159278
R7502 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 0.159278
R7503 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 0.159278
R7504 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 0.159278
R7505 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 0.159278
R7506 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 0.159278
R7507 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 0.159278
R7508 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 0.159278
R7509 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 0.159278
R7510 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 0.159278
R7511 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 0.159278
R7512 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 0.159278
R7513 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 0.159278
R7514 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 0.159278
R7515 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 0.137822
R7516 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 0.1368
R7517 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 0.1368
R7518 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 0.1368
R7519 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 0.1368
R7520 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 0.1368
R7521 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 0.1368
R7522 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 0.1368
R7523 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 0.1368
R7524 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 0.1368
R7525 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 0.1368
R7526 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 0.1368
R7527 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 0.1368
R7528 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 0.1368
R7529 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 0.1368
R7530 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 0.1368
R7531 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 0.1368
R7532 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 0.1368
R7533 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 0.1368
R7534 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 0.1368
R7535 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 0.1368
R7536 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 0.1368
R7537 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 0.1368
R7538 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 0.1368
R7539 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 0.1368
R7540 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 0.1368
R7541 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 0.1368
R7542 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 0.1368
R7543 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 0.1368
R7544 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 0.1368
R7545 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 0.1368
R7546 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 0.1368
R7547 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 0.114322
R7548 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 0.1133
R7549 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 0.1133
R7550 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 0.1133
R7551 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 0.1133
R7552 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 0.1133
R7553 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 0.1133
R7554 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 0.1133
R7555 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 0.1133
R7556 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 0.1133
R7557 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 0.1133
R7558 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 0.1133
R7559 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 0.1133
R7560 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 0.1133
R7561 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 0.1133
R7562 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 0.1133
R7563 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 0.1133
R7564 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 0.1133
R7565 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 0.1133
R7566 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 0.1133
R7567 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 0.00152174
R7568 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 0.00152174
R7569 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 0.00152174
R7570 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 0.00152174
R7571 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 0.00152174
R7572 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 0.00152174
R7573 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 0.00152174
R7574 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 0.00152174
R7575 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 0.00152174
R7576 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 0.00152174
R7577 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 0.00152174
R7578 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 0.00152174
R7579 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 0.00152174
R7580 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 0.00152174
R7581 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 0.00152174
R7582 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 0.00152174
R7583 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 0.00152174
R7584 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 0.00152174
R7585 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 0.00152174
R7586 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 0.00152174
R7587 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 0.00152174
R7588 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 0.00152174
R7589 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 0.00152174
R7590 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 0.00152174
R7591 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 0.00152174
R7592 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 0.00152174
R7593 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 0.00152174
R7594 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 0.00152174
R7595 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 0.00152174
R7596 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 0.00152174
R7597 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 0.00152174
R7598 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 0.00152174
R7599 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 0.00152174
R7600 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 0.00152174
R7601 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 0.00152174
R7602 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 0.00152174
R7603 bgr_0.START_UP_NFET1 bgr_0.START_UP_NFET1.t0 141.653
R7604 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 525.38
R7605 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 525.38
R7606 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 366.856
R7607 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 366.856
R7608 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 281.168
R7609 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 281.168
R7610 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 281.168
R7611 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 281.168
R7612 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 244.214
R7613 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 244.214
R7614 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 166.03
R7615 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 166.03
R7616 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 117.849
R7617 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 117.849
R7618 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 85.6894
R7619 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 85.6894
R7620 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 39.5005
R7621 a_5750_2946.t0 a_5750_2946.t1 169.905
R7622 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n16 4020
R7623 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n17 4020
R7624 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n17 4020
R7625 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n16 4020
R7626 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.t13 660.109
R7627 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.t10 660.109
R7628 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.n14 428.8
R7629 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.n15 428.8
R7630 two_stage_opamp_dummy_magic_0.VD3.t14 two_stage_opamp_dummy_magic_0.VD3.n16 239.915
R7631 two_stage_opamp_dummy_magic_0.VD3.t11 two_stage_opamp_dummy_magic_0.VD3.n17 239.915
R7632 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.n19 230.4
R7633 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.n21 230.4
R7634 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.n14 198.4
R7635 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.n15 198.4
R7636 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.n11 160.428
R7637 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n7 160.427
R7638 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.n0 160.427
R7639 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.n32 160.053
R7640 two_stage_opamp_dummy_magic_0.VD3.n31 two_stage_opamp_dummy_magic_0.VD3.n30 159.803
R7641 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.n12 159.803
R7642 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.n5 159.802
R7643 two_stage_opamp_dummy_magic_0.VD3.n4 two_stage_opamp_dummy_magic_0.VD3.n3 159.802
R7644 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.n1 159.802
R7645 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.n9 155.302
R7646 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.t12 155.125
R7647 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.t15 155.125
R7648 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.n27 146.002
R7649 two_stage_opamp_dummy_magic_0.VD3.t26 two_stage_opamp_dummy_magic_0.VD3.t14 98.2764
R7650 two_stage_opamp_dummy_magic_0.VD3.t7 two_stage_opamp_dummy_magic_0.VD3.t26 98.2764
R7651 two_stage_opamp_dummy_magic_0.VD3.t0 two_stage_opamp_dummy_magic_0.VD3.t7 98.2764
R7652 two_stage_opamp_dummy_magic_0.VD3.t24 two_stage_opamp_dummy_magic_0.VD3.t0 98.2764
R7653 two_stage_opamp_dummy_magic_0.VD3.t17 two_stage_opamp_dummy_magic_0.VD3.t24 98.2764
R7654 two_stage_opamp_dummy_magic_0.VD3.t28 two_stage_opamp_dummy_magic_0.VD3.t2 98.2764
R7655 two_stage_opamp_dummy_magic_0.VD3.t2 two_stage_opamp_dummy_magic_0.VD3.t4 98.2764
R7656 two_stage_opamp_dummy_magic_0.VD3.t4 two_stage_opamp_dummy_magic_0.VD3.t33 98.2764
R7657 two_stage_opamp_dummy_magic_0.VD3.t33 two_stage_opamp_dummy_magic_0.VD3.t22 98.2764
R7658 two_stage_opamp_dummy_magic_0.VD3.t22 two_stage_opamp_dummy_magic_0.VD3.t11 98.2764
R7659 two_stage_opamp_dummy_magic_0.VD3.n16 two_stage_opamp_dummy_magic_0.VD3.n14 92.5005
R7660 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.n25 92.5005
R7661 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n24 92.5005
R7662 two_stage_opamp_dummy_magic_0.VD3.n17 two_stage_opamp_dummy_magic_0.VD3.n15 92.5005
R7663 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n22 92.5005
R7664 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.n23 92.5005
R7665 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.t17 49.1384
R7666 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.t28 49.1384
R7667 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.n20 21.3338
R7668 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.n18 21.3338
R7669 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.n26 19.2005
R7670 two_stage_opamp_dummy_magic_0.VD3.n29 two_stage_opamp_dummy_magic_0.VD3.n28 13.8005
R7671 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.t3 11.2576
R7672 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.t5 11.2576
R7673 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.t19 11.2576
R7674 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.t21 11.2576
R7675 two_stage_opamp_dummy_magic_0.VD3.n7 two_stage_opamp_dummy_magic_0.VD3.t6 11.2576
R7676 two_stage_opamp_dummy_magic_0.VD3.n7 two_stage_opamp_dummy_magic_0.VD3.t31 11.2576
R7677 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.t36 11.2576
R7678 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.t35 11.2576
R7679 two_stage_opamp_dummy_magic_0.VD3.n3 two_stage_opamp_dummy_magic_0.VD3.t37 11.2576
R7680 two_stage_opamp_dummy_magic_0.VD3.n3 two_stage_opamp_dummy_magic_0.VD3.t9 11.2576
R7681 two_stage_opamp_dummy_magic_0.VD3.n1 two_stage_opamp_dummy_magic_0.VD3.t20 11.2576
R7682 two_stage_opamp_dummy_magic_0.VD3.n1 two_stage_opamp_dummy_magic_0.VD3.t16 11.2576
R7683 two_stage_opamp_dummy_magic_0.VD3.n0 two_stage_opamp_dummy_magic_0.VD3.t32 11.2576
R7684 two_stage_opamp_dummy_magic_0.VD3.n0 two_stage_opamp_dummy_magic_0.VD3.t30 11.2576
R7685 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.t34 11.2576
R7686 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.t23 11.2576
R7687 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.t1 11.2576
R7688 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.t25 11.2576
R7689 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.t27 11.2576
R7690 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.t8 11.2576
R7691 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.t18 11.2576
R7692 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.t29 11.2576
R7693 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.VD3.n33 5.40675
R7694 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.n8 4.5005
R7695 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.VD3.n10 0.78175
R7696 two_stage_opamp_dummy_magic_0.VD3.n4 two_stage_opamp_dummy_magic_0.VD3.n2 0.6255
R7697 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.n4 0.6255
R7698 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n6 0.6255
R7699 two_stage_opamp_dummy_magic_0.VD3.n31 two_stage_opamp_dummy_magic_0.VD3.n29 0.6255
R7700 two_stage_opamp_dummy_magic_0.VD3.n29 two_stage_opamp_dummy_magic_0.VD3.n13 0.6255
R7701 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.n31 0.2505
R7702 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 628.034
R7703 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 626.784
R7704 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 626.784
R7705 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 289.2
R7706 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 289.2
R7707 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 228.252
R7708 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 212.733
R7709 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 212.733
R7710 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 176.733
R7711 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 176.733
R7712 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 176.733
R7713 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 176.733
R7714 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 176.733
R7715 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 152
R7716 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 152
R7717 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 112.468
R7718 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 112.468
R7719 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 112.468
R7720 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 112.468
R7721 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 112.468
R7722 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 112.468
R7723 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 112.468
R7724 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 112.468
R7725 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 78.8005
R7726 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 78.8005
R7727 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 78.8005
R7728 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 78.8005
R7729 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 78.8005
R7730 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 78.8005
R7731 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 48.0005
R7732 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 48.0005
R7733 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 48.0005
R7734 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 48.0005
R7735 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 48.0005
R7736 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 48.0005
R7737 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 45.5227
R7738 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 45.5227
R7739 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 45.5227
R7740 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 45.5227
R7741 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 33.8443
R7742 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 14.2693
R7743 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 14.2693
R7744 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 1.2505
R7745 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 1.2505
R7746 bgr_0.V_p_2.n0 bgr_0.V_p_2.n2 229.562
R7747 bgr_0.V_p_2.n1 bgr_0.V_p_2.n5 228.939
R7748 bgr_0.V_p_2.n0 bgr_0.V_p_2.n4 228.939
R7749 bgr_0.V_p_2.n0 bgr_0.V_p_2.n3 228.939
R7750 bgr_0.V_p_2.n6 bgr_0.V_p_2.n1 228.938
R7751 bgr_0.V_p_2.n1 bgr_0.V_p_2.t9 98.2279
R7752 bgr_0.V_p_2.n5 bgr_0.V_p_2.t0 48.0005
R7753 bgr_0.V_p_2.n5 bgr_0.V_p_2.t4 48.0005
R7754 bgr_0.V_p_2.n4 bgr_0.V_p_2.t1 48.0005
R7755 bgr_0.V_p_2.n4 bgr_0.V_p_2.t10 48.0005
R7756 bgr_0.V_p_2.n3 bgr_0.V_p_2.t7 48.0005
R7757 bgr_0.V_p_2.n3 bgr_0.V_p_2.t3 48.0005
R7758 bgr_0.V_p_2.n2 bgr_0.V_p_2.t2 48.0005
R7759 bgr_0.V_p_2.n2 bgr_0.V_p_2.t8 48.0005
R7760 bgr_0.V_p_2.t5 bgr_0.V_p_2.n6 48.0005
R7761 bgr_0.V_p_2.n6 bgr_0.V_p_2.t6 48.0005
R7762 bgr_0.V_p_2.n1 bgr_0.V_p_2.n0 1.8755
R7763 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.t16 673.346
R7764 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.n19 619.134
R7765 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.t24 611.739
R7766 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.t12 611.739
R7767 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.t18 611.739
R7768 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t27 611.739
R7769 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.t28 421.75
R7770 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.t30 421.75
R7771 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.t11 421.75
R7772 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.t14 421.75
R7773 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.t31 421.75
R7774 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.t29 421.75
R7775 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.t25 421.75
R7776 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.t20 421.75
R7777 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.t23 421.75
R7778 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.t21 421.75
R7779 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.t26 421.75
R7780 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.t13 421.75
R7781 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t22 421.75
R7782 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.t17 421.75
R7783 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.t19 421.75
R7784 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.t15 421.75
R7785 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.t9 288.166
R7786 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.n17 169.125
R7787 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.n8 169.125
R7788 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.n13 167.094
R7789 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.n14 167.094
R7790 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.n15 167.094
R7791 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.n9 167.094
R7792 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.n10 167.094
R7793 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.n11 167.094
R7794 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.n4 167.094
R7795 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.n5 167.094
R7796 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.n6 167.094
R7797 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.n0 167.094
R7798 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.n1 167.094
R7799 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.n2 167.094
R7800 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.n23 140.547
R7801 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n26 140.546
R7802 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n27 139.297
R7803 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.n24 139.297
R7804 bgr_0.VB2_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb2.n22 108.531
R7805 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.t6 62.5402
R7806 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.t10 62.5402
R7807 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.n16 47.1294
R7808 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.n12 47.1294
R7809 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.n7 47.1294
R7810 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.n3 47.1294
R7811 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.n18 38.7817
R7812 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.t4 24.0005
R7813 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.t2 24.0005
R7814 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.t3 24.0005
R7815 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.t1 24.0005
R7816 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.t8 24.0005
R7817 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.t0 24.0005
R7818 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.t5 24.0005
R7819 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.t7 24.0005
R7820 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.n20 14.6443
R7821 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.n21 7.78175
R7822 bgr_0.VB2_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb2.n29 5.6255
R7823 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n25 3.71925
R7824 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n28 3.71925
R7825 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.t16 623.701
R7826 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.t23 611.739
R7827 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.t11 611.739
R7828 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.t17 611.739
R7829 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t26 611.739
R7830 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.t27 421.75
R7831 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.t8 421.75
R7832 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.t10 421.75
R7833 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.t13 421.75
R7834 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.t9 421.75
R7835 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.t28 421.75
R7836 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.t24 421.75
R7837 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.t19 421.75
R7838 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.t22 421.75
R7839 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.t20 421.75
R7840 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.t25 421.75
R7841 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.t12 421.75
R7842 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t21 421.75
R7843 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.t15 421.75
R7844 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.t18 421.75
R7845 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.t14 421.75
R7846 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.n14 176.964
R7847 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.n13 169.343
R7848 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.n20 167.094
R7849 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.n21 167.094
R7850 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.n22 167.094
R7851 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.n16 167.094
R7852 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.n17 167.094
R7853 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.n18 167.094
R7854 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.n9 167.094
R7855 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.n10 167.094
R7856 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.n11 167.094
R7857 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.n5 167.094
R7858 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.n6 167.094
R7859 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.n7 167.094
R7860 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.n24 166.25
R7861 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.n1 139.639
R7862 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.n2 139.638
R7863 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.n0 134.577
R7864 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb3.n26 128.439
R7865 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.n23 47.1294
R7866 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.n19 47.1294
R7867 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.n12 47.1294
R7868 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.n8 47.1294
R7869 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.n15 27.9067
R7870 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t1 24.0005
R7871 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t4 24.0005
R7872 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.t2 24.0005
R7873 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.t6 24.0005
R7874 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.t5 24.0005
R7875 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.t3 24.0005
R7876 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.t0 10.9449
R7877 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.t7 10.9449
R7878 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.n3 4.5005
R7879 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.n25 3.09425
R7880 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb3.n4 0.96925
R7881 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.t13 449.868
R7882 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.t17 449.868
R7883 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.t14 449.868
R7884 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.t18 449.868
R7885 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.n0 339.961
R7886 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.n1 339.272
R7887 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.t24 273.134
R7888 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.t19 273.134
R7889 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.t7 273.134
R7890 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.t16 273.134
R7891 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.t22 273.134
R7892 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.t10 273.134
R7893 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.t20 273.134
R7894 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.t8 273.134
R7895 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.t25 273.134
R7896 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.t12 273.134
R7897 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.t23 273.134
R7898 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.t11 273.134
R7899 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.t21 273.134
R7900 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.t9 273.134
R7901 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.t6 273.134
R7902 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.t15 273.134
R7903 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t3 184.625
R7904 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.n19 176.733
R7905 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.n18 176.733
R7906 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.n17 176.733
R7907 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.n13 176.733
R7908 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.n14 176.733
R7909 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.n15 176.733
R7910 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.n10 176.733
R7911 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.n9 176.733
R7912 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.n8 176.733
R7913 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.n4 176.733
R7914 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.n5 176.733
R7915 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.n6 176.733
R7916 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.n12 170.269
R7917 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.n21 165.8
R7918 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb1.n23 89.8443
R7919 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t2 61.1914
R7920 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.n20 56.2338
R7921 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.n16 56.2338
R7922 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.n11 56.2338
R7923 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.n7 56.2338
R7924 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t0 39.4005
R7925 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t4 39.4005
R7926 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t5 39.4005
R7927 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t1 39.4005
R7928 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.n22 22.3599
R7929 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.n3 6.81097
R7930 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb1.n2 4.46925
R7931 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.n7 114.719
R7932 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n4 114.719
R7933 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.n8 114.156
R7934 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n5 114.156
R7935 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n0 113.081
R7936 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n15 111.769
R7937 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n17 111.769
R7938 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VD1.n19 111.769
R7939 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n1 111.769
R7940 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n3 109.656
R7941 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n12 107.269
R7942 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t8 16.0005
R7943 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t13 16.0005
R7944 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.t18 16.0005
R7945 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.t2 16.0005
R7946 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t20 16.0005
R7947 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t0 16.0005
R7948 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.t1 16.0005
R7949 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.t4 16.0005
R7950 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t5 16.0005
R7951 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t16 16.0005
R7952 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t19 16.0005
R7953 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t21 16.0005
R7954 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t17 16.0005
R7955 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t3 16.0005
R7956 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.t7 16.0005
R7957 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.t12 16.0005
R7958 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t6 16.0005
R7959 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t11 16.0005
R7960 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t9 16.0005
R7961 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t10 16.0005
R7962 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t15 16.0005
R7963 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t14 16.0005
R7964 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n13 4.5005
R7965 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n10 4.5005
R7966 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n14 3.563
R7967 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n16 1.313
R7968 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n2 1.2505
R7969 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VD1.n18 1.2505
R7970 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.n9 0.563
R7971 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.n6 0.563
R7972 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n11 0.21925
R7973 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n3 630.827
R7974 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n8 630.264
R7975 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n6 630.264
R7976 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n4 630.264
R7977 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n13 627.784
R7978 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n0 627.784
R7979 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.n2 627.168
R7980 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n16 626.534
R7981 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n14 626.534
R7982 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.n18 626.534
R7983 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n1 622.034
R7984 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.t9 78.8005
R7985 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.t14 78.8005
R7986 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t6 78.8005
R7987 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t11 78.8005
R7988 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t13 78.8005
R7989 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t17 78.8005
R7990 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t12 78.8005
R7991 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t7 78.8005
R7992 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.t21 78.8005
R7993 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.t5 78.8005
R7994 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t4 78.8005
R7995 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t20 78.8005
R7996 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t19 78.8005
R7997 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t1 78.8005
R7998 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.t2 78.8005
R7999 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.t0 78.8005
R8000 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t3 78.8005
R8001 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t16 78.8005
R8002 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t18 78.8005
R8003 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t8 78.8005
R8004 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.t10 78.8005
R8005 two_stage_opamp_dummy_magic_0.V_err_p.t15 two_stage_opamp_dummy_magic_0.V_err_p.n19 78.8005
R8006 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.n9 5.0005
R8007 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n11 4.5005
R8008 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n10 1.3272
R8009 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n15 1.2505
R8010 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n17 1.2505
R8011 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n12 1.2505
R8012 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n5 0.563
R8013 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n7 0.563
R8014 bgr_0.Vin+.n3 bgr_0.Vin+.n2 526.183
R8015 bgr_0.Vin+.n1 bgr_0.Vin+.n0 514.134
R8016 bgr_0.Vin+.n0 bgr_0.Vin+.t6 303.259
R8017 bgr_0.Vin+.n7 bgr_0.Vin+.n3 215.732
R8018 bgr_0.Vin+.n0 bgr_0.Vin+.t8 174.726
R8019 bgr_0.Vin+.n1 bgr_0.Vin+.t10 174.726
R8020 bgr_0.Vin+.n2 bgr_0.Vin+.t7 174.726
R8021 bgr_0.Vin+.n6 bgr_0.Vin+.n4 170.56
R8022 bgr_0.Vin+.n6 bgr_0.Vin+.n5 168.435
R8023 bgr_0.Vin+.t0 bgr_0.Vin+.n8 158.796
R8024 bgr_0.Vin+.n8 bgr_0.Vin+.t1 147.981
R8025 bgr_0.Vin+.n2 bgr_0.Vin+.n1 128.534
R8026 bgr_0.Vin+.n3 bgr_0.Vin+.t9 96.4005
R8027 bgr_0.Vin+.n7 bgr_0.Vin+.n6 13.5005
R8028 bgr_0.Vin+.n5 bgr_0.Vin+.t2 13.1338
R8029 bgr_0.Vin+.n5 bgr_0.Vin+.t5 13.1338
R8030 bgr_0.Vin+.n4 bgr_0.Vin+.t4 13.1338
R8031 bgr_0.Vin+.n4 bgr_0.Vin+.t3 13.1338
R8032 bgr_0.Vin+.n8 bgr_0.Vin+.n7 1.438
R8033 bgr_0.V_p_1.n6 bgr_0.V_p_1.n1 229.562
R8034 bgr_0.V_p_1.n1 bgr_0.V_p_1.n5 228.939
R8035 bgr_0.V_p_1.n1 bgr_0.V_p_1.n4 228.939
R8036 bgr_0.V_p_1.n0 bgr_0.V_p_1.n3 228.939
R8037 bgr_0.V_p_1.n0 bgr_0.V_p_1.n2 228.939
R8038 bgr_0.V_p_1.n0 bgr_0.V_p_1.t10 98.2279
R8039 bgr_0.V_p_1.n5 bgr_0.V_p_1.t5 48.0005
R8040 bgr_0.V_p_1.n5 bgr_0.V_p_1.t2 48.0005
R8041 bgr_0.V_p_1.n4 bgr_0.V_p_1.t0 48.0005
R8042 bgr_0.V_p_1.n4 bgr_0.V_p_1.t9 48.0005
R8043 bgr_0.V_p_1.n3 bgr_0.V_p_1.t6 48.0005
R8044 bgr_0.V_p_1.n3 bgr_0.V_p_1.t3 48.0005
R8045 bgr_0.V_p_1.n2 bgr_0.V_p_1.t1 48.0005
R8046 bgr_0.V_p_1.n2 bgr_0.V_p_1.t8 48.0005
R8047 bgr_0.V_p_1.t4 bgr_0.V_p_1.n6 48.0005
R8048 bgr_0.V_p_1.n6 bgr_0.V_p_1.t7 48.0005
R8049 bgr_0.V_p_1.n1 bgr_0.V_p_1.n0 1.8755
R8050 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.t6 327.623
R8051 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.t4 326.365
R8052 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t10 168.701
R8053 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t9 168.701
R8054 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.n7 165.8
R8055 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.n5 165.8
R8056 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.n2 165.8
R8057 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.n0 165.8
R8058 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.t5 157.989
R8059 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.t11 157.989
R8060 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t8 157.989
R8061 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t12 157.989
R8062 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.t13 157.989
R8063 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.t7 157.989
R8064 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.t2 117.591
R8065 two_stage_opamp_dummy_magic_0.V_tot.t0 two_stage_opamp_dummy_magic_0.V_tot.n11 117.591
R8066 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.t1 108.424
R8067 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.t3 108.424
R8068 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.n10 42.6121
R8069 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n9 21.2996
R8070 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n8 17.0005
R8071 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.n3 3.31612
R8072 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.n1 1.26612
R8073 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.n6 1.2505
R8074 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.n4 1.15363
R8075 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t13 355.293
R8076 bgr_0.1st_Vout_2.n19 bgr_0.1st_Vout_2.t14 346.8
R8077 bgr_0.1st_Vout_2.n21 bgr_0.1st_Vout_2.n20 339.522
R8078 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.n6 339.522
R8079 bgr_0.1st_Vout_2.n15 bgr_0.1st_Vout_2.n14 335.022
R8080 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.t1 275.909
R8081 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.n10 227.909
R8082 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.n12 222.034
R8083 bgr_0.1st_Vout_2.n17 bgr_0.1st_Vout_2.t26 184.097
R8084 bgr_0.1st_Vout_2.n17 bgr_0.1st_Vout_2.t36 184.097
R8085 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t19 184.097
R8086 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t32 184.097
R8087 bgr_0.1st_Vout_2.n18 bgr_0.1st_Vout_2.n17 166.05
R8088 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.n8 166.05
R8089 bgr_0.1st_Vout_2.n19 bgr_0.1st_Vout_2.n4 57.7228
R8090 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.t10 48.0005
R8091 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.t0 48.0005
R8092 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t9 48.0005
R8093 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t8 48.0005
R8094 bgr_0.1st_Vout_2.n14 bgr_0.1st_Vout_2.t2 39.4005
R8095 bgr_0.1st_Vout_2.n14 bgr_0.1st_Vout_2.t5 39.4005
R8096 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t4 39.4005
R8097 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t6 39.4005
R8098 bgr_0.1st_Vout_2.t7 bgr_0.1st_Vout_2.n21 39.4005
R8099 bgr_0.1st_Vout_2.n21 bgr_0.1st_Vout_2.t3 39.4005
R8100 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t17 4.8295
R8101 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t16 4.8295
R8102 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t27 4.8295
R8103 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t23 4.8295
R8104 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.t35 4.8295
R8105 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t34 4.8295
R8106 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t28 4.8295
R8107 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t21 4.5005
R8108 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t15 4.5005
R8109 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t12 4.5005
R8110 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t30 4.5005
R8111 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t22 4.5005
R8112 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t18 4.5005
R8113 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.t11 4.5005
R8114 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t31 4.5005
R8115 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t29 4.5005
R8116 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t33 4.5005
R8117 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t24 4.5005
R8118 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t20 4.5005
R8119 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t25 4.5005
R8120 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.n11 4.5005
R8121 bgr_0.1st_Vout_2.n16 bgr_0.1st_Vout_2.n15 4.5005
R8122 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.n7 1.3755
R8123 bgr_0.1st_Vout_2.n18 bgr_0.1st_Vout_2.n16 1.3755
R8124 bgr_0.1st_Vout_2.n20 bgr_0.1st_Vout_2.n19 1.188
R8125 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n5 0.9405
R8126 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.n0 0.8935
R8127 bgr_0.1st_Vout_2.n15 bgr_0.1st_Vout_2.n13 0.78175
R8128 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.n2 0.6585
R8129 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.n3 0.6585
R8130 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n1 0.6585
R8131 bgr_0.1st_Vout_2.n16 bgr_0.1st_Vout_2.n9 0.6255
R8132 bgr_0.1st_Vout_2.n20 bgr_0.1st_Vout_2.n18 0.6255
R8133 bgr_0.cap_res2 bgr_0.cap_res2.t20 188.315
R8134 bgr_0.cap_res2 bgr_0.cap_res2.t9 0.259
R8135 bgr_0.cap_res2.t13 bgr_0.cap_res2.t8 0.1603
R8136 bgr_0.cap_res2.t2 bgr_0.cap_res2.t6 0.1603
R8137 bgr_0.cap_res2.t5 bgr_0.cap_res2.t1 0.1603
R8138 bgr_0.cap_res2.t19 bgr_0.cap_res2.t0 0.1603
R8139 bgr_0.cap_res2.t14 bgr_0.cap_res2.t10 0.1603
R8140 bgr_0.cap_res2.t4 bgr_0.cap_res2.t7 0.1603
R8141 bgr_0.cap_res2.t18 bgr_0.cap_res2.t16 0.1603
R8142 bgr_0.cap_res2.t12 bgr_0.cap_res2.t15 0.1603
R8143 bgr_0.cap_res2.n1 bgr_0.cap_res2.t17 0.159278
R8144 bgr_0.cap_res2.n2 bgr_0.cap_res2.t11 0.159278
R8145 bgr_0.cap_res2.n3 bgr_0.cap_res2.t3 0.159278
R8146 bgr_0.cap_res2.n3 bgr_0.cap_res2.t13 0.1368
R8147 bgr_0.cap_res2.n3 bgr_0.cap_res2.t2 0.1368
R8148 bgr_0.cap_res2.n2 bgr_0.cap_res2.t5 0.1368
R8149 bgr_0.cap_res2.n2 bgr_0.cap_res2.t19 0.1368
R8150 bgr_0.cap_res2.n1 bgr_0.cap_res2.t14 0.1368
R8151 bgr_0.cap_res2.n1 bgr_0.cap_res2.t4 0.1368
R8152 bgr_0.cap_res2.n0 bgr_0.cap_res2.t18 0.1368
R8153 bgr_0.cap_res2.n0 bgr_0.cap_res2.t12 0.1368
R8154 bgr_0.cap_res2.t17 bgr_0.cap_res2.n0 0.00152174
R8155 bgr_0.cap_res2.t11 bgr_0.cap_res2.n1 0.00152174
R8156 bgr_0.cap_res2.t3 bgr_0.cap_res2.n2 0.00152174
R8157 bgr_0.cap_res2.t9 bgr_0.cap_res2.n3 0.00152174
R8158 VIN-.n4 VIN-.t8 485.021
R8159 VIN-.n1 VIN-.t6 484.159
R8160 VIN-.n5 VIN-.t7 483.358
R8161 VIN-.n8 VIN-.t10 431.536
R8162 VIN-.n2 VIN-.t9 431.536
R8163 VIN-.n6 VIN-.t1 431.257
R8164 VIN-.n0 VIN-.t0 431.257
R8165 VIN-.n6 VIN-.t2 289.908
R8166 VIN-.n0 VIN-.t5 289.908
R8167 VIN-.n8 VIN-.t4 279.183
R8168 VIN-.n2 VIN-.t3 279.183
R8169 VIN-.n7 VIN-.n6 233.374
R8170 VIN-.n1 VIN-.n0 233.374
R8171 VIN-.n9 VIN-.n8 188.989
R8172 VIN-.n3 VIN-.n2 188.989
R8173 VIN-.n4 VIN-.n3 2.463
R8174 VIN- VIN-.n9 2.03175
R8175 VIN-.n5 VIN-.n4 1.563
R8176 VIN-.n3 VIN-.n1 1.2755
R8177 VIN-.n9 VIN-.n7 1.2755
R8178 VIN-.n7 VIN-.n5 0.8005
R8179 two_stage_opamp_dummy_magic_0.V_p.n20 two_stage_opamp_dummy_magic_0.V_p.t29 202.595
R8180 two_stage_opamp_dummy_magic_0.V_p.n5 two_stage_opamp_dummy_magic_0.V_p.n3 118.168
R8181 two_stage_opamp_dummy_magic_0.V_p.n2 two_stage_opamp_dummy_magic_0.V_p.n0 117.831
R8182 two_stage_opamp_dummy_magic_0.V_p.n36 two_stage_opamp_dummy_magic_0.V_p.n35 117.269
R8183 two_stage_opamp_dummy_magic_0.V_p.n11 two_stage_opamp_dummy_magic_0.V_p.n10 117.269
R8184 two_stage_opamp_dummy_magic_0.V_p.n9 two_stage_opamp_dummy_magic_0.V_p.n8 117.269
R8185 two_stage_opamp_dummy_magic_0.V_p.n7 two_stage_opamp_dummy_magic_0.V_p.n6 117.269
R8186 two_stage_opamp_dummy_magic_0.V_p.n5 two_stage_opamp_dummy_magic_0.V_p.n4 117.269
R8187 two_stage_opamp_dummy_magic_0.V_p.n2 two_stage_opamp_dummy_magic_0.V_p.n1 117.269
R8188 two_stage_opamp_dummy_magic_0.V_p.n38 two_stage_opamp_dummy_magic_0.V_p.n37 117.267
R8189 two_stage_opamp_dummy_magic_0.V_p.n33 two_stage_opamp_dummy_magic_0.V_p.n12 113.136
R8190 two_stage_opamp_dummy_magic_0.V_p.n30 two_stage_opamp_dummy_magic_0.V_p.n13 101.335
R8191 two_stage_opamp_dummy_magic_0.V_p.n16 two_stage_opamp_dummy_magic_0.V_p.n14 99.647
R8192 two_stage_opamp_dummy_magic_0.V_p.n29 two_stage_opamp_dummy_magic_0.V_p.n28 99.0845
R8193 two_stage_opamp_dummy_magic_0.V_p.n27 two_stage_opamp_dummy_magic_0.V_p.n26 99.0845
R8194 two_stage_opamp_dummy_magic_0.V_p.n25 two_stage_opamp_dummy_magic_0.V_p.n24 99.0845
R8195 two_stage_opamp_dummy_magic_0.V_p.n23 two_stage_opamp_dummy_magic_0.V_p.n22 99.0845
R8196 two_stage_opamp_dummy_magic_0.V_p.n18 two_stage_opamp_dummy_magic_0.V_p.n17 99.0845
R8197 two_stage_opamp_dummy_magic_0.V_p.n16 two_stage_opamp_dummy_magic_0.V_p.n15 99.0845
R8198 two_stage_opamp_dummy_magic_0.V_p.n32 two_stage_opamp_dummy_magic_0.V_p.n31 94.5845
R8199 two_stage_opamp_dummy_magic_0.V_p.n20 two_stage_opamp_dummy_magic_0.V_p.n19 94.5845
R8200 two_stage_opamp_dummy_magic_0.V_p.n35 two_stage_opamp_dummy_magic_0.V_p.t13 16.0005
R8201 two_stage_opamp_dummy_magic_0.V_p.n35 two_stage_opamp_dummy_magic_0.V_p.t22 16.0005
R8202 two_stage_opamp_dummy_magic_0.V_p.n12 two_stage_opamp_dummy_magic_0.V_p.t17 16.0005
R8203 two_stage_opamp_dummy_magic_0.V_p.n12 two_stage_opamp_dummy_magic_0.V_p.t5 16.0005
R8204 two_stage_opamp_dummy_magic_0.V_p.n10 two_stage_opamp_dummy_magic_0.V_p.t18 16.0005
R8205 two_stage_opamp_dummy_magic_0.V_p.n10 two_stage_opamp_dummy_magic_0.V_p.t4 16.0005
R8206 two_stage_opamp_dummy_magic_0.V_p.n8 two_stage_opamp_dummy_magic_0.V_p.t26 16.0005
R8207 two_stage_opamp_dummy_magic_0.V_p.n8 two_stage_opamp_dummy_magic_0.V_p.t23 16.0005
R8208 two_stage_opamp_dummy_magic_0.V_p.n6 two_stage_opamp_dummy_magic_0.V_p.t24 16.0005
R8209 two_stage_opamp_dummy_magic_0.V_p.n6 two_stage_opamp_dummy_magic_0.V_p.t15 16.0005
R8210 two_stage_opamp_dummy_magic_0.V_p.n4 two_stage_opamp_dummy_magic_0.V_p.t8 16.0005
R8211 two_stage_opamp_dummy_magic_0.V_p.n4 two_stage_opamp_dummy_magic_0.V_p.t21 16.0005
R8212 two_stage_opamp_dummy_magic_0.V_p.n3 two_stage_opamp_dummy_magic_0.V_p.t16 16.0005
R8213 two_stage_opamp_dummy_magic_0.V_p.n3 two_stage_opamp_dummy_magic_0.V_p.t34 16.0005
R8214 two_stage_opamp_dummy_magic_0.V_p.n1 two_stage_opamp_dummy_magic_0.V_p.t12 16.0005
R8215 two_stage_opamp_dummy_magic_0.V_p.n1 two_stage_opamp_dummy_magic_0.V_p.t20 16.0005
R8216 two_stage_opamp_dummy_magic_0.V_p.n0 two_stage_opamp_dummy_magic_0.V_p.t19 16.0005
R8217 two_stage_opamp_dummy_magic_0.V_p.n0 two_stage_opamp_dummy_magic_0.V_p.t3 16.0005
R8218 two_stage_opamp_dummy_magic_0.V_p.t25 two_stage_opamp_dummy_magic_0.V_p.n38 16.0005
R8219 two_stage_opamp_dummy_magic_0.V_p.n38 two_stage_opamp_dummy_magic_0.V_p.t36 16.0005
R8220 two_stage_opamp_dummy_magic_0.V_p.n31 two_stage_opamp_dummy_magic_0.V_p.t14 9.6005
R8221 two_stage_opamp_dummy_magic_0.V_p.n31 two_stage_opamp_dummy_magic_0.V_p.t0 9.6005
R8222 two_stage_opamp_dummy_magic_0.V_p.n28 two_stage_opamp_dummy_magic_0.V_p.t33 9.6005
R8223 two_stage_opamp_dummy_magic_0.V_p.n28 two_stage_opamp_dummy_magic_0.V_p.t39 9.6005
R8224 two_stage_opamp_dummy_magic_0.V_p.n26 two_stage_opamp_dummy_magic_0.V_p.t30 9.6005
R8225 two_stage_opamp_dummy_magic_0.V_p.n26 two_stage_opamp_dummy_magic_0.V_p.t9 9.6005
R8226 two_stage_opamp_dummy_magic_0.V_p.n24 two_stage_opamp_dummy_magic_0.V_p.t11 9.6005
R8227 two_stage_opamp_dummy_magic_0.V_p.n24 two_stage_opamp_dummy_magic_0.V_p.t7 9.6005
R8228 two_stage_opamp_dummy_magic_0.V_p.n22 two_stage_opamp_dummy_magic_0.V_p.t28 9.6005
R8229 two_stage_opamp_dummy_magic_0.V_p.n22 two_stage_opamp_dummy_magic_0.V_p.t32 9.6005
R8230 two_stage_opamp_dummy_magic_0.V_p.n19 two_stage_opamp_dummy_magic_0.V_p.t27 9.6005
R8231 two_stage_opamp_dummy_magic_0.V_p.n19 two_stage_opamp_dummy_magic_0.V_p.t10 9.6005
R8232 two_stage_opamp_dummy_magic_0.V_p.n17 two_stage_opamp_dummy_magic_0.V_p.t40 9.6005
R8233 two_stage_opamp_dummy_magic_0.V_p.n17 two_stage_opamp_dummy_magic_0.V_p.t31 9.6005
R8234 two_stage_opamp_dummy_magic_0.V_p.n15 two_stage_opamp_dummy_magic_0.V_p.t35 9.6005
R8235 two_stage_opamp_dummy_magic_0.V_p.n15 two_stage_opamp_dummy_magic_0.V_p.t6 9.6005
R8236 two_stage_opamp_dummy_magic_0.V_p.n14 two_stage_opamp_dummy_magic_0.V_p.t2 9.6005
R8237 two_stage_opamp_dummy_magic_0.V_p.n14 two_stage_opamp_dummy_magic_0.V_p.t1 9.6005
R8238 two_stage_opamp_dummy_magic_0.V_p.n13 two_stage_opamp_dummy_magic_0.V_p.t38 9.6005
R8239 two_stage_opamp_dummy_magic_0.V_p.n13 two_stage_opamp_dummy_magic_0.V_p.t37 9.6005
R8240 two_stage_opamp_dummy_magic_0.V_p.n21 two_stage_opamp_dummy_magic_0.V_p.n20 4.5005
R8241 two_stage_opamp_dummy_magic_0.V_p.n32 two_stage_opamp_dummy_magic_0.V_p.n30 4.5005
R8242 two_stage_opamp_dummy_magic_0.V_p.n34 two_stage_opamp_dummy_magic_0.V_p.n33 4.5005
R8243 two_stage_opamp_dummy_magic_0.V_p.n34 two_stage_opamp_dummy_magic_0.V_p.n11 3.65675
R8244 two_stage_opamp_dummy_magic_0.V_p.n33 two_stage_opamp_dummy_magic_0.V_p.n32 1.28175
R8245 two_stage_opamp_dummy_magic_0.V_p.n18 two_stage_opamp_dummy_magic_0.V_p.n16 0.563
R8246 two_stage_opamp_dummy_magic_0.V_p.n21 two_stage_opamp_dummy_magic_0.V_p.n18 0.563
R8247 two_stage_opamp_dummy_magic_0.V_p.n23 two_stage_opamp_dummy_magic_0.V_p.n21 0.563
R8248 two_stage_opamp_dummy_magic_0.V_p.n25 two_stage_opamp_dummy_magic_0.V_p.n23 0.563
R8249 two_stage_opamp_dummy_magic_0.V_p.n27 two_stage_opamp_dummy_magic_0.V_p.n25 0.563
R8250 two_stage_opamp_dummy_magic_0.V_p.n29 two_stage_opamp_dummy_magic_0.V_p.n27 0.563
R8251 two_stage_opamp_dummy_magic_0.V_p.n30 two_stage_opamp_dummy_magic_0.V_p.n29 0.563
R8252 two_stage_opamp_dummy_magic_0.V_p.n7 two_stage_opamp_dummy_magic_0.V_p.n5 0.563
R8253 two_stage_opamp_dummy_magic_0.V_p.n9 two_stage_opamp_dummy_magic_0.V_p.n7 0.563
R8254 two_stage_opamp_dummy_magic_0.V_p.n11 two_stage_opamp_dummy_magic_0.V_p.n9 0.563
R8255 two_stage_opamp_dummy_magic_0.V_p.n37 two_stage_opamp_dummy_magic_0.V_p.n36 0.563
R8256 two_stage_opamp_dummy_magic_0.V_p.n37 two_stage_opamp_dummy_magic_0.V_p.n2 0.563
R8257 two_stage_opamp_dummy_magic_0.V_p.n36 two_stage_opamp_dummy_magic_0.V_p.n34 0.53175
R8258 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 610.534
R8259 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 610.534
R8260 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 433.8
R8261 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 433.8
R8262 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 433.8
R8263 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 433.8
R8264 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 433.8
R8265 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 433.8
R8266 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 433.8
R8267 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 433.8
R8268 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 433.8
R8269 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 433.8
R8270 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 433.8
R8271 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 433.8
R8272 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 433.8
R8273 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 433.8
R8274 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 433.8
R8275 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 433.8
R8276 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 433.8
R8277 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 433.8
R8278 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 339.836
R8279 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 339.834
R8280 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 339.272
R8281 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 334.772
R8282 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 221.293
R8283 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 176.733
R8284 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 176.733
R8285 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 176.733
R8286 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 176.733
R8287 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 176.733
R8288 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 176.733
R8289 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 176.733
R8290 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 176.733
R8291 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 176.733
R8292 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 176.733
R8293 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 176.733
R8294 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 176.733
R8295 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 176.733
R8296 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 176.733
R8297 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 176.733
R8298 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 176.733
R8299 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 118.45
R8300 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.V_tail_gate.n29 86.7036
R8301 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 64.5795
R8302 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 56.2338
R8303 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 56.2338
R8304 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 53.2453
R8305 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 39.4005
R8306 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 39.4005
R8307 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 39.4005
R8308 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 39.4005
R8309 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 39.4005
R8310 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 39.4005
R8311 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 39.4005
R8312 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 39.4005
R8313 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.V_tail_gate.n6 18.3599
R8314 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 16.0005
R8315 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 16.0005
R8316 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 16.0005
R8317 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 16.0005
R8318 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 4.5005
R8319 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 0.563
R8320 a_11220_17410.t0 a_11220_17410.t1 258.591
R8321 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 144.827
R8322 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 134.577
R8323 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 120.66
R8324 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 97.4009
R8325 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 96.8384
R8326 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 96.8384
R8327 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 96.8384
R8328 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 96.8384
R8329 bgr_0.V_CMFB_S2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 95.9693
R8330 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 24.0005
R8331 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 24.0005
R8332 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 24.0005
R8333 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 24.0005
R8334 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 8.0005
R8335 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 8.0005
R8336 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 8.0005
R8337 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 8.0005
R8338 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 8.0005
R8339 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 8.0005
R8340 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 8.0005
R8341 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 8.0005
R8342 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 8.0005
R8343 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 8.0005
R8344 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 5.813
R8345 bgr_0.V_CMFB_S2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 1.46925
R8346 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 0.563
R8347 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 0.563
R8348 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 0.563
R8349 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n1 4020
R8350 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.n1 4020
R8351 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n7 4020
R8352 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.n7 4020
R8353 two_stage_opamp_dummy_magic_0.VD4.n4 two_stage_opamp_dummy_magic_0.VD4.t22 660.109
R8354 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.t25 660.109
R8355 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n11 428.8
R8356 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n0 428.8
R8357 two_stage_opamp_dummy_magic_0.VD4.t23 two_stage_opamp_dummy_magic_0.VD4.n8 239.915
R8358 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.t26 239.915
R8359 two_stage_opamp_dummy_magic_0.VD4.n6 two_stage_opamp_dummy_magic_0.VD4.n5 230.4
R8360 two_stage_opamp_dummy_magic_0.VD4.n6 two_stage_opamp_dummy_magic_0.VD4.n3 230.4
R8361 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n3 198.4
R8362 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.n0 198.4
R8363 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.n28 160.428
R8364 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.n15 160.427
R8365 two_stage_opamp_dummy_magic_0.VD4.n22 two_stage_opamp_dummy_magic_0.VD4.n14 160.427
R8366 two_stage_opamp_dummy_magic_0.VD4.n25 two_stage_opamp_dummy_magic_0.VD4.n13 160.053
R8367 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.n29 159.803
R8368 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n26 159.803
R8369 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.n20 159.802
R8370 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.n18 159.802
R8371 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.n16 159.802
R8372 two_stage_opamp_dummy_magic_0.VD4.n24 two_stage_opamp_dummy_magic_0.VD4.n23 155.302
R8373 two_stage_opamp_dummy_magic_0.VD4.n4 two_stage_opamp_dummy_magic_0.VD4.t24 155.125
R8374 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.t27 155.125
R8375 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.n32 146.004
R8376 two_stage_opamp_dummy_magic_0.VD4.t2 two_stage_opamp_dummy_magic_0.VD4.t23 98.2764
R8377 two_stage_opamp_dummy_magic_0.VD4.t8 two_stage_opamp_dummy_magic_0.VD4.t2 98.2764
R8378 two_stage_opamp_dummy_magic_0.VD4.t16 two_stage_opamp_dummy_magic_0.VD4.t8 98.2764
R8379 two_stage_opamp_dummy_magic_0.VD4.t12 two_stage_opamp_dummy_magic_0.VD4.t16 98.2764
R8380 two_stage_opamp_dummy_magic_0.VD4.t18 two_stage_opamp_dummy_magic_0.VD4.t12 98.2764
R8381 two_stage_opamp_dummy_magic_0.VD4.t4 two_stage_opamp_dummy_magic_0.VD4.t20 98.2764
R8382 two_stage_opamp_dummy_magic_0.VD4.t10 two_stage_opamp_dummy_magic_0.VD4.t4 98.2764
R8383 two_stage_opamp_dummy_magic_0.VD4.t6 two_stage_opamp_dummy_magic_0.VD4.t10 98.2764
R8384 two_stage_opamp_dummy_magic_0.VD4.t14 two_stage_opamp_dummy_magic_0.VD4.t6 98.2764
R8385 two_stage_opamp_dummy_magic_0.VD4.t26 two_stage_opamp_dummy_magic_0.VD4.t14 98.2764
R8386 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n10 92.5005
R8387 two_stage_opamp_dummy_magic_0.VD4.n7 two_stage_opamp_dummy_magic_0.VD4.n6 92.5005
R8388 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.n7 92.5005
R8389 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n0 92.5005
R8390 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n1 92.5005
R8391 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.n1 92.5005
R8392 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.t18 49.1384
R8393 two_stage_opamp_dummy_magic_0.VD4.t20 two_stage_opamp_dummy_magic_0.VD4.n9 49.1384
R8394 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.n4 21.3338
R8395 two_stage_opamp_dummy_magic_0.VD4.n3 two_stage_opamp_dummy_magic_0.VD4.n2 21.3338
R8396 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.n12 19.2005
R8397 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.n31 13.8005
R8398 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.t5 11.2576
R8399 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.t11 11.2576
R8400 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.t7 11.2576
R8401 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.t15 11.2576
R8402 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.t17 11.2576
R8403 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.t13 11.2576
R8404 two_stage_opamp_dummy_magic_0.VD4.n23 two_stage_opamp_dummy_magic_0.VD4.t31 11.2576
R8405 two_stage_opamp_dummy_magic_0.VD4.n23 two_stage_opamp_dummy_magic_0.VD4.t35 11.2576
R8406 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.t33 11.2576
R8407 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.t36 11.2576
R8408 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.t37 11.2576
R8409 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.t29 11.2576
R8410 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.t32 11.2576
R8411 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.t30 11.2576
R8412 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.t34 11.2576
R8413 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.t1 11.2576
R8414 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.t0 11.2576
R8415 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.t28 11.2576
R8416 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.t3 11.2576
R8417 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.t9 11.2576
R8418 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.t19 11.2576
R8419 two_stage_opamp_dummy_magic_0.VD4.t21 two_stage_opamp_dummy_magic_0.VD4.n33 11.2576
R8420 two_stage_opamp_dummy_magic_0.VD4.n25 two_stage_opamp_dummy_magic_0.VD4.n24 6.188
R8421 two_stage_opamp_dummy_magic_0.VD4.n24 two_stage_opamp_dummy_magic_0.VD4.n22 4.5005
R8422 two_stage_opamp_dummy_magic_0.VD4.n31 two_stage_opamp_dummy_magic_0.VD4.n30 0.6255
R8423 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.n17 0.6255
R8424 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.n19 0.6255
R8425 two_stage_opamp_dummy_magic_0.VD4.n22 two_stage_opamp_dummy_magic_0.VD4.n21 0.6255
R8426 two_stage_opamp_dummy_magic_0.VD4.n31 two_stage_opamp_dummy_magic_0.VD4.n27 0.6255
R8427 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n25 0.2505
R8428 VIN+.n9 VIN+.t5 485.127
R8429 VIN+.n4 VIN+.t3 485.127
R8430 VIN+.n3 VIN+.t4 485.127
R8431 VIN+.n7 VIN+.t9 318.656
R8432 VIN+.n7 VIN+.t2 318.656
R8433 VIN+.n5 VIN+.t7 318.656
R8434 VIN+.n5 VIN+.t1 318.656
R8435 VIN+.n1 VIN+.t8 318.656
R8436 VIN+.n1 VIN+.t6 318.656
R8437 VIN+.n0 VIN+.t10 318.656
R8438 VIN+.n0 VIN+.t0 318.656
R8439 VIN+.n2 VIN+.n0 167.05
R8440 VIN+.n8 VIN+.n7 165.8
R8441 VIN+.n6 VIN+.n5 165.8
R8442 VIN+.n2 VIN+.n1 165.8
R8443 VIN+.n6 VIN+.n4 2.34425
R8444 VIN+.n4 VIN+.n3 1.3005
R8445 VIN+.n8 VIN+.n6 1.2505
R8446 VIN+ VIN+.n9 1.213
R8447 VIN+.n3 VIN+.n2 1.15675
R8448 VIN+.n9 VIN+.n8 1.15675
R8449 a_13730_17020.t0 a_13730_17020.t1 258.591
R8450 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.n2 526.183
R8451 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.n0 514.134
R8452 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t3 303.259
R8453 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n4 287.264
R8454 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n3 283.961
R8455 bgr_0.V_CUR_REF_REG.t0 bgr_0.V_CUR_REF_REG.n5 245.284
R8456 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t7 174.726
R8457 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t5 174.726
R8458 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.t6 174.726
R8459 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.n1 128.534
R8460 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.t4 96.4005
R8461 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t1 39.4005
R8462 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t2 39.4005
R8463 a_12828_17530.t0 a_12828_17530.t1 376.99
R8464 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.t12 650.729
R8465 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.n6 630.607
R8466 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n8 627.128
R8467 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n10 627.128
R8468 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.n0 227.784
R8469 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.n1 226.534
R8470 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.n3 226.534
R8471 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.t10 78.8005
R8472 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.t4 78.8005
R8473 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.t1 78.8005
R8474 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.t3 78.8005
R8475 two_stage_opamp_dummy_magic_0.err_amp_out.n10 two_stage_opamp_dummy_magic_0.err_amp_out.t0 78.8005
R8476 two_stage_opamp_dummy_magic_0.err_amp_out.n10 two_stage_opamp_dummy_magic_0.err_amp_out.t2 78.8005
R8477 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t6 48.0005
R8478 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t8 48.0005
R8479 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t5 48.0005
R8480 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t7 48.0005
R8481 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t11 48.0005
R8482 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t9 48.0005
R8483 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.n5 21.1255
R8484 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.n4 10.8755
R8485 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n7 1.3755
R8486 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.n2 1.2505
R8487 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n9 1.2505
R8488 bgr_0.START_UP.n4 bgr_0.START_UP.t6 238.322
R8489 bgr_0.START_UP.n4 bgr_0.START_UP.t7 238.322
R8490 bgr_0.START_UP.n3 bgr_0.START_UP.n1 175.56
R8491 bgr_0.START_UP.n3 bgr_0.START_UP.n2 168.936
R8492 bgr_0.START_UP.n5 bgr_0.START_UP.n4 166.925
R8493 bgr_0.START_UP.n0 bgr_0.START_UP.t5 130.001
R8494 bgr_0.START_UP.n0 bgr_0.START_UP.t4 81.7074
R8495 bgr_0.START_UP bgr_0.START_UP.n0 38.2614
R8496 bgr_0.START_UP bgr_0.START_UP.n5 14.7817
R8497 bgr_0.START_UP.n1 bgr_0.START_UP.t0 13.1338
R8498 bgr_0.START_UP.n1 bgr_0.START_UP.t1 13.1338
R8499 bgr_0.START_UP.n2 bgr_0.START_UP.t2 13.1338
R8500 bgr_0.START_UP.n2 bgr_0.START_UP.t3 13.1338
R8501 bgr_0.START_UP.n5 bgr_0.START_UP.n3 4.21925
R8502 a_5230_5738.t0 a_5230_5738.t1 294.339
R8503 a_11220_17290.t0 a_11220_17290.t1 376.99
R8504 a_12828_17650.t0 a_12828_17650.t1 258.591
R8505 a_14520_5738.t0 a_14520_5738.t1 294.339
R8506 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 2655
R8507 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 2595
R8508 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 2280
R8509 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 2250
R8510 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 672.159
R8511 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 672.159
R8512 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 276.8
R8513 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 240
R8514 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 206.4
R8515 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 204.8
R8516 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 180.904
R8517 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 170.3
R8518 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 160.517
R8519 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 160.517
R8520 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 110.425
R8521 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 110.05
R8522 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 95.7988
R8523 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 92.5005
R8524 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 92.5005
R8525 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 92.5005
R8526 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 92.5005
R8527 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 89.6005
R8528 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 89.6005
R8529 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 76.8005
R8530 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 75.9449
R8531 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 75.9449
R8532 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 47.8997
R8533 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 47.8997
R8534 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 38.4005
R8535 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 24.5338
R8536 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 24.5338
R8537 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 16.8187
R8538 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 16.8187
R8539 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 12.313
R8540 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 12.313
R8541 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 10.9449
R8542 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 10.9449
R8543 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 6.21925
R8544 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 4.5005
R8545 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.n0 220.678
R8546 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t0 16.0005
R8547 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t1 16.0005
R8548 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.t3 9.6005
R8549 two_stage_opamp_dummy_magic_0.V_p_mir.t2 two_stage_opamp_dummy_magic_0.V_p_mir.n1 9.6005
R8550 a_5350_5738.t0 a_5350_5738.t1 169.905
R8551 a_14240_2946.t0 a_14240_2946.t1 169.905
R8552 a_13790_17550.t0 a_13790_17550.t1 258.591
C0 two_stage_opamp_dummy_magic_0.Y VOUT+ 2.10995f
C1 bgr_0.PFET_GATE_10uA bgr_0.V_TOP 2.47368f
C2 VIN- VIN+ 0.555219f
C3 bgr_0.Vbe2 bgr_0.PFET_GATE_10uA 0.242909f
C4 VDDA bgr_0.PFET_GATE_10uA 10.3925f
C5 VOUT- VOUT+ 0.210644f
C6 VIN+ two_stage_opamp_dummy_magic_0.VD1 0.057219f
C7 bgr_0.PFET_GATE_10uA bgr_0.1st_Vout_1 0.035393f
C8 li_10610_16720# bgr_0.cap_res2 0.020538f
C9 bgr_0.cap_res2 bgr_0.PFET_GATE_10uA 0.018633f
C10 bgr_0.NFET_GATE_10uA bgr_0.PFET_GATE_10uA 0.050552f
C11 li_12710_16610# bgr_0.1st_Vout_1 0.020439f
C12 VDDA two_stage_opamp_dummy_magic_0.V_err_gate 4.21536f
C13 m2_7180_19780# bgr_0.PFET_GATE_10uA 0.012f
C14 bgr_0.START_UP bgr_0.V_TOP 0.815644f
C15 li_7110_16510# VDDA 0.021911f
C16 bgr_0.START_UP bgr_0.Vbe2 0.193132f
C17 VDDA bgr_0.START_UP 1.37392f
C18 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_gate 0.136183f
C19 bgr_0.START_UP bgr_0.1st_Vout_1 0.030647f
C20 bgr_0.START_UP_NFET1 bgr_0.START_UP 0.145663f
C21 m2_8540_19780# bgr_0.V_TOP 0.012f
C22 m2_8540_19780# VDDA 0.010446f
C23 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.V_err_gate 0.011317f
C24 bgr_0.NFET_GATE_10uA bgr_0.START_UP 0.518732f
C25 m2_8540_19780# bgr_0.1st_Vout_1 0.075543f
C26 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.V_err_gate 0.03991f
C27 two_stage_opamp_dummy_magic_0.cap_res_X VDDA 0.770449f
C28 two_stage_opamp_dummy_magic_0.err_amp_out VDDA 1.00936f
C29 bgr_0.V_TOP two_stage_opamp_dummy_magic_0.V_err_amp_ref 1.13839f
C30 bgr_0.Vbe2 two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.014154f
C31 VDDA two_stage_opamp_dummy_magic_0.V_err_amp_ref 4.30887f
C32 two_stage_opamp_dummy_magic_0.cap_res_X bgr_0.cap_res2 0.048779f
C33 two_stage_opamp_dummy_magic_0.V_err_amp_ref bgr_0.1st_Vout_1 0.477103f
C34 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.Y 1.06369f
C35 bgr_0.cap_res2 two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.551434f
C36 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.559544f
C37 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.Vb2_Vb3 0.04831f
C38 VOUT+ two_stage_opamp_dummy_magic_0.V_err_gate 0.037082f
C39 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.Y 0.040365f
C40 two_stage_opamp_dummy_magic_0.cap_res_X VOUT- 50.7533f
C41 VOUT- two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.055846f
C42 two_stage_opamp_dummy_magic_0.cap_res_X VOUT+ 0.020189f
C43 li_5710_16610# bgr_0.V_TOP 0.020062f
C44 bgr_0.Vbe2 bgr_0.V_TOP 0.285619f
C45 VDDA bgr_0.V_TOP 16.1354f
C46 VDDA bgr_0.Vbe2 0.016701f
C47 bgr_0.V_TOP bgr_0.1st_Vout_1 0.925484f
C48 VDDA bgr_0.1st_Vout_1 2.06087f
C49 bgr_0.START_UP bgr_0.PFET_GATE_10uA 0.166283f
C50 VDDA bgr_0.START_UP_NFET1 0.150608f
C51 bgr_0.NFET_GATE_10uA bgr_0.V_TOP 0.080353f
C52 VDDA bgr_0.cap_res2 0.58582f
C53 bgr_0.NFET_GATE_10uA bgr_0.Vbe2 0.021455f
C54 VDDA bgr_0.NFET_GATE_10uA 1.04958f
C55 bgr_0.cap_res2 bgr_0.1st_Vout_1 0.822981f
C56 bgr_0.NFET_GATE_10uA bgr_0.1st_Vout_1 1.02268f
C57 m2_7180_19780# VDDA 0.010446f
C58 bgr_0.NFET_GATE_10uA bgr_0.START_UP_NFET1 0.318695f
C59 VDDA two_stage_opamp_dummy_magic_0.VD3 3.69967f
C60 VDDA two_stage_opamp_dummy_magic_0.Vb2_Vb3 0.953371f
C61 two_stage_opamp_dummy_magic_0.Y VDDA 4.15025f
C62 bgr_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_amp_ref 2.46518f
C63 VIN- two_stage_opamp_dummy_magic_0.VD1 0.881219f
C64 VDDA VOUT- 6.78204f
C65 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_amp_ref 1.3653f
C66 VDDA VOUT+ 6.69227f
C67 bgr_0.START_UP two_stage_opamp_dummy_magic_0.V_err_amp_ref 2.09763f
C68 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.err_amp_out 0.017583f
C69 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.V_err_amp_ref 1.03641f
C70 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.406563f
C71 VOUT+ two_stage_opamp_dummy_magic_0.Vb2_Vb3 0.059472f
C72 VIN+ GNDA 2.09083f
C73 VIN- GNDA 2.156752f
C74 VOUT+ GNDA 17.68936f
C75 VOUT- GNDA 17.676865f
C76 VDDA GNDA 0.149176p
C77 li_7110_16510# GNDA 0.050654f $ **FLOATING
C78 li_14110_16610# GNDA 0.050514f $ **FLOATING
C79 li_12710_16610# GNDA 0.049721f $ **FLOATING
C80 li_5710_16610# GNDA 0.047034f $ **FLOATING
C81 li_10610_16720# GNDA 0.049096f $ **FLOATING
C82 li_9210_16720# GNDA 0.043891f $ **FLOATING
C83 two_stage_opamp_dummy_magic_0.VD1 GNDA 2.38758f
C84 two_stage_opamp_dummy_magic_0.Y GNDA 4.953576f
C85 two_stage_opamp_dummy_magic_0.cap_res_X GNDA 33.10225f
C86 two_stage_opamp_dummy_magic_0.err_amp_out GNDA 2.932267f
C87 bgr_0.cap_res2 GNDA 7.936877f
C88 bgr_0.1st_Vout_1 GNDA 4.986571f
C89 two_stage_opamp_dummy_magic_0.V_err_amp_ref GNDA 13.86926f
C90 bgr_0.V_TOP GNDA 6.838887f
C91 bgr_0.PFET_GATE_10uA GNDA 5.13254f
C92 bgr_0.Vbe2 GNDA 17.0659f
C93 bgr_0.START_UP GNDA 7.190383f
C94 bgr_0.START_UP_NFET1 GNDA 5.28339f
C95 two_stage_opamp_dummy_magic_0.V_err_gate GNDA 14.820534f
C96 bgr_0.NFET_GATE_10uA GNDA 7.08898f
C97 two_stage_opamp_dummy_magic_0.VD3 GNDA 6.533089f
C98 two_stage_opamp_dummy_magic_0.Vb2_Vb3 GNDA 3.53474f
C99 bgr_0.START_UP.t4 GNDA 1.6623f
C100 bgr_0.START_UP.t5 GNDA 0.043697f
C101 bgr_0.START_UP.n0 GNDA 1.12862f
C102 bgr_0.START_UP.t0 GNDA 0.041701f
C103 bgr_0.START_UP.t1 GNDA 0.041701f
C104 bgr_0.START_UP.n1 GNDA 0.151283f
C105 bgr_0.START_UP.t2 GNDA 0.041701f
C106 bgr_0.START_UP.t3 GNDA 0.041701f
C107 bgr_0.START_UP.n2 GNDA 0.139173f
C108 bgr_0.START_UP.n3 GNDA 0.720787f
C109 bgr_0.START_UP.t7 GNDA 0.01567f
C110 bgr_0.START_UP.t6 GNDA 0.01567f
C111 bgr_0.START_UP.n4 GNDA 0.044238f
C112 bgr_0.START_UP.n5 GNDA 0.445182f
C113 two_stage_opamp_dummy_magic_0.err_amp_out.t5 GNDA 0.013381f
C114 two_stage_opamp_dummy_magic_0.err_amp_out.t7 GNDA 0.013381f
C115 two_stage_opamp_dummy_magic_0.err_amp_out.n0 GNDA 0.038511f
C116 two_stage_opamp_dummy_magic_0.err_amp_out.t6 GNDA 0.013381f
C117 two_stage_opamp_dummy_magic_0.err_amp_out.t8 GNDA 0.013381f
C118 two_stage_opamp_dummy_magic_0.err_amp_out.n1 GNDA 0.037365f
C119 two_stage_opamp_dummy_magic_0.err_amp_out.n2 GNDA 0.464702f
C120 two_stage_opamp_dummy_magic_0.err_amp_out.t11 GNDA 0.013381f
C121 two_stage_opamp_dummy_magic_0.err_amp_out.t9 GNDA 0.013381f
C122 two_stage_opamp_dummy_magic_0.err_amp_out.n3 GNDA 0.037365f
C123 two_stage_opamp_dummy_magic_0.err_amp_out.n4 GNDA 0.496077f
C124 two_stage_opamp_dummy_magic_0.err_amp_out.t12 GNDA 0.095614f
C125 two_stage_opamp_dummy_magic_0.err_amp_out.n5 GNDA 1.60863f
C126 two_stage_opamp_dummy_magic_0.err_amp_out.t10 GNDA 0.013381f
C127 two_stage_opamp_dummy_magic_0.err_amp_out.t4 GNDA 0.013381f
C128 two_stage_opamp_dummy_magic_0.err_amp_out.n6 GNDA 0.031078f
C129 two_stage_opamp_dummy_magic_0.err_amp_out.n7 GNDA 0.918238f
C130 two_stage_opamp_dummy_magic_0.err_amp_out.t1 GNDA 0.013381f
C131 two_stage_opamp_dummy_magic_0.err_amp_out.t3 GNDA 0.013381f
C132 two_stage_opamp_dummy_magic_0.err_amp_out.n8 GNDA 0.031328f
C133 two_stage_opamp_dummy_magic_0.err_amp_out.n9 GNDA 0.351359f
C134 two_stage_opamp_dummy_magic_0.err_amp_out.t0 GNDA 0.013381f
C135 two_stage_opamp_dummy_magic_0.err_amp_out.t2 GNDA 0.013381f
C136 two_stage_opamp_dummy_magic_0.err_amp_out.n10 GNDA 0.031328f
C137 bgr_0.V_CUR_REF_REG.t3 GNDA 0.014208f
C138 bgr_0.V_CUR_REF_REG.n0 GNDA 0.030473f
C139 bgr_0.V_CUR_REF_REG.n1 GNDA 0.023714f
C140 bgr_0.V_CUR_REF_REG.n2 GNDA 0.024034f
C141 bgr_0.V_CUR_REF_REG.n3 GNDA 0.231183f
C142 bgr_0.V_CUR_REF_REG.n4 GNDA 0.01997f
C143 bgr_0.V_CUR_REF_REG.n5 GNDA 1.47498f
C144 bgr_0.V_CUR_REF_REG.t0 GNDA 0.42777f
C145 VIN+.t0 GNDA 0.041803f
C146 VIN+.t10 GNDA 0.041803f
C147 VIN+.n0 GNDA 0.086391f
C148 VIN+.t6 GNDA 0.041803f
C149 VIN+.t8 GNDA 0.041803f
C150 VIN+.n1 GNDA 0.085194f
C151 VIN+.n2 GNDA 0.359761f
C152 VIN+.t4 GNDA 0.058811f
C153 VIN+.n3 GNDA 0.215335f
C154 VIN+.t3 GNDA 0.058811f
C155 VIN+.n4 GNDA 0.262589f
C156 VIN+.t1 GNDA 0.041803f
C157 VIN+.t7 GNDA 0.041803f
C158 VIN+.n5 GNDA 0.085194f
C159 VIN+.n6 GNDA 0.248358f
C160 VIN+.t2 GNDA 0.041803f
C161 VIN+.t9 GNDA 0.041803f
C162 VIN+.n7 GNDA 0.085194f
C163 VIN+.n8 GNDA 0.200956f
C164 VIN+.t5 GNDA 0.058811f
C165 VIN+.n9 GNDA 0.211601f
C166 two_stage_opamp_dummy_magic_0.VD4.t19 GNDA 0.024416f
C167 two_stage_opamp_dummy_magic_0.VD4.n0 GNDA 0.069509f
C168 two_stage_opamp_dummy_magic_0.VD4.n1 GNDA 0.094519f
C169 two_stage_opamp_dummy_magic_0.VD4.t27 GNDA 0.120449f
C170 two_stage_opamp_dummy_magic_0.VD4.t25 GNDA 0.042516f
C171 two_stage_opamp_dummy_magic_0.VD4.n2 GNDA 0.078578f
C172 two_stage_opamp_dummy_magic_0.VD4.n3 GNDA 0.050655f
C173 two_stage_opamp_dummy_magic_0.VD4.t24 GNDA 0.120449f
C174 two_stage_opamp_dummy_magic_0.VD4.t22 GNDA 0.042516f
C175 two_stage_opamp_dummy_magic_0.VD4.n4 GNDA 0.078578f
C176 two_stage_opamp_dummy_magic_0.VD4.n5 GNDA 0.050655f
C177 two_stage_opamp_dummy_magic_0.VD4.n6 GNDA 0.050227f
C178 two_stage_opamp_dummy_magic_0.VD4.n7 GNDA 0.094519f
C179 two_stage_opamp_dummy_magic_0.VD4.n8 GNDA 0.281683f
C180 two_stage_opamp_dummy_magic_0.VD4.t23 GNDA 0.420453f
C181 two_stage_opamp_dummy_magic_0.VD4.t2 GNDA 0.242764f
C182 two_stage_opamp_dummy_magic_0.VD4.t8 GNDA 0.242764f
C183 two_stage_opamp_dummy_magic_0.VD4.t16 GNDA 0.242764f
C184 two_stage_opamp_dummy_magic_0.VD4.t12 GNDA 0.242764f
C185 two_stage_opamp_dummy_magic_0.VD4.t18 GNDA 0.182073f
C186 two_stage_opamp_dummy_magic_0.VD4.n9 GNDA 0.121382f
C187 two_stage_opamp_dummy_magic_0.VD4.t20 GNDA 0.182073f
C188 two_stage_opamp_dummy_magic_0.VD4.t4 GNDA 0.242764f
C189 two_stage_opamp_dummy_magic_0.VD4.t10 GNDA 0.242764f
C190 two_stage_opamp_dummy_magic_0.VD4.t6 GNDA 0.242764f
C191 two_stage_opamp_dummy_magic_0.VD4.t14 GNDA 0.242764f
C192 two_stage_opamp_dummy_magic_0.VD4.t26 GNDA 0.420453f
C193 two_stage_opamp_dummy_magic_0.VD4.n10 GNDA 0.281683f
C194 two_stage_opamp_dummy_magic_0.VD4.n11 GNDA 0.069509f
C195 two_stage_opamp_dummy_magic_0.VD4.n12 GNDA 0.097309f
C196 two_stage_opamp_dummy_magic_0.VD4.t3 GNDA 0.024416f
C197 two_stage_opamp_dummy_magic_0.VD4.t9 GNDA 0.024416f
C198 two_stage_opamp_dummy_magic_0.VD4.n13 GNDA 0.084727f
C199 two_stage_opamp_dummy_magic_0.VD4.t0 GNDA 0.024416f
C200 two_stage_opamp_dummy_magic_0.VD4.t28 GNDA 0.024416f
C201 two_stage_opamp_dummy_magic_0.VD4.n14 GNDA 0.084913f
C202 two_stage_opamp_dummy_magic_0.VD4.t34 GNDA 0.024416f
C203 two_stage_opamp_dummy_magic_0.VD4.t1 GNDA 0.024416f
C204 two_stage_opamp_dummy_magic_0.VD4.n15 GNDA 0.084913f
C205 two_stage_opamp_dummy_magic_0.VD4.t32 GNDA 0.024416f
C206 two_stage_opamp_dummy_magic_0.VD4.t30 GNDA 0.024416f
C207 two_stage_opamp_dummy_magic_0.VD4.n16 GNDA 0.084613f
C208 two_stage_opamp_dummy_magic_0.VD4.n17 GNDA 0.15974f
C209 two_stage_opamp_dummy_magic_0.VD4.t37 GNDA 0.024416f
C210 two_stage_opamp_dummy_magic_0.VD4.t29 GNDA 0.024416f
C211 two_stage_opamp_dummy_magic_0.VD4.n18 GNDA 0.084613f
C212 two_stage_opamp_dummy_magic_0.VD4.n19 GNDA 0.082811f
C213 two_stage_opamp_dummy_magic_0.VD4.t33 GNDA 0.024416f
C214 two_stage_opamp_dummy_magic_0.VD4.t36 GNDA 0.024416f
C215 two_stage_opamp_dummy_magic_0.VD4.n20 GNDA 0.084613f
C216 two_stage_opamp_dummy_magic_0.VD4.n21 GNDA 0.082811f
C217 two_stage_opamp_dummy_magic_0.VD4.n22 GNDA 0.099252f
C218 two_stage_opamp_dummy_magic_0.VD4.t31 GNDA 0.024416f
C219 two_stage_opamp_dummy_magic_0.VD4.t35 GNDA 0.024416f
C220 two_stage_opamp_dummy_magic_0.VD4.n23 GNDA 0.08286f
C221 two_stage_opamp_dummy_magic_0.VD4.n24 GNDA 0.100481f
C222 two_stage_opamp_dummy_magic_0.VD4.n25 GNDA 0.094683f
C223 two_stage_opamp_dummy_magic_0.VD4.t17 GNDA 0.024416f
C224 two_stage_opamp_dummy_magic_0.VD4.t13 GNDA 0.024416f
C225 two_stage_opamp_dummy_magic_0.VD4.n26 GNDA 0.084612f
C226 two_stage_opamp_dummy_magic_0.VD4.n27 GNDA 0.078625f
C227 two_stage_opamp_dummy_magic_0.VD4.t7 GNDA 0.024416f
C228 two_stage_opamp_dummy_magic_0.VD4.t15 GNDA 0.024416f
C229 two_stage_opamp_dummy_magic_0.VD4.n28 GNDA 0.084913f
C230 two_stage_opamp_dummy_magic_0.VD4.t5 GNDA 0.024416f
C231 two_stage_opamp_dummy_magic_0.VD4.t11 GNDA 0.024416f
C232 two_stage_opamp_dummy_magic_0.VD4.n29 GNDA 0.084612f
C233 two_stage_opamp_dummy_magic_0.VD4.n30 GNDA 0.15974f
C234 two_stage_opamp_dummy_magic_0.VD4.n31 GNDA 0.029845f
C235 two_stage_opamp_dummy_magic_0.VD4.n32 GNDA 0.057972f
C236 two_stage_opamp_dummy_magic_0.VD4.n33 GNDA 0.079606f
C237 two_stage_opamp_dummy_magic_0.VD4.t21 GNDA 0.024416f
C238 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 GNDA 0.418194f
C239 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA 0.100765f
C240 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 GNDA 0.100765f
C241 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 GNDA 0.416703f
C242 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA 0.100765f
C243 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 GNDA 0.100765f
C244 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 GNDA 0.415104f
C245 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 GNDA 0.575542f
C246 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 GNDA 0.100765f
C247 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 GNDA 0.100765f
C248 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 GNDA 0.415104f
C249 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 GNDA 0.300326f
C250 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 GNDA 0.100765f
C251 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 GNDA 0.100765f
C252 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 GNDA 0.415104f
C253 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 GNDA 0.300326f
C254 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 GNDA 0.100765f
C255 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 GNDA 0.100765f
C256 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 GNDA 0.415104f
C257 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 GNDA 0.431646f
C258 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 GNDA 5.28083f
C259 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 GNDA 0.033588f
C260 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 GNDA 0.033588f
C261 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 GNDA 0.122084f
C262 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 GNDA 0.033588f
C263 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 GNDA 0.033588f
C264 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 GNDA 0.101451f
C265 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 GNDA 0.634217f
C266 bgr_0.V_CMFB_S2 GNDA 4.31626f
C267 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 GNDA 0.027366f
C268 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 GNDA 0.027366f
C269 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 GNDA 0.066f
C270 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 GNDA 0.027366f
C271 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 GNDA 0.027366f
C272 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 GNDA 0.068505f
C273 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 GNDA 0.027366f
C274 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 GNDA 0.027366f
C275 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 GNDA 0.068137f
C276 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 GNDA 0.462666f
C277 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 GNDA 0.027366f
C278 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 GNDA 0.027366f
C279 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 GNDA 0.068505f
C280 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 GNDA 0.303668f
C281 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 GNDA 0.704212f
C282 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 GNDA 0.041049f
C283 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 GNDA 0.041049f
C284 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 GNDA 0.148551f
C285 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 GNDA 0.072861f
C286 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 GNDA 0.072861f
C287 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 GNDA 0.072861f
C288 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 GNDA 0.072861f
C289 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 GNDA 0.072861f
C290 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 GNDA 0.072861f
C291 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 GNDA 0.072861f
C292 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 GNDA 0.085041f
C293 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 GNDA 0.08018f
C294 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 GNDA 0.050284f
C295 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 GNDA 0.050284f
C296 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 GNDA 0.050284f
C297 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 GNDA 0.050284f
C298 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 GNDA 0.050284f
C299 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 GNDA 0.044933f
C300 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 GNDA 0.072861f
C301 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 GNDA 0.072861f
C302 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 GNDA 0.072861f
C303 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 GNDA 0.072861f
C304 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 GNDA 0.072861f
C305 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 GNDA 0.072861f
C306 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 GNDA 0.072861f
C307 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 GNDA 0.072861f
C308 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 GNDA 0.072861f
C309 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 GNDA 0.072861f
C310 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 GNDA 0.072861f
C311 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 GNDA 0.085041f
C312 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 GNDA 0.08018f
C313 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 GNDA 0.050284f
C314 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 GNDA 0.050284f
C315 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 GNDA 0.050284f
C316 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 GNDA 0.050284f
C317 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 GNDA 0.050284f
C318 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 GNDA 0.050284f
C319 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 GNDA 0.050284f
C320 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 GNDA 0.050284f
C321 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 GNDA 0.050284f
C322 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 GNDA 0.044933f
C323 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 GNDA 0.112294f
C324 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 GNDA 0.041049f
C325 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 GNDA 0.041049f
C326 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 GNDA 0.082097f
C327 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 GNDA 0.318224f
C328 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 GNDA 3.34383f
C329 bgr_0.TAIL_CUR_MIR_BIAS GNDA 3.53441f
C330 two_stage_opamp_dummy_magic_0.V_p.t36 GNDA 0.014624f
C331 two_stage_opamp_dummy_magic_0.V_p.t19 GNDA 0.014624f
C332 two_stage_opamp_dummy_magic_0.V_p.t3 GNDA 0.014624f
C333 two_stage_opamp_dummy_magic_0.V_p.n0 GNDA 0.052539f
C334 two_stage_opamp_dummy_magic_0.V_p.t12 GNDA 0.014624f
C335 two_stage_opamp_dummy_magic_0.V_p.t20 GNDA 0.014624f
C336 two_stage_opamp_dummy_magic_0.V_p.n1 GNDA 0.052133f
C337 two_stage_opamp_dummy_magic_0.V_p.n2 GNDA 0.176305f
C338 two_stage_opamp_dummy_magic_0.V_p.t16 GNDA 0.014624f
C339 two_stage_opamp_dummy_magic_0.V_p.t34 GNDA 0.014624f
C340 two_stage_opamp_dummy_magic_0.V_p.n3 GNDA 0.052516f
C341 two_stage_opamp_dummy_magic_0.V_p.t8 GNDA 0.014624f
C342 two_stage_opamp_dummy_magic_0.V_p.t21 GNDA 0.014624f
C343 two_stage_opamp_dummy_magic_0.V_p.n4 GNDA 0.052133f
C344 two_stage_opamp_dummy_magic_0.V_p.n5 GNDA 0.174572f
C345 two_stage_opamp_dummy_magic_0.V_p.t24 GNDA 0.014624f
C346 two_stage_opamp_dummy_magic_0.V_p.t15 GNDA 0.014624f
C347 two_stage_opamp_dummy_magic_0.V_p.n6 GNDA 0.052133f
C348 two_stage_opamp_dummy_magic_0.V_p.n7 GNDA 0.091767f
C349 two_stage_opamp_dummy_magic_0.V_p.t26 GNDA 0.014624f
C350 two_stage_opamp_dummy_magic_0.V_p.t23 GNDA 0.014624f
C351 two_stage_opamp_dummy_magic_0.V_p.n8 GNDA 0.052133f
C352 two_stage_opamp_dummy_magic_0.V_p.n9 GNDA 0.091767f
C353 two_stage_opamp_dummy_magic_0.V_p.t18 GNDA 0.014624f
C354 two_stage_opamp_dummy_magic_0.V_p.t4 GNDA 0.014624f
C355 two_stage_opamp_dummy_magic_0.V_p.n10 GNDA 0.052133f
C356 two_stage_opamp_dummy_magic_0.V_p.n11 GNDA 0.140027f
C357 two_stage_opamp_dummy_magic_0.V_p.t17 GNDA 0.014624f
C358 two_stage_opamp_dummy_magic_0.V_p.t5 GNDA 0.014624f
C359 two_stage_opamp_dummy_magic_0.V_p.n12 GNDA 0.049685f
C360 two_stage_opamp_dummy_magic_0.V_p.t38 GNDA 0.024373f
C361 two_stage_opamp_dummy_magic_0.V_p.t37 GNDA 0.024373f
C362 two_stage_opamp_dummy_magic_0.V_p.n13 GNDA 0.099127f
C363 two_stage_opamp_dummy_magic_0.V_p.t2 GNDA 0.024373f
C364 two_stage_opamp_dummy_magic_0.V_p.t1 GNDA 0.024373f
C365 two_stage_opamp_dummy_magic_0.V_p.n14 GNDA 0.097223f
C366 two_stage_opamp_dummy_magic_0.V_p.t35 GNDA 0.024373f
C367 two_stage_opamp_dummy_magic_0.V_p.t6 GNDA 0.024373f
C368 two_stage_opamp_dummy_magic_0.V_p.n15 GNDA 0.096773f
C369 two_stage_opamp_dummy_magic_0.V_p.n16 GNDA 0.165755f
C370 two_stage_opamp_dummy_magic_0.V_p.t40 GNDA 0.024373f
C371 two_stage_opamp_dummy_magic_0.V_p.t31 GNDA 0.024373f
C372 two_stage_opamp_dummy_magic_0.V_p.n17 GNDA 0.096773f
C373 two_stage_opamp_dummy_magic_0.V_p.n18 GNDA 0.086515f
C374 two_stage_opamp_dummy_magic_0.V_p.t29 GNDA 0.085877f
C375 two_stage_opamp_dummy_magic_0.V_p.t27 GNDA 0.024373f
C376 two_stage_opamp_dummy_magic_0.V_p.t10 GNDA 0.024373f
C377 two_stage_opamp_dummy_magic_0.V_p.n19 GNDA 0.094049f
C378 two_stage_opamp_dummy_magic_0.V_p.n20 GNDA 0.56785f
C379 two_stage_opamp_dummy_magic_0.V_p.n21 GNDA 0.029248f
C380 two_stage_opamp_dummy_magic_0.V_p.t28 GNDA 0.024373f
C381 two_stage_opamp_dummy_magic_0.V_p.t32 GNDA 0.024373f
C382 two_stage_opamp_dummy_magic_0.V_p.n22 GNDA 0.096773f
C383 two_stage_opamp_dummy_magic_0.V_p.n23 GNDA 0.086515f
C384 two_stage_opamp_dummy_magic_0.V_p.t11 GNDA 0.024373f
C385 two_stage_opamp_dummy_magic_0.V_p.t7 GNDA 0.024373f
C386 two_stage_opamp_dummy_magic_0.V_p.n24 GNDA 0.096773f
C387 two_stage_opamp_dummy_magic_0.V_p.n25 GNDA 0.086515f
C388 two_stage_opamp_dummy_magic_0.V_p.t30 GNDA 0.024373f
C389 two_stage_opamp_dummy_magic_0.V_p.t9 GNDA 0.024373f
C390 two_stage_opamp_dummy_magic_0.V_p.n26 GNDA 0.096773f
C391 two_stage_opamp_dummy_magic_0.V_p.n27 GNDA 0.086515f
C392 two_stage_opamp_dummy_magic_0.V_p.t33 GNDA 0.024373f
C393 two_stage_opamp_dummy_magic_0.V_p.t39 GNDA 0.024373f
C394 two_stage_opamp_dummy_magic_0.V_p.n28 GNDA 0.096773f
C395 two_stage_opamp_dummy_magic_0.V_p.n29 GNDA 0.086515f
C396 two_stage_opamp_dummy_magic_0.V_p.n30 GNDA 0.159231f
C397 two_stage_opamp_dummy_magic_0.V_p.t14 GNDA 0.024373f
C398 two_stage_opamp_dummy_magic_0.V_p.t0 GNDA 0.024373f
C399 two_stage_opamp_dummy_magic_0.V_p.n31 GNDA 0.094049f
C400 two_stage_opamp_dummy_magic_0.V_p.n32 GNDA 0.078027f
C401 two_stage_opamp_dummy_magic_0.V_p.n33 GNDA 0.082224f
C402 two_stage_opamp_dummy_magic_0.V_p.n34 GNDA 0.07702f
C403 two_stage_opamp_dummy_magic_0.V_p.t13 GNDA 0.014624f
C404 two_stage_opamp_dummy_magic_0.V_p.t22 GNDA 0.014624f
C405 two_stage_opamp_dummy_magic_0.V_p.n35 GNDA 0.052133f
C406 two_stage_opamp_dummy_magic_0.V_p.n36 GNDA 0.09128f
C407 two_stage_opamp_dummy_magic_0.V_p.n37 GNDA 0.091767f
C408 two_stage_opamp_dummy_magic_0.V_p.n38 GNDA 0.052133f
C409 two_stage_opamp_dummy_magic_0.V_p.t25 GNDA 0.014624f
C410 VIN-.t6 GNDA 0.050642f
C411 VIN-.t5 GNDA 0.033412f
C412 VIN-.t0 GNDA 0.041251f
C413 VIN-.n0 GNDA 0.059274f
C414 VIN-.n1 GNDA 0.280478f
C415 VIN-.t3 GNDA 0.032863f
C416 VIN-.t9 GNDA 0.041265f
C417 VIN-.n2 GNDA 0.064892f
C418 VIN-.n3 GNDA 0.200879f
C419 VIN-.t8 GNDA 0.050078f
C420 VIN-.n4 GNDA 0.236241f
C421 VIN-.t7 GNDA 0.050425f
C422 VIN-.n5 GNDA 0.180621f
C423 VIN-.t2 GNDA 0.033412f
C424 VIN-.t1 GNDA 0.041251f
C425 VIN-.n6 GNDA 0.059274f
C426 VIN-.n7 GNDA 0.149629f
C427 VIN-.t4 GNDA 0.032863f
C428 VIN-.t10 GNDA 0.041265f
C429 VIN-.n8 GNDA 0.064892f
C430 VIN-.n9 GNDA 0.186141f
C431 bgr_0.cap_res2.t6 GNDA 0.406156f
C432 bgr_0.cap_res2.t2 GNDA 0.407628f
C433 bgr_0.cap_res2.t8 GNDA 0.406156f
C434 bgr_0.cap_res2.t13 GNDA 0.407628f
C435 bgr_0.cap_res2.t0 GNDA 0.406156f
C436 bgr_0.cap_res2.t19 GNDA 0.407628f
C437 bgr_0.cap_res2.t1 GNDA 0.406156f
C438 bgr_0.cap_res2.t5 GNDA 0.407628f
C439 bgr_0.cap_res2.t7 GNDA 0.406156f
C440 bgr_0.cap_res2.t4 GNDA 0.407628f
C441 bgr_0.cap_res2.t10 GNDA 0.406156f
C442 bgr_0.cap_res2.t14 GNDA 0.407628f
C443 bgr_0.cap_res2.t15 GNDA 0.406156f
C444 bgr_0.cap_res2.t12 GNDA 0.407628f
C445 bgr_0.cap_res2.t16 GNDA 0.406156f
C446 bgr_0.cap_res2.t18 GNDA 0.407628f
C447 bgr_0.cap_res2.n0 GNDA 0.272247f
C448 bgr_0.cap_res2.t17 GNDA 0.216805f
C449 bgr_0.cap_res2.n1 GNDA 0.295394f
C450 bgr_0.cap_res2.t11 GNDA 0.216805f
C451 bgr_0.cap_res2.n2 GNDA 0.295394f
C452 bgr_0.cap_res2.t3 GNDA 0.216805f
C453 bgr_0.cap_res2.n3 GNDA 0.295394f
C454 bgr_0.cap_res2.t9 GNDA 0.214043f
C455 bgr_0.cap_res2.t20 GNDA 0.133038f
C456 bgr_0.1st_Vout_2.n0 GNDA 0.995956f
C457 bgr_0.1st_Vout_2.n1 GNDA 0.240335f
C458 bgr_0.1st_Vout_2.n2 GNDA 0.995956f
C459 bgr_0.1st_Vout_2.n3 GNDA 0.240335f
C460 bgr_0.1st_Vout_2.n4 GNDA 0.805677f
C461 bgr_0.1st_Vout_2.n5 GNDA 0.240335f
C462 bgr_0.1st_Vout_2.t13 GNDA 0.021508f
C463 bgr_0.1st_Vout_2.n6 GNDA 0.02259f
C464 bgr_0.1st_Vout_2.n7 GNDA 0.171874f
C465 bgr_0.1st_Vout_2.t32 GNDA 0.013652f
C466 bgr_0.1st_Vout_2.t19 GNDA 0.013652f
C467 bgr_0.1st_Vout_2.n8 GNDA 0.03037f
C468 bgr_0.1st_Vout_2.n9 GNDA 0.083918f
C469 bgr_0.1st_Vout_2.n10 GNDA 0.012945f
C470 bgr_0.1st_Vout_2.t1 GNDA 0.018875f
C471 bgr_0.1st_Vout_2.n11 GNDA 0.195802f
C472 bgr_0.1st_Vout_2.n12 GNDA 0.011712f
C473 bgr_0.1st_Vout_2.n13 GNDA 0.049674f
C474 bgr_0.1st_Vout_2.n14 GNDA 0.021654f
C475 bgr_0.1st_Vout_2.n15 GNDA 0.080059f
C476 bgr_0.1st_Vout_2.n16 GNDA 0.03943f
C477 bgr_0.1st_Vout_2.t36 GNDA 0.013652f
C478 bgr_0.1st_Vout_2.t26 GNDA 0.013652f
C479 bgr_0.1st_Vout_2.n17 GNDA 0.03037f
C480 bgr_0.1st_Vout_2.n18 GNDA 0.083918f
C481 bgr_0.1st_Vout_2.t17 GNDA 0.364565f
C482 bgr_0.1st_Vout_2.t21 GNDA 0.358459f
C483 bgr_0.1st_Vout_2.t15 GNDA 0.358459f
C484 bgr_0.1st_Vout_2.t16 GNDA 0.364565f
C485 bgr_0.1st_Vout_2.t12 GNDA 0.358459f
C486 bgr_0.1st_Vout_2.t27 GNDA 0.364565f
C487 bgr_0.1st_Vout_2.t30 GNDA 0.358459f
C488 bgr_0.1st_Vout_2.t22 GNDA 0.358459f
C489 bgr_0.1st_Vout_2.t23 GNDA 0.364565f
C490 bgr_0.1st_Vout_2.t18 GNDA 0.358459f
C491 bgr_0.1st_Vout_2.t35 GNDA 0.364565f
C492 bgr_0.1st_Vout_2.t11 GNDA 0.358459f
C493 bgr_0.1st_Vout_2.t31 GNDA 0.358459f
C494 bgr_0.1st_Vout_2.t34 GNDA 0.364565f
C495 bgr_0.1st_Vout_2.t29 GNDA 0.358459f
C496 bgr_0.1st_Vout_2.t28 GNDA 0.364565f
C497 bgr_0.1st_Vout_2.t33 GNDA 0.358459f
C498 bgr_0.1st_Vout_2.t24 GNDA 0.358459f
C499 bgr_0.1st_Vout_2.t20 GNDA 0.358459f
C500 bgr_0.1st_Vout_2.t25 GNDA 0.358459f
C501 bgr_0.1st_Vout_2.t14 GNDA 0.023417f
C502 bgr_0.1st_Vout_2.n19 GNDA 0.516024f
C503 bgr_0.1st_Vout_2.n20 GNDA 0.106455f
C504 bgr_0.1st_Vout_2.n21 GNDA 0.02259f
C505 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA 0.092891f
C506 two_stage_opamp_dummy_magic_0.V_tot.t6 GNDA 0.011218f
C507 two_stage_opamp_dummy_magic_0.V_tot.n0 GNDA 0.018267f
C508 two_stage_opamp_dummy_magic_0.V_tot.n1 GNDA 0.106822f
C509 two_stage_opamp_dummy_magic_0.V_tot.n2 GNDA 0.021464f
C510 two_stage_opamp_dummy_magic_0.V_tot.n3 GNDA 0.095301f
C511 two_stage_opamp_dummy_magic_0.V_tot.t4 GNDA 0.011144f
C512 two_stage_opamp_dummy_magic_0.V_tot.n4 GNDA 0.091464f
C513 two_stage_opamp_dummy_magic_0.V_tot.n5 GNDA 0.021464f
C514 two_stage_opamp_dummy_magic_0.V_tot.n6 GNDA 0.066547f
C515 two_stage_opamp_dummy_magic_0.V_tot.n7 GNDA 0.021464f
C516 two_stage_opamp_dummy_magic_0.V_tot.n8 GNDA 0.204094f
C517 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA 0.098951f
C518 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA 0.092891f
C519 two_stage_opamp_dummy_magic_0.V_tot.n9 GNDA 0.321853f
C520 two_stage_opamp_dummy_magic_0.V_tot.n10 GNDA 0.772935f
C521 two_stage_opamp_dummy_magic_0.V_tot.n11 GNDA 0.513063f
C522 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA 0.098962f
C523 bgr_0.Vin+.t6 GNDA 0.020459f
C524 bgr_0.Vin+.t8 GNDA 0.013299f
C525 bgr_0.Vin+.n0 GNDA 0.04388f
C526 bgr_0.Vin+.t10 GNDA 0.013299f
C527 bgr_0.Vin+.n1 GNDA 0.034146f
C528 bgr_0.Vin+.t7 GNDA 0.013299f
C529 bgr_0.Vin+.n2 GNDA 0.034607f
C530 bgr_0.Vin+.n3 GNDA 0.074523f
C531 bgr_0.Vin+.t4 GNDA 0.043132f
C532 bgr_0.Vin+.t3 GNDA 0.043132f
C533 bgr_0.Vin+.n4 GNDA 0.144858f
C534 bgr_0.Vin+.t2 GNDA 0.043132f
C535 bgr_0.Vin+.t5 GNDA 0.043132f
C536 bgr_0.Vin+.n5 GNDA 0.142495f
C537 bgr_0.Vin+.n6 GNDA 0.656763f
C538 bgr_0.Vin+.n7 GNDA 0.71769f
C539 bgr_0.Vin+.t1 GNDA 0.125873f
C540 bgr_0.Vin+.n8 GNDA 0.446219f
C541 bgr_0.Vin+.t0 GNDA 0.137433f
C542 two_stage_opamp_dummy_magic_0.V_err_p.n0 GNDA 0.02127f
C543 two_stage_opamp_dummy_magic_0.V_err_p.n1 GNDA 0.020358f
C544 two_stage_opamp_dummy_magic_0.V_err_p.n2 GNDA 0.020407f
C545 two_stage_opamp_dummy_magic_0.V_err_p.n3 GNDA 0.021244f
C546 two_stage_opamp_dummy_magic_0.V_err_p.n4 GNDA 0.021116f
C547 two_stage_opamp_dummy_magic_0.V_err_p.n5 GNDA 0.299998f
C548 two_stage_opamp_dummy_magic_0.V_err_p.n6 GNDA 0.021116f
C549 two_stage_opamp_dummy_magic_0.V_err_p.n7 GNDA 0.156484f
C550 two_stage_opamp_dummy_magic_0.V_err_p.n8 GNDA 0.021116f
C551 two_stage_opamp_dummy_magic_0.V_err_p.n9 GNDA 0.190977f
C552 two_stage_opamp_dummy_magic_0.V_err_p.n10 GNDA 0.153542f
C553 two_stage_opamp_dummy_magic_0.V_err_p.n11 GNDA 0.133374f
C554 two_stage_opamp_dummy_magic_0.V_err_p.n12 GNDA 0.242929f
C555 two_stage_opamp_dummy_magic_0.V_err_p.n13 GNDA 0.02127f
C556 two_stage_opamp_dummy_magic_0.V_err_p.n14 GNDA 0.020976f
C557 two_stage_opamp_dummy_magic_0.V_err_p.n15 GNDA 0.328367f
C558 two_stage_opamp_dummy_magic_0.V_err_p.n16 GNDA 0.020976f
C559 two_stage_opamp_dummy_magic_0.V_err_p.n17 GNDA 0.180843f
C560 two_stage_opamp_dummy_magic_0.V_err_p.n18 GNDA 0.180843f
C561 two_stage_opamp_dummy_magic_0.V_err_p.n19 GNDA 0.020976f
C562 bgr_0.VB3_CUR_BIAS GNDA 6.0158f
C563 two_stage_opamp_dummy_magic_0.Vb3.t1 GNDA 0.034262f
C564 two_stage_opamp_dummy_magic_0.Vb3.t4 GNDA 0.034262f
C565 two_stage_opamp_dummy_magic_0.Vb3.n0 GNDA 0.103485f
C566 two_stage_opamp_dummy_magic_0.Vb3.t5 GNDA 0.034262f
C567 two_stage_opamp_dummy_magic_0.Vb3.t3 GNDA 0.034262f
C568 two_stage_opamp_dummy_magic_0.Vb3.n1 GNDA 0.11036f
C569 two_stage_opamp_dummy_magic_0.Vb3.t2 GNDA 0.034262f
C570 two_stage_opamp_dummy_magic_0.Vb3.t6 GNDA 0.034262f
C571 two_stage_opamp_dummy_magic_0.Vb3.n2 GNDA 0.11036f
C572 two_stage_opamp_dummy_magic_0.Vb3.n3 GNDA 0.608411f
C573 two_stage_opamp_dummy_magic_0.Vb3.n4 GNDA 0.22714f
C574 two_stage_opamp_dummy_magic_0.Vb3.t14 GNDA 0.169595f
C575 two_stage_opamp_dummy_magic_0.Vb3.t18 GNDA 0.169595f
C576 two_stage_opamp_dummy_magic_0.Vb3.t15 GNDA 0.169595f
C577 two_stage_opamp_dummy_magic_0.Vb3.t21 GNDA 0.169595f
C578 two_stage_opamp_dummy_magic_0.Vb3.t26 GNDA 0.195711f
C579 two_stage_opamp_dummy_magic_0.Vb3.n5 GNDA 0.158896f
C580 two_stage_opamp_dummy_magic_0.Vb3.n6 GNDA 0.097646f
C581 two_stage_opamp_dummy_magic_0.Vb3.n7 GNDA 0.097646f
C582 two_stage_opamp_dummy_magic_0.Vb3.n8 GNDA 0.091432f
C583 two_stage_opamp_dummy_magic_0.Vb3.t12 GNDA 0.169595f
C584 two_stage_opamp_dummy_magic_0.Vb3.t25 GNDA 0.169595f
C585 two_stage_opamp_dummy_magic_0.Vb3.t20 GNDA 0.169595f
C586 two_stage_opamp_dummy_magic_0.Vb3.t22 GNDA 0.169595f
C587 two_stage_opamp_dummy_magic_0.Vb3.t17 GNDA 0.195711f
C588 two_stage_opamp_dummy_magic_0.Vb3.n9 GNDA 0.158896f
C589 two_stage_opamp_dummy_magic_0.Vb3.n10 GNDA 0.097646f
C590 two_stage_opamp_dummy_magic_0.Vb3.n11 GNDA 0.097646f
C591 two_stage_opamp_dummy_magic_0.Vb3.n12 GNDA 0.091432f
C592 two_stage_opamp_dummy_magic_0.Vb3.n13 GNDA 0.062373f
C593 two_stage_opamp_dummy_magic_0.Vb3.t0 GNDA 0.123342f
C594 two_stage_opamp_dummy_magic_0.Vb3.t7 GNDA 0.123342f
C595 two_stage_opamp_dummy_magic_0.Vb3.n14 GNDA 0.454379f
C596 two_stage_opamp_dummy_magic_0.Vb3.t16 GNDA 0.196517f
C597 two_stage_opamp_dummy_magic_0.Vb3.n15 GNDA 2.15298f
C598 two_stage_opamp_dummy_magic_0.Vb3.t19 GNDA 0.169595f
C599 two_stage_opamp_dummy_magic_0.Vb3.t24 GNDA 0.169595f
C600 two_stage_opamp_dummy_magic_0.Vb3.t28 GNDA 0.169595f
C601 two_stage_opamp_dummy_magic_0.Vb3.t9 GNDA 0.169595f
C602 two_stage_opamp_dummy_magic_0.Vb3.t11 GNDA 0.195711f
C603 two_stage_opamp_dummy_magic_0.Vb3.n16 GNDA 0.158896f
C604 two_stage_opamp_dummy_magic_0.Vb3.n17 GNDA 0.097646f
C605 two_stage_opamp_dummy_magic_0.Vb3.n18 GNDA 0.097646f
C606 two_stage_opamp_dummy_magic_0.Vb3.n19 GNDA 0.091432f
C607 two_stage_opamp_dummy_magic_0.Vb3.t13 GNDA 0.169595f
C608 two_stage_opamp_dummy_magic_0.Vb3.t10 GNDA 0.169595f
C609 two_stage_opamp_dummy_magic_0.Vb3.t8 GNDA 0.169595f
C610 two_stage_opamp_dummy_magic_0.Vb3.t27 GNDA 0.169595f
C611 two_stage_opamp_dummy_magic_0.Vb3.t23 GNDA 0.195711f
C612 two_stage_opamp_dummy_magic_0.Vb3.n20 GNDA 0.158896f
C613 two_stage_opamp_dummy_magic_0.Vb3.n21 GNDA 0.097646f
C614 two_stage_opamp_dummy_magic_0.Vb3.n22 GNDA 0.097646f
C615 two_stage_opamp_dummy_magic_0.Vb3.n23 GNDA 0.091432f
C616 two_stage_opamp_dummy_magic_0.Vb3.n24 GNDA 0.055211f
C617 two_stage_opamp_dummy_magic_0.Vb3.n25 GNDA 1.48367f
C618 two_stage_opamp_dummy_magic_0.Vb3.n26 GNDA 6.08823f
C619 two_stage_opamp_dummy_magic_0.Vb2.t15 GNDA 0.093589f
C620 two_stage_opamp_dummy_magic_0.Vb2.t19 GNDA 0.093589f
C621 two_stage_opamp_dummy_magic_0.Vb2.t17 GNDA 0.093589f
C622 two_stage_opamp_dummy_magic_0.Vb2.t22 GNDA 0.093589f
C623 two_stage_opamp_dummy_magic_0.Vb2.t27 GNDA 0.108001f
C624 two_stage_opamp_dummy_magic_0.Vb2.n0 GNDA 0.087685f
C625 two_stage_opamp_dummy_magic_0.Vb2.n1 GNDA 0.053884f
C626 two_stage_opamp_dummy_magic_0.Vb2.n2 GNDA 0.053884f
C627 two_stage_opamp_dummy_magic_0.Vb2.n3 GNDA 0.050455f
C628 two_stage_opamp_dummy_magic_0.Vb2.t13 GNDA 0.093589f
C629 two_stage_opamp_dummy_magic_0.Vb2.t26 GNDA 0.093589f
C630 two_stage_opamp_dummy_magic_0.Vb2.t21 GNDA 0.093589f
C631 two_stage_opamp_dummy_magic_0.Vb2.t23 GNDA 0.093589f
C632 two_stage_opamp_dummy_magic_0.Vb2.t18 GNDA 0.108001f
C633 two_stage_opamp_dummy_magic_0.Vb2.n4 GNDA 0.087685f
C634 two_stage_opamp_dummy_magic_0.Vb2.n5 GNDA 0.053884f
C635 two_stage_opamp_dummy_magic_0.Vb2.n6 GNDA 0.053884f
C636 two_stage_opamp_dummy_magic_0.Vb2.n7 GNDA 0.050455f
C637 two_stage_opamp_dummy_magic_0.Vb2.n8 GNDA 0.033749f
C638 two_stage_opamp_dummy_magic_0.Vb2.t20 GNDA 0.093589f
C639 two_stage_opamp_dummy_magic_0.Vb2.t25 GNDA 0.093589f
C640 two_stage_opamp_dummy_magic_0.Vb2.t29 GNDA 0.093589f
C641 two_stage_opamp_dummy_magic_0.Vb2.t31 GNDA 0.093589f
C642 two_stage_opamp_dummy_magic_0.Vb2.t12 GNDA 0.108001f
C643 two_stage_opamp_dummy_magic_0.Vb2.n9 GNDA 0.087685f
C644 two_stage_opamp_dummy_magic_0.Vb2.n10 GNDA 0.053884f
C645 two_stage_opamp_dummy_magic_0.Vb2.n11 GNDA 0.053884f
C646 two_stage_opamp_dummy_magic_0.Vb2.n12 GNDA 0.050455f
C647 two_stage_opamp_dummy_magic_0.Vb2.t14 GNDA 0.093589f
C648 two_stage_opamp_dummy_magic_0.Vb2.t11 GNDA 0.093589f
C649 two_stage_opamp_dummy_magic_0.Vb2.t30 GNDA 0.093589f
C650 two_stage_opamp_dummy_magic_0.Vb2.t28 GNDA 0.093589f
C651 two_stage_opamp_dummy_magic_0.Vb2.t24 GNDA 0.108001f
C652 two_stage_opamp_dummy_magic_0.Vb2.n13 GNDA 0.087685f
C653 two_stage_opamp_dummy_magic_0.Vb2.n14 GNDA 0.053884f
C654 two_stage_opamp_dummy_magic_0.Vb2.n15 GNDA 0.053884f
C655 two_stage_opamp_dummy_magic_0.Vb2.n16 GNDA 0.050455f
C656 two_stage_opamp_dummy_magic_0.Vb2.n17 GNDA 0.033749f
C657 two_stage_opamp_dummy_magic_0.Vb2.n18 GNDA 1.26875f
C658 two_stage_opamp_dummy_magic_0.Vb2.t6 GNDA 0.011911f
C659 two_stage_opamp_dummy_magic_0.Vb2.t10 GNDA 0.011911f
C660 two_stage_opamp_dummy_magic_0.Vb2.n19 GNDA 0.025812f
C661 two_stage_opamp_dummy_magic_0.Vb2.t9 GNDA 0.036993f
C662 two_stage_opamp_dummy_magic_0.Vb2.n20 GNDA 0.12548f
C663 two_stage_opamp_dummy_magic_0.Vb2.n21 GNDA 1.11042f
C664 two_stage_opamp_dummy_magic_0.Vb2.t16 GNDA 0.1131f
C665 two_stage_opamp_dummy_magic_0.Vb2.n22 GNDA 3.08838f
C666 two_stage_opamp_dummy_magic_0.Vb2.t8 GNDA 0.018907f
C667 two_stage_opamp_dummy_magic_0.Vb2.t0 GNDA 0.018907f
C668 two_stage_opamp_dummy_magic_0.Vb2.n23 GNDA 0.063392f
C669 two_stage_opamp_dummy_magic_0.Vb2.t3 GNDA 0.018907f
C670 two_stage_opamp_dummy_magic_0.Vb2.t1 GNDA 0.018907f
C671 two_stage_opamp_dummy_magic_0.Vb2.n24 GNDA 0.061653f
C672 two_stage_opamp_dummy_magic_0.Vb2.n25 GNDA 0.497935f
C673 two_stage_opamp_dummy_magic_0.Vb2.t5 GNDA 0.018907f
C674 two_stage_opamp_dummy_magic_0.Vb2.t7 GNDA 0.018907f
C675 two_stage_opamp_dummy_magic_0.Vb2.n26 GNDA 0.063392f
C676 two_stage_opamp_dummy_magic_0.Vb2.t4 GNDA 0.018907f
C677 two_stage_opamp_dummy_magic_0.Vb2.t2 GNDA 0.018907f
C678 two_stage_opamp_dummy_magic_0.Vb2.n27 GNDA 0.061653f
C679 two_stage_opamp_dummy_magic_0.Vb2.n28 GNDA 0.497935f
C680 two_stage_opamp_dummy_magic_0.Vb2.n29 GNDA 0.259717f
C681 bgr_0.VB2_CUR_BIAS GNDA 2.86975f
C682 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 GNDA 0.020233f
C683 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 GNDA 0.020233f
C684 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 GNDA 0.020233f
C685 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 GNDA 0.047731f
C686 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 GNDA 0.020233f
C687 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 GNDA 0.020233f
C688 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 GNDA 0.046922f
C689 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 GNDA 0.884615f
C690 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 GNDA 0.020233f
C691 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 GNDA 0.020233f
C692 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 GNDA 0.046922f
C693 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 GNDA 2.10658f
C694 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 GNDA 1.98101f
C695 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 GNDA 0.020233f
C696 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 GNDA 0.020233f
C697 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 GNDA 0.04777f
C698 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 GNDA 0.016692f
C699 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 GNDA 0.016692f
C700 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 GNDA 0.016692f
C701 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 GNDA 0.016692f
C702 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 GNDA 0.016692f
C703 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 GNDA 0.036166f
C704 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 GNDA 0.051623f
C705 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 GNDA 0.020233f
C706 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 GNDA 0.020233f
C707 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 GNDA 0.04777f
C708 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 GNDA 0.17992f
C709 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 GNDA 0.05811f
C710 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 GNDA 0.039231f
C711 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 GNDA 0.044006f
C712 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 GNDA 0.044006f
C713 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 GNDA 0.039231f
C714 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 GNDA 0.016692f
C715 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 GNDA 0.016692f
C716 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 GNDA 0.016692f
C717 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 GNDA 0.036166f
C718 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 GNDA 0.056399f
C719 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 GNDA 0.044006f
C720 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 GNDA 0.039231f
C721 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 GNDA 0.05811f
C722 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 GNDA 0.17992f
C723 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 GNDA 0.746838f
C724 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 GNDA 0.061393f
C725 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 GNDA 0.020233f
C726 two_stage_opamp_dummy_magic_0.VD3.t32 GNDA 0.03144f
C727 two_stage_opamp_dummy_magic_0.VD3.t30 GNDA 0.03144f
C728 two_stage_opamp_dummy_magic_0.VD3.n0 GNDA 0.10934f
C729 two_stage_opamp_dummy_magic_0.VD3.t20 GNDA 0.03144f
C730 two_stage_opamp_dummy_magic_0.VD3.t16 GNDA 0.03144f
C731 two_stage_opamp_dummy_magic_0.VD3.n1 GNDA 0.108953f
C732 two_stage_opamp_dummy_magic_0.VD3.n2 GNDA 0.205692f
C733 two_stage_opamp_dummy_magic_0.VD3.t37 GNDA 0.03144f
C734 two_stage_opamp_dummy_magic_0.VD3.t9 GNDA 0.03144f
C735 two_stage_opamp_dummy_magic_0.VD3.n3 GNDA 0.108953f
C736 two_stage_opamp_dummy_magic_0.VD3.n4 GNDA 0.106633f
C737 two_stage_opamp_dummy_magic_0.VD3.t36 GNDA 0.03144f
C738 two_stage_opamp_dummy_magic_0.VD3.t35 GNDA 0.03144f
C739 two_stage_opamp_dummy_magic_0.VD3.n5 GNDA 0.108953f
C740 two_stage_opamp_dummy_magic_0.VD3.n6 GNDA 0.106633f
C741 two_stage_opamp_dummy_magic_0.VD3.t6 GNDA 0.03144f
C742 two_stage_opamp_dummy_magic_0.VD3.t31 GNDA 0.03144f
C743 two_stage_opamp_dummy_magic_0.VD3.n7 GNDA 0.10934f
C744 two_stage_opamp_dummy_magic_0.VD3.n8 GNDA 0.127804f
C745 two_stage_opamp_dummy_magic_0.VD3.t19 GNDA 0.03144f
C746 two_stage_opamp_dummy_magic_0.VD3.t21 GNDA 0.03144f
C747 two_stage_opamp_dummy_magic_0.VD3.n9 GNDA 0.106696f
C748 two_stage_opamp_dummy_magic_0.VD3.n10 GNDA 0.089361f
C749 two_stage_opamp_dummy_magic_0.VD3.t27 GNDA 0.03144f
C750 two_stage_opamp_dummy_magic_0.VD3.t8 GNDA 0.03144f
C751 two_stage_opamp_dummy_magic_0.VD3.n11 GNDA 0.10934f
C752 two_stage_opamp_dummy_magic_0.VD3.t1 GNDA 0.03144f
C753 two_stage_opamp_dummy_magic_0.VD3.t25 GNDA 0.03144f
C754 two_stage_opamp_dummy_magic_0.VD3.n12 GNDA 0.108953f
C755 two_stage_opamp_dummy_magic_0.VD3.n13 GNDA 0.205693f
C756 two_stage_opamp_dummy_magic_0.VD3.n14 GNDA 0.089505f
C757 two_stage_opamp_dummy_magic_0.VD3.n15 GNDA 0.089505f
C758 two_stage_opamp_dummy_magic_0.VD3.n16 GNDA 0.362715f
C759 two_stage_opamp_dummy_magic_0.VD3.n17 GNDA 0.362715f
C760 two_stage_opamp_dummy_magic_0.VD3.t14 GNDA 0.541405f
C761 two_stage_opamp_dummy_magic_0.VD3.t26 GNDA 0.3126f
C762 two_stage_opamp_dummy_magic_0.VD3.t7 GNDA 0.3126f
C763 two_stage_opamp_dummy_magic_0.VD3.t0 GNDA 0.3126f
C764 two_stage_opamp_dummy_magic_0.VD3.t24 GNDA 0.3126f
C765 two_stage_opamp_dummy_magic_0.VD3.t17 GNDA 0.23445f
C766 two_stage_opamp_dummy_magic_0.VD3.t15 GNDA 0.155099f
C767 two_stage_opamp_dummy_magic_0.VD3.t13 GNDA 0.054747f
C768 two_stage_opamp_dummy_magic_0.VD3.n18 GNDA 0.101182f
C769 two_stage_opamp_dummy_magic_0.VD3.n19 GNDA 0.065226f
C770 two_stage_opamp_dummy_magic_0.VD3.t12 GNDA 0.155099f
C771 two_stage_opamp_dummy_magic_0.VD3.t10 GNDA 0.054747f
C772 two_stage_opamp_dummy_magic_0.VD3.n20 GNDA 0.101182f
C773 two_stage_opamp_dummy_magic_0.VD3.n21 GNDA 0.065226f
C774 two_stage_opamp_dummy_magic_0.VD3.n22 GNDA 0.064676f
C775 two_stage_opamp_dummy_magic_0.VD3.n23 GNDA 0.12171f
C776 two_stage_opamp_dummy_magic_0.VD3.t11 GNDA 0.541405f
C777 two_stage_opamp_dummy_magic_0.VD3.t22 GNDA 0.3126f
C778 two_stage_opamp_dummy_magic_0.VD3.t33 GNDA 0.3126f
C779 two_stage_opamp_dummy_magic_0.VD3.t4 GNDA 0.3126f
C780 two_stage_opamp_dummy_magic_0.VD3.t2 GNDA 0.3126f
C781 two_stage_opamp_dummy_magic_0.VD3.t28 GNDA 0.23445f
C782 two_stage_opamp_dummy_magic_0.VD3.n24 GNDA 0.1563f
C783 two_stage_opamp_dummy_magic_0.VD3.n25 GNDA 0.12171f
C784 two_stage_opamp_dummy_magic_0.VD3.n26 GNDA 0.125303f
C785 two_stage_opamp_dummy_magic_0.VD3.t18 GNDA 0.03144f
C786 two_stage_opamp_dummy_magic_0.VD3.t29 GNDA 0.03144f
C787 two_stage_opamp_dummy_magic_0.VD3.n27 GNDA 0.102506f
C788 two_stage_opamp_dummy_magic_0.VD3.n28 GNDA 0.074649f
C789 two_stage_opamp_dummy_magic_0.VD3.n29 GNDA 0.038431f
C790 two_stage_opamp_dummy_magic_0.VD3.t3 GNDA 0.03144f
C791 two_stage_opamp_dummy_magic_0.VD3.t5 GNDA 0.03144f
C792 two_stage_opamp_dummy_magic_0.VD3.n30 GNDA 0.108953f
C793 two_stage_opamp_dummy_magic_0.VD3.n31 GNDA 0.101243f
C794 two_stage_opamp_dummy_magic_0.VD3.t34 GNDA 0.03144f
C795 two_stage_opamp_dummy_magic_0.VD3.t23 GNDA 0.03144f
C796 two_stage_opamp_dummy_magic_0.VD3.n32 GNDA 0.1091f
C797 two_stage_opamp_dummy_magic_0.VD3.n33 GNDA 0.116136f
C798 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 GNDA 0.163765f
C799 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 GNDA 0.409099f
C800 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 GNDA 0.409099f
C801 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 GNDA 0.485537f
C802 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 GNDA 0.256456f
C803 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 GNDA 0.162306f
C804 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 GNDA 0.446073f
C805 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 GNDA 0.149996f
C806 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 GNDA 0.917914f
C807 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 GNDA 0.446073f
C808 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 GNDA 0.409099f
C809 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 GNDA 0.409099f
C810 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 GNDA 0.485537f
C811 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 GNDA 0.256456f
C812 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 GNDA 0.162306f
C813 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 GNDA 0.149996f
C814 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 GNDA 0.917423f
C815 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 GNDA 0.163765f
C816 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 GNDA 0.345114f
C817 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 GNDA 0.346365f
C818 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 GNDA 0.345114f
C819 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 GNDA 0.34782f
C820 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 GNDA 0.378304f
C821 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 GNDA 0.345114f
C822 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 GNDA 0.346365f
C823 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 GNDA 0.345114f
C824 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 GNDA 0.346365f
C825 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 GNDA 0.345114f
C826 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 GNDA 0.346365f
C827 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 GNDA 0.345114f
C828 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 GNDA 0.346365f
C829 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 GNDA 0.345114f
C830 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 GNDA 0.346365f
C831 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 GNDA 0.345114f
C832 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 GNDA 0.346365f
C833 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 GNDA 0.345114f
C834 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 GNDA 0.346365f
C835 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 GNDA 0.345114f
C836 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 GNDA 0.346365f
C837 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 GNDA 0.345114f
C838 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 GNDA 0.346365f
C839 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 GNDA 0.345114f
C840 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 GNDA 0.346365f
C841 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 GNDA 0.345114f
C842 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 GNDA 0.346365f
C843 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 GNDA 0.345114f
C844 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 GNDA 0.346365f
C845 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 GNDA 0.345114f
C846 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 GNDA 0.346365f
C847 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 GNDA 0.345114f
C848 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 GNDA 0.346365f
C849 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 GNDA 0.345114f
C850 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 GNDA 0.346365f
C851 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 GNDA 0.345114f
C852 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 GNDA 0.346365f
C853 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 GNDA 0.345114f
C854 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 GNDA 0.346365f
C855 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 GNDA 0.345114f
C856 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 GNDA 0.346365f
C857 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 GNDA 0.345114f
C858 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 GNDA 0.346365f
C859 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 GNDA 0.345114f
C860 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 GNDA 0.346365f
C861 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 GNDA 0.345114f
C862 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 GNDA 0.346365f
C863 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 GNDA 0.345114f
C864 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 GNDA 0.346365f
C865 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 GNDA 0.345114f
C866 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 GNDA 0.346365f
C867 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 GNDA 0.345114f
C868 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 GNDA 0.346365f
C869 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 GNDA 0.345114f
C870 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 GNDA 0.346365f
C871 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 GNDA 0.345114f
C872 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 GNDA 0.346365f
C873 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 GNDA 0.345114f
C874 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 GNDA 0.346365f
C875 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 GNDA 0.345114f
C876 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 GNDA 0.346365f
C877 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 GNDA 0.345114f
C878 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 GNDA 0.346365f
C879 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 GNDA 0.345114f
C880 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 GNDA 0.362035f
C881 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 GNDA 0.345114f
C882 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 GNDA 0.185368f
C883 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 GNDA 0.198389f
C884 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 GNDA 0.345114f
C885 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 GNDA 0.185368f
C886 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 GNDA 0.196789f
C887 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 GNDA 0.345114f
C888 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 GNDA 0.185368f
C889 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 GNDA 0.196789f
C890 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 GNDA 0.345114f
C891 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 GNDA 0.185368f
C892 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 GNDA 0.196789f
C893 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 GNDA 0.345114f
C894 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 GNDA 0.185368f
C895 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 GNDA 0.196789f
C896 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 GNDA 0.345114f
C897 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 GNDA 0.185368f
C898 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 GNDA 0.196789f
C899 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 GNDA 0.345114f
C900 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 GNDA 0.185368f
C901 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 GNDA 0.196789f
C902 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 GNDA 0.345114f
C903 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 GNDA 0.185368f
C904 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 GNDA 0.196789f
C905 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 GNDA 0.345114f
C906 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 GNDA 0.185368f
C907 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 GNDA 0.196789f
C908 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 GNDA 0.345114f
C909 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 GNDA 0.346365f
C910 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 GNDA 0.166846f
C911 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 GNDA 0.215207f
C912 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 GNDA 0.18422f
C913 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 GNDA 0.233728f
C914 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 GNDA 0.18422f
C915 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 GNDA 0.250999f
C916 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 GNDA 0.18422f
C917 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 GNDA 0.250999f
C918 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 GNDA 0.18422f
C919 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 GNDA 0.250999f
C920 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 GNDA 0.18422f
C921 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 GNDA 0.250999f
C922 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 GNDA 0.18422f
C923 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 GNDA 0.250999f
C924 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 GNDA 0.18422f
C925 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 GNDA 0.250999f
C926 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 GNDA 0.18422f
C927 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 GNDA 0.250999f
C928 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 GNDA 0.18422f
C929 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 GNDA 0.250999f
C930 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 GNDA 0.18422f
C931 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 GNDA 0.250999f
C932 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 GNDA 0.18422f
C933 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 GNDA 0.250999f
C934 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 GNDA 0.18422f
C935 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 GNDA 0.250999f
C936 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 GNDA 0.18422f
C937 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 GNDA 0.250999f
C938 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 GNDA 0.18422f
C939 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 GNDA 0.250999f
C940 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 GNDA 0.18422f
C941 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 GNDA 0.250999f
C942 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 GNDA 0.18422f
C943 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 GNDA 0.233728f
C944 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 GNDA 0.343967f
C945 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 GNDA 0.166846f
C946 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 GNDA 0.216458f
C947 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 GNDA 0.343967f
C948 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 GNDA 0.166846f
C949 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 GNDA 0.216458f
C950 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 GNDA 0.343967f
C951 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 GNDA 0.345114f
C952 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 GNDA 0.363635f
C953 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 GNDA 0.363635f
C954 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 GNDA 0.363635f
C955 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 GNDA 0.185368f
C956 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 GNDA 0.216458f
C957 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 GNDA 0.343967f
C958 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 GNDA 0.166846f
C959 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 GNDA 0.197936f
C960 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 GNDA 0.343967f
C961 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 GNDA 0.166846f
C962 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 GNDA 0.216458f
C963 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 GNDA 0.343967f
C964 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 GNDA 0.166846f
C965 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 GNDA 0.216458f
C966 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 GNDA 0.343967f
C967 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 GNDA 0.166846f
C968 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 GNDA 0.216458f
C969 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 GNDA 0.343967f
C970 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 GNDA 0.345114f
C971 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 GNDA 0.363635f
C972 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 GNDA 0.363635f
C973 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 GNDA 0.363635f
C974 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 GNDA 0.185368f
C975 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 GNDA 0.216458f
C976 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 GNDA 0.343967f
C977 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 GNDA 0.345114f
C978 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 GNDA 0.363635f
C979 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 GNDA 0.363635f
C980 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 GNDA 0.363635f
C981 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 GNDA 0.185368f
C982 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 GNDA 0.216458f
C983 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 GNDA 0.343967f
C984 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 GNDA 0.216458f
C985 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 GNDA 0.185368f
C986 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 GNDA 0.363635f
C987 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 GNDA 0.363635f
C988 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 GNDA 0.363635f
C989 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 GNDA 0.602274f
C990 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 GNDA 0.298233f
C991 VOUT+.t5 GNDA 0.043577f
C992 VOUT+.t18 GNDA 0.043577f
C993 VOUT+.n0 GNDA 0.175148f
C994 VOUT+.t13 GNDA 0.043577f
C995 VOUT+.t17 GNDA 0.043577f
C996 VOUT+.n1 GNDA 0.174825f
C997 VOUT+.n2 GNDA 0.172223f
C998 VOUT+.t12 GNDA 0.043577f
C999 VOUT+.t16 GNDA 0.043577f
C1000 VOUT+.n3 GNDA 0.174825f
C1001 VOUT+.n4 GNDA 0.088815f
C1002 VOUT+.t10 GNDA 0.043577f
C1003 VOUT+.t14 GNDA 0.043577f
C1004 VOUT+.n5 GNDA 0.174825f
C1005 VOUT+.n6 GNDA 0.088815f
C1006 VOUT+.t9 GNDA 0.043577f
C1007 VOUT+.t6 GNDA 0.043577f
C1008 VOUT+.n7 GNDA 0.175148f
C1009 VOUT+.n8 GNDA 0.105197f
C1010 VOUT+.t11 GNDA 0.043577f
C1011 VOUT+.t15 GNDA 0.043577f
C1012 VOUT+.n9 GNDA 0.172685f
C1013 VOUT+.n10 GNDA 0.210763f
C1014 VOUT+.t117 GNDA 0.295461f
C1015 VOUT+.t26 GNDA 0.290513f
C1016 VOUT+.n11 GNDA 0.194779f
C1017 VOUT+.t124 GNDA 0.290513f
C1018 VOUT+.n12 GNDA 0.127099f
C1019 VOUT+.t72 GNDA 0.295461f
C1020 VOUT+.t39 GNDA 0.290513f
C1021 VOUT+.n13 GNDA 0.194779f
C1022 VOUT+.t127 GNDA 0.290513f
C1023 VOUT+.t35 GNDA 0.294841f
C1024 VOUT+.t87 GNDA 0.294841f
C1025 VOUT+.t43 GNDA 0.294841f
C1026 VOUT+.t96 GNDA 0.294841f
C1027 VOUT+.t143 GNDA 0.294841f
C1028 VOUT+.t106 GNDA 0.294841f
C1029 VOUT+.t154 GNDA 0.294841f
C1030 VOUT+.t65 GNDA 0.294841f
C1031 VOUT+.t116 GNDA 0.294841f
C1032 VOUT+.t73 GNDA 0.294841f
C1033 VOUT+.t149 GNDA 0.290513f
C1034 VOUT+.n14 GNDA 0.195399f
C1035 VOUT+.t59 GNDA 0.290513f
C1036 VOUT+.n15 GNDA 0.24987f
C1037 VOUT+.t97 GNDA 0.290513f
C1038 VOUT+.n16 GNDA 0.24987f
C1039 VOUT+.t131 GNDA 0.290513f
C1040 VOUT+.n17 GNDA 0.24987f
C1041 VOUT+.t24 GNDA 0.290513f
C1042 VOUT+.n18 GNDA 0.24987f
C1043 VOUT+.t75 GNDA 0.290513f
C1044 VOUT+.n19 GNDA 0.24987f
C1045 VOUT+.t112 GNDA 0.290513f
C1046 VOUT+.n20 GNDA 0.24987f
C1047 VOUT+.t144 GNDA 0.290513f
C1048 VOUT+.n21 GNDA 0.24987f
C1049 VOUT+.t55 GNDA 0.290513f
C1050 VOUT+.n22 GNDA 0.24987f
C1051 VOUT+.t95 GNDA 0.290513f
C1052 VOUT+.n23 GNDA 0.24987f
C1053 VOUT+.n24 GNDA 0.236042f
C1054 VOUT+.t38 GNDA 0.295461f
C1055 VOUT+.t142 GNDA 0.290513f
C1056 VOUT+.n25 GNDA 0.194779f
C1057 VOUT+.t94 GNDA 0.290513f
C1058 VOUT+.t20 GNDA 0.295461f
C1059 VOUT+.t58 GNDA 0.290513f
C1060 VOUT+.n26 GNDA 0.194779f
C1061 VOUT+.n27 GNDA 0.236042f
C1062 VOUT+.t80 GNDA 0.295461f
C1063 VOUT+.t42 GNDA 0.290513f
C1064 VOUT+.n28 GNDA 0.194779f
C1065 VOUT+.t133 GNDA 0.290513f
C1066 VOUT+.t61 GNDA 0.295461f
C1067 VOUT+.t100 GNDA 0.290513f
C1068 VOUT+.n29 GNDA 0.194779f
C1069 VOUT+.n30 GNDA 0.236042f
C1070 VOUT+.t121 GNDA 0.295461f
C1071 VOUT+.t84 GNDA 0.290513f
C1072 VOUT+.n31 GNDA 0.194779f
C1073 VOUT+.t32 GNDA 0.290513f
C1074 VOUT+.t104 GNDA 0.295461f
C1075 VOUT+.t137 GNDA 0.290513f
C1076 VOUT+.n32 GNDA 0.194779f
C1077 VOUT+.n33 GNDA 0.236042f
C1078 VOUT+.t85 GNDA 0.295461f
C1079 VOUT+.t50 GNDA 0.290513f
C1080 VOUT+.n34 GNDA 0.194779f
C1081 VOUT+.t138 GNDA 0.290513f
C1082 VOUT+.t67 GNDA 0.295461f
C1083 VOUT+.t103 GNDA 0.290513f
C1084 VOUT+.n35 GNDA 0.194779f
C1085 VOUT+.n36 GNDA 0.236042f
C1086 VOUT+.t123 GNDA 0.295461f
C1087 VOUT+.t90 GNDA 0.290513f
C1088 VOUT+.n37 GNDA 0.194779f
C1089 VOUT+.t36 GNDA 0.290513f
C1090 VOUT+.t107 GNDA 0.295337f
C1091 VOUT+.t141 GNDA 0.290513f
C1092 VOUT+.n38 GNDA 0.193087f
C1093 VOUT+.n39 GNDA 0.236042f
C1094 VOUT+.t108 GNDA 0.295461f
C1095 VOUT+.t70 GNDA 0.290513f
C1096 VOUT+.n40 GNDA 0.194779f
C1097 VOUT+.t91 GNDA 0.290513f
C1098 VOUT+.n41 GNDA 0.127099f
C1099 VOUT+.t68 GNDA 0.295461f
C1100 VOUT+.t31 GNDA 0.290513f
C1101 VOUT+.n42 GNDA 0.194779f
C1102 VOUT+.t52 GNDA 0.290513f
C1103 VOUT+.t54 GNDA 0.294841f
C1104 VOUT+.t156 GNDA 0.294841f
C1105 VOUT+.t145 GNDA 0.295461f
C1106 VOUT+.t45 GNDA 0.290513f
C1107 VOUT+.n43 GNDA 0.194779f
C1108 VOUT+.t136 GNDA 0.290513f
C1109 VOUT+.n44 GNDA 0.127099f
C1110 VOUT+.t101 GNDA 0.290513f
C1111 VOUT+.n45 GNDA 0.12256f
C1112 VOUT+.t37 GNDA 0.294841f
C1113 VOUT+.t113 GNDA 0.295461f
C1114 VOUT+.t151 GNDA 0.290513f
C1115 VOUT+.n46 GNDA 0.194779f
C1116 VOUT+.t98 GNDA 0.290513f
C1117 VOUT+.n47 GNDA 0.127099f
C1118 VOUT+.t60 GNDA 0.290513f
C1119 VOUT+.n48 GNDA 0.12256f
C1120 VOUT+.t140 GNDA 0.294841f
C1121 VOUT+.t76 GNDA 0.295461f
C1122 VOUT+.t118 GNDA 0.290513f
C1123 VOUT+.n49 GNDA 0.194779f
C1124 VOUT+.t57 GNDA 0.290513f
C1125 VOUT+.n50 GNDA 0.127099f
C1126 VOUT+.t21 GNDA 0.290513f
C1127 VOUT+.n51 GNDA 0.12256f
C1128 VOUT+.t105 GNDA 0.294841f
C1129 VOUT+.t25 GNDA 0.295461f
C1130 VOUT+.t66 GNDA 0.290513f
C1131 VOUT+.n52 GNDA 0.194779f
C1132 VOUT+.t81 GNDA 0.290513f
C1133 VOUT+.n53 GNDA 0.127099f
C1134 VOUT+.t44 GNDA 0.290513f
C1135 VOUT+.n54 GNDA 0.12256f
C1136 VOUT+.t125 GNDA 0.294841f
C1137 VOUT+.t88 GNDA 0.294841f
C1138 VOUT+.t51 GNDA 0.294841f
C1139 VOUT+.t150 GNDA 0.294841f
C1140 VOUT+.t33 GNDA 0.294841f
C1141 VOUT+.t134 GNDA 0.290513f
C1142 VOUT+.n55 GNDA 0.195399f
C1143 VOUT+.t110 GNDA 0.290513f
C1144 VOUT+.n56 GNDA 0.24987f
C1145 VOUT+.t147 GNDA 0.290513f
C1146 VOUT+.n57 GNDA 0.24987f
C1147 VOUT+.t46 GNDA 0.290513f
C1148 VOUT+.n58 GNDA 0.24987f
C1149 VOUT+.t86 GNDA 0.290513f
C1150 VOUT+.n59 GNDA 0.30888f
C1151 VOUT+.t62 GNDA 0.290513f
C1152 VOUT+.n60 GNDA 0.30888f
C1153 VOUT+.t102 GNDA 0.290513f
C1154 VOUT+.n61 GNDA 0.30888f
C1155 VOUT+.t139 GNDA 0.290513f
C1156 VOUT+.n62 GNDA 0.30888f
C1157 VOUT+.t119 GNDA 0.290513f
C1158 VOUT+.n63 GNDA 0.24987f
C1159 VOUT+.t155 GNDA 0.290513f
C1160 VOUT+.n64 GNDA 0.24987f
C1161 VOUT+.n65 GNDA 0.236042f
C1162 VOUT+.t28 GNDA 0.295461f
C1163 VOUT+.t130 GNDA 0.290513f
C1164 VOUT+.n66 GNDA 0.194779f
C1165 VOUT+.t152 GNDA 0.290513f
C1166 VOUT+.t77 GNDA 0.295461f
C1167 VOUT+.t115 GNDA 0.290513f
C1168 VOUT+.n67 GNDA 0.194779f
C1169 VOUT+.n68 GNDA 0.236042f
C1170 VOUT+.t63 GNDA 0.295461f
C1171 VOUT+.t23 GNDA 0.290513f
C1172 VOUT+.n69 GNDA 0.194779f
C1173 VOUT+.t48 GNDA 0.290513f
C1174 VOUT+.t111 GNDA 0.295461f
C1175 VOUT+.t148 GNDA 0.290513f
C1176 VOUT+.n70 GNDA 0.194779f
C1177 VOUT+.n71 GNDA 0.236042f
C1178 VOUT+.t114 GNDA 0.295461f
C1179 VOUT+.t79 GNDA 0.290513f
C1180 VOUT+.n72 GNDA 0.194779f
C1181 VOUT+.t27 GNDA 0.290513f
C1182 VOUT+.t99 GNDA 0.295461f
C1183 VOUT+.t132 GNDA 0.290513f
C1184 VOUT+.n73 GNDA 0.194779f
C1185 VOUT+.n74 GNDA 0.236042f
C1186 VOUT+.t74 GNDA 0.295461f
C1187 VOUT+.t40 GNDA 0.290513f
C1188 VOUT+.n75 GNDA 0.194779f
C1189 VOUT+.t128 GNDA 0.290513f
C1190 VOUT+.t56 GNDA 0.295461f
C1191 VOUT+.t93 GNDA 0.290513f
C1192 VOUT+.n76 GNDA 0.194779f
C1193 VOUT+.n77 GNDA 0.236042f
C1194 VOUT+.t109 GNDA 0.295461f
C1195 VOUT+.t71 GNDA 0.290513f
C1196 VOUT+.n78 GNDA 0.194779f
C1197 VOUT+.t19 GNDA 0.290513f
C1198 VOUT+.t92 GNDA 0.295461f
C1199 VOUT+.t126 GNDA 0.290513f
C1200 VOUT+.n79 GNDA 0.194779f
C1201 VOUT+.n80 GNDA 0.236042f
C1202 VOUT+.t69 GNDA 0.295461f
C1203 VOUT+.t34 GNDA 0.290513f
C1204 VOUT+.n81 GNDA 0.194779f
C1205 VOUT+.t122 GNDA 0.290513f
C1206 VOUT+.t53 GNDA 0.295461f
C1207 VOUT+.t89 GNDA 0.290513f
C1208 VOUT+.n82 GNDA 0.194779f
C1209 VOUT+.n83 GNDA 0.236042f
C1210 VOUT+.t30 GNDA 0.295461f
C1211 VOUT+.t135 GNDA 0.290513f
C1212 VOUT+.n84 GNDA 0.194779f
C1213 VOUT+.t83 GNDA 0.290513f
C1214 VOUT+.t153 GNDA 0.295461f
C1215 VOUT+.t49 GNDA 0.290513f
C1216 VOUT+.n85 GNDA 0.194779f
C1217 VOUT+.n86 GNDA 0.236042f
C1218 VOUT+.t64 GNDA 0.295461f
C1219 VOUT+.t29 GNDA 0.290513f
C1220 VOUT+.n87 GNDA 0.194779f
C1221 VOUT+.t120 GNDA 0.290513f
C1222 VOUT+.t47 GNDA 0.295461f
C1223 VOUT+.t82 GNDA 0.290513f
C1224 VOUT+.n88 GNDA 0.194779f
C1225 VOUT+.n89 GNDA 0.236042f
C1226 VOUT+.t22 GNDA 0.295461f
C1227 VOUT+.t129 GNDA 0.290513f
C1228 VOUT+.n90 GNDA 0.194779f
C1229 VOUT+.t78 GNDA 0.290513f
C1230 VOUT+.n91 GNDA 0.236042f
C1231 VOUT+.t41 GNDA 0.290513f
C1232 VOUT+.n92 GNDA 0.127099f
C1233 VOUT+.t146 GNDA 0.290513f
C1234 VOUT+.n93 GNDA 0.238016f
C1235 VOUT+.n94 GNDA 0.268648f
C1236 VOUT+.t0 GNDA 0.05084f
C1237 VOUT+.t7 GNDA 0.05084f
C1238 VOUT+.n95 GNDA 0.235187f
C1239 VOUT+.t3 GNDA 0.05084f
C1240 VOUT+.t2 GNDA 0.05084f
C1241 VOUT+.n96 GNDA 0.2344f
C1242 VOUT+.n97 GNDA 0.144847f
C1243 VOUT+.t8 GNDA 0.05084f
C1244 VOUT+.t4 GNDA 0.05084f
C1245 VOUT+.n98 GNDA 0.2344f
C1246 VOUT+.n99 GNDA 0.089159f
C1247 VOUT+.t1 GNDA 0.084056f
C1248 VOUT+.n100 GNDA 0.119121f
C1249 bgr_0.V_mir1.t8 GNDA 0.053881f
C1250 bgr_0.V_mir1.t6 GNDA 0.042444f
C1251 bgr_0.V_mir1.t17 GNDA 0.042444f
C1252 bgr_0.V_mir1.t20 GNDA 0.06851f
C1253 bgr_0.V_mir1.n0 GNDA 0.076506f
C1254 bgr_0.V_mir1.n1 GNDA 0.052264f
C1255 bgr_0.V_mir1.n2 GNDA 0.081315f
C1256 bgr_0.V_mir1.t9 GNDA 0.03537f
C1257 bgr_0.V_mir1.t7 GNDA 0.03537f
C1258 bgr_0.V_mir1.n3 GNDA 0.08097f
C1259 bgr_0.V_mir1.n4 GNDA 0.203577f
C1260 bgr_0.V_mir1.t13 GNDA 0.017685f
C1261 bgr_0.V_mir1.t14 GNDA 0.017685f
C1262 bgr_0.V_mir1.n5 GNDA 0.046242f
C1263 bgr_0.V_mir1.t15 GNDA 0.075466f
C1264 bgr_0.V_mir1.t16 GNDA 0.017685f
C1265 bgr_0.V_mir1.t12 GNDA 0.017685f
C1266 bgr_0.V_mir1.n6 GNDA 0.050199f
C1267 bgr_0.V_mir1.n7 GNDA 0.827814f
C1268 bgr_0.V_mir1.n8 GNDA 0.268286f
C1269 bgr_0.V_mir1.t0 GNDA 0.053881f
C1270 bgr_0.V_mir1.t4 GNDA 0.042444f
C1271 bgr_0.V_mir1.t18 GNDA 0.042444f
C1272 bgr_0.V_mir1.t21 GNDA 0.06851f
C1273 bgr_0.V_mir1.n9 GNDA 0.076506f
C1274 bgr_0.V_mir1.n10 GNDA 0.052264f
C1275 bgr_0.V_mir1.n11 GNDA 0.081315f
C1276 bgr_0.V_mir1.t1 GNDA 0.03537f
C1277 bgr_0.V_mir1.t5 GNDA 0.03537f
C1278 bgr_0.V_mir1.n12 GNDA 0.08097f
C1279 bgr_0.V_mir1.n13 GNDA 0.156007f
C1280 bgr_0.V_mir1.n14 GNDA 0.09373f
C1281 bgr_0.V_mir1.n15 GNDA 0.699157f
C1282 bgr_0.V_mir1.t10 GNDA 0.053881f
C1283 bgr_0.V_mir1.t2 GNDA 0.042444f
C1284 bgr_0.V_mir1.t19 GNDA 0.042444f
C1285 bgr_0.V_mir1.t22 GNDA 0.06851f
C1286 bgr_0.V_mir1.n16 GNDA 0.076506f
C1287 bgr_0.V_mir1.n17 GNDA 0.052264f
C1288 bgr_0.V_mir1.n18 GNDA 0.081315f
C1289 bgr_0.V_mir1.n19 GNDA 0.201563f
C1290 bgr_0.V_mir1.t3 GNDA 0.03537f
C1291 bgr_0.V_mir1.n20 GNDA 0.08097f
C1292 bgr_0.V_mir1.t11 GNDA 0.03537f
C1293 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 GNDA 0.472073f
C1294 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 GNDA 0.113823f
C1295 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 GNDA 0.113823f
C1296 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 GNDA 0.470705f
C1297 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 GNDA 0.113823f
C1298 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 GNDA 0.113823f
C1299 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 GNDA 0.468899f
C1300 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 GNDA 0.65013f
C1301 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 GNDA 0.113823f
C1302 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 GNDA 0.113823f
C1303 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 GNDA 0.468899f
C1304 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 GNDA 0.339247f
C1305 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 GNDA 0.113823f
C1306 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 GNDA 0.113823f
C1307 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 GNDA 0.468899f
C1308 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 GNDA 0.339247f
C1309 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 GNDA 0.113823f
C1310 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 GNDA 0.113823f
C1311 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 GNDA 0.468899f
C1312 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 GNDA 0.490393f
C1313 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 GNDA 7.05f
C1314 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 GNDA 0.037941f
C1315 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 GNDA 0.037941f
C1316 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 GNDA 0.137905f
C1317 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 GNDA 0.037941f
C1318 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 GNDA 0.037941f
C1319 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 GNDA 0.114599f
C1320 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 GNDA 0.716408f
C1321 bgr_0.V_CMFB_S4 GNDA 5.75369f
C1322 two_stage_opamp_dummy_magic_0.Y.t14 GNDA 0.053187f
C1323 two_stage_opamp_dummy_magic_0.Y.t24 GNDA 0.053187f
C1324 two_stage_opamp_dummy_magic_0.Y.n0 GNDA 0.184972f
C1325 two_stage_opamp_dummy_magic_0.Y.t12 GNDA 0.053187f
C1326 two_stage_opamp_dummy_magic_0.Y.t7 GNDA 0.053187f
C1327 two_stage_opamp_dummy_magic_0.Y.n1 GNDA 0.184316f
C1328 two_stage_opamp_dummy_magic_0.Y.n2 GNDA 0.347971f
C1329 two_stage_opamp_dummy_magic_0.Y.t13 GNDA 0.053187f
C1330 two_stage_opamp_dummy_magic_0.Y.t18 GNDA 0.053187f
C1331 two_stage_opamp_dummy_magic_0.Y.n3 GNDA 0.184316f
C1332 two_stage_opamp_dummy_magic_0.Y.n4 GNDA 0.180392f
C1333 two_stage_opamp_dummy_magic_0.Y.t8 GNDA 0.053187f
C1334 two_stage_opamp_dummy_magic_0.Y.t9 GNDA 0.053187f
C1335 two_stage_opamp_dummy_magic_0.Y.n5 GNDA 0.184316f
C1336 two_stage_opamp_dummy_magic_0.Y.n6 GNDA 0.180392f
C1337 two_stage_opamp_dummy_magic_0.Y.t23 GNDA 0.053187f
C1338 two_stage_opamp_dummy_magic_0.Y.t10 GNDA 0.053187f
C1339 two_stage_opamp_dummy_magic_0.Y.n7 GNDA 0.184316f
C1340 two_stage_opamp_dummy_magic_0.Y.n8 GNDA 0.212415f
C1341 two_stage_opamp_dummy_magic_0.Y.t5 GNDA 0.053187f
C1342 two_stage_opamp_dummy_magic_0.Y.t3 GNDA 0.053187f
C1343 two_stage_opamp_dummy_magic_0.Y.n9 GNDA 0.180498f
C1344 two_stage_opamp_dummy_magic_0.Y.n10 GNDA 0.149147f
C1345 two_stage_opamp_dummy_magic_0.Y.t4 GNDA 0.022794f
C1346 two_stage_opamp_dummy_magic_0.Y.t6 GNDA 0.022794f
C1347 two_stage_opamp_dummy_magic_0.Y.n11 GNDA 0.076959f
C1348 two_stage_opamp_dummy_magic_0.Y.t21 GNDA 0.022794f
C1349 two_stage_opamp_dummy_magic_0.Y.t19 GNDA 0.022794f
C1350 two_stage_opamp_dummy_magic_0.Y.n12 GNDA 0.082252f
C1351 two_stage_opamp_dummy_magic_0.Y.t0 GNDA 0.022794f
C1352 two_stage_opamp_dummy_magic_0.Y.t1 GNDA 0.022794f
C1353 two_stage_opamp_dummy_magic_0.Y.n13 GNDA 0.081534f
C1354 two_stage_opamp_dummy_magic_0.Y.n14 GNDA 0.302737f
C1355 two_stage_opamp_dummy_magic_0.Y.t20 GNDA 0.022794f
C1356 two_stage_opamp_dummy_magic_0.Y.t15 GNDA 0.022794f
C1357 two_stage_opamp_dummy_magic_0.Y.n15 GNDA 0.081534f
C1358 two_stage_opamp_dummy_magic_0.Y.n16 GNDA 0.157046f
C1359 two_stage_opamp_dummy_magic_0.Y.t17 GNDA 0.022794f
C1360 two_stage_opamp_dummy_magic_0.Y.t2 GNDA 0.022794f
C1361 two_stage_opamp_dummy_magic_0.Y.n17 GNDA 0.081534f
C1362 two_stage_opamp_dummy_magic_0.Y.n18 GNDA 0.157046f
C1363 two_stage_opamp_dummy_magic_0.Y.t16 GNDA 0.022794f
C1364 two_stage_opamp_dummy_magic_0.Y.t22 GNDA 0.022794f
C1365 two_stage_opamp_dummy_magic_0.Y.n19 GNDA 0.082252f
C1366 two_stage_opamp_dummy_magic_0.Y.n20 GNDA 0.191279f
C1367 two_stage_opamp_dummy_magic_0.Y.n21 GNDA 0.123631f
C1368 two_stage_opamp_dummy_magic_0.Y.t46 GNDA 0.031912f
C1369 two_stage_opamp_dummy_magic_0.Y.t35 GNDA 0.031912f
C1370 two_stage_opamp_dummy_magic_0.Y.t47 GNDA 0.031912f
C1371 two_stage_opamp_dummy_magic_0.Y.t31 GNDA 0.031912f
C1372 two_stage_opamp_dummy_magic_0.Y.t43 GNDA 0.031912f
C1373 two_stage_opamp_dummy_magic_0.Y.t28 GNDA 0.031912f
C1374 two_stage_opamp_dummy_magic_0.Y.t41 GNDA 0.031912f
C1375 two_stage_opamp_dummy_magic_0.Y.t26 GNDA 0.03875f
C1376 two_stage_opamp_dummy_magic_0.Y.n22 GNDA 0.03875f
C1377 two_stage_opamp_dummy_magic_0.Y.n23 GNDA 0.025074f
C1378 two_stage_opamp_dummy_magic_0.Y.n24 GNDA 0.025074f
C1379 two_stage_opamp_dummy_magic_0.Y.n25 GNDA 0.025074f
C1380 two_stage_opamp_dummy_magic_0.Y.n26 GNDA 0.025074f
C1381 two_stage_opamp_dummy_magic_0.Y.n27 GNDA 0.025074f
C1382 two_stage_opamp_dummy_magic_0.Y.n28 GNDA 0.022459f
C1383 two_stage_opamp_dummy_magic_0.Y.t34 GNDA 0.031912f
C1384 two_stage_opamp_dummy_magic_0.Y.t51 GNDA 0.03875f
C1385 two_stage_opamp_dummy_magic_0.Y.n29 GNDA 0.036135f
C1386 two_stage_opamp_dummy_magic_0.Y.n30 GNDA 0.022101f
C1387 two_stage_opamp_dummy_magic_0.Y.t53 GNDA 0.049008f
C1388 two_stage_opamp_dummy_magic_0.Y.t40 GNDA 0.049008f
C1389 two_stage_opamp_dummy_magic_0.Y.t54 GNDA 0.049008f
C1390 two_stage_opamp_dummy_magic_0.Y.t38 GNDA 0.049008f
C1391 two_stage_opamp_dummy_magic_0.Y.t50 GNDA 0.049008f
C1392 two_stage_opamp_dummy_magic_0.Y.t33 GNDA 0.049008f
C1393 two_stage_opamp_dummy_magic_0.Y.t45 GNDA 0.049008f
C1394 two_stage_opamp_dummy_magic_0.Y.t30 GNDA 0.055713f
C1395 two_stage_opamp_dummy_magic_0.Y.n31 GNDA 0.05028f
C1396 two_stage_opamp_dummy_magic_0.Y.n32 GNDA 0.030772f
C1397 two_stage_opamp_dummy_magic_0.Y.n33 GNDA 0.030772f
C1398 two_stage_opamp_dummy_magic_0.Y.n34 GNDA 0.030772f
C1399 two_stage_opamp_dummy_magic_0.Y.n35 GNDA 0.030772f
C1400 two_stage_opamp_dummy_magic_0.Y.n36 GNDA 0.030772f
C1401 two_stage_opamp_dummy_magic_0.Y.n37 GNDA 0.028157f
C1402 two_stage_opamp_dummy_magic_0.Y.t39 GNDA 0.049008f
C1403 two_stage_opamp_dummy_magic_0.Y.t25 GNDA 0.055713f
C1404 two_stage_opamp_dummy_magic_0.Y.n38 GNDA 0.047665f
C1405 two_stage_opamp_dummy_magic_0.Y.n39 GNDA 0.022031f
C1406 two_stage_opamp_dummy_magic_0.Y.n40 GNDA 0.153015f
C1407 two_stage_opamp_dummy_magic_0.Y.t11 GNDA 0.741299f
C1408 two_stage_opamp_dummy_magic_0.Y.t29 GNDA 0.100295f
C1409 two_stage_opamp_dummy_magic_0.Y.t42 GNDA 0.100295f
C1410 two_stage_opamp_dummy_magic_0.Y.t27 GNDA 0.106821f
C1411 two_stage_opamp_dummy_magic_0.Y.n41 GNDA 0.084651f
C1412 two_stage_opamp_dummy_magic_0.Y.n42 GNDA 0.045253f
C1413 two_stage_opamp_dummy_magic_0.Y.t44 GNDA 0.100295f
C1414 two_stage_opamp_dummy_magic_0.Y.t32 GNDA 0.100295f
C1415 two_stage_opamp_dummy_magic_0.Y.t49 GNDA 0.100295f
C1416 two_stage_opamp_dummy_magic_0.Y.t37 GNDA 0.100295f
C1417 two_stage_opamp_dummy_magic_0.Y.t48 GNDA 0.100295f
C1418 two_stage_opamp_dummy_magic_0.Y.t36 GNDA 0.100295f
C1419 two_stage_opamp_dummy_magic_0.Y.t52 GNDA 0.106821f
C1420 two_stage_opamp_dummy_magic_0.Y.n43 GNDA 0.084651f
C1421 two_stage_opamp_dummy_magic_0.Y.n44 GNDA 0.047868f
C1422 two_stage_opamp_dummy_magic_0.Y.n45 GNDA 0.047868f
C1423 two_stage_opamp_dummy_magic_0.Y.n46 GNDA 0.047868f
C1424 two_stage_opamp_dummy_magic_0.Y.n47 GNDA 0.047868f
C1425 two_stage_opamp_dummy_magic_0.Y.n48 GNDA 0.045253f
C1426 two_stage_opamp_dummy_magic_0.Y.n49 GNDA 0.024415f
C1427 two_stage_opamp_dummy_magic_0.Y.n50 GNDA 1.03694f
C1428 two_stage_opamp_dummy_magic_0.Y.n51 GNDA 0.458663f
C1429 bgr_0.PFET_GATE_10uA.t23 GNDA 0.039179f
C1430 bgr_0.PFET_GATE_10uA.t16 GNDA 0.057916f
C1431 bgr_0.PFET_GATE_10uA.n0 GNDA 0.063817f
C1432 bgr_0.PFET_GATE_10uA.t29 GNDA 0.039179f
C1433 bgr_0.PFET_GATE_10uA.t17 GNDA 0.057916f
C1434 bgr_0.PFET_GATE_10uA.n1 GNDA 0.063817f
C1435 bgr_0.PFET_GATE_10uA.n2 GNDA 0.076791f
C1436 bgr_0.PFET_GATE_10uA.t10 GNDA 0.039179f
C1437 bgr_0.PFET_GATE_10uA.t24 GNDA 0.057916f
C1438 bgr_0.PFET_GATE_10uA.n3 GNDA 0.063817f
C1439 bgr_0.PFET_GATE_10uA.t18 GNDA 0.039179f
C1440 bgr_0.PFET_GATE_10uA.t25 GNDA 0.057916f
C1441 bgr_0.PFET_GATE_10uA.n4 GNDA 0.063817f
C1442 bgr_0.PFET_GATE_10uA.n5 GNDA 0.064022f
C1443 bgr_0.PFET_GATE_10uA.t3 GNDA 0.781422f
C1444 bgr_0.PFET_GATE_10uA.t8 GNDA 0.586977f
C1445 bgr_0.PFET_GATE_10uA.t1 GNDA 0.040183f
C1446 bgr_0.PFET_GATE_10uA.t7 GNDA 0.040183f
C1447 bgr_0.PFET_GATE_10uA.n6 GNDA 0.102705f
C1448 bgr_0.PFET_GATE_10uA.t0 GNDA 0.040183f
C1449 bgr_0.PFET_GATE_10uA.t4 GNDA 0.040183f
C1450 bgr_0.PFET_GATE_10uA.n7 GNDA 0.100051f
C1451 bgr_0.PFET_GATE_10uA.n8 GNDA 0.978629f
C1452 bgr_0.PFET_GATE_10uA.t2 GNDA 0.040183f
C1453 bgr_0.PFET_GATE_10uA.t9 GNDA 0.040183f
C1454 bgr_0.PFET_GATE_10uA.n9 GNDA 0.100051f
C1455 bgr_0.PFET_GATE_10uA.n10 GNDA 0.554934f
C1456 bgr_0.PFET_GATE_10uA.n11 GNDA 1.13286f
C1457 bgr_0.PFET_GATE_10uA.t6 GNDA 0.040183f
C1458 bgr_0.PFET_GATE_10uA.t5 GNDA 0.040183f
C1459 bgr_0.PFET_GATE_10uA.n12 GNDA 0.096913f
C1460 bgr_0.PFET_GATE_10uA.n13 GNDA 0.356682f
C1461 bgr_0.PFET_GATE_10uA.n14 GNDA 3.84996f
C1462 bgr_0.PFET_GATE_10uA.t13 GNDA 0.045299f
C1463 bgr_0.PFET_GATE_10uA.t21 GNDA 0.045299f
C1464 bgr_0.PFET_GATE_10uA.n15 GNDA 0.137138f
C1465 bgr_0.PFET_GATE_10uA.n16 GNDA 1.78858f
C1466 bgr_0.PFET_GATE_10uA.n17 GNDA 1.41725f
C1467 bgr_0.PFET_GATE_10uA.t27 GNDA 0.039179f
C1468 bgr_0.PFET_GATE_10uA.t20 GNDA 0.039179f
C1469 bgr_0.PFET_GATE_10uA.t12 GNDA 0.039179f
C1470 bgr_0.PFET_GATE_10uA.t26 GNDA 0.039179f
C1471 bgr_0.PFET_GATE_10uA.t19 GNDA 0.039179f
C1472 bgr_0.PFET_GATE_10uA.t11 GNDA 0.057916f
C1473 bgr_0.PFET_GATE_10uA.n18 GNDA 0.071675f
C1474 bgr_0.PFET_GATE_10uA.n19 GNDA 0.051234f
C1475 bgr_0.PFET_GATE_10uA.n20 GNDA 0.051234f
C1476 bgr_0.PFET_GATE_10uA.n21 GNDA 0.051234f
C1477 bgr_0.PFET_GATE_10uA.n22 GNDA 0.043376f
C1478 bgr_0.PFET_GATE_10uA.t14 GNDA 0.039179f
C1479 bgr_0.PFET_GATE_10uA.t22 GNDA 0.039179f
C1480 bgr_0.PFET_GATE_10uA.t28 GNDA 0.039179f
C1481 bgr_0.PFET_GATE_10uA.t15 GNDA 0.057916f
C1482 bgr_0.PFET_GATE_10uA.n23 GNDA 0.071675f
C1483 bgr_0.PFET_GATE_10uA.n24 GNDA 0.051234f
C1484 bgr_0.PFET_GATE_10uA.n25 GNDA 0.043376f
C1485 bgr_0.PFET_GATE_10uA.n26 GNDA 0.05954f
C1486 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 GNDA 0.025048f
C1487 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 GNDA 0.025048f
C1488 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 GNDA 0.062786f
C1489 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 GNDA 0.025048f
C1490 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 GNDA 0.025048f
C1491 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 GNDA 0.062455f
C1492 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 GNDA 0.555098f
C1493 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 GNDA 0.025048f
C1494 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 GNDA 0.025048f
C1495 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 GNDA 0.050096f
C1496 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 GNDA 0.279975f
C1497 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 GNDA 0.320788f
C1498 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 GNDA 0.050096f
C1499 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 GNDA 0.050096f
C1500 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 GNDA 0.146978f
C1501 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 GNDA 0.050096f
C1502 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 GNDA 0.050096f
C1503 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 GNDA 0.146311f
C1504 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 GNDA 0.505735f
C1505 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 GNDA 0.050096f
C1506 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 GNDA 0.050096f
C1507 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 GNDA 0.146311f
C1508 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 GNDA 0.261968f
C1509 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 GNDA 0.050096f
C1510 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 GNDA 0.050096f
C1511 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 GNDA 0.146311f
C1512 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 GNDA 0.261968f
C1513 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 GNDA 0.050096f
C1514 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 GNDA 0.050096f
C1515 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 GNDA 0.146311f
C1516 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 GNDA 0.376359f
C1517 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 GNDA 2.53757f
C1518 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 GNDA 2.79499f
C1519 bgr_0.V_CMFB_S1 GNDA 0.046745f
C1520 two_stage_opamp_dummy_magic_0.X.t14 GNDA 0.052601f
C1521 two_stage_opamp_dummy_magic_0.X.t7 GNDA 0.052601f
C1522 two_stage_opamp_dummy_magic_0.X.n0 GNDA 0.182935f
C1523 two_stage_opamp_dummy_magic_0.X.t2 GNDA 0.052601f
C1524 two_stage_opamp_dummy_magic_0.X.t20 GNDA 0.052601f
C1525 two_stage_opamp_dummy_magic_0.X.n1 GNDA 0.182287f
C1526 two_stage_opamp_dummy_magic_0.X.n2 GNDA 0.344139f
C1527 two_stage_opamp_dummy_magic_0.X.t18 GNDA 0.052601f
C1528 two_stage_opamp_dummy_magic_0.X.t1 GNDA 0.052601f
C1529 two_stage_opamp_dummy_magic_0.X.n3 GNDA 0.182287f
C1530 two_stage_opamp_dummy_magic_0.X.n4 GNDA 0.178405f
C1531 two_stage_opamp_dummy_magic_0.X.t16 GNDA 0.052601f
C1532 two_stage_opamp_dummy_magic_0.X.t12 GNDA 0.052601f
C1533 two_stage_opamp_dummy_magic_0.X.n5 GNDA 0.182287f
C1534 two_stage_opamp_dummy_magic_0.X.n6 GNDA 0.178405f
C1535 two_stage_opamp_dummy_magic_0.X.t6 GNDA 0.052601f
C1536 two_stage_opamp_dummy_magic_0.X.t0 GNDA 0.052601f
C1537 two_stage_opamp_dummy_magic_0.X.n7 GNDA 0.182287f
C1538 two_stage_opamp_dummy_magic_0.X.n8 GNDA 0.210076f
C1539 two_stage_opamp_dummy_magic_0.X.t13 GNDA 0.052601f
C1540 two_stage_opamp_dummy_magic_0.X.t17 GNDA 0.052601f
C1541 two_stage_opamp_dummy_magic_0.X.n9 GNDA 0.178511f
C1542 two_stage_opamp_dummy_magic_0.X.n10 GNDA 0.147505f
C1543 two_stage_opamp_dummy_magic_0.X.t19 GNDA 0.022543f
C1544 two_stage_opamp_dummy_magic_0.X.t10 GNDA 0.022543f
C1545 two_stage_opamp_dummy_magic_0.X.n11 GNDA 0.076111f
C1546 two_stage_opamp_dummy_magic_0.X.t21 GNDA 0.022543f
C1547 two_stage_opamp_dummy_magic_0.X.t5 GNDA 0.022543f
C1548 two_stage_opamp_dummy_magic_0.X.n12 GNDA 0.081346f
C1549 two_stage_opamp_dummy_magic_0.X.t8 GNDA 0.022543f
C1550 two_stage_opamp_dummy_magic_0.X.t22 GNDA 0.022543f
C1551 two_stage_opamp_dummy_magic_0.X.n13 GNDA 0.081346f
C1552 two_stage_opamp_dummy_magic_0.X.t15 GNDA 0.022543f
C1553 two_stage_opamp_dummy_magic_0.X.t3 GNDA 0.022543f
C1554 two_stage_opamp_dummy_magic_0.X.n14 GNDA 0.080636f
C1555 two_stage_opamp_dummy_magic_0.X.n15 GNDA 0.299403f
C1556 two_stage_opamp_dummy_magic_0.X.t4 GNDA 0.022543f
C1557 two_stage_opamp_dummy_magic_0.X.t23 GNDA 0.022543f
C1558 two_stage_opamp_dummy_magic_0.X.n16 GNDA 0.080636f
C1559 two_stage_opamp_dummy_magic_0.X.n17 GNDA 0.155317f
C1560 two_stage_opamp_dummy_magic_0.X.t9 GNDA 0.022543f
C1561 two_stage_opamp_dummy_magic_0.X.t24 GNDA 0.022543f
C1562 two_stage_opamp_dummy_magic_0.X.n18 GNDA 0.080636f
C1563 two_stage_opamp_dummy_magic_0.X.n19 GNDA 0.155317f
C1564 two_stage_opamp_dummy_magic_0.X.n20 GNDA 0.189173f
C1565 two_stage_opamp_dummy_magic_0.X.n21 GNDA 0.122269f
C1566 two_stage_opamp_dummy_magic_0.X.n22 GNDA 0.128676f
C1567 two_stage_opamp_dummy_magic_0.X.t47 GNDA 0.03156f
C1568 two_stage_opamp_dummy_magic_0.X.t33 GNDA 0.038324f
C1569 two_stage_opamp_dummy_magic_0.X.n23 GNDA 0.035737f
C1570 two_stage_opamp_dummy_magic_0.X.t37 GNDA 0.03156f
C1571 two_stage_opamp_dummy_magic_0.X.t50 GNDA 0.03156f
C1572 two_stage_opamp_dummy_magic_0.X.t25 GNDA 0.03156f
C1573 two_stage_opamp_dummy_magic_0.X.t42 GNDA 0.03156f
C1574 two_stage_opamp_dummy_magic_0.X.t28 GNDA 0.03156f
C1575 two_stage_opamp_dummy_magic_0.X.t44 GNDA 0.03156f
C1576 two_stage_opamp_dummy_magic_0.X.t32 GNDA 0.03156f
C1577 two_stage_opamp_dummy_magic_0.X.t54 GNDA 0.038324f
C1578 two_stage_opamp_dummy_magic_0.X.n24 GNDA 0.038324f
C1579 two_stage_opamp_dummy_magic_0.X.n25 GNDA 0.024798f
C1580 two_stage_opamp_dummy_magic_0.X.n26 GNDA 0.024798f
C1581 two_stage_opamp_dummy_magic_0.X.n27 GNDA 0.024798f
C1582 two_stage_opamp_dummy_magic_0.X.n28 GNDA 0.024798f
C1583 two_stage_opamp_dummy_magic_0.X.n29 GNDA 0.024798f
C1584 two_stage_opamp_dummy_magic_0.X.n30 GNDA 0.022211f
C1585 two_stage_opamp_dummy_magic_0.X.n31 GNDA 0.021857f
C1586 two_stage_opamp_dummy_magic_0.X.t52 GNDA 0.048468f
C1587 two_stage_opamp_dummy_magic_0.X.t40 GNDA 0.0551f
C1588 two_stage_opamp_dummy_magic_0.X.n32 GNDA 0.04714f
C1589 two_stage_opamp_dummy_magic_0.X.t41 GNDA 0.048468f
C1590 two_stage_opamp_dummy_magic_0.X.t53 GNDA 0.048468f
C1591 two_stage_opamp_dummy_magic_0.X.t31 GNDA 0.048468f
C1592 two_stage_opamp_dummy_magic_0.X.t46 GNDA 0.048468f
C1593 two_stage_opamp_dummy_magic_0.X.t36 GNDA 0.048468f
C1594 two_stage_opamp_dummy_magic_0.X.t49 GNDA 0.048468f
C1595 two_stage_opamp_dummy_magic_0.X.t39 GNDA 0.048468f
C1596 two_stage_opamp_dummy_magic_0.X.t29 GNDA 0.0551f
C1597 two_stage_opamp_dummy_magic_0.X.n33 GNDA 0.049726f
C1598 two_stage_opamp_dummy_magic_0.X.n34 GNDA 0.030433f
C1599 two_stage_opamp_dummy_magic_0.X.n35 GNDA 0.030433f
C1600 two_stage_opamp_dummy_magic_0.X.n36 GNDA 0.030433f
C1601 two_stage_opamp_dummy_magic_0.X.n37 GNDA 0.030433f
C1602 two_stage_opamp_dummy_magic_0.X.n38 GNDA 0.030433f
C1603 two_stage_opamp_dummy_magic_0.X.n39 GNDA 0.027847f
C1604 two_stage_opamp_dummy_magic_0.X.n40 GNDA 0.021789f
C1605 two_stage_opamp_dummy_magic_0.X.n41 GNDA 0.153028f
C1606 two_stage_opamp_dummy_magic_0.X.n42 GNDA 0.454714f
C1607 two_stage_opamp_dummy_magic_0.X.t30 GNDA 0.09919f
C1608 two_stage_opamp_dummy_magic_0.X.t43 GNDA 0.09919f
C1609 two_stage_opamp_dummy_magic_0.X.t27 GNDA 0.09919f
C1610 two_stage_opamp_dummy_magic_0.X.t51 GNDA 0.09919f
C1611 two_stage_opamp_dummy_magic_0.X.t38 GNDA 0.09919f
C1612 two_stage_opamp_dummy_magic_0.X.t48 GNDA 0.09919f
C1613 two_stage_opamp_dummy_magic_0.X.t35 GNDA 0.105644f
C1614 two_stage_opamp_dummy_magic_0.X.n43 GNDA 0.083719f
C1615 two_stage_opamp_dummy_magic_0.X.n44 GNDA 0.047341f
C1616 two_stage_opamp_dummy_magic_0.X.n45 GNDA 0.047341f
C1617 two_stage_opamp_dummy_magic_0.X.n46 GNDA 0.047341f
C1618 two_stage_opamp_dummy_magic_0.X.n47 GNDA 0.047341f
C1619 two_stage_opamp_dummy_magic_0.X.n48 GNDA 0.044755f
C1620 two_stage_opamp_dummy_magic_0.X.t45 GNDA 0.09919f
C1621 two_stage_opamp_dummy_magic_0.X.t34 GNDA 0.09919f
C1622 two_stage_opamp_dummy_magic_0.X.t26 GNDA 0.105644f
C1623 two_stage_opamp_dummy_magic_0.X.n49 GNDA 0.083719f
C1624 two_stage_opamp_dummy_magic_0.X.n50 GNDA 0.044755f
C1625 two_stage_opamp_dummy_magic_0.X.n51 GNDA 0.024251f
C1626 two_stage_opamp_dummy_magic_0.X.n52 GNDA 1.03308f
C1627 two_stage_opamp_dummy_magic_0.X.t11 GNDA 0.734227f
C1628 two_stage_opamp_dummy_magic_0.V_err_gate.n0 GNDA 1.91359f
C1629 two_stage_opamp_dummy_magic_0.V_err_gate.n1 GNDA 8.98709f
C1630 two_stage_opamp_dummy_magic_0.V_err_gate.t10 GNDA 0.026899f
C1631 two_stage_opamp_dummy_magic_0.V_err_gate.t11 GNDA 0.026899f
C1632 two_stage_opamp_dummy_magic_0.V_err_gate.n2 GNDA 0.062787f
C1633 two_stage_opamp_dummy_magic_0.V_err_gate.t3 GNDA 0.026899f
C1634 two_stage_opamp_dummy_magic_0.V_err_gate.t0 GNDA 0.026899f
C1635 two_stage_opamp_dummy_magic_0.V_err_gate.n3 GNDA 0.062382f
C1636 two_stage_opamp_dummy_magic_0.V_err_gate.t7 GNDA 0.026899f
C1637 two_stage_opamp_dummy_magic_0.V_err_gate.t8 GNDA 0.026899f
C1638 two_stage_opamp_dummy_magic_0.V_err_gate.n4 GNDA 0.062382f
C1639 two_stage_opamp_dummy_magic_0.V_err_gate.t23 GNDA 0.022191f
C1640 two_stage_opamp_dummy_magic_0.V_err_gate.t32 GNDA 0.022191f
C1641 two_stage_opamp_dummy_magic_0.V_err_gate.t21 GNDA 0.022191f
C1642 two_stage_opamp_dummy_magic_0.V_err_gate.t30 GNDA 0.022191f
C1643 two_stage_opamp_dummy_magic_0.V_err_gate.t16 GNDA 0.022191f
C1644 two_stage_opamp_dummy_magic_0.V_err_gate.t25 GNDA 0.022191f
C1645 two_stage_opamp_dummy_magic_0.V_err_gate.t18 GNDA 0.022191f
C1646 two_stage_opamp_dummy_magic_0.V_err_gate.t28 GNDA 0.022191f
C1647 two_stage_opamp_dummy_magic_0.V_err_gate.t15 GNDA 0.022191f
C1648 two_stage_opamp_dummy_magic_0.V_err_gate.t24 GNDA 0.022191f
C1649 two_stage_opamp_dummy_magic_0.V_err_gate.t33 GNDA 0.022191f
C1650 two_stage_opamp_dummy_magic_0.V_err_gate.t22 GNDA 0.022191f
C1651 two_stage_opamp_dummy_magic_0.V_err_gate.t31 GNDA 0.022191f
C1652 two_stage_opamp_dummy_magic_0.V_err_gate.t19 GNDA 0.022191f
C1653 two_stage_opamp_dummy_magic_0.V_err_gate.t26 GNDA 0.022191f
C1654 two_stage_opamp_dummy_magic_0.V_err_gate.t20 GNDA 0.022191f
C1655 two_stage_opamp_dummy_magic_0.V_err_gate.t29 GNDA 0.048082f
C1656 two_stage_opamp_dummy_magic_0.V_err_gate.n5 GNDA 0.07498f
C1657 two_stage_opamp_dummy_magic_0.V_err_gate.n6 GNDA 0.058505f
C1658 two_stage_opamp_dummy_magic_0.V_err_gate.n7 GNDA 0.058505f
C1659 two_stage_opamp_dummy_magic_0.V_err_gate.n8 GNDA 0.058505f
C1660 two_stage_opamp_dummy_magic_0.V_err_gate.n9 GNDA 0.058505f
C1661 two_stage_opamp_dummy_magic_0.V_err_gate.n10 GNDA 0.058505f
C1662 two_stage_opamp_dummy_magic_0.V_err_gate.n11 GNDA 0.058505f
C1663 two_stage_opamp_dummy_magic_0.V_err_gate.n12 GNDA 0.058505f
C1664 two_stage_opamp_dummy_magic_0.V_err_gate.n13 GNDA 0.058505f
C1665 two_stage_opamp_dummy_magic_0.V_err_gate.n14 GNDA 0.058505f
C1666 two_stage_opamp_dummy_magic_0.V_err_gate.n15 GNDA 0.058505f
C1667 two_stage_opamp_dummy_magic_0.V_err_gate.n16 GNDA 0.058505f
C1668 two_stage_opamp_dummy_magic_0.V_err_gate.n17 GNDA 0.058505f
C1669 two_stage_opamp_dummy_magic_0.V_err_gate.n18 GNDA 0.058505f
C1670 two_stage_opamp_dummy_magic_0.V_err_gate.n19 GNDA 0.058505f
C1671 two_stage_opamp_dummy_magic_0.V_err_gate.n20 GNDA 0.050064f
C1672 two_stage_opamp_dummy_magic_0.V_err_gate.t14 GNDA 0.022191f
C1673 two_stage_opamp_dummy_magic_0.V_err_gate.t27 GNDA 0.022191f
C1674 two_stage_opamp_dummy_magic_0.V_err_gate.t17 GNDA 0.048082f
C1675 two_stage_opamp_dummy_magic_0.V_err_gate.n21 GNDA 0.07498f
C1676 two_stage_opamp_dummy_magic_0.V_err_gate.n22 GNDA 0.050064f
C1677 two_stage_opamp_dummy_magic_0.V_err_gate.n23 GNDA 0.080671f
C1678 two_stage_opamp_dummy_magic_0.V_err_gate.t2 GNDA 0.026899f
C1679 two_stage_opamp_dummy_magic_0.V_err_gate.t4 GNDA 0.026899f
C1680 two_stage_opamp_dummy_magic_0.V_err_gate.n24 GNDA 0.053798f
C1681 two_stage_opamp_dummy_magic_0.V_err_gate.n25 GNDA 0.160251f
C1682 two_stage_opamp_dummy_magic_0.V_err_gate.t9 GNDA 0.026899f
C1683 two_stage_opamp_dummy_magic_0.V_err_gate.t13 GNDA 0.026899f
C1684 two_stage_opamp_dummy_magic_0.V_err_gate.n26 GNDA 0.062382f
C1685 two_stage_opamp_dummy_magic_0.V_err_gate.t12 GNDA 0.026899f
C1686 two_stage_opamp_dummy_magic_0.V_err_gate.t1 GNDA 0.026899f
C1687 two_stage_opamp_dummy_magic_0.V_err_gate.n27 GNDA 0.061917f
C1688 two_stage_opamp_dummy_magic_0.V_err_gate.t6 GNDA 0.053798f
C1689 two_stage_opamp_dummy_magic_0.V_err_gate.t5 GNDA 0.053798f
C1690 two_stage_opamp_dummy_magic_0.V_err_gate.n28 GNDA 0.165934f
C1691 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 GNDA 0.067041f
C1692 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 GNDA 0.025069f
C1693 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 GNDA 0.078631f
C1694 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 GNDA 0.025069f
C1695 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 GNDA 0.064367f
C1696 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 GNDA 0.025069f
C1697 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 GNDA 0.064367f
C1698 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 GNDA 0.025069f
C1699 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 GNDA 0.09875f
C1700 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 GNDA 0.640196f
C1701 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 GNDA 0.081305f
C1702 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 GNDA 0.081305f
C1703 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 GNDA 0.272455f
C1704 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 GNDA 3.06995f
C1705 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 GNDA 0.081305f
C1706 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 GNDA 0.081305f
C1707 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 GNDA 0.272455f
C1708 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 GNDA 0.73573f
C1709 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 GNDA 0.081305f
C1710 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 GNDA 0.081305f
C1711 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 GNDA 0.272455f
C1712 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 GNDA 1.05185f
C1713 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 GNDA 0.914983f
C1714 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 GNDA 0.039179f
C1715 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 GNDA 0.012307f
C1716 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 GNDA 0.022965f
C1717 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 GNDA 0.054829f
C1718 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 GNDA 0.342833f
C1719 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 GNDA 0.012307f
C1720 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 GNDA 0.022965f
C1721 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 GNDA 0.054829f
C1722 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 GNDA 0.316697f
C1723 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 GNDA 0.038804f
C1724 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 GNDA 0.30837f
C1725 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 GNDA 0.012307f
C1726 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 GNDA 0.022965f
C1727 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 GNDA 0.054829f
C1728 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 GNDA 0.191487f
C1729 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 GNDA 0.012307f
C1730 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 GNDA 0.022965f
C1731 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 GNDA 0.054829f
C1732 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 GNDA 0.297626f
C1733 bgr_0.V_mir2.t2 GNDA 0.017685f
C1734 bgr_0.V_mir2.t1 GNDA 0.017685f
C1735 bgr_0.V_mir2.n0 GNDA 0.046242f
C1736 bgr_0.V_mir2.t0 GNDA 0.075466f
C1737 bgr_0.V_mir2.t3 GNDA 0.017685f
C1738 bgr_0.V_mir2.t4 GNDA 0.017685f
C1739 bgr_0.V_mir2.n1 GNDA 0.050199f
C1740 bgr_0.V_mir2.n2 GNDA 0.827814f
C1741 bgr_0.V_mir2.n3 GNDA 0.268286f
C1742 bgr_0.V_mir2.t5 GNDA 0.042444f
C1743 bgr_0.V_mir2.t18 GNDA 0.042444f
C1744 bgr_0.V_mir2.t20 GNDA 0.06851f
C1745 bgr_0.V_mir2.n4 GNDA 0.076506f
C1746 bgr_0.V_mir2.n5 GNDA 0.052264f
C1747 bgr_0.V_mir2.t9 GNDA 0.053881f
C1748 bgr_0.V_mir2.n6 GNDA 0.081315f
C1749 bgr_0.V_mir2.t6 GNDA 0.03537f
C1750 bgr_0.V_mir2.t10 GNDA 0.03537f
C1751 bgr_0.V_mir2.n7 GNDA 0.08097f
C1752 bgr_0.V_mir2.n8 GNDA 0.201563f
C1753 bgr_0.V_mir2.t15 GNDA 0.042444f
C1754 bgr_0.V_mir2.t21 GNDA 0.042444f
C1755 bgr_0.V_mir2.t17 GNDA 0.06851f
C1756 bgr_0.V_mir2.n9 GNDA 0.076506f
C1757 bgr_0.V_mir2.n10 GNDA 0.052264f
C1758 bgr_0.V_mir2.t7 GNDA 0.053881f
C1759 bgr_0.V_mir2.n11 GNDA 0.081315f
C1760 bgr_0.V_mir2.t16 GNDA 0.03537f
C1761 bgr_0.V_mir2.t8 GNDA 0.03537f
C1762 bgr_0.V_mir2.n12 GNDA 0.08097f
C1763 bgr_0.V_mir2.n13 GNDA 0.203577f
C1764 bgr_0.V_mir2.n14 GNDA 0.699157f
C1765 bgr_0.V_mir2.n15 GNDA 0.09373f
C1766 bgr_0.V_mir2.t13 GNDA 0.042444f
C1767 bgr_0.V_mir2.t19 GNDA 0.042444f
C1768 bgr_0.V_mir2.t22 GNDA 0.06851f
C1769 bgr_0.V_mir2.n16 GNDA 0.076506f
C1770 bgr_0.V_mir2.n17 GNDA 0.052264f
C1771 bgr_0.V_mir2.t11 GNDA 0.053881f
C1772 bgr_0.V_mir2.n18 GNDA 0.081315f
C1773 bgr_0.V_mir2.n19 GNDA 0.156007f
C1774 bgr_0.V_mir2.t12 GNDA 0.03537f
C1775 bgr_0.V_mir2.n20 GNDA 0.08097f
C1776 bgr_0.V_mir2.t14 GNDA 0.03537f
C1777 two_stage_opamp_dummy_magic_0.cap_res_X.t2 GNDA 0.344645f
C1778 two_stage_opamp_dummy_magic_0.cap_res_X.t39 GNDA 0.167175f
C1779 two_stage_opamp_dummy_magic_0.cap_res_X.n0 GNDA 0.198327f
C1780 two_stage_opamp_dummy_magic_0.cap_res_X.t38 GNDA 0.344645f
C1781 two_stage_opamp_dummy_magic_0.cap_res_X.t77 GNDA 0.167175f
C1782 two_stage_opamp_dummy_magic_0.cap_res_X.n1 GNDA 0.216884f
C1783 two_stage_opamp_dummy_magic_0.cap_res_X.t23 GNDA 0.344645f
C1784 two_stage_opamp_dummy_magic_0.cap_res_X.t61 GNDA 0.167175f
C1785 two_stage_opamp_dummy_magic_0.cap_res_X.n2 GNDA 0.216884f
C1786 two_stage_opamp_dummy_magic_0.cap_res_X.t56 GNDA 0.344645f
C1787 two_stage_opamp_dummy_magic_0.cap_res_X.t96 GNDA 0.167175f
C1788 two_stage_opamp_dummy_magic_0.cap_res_X.n3 GNDA 0.216884f
C1789 two_stage_opamp_dummy_magic_0.cap_res_X.t94 GNDA 0.344645f
C1790 two_stage_opamp_dummy_magic_0.cap_res_X.t83 GNDA 0.345795f
C1791 two_stage_opamp_dummy_magic_0.cap_res_X.t44 GNDA 0.364353f
C1792 two_stage_opamp_dummy_magic_0.cap_res_X.t136 GNDA 0.364353f
C1793 two_stage_opamp_dummy_magic_0.cap_res_X.t32 GNDA 0.364353f
C1794 two_stage_opamp_dummy_magic_0.cap_res_X.t130 GNDA 0.185733f
C1795 two_stage_opamp_dummy_magic_0.cap_res_X.n4 GNDA 0.216884f
C1796 two_stage_opamp_dummy_magic_0.cap_res_X.t72 GNDA 0.344645f
C1797 two_stage_opamp_dummy_magic_0.cap_res_X.t131 GNDA 0.345795f
C1798 two_stage_opamp_dummy_magic_0.cap_res_X.t97 GNDA 0.364353f
C1799 two_stage_opamp_dummy_magic_0.cap_res_X.t117 GNDA 0.364353f
C1800 two_stage_opamp_dummy_magic_0.cap_res_X.t14 GNDA 0.364353f
C1801 two_stage_opamp_dummy_magic_0.cap_res_X.t113 GNDA 0.185733f
C1802 two_stage_opamp_dummy_magic_0.cap_res_X.n5 GNDA 0.216884f
C1803 two_stage_opamp_dummy_magic_0.cap_res_X.t118 GNDA 0.345795f
C1804 two_stage_opamp_dummy_magic_0.cap_res_X.t138 GNDA 0.347048f
C1805 two_stage_opamp_dummy_magic_0.cap_res_X.t74 GNDA 0.345795f
C1806 two_stage_opamp_dummy_magic_0.cap_res_X.t101 GNDA 0.348506f
C1807 two_stage_opamp_dummy_magic_0.cap_res_X.t62 GNDA 0.37905f
C1808 two_stage_opamp_dummy_magic_0.cap_res_X.t123 GNDA 0.345795f
C1809 two_stage_opamp_dummy_magic_0.cap_res_X.t106 GNDA 0.347048f
C1810 two_stage_opamp_dummy_magic_0.cap_res_X.t21 GNDA 0.345795f
C1811 two_stage_opamp_dummy_magic_0.cap_res_X.t37 GNDA 0.347048f
C1812 two_stage_opamp_dummy_magic_0.cap_res_X.t89 GNDA 0.345795f
C1813 two_stage_opamp_dummy_magic_0.cap_res_X.t70 GNDA 0.347048f
C1814 two_stage_opamp_dummy_magic_0.cap_res_X.t121 GNDA 0.345795f
C1815 two_stage_opamp_dummy_magic_0.cap_res_X.t6 GNDA 0.347048f
C1816 two_stage_opamp_dummy_magic_0.cap_res_X.t63 GNDA 0.345795f
C1817 two_stage_opamp_dummy_magic_0.cap_res_X.t115 GNDA 0.347048f
C1818 two_stage_opamp_dummy_magic_0.cap_res_X.t93 GNDA 0.345795f
C1819 two_stage_opamp_dummy_magic_0.cap_res_X.t40 GNDA 0.347048f
C1820 two_stage_opamp_dummy_magic_0.cap_res_X.t103 GNDA 0.345795f
C1821 two_stage_opamp_dummy_magic_0.cap_res_X.t16 GNDA 0.347048f
C1822 two_stage_opamp_dummy_magic_0.cap_res_X.t128 GNDA 0.345795f
C1823 two_stage_opamp_dummy_magic_0.cap_res_X.t78 GNDA 0.347048f
C1824 two_stage_opamp_dummy_magic_0.cap_res_X.t68 GNDA 0.345795f
C1825 two_stage_opamp_dummy_magic_0.cap_res_X.t119 GNDA 0.347048f
C1826 two_stage_opamp_dummy_magic_0.cap_res_X.t100 GNDA 0.345795f
C1827 two_stage_opamp_dummy_magic_0.cap_res_X.t49 GNDA 0.347048f
C1828 two_stage_opamp_dummy_magic_0.cap_res_X.t109 GNDA 0.345795f
C1829 two_stage_opamp_dummy_magic_0.cap_res_X.t22 GNDA 0.347048f
C1830 two_stage_opamp_dummy_magic_0.cap_res_X.t137 GNDA 0.345795f
C1831 two_stage_opamp_dummy_magic_0.cap_res_X.t87 GNDA 0.347048f
C1832 two_stage_opamp_dummy_magic_0.cap_res_X.t9 GNDA 0.345795f
C1833 two_stage_opamp_dummy_magic_0.cap_res_X.t59 GNDA 0.347048f
C1834 two_stage_opamp_dummy_magic_0.cap_res_X.t36 GNDA 0.345795f
C1835 two_stage_opamp_dummy_magic_0.cap_res_X.t124 GNDA 0.347048f
C1836 two_stage_opamp_dummy_magic_0.cap_res_X.t114 GNDA 0.345795f
C1837 two_stage_opamp_dummy_magic_0.cap_res_X.t24 GNDA 0.347048f
C1838 two_stage_opamp_dummy_magic_0.cap_res_X.t5 GNDA 0.345795f
C1839 two_stage_opamp_dummy_magic_0.cap_res_X.t92 GNDA 0.347048f
C1840 two_stage_opamp_dummy_magic_0.cap_res_X.t15 GNDA 0.345795f
C1841 two_stage_opamp_dummy_magic_0.cap_res_X.t64 GNDA 0.347048f
C1842 two_stage_opamp_dummy_magic_0.cap_res_X.t42 GNDA 0.345795f
C1843 two_stage_opamp_dummy_magic_0.cap_res_X.t127 GNDA 0.347048f
C1844 two_stage_opamp_dummy_magic_0.cap_res_X.t53 GNDA 0.345795f
C1845 two_stage_opamp_dummy_magic_0.cap_res_X.t105 GNDA 0.347048f
C1846 two_stage_opamp_dummy_magic_0.cap_res_X.t81 GNDA 0.345795f
C1847 two_stage_opamp_dummy_magic_0.cap_res_X.t31 GNDA 0.347048f
C1848 two_stage_opamp_dummy_magic_0.cap_res_X.t90 GNDA 0.345795f
C1849 two_stage_opamp_dummy_magic_0.cap_res_X.t3 GNDA 0.347048f
C1850 two_stage_opamp_dummy_magic_0.cap_res_X.t122 GNDA 0.345795f
C1851 two_stage_opamp_dummy_magic_0.cap_res_X.t73 GNDA 0.347048f
C1852 two_stage_opamp_dummy_magic_0.cap_res_X.t58 GNDA 0.345795f
C1853 two_stage_opamp_dummy_magic_0.cap_res_X.t111 GNDA 0.347048f
C1854 two_stage_opamp_dummy_magic_0.cap_res_X.t88 GNDA 0.345795f
C1855 two_stage_opamp_dummy_magic_0.cap_res_X.t35 GNDA 0.347048f
C1856 two_stage_opamp_dummy_magic_0.cap_res_X.t98 GNDA 0.345795f
C1857 two_stage_opamp_dummy_magic_0.cap_res_X.t10 GNDA 0.347048f
C1858 two_stage_opamp_dummy_magic_0.cap_res_X.t125 GNDA 0.345795f
C1859 two_stage_opamp_dummy_magic_0.cap_res_X.t76 GNDA 0.347048f
C1860 two_stage_opamp_dummy_magic_0.cap_res_X.t133 GNDA 0.345795f
C1861 two_stage_opamp_dummy_magic_0.cap_res_X.t45 GNDA 0.347048f
C1862 two_stage_opamp_dummy_magic_0.cap_res_X.t28 GNDA 0.345795f
C1863 two_stage_opamp_dummy_magic_0.cap_res_X.t120 GNDA 0.347048f
C1864 two_stage_opamp_dummy_magic_0.cap_res_X.t7 GNDA 0.345795f
C1865 two_stage_opamp_dummy_magic_0.cap_res_X.t71 GNDA 0.362749f
C1866 two_stage_opamp_dummy_magic_0.cap_res_X.t95 GNDA 0.345795f
C1867 two_stage_opamp_dummy_magic_0.cap_res_X.t107 GNDA 0.185733f
C1868 two_stage_opamp_dummy_magic_0.cap_res_X.n6 GNDA 0.198781f
C1869 two_stage_opamp_dummy_magic_0.cap_res_X.t134 GNDA 0.345795f
C1870 two_stage_opamp_dummy_magic_0.cap_res_X.t20 GNDA 0.185733f
C1871 two_stage_opamp_dummy_magic_0.cap_res_X.n7 GNDA 0.197177f
C1872 two_stage_opamp_dummy_magic_0.cap_res_X.t85 GNDA 0.345795f
C1873 two_stage_opamp_dummy_magic_0.cap_res_X.t52 GNDA 0.185733f
C1874 two_stage_opamp_dummy_magic_0.cap_res_X.n8 GNDA 0.197177f
C1875 two_stage_opamp_dummy_magic_0.cap_res_X.t33 GNDA 0.345795f
C1876 two_stage_opamp_dummy_magic_0.cap_res_X.t84 GNDA 0.185733f
C1877 two_stage_opamp_dummy_magic_0.cap_res_X.n9 GNDA 0.197177f
C1878 two_stage_opamp_dummy_magic_0.cap_res_X.t75 GNDA 0.345795f
C1879 two_stage_opamp_dummy_magic_0.cap_res_X.t132 GNDA 0.185733f
C1880 two_stage_opamp_dummy_magic_0.cap_res_X.n10 GNDA 0.197177f
C1881 two_stage_opamp_dummy_magic_0.cap_res_X.t27 GNDA 0.345795f
C1882 two_stage_opamp_dummy_magic_0.cap_res_X.t30 GNDA 0.185733f
C1883 two_stage_opamp_dummy_magic_0.cap_res_X.n11 GNDA 0.197177f
C1884 two_stage_opamp_dummy_magic_0.cap_res_X.t116 GNDA 0.345795f
C1885 two_stage_opamp_dummy_magic_0.cap_res_X.t69 GNDA 0.185733f
C1886 two_stage_opamp_dummy_magic_0.cap_res_X.n12 GNDA 0.197177f
C1887 two_stage_opamp_dummy_magic_0.cap_res_X.t66 GNDA 0.345795f
C1888 two_stage_opamp_dummy_magic_0.cap_res_X.t104 GNDA 0.185733f
C1889 two_stage_opamp_dummy_magic_0.cap_res_X.n13 GNDA 0.197177f
C1890 two_stage_opamp_dummy_magic_0.cap_res_X.t110 GNDA 0.345795f
C1891 two_stage_opamp_dummy_magic_0.cap_res_X.t17 GNDA 0.185733f
C1892 two_stage_opamp_dummy_magic_0.cap_res_X.n14 GNDA 0.197177f
C1893 two_stage_opamp_dummy_magic_0.cap_res_X.t129 GNDA 0.345795f
C1894 two_stage_opamp_dummy_magic_0.cap_res_X.t79 GNDA 0.347048f
C1895 two_stage_opamp_dummy_magic_0.cap_res_X.t50 GNDA 0.345795f
C1896 two_stage_opamp_dummy_magic_0.cap_res_X.t8 GNDA 0.347048f
C1897 two_stage_opamp_dummy_magic_0.cap_res_X.t57 GNDA 0.167175f
C1898 two_stage_opamp_dummy_magic_0.cap_res_X.n15 GNDA 0.215631f
C1899 two_stage_opamp_dummy_magic_0.cap_res_X.t48 GNDA 0.184584f
C1900 two_stage_opamp_dummy_magic_0.cap_res_X.n16 GNDA 0.234189f
C1901 two_stage_opamp_dummy_magic_0.cap_res_X.t80 GNDA 0.184584f
C1902 two_stage_opamp_dummy_magic_0.cap_res_X.n17 GNDA 0.251494f
C1903 two_stage_opamp_dummy_magic_0.cap_res_X.t41 GNDA 0.184584f
C1904 two_stage_opamp_dummy_magic_0.cap_res_X.n18 GNDA 0.251494f
C1905 two_stage_opamp_dummy_magic_0.cap_res_X.t4 GNDA 0.184584f
C1906 two_stage_opamp_dummy_magic_0.cap_res_X.n19 GNDA 0.251494f
C1907 two_stage_opamp_dummy_magic_0.cap_res_X.t34 GNDA 0.184584f
C1908 two_stage_opamp_dummy_magic_0.cap_res_X.n20 GNDA 0.251494f
C1909 two_stage_opamp_dummy_magic_0.cap_res_X.t135 GNDA 0.184584f
C1910 two_stage_opamp_dummy_magic_0.cap_res_X.n21 GNDA 0.251494f
C1911 two_stage_opamp_dummy_magic_0.cap_res_X.t99 GNDA 0.184584f
C1912 two_stage_opamp_dummy_magic_0.cap_res_X.n22 GNDA 0.251494f
C1913 two_stage_opamp_dummy_magic_0.cap_res_X.t60 GNDA 0.184584f
C1914 two_stage_opamp_dummy_magic_0.cap_res_X.n23 GNDA 0.251494f
C1915 two_stage_opamp_dummy_magic_0.cap_res_X.t91 GNDA 0.184584f
C1916 two_stage_opamp_dummy_magic_0.cap_res_X.n24 GNDA 0.251494f
C1917 two_stage_opamp_dummy_magic_0.cap_res_X.t55 GNDA 0.184584f
C1918 two_stage_opamp_dummy_magic_0.cap_res_X.n25 GNDA 0.251494f
C1919 two_stage_opamp_dummy_magic_0.cap_res_X.t18 GNDA 0.184584f
C1920 two_stage_opamp_dummy_magic_0.cap_res_X.n26 GNDA 0.251494f
C1921 two_stage_opamp_dummy_magic_0.cap_res_X.t47 GNDA 0.184584f
C1922 two_stage_opamp_dummy_magic_0.cap_res_X.n27 GNDA 0.251494f
C1923 two_stage_opamp_dummy_magic_0.cap_res_X.t12 GNDA 0.184584f
C1924 two_stage_opamp_dummy_magic_0.cap_res_X.n28 GNDA 0.251494f
C1925 two_stage_opamp_dummy_magic_0.cap_res_X.t108 GNDA 0.184584f
C1926 two_stage_opamp_dummy_magic_0.cap_res_X.n29 GNDA 0.251494f
C1927 two_stage_opamp_dummy_magic_0.cap_res_X.t1 GNDA 0.184584f
C1928 two_stage_opamp_dummy_magic_0.cap_res_X.n30 GNDA 0.251494f
C1929 two_stage_opamp_dummy_magic_0.cap_res_X.t102 GNDA 0.184584f
C1930 two_stage_opamp_dummy_magic_0.cap_res_X.n31 GNDA 0.234189f
C1931 two_stage_opamp_dummy_magic_0.cap_res_X.t25 GNDA 0.344645f
C1932 two_stage_opamp_dummy_magic_0.cap_res_X.t65 GNDA 0.167175f
C1933 two_stage_opamp_dummy_magic_0.cap_res_X.n32 GNDA 0.216884f
C1934 two_stage_opamp_dummy_magic_0.cap_res_X.t43 GNDA 0.344645f
C1935 two_stage_opamp_dummy_magic_0.cap_res_X.t82 GNDA 0.167175f
C1936 two_stage_opamp_dummy_magic_0.cap_res_X.n33 GNDA 0.216884f
C1937 two_stage_opamp_dummy_magic_0.cap_res_X.t11 GNDA 0.344645f
C1938 two_stage_opamp_dummy_magic_0.cap_res_X.t67 GNDA 0.345795f
C1939 two_stage_opamp_dummy_magic_0.cap_res_X.t26 GNDA 0.364353f
C1940 two_stage_opamp_dummy_magic_0.cap_res_X.t54 GNDA 0.364353f
C1941 two_stage_opamp_dummy_magic_0.cap_res_X.t86 GNDA 0.364353f
C1942 two_stage_opamp_dummy_magic_0.cap_res_X.t46 GNDA 0.185733f
C1943 two_stage_opamp_dummy_magic_0.cap_res_X.n34 GNDA 0.216884f
C1944 two_stage_opamp_dummy_magic_0.cap_res_X.t112 GNDA 0.344645f
C1945 two_stage_opamp_dummy_magic_0.cap_res_X.n35 GNDA 0.216884f
C1946 two_stage_opamp_dummy_magic_0.cap_res_X.t13 GNDA 0.185733f
C1947 two_stage_opamp_dummy_magic_0.cap_res_X.t51 GNDA 0.364353f
C1948 two_stage_opamp_dummy_magic_0.cap_res_X.t19 GNDA 0.364353f
C1949 two_stage_opamp_dummy_magic_0.cap_res_X.t126 GNDA 0.364353f
C1950 two_stage_opamp_dummy_magic_0.cap_res_X.t29 GNDA 0.337351f
C1951 two_stage_opamp_dummy_magic_0.cap_res_X.t0 GNDA 0.298183f
C1952 VOUT-.t17 GNDA 0.051003f
C1953 VOUT-.t9 GNDA 0.051003f
C1954 VOUT-.n0 GNDA 0.235943f
C1955 VOUT-.t13 GNDA 0.051003f
C1956 VOUT-.t18 GNDA 0.051003f
C1957 VOUT-.n1 GNDA 0.235153f
C1958 VOUT-.n2 GNDA 0.145313f
C1959 VOUT-.t0 GNDA 0.051003f
C1960 VOUT-.t16 GNDA 0.051003f
C1961 VOUT-.n3 GNDA 0.235153f
C1962 VOUT-.n4 GNDA 0.089445f
C1963 VOUT-.t12 GNDA 0.084326f
C1964 VOUT-.n5 GNDA 0.119504f
C1965 VOUT-.t14 GNDA 0.043717f
C1966 VOUT-.t11 GNDA 0.043717f
C1967 VOUT-.n6 GNDA 0.175711f
C1968 VOUT-.t2 GNDA 0.043717f
C1969 VOUT-.t15 GNDA 0.043717f
C1970 VOUT-.n7 GNDA 0.17571f
C1971 VOUT-.t5 GNDA 0.043717f
C1972 VOUT-.t10 GNDA 0.043717f
C1973 VOUT-.n8 GNDA 0.175387f
C1974 VOUT-.n9 GNDA 0.172777f
C1975 VOUT-.t1 GNDA 0.043717f
C1976 VOUT-.t7 GNDA 0.043717f
C1977 VOUT-.n10 GNDA 0.175387f
C1978 VOUT-.n11 GNDA 0.0891f
C1979 VOUT-.t6 GNDA 0.043717f
C1980 VOUT-.t3 GNDA 0.043717f
C1981 VOUT-.n12 GNDA 0.175387f
C1982 VOUT-.n13 GNDA 0.0891f
C1983 VOUT-.n14 GNDA 0.105535f
C1984 VOUT-.t8 GNDA 0.043717f
C1985 VOUT-.t4 GNDA 0.043717f
C1986 VOUT-.n15 GNDA 0.17324f
C1987 VOUT-.n16 GNDA 0.211953f
C1988 VOUT-.t100 GNDA 0.291446f
C1989 VOUT-.t107 GNDA 0.29641f
C1990 VOUT-.t149 GNDA 0.291446f
C1991 VOUT-.n17 GNDA 0.195405f
C1992 VOUT-.n18 GNDA 0.127508f
C1993 VOUT-.t47 GNDA 0.295788f
C1994 VOUT-.t91 GNDA 0.295788f
C1995 VOUT-.t41 GNDA 0.295788f
C1996 VOUT-.t130 GNDA 0.295788f
C1997 VOUT-.t82 GNDA 0.295788f
C1998 VOUT-.t124 GNDA 0.295788f
C1999 VOUT-.t72 GNDA 0.295788f
C2000 VOUT-.t23 GNDA 0.295788f
C2001 VOUT-.t62 GNDA 0.295788f
C2002 VOUT-.t150 GNDA 0.295788f
C2003 VOUT-.t86 GNDA 0.291446f
C2004 VOUT-.n19 GNDA 0.196026f
C2005 VOUT-.t50 GNDA 0.291446f
C2006 VOUT-.n20 GNDA 0.250673f
C2007 VOUT-.t137 GNDA 0.291446f
C2008 VOUT-.n21 GNDA 0.250673f
C2009 VOUT-.t105 GNDA 0.291446f
C2010 VOUT-.n22 GNDA 0.250673f
C2011 VOUT-.t73 GNDA 0.291446f
C2012 VOUT-.n23 GNDA 0.250673f
C2013 VOUT-.t25 GNDA 0.291446f
C2014 VOUT-.n24 GNDA 0.250673f
C2015 VOUT-.t127 GNDA 0.291446f
C2016 VOUT-.n25 GNDA 0.250673f
C2017 VOUT-.t88 GNDA 0.291446f
C2018 VOUT-.n26 GNDA 0.250673f
C2019 VOUT-.t53 GNDA 0.291446f
C2020 VOUT-.n27 GNDA 0.250673f
C2021 VOUT-.t140 GNDA 0.291446f
C2022 VOUT-.n28 GNDA 0.250673f
C2023 VOUT-.t109 GNDA 0.291446f
C2024 VOUT-.t28 GNDA 0.29641f
C2025 VOUT-.t78 GNDA 0.291446f
C2026 VOUT-.n29 GNDA 0.195405f
C2027 VOUT-.n30 GNDA 0.2368f
C2028 VOUT-.t24 GNDA 0.29641f
C2029 VOUT-.t112 GNDA 0.291446f
C2030 VOUT-.n31 GNDA 0.195405f
C2031 VOUT-.t77 GNDA 0.291446f
C2032 VOUT-.t129 GNDA 0.29641f
C2033 VOUT-.t37 GNDA 0.291446f
C2034 VOUT-.n32 GNDA 0.195405f
C2035 VOUT-.n33 GNDA 0.2368f
C2036 VOUT-.t59 GNDA 0.29641f
C2037 VOUT-.t147 GNDA 0.291446f
C2038 VOUT-.n34 GNDA 0.195405f
C2039 VOUT-.t116 GNDA 0.291446f
C2040 VOUT-.t32 GNDA 0.29641f
C2041 VOUT-.t81 GNDA 0.291446f
C2042 VOUT-.n35 GNDA 0.195405f
C2043 VOUT-.n36 GNDA 0.2368f
C2044 VOUT-.t99 GNDA 0.29641f
C2045 VOUT-.t46 GNDA 0.291446f
C2046 VOUT-.n37 GNDA 0.195405f
C2047 VOUT-.t153 GNDA 0.291446f
C2048 VOUT-.t69 GNDA 0.29641f
C2049 VOUT-.t122 GNDA 0.291446f
C2050 VOUT-.n38 GNDA 0.195405f
C2051 VOUT-.n39 GNDA 0.2368f
C2052 VOUT-.t67 GNDA 0.29641f
C2053 VOUT-.t154 GNDA 0.291446f
C2054 VOUT-.n40 GNDA 0.195405f
C2055 VOUT-.t123 GNDA 0.291446f
C2056 VOUT-.t35 GNDA 0.29641f
C2057 VOUT-.t84 GNDA 0.291446f
C2058 VOUT-.n41 GNDA 0.195405f
C2059 VOUT-.n42 GNDA 0.2368f
C2060 VOUT-.t104 GNDA 0.29641f
C2061 VOUT-.t52 GNDA 0.291446f
C2062 VOUT-.n43 GNDA 0.195405f
C2063 VOUT-.t22 GNDA 0.291446f
C2064 VOUT-.t76 GNDA 0.29641f
C2065 VOUT-.t126 GNDA 0.291446f
C2066 VOUT-.n44 GNDA 0.195405f
C2067 VOUT-.n45 GNDA 0.2368f
C2068 VOUT-.t95 GNDA 0.291446f
C2069 VOUT-.t83 GNDA 0.29641f
C2070 VOUT-.t56 GNDA 0.291446f
C2071 VOUT-.n46 GNDA 0.195405f
C2072 VOUT-.n47 GNDA 0.127508f
C2073 VOUT-.t132 GNDA 0.295788f
C2074 VOUT-.t114 GNDA 0.295788f
C2075 VOUT-.t90 GNDA 0.29641f
C2076 VOUT-.t131 GNDA 0.291446f
C2077 VOUT-.n48 GNDA 0.195405f
C2078 VOUT-.t103 GNDA 0.291446f
C2079 VOUT-.n49 GNDA 0.127508f
C2080 VOUT-.t71 GNDA 0.291446f
C2081 VOUT-.n50 GNDA 0.122954f
C2082 VOUT-.t146 GNDA 0.295788f
C2083 VOUT-.t128 GNDA 0.29641f
C2084 VOUT-.t31 GNDA 0.291446f
C2085 VOUT-.n51 GNDA 0.195405f
C2086 VOUT-.t138 GNDA 0.291446f
C2087 VOUT-.n52 GNDA 0.127508f
C2088 VOUT-.t106 GNDA 0.291446f
C2089 VOUT-.n53 GNDA 0.122954f
C2090 VOUT-.t45 GNDA 0.295788f
C2091 VOUT-.t26 GNDA 0.29641f
C2092 VOUT-.t60 GNDA 0.291446f
C2093 VOUT-.n54 GNDA 0.195405f
C2094 VOUT-.t40 GNDA 0.291446f
C2095 VOUT-.n55 GNDA 0.127508f
C2096 VOUT-.t143 GNDA 0.291446f
C2097 VOUT-.n56 GNDA 0.122954f
C2098 VOUT-.t85 GNDA 0.295788f
C2099 VOUT-.t74 GNDA 0.29641f
C2100 VOUT-.t113 GNDA 0.291446f
C2101 VOUT-.n57 GNDA 0.195405f
C2102 VOUT-.t21 GNDA 0.291446f
C2103 VOUT-.n58 GNDA 0.127508f
C2104 VOUT-.t125 GNDA 0.291446f
C2105 VOUT-.n59 GNDA 0.122954f
C2106 VOUT-.t63 GNDA 0.295788f
C2107 VOUT-.t101 GNDA 0.295788f
C2108 VOUT-.t134 GNDA 0.295788f
C2109 VOUT-.t119 GNDA 0.295788f
C2110 VOUT-.t155 GNDA 0.295788f
C2111 VOUT-.t118 GNDA 0.291446f
C2112 VOUT-.n60 GNDA 0.196026f
C2113 VOUT-.t80 GNDA 0.291446f
C2114 VOUT-.n61 GNDA 0.250673f
C2115 VOUT-.t96 GNDA 0.291446f
C2116 VOUT-.n62 GNDA 0.250673f
C2117 VOUT-.t61 GNDA 0.291446f
C2118 VOUT-.n63 GNDA 0.250673f
C2119 VOUT-.t27 GNDA 0.291446f
C2120 VOUT-.n64 GNDA 0.309872f
C2121 VOUT-.t44 GNDA 0.291446f
C2122 VOUT-.n65 GNDA 0.309872f
C2123 VOUT-.t144 GNDA 0.291446f
C2124 VOUT-.n66 GNDA 0.309872f
C2125 VOUT-.t111 GNDA 0.291446f
C2126 VOUT-.n67 GNDA 0.309872f
C2127 VOUT-.t75 GNDA 0.291446f
C2128 VOUT-.n68 GNDA 0.250673f
C2129 VOUT-.t92 GNDA 0.291446f
C2130 VOUT-.n69 GNDA 0.250673f
C2131 VOUT-.t55 GNDA 0.291446f
C2132 VOUT-.t39 GNDA 0.29641f
C2133 VOUT-.t19 GNDA 0.291446f
C2134 VOUT-.n70 GNDA 0.195405f
C2135 VOUT-.n71 GNDA 0.2368f
C2136 VOUT-.t34 GNDA 0.29641f
C2137 VOUT-.t51 GNDA 0.291446f
C2138 VOUT-.n72 GNDA 0.195405f
C2139 VOUT-.t156 GNDA 0.291446f
C2140 VOUT-.t136 GNDA 0.29641f
C2141 VOUT-.t120 GNDA 0.291446f
C2142 VOUT-.n73 GNDA 0.195405f
C2143 VOUT-.n74 GNDA 0.2368f
C2144 VOUT-.t68 GNDA 0.29641f
C2145 VOUT-.t87 GNDA 0.291446f
C2146 VOUT-.n75 GNDA 0.195405f
C2147 VOUT-.t49 GNDA 0.291446f
C2148 VOUT-.t36 GNDA 0.29641f
C2149 VOUT-.t151 GNDA 0.291446f
C2150 VOUT-.n76 GNDA 0.195405f
C2151 VOUT-.n77 GNDA 0.2368f
C2152 VOUT-.t94 GNDA 0.29641f
C2153 VOUT-.t42 GNDA 0.291446f
C2154 VOUT-.n78 GNDA 0.195405f
C2155 VOUT-.t145 GNDA 0.291446f
C2156 VOUT-.t64 GNDA 0.29641f
C2157 VOUT-.t117 GNDA 0.291446f
C2158 VOUT-.n79 GNDA 0.195405f
C2159 VOUT-.n80 GNDA 0.2368f
C2160 VOUT-.t54 GNDA 0.29641f
C2161 VOUT-.t141 GNDA 0.291446f
C2162 VOUT-.n81 GNDA 0.195405f
C2163 VOUT-.t110 GNDA 0.291446f
C2164 VOUT-.t29 GNDA 0.29641f
C2165 VOUT-.t79 GNDA 0.291446f
C2166 VOUT-.n82 GNDA 0.195405f
C2167 VOUT-.n83 GNDA 0.2368f
C2168 VOUT-.t89 GNDA 0.29641f
C2169 VOUT-.t38 GNDA 0.291446f
C2170 VOUT-.n84 GNDA 0.195405f
C2171 VOUT-.t139 GNDA 0.291446f
C2172 VOUT-.t57 GNDA 0.29641f
C2173 VOUT-.t108 GNDA 0.291446f
C2174 VOUT-.n85 GNDA 0.195405f
C2175 VOUT-.n86 GNDA 0.2368f
C2176 VOUT-.t48 GNDA 0.29641f
C2177 VOUT-.t135 GNDA 0.291446f
C2178 VOUT-.n87 GNDA 0.195405f
C2179 VOUT-.t102 GNDA 0.291446f
C2180 VOUT-.t20 GNDA 0.29641f
C2181 VOUT-.t70 GNDA 0.291446f
C2182 VOUT-.n88 GNDA 0.195405f
C2183 VOUT-.n89 GNDA 0.2368f
C2184 VOUT-.t148 GNDA 0.29641f
C2185 VOUT-.t98 GNDA 0.291446f
C2186 VOUT-.n90 GNDA 0.195405f
C2187 VOUT-.t66 GNDA 0.291446f
C2188 VOUT-.t121 GNDA 0.29641f
C2189 VOUT-.t33 GNDA 0.291446f
C2190 VOUT-.n91 GNDA 0.195405f
C2191 VOUT-.n92 GNDA 0.2368f
C2192 VOUT-.t43 GNDA 0.29641f
C2193 VOUT-.t133 GNDA 0.291446f
C2194 VOUT-.n93 GNDA 0.195405f
C2195 VOUT-.t97 GNDA 0.291446f
C2196 VOUT-.t152 GNDA 0.29641f
C2197 VOUT-.t65 GNDA 0.291446f
C2198 VOUT-.n94 GNDA 0.195405f
C2199 VOUT-.n95 GNDA 0.2368f
C2200 VOUT-.t115 GNDA 0.29641f
C2201 VOUT-.t30 GNDA 0.291446f
C2202 VOUT-.n96 GNDA 0.195405f
C2203 VOUT-.t58 GNDA 0.291446f
C2204 VOUT-.n97 GNDA 0.2368f
C2205 VOUT-.t93 GNDA 0.291446f
C2206 VOUT-.n98 GNDA 0.127508f
C2207 VOUT-.t142 GNDA 0.291446f
C2208 VOUT-.n99 GNDA 0.23878f
C2209 VOUT-.n100 GNDA 0.268998f
C2210 two_stage_opamp_dummy_magic_0.VD2.t15 GNDA 0.013877f
C2211 two_stage_opamp_dummy_magic_0.VD2.t1 GNDA 0.013877f
C2212 two_stage_opamp_dummy_magic_0.VD2.t7 GNDA 0.013877f
C2213 two_stage_opamp_dummy_magic_0.VD2.n0 GNDA 0.048872f
C2214 two_stage_opamp_dummy_magic_0.VD2.t17 GNDA 0.013877f
C2215 two_stage_opamp_dummy_magic_0.VD2.t8 GNDA 0.013877f
C2216 two_stage_opamp_dummy_magic_0.VD2.n1 GNDA 0.047884f
C2217 two_stage_opamp_dummy_magic_0.VD2.n2 GNDA 0.193373f
C2218 two_stage_opamp_dummy_magic_0.VD2.t3 GNDA 0.013877f
C2219 two_stage_opamp_dummy_magic_0.VD2.t18 GNDA 0.013877f
C2220 two_stage_opamp_dummy_magic_0.VD2.n3 GNDA 0.047884f
C2221 two_stage_opamp_dummy_magic_0.VD2.n4 GNDA 0.140662f
C2222 two_stage_opamp_dummy_magic_0.VD2.t21 GNDA 0.013877f
C2223 two_stage_opamp_dummy_magic_0.VD2.t4 GNDA 0.013877f
C2224 two_stage_opamp_dummy_magic_0.VD2.n5 GNDA 0.04687f
C2225 two_stage_opamp_dummy_magic_0.VD2.t5 GNDA 0.013877f
C2226 two_stage_opamp_dummy_magic_0.VD2.t16 GNDA 0.013877f
C2227 two_stage_opamp_dummy_magic_0.VD2.n6 GNDA 0.050131f
C2228 two_stage_opamp_dummy_magic_0.VD2.t13 GNDA 0.013877f
C2229 two_stage_opamp_dummy_magic_0.VD2.t10 GNDA 0.013877f
C2230 two_stage_opamp_dummy_magic_0.VD2.n7 GNDA 0.04969f
C2231 two_stage_opamp_dummy_magic_0.VD2.n8 GNDA 0.186051f
C2232 two_stage_opamp_dummy_magic_0.VD2.t0 GNDA 0.013877f
C2233 two_stage_opamp_dummy_magic_0.VD2.t9 GNDA 0.013877f
C2234 two_stage_opamp_dummy_magic_0.VD2.n9 GNDA 0.050131f
C2235 two_stage_opamp_dummy_magic_0.VD2.t20 GNDA 0.013877f
C2236 two_stage_opamp_dummy_magic_0.VD2.t14 GNDA 0.013877f
C2237 two_stage_opamp_dummy_magic_0.VD2.n10 GNDA 0.04969f
C2238 two_stage_opamp_dummy_magic_0.VD2.n11 GNDA 0.186051f
C2239 two_stage_opamp_dummy_magic_0.VD2.n12 GNDA 0.027755f
C2240 two_stage_opamp_dummy_magic_0.VD2.n13 GNDA 0.081264f
C2241 two_stage_opamp_dummy_magic_0.VD2.t2 GNDA 0.013877f
C2242 two_stage_opamp_dummy_magic_0.VD2.t12 GNDA 0.013877f
C2243 two_stage_opamp_dummy_magic_0.VD2.n14 GNDA 0.045463f
C2244 two_stage_opamp_dummy_magic_0.VD2.n15 GNDA 0.069533f
C2245 two_stage_opamp_dummy_magic_0.VD2.n16 GNDA 0.083264f
C2246 two_stage_opamp_dummy_magic_0.VD2.t11 GNDA 0.013877f
C2247 two_stage_opamp_dummy_magic_0.VD2.t6 GNDA 0.013877f
C2248 two_stage_opamp_dummy_magic_0.VD2.n17 GNDA 0.047884f
C2249 two_stage_opamp_dummy_magic_0.VD2.n18 GNDA 0.193373f
C2250 two_stage_opamp_dummy_magic_0.VD2.n19 GNDA 0.048872f
C2251 two_stage_opamp_dummy_magic_0.VD2.t19 GNDA 0.013877f
C2252 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 GNDA 0.033498f
C2253 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 GNDA 0.033498f
C2254 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 GNDA 0.084004f
C2255 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 GNDA 0.033498f
C2256 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 GNDA 0.033498f
C2257 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 GNDA 0.083562f
C2258 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 GNDA 0.566043f
C2259 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 GNDA 0.033498f
C2260 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 GNDA 0.033498f
C2261 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 GNDA 0.083562f
C2262 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 GNDA 0.594775f
C2263 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 GNDA 0.428693f
C2264 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 GNDA 0.066996f
C2265 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 GNDA 0.066996f
C2266 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 GNDA 0.196564f
C2267 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 GNDA 0.066996f
C2268 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 GNDA 0.066996f
C2269 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 GNDA 0.195672f
C2270 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 GNDA 0.676354f
C2271 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 GNDA 0.066996f
C2272 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 GNDA 0.066996f
C2273 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 GNDA 0.195672f
C2274 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 GNDA 0.350348f
C2275 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 GNDA 0.066996f
C2276 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 GNDA 0.066996f
C2277 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 GNDA 0.195672f
C2278 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 GNDA 0.350348f
C2279 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 GNDA 0.066996f
C2280 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 GNDA 0.066996f
C2281 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 GNDA 0.195672f
C2282 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 GNDA 0.505738f
C2283 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 GNDA 4.90775f
C2284 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 GNDA 3.90403f
C2285 bgr_0.V_CMFB_S3 GNDA 0.014596f
C2286 bgr_0.cap_res1.t7 GNDA 0.417173f
C2287 bgr_0.cap_res1.t11 GNDA 0.418684f
C2288 bgr_0.cap_res1.t1 GNDA 0.417173f
C2289 bgr_0.cap_res1.t15 GNDA 0.418684f
C2290 bgr_0.cap_res1.t4 GNDA 0.417173f
C2291 bgr_0.cap_res1.t8 GNDA 0.418684f
C2292 bgr_0.cap_res1.t16 GNDA 0.417173f
C2293 bgr_0.cap_res1.t10 GNDA 0.418684f
C2294 bgr_0.cap_res1.t9 GNDA 0.417173f
C2295 bgr_0.cap_res1.t13 GNDA 0.418684f
C2296 bgr_0.cap_res1.t2 GNDA 0.417173f
C2297 bgr_0.cap_res1.t17 GNDA 0.418684f
C2298 bgr_0.cap_res1.t14 GNDA 0.417173f
C2299 bgr_0.cap_res1.t20 GNDA 0.418684f
C2300 bgr_0.cap_res1.t6 GNDA 0.417173f
C2301 bgr_0.cap_res1.t3 GNDA 0.418684f
C2302 bgr_0.cap_res1.n0 GNDA 0.279631f
C2303 bgr_0.cap_res1.t5 GNDA 0.222685f
C2304 bgr_0.cap_res1.n1 GNDA 0.303406f
C2305 bgr_0.cap_res1.t19 GNDA 0.222685f
C2306 bgr_0.cap_res1.n2 GNDA 0.303406f
C2307 bgr_0.cap_res1.t12 GNDA 0.222685f
C2308 bgr_0.cap_res1.n3 GNDA 0.303406f
C2309 bgr_0.cap_res1.t18 GNDA 0.649059f
C2310 bgr_0.cap_res1.t0 GNDA 0.10618f
C2311 bgr_0.1st_Vout_1.n0 GNDA 0.573726f
C2312 bgr_0.1st_Vout_1.n1 GNDA 1.42916f
C2313 bgr_0.1st_Vout_1.n2 GNDA 1.78489f
C2314 bgr_0.1st_Vout_1.n3 GNDA 0.125562f
C2315 bgr_0.1st_Vout_1.t20 GNDA 0.352846f
C2316 bgr_0.1st_Vout_1.t11 GNDA 0.346937f
C2317 bgr_0.1st_Vout_1.t32 GNDA 0.346937f
C2318 bgr_0.1st_Vout_1.t29 GNDA 0.352846f
C2319 bgr_0.1st_Vout_1.t34 GNDA 0.346937f
C2320 bgr_0.1st_Vout_1.t25 GNDA 0.352846f
C2321 bgr_0.1st_Vout_1.t21 GNDA 0.346937f
C2322 bgr_0.1st_Vout_1.t12 GNDA 0.346937f
C2323 bgr_0.1st_Vout_1.t35 GNDA 0.352846f
C2324 bgr_0.1st_Vout_1.t16 GNDA 0.346937f
C2325 bgr_0.1st_Vout_1.t33 GNDA 0.352846f
C2326 bgr_0.1st_Vout_1.t26 GNDA 0.346937f
C2327 bgr_0.1st_Vout_1.t22 GNDA 0.346937f
C2328 bgr_0.1st_Vout_1.t17 GNDA 0.352846f
C2329 bgr_0.1st_Vout_1.t24 GNDA 0.346937f
C2330 bgr_0.1st_Vout_1.t28 GNDA 0.352846f
C2331 bgr_0.1st_Vout_1.t23 GNDA 0.346937f
C2332 bgr_0.1st_Vout_1.t13 GNDA 0.346937f
C2333 bgr_0.1st_Vout_1.t18 GNDA 0.346937f
C2334 bgr_0.1st_Vout_1.t36 GNDA 0.346937f
C2335 bgr_0.1st_Vout_1.t30 GNDA 0.022665f
C2336 bgr_0.1st_Vout_1.n4 GNDA 0.021864f
C2337 bgr_0.1st_Vout_1.t14 GNDA 0.013213f
C2338 bgr_0.1st_Vout_1.t31 GNDA 0.013213f
C2339 bgr_0.1st_Vout_1.n5 GNDA 0.029393f
C2340 bgr_0.1st_Vout_1.t7 GNDA 0.018268f
C2341 bgr_0.1st_Vout_1.n6 GNDA 0.012529f
C2342 bgr_0.1st_Vout_1.n7 GNDA 0.189508f
C2343 bgr_0.1st_Vout_1.n8 GNDA 0.011336f
C2344 bgr_0.1st_Vout_1.n9 GNDA 0.020958f
C2345 bgr_0.1st_Vout_1.t19 GNDA 0.013213f
C2346 bgr_0.1st_Vout_1.t27 GNDA 0.013213f
C2347 bgr_0.1st_Vout_1.n10 GNDA 0.029393f
C2348 bgr_0.1st_Vout_1.n11 GNDA 0.021864f
C2349 bgr_0.1st_Vout_1.t15 GNDA 0.020738f
C2350 VDDA.t87 GNDA 0.019992f
C2351 VDDA.t232 GNDA 0.019992f
C2352 VDDA.n0 GNDA 0.082674f
C2353 VDDA.t137 GNDA 0.019992f
C2354 VDDA.t78 GNDA 0.019992f
C2355 VDDA.n1 GNDA 0.082357f
C2356 VDDA.n2 GNDA 0.114184f
C2357 VDDA.t140 GNDA 0.019992f
C2358 VDDA.t79 GNDA 0.019992f
C2359 VDDA.n3 GNDA 0.082357f
C2360 VDDA.n4 GNDA 0.059583f
C2361 VDDA.t139 GNDA 0.019992f
C2362 VDDA.t95 GNDA 0.019992f
C2363 VDDA.n5 GNDA 0.082357f
C2364 VDDA.n6 GNDA 0.059583f
C2365 VDDA.t138 GNDA 0.019992f
C2366 VDDA.t44 GNDA 0.019992f
C2367 VDDA.n7 GNDA 0.082357f
C2368 VDDA.n8 GNDA 0.059583f
C2369 VDDA.t241 GNDA 0.019992f
C2370 VDDA.t43 GNDA 0.019992f
C2371 VDDA.n9 GNDA 0.082357f
C2372 VDDA.n10 GNDA 0.172082f
C2373 VDDA.t143 GNDA 0.039983f
C2374 VDDA.t82 GNDA 0.039983f
C2375 VDDA.n11 GNDA 0.160407f
C2376 VDDA.n12 GNDA 0.081491f
C2377 VDDA.t375 GNDA 0.03983f
C2378 VDDA.n13 GNDA 0.053933f
C2379 VDDA.n14 GNDA 0.076127f
C2380 VDDA.t382 GNDA 0.044236f
C2381 VDDA.t380 GNDA 0.019371f
C2382 VDDA.n15 GNDA 0.07017f
C2383 VDDA.n16 GNDA 0.041309f
C2384 VDDA.t369 GNDA 0.044236f
C2385 VDDA.t367 GNDA 0.019371f
C2386 VDDA.n17 GNDA 0.07017f
C2387 VDDA.n18 GNDA 0.041309f
C2388 VDDA.n19 GNDA 0.043981f
C2389 VDDA.n20 GNDA 0.076127f
C2390 VDDA.n21 GNDA 0.220076f
C2391 VDDA.t368 GNDA 0.272557f
C2392 VDDA.t226 GNDA 0.1576f
C2393 VDDA.t147 GNDA 0.1576f
C2394 VDDA.t216 GNDA 0.1576f
C2395 VDDA.t46 GNDA 0.1576f
C2396 VDDA.t225 GNDA 0.1182f
C2397 VDDA.n22 GNDA 0.0788f
C2398 VDDA.t161 GNDA 0.1182f
C2399 VDDA.t75 GNDA 0.1576f
C2400 VDDA.t217 GNDA 0.1576f
C2401 VDDA.t183 GNDA 0.1576f
C2402 VDDA.t144 GNDA 0.1576f
C2403 VDDA.t381 GNDA 0.272557f
C2404 VDDA.n23 GNDA 0.220076f
C2405 VDDA.n24 GNDA 0.053933f
C2406 VDDA.n25 GNDA 0.102059f
C2407 VDDA.n26 GNDA 0.069846f
C2408 VDDA.n27 GNDA 0.103601f
C2409 VDDA.n28 GNDA 0.103601f
C2410 VDDA.n29 GNDA 0.102926f
C2411 VDDA.t363 GNDA 0.03983f
C2412 VDDA.t219 GNDA 0.039983f
C2413 VDDA.t215 GNDA 0.039983f
C2414 VDDA.n30 GNDA 0.160407f
C2415 VDDA.n31 GNDA 0.081491f
C2416 VDDA.t133 GNDA 0.039983f
C2417 VDDA.t160 GNDA 0.039983f
C2418 VDDA.n32 GNDA 0.160407f
C2419 VDDA.n33 GNDA 0.081491f
C2420 VDDA.t157 GNDA 0.039983f
C2421 VDDA.t52 GNDA 0.039983f
C2422 VDDA.n34 GNDA 0.160407f
C2423 VDDA.n35 GNDA 0.081491f
C2424 VDDA.t121 GNDA 0.039983f
C2425 VDDA.t236 GNDA 0.039983f
C2426 VDDA.n36 GNDA 0.160407f
C2427 VDDA.n37 GNDA 0.171241f
C2428 VDDA.n38 GNDA 0.12929f
C2429 VDDA.t361 GNDA 0.048328f
C2430 VDDA.n39 GNDA 0.092466f
C2431 VDDA.n40 GNDA 0.054021f
C2432 VDDA.n41 GNDA 0.080828f
C2433 VDDA.n42 GNDA 0.355777f
C2434 VDDA.t362 GNDA 0.549534f
C2435 VDDA.t120 GNDA 0.304205f
C2436 VDDA.t235 GNDA 0.304205f
C2437 VDDA.t156 GNDA 0.304205f
C2438 VDDA.t51 GNDA 0.304205f
C2439 VDDA.t132 GNDA 0.228154f
C2440 VDDA.n43 GNDA 0.152103f
C2441 VDDA.t159 GNDA 0.228154f
C2442 VDDA.t218 GNDA 0.304205f
C2443 VDDA.t214 GNDA 0.304205f
C2444 VDDA.t142 GNDA 0.304205f
C2445 VDDA.t81 GNDA 0.304205f
C2446 VDDA.t374 GNDA 0.549534f
C2447 VDDA.n44 GNDA 0.355777f
C2448 VDDA.n45 GNDA 0.080828f
C2449 VDDA.n46 GNDA 0.054021f
C2450 VDDA.t373 GNDA 0.048328f
C2451 VDDA.n47 GNDA 0.092466f
C2452 VDDA.n48 GNDA 0.128957f
C2453 VDDA.n49 GNDA 0.096748f
C2454 VDDA.t222 GNDA 0.019992f
C2455 VDDA.t227 GNDA 0.019992f
C2456 VDDA.n50 GNDA 0.082674f
C2457 VDDA.t458 GNDA 0.019992f
C2458 VDDA.t459 GNDA 0.019992f
C2459 VDDA.n51 GNDA 0.082357f
C2460 VDDA.n52 GNDA 0.114184f
C2461 VDDA.t158 GNDA 0.019992f
C2462 VDDA.t184 GNDA 0.019992f
C2463 VDDA.n53 GNDA 0.082357f
C2464 VDDA.n54 GNDA 0.059583f
C2465 VDDA.t468 GNDA 0.019992f
C2466 VDDA.t98 GNDA 0.019992f
C2467 VDDA.n55 GNDA 0.082357f
C2468 VDDA.n56 GNDA 0.059583f
C2469 VDDA.t146 GNDA 0.019992f
C2470 VDDA.t164 GNDA 0.019992f
C2471 VDDA.n57 GNDA 0.082357f
C2472 VDDA.n58 GNDA 0.059583f
C2473 VDDA.t145 GNDA 0.019992f
C2474 VDDA.t30 GNDA 0.019992f
C2475 VDDA.n59 GNDA 0.082357f
C2476 VDDA.n60 GNDA 0.205853f
C2477 VDDA.n61 GNDA 0.190255f
C2478 VDDA.t419 GNDA 0.023323f
C2479 VDDA.t119 GNDA 0.023323f
C2480 VDDA.n62 GNDA 0.081114f
C2481 VDDA.t3 GNDA 0.023323f
C2482 VDDA.t42 GNDA 0.023323f
C2483 VDDA.n63 GNDA 0.080827f
C2484 VDDA.n64 GNDA 0.152593f
C2485 VDDA.t60 GNDA 0.023323f
C2486 VDDA.t54 GNDA 0.023323f
C2487 VDDA.n65 GNDA 0.081114f
C2488 VDDA.t224 GNDA 0.023323f
C2489 VDDA.t248 GNDA 0.023323f
C2490 VDDA.n66 GNDA 0.080827f
C2491 VDDA.n67 GNDA 0.152593f
C2492 VDDA.n68 GNDA 0.021324f
C2493 VDDA.n69 GNDA 0.066399f
C2494 VDDA.n70 GNDA 0.09029f
C2495 VDDA.t385 GNDA 0.11506f
C2496 VDDA.t383 GNDA 0.040614f
C2497 VDDA.n71 GNDA 0.075062f
C2498 VDDA.n72 GNDA 0.048388f
C2499 VDDA.t303 GNDA 0.11506f
C2500 VDDA.t301 GNDA 0.040614f
C2501 VDDA.n73 GNDA 0.075062f
C2502 VDDA.n74 GNDA 0.048388f
C2503 VDDA.n75 GNDA 0.04798f
C2504 VDDA.n76 GNDA 0.09029f
C2505 VDDA.n77 GNDA 0.269081f
C2506 VDDA.t302 GNDA 0.401642f
C2507 VDDA.t418 GNDA 0.231902f
C2508 VDDA.t118 GNDA 0.231902f
C2509 VDDA.t2 GNDA 0.231902f
C2510 VDDA.t41 GNDA 0.231902f
C2511 VDDA.t69 GNDA 0.173927f
C2512 VDDA.n78 GNDA 0.115951f
C2513 VDDA.t181 GNDA 0.173927f
C2514 VDDA.t223 GNDA 0.231902f
C2515 VDDA.t247 GNDA 0.231902f
C2516 VDDA.t59 GNDA 0.231902f
C2517 VDDA.t53 GNDA 0.231902f
C2518 VDDA.t384 GNDA 0.401642f
C2519 VDDA.n79 GNDA 0.269081f
C2520 VDDA.n80 GNDA 0.066399f
C2521 VDDA.n81 GNDA 0.092956f
C2522 VDDA.t70 GNDA 0.023323f
C2523 VDDA.t182 GNDA 0.023323f
C2524 VDDA.n82 GNDA 0.076044f
C2525 VDDA.n83 GNDA 0.051902f
C2526 VDDA.n84 GNDA 0.028951f
C2527 VDDA.n85 GNDA 0.116321f
C2528 VDDA.t243 GNDA 0.023323f
C2529 VDDA.t195 GNDA 0.023323f
C2530 VDDA.n86 GNDA 0.081114f
C2531 VDDA.t127 GNDA 0.023323f
C2532 VDDA.t432 GNDA 0.023323f
C2533 VDDA.n87 GNDA 0.080827f
C2534 VDDA.n88 GNDA 0.152593f
C2535 VDDA.t197 GNDA 0.023323f
C2536 VDDA.t9 GNDA 0.023323f
C2537 VDDA.n89 GNDA 0.081114f
C2538 VDDA.t421 GNDA 0.023323f
C2539 VDDA.t166 GNDA 0.023323f
C2540 VDDA.n90 GNDA 0.080827f
C2541 VDDA.n91 GNDA 0.152593f
C2542 VDDA.n92 GNDA 0.021324f
C2543 VDDA.n93 GNDA 0.066399f
C2544 VDDA.n94 GNDA 0.09029f
C2545 VDDA.t318 GNDA 0.11506f
C2546 VDDA.t316 GNDA 0.040614f
C2547 VDDA.n95 GNDA 0.075062f
C2548 VDDA.n96 GNDA 0.048388f
C2549 VDDA.t406 GNDA 0.11506f
C2550 VDDA.t404 GNDA 0.040614f
C2551 VDDA.n97 GNDA 0.075062f
C2552 VDDA.n98 GNDA 0.048388f
C2553 VDDA.n99 GNDA 0.04798f
C2554 VDDA.n100 GNDA 0.09029f
C2555 VDDA.n101 GNDA 0.269081f
C2556 VDDA.t405 GNDA 0.401642f
C2557 VDDA.t242 GNDA 0.231902f
C2558 VDDA.t194 GNDA 0.231902f
C2559 VDDA.t126 GNDA 0.231902f
C2560 VDDA.t431 GNDA 0.231902f
C2561 VDDA.t55 GNDA 0.173927f
C2562 VDDA.n102 GNDA 0.115951f
C2563 VDDA.t429 GNDA 0.173927f
C2564 VDDA.t420 GNDA 0.231902f
C2565 VDDA.t165 GNDA 0.231902f
C2566 VDDA.t196 GNDA 0.231902f
C2567 VDDA.t8 GNDA 0.231902f
C2568 VDDA.t317 GNDA 0.401642f
C2569 VDDA.n103 GNDA 0.269081f
C2570 VDDA.n104 GNDA 0.066399f
C2571 VDDA.n105 GNDA 0.092956f
C2572 VDDA.t56 GNDA 0.023323f
C2573 VDDA.t430 GNDA 0.023323f
C2574 VDDA.n106 GNDA 0.076044f
C2575 VDDA.n107 GNDA 0.051902f
C2576 VDDA.n108 GNDA 0.028951f
C2577 VDDA.n109 GNDA 0.114322f
C2578 VDDA.t170 GNDA 0.039983f
C2579 VDDA.t136 GNDA 0.039983f
C2580 VDDA.n110 GNDA 0.160407f
C2581 VDDA.n111 GNDA 0.081491f
C2582 VDDA.t345 GNDA 0.03983f
C2583 VDDA.n112 GNDA 0.080828f
C2584 VDDA.n113 GNDA 0.053933f
C2585 VDDA.n114 GNDA 0.076127f
C2586 VDDA.t372 GNDA 0.044236f
C2587 VDDA.t370 GNDA 0.019371f
C2588 VDDA.n115 GNDA 0.07017f
C2589 VDDA.n116 GNDA 0.041309f
C2590 VDDA.t348 GNDA 0.044236f
C2591 VDDA.t346 GNDA 0.019371f
C2592 VDDA.n117 GNDA 0.07017f
C2593 VDDA.n118 GNDA 0.041309f
C2594 VDDA.n119 GNDA 0.043981f
C2595 VDDA.n120 GNDA 0.076127f
C2596 VDDA.n121 GNDA 0.220076f
C2597 VDDA.t347 GNDA 0.272557f
C2598 VDDA.t153 GNDA 0.1576f
C2599 VDDA.t141 GNDA 0.1576f
C2600 VDDA.t80 GNDA 0.1576f
C2601 VDDA.t90 GNDA 0.1576f
C2602 VDDA.t45 GNDA 0.1182f
C2603 VDDA.n122 GNDA 0.0788f
C2604 VDDA.t13 GNDA 0.1182f
C2605 VDDA.t86 GNDA 0.1576f
C2606 VDDA.t83 GNDA 0.1576f
C2607 VDDA.t152 GNDA 0.1576f
C2608 VDDA.t134 GNDA 0.1576f
C2609 VDDA.t371 GNDA 0.272557f
C2610 VDDA.n123 GNDA 0.220076f
C2611 VDDA.n124 GNDA 0.053933f
C2612 VDDA.n125 GNDA 0.102059f
C2613 VDDA.t366 GNDA 0.03983f
C2614 VDDA.t77 GNDA 0.039983f
C2615 VDDA.t92 GNDA 0.039983f
C2616 VDDA.n126 GNDA 0.160407f
C2617 VDDA.n127 GNDA 0.081491f
C2618 VDDA.t19 GNDA 0.039983f
C2619 VDDA.t15 GNDA 0.039983f
C2620 VDDA.n128 GNDA 0.160407f
C2621 VDDA.n129 GNDA 0.081491f
C2622 VDDA.t94 GNDA 0.039983f
C2623 VDDA.t85 GNDA 0.039983f
C2624 VDDA.n130 GNDA 0.160407f
C2625 VDDA.n131 GNDA 0.081491f
C2626 VDDA.t168 GNDA 0.039983f
C2627 VDDA.t17 GNDA 0.039983f
C2628 VDDA.n132 GNDA 0.160407f
C2629 VDDA.n133 GNDA 0.171241f
C2630 VDDA.n134 GNDA 0.12929f
C2631 VDDA.t364 GNDA 0.048328f
C2632 VDDA.n135 GNDA 0.092466f
C2633 VDDA.n136 GNDA 0.054021f
C2634 VDDA.n137 GNDA 0.355777f
C2635 VDDA.n138 GNDA 0.355777f
C2636 VDDA.t344 GNDA 0.549534f
C2637 VDDA.t169 GNDA 0.304205f
C2638 VDDA.t135 GNDA 0.304205f
C2639 VDDA.t76 GNDA 0.304205f
C2640 VDDA.t91 GNDA 0.304205f
C2641 VDDA.t18 GNDA 0.228154f
C2642 VDDA.n139 GNDA 0.080828f
C2643 VDDA.n140 GNDA 0.103601f
C2644 VDDA.n141 GNDA 0.103601f
C2645 VDDA.t365 GNDA 0.549534f
C2646 VDDA.t16 GNDA 0.304205f
C2647 VDDA.t167 GNDA 0.304205f
C2648 VDDA.t84 GNDA 0.304205f
C2649 VDDA.t93 GNDA 0.304205f
C2650 VDDA.t14 GNDA 0.228154f
C2651 VDDA.n142 GNDA 0.152103f
C2652 VDDA.n143 GNDA 0.102926f
C2653 VDDA.n144 GNDA 0.069846f
C2654 VDDA.n145 GNDA 0.054021f
C2655 VDDA.t343 GNDA 0.048328f
C2656 VDDA.n146 GNDA 0.092466f
C2657 VDDA.n147 GNDA 0.128957f
C2658 VDDA.n148 GNDA 0.098747f
C2659 VDDA.n149 GNDA 0.05531f
C2660 VDDA.n150 GNDA 0.187042f
C2661 VDDA.n151 GNDA 0.064556f
C2662 VDDA.n152 GNDA 0.172346f
C2663 VDDA.t312 GNDA 0.012556f
C2664 VDDA.n153 GNDA 0.026718f
C2665 VDDA.t415 GNDA 0.012556f
C2666 VDDA.n154 GNDA 0.026718f
C2667 VDDA.n155 GNDA 0.038793f
C2668 VDDA.n156 GNDA 0.065203f
C2669 VDDA.n157 GNDA 0.173768f
C2670 VDDA.t357 GNDA 0.012556f
C2671 VDDA.n158 GNDA 0.026718f
C2672 VDDA.t339 GNDA 0.012556f
C2673 VDDA.n159 GNDA 0.026718f
C2674 VDDA.n160 GNDA 0.036151f
C2675 VDDA.n161 GNDA 0.044876f
C2676 VDDA.n162 GNDA 0.173768f
C2677 VDDA.t338 GNDA 0.169043f
C2678 VDDA.t7 GNDA 0.104456f
C2679 VDDA.t61 GNDA 0.104456f
C2680 VDDA.t426 GNDA 0.104456f
C2681 VDDA.t31 GNDA 0.104456f
C2682 VDDA.t199 GNDA 0.078342f
C2683 VDDA.t356 GNDA 0.169043f
C2684 VDDA.t228 GNDA 0.104456f
C2685 VDDA.t35 GNDA 0.104456f
C2686 VDDA.t32 GNDA 0.104456f
C2687 VDDA.t441 GNDA 0.104456f
C2688 VDDA.t427 GNDA 0.078342f
C2689 VDDA.n163 GNDA 0.06585f
C2690 VDDA.n164 GNDA 0.052228f
C2691 VDDA.n165 GNDA 0.06585f
C2692 VDDA.n166 GNDA 0.043981f
C2693 VDDA.n167 GNDA 0.035585f
C2694 VDDA.n168 GNDA 0.08274f
C2695 VDDA.n169 GNDA 0.08274f
C2696 VDDA.n170 GNDA 0.172346f
C2697 VDDA.t414 GNDA 0.165634f
C2698 VDDA.t6 GNDA 0.102623f
C2699 VDDA.t209 GNDA 0.102623f
C2700 VDDA.t428 GNDA 0.102623f
C2701 VDDA.t12 GNDA 0.102623f
C2702 VDDA.t36 GNDA 0.076968f
C2703 VDDA.t311 GNDA 0.165634f
C2704 VDDA.t229 GNDA 0.102623f
C2705 VDDA.t68 GNDA 0.102623f
C2706 VDDA.t198 GNDA 0.102623f
C2707 VDDA.t200 GNDA 0.102623f
C2708 VDDA.t117 GNDA 0.076968f
C2709 VDDA.n171 GNDA 0.06585f
C2710 VDDA.n172 GNDA 0.051312f
C2711 VDDA.n173 GNDA 0.06585f
C2712 VDDA.n174 GNDA 0.043772f
C2713 VDDA.n175 GNDA 0.035585f
C2714 VDDA.n176 GNDA 0.068889f
C2715 VDDA.n177 GNDA 0.092151f
C2716 VDDA.n179 GNDA 0.051023f
C2717 VDDA.n180 GNDA 0.080633f
C2718 VDDA.n181 GNDA 0.102305f
C2719 VDDA.n182 GNDA 0.102305f
C2720 VDDA.n183 GNDA 0.102305f
C2721 VDDA.n185 GNDA 0.051023f
C2722 VDDA.n187 GNDA 0.051023f
C2723 VDDA.n189 GNDA 0.051023f
C2724 VDDA.n191 GNDA 0.051023f
C2725 VDDA.n193 GNDA 0.051023f
C2726 VDDA.n195 GNDA 0.051023f
C2727 VDDA.n197 GNDA 0.051023f
C2728 VDDA.n199 GNDA 0.051023f
C2729 VDDA.n201 GNDA 0.083495f
C2730 VDDA.t397 GNDA 0.012141f
C2731 VDDA.n202 GNDA 0.018027f
C2732 VDDA.n203 GNDA 0.01595f
C2733 VDDA.n204 GNDA 0.054477f
C2734 VDDA.n205 GNDA 0.063299f
C2735 VDDA.n206 GNDA 0.209192f
C2736 VDDA.t396 GNDA 0.165634f
C2737 VDDA.t179 GNDA 0.102623f
C2738 VDDA.t115 GNDA 0.102623f
C2739 VDDA.t237 GNDA 0.102623f
C2740 VDDA.t49 GNDA 0.102623f
C2741 VDDA.t20 GNDA 0.102623f
C2742 VDDA.t64 GNDA 0.102623f
C2743 VDDA.t88 GNDA 0.102623f
C2744 VDDA.t33 GNDA 0.102623f
C2745 VDDA.t442 GNDA 0.102623f
C2746 VDDA.t62 GNDA 0.076968f
C2747 VDDA.n207 GNDA 0.051312f
C2748 VDDA.t191 GNDA 0.076968f
C2749 VDDA.t239 GNDA 0.102623f
C2750 VDDA.t39 GNDA 0.102623f
C2751 VDDA.t187 GNDA 0.102623f
C2752 VDDA.t439 GNDA 0.102623f
C2753 VDDA.t230 GNDA 0.102623f
C2754 VDDA.t4 GNDA 0.102623f
C2755 VDDA.t189 GNDA 0.102623f
C2756 VDDA.t37 GNDA 0.102623f
C2757 VDDA.t66 GNDA 0.102623f
C2758 VDDA.t390 GNDA 0.165634f
C2759 VDDA.n208 GNDA 0.209192f
C2760 VDDA.n209 GNDA 0.063299f
C2761 VDDA.n210 GNDA 0.054477f
C2762 VDDA.n211 GNDA 0.01595f
C2763 VDDA.t391 GNDA 0.012141f
C2764 VDDA.n212 GNDA 0.017587f
C2765 VDDA.n213 GNDA 0.087494f
C2766 VDDA.n214 GNDA 0.081361f
C2767 VDDA.n216 GNDA 0.065024f
C2768 VDDA.n217 GNDA 0.011995f
C2769 VDDA.n218 GNDA 0.035432f
C2770 VDDA.n219 GNDA 0.035432f
C2771 VDDA.n220 GNDA 0.036128f
C2772 VDDA.n221 GNDA 0.090779f
C2773 VDDA.n222 GNDA 0.011995f
C2774 VDDA.n223 GNDA 0.05328f
C2775 VDDA.n224 GNDA 0.05328f
C2776 VDDA.n225 GNDA 0.05328f
C2777 VDDA.t100 GNDA 0.021324f
C2778 VDDA.n226 GNDA 0.073999f
C2779 VDDA.t309 GNDA 0.097402f
C2780 VDDA.n227 GNDA 0.0483f
C2781 VDDA.n228 GNDA 0.046368f
C2782 VDDA.t307 GNDA 0.03701f
C2783 VDDA.n229 GNDA 0.039183f
C2784 VDDA.n230 GNDA 0.02933f
C2785 VDDA.n231 GNDA 0.045573f
C2786 VDDA.n232 GNDA 0.298773f
C2787 VDDA.t308 GNDA 0.284007f
C2788 VDDA.n233 GNDA 0.092461f
C2789 VDDA.n234 GNDA 0.023115f
C2790 VDDA.t99 GNDA 0.129445f
C2791 VDDA.t329 GNDA 0.307122f
C2792 VDDA.n235 GNDA 0.301866f
C2793 VDDA.n236 GNDA 0.04729f
C2794 VDDA.n237 GNDA 0.030325f
C2795 VDDA.t328 GNDA 0.037675f
C2796 VDDA.n238 GNDA 0.039183f
C2797 VDDA.t330 GNDA 0.076078f
C2798 VDDA.n239 GNDA 0.052212f
C2799 VDDA.n240 GNDA 0.103903f
C2800 VDDA.n241 GNDA 0.069119f
C2801 VDDA.t351 GNDA 0.015576f
C2802 VDDA.n242 GNDA 0.016922f
C2803 VDDA.t349 GNDA 0.013068f
C2804 VDDA.n243 GNDA 0.016545f
C2805 VDDA.n244 GNDA 0.021303f
C2806 VDDA.n245 GNDA 0.029894f
C2807 VDDA.n246 GNDA 0.159455f
C2808 VDDA.t350 GNDA 0.176608f
C2809 VDDA.t422 GNDA 0.119949f
C2810 VDDA.t377 GNDA 0.176608f
C2811 VDDA.n247 GNDA 0.159455f
C2812 VDDA.n248 GNDA 0.029894f
C2813 VDDA.n249 GNDA 0.021303f
C2814 VDDA.t376 GNDA 0.013068f
C2815 VDDA.n250 GNDA 0.016545f
C2816 VDDA.t379 GNDA 0.015576f
C2817 VDDA.n251 GNDA 0.01889f
C2818 VDDA.n252 GNDA 0.064825f
C2819 VDDA.n253 GNDA 0.190377f
C2820 VDDA.n254 GNDA 4.39288f
C2821 VDDA.t470 GNDA 0.736718f
C2822 VDDA.t471 GNDA 0.7852f
C2823 VDDA.t469 GNDA 0.7852f
C2824 VDDA.t472 GNDA 0.752935f
C2825 VDDA.n255 GNDA 0.526323f
C2826 VDDA.n256 GNDA 0.255528f
C2827 VDDA.n257 GNDA 0.327604f
C2828 VDDA.n258 GNDA 2.34056f
C2829 VDDA.n259 GNDA 0.021324f
C2830 VDDA.n260 GNDA 0.01614f
C2831 VDDA.n261 GNDA 0.01614f
C2832 VDDA.n262 GNDA 0.047167f
C2833 VDDA.n263 GNDA 0.021324f
C2834 VDDA.t336 GNDA 0.025033f
C2835 VDDA.t334 GNDA 0.016495f
C2836 VDDA.n264 GNDA 0.039271f
C2837 VDDA.n265 GNDA 0.055877f
C2838 VDDA.n266 GNDA 0.105047f
C2839 VDDA.n267 GNDA 0.105047f
C2840 VDDA.t315 GNDA 0.025033f
C2841 VDDA.t313 GNDA 0.016495f
C2842 VDDA.n268 GNDA 0.039271f
C2843 VDDA.n269 GNDA 0.079966f
C2844 VDDA.n270 GNDA 0.055877f
C2845 VDDA.n271 GNDA 0.021324f
C2846 VDDA.n272 GNDA 0.01614f
C2847 VDDA.n273 GNDA 0.016875f
C2848 VDDA.n274 GNDA 0.016761f
C2849 VDDA.n275 GNDA 0.130295f
C2850 VDDA.n276 GNDA 0.016761f
C2851 VDDA.n277 GNDA 0.06787f
C2852 VDDA.n278 GNDA 0.016761f
C2853 VDDA.n279 GNDA 0.06787f
C2854 VDDA.n280 GNDA 0.01614f
C2855 VDDA.n281 GNDA 0.065549f
C2856 VDDA.n282 GNDA 0.105047f
C2857 VDDA.t342 GNDA 0.025033f
C2858 VDDA.t340 GNDA 0.016495f
C2859 VDDA.n283 GNDA 0.039271f
C2860 VDDA.n284 GNDA 0.055877f
C2861 VDDA.t412 GNDA 0.025033f
C2862 VDDA.t410 GNDA 0.016495f
C2863 VDDA.n285 GNDA 0.039271f
C2864 VDDA.n286 GNDA 0.055877f
C2865 VDDA.n287 GNDA 0.079966f
C2866 VDDA.n288 GNDA 0.105047f
C2867 VDDA.n289 GNDA 0.228403f
C2868 VDDA.t411 GNDA 0.208322f
C2869 VDDA.t47 GNDA 0.131944f
C2870 VDDA.t0 GNDA 0.131944f
C2871 VDDA.t435 GNDA 0.131944f
C2872 VDDA.t437 GNDA 0.131944f
C2873 VDDA.t460 GNDA 0.131944f
C2874 VDDA.t205 GNDA 0.131944f
C2875 VDDA.t433 GNDA 0.131944f
C2876 VDDA.t220 GNDA 0.131944f
C2877 VDDA.t73 GNDA 0.098958f
C2878 VDDA.n290 GNDA 0.065972f
C2879 VDDA.t128 GNDA 0.098958f
C2880 VDDA.t444 GNDA 0.131944f
C2881 VDDA.t416 GNDA 0.131944f
C2882 VDDA.t233 GNDA 0.131944f
C2883 VDDA.t22 GNDA 0.131944f
C2884 VDDA.t185 GNDA 0.131944f
C2885 VDDA.t124 GNDA 0.131944f
C2886 VDDA.t171 GNDA 0.131944f
C2887 VDDA.t207 GNDA 0.131944f
C2888 VDDA.t341 GNDA 0.208322f
C2889 VDDA.n291 GNDA 0.228403f
C2890 VDDA.n292 GNDA 0.065549f
C2891 VDDA.n293 GNDA 0.111665f
C2892 VDDA.n294 GNDA 0.047167f
C2893 VDDA.n295 GNDA 0.021324f
C2894 VDDA.n296 GNDA 0.016761f
C2895 VDDA.n297 GNDA 0.06787f
C2896 VDDA.n298 GNDA 0.016761f
C2897 VDDA.n299 GNDA 0.06787f
C2898 VDDA.n300 GNDA 0.016761f
C2899 VDDA.n301 GNDA 0.06787f
C2900 VDDA.n302 GNDA 0.016761f
C2901 VDDA.n303 GNDA 0.097191f
C2902 VDDA.n304 GNDA 0.021324f
C2903 VDDA.n305 GNDA 0.01614f
C2904 VDDA.n306 GNDA 0.01614f
C2905 VDDA.n307 GNDA 0.047167f
C2906 VDDA.n308 GNDA 0.021324f
C2907 VDDA.n309 GNDA 0.01614f
C2908 VDDA.n310 GNDA 0.021324f
C2909 VDDA.n311 GNDA 0.01614f
C2910 VDDA.n312 GNDA 0.047167f
C2911 VDDA.n313 GNDA 0.021324f
C2912 VDDA.n314 GNDA 0.021324f
C2913 VDDA.n315 GNDA 0.047167f
C2914 VDDA.n316 GNDA 0.021324f
C2915 VDDA.n317 GNDA 0.021324f
C2916 VDDA.n318 GNDA 0.01614f
C2917 VDDA.n319 GNDA 0.047167f
C2918 VDDA.n320 GNDA 0.021324f
C2919 VDDA.n321 GNDA 0.021324f
C2920 VDDA.n322 GNDA 0.047167f
C2921 VDDA.n323 GNDA 0.021324f
C2922 VDDA.n324 GNDA 0.01614f
C2923 VDDA.n325 GNDA 0.047167f
C2924 VDDA.n326 GNDA 0.021324f
C2925 VDDA.n327 GNDA 0.050645f
C2926 VDDA.n328 GNDA 0.047167f
C2927 VDDA.n329 GNDA 0.034816f
C2928 VDDA.n330 GNDA 0.033255f
C2929 VDDA.n331 GNDA 0.228403f
C2930 VDDA.t314 GNDA 0.208322f
C2931 VDDA.t245 GNDA 0.131944f
C2932 VDDA.t148 GNDA 0.131944f
C2933 VDDA.t111 GNDA 0.131944f
C2934 VDDA.t122 GNDA 0.131944f
C2935 VDDA.t105 GNDA 0.131944f
C2936 VDDA.t71 GNDA 0.131944f
C2937 VDDA.t424 GNDA 0.131944f
C2938 VDDA.t162 GNDA 0.131944f
C2939 VDDA.t113 GNDA 0.098958f
C2940 VDDA.n332 GNDA 0.065972f
C2941 VDDA.t203 GNDA 0.098958f
C2942 VDDA.t464 GNDA 0.131944f
C2943 VDDA.t10 GNDA 0.131944f
C2944 VDDA.t154 GNDA 0.131944f
C2945 VDDA.t96 GNDA 0.131944f
C2946 VDDA.t150 GNDA 0.131944f
C2947 VDDA.t456 GNDA 0.131944f
C2948 VDDA.t57 GNDA 0.131944f
C2949 VDDA.t28 GNDA 0.131944f
C2950 VDDA.t335 GNDA 0.208322f
C2951 VDDA.n333 GNDA 0.228403f
C2952 VDDA.n334 GNDA 0.033255f
C2953 VDDA.n335 GNDA 0.034816f
C2954 VDDA.n336 GNDA 0.047167f
C2955 VDDA.n337 GNDA 0.064558f
C2956 VDDA.n338 GNDA 0.195999f
C2957 VDDA.t276 GNDA 0.019992f
C2958 VDDA.t274 GNDA 0.019992f
C2959 VDDA.n339 GNDA 0.066046f
C2960 VDDA.n340 GNDA 0.085224f
C2961 VDDA.t394 GNDA 0.061266f
C2962 VDDA.n341 GNDA 0.107955f
C2963 VDDA.n342 GNDA 0.147162f
C2964 VDDA.n343 GNDA 0.147162f
C2965 VDDA.n344 GNDA 0.146486f
C2966 VDDA.t333 GNDA 0.061266f
C2967 VDDA.t331 GNDA 0.095328f
C2968 VDDA.t360 GNDA 0.025033f
C2969 VDDA.t358 GNDA 0.012633f
C2970 VDDA.n345 GNDA 0.039468f
C2971 VDDA.n346 GNDA 0.022758f
C2972 VDDA.n347 GNDA 0.040446f
C2973 VDDA.t400 GNDA 0.025033f
C2974 VDDA.t398 GNDA 0.012633f
C2975 VDDA.n348 GNDA 0.039468f
C2976 VDDA.n349 GNDA 0.040446f
C2977 VDDA.n350 GNDA 0.040446f
C2978 VDDA.n351 GNDA 0.033187f
C2979 VDDA.n352 GNDA 0.159475f
C2980 VDDA.t359 GNDA 0.200244f
C2981 VDDA.t244 GNDA 0.090712f
C2982 VDDA.n353 GNDA 0.060475f
C2983 VDDA.t193 GNDA 0.090712f
C2984 VDDA.t399 GNDA 0.203197f
C2985 VDDA.n354 GNDA 0.167517f
C2986 VDDA.n355 GNDA 0.033187f
C2987 VDDA.n356 GNDA 0.022758f
C2988 VDDA.n357 GNDA 0.031972f
C2989 VDDA.t295 GNDA 0.019992f
C2990 VDDA.t256 GNDA 0.019992f
C2991 VDDA.n358 GNDA 0.066046f
C2992 VDDA.n359 GNDA 0.085224f
C2993 VDDA.t267 GNDA 0.019992f
C2994 VDDA.t286 GNDA 0.019992f
C2995 VDDA.n360 GNDA 0.066046f
C2996 VDDA.n361 GNDA 0.085224f
C2997 VDDA.t251 GNDA 0.019992f
C2998 VDDA.t270 GNDA 0.019992f
C2999 VDDA.n362 GNDA 0.066046f
C3000 VDDA.n363 GNDA 0.085224f
C3001 VDDA.t284 GNDA 0.019992f
C3002 VDDA.t292 GNDA 0.019992f
C3003 VDDA.n364 GNDA 0.066046f
C3004 VDDA.n365 GNDA 0.085224f
C3005 VDDA.t265 GNDA 0.019992f
C3006 VDDA.t261 GNDA 0.019992f
C3007 VDDA.n366 GNDA 0.066046f
C3008 VDDA.n367 GNDA 0.085224f
C3009 VDDA.t290 GNDA 0.019992f
C3010 VDDA.t300 GNDA 0.019992f
C3011 VDDA.n368 GNDA 0.066046f
C3012 VDDA.n369 GNDA 0.085224f
C3013 VDDA.t258 GNDA 0.019992f
C3014 VDDA.t279 GNDA 0.019992f
C3015 VDDA.n370 GNDA 0.066046f
C3016 VDDA.n371 GNDA 0.085224f
C3017 VDDA.n372 GNDA 0.094096f
C3018 VDDA.n373 GNDA 0.113771f
C3019 VDDA.n374 GNDA 0.076687f
C3020 VDDA.n375 GNDA 0.093629f
C3021 VDDA.n376 GNDA 0.344978f
C3022 VDDA.t332 GNDA 0.445136f
C3023 VDDA.t257 GNDA 0.320865f
C3024 VDDA.t278 GNDA 0.320865f
C3025 VDDA.t289 GNDA 0.320865f
C3026 VDDA.t299 GNDA 0.320865f
C3027 VDDA.t264 GNDA 0.320865f
C3028 VDDA.t260 GNDA 0.320865f
C3029 VDDA.t283 GNDA 0.320865f
C3030 VDDA.t291 GNDA 0.240649f
C3031 VDDA.n377 GNDA 0.160432f
C3032 VDDA.t250 GNDA 0.240649f
C3033 VDDA.t269 GNDA 0.320865f
C3034 VDDA.t266 GNDA 0.320865f
C3035 VDDA.t285 GNDA 0.320865f
C3036 VDDA.t294 GNDA 0.320865f
C3037 VDDA.t255 GNDA 0.320865f
C3038 VDDA.t275 GNDA 0.320865f
C3039 VDDA.t273 GNDA 0.320865f
C3040 VDDA.t393 GNDA 0.445136f
C3041 VDDA.n378 GNDA 0.344978f
C3042 VDDA.n379 GNDA 0.093629f
C3043 VDDA.n380 GNDA 0.076687f
C3044 VDDA.t392 GNDA 0.095328f
C3045 VDDA.n381 GNDA 0.113771f
C3046 VDDA.n382 GNDA 0.052225f
C3047 VDDA.n383 GNDA 0.016094f
C3048 VDDA.t324 GNDA 0.025219f
C3049 VDDA.t322 GNDA 0.012306f
C3050 VDDA.n384 GNDA 0.037776f
C3051 VDDA.n385 GNDA 0.022653f
C3052 VDDA.n386 GNDA 0.040446f
C3053 VDDA.t321 GNDA 0.025219f
C3054 VDDA.t319 GNDA 0.012306f
C3055 VDDA.n387 GNDA 0.037776f
C3056 VDDA.n388 GNDA 0.040446f
C3057 VDDA.n389 GNDA 0.040446f
C3058 VDDA.n390 GNDA 0.033187f
C3059 VDDA.n391 GNDA 0.159475f
C3060 VDDA.t323 GNDA 0.200244f
C3061 VDDA.t26 GNDA 0.090712f
C3062 VDDA.n392 GNDA 0.060475f
C3063 VDDA.t107 GNDA 0.090712f
C3064 VDDA.t320 GNDA 0.200244f
C3065 VDDA.n393 GNDA 0.159475f
C3066 VDDA.n394 GNDA 0.033187f
C3067 VDDA.n395 GNDA 0.022653f
C3068 VDDA.n396 GNDA 0.023799f
C3069 VDDA.n397 GNDA 0.044547f
C3070 VDDA.n398 GNDA 0.093855f
C3071 VDDA.n399 GNDA 0.162977f
C3072 VDDA.n400 GNDA 0.016623f
C3073 VDDA.n401 GNDA 0.058679f
C3074 VDDA.t327 GNDA 0.026299f
C3075 VDDA.n402 GNDA 0.021991f
C3076 VDDA.n403 GNDA 0.047599f
C3077 VDDA.n404 GNDA 0.047599f
C3078 VDDA.n405 GNDA 0.047599f
C3079 VDDA.t388 GNDA 0.026299f
C3080 VDDA.t386 GNDA 0.013124f
C3081 VDDA.n406 GNDA 0.016592f
C3082 VDDA.n407 GNDA 0.058709f
C3083 VDDA.t403 GNDA 0.025097f
C3084 VDDA.n408 GNDA 0.043981f
C3085 VDDA.n409 GNDA 0.069292f
C3086 VDDA.n410 GNDA 0.069292f
C3087 VDDA.n411 GNDA 0.069292f
C3088 VDDA.t409 GNDA 0.025097f
C3089 VDDA.t407 GNDA 0.013124f
C3090 VDDA.n412 GNDA 0.01663f
C3091 VDDA.n413 GNDA 0.058672f
C3092 VDDA.t354 GNDA 0.02631f
C3093 VDDA.n414 GNDA 0.021991f
C3094 VDDA.n415 GNDA 0.047599f
C3095 VDDA.n416 GNDA 0.047599f
C3096 VDDA.n417 GNDA 0.047599f
C3097 VDDA.t306 GNDA 0.02631f
C3098 VDDA.t304 GNDA 0.013124f
C3099 VDDA.n418 GNDA 0.01663f
C3100 VDDA.n419 GNDA 0.080302f
C3101 VDDA.n420 GNDA 0.045058f
C3102 VDDA.n421 GNDA 0.02689f
C3103 VDDA.n422 GNDA 0.036941f
C3104 VDDA.n423 GNDA 0.168291f
C3105 VDDA.t305 GNDA 0.203766f
C3106 VDDA.t201 GNDA 0.122782f
C3107 VDDA.t24 GNDA 0.092086f
C3108 VDDA.n424 GNDA 0.061391f
C3109 VDDA.t130 GNDA 0.092086f
C3110 VDDA.t452 GNDA 0.122782f
C3111 VDDA.t353 GNDA 0.203766f
C3112 VDDA.n425 GNDA 0.168291f
C3113 VDDA.n426 GNDA 0.036941f
C3114 VDDA.n427 GNDA 0.02689f
C3115 VDDA.t352 GNDA 0.01354f
C3116 VDDA.n428 GNDA 0.044593f
C3117 VDDA.n429 GNDA 0.040505f
C3118 VDDA.n430 GNDA 0.016592f
C3119 VDDA.n431 GNDA 0.058709f
C3120 VDDA.n432 GNDA 0.016592f
C3121 VDDA.n433 GNDA 0.058709f
C3122 VDDA.n434 GNDA 0.016592f
C3123 VDDA.n435 GNDA 0.058709f
C3124 VDDA.n436 GNDA 0.016592f
C3125 VDDA.n437 GNDA 0.058709f
C3126 VDDA.n438 GNDA 0.040505f
C3127 VDDA.n439 GNDA 0.045389f
C3128 VDDA.n440 GNDA 0.04155f
C3129 VDDA.n441 GNDA 0.051785f
C3130 VDDA.n442 GNDA 0.19798f
C3131 VDDA.t408 GNDA 0.203766f
C3132 VDDA.t109 GNDA 0.122782f
C3133 VDDA.t175 GNDA 0.122782f
C3134 VDDA.t448 GNDA 0.122782f
C3135 VDDA.t454 GNDA 0.122782f
C3136 VDDA.t101 GNDA 0.122782f
C3137 VDDA.t446 GNDA 0.092086f
C3138 VDDA.n443 GNDA 0.061391f
C3139 VDDA.t177 GNDA 0.092086f
C3140 VDDA.t450 GNDA 0.122782f
C3141 VDDA.t462 GNDA 0.122782f
C3142 VDDA.t212 GNDA 0.122782f
C3143 VDDA.t402 GNDA 0.203766f
C3144 VDDA.n444 GNDA 0.18318f
C3145 VDDA.n445 GNDA 0.044385f
C3146 VDDA.n446 GNDA 0.03422f
C3147 VDDA.t401 GNDA 0.013124f
C3148 VDDA.n447 GNDA 0.045389f
C3149 VDDA.n448 GNDA 0.047835f
C3150 VDDA.n449 GNDA 0.016623f
C3151 VDDA.n450 GNDA 0.058679f
C3152 VDDA.n451 GNDA 0.047835f
C3153 VDDA.n452 GNDA 0.044187f
C3154 VDDA.n453 GNDA 0.02689f
C3155 VDDA.n454 GNDA 0.036431f
C3156 VDDA.n455 GNDA 0.166472f
C3157 VDDA.t387 GNDA 0.200244f
C3158 VDDA.t173 GNDA 0.120949f
C3159 VDDA.t103 GNDA 0.082465f
C3160 VDDA.n456 GNDA 0.030237f
C3161 VDDA.n457 GNDA 0.038484f
C3162 VDDA.t466 GNDA 0.090712f
C3163 VDDA.t210 GNDA 0.120949f
C3164 VDDA.t326 GNDA 0.200244f
C3165 VDDA.n458 GNDA 0.167492f
C3166 VDDA.n459 GNDA 0.03745f
C3167 VDDA.n460 GNDA 0.02689f
C3168 VDDA.t325 GNDA 0.013124f
C3169 VDDA.n461 GNDA 0.044187f
C3170 VDDA.n462 GNDA 0.088133f
C3171 VDDA.n463 GNDA 0.132296f
C3172 VDDA.t288 GNDA 0.37251f
C3173 VDDA.t296 GNDA 0.37386f
C3174 VDDA.t268 GNDA 0.37251f
C3175 VDDA.t252 GNDA 0.37386f
C3176 VDDA.t277 GNDA 0.37251f
C3177 VDDA.t281 GNDA 0.37386f
C3178 VDDA.t253 GNDA 0.37251f
C3179 VDDA.t293 GNDA 0.37386f
C3180 VDDA.t282 GNDA 0.37251f
C3181 VDDA.t298 GNDA 0.37386f
C3182 VDDA.t271 GNDA 0.37251f
C3183 VDDA.t254 GNDA 0.37386f
C3184 VDDA.t249 GNDA 0.37251f
C3185 VDDA.t263 GNDA 0.37386f
C3186 VDDA.t287 GNDA 0.37251f
C3187 VDDA.t272 GNDA 0.37386f
C3188 VDDA.n464 GNDA 0.249694f
C3189 VDDA.t280 GNDA 0.198844f
C3190 VDDA.n465 GNDA 0.270923f
C3191 VDDA.t262 GNDA 0.198844f
C3192 VDDA.n466 GNDA 0.270923f
C3193 VDDA.t297 GNDA 0.198844f
C3194 VDDA.n467 GNDA 0.270923f
C3195 VDDA.t259 GNDA 0.296715f
C3196 VDDA.n468 GNDA 0.258551f
C3197 VDDA.n469 GNDA 0.803512f
C3198 bgr_0.Vin-.n0 GNDA 0.073641f
C3199 bgr_0.Vin-.n1 GNDA 0.338979f
C3200 bgr_0.Vin-.n2 GNDA 0.510703f
C3201 bgr_0.Vin-.t2 GNDA 0.276239f
C3202 bgr_0.Vin-.n3 GNDA 0.331333f
C3203 bgr_0.Vin-.n4 GNDA 0.073776f
C3204 bgr_0.Vin-.n5 GNDA 0.12627f
C3205 bgr_0.Vin-.n6 GNDA 0.074468f
C3206 bgr_0.Vin-.n7 GNDA 0.998981f
C3207 bgr_0.Vin-.t4 GNDA 0.028614f
C3208 bgr_0.Vin-.t5 GNDA 0.028614f
C3209 bgr_0.Vin-.n8 GNDA 0.099613f
C3210 bgr_0.Vin-.t7 GNDA 0.028614f
C3211 bgr_0.Vin-.t6 GNDA 0.028614f
C3212 bgr_0.Vin-.n9 GNDA 0.095121f
C3213 bgr_0.Vin-.n10 GNDA 0.408067f
C3214 bgr_0.Vin-.t0 GNDA 0.098662f
C3215 bgr_0.Vin-.n11 GNDA 0.025702f
C3216 bgr_0.Vin-.n12 GNDA 0.469862f
C3217 bgr_0.Vin-.n13 GNDA 0.222852f
C3218 bgr_0.Vin-.t10 GNDA 0.023594f
C3219 bgr_0.Vin-.n14 GNDA 0.027673f
C3220 bgr_0.Vin-.n15 GNDA 0.022653f
C3221 bgr_0.Vin-.n16 GNDA 0.022653f
C3222 bgr_0.Vin-.n17 GNDA 0.040466f
C3223 bgr_0.Vin-.n18 GNDA 0.524007f
C3224 bgr_0.Vin-.n19 GNDA 0.461299f
C3225 bgr_0.Vin-.n20 GNDA 0.166915f
C3226 bgr_0.Vin-.n21 GNDA 0.074625f
C3227 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter GNDA 0.043026f
C3228 bgr_0.V_TOP.t31 GNDA 0.115045f
C3229 bgr_0.V_TOP.t44 GNDA 0.115045f
C3230 bgr_0.V_TOP.t18 GNDA 0.115045f
C3231 bgr_0.V_TOP.t26 GNDA 0.115045f
C3232 bgr_0.V_TOP.t37 GNDA 0.115045f
C3233 bgr_0.V_TOP.t35 GNDA 0.115045f
C3234 bgr_0.V_TOP.t48 GNDA 0.115045f
C3235 bgr_0.V_TOP.t20 GNDA 0.115045f
C3236 bgr_0.V_TOP.t27 GNDA 0.115045f
C3237 bgr_0.V_TOP.t41 GNDA 0.115045f
C3238 bgr_0.V_TOP.t38 GNDA 0.115045f
C3239 bgr_0.V_TOP.t14 GNDA 0.115045f
C3240 bgr_0.V_TOP.t23 GNDA 0.115045f
C3241 bgr_0.V_TOP.t29 GNDA 0.115045f
C3242 bgr_0.V_TOP.t43 GNDA 0.150392f
C3243 bgr_0.V_TOP.n0 GNDA 0.084081f
C3244 bgr_0.V_TOP.n1 GNDA 0.061357f
C3245 bgr_0.V_TOP.n2 GNDA 0.061357f
C3246 bgr_0.V_TOP.n3 GNDA 0.061357f
C3247 bgr_0.V_TOP.n4 GNDA 0.061357f
C3248 bgr_0.V_TOP.n5 GNDA 0.057217f
C3249 bgr_0.V_TOP.t2 GNDA 0.147947f
C3250 bgr_0.V_TOP.t4 GNDA 0.155772f
C3251 bgr_0.V_TOP.t1 GNDA 0.010957f
C3252 bgr_0.V_TOP.t0 GNDA 0.010957f
C3253 bgr_0.V_TOP.n6 GNDA 0.027281f
C3254 bgr_0.V_TOP.n7 GNDA 0.726844f
C3255 bgr_0.V_TOP.t5 GNDA 0.010957f
C3256 bgr_0.V_TOP.t12 GNDA 0.010957f
C3257 bgr_0.V_TOP.n8 GNDA 0.026425f
C3258 bgr_0.V_TOP.t9 GNDA 0.010957f
C3259 bgr_0.V_TOP.t10 GNDA 0.010957f
C3260 bgr_0.V_TOP.n9 GNDA 0.027465f
C3261 bgr_0.V_TOP.t3 GNDA 0.010957f
C3262 bgr_0.V_TOP.t13 GNDA 0.010957f
C3263 bgr_0.V_TOP.n10 GNDA 0.027281f
C3264 bgr_0.V_TOP.n11 GNDA 0.252824f
C3265 bgr_0.V_TOP.n12 GNDA 0.153577f
C3266 bgr_0.V_TOP.n13 GNDA 0.087653f
C3267 bgr_0.V_TOP.t11 GNDA 0.010957f
C3268 bgr_0.V_TOP.t8 GNDA 0.010957f
C3269 bgr_0.V_TOP.n14 GNDA 0.027281f
C3270 bgr_0.V_TOP.n15 GNDA 0.151313f
C3271 bgr_0.V_TOP.t6 GNDA 0.010957f
C3272 bgr_0.V_TOP.t7 GNDA 0.010957f
C3273 bgr_0.V_TOP.n16 GNDA 0.027281f
C3274 bgr_0.V_TOP.n17 GNDA 0.149874f
C3275 bgr_0.V_TOP.n18 GNDA 0.329448f
C3276 bgr_0.V_TOP.n19 GNDA 0.023183f
C3277 bgr_0.V_TOP.n20 GNDA 0.057217f
C3278 bgr_0.V_TOP.n21 GNDA 0.061357f
C3279 bgr_0.V_TOP.n22 GNDA 0.061357f
C3280 bgr_0.V_TOP.n23 GNDA 0.061357f
C3281 bgr_0.V_TOP.n24 GNDA 0.061357f
C3282 bgr_0.V_TOP.n25 GNDA 0.061357f
C3283 bgr_0.V_TOP.n26 GNDA 0.061357f
C3284 bgr_0.V_TOP.n27 GNDA 0.057217f
C3285 bgr_0.V_TOP.t32 GNDA 0.132572f
C3286 bgr_0.V_TOP.t49 GNDA 0.445732f
C3287 bgr_0.V_TOP.t39 GNDA 0.438267f
C3288 bgr_0.V_TOP.n28 GNDA 0.293844f
C3289 bgr_0.V_TOP.t28 GNDA 0.438267f
C3290 bgr_0.V_TOP.t25 GNDA 0.445732f
C3291 bgr_0.V_TOP.t33 GNDA 0.438267f
C3292 bgr_0.V_TOP.n29 GNDA 0.293844f
C3293 bgr_0.V_TOP.n30 GNDA 0.273917f
C3294 bgr_0.V_TOP.t21 GNDA 0.445732f
C3295 bgr_0.V_TOP.t15 GNDA 0.438267f
C3296 bgr_0.V_TOP.n31 GNDA 0.293844f
C3297 bgr_0.V_TOP.t40 GNDA 0.438267f
C3298 bgr_0.V_TOP.t34 GNDA 0.445732f
C3299 bgr_0.V_TOP.t45 GNDA 0.438267f
C3300 bgr_0.V_TOP.n32 GNDA 0.293844f
C3301 bgr_0.V_TOP.n33 GNDA 0.356092f
C3302 bgr_0.V_TOP.t30 GNDA 0.445732f
C3303 bgr_0.V_TOP.t22 GNDA 0.438267f
C3304 bgr_0.V_TOP.n34 GNDA 0.293844f
C3305 bgr_0.V_TOP.t16 GNDA 0.438267f
C3306 bgr_0.V_TOP.t46 GNDA 0.445732f
C3307 bgr_0.V_TOP.t19 GNDA 0.438267f
C3308 bgr_0.V_TOP.n35 GNDA 0.293844f
C3309 bgr_0.V_TOP.n36 GNDA 0.356092f
C3310 bgr_0.V_TOP.t24 GNDA 0.445732f
C3311 bgr_0.V_TOP.t17 GNDA 0.438267f
C3312 bgr_0.V_TOP.n37 GNDA 0.293844f
C3313 bgr_0.V_TOP.t42 GNDA 0.438267f
C3314 bgr_0.V_TOP.n38 GNDA 0.273917f
C3315 bgr_0.V_TOP.t47 GNDA 0.438267f
C3316 bgr_0.V_TOP.n39 GNDA 0.191742f
C3317 bgr_0.V_TOP.t36 GNDA 0.438267f
C3318 bgr_0.V_TOP.n40 GNDA 0.893239f
.ends

