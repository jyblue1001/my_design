* NGSPICE file created from opamp_cell.ext - technology: sky130A

**.subckt opamp_cell
X0 w_8020_4460# p_bias p_bias w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=1.25 ps=6 w=2.5 l=0.5
X1 w_8020_4460# n_left n_left w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X2 v_common_n a_7320_4730# n_left a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X3 w_8020_4460# p_bias v_common_p w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X4 w_8020_4460# p_bias p_bias w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X5 n_left a_7320_4730# v_common_n a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X6 a_7760_2448# p_right a_8190_3850# sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X7 a_9460_3850# n_right w_8020_4460# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X8 a_9460_3850# a_10686_2448# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X9 v_common_p a_7320_4730# p_left w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X10 a_9460_3850# p_right a_8190_3850# a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X11 w_8020_4460# n_right a_9460_3850# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X12 p_right p_left a_8190_3850# a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X13 p_left a_7320_4730# v_common_p w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X14 a_8190_3850# p_right a_9460_3850# a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X15 a_8190_3850# p_left p_left a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X16 w_8020_4460# p_bias v_common_p w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X17 v_common_n n_bias a_8190_3850# a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X18 n_bias n_bias a_8190_3850# a_8190_3850# sky130_fd_pr__nfet_01v8 ad=1.25 pd=6 as=0.625 ps=3 w=2.5 l=0.5
X19 v_common_p p_bias w_8020_4460# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X20 n_right a_10686_2448# a_8190_3850# sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X21 p_bias p_bias w_8020_4460# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X22 a_9460_3850# n_right w_8020_4460# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X23 a_9460_3850# a_7760_2448# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X24 v_common_p a_7750_4400# p_right w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X25 a_9460_3850# p_right a_8190_3850# a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X26 n_left n_left w_8020_4460# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X27 w_8020_4460# n_right a_9460_3850# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X28 p_left p_left a_8190_3850# a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X29 v_common_n a_7750_4400# n_right a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X30 p_right a_7750_4400# v_common_p w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X31 w_8020_4460# n_left n_right w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X32 a_8190_3850# p_right a_9460_3850# a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X33 a_8190_3850# p_left p_right a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X34 n_right a_7750_4400# v_common_n a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X35 p_bias n_bias a_8190_3850# sky130_fd_pr__res_xhigh_po_2p85 l=0.51
X36 v_common_p p_bias w_8020_4460# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X37 a_8190_3850# n_bias n_bias a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=1.25 ps=6 w=2.5 l=0.5
X38 p_bias p_bias w_8020_4460# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0.625 ps=3 w=2.5 l=0.5
X39 n_right n_left w_8020_4460# w_8020_4460# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X40 a_8190_3850# n_bias v_common_n a_8190_3850# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
**.ends

