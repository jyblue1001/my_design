magic
tech sky130A
timestamp 1738218882
<< nwell >>
rect -1545 620 385 1205
<< pwell >>
rect -865 520 -850 525
rect -1370 390 -55 515
rect -805 385 -55 390
rect -805 380 -440 385
rect -805 320 -640 380
rect -525 345 -440 380
rect -525 330 -475 345
rect -455 330 -440 345
rect -525 320 -440 330
rect -495 315 -455 320
rect -445 290 -405 315
<< nmos >>
rect -1300 410 -1285 510
rect -1155 410 -1140 510
rect -1010 410 -995 510
rect -865 410 -850 510
rect -720 410 -705 510
rect -575 410 -560 510
rect -430 410 -415 510
rect -285 410 -270 510
rect -140 410 -125 510
rect -1455 155 -1395 255
rect -1345 155 -1285 255
rect -1235 155 -1175 255
rect -1125 155 -1065 255
rect -795 155 -735 255
rect -685 155 -625 255
rect -575 155 -515 255
rect -465 155 -405 255
rect -75 155 -15 255
rect 35 155 95 255
rect 145 155 205 255
rect 255 155 315 255
<< pmos >>
rect -1475 1085 -1415 1185
rect -1365 1085 -1305 1185
rect -1255 1085 -1195 1185
rect -1145 1085 -1085 1185
rect -1035 1085 -975 1185
rect -925 1085 -865 1185
rect -815 1085 -755 1185
rect -705 1085 -645 1185
rect -515 1085 -455 1185
rect -405 1085 -345 1185
rect -295 1085 -235 1185
rect -185 1085 -125 1185
rect -75 1085 -15 1185
rect 35 1085 95 1185
rect 145 1085 205 1185
rect 255 1085 315 1185
rect -1300 640 -1285 840
rect -1155 640 -1140 840
rect -1010 640 -995 840
rect -865 640 -850 840
rect -720 640 -705 840
rect -575 640 -560 840
rect -430 640 -415 840
rect -285 640 -270 840
rect -140 640 -125 840
<< ndiff >>
rect -1350 495 -1300 510
rect -1350 425 -1335 495
rect -1315 425 -1300 495
rect -1350 410 -1300 425
rect -1285 495 -1235 510
rect -1285 425 -1270 495
rect -1250 425 -1235 495
rect -1285 410 -1235 425
rect -1205 495 -1155 510
rect -1205 425 -1190 495
rect -1170 425 -1155 495
rect -1205 410 -1155 425
rect -1140 495 -1090 510
rect -1140 425 -1125 495
rect -1105 425 -1090 495
rect -1140 410 -1090 425
rect -1060 495 -1010 510
rect -1060 425 -1045 495
rect -1025 425 -1010 495
rect -1060 410 -1010 425
rect -995 495 -945 510
rect -995 425 -980 495
rect -960 425 -945 495
rect -995 410 -945 425
rect -915 495 -865 510
rect -915 425 -900 495
rect -880 425 -865 495
rect -915 410 -865 425
rect -850 495 -800 510
rect -850 425 -835 495
rect -815 425 -800 495
rect -850 410 -800 425
rect -770 495 -720 510
rect -770 425 -755 495
rect -735 425 -720 495
rect -770 410 -720 425
rect -705 495 -655 510
rect -705 425 -690 495
rect -670 425 -655 495
rect -705 410 -655 425
rect -625 495 -575 510
rect -625 425 -610 495
rect -590 425 -575 495
rect -625 410 -575 425
rect -560 495 -510 510
rect -560 425 -545 495
rect -525 425 -510 495
rect -560 410 -510 425
rect -480 495 -430 510
rect -480 425 -465 495
rect -445 425 -430 495
rect -480 410 -430 425
rect -415 495 -365 510
rect -415 425 -400 495
rect -380 425 -365 495
rect -415 410 -365 425
rect -335 495 -285 510
rect -335 425 -320 495
rect -300 425 -285 495
rect -335 410 -285 425
rect -270 495 -220 510
rect -270 425 -255 495
rect -235 425 -220 495
rect -270 410 -220 425
rect -190 495 -140 510
rect -190 425 -175 495
rect -155 425 -140 495
rect -190 410 -140 425
rect -125 495 -75 510
rect -125 425 -110 495
rect -90 425 -75 495
rect -125 410 -75 425
rect -1505 240 -1455 255
rect -1505 170 -1490 240
rect -1470 170 -1455 240
rect -1505 155 -1455 170
rect -1395 240 -1345 255
rect -1395 170 -1380 240
rect -1360 170 -1345 240
rect -1395 155 -1345 170
rect -1285 240 -1235 255
rect -1285 170 -1270 240
rect -1250 170 -1235 240
rect -1285 155 -1235 170
rect -1175 240 -1125 255
rect -1175 170 -1160 240
rect -1140 170 -1125 240
rect -1175 155 -1125 170
rect -1065 240 -1015 255
rect -1065 170 -1050 240
rect -1030 170 -1015 240
rect -1065 155 -1015 170
rect -845 240 -795 255
rect -845 170 -830 240
rect -810 170 -795 240
rect -845 155 -795 170
rect -735 240 -685 255
rect -735 170 -720 240
rect -700 170 -685 240
rect -735 155 -685 170
rect -625 240 -575 255
rect -625 170 -610 240
rect -590 170 -575 240
rect -625 155 -575 170
rect -515 240 -465 255
rect -515 170 -500 240
rect -480 170 -465 240
rect -515 155 -465 170
rect -405 240 -355 255
rect -405 170 -390 240
rect -370 170 -355 240
rect -405 155 -355 170
rect -125 240 -75 255
rect -125 170 -110 240
rect -90 170 -75 240
rect -125 155 -75 170
rect -15 240 35 255
rect -15 170 0 240
rect 20 170 35 240
rect -15 155 35 170
rect 95 240 145 255
rect 95 170 110 240
rect 130 170 145 240
rect 95 155 145 170
rect 205 240 255 255
rect 205 170 220 240
rect 240 170 255 240
rect 205 155 255 170
rect 315 240 365 255
rect 315 170 330 240
rect 350 170 365 240
rect 315 155 365 170
<< pdiff >>
rect -1525 1170 -1475 1185
rect -1525 1100 -1510 1170
rect -1490 1100 -1475 1170
rect -1525 1085 -1475 1100
rect -1415 1170 -1365 1185
rect -1415 1100 -1400 1170
rect -1380 1100 -1365 1170
rect -1415 1085 -1365 1100
rect -1305 1170 -1255 1185
rect -1305 1100 -1290 1170
rect -1270 1100 -1255 1170
rect -1305 1085 -1255 1100
rect -1195 1170 -1145 1185
rect -1195 1100 -1180 1170
rect -1160 1100 -1145 1170
rect -1195 1085 -1145 1100
rect -1085 1170 -1035 1185
rect -1085 1100 -1070 1170
rect -1050 1100 -1035 1170
rect -1085 1085 -1035 1100
rect -975 1170 -925 1185
rect -975 1100 -960 1170
rect -940 1100 -925 1170
rect -975 1085 -925 1100
rect -865 1170 -815 1185
rect -865 1100 -850 1170
rect -830 1100 -815 1170
rect -865 1085 -815 1100
rect -755 1170 -705 1185
rect -755 1100 -740 1170
rect -720 1100 -705 1170
rect -755 1085 -705 1100
rect -645 1170 -595 1185
rect -645 1100 -630 1170
rect -610 1100 -595 1170
rect -645 1085 -595 1100
rect -565 1170 -515 1185
rect -565 1100 -550 1170
rect -530 1100 -515 1170
rect -565 1085 -515 1100
rect -455 1170 -405 1185
rect -455 1100 -440 1170
rect -420 1100 -405 1170
rect -455 1085 -405 1100
rect -345 1170 -295 1185
rect -345 1100 -330 1170
rect -310 1100 -295 1170
rect -345 1085 -295 1100
rect -235 1170 -185 1185
rect -235 1100 -220 1170
rect -200 1100 -185 1170
rect -235 1085 -185 1100
rect -125 1170 -75 1185
rect -125 1100 -110 1170
rect -90 1100 -75 1170
rect -125 1085 -75 1100
rect -15 1170 35 1185
rect -15 1100 0 1170
rect 20 1100 35 1170
rect -15 1085 35 1100
rect 95 1170 145 1185
rect 95 1100 110 1170
rect 130 1100 145 1170
rect 95 1085 145 1100
rect 205 1170 255 1185
rect 205 1100 220 1170
rect 240 1100 255 1170
rect 205 1085 255 1100
rect 315 1170 365 1185
rect 315 1100 330 1170
rect 350 1100 365 1170
rect 315 1085 365 1100
rect -1350 825 -1300 840
rect -1350 655 -1335 825
rect -1315 655 -1300 825
rect -1350 640 -1300 655
rect -1285 825 -1235 840
rect -1285 655 -1270 825
rect -1250 655 -1235 825
rect -1285 640 -1235 655
rect -1205 825 -1155 840
rect -1205 655 -1190 825
rect -1170 655 -1155 825
rect -1205 640 -1155 655
rect -1140 825 -1090 840
rect -1140 655 -1125 825
rect -1105 655 -1090 825
rect -1140 640 -1090 655
rect -1060 825 -1010 840
rect -1060 655 -1045 825
rect -1025 655 -1010 825
rect -1060 640 -1010 655
rect -995 825 -945 840
rect -995 655 -980 825
rect -960 655 -945 825
rect -995 640 -945 655
rect -915 825 -865 840
rect -915 655 -900 825
rect -880 655 -865 825
rect -915 640 -865 655
rect -850 825 -800 840
rect -850 655 -835 825
rect -815 655 -800 825
rect -850 640 -800 655
rect -770 825 -720 840
rect -770 655 -755 825
rect -735 655 -720 825
rect -770 640 -720 655
rect -705 825 -655 840
rect -705 655 -690 825
rect -670 655 -655 825
rect -705 640 -655 655
rect -625 825 -575 840
rect -625 655 -610 825
rect -590 655 -575 825
rect -625 640 -575 655
rect -560 825 -510 840
rect -560 655 -545 825
rect -525 655 -510 825
rect -560 640 -510 655
rect -480 825 -430 840
rect -480 655 -465 825
rect -445 655 -430 825
rect -480 640 -430 655
rect -415 825 -365 840
rect -415 655 -400 825
rect -380 655 -365 825
rect -415 640 -365 655
rect -335 825 -285 840
rect -335 655 -320 825
rect -300 655 -285 825
rect -335 640 -285 655
rect -270 825 -220 840
rect -270 655 -255 825
rect -235 655 -220 825
rect -270 640 -220 655
rect -190 825 -140 840
rect -190 655 -175 825
rect -155 655 -140 825
rect -190 640 -140 655
rect -125 825 -75 840
rect -125 655 -110 825
rect -90 655 -75 825
rect -125 640 -75 655
<< ndiffc >>
rect -1335 425 -1315 495
rect -1270 425 -1250 495
rect -1190 425 -1170 495
rect -1125 425 -1105 495
rect -1045 425 -1025 495
rect -980 425 -960 495
rect -900 425 -880 495
rect -835 425 -815 495
rect -755 425 -735 495
rect -690 425 -670 495
rect -610 425 -590 495
rect -545 425 -525 495
rect -465 425 -445 495
rect -400 425 -380 495
rect -320 425 -300 495
rect -255 425 -235 495
rect -175 425 -155 495
rect -110 425 -90 495
rect -1490 170 -1470 240
rect -1380 170 -1360 240
rect -1270 170 -1250 240
rect -1160 170 -1140 240
rect -1050 170 -1030 240
rect -830 170 -810 240
rect -720 170 -700 240
rect -610 170 -590 240
rect -500 170 -480 240
rect -390 170 -370 240
rect -110 170 -90 240
rect 0 170 20 240
rect 110 170 130 240
rect 220 170 240 240
rect 330 170 350 240
<< pdiffc >>
rect -1510 1100 -1490 1170
rect -1400 1100 -1380 1170
rect -1290 1100 -1270 1170
rect -1180 1100 -1160 1170
rect -1070 1100 -1050 1170
rect -960 1100 -940 1170
rect -850 1100 -830 1170
rect -740 1100 -720 1170
rect -630 1100 -610 1170
rect -550 1100 -530 1170
rect -440 1100 -420 1170
rect -330 1100 -310 1170
rect -220 1100 -200 1170
rect -110 1100 -90 1170
rect 0 1100 20 1170
rect 110 1100 130 1170
rect 220 1100 240 1170
rect 330 1100 350 1170
rect -1335 655 -1315 825
rect -1270 655 -1250 825
rect -1190 655 -1170 825
rect -1125 655 -1105 825
rect -1045 655 -1025 825
rect -980 655 -960 825
rect -900 655 -880 825
rect -835 655 -815 825
rect -755 655 -735 825
rect -690 655 -670 825
rect -610 655 -590 825
rect -545 655 -525 825
rect -465 655 -445 825
rect -400 655 -380 825
rect -320 655 -300 825
rect -255 655 -235 825
rect -175 655 -155 825
rect -110 655 -90 825
<< psubdiff >>
rect -45 495 5 510
rect -45 425 -30 495
rect -10 425 5 495
rect -45 410 5 425
<< nsubdiff >>
rect -45 825 5 840
rect -45 655 -30 825
rect -10 655 5 825
rect -45 640 5 655
<< psubdiffcont >>
rect -30 425 -10 495
<< nsubdiffcont >>
rect -30 655 -10 825
<< poly >>
rect -1475 1185 -1415 1200
rect -1365 1185 -1305 1200
rect -1255 1185 -1195 1200
rect -1145 1185 -1085 1200
rect -1035 1185 -975 1200
rect -925 1185 -865 1200
rect -815 1185 -755 1200
rect -705 1185 -645 1200
rect -515 1185 -455 1200
rect -405 1185 -345 1200
rect -295 1185 -235 1200
rect -185 1185 -125 1200
rect -75 1185 -15 1200
rect 35 1185 95 1200
rect 145 1185 205 1200
rect 255 1185 315 1200
rect -1475 1075 -1415 1085
rect -1365 1075 -1305 1085
rect -1255 1075 -1195 1085
rect -1145 1075 -1085 1085
rect -1035 1075 -975 1085
rect -925 1075 -865 1085
rect -815 1075 -755 1085
rect -705 1075 -645 1085
rect -1475 1055 -645 1075
rect -515 1075 -455 1085
rect -405 1075 -345 1085
rect -295 1075 -235 1085
rect -185 1075 -125 1085
rect -75 1075 -15 1085
rect 35 1075 95 1085
rect 145 1075 205 1085
rect 255 1075 315 1085
rect -515 1060 315 1075
rect 340 1060 380 1070
rect -895 970 -880 1055
rect -910 960 -870 970
rect -910 940 -900 960
rect -880 940 -870 960
rect -910 930 -870 940
rect -1010 890 -125 905
rect 50 895 65 1060
rect 340 1040 350 1060
rect 370 1040 380 1060
rect 340 1030 380 1040
rect -1300 840 -1285 855
rect -1155 840 -1140 855
rect -1010 840 -995 890
rect -865 840 -850 855
rect -720 840 -705 855
rect -575 840 -560 855
rect -430 840 -415 855
rect -285 840 -270 855
rect -140 840 -125 890
rect 35 885 75 895
rect 35 865 45 885
rect 65 865 75 885
rect 35 855 75 865
rect 340 665 355 1030
rect 340 650 1245 665
rect -1300 585 -1285 640
rect -1155 600 -1140 640
rect -1010 600 -995 640
rect -865 625 -850 640
rect -1665 570 -1285 585
rect -1300 510 -1285 570
rect -1180 590 -1140 600
rect -1180 570 -1170 590
rect -1150 570 -1140 590
rect -1180 560 -1140 570
rect -1035 590 -995 600
rect -1035 570 -1025 590
rect -1005 570 -995 590
rect -970 615 -850 625
rect -970 595 -960 615
rect -940 610 -850 615
rect -940 595 -930 610
rect -970 585 -930 595
rect -1035 560 -995 570
rect -1155 510 -1140 560
rect -1010 535 -995 560
rect -1010 520 -850 535
rect -1010 510 -995 520
rect -865 510 -850 520
rect -720 510 -705 640
rect -575 630 -560 640
rect -655 615 -560 630
rect -535 615 -495 625
rect -430 615 -415 640
rect -285 615 -270 640
rect -140 625 -125 640
rect -655 565 -640 615
rect -535 595 -525 615
rect -505 600 -160 615
rect -505 595 -495 600
rect -535 590 -495 595
rect -680 555 -640 565
rect -495 560 -455 565
rect -680 535 -670 555
rect -650 535 -640 555
rect -680 525 -640 535
rect -575 555 -455 560
rect -575 545 -485 555
rect -575 510 -560 545
rect -495 535 -485 545
rect -465 535 -455 555
rect -495 525 -455 535
rect -430 510 -415 600
rect -175 580 -160 600
rect -175 565 -125 580
rect -390 550 -350 560
rect -390 530 -380 550
rect -360 535 -350 550
rect -360 530 -270 535
rect -390 520 -270 530
rect -285 510 -270 520
rect -140 510 -125 565
rect 50 555 90 565
rect 50 535 60 555
rect 80 535 90 555
rect 50 525 90 535
rect -1300 395 -1285 410
rect -1155 395 -1140 410
rect -1010 395 -995 410
rect -865 395 -850 410
rect -720 370 -705 410
rect -575 395 -560 410
rect -1665 355 -705 370
rect -430 330 -415 410
rect -285 395 -270 410
rect -285 385 -230 395
rect -285 365 -260 385
rect -240 365 -230 385
rect -285 355 -230 365
rect -140 330 -125 410
rect -495 320 -455 330
rect -1500 300 -1460 310
rect -1500 280 -1490 300
rect -1470 290 -1460 300
rect -1280 300 -1240 310
rect -1280 290 -1270 300
rect -1470 280 -1270 290
rect -1250 290 -1240 300
rect -1060 300 -1020 310
rect -1060 290 -1050 300
rect -1250 280 -1050 290
rect -1030 290 -1020 300
rect -495 300 -485 320
rect -465 300 -455 320
rect -430 315 -125 330
rect -495 290 -455 300
rect -1030 280 -405 290
rect 75 280 90 525
rect 340 305 355 650
rect 340 295 380 305
rect -1500 265 -405 280
rect -1455 255 -1395 265
rect -1345 255 -1285 265
rect -1235 255 -1175 265
rect -1125 255 -1065 265
rect -795 255 -735 265
rect -685 255 -625 265
rect -575 255 -515 265
rect -465 255 -405 265
rect -75 265 315 280
rect 340 275 350 295
rect 370 275 380 295
rect 340 265 380 275
rect -75 255 -15 265
rect 35 255 95 265
rect 145 255 205 265
rect 255 255 315 265
rect -1455 140 -1395 155
rect -1345 140 -1285 155
rect -1235 140 -1175 155
rect -1125 140 -1065 155
rect -795 140 -735 155
rect -685 140 -625 155
rect -575 140 -515 155
rect -465 140 -405 155
rect -75 140 -15 155
rect 35 140 95 155
rect 145 140 205 155
rect 255 140 315 155
<< polycont >>
rect -900 940 -880 960
rect 350 1040 370 1060
rect 45 865 65 885
rect -1170 570 -1150 590
rect -1025 570 -1005 590
rect -960 595 -940 615
rect -525 595 -505 615
rect -670 535 -650 555
rect -485 535 -465 555
rect -380 530 -360 550
rect 60 535 80 555
rect -260 365 -240 385
rect -1490 280 -1470 300
rect -1270 280 -1250 300
rect -1050 280 -1030 300
rect -485 300 -465 320
rect 350 275 370 295
<< locali >>
rect -1510 1200 -610 1220
rect -1510 1180 -1490 1200
rect -1290 1180 -1270 1200
rect -1070 1180 -1050 1200
rect -850 1180 -830 1200
rect -630 1180 -610 1200
rect -550 1200 350 1220
rect -550 1180 -530 1200
rect -330 1180 -310 1200
rect -110 1180 -90 1200
rect 110 1180 130 1200
rect 330 1180 350 1200
rect -1520 1170 -1480 1180
rect -1520 1100 -1510 1170
rect -1490 1100 -1480 1170
rect -1520 1090 -1480 1100
rect -1410 1170 -1370 1180
rect -1410 1100 -1400 1170
rect -1380 1100 -1370 1170
rect -1410 1090 -1370 1100
rect -1300 1170 -1260 1180
rect -1300 1100 -1290 1170
rect -1270 1100 -1260 1170
rect -1300 1090 -1260 1100
rect -1190 1170 -1150 1180
rect -1190 1100 -1180 1170
rect -1160 1100 -1150 1170
rect -1190 1090 -1150 1100
rect -1080 1170 -1040 1180
rect -1080 1100 -1070 1170
rect -1050 1100 -1040 1170
rect -1080 1090 -1040 1100
rect -970 1170 -930 1180
rect -970 1100 -960 1170
rect -940 1100 -930 1170
rect -970 1090 -930 1100
rect -860 1170 -820 1180
rect -860 1100 -850 1170
rect -830 1100 -820 1170
rect -860 1090 -820 1100
rect -750 1170 -710 1180
rect -750 1100 -740 1170
rect -720 1100 -710 1170
rect -750 1090 -710 1100
rect -640 1170 -600 1180
rect -640 1100 -630 1170
rect -610 1100 -600 1170
rect -640 1090 -600 1100
rect -560 1170 -520 1180
rect -560 1100 -550 1170
rect -530 1100 -520 1170
rect -560 1090 -520 1100
rect -450 1170 -410 1180
rect -450 1100 -440 1170
rect -420 1100 -410 1170
rect -450 1090 -410 1100
rect -340 1170 -300 1180
rect -340 1100 -330 1170
rect -310 1100 -300 1170
rect -340 1090 -300 1100
rect -230 1170 -190 1180
rect -230 1100 -220 1170
rect -200 1100 -190 1170
rect -230 1090 -190 1100
rect -120 1170 -80 1180
rect -120 1100 -110 1170
rect -90 1100 -80 1170
rect -120 1090 -80 1100
rect -10 1170 30 1180
rect -10 1100 0 1170
rect 20 1100 30 1170
rect -10 1090 30 1100
rect 100 1170 140 1180
rect 100 1100 110 1170
rect 130 1100 140 1170
rect 100 1090 140 1100
rect 210 1170 250 1180
rect 210 1100 220 1170
rect 240 1100 250 1170
rect 210 1090 250 1100
rect 320 1170 360 1180
rect 320 1100 330 1170
rect 350 1100 360 1170
rect 395 1175 450 1185
rect 395 1140 405 1175
rect 440 1140 450 1175
rect 395 1130 450 1140
rect 320 1090 360 1100
rect -1510 1070 -1490 1090
rect -630 1085 -610 1090
rect -1565 1050 -1490 1070
rect 340 1070 360 1090
rect 340 1060 380 1070
rect -1565 395 -1545 1050
rect 340 1040 350 1060
rect 370 1040 380 1060
rect 340 1030 380 1040
rect 400 1010 420 1130
rect -980 990 420 1010
rect -980 835 -960 990
rect -910 960 -870 970
rect -910 940 -900 960
rect -880 940 -870 960
rect -910 930 -870 940
rect -900 835 -880 930
rect 35 885 75 895
rect 35 875 45 885
rect -835 865 45 875
rect 65 875 75 885
rect 65 865 420 875
rect -835 855 420 865
rect -835 835 -815 855
rect -110 835 -90 855
rect -1345 825 -1305 835
rect -1345 655 -1335 825
rect -1315 655 -1305 825
rect -1345 645 -1305 655
rect -1280 825 -1240 835
rect -1280 655 -1270 825
rect -1250 655 -1240 825
rect -1280 645 -1240 655
rect -1200 825 -1160 835
rect -1200 655 -1190 825
rect -1170 655 -1160 825
rect -1200 645 -1160 655
rect -1135 825 -1095 835
rect -1135 655 -1125 825
rect -1105 655 -1095 825
rect -1135 645 -1095 655
rect -1055 825 -1015 835
rect -1055 655 -1045 825
rect -1025 655 -1015 825
rect -1055 645 -1015 655
rect -990 825 -950 835
rect -990 655 -980 825
rect -960 655 -950 825
rect -990 645 -950 655
rect -910 825 -870 835
rect -910 655 -900 825
rect -880 655 -870 825
rect -910 645 -870 655
rect -845 825 -805 835
rect -845 655 -835 825
rect -815 655 -805 825
rect -845 645 -805 655
rect -765 825 -725 835
rect -765 655 -755 825
rect -735 655 -725 825
rect -765 645 -725 655
rect -700 825 -660 835
rect -700 655 -690 825
rect -670 675 -660 825
rect -620 825 -580 835
rect -670 655 -655 675
rect -700 645 -655 655
rect -620 655 -610 825
rect -590 655 -580 825
rect -620 645 -580 655
rect -555 825 -515 835
rect -555 655 -545 825
rect -525 655 -515 825
rect -555 645 -515 655
rect -475 825 -435 835
rect -475 655 -465 825
rect -445 655 -435 825
rect -475 645 -435 655
rect -410 825 -370 835
rect -410 655 -400 825
rect -380 655 -370 825
rect -410 645 -370 655
rect -330 825 -290 835
rect -330 655 -320 825
rect -300 655 -290 825
rect -330 645 -290 655
rect -265 825 -225 835
rect -265 655 -255 825
rect -235 655 -225 825
rect -265 645 -225 655
rect -185 825 -145 835
rect -185 655 -175 825
rect -155 655 -145 825
rect -185 645 -145 655
rect -120 825 -80 835
rect -120 655 -110 825
rect -90 655 -80 825
rect -120 645 -80 655
rect -40 825 0 835
rect -40 655 -30 825
rect -10 655 0 825
rect 400 805 420 855
rect 395 795 450 805
rect 395 760 405 795
rect 440 760 450 795
rect 395 750 450 760
rect -40 645 0 655
rect -1260 590 -1240 645
rect -1180 590 -1140 600
rect -1260 570 -1170 590
rect -1150 570 -1140 590
rect -1260 505 -1240 570
rect -1180 560 -1140 570
rect -1115 590 -1095 645
rect -970 625 -950 645
rect -970 615 -930 625
rect -1035 590 -995 600
rect -1115 570 -1025 590
rect -1005 570 -995 590
rect -1115 505 -1095 570
rect -1035 560 -995 570
rect -970 595 -960 615
rect -940 595 -930 615
rect -970 585 -930 595
rect -970 505 -950 585
rect -900 505 -880 645
rect -845 505 -825 645
rect -745 625 -725 645
rect -610 625 -590 645
rect -745 605 -590 625
rect -745 505 -725 605
rect -680 555 -640 565
rect -680 535 -670 555
rect -650 535 -640 555
rect -680 525 -640 535
rect -680 505 -660 525
rect -610 505 -590 605
rect -545 625 -525 645
rect -545 615 -495 625
rect -545 595 -525 615
rect -505 595 -495 615
rect -545 590 -495 595
rect -545 505 -525 590
rect -470 565 -450 645
rect -495 555 -450 565
rect -495 535 -485 555
rect -465 535 -450 555
rect -495 525 -450 535
rect -390 560 -370 645
rect -390 550 -350 560
rect -390 530 -380 550
rect -360 530 -350 550
rect -390 520 -350 530
rect -390 505 -370 520
rect -320 505 -300 645
rect -255 565 -235 645
rect 395 590 450 600
rect 395 565 405 590
rect -255 555 405 565
rect 440 555 450 590
rect -255 545 60 555
rect -255 505 -235 545
rect -110 505 -90 545
rect 50 535 60 545
rect 80 545 450 555
rect 80 535 90 545
rect 50 525 90 535
rect -1345 495 -1305 505
rect -1345 425 -1335 495
rect -1315 425 -1305 495
rect -1345 415 -1305 425
rect -1280 495 -1240 505
rect -1280 425 -1270 495
rect -1250 425 -1240 495
rect -1280 415 -1240 425
rect -1200 495 -1160 505
rect -1200 425 -1190 495
rect -1170 425 -1160 495
rect -1200 415 -1160 425
rect -1135 495 -1095 505
rect -1135 425 -1125 495
rect -1105 425 -1095 495
rect -1135 415 -1095 425
rect -1055 495 -1015 505
rect -1055 425 -1045 495
rect -1025 425 -1015 495
rect -1055 415 -1015 425
rect -990 495 -950 505
rect -990 425 -980 495
rect -960 425 -950 495
rect -990 415 -950 425
rect -910 495 -870 505
rect -910 425 -900 495
rect -880 425 -870 495
rect -910 415 -870 425
rect -845 495 -805 505
rect -845 425 -835 495
rect -815 425 -805 495
rect -845 415 -805 425
rect -765 495 -725 505
rect -765 425 -755 495
rect -735 425 -725 495
rect -765 415 -725 425
rect -700 495 -660 505
rect -700 425 -690 495
rect -670 425 -660 495
rect -700 415 -660 425
rect -620 495 -580 505
rect -620 425 -610 495
rect -590 425 -580 495
rect -620 415 -580 425
rect -555 495 -515 505
rect -555 425 -545 495
rect -525 425 -515 495
rect -555 415 -515 425
rect -475 495 -435 505
rect -475 425 -465 495
rect -445 425 -435 495
rect -475 415 -435 425
rect -410 495 -370 505
rect -410 425 -400 495
rect -380 425 -370 495
rect -410 415 -370 425
rect -330 495 -290 505
rect -330 425 -320 495
rect -300 425 -290 495
rect -330 415 -290 425
rect -265 495 -220 505
rect -265 425 -255 495
rect -235 425 -220 495
rect -265 415 -220 425
rect -185 495 -145 505
rect -185 425 -175 495
rect -155 425 -145 495
rect -185 415 -145 425
rect -120 495 -80 505
rect -120 425 -110 495
rect -90 425 -80 495
rect -120 415 -80 425
rect -40 495 0 505
rect -40 425 -30 495
rect -10 425 0 495
rect -40 415 0 425
rect -1565 375 -810 395
rect -320 380 -300 415
rect -1500 300 -1460 310
rect -1500 280 -1490 300
rect -1470 280 -1460 300
rect -1500 270 -1460 280
rect -1280 300 -1240 310
rect -1280 280 -1270 300
rect -1250 280 -1240 300
rect -1280 270 -1240 280
rect -1060 300 -1020 310
rect -1060 280 -1050 300
rect -1030 280 -1020 300
rect -1060 270 -1020 280
rect -1490 250 -1470 270
rect -1270 250 -1250 270
rect -1050 250 -1030 270
rect -830 250 -810 375
rect -475 360 -300 380
rect -270 385 -230 395
rect -270 365 -260 385
rect -240 375 -230 385
rect 395 375 450 380
rect -240 370 450 375
rect -240 365 405 370
rect -475 330 -455 360
rect -270 355 405 365
rect -495 320 -455 330
rect 395 335 405 355
rect 440 335 450 370
rect 395 325 450 335
rect -495 300 -485 320
rect -465 300 -455 320
rect -495 290 -455 300
rect 340 295 380 305
rect 340 275 350 295
rect 370 275 380 295
rect 340 265 380 275
rect -610 250 -590 255
rect 340 250 360 265
rect -1500 240 -1460 250
rect -1500 170 -1490 240
rect -1470 170 -1460 240
rect -1500 160 -1460 170
rect -1390 240 -1350 250
rect -1390 170 -1380 240
rect -1360 170 -1350 240
rect -1390 160 -1350 170
rect -1280 240 -1240 250
rect -1280 170 -1270 240
rect -1250 170 -1240 240
rect -1280 160 -1240 170
rect -1170 240 -1130 250
rect -1170 170 -1160 240
rect -1140 170 -1130 240
rect -1170 160 -1130 170
rect -1060 240 -1020 250
rect -1060 170 -1050 240
rect -1030 170 -1020 240
rect -1060 160 -1020 170
rect -840 240 -800 250
rect -840 170 -830 240
rect -810 170 -800 240
rect -840 160 -800 170
rect -730 240 -690 250
rect -730 170 -720 240
rect -700 170 -690 240
rect -730 160 -690 170
rect -620 240 -580 250
rect -620 170 -610 240
rect -590 170 -580 240
rect -620 160 -580 170
rect -510 240 -470 250
rect -510 170 -500 240
rect -480 170 -470 240
rect -510 160 -470 170
rect -400 240 -360 250
rect -400 170 -390 240
rect -370 170 -360 240
rect -400 160 -360 170
rect -120 240 -80 250
rect -120 170 -110 240
rect -90 170 -80 240
rect -120 160 -80 170
rect -10 240 30 250
rect -10 170 0 240
rect 20 170 30 240
rect -10 160 30 170
rect 100 240 140 250
rect 100 170 110 240
rect 130 170 140 240
rect 100 160 140 170
rect 210 240 250 250
rect 210 170 220 240
rect 240 170 250 240
rect 210 160 250 170
rect 320 240 360 250
rect 320 170 330 240
rect 350 170 360 240
rect 320 160 360 170
rect -1490 140 -1470 160
rect -1270 140 -1250 160
rect -1050 140 -1030 160
rect -1640 120 -1030 140
rect -830 140 -810 160
rect -610 140 -590 160
rect -390 140 -370 160
rect -830 120 -370 140
rect -110 140 -90 160
rect 110 140 130 160
rect 330 140 350 160
rect -110 120 350 140
<< viali >>
rect -1400 1100 -1380 1170
rect -1180 1100 -1160 1170
rect -960 1100 -940 1170
rect -740 1100 -720 1170
rect -440 1100 -420 1170
rect -220 1100 -200 1170
rect 0 1100 20 1170
rect 220 1100 240 1170
rect 405 1140 440 1175
rect -1335 655 -1315 825
rect -1190 655 -1170 825
rect -1045 655 -1025 825
rect -690 655 -670 825
rect -465 655 -445 825
rect -175 655 -155 825
rect -30 655 -10 825
rect 405 760 440 795
rect 405 555 440 590
rect -1335 425 -1315 495
rect -1190 425 -1170 495
rect -1045 425 -1025 495
rect -690 425 -670 495
rect -465 425 -445 495
rect -175 425 -155 495
rect -30 425 -10 495
rect 405 335 440 370
rect -1380 170 -1360 240
rect -1160 170 -1140 240
rect -720 170 -700 240
rect -500 170 -480 240
rect 0 170 20 240
rect 220 170 240 240
<< metal1 >>
rect -1520 1170 365 1275
rect -1520 1100 -1400 1170
rect -1380 1100 -1180 1170
rect -1160 1100 -960 1170
rect -940 1100 -740 1170
rect -720 1100 -440 1170
rect -420 1100 -220 1170
rect -200 1100 0 1170
rect 20 1100 220 1170
rect 240 1100 365 1170
rect 395 1175 450 1185
rect 395 1140 405 1175
rect 440 1140 450 1175
rect 395 1130 450 1140
rect -1520 825 365 1100
rect -1520 655 -1335 825
rect -1315 655 -1190 825
rect -1170 655 -1045 825
rect -1025 655 -690 825
rect -670 655 -465 825
rect -445 655 -175 825
rect -155 655 -30 825
rect -10 655 365 825
rect 395 795 450 805
rect 395 760 405 795
rect 440 760 450 795
rect 395 750 450 760
rect -1520 640 365 655
rect 395 590 450 600
rect 395 555 405 590
rect 440 555 450 590
rect 395 545 450 555
rect -1520 495 365 510
rect -1520 425 -1335 495
rect -1315 425 -1190 495
rect -1170 425 -1045 495
rect -1025 425 -690 495
rect -670 425 -465 495
rect -445 425 -175 495
rect -155 425 -30 495
rect -10 425 365 495
rect -1520 240 365 425
rect 395 370 450 380
rect 395 335 405 370
rect 440 335 450 370
rect 395 325 450 335
rect -1520 170 -1380 240
rect -1360 170 -1160 240
rect -1140 170 -720 240
rect -700 170 -500 240
rect -480 170 0 240
rect 20 170 220 240
rect 240 170 365 240
rect -1520 155 365 170
<< via1 >>
rect 405 1140 440 1175
rect 405 760 440 795
rect 405 555 440 590
rect 405 335 440 370
<< metal2 >>
rect 395 1175 450 1185
rect 395 1140 405 1175
rect 440 1140 450 1175
rect 395 1130 450 1140
rect 395 795 450 805
rect 395 760 405 795
rect 440 760 450 795
rect 395 750 450 760
rect 395 590 450 600
rect 395 555 405 590
rect 440 555 450 590
rect 395 545 450 555
rect 395 370 450 380
rect 395 335 405 370
rect 440 335 450 370
rect 395 325 450 335
<< via2 >>
rect 405 1140 440 1175
rect 405 760 440 795
rect 405 555 440 590
rect 405 335 440 370
<< metal3 >>
rect 395 1175 1200 1185
rect 395 1140 405 1175
rect 440 1140 1200 1175
rect 395 1130 1200 1140
rect 395 795 450 805
rect 395 760 405 795
rect 440 760 450 795
rect 395 750 450 760
rect 570 735 1200 1130
rect 395 590 450 600
rect 395 555 405 590
rect 440 555 450 590
rect 395 545 450 555
rect 570 380 860 615
rect 395 370 860 380
rect 395 335 405 370
rect 440 335 860 370
rect 395 325 860 335
<< via3 >>
rect 405 760 440 795
rect 405 555 440 590
<< mimcap >>
rect 585 795 1185 1170
rect 585 760 595 795
rect 630 760 1185 795
rect 585 750 1185 760
rect 585 590 845 600
rect 585 555 595 590
rect 630 555 845 590
rect 585 340 845 555
<< mimcapcontact >>
rect 595 760 630 795
rect 595 555 630 590
<< metal4 >>
rect 395 795 640 805
rect 395 760 405 795
rect 440 760 595 795
rect 630 760 640 795
rect 395 750 640 760
rect 395 590 640 600
rect 395 555 405 590
rect 440 555 595 590
rect 630 555 640 590
rect 395 545 640 555
<< labels >>
flabel locali -745 585 -745 585 7 FreeSans 160 0 -80 0 DOWN_b_b
flabel locali -1240 610 -1240 610 3 FreeSans 160 0 80 0 UP_PFD_b
flabel poly 65 940 65 940 3 FreeSans 160 0 80 0 UP_input
flabel poly -1010 905 -1010 905 7 FreeSans 160 0 -80 0 UP
flabel locali -295 990 -295 990 5 FreeSans 160 0 0 -80 UP_b
flabel locali 175 355 175 355 5 FreeSans 160 0 0 -80 DOWN
flabel poly -265 325 -265 325 5 FreeSans 160 0 0 -80 DOWN_b
flabel poly 75 320 75 320 7 FreeSans 160 0 -80 0 DOWN_input
flabel metal1 -1520 285 -1520 285 7 FreeSans 160 0 -80 0 GNDA
flabel locali -1640 130 -1640 130 7 FreeSans 160 0 -80 0 I_IN
flabel metal1 -1520 875 -1520 875 7 FreeSans 160 0 -80 0 VDDA
flabel poly -1665 575 -1665 575 7 FreeSans 160 0 -80 0 UP_PFD
flabel poly -1665 365 -1665 365 7 FreeSans 160 0 -80 0 DOWN_PFD
flabel poly 1245 660 1245 660 3 FreeSans 400 0 200 0 VOUT
<< end >>
