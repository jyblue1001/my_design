magic
tech sky130A
timestamp 1746520359
<< nwell >>
rect 2150 1850 4655 2750
<< pwell >>
rect 2810 1560 3650 1660
<< nmos >>
rect 2850 1560 2910 1660
rect 2950 1560 3010 1660
rect 3050 1560 3110 1660
rect 3150 1560 3210 1660
rect 3250 1560 3310 1660
rect 3350 1560 3410 1660
rect 3450 1560 3510 1660
rect 3550 1560 3610 1660
rect 2770 985 3170 1385
rect 3290 985 3690 1385
rect 2720 755 3720 855
<< pmos >>
rect 2650 2330 2710 2730
rect 2750 2330 2810 2730
rect 2850 2330 2910 2730
rect 2950 2330 3010 2730
rect 3050 2330 3110 2730
rect 3150 2330 3210 2730
rect 3250 2330 3310 2730
rect 3350 2330 3410 2730
rect 3450 2330 3510 2730
rect 3550 2330 3610 2730
rect 3650 2330 3710 2730
rect 3750 2330 3810 2730
rect 2650 1910 2710 2110
rect 2750 1910 2810 2110
rect 2850 1910 2910 2110
rect 2950 1910 3010 2110
rect 3050 1910 3110 2110
rect 3150 1910 3210 2110
rect 3250 1910 3310 2110
rect 3350 1910 3410 2110
rect 3450 1910 3510 2110
rect 3550 1910 3610 2110
rect 3650 1910 3710 2110
rect 3750 1910 3810 2110
rect 4415 1910 4430 2110
rect 4540 1910 4555 2110
<< ndiff >>
rect 2810 1645 2850 1660
rect 2810 1625 2820 1645
rect 2840 1625 2850 1645
rect 2810 1595 2850 1625
rect 2810 1575 2820 1595
rect 2840 1575 2850 1595
rect 2810 1560 2850 1575
rect 2910 1645 2950 1660
rect 2910 1625 2920 1645
rect 2940 1625 2950 1645
rect 2910 1595 2950 1625
rect 2910 1575 2920 1595
rect 2940 1575 2950 1595
rect 2910 1560 2950 1575
rect 3010 1645 3050 1660
rect 3010 1625 3020 1645
rect 3040 1625 3050 1645
rect 3010 1595 3050 1625
rect 3010 1575 3020 1595
rect 3040 1575 3050 1595
rect 3010 1560 3050 1575
rect 3110 1645 3150 1660
rect 3110 1625 3120 1645
rect 3140 1625 3150 1645
rect 3110 1595 3150 1625
rect 3110 1575 3120 1595
rect 3140 1575 3150 1595
rect 3110 1560 3150 1575
rect 3210 1645 3250 1660
rect 3210 1625 3220 1645
rect 3240 1625 3250 1645
rect 3210 1595 3250 1625
rect 3210 1575 3220 1595
rect 3240 1575 3250 1595
rect 3210 1560 3250 1575
rect 3310 1645 3350 1660
rect 3310 1625 3320 1645
rect 3340 1625 3350 1645
rect 3310 1595 3350 1625
rect 3310 1575 3320 1595
rect 3340 1575 3350 1595
rect 3310 1560 3350 1575
rect 3410 1645 3450 1660
rect 3410 1625 3420 1645
rect 3440 1625 3450 1645
rect 3410 1595 3450 1625
rect 3410 1575 3420 1595
rect 3440 1575 3450 1595
rect 3410 1560 3450 1575
rect 3510 1645 3550 1660
rect 3510 1625 3520 1645
rect 3540 1625 3550 1645
rect 3510 1595 3550 1625
rect 3510 1575 3520 1595
rect 3540 1575 3550 1595
rect 3510 1560 3550 1575
rect 3610 1645 3650 1660
rect 3610 1625 3620 1645
rect 3640 1625 3650 1645
rect 3610 1595 3650 1625
rect 3610 1575 3620 1595
rect 3640 1575 3650 1595
rect 3610 1560 3650 1575
rect 2730 1370 2770 1385
rect 2730 1350 2740 1370
rect 2760 1350 2770 1370
rect 2730 1320 2770 1350
rect 2730 1300 2740 1320
rect 2760 1300 2770 1320
rect 2730 1270 2770 1300
rect 2730 1250 2740 1270
rect 2760 1250 2770 1270
rect 2730 1220 2770 1250
rect 2730 1200 2740 1220
rect 2760 1200 2770 1220
rect 2730 1170 2770 1200
rect 2730 1150 2740 1170
rect 2760 1150 2770 1170
rect 2730 1120 2770 1150
rect 2730 1100 2740 1120
rect 2760 1100 2770 1120
rect 2730 1070 2770 1100
rect 2730 1050 2740 1070
rect 2760 1050 2770 1070
rect 2730 1020 2770 1050
rect 2730 1000 2740 1020
rect 2760 1000 2770 1020
rect 2730 985 2770 1000
rect 3170 1370 3210 1385
rect 3250 1370 3290 1385
rect 3170 1350 3180 1370
rect 3200 1350 3210 1370
rect 3250 1350 3260 1370
rect 3280 1350 3290 1370
rect 3170 1320 3210 1350
rect 3250 1320 3290 1350
rect 3170 1300 3180 1320
rect 3200 1300 3210 1320
rect 3250 1300 3260 1320
rect 3280 1300 3290 1320
rect 3170 1270 3210 1300
rect 3250 1270 3290 1300
rect 3170 1250 3180 1270
rect 3200 1250 3210 1270
rect 3250 1250 3260 1270
rect 3280 1250 3290 1270
rect 3170 1220 3210 1250
rect 3250 1220 3290 1250
rect 3170 1200 3180 1220
rect 3200 1200 3210 1220
rect 3250 1200 3260 1220
rect 3280 1200 3290 1220
rect 3170 1170 3210 1200
rect 3250 1170 3290 1200
rect 3170 1150 3180 1170
rect 3200 1150 3210 1170
rect 3250 1150 3260 1170
rect 3280 1150 3290 1170
rect 3170 1120 3210 1150
rect 3250 1120 3290 1150
rect 3170 1100 3180 1120
rect 3200 1100 3210 1120
rect 3250 1100 3260 1120
rect 3280 1100 3290 1120
rect 3170 1070 3210 1100
rect 3250 1070 3290 1100
rect 3170 1050 3180 1070
rect 3200 1050 3210 1070
rect 3250 1050 3260 1070
rect 3280 1050 3290 1070
rect 3170 1020 3210 1050
rect 3250 1020 3290 1050
rect 3170 1000 3180 1020
rect 3200 1000 3210 1020
rect 3250 1000 3260 1020
rect 3280 1000 3290 1020
rect 3170 985 3210 1000
rect 3250 985 3290 1000
rect 3690 1370 3730 1385
rect 3690 1350 3700 1370
rect 3720 1350 3730 1370
rect 3690 1320 3730 1350
rect 3690 1300 3700 1320
rect 3720 1300 3730 1320
rect 3690 1270 3730 1300
rect 3690 1250 3700 1270
rect 3720 1250 3730 1270
rect 3690 1220 3730 1250
rect 3690 1200 3700 1220
rect 3720 1200 3730 1220
rect 3690 1170 3730 1200
rect 3690 1150 3700 1170
rect 3720 1150 3730 1170
rect 3690 1120 3730 1150
rect 3690 1100 3700 1120
rect 3720 1100 3730 1120
rect 3690 1070 3730 1100
rect 3690 1050 3700 1070
rect 3720 1050 3730 1070
rect 3690 1020 3730 1050
rect 3690 1000 3700 1020
rect 3720 1000 3730 1020
rect 3690 985 3730 1000
rect 2680 840 2720 855
rect 2680 820 2690 840
rect 2710 820 2720 840
rect 2680 790 2720 820
rect 2680 770 2690 790
rect 2710 770 2720 790
rect 2680 755 2720 770
rect 3720 840 3760 855
rect 3720 820 3730 840
rect 3750 820 3760 840
rect 3720 790 3760 820
rect 3720 770 3730 790
rect 3750 770 3760 790
rect 3720 755 3760 770
<< pdiff >>
rect 2610 2715 2650 2730
rect 2610 2695 2620 2715
rect 2640 2695 2650 2715
rect 2610 2665 2650 2695
rect 2610 2645 2620 2665
rect 2640 2645 2650 2665
rect 2610 2615 2650 2645
rect 2610 2595 2620 2615
rect 2640 2595 2650 2615
rect 2610 2565 2650 2595
rect 2610 2545 2620 2565
rect 2640 2545 2650 2565
rect 2610 2515 2650 2545
rect 2610 2495 2620 2515
rect 2640 2495 2650 2515
rect 2610 2465 2650 2495
rect 2610 2445 2620 2465
rect 2640 2445 2650 2465
rect 2610 2415 2650 2445
rect 2610 2395 2620 2415
rect 2640 2395 2650 2415
rect 2610 2365 2650 2395
rect 2610 2345 2620 2365
rect 2640 2345 2650 2365
rect 2610 2330 2650 2345
rect 2710 2715 2750 2730
rect 2710 2695 2720 2715
rect 2740 2695 2750 2715
rect 2710 2665 2750 2695
rect 2710 2645 2720 2665
rect 2740 2645 2750 2665
rect 2710 2615 2750 2645
rect 2710 2595 2720 2615
rect 2740 2595 2750 2615
rect 2710 2565 2750 2595
rect 2710 2545 2720 2565
rect 2740 2545 2750 2565
rect 2710 2515 2750 2545
rect 2710 2495 2720 2515
rect 2740 2495 2750 2515
rect 2710 2465 2750 2495
rect 2710 2445 2720 2465
rect 2740 2445 2750 2465
rect 2710 2415 2750 2445
rect 2710 2395 2720 2415
rect 2740 2395 2750 2415
rect 2710 2365 2750 2395
rect 2710 2345 2720 2365
rect 2740 2345 2750 2365
rect 2710 2330 2750 2345
rect 2810 2715 2850 2730
rect 2810 2695 2820 2715
rect 2840 2695 2850 2715
rect 2810 2665 2850 2695
rect 2810 2645 2820 2665
rect 2840 2645 2850 2665
rect 2810 2615 2850 2645
rect 2810 2595 2820 2615
rect 2840 2595 2850 2615
rect 2810 2565 2850 2595
rect 2810 2545 2820 2565
rect 2840 2545 2850 2565
rect 2810 2515 2850 2545
rect 2810 2495 2820 2515
rect 2840 2495 2850 2515
rect 2810 2465 2850 2495
rect 2810 2445 2820 2465
rect 2840 2445 2850 2465
rect 2810 2415 2850 2445
rect 2810 2395 2820 2415
rect 2840 2395 2850 2415
rect 2810 2365 2850 2395
rect 2810 2345 2820 2365
rect 2840 2345 2850 2365
rect 2810 2330 2850 2345
rect 2910 2715 2950 2730
rect 2910 2695 2920 2715
rect 2940 2695 2950 2715
rect 2910 2665 2950 2695
rect 2910 2645 2920 2665
rect 2940 2645 2950 2665
rect 2910 2615 2950 2645
rect 2910 2595 2920 2615
rect 2940 2595 2950 2615
rect 2910 2565 2950 2595
rect 2910 2545 2920 2565
rect 2940 2545 2950 2565
rect 2910 2515 2950 2545
rect 2910 2495 2920 2515
rect 2940 2495 2950 2515
rect 2910 2465 2950 2495
rect 2910 2445 2920 2465
rect 2940 2445 2950 2465
rect 2910 2415 2950 2445
rect 2910 2395 2920 2415
rect 2940 2395 2950 2415
rect 2910 2365 2950 2395
rect 2910 2345 2920 2365
rect 2940 2345 2950 2365
rect 2910 2330 2950 2345
rect 3010 2715 3050 2730
rect 3010 2695 3020 2715
rect 3040 2695 3050 2715
rect 3010 2665 3050 2695
rect 3010 2645 3020 2665
rect 3040 2645 3050 2665
rect 3010 2615 3050 2645
rect 3010 2595 3020 2615
rect 3040 2595 3050 2615
rect 3010 2565 3050 2595
rect 3010 2545 3020 2565
rect 3040 2545 3050 2565
rect 3010 2515 3050 2545
rect 3010 2495 3020 2515
rect 3040 2495 3050 2515
rect 3010 2465 3050 2495
rect 3010 2445 3020 2465
rect 3040 2445 3050 2465
rect 3010 2415 3050 2445
rect 3010 2395 3020 2415
rect 3040 2395 3050 2415
rect 3010 2365 3050 2395
rect 3010 2345 3020 2365
rect 3040 2345 3050 2365
rect 3010 2330 3050 2345
rect 3110 2715 3150 2730
rect 3110 2695 3120 2715
rect 3140 2695 3150 2715
rect 3110 2665 3150 2695
rect 3110 2645 3120 2665
rect 3140 2645 3150 2665
rect 3110 2615 3150 2645
rect 3110 2595 3120 2615
rect 3140 2595 3150 2615
rect 3110 2565 3150 2595
rect 3110 2545 3120 2565
rect 3140 2545 3150 2565
rect 3110 2515 3150 2545
rect 3110 2495 3120 2515
rect 3140 2495 3150 2515
rect 3110 2465 3150 2495
rect 3110 2445 3120 2465
rect 3140 2445 3150 2465
rect 3110 2415 3150 2445
rect 3110 2395 3120 2415
rect 3140 2395 3150 2415
rect 3110 2365 3150 2395
rect 3110 2345 3120 2365
rect 3140 2345 3150 2365
rect 3110 2330 3150 2345
rect 3210 2715 3250 2730
rect 3210 2695 3220 2715
rect 3240 2695 3250 2715
rect 3210 2665 3250 2695
rect 3210 2645 3220 2665
rect 3240 2645 3250 2665
rect 3210 2615 3250 2645
rect 3210 2595 3220 2615
rect 3240 2595 3250 2615
rect 3210 2565 3250 2595
rect 3210 2545 3220 2565
rect 3240 2545 3250 2565
rect 3210 2515 3250 2545
rect 3210 2495 3220 2515
rect 3240 2495 3250 2515
rect 3210 2465 3250 2495
rect 3210 2445 3220 2465
rect 3240 2445 3250 2465
rect 3210 2415 3250 2445
rect 3210 2395 3220 2415
rect 3240 2395 3250 2415
rect 3210 2365 3250 2395
rect 3210 2345 3220 2365
rect 3240 2345 3250 2365
rect 3210 2330 3250 2345
rect 3310 2715 3350 2730
rect 3310 2695 3320 2715
rect 3340 2695 3350 2715
rect 3310 2665 3350 2695
rect 3310 2645 3320 2665
rect 3340 2645 3350 2665
rect 3310 2615 3350 2645
rect 3310 2595 3320 2615
rect 3340 2595 3350 2615
rect 3310 2565 3350 2595
rect 3310 2545 3320 2565
rect 3340 2545 3350 2565
rect 3310 2515 3350 2545
rect 3310 2495 3320 2515
rect 3340 2495 3350 2515
rect 3310 2465 3350 2495
rect 3310 2445 3320 2465
rect 3340 2445 3350 2465
rect 3310 2415 3350 2445
rect 3310 2395 3320 2415
rect 3340 2395 3350 2415
rect 3310 2365 3350 2395
rect 3310 2345 3320 2365
rect 3340 2345 3350 2365
rect 3310 2330 3350 2345
rect 3410 2715 3450 2730
rect 3410 2695 3420 2715
rect 3440 2695 3450 2715
rect 3410 2665 3450 2695
rect 3410 2645 3420 2665
rect 3440 2645 3450 2665
rect 3410 2615 3450 2645
rect 3410 2595 3420 2615
rect 3440 2595 3450 2615
rect 3410 2565 3450 2595
rect 3410 2545 3420 2565
rect 3440 2545 3450 2565
rect 3410 2515 3450 2545
rect 3410 2495 3420 2515
rect 3440 2495 3450 2515
rect 3410 2465 3450 2495
rect 3410 2445 3420 2465
rect 3440 2445 3450 2465
rect 3410 2415 3450 2445
rect 3410 2395 3420 2415
rect 3440 2395 3450 2415
rect 3410 2365 3450 2395
rect 3410 2345 3420 2365
rect 3440 2345 3450 2365
rect 3410 2330 3450 2345
rect 3510 2715 3550 2730
rect 3510 2695 3520 2715
rect 3540 2695 3550 2715
rect 3510 2665 3550 2695
rect 3510 2645 3520 2665
rect 3540 2645 3550 2665
rect 3510 2615 3550 2645
rect 3510 2595 3520 2615
rect 3540 2595 3550 2615
rect 3510 2565 3550 2595
rect 3510 2545 3520 2565
rect 3540 2545 3550 2565
rect 3510 2515 3550 2545
rect 3510 2495 3520 2515
rect 3540 2495 3550 2515
rect 3510 2465 3550 2495
rect 3510 2445 3520 2465
rect 3540 2445 3550 2465
rect 3510 2415 3550 2445
rect 3510 2395 3520 2415
rect 3540 2395 3550 2415
rect 3510 2365 3550 2395
rect 3510 2345 3520 2365
rect 3540 2345 3550 2365
rect 3510 2330 3550 2345
rect 3610 2715 3650 2730
rect 3610 2695 3620 2715
rect 3640 2695 3650 2715
rect 3610 2665 3650 2695
rect 3610 2645 3620 2665
rect 3640 2645 3650 2665
rect 3610 2615 3650 2645
rect 3610 2595 3620 2615
rect 3640 2595 3650 2615
rect 3610 2565 3650 2595
rect 3610 2545 3620 2565
rect 3640 2545 3650 2565
rect 3610 2515 3650 2545
rect 3610 2495 3620 2515
rect 3640 2495 3650 2515
rect 3610 2465 3650 2495
rect 3610 2445 3620 2465
rect 3640 2445 3650 2465
rect 3610 2415 3650 2445
rect 3610 2395 3620 2415
rect 3640 2395 3650 2415
rect 3610 2365 3650 2395
rect 3610 2345 3620 2365
rect 3640 2345 3650 2365
rect 3610 2330 3650 2345
rect 3710 2715 3750 2730
rect 3710 2695 3720 2715
rect 3740 2695 3750 2715
rect 3710 2665 3750 2695
rect 3710 2645 3720 2665
rect 3740 2645 3750 2665
rect 3710 2615 3750 2645
rect 3710 2595 3720 2615
rect 3740 2595 3750 2615
rect 3710 2565 3750 2595
rect 3710 2545 3720 2565
rect 3740 2545 3750 2565
rect 3710 2515 3750 2545
rect 3710 2495 3720 2515
rect 3740 2495 3750 2515
rect 3710 2465 3750 2495
rect 3710 2445 3720 2465
rect 3740 2445 3750 2465
rect 3710 2415 3750 2445
rect 3710 2395 3720 2415
rect 3740 2395 3750 2415
rect 3710 2365 3750 2395
rect 3710 2345 3720 2365
rect 3740 2345 3750 2365
rect 3710 2330 3750 2345
rect 3810 2715 3850 2730
rect 3810 2695 3820 2715
rect 3840 2695 3850 2715
rect 3810 2665 3850 2695
rect 3810 2645 3820 2665
rect 3840 2645 3850 2665
rect 3810 2615 3850 2645
rect 3810 2595 3820 2615
rect 3840 2595 3850 2615
rect 3810 2565 3850 2595
rect 3810 2545 3820 2565
rect 3840 2545 3850 2565
rect 3810 2515 3850 2545
rect 3810 2495 3820 2515
rect 3840 2495 3850 2515
rect 3810 2465 3850 2495
rect 3810 2445 3820 2465
rect 3840 2445 3850 2465
rect 3810 2415 3850 2445
rect 3810 2395 3820 2415
rect 3840 2395 3850 2415
rect 3810 2365 3850 2395
rect 3810 2345 3820 2365
rect 3840 2345 3850 2365
rect 3810 2330 3850 2345
rect 2610 2095 2650 2110
rect 2610 2075 2620 2095
rect 2640 2075 2650 2095
rect 2610 2045 2650 2075
rect 2610 2025 2620 2045
rect 2640 2025 2650 2045
rect 2610 1995 2650 2025
rect 2610 1975 2620 1995
rect 2640 1975 2650 1995
rect 2610 1945 2650 1975
rect 2610 1925 2620 1945
rect 2640 1925 2650 1945
rect 2610 1910 2650 1925
rect 2710 2095 2750 2110
rect 2710 2075 2720 2095
rect 2740 2075 2750 2095
rect 2710 2045 2750 2075
rect 2710 2025 2720 2045
rect 2740 2025 2750 2045
rect 2710 1995 2750 2025
rect 2710 1975 2720 1995
rect 2740 1975 2750 1995
rect 2710 1945 2750 1975
rect 2710 1925 2720 1945
rect 2740 1925 2750 1945
rect 2710 1910 2750 1925
rect 2810 2095 2850 2110
rect 2810 2075 2820 2095
rect 2840 2075 2850 2095
rect 2810 2045 2850 2075
rect 2810 2025 2820 2045
rect 2840 2025 2850 2045
rect 2810 1995 2850 2025
rect 2810 1975 2820 1995
rect 2840 1975 2850 1995
rect 2810 1945 2850 1975
rect 2810 1925 2820 1945
rect 2840 1925 2850 1945
rect 2810 1910 2850 1925
rect 2910 2095 2950 2110
rect 2910 2075 2920 2095
rect 2940 2075 2950 2095
rect 2910 2045 2950 2075
rect 2910 2025 2920 2045
rect 2940 2025 2950 2045
rect 2910 1995 2950 2025
rect 2910 1975 2920 1995
rect 2940 1975 2950 1995
rect 2910 1945 2950 1975
rect 2910 1925 2920 1945
rect 2940 1925 2950 1945
rect 2910 1910 2950 1925
rect 3010 2095 3050 2110
rect 3010 2075 3020 2095
rect 3040 2075 3050 2095
rect 3010 2045 3050 2075
rect 3010 2025 3020 2045
rect 3040 2025 3050 2045
rect 3010 1995 3050 2025
rect 3010 1975 3020 1995
rect 3040 1975 3050 1995
rect 3010 1945 3050 1975
rect 3010 1925 3020 1945
rect 3040 1925 3050 1945
rect 3010 1910 3050 1925
rect 3110 2095 3150 2110
rect 3110 2075 3120 2095
rect 3140 2075 3150 2095
rect 3110 2045 3150 2075
rect 3110 2025 3120 2045
rect 3140 2025 3150 2045
rect 3110 1995 3150 2025
rect 3110 1975 3120 1995
rect 3140 1975 3150 1995
rect 3110 1945 3150 1975
rect 3110 1925 3120 1945
rect 3140 1925 3150 1945
rect 3110 1910 3150 1925
rect 3210 2095 3250 2110
rect 3210 2075 3220 2095
rect 3240 2075 3250 2095
rect 3210 2045 3250 2075
rect 3210 2025 3220 2045
rect 3240 2025 3250 2045
rect 3210 1995 3250 2025
rect 3210 1975 3220 1995
rect 3240 1975 3250 1995
rect 3210 1945 3250 1975
rect 3210 1925 3220 1945
rect 3240 1925 3250 1945
rect 3210 1910 3250 1925
rect 3310 2095 3350 2110
rect 3310 2075 3320 2095
rect 3340 2075 3350 2095
rect 3310 2045 3350 2075
rect 3310 2025 3320 2045
rect 3340 2025 3350 2045
rect 3310 1995 3350 2025
rect 3310 1975 3320 1995
rect 3340 1975 3350 1995
rect 3310 1945 3350 1975
rect 3310 1925 3320 1945
rect 3340 1925 3350 1945
rect 3310 1910 3350 1925
rect 3410 2095 3450 2110
rect 3410 2075 3420 2095
rect 3440 2075 3450 2095
rect 3410 2045 3450 2075
rect 3410 2025 3420 2045
rect 3440 2025 3450 2045
rect 3410 1995 3450 2025
rect 3410 1975 3420 1995
rect 3440 1975 3450 1995
rect 3410 1945 3450 1975
rect 3410 1925 3420 1945
rect 3440 1925 3450 1945
rect 3410 1910 3450 1925
rect 3510 2095 3550 2110
rect 3510 2075 3520 2095
rect 3540 2075 3550 2095
rect 3510 2045 3550 2075
rect 3510 2025 3520 2045
rect 3540 2025 3550 2045
rect 3510 1995 3550 2025
rect 3510 1975 3520 1995
rect 3540 1975 3550 1995
rect 3510 1945 3550 1975
rect 3510 1925 3520 1945
rect 3540 1925 3550 1945
rect 3510 1910 3550 1925
rect 3610 2095 3650 2110
rect 3610 2075 3620 2095
rect 3640 2075 3650 2095
rect 3610 2045 3650 2075
rect 3610 2025 3620 2045
rect 3640 2025 3650 2045
rect 3610 1995 3650 2025
rect 3610 1975 3620 1995
rect 3640 1975 3650 1995
rect 3610 1945 3650 1975
rect 3610 1925 3620 1945
rect 3640 1925 3650 1945
rect 3610 1910 3650 1925
rect 3710 2095 3750 2110
rect 3710 2075 3720 2095
rect 3740 2075 3750 2095
rect 3710 2045 3750 2075
rect 3710 2025 3720 2045
rect 3740 2025 3750 2045
rect 3710 1995 3750 2025
rect 3710 1975 3720 1995
rect 3740 1975 3750 1995
rect 3710 1945 3750 1975
rect 3710 1925 3720 1945
rect 3740 1925 3750 1945
rect 3710 1910 3750 1925
rect 3810 2095 3850 2110
rect 3810 2075 3820 2095
rect 3840 2075 3850 2095
rect 3810 2045 3850 2075
rect 3810 2025 3820 2045
rect 3840 2025 3850 2045
rect 3810 1995 3850 2025
rect 3810 1975 3820 1995
rect 3840 1975 3850 1995
rect 3810 1945 3850 1975
rect 3810 1925 3820 1945
rect 3840 1925 3850 1945
rect 3810 1910 3850 1925
rect 4375 2095 4415 2110
rect 4375 2075 4385 2095
rect 4405 2075 4415 2095
rect 4375 2045 4415 2075
rect 4375 2025 4385 2045
rect 4405 2025 4415 2045
rect 4375 1995 4415 2025
rect 4375 1975 4385 1995
rect 4405 1975 4415 1995
rect 4375 1945 4415 1975
rect 4375 1925 4385 1945
rect 4405 1925 4415 1945
rect 4375 1910 4415 1925
rect 4430 2095 4470 2110
rect 4430 2075 4440 2095
rect 4460 2075 4470 2095
rect 4430 2045 4470 2075
rect 4430 2025 4440 2045
rect 4460 2025 4470 2045
rect 4430 1995 4470 2025
rect 4430 1975 4440 1995
rect 4460 1975 4470 1995
rect 4430 1945 4470 1975
rect 4430 1925 4440 1945
rect 4460 1925 4470 1945
rect 4430 1910 4470 1925
rect 4500 2095 4540 2110
rect 4500 2075 4510 2095
rect 4530 2075 4540 2095
rect 4500 2045 4540 2075
rect 4500 2025 4510 2045
rect 4530 2025 4540 2045
rect 4500 1995 4540 2025
rect 4500 1975 4510 1995
rect 4530 1975 4540 1995
rect 4500 1945 4540 1975
rect 4500 1925 4510 1945
rect 4530 1925 4540 1945
rect 4500 1910 4540 1925
rect 4555 2095 4595 2110
rect 4555 2075 4565 2095
rect 4585 2075 4595 2095
rect 4555 2045 4595 2075
rect 4555 2025 4565 2045
rect 4585 2025 4595 2045
rect 4555 1995 4595 2025
rect 4555 1975 4565 1995
rect 4585 1975 4595 1995
rect 4555 1945 4595 1975
rect 4555 1925 4565 1945
rect 4585 1925 4595 1945
rect 4555 1910 4595 1925
<< ndiffc >>
rect 2820 1625 2840 1645
rect 2820 1575 2840 1595
rect 2920 1625 2940 1645
rect 2920 1575 2940 1595
rect 3020 1625 3040 1645
rect 3020 1575 3040 1595
rect 3120 1625 3140 1645
rect 3120 1575 3140 1595
rect 3220 1625 3240 1645
rect 3220 1575 3240 1595
rect 3320 1625 3340 1645
rect 3320 1575 3340 1595
rect 3420 1625 3440 1645
rect 3420 1575 3440 1595
rect 3520 1625 3540 1645
rect 3520 1575 3540 1595
rect 3620 1625 3640 1645
rect 3620 1575 3640 1595
rect 2740 1350 2760 1370
rect 2740 1300 2760 1320
rect 2740 1250 2760 1270
rect 2740 1200 2760 1220
rect 2740 1150 2760 1170
rect 2740 1100 2760 1120
rect 2740 1050 2760 1070
rect 2740 1000 2760 1020
rect 3180 1350 3200 1370
rect 3260 1350 3280 1370
rect 3180 1300 3200 1320
rect 3260 1300 3280 1320
rect 3180 1250 3200 1270
rect 3260 1250 3280 1270
rect 3180 1200 3200 1220
rect 3260 1200 3280 1220
rect 3180 1150 3200 1170
rect 3260 1150 3280 1170
rect 3180 1100 3200 1120
rect 3260 1100 3280 1120
rect 3180 1050 3200 1070
rect 3260 1050 3280 1070
rect 3180 1000 3200 1020
rect 3260 1000 3280 1020
rect 3700 1350 3720 1370
rect 3700 1300 3720 1320
rect 3700 1250 3720 1270
rect 3700 1200 3720 1220
rect 3700 1150 3720 1170
rect 3700 1100 3720 1120
rect 3700 1050 3720 1070
rect 3700 1000 3720 1020
rect 2690 820 2710 840
rect 2690 770 2710 790
rect 3730 820 3750 840
rect 3730 770 3750 790
<< pdiffc >>
rect 2620 2695 2640 2715
rect 2620 2645 2640 2665
rect 2620 2595 2640 2615
rect 2620 2545 2640 2565
rect 2620 2495 2640 2515
rect 2620 2445 2640 2465
rect 2620 2395 2640 2415
rect 2620 2345 2640 2365
rect 2720 2695 2740 2715
rect 2720 2645 2740 2665
rect 2720 2595 2740 2615
rect 2720 2545 2740 2565
rect 2720 2495 2740 2515
rect 2720 2445 2740 2465
rect 2720 2395 2740 2415
rect 2720 2345 2740 2365
rect 2820 2695 2840 2715
rect 2820 2645 2840 2665
rect 2820 2595 2840 2615
rect 2820 2545 2840 2565
rect 2820 2495 2840 2515
rect 2820 2445 2840 2465
rect 2820 2395 2840 2415
rect 2820 2345 2840 2365
rect 2920 2695 2940 2715
rect 2920 2645 2940 2665
rect 2920 2595 2940 2615
rect 2920 2545 2940 2565
rect 2920 2495 2940 2515
rect 2920 2445 2940 2465
rect 2920 2395 2940 2415
rect 2920 2345 2940 2365
rect 3020 2695 3040 2715
rect 3020 2645 3040 2665
rect 3020 2595 3040 2615
rect 3020 2545 3040 2565
rect 3020 2495 3040 2515
rect 3020 2445 3040 2465
rect 3020 2395 3040 2415
rect 3020 2345 3040 2365
rect 3120 2695 3140 2715
rect 3120 2645 3140 2665
rect 3120 2595 3140 2615
rect 3120 2545 3140 2565
rect 3120 2495 3140 2515
rect 3120 2445 3140 2465
rect 3120 2395 3140 2415
rect 3120 2345 3140 2365
rect 3220 2695 3240 2715
rect 3220 2645 3240 2665
rect 3220 2595 3240 2615
rect 3220 2545 3240 2565
rect 3220 2495 3240 2515
rect 3220 2445 3240 2465
rect 3220 2395 3240 2415
rect 3220 2345 3240 2365
rect 3320 2695 3340 2715
rect 3320 2645 3340 2665
rect 3320 2595 3340 2615
rect 3320 2545 3340 2565
rect 3320 2495 3340 2515
rect 3320 2445 3340 2465
rect 3320 2395 3340 2415
rect 3320 2345 3340 2365
rect 3420 2695 3440 2715
rect 3420 2645 3440 2665
rect 3420 2595 3440 2615
rect 3420 2545 3440 2565
rect 3420 2495 3440 2515
rect 3420 2445 3440 2465
rect 3420 2395 3440 2415
rect 3420 2345 3440 2365
rect 3520 2695 3540 2715
rect 3520 2645 3540 2665
rect 3520 2595 3540 2615
rect 3520 2545 3540 2565
rect 3520 2495 3540 2515
rect 3520 2445 3540 2465
rect 3520 2395 3540 2415
rect 3520 2345 3540 2365
rect 3620 2695 3640 2715
rect 3620 2645 3640 2665
rect 3620 2595 3640 2615
rect 3620 2545 3640 2565
rect 3620 2495 3640 2515
rect 3620 2445 3640 2465
rect 3620 2395 3640 2415
rect 3620 2345 3640 2365
rect 3720 2695 3740 2715
rect 3720 2645 3740 2665
rect 3720 2595 3740 2615
rect 3720 2545 3740 2565
rect 3720 2495 3740 2515
rect 3720 2445 3740 2465
rect 3720 2395 3740 2415
rect 3720 2345 3740 2365
rect 3820 2695 3840 2715
rect 3820 2645 3840 2665
rect 3820 2595 3840 2615
rect 3820 2545 3840 2565
rect 3820 2495 3840 2515
rect 3820 2445 3840 2465
rect 3820 2395 3840 2415
rect 3820 2345 3840 2365
rect 2620 2075 2640 2095
rect 2620 2025 2640 2045
rect 2620 1975 2640 1995
rect 2620 1925 2640 1945
rect 2720 2075 2740 2095
rect 2720 2025 2740 2045
rect 2720 1975 2740 1995
rect 2720 1925 2740 1945
rect 2820 2075 2840 2095
rect 2820 2025 2840 2045
rect 2820 1975 2840 1995
rect 2820 1925 2840 1945
rect 2920 2075 2940 2095
rect 2920 2025 2940 2045
rect 2920 1975 2940 1995
rect 2920 1925 2940 1945
rect 3020 2075 3040 2095
rect 3020 2025 3040 2045
rect 3020 1975 3040 1995
rect 3020 1925 3040 1945
rect 3120 2075 3140 2095
rect 3120 2025 3140 2045
rect 3120 1975 3140 1995
rect 3120 1925 3140 1945
rect 3220 2075 3240 2095
rect 3220 2025 3240 2045
rect 3220 1975 3240 1995
rect 3220 1925 3240 1945
rect 3320 2075 3340 2095
rect 3320 2025 3340 2045
rect 3320 1975 3340 1995
rect 3320 1925 3340 1945
rect 3420 2075 3440 2095
rect 3420 2025 3440 2045
rect 3420 1975 3440 1995
rect 3420 1925 3440 1945
rect 3520 2075 3540 2095
rect 3520 2025 3540 2045
rect 3520 1975 3540 1995
rect 3520 1925 3540 1945
rect 3620 2075 3640 2095
rect 3620 2025 3640 2045
rect 3620 1975 3640 1995
rect 3620 1925 3640 1945
rect 3720 2075 3740 2095
rect 3720 2025 3740 2045
rect 3720 1975 3740 1995
rect 3720 1925 3740 1945
rect 3820 2075 3840 2095
rect 3820 2025 3840 2045
rect 3820 1975 3840 1995
rect 3820 1925 3840 1945
rect 4385 2075 4405 2095
rect 4385 2025 4405 2045
rect 4385 1975 4405 1995
rect 4385 1925 4405 1945
rect 4440 2075 4460 2095
rect 4440 2025 4460 2045
rect 4440 1975 4460 1995
rect 4440 1925 4460 1945
rect 4510 2075 4530 2095
rect 4510 2025 4530 2045
rect 4510 1975 4530 1995
rect 4510 1925 4530 1945
rect 4565 2075 4585 2095
rect 4565 2025 4585 2045
rect 4565 1975 4585 1995
rect 4565 1925 4585 1945
<< psubdiff >>
rect 3210 1370 3250 1385
rect 3210 1350 3220 1370
rect 3240 1350 3250 1370
rect 3210 1320 3250 1350
rect 3210 1300 3220 1320
rect 3240 1300 3250 1320
rect 3210 1270 3250 1300
rect 3210 1250 3220 1270
rect 3240 1250 3250 1270
rect 3210 1220 3250 1250
rect 3210 1200 3220 1220
rect 3240 1200 3250 1220
rect 3210 1170 3250 1200
rect 3210 1150 3220 1170
rect 3240 1150 3250 1170
rect 3210 1120 3250 1150
rect 3210 1100 3220 1120
rect 3240 1100 3250 1120
rect 3210 1070 3250 1100
rect 3210 1050 3220 1070
rect 3240 1050 3250 1070
rect 3210 1020 3250 1050
rect 3210 1000 3220 1020
rect 3240 1000 3250 1020
rect 3210 985 3250 1000
rect 645 820 695 835
rect 645 800 660 820
rect 680 800 695 820
rect 645 770 695 800
rect 645 750 660 770
rect 680 750 695 770
rect 3760 840 3800 855
rect 3760 820 3770 840
rect 3790 820 3800 840
rect 3760 790 3800 820
rect 3760 770 3770 790
rect 3790 770 3800 790
rect 3760 755 3800 770
rect 645 720 695 750
rect 645 700 660 720
rect 680 700 695 720
rect 645 685 695 700
<< nsubdiff >>
rect 2570 2715 2610 2730
rect 2570 2695 2580 2715
rect 2600 2695 2610 2715
rect 2570 2665 2610 2695
rect 2570 2645 2580 2665
rect 2600 2645 2610 2665
rect 2570 2615 2610 2645
rect 2570 2595 2580 2615
rect 2600 2595 2610 2615
rect 2570 2565 2610 2595
rect 2570 2545 2580 2565
rect 2600 2545 2610 2565
rect 2570 2515 2610 2545
rect 2570 2495 2580 2515
rect 2600 2495 2610 2515
rect 2570 2465 2610 2495
rect 2570 2445 2580 2465
rect 2600 2445 2610 2465
rect 2570 2415 2610 2445
rect 2570 2395 2580 2415
rect 2600 2395 2610 2415
rect 2570 2365 2610 2395
rect 2570 2345 2580 2365
rect 2600 2345 2610 2365
rect 2570 2330 2610 2345
rect 3850 2715 3890 2730
rect 3850 2695 3860 2715
rect 3880 2695 3890 2715
rect 3850 2665 3890 2695
rect 3850 2645 3860 2665
rect 3880 2645 3890 2665
rect 3850 2615 3890 2645
rect 3850 2595 3860 2615
rect 3880 2595 3890 2615
rect 3850 2565 3890 2595
rect 3850 2545 3860 2565
rect 3880 2545 3890 2565
rect 3850 2515 3890 2545
rect 3850 2495 3860 2515
rect 3880 2495 3890 2515
rect 3850 2465 3890 2495
rect 3850 2445 3860 2465
rect 3880 2445 3890 2465
rect 3850 2415 3890 2445
rect 3850 2395 3860 2415
rect 3880 2395 3890 2415
rect 3850 2365 3890 2395
rect 3850 2345 3860 2365
rect 3880 2345 3890 2365
rect 3850 2330 3890 2345
rect 2570 2095 2610 2110
rect 2570 2075 2580 2095
rect 2600 2075 2610 2095
rect 2570 2045 2610 2075
rect 2570 2025 2580 2045
rect 2600 2025 2610 2045
rect 2570 1995 2610 2025
rect 2570 1975 2580 1995
rect 2600 1975 2610 1995
rect 2570 1945 2610 1975
rect 2570 1925 2580 1945
rect 2600 1925 2610 1945
rect 2570 1910 2610 1925
rect 3850 2095 3890 2110
rect 3850 2075 3860 2095
rect 3880 2075 3890 2095
rect 3850 2045 3890 2075
rect 3850 2025 3860 2045
rect 3880 2025 3890 2045
rect 3850 1995 3890 2025
rect 3850 1975 3860 1995
rect 3880 1975 3890 1995
rect 3850 1945 3890 1975
rect 3850 1925 3860 1945
rect 3880 1925 3890 1945
rect 3850 1910 3890 1925
<< psubdiffcont >>
rect 3220 1350 3240 1370
rect 3220 1300 3240 1320
rect 3220 1250 3240 1270
rect 3220 1200 3240 1220
rect 3220 1150 3240 1170
rect 3220 1100 3240 1120
rect 3220 1050 3240 1070
rect 3220 1000 3240 1020
rect 660 800 680 820
rect 660 750 680 770
rect 3770 820 3790 840
rect 3770 770 3790 790
rect 660 700 680 720
<< nsubdiffcont >>
rect 2580 2695 2600 2715
rect 2580 2645 2600 2665
rect 2580 2595 2600 2615
rect 2580 2545 2600 2565
rect 2580 2495 2600 2515
rect 2580 2445 2600 2465
rect 2580 2395 2600 2415
rect 2580 2345 2600 2365
rect 3860 2695 3880 2715
rect 3860 2645 3880 2665
rect 3860 2595 3880 2615
rect 3860 2545 3880 2565
rect 3860 2495 3880 2515
rect 3860 2445 3880 2465
rect 3860 2395 3880 2415
rect 3860 2345 3880 2365
rect 2580 2075 2600 2095
rect 2580 2025 2600 2045
rect 2580 1975 2600 1995
rect 2580 1925 2600 1945
rect 3860 2075 3880 2095
rect 3860 2025 3880 2045
rect 3860 1975 3880 1995
rect 3860 1925 3880 1945
<< poly >>
rect 2650 2730 2710 2745
rect 2750 2730 2810 2745
rect 2850 2730 2910 2745
rect 2950 2730 3010 2745
rect 3050 2730 3110 2745
rect 3150 2730 3210 2745
rect 3250 2730 3310 2745
rect 3350 2730 3410 2745
rect 3450 2730 3510 2745
rect 3550 2730 3610 2745
rect 3650 2730 3710 2745
rect 3750 2730 3810 2745
rect 2650 2320 2710 2330
rect 2750 2320 2810 2330
rect 2850 2320 2910 2330
rect 2950 2320 3010 2330
rect 3050 2320 3110 2330
rect 3150 2320 3210 2330
rect 3250 2320 3310 2330
rect 3350 2320 3410 2330
rect 3450 2320 3510 2330
rect 3550 2320 3610 2330
rect 3650 2320 3710 2330
rect 3750 2320 3810 2330
rect 2650 2305 3810 2320
rect 4515 2195 4555 2205
rect 4515 2175 4525 2195
rect 4545 2175 4555 2195
rect 4515 2165 4555 2175
rect 2650 2110 2710 2125
rect 2750 2110 2810 2125
rect 2850 2110 2910 2125
rect 2950 2110 3010 2125
rect 3050 2110 3110 2125
rect 3150 2110 3210 2125
rect 3250 2110 3310 2125
rect 3350 2110 3410 2125
rect 3450 2110 3510 2125
rect 3550 2110 3610 2125
rect 3650 2110 3710 2125
rect 3750 2110 3810 2125
rect 4415 2110 4430 2125
rect 4540 2110 4555 2165
rect 2650 1900 2710 1910
rect 2750 1900 2810 1910
rect 2850 1900 2910 1910
rect 2950 1900 3010 1910
rect 2650 1885 3010 1900
rect 3050 1900 3110 1910
rect 3150 1900 3210 1910
rect 3250 1900 3310 1910
rect 3350 1900 3410 1910
rect 3050 1885 3410 1900
rect 3450 1900 3510 1910
rect 3550 1900 3610 1910
rect 3650 1900 3710 1910
rect 3750 1900 3810 1910
rect 3450 1885 3810 1900
rect 2910 1865 2920 1885
rect 2940 1865 2950 1885
rect 2910 1855 2950 1865
rect 3175 1850 3195 1885
rect 3510 1865 3520 1885
rect 3540 1865 3550 1885
rect 3510 1855 3550 1865
rect 4415 1870 4430 1910
rect 4540 1895 4555 1910
rect 4485 1870 4525 1880
rect 4415 1850 4495 1870
rect 4515 1850 4525 1870
rect 3165 1840 3205 1850
rect 4485 1840 4525 1850
rect 3165 1820 3175 1840
rect 3195 1820 3205 1840
rect 3165 1810 3205 1820
rect 3050 1705 3090 1715
rect 3050 1685 3060 1705
rect 3080 1685 3090 1705
rect 3370 1705 3410 1715
rect 3370 1685 3380 1705
rect 3400 1685 3410 1705
rect 2850 1660 2910 1675
rect 2950 1660 3010 1675
rect 3050 1670 3410 1685
rect 3050 1660 3110 1670
rect 3150 1660 3210 1670
rect 3250 1660 3310 1670
rect 3350 1660 3410 1670
rect 3450 1660 3510 1675
rect 3550 1660 3610 1675
rect 2850 1550 2910 1560
rect 2950 1550 3010 1560
rect 2850 1535 3010 1550
rect 3050 1545 3110 1560
rect 3150 1545 3210 1560
rect 3250 1545 3310 1560
rect 3350 1545 3410 1560
rect 3450 1550 3510 1560
rect 3550 1550 3610 1560
rect 3450 1535 3610 1550
rect 2910 1515 2920 1535
rect 2940 1515 2950 1535
rect 2910 1505 2950 1515
rect 3510 1515 3520 1535
rect 3540 1515 3550 1535
rect 3510 1505 3550 1515
rect 2770 1430 3170 1440
rect 2770 1410 2780 1430
rect 2800 1410 2820 1430
rect 2840 1410 2860 1430
rect 2880 1410 2900 1430
rect 2920 1410 2940 1430
rect 2960 1410 2980 1430
rect 3000 1410 3020 1430
rect 3040 1410 3060 1430
rect 3080 1410 3100 1430
rect 3120 1410 3140 1430
rect 3160 1410 3170 1430
rect 2770 1385 3170 1410
rect 3290 1430 3690 1440
rect 3290 1410 3300 1430
rect 3320 1410 3340 1430
rect 3360 1410 3380 1430
rect 3400 1410 3420 1430
rect 3440 1410 3460 1430
rect 3480 1410 3500 1430
rect 3520 1410 3540 1430
rect 3560 1410 3580 1430
rect 3600 1410 3620 1430
rect 3640 1410 3660 1430
rect 3680 1410 3690 1430
rect 3290 1385 3690 1410
rect 2770 970 3170 985
rect 3290 970 3690 985
rect 2720 900 2760 910
rect 2720 880 2730 900
rect 2750 880 2760 900
rect 2720 870 2760 880
rect 2800 900 2840 910
rect 2800 880 2810 900
rect 2830 880 2840 900
rect 2800 870 2840 880
rect 2880 900 2920 910
rect 2880 880 2890 900
rect 2910 880 2920 900
rect 2880 870 2920 880
rect 2960 900 3000 910
rect 2960 880 2970 900
rect 2990 880 3000 900
rect 2960 870 3000 880
rect 3040 900 3080 910
rect 3040 880 3050 900
rect 3070 880 3080 900
rect 3040 870 3080 880
rect 3120 900 3160 910
rect 3120 880 3130 900
rect 3150 880 3160 900
rect 3120 870 3160 880
rect 3200 900 3240 910
rect 3200 880 3210 900
rect 3230 880 3240 900
rect 3200 870 3240 880
rect 3280 900 3320 910
rect 3280 880 3290 900
rect 3310 880 3320 900
rect 3280 870 3320 880
rect 3360 900 3400 910
rect 3360 880 3370 900
rect 3390 880 3400 900
rect 3360 870 3400 880
rect 3440 900 3480 910
rect 3440 880 3450 900
rect 3470 880 3480 900
rect 3440 870 3480 880
rect 3520 900 3560 910
rect 3520 880 3530 900
rect 3550 880 3560 900
rect 3520 870 3560 880
rect 3600 900 3640 910
rect 3600 880 3610 900
rect 3630 880 3640 900
rect 3600 870 3640 880
rect 3680 900 3720 910
rect 3680 880 3690 900
rect 3710 880 3720 900
rect 3680 870 3720 880
rect 2720 855 3720 870
rect 2720 740 3720 755
<< polycont >>
rect 4525 2175 4545 2195
rect 2920 1865 2940 1885
rect 3520 1865 3540 1885
rect 4495 1850 4515 1870
rect 3175 1820 3195 1840
rect 3060 1685 3080 1705
rect 3380 1685 3400 1705
rect 2920 1515 2940 1535
rect 3520 1515 3540 1535
rect 2780 1410 2800 1430
rect 2820 1410 2840 1430
rect 2860 1410 2880 1430
rect 2900 1410 2920 1430
rect 2940 1410 2960 1430
rect 2980 1410 3000 1430
rect 3020 1410 3040 1430
rect 3060 1410 3080 1430
rect 3100 1410 3120 1430
rect 3140 1410 3160 1430
rect 3300 1410 3320 1430
rect 3340 1410 3360 1430
rect 3380 1410 3400 1430
rect 3420 1410 3440 1430
rect 3460 1410 3480 1430
rect 3500 1410 3520 1430
rect 3540 1410 3560 1430
rect 3580 1410 3600 1430
rect 3620 1410 3640 1430
rect 3660 1410 3680 1430
rect 2730 880 2750 900
rect 2810 880 2830 900
rect 2890 880 2910 900
rect 2970 880 2990 900
rect 3050 880 3070 900
rect 3130 880 3150 900
rect 3210 880 3230 900
rect 3290 880 3310 900
rect 3370 880 3390 900
rect 3450 880 3470 900
rect 3530 880 3550 900
rect 3610 880 3630 900
rect 3690 880 3710 900
<< xpolycontact >>
rect 1005 2490 1225 2525
rect 1895 2490 2115 2525
rect 1005 2430 1225 2465
rect 1895 2430 2115 2465
rect 1005 2370 1225 2405
rect 1895 2370 2115 2405
rect 1005 2310 1225 2345
rect 1895 2310 2115 2345
rect 1005 2250 1225 2285
rect 1895 2250 2115 2285
rect 1005 1980 1225 2015
rect 1895 1980 2115 2015
rect 1005 1920 1225 1955
rect 1895 1920 2115 1955
rect 1005 1860 1225 1895
rect 1895 1860 2115 1895
rect 1005 1800 1225 1835
rect 1895 1800 2115 1835
rect 1005 1740 1225 1775
rect 1895 1740 2115 1775
rect 1005 1505 1225 1540
rect 1575 1505 1795 1540
rect 1005 1445 1225 1480
rect 1895 1445 2115 1480
rect 1005 1385 1225 1420
rect 1895 1385 2115 1420
rect 1005 1325 1225 1360
rect 1895 1325 2115 1360
rect 1005 1265 1225 1300
rect 1895 1265 2115 1300
rect 1005 1205 1225 1240
rect 1895 1205 2115 1240
<< xpolyres >>
rect 1225 2490 1895 2525
rect 1225 2430 1895 2465
rect 1225 2370 1895 2405
rect 1225 2310 1895 2345
rect 1225 2250 1895 2285
rect 1225 1980 1895 2015
rect 1225 1920 1895 1955
rect 1225 1860 1895 1895
rect 1225 1800 1895 1835
rect 1225 1740 1895 1775
rect 1225 1505 1575 1540
rect 1225 1445 1895 1480
rect 1225 1385 1895 1420
rect 1225 1325 1895 1360
rect 1225 1265 1895 1300
rect 1225 1205 1895 1240
<< locali >>
rect 2610 2775 2650 2785
rect 2610 2755 2620 2775
rect 2640 2755 2650 2775
rect 2610 2745 2650 2755
rect 2810 2775 2850 2785
rect 2810 2755 2820 2775
rect 2840 2755 2850 2775
rect 2810 2745 2850 2755
rect 3010 2775 3050 2785
rect 3010 2755 3020 2775
rect 3040 2755 3050 2775
rect 3010 2745 3050 2755
rect 3210 2775 3250 2785
rect 3210 2755 3220 2775
rect 3240 2755 3250 2775
rect 3210 2745 3250 2755
rect 3410 2775 3450 2785
rect 3410 2755 3420 2775
rect 3440 2755 3450 2775
rect 3410 2745 3450 2755
rect 3610 2775 3650 2785
rect 3610 2755 3620 2775
rect 3640 2755 3650 2775
rect 3610 2745 3650 2755
rect 3810 2775 3850 2785
rect 3810 2755 3820 2775
rect 3840 2755 3850 2775
rect 3810 2745 3850 2755
rect 2620 2725 2640 2745
rect 2820 2725 2840 2745
rect 3020 2725 3040 2745
rect 2575 2715 2645 2725
rect 2575 2695 2580 2715
rect 2600 2695 2620 2715
rect 2640 2695 2645 2715
rect 2575 2665 2645 2695
rect 2575 2645 2580 2665
rect 2600 2645 2620 2665
rect 2640 2645 2645 2665
rect 2575 2615 2645 2645
rect 2575 2595 2580 2615
rect 2600 2595 2620 2615
rect 2640 2595 2645 2615
rect 2575 2565 2645 2595
rect 2575 2545 2580 2565
rect 2600 2545 2620 2565
rect 2640 2545 2645 2565
rect 945 2515 1005 2525
rect 945 2495 955 2515
rect 975 2495 1005 2515
rect 945 2490 1005 2495
rect 945 2485 985 2490
rect 1895 2465 2115 2490
rect 2575 2515 2645 2545
rect 2575 2495 2580 2515
rect 2600 2495 2620 2515
rect 2640 2495 2645 2515
rect 2575 2465 2645 2495
rect 2575 2445 2580 2465
rect 2600 2445 2620 2465
rect 2640 2445 2645 2465
rect 1005 2405 1225 2430
rect 2575 2415 2645 2445
rect 1895 2345 2115 2370
rect 2575 2395 2580 2415
rect 2600 2395 2620 2415
rect 2640 2395 2645 2415
rect 2575 2365 2645 2395
rect 2575 2345 2580 2365
rect 2600 2345 2620 2365
rect 2640 2345 2645 2365
rect 2575 2335 2645 2345
rect 2715 2715 2745 2725
rect 2715 2695 2720 2715
rect 2740 2695 2745 2715
rect 2715 2665 2745 2695
rect 2715 2645 2720 2665
rect 2740 2645 2745 2665
rect 2715 2615 2745 2645
rect 2715 2595 2720 2615
rect 2740 2595 2745 2615
rect 2715 2565 2745 2595
rect 2715 2545 2720 2565
rect 2740 2545 2745 2565
rect 2715 2515 2745 2545
rect 2715 2495 2720 2515
rect 2740 2495 2745 2515
rect 2715 2465 2745 2495
rect 2715 2445 2720 2465
rect 2740 2445 2745 2465
rect 2715 2415 2745 2445
rect 2715 2395 2720 2415
rect 2740 2395 2745 2415
rect 2715 2365 2745 2395
rect 2715 2345 2720 2365
rect 2740 2345 2745 2365
rect 2715 2335 2745 2345
rect 2815 2715 2845 2725
rect 2815 2695 2820 2715
rect 2840 2695 2845 2715
rect 2815 2665 2845 2695
rect 2815 2645 2820 2665
rect 2840 2645 2845 2665
rect 2815 2615 2845 2645
rect 2815 2595 2820 2615
rect 2840 2595 2845 2615
rect 2815 2565 2845 2595
rect 2815 2545 2820 2565
rect 2840 2545 2845 2565
rect 2815 2515 2845 2545
rect 2815 2495 2820 2515
rect 2840 2495 2845 2515
rect 2815 2465 2845 2495
rect 2815 2445 2820 2465
rect 2840 2445 2845 2465
rect 2815 2415 2845 2445
rect 2815 2395 2820 2415
rect 2840 2395 2845 2415
rect 2815 2365 2845 2395
rect 2815 2345 2820 2365
rect 2840 2345 2845 2365
rect 2815 2335 2845 2345
rect 2915 2715 2945 2725
rect 2915 2695 2920 2715
rect 2940 2695 2945 2715
rect 2915 2665 2945 2695
rect 2915 2645 2920 2665
rect 2940 2645 2945 2665
rect 2915 2615 2945 2645
rect 2915 2595 2920 2615
rect 2940 2595 2945 2615
rect 2915 2565 2945 2595
rect 2915 2545 2920 2565
rect 2940 2545 2945 2565
rect 2915 2515 2945 2545
rect 2915 2495 2920 2515
rect 2940 2495 2945 2515
rect 2915 2465 2945 2495
rect 2915 2445 2920 2465
rect 2940 2445 2945 2465
rect 2915 2415 2945 2445
rect 2915 2395 2920 2415
rect 2940 2395 2945 2415
rect 2915 2365 2945 2395
rect 2915 2345 2920 2365
rect 2940 2345 2945 2365
rect 2915 2335 2945 2345
rect 3015 2715 3045 2725
rect 3015 2695 3020 2715
rect 3040 2695 3045 2715
rect 3015 2665 3045 2695
rect 3015 2645 3020 2665
rect 3040 2645 3045 2665
rect 3015 2615 3045 2645
rect 3015 2595 3020 2615
rect 3040 2595 3045 2615
rect 3015 2565 3045 2595
rect 3015 2545 3020 2565
rect 3040 2545 3045 2565
rect 3015 2515 3045 2545
rect 3015 2495 3020 2515
rect 3040 2495 3045 2515
rect 3015 2465 3045 2495
rect 3015 2445 3020 2465
rect 3040 2445 3045 2465
rect 3015 2415 3045 2445
rect 3015 2395 3020 2415
rect 3040 2395 3045 2415
rect 3015 2365 3045 2395
rect 3015 2345 3020 2365
rect 3040 2345 3045 2365
rect 3015 2335 3045 2345
rect 3115 2715 3145 2725
rect 3115 2695 3120 2715
rect 3140 2695 3145 2715
rect 3115 2665 3145 2695
rect 3115 2645 3120 2665
rect 3140 2645 3145 2665
rect 3115 2615 3145 2645
rect 3115 2595 3120 2615
rect 3140 2595 3145 2615
rect 3115 2565 3145 2595
rect 3115 2545 3120 2565
rect 3140 2545 3145 2565
rect 3115 2515 3145 2545
rect 3115 2495 3120 2515
rect 3140 2495 3145 2515
rect 3115 2465 3145 2495
rect 3115 2445 3120 2465
rect 3140 2445 3145 2465
rect 3115 2415 3145 2445
rect 3115 2395 3120 2415
rect 3140 2395 3145 2415
rect 3115 2365 3145 2395
rect 3115 2345 3120 2365
rect 3140 2345 3145 2365
rect 3115 2335 3145 2345
rect 3215 2715 3245 2745
rect 3420 2725 3440 2745
rect 3620 2725 3640 2745
rect 3820 2725 3840 2745
rect 3215 2695 3220 2715
rect 3240 2695 3245 2715
rect 3215 2665 3245 2695
rect 3215 2645 3220 2665
rect 3240 2645 3245 2665
rect 3215 2615 3245 2645
rect 3215 2595 3220 2615
rect 3240 2595 3245 2615
rect 3215 2565 3245 2595
rect 3215 2545 3220 2565
rect 3240 2545 3245 2565
rect 3215 2515 3245 2545
rect 3215 2495 3220 2515
rect 3240 2495 3245 2515
rect 3215 2465 3245 2495
rect 3215 2445 3220 2465
rect 3240 2445 3245 2465
rect 3215 2415 3245 2445
rect 3215 2395 3220 2415
rect 3240 2395 3245 2415
rect 3215 2365 3245 2395
rect 3215 2345 3220 2365
rect 3240 2345 3245 2365
rect 3215 2335 3245 2345
rect 3315 2715 3345 2725
rect 3315 2695 3320 2715
rect 3340 2695 3345 2715
rect 3315 2665 3345 2695
rect 3315 2645 3320 2665
rect 3340 2645 3345 2665
rect 3315 2615 3345 2645
rect 3315 2595 3320 2615
rect 3340 2595 3345 2615
rect 3315 2565 3345 2595
rect 3315 2545 3320 2565
rect 3340 2545 3345 2565
rect 3315 2515 3345 2545
rect 3315 2495 3320 2515
rect 3340 2495 3345 2515
rect 3315 2465 3345 2495
rect 3315 2445 3320 2465
rect 3340 2445 3345 2465
rect 3315 2415 3345 2445
rect 3315 2395 3320 2415
rect 3340 2395 3345 2415
rect 3315 2365 3345 2395
rect 3315 2345 3320 2365
rect 3340 2345 3345 2365
rect 3315 2335 3345 2345
rect 3415 2715 3445 2725
rect 3415 2695 3420 2715
rect 3440 2695 3445 2715
rect 3415 2665 3445 2695
rect 3415 2645 3420 2665
rect 3440 2645 3445 2665
rect 3415 2615 3445 2645
rect 3415 2595 3420 2615
rect 3440 2595 3445 2615
rect 3415 2565 3445 2595
rect 3415 2545 3420 2565
rect 3440 2545 3445 2565
rect 3415 2515 3445 2545
rect 3415 2495 3420 2515
rect 3440 2495 3445 2515
rect 3415 2465 3445 2495
rect 3415 2445 3420 2465
rect 3440 2445 3445 2465
rect 3415 2415 3445 2445
rect 3415 2395 3420 2415
rect 3440 2395 3445 2415
rect 3415 2365 3445 2395
rect 3415 2345 3420 2365
rect 3440 2345 3445 2365
rect 3415 2335 3445 2345
rect 3515 2715 3545 2725
rect 3515 2695 3520 2715
rect 3540 2695 3545 2715
rect 3515 2665 3545 2695
rect 3515 2645 3520 2665
rect 3540 2645 3545 2665
rect 3515 2615 3545 2645
rect 3515 2595 3520 2615
rect 3540 2595 3545 2615
rect 3515 2565 3545 2595
rect 3515 2545 3520 2565
rect 3540 2545 3545 2565
rect 3515 2515 3545 2545
rect 3515 2495 3520 2515
rect 3540 2495 3545 2515
rect 3515 2465 3545 2495
rect 3515 2445 3520 2465
rect 3540 2445 3545 2465
rect 3515 2415 3545 2445
rect 3515 2395 3520 2415
rect 3540 2395 3545 2415
rect 3515 2365 3545 2395
rect 3515 2345 3520 2365
rect 3540 2345 3545 2365
rect 3515 2335 3545 2345
rect 3615 2715 3645 2725
rect 3615 2695 3620 2715
rect 3640 2695 3645 2715
rect 3615 2665 3645 2695
rect 3615 2645 3620 2665
rect 3640 2645 3645 2665
rect 3615 2615 3645 2645
rect 3615 2595 3620 2615
rect 3640 2595 3645 2615
rect 3615 2565 3645 2595
rect 3615 2545 3620 2565
rect 3640 2545 3645 2565
rect 3615 2515 3645 2545
rect 3615 2495 3620 2515
rect 3640 2495 3645 2515
rect 3615 2465 3645 2495
rect 3615 2445 3620 2465
rect 3640 2445 3645 2465
rect 3615 2415 3645 2445
rect 3615 2395 3620 2415
rect 3640 2395 3645 2415
rect 3615 2365 3645 2395
rect 3615 2345 3620 2365
rect 3640 2345 3645 2365
rect 3615 2335 3645 2345
rect 3715 2715 3745 2725
rect 3715 2695 3720 2715
rect 3740 2695 3745 2715
rect 3715 2665 3745 2695
rect 3715 2645 3720 2665
rect 3740 2645 3745 2665
rect 3715 2615 3745 2645
rect 3715 2595 3720 2615
rect 3740 2595 3745 2615
rect 3715 2565 3745 2595
rect 3715 2545 3720 2565
rect 3740 2545 3745 2565
rect 3715 2515 3745 2545
rect 3715 2495 3720 2515
rect 3740 2495 3745 2515
rect 3715 2465 3745 2495
rect 3715 2445 3720 2465
rect 3740 2445 3745 2465
rect 3715 2415 3745 2445
rect 3715 2395 3720 2415
rect 3740 2395 3745 2415
rect 3715 2365 3745 2395
rect 3715 2345 3720 2365
rect 3740 2345 3745 2365
rect 3715 2335 3745 2345
rect 3815 2715 3885 2725
rect 3815 2695 3820 2715
rect 3840 2695 3860 2715
rect 3880 2695 3885 2715
rect 3815 2665 3885 2695
rect 3815 2645 3820 2665
rect 3840 2645 3860 2665
rect 3880 2645 3885 2665
rect 3815 2615 3885 2645
rect 3815 2595 3820 2615
rect 3840 2595 3860 2615
rect 3880 2595 3885 2615
rect 3815 2565 3885 2595
rect 3815 2545 3820 2565
rect 3840 2545 3860 2565
rect 3880 2545 3885 2565
rect 3815 2515 3885 2545
rect 3815 2495 3820 2515
rect 3840 2495 3860 2515
rect 3880 2495 3885 2515
rect 3815 2465 3885 2495
rect 3815 2445 3820 2465
rect 3840 2445 3860 2465
rect 3880 2445 3885 2465
rect 3815 2415 3885 2445
rect 3815 2395 3820 2415
rect 3840 2395 3860 2415
rect 3880 2395 3885 2415
rect 3815 2365 3885 2395
rect 3815 2345 3820 2365
rect 3840 2345 3860 2365
rect 3880 2345 3885 2365
rect 3815 2335 3885 2345
rect 2720 2315 2740 2335
rect 1005 2285 1225 2310
rect 2710 2305 2750 2315
rect 2710 2285 2720 2305
rect 2740 2285 2750 2305
rect 2710 2275 2750 2285
rect 2920 2270 2940 2335
rect 1895 2220 2115 2250
rect 2910 2260 2950 2270
rect 2910 2240 2920 2260
rect 2940 2240 2950 2260
rect 2910 2230 2950 2240
rect 3120 2225 3140 2335
rect 3320 2225 3340 2335
rect 3520 2270 3540 2335
rect 3720 2315 3740 2335
rect 3710 2305 3750 2315
rect 3710 2285 3720 2305
rect 3740 2285 3750 2305
rect 3710 2275 3750 2285
rect 3510 2260 3550 2270
rect 3510 2240 3520 2260
rect 3540 2240 3550 2260
rect 3510 2230 3550 2240
rect 1895 2200 1905 2220
rect 1925 2200 1950 2220
rect 1970 2200 1995 2220
rect 2015 2200 2040 2220
rect 2060 2200 2085 2220
rect 2105 2200 2115 2220
rect 1895 2190 2115 2200
rect 3110 2215 3150 2225
rect 3110 2195 3120 2215
rect 3140 2195 3150 2215
rect 3110 2185 3150 2195
rect 3310 2215 3350 2225
rect 3310 2195 3320 2215
rect 3340 2195 3350 2215
rect 3310 2185 3350 2195
rect 4375 2205 4415 2210
rect 4375 2185 4385 2205
rect 4405 2195 4555 2205
rect 4405 2185 4525 2195
rect 4375 2175 4415 2185
rect 4515 2175 4525 2185
rect 4545 2175 4555 2195
rect 2610 2155 2650 2165
rect 2610 2135 2620 2155
rect 2640 2135 2650 2155
rect 2610 2125 2650 2135
rect 2810 2155 2850 2165
rect 2810 2135 2820 2155
rect 2840 2135 2850 2155
rect 2810 2125 2850 2135
rect 3010 2155 3050 2165
rect 3010 2135 3020 2155
rect 3040 2135 3050 2155
rect 3010 2125 3050 2135
rect 3110 2155 3150 2165
rect 3110 2135 3120 2155
rect 3140 2135 3150 2155
rect 3110 2125 3150 2135
rect 3210 2155 3250 2165
rect 3210 2135 3220 2155
rect 3240 2135 3250 2155
rect 3210 2125 3250 2135
rect 3310 2155 3350 2165
rect 3310 2135 3320 2155
rect 3340 2135 3350 2155
rect 3310 2125 3350 2135
rect 3410 2155 3450 2165
rect 3410 2135 3420 2155
rect 3440 2135 3450 2155
rect 3410 2125 3450 2135
rect 3610 2155 3650 2165
rect 3610 2135 3620 2155
rect 3640 2135 3650 2155
rect 3610 2125 3650 2135
rect 3810 2155 3850 2165
rect 3810 2135 3820 2155
rect 3840 2135 3850 2155
rect 3810 2125 3850 2135
rect 2620 2105 2640 2125
rect 2820 2105 2840 2125
rect 3020 2105 3040 2125
rect 3120 2105 3140 2125
rect 3220 2105 3240 2125
rect 3320 2105 3340 2125
rect 3420 2105 3440 2125
rect 3620 2105 3640 2125
rect 3820 2105 3840 2125
rect 4385 2105 4405 2175
rect 4515 2165 4555 2175
rect 4585 2155 4625 2165
rect 4585 2135 4595 2155
rect 4615 2135 4625 2155
rect 4585 2125 4625 2135
rect 4595 2105 4615 2125
rect 2575 2095 2645 2105
rect 2575 2075 2580 2095
rect 2600 2075 2620 2095
rect 2640 2075 2645 2095
rect 2575 2045 2645 2075
rect 2575 2025 2580 2045
rect 2600 2025 2620 2045
rect 2640 2025 2645 2045
rect 945 2005 1005 2015
rect 945 1985 955 2005
rect 975 1985 1005 2005
rect 945 1980 1005 1985
rect 945 1975 985 1980
rect 1895 1955 2115 1980
rect 2575 1995 2645 2025
rect 2575 1975 2580 1995
rect 2600 1975 2620 1995
rect 2640 1975 2645 1995
rect 2575 1945 2645 1975
rect 2575 1925 2580 1945
rect 2600 1925 2620 1945
rect 2640 1925 2645 1945
rect 1005 1895 1225 1920
rect 2575 1915 2645 1925
rect 2715 2095 2745 2105
rect 2715 2075 2720 2095
rect 2740 2075 2745 2095
rect 2715 2045 2745 2075
rect 2715 2025 2720 2045
rect 2740 2025 2745 2045
rect 2715 1995 2745 2025
rect 2715 1975 2720 1995
rect 2740 1975 2745 1995
rect 2715 1945 2745 1975
rect 2715 1925 2720 1945
rect 2740 1925 2745 1945
rect 2715 1915 2745 1925
rect 2815 2095 2845 2105
rect 2815 2075 2820 2095
rect 2840 2075 2845 2095
rect 2815 2045 2845 2075
rect 2815 2025 2820 2045
rect 2840 2025 2845 2045
rect 2815 1995 2845 2025
rect 2815 1975 2820 1995
rect 2840 1975 2845 1995
rect 2815 1945 2845 1975
rect 2815 1925 2820 1945
rect 2840 1925 2845 1945
rect 2815 1915 2845 1925
rect 2915 2095 2945 2105
rect 2915 2075 2920 2095
rect 2940 2075 2945 2095
rect 2915 2045 2945 2075
rect 2915 2025 2920 2045
rect 2940 2025 2945 2045
rect 2915 1995 2945 2025
rect 2915 1975 2920 1995
rect 2940 1975 2945 1995
rect 2915 1945 2945 1975
rect 2915 1925 2920 1945
rect 2940 1925 2945 1945
rect 2915 1915 2945 1925
rect 3015 2095 3045 2105
rect 3015 2075 3020 2095
rect 3040 2075 3045 2095
rect 3015 2045 3045 2075
rect 3015 2025 3020 2045
rect 3040 2025 3045 2045
rect 3015 1995 3045 2025
rect 3015 1975 3020 1995
rect 3040 1975 3045 1995
rect 3015 1945 3045 1975
rect 3015 1925 3020 1945
rect 3040 1925 3045 1945
rect 3015 1915 3045 1925
rect 3115 2095 3145 2105
rect 3115 2075 3120 2095
rect 3140 2075 3145 2095
rect 3115 2045 3145 2075
rect 3115 2025 3120 2045
rect 3140 2025 3145 2045
rect 3115 1995 3145 2025
rect 3115 1975 3120 1995
rect 3140 1975 3145 1995
rect 3115 1945 3145 1975
rect 3115 1925 3120 1945
rect 3140 1925 3145 1945
rect 3115 1915 3145 1925
rect 3215 2095 3245 2105
rect 3215 2075 3220 2095
rect 3240 2075 3245 2095
rect 3215 2045 3245 2075
rect 3215 2025 3220 2045
rect 3240 2025 3245 2045
rect 3215 1995 3245 2025
rect 3215 1975 3220 1995
rect 3240 1975 3245 1995
rect 3215 1945 3245 1975
rect 3215 1925 3220 1945
rect 3240 1925 3245 1945
rect 3215 1915 3245 1925
rect 3315 2095 3345 2105
rect 3315 2075 3320 2095
rect 3340 2075 3345 2095
rect 3315 2045 3345 2075
rect 3315 2025 3320 2045
rect 3340 2025 3345 2045
rect 3315 1995 3345 2025
rect 3315 1975 3320 1995
rect 3340 1975 3345 1995
rect 3315 1945 3345 1975
rect 3315 1925 3320 1945
rect 3340 1925 3345 1945
rect 3315 1915 3345 1925
rect 3415 2095 3445 2105
rect 3415 2075 3420 2095
rect 3440 2075 3445 2095
rect 3415 2045 3445 2075
rect 3415 2025 3420 2045
rect 3440 2025 3445 2045
rect 3415 1995 3445 2025
rect 3415 1975 3420 1995
rect 3440 1975 3445 1995
rect 3415 1945 3445 1975
rect 3415 1925 3420 1945
rect 3440 1925 3445 1945
rect 3415 1915 3445 1925
rect 3515 2095 3545 2105
rect 3515 2075 3520 2095
rect 3540 2075 3545 2095
rect 3515 2045 3545 2075
rect 3515 2025 3520 2045
rect 3540 2025 3545 2045
rect 3515 1995 3545 2025
rect 3515 1975 3520 1995
rect 3540 1975 3545 1995
rect 3515 1945 3545 1975
rect 3515 1925 3520 1945
rect 3540 1925 3545 1945
rect 3515 1915 3545 1925
rect 3615 2095 3645 2105
rect 3615 2075 3620 2095
rect 3640 2075 3645 2095
rect 3615 2045 3645 2075
rect 3615 2025 3620 2045
rect 3640 2025 3645 2045
rect 3615 1995 3645 2025
rect 3615 1975 3620 1995
rect 3640 1975 3645 1995
rect 3615 1945 3645 1975
rect 3615 1925 3620 1945
rect 3640 1925 3645 1945
rect 3615 1915 3645 1925
rect 3715 2095 3745 2105
rect 3715 2075 3720 2095
rect 3740 2075 3745 2095
rect 3715 2045 3745 2075
rect 3715 2025 3720 2045
rect 3740 2025 3745 2045
rect 3715 1995 3745 2025
rect 3715 1975 3720 1995
rect 3740 1975 3745 1995
rect 3715 1945 3745 1975
rect 3715 1925 3720 1945
rect 3740 1925 3745 1945
rect 3715 1915 3745 1925
rect 3815 2095 3885 2105
rect 3815 2075 3820 2095
rect 3840 2075 3860 2095
rect 3880 2075 3885 2095
rect 3815 2045 3885 2075
rect 3815 2025 3820 2045
rect 3840 2025 3860 2045
rect 3880 2025 3885 2045
rect 3815 1995 3885 2025
rect 3815 1975 3820 1995
rect 3840 1975 3860 1995
rect 3880 1975 3885 1995
rect 3815 1945 3885 1975
rect 3815 1925 3820 1945
rect 3840 1925 3860 1945
rect 3880 1925 3885 1945
rect 3815 1915 3885 1925
rect 4380 2095 4410 2105
rect 4380 2075 4385 2095
rect 4405 2075 4410 2095
rect 4380 2045 4410 2075
rect 4380 2025 4385 2045
rect 4405 2025 4410 2045
rect 4380 1995 4410 2025
rect 4380 1975 4385 1995
rect 4405 1975 4410 1995
rect 4380 1945 4410 1975
rect 4380 1925 4385 1945
rect 4405 1925 4410 1945
rect 4380 1915 4410 1925
rect 4435 2095 4465 2105
rect 4435 2075 4440 2095
rect 4460 2075 4465 2095
rect 4435 2045 4465 2075
rect 4435 2025 4440 2045
rect 4460 2025 4465 2045
rect 4435 1995 4465 2025
rect 4435 1975 4440 1995
rect 4460 1975 4465 1995
rect 4435 1945 4465 1975
rect 4435 1925 4440 1945
rect 4460 1925 4465 1945
rect 4435 1915 4465 1925
rect 4505 2095 4535 2105
rect 4505 2075 4510 2095
rect 4530 2075 4535 2095
rect 4505 2045 4535 2075
rect 4505 2025 4510 2045
rect 4530 2025 4535 2045
rect 4505 1995 4535 2025
rect 4505 1975 4510 1995
rect 4530 1975 4535 1995
rect 4505 1945 4535 1975
rect 4505 1925 4510 1945
rect 4530 1925 4535 1945
rect 4505 1915 4535 1925
rect 4560 2095 4615 2105
rect 4560 2075 4565 2095
rect 4585 2075 4615 2095
rect 4560 2045 4595 2075
rect 4560 2025 4565 2045
rect 4585 2025 4595 2045
rect 4560 1995 4595 2025
rect 4560 1975 4565 1995
rect 4585 1975 4595 1995
rect 4560 1945 4595 1975
rect 4560 1925 4565 1945
rect 4585 1925 4595 1945
rect 4560 1915 4595 1925
rect 1895 1835 2115 1860
rect 2720 1850 2740 1915
rect 2920 1895 2940 1915
rect 3120 1895 3140 1915
rect 3320 1895 3340 1915
rect 3520 1895 3540 1915
rect 2910 1885 2950 1895
rect 2910 1865 2920 1885
rect 2940 1865 2950 1885
rect 3120 1885 3340 1895
rect 3120 1875 3240 1885
rect 2910 1855 2950 1865
rect 3230 1865 3240 1875
rect 3260 1875 3340 1885
rect 3510 1885 3550 1895
rect 3260 1865 3270 1875
rect 3230 1855 3270 1865
rect 3510 1865 3520 1885
rect 3540 1865 3550 1885
rect 3510 1855 3550 1865
rect 3720 1850 3740 1915
rect 2710 1840 2750 1850
rect 2710 1820 2720 1840
rect 2740 1820 2750 1840
rect 2710 1810 2750 1820
rect 3165 1840 3205 1850
rect 3165 1820 3175 1840
rect 3195 1820 3205 1840
rect 3165 1810 3205 1820
rect 3710 1840 3750 1850
rect 3710 1820 3720 1840
rect 3740 1820 3750 1840
rect 3710 1810 3750 1820
rect 1005 1775 1225 1800
rect 3230 1795 3270 1805
rect 3230 1775 3240 1795
rect 3260 1775 3270 1795
rect 3230 1765 3270 1775
rect 1895 1710 2115 1740
rect 2910 1750 2950 1760
rect 2910 1730 2920 1750
rect 2940 1730 2950 1750
rect 2910 1720 2950 1730
rect 3510 1750 3550 1760
rect 3510 1730 3520 1750
rect 3540 1730 3550 1750
rect 3510 1720 3550 1730
rect 1895 1690 1905 1710
rect 1925 1690 1950 1710
rect 1970 1690 1995 1710
rect 2015 1690 2040 1710
rect 2060 1690 2085 1710
rect 2105 1690 2115 1710
rect 1895 1680 2115 1690
rect 2920 1655 2940 1720
rect 3050 1705 3090 1715
rect 3050 1685 3060 1705
rect 3080 1685 3090 1705
rect 3050 1675 3090 1685
rect 3110 1705 3150 1715
rect 3110 1685 3120 1705
rect 3140 1685 3150 1705
rect 3110 1675 3150 1685
rect 3310 1705 3350 1715
rect 3310 1685 3320 1705
rect 3340 1685 3350 1705
rect 3310 1675 3350 1685
rect 3370 1705 3410 1715
rect 3370 1685 3380 1705
rect 3400 1685 3410 1705
rect 3370 1675 3410 1685
rect 3120 1655 3140 1675
rect 3320 1655 3340 1675
rect 3520 1655 3540 1720
rect 4440 1715 4460 1915
rect 4505 1880 4525 1915
rect 4485 1870 4525 1880
rect 4485 1850 4495 1870
rect 4515 1850 4525 1870
rect 4485 1840 4525 1850
rect 4430 1705 4470 1715
rect 4430 1685 4440 1705
rect 4460 1685 4470 1705
rect 4430 1675 4470 1685
rect 2810 1645 2845 1655
rect 2810 1625 2820 1645
rect 2840 1625 2845 1645
rect 2810 1595 2845 1625
rect 2810 1575 2820 1595
rect 2840 1575 2845 1595
rect 2810 1565 2845 1575
rect 2915 1645 2945 1655
rect 2915 1625 2920 1645
rect 2940 1625 2945 1645
rect 2915 1595 2945 1625
rect 2915 1575 2920 1595
rect 2940 1575 2945 1595
rect 2915 1565 2945 1575
rect 3015 1645 3045 1655
rect 3015 1625 3020 1645
rect 3040 1625 3045 1645
rect 3015 1595 3045 1625
rect 3015 1575 3020 1595
rect 3040 1575 3045 1595
rect 3015 1565 3045 1575
rect 3115 1645 3145 1655
rect 3115 1625 3120 1645
rect 3140 1625 3145 1645
rect 3115 1595 3145 1625
rect 3115 1575 3120 1595
rect 3140 1575 3145 1595
rect 3115 1565 3145 1575
rect 3215 1645 3245 1655
rect 3215 1625 3220 1645
rect 3240 1625 3245 1645
rect 3215 1595 3245 1625
rect 3215 1575 3220 1595
rect 3240 1575 3245 1595
rect 3215 1565 3245 1575
rect 3315 1645 3345 1655
rect 3315 1625 3320 1645
rect 3340 1625 3345 1645
rect 3315 1595 3345 1625
rect 3315 1575 3320 1595
rect 3340 1575 3345 1595
rect 3315 1565 3345 1575
rect 3415 1645 3445 1655
rect 3415 1625 3420 1645
rect 3440 1625 3445 1645
rect 3415 1595 3445 1625
rect 3415 1575 3420 1595
rect 3440 1575 3445 1595
rect 3415 1565 3445 1575
rect 3515 1645 3545 1655
rect 3515 1625 3520 1645
rect 3540 1625 3545 1645
rect 3515 1595 3545 1625
rect 3515 1575 3520 1595
rect 3540 1575 3545 1595
rect 3515 1565 3545 1575
rect 3615 1645 3650 1655
rect 3615 1625 3620 1645
rect 3640 1625 3650 1645
rect 3615 1595 3650 1625
rect 3615 1575 3620 1595
rect 3640 1575 3650 1595
rect 3615 1565 3650 1575
rect 945 1530 1005 1540
rect 945 1510 955 1530
rect 975 1510 1005 1530
rect 945 1505 1005 1510
rect 1795 1530 2115 1540
rect 1795 1510 1905 1530
rect 1925 1510 1950 1530
rect 1970 1510 1995 1530
rect 2015 1510 2040 1530
rect 2060 1510 2085 1530
rect 2105 1510 2115 1530
rect 1795 1505 2115 1510
rect 945 1500 985 1505
rect 1895 1480 2115 1505
rect 2820 1500 2840 1565
rect 2910 1535 2950 1545
rect 2910 1515 2920 1535
rect 2940 1515 2950 1535
rect 2910 1505 2950 1515
rect 3020 1500 3040 1565
rect 3220 1500 3240 1565
rect 3420 1500 3440 1565
rect 3510 1535 3550 1545
rect 3510 1515 3520 1535
rect 3540 1515 3550 1535
rect 3510 1505 3550 1515
rect 3620 1500 3640 1565
rect 2810 1490 2850 1500
rect 2810 1470 2820 1490
rect 2840 1470 2850 1490
rect 2810 1460 2850 1470
rect 3010 1490 3050 1500
rect 3010 1470 3020 1490
rect 3040 1470 3050 1490
rect 3010 1460 3050 1470
rect 3210 1490 3250 1500
rect 3210 1470 3220 1490
rect 3240 1470 3250 1490
rect 3210 1460 3250 1470
rect 3410 1490 3450 1500
rect 3410 1470 3420 1490
rect 3440 1470 3450 1490
rect 3410 1460 3450 1470
rect 3610 1490 3650 1500
rect 3610 1470 3620 1490
rect 3640 1470 3650 1490
rect 3610 1460 3650 1470
rect 1005 1420 1225 1445
rect 2820 1440 2840 1460
rect 3020 1440 3040 1460
rect 2735 1430 3170 1440
rect 1895 1360 2115 1385
rect 2735 1410 2780 1430
rect 2800 1410 2820 1430
rect 2840 1410 2860 1430
rect 2880 1410 2900 1430
rect 2920 1410 2940 1430
rect 2960 1410 2980 1430
rect 3000 1410 3020 1430
rect 3040 1410 3060 1430
rect 3080 1410 3100 1430
rect 3120 1410 3140 1430
rect 3160 1410 3170 1430
rect 2735 1400 3170 1410
rect 3290 1430 3730 1440
rect 3290 1410 3300 1430
rect 3320 1410 3340 1430
rect 3360 1410 3380 1430
rect 3400 1410 3420 1430
rect 3440 1410 3460 1430
rect 3480 1410 3500 1430
rect 3520 1410 3540 1430
rect 3560 1410 3580 1430
rect 3600 1410 3620 1430
rect 3640 1410 3660 1430
rect 3680 1410 3700 1430
rect 3720 1410 3730 1430
rect 3290 1400 3730 1410
rect 2735 1370 2765 1400
rect 2735 1350 2740 1370
rect 2760 1350 2765 1370
rect 1005 1300 1225 1325
rect 2735 1320 2765 1350
rect 2735 1300 2740 1320
rect 2760 1300 2765 1320
rect 945 1240 985 1245
rect 1895 1240 2115 1265
rect 945 1235 1005 1240
rect 945 1215 955 1235
rect 975 1215 1005 1235
rect 945 1205 1005 1215
rect 2735 1270 2765 1300
rect 2735 1250 2740 1270
rect 2760 1250 2765 1270
rect 2735 1220 2765 1250
rect 2735 1200 2740 1220
rect 2760 1200 2765 1220
rect 2735 1170 2765 1200
rect 2735 1150 2740 1170
rect 2760 1150 2765 1170
rect 2735 1120 2765 1150
rect 2735 1100 2740 1120
rect 2760 1100 2765 1120
rect 2735 1070 2765 1100
rect 2735 1050 2740 1070
rect 2760 1050 2765 1070
rect 2735 1020 2765 1050
rect 2735 1000 2740 1020
rect 2760 1000 2765 1020
rect 2735 990 2765 1000
rect 3175 1370 3285 1380
rect 3175 1350 3180 1370
rect 3200 1350 3220 1370
rect 3240 1350 3260 1370
rect 3280 1350 3285 1370
rect 3175 1320 3285 1350
rect 3175 1300 3180 1320
rect 3200 1300 3220 1320
rect 3240 1300 3260 1320
rect 3280 1300 3285 1320
rect 3175 1270 3285 1300
rect 3175 1250 3180 1270
rect 3200 1250 3220 1270
rect 3240 1250 3260 1270
rect 3280 1250 3285 1270
rect 3175 1220 3285 1250
rect 3175 1200 3180 1220
rect 3200 1200 3220 1220
rect 3240 1200 3260 1220
rect 3280 1200 3285 1220
rect 3175 1170 3285 1200
rect 3175 1150 3180 1170
rect 3200 1150 3220 1170
rect 3240 1150 3260 1170
rect 3280 1150 3285 1170
rect 3175 1120 3285 1150
rect 3175 1100 3180 1120
rect 3200 1100 3220 1120
rect 3240 1100 3260 1120
rect 3280 1100 3285 1120
rect 3175 1070 3285 1100
rect 3175 1050 3180 1070
rect 3200 1050 3220 1070
rect 3240 1050 3260 1070
rect 3280 1050 3285 1070
rect 3175 1020 3285 1050
rect 3175 1000 3180 1020
rect 3200 1000 3220 1020
rect 3240 1000 3260 1020
rect 3280 1000 3285 1020
rect 3175 990 3285 1000
rect 3695 1370 3725 1400
rect 3695 1350 3700 1370
rect 3720 1350 3725 1370
rect 3695 1320 3725 1350
rect 3695 1300 3700 1320
rect 3720 1300 3725 1320
rect 3695 1270 3725 1300
rect 3695 1250 3700 1270
rect 3720 1250 3725 1270
rect 3695 1220 3725 1250
rect 3695 1200 3700 1220
rect 3720 1200 3725 1220
rect 3695 1170 3725 1200
rect 3695 1150 3700 1170
rect 3720 1150 3725 1170
rect 3695 1120 3725 1150
rect 3695 1100 3700 1120
rect 3720 1100 3725 1120
rect 3695 1070 3725 1100
rect 3695 1050 3700 1070
rect 3720 1050 3725 1070
rect 3695 1020 3725 1050
rect 3695 1000 3700 1020
rect 3720 1000 3725 1020
rect 3695 990 3725 1000
rect 3180 970 3200 990
rect 3220 970 3240 990
rect 3260 970 3280 990
rect 3170 960 3290 970
rect 3170 940 3180 960
rect 3200 940 3220 960
rect 3240 940 3260 960
rect 3280 940 3290 960
rect 3170 930 3290 940
rect 2690 900 3760 910
rect 2690 880 2730 900
rect 2750 880 2810 900
rect 2830 880 2890 900
rect 2910 880 2970 900
rect 2990 880 3050 900
rect 3070 880 3130 900
rect 3150 880 3210 900
rect 3230 880 3290 900
rect 3310 880 3370 900
rect 3390 880 3450 900
rect 3470 880 3530 900
rect 3550 880 3610 900
rect 3630 880 3690 900
rect 3710 880 3730 900
rect 3750 880 3760 900
rect 2690 870 3760 880
rect 2690 850 2710 870
rect 2685 840 2715 850
rect 650 820 690 830
rect 650 800 660 820
rect 680 800 690 820
rect 650 770 690 800
rect 650 750 660 770
rect 680 750 690 770
rect 2685 820 2690 840
rect 2710 820 2715 840
rect 2685 790 2715 820
rect 2685 770 2690 790
rect 2710 770 2715 790
rect 2685 760 2715 770
rect 3725 840 3795 850
rect 3725 820 3730 840
rect 3750 820 3770 840
rect 3790 825 3795 840
rect 3790 820 3835 825
rect 3725 815 3835 820
rect 3725 795 3805 815
rect 3825 795 3835 815
rect 3725 790 3835 795
rect 3725 770 3730 790
rect 3750 770 3770 790
rect 3790 785 3835 790
rect 3790 770 3795 785
rect 3725 760 3795 770
rect 650 720 690 750
rect 650 700 660 720
rect 680 700 690 720
rect 650 660 690 700
rect 5 535 4740 660
rect 650 10 690 535
rect 1330 10 1370 535
rect 2010 10 2050 535
rect 2690 10 2730 535
rect 3370 10 3410 535
rect 4050 10 4090 535
<< viali >>
rect 2620 2755 2640 2775
rect 2820 2755 2840 2775
rect 3020 2755 3040 2775
rect 3220 2755 3240 2775
rect 3420 2755 3440 2775
rect 3620 2755 3640 2775
rect 3820 2755 3840 2775
rect 955 2495 975 2515
rect 2720 2285 2740 2305
rect 2920 2240 2940 2260
rect 3720 2285 3740 2305
rect 3520 2240 3540 2260
rect 1905 2200 1925 2220
rect 1950 2200 1970 2220
rect 1995 2200 2015 2220
rect 2040 2200 2060 2220
rect 2085 2200 2105 2220
rect 3120 2195 3140 2215
rect 3320 2195 3340 2215
rect 4385 2185 4405 2205
rect 2620 2135 2640 2155
rect 2820 2135 2840 2155
rect 3020 2135 3040 2155
rect 3120 2135 3140 2155
rect 3220 2135 3240 2155
rect 3320 2135 3340 2155
rect 3420 2135 3440 2155
rect 3620 2135 3640 2155
rect 3820 2135 3840 2155
rect 4595 2135 4615 2155
rect 955 1985 975 2005
rect 2920 1865 2940 1885
rect 3240 1865 3260 1885
rect 3520 1865 3540 1885
rect 2720 1820 2740 1840
rect 3175 1820 3195 1840
rect 3720 1820 3740 1840
rect 3240 1775 3260 1795
rect 2920 1730 2940 1750
rect 3520 1730 3540 1750
rect 1905 1690 1925 1710
rect 1950 1690 1970 1710
rect 1995 1690 2015 1710
rect 2040 1690 2060 1710
rect 2085 1690 2105 1710
rect 3060 1685 3080 1705
rect 3120 1685 3140 1705
rect 3320 1685 3340 1705
rect 3380 1685 3400 1705
rect 4495 1850 4515 1870
rect 4440 1685 4460 1705
rect 955 1510 975 1530
rect 1905 1510 1925 1530
rect 1950 1510 1970 1530
rect 1995 1510 2015 1530
rect 2040 1510 2060 1530
rect 2085 1510 2105 1530
rect 2920 1515 2940 1535
rect 3520 1515 3540 1535
rect 2820 1470 2840 1490
rect 3020 1470 3040 1490
rect 3220 1470 3240 1490
rect 3420 1470 3440 1490
rect 3620 1470 3640 1490
rect 3700 1410 3720 1430
rect 955 1215 975 1235
rect 3180 940 3200 960
rect 3220 940 3240 960
rect 3260 940 3280 960
rect 3730 880 3750 900
rect 660 800 680 820
rect 3805 795 3825 815
<< metal1 >>
rect 3220 2785 3240 3150
rect 2610 2780 2650 2785
rect 2610 2750 2615 2780
rect 2645 2750 2650 2780
rect 2610 2745 2650 2750
rect 2810 2780 2850 2785
rect 2810 2750 2815 2780
rect 2845 2750 2850 2780
rect 2810 2745 2850 2750
rect 3010 2780 3050 2785
rect 3010 2750 3015 2780
rect 3045 2750 3050 2780
rect 3010 2745 3050 2750
rect 3210 2775 3250 2785
rect 3210 2755 3220 2775
rect 3240 2755 3250 2775
rect 3210 2745 3250 2755
rect 3410 2780 3450 2785
rect 3410 2750 3415 2780
rect 3445 2750 3450 2780
rect 3410 2745 3450 2750
rect 3610 2780 3650 2785
rect 3610 2750 3615 2780
rect 3645 2750 3650 2780
rect 3610 2745 3650 2750
rect 3810 2780 3850 2785
rect 3810 2750 3815 2780
rect 3845 2750 3850 2780
rect 3810 2745 3850 2750
rect 945 2520 985 2525
rect 945 2490 950 2520
rect 980 2490 985 2520
rect 945 2485 985 2490
rect 2150 2310 2190 2315
rect 2150 2280 2155 2310
rect 2185 2280 2190 2310
rect 2150 2275 2190 2280
rect 2710 2310 2750 2315
rect 2710 2280 2715 2310
rect 2745 2280 2750 2310
rect 2710 2275 2750 2280
rect 3710 2310 3750 2315
rect 3710 2280 3715 2310
rect 3745 2280 3750 2310
rect 3710 2275 3750 2280
rect 4375 2310 4415 2315
rect 4375 2280 4380 2310
rect 4410 2280 4415 2310
rect 4375 2275 4415 2280
rect 1895 2225 2115 2230
rect 1895 2195 1900 2225
rect 2110 2195 2115 2225
rect 1895 2190 2115 2195
rect 945 2010 985 2015
rect 945 1980 950 2010
rect 980 1980 985 2010
rect 945 1975 985 1980
rect 2160 1720 2180 2275
rect 2910 2265 2950 2270
rect 2910 2235 2915 2265
rect 2945 2235 2950 2265
rect 2910 2230 2950 2235
rect 3510 2265 3550 2270
rect 3510 2235 3515 2265
rect 3545 2235 3550 2265
rect 3510 2230 3550 2235
rect 4315 2265 4355 2270
rect 4315 2235 4320 2265
rect 4350 2235 4355 2265
rect 4315 2230 4355 2235
rect 3110 2220 3150 2225
rect 3110 2190 3115 2220
rect 3145 2190 3150 2220
rect 3110 2185 3150 2190
rect 3310 2220 3350 2225
rect 3310 2190 3315 2220
rect 3345 2190 3350 2220
rect 3310 2185 3350 2190
rect 2610 2160 2650 2165
rect 2610 2130 2615 2160
rect 2645 2130 2650 2160
rect 2610 2125 2650 2130
rect 2810 2160 2850 2165
rect 2810 2130 2815 2160
rect 2845 2130 2850 2160
rect 2810 2125 2850 2130
rect 3010 2160 3050 2165
rect 3010 2130 3015 2160
rect 3045 2130 3050 2160
rect 3010 2125 3050 2130
rect 3110 2155 3150 2165
rect 3110 2135 3120 2155
rect 3140 2135 3150 2155
rect 3110 2125 3150 2135
rect 3210 2160 3250 2165
rect 3210 2130 3215 2160
rect 3245 2130 3250 2160
rect 3210 2125 3250 2130
rect 3310 2155 3350 2165
rect 3310 2135 3320 2155
rect 3340 2135 3350 2155
rect 3310 2125 3350 2135
rect 3410 2160 3450 2165
rect 3410 2130 3415 2160
rect 3445 2130 3450 2160
rect 3410 2125 3450 2130
rect 3610 2160 3650 2165
rect 3610 2130 3615 2160
rect 3645 2130 3650 2160
rect 3610 2125 3650 2130
rect 3810 2160 3850 2165
rect 3810 2130 3815 2160
rect 3845 2130 3850 2160
rect 3810 2125 3850 2130
rect 2910 1890 2950 1895
rect 2910 1860 2915 1890
rect 2945 1860 2950 1890
rect 2910 1855 2950 1860
rect 3110 1890 3150 1895
rect 3110 1860 3115 1890
rect 3145 1860 3150 1890
rect 3110 1855 3150 1860
rect 3230 1885 3270 1895
rect 3230 1865 3240 1885
rect 3260 1865 3270 1885
rect 3230 1855 3270 1865
rect 3310 1890 3350 1895
rect 3310 1860 3315 1890
rect 3345 1860 3350 1890
rect 3310 1855 3350 1860
rect 3510 1890 3550 1895
rect 3510 1860 3515 1890
rect 3545 1860 3550 1890
rect 3510 1855 3550 1860
rect 2710 1845 2750 1850
rect 2710 1815 2715 1845
rect 2745 1815 2750 1845
rect 2710 1810 2750 1815
rect 2990 1845 3030 1850
rect 2990 1815 2995 1845
rect 3025 1815 3030 1845
rect 2990 1810 3030 1815
rect 3000 1760 3020 1810
rect 2910 1755 2950 1760
rect 2910 1725 2915 1755
rect 2945 1725 2950 1755
rect 2910 1720 2950 1725
rect 2990 1755 3030 1760
rect 2990 1725 2995 1755
rect 3025 1725 3030 1755
rect 2990 1720 3030 1725
rect 465 1715 505 1720
rect 465 1685 470 1715
rect 500 1685 505 1715
rect 465 725 505 1685
rect 1895 1715 2115 1720
rect 1895 1685 1900 1715
rect 2110 1685 2115 1715
rect 1895 1680 2115 1685
rect 2150 1710 2190 1720
rect 3120 1715 3140 1855
rect 3165 1845 3205 1850
rect 3165 1815 3170 1845
rect 3200 1815 3205 1845
rect 3165 1810 3205 1815
rect 3240 1805 3260 1855
rect 3230 1800 3270 1805
rect 3230 1770 3235 1800
rect 3265 1770 3270 1800
rect 3230 1765 3270 1770
rect 3320 1715 3340 1855
rect 3430 1845 3470 1850
rect 3430 1815 3435 1845
rect 3465 1815 3470 1845
rect 3430 1810 3470 1815
rect 3710 1845 3750 1850
rect 3710 1815 3715 1845
rect 3745 1815 3750 1845
rect 3710 1810 3750 1815
rect 3440 1760 3460 1810
rect 4220 1800 4260 1805
rect 4220 1770 4225 1800
rect 4255 1770 4260 1800
rect 4220 1765 4260 1770
rect 3430 1755 3470 1760
rect 3430 1725 3435 1755
rect 3465 1725 3470 1755
rect 3430 1720 3470 1725
rect 3510 1755 3550 1760
rect 3510 1725 3515 1755
rect 3545 1725 3550 1755
rect 3510 1720 3550 1725
rect 2150 1680 2155 1710
rect 2185 1680 2190 1710
rect 2150 1675 2190 1680
rect 3050 1710 3090 1715
rect 3050 1680 3055 1710
rect 3085 1680 3090 1710
rect 3050 1675 3090 1680
rect 3110 1705 3150 1715
rect 3110 1685 3120 1705
rect 3140 1685 3150 1705
rect 3110 1675 3150 1685
rect 3310 1705 3350 1715
rect 3310 1685 3320 1705
rect 3340 1685 3350 1705
rect 3310 1675 3350 1685
rect 3370 1710 3410 1715
rect 3370 1680 3375 1710
rect 3405 1680 3410 1710
rect 3370 1675 3410 1680
rect 2910 1540 2950 1545
rect 835 1535 875 1540
rect 835 1505 840 1535
rect 870 1505 875 1535
rect 650 825 690 830
rect 650 795 655 825
rect 685 795 690 825
rect 650 790 690 795
rect 155 160 505 725
rect 835 725 875 1505
rect 945 1535 985 1540
rect 945 1505 950 1535
rect 980 1505 985 1535
rect 945 1500 985 1505
rect 1895 1535 2115 1540
rect 1895 1505 1900 1535
rect 2110 1505 2115 1535
rect 2910 1510 2915 1540
rect 2945 1510 2950 1540
rect 2910 1505 2950 1510
rect 3510 1540 3550 1545
rect 3510 1510 3515 1540
rect 3545 1510 3550 1540
rect 3510 1505 3550 1510
rect 1895 1500 2115 1505
rect 2810 1495 2850 1500
rect 2810 1465 2815 1495
rect 2845 1465 2850 1495
rect 2810 1460 2850 1465
rect 3010 1495 3050 1500
rect 3010 1465 3015 1495
rect 3045 1465 3050 1495
rect 3010 1460 3050 1465
rect 3210 1495 3250 1500
rect 3210 1465 3215 1495
rect 3245 1465 3250 1495
rect 3210 1460 3250 1465
rect 3410 1495 3450 1500
rect 3410 1465 3415 1495
rect 3445 1465 3450 1495
rect 3410 1460 3450 1465
rect 3610 1495 3650 1500
rect 3610 1465 3615 1495
rect 3645 1465 3650 1495
rect 3610 1460 3650 1465
rect 4230 1440 4250 1765
rect 4325 1545 4345 2230
rect 4385 2210 4405 2275
rect 4375 2205 4415 2210
rect 4375 2185 4385 2205
rect 4405 2185 4415 2205
rect 4375 2175 4415 2185
rect 4585 2160 4625 2165
rect 4585 2130 4590 2160
rect 4620 2130 4625 2160
rect 4585 2125 4625 2130
rect 4485 1870 4525 1880
rect 4485 1850 4495 1870
rect 4515 1850 4525 1870
rect 4485 1840 4525 1850
rect 4430 1710 4470 1715
rect 4430 1680 4435 1710
rect 4465 1680 4470 1710
rect 4430 1675 4470 1680
rect 4315 1540 4355 1545
rect 4315 1510 4320 1540
rect 4350 1510 4355 1540
rect 4315 1505 4355 1510
rect 3690 1435 3730 1440
rect 3690 1405 3695 1435
rect 3725 1405 3730 1435
rect 3690 1400 3730 1405
rect 4220 1435 4260 1440
rect 4220 1405 4225 1435
rect 4255 1405 4260 1435
rect 4220 1400 4260 1405
rect 945 1240 985 1245
rect 945 1210 950 1240
rect 980 1210 985 1240
rect 945 1205 985 1210
rect 3170 965 3290 970
rect 3170 935 3175 965
rect 3205 935 3215 965
rect 3245 935 3255 965
rect 3285 935 3290 965
rect 3170 930 3290 935
rect 4505 910 4525 1840
rect 3720 905 3760 910
rect 3720 875 3725 905
rect 3755 875 3760 905
rect 3720 870 3760 875
rect 4495 905 4535 910
rect 4495 875 4500 905
rect 4530 875 4535 905
rect 4495 870 4535 875
rect 3795 820 3835 825
rect 3795 790 3800 820
rect 3830 790 3835 820
rect 3795 785 3835 790
rect 835 690 4585 725
rect 835 160 1185 690
rect 1515 160 1865 690
rect 2195 160 2545 690
rect 2875 160 3225 690
rect 3555 160 3905 690
rect 4235 160 4585 690
<< via1 >>
rect 2615 2775 2645 2780
rect 2615 2755 2620 2775
rect 2620 2755 2640 2775
rect 2640 2755 2645 2775
rect 2615 2750 2645 2755
rect 2815 2775 2845 2780
rect 2815 2755 2820 2775
rect 2820 2755 2840 2775
rect 2840 2755 2845 2775
rect 2815 2750 2845 2755
rect 3015 2775 3045 2780
rect 3015 2755 3020 2775
rect 3020 2755 3040 2775
rect 3040 2755 3045 2775
rect 3015 2750 3045 2755
rect 3415 2775 3445 2780
rect 3415 2755 3420 2775
rect 3420 2755 3440 2775
rect 3440 2755 3445 2775
rect 3415 2750 3445 2755
rect 3615 2775 3645 2780
rect 3615 2755 3620 2775
rect 3620 2755 3640 2775
rect 3640 2755 3645 2775
rect 3615 2750 3645 2755
rect 3815 2775 3845 2780
rect 3815 2755 3820 2775
rect 3820 2755 3840 2775
rect 3840 2755 3845 2775
rect 3815 2750 3845 2755
rect 950 2515 980 2520
rect 950 2495 955 2515
rect 955 2495 975 2515
rect 975 2495 980 2515
rect 950 2490 980 2495
rect 2155 2280 2185 2310
rect 2715 2305 2745 2310
rect 2715 2285 2720 2305
rect 2720 2285 2740 2305
rect 2740 2285 2745 2305
rect 2715 2280 2745 2285
rect 3715 2305 3745 2310
rect 3715 2285 3720 2305
rect 3720 2285 3740 2305
rect 3740 2285 3745 2305
rect 3715 2280 3745 2285
rect 4380 2280 4410 2310
rect 1900 2220 2110 2225
rect 1900 2200 1905 2220
rect 1905 2200 1925 2220
rect 1925 2200 1950 2220
rect 1950 2200 1970 2220
rect 1970 2200 1995 2220
rect 1995 2200 2015 2220
rect 2015 2200 2040 2220
rect 2040 2200 2060 2220
rect 2060 2200 2085 2220
rect 2085 2200 2105 2220
rect 2105 2200 2110 2220
rect 1900 2195 2110 2200
rect 950 2005 980 2010
rect 950 1985 955 2005
rect 955 1985 975 2005
rect 975 1985 980 2005
rect 950 1980 980 1985
rect 2915 2260 2945 2265
rect 2915 2240 2920 2260
rect 2920 2240 2940 2260
rect 2940 2240 2945 2260
rect 2915 2235 2945 2240
rect 3515 2260 3545 2265
rect 3515 2240 3520 2260
rect 3520 2240 3540 2260
rect 3540 2240 3545 2260
rect 3515 2235 3545 2240
rect 4320 2235 4350 2265
rect 3115 2215 3145 2220
rect 3115 2195 3120 2215
rect 3120 2195 3140 2215
rect 3140 2195 3145 2215
rect 3115 2190 3145 2195
rect 3315 2215 3345 2220
rect 3315 2195 3320 2215
rect 3320 2195 3340 2215
rect 3340 2195 3345 2215
rect 3315 2190 3345 2195
rect 2615 2155 2645 2160
rect 2615 2135 2620 2155
rect 2620 2135 2640 2155
rect 2640 2135 2645 2155
rect 2615 2130 2645 2135
rect 2815 2155 2845 2160
rect 2815 2135 2820 2155
rect 2820 2135 2840 2155
rect 2840 2135 2845 2155
rect 2815 2130 2845 2135
rect 3015 2155 3045 2160
rect 3015 2135 3020 2155
rect 3020 2135 3040 2155
rect 3040 2135 3045 2155
rect 3015 2130 3045 2135
rect 3215 2155 3245 2160
rect 3215 2135 3220 2155
rect 3220 2135 3240 2155
rect 3240 2135 3245 2155
rect 3215 2130 3245 2135
rect 3415 2155 3445 2160
rect 3415 2135 3420 2155
rect 3420 2135 3440 2155
rect 3440 2135 3445 2155
rect 3415 2130 3445 2135
rect 3615 2155 3645 2160
rect 3615 2135 3620 2155
rect 3620 2135 3640 2155
rect 3640 2135 3645 2155
rect 3615 2130 3645 2135
rect 3815 2155 3845 2160
rect 3815 2135 3820 2155
rect 3820 2135 3840 2155
rect 3840 2135 3845 2155
rect 3815 2130 3845 2135
rect 2915 1885 2945 1890
rect 2915 1865 2920 1885
rect 2920 1865 2940 1885
rect 2940 1865 2945 1885
rect 2915 1860 2945 1865
rect 3115 1860 3145 1890
rect 3315 1860 3345 1890
rect 3515 1885 3545 1890
rect 3515 1865 3520 1885
rect 3520 1865 3540 1885
rect 3540 1865 3545 1885
rect 3515 1860 3545 1865
rect 2715 1840 2745 1845
rect 2715 1820 2720 1840
rect 2720 1820 2740 1840
rect 2740 1820 2745 1840
rect 2715 1815 2745 1820
rect 2995 1815 3025 1845
rect 2915 1750 2945 1755
rect 2915 1730 2920 1750
rect 2920 1730 2940 1750
rect 2940 1730 2945 1750
rect 2915 1725 2945 1730
rect 2995 1725 3025 1755
rect 470 1685 500 1715
rect 1900 1710 2110 1715
rect 1900 1690 1905 1710
rect 1905 1690 1925 1710
rect 1925 1690 1950 1710
rect 1950 1690 1970 1710
rect 1970 1690 1995 1710
rect 1995 1690 2015 1710
rect 2015 1690 2040 1710
rect 2040 1690 2060 1710
rect 2060 1690 2085 1710
rect 2085 1690 2105 1710
rect 2105 1690 2110 1710
rect 1900 1685 2110 1690
rect 3170 1840 3200 1845
rect 3170 1820 3175 1840
rect 3175 1820 3195 1840
rect 3195 1820 3200 1840
rect 3170 1815 3200 1820
rect 3235 1795 3265 1800
rect 3235 1775 3240 1795
rect 3240 1775 3260 1795
rect 3260 1775 3265 1795
rect 3235 1770 3265 1775
rect 3435 1815 3465 1845
rect 3715 1840 3745 1845
rect 3715 1820 3720 1840
rect 3720 1820 3740 1840
rect 3740 1820 3745 1840
rect 3715 1815 3745 1820
rect 4225 1770 4255 1800
rect 3435 1725 3465 1755
rect 3515 1750 3545 1755
rect 3515 1730 3520 1750
rect 3520 1730 3540 1750
rect 3540 1730 3545 1750
rect 3515 1725 3545 1730
rect 2155 1680 2185 1710
rect 3055 1705 3085 1710
rect 3055 1685 3060 1705
rect 3060 1685 3080 1705
rect 3080 1685 3085 1705
rect 3055 1680 3085 1685
rect 3375 1705 3405 1710
rect 3375 1685 3380 1705
rect 3380 1685 3400 1705
rect 3400 1685 3405 1705
rect 3375 1680 3405 1685
rect 840 1505 870 1535
rect 655 820 685 825
rect 655 800 660 820
rect 660 800 680 820
rect 680 800 685 820
rect 655 795 685 800
rect 950 1530 980 1535
rect 950 1510 955 1530
rect 955 1510 975 1530
rect 975 1510 980 1530
rect 950 1505 980 1510
rect 1900 1530 2110 1535
rect 1900 1510 1905 1530
rect 1905 1510 1925 1530
rect 1925 1510 1950 1530
rect 1950 1510 1970 1530
rect 1970 1510 1995 1530
rect 1995 1510 2015 1530
rect 2015 1510 2040 1530
rect 2040 1510 2060 1530
rect 2060 1510 2085 1530
rect 2085 1510 2105 1530
rect 2105 1510 2110 1530
rect 1900 1505 2110 1510
rect 2915 1535 2945 1540
rect 2915 1515 2920 1535
rect 2920 1515 2940 1535
rect 2940 1515 2945 1535
rect 2915 1510 2945 1515
rect 3515 1535 3545 1540
rect 3515 1515 3520 1535
rect 3520 1515 3540 1535
rect 3540 1515 3545 1535
rect 3515 1510 3545 1515
rect 2815 1490 2845 1495
rect 2815 1470 2820 1490
rect 2820 1470 2840 1490
rect 2840 1470 2845 1490
rect 2815 1465 2845 1470
rect 3015 1490 3045 1495
rect 3015 1470 3020 1490
rect 3020 1470 3040 1490
rect 3040 1470 3045 1490
rect 3015 1465 3045 1470
rect 3215 1490 3245 1495
rect 3215 1470 3220 1490
rect 3220 1470 3240 1490
rect 3240 1470 3245 1490
rect 3215 1465 3245 1470
rect 3415 1490 3445 1495
rect 3415 1470 3420 1490
rect 3420 1470 3440 1490
rect 3440 1470 3445 1490
rect 3415 1465 3445 1470
rect 3615 1490 3645 1495
rect 3615 1470 3620 1490
rect 3620 1470 3640 1490
rect 3640 1470 3645 1490
rect 3615 1465 3645 1470
rect 4590 2155 4620 2160
rect 4590 2135 4595 2155
rect 4595 2135 4615 2155
rect 4615 2135 4620 2155
rect 4590 2130 4620 2135
rect 4435 1705 4465 1710
rect 4435 1685 4440 1705
rect 4440 1685 4460 1705
rect 4460 1685 4465 1705
rect 4435 1680 4465 1685
rect 4320 1510 4350 1540
rect 3695 1430 3725 1435
rect 3695 1410 3700 1430
rect 3700 1410 3720 1430
rect 3720 1410 3725 1430
rect 3695 1405 3725 1410
rect 4225 1405 4255 1435
rect 950 1235 980 1240
rect 950 1215 955 1235
rect 955 1215 975 1235
rect 975 1215 980 1235
rect 950 1210 980 1215
rect 3175 960 3205 965
rect 3175 940 3180 960
rect 3180 940 3200 960
rect 3200 940 3205 960
rect 3175 935 3205 940
rect 3215 960 3245 965
rect 3215 940 3220 960
rect 3220 940 3240 960
rect 3240 940 3245 960
rect 3215 935 3245 940
rect 3255 960 3285 965
rect 3255 940 3260 960
rect 3260 940 3280 960
rect 3280 940 3285 960
rect 3255 935 3285 940
rect 3725 900 3755 905
rect 3725 880 3730 900
rect 3730 880 3750 900
rect 3750 880 3755 900
rect 3725 875 3755 880
rect 4500 875 4530 905
rect 3800 815 3830 820
rect 3800 795 3805 815
rect 3805 795 3825 815
rect 3825 795 3830 815
rect 3800 790 3830 795
<< metal2 >>
rect -130 2905 -90 2910
rect -130 2875 -125 2905
rect -95 2875 -90 2905
rect -130 2870 -90 2875
rect 4830 2905 4870 2910
rect 4830 2875 4835 2905
rect 4865 2875 4870 2905
rect 4830 2870 4870 2875
rect -130 2780 -90 2785
rect -130 2750 -125 2780
rect -95 2775 -90 2780
rect 2610 2780 2650 2785
rect 2610 2775 2615 2780
rect -95 2755 2615 2775
rect -95 2750 -90 2755
rect -130 2745 -90 2750
rect 2610 2750 2615 2755
rect 2645 2775 2650 2780
rect 2810 2780 2850 2785
rect 2810 2775 2815 2780
rect 2645 2755 2815 2775
rect 2645 2750 2650 2755
rect 2610 2745 2650 2750
rect 2810 2750 2815 2755
rect 2845 2775 2850 2780
rect 3010 2780 3050 2785
rect 3010 2775 3015 2780
rect 2845 2755 3015 2775
rect 2845 2750 2850 2755
rect 2810 2745 2850 2750
rect 3010 2750 3015 2755
rect 3045 2775 3050 2780
rect 3410 2780 3450 2785
rect 3410 2775 3415 2780
rect 3045 2755 3415 2775
rect 3045 2750 3050 2755
rect 3010 2745 3050 2750
rect 3410 2750 3415 2755
rect 3445 2775 3450 2780
rect 3610 2780 3650 2785
rect 3610 2775 3615 2780
rect 3445 2755 3615 2775
rect 3445 2750 3450 2755
rect 3410 2745 3450 2750
rect 3610 2750 3615 2755
rect 3645 2775 3650 2780
rect 3810 2780 3850 2785
rect 3810 2775 3815 2780
rect 3645 2755 3815 2775
rect 3645 2750 3650 2755
rect 3610 2745 3650 2750
rect 3810 2750 3815 2755
rect 3845 2775 3850 2780
rect 4830 2780 4870 2785
rect 4830 2775 4835 2780
rect 3845 2755 4835 2775
rect 3845 2750 3850 2755
rect 3810 2745 3850 2750
rect 4830 2750 4835 2755
rect 4865 2750 4870 2780
rect 4830 2745 4870 2750
rect -55 2520 985 2525
rect -55 2490 -50 2520
rect -20 2490 950 2520
rect 980 2490 985 2520
rect -55 2485 985 2490
rect 2150 2310 2190 2315
rect 2150 2280 2155 2310
rect 2185 2305 2190 2310
rect 2710 2310 2750 2315
rect 2710 2305 2715 2310
rect 2185 2285 2715 2305
rect 2185 2280 2190 2285
rect 2150 2275 2190 2280
rect 2710 2280 2715 2285
rect 2745 2305 2750 2310
rect 3710 2310 3750 2315
rect 3710 2305 3715 2310
rect 2745 2285 3715 2305
rect 2745 2280 2750 2285
rect 2710 2275 2750 2280
rect 3710 2280 3715 2285
rect 3745 2305 3750 2310
rect 4375 2310 4415 2315
rect 4375 2305 4380 2310
rect 3745 2285 4380 2305
rect 3745 2280 3750 2285
rect 3710 2275 3750 2280
rect 4375 2280 4380 2285
rect 4410 2280 4415 2310
rect 4375 2275 4415 2280
rect 2910 2265 2950 2270
rect 2910 2235 2915 2265
rect 2945 2260 2950 2265
rect 3510 2265 3550 2270
rect 3510 2260 3515 2265
rect 2945 2240 3515 2260
rect 2945 2235 2950 2240
rect 2910 2230 2950 2235
rect 3510 2235 3515 2240
rect 3545 2260 3550 2265
rect 4315 2265 4355 2270
rect 4315 2260 4320 2265
rect 3545 2240 4320 2260
rect 3545 2235 3550 2240
rect 3510 2230 3550 2235
rect 4315 2235 4320 2240
rect 4350 2235 4355 2265
rect 4315 2230 4355 2235
rect 1895 2225 2115 2230
rect 1895 2195 1900 2225
rect 2110 2215 2115 2225
rect 3110 2220 3150 2225
rect 3110 2215 3115 2220
rect 2110 2195 3115 2215
rect 1895 2190 2115 2195
rect 3110 2190 3115 2195
rect 3145 2215 3150 2220
rect 3310 2220 3350 2225
rect 3310 2215 3315 2220
rect 3145 2195 3315 2215
rect 3145 2190 3150 2195
rect 3110 2185 3150 2190
rect 3310 2190 3315 2195
rect 3345 2190 3350 2220
rect 3310 2185 3350 2190
rect -130 2160 -90 2165
rect -130 2130 -125 2160
rect -95 2155 -90 2160
rect 2610 2160 2650 2165
rect 2610 2155 2615 2160
rect -95 2135 2615 2155
rect -95 2130 -90 2135
rect -130 2125 -90 2130
rect 2610 2130 2615 2135
rect 2645 2155 2650 2160
rect 2810 2160 2850 2165
rect 2810 2155 2815 2160
rect 2645 2135 2815 2155
rect 2645 2130 2650 2135
rect 2610 2125 2650 2130
rect 2810 2130 2815 2135
rect 2845 2155 2850 2160
rect 3010 2160 3050 2165
rect 3010 2155 3015 2160
rect 2845 2135 3015 2155
rect 2845 2130 2850 2135
rect 2810 2125 2850 2130
rect 3010 2130 3015 2135
rect 3045 2155 3050 2160
rect 3210 2160 3250 2165
rect 3210 2155 3215 2160
rect 3045 2135 3215 2155
rect 3045 2130 3050 2135
rect 3010 2125 3050 2130
rect 3210 2130 3215 2135
rect 3245 2155 3250 2160
rect 3410 2160 3450 2165
rect 3410 2155 3415 2160
rect 3245 2135 3415 2155
rect 3245 2130 3250 2135
rect 3210 2125 3250 2130
rect 3410 2130 3415 2135
rect 3445 2155 3450 2160
rect 3610 2160 3650 2165
rect 3610 2155 3615 2160
rect 3445 2135 3615 2155
rect 3445 2130 3450 2135
rect 3410 2125 3450 2130
rect 3610 2130 3615 2135
rect 3645 2155 3650 2160
rect 3810 2160 3850 2165
rect 3810 2155 3815 2160
rect 3645 2135 3815 2155
rect 3645 2130 3650 2135
rect 3610 2125 3650 2130
rect 3810 2130 3815 2135
rect 3845 2155 3850 2160
rect 4585 2160 4625 2165
rect 4585 2155 4590 2160
rect 3845 2135 4590 2155
rect 3845 2130 3850 2135
rect 3810 2125 3850 2130
rect 4585 2130 4590 2135
rect 4620 2155 4625 2160
rect 4830 2160 4870 2165
rect 4830 2155 4835 2160
rect 4620 2135 4835 2155
rect 4620 2130 4625 2135
rect 4585 2125 4625 2130
rect 4830 2130 4835 2135
rect 4865 2130 4870 2160
rect 4830 2125 4870 2130
rect -55 2010 985 2015
rect -55 1980 -50 2010
rect -20 1980 950 2010
rect 980 1980 985 2010
rect -55 1975 985 1980
rect 2910 1890 2950 1895
rect 2910 1860 2915 1890
rect 2945 1885 2950 1890
rect 3110 1890 3150 1895
rect 3110 1885 3115 1890
rect 2945 1865 3115 1885
rect 2945 1860 2950 1865
rect 2910 1855 2950 1860
rect 3110 1860 3115 1865
rect 3145 1885 3150 1890
rect 3310 1890 3350 1895
rect 3310 1885 3315 1890
rect 3145 1865 3315 1885
rect 3145 1860 3150 1865
rect 3110 1855 3150 1860
rect 3310 1860 3315 1865
rect 3345 1885 3350 1890
rect 3510 1890 3550 1895
rect 3510 1885 3515 1890
rect 3345 1865 3515 1885
rect 3345 1860 3350 1865
rect 3310 1855 3350 1860
rect 3510 1860 3515 1865
rect 3545 1860 3550 1890
rect 3510 1855 3550 1860
rect 2710 1845 2750 1850
rect 2710 1815 2715 1845
rect 2745 1840 2750 1845
rect 2990 1845 3030 1850
rect 2990 1840 2995 1845
rect 2745 1820 2995 1840
rect 2745 1815 2750 1820
rect 2710 1810 2750 1815
rect 2990 1815 2995 1820
rect 3025 1840 3030 1845
rect 3165 1845 3205 1850
rect 3165 1840 3170 1845
rect 3025 1820 3170 1840
rect 3025 1815 3030 1820
rect 2990 1810 3030 1815
rect 3165 1815 3170 1820
rect 3200 1840 3205 1845
rect 3430 1845 3470 1850
rect 3430 1840 3435 1845
rect 3200 1820 3435 1840
rect 3200 1815 3205 1820
rect 3165 1810 3205 1815
rect 3430 1815 3435 1820
rect 3465 1840 3470 1845
rect 3710 1845 3750 1850
rect 3710 1840 3715 1845
rect 3465 1820 3715 1840
rect 3465 1815 3470 1820
rect 3430 1810 3470 1815
rect 3710 1815 3715 1820
rect 3745 1815 3750 1845
rect 3710 1810 3750 1815
rect 3230 1800 3270 1805
rect 3230 1770 3235 1800
rect 3265 1795 3270 1800
rect 4220 1800 4260 1805
rect 4220 1795 4225 1800
rect 3265 1775 4225 1795
rect 3265 1770 3270 1775
rect 3230 1765 3270 1770
rect 4220 1770 4225 1775
rect 4255 1770 4260 1800
rect 4220 1765 4260 1770
rect 2910 1755 2950 1760
rect 2910 1725 2915 1755
rect 2945 1750 2950 1755
rect 2990 1755 3030 1760
rect 2990 1750 2995 1755
rect 2945 1730 2995 1750
rect 2945 1725 2950 1730
rect 2910 1720 2950 1725
rect 2990 1725 2995 1730
rect 3025 1750 3030 1755
rect 3430 1755 3470 1760
rect 3430 1750 3435 1755
rect 3025 1730 3435 1750
rect 3025 1725 3030 1730
rect 2990 1720 3030 1725
rect 3430 1725 3435 1730
rect 3465 1750 3470 1755
rect 3510 1755 3550 1760
rect 3510 1750 3515 1755
rect 3465 1730 3515 1750
rect 3465 1725 3470 1730
rect 3430 1720 3470 1725
rect 3510 1725 3515 1730
rect 3545 1725 3550 1755
rect 3510 1720 3550 1725
rect 465 1715 2115 1720
rect 465 1685 470 1715
rect 500 1685 1900 1715
rect 2110 1705 2115 1715
rect 2150 1710 2190 1720
rect 2150 1705 2155 1710
rect 2110 1685 2155 1705
rect 465 1680 2115 1685
rect 2150 1680 2155 1685
rect 2185 1705 2190 1710
rect 3050 1710 3090 1715
rect 3050 1705 3055 1710
rect 2185 1685 3055 1705
rect 2185 1680 2190 1685
rect 2150 1675 2190 1680
rect 3050 1680 3055 1685
rect 3085 1705 3090 1710
rect 3370 1710 3410 1715
rect 3370 1705 3375 1710
rect 3085 1685 3375 1705
rect 3085 1680 3090 1685
rect 3050 1675 3090 1680
rect 3370 1680 3375 1685
rect 3405 1705 3410 1710
rect 4430 1710 4470 1715
rect 4430 1705 4435 1710
rect 3405 1685 4435 1705
rect 3405 1680 3410 1685
rect 3370 1675 3410 1680
rect 4430 1680 4435 1685
rect 4465 1680 4470 1710
rect 4430 1675 4470 1680
rect 2910 1540 2950 1545
rect 835 1535 985 1540
rect 835 1505 840 1535
rect 870 1505 950 1535
rect 980 1505 985 1535
rect 835 1500 985 1505
rect 1895 1535 2115 1540
rect 2910 1535 2915 1540
rect 1895 1505 1900 1535
rect 2110 1515 2915 1535
rect 2110 1505 2115 1515
rect 2910 1510 2915 1515
rect 2945 1535 2950 1540
rect 3510 1540 3550 1545
rect 3510 1535 3515 1540
rect 2945 1515 3515 1535
rect 2945 1510 2950 1515
rect 2910 1505 2950 1510
rect 3510 1510 3515 1515
rect 3545 1535 3550 1540
rect 4315 1540 4355 1545
rect 4315 1535 4320 1540
rect 3545 1515 4320 1535
rect 3545 1510 3550 1515
rect 3510 1505 3550 1510
rect 4315 1510 4320 1515
rect 4350 1510 4355 1540
rect 4315 1505 4355 1510
rect 1895 1500 2115 1505
rect 2810 1495 2850 1500
rect 2810 1465 2815 1495
rect 2845 1490 2850 1495
rect 3010 1495 3050 1500
rect 3010 1490 3015 1495
rect 2845 1470 3015 1490
rect 2845 1465 2850 1470
rect 2810 1460 2850 1465
rect 3010 1465 3015 1470
rect 3045 1490 3050 1495
rect 3210 1495 3250 1500
rect 3210 1490 3215 1495
rect 3045 1470 3215 1490
rect 3045 1465 3050 1470
rect 3010 1460 3050 1465
rect 3210 1465 3215 1470
rect 3245 1490 3250 1495
rect 3410 1495 3450 1500
rect 3410 1490 3415 1495
rect 3245 1470 3415 1490
rect 3245 1465 3250 1470
rect 3210 1460 3250 1465
rect 3410 1465 3415 1470
rect 3445 1490 3450 1495
rect 3610 1495 3650 1500
rect 3610 1490 3615 1495
rect 3445 1470 3615 1490
rect 3445 1465 3450 1470
rect 3410 1460 3450 1465
rect 3610 1465 3615 1470
rect 3645 1465 3650 1495
rect 3610 1460 3650 1465
rect 3690 1435 3730 1440
rect 3690 1405 3695 1435
rect 3725 1430 3730 1435
rect 4220 1435 4260 1440
rect 4220 1430 4225 1435
rect 3725 1410 4225 1430
rect 3725 1405 3730 1410
rect 3690 1400 3730 1405
rect 4220 1405 4225 1410
rect 4255 1405 4260 1435
rect 4220 1400 4260 1405
rect -55 1240 985 1245
rect -55 1210 -50 1240
rect -20 1210 950 1240
rect 980 1210 985 1240
rect -55 1205 985 1210
rect -55 965 -15 970
rect -55 935 -50 965
rect -20 960 -15 965
rect 3170 965 3290 970
rect 3170 960 3175 965
rect -20 940 3175 960
rect -20 935 -15 940
rect -55 930 -15 935
rect 3170 935 3175 940
rect 3205 935 3215 965
rect 3245 935 3255 965
rect 3285 960 3290 965
rect 4755 965 4795 970
rect 4755 960 4760 965
rect 3285 940 4760 960
rect 3285 935 3290 940
rect 3170 930 3290 935
rect 4755 935 4760 940
rect 4790 935 4795 965
rect 4755 930 4795 935
rect 3720 905 3760 910
rect 3720 875 3725 905
rect 3755 900 3760 905
rect 4495 905 4535 910
rect 4495 900 4500 905
rect 3755 880 4500 900
rect 3755 875 3760 880
rect 3720 870 3760 875
rect 4495 875 4500 880
rect 4530 875 4535 905
rect 4495 870 4535 875
rect -55 825 -15 830
rect -55 795 -50 825
rect -20 820 -15 825
rect 650 825 690 830
rect 650 820 655 825
rect -20 800 655 820
rect -20 795 -15 800
rect -55 790 -15 795
rect 650 795 655 800
rect 685 795 690 825
rect 650 790 690 795
rect 3795 820 3835 825
rect 3795 790 3800 820
rect 3830 815 3835 820
rect 4755 820 4795 825
rect 4755 815 4760 820
rect 3830 795 4760 815
rect 3830 790 3835 795
rect 3795 785 3835 790
rect 4755 790 4760 795
rect 4790 790 4795 820
rect 4755 785 4795 790
rect -130 -90 -90 -85
rect -130 -120 -125 -90
rect -95 -120 -90 -90
rect -130 -125 -90 -120
<< via2 >>
rect -125 2875 -95 2905
rect 4835 2875 4865 2905
rect -125 2750 -95 2780
rect 4835 2750 4865 2780
rect -50 2490 -20 2520
rect -125 2130 -95 2160
rect 4835 2130 4865 2160
rect -50 1980 -20 2010
rect -50 1210 -20 1240
rect -50 935 -20 965
rect 4760 935 4790 965
rect -50 795 -20 825
rect 4760 790 4790 820
rect -125 -120 -95 -90
<< metal3 >>
rect -135 2910 -85 2915
rect -135 2870 -130 2910
rect -90 2870 -85 2910
rect -135 2865 -85 2870
rect 4825 2910 4875 2915
rect 4825 2870 4830 2910
rect 4870 2870 4875 2910
rect 4825 2865 4875 2870
rect -130 2780 -90 2865
rect -60 2835 -10 2840
rect -60 2795 -55 2835
rect -15 2795 -10 2835
rect -60 2790 -10 2795
rect 4750 2835 4800 2840
rect 4750 2795 4755 2835
rect 4795 2795 4800 2835
rect 4750 2790 4800 2795
rect -130 2750 -125 2780
rect -95 2750 -90 2780
rect -130 2160 -90 2750
rect -130 2130 -125 2160
rect -95 2130 -90 2160
rect -130 -80 -90 2130
rect -55 2520 -15 2790
rect -55 2490 -50 2520
rect -20 2490 -15 2520
rect -55 2010 -15 2490
rect -55 1980 -50 2010
rect -20 1980 -15 2010
rect -55 1240 -15 1980
rect -55 1210 -50 1240
rect -20 1210 -15 1240
rect -55 965 -15 1210
rect -55 935 -50 965
rect -20 935 -15 965
rect -55 825 -15 935
rect -55 795 -50 825
rect -20 795 -15 825
rect -55 -5 -15 795
rect 4755 965 4795 2790
rect 4755 935 4760 965
rect 4790 935 4795 965
rect 4755 820 4795 935
rect 4755 790 4760 820
rect 4790 790 4795 820
rect 4755 -5 4795 790
rect 4830 2780 4870 2865
rect 4830 2750 4835 2780
rect 4865 2750 4870 2780
rect 4830 2160 4870 2750
rect 4830 2130 4835 2160
rect 4865 2130 4870 2160
rect -60 -10 -10 -5
rect -60 -50 -55 -10
rect -15 -50 -10 -10
rect -60 -55 -10 -50
rect 4750 -10 4800 -5
rect 4750 -50 4755 -10
rect 4795 -50 4800 -10
rect 4750 -55 4800 -50
rect 4830 -80 4870 2130
rect -135 -85 -85 -80
rect -135 -125 -130 -85
rect -90 -125 -85 -85
rect -135 -130 -85 -125
rect 4825 -85 4875 -80
rect 4825 -125 4830 -85
rect 4870 -125 4875 -85
rect 4825 -130 4875 -125
<< via3 >>
rect -130 2905 -90 2910
rect -130 2875 -125 2905
rect -125 2875 -95 2905
rect -95 2875 -90 2905
rect -130 2870 -90 2875
rect 4830 2905 4870 2910
rect 4830 2875 4835 2905
rect 4835 2875 4865 2905
rect 4865 2875 4870 2905
rect 4830 2870 4870 2875
rect -55 2795 -15 2835
rect 4755 2795 4795 2835
rect -55 -50 -15 -10
rect 4755 -50 4795 -10
rect -130 -90 -90 -85
rect -130 -120 -125 -90
rect -125 -120 -95 -90
rect -95 -120 -90 -90
rect -130 -125 -90 -120
rect 4830 -125 4870 -85
<< metal4 >>
rect -135 2910 -85 2915
rect 4825 2910 4875 2915
rect -135 2870 -130 2910
rect -90 2870 4830 2910
rect 4870 2870 4875 2910
rect -135 2865 -85 2870
rect 4825 2865 4875 2870
rect -60 2835 -10 2840
rect 4750 2835 4800 2840
rect -60 2795 -55 2835
rect -15 2795 4755 2835
rect 4795 2795 4800 2835
rect -60 2790 -10 2795
rect 4750 2790 4800 2795
rect -60 -10 -10 -5
rect 4750 -10 4800 -5
rect -60 -50 -55 -10
rect -15 -50 4755 -10
rect 4795 -50 4800 -10
rect -60 -55 -10 -50
rect 4750 -55 4800 -50
rect -135 -85 -85 -80
rect 4825 -85 4875 -80
rect -135 -125 -130 -85
rect -90 -125 4830 -85
rect 4870 -125 4875 -85
rect -135 -130 -85 -125
rect 4825 -130 4875 -125
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 675 0 1 0
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1723858470
transform 1 0 -5 0 1 0
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1723858470
transform 1 0 1355 0 1 0
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1723858470
transform 1 0 2035 0 1 0
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1723858470
transform 1 0 2715 0 1 0
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1723858470
transform 1 0 3395 0 1 0
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1723858470
transform 1 0 4075 0 1 0
box 0 0 670 670
<< labels >>
flabel metal3 4870 1400 4870 1400 3 FreeSans 800 0 80 0 VDDA
port 1 e
flabel metal3 4795 1175 4795 1175 3 FreeSans 800 0 80 0 GNDA
port 6 e
flabel metal1 3230 3150 3230 3150 1 FreeSans 800 0 0 400 V_out
port 5 n
flabel metal1 4525 1615 4525 1615 3 FreeSans 400 0 80 0 start_up
flabel locali 2820 1450 2820 1450 7 FreeSans 400 0 -80 0 V_p
flabel metal2 2285 1685 2285 1685 5 FreeSans 400 0 0 -80 Vin-
flabel metal2 2285 1515 2285 1515 5 FreeSans 400 0 0 -80 Vin+
flabel metal1 4415 2295 4415 2295 3 FreeSans 400 0 80 0 V_TOP
flabel metal2 3750 1830 3750 1830 3 FreeSans 400 0 80 0 1st_Vout
flabel metal1 3120 1790 3120 1790 7 FreeSans 400 0 -80 0 V_mirror
flabel metal1 875 1040 875 1040 3 FreeSans 400 0 80 0 Vbe2
<< end >>
