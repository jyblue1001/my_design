* PEX produced on Sun Jul 20 03:56:35 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 bgr_0.Vin+.t5 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 GNDA.t288 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 two_stage_opamp_dummy_magic_0.Y.t25 GNDA.t303 VDDA.t415 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X2 GNDA.t62 VDDA.t204 VDDA.t206 VDDA.t205 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X3 two_stage_opamp_dummy_magic_0.err_amp_out.t10 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 GNDA.t139 GNDA.t138 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X4 two_stage_opamp_dummy_magic_0.V_p_mir.t2 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 GNDA.t69 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X5 two_stage_opamp_dummy_magic_0.VD2.t16 GNDA.t266 GNDA.t267 GNDA.t259 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X6 VOUT+.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 VDDA.t91 bgr_0.V_mir1.t17 bgr_0.1st_Vout_1.t5 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X8 VDDA.t203 VDDA.t201 VOUT-.t6 VDDA.t202 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X9 VOUT+.t20 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 VOUT+.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X11 GNDA.t57 VDDA.t469 bgr_0.V_TOP.t6 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X12 VOUT+.t22 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 bgr_0.1st_Vout_2.t11 bgr_0.cap_res2.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X14 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 GNDA.t263 GNDA.t265 GNDA.t264 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X15 VOUT+.t23 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 GNDA.t71 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 two_stage_opamp_dummy_magic_0.V_source.t24 GNDA.t70 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X17 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 bgr_0.NFET_GATE_10uA.t5 GNDA.t313 GNDA.t312 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X18 two_stage_opamp_dummy_magic_0.Y.t22 two_stage_opamp_dummy_magic_0.Vb2.t11 two_stage_opamp_dummy_magic_0.VD4.t21 two_stage_opamp_dummy_magic_0.VD4.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X19 VOUT+.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 VOUT+.t25 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 GNDA.t119 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 two_stage_opamp_dummy_magic_0.V_source.t23 GNDA.t118 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X22 a_7460_23988.t0 bgr_0.Vin+.t4 GNDA.t133 sky130_fd_pr__res_xhigh_po_0p35 l=6
X23 bgr_0.V_mir2.t4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 bgr_0.V_p_2.t6 GNDA.t144 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X24 VDDA.t200 VDDA.t198 VDDA.t200 VDDA.t199 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X25 VOUT+.t26 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X26 bgr_0.1st_Vout_2.t12 bgr_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 two_stage_opamp_dummy_magic_0.Vb1.t13 bgr_0.PFET_GATE_10uA.t10 VDDA.t276 VDDA.t275 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X28 two_stage_opamp_dummy_magic_0.V_err_p.t20 two_stage_opamp_dummy_magic_0.V_err_gate.t14 VDDA.t269 VDDA.t268 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X29 two_stage_opamp_dummy_magic_0.X.t23 GNDA.t261 GNDA.t262 GNDA.t173 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X30 two_stage_opamp_dummy_magic_0.X.t14 two_stage_opamp_dummy_magic_0.Vb1.t14 two_stage_opamp_dummy_magic_0.VD1.t14 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X31 GNDA.t137 a_6930_22564.t0 GNDA.t36 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X32 VDDA.t197 VDDA.t195 bgr_0.V_TOP.t5 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X33 VOUT-.t19 two_stage_opamp_dummy_magic_0.cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 VOUT-.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 VOUT-.t21 two_stage_opamp_dummy_magic_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 VOUT+.t27 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 bgr_0.1st_Vout_1.t11 bgr_0.cap_res1.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 VOUT+.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 VOUT+.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 bgr_0.PFET_GATE_10uA.t11 VDDA.t338 VDDA.t337 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X41 VDDA.t414 two_stage_opamp_dummy_magic_0.Y.t26 VOUT+.t16 VDDA.t413 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X42 VOUT-.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 VDDA.t443 bgr_0.PFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 VDDA.t442 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X44 two_stage_opamp_dummy_magic_0.Y.t21 GNDA.t258 GNDA.t260 GNDA.t259 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X45 VOUT+.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 bgr_0.cap_res2.t0 bgr_0.PFET_GATE_10uA.t0 GNDA.t55 sky130_fd_pr__res_high_po_0p35 l=2.05
X47 VDDA.t73 bgr_0.V_mir2.t17 bgr_0.1st_Vout_2.t3 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X48 bgr_0.1st_Vout_1.t12 bgr_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 VDDA.t412 two_stage_opamp_dummy_magic_0.Y.t27 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 GNDA.t304 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X50 VDDA.t85 bgr_0.1st_Vout_1.t13 bgr_0.V_TOP.t12 VDDA.t84 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X51 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 two_stage_opamp_dummy_magic_0.V_tot.t4 two_stage_opamp_dummy_magic_0.V_err_p.t1 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X52 VOUT+.t31 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X53 VOUT-.t23 two_stage_opamp_dummy_magic_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X54 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 two_stage_opamp_dummy_magic_0.X.t25 VDDA.t240 GNDA.t140 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X55 bgr_0.START_UP.t1 bgr_0.START_UP.t0 bgr_0.START_UP_NFET1.t0 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X56 two_stage_opamp_dummy_magic_0.Y.t16 two_stage_opamp_dummy_magic_0.Vb2.t12 two_stage_opamp_dummy_magic_0.VD4.t19 two_stage_opamp_dummy_magic_0.VD4.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X57 VOUT-.t24 two_stage_opamp_dummy_magic_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X58 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 GNDA.t128 GNDA.t127 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X59 bgr_0.V_TOP.t14 VDDA.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X60 VOUT-.t25 two_stage_opamp_dummy_magic_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 two_stage_opamp_dummy_magic_0.V_err_gate.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 two_stage_opamp_dummy_magic_0.V_er_mir_p.t4 VDDA.t433 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X62 two_stage_opamp_dummy_magic_0.VD1.t17 VIN-.t0 two_stage_opamp_dummy_magic_0.V_source.t33 GNDA.t167 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X63 VOUT-.t26 two_stage_opamp_dummy_magic_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X64 VOUT+.t32 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X65 VOUT-.t27 two_stage_opamp_dummy_magic_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 VOUT-.t28 two_stage_opamp_dummy_magic_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 VOUT-.t29 two_stage_opamp_dummy_magic_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 VOUT+.t15 two_stage_opamp_dummy_magic_0.Y.t28 VDDA.t411 VDDA.t410 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X69 two_stage_opamp_dummy_magic_0.V_source.t22 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 GNDA.t121 GNDA.t120 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X70 bgr_0.V_mir2.t16 bgr_0.V_mir2.t15 VDDA.t19 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X71 two_stage_opamp_dummy_magic_0.VD3.t31 two_stage_opamp_dummy_magic_0.Vb3.t8 VDDA.t375 VDDA.t374 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X72 VOUT+.t33 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X73 VDDA.t285 bgr_0.V_mir1.t14 bgr_0.V_mir1.t15 VDDA.t284 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X74 bgr_0.1st_Vout_1.t14 bgr_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 VDDA.t239 two_stage_opamp_dummy_magic_0.X.t26 VOUT-.t8 VDDA.t238 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X76 two_stage_opamp_dummy_magic_0.VD2.t9 VIN+.t0 two_stage_opamp_dummy_magic_0.V_source.t26 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X77 VDDA.t298 two_stage_opamp_dummy_magic_0.V_err_gate.t15 two_stage_opamp_dummy_magic_0.V_er_mir_p.t19 VDDA.t297 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X78 bgr_0.V_TOP.t15 VDDA.t246 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 VOUT-.t30 two_stage_opamp_dummy_magic_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X80 bgr_0.1st_Vout_2.t2 bgr_0.V_CUR_REF_REG.t3 bgr_0.V_p_2.t2 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X81 two_stage_opamp_dummy_magic_0.Vb2_2.t2 two_stage_opamp_dummy_magic_0.Vb2.t13 VDDA.t242 VDDA.t241 sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.36 ps=2.2 w=1.8 l=0.2
X82 VOUT+.t34 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 bgr_0.V_TOP.t16 VDDA.t247 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 GNDA.t154 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 two_stage_opamp_dummy_magic_0.V_source.t21 GNDA.t153 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X85 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 bgr_0.PFET_GATE_10uA.t13 VDDA.t458 VDDA.t457 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X86 VDDA.t263 bgr_0.PFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 VDDA.t262 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X87 GNDA.t257 GNDA.t256 two_stage_opamp_dummy_magic_0.VD1.t19 GNDA.t249 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X88 VOUT-.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 two_stage_opamp_dummy_magic_0.V_err_p.t19 two_stage_opamp_dummy_magic_0.V_err_gate.t16 VDDA.t447 VDDA.t446 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X90 VOUT-.t32 two_stage_opamp_dummy_magic_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X91 GNDA.t255 GNDA.t253 VOUT+.t5 GNDA.t254 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X92 bgr_0.Vin-.t5 bgr_0.V_TOP.t17 VDDA.t46 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X93 bgr_0.PFET_GATE_10uA.t9 bgr_0.1st_Vout_2.t13 VDDA.t314 VDDA.t313 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X94 VOUT+.t35 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 VOUT-.t33 two_stage_opamp_dummy_magic_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X96 two_stage_opamp_dummy_magic_0.X.t17 two_stage_opamp_dummy_magic_0.Vb1.t15 two_stage_opamp_dummy_magic_0.VD1.t13 GNDA.t167 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X97 two_stage_opamp_dummy_magic_0.VD3.t37 two_stage_opamp_dummy_magic_0.VD3.t35 two_stage_opamp_dummy_magic_0.X.t10 two_stage_opamp_dummy_magic_0.VD3.t36 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X98 bgr_0.1st_Vout_1.t10 bgr_0.Vin+.t6 bgr_0.V_p_1.t10 GNDA.t293 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X99 VDDA.t194 VDDA.t192 GNDA.t63 VDDA.t193 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X100 VOUT+.t36 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X101 GNDA.t59 VDDA.t470 bgr_0.V_p_2.t8 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X102 two_stage_opamp_dummy_magic_0.VD3.t30 two_stage_opamp_dummy_magic_0.Vb3.t9 VDDA.t366 VDDA.t365 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X103 GNDA.t252 GNDA.t251 two_stage_opamp_dummy_magic_0.VD2.t15 GNDA.t246 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X104 a_5310_4968.t0 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA.t54 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X105 VOUT-.t34 two_stage_opamp_dummy_magic_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X106 bgr_0.V_TOP.t18 VDDA.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 VDDA.t316 bgr_0.1st_Vout_2.t14 bgr_0.PFET_GATE_10uA.t8 VDDA.t315 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X108 two_stage_opamp_dummy_magic_0.Y.t1 two_stage_opamp_dummy_magic_0.Vb1.t16 two_stage_opamp_dummy_magic_0.VD2.t3 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X109 two_stage_opamp_dummy_magic_0.err_amp_out.t11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 two_stage_opamp_dummy_magic_0.V_err_p.t6 VDDA.t450 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X110 VDDA.t408 two_stage_opamp_dummy_magic_0.Y.t29 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 GNDA.t305 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X111 a_14560_4968.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 GNDA.t136 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X112 VOUT+.t37 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 two_stage_opamp_dummy_magic_0.X.t27 VDDA.t16 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X114 bgr_0.V_TOP.t19 VDDA.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 bgr_0.V_TOP.t4 VDDA.t189 VDDA.t191 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X116 VOUT-.t35 two_stage_opamp_dummy_magic_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X117 GNDA.t123 bgr_0.NFET_GATE_10uA.t6 two_stage_opamp_dummy_magic_0.Vb3.t5 GNDA.t122 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X118 VOUT-.t36 two_stage_opamp_dummy_magic_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 bgr_0.1st_Vout_1.t7 bgr_0.Vin+.t7 bgr_0.V_p_1.t9 GNDA.t292 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X120 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 bgr_0.V_TOP.t20 VDDA.t44 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X121 VOUT-.t37 two_stage_opamp_dummy_magic_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 VOUT-.t38 two_stage_opamp_dummy_magic_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 VOUT-.t39 two_stage_opamp_dummy_magic_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 bgr_0.1st_Vout_2.t15 bgr_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 two_stage_opamp_dummy_magic_0.V_err_gate.t0 two_stage_opamp_dummy_magic_0.V_tot.t5 two_stage_opamp_dummy_magic_0.V_er_mir_p.t9 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X126 GNDA.t250 GNDA.t248 two_stage_opamp_dummy_magic_0.X.t22 GNDA.t249 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X127 VOUT+.t38 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 VOUT+.t39 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 VDDA.t68 bgr_0.1st_Vout_1.t15 bgr_0.V_TOP.t11 VDDA.t67 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X130 VOUT+.t40 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 two_stage_opamp_dummy_magic_0.Y.t30 GNDA.t306 VDDA.t409 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X132 VOUT+.t41 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 VOUT-.t18 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 GNDA.t296 GNDA.t295 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X134 VOUT+.t42 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X135 a_12530_23988.t0 bgr_0.Vin-.t6 GNDA.t135 sky130_fd_pr__res_xhigh_po_0p35 l=6
X136 VOUT+.t14 two_stage_opamp_dummy_magic_0.Y.t31 VDDA.t407 VDDA.t406 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X137 two_stage_opamp_dummy_magic_0.V_source.t20 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 GNDA.t156 GNDA.t155 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X138 VDDA.t51 two_stage_opamp_dummy_magic_0.X.t28 VOUT-.t2 VDDA.t50 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X139 GNDA.t247 GNDA.t245 two_stage_opamp_dummy_magic_0.Y.t20 GNDA.t246 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X140 two_stage_opamp_dummy_magic_0.VD4.t23 VDDA.t179 VDDA.t181 VDDA.t180 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X141 GNDA.t300 bgr_0.NFET_GATE_10uA.t7 two_stage_opamp_dummy_magic_0.Vb2.t8 GNDA.t299 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X142 GNDA.t77 bgr_0.NFET_GATE_10uA.t8 two_stage_opamp_dummy_magic_0.Vb2.t7 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X143 bgr_0.1st_Vout_2.t1 bgr_0.V_CUR_REF_REG.t4 bgr_0.V_p_2.t1 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X144 VDDA.t460 two_stage_opamp_dummy_magic_0.V_err_gate.t17 two_stage_opamp_dummy_magic_0.V_err_p.t18 VDDA.t459 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X145 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 bgr_0.NFET_GATE_10uA.t9 GNDA.t281 GNDA.t280 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X146 two_stage_opamp_dummy_magic_0.VD4.t17 two_stage_opamp_dummy_magic_0.Vb2.t14 two_stage_opamp_dummy_magic_0.Y.t6 two_stage_opamp_dummy_magic_0.VD4.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X147 VDDA.t188 VDDA.t186 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 VDDA.t187 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X148 VOUT-.t40 two_stage_opamp_dummy_magic_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 GNDA.t47 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 two_stage_opamp_dummy_magic_0.V_source.t19 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X150 VDDA.t213 bgr_0.PFET_GATE_10uA.t15 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X151 VOUT-.t41 two_stage_opamp_dummy_magic_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 bgr_0.1st_Vout_2.t16 bgr_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X153 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 bgr_0.PFET_GATE_10uA.t16 VDDA.t220 VDDA.t219 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X154 two_stage_opamp_dummy_magic_0.VD3.t29 two_stage_opamp_dummy_magic_0.Vb3.t10 VDDA.t216 VDDA.t215 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X155 VOUT-.t17 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 GNDA.t287 GNDA.t286 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X156 VDDA.t185 VDDA.t182 VDDA.t184 VDDA.t183 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0 ps=0 w=1.8 l=0.2
X157 VOUT-.t42 two_stage_opamp_dummy_magic_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 VOUT+.t43 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 two_stage_opamp_dummy_magic_0.V_source.t38 VIN-.t1 two_stage_opamp_dummy_magic_0.VD1.t20 GNDA.t147 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X160 two_stage_opamp_dummy_magic_0.V_er_mir_p.t18 two_stage_opamp_dummy_magic_0.V_err_gate.t18 VDDA.t267 VDDA.t266 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X161 VOUT-.t43 two_stage_opamp_dummy_magic_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 VOUT+.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X163 VOUT+.t45 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 bgr_0.1st_Vout_1.t16 bgr_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 GNDA.t307 two_stage_opamp_dummy_magic_0.Y.t32 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 VDDA.t405 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X166 VOUT+.t4 GNDA.t242 GNDA.t244 GNDA.t243 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X167 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 two_stage_opamp_dummy_magic_0.X.t29 GNDA.t323 VDDA.t428 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X168 GNDA.t49 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 two_stage_opamp_dummy_magic_0.V_source.t18 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X169 a_14680_4968.t0 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA.t20 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X170 VDDA.t66 bgr_0.V_mir1.t12 bgr_0.V_mir1.t13 VDDA.t65 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X171 GNDA.t134 a_7580_22380.t0 GNDA.t133 sky130_fd_pr__res_xhigh_po_0p35 l=6
X172 two_stage_opamp_dummy_magic_0.V_source.t4 VIN+.t1 two_stage_opamp_dummy_magic_0.VD2.t4 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X173 VOUT-.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 VOUT-.t45 two_stage_opamp_dummy_magic_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 VOUT+.t46 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 VOUT-.t46 two_stage_opamp_dummy_magic_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 VOUT-.t47 two_stage_opamp_dummy_magic_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X178 VOUT-.t48 two_stage_opamp_dummy_magic_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X179 two_stage_opamp_dummy_magic_0.VD4.t15 two_stage_opamp_dummy_magic_0.Vb2.t15 two_stage_opamp_dummy_magic_0.Y.t8 two_stage_opamp_dummy_magic_0.VD4.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X180 two_stage_opamp_dummy_magic_0.Vb1.t3 two_stage_opamp_dummy_magic_0.Vb1.t2 two_stage_opamp_dummy_magic_0.Vb1_2.t4 GNDA.t132 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X181 bgr_0.V_TOP.t21 VDDA.t350 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 VDDA.t176 VDDA.t178 VDDA.t177 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X183 a_5190_4968.t0 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA.t19 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X184 VDDA.t376 two_stage_opamp_dummy_magic_0.Y.t33 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 GNDA.t308 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X185 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 two_stage_opamp_dummy_magic_0.V_tot.t6 two_stage_opamp_dummy_magic_0.V_err_p.t10 VDDA.t237 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X186 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 two_stage_opamp_dummy_magic_0.X.t30 VDDA.t430 GNDA.t326 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X187 VOUT-.t49 two_stage_opamp_dummy_magic_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 VOUT-.t50 two_stage_opamp_dummy_magic_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 two_stage_opamp_dummy_magic_0.V_source.t17 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 GNDA.t33 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X190 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 two_stage_opamp_dummy_magic_0.X.t31 VDDA.t364 GNDA.t283 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X191 GNDA.t241 GNDA.t239 bgr_0.NFET_GATE_10uA.t3 GNDA.t240 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X192 VOUT+.t47 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X193 VOUT+.t48 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X194 two_stage_opamp_dummy_magic_0.V_err_gate.t10 bgr_0.NFET_GATE_10uA.t10 GNDA.t42 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X195 VOUT+.t3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 GNDA.t94 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X196 VOUT+.t49 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 two_stage_opamp_dummy_magic_0.Vb2.t0 two_stage_opamp_dummy_magic_0.Vb2_2.t7 two_stage_opamp_dummy_magic_0.Vb2_2.t9 two_stage_opamp_dummy_magic_0.Vb2_2.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X198 VOUT+.t50 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 two_stage_opamp_dummy_magic_0.Vb2.t6 bgr_0.NFET_GATE_10uA.t11 GNDA.t125 GNDA.t124 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X200 VDDA.t59 bgr_0.V_mir1.t18 bgr_0.1st_Vout_1.t4 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X201 two_stage_opamp_dummy_magic_0.V_err_gate.t8 VDDA.t173 VDDA.t175 VDDA.t174 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X202 two_stage_opamp_dummy_magic_0.VD1.t12 two_stage_opamp_dummy_magic_0.Vb1.t17 two_stage_opamp_dummy_magic_0.X.t13 GNDA.t147 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X203 VDDA.t280 two_stage_opamp_dummy_magic_0.Vb3.t11 two_stage_opamp_dummy_magic_0.VD3.t28 VDDA.t279 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X204 VOUT+.t51 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X205 VDDA.t172 VDDA.t170 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 VDDA.t171 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X206 VOUT-.t51 two_stage_opamp_dummy_magic_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 bgr_0.PFET_GATE_10uA.t17 VDDA.t441 VDDA.t440 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X208 VOUT+.t13 two_stage_opamp_dummy_magic_0.Y.t34 VDDA.t404 VDDA.t403 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X209 VOUT-.t52 two_stage_opamp_dummy_magic_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 two_stage_opamp_dummy_magic_0.V_source.t16 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 GNDA.t35 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X211 two_stage_opamp_dummy_magic_0.VD2.t5 two_stage_opamp_dummy_magic_0.Vb1.t18 two_stage_opamp_dummy_magic_0.Y.t4 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X212 VDDA.t169 VDDA.t167 two_stage_opamp_dummy_magic_0.Vb2_2.t3 VDDA.t168 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.36 ps=2.2 w=1.8 l=0.2
X213 VDDA.t49 two_stage_opamp_dummy_magic_0.X.t32 VOUT-.t1 VDDA.t48 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X214 VOUT+.t52 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X215 bgr_0.V_TOP.t22 VDDA.t351 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 VDDA.t445 two_stage_opamp_dummy_magic_0.V_err_gate.t19 two_stage_opamp_dummy_magic_0.V_er_mir_p.t17 VDDA.t444 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X217 VOUT+.t53 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X218 VOUT-.t53 two_stage_opamp_dummy_magic_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X219 bgr_0.1st_Vout_2.t4 bgr_0.V_mir2.t18 VDDA.t75 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X220 VOUT+.t54 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X221 VOUT+.t55 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 VOUT+.t56 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 GNDA.t97 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 two_stage_opamp_dummy_magic_0.V_source.t15 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X224 VOUT-.t15 a_14240_1956.t0 GNDA.t270 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X225 bgr_0.V_mir1.t3 bgr_0.Vin-.t8 bgr_0.V_p_1.t4 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X226 bgr_0.Vin-.t4 bgr_0.V_TOP.t23 VDDA.t353 VDDA.t352 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X227 VDDA.t468 two_stage_opamp_dummy_magic_0.Vb3.t12 two_stage_opamp_dummy_magic_0.VD3.t27 VDDA.t467 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X228 two_stage_opamp_dummy_magic_0.V_err_p.t17 two_stage_opamp_dummy_magic_0.V_err_gate.t20 VDDA.t454 VDDA.t453 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X229 GNDA.t309 two_stage_opamp_dummy_magic_0.Y.t35 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 VDDA.t402 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X230 two_stage_opamp_dummy_magic_0.VD4.t29 two_stage_opamp_dummy_magic_0.VD4.t27 two_stage_opamp_dummy_magic_0.Y.t18 two_stage_opamp_dummy_magic_0.VD4.t28 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X231 a_5310_4968.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 GNDA.t320 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X232 VOUT-.t54 two_stage_opamp_dummy_magic_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X233 VOUT-.t55 two_stage_opamp_dummy_magic_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X234 VOUT-.t56 two_stage_opamp_dummy_magic_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X235 VOUT+.t57 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 VDDA.t70 bgr_0.1st_Vout_1.t17 bgr_0.V_TOP.t10 VDDA.t69 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X237 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 two_stage_opamp_dummy_magic_0.X.t33 GNDA.t282 VDDA.t363 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X238 VOUT-.t57 two_stage_opamp_dummy_magic_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 two_stage_opamp_dummy_magic_0.V_source.t2 VIN+.t2 two_stage_opamp_dummy_magic_0.VD2.t1 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X240 VOUT+.t58 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 two_stage_opamp_dummy_magic_0.V_source.t36 VIN+.t3 two_stage_opamp_dummy_magic_0.VD2.t18 GNDA.t165 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X242 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 GNDA.t237 GNDA.t238 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X243 VOUT+.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 two_stage_opamp_dummy_magic_0.V_err_p.t16 two_stage_opamp_dummy_magic_0.V_err_gate.t21 VDDA.t232 VDDA.t231 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X245 a_14680_4968.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 GNDA.t166 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X246 VOUT+.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 bgr_0.1st_Vout_2.t17 bgr_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X248 a_6810_23838.t0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 GNDA.t36 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X249 two_stage_opamp_dummy_magic_0.Vb1.t5 two_stage_opamp_dummy_magic_0.Vb1.t4 two_stage_opamp_dummy_magic_0.Vb1_2.t3 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X250 bgr_0.V_mir1.t0 bgr_0.Vin-.t9 bgr_0.V_p_1.t3 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X251 VOUT+.t61 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X252 VOUT+.t62 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 two_stage_opamp_dummy_magic_0.err_amp_out.t2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 two_stage_opamp_dummy_magic_0.V_err_p.t5 VDDA.t230 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X254 VOUT-.t58 two_stage_opamp_dummy_magic_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X255 VOUT-.t59 two_stage_opamp_dummy_magic_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 bgr_0.1st_Vout_2.t18 bgr_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X257 GNDA.t96 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 VOUT-.t7 GNDA.t95 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X258 VOUT+.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X259 VOUT+.t64 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X260 bgr_0.V_mir2.t14 bgr_0.V_mir2.t13 VDDA.t421 VDDA.t420 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X261 bgr_0.1st_Vout_1.t18 bgr_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 GNDA.t338 a_12410_22380.t1 GNDA.t337 sky130_fd_pr__res_xhigh_po_0p35 l=6
X263 two_stage_opamp_dummy_magic_0.V_err_gate.t12 two_stage_opamp_dummy_magic_0.V_tot.t7 two_stage_opamp_dummy_magic_0.V_er_mir_p.t8 VDDA.t288 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X264 VOUT-.t60 two_stage_opamp_dummy_magic_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 VOUT-.t61 two_stage_opamp_dummy_magic_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 VOUT+.t65 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X267 VOUT+.t66 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X268 VOUT-.t62 two_stage_opamp_dummy_magic_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 bgr_0.cap_res1.t0 bgr_0.V_TOP.t1 GNDA.t45 sky130_fd_pr__res_high_po_0p35 l=2.05
X270 VOUT-.t63 two_stage_opamp_dummy_magic_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 VDDA.t462 two_stage_opamp_dummy_magic_0.Vb3.t13 two_stage_opamp_dummy_magic_0.VD4.t37 VDDA.t461 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X272 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 GNDA.t279 GNDA.t278 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X273 VOUT+.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X274 VOUT+.t68 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X275 two_stage_opamp_dummy_magic_0.VD2.t2 two_stage_opamp_dummy_magic_0.Vb1.t19 two_stage_opamp_dummy_magic_0.Y.t0 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X276 bgr_0.1st_Vout_1.t19 bgr_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 two_stage_opamp_dummy_magic_0.Y.t2 two_stage_opamp_dummy_magic_0.Vb2.t16 two_stage_opamp_dummy_magic_0.VD4.t13 two_stage_opamp_dummy_magic_0.VD4.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X278 VOUT+.t12 two_stage_opamp_dummy_magic_0.Y.t36 VDDA.t401 VDDA.t400 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X279 VDDA.t64 two_stage_opamp_dummy_magic_0.X.t34 VOUT-.t4 VDDA.t63 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X280 two_stage_opamp_dummy_magic_0.VD2.t13 two_stage_opamp_dummy_magic_0.Vb1.t20 two_stage_opamp_dummy_magic_0.Y.t17 GNDA.t165 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X281 VOUT-.t64 two_stage_opamp_dummy_magic_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X282 VDDA.t283 two_stage_opamp_dummy_magic_0.X.t35 VOUT-.t9 VDDA.t282 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X283 VOUT+.t69 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 bgr_0.1st_Vout_2.t19 bgr_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X285 VDDA.t236 two_stage_opamp_dummy_magic_0.V_err_gate.t22 two_stage_opamp_dummy_magic_0.V_err_p.t15 VDDA.t235 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X286 VDDA.t166 VDDA.t164 two_stage_opamp_dummy_magic_0.err_amp_out.t1 VDDA.t165 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X287 VOUT-.t65 two_stage_opamp_dummy_magic_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X288 GNDA.t44 a_13060_22630.t0 GNDA.t43 sky130_fd_pr__res_xhigh_po_0p35 l=4
X289 VDDA.t163 VDDA.t161 two_stage_opamp_dummy_magic_0.VD3.t21 VDDA.t162 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X290 VOUT+.t70 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X291 bgr_0.PFET_GATE_10uA.t7 bgr_0.1st_Vout_2.t20 VDDA.t304 VDDA.t303 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X292 GNDA.t236 GNDA.t234 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 GNDA.t235 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X293 GNDA.t335 bgr_0.NFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_0.Vb2.t5 GNDA.t334 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X294 bgr_0.1st_Vout_1.t20 bgr_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 VIN-.t2 two_stage_opamp_dummy_magic_0.V_p_mir.t0 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X296 two_stage_opamp_dummy_magic_0.V_source.t39 VIN-.t3 two_stage_opamp_dummy_magic_0.VD1.t21 GNDA.t329 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X297 VOUT-.t66 two_stage_opamp_dummy_magic_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X298 VDDA.t160 VDDA.t158 two_stage_opamp_dummy_magic_0.V_err_gate.t7 VDDA.t159 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X299 VOUT+.t71 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 VOUT-.t67 two_stage_opamp_dummy_magic_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 VDDA.t23 bgr_0.PFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_0.Vb1.t12 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X302 two_stage_opamp_dummy_magic_0.V_er_mir_p.t16 two_stage_opamp_dummy_magic_0.V_err_gate.t23 VDDA.t425 VDDA.t424 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X303 VOUT-.t68 two_stage_opamp_dummy_magic_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 a_14560_4968.t0 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA.t92 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X305 GNDA.t302 two_stage_opamp_dummy_magic_0.Y.t37 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 VDDA.t399 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X306 VOUT+.t72 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X307 VOUT+.t73 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X308 bgr_0.1st_Vout_1.t21 bgr_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 VDDA.t345 two_stage_opamp_dummy_magic_0.Vb3.t14 two_stage_opamp_dummy_magic_0.VD4.t32 VDDA.t344 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X310 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 two_stage_opamp_dummy_magic_0.X.t36 GNDA.t158 VDDA.t281 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X311 two_stage_opamp_dummy_magic_0.V_source.t28 VIN+.t4 two_stage_opamp_dummy_magic_0.VD2.t10 GNDA.t114 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X312 two_stage_opamp_dummy_magic_0.Y.t7 two_stage_opamp_dummy_magic_0.Vb2.t17 two_stage_opamp_dummy_magic_0.VD4.t11 two_stage_opamp_dummy_magic_0.VD4.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X313 VDDA.t261 bgr_0.PFET_GATE_10uA.t19 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 VDDA.t260 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X314 VOUT+.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 VOUT-.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 VDDA.t155 VDDA.t157 VDDA.t156 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X317 VOUT-.t70 two_stage_opamp_dummy_magic_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 VOUT+.t75 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 VOUT+.t76 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 bgr_0.V_TOP.t24 VDDA.t354 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X321 VDDA.t397 two_stage_opamp_dummy_magic_0.Y.t38 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 GNDA.t317 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X322 two_stage_opamp_dummy_magic_0.Vb1.t11 GNDA.t231 GNDA.t233 GNDA.t232 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X323 two_stage_opamp_dummy_magic_0.Vb2_2.t1 two_stage_opamp_dummy_magic_0.Vb2.t1 two_stage_opamp_dummy_magic_0.Vb2.t2 two_stage_opamp_dummy_magic_0.Vb2_2.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X324 VOUT+.t77 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X325 VOUT-.t71 two_stage_opamp_dummy_magic_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X326 bgr_0.1st_Vout_2.t7 bgr_0.V_mir2.t19 VDDA.t272 VDDA.t271 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X327 VOUT-.t72 two_stage_opamp_dummy_magic_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 VOUT-.t73 two_stage_opamp_dummy_magic_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X329 VOUT-.t74 two_stage_opamp_dummy_magic_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 two_stage_opamp_dummy_magic_0.VD1.t11 two_stage_opamp_dummy_magic_0.Vb1.t21 two_stage_opamp_dummy_magic_0.X.t18 GNDA.t329 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X331 VOUT+.t78 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X332 VOUT+.t79 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X333 VOUT+.t80 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X334 VOUT+.t81 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X335 bgr_0.V_TOP.t25 VDDA.t227 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X336 two_stage_opamp_dummy_magic_0.err_amp_out.t4 GNDA.t228 GNDA.t230 GNDA.t229 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X337 VDDA.t229 bgr_0.V_TOP.t26 bgr_0.Vin-.t3 VDDA.t228 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X338 two_stage_opamp_dummy_magic_0.VD3.t19 two_stage_opamp_dummy_magic_0.Vb2.t18 two_stage_opamp_dummy_magic_0.X.t6 two_stage_opamp_dummy_magic_0.VD3.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X339 two_stage_opamp_dummy_magic_0.VD2.t8 two_stage_opamp_dummy_magic_0.Vb1.t22 two_stage_opamp_dummy_magic_0.Y.t11 GNDA.t114 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X340 bgr_0.1st_Vout_2.t21 bgr_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X341 VOUT-.t75 two_stage_opamp_dummy_magic_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X342 VOUT-.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X343 bgr_0.V_mir1.t11 bgr_0.V_mir1.t10 VDDA.t13 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X344 VOUT+.t82 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 two_stage_opamp_dummy_magic_0.V_err_p.t9 two_stage_opamp_dummy_magic_0.V_tot.t8 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 VDDA.t214 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X346 VDDA.t341 two_stage_opamp_dummy_magic_0.X.t37 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 GNDA.t271 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X347 VOUT-.t77 two_stage_opamp_dummy_magic_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X348 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 a_14240_1956.t1 GNDA.t332 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X349 bgr_0.1st_Vout_1.t22 bgr_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 GNDA.t106 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 two_stage_opamp_dummy_magic_0.err_amp_out.t9 GNDA.t105 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X351 VDDA.t320 bgr_0.PFET_GATE_10uA.t20 bgr_0.V_CUR_REF_REG.t2 VDDA.t319 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X352 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_0.Y.t23 GNDA.t325 sky130_fd_pr__res_high_po_1p41 l=1.41
X353 VOUT-.t78 two_stage_opamp_dummy_magic_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X354 bgr_0.1st_Vout_2.t22 bgr_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X355 VDDA.t347 two_stage_opamp_dummy_magic_0.Vb3.t15 two_stage_opamp_dummy_magic_0.VD4.t33 VDDA.t346 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X356 VOUT-.t79 two_stage_opamp_dummy_magic_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X357 VOUT+.t83 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X358 VOUT+.t84 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 two_stage_opamp_dummy_magic_0.V_source.t3 VIN-.t4 two_stage_opamp_dummy_magic_0.VD1.t1 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X360 VOUT+.t85 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X361 a_7460_23988.t1 a_7580_22380.t1 GNDA.t133 sky130_fd_pr__res_xhigh_po_0p35 l=6
X362 VOUT-.t80 two_stage_opamp_dummy_magic_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 bgr_0.V_p_2.t5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 bgr_0.V_mir2.t3 GNDA.t126 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X364 two_stage_opamp_dummy_magic_0.V_er_mir_p.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 two_stage_opamp_dummy_magic_0.V_err_gate.t6 VDDA.t419 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X365 a_5190_4968.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 GNDA.t130 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X366 GNDA.t318 two_stage_opamp_dummy_magic_0.Y.t39 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 VDDA.t398 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X367 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 two_stage_opamp_dummy_magic_0.X.t38 GNDA.t56 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X368 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 two_stage_opamp_dummy_magic_0.X.t39 GNDA.t30 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X369 two_stage_opamp_dummy_magic_0.V_source.t37 VIN+.t5 two_stage_opamp_dummy_magic_0.VD2.t19 GNDA.t131 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X370 bgr_0.1st_Vout_2.t23 bgr_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X371 VOUT-.t81 two_stage_opamp_dummy_magic_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 VOUT-.t82 two_stage_opamp_dummy_magic_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 a_5760_1956.t0 GNDA.t91 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X374 bgr_0.1st_Vout_1.t23 bgr_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 GNDA.t182 GNDA.t227 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X376 VDDA.t335 GNDA.t224 GNDA.t226 GNDA.t225 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X377 VOUT-.t83 two_stage_opamp_dummy_magic_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X378 bgr_0.1st_Vout_2.t24 bgr_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 bgr_0.PFET_GATE_10uA.t6 bgr_0.1st_Vout_2.t25 VDDA.t373 VDDA.t372 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X380 VDDA.t61 bgr_0.V_mir1.t19 bgr_0.1st_Vout_1.t3 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X381 VOUT-.t84 two_stage_opamp_dummy_magic_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 VDDA.t40 bgr_0.V_TOP.t27 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X383 GNDA.t331 bgr_0.NFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_0.Vb3.t4 GNDA.t330 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X384 VOUT+.t86 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X385 two_stage_opamp_dummy_magic_0.V_source.t27 two_stage_opamp_dummy_magic_0.err_amp_out.t12 GNDA.t53 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X386 GNDA.t182 GNDA.t223 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X387 VOUT-.t85 two_stage_opamp_dummy_magic_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 VDDA.t154 VDDA.t152 bgr_0.V_TOP.t3 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X389 VOUT+.t87 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X390 two_stage_opamp_dummy_magic_0.Vb3.t3 bgr_0.NFET_GATE_10uA.t14 GNDA.t88 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X391 VDDA.t151 VDDA.t149 two_stage_opamp_dummy_magic_0.V_err_p.t8 VDDA.t150 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X392 two_stage_opamp_dummy_magic_0.VD1.t10 two_stage_opamp_dummy_magic_0.Vb1.t23 two_stage_opamp_dummy_magic_0.X.t15 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X393 VOUT-.t86 two_stage_opamp_dummy_magic_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 two_stage_opamp_dummy_magic_0.VD4.t31 two_stage_opamp_dummy_magic_0.Vb3.t16 VDDA.t343 VDDA.t342 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X395 two_stage_opamp_dummy_magic_0.VD4.t9 two_stage_opamp_dummy_magic_0.Vb2.t19 two_stage_opamp_dummy_magic_0.Y.t5 two_stage_opamp_dummy_magic_0.VD4.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X396 VOUT-.t87 two_stage_opamp_dummy_magic_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X397 VOUT+.t88 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X398 GNDA.t182 GNDA.t222 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X399 VOUT+.t11 two_stage_opamp_dummy_magic_0.Y.t40 VDDA.t396 VDDA.t395 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X400 VOUT-.t88 two_stage_opamp_dummy_magic_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 bgr_0.1st_Vout_2.t8 bgr_0.V_mir2.t20 VDDA.t274 VDDA.t273 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X402 two_stage_opamp_dummy_magic_0.VD2.t11 two_stage_opamp_dummy_magic_0.Vb1.t24 two_stage_opamp_dummy_magic_0.Y.t12 GNDA.t131 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X403 VOUT+.t89 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 bgr_0.V_TOP.t9 bgr_0.1st_Vout_1.t24 VDDA.t318 VDDA.t317 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X405 GNDA.t182 GNDA.t221 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X406 GNDA.t220 GNDA.t218 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 GNDA.t219 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X407 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 two_stage_opamp_dummy_magic_0.Y.t41 VDDA.t382 GNDA.t294 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X408 VOUT-.t89 two_stage_opamp_dummy_magic_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X409 two_stage_opamp_dummy_magic_0.Vb2.t4 bgr_0.NFET_GATE_10uA.t15 GNDA.t162 GNDA.t161 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X410 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 VDDA.t143 VDDA.t145 VDDA.t144 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X411 bgr_0.START_UP_NFET1.t0 bgr_0.START_UP_NFET1.t1 GNDA.t277 GNDA.t276 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X412 VDDA.t6 two_stage_opamp_dummy_magic_0.X.t40 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X413 bgr_0.V_p_2.t10 bgr_0.V_CUR_REF_REG.t5 bgr_0.1st_Vout_2.t10 GNDA.t275 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X414 VDDA.t148 VDDA.t146 bgr_0.NFET_GATE_10uA.t0 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X415 VOUT+.t90 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 VOUT+.t91 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 bgr_0.PFET_GATE_10uA.t21 VDDA.t300 VDDA.t299 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X418 GNDA.t16 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X419 VDDA.t439 bgr_0.PFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 VDDA.t438 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X420 two_stage_opamp_dummy_magic_0.V_er_mir_p.t2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 two_stage_opamp_dummy_magic_0.V_err_gate.t5 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X421 VOUT+.t92 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X422 two_stage_opamp_dummy_magic_0.V_source.t5 VIN-.t5 two_stage_opamp_dummy_magic_0.VD1.t2 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X423 a_13180_23838.t1 bgr_0.V_CUR_REF_REG.t1 GNDA.t163 sky130_fd_pr__res_xhigh_po_0p35 l=4
X424 two_stage_opamp_dummy_magic_0.VD4.t30 two_stage_opamp_dummy_magic_0.Vb3.t17 VDDA.t302 VDDA.t301 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X425 two_stage_opamp_dummy_magic_0.V_er_mir_p.t7 two_stage_opamp_dummy_magic_0.V_tot.t9 two_stage_opamp_dummy_magic_0.V_err_gate.t11 VDDA.t209 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X426 VOUT-.t90 two_stage_opamp_dummy_magic_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 bgr_0.V_TOP.t28 VDDA.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 two_stage_opamp_dummy_magic_0.X.t24 two_stage_opamp_dummy_magic_0.VD3.t32 two_stage_opamp_dummy_magic_0.VD3.t34 two_stage_opamp_dummy_magic_0.VD3.t33 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X429 VOUT-.t91 two_stage_opamp_dummy_magic_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X430 VOUT-.t92 two_stage_opamp_dummy_magic_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 VDDA.t142 VDDA.t140 bgr_0.PFET_GATE_10uA.t2 VDDA.t141 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X432 VDDA.t10 bgr_0.V_TOP.t29 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X433 GNDA.t169 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 GNDA.t168 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X434 VOUT-.t93 two_stage_opamp_dummy_magic_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 VOUT-.t94 two_stage_opamp_dummy_magic_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 GNDA.t217 GNDA.t214 GNDA.t216 GNDA.t215 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X437 VOUT-.t95 two_stage_opamp_dummy_magic_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 GNDA.t99 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 two_stage_opamp_dummy_magic_0.V_source.t14 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X439 bgr_0.1st_Vout_1.t8 bgr_0.Vin+.t8 bgr_0.V_p_1.t8 GNDA.t291 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X440 VOUT+.t93 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 bgr_0.V_TOP.t30 VDDA.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X442 bgr_0.Vin+.t3 bgr_0.V_TOP.t31 VDDA.t244 VDDA.t243 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X443 VOUT-.t16 two_stage_opamp_dummy_magic_0.X.t41 VDDA.t362 VDDA.t361 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X444 two_stage_opamp_dummy_magic_0.V_err_p.t7 VDDA.t137 VDDA.t139 VDDA.t138 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X445 VOUT+.t94 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X446 two_stage_opamp_dummy_magic_0.Vb2_2.t6 two_stage_opamp_dummy_magic_0.Vb2_2.t4 two_stage_opamp_dummy_magic_0.Vb2_2.t6 two_stage_opamp_dummy_magic_0.Vb2_2.t5 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X447 VOUT-.t96 two_stage_opamp_dummy_magic_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X448 VOUT+.t95 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X449 bgr_0.V_mir2.t12 bgr_0.V_mir2.t11 VDDA.t234 VDDA.t233 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X450 two_stage_opamp_dummy_magic_0.VD4.t35 two_stage_opamp_dummy_magic_0.Vb3.t18 VDDA.t368 VDDA.t367 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X451 VOUT+.t96 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 VOUT-.t97 two_stage_opamp_dummy_magic_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X453 VOUT-.t98 two_stage_opamp_dummy_magic_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X454 two_stage_opamp_dummy_magic_0.V_source.t13 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 GNDA.t110 GNDA.t109 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X455 bgr_0.NFET_GATE_10uA.t2 bgr_0.NFET_GATE_10uA.t1 GNDA.t29 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X456 GNDA.t340 bgr_0.NFET_GATE_10uA.t16 two_stage_opamp_dummy_magic_0.Vb3.t2 GNDA.t339 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X457 bgr_0.V_p_2.t9 bgr_0.V_CUR_REF_REG.t6 bgr_0.1st_Vout_2.t9 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X458 VDDA.t27 two_stage_opamp_dummy_magic_0.V_err_gate.t24 two_stage_opamp_dummy_magic_0.V_err_p.t14 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X459 VOUT-.t99 two_stage_opamp_dummy_magic_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 bgr_0.V_TOP.t32 VDDA.t245 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 VDDA.t77 two_stage_opamp_dummy_magic_0.V_err_gate.t25 two_stage_opamp_dummy_magic_0.V_er_mir_p.t15 VDDA.t76 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X462 VOUT-.t100 two_stage_opamp_dummy_magic_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 two_stage_opamp_dummy_magic_0.X.t0 two_stage_opamp_dummy_magic_0.Vb2.t20 two_stage_opamp_dummy_magic_0.VD3.t17 two_stage_opamp_dummy_magic_0.VD3.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X464 two_stage_opamp_dummy_magic_0.VD1.t9 two_stage_opamp_dummy_magic_0.Vb1.t25 two_stage_opamp_dummy_magic_0.X.t16 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X465 bgr_0.1st_Vout_1.t2 bgr_0.V_mir1.t20 VDDA.t87 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X466 VDDA.t249 bgr_0.V_TOP.t33 bgr_0.Vin-.t2 VDDA.t248 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X467 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 VDDA.t134 VDDA.t136 VDDA.t135 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X468 VOUT-.t101 two_stage_opamp_dummy_magic_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X469 VOUT+.t97 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 bgr_0.PFET_GATE_10uA.t23 VDDA.t456 VDDA.t455 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X471 VOUT+.t98 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 VDDA.t259 bgr_0.PFET_GATE_10uA.t24 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 VDDA.t258 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X473 VOUT+.t2 VDDA.t131 VDDA.t133 VDDA.t132 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X474 VOUT+.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X475 VOUT+.t100 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X476 VOUT+.t101 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X477 bgr_0.1st_Vout_1.t25 bgr_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X478 VOUT-.t102 two_stage_opamp_dummy_magic_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X479 bgr_0.1st_Vout_2.t26 bgr_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X480 two_stage_opamp_dummy_magic_0.V_err_p.t4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 two_stage_opamp_dummy_magic_0.err_amp_out.t0 VDDA.t71 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X481 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 two_stage_opamp_dummy_magic_0.Y.t42 VDDA.t390 GNDA.t82 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X482 GNDA.t213 GNDA.t211 VDDA.t334 GNDA.t212 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X483 two_stage_opamp_dummy_magic_0.VD4.t36 two_stage_opamp_dummy_magic_0.Vb3.t19 VDDA.t449 VDDA.t448 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X484 VOUT+.t102 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X485 VOUT+.t17 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 GNDA.t322 GNDA.t321 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X486 bgr_0.V_p_2.t0 bgr_0.V_CUR_REF_REG.t7 bgr_0.1st_Vout_2.t0 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X487 VDDA.t223 two_stage_opamp_dummy_magic_0.X.t42 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA.t117 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X488 GNDA.t108 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 two_stage_opamp_dummy_magic_0.err_amp_out.t8 GNDA.t107 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X489 bgr_0.1st_Vout_1.t26 bgr_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 bgr_0.START_UP.t5 bgr_0.V_TOP.t34 VDDA.t251 VDDA.t250 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X491 VOUT-.t103 two_stage_opamp_dummy_magic_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X492 VOUT-.t104 two_stage_opamp_dummy_magic_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 VOUT-.t105 two_stage_opamp_dummy_magic_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X494 bgr_0.V_TOP.t8 bgr_0.1st_Vout_1.t27 VDDA.t57 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X495 two_stage_opamp_dummy_magic_0.V_er_mir_p.t6 two_stage_opamp_dummy_magic_0.V_tot.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t13 VDDA.t432 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X496 two_stage_opamp_dummy_magic_0.V_source.t30 VIN-.t6 two_stage_opamp_dummy_magic_0.VD1.t15 GNDA.t84 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X497 VOUT-.t106 two_stage_opamp_dummy_magic_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 GNDA.t83 two_stage_opamp_dummy_magic_0.Y.t43 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 VDDA.t394 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X499 VOUT+.t103 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X500 two_stage_opamp_dummy_magic_0.Vb2.t10 GNDA.t208 GNDA.t210 GNDA.t209 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X501 VOUT+.t104 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X502 VDDA.t393 two_stage_opamp_dummy_magic_0.Y.t44 VOUT+.t10 VDDA.t392 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X503 GNDA.t112 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 two_stage_opamp_dummy_magic_0.V_source.t12 GNDA.t111 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X504 VOUT+.t105 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X505 bgr_0.1st_Vout_1.t28 bgr_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X506 VOUT+.t18 a_5760_1956.t1 GNDA.t327 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X507 bgr_0.1st_Vout_2.t27 bgr_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X508 bgr_0.V_TOP.t7 bgr_0.1st_Vout_1.t29 VDDA.t370 VDDA.t369 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X509 VOUT-.t12 two_stage_opamp_dummy_magic_0.X.t43 VDDA.t326 VDDA.t325 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X510 two_stage_opamp_dummy_magic_0.V_er_mir_p.t14 two_stage_opamp_dummy_magic_0.V_err_gate.t26 VDDA.t278 VDDA.t277 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X511 VOUT+.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X512 two_stage_opamp_dummy_magic_0.X.t8 two_stage_opamp_dummy_magic_0.Vb2.t21 two_stage_opamp_dummy_magic_0.VD3.t15 two_stage_opamp_dummy_magic_0.VD3.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X513 VOUT+.t107 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X514 bgr_0.1st_Vout_1.t30 bgr_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X515 VOUT-.t107 two_stage_opamp_dummy_magic_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X516 two_stage_opamp_dummy_magic_0.V_source.t11 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 GNDA.t65 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X517 VDDA.t466 two_stage_opamp_dummy_magic_0.Vb3.t20 two_stage_opamp_dummy_magic_0.VD3.t26 VDDA.t465 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X518 VOUT-.t108 two_stage_opamp_dummy_magic_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X519 VDDA.t8 two_stage_opamp_dummy_magic_0.Vb3.t21 two_stage_opamp_dummy_magic_0.VD4.t1 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X520 VOUT-.t109 two_stage_opamp_dummy_magic_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X521 two_stage_opamp_dummy_magic_0.VD1.t16 VIN-.t7 two_stage_opamp_dummy_magic_0.V_source.t31 GNDA.t164 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X522 VDDA.t265 two_stage_opamp_dummy_magic_0.V_err_gate.t27 two_stage_opamp_dummy_magic_0.V_er_mir_p.t13 VDDA.t264 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X523 VOUT+.t108 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X524 VOUT+.t109 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 VOUT-.t110 two_stage_opamp_dummy_magic_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X526 VOUT+.t110 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X527 VOUT+.t111 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 VOUT+.t112 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X529 bgr_0.1st_Vout_1.t31 bgr_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X530 VOUT+.t113 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X531 two_stage_opamp_dummy_magic_0.VD1.t8 two_stage_opamp_dummy_magic_0.Vb1.t26 two_stage_opamp_dummy_magic_0.X.t19 GNDA.t84 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X532 bgr_0.V_mir1.t9 bgr_0.V_mir1.t8 VDDA.t38 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X533 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0 ps=0 w=3.5 l=0.2
X534 GNDA.t116 two_stage_opamp_dummy_magic_0.X.t44 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 VDDA.t222 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X535 two_stage_opamp_dummy_magic_0.VD2.t17 VIN+.t6 two_stage_opamp_dummy_magic_0.V_source.t35 GNDA.t72 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X536 VOUT-.t111 two_stage_opamp_dummy_magic_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X537 VOUT+.t114 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X538 VOUT+.t115 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X539 VOUT-.t112 two_stage_opamp_dummy_magic_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X540 VOUT-.t113 two_stage_opamp_dummy_magic_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X541 GNDA.t8 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 VOUT-.t0 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X542 GNDA.t182 GNDA.t207 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X543 GNDA.t180 GNDA.t178 two_stage_opamp_dummy_magic_0.Vb1.t10 GNDA.t179 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X544 two_stage_opamp_dummy_magic_0.V_err_p.t21 two_stage_opamp_dummy_magic_0.V_tot.t11 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 VDDA.t416 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X545 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 two_stage_opamp_dummy_magic_0.Y.t45 VDDA.t391 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X546 VDDA.t429 two_stage_opamp_dummy_magic_0.X.t45 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA.t324 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X547 GNDA.t152 bgr_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 GNDA.t151 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X548 two_stage_opamp_dummy_magic_0.cap_res_X.t0 two_stage_opamp_dummy_magic_0.X.t11 GNDA.t129 sky130_fd_pr__res_high_po_1p41 l=1.41
X549 GNDA.t142 bgr_0.NFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 GNDA.t141 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X550 VDDA.t431 two_stage_opamp_dummy_magic_0.X.t46 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 GNDA.t328 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X551 VOUT+.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X552 two_stage_opamp_dummy_magic_0.Vb2.t3 bgr_0.NFET_GATE_10uA.t19 GNDA.t316 GNDA.t315 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X553 VOUT-.t114 two_stage_opamp_dummy_magic_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X554 VOUT+.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X555 VOUT+.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X556 VDDA.t253 bgr_0.V_mir2.t21 bgr_0.1st_Vout_2.t5 VDDA.t252 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X557 VOUT-.t115 two_stage_opamp_dummy_magic_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X558 bgr_0.1st_Vout_2.t28 bgr_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X559 two_stage_opamp_dummy_magic_0.VD3.t13 two_stage_opamp_dummy_magic_0.Vb2.t22 two_stage_opamp_dummy_magic_0.X.t4 two_stage_opamp_dummy_magic_0.VD3.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X560 two_stage_opamp_dummy_magic_0.V_er_mir_p.t1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 two_stage_opamp_dummy_magic_0.V_err_gate.t4 VDDA.t270 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X561 VDDA.t130 VDDA.t128 two_stage_opamp_dummy_magic_0.Vb1.t1 VDDA.t129 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X562 two_stage_opamp_dummy_magic_0.X.t20 two_stage_opamp_dummy_magic_0.Vb1.t27 two_stage_opamp_dummy_magic_0.VD1.t7 GNDA.t164 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X563 VOUT+.t119 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X564 bgr_0.V_p_1.t2 bgr_0.Vin-.t10 bgr_0.V_mir1.t16 GNDA.t148 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X565 two_stage_opamp_dummy_magic_0.Vb1.t0 VDDA.t125 VDDA.t127 VDDA.t126 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X566 GNDA.t145 VDDA.t122 VDDA.t124 VDDA.t123 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X567 VOUT-.t116 two_stage_opamp_dummy_magic_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X568 VOUT-.t117 two_stage_opamp_dummy_magic_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X569 GNDA.t206 GNDA.t204 VOUT-.t14 GNDA.t205 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X570 GNDA.t182 GNDA.t194 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X571 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 VDDA.t119 VDDA.t121 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X572 bgr_0.1st_Vout_2.t29 bgr_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X573 bgr_0.PFET_GATE_10uA.t1 VDDA.t116 VDDA.t118 VDDA.t117 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X574 VDDA.t389 two_stage_opamp_dummy_magic_0.Y.t46 VOUT+.t9 VDDA.t388 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X575 VOUT-.t118 two_stage_opamp_dummy_magic_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X576 VOUT-.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X577 GNDA.t67 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 two_stage_opamp_dummy_magic_0.V_source.t10 GNDA.t66 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X578 VDDA.t115 VDDA.t113 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 VDDA.t114 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X579 VDDA.t112 VDDA.t110 VOUT+.t1 VDDA.t111 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X580 VOUT+.t120 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X581 bgr_0.1st_Vout_1.t1 bgr_0.V_mir1.t21 VDDA.t89 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X582 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 bgr_0.PFET_GATE_10uA.t25 VDDA.t211 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X583 two_stage_opamp_dummy_magic_0.Y.t9 two_stage_opamp_dummy_magic_0.Vb1.t28 two_stage_opamp_dummy_magic_0.VD2.t6 GNDA.t72 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X584 VOUT-.t3 two_stage_opamp_dummy_magic_0.X.t47 VDDA.t55 VDDA.t54 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X585 VDDA.t4 two_stage_opamp_dummy_magic_0.Vb3.t22 two_stage_opamp_dummy_magic_0.VD4.t0 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X586 VOUT-.t120 two_stage_opamp_dummy_magic_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X587 VOUT+.t121 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X588 GNDA.t24 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 VOUT+.t0 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X589 two_stage_opamp_dummy_magic_0.V_err_p.t13 two_stage_opamp_dummy_magic_0.V_err_gate.t28 VDDA.t340 VDDA.t339 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X590 bgr_0.1st_Vout_1.t32 bgr_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X591 GNDA.t203 GNDA.t202 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X592 VOUT+.t122 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X593 a_6810_23838.t1 a_6930_22564.t1 GNDA.t36 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X594 VOUT-.t121 two_stage_opamp_dummy_magic_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X595 VOUT+.t123 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X596 GNDA.t182 GNDA.t201 bgr_0.Vin-.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X597 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 two_stage_opamp_dummy_magic_0.Vb3.t6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X598 VOUT+.t124 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X599 bgr_0.1st_Vout_2.t30 bgr_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X600 two_stage_opamp_dummy_magic_0.V_source.t9 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 GNDA.t79 GNDA.t78 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X601 bgr_0.V_p_1.t1 bgr_0.Vin-.t11 bgr_0.V_mir1.t1 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X602 two_stage_opamp_dummy_magic_0.VD3.t11 two_stage_opamp_dummy_magic_0.Vb2.t23 two_stage_opamp_dummy_magic_0.X.t9 two_stage_opamp_dummy_magic_0.VD3.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X603 VDDA.t296 two_stage_opamp_dummy_magic_0.V_err_gate.t29 two_stage_opamp_dummy_magic_0.V_err_p.t12 VDDA.t295 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X604 two_stage_opamp_dummy_magic_0.VD3.t25 two_stage_opamp_dummy_magic_0.Vb3.t23 VDDA.t290 VDDA.t289 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X605 VOUT+.t125 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X606 two_stage_opamp_dummy_magic_0.Y.t19 two_stage_opamp_dummy_magic_0.Vb2.t24 two_stage_opamp_dummy_magic_0.VD4.t7 two_stage_opamp_dummy_magic_0.VD4.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X607 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 two_stage_opamp_dummy_magic_0.Y.t47 GNDA.t301 VDDA.t387 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X608 a_12530_23988.t1 a_12410_22380.t0 GNDA.t319 sky130_fd_pr__res_xhigh_po_0p35 l=6
X609 VDDA.t452 bgr_0.V_mir2.t9 bgr_0.V_mir2.t10 VDDA.t451 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X610 bgr_0.1st_Vout_2.t31 bgr_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X611 GNDA.t285 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 VOUT+.t6 GNDA.t284 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X612 GNDA.t75 two_stage_opamp_dummy_magic_0.X.t48 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 VDDA.t80 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X613 two_stage_opamp_dummy_magic_0.V_source.t8 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 GNDA.t81 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X614 two_stage_opamp_dummy_magic_0.VD2.t21 VIN+.t7 two_stage_opamp_dummy_magic_0.V_source.t40 GNDA.t157 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X615 VOUT-.t122 two_stage_opamp_dummy_magic_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X616 bgr_0.V_p_2.t4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 bgr_0.V_mir2.t2 GNDA.t143 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X617 VDDA.t109 VDDA.t107 two_stage_opamp_dummy_magic_0.VD4.t22 VDDA.t108 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X618 VOUT+.t126 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X619 bgr_0.1st_Vout_1.t33 bgr_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X620 VDDA.t25 two_stage_opamp_dummy_magic_0.V_err_gate.t30 two_stage_opamp_dummy_magic_0.V_err_p.t11 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X621 bgr_0.1st_Vout_2.t32 bgr_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X622 VOUT-.t123 two_stage_opamp_dummy_magic_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X623 two_stage_opamp_dummy_magic_0.VD3.t9 two_stage_opamp_dummy_magic_0.Vb2.t25 two_stage_opamp_dummy_magic_0.X.t3 two_stage_opamp_dummy_magic_0.VD3.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X624 two_stage_opamp_dummy_magic_0.Vb1_2.t2 two_stage_opamp_dummy_magic_0.Vb1.t6 two_stage_opamp_dummy_magic_0.Vb1.t7 GNDA.t336 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X625 VOUT+.t127 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X626 two_stage_opamp_dummy_magic_0.VD3.t20 VDDA.t104 VDDA.t106 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X627 two_stage_opamp_dummy_magic_0.V_err_p.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 two_stage_opamp_dummy_magic_0.err_amp_out.t5 VDDA.t336 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X628 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 two_stage_opamp_dummy_magic_0.Y.t48 VDDA.t386 GNDA.t298 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X629 VDDA.t333 GNDA.t198 GNDA.t200 GNDA.t199 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X630 VOUT-.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X631 VOUT-.t125 two_stage_opamp_dummy_magic_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X632 a_13180_23838.t0 a_13060_22630.t1 GNDA.t100 sky130_fd_pr__res_xhigh_po_0p35 l=4
X633 bgr_0.V_CUR_REF_REG.t0 VDDA.t101 VDDA.t103 VDDA.t102 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X634 VOUT+.t128 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X635 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 bgr_0.PFET_GATE_10uA.t26 VDDA.t218 VDDA.t217 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X636 VDDA.t356 bgr_0.1st_Vout_2.t33 bgr_0.PFET_GATE_10uA.t5 VDDA.t355 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X637 two_stage_opamp_dummy_magic_0.V_er_mir_p.t12 two_stage_opamp_dummy_magic_0.V_err_gate.t31 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X638 bgr_0.V_p_1.t0 bgr_0.Vin-.t12 bgr_0.V_mir1.t2 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X639 bgr_0.START_UP.t4 bgr_0.V_TOP.t35 VDDA.t330 VDDA.t329 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X640 bgr_0.V_TOP.t36 VDDA.t331 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X641 VOUT-.t126 two_stage_opamp_dummy_magic_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X642 VOUT-.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X643 VOUT-.t128 two_stage_opamp_dummy_magic_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X644 VOUT+.t129 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X645 GNDA.t273 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 two_stage_opamp_dummy_magic_0.V_p_mir.t1 GNDA.t272 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X646 VDDA.t385 two_stage_opamp_dummy_magic_0.Y.t49 VOUT+.t8 VDDA.t384 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X647 VOUT-.t11 two_stage_opamp_dummy_magic_0.X.t49 VDDA.t324 VDDA.t323 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X648 VOUT-.t129 two_stage_opamp_dummy_magic_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X649 VOUT-.t13 GNDA.t195 GNDA.t197 GNDA.t196 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X650 two_stage_opamp_dummy_magic_0.Y.t15 two_stage_opamp_dummy_magic_0.Vb1.t29 two_stage_opamp_dummy_magic_0.VD2.t12 GNDA.t157 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X651 VOUT-.t10 two_stage_opamp_dummy_magic_0.X.t50 VDDA.t322 VDDA.t321 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X652 two_stage_opamp_dummy_magic_0.VD3.t7 two_stage_opamp_dummy_magic_0.Vb2.t26 two_stage_opamp_dummy_magic_0.X.t7 two_stage_opamp_dummy_magic_0.VD3.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X653 two_stage_opamp_dummy_magic_0.V_er_mir_p.t11 two_stage_opamp_dummy_magic_0.V_err_gate.t32 VDDA.t294 VDDA.t293 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X654 VOUT+.t130 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X655 VOUT+.t131 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X656 two_stage_opamp_dummy_magic_0.VD3.t24 two_stage_opamp_dummy_magic_0.Vb3.t24 VDDA.t30 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X657 bgr_0.V_TOP.t37 VDDA.t224 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X658 VDDA.t226 bgr_0.V_TOP.t38 bgr_0.Vin+.t2 VDDA.t225 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X659 VOUT-.t130 two_stage_opamp_dummy_magic_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X660 bgr_0.Vin-.t1 bgr_0.START_UP.t6 bgr_0.V_TOP.t0 VDDA.t52 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X661 VOUT-.t131 two_stage_opamp_dummy_magic_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X662 two_stage_opamp_dummy_magic_0.Vb3.t7 GNDA.t191 GNDA.t193 GNDA.t192 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X663 two_stage_opamp_dummy_magic_0.V_source.t7 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 GNDA.t274 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X664 bgr_0.V_TOP.t39 VDDA.t327 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X665 bgr_0.1st_Vout_1.t0 bgr_0.V_mir1.t22 VDDA.t349 VDDA.t348 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X666 bgr_0.V_TOP.t13 bgr_0.START_UP.t7 bgr_0.Vin-.t0 VDDA.t305 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X667 two_stage_opamp_dummy_magic_0.VD1.t4 VIN-.t8 two_stage_opamp_dummy_magic_0.V_source.t25 GNDA.t86 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X668 GNDA.t190 GNDA.t189 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 GNDA.t78 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X669 two_stage_opamp_dummy_magic_0.Vb3.t0 two_stage_opamp_dummy_magic_0.Vb2.t27 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X670 bgr_0.V_TOP.t40 VDDA.t328 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X671 VDDA.t423 two_stage_opamp_dummy_magic_0.V_err_gate.t33 two_stage_opamp_dummy_magic_0.V_er_mir_p.t10 VDDA.t422 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X672 VOUT-.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X673 VOUT-.t133 two_stage_opamp_dummy_magic_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X674 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 two_stage_opamp_dummy_magic_0.Y.t50 GNDA.t297 VDDA.t383 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X675 VOUT-.t134 two_stage_opamp_dummy_magic_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X676 VDDA.t100 VDDA.t98 GNDA.t170 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X677 VOUT+.t132 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X678 VOUT-.t135 two_stage_opamp_dummy_magic_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X679 VOUT-.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X680 GNDA.t115 two_stage_opamp_dummy_magic_0.X.t51 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 VDDA.t221 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X681 two_stage_opamp_dummy_magic_0.VD2.t0 VIN+.t8 two_stage_opamp_dummy_magic_0.V_source.t1 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X682 bgr_0.V_p_1.t5 VDDA.t471 GNDA.t61 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X683 VOUT+.t133 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X684 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 bgr_0.NFET_GATE_10uA.t20 GNDA.t90 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X685 bgr_0.Vin+.t0 bgr_0.V_TOP.t41 VDDA.t33 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X686 bgr_0.V_TOP.t42 VDDA.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X687 GNDA.t160 bgr_0.NFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X688 two_stage_opamp_dummy_magic_0.Vb1_2.t1 two_stage_opamp_dummy_magic_0.Vb1.t8 two_stage_opamp_dummy_magic_0.Vb1.t9 GNDA.t333 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X689 VDDA.t435 bgr_0.V_mir2.t7 bgr_0.V_mir2.t8 VDDA.t434 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X690 VDDA.t287 bgr_0.V_mir1.t6 bgr_0.V_mir1.t7 VDDA.t286 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X691 VDDA.t82 bgr_0.V_TOP.t43 bgr_0.Vin+.t1 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X692 bgr_0.V_p_1.t7 bgr_0.Vin+.t9 bgr_0.1st_Vout_1.t9 GNDA.t290 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X693 two_stage_opamp_dummy_magic_0.V_err_p.t0 two_stage_opamp_dummy_magic_0.V_tot.t12 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X694 bgr_0.NFET_GATE_10uA.t4 bgr_0.PFET_GATE_10uA.t27 VDDA.t437 VDDA.t436 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X695 two_stage_opamp_dummy_magic_0.X.t2 two_stage_opamp_dummy_magic_0.Vb2.t28 two_stage_opamp_dummy_magic_0.VD3.t5 two_stage_opamp_dummy_magic_0.VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X696 VDDA.t21 bgr_0.PFET_GATE_10uA.t28 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X697 bgr_0.V_TOP.t44 VDDA.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X698 VOUT-.t137 two_stage_opamp_dummy_magic_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X699 two_stage_opamp_dummy_magic_0.VD4.t5 two_stage_opamp_dummy_magic_0.Vb2.t29 two_stage_opamp_dummy_magic_0.Y.t3 two_stage_opamp_dummy_magic_0.VD4.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X700 VOUT-.t138 two_stage_opamp_dummy_magic_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X701 two_stage_opamp_dummy_magic_0.X.t21 two_stage_opamp_dummy_magic_0.Vb1.t30 two_stage_opamp_dummy_magic_0.VD1.t6 GNDA.t86 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X702 VDDA.t15 two_stage_opamp_dummy_magic_0.Vb3.t25 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X703 VOUT-.t139 two_stage_opamp_dummy_magic_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X704 bgr_0.V_TOP.t2 VDDA.t95 VDDA.t97 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X705 VOUT+.t134 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X706 VOUT+.t135 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X707 VOUT+.t136 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X708 two_stage_opamp_dummy_magic_0.VD4.t34 two_stage_opamp_dummy_magic_0.Vb3.t26 VDDA.t360 VDDA.t359 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X709 GNDA.t102 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 two_stage_opamp_dummy_magic_0.err_amp_out.t7 GNDA.t101 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X710 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 bgr_0.V_TOP.t45 VDDA.t310 VDDA.t309 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X711 bgr_0.1st_Vout_1.t34 bgr_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X712 VDDA.t381 two_stage_opamp_dummy_magic_0.Y.t51 VOUT+.t7 VDDA.t380 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X713 two_stage_opamp_dummy_magic_0.Y.t24 two_stage_opamp_dummy_magic_0.Vb1.t31 two_stage_opamp_dummy_magic_0.VD2.t20 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X714 VOUT-.t5 VDDA.t92 VDDA.t94 VDDA.t93 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X715 VOUT-.t140 two_stage_opamp_dummy_magic_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X716 bgr_0.V_p_1.t6 bgr_0.Vin+.t10 bgr_0.1st_Vout_1.t6 GNDA.t289 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X717 VOUT+.t137 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X718 two_stage_opamp_dummy_magic_0.err_amp_out.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 two_stage_opamp_dummy_magic_0.V_err_p.t2 VDDA.t292 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X719 GNDA.t188 GNDA.t186 VDDA.t332 GNDA.t187 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X720 VOUT+.t138 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X721 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 GNDA.t51 GNDA.t50 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X722 VOUT-.t141 two_stage_opamp_dummy_magic_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X723 GNDA.t150 bgr_0.NFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_0.V_err_gate.t9 GNDA.t149 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X724 VDDA.t358 bgr_0.1st_Vout_2.t34 bgr_0.PFET_GATE_10uA.t4 VDDA.t357 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X725 two_stage_opamp_dummy_magic_0.Vb3.t1 bgr_0.NFET_GATE_10uA.t23 GNDA.t269 GNDA.t268 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X726 bgr_0.V_mir1.t5 bgr_0.V_mir1.t4 VDDA.t418 VDDA.t417 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X727 two_stage_opamp_dummy_magic_0.VD4.t3 two_stage_opamp_dummy_magic_0.Vb2.t30 two_stage_opamp_dummy_magic_0.Y.t13 two_stage_opamp_dummy_magic_0.VD4.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X728 two_stage_opamp_dummy_magic_0.V_p_mir.t3 VIN+.t9 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X729 two_stage_opamp_dummy_magic_0.VD1.t0 VIN-.t9 two_stage_opamp_dummy_magic_0.V_source.t0 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X730 VOUT-.t142 two_stage_opamp_dummy_magic_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X731 GNDA.t185 GNDA.t183 two_stage_opamp_dummy_magic_0.Vb2.t9 GNDA.t184 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X732 two_stage_opamp_dummy_magic_0.V_err_gate.t1 two_stage_opamp_dummy_magic_0.V_tot.t13 two_stage_opamp_dummy_magic_0.V_er_mir_p.t5 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X733 VOUT+.t139 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X734 VOUT+.t140 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X735 VOUT+.t141 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X736 VDDA.t312 bgr_0.V_TOP.t46 bgr_0.START_UP.t3 VDDA.t311 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X737 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 two_stage_opamp_dummy_magic_0.Y.t52 GNDA.t310 VDDA.t379 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X738 GNDA.t74 two_stage_opamp_dummy_magic_0.X.t52 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X739 VOUT+.t142 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X740 VOUT+.t143 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X741 bgr_0.1st_Vout_1.t35 bgr_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X742 bgr_0.1st_Vout_2.t35 bgr_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X743 GNDA.t73 two_stage_opamp_dummy_magic_0.X.t53 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 VDDA.t78 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X744 VOUT-.t143 two_stage_opamp_dummy_magic_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X745 VDDA.t257 bgr_0.PFET_GATE_10uA.t29 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 VDDA.t256 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X746 two_stage_opamp_dummy_magic_0.VD2.t14 VIN+.t10 two_stage_opamp_dummy_magic_0.V_source.t32 GNDA.t113 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X747 two_stage_opamp_dummy_magic_0.X.t1 two_stage_opamp_dummy_magic_0.Vb2.t31 two_stage_opamp_dummy_magic_0.VD3.t3 two_stage_opamp_dummy_magic_0.VD3.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X748 VOUT-.t144 two_stage_opamp_dummy_magic_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X749 GNDA.t182 GNDA.t181 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X750 VDDA.t208 two_stage_opamp_dummy_magic_0.Vb3.t27 two_stage_opamp_dummy_magic_0.VD3.t23 VDDA.t207 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X751 VOUT-.t145 two_stage_opamp_dummy_magic_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X752 VDDA.t255 bgr_0.V_mir2.t22 bgr_0.1st_Vout_2.t6 VDDA.t254 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X753 VOUT+.t144 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X754 bgr_0.1st_Vout_1.t36 bgr_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X755 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 two_stage_opamp_dummy_magic_0.Y.t53 VDDA.t377 GNDA.t311 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X756 VOUT-.t146 two_stage_opamp_dummy_magic_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X757 bgr_0.V_TOP.t47 VDDA.t306 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X758 GNDA.t177 GNDA.t175 two_stage_opamp_dummy_magic_0.V_source.t34 GNDA.t176 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X759 VOUT-.t147 two_stage_opamp_dummy_magic_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X760 bgr_0.V_mir2.t1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 bgr_0.V_p_2.t3 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X761 VOUT+.t145 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X762 VOUT+.t146 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X763 VOUT+.t147 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X764 VOUT-.t148 two_stage_opamp_dummy_magic_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X765 VOUT-.t149 two_stage_opamp_dummy_magic_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X766 bgr_0.PFET_GATE_10uA.t3 VDDA.t472 GNDA.t39 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X767 two_stage_opamp_dummy_magic_0.X.t12 two_stage_opamp_dummy_magic_0.Vb1.t32 two_stage_opamp_dummy_magic_0.VD1.t5 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X768 VOUT+.t148 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X769 two_stage_opamp_dummy_magic_0.V_source.t29 two_stage_opamp_dummy_magic_0.Vb1.t33 two_stage_opamp_dummy_magic_0.Vb1_2.t0 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.6 ps=3.8 w=1.5 l=3
X770 two_stage_opamp_dummy_magic_0.Y.t14 two_stage_opamp_dummy_magic_0.VD4.t24 two_stage_opamp_dummy_magic_0.VD4.t26 two_stage_opamp_dummy_magic_0.VD4.t25 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X771 VOUT+.t149 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X772 VOUT-.t150 two_stage_opamp_dummy_magic_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X773 VOUT+.t150 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X774 two_stage_opamp_dummy_magic_0.X.t5 two_stage_opamp_dummy_magic_0.Vb2.t32 two_stage_opamp_dummy_magic_0.VD3.t1 two_stage_opamp_dummy_magic_0.VD3.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X775 VOUT-.t151 two_stage_opamp_dummy_magic_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X776 two_stage_opamp_dummy_magic_0.Y.t10 two_stage_opamp_dummy_magic_0.Vb1.t34 two_stage_opamp_dummy_magic_0.VD2.t7 GNDA.t113 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X777 VDDA.t427 two_stage_opamp_dummy_magic_0.Vb3.t28 two_stage_opamp_dummy_magic_0.VD3.t22 VDDA.t426 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X778 VOUT+.t151 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X779 VOUT-.t152 two_stage_opamp_dummy_magic_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X780 VOUT-.t153 two_stage_opamp_dummy_magic_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X781 VDDA.t378 two_stage_opamp_dummy_magic_0.Y.t54 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 GNDA.t314 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X782 VDDA.t308 bgr_0.V_TOP.t48 bgr_0.START_UP.t2 VDDA.t307 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X783 VOUT+.t152 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X784 bgr_0.V_TOP.t49 VDDA.t371 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X785 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 two_stage_opamp_dummy_magic_0.X.t54 VDDA.t28 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X786 VOUT+.t153 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X787 VDDA.t464 bgr_0.V_mir2.t5 bgr_0.V_mir2.t6 VDDA.t463 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X788 two_stage_opamp_dummy_magic_0.err_amp_out.t6 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 GNDA.t104 GNDA.t103 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X789 VOUT+.t154 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X790 VOUT-.t154 two_stage_opamp_dummy_magic_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X791 VOUT-.t155 two_stage_opamp_dummy_magic_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X792 bgr_0.1st_Vout_2.t36 bgr_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X793 VOUT+.t155 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X794 two_stage_opamp_dummy_magic_0.VD1.t18 GNDA.t172 GNDA.t174 GNDA.t173 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X795 VOUT+.t156 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X796 two_stage_opamp_dummy_magic_0.V_err_gate.t2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 two_stage_opamp_dummy_magic_0.V_er_mir_p.t0 VDDA.t291 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X797 two_stage_opamp_dummy_magic_0.VD1.t3 VIN-.t10 two_stage_opamp_dummy_magic_0.V_source.t6 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X798 bgr_0.V_mir2.t0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 bgr_0.V_p_2.t7 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X799 VOUT-.t156 two_stage_opamp_dummy_magic_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 bgr_0.Vin+.n1 bgr_0.Vin+.n0 514.134
R1 bgr_0.Vin+.n3 bgr_0.Vin+.n2 514.134
R2 bgr_0.Vin+.n4 bgr_0.Vin+.n3 402.817
R3 bgr_0.Vin+.n0 bgr_0.Vin+.t8 303.259
R4 bgr_0.Vin+.n0 bgr_0.Vin+.t9 174.726
R5 bgr_0.Vin+.n1 bgr_0.Vin+.t6 174.726
R6 bgr_0.Vin+.n2 bgr_0.Vin+.t10 174.726
R7 bgr_0.Vin+.n3 bgr_0.Vin+.t7 174.726
R8 bgr_0.Vin+.n10 bgr_0.Vin+.t5 158.989
R9 bgr_0.Vin+.n2 bgr_0.Vin+.n1 128.534
R10 bgr_0.Vin+.t4 bgr_0.Vin+.n10 118.754
R11 bgr_0.Vin+.n6 bgr_0.Vin+.n5 74.288
R12 bgr_0.Vin+.n8 bgr_0.Vin+.n7 74.288
R13 bgr_0.Vin+.n10 bgr_0.Vin+.n9 35.5943
R14 bgr_0.Vin+.n8 bgr_0.Vin+.n6 14.1255
R15 bgr_0.Vin+.n5 bgr_0.Vin+.t2 13.1338
R16 bgr_0.Vin+.n5 bgr_0.Vin+.t0 13.1338
R17 bgr_0.Vin+.n7 bgr_0.Vin+.t1 13.1338
R18 bgr_0.Vin+.n7 bgr_0.Vin+.t3 13.1338
R19 bgr_0.Vin+.n9 bgr_0.Vin+.n8 5.188
R20 bgr_0.Vin+.n6 bgr_0.Vin+.n4 5.188
R21 bgr_0.Vin+.n9 bgr_0.Vin+.n4 2.1255
R22 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 807.99
R23 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 195.296
R24 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n142 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 84.0884
R25 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 83.5719
R26 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 83.5719
R27 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 83.5719
R28 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 83.5719
R29 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 83.5719
R30 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 83.5719
R31 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 83.5719
R32 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 83.5719
R33 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 83.5719
R34 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 83.5719
R35 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 83.5719
R36 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 83.5719
R37 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 83.5719
R38 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 83.5719
R39 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 83.5719
R40 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 83.5719
R41 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 83.5719
R42 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 83.5719
R43 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 83.5719
R44 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 83.5719
R45 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 83.5719
R46 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R47 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 83.5719
R48 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 73.8495
R49 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 73.8495
R50 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 73.3165
R51 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 73.3165
R52 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 73.3165
R53 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 73.3165
R54 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 73.3165
R55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 73.19
R56 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 73.19
R57 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 73.19
R58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 73.19
R59 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 73.19
R60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 73.19
R61 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 65.0299
R62 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 65.0299
R63 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 26.074
R64 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 26.074
R65 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 26.074
R66 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 26.074
R67 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 26.074
R68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 26.074
R69 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 26.074
R70 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 26.074
R71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 26.074
R72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 26.074
R73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 25.7843
R74 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 25.7843
R75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 25.7843
R76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 25.7843
R77 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 25.7843
R78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 25.7843
R79 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 9.3005
R80 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R81 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 9.3005
R82 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R83 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 9.3005
R84 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R85 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 9.3005
R86 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R87 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 9.3005
R88 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R89 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 9.3005
R90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R91 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 9.3005
R92 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 9.3005
R93 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 9.3005
R94 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 9.3005
R95 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R96 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 9.3005
R97 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 9.3005
R98 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 9.3005
R99 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R100 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 9.3005
R101 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 9.3005
R102 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R103 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 9.3005
R104 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R105 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 9.3005
R106 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 9.3005
R107 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 9.3005
R108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 9.3005
R109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 9.3005
R110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 9.3005
R111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 9.3005
R112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 9.3005
R113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 9.3005
R114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 9.3005
R115 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 9.3005
R116 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R117 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 9.3005
R118 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 9.3005
R119 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 9.3005
R120 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 9.3005
R121 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 9.3005
R122 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 9.3005
R123 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R124 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 9.3005
R125 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 9.3005
R126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 9.3005
R127 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R128 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 9.3005
R129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 9.3005
R130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R131 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 9.3005
R132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 9.3005
R133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 4.64654
R134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 4.64654
R135 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 4.64654
R136 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 4.64654
R137 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 4.64654
R138 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 4.64654
R139 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 4.64654
R140 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 4.64654
R141 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 4.64654
R142 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 2.36206
R143 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 2.36206
R144 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 2.36206
R145 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 2.36206
R146 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 2.19742
R147 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 2.19742
R148 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 2.19742
R149 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 1.56363
R150 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 1.56363
R151 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 1.5505
R152 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 1.5505
R153 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 1.5505
R154 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 1.5505
R155 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 1.5505
R156 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 1.5505
R157 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 1.5505
R158 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 1.5505
R159 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 1.5505
R160 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.5505
R161 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 1.5505
R162 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 1.5505
R163 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 1.5505
R164 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 1.5505
R165 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 1.5505
R166 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 1.5505
R167 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n143 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n142 1.5505
R168 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n145 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n144 1.5505
R169 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R170 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 1.25468
R171 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 1.25468
R172 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 1.25468
R173 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 1.25468
R174 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 1.25468
R175 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 1.25468
R176 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 1.19225
R177 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 1.19225
R178 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 1.19225
R179 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 1.19225
R180 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 1.19225
R181 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n142 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.14402
R182 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 1.07024
R183 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 1.07024
R184 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.07024
R185 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 1.07024
R186 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 1.07024
R187 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 1.07024
R188 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 1.0237
R189 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 1.0237
R190 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 1.0237
R191 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 1.0237
R192 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 1.0237
R193 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 1.0237
R194 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 0.885803
R195 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.885803
R196 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 0.885803
R197 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 0.885803
R198 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 0.885803
R199 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 0.885803
R200 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 0.885803
R201 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.885803
R202 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.812055
R203 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 0.812055
R204 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.77514
R205 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.77514
R206 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 0.77514
R207 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.77514
R208 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 0.77514
R209 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 0.77514
R210 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 0.77514
R211 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 0.77514
R212 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R213 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 0.756696
R214 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.756696
R215 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R216 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R217 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R218 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R219 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.756696
R220 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.711459
R221 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 0.711459
R222 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n145 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 0.701365
R223 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.647417
R224 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 0.647417
R225 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 0.590702
R226 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 0.590702
R227 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 0.590702
R228 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 0.590702
R229 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 0.590702
R230 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.590702
R231 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 0.576566
R232 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.576566
R233 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.530034
R234 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 0.530034
R235 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 0.290206
R236 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 0.290206
R237 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 0.290206
R238 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 0.290206
R239 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 0.290206
R240 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 0.290206
R241 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 0.290206
R242 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 0.290206
R243 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R244 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R245 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R246 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R247 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 0.203382
R248 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n145 0.203382
R249 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 0.154071
R250 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 0.154071
R251 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n143 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.154071
R252 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 0.154071
R253 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 0.137464
R254 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 0.137464
R255 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 0.134964
R256 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 0.134964
R257 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.0183571
R258 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.0183571
R259 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 0.0183571
R260 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 0.0183571
R261 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 0.0183571
R262 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 0.0183571
R263 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 0.0183571
R264 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0183571
R265 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0183571
R266 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n144 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R267 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n144 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n143 0.0183571
R268 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R269 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 0.0183571
R270 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 0.0183571
R271 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 0.0183571
R272 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 0.0183571
R273 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 0.0183571
R274 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R275 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 0.0106786
R276 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 0.0106786
R277 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0106786
R278 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 0.00992001
R279 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.00992001
R280 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 0.00992001
R281 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 0.00992001
R282 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 0.00992001
R283 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 0.00992001
R284 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 0.00992001
R285 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 0.00992001
R286 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 0.00992001
R287 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.00992001
R288 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R289 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.00992001
R290 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 0.00992001
R291 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.00992001
R292 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 0.00992001
R293 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.00992001
R294 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 0.00992001
R295 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R296 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 0.00817857
R297 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 0.00817857
R298 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 0.00817857
R299 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.00817857
R300 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 0.00817857
R301 GNDA.n2274 GNDA.n45 183150
R302 GNDA.n393 GNDA.n45 156825
R303 GNDA.n2274 GNDA.n46 137500
R304 GNDA.n315 GNDA.n245 13230.3
R305 GNDA.n2275 GNDA.n44 13230.3
R306 GNDA.n387 GNDA.n240 13200
R307 GNDA.n384 GNDA.n244 12026.7
R308 GNDA.n2275 GNDA.n43 12026.7
R309 GNDA.n398 GNDA.n397 11535.1
R310 GNDA.n388 GNDA.n243 11440
R311 GNDA.n383 GNDA.n382 11163
R312 GNDA.n382 GNDA.n246 11163
R313 GNDA.n242 GNDA.n241 10995.4
R314 GNDA.n386 GNDA.n385 10775.9
R315 GNDA.n392 GNDA.n237 10458.6
R316 GNDA.n393 GNDA.n392 10437.1
R317 GNDA.n396 GNDA.n393 10431.7
R318 GNDA.n239 GNDA.n237 10299.2
R319 GNDA.n385 GNDA.n243 10217
R320 GNDA.n243 GNDA.n242 10217
R321 GNDA.n389 GNDA.n241 9265.27
R322 GNDA.n241 GNDA.n46 8214.68
R323 GNDA.n386 GNDA.n238 8140
R324 GNDA.n388 GNDA.n387 7385.71
R325 GNDA.n395 GNDA.n394 6640.37
R326 GNDA.n401 GNDA.n400 6580
R327 GNDA.n387 GNDA.n386 6364.29
R328 GNDA.n397 GNDA.n396 6053.72
R329 GNDA.n398 GNDA.n239 6053.72
R330 GNDA.n390 GNDA.n389 5313.76
R331 GNDA.n355 GNDA.n245 4187.59
R332 GNDA.n380 GNDA.n44 4187.59
R333 GNDA.n397 GNDA.n391 4106.67
R334 GNDA.n392 GNDA.t182 4106.67
R335 GNDA.n399 GNDA.n398 4106.67
R336 GNDA.n403 GNDA.n237 3947.06
R337 GNDA.t19 GNDA.n2274 3899.06
R338 GNDA.n384 GNDA.n383 3223.76
R339 GNDA.n246 GNDA.n43 3223.76
R340 GNDA.n2274 GNDA.t58 3182.21
R341 GNDA.n389 GNDA.n388 2900.98
R342 GNDA.n394 GNDA.n46 2704.59
R343 GNDA.n383 GNDA.n245 2699.31
R344 GNDA.n246 GNDA.n44 2699.31
R345 GNDA.n400 GNDA.n238 2680
R346 GNDA.n244 GNDA.n238 2453.69
R347 GNDA.t92 GNDA.n315 2097.43
R348 GNDA.n402 GNDA.n238 1964.17
R349 GNDA.n390 GNDA.n240 1885.71
R350 GNDA.n382 GNDA.n381 1800
R351 GNDA.t45 GNDA.n403 1404.35
R352 GNDA.n402 GNDA.n401 1375
R353 GNDA.n401 GNDA.n239 1375
R354 GNDA.n396 GNDA.n395 1356.67
R355 GNDA.n395 GNDA.n45 1356.67
R356 GNDA.n1493 GNDA.n1291 1224.73
R357 GNDA.n1359 GNDA.n1324 1214.72
R358 GNDA.n1359 GNDA.n1358 1214.72
R359 GNDA.n1358 GNDA.n1357 1214.72
R360 GNDA.n1357 GNDA.n1332 1214.72
R361 GNDA.n1332 GNDA.n416 1214.72
R362 GNDA.n1349 GNDA.n415 1214.72
R363 GNDA.n1349 GNDA.n1348 1214.72
R364 GNDA.n1348 GNDA.n1347 1214.72
R365 GNDA.n1347 GNDA.n1343 1214.72
R366 GNDA.n1343 GNDA.n414 1214.72
R367 GNDA.n2198 GNDA.n96 1185.07
R368 GNDA.n2198 GNDA.n2197 1185.07
R369 GNDA.n380 GNDA.n379 1182.8
R370 GNDA.n356 GNDA.n355 1182.8
R371 GNDA.n400 GNDA.n399 1043.16
R372 GNDA.n394 GNDA.n391 1043.16
R373 GNDA.n2264 GNDA.t276 1029.15
R374 GNDA.n703 GNDA.n702 979.201
R375 GNDA.n403 GNDA.n402 936.601
R376 GNDA.t129 GNDA.n244 849.628
R377 GNDA.t182 GNDA.n416 823.313
R378 GNDA.n289 GNDA.t186 749.742
R379 GNDA.n336 GNDA.t198 749.742
R380 GNDA.n7 GNDA.t224 749.742
R381 GNDA.n2296 GNDA.t211 749.742
R382 GNDA.n315 GNDA.t129 685.448
R383 GNDA.n1316 GNDA.n1312 669.307
R384 GNDA.n391 GNDA.n390 668.693
R385 GNDA.n259 GNDA.t214 659.367
R386 GNDA.n284 GNDA.t175 659.367
R387 GNDA.n2157 GNDA.n2156 590.689
R388 GNDA.n2182 GNDA.n2181 590.689
R389 GNDA.n2163 GNDA.n180 590.689
R390 GNDA.n2211 GNDA.n47 590.689
R391 GNDA.n2227 GNDA.n2226 590.689
R392 GNDA.n545 GNDA.n544 590.689
R393 GNDA.n2206 GNDA.t276 586.76
R394 GNDA.n2153 GNDA.n192 585
R395 GNDA.n2151 GNDA.n2150 585
R396 GNDA.n194 GNDA.n193 585
R397 GNDA.n200 GNDA.n196 585
R398 GNDA.n2143 GNDA.n2142 585
R399 GNDA.n2140 GNDA.n198 585
R400 GNDA.n2139 GNDA.n201 585
R401 GNDA.n2137 GNDA.n2136 585
R402 GNDA.n203 GNDA.n202 585
R403 GNDA.n2131 GNDA.n2130 585
R404 GNDA.n2128 GNDA.n207 585
R405 GNDA.n2126 GNDA.n2125 585
R406 GNDA.n2125 GNDA.n2124 585
R407 GNDA.n207 GNDA.n206 585
R408 GNDA.n2132 GNDA.n2131 585
R409 GNDA.n2132 GNDA.n181 585
R410 GNDA.n2133 GNDA.n203 585
R411 GNDA.n2136 GNDA.n2135 585
R412 GNDA.n205 GNDA.n201 585
R413 GNDA.n198 GNDA.n197 585
R414 GNDA.n2144 GNDA.n2143 585
R415 GNDA.n2146 GNDA.n196 585
R416 GNDA.n2147 GNDA.n194 585
R417 GNDA.n2150 GNDA.n2149 585
R418 GNDA.n195 GNDA.n192 585
R419 GNDA.n195 GNDA.n181 585
R420 GNDA.n2009 GNDA.n463 585
R421 GNDA.n2010 GNDA.n461 585
R422 GNDA.n460 GNDA.n457 585
R423 GNDA.n2016 GNDA.n456 585
R424 GNDA.n2017 GNDA.n455 585
R425 GNDA.n2018 GNDA.n453 585
R426 GNDA.n452 GNDA.n449 585
R427 GNDA.n2024 GNDA.n448 585
R428 GNDA.n2025 GNDA.n447 585
R429 GNDA.n2026 GNDA.n445 585
R430 GNDA.n444 GNDA.n440 585
R431 GNDA.n2031 GNDA.n436 585
R432 GNDA.n2031 GNDA.n2030 585
R433 GNDA.n2028 GNDA.n440 585
R434 GNDA.n2027 GNDA.n2026 585
R435 GNDA.n2027 GNDA.n417 585
R436 GNDA.n2025 GNDA.n442 585
R437 GNDA.n2024 GNDA.n2023 585
R438 GNDA.n2021 GNDA.n449 585
R439 GNDA.n2019 GNDA.n2018 585
R440 GNDA.n2017 GNDA.n450 585
R441 GNDA.n2016 GNDA.n2015 585
R442 GNDA.n2013 GNDA.n457 585
R443 GNDA.n2011 GNDA.n2010 585
R444 GNDA.n2009 GNDA.n458 585
R445 GNDA.n458 GNDA.n417 585
R446 GNDA.n1718 GNDA.n1717 585
R447 GNDA.n1718 GNDA.n414 585
R448 GNDA.n869 GNDA.n868 585
R449 GNDA.n1343 GNDA.n868 585
R450 GNDA.n1345 GNDA.n1342 585
R451 GNDA.n1347 GNDA.n1342 585
R452 GNDA.n1344 GNDA.n1341 585
R453 GNDA.n1348 GNDA.n1341 585
R454 GNDA.n1340 GNDA.n1338 585
R455 GNDA.n1349 GNDA.n1340 585
R456 GNDA.n1339 GNDA.n1336 585
R457 GNDA.n1339 GNDA.n415 585
R458 GNDA.n1353 GNDA.n1335 585
R459 GNDA.n1335 GNDA.n416 585
R460 GNDA.n1354 GNDA.n1334 585
R461 GNDA.n1334 GNDA.n1332 585
R462 GNDA.n1355 GNDA.n1331 585
R463 GNDA.n1357 GNDA.n1331 585
R464 GNDA.n1330 GNDA.n1328 585
R465 GNDA.n1358 GNDA.n1330 585
R466 GNDA.n1361 GNDA.n1327 585
R467 GNDA.n1359 GNDA.n1327 585
R468 GNDA.n1363 GNDA.n1362 585
R469 GNDA.n1363 GNDA.n1324 585
R470 GNDA.n1362 GNDA.n1323 585
R471 GNDA.n1324 GNDA.n1323 585
R472 GNDA.n1361 GNDA.n1360 585
R473 GNDA.n1360 GNDA.n1359 585
R474 GNDA.n1329 GNDA.n1328 585
R475 GNDA.n1358 GNDA.n1329 585
R476 GNDA.n1356 GNDA.n1355 585
R477 GNDA.n1357 GNDA.n1356 585
R478 GNDA.n1354 GNDA.n1333 585
R479 GNDA.n1333 GNDA.n1332 585
R480 GNDA.n1353 GNDA.n1352 585
R481 GNDA.n1352 GNDA.n416 585
R482 GNDA.n1351 GNDA.n1336 585
R483 GNDA.n1351 GNDA.n415 585
R484 GNDA.n1350 GNDA.n1338 585
R485 GNDA.n1350 GNDA.n1349 585
R486 GNDA.n1344 GNDA.n1337 585
R487 GNDA.n1348 GNDA.n1337 585
R488 GNDA.n1346 GNDA.n1345 585
R489 GNDA.n1347 GNDA.n1346 585
R490 GNDA.n870 GNDA.n869 585
R491 GNDA.n1343 GNDA.n870 585
R492 GNDA.n1717 GNDA.n1716 585
R493 GNDA.n1716 GNDA.n414 585
R494 GNDA.n1393 GNDA.n1392 585
R495 GNDA.n1394 GNDA.n1393 585
R496 GNDA.n1391 GNDA.n1326 585
R497 GNDA.n1326 GNDA.n1325 585
R498 GNDA.n1390 GNDA.n1389 585
R499 GNDA.n1389 GNDA.n1388 585
R500 GNDA.n1365 GNDA.n1364 585
R501 GNDA.n1387 GNDA.n1365 585
R502 GNDA.n1385 GNDA.n1384 585
R503 GNDA.n1386 GNDA.n1385 585
R504 GNDA.n1383 GNDA.n1367 585
R505 GNDA.n1367 GNDA.n1366 585
R506 GNDA.n1382 GNDA.n1381 585
R507 GNDA.n1381 GNDA.n1380 585
R508 GNDA.n1369 GNDA.n1368 585
R509 GNDA.n1379 GNDA.n1369 585
R510 GNDA.n1377 GNDA.n1376 585
R511 GNDA.n1378 GNDA.n1377 585
R512 GNDA.n1375 GNDA.n1371 585
R513 GNDA.n1371 GNDA.n1370 585
R514 GNDA.n1374 GNDA.n1373 585
R515 GNDA.n1373 GNDA.n1372 585
R516 GNDA.n825 GNDA.n824 585
R517 GNDA.n824 GNDA.n413 585
R518 GNDA.n1317 GNDA.n1313 585
R519 GNDA.n1411 GNDA.n1410 585
R520 GNDA.t182 GNDA.n1411 585
R521 GNDA.n2034 GNDA.n2033 585
R522 GNDA.n437 GNDA.n435 585
R523 GNDA.n1847 GNDA.n1846 585
R524 GNDA.n1849 GNDA.n1848 585
R525 GNDA.n1851 GNDA.n1850 585
R526 GNDA.n1853 GNDA.n1852 585
R527 GNDA.n1855 GNDA.n1854 585
R528 GNDA.n1857 GNDA.n1856 585
R529 GNDA.n1859 GNDA.n1858 585
R530 GNDA.n1861 GNDA.n1860 585
R531 GNDA.n1863 GNDA.n1862 585
R532 GNDA.n1864 GNDA.n1845 585
R533 GNDA.n916 GNDA.n915 585
R534 GNDA.n914 GNDA.n913 585
R535 GNDA.n912 GNDA.n911 585
R536 GNDA.n910 GNDA.n909 585
R537 GNDA.n908 GNDA.n907 585
R538 GNDA.n906 GNDA.n905 585
R539 GNDA.n904 GNDA.n903 585
R540 GNDA.n902 GNDA.n901 585
R541 GNDA.n900 GNDA.n899 585
R542 GNDA.n898 GNDA.n897 585
R543 GNDA.n896 GNDA.n895 585
R544 GNDA.n441 GNDA.n438 585
R545 GNDA.n1112 GNDA.n1111 585
R546 GNDA.n1110 GNDA.n1109 585
R547 GNDA.n1108 GNDA.n1107 585
R548 GNDA.n1106 GNDA.n1105 585
R549 GNDA.n1104 GNDA.n1103 585
R550 GNDA.n1102 GNDA.n1101 585
R551 GNDA.n1100 GNDA.n1099 585
R552 GNDA.n1098 GNDA.n1097 585
R553 GNDA.n1096 GNDA.n1095 585
R554 GNDA.n1094 GNDA.n1093 585
R555 GNDA.n1092 GNDA.n1091 585
R556 GNDA.n919 GNDA.n894 585
R557 GNDA.n1719 GNDA.n439 585
R558 GNDA.n1719 GNDA.n867 585
R559 GNDA.n1814 GNDA.n826 585
R560 GNDA.n1801 GNDA.n827 585
R561 GNDA.n1810 GNDA.n1809 585
R562 GNDA.n846 GNDA.n844 585
R563 GNDA.n1726 GNDA.n1725 585
R564 GNDA.n1730 GNDA.n1729 585
R565 GNDA.n1732 GNDA.n1731 585
R566 GNDA.n1739 GNDA.n1738 585
R567 GNDA.n1737 GNDA.n1723 585
R568 GNDA.n1745 GNDA.n1744 585
R569 GNDA.n1747 GNDA.n1746 585
R570 GNDA.n1721 GNDA.n1720 585
R571 GNDA.n1715 GNDA.n439 585
R572 GNDA.n1715 GNDA.n867 585
R573 GNDA.n1714 GNDA.n1713 585
R574 GNDA.n1711 GNDA.n1710 585
R575 GNDA.n1709 GNDA.n1708 585
R576 GNDA.n1625 GNDA.n873 585
R577 GNDA.n1627 GNDA.n1626 585
R578 GNDA.n1631 GNDA.n1630 585
R579 GNDA.n1633 GNDA.n1632 585
R580 GNDA.n1640 GNDA.n1639 585
R581 GNDA.n1638 GNDA.n1623 585
R582 GNDA.n1646 GNDA.n1645 585
R583 GNDA.n1648 GNDA.n1647 585
R584 GNDA.n1621 GNDA.n1620 585
R585 GNDA.n508 GNDA.n208 585
R586 GNDA.n512 GNDA.n509 585
R587 GNDA.n514 GNDA.n513 585
R588 GNDA.n515 GNDA.n507 585
R589 GNDA.n517 GNDA.n516 585
R590 GNDA.n519 GNDA.n505 585
R591 GNDA.n521 GNDA.n520 585
R592 GNDA.n522 GNDA.n504 585
R593 GNDA.n524 GNDA.n523 585
R594 GNDA.n526 GNDA.n502 585
R595 GNDA.n528 GNDA.n527 585
R596 GNDA.n529 GNDA.n501 585
R597 GNDA.n2103 GNDA.n2102 585
R598 GNDA.n2104 GNDA.n217 585
R599 GNDA.n2106 GNDA.n2105 585
R600 GNDA.n2108 GNDA.n215 585
R601 GNDA.n2110 GNDA.n2109 585
R602 GNDA.n2111 GNDA.n214 585
R603 GNDA.n2113 GNDA.n2112 585
R604 GNDA.n2115 GNDA.n212 585
R605 GNDA.n2117 GNDA.n2116 585
R606 GNDA.n2118 GNDA.n211 585
R607 GNDA.n2120 GNDA.n2119 585
R608 GNDA.n2122 GNDA.n210 585
R609 GNDA.n2051 GNDA.n2050 585
R610 GNDA.n2052 GNDA.n228 585
R611 GNDA.n2054 GNDA.n2053 585
R612 GNDA.n2056 GNDA.n226 585
R613 GNDA.n2058 GNDA.n2057 585
R614 GNDA.n2059 GNDA.n225 585
R615 GNDA.n2061 GNDA.n2060 585
R616 GNDA.n2063 GNDA.n223 585
R617 GNDA.n2065 GNDA.n2064 585
R618 GNDA.n2066 GNDA.n222 585
R619 GNDA.n2068 GNDA.n2067 585
R620 GNDA.n2070 GNDA.n221 585
R621 GNDA.n2007 GNDA.n466 585
R622 GNDA.n467 GNDA.n466 585
R623 GNDA.n2001 GNDA.n2000 585
R624 GNDA.n1998 GNDA.n486 585
R625 GNDA.n1891 GNDA.n1890 585
R626 GNDA.n1993 GNDA.n1992 585
R627 GNDA.n1991 GNDA.n1990 585
R628 GNDA.n1917 GNDA.n1895 585
R629 GNDA.n1919 GNDA.n1918 585
R630 GNDA.n1924 GNDA.n1923 585
R631 GNDA.n1922 GNDA.n1915 585
R632 GNDA.n1930 GNDA.n1929 585
R633 GNDA.n1932 GNDA.n1931 585
R634 GNDA.n480 GNDA.n465 585
R635 GNDA.n2007 GNDA.n2006 585
R636 GNDA.n2006 GNDA.n467 585
R637 GNDA.n2005 GNDA.n464 585
R638 GNDA.n1021 GNDA.n468 585
R639 GNDA.n1044 GNDA.n1043 585
R640 GNDA.n1041 GNDA.n1040 585
R641 GNDA.n1039 GNDA.n1038 585
R642 GNDA.n1034 GNDA.n1033 585
R643 GNDA.n1032 GNDA.n1031 585
R644 GNDA.n1027 GNDA.n1026 585
R645 GNDA.n1025 GNDA.n947 585
R646 GNDA.n1052 GNDA.n1051 585
R647 GNDA.n1054 GNDA.n1053 585
R648 GNDA.n1057 GNDA.n1056 585
R649 GNDA.n1233 GNDA.n1232 585
R650 GNDA.n1230 GNDA.n1229 585
R651 GNDA.n1228 GNDA.n1227 585
R652 GNDA.n1144 GNDA.n1062 585
R653 GNDA.n1146 GNDA.n1145 585
R654 GNDA.n1150 GNDA.n1149 585
R655 GNDA.n1152 GNDA.n1151 585
R656 GNDA.n1159 GNDA.n1158 585
R657 GNDA.n1157 GNDA.n1142 585
R658 GNDA.n1165 GNDA.n1164 585
R659 GNDA.n1167 GNDA.n1166 585
R660 GNDA.n1140 GNDA.n1139 585
R661 GNDA.n820 GNDA.n819 585
R662 GNDA.n818 GNDA.n500 585
R663 GNDA.n817 GNDA.n816 585
R664 GNDA.n815 GNDA.n814 585
R665 GNDA.n813 GNDA.n812 585
R666 GNDA.n811 GNDA.n810 585
R667 GNDA.n809 GNDA.n808 585
R668 GNDA.n807 GNDA.n806 585
R669 GNDA.n805 GNDA.n804 585
R670 GNDA.n803 GNDA.n802 585
R671 GNDA.n801 GNDA.n800 585
R672 GNDA.n1839 GNDA.n494 585
R673 GNDA.n1866 GNDA.n1865 585
R674 GNDA.n1868 GNDA.n1844 585
R675 GNDA.n1871 GNDA.n1870 585
R676 GNDA.n1872 GNDA.n1843 585
R677 GNDA.n1874 GNDA.n1873 585
R678 GNDA.n1876 GNDA.n1842 585
R679 GNDA.n1879 GNDA.n1878 585
R680 GNDA.n1880 GNDA.n1841 585
R681 GNDA.n1882 GNDA.n1881 585
R682 GNDA.n1884 GNDA.n1840 585
R683 GNDA.n1885 GNDA.n488 585
R684 GNDA.n1839 GNDA.n487 585
R685 GNDA.n1837 GNDA.n1836 585
R686 GNDA.n1835 GNDA.n823 585
R687 GNDA.n1834 GNDA.n822 585
R688 GNDA.n1839 GNDA.n822 585
R689 GNDA.n1833 GNDA.n1832 585
R690 GNDA.n1831 GNDA.n1830 585
R691 GNDA.n1829 GNDA.n1828 585
R692 GNDA.n1827 GNDA.n1826 585
R693 GNDA.n1825 GNDA.n1824 585
R694 GNDA.n1823 GNDA.n1822 585
R695 GNDA.n1821 GNDA.n1820 585
R696 GNDA.n1819 GNDA.n1818 585
R697 GNDA.n1817 GNDA.n1816 585
R698 GNDA.n1816 GNDA.n1815 585
R699 GNDA.n2265 GNDA.n54 585
R700 GNDA.n2268 GNDA.n2267 585
R701 GNDA.n2267 GNDA.n2266 585
R702 GNDA.n53 GNDA.n52 585
R703 GNDA.n2263 GNDA.n53 585
R704 GNDA.n2261 GNDA.n2260 585
R705 GNDA.n2262 GNDA.n2261 585
R706 GNDA.n2259 GNDA.n56 585
R707 GNDA.n56 GNDA.n55 585
R708 GNDA.n2258 GNDA.n2257 585
R709 GNDA.n2257 GNDA.n2256 585
R710 GNDA.n58 GNDA.n57 585
R711 GNDA.n59 GNDA.n58 585
R712 GNDA.n2042 GNDA.n2041 585
R713 GNDA.n2041 GNDA.n2040 585
R714 GNDA.n2043 GNDA.n2038 585
R715 GNDA.n2038 GNDA.n2037 585
R716 GNDA.n2045 GNDA.n2044 585
R717 GNDA.n2046 GNDA.n2045 585
R718 GNDA.n2039 GNDA.n231 585
R719 GNDA.n2047 GNDA.n231 585
R720 GNDA.n2049 GNDA.n229 585
R721 GNDA.n2049 GNDA.n2048 585
R722 GNDA.n2264 GNDA.n49 585
R723 GNDA.n1136 GNDA.n1135 585
R724 GNDA.n1130 GNDA.n1082 585
R725 GNDA.n1134 GNDA.n1082 585
R726 GNDA.n1132 GNDA.n1131 585
R727 GNDA.n1133 GNDA.n1132 585
R728 GNDA.n1129 GNDA.n1084 585
R729 GNDA.n1084 GNDA.n1083 585
R730 GNDA.n1128 GNDA.n1127 585
R731 GNDA.n1127 GNDA.n1126 585
R732 GNDA.n1125 GNDA.n1085 585
R733 GNDA.n1125 GNDA.n408 585
R734 GNDA.n1124 GNDA.n1123 585
R735 GNDA.n1124 GNDA.n409 585
R736 GNDA.n1122 GNDA.n1086 585
R737 GNDA.n1118 GNDA.n1086 585
R738 GNDA.n1121 GNDA.n1120 585
R739 GNDA.n1120 GNDA.n1119 585
R740 GNDA.n1088 GNDA.n1087 585
R741 GNDA.n1117 GNDA.n1088 585
R742 GNDA.n1115 GNDA.n1114 585
R743 GNDA.n1116 GNDA.n1115 585
R744 GNDA.n1113 GNDA.n1090 585
R745 GNDA.n1090 GNDA.n1089 585
R746 GNDA.n1138 GNDA.n406 585
R747 GNDA.n1519 GNDA.n1518 585
R748 GNDA.n1521 GNDA.n1283 585
R749 GNDA.n1616 GNDA.n1615 585
R750 GNDA.n1613 GNDA.n1612 585
R751 GNDA.n1611 GNDA.n1610 585
R752 GNDA.n1527 GNDA.n1263 585
R753 GNDA.n1529 GNDA.n1528 585
R754 GNDA.n1533 GNDA.n1532 585
R755 GNDA.n1535 GNDA.n1534 585
R756 GNDA.n1542 GNDA.n1541 585
R757 GNDA.n1540 GNDA.n1525 585
R758 GNDA.n1548 GNDA.n1547 585
R759 GNDA.n1550 GNDA.n1549 585
R760 GNDA.n1523 GNDA.n1522 585
R761 GNDA.n1513 GNDA.n1284 585
R762 GNDA.n1517 GNDA.n1284 585
R763 GNDA.n1515 GNDA.n1514 585
R764 GNDA.n1516 GNDA.n1515 585
R765 GNDA.n1512 GNDA.n1286 585
R766 GNDA.n1286 GNDA.n1285 585
R767 GNDA.n1511 GNDA.n1510 585
R768 GNDA.n1510 GNDA.n1509 585
R769 GNDA.n1508 GNDA.n1287 585
R770 GNDA.n1508 GNDA.n411 585
R771 GNDA.n1507 GNDA.n1506 585
R772 GNDA.n1507 GNDA.n412 585
R773 GNDA.n1505 GNDA.n1288 585
R774 GNDA.n1501 GNDA.n1288 585
R775 GNDA.n1504 GNDA.n1503 585
R776 GNDA.n1503 GNDA.n1502 585
R777 GNDA.n1290 GNDA.n1289 585
R778 GNDA.n1500 GNDA.n1290 585
R779 GNDA.n1498 GNDA.n1497 585
R780 GNDA.n1499 GNDA.n1498 585
R781 GNDA.n1496 GNDA.n1292 585
R782 GNDA.n1292 GNDA.n1291 585
R783 GNDA.n1495 GNDA.n1494 585
R784 GNDA.n1494 GNDA.n1493 585
R785 GNDA.n1294 GNDA.n1293 585
R786 GNDA.n1492 GNDA.n1294 585
R787 GNDA.n1490 GNDA.n1489 585
R788 GNDA.n1491 GNDA.n1490 585
R789 GNDA.n1488 GNDA.n1296 585
R790 GNDA.n1296 GNDA.n1295 585
R791 GNDA.n1487 GNDA.n1486 585
R792 GNDA.n1486 GNDA.n1485 585
R793 GNDA.n1298 GNDA.n1297 585
R794 GNDA.n1484 GNDA.n1298 585
R795 GNDA.n1482 GNDA.n1481 585
R796 GNDA.n1483 GNDA.n1482 585
R797 GNDA.n1480 GNDA.n1300 585
R798 GNDA.n1300 GNDA.n1299 585
R799 GNDA.n1479 GNDA.n1478 585
R800 GNDA.n1478 GNDA.n1477 585
R801 GNDA.n1302 GNDA.n1301 585
R802 GNDA.n1476 GNDA.n1302 585
R803 GNDA.n1474 GNDA.n1473 585
R804 GNDA.n1475 GNDA.n1474 585
R805 GNDA.n1472 GNDA.n1304 585
R806 GNDA.n1304 GNDA.n1303 585
R807 GNDA.n1424 GNDA.n1305 585
R808 GNDA.n1424 GNDA.n1423 585
R809 GNDA.n1417 GNDA.n1306 585
R810 GNDA.n1421 GNDA.n1306 585
R811 GNDA.n1419 GNDA.n1418 585
R812 GNDA.n1420 GNDA.n1419 585
R813 GNDA.n1416 GNDA.n1308 585
R814 GNDA.n1308 GNDA.n1307 585
R815 GNDA.n1415 GNDA.n1414 585
R816 GNDA.n1414 GNDA.n1413 585
R817 GNDA.n1310 GNDA.n1309 585
R818 GNDA.n1412 GNDA.n1310 585
R819 GNDA.n1408 GNDA.n1407 585
R820 GNDA.n1407 GNDA.n1311 585
R821 GNDA.n1406 GNDA.n1318 585
R822 GNDA.n1406 GNDA.n1405 585
R823 GNDA.n1400 GNDA.n1319 585
R824 GNDA.n1404 GNDA.n1319 585
R825 GNDA.n1402 GNDA.n1401 585
R826 GNDA.n1403 GNDA.n1402 585
R827 GNDA.n1399 GNDA.n1321 585
R828 GNDA.n1321 GNDA.n1320 585
R829 GNDA.n1398 GNDA.n1397 585
R830 GNDA.n1397 GNDA.n1396 585
R831 GNDA.n1449 GNDA.n893 585
R832 GNDA.n1450 GNDA.n1448 585
R833 GNDA.n1451 GNDA.n1446 585
R834 GNDA.n1444 GNDA.n1441 585
R835 GNDA.n1457 GNDA.n1440 585
R836 GNDA.n1458 GNDA.n1438 585
R837 GNDA.n1459 GNDA.n1437 585
R838 GNDA.n1435 GNDA.n1433 585
R839 GNDA.n1464 GNDA.n1432 585
R840 GNDA.n1465 GNDA.n1430 585
R841 GNDA.n1429 GNDA.n1426 585
R842 GNDA.n1470 GNDA.n1425 585
R843 GNDA.n1619 GNDA.n1618 585
R844 GNDA.n1619 GNDA.n867 585
R845 GNDA.n1470 GNDA.n1469 585
R846 GNDA.n1467 GNDA.n1426 585
R847 GNDA.n1466 GNDA.n1465 585
R848 GNDA.n1464 GNDA.n1463 585
R849 GNDA.n1462 GNDA.n1433 585
R850 GNDA.n1460 GNDA.n1459 585
R851 GNDA.n1458 GNDA.n1434 585
R852 GNDA.n1457 GNDA.n1456 585
R853 GNDA.n1454 GNDA.n1441 585
R854 GNDA.n1452 GNDA.n1451 585
R855 GNDA.n1450 GNDA.n1443 585
R856 GNDA.n1449 GNDA.n1260 585
R857 GNDA.n1618 GNDA.n1617 585
R858 GNDA.n1617 GNDA.n867 585
R859 GNDA.n1236 GNDA.n943 585
R860 GNDA.n1237 GNDA.n934 585
R861 GNDA.n1240 GNDA.n933 585
R862 GNDA.n1241 GNDA.n932 585
R863 GNDA.n1244 GNDA.n931 585
R864 GNDA.n1245 GNDA.n930 585
R865 GNDA.n1248 GNDA.n929 585
R866 GNDA.n1250 GNDA.n928 585
R867 GNDA.n1251 GNDA.n927 585
R868 GNDA.n1252 GNDA.n926 585
R869 GNDA.n935 GNDA.n918 585
R870 GNDA.n1258 GNDA.n917 585
R871 GNDA.n1059 GNDA.n1058 585
R872 GNDA.n1058 GNDA.n467 585
R873 GNDA.n1258 GNDA.n1257 585
R874 GNDA.n920 GNDA.n918 585
R875 GNDA.n1253 GNDA.n1252 585
R876 GNDA.n1251 GNDA.n925 585
R877 GNDA.n1250 GNDA.n1249 585
R878 GNDA.n1248 GNDA.n1247 585
R879 GNDA.n1246 GNDA.n1245 585
R880 GNDA.n1244 GNDA.n1243 585
R881 GNDA.n1242 GNDA.n1241 585
R882 GNDA.n1240 GNDA.n1239 585
R883 GNDA.n1238 GNDA.n1237 585
R884 GNDA.n1236 GNDA.n1235 585
R885 GNDA.n1234 GNDA.n1059 585
R886 GNDA.n1234 GNDA.n467 585
R887 GNDA.n2184 GNDA.n170 585
R888 GNDA.n2187 GNDA.n2186 585
R889 GNDA.n173 GNDA.n172 585
R890 GNDA.n2082 GNDA.n2081 585
R891 GNDA.n2087 GNDA.n2080 585
R892 GNDA.n2088 GNDA.n2079 585
R893 GNDA.n2089 GNDA.n2078 585
R894 GNDA.n2076 GNDA.n2075 585
R895 GNDA.n2094 GNDA.n2074 585
R896 GNDA.n2095 GNDA.n2073 585
R897 GNDA.n2072 GNDA.n220 585
R898 GNDA.n2101 GNDA.n2100 585
R899 GNDA.n2100 GNDA.n2099 585
R900 GNDA.n2097 GNDA.n220 585
R901 GNDA.n2096 GNDA.n2095 585
R902 GNDA.n2094 GNDA.n2093 585
R903 GNDA.n2092 GNDA.n2076 585
R904 GNDA.n2090 GNDA.n2089 585
R905 GNDA.n2088 GNDA.n2077 585
R906 GNDA.n2087 GNDA.n2086 585
R907 GNDA.n2084 GNDA.n2082 585
R908 GNDA.n172 GNDA.n171 585
R909 GNDA.n2188 GNDA.n2187 585
R910 GNDA.n2190 GNDA.n170 585
R911 GNDA.n2154 GNDA.n191 585
R912 GNDA.n2155 GNDA.n2154 585
R913 GNDA.n798 GNDA.n797 585
R914 GNDA.n797 GNDA.n236 585
R915 GNDA.n796 GNDA.n533 585
R916 GNDA.n796 GNDA.n795 585
R917 GNDA.n784 GNDA.n532 585
R918 GNDA.n794 GNDA.n532 585
R919 GNDA.n792 GNDA.n791 585
R920 GNDA.n793 GNDA.n792 585
R921 GNDA.n549 GNDA.n547 585
R922 GNDA.n547 GNDA.n546 585
R923 GNDA.n711 GNDA.n710 585
R924 GNDA.n710 GNDA.n405 585
R925 GNDA.n712 GNDA.n708 585
R926 GNDA.n708 GNDA.n707 585
R927 GNDA.n721 GNDA.n720 585
R928 GNDA.n722 GNDA.n721 585
R929 GNDA.n696 GNDA.n695 585
R930 GNDA.n723 GNDA.n696 585
R931 GNDA.n726 GNDA.n725 585
R932 GNDA.n725 GNDA.n724 585
R933 GNDA.n700 GNDA.n697 585
R934 GNDA.n700 GNDA.n699 585
R935 GNDA.n690 GNDA.n190 585
R936 GNDA.n698 GNDA.n190 585
R937 GNDA.n2192 GNDA.n99 585
R938 GNDA.n183 GNDA.n99 585
R939 GNDA.n566 GNDA.n191 585
R940 GNDA.n685 GNDA.n566 585
R941 GNDA.n688 GNDA.n687 585
R942 GNDA.n687 GNDA.n686 585
R943 GNDA.n684 GNDA.n568 585
R944 GNDA.n684 GNDA.n683 585
R945 GNDA.n672 GNDA.n567 585
R946 GNDA.n682 GNDA.n567 585
R947 GNDA.n680 GNDA.n679 585
R948 GNDA.n681 GNDA.n680 585
R949 GNDA.n571 GNDA.n569 585
R950 GNDA.n596 GNDA.n569 585
R951 GNDA.n599 GNDA.n598 585
R952 GNDA.n598 GNDA.n597 585
R953 GNDA.n600 GNDA.n594 585
R954 GNDA.n594 GNDA.n593 585
R955 GNDA.n609 GNDA.n608 585
R956 GNDA.n610 GNDA.n609 585
R957 GNDA.n592 GNDA.n591 585
R958 GNDA.n611 GNDA.n592 585
R959 GNDA.n614 GNDA.n613 585
R960 GNDA.n613 GNDA.n612 585
R961 GNDA.n588 GNDA.n98 585
R962 GNDA.n98 GNDA.n97 585
R963 GNDA.n2195 GNDA.n2194 585
R964 GNDA.n2196 GNDA.n2195 585
R965 GNDA.n2192 GNDA.n2191 585
R966 GNDA.n2191 GNDA.n88 585
R967 GNDA.n169 GNDA.n87 585
R968 GNDA.n2228 GNDA.n87 585
R969 GNDA.n2230 GNDA.n85 585
R970 GNDA.n2230 GNDA.n2229 585
R971 GNDA.n2246 GNDA.n2245 585
R972 GNDA.n2245 GNDA.n2244 585
R973 GNDA.n2233 GNDA.n2231 585
R974 GNDA.n2243 GNDA.n2231 585
R975 GNDA.n2241 GNDA.n2240 585
R976 GNDA.n2242 GNDA.n2241 585
R977 GNDA.n2236 GNDA.n62 585
R978 GNDA.n2232 GNDA.n62 585
R979 GNDA.n2254 GNDA.n2253 585
R980 GNDA.n2255 GNDA.n2254 585
R981 GNDA.n64 GNDA.n63 585
R982 GNDA.n106 GNDA.n63 585
R983 GNDA.n105 GNDA.n104 585
R984 GNDA.n107 GNDA.n105 585
R985 GNDA.n111 GNDA.n110 585
R986 GNDA.n110 GNDA.n109 585
R987 GNDA.n112 GNDA.n48 585
R988 GNDA.n108 GNDA.n48 585
R989 GNDA.n2271 GNDA.n2270 585
R990 GNDA.n2272 GNDA.n2271 585
R991 GNDA.n333 GNDA.n252 543.014
R992 GNDA.n2293 GNDA.n17 543.014
R993 GNDA.n42 GNDA.t242 524.808
R994 GNDA.n2289 GNDA.t253 524.808
R995 GNDA.n314 GNDA.t204 524.808
R996 GNDA.n329 GNDA.t195 524.808
R997 GNDA.t182 GNDA.n414 512.884
R998 GNDA.n251 GNDA.t261 508.743
R999 GNDA.n2308 GNDA.t178 508.743
R1000 GNDA.n254 GNDA.t231 508.743
R1001 GNDA.n14 GNDA.t266 508.743
R1002 GNDA.n2302 GNDA.t245 508.743
R1003 GNDA.n352 GNDA.t248 499.442
R1004 GNDA.n340 GNDA.t256 499.442
R1005 GNDA.n2300 GNDA.t258 499.442
R1006 GNDA.n343 GNDA.t189 475.976
R1007 GNDA.n343 GNDA.t172 475.976
R1008 GNDA.n10 GNDA.t251 475.976
R1009 GNDA.n10 GNDA.t237 475.976
R1010 GNDA.n542 GNDA.t218 418.368
R1011 GNDA.n2159 GNDA.t208 418.368
R1012 GNDA.n2179 GNDA.t191 418.368
R1013 GNDA.n2162 GNDA.t239 418.368
R1014 GNDA.n2210 GNDA.t263 418.368
R1015 GNDA.n2224 GNDA.t183 418.368
R1016 GNDA.n355 GNDA.t235 409.656
R1017 GNDA.t229 GNDA.n380 409.656
R1018 GNDA.t182 GNDA.n415 391.411
R1019 GNDA.n1422 GNDA.n234 370.214
R1020 GNDA.n1422 GNDA.n233 365.957
R1021 GNDA.n358 GNDA.t234 338.034
R1022 GNDA.n377 GNDA.t228 338.034
R1023 GNDA.t235 GNDA.t50 333.793
R1024 GNDA.t50 GNDA.t105 333.793
R1025 GNDA.t105 GNDA.t103 333.793
R1026 GNDA.t103 GNDA.t15 333.793
R1027 GNDA.t15 GNDA.t127 333.793
R1028 GNDA.t107 GNDA.t138 333.793
R1029 GNDA.t138 GNDA.t168 333.793
R1030 GNDA.t168 GNDA.t278 333.793
R1031 GNDA.t278 GNDA.t101 333.793
R1032 GNDA.t101 GNDA.t229 333.793
R1033 GNDA.t182 GNDA.n233 327.661
R1034 GNDA.t182 GNDA.n179 172.876
R1035 GNDA.n2183 GNDA.t182 172.876
R1036 GNDA.t182 GNDA.n234 323.404
R1037 GNDA.n181 GNDA.t182 172.615
R1038 GNDA.t182 GNDA.n60 172.615
R1039 GNDA.n349 GNDA.n348 296.158
R1040 GNDA.n2307 GNDA.n2306 296.158
R1041 GNDA.n256 GNDA.n255 296.158
R1042 GNDA.n17 GNDA.n16 296.158
R1043 GNDA.n2305 GNDA.n2304 296.158
R1044 GNDA.t182 GNDA.t21 295.808
R1045 GNDA.n339 GNDA.n252 292.5
R1046 GNDA.n348 GNDA.n347 292.5
R1047 GNDA.n2305 GNDA.n3 292.5
R1048 GNDA.n351 GNDA.n252 292.5
R1049 GNDA.n17 GNDA.n4 292.5
R1050 GNDA.n1839 GNDA.n493 264.301
R1051 GNDA.n799 GNDA.n530 264.301
R1052 GNDA.n1888 GNDA.n1887 264.301
R1053 GNDA.n2269 GNDA.n51 264.301
R1054 GNDA.n1137 GNDA.n1081 264.301
R1055 GNDA.n1520 GNDA.n1282 264.301
R1056 GNDA.n2050 GNDA.n2049 259.416
R1057 GNDA.n1111 GNDA.n1090 259.416
R1058 GNDA.n1425 GNDA.n1424 259.416
R1059 GNDA.n1393 GNDA.n1363 259.416
R1060 GNDA.n917 GNDA.n916 259.416
R1061 GNDA.n2034 GNDA.n436 259.416
R1062 GNDA.n2102 GNDA.n2101 259.416
R1063 GNDA.n2126 GNDA.n208 259.416
R1064 GNDA.n1494 GNDA.n1292 259.416
R1065 GNDA.n151 GNDA.n150 258.334
R1066 GNDA.n1206 GNDA.n1205 258.334
R1067 GNDA.n1786 GNDA.n1785 258.334
R1068 GNDA.n1687 GNDA.n1686 258.334
R1069 GNDA.n1003 GNDA.n1002 258.334
R1070 GNDA.n1969 GNDA.n1912 258.334
R1071 GNDA.n654 GNDA.n577 258.334
R1072 GNDA.n766 GNDA.n555 258.334
R1073 GNDA.n1589 GNDA.n1588 258.334
R1074 GNDA.n2152 GNDA.n179 254.34
R1075 GNDA.n199 GNDA.n179 254.34
R1076 GNDA.n2141 GNDA.n179 254.34
R1077 GNDA.n2138 GNDA.n179 254.34
R1078 GNDA.n2129 GNDA.n179 254.34
R1079 GNDA.n2127 GNDA.n179 254.34
R1080 GNDA.n2123 GNDA.n181 254.34
R1081 GNDA.n2134 GNDA.n181 254.34
R1082 GNDA.n204 GNDA.n181 254.34
R1083 GNDA.n2145 GNDA.n181 254.34
R1084 GNDA.n2148 GNDA.n181 254.34
R1085 GNDA.n462 GNDA.n235 254.34
R1086 GNDA.n459 GNDA.n235 254.34
R1087 GNDA.n454 GNDA.n235 254.34
R1088 GNDA.n451 GNDA.n235 254.34
R1089 GNDA.n446 GNDA.n235 254.34
R1090 GNDA.n443 GNDA.n235 254.34
R1091 GNDA.n2029 GNDA.n417 254.34
R1092 GNDA.n2022 GNDA.n417 254.34
R1093 GNDA.n2020 GNDA.n417 254.34
R1094 GNDA.n2014 GNDA.n417 254.34
R1095 GNDA.n2012 GNDA.n417 254.34
R1096 GNDA.n2036 GNDA.n2035 254.34
R1097 GNDA.n2036 GNDA.n434 254.34
R1098 GNDA.n2036 GNDA.n433 254.34
R1099 GNDA.n2036 GNDA.n432 254.34
R1100 GNDA.n2036 GNDA.n431 254.34
R1101 GNDA.n2036 GNDA.n430 254.34
R1102 GNDA.n2036 GNDA.n429 254.34
R1103 GNDA.n2036 GNDA.n428 254.34
R1104 GNDA.n2036 GNDA.n427 254.34
R1105 GNDA.n2036 GNDA.n426 254.34
R1106 GNDA.n2036 GNDA.n425 254.34
R1107 GNDA.n2036 GNDA.n424 254.34
R1108 GNDA.n2036 GNDA.n423 254.34
R1109 GNDA.n2036 GNDA.n422 254.34
R1110 GNDA.n2036 GNDA.n421 254.34
R1111 GNDA.n2036 GNDA.n420 254.34
R1112 GNDA.n2036 GNDA.n419 254.34
R1113 GNDA.n2036 GNDA.n418 254.34
R1114 GNDA.n1813 GNDA.n1812 254.34
R1115 GNDA.n1812 GNDA.n1811 254.34
R1116 GNDA.n1812 GNDA.n843 254.34
R1117 GNDA.n1812 GNDA.n842 254.34
R1118 GNDA.n1812 GNDA.n841 254.34
R1119 GNDA.n1812 GNDA.n840 254.34
R1120 GNDA.n1812 GNDA.n839 254.34
R1121 GNDA.n1812 GNDA.n838 254.34
R1122 GNDA.n1812 GNDA.n837 254.34
R1123 GNDA.n1812 GNDA.n836 254.34
R1124 GNDA.n1812 GNDA.n835 254.34
R1125 GNDA.n1812 GNDA.n834 254.34
R1126 GNDA.n511 GNDA.n182 254.34
R1127 GNDA.n510 GNDA.n182 254.34
R1128 GNDA.n518 GNDA.n182 254.34
R1129 GNDA.n506 GNDA.n182 254.34
R1130 GNDA.n525 GNDA.n182 254.34
R1131 GNDA.n503 GNDA.n182 254.34
R1132 GNDA.n219 GNDA.n182 254.34
R1133 GNDA.n2107 GNDA.n182 254.34
R1134 GNDA.n216 GNDA.n182 254.34
R1135 GNDA.n2114 GNDA.n182 254.34
R1136 GNDA.n213 GNDA.n182 254.34
R1137 GNDA.n2121 GNDA.n182 254.34
R1138 GNDA.n230 GNDA.n182 254.34
R1139 GNDA.n2055 GNDA.n182 254.34
R1140 GNDA.n227 GNDA.n182 254.34
R1141 GNDA.n2062 GNDA.n182 254.34
R1142 GNDA.n224 GNDA.n182 254.34
R1143 GNDA.n2069 GNDA.n182 254.34
R1144 GNDA.n2003 GNDA.n2002 254.34
R1145 GNDA.n2003 GNDA.n485 254.34
R1146 GNDA.n2003 GNDA.n484 254.34
R1147 GNDA.n2003 GNDA.n483 254.34
R1148 GNDA.n2003 GNDA.n482 254.34
R1149 GNDA.n2003 GNDA.n481 254.34
R1150 GNDA.n2004 GNDA.n2003 254.34
R1151 GNDA.n2003 GNDA.n479 254.34
R1152 GNDA.n2003 GNDA.n478 254.34
R1153 GNDA.n2003 GNDA.n477 254.34
R1154 GNDA.n2003 GNDA.n476 254.34
R1155 GNDA.n2003 GNDA.n475 254.34
R1156 GNDA.n2003 GNDA.n474 254.34
R1157 GNDA.n2003 GNDA.n473 254.34
R1158 GNDA.n2003 GNDA.n472 254.34
R1159 GNDA.n2003 GNDA.n471 254.34
R1160 GNDA.n2003 GNDA.n470 254.34
R1161 GNDA.n2003 GNDA.n469 254.34
R1162 GNDA.n1839 GNDA.n821 254.34
R1163 GNDA.n1839 GNDA.n499 254.34
R1164 GNDA.n1839 GNDA.n498 254.34
R1165 GNDA.n1839 GNDA.n497 254.34
R1166 GNDA.n1839 GNDA.n496 254.34
R1167 GNDA.n1839 GNDA.n495 254.34
R1168 GNDA.n1867 GNDA.n1839 254.34
R1169 GNDA.n1869 GNDA.n1839 254.34
R1170 GNDA.n1875 GNDA.n1839 254.34
R1171 GNDA.n1877 GNDA.n1839 254.34
R1172 GNDA.n1883 GNDA.n1839 254.34
R1173 GNDA.n1886 GNDA.n1839 254.34
R1174 GNDA.n1839 GNDA.n1838 254.34
R1175 GNDA.n1839 GNDA.n489 254.34
R1176 GNDA.n1839 GNDA.n490 254.34
R1177 GNDA.n1839 GNDA.n491 254.34
R1178 GNDA.n1839 GNDA.n492 254.34
R1179 GNDA.n1812 GNDA.n833 254.34
R1180 GNDA.n1812 GNDA.n832 254.34
R1181 GNDA.n1812 GNDA.n831 254.34
R1182 GNDA.n1812 GNDA.n830 254.34
R1183 GNDA.n1812 GNDA.n829 254.34
R1184 GNDA.n1812 GNDA.n828 254.34
R1185 GNDA.n1447 GNDA.n233 254.34
R1186 GNDA.n1445 GNDA.n233 254.34
R1187 GNDA.n1439 GNDA.n233 254.34
R1188 GNDA.n1436 GNDA.n233 254.34
R1189 GNDA.n1431 GNDA.n233 254.34
R1190 GNDA.n1428 GNDA.n233 254.34
R1191 GNDA.n1468 GNDA.n234 254.34
R1192 GNDA.n1427 GNDA.n234 254.34
R1193 GNDA.n1461 GNDA.n234 254.34
R1194 GNDA.n1455 GNDA.n234 254.34
R1195 GNDA.n1453 GNDA.n234 254.34
R1196 GNDA.n1442 GNDA.n234 254.34
R1197 GNDA.n942 GNDA.n941 254.34
R1198 GNDA.n941 GNDA.n940 254.34
R1199 GNDA.n941 GNDA.n939 254.34
R1200 GNDA.n941 GNDA.n938 254.34
R1201 GNDA.n941 GNDA.n937 254.34
R1202 GNDA.n941 GNDA.n936 254.34
R1203 GNDA.n1256 GNDA.n1255 254.34
R1204 GNDA.n1255 GNDA.n1254 254.34
R1205 GNDA.n1255 GNDA.n924 254.34
R1206 GNDA.n1255 GNDA.n923 254.34
R1207 GNDA.n1255 GNDA.n922 254.34
R1208 GNDA.n1255 GNDA.n921 254.34
R1209 GNDA.n2185 GNDA.n2183 254.34
R1210 GNDA.n2183 GNDA.n178 254.34
R1211 GNDA.n2183 GNDA.n177 254.34
R1212 GNDA.n2183 GNDA.n176 254.34
R1213 GNDA.n2183 GNDA.n175 254.34
R1214 GNDA.n2183 GNDA.n174 254.34
R1215 GNDA.n2098 GNDA.n60 254.34
R1216 GNDA.n2071 GNDA.n60 254.34
R1217 GNDA.n2091 GNDA.n60 254.34
R1218 GNDA.n2085 GNDA.n60 254.34
R1219 GNDA.n2083 GNDA.n60 254.34
R1220 GNDA.n2189 GNDA.n60 254.34
R1221 GNDA.t182 GNDA.n1312 250.349
R1222 GNDA.n2099 GNDA.n2070 249.663
R1223 GNDA.n1257 GNDA.n919 249.663
R1224 GNDA.n1397 GNDA.n1323 249.663
R1225 GNDA.n1837 GNDA.n824 249.663
R1226 GNDA.n2030 GNDA.n441 249.663
R1227 GNDA.n1866 GNDA.n1845 249.663
R1228 GNDA.n2124 GNDA.n2122 249.663
R1229 GNDA.n820 GNDA.n501 249.663
R1230 GNDA.n1469 GNDA.n1304 249.663
R1231 GNDA.n356 GNDA.t236 233
R1232 GNDA.n379 GNDA.t230 233
R1233 GNDA.n258 GNDA.n257 197.133
R1234 GNDA.n286 GNDA.n285 197.133
R1235 GNDA.n2271 GNDA.n49 197
R1236 GNDA.n1139 GNDA.n1138 197
R1237 GNDA.n1411 GNDA.n1313 197
R1238 GNDA.n1620 GNDA.n1619 197
R1239 GNDA.n1720 GNDA.n1719 197
R1240 GNDA.n1058 GNDA.n1057 197
R1241 GNDA.n480 GNDA.n466 197
R1242 GNDA.n2195 GNDA.n99 197
R1243 GNDA.n2154 GNDA.n190 197
R1244 GNDA.n1522 GNDA.n1521 197
R1245 GNDA.n317 GNDA.t270 195.644
R1246 GNDA.n2201 GNDA.n61 195
R1247 GNDA.n706 GNDA.n705 195
R1248 GNDA.n375 GNDA.n374 194.3
R1249 GNDA.n372 GNDA.n371 194.3
R1250 GNDA.n368 GNDA.n367 194.3
R1251 GNDA.n365 GNDA.n364 194.3
R1252 GNDA.n361 GNDA.n360 194.3
R1253 GNDA.n2191 GNDA.n87 187.249
R1254 GNDA.n1234 GNDA.n1233 187.249
R1255 GNDA.n1715 GNDA.n1714 187.249
R1256 GNDA.n1815 GNDA.n1814 187.249
R1257 GNDA.n2006 GNDA.n2005 187.249
R1258 GNDA.n2001 GNDA.n487 187.249
R1259 GNDA.n687 GNDA.n566 187.249
R1260 GNDA.n797 GNDA.n494 187.249
R1261 GNDA.n1617 GNDA.n1616 187.249
R1262 GNDA.n152 GNDA.n151 185
R1263 GNDA.n154 GNDA.n153 185
R1264 GNDA.n156 GNDA.n155 185
R1265 GNDA.n158 GNDA.n157 185
R1266 GNDA.n160 GNDA.n159 185
R1267 GNDA.n162 GNDA.n161 185
R1268 GNDA.n164 GNDA.n163 185
R1269 GNDA.n166 GNDA.n165 185
R1270 GNDA.n167 GNDA.n83 185
R1271 GNDA.n134 GNDA.n133 185
R1272 GNDA.n136 GNDA.n135 185
R1273 GNDA.n138 GNDA.n137 185
R1274 GNDA.n140 GNDA.n139 185
R1275 GNDA.n142 GNDA.n141 185
R1276 GNDA.n144 GNDA.n143 185
R1277 GNDA.n146 GNDA.n145 185
R1278 GNDA.n148 GNDA.n147 185
R1279 GNDA.n150 GNDA.n149 185
R1280 GNDA.n116 GNDA.n115 185
R1281 GNDA.n118 GNDA.n117 185
R1282 GNDA.n120 GNDA.n119 185
R1283 GNDA.n122 GNDA.n121 185
R1284 GNDA.n124 GNDA.n123 185
R1285 GNDA.n126 GNDA.n125 185
R1286 GNDA.n128 GNDA.n127 185
R1287 GNDA.n130 GNDA.n129 185
R1288 GNDA.n132 GNDA.n131 185
R1289 GNDA.n114 GNDA.n113 185
R1290 GNDA.n102 GNDA.n101 185
R1291 GNDA.n103 GNDA.n66 185
R1292 GNDA.n2252 GNDA.n2251 185
R1293 GNDA.n2235 GNDA.n65 185
R1294 GNDA.n2239 GNDA.n2238 185
R1295 GNDA.n2237 GNDA.n2234 185
R1296 GNDA.n86 GNDA.n84 185
R1297 GNDA.n2248 GNDA.n2247 185
R1298 GNDA.n1207 GNDA.n1206 185
R1299 GNDA.n1209 GNDA.n1208 185
R1300 GNDA.n1211 GNDA.n1210 185
R1301 GNDA.n1213 GNDA.n1212 185
R1302 GNDA.n1215 GNDA.n1214 185
R1303 GNDA.n1217 GNDA.n1216 185
R1304 GNDA.n1219 GNDA.n1218 185
R1305 GNDA.n1221 GNDA.n1220 185
R1306 GNDA.n1222 GNDA.n1060 185
R1307 GNDA.n1189 GNDA.n1188 185
R1308 GNDA.n1191 GNDA.n1190 185
R1309 GNDA.n1193 GNDA.n1192 185
R1310 GNDA.n1195 GNDA.n1194 185
R1311 GNDA.n1197 GNDA.n1196 185
R1312 GNDA.n1199 GNDA.n1198 185
R1313 GNDA.n1201 GNDA.n1200 185
R1314 GNDA.n1203 GNDA.n1202 185
R1315 GNDA.n1205 GNDA.n1204 185
R1316 GNDA.n1171 GNDA.n1170 185
R1317 GNDA.n1173 GNDA.n1172 185
R1318 GNDA.n1175 GNDA.n1174 185
R1319 GNDA.n1177 GNDA.n1176 185
R1320 GNDA.n1179 GNDA.n1178 185
R1321 GNDA.n1181 GNDA.n1180 185
R1322 GNDA.n1183 GNDA.n1182 185
R1323 GNDA.n1185 GNDA.n1184 185
R1324 GNDA.n1187 GNDA.n1186 185
R1325 GNDA.n1169 GNDA.n1168 185
R1326 GNDA.n1163 GNDA.n1162 185
R1327 GNDA.n1161 GNDA.n1160 185
R1328 GNDA.n1156 GNDA.n1155 185
R1329 GNDA.n1154 GNDA.n1153 185
R1330 GNDA.n1148 GNDA.n1147 185
R1331 GNDA.n1143 GNDA.n1064 185
R1332 GNDA.n1226 GNDA.n1225 185
R1333 GNDA.n1063 GNDA.n1061 185
R1334 GNDA.n1787 GNDA.n1786 185
R1335 GNDA.n1789 GNDA.n1788 185
R1336 GNDA.n1791 GNDA.n1790 185
R1337 GNDA.n1793 GNDA.n1792 185
R1338 GNDA.n1795 GNDA.n1794 185
R1339 GNDA.n1797 GNDA.n1796 185
R1340 GNDA.n1799 GNDA.n1798 185
R1341 GNDA.n1800 GNDA.n865 185
R1342 GNDA.n1804 GNDA.n1803 185
R1343 GNDA.n1769 GNDA.n1768 185
R1344 GNDA.n1771 GNDA.n1770 185
R1345 GNDA.n1773 GNDA.n1772 185
R1346 GNDA.n1775 GNDA.n1774 185
R1347 GNDA.n1777 GNDA.n1776 185
R1348 GNDA.n1779 GNDA.n1778 185
R1349 GNDA.n1781 GNDA.n1780 185
R1350 GNDA.n1783 GNDA.n1782 185
R1351 GNDA.n1785 GNDA.n1784 185
R1352 GNDA.n1751 GNDA.n1750 185
R1353 GNDA.n1753 GNDA.n1752 185
R1354 GNDA.n1755 GNDA.n1754 185
R1355 GNDA.n1757 GNDA.n1756 185
R1356 GNDA.n1759 GNDA.n1758 185
R1357 GNDA.n1761 GNDA.n1760 185
R1358 GNDA.n1763 GNDA.n1762 185
R1359 GNDA.n1765 GNDA.n1764 185
R1360 GNDA.n1767 GNDA.n1766 185
R1361 GNDA.n1688 GNDA.n1687 185
R1362 GNDA.n1690 GNDA.n1689 185
R1363 GNDA.n1692 GNDA.n1691 185
R1364 GNDA.n1694 GNDA.n1693 185
R1365 GNDA.n1696 GNDA.n1695 185
R1366 GNDA.n1698 GNDA.n1697 185
R1367 GNDA.n1700 GNDA.n1699 185
R1368 GNDA.n1702 GNDA.n1701 185
R1369 GNDA.n1703 GNDA.n871 185
R1370 GNDA.n1670 GNDA.n1669 185
R1371 GNDA.n1672 GNDA.n1671 185
R1372 GNDA.n1674 GNDA.n1673 185
R1373 GNDA.n1676 GNDA.n1675 185
R1374 GNDA.n1678 GNDA.n1677 185
R1375 GNDA.n1680 GNDA.n1679 185
R1376 GNDA.n1682 GNDA.n1681 185
R1377 GNDA.n1684 GNDA.n1683 185
R1378 GNDA.n1686 GNDA.n1685 185
R1379 GNDA.n1652 GNDA.n1651 185
R1380 GNDA.n1654 GNDA.n1653 185
R1381 GNDA.n1656 GNDA.n1655 185
R1382 GNDA.n1658 GNDA.n1657 185
R1383 GNDA.n1660 GNDA.n1659 185
R1384 GNDA.n1662 GNDA.n1661 185
R1385 GNDA.n1664 GNDA.n1663 185
R1386 GNDA.n1666 GNDA.n1665 185
R1387 GNDA.n1668 GNDA.n1667 185
R1388 GNDA.n1650 GNDA.n1649 185
R1389 GNDA.n1644 GNDA.n1643 185
R1390 GNDA.n1642 GNDA.n1641 185
R1391 GNDA.n1637 GNDA.n1636 185
R1392 GNDA.n1635 GNDA.n1634 185
R1393 GNDA.n1629 GNDA.n1628 185
R1394 GNDA.n1624 GNDA.n875 185
R1395 GNDA.n1707 GNDA.n1706 185
R1396 GNDA.n874 GNDA.n872 185
R1397 GNDA.n1749 GNDA.n1748 185
R1398 GNDA.n1743 GNDA.n1742 185
R1399 GNDA.n1741 GNDA.n1740 185
R1400 GNDA.n1736 GNDA.n1735 185
R1401 GNDA.n1734 GNDA.n1733 185
R1402 GNDA.n1728 GNDA.n1727 185
R1403 GNDA.n1724 GNDA.n848 185
R1404 GNDA.n1808 GNDA.n1807 185
R1405 GNDA.n847 GNDA.n845 185
R1406 GNDA.n1004 GNDA.n1003 185
R1407 GNDA.n1006 GNDA.n1005 185
R1408 GNDA.n1008 GNDA.n1007 185
R1409 GNDA.n1010 GNDA.n1009 185
R1410 GNDA.n1012 GNDA.n1011 185
R1411 GNDA.n1014 GNDA.n1013 185
R1412 GNDA.n1016 GNDA.n1015 185
R1413 GNDA.n1018 GNDA.n1017 185
R1414 GNDA.n1019 GNDA.n967 185
R1415 GNDA.n986 GNDA.n985 185
R1416 GNDA.n988 GNDA.n987 185
R1417 GNDA.n990 GNDA.n989 185
R1418 GNDA.n992 GNDA.n991 185
R1419 GNDA.n994 GNDA.n993 185
R1420 GNDA.n996 GNDA.n995 185
R1421 GNDA.n998 GNDA.n997 185
R1422 GNDA.n1000 GNDA.n999 185
R1423 GNDA.n1002 GNDA.n1001 185
R1424 GNDA.n959 GNDA.n945 185
R1425 GNDA.n970 GNDA.n969 185
R1426 GNDA.n972 GNDA.n971 185
R1427 GNDA.n974 GNDA.n973 185
R1428 GNDA.n976 GNDA.n975 185
R1429 GNDA.n978 GNDA.n977 185
R1430 GNDA.n980 GNDA.n979 185
R1431 GNDA.n982 GNDA.n981 185
R1432 GNDA.n984 GNDA.n983 185
R1433 GNDA.n949 GNDA.n946 185
R1434 GNDA.n1050 GNDA.n1049 185
R1435 GNDA.n1024 GNDA.n948 185
R1436 GNDA.n1030 GNDA.n1029 185
R1437 GNDA.n1028 GNDA.n1023 185
R1438 GNDA.n1037 GNDA.n1036 185
R1439 GNDA.n1035 GNDA.n1022 185
R1440 GNDA.n1042 GNDA.n968 185
R1441 GNDA.n1046 GNDA.n1045 185
R1442 GNDA.n1971 GNDA.n1912 185
R1443 GNDA.n1985 GNDA.n1984 185
R1444 GNDA.n1983 GNDA.n1913 185
R1445 GNDA.n1982 GNDA.n1981 185
R1446 GNDA.n1980 GNDA.n1979 185
R1447 GNDA.n1978 GNDA.n1977 185
R1448 GNDA.n1976 GNDA.n1975 185
R1449 GNDA.n1974 GNDA.n1973 185
R1450 GNDA.n1972 GNDA.n1889 185
R1451 GNDA.n1954 GNDA.n1953 185
R1452 GNDA.n1956 GNDA.n1955 185
R1453 GNDA.n1958 GNDA.n1957 185
R1454 GNDA.n1960 GNDA.n1959 185
R1455 GNDA.n1962 GNDA.n1961 185
R1456 GNDA.n1964 GNDA.n1963 185
R1457 GNDA.n1966 GNDA.n1965 185
R1458 GNDA.n1968 GNDA.n1967 185
R1459 GNDA.n1970 GNDA.n1969 185
R1460 GNDA.n1936 GNDA.n1935 185
R1461 GNDA.n1938 GNDA.n1937 185
R1462 GNDA.n1940 GNDA.n1939 185
R1463 GNDA.n1942 GNDA.n1941 185
R1464 GNDA.n1944 GNDA.n1943 185
R1465 GNDA.n1946 GNDA.n1945 185
R1466 GNDA.n1948 GNDA.n1947 185
R1467 GNDA.n1950 GNDA.n1949 185
R1468 GNDA.n1952 GNDA.n1951 185
R1469 GNDA.n1934 GNDA.n1933 185
R1470 GNDA.n1928 GNDA.n1927 185
R1471 GNDA.n1926 GNDA.n1925 185
R1472 GNDA.n1921 GNDA.n1920 185
R1473 GNDA.n1916 GNDA.n1897 185
R1474 GNDA.n1989 GNDA.n1988 185
R1475 GNDA.n1896 GNDA.n1894 185
R1476 GNDA.n1995 GNDA.n1994 185
R1477 GNDA.n1997 GNDA.n1996 185
R1478 GNDA.n654 GNDA.n653 185
R1479 GNDA.n656 GNDA.n576 185
R1480 GNDA.n659 GNDA.n658 185
R1481 GNDA.n660 GNDA.n575 185
R1482 GNDA.n662 GNDA.n661 185
R1483 GNDA.n664 GNDA.n574 185
R1484 GNDA.n667 GNDA.n666 185
R1485 GNDA.n668 GNDA.n573 185
R1486 GNDA.n670 GNDA.n669 185
R1487 GNDA.n636 GNDA.n581 185
R1488 GNDA.n638 GNDA.n637 185
R1489 GNDA.n640 GNDA.n580 185
R1490 GNDA.n643 GNDA.n642 185
R1491 GNDA.n644 GNDA.n579 185
R1492 GNDA.n646 GNDA.n645 185
R1493 GNDA.n648 GNDA.n578 185
R1494 GNDA.n651 GNDA.n650 185
R1495 GNDA.n652 GNDA.n577 185
R1496 GNDA.n620 GNDA.n619 185
R1497 GNDA.n621 GNDA.n586 185
R1498 GNDA.n623 GNDA.n622 185
R1499 GNDA.n625 GNDA.n584 185
R1500 GNDA.n627 GNDA.n626 185
R1501 GNDA.n628 GNDA.n583 185
R1502 GNDA.n630 GNDA.n629 185
R1503 GNDA.n632 GNDA.n582 185
R1504 GNDA.n635 GNDA.n634 185
R1505 GNDA.n618 GNDA.n589 185
R1506 GNDA.n616 GNDA.n615 185
R1507 GNDA.n607 GNDA.n590 185
R1508 GNDA.n606 GNDA.n605 185
R1509 GNDA.n603 GNDA.n601 185
R1510 GNDA.n595 GNDA.n572 185
R1511 GNDA.n678 GNDA.n677 185
R1512 GNDA.n675 GNDA.n570 185
R1513 GNDA.n674 GNDA.n673 185
R1514 GNDA.n766 GNDA.n765 185
R1515 GNDA.n768 GNDA.n554 185
R1516 GNDA.n771 GNDA.n770 185
R1517 GNDA.n772 GNDA.n553 185
R1518 GNDA.n774 GNDA.n773 185
R1519 GNDA.n776 GNDA.n552 185
R1520 GNDA.n779 GNDA.n778 185
R1521 GNDA.n780 GNDA.n551 185
R1522 GNDA.n782 GNDA.n781 185
R1523 GNDA.n748 GNDA.n559 185
R1524 GNDA.n750 GNDA.n749 185
R1525 GNDA.n752 GNDA.n558 185
R1526 GNDA.n755 GNDA.n754 185
R1527 GNDA.n756 GNDA.n557 185
R1528 GNDA.n758 GNDA.n757 185
R1529 GNDA.n760 GNDA.n556 185
R1530 GNDA.n763 GNDA.n762 185
R1531 GNDA.n764 GNDA.n555 185
R1532 GNDA.n732 GNDA.n731 185
R1533 GNDA.n733 GNDA.n564 185
R1534 GNDA.n735 GNDA.n734 185
R1535 GNDA.n737 GNDA.n562 185
R1536 GNDA.n739 GNDA.n738 185
R1537 GNDA.n740 GNDA.n561 185
R1538 GNDA.n742 GNDA.n741 185
R1539 GNDA.n744 GNDA.n560 185
R1540 GNDA.n747 GNDA.n746 185
R1541 GNDA.n730 GNDA.n693 185
R1542 GNDA.n728 GNDA.n727 185
R1543 GNDA.n719 GNDA.n694 185
R1544 GNDA.n718 GNDA.n717 185
R1545 GNDA.n715 GNDA.n713 185
R1546 GNDA.n709 GNDA.n550 185
R1547 GNDA.n790 GNDA.n789 185
R1548 GNDA.n787 GNDA.n548 185
R1549 GNDA.n786 GNDA.n785 185
R1550 GNDA.n1590 GNDA.n1589 185
R1551 GNDA.n1592 GNDA.n1591 185
R1552 GNDA.n1594 GNDA.n1593 185
R1553 GNDA.n1596 GNDA.n1595 185
R1554 GNDA.n1598 GNDA.n1597 185
R1555 GNDA.n1600 GNDA.n1599 185
R1556 GNDA.n1602 GNDA.n1601 185
R1557 GNDA.n1604 GNDA.n1603 185
R1558 GNDA.n1605 GNDA.n1261 185
R1559 GNDA.n1572 GNDA.n1571 185
R1560 GNDA.n1574 GNDA.n1573 185
R1561 GNDA.n1576 GNDA.n1575 185
R1562 GNDA.n1578 GNDA.n1577 185
R1563 GNDA.n1580 GNDA.n1579 185
R1564 GNDA.n1582 GNDA.n1581 185
R1565 GNDA.n1584 GNDA.n1583 185
R1566 GNDA.n1586 GNDA.n1585 185
R1567 GNDA.n1588 GNDA.n1587 185
R1568 GNDA.n1554 GNDA.n1553 185
R1569 GNDA.n1556 GNDA.n1555 185
R1570 GNDA.n1558 GNDA.n1557 185
R1571 GNDA.n1560 GNDA.n1559 185
R1572 GNDA.n1562 GNDA.n1561 185
R1573 GNDA.n1564 GNDA.n1563 185
R1574 GNDA.n1566 GNDA.n1565 185
R1575 GNDA.n1568 GNDA.n1567 185
R1576 GNDA.n1570 GNDA.n1569 185
R1577 GNDA.n1552 GNDA.n1551 185
R1578 GNDA.n1546 GNDA.n1545 185
R1579 GNDA.n1544 GNDA.n1543 185
R1580 GNDA.n1539 GNDA.n1538 185
R1581 GNDA.n1537 GNDA.n1536 185
R1582 GNDA.n1531 GNDA.n1530 185
R1583 GNDA.n1526 GNDA.n1265 185
R1584 GNDA.n1609 GNDA.n1608 185
R1585 GNDA.n1264 GNDA.n1262 185
R1586 GNDA.n1395 GNDA.n1394 183.948
R1587 GNDA.n1423 GNDA.n1422 183.948
R1588 GNDA.n1396 GNDA.n1395 180.013
R1589 GNDA.n1422 GNDA.n1303 180.013
R1590 GNDA.n2049 GNDA.n231 175.546
R1591 GNDA.n2045 GNDA.n231 175.546
R1592 GNDA.n2045 GNDA.n2038 175.546
R1593 GNDA.n2041 GNDA.n2038 175.546
R1594 GNDA.n2041 GNDA.n58 175.546
R1595 GNDA.n2257 GNDA.n58 175.546
R1596 GNDA.n2257 GNDA.n56 175.546
R1597 GNDA.n2261 GNDA.n56 175.546
R1598 GNDA.n2261 GNDA.n53 175.546
R1599 GNDA.n2267 GNDA.n53 175.546
R1600 GNDA.n2267 GNDA.n54 175.546
R1601 GNDA.n2230 GNDA.n87 175.546
R1602 GNDA.n2245 GNDA.n2230 175.546
R1603 GNDA.n2245 GNDA.n2231 175.546
R1604 GNDA.n2241 GNDA.n2231 175.546
R1605 GNDA.n2241 GNDA.n62 175.546
R1606 GNDA.n2254 GNDA.n62 175.546
R1607 GNDA.n2254 GNDA.n63 175.546
R1608 GNDA.n105 GNDA.n63 175.546
R1609 GNDA.n110 GNDA.n105 175.546
R1610 GNDA.n110 GNDA.n48 175.546
R1611 GNDA.n2271 GNDA.n48 175.546
R1612 GNDA.n2097 GNDA.n2096 175.546
R1613 GNDA.n2093 GNDA.n2092 175.546
R1614 GNDA.n2090 GNDA.n2077 175.546
R1615 GNDA.n2086 GNDA.n2084 175.546
R1616 GNDA.n2188 GNDA.n171 175.546
R1617 GNDA.n2068 GNDA.n222 175.546
R1618 GNDA.n2064 GNDA.n2063 175.546
R1619 GNDA.n2061 GNDA.n225 175.546
R1620 GNDA.n2057 GNDA.n2056 175.546
R1621 GNDA.n2054 GNDA.n228 175.546
R1622 GNDA.n1115 GNDA.n1090 175.546
R1623 GNDA.n1115 GNDA.n1088 175.546
R1624 GNDA.n1120 GNDA.n1088 175.546
R1625 GNDA.n1120 GNDA.n1086 175.546
R1626 GNDA.n1124 GNDA.n1086 175.546
R1627 GNDA.n1125 GNDA.n1124 175.546
R1628 GNDA.n1127 GNDA.n1125 175.546
R1629 GNDA.n1127 GNDA.n1084 175.546
R1630 GNDA.n1132 GNDA.n1084 175.546
R1631 GNDA.n1132 GNDA.n1082 175.546
R1632 GNDA.n1136 GNDA.n1082 175.546
R1633 GNDA.n1229 GNDA.n1228 175.546
R1634 GNDA.n1145 GNDA.n1144 175.546
R1635 GNDA.n1151 GNDA.n1150 175.546
R1636 GNDA.n1158 GNDA.n1157 175.546
R1637 GNDA.n1166 GNDA.n1165 175.546
R1638 GNDA.n1253 GNDA.n920 175.546
R1639 GNDA.n1249 GNDA.n925 175.546
R1640 GNDA.n1247 GNDA.n1246 175.546
R1641 GNDA.n1243 GNDA.n1242 175.546
R1642 GNDA.n1239 GNDA.n1238 175.546
R1643 GNDA.n1093 GNDA.n1092 175.546
R1644 GNDA.n1097 GNDA.n1096 175.546
R1645 GNDA.n1101 GNDA.n1100 175.546
R1646 GNDA.n1105 GNDA.n1104 175.546
R1647 GNDA.n1109 GNDA.n1108 175.546
R1648 GNDA.n1430 GNDA.n1429 175.546
R1649 GNDA.n1435 GNDA.n1432 175.546
R1650 GNDA.n1438 GNDA.n1437 175.546
R1651 GNDA.n1444 GNDA.n1440 175.546
R1652 GNDA.n1448 GNDA.n1446 175.546
R1653 GNDA.n1397 GNDA.n1321 175.546
R1654 GNDA.n1402 GNDA.n1321 175.546
R1655 GNDA.n1402 GNDA.n1319 175.546
R1656 GNDA.n1406 GNDA.n1319 175.546
R1657 GNDA.n1407 GNDA.n1406 175.546
R1658 GNDA.n1407 GNDA.n1310 175.546
R1659 GNDA.n1414 GNDA.n1310 175.546
R1660 GNDA.n1414 GNDA.n1308 175.546
R1661 GNDA.n1419 GNDA.n1308 175.546
R1662 GNDA.n1419 GNDA.n1306 175.546
R1663 GNDA.n1424 GNDA.n1306 175.546
R1664 GNDA.n1710 GNDA.n1709 175.546
R1665 GNDA.n1626 GNDA.n1625 175.546
R1666 GNDA.n1632 GNDA.n1631 175.546
R1667 GNDA.n1639 GNDA.n1638 175.546
R1668 GNDA.n1647 GNDA.n1646 175.546
R1669 GNDA.n1360 GNDA.n1323 175.546
R1670 GNDA.n1360 GNDA.n1329 175.546
R1671 GNDA.n1356 GNDA.n1329 175.546
R1672 GNDA.n1356 GNDA.n1333 175.546
R1673 GNDA.n1352 GNDA.n1333 175.546
R1674 GNDA.n1352 GNDA.n1351 175.546
R1675 GNDA.n1351 GNDA.n1350 175.546
R1676 GNDA.n1350 GNDA.n1337 175.546
R1677 GNDA.n1346 GNDA.n1337 175.546
R1678 GNDA.n1346 GNDA.n870 175.546
R1679 GNDA.n1716 GNDA.n870 175.546
R1680 GNDA.n823 GNDA.n822 175.546
R1681 GNDA.n1832 GNDA.n822 175.546
R1682 GNDA.n1830 GNDA.n1829 175.546
R1683 GNDA.n1826 GNDA.n1825 175.546
R1684 GNDA.n1822 GNDA.n1821 175.546
R1685 GNDA.n1818 GNDA.n1817 175.546
R1686 GNDA.n1373 GNDA.n824 175.546
R1687 GNDA.n1373 GNDA.n1371 175.546
R1688 GNDA.n1377 GNDA.n1371 175.546
R1689 GNDA.n1377 GNDA.n1369 175.546
R1690 GNDA.n1381 GNDA.n1369 175.546
R1691 GNDA.n1381 GNDA.n1367 175.546
R1692 GNDA.n1385 GNDA.n1367 175.546
R1693 GNDA.n1385 GNDA.n1365 175.546
R1694 GNDA.n1389 GNDA.n1365 175.546
R1695 GNDA.n1389 GNDA.n1326 175.546
R1696 GNDA.n1393 GNDA.n1326 175.546
R1697 GNDA.n1810 GNDA.n827 175.546
R1698 GNDA.n1725 GNDA.n844 175.546
R1699 GNDA.n1731 GNDA.n1730 175.546
R1700 GNDA.n1738 GNDA.n1737 175.546
R1701 GNDA.n1746 GNDA.n1745 175.546
R1702 GNDA.n1363 GNDA.n1327 175.546
R1703 GNDA.n1330 GNDA.n1327 175.546
R1704 GNDA.n1331 GNDA.n1330 175.546
R1705 GNDA.n1334 GNDA.n1331 175.546
R1706 GNDA.n1335 GNDA.n1334 175.546
R1707 GNDA.n1339 GNDA.n1335 175.546
R1708 GNDA.n1340 GNDA.n1339 175.546
R1709 GNDA.n1341 GNDA.n1340 175.546
R1710 GNDA.n1342 GNDA.n1341 175.546
R1711 GNDA.n1342 GNDA.n868 175.546
R1712 GNDA.n1718 GNDA.n868 175.546
R1713 GNDA.n935 GNDA.n926 175.546
R1714 GNDA.n928 GNDA.n927 175.546
R1715 GNDA.n930 GNDA.n929 175.546
R1716 GNDA.n932 GNDA.n931 175.546
R1717 GNDA.n934 GNDA.n933 175.546
R1718 GNDA.n897 GNDA.n896 175.546
R1719 GNDA.n901 GNDA.n900 175.546
R1720 GNDA.n905 GNDA.n904 175.546
R1721 GNDA.n909 GNDA.n908 175.546
R1722 GNDA.n913 GNDA.n912 175.546
R1723 GNDA.n1043 GNDA.n468 175.546
R1724 GNDA.n1040 GNDA.n1039 175.546
R1725 GNDA.n1033 GNDA.n1032 175.546
R1726 GNDA.n1026 GNDA.n1025 175.546
R1727 GNDA.n1053 GNDA.n1052 175.546
R1728 GNDA.n2028 GNDA.n2027 175.546
R1729 GNDA.n2027 GNDA.n442 175.546
R1730 GNDA.n2023 GNDA.n2021 175.546
R1731 GNDA.n2019 GNDA.n450 175.546
R1732 GNDA.n2015 GNDA.n2013 175.546
R1733 GNDA.n2011 GNDA.n458 175.546
R1734 GNDA.n1870 GNDA.n1868 175.546
R1735 GNDA.n1874 GNDA.n1843 175.546
R1736 GNDA.n1878 GNDA.n1876 175.546
R1737 GNDA.n1882 GNDA.n1841 175.546
R1738 GNDA.n1885 GNDA.n1884 175.546
R1739 GNDA.n1862 GNDA.n1861 175.546
R1740 GNDA.n1858 GNDA.n1857 175.546
R1741 GNDA.n1854 GNDA.n1853 175.546
R1742 GNDA.n1850 GNDA.n1849 175.546
R1743 GNDA.n1846 GNDA.n435 175.546
R1744 GNDA.n1890 GNDA.n486 175.546
R1745 GNDA.n1992 GNDA.n1991 175.546
R1746 GNDA.n1918 GNDA.n1917 175.546
R1747 GNDA.n1923 GNDA.n1922 175.546
R1748 GNDA.n1931 GNDA.n1930 175.546
R1749 GNDA.n445 GNDA.n444 175.546
R1750 GNDA.n448 GNDA.n447 175.546
R1751 GNDA.n453 GNDA.n452 175.546
R1752 GNDA.n456 GNDA.n455 175.546
R1753 GNDA.n461 GNDA.n460 175.546
R1754 GNDA.n2073 GNDA.n2072 175.546
R1755 GNDA.n2075 GNDA.n2074 175.546
R1756 GNDA.n2079 GNDA.n2078 175.546
R1757 GNDA.n2081 GNDA.n2080 175.546
R1758 GNDA.n2186 GNDA.n173 175.546
R1759 GNDA.n2120 GNDA.n211 175.546
R1760 GNDA.n2116 GNDA.n2115 175.546
R1761 GNDA.n2113 GNDA.n214 175.546
R1762 GNDA.n2109 GNDA.n2108 175.546
R1763 GNDA.n2106 GNDA.n217 175.546
R1764 GNDA.n687 GNDA.n684 175.546
R1765 GNDA.n684 GNDA.n567 175.546
R1766 GNDA.n680 GNDA.n567 175.546
R1767 GNDA.n680 GNDA.n569 175.546
R1768 GNDA.n598 GNDA.n569 175.546
R1769 GNDA.n598 GNDA.n594 175.546
R1770 GNDA.n609 GNDA.n594 175.546
R1771 GNDA.n609 GNDA.n592 175.546
R1772 GNDA.n613 GNDA.n592 175.546
R1773 GNDA.n613 GNDA.n98 175.546
R1774 GNDA.n2195 GNDA.n98 175.546
R1775 GNDA.n2132 GNDA.n206 175.546
R1776 GNDA.n2133 GNDA.n2132 175.546
R1777 GNDA.n2135 GNDA.n205 175.546
R1778 GNDA.n2144 GNDA.n197 175.546
R1779 GNDA.n2147 GNDA.n2146 175.546
R1780 GNDA.n2149 GNDA.n195 175.546
R1781 GNDA.n816 GNDA.n500 175.546
R1782 GNDA.n814 GNDA.n813 175.546
R1783 GNDA.n810 GNDA.n809 175.546
R1784 GNDA.n806 GNDA.n805 175.546
R1785 GNDA.n802 GNDA.n801 175.546
R1786 GNDA.n527 GNDA.n526 175.546
R1787 GNDA.n524 GNDA.n504 175.546
R1788 GNDA.n520 GNDA.n519 175.546
R1789 GNDA.n517 GNDA.n507 175.546
R1790 GNDA.n513 GNDA.n512 175.546
R1791 GNDA.n797 GNDA.n796 175.546
R1792 GNDA.n796 GNDA.n532 175.546
R1793 GNDA.n792 GNDA.n532 175.546
R1794 GNDA.n792 GNDA.n547 175.546
R1795 GNDA.n710 GNDA.n547 175.546
R1796 GNDA.n710 GNDA.n708 175.546
R1797 GNDA.n721 GNDA.n708 175.546
R1798 GNDA.n721 GNDA.n696 175.546
R1799 GNDA.n725 GNDA.n696 175.546
R1800 GNDA.n725 GNDA.n700 175.546
R1801 GNDA.n700 GNDA.n190 175.546
R1802 GNDA.n2130 GNDA.n2128 175.546
R1803 GNDA.n2137 GNDA.n202 175.546
R1804 GNDA.n2140 GNDA.n2139 175.546
R1805 GNDA.n2142 GNDA.n200 175.546
R1806 GNDA.n2151 GNDA.n193 175.546
R1807 GNDA.n1467 GNDA.n1466 175.546
R1808 GNDA.n1463 GNDA.n1462 175.546
R1809 GNDA.n1460 GNDA.n1434 175.546
R1810 GNDA.n1456 GNDA.n1454 175.546
R1811 GNDA.n1452 GNDA.n1443 175.546
R1812 GNDA.n1474 GNDA.n1304 175.546
R1813 GNDA.n1474 GNDA.n1302 175.546
R1814 GNDA.n1478 GNDA.n1302 175.546
R1815 GNDA.n1478 GNDA.n1300 175.546
R1816 GNDA.n1482 GNDA.n1300 175.546
R1817 GNDA.n1482 GNDA.n1298 175.546
R1818 GNDA.n1486 GNDA.n1298 175.546
R1819 GNDA.n1486 GNDA.n1296 175.546
R1820 GNDA.n1490 GNDA.n1296 175.546
R1821 GNDA.n1490 GNDA.n1294 175.546
R1822 GNDA.n1494 GNDA.n1294 175.546
R1823 GNDA.n1612 GNDA.n1611 175.546
R1824 GNDA.n1528 GNDA.n1527 175.546
R1825 GNDA.n1534 GNDA.n1533 175.546
R1826 GNDA.n1541 GNDA.n1540 175.546
R1827 GNDA.n1549 GNDA.n1548 175.546
R1828 GNDA.n1498 GNDA.n1292 175.546
R1829 GNDA.n1498 GNDA.n1290 175.546
R1830 GNDA.n1503 GNDA.n1290 175.546
R1831 GNDA.n1503 GNDA.n1288 175.546
R1832 GNDA.n1507 GNDA.n1288 175.546
R1833 GNDA.n1508 GNDA.n1507 175.546
R1834 GNDA.n1510 GNDA.n1508 175.546
R1835 GNDA.n1510 GNDA.n1286 175.546
R1836 GNDA.n1515 GNDA.n1286 175.546
R1837 GNDA.n1515 GNDA.n1284 175.546
R1838 GNDA.n1519 GNDA.n1284 175.546
R1839 GNDA.n941 GNDA.n232 173.881
R1840 GNDA.t182 GNDA.n235 172.876
R1841 GNDA.t182 GNDA.n417 172.615
R1842 GNDA.n1255 GNDA.n232 171.624
R1843 GNDA.n381 GNDA.t127 166.898
R1844 GNDA.n381 GNDA.t107 166.898
R1845 GNDA.n115 GNDA.n114 163.333
R1846 GNDA.n1170 GNDA.n1169 163.333
R1847 GNDA.n1750 GNDA.n1749 163.333
R1848 GNDA.n1651 GNDA.n1650 163.333
R1849 GNDA.n959 GNDA.n949 163.333
R1850 GNDA.n1935 GNDA.n1934 163.333
R1851 GNDA.n619 GNDA.n618 163.333
R1852 GNDA.n731 GNDA.n730 163.333
R1853 GNDA.n1553 GNDA.n1552 163.333
R1854 GNDA.n344 GNDA.n343 161.3
R1855 GNDA.n11 GNDA.n10 161.3
R1856 GNDA.t332 GNDA.t136 159.71
R1857 GNDA.n147 GNDA.n146 150
R1858 GNDA.n143 GNDA.n142 150
R1859 GNDA.n139 GNDA.n138 150
R1860 GNDA.n135 GNDA.n134 150
R1861 GNDA.n131 GNDA.n130 150
R1862 GNDA.n127 GNDA.n126 150
R1863 GNDA.n123 GNDA.n122 150
R1864 GNDA.n119 GNDA.n118 150
R1865 GNDA.n2248 GNDA.n84 150
R1866 GNDA.n2238 GNDA.n2237 150
R1867 GNDA.n2251 GNDA.n65 150
R1868 GNDA.n101 GNDA.n66 150
R1869 GNDA.n155 GNDA.n154 150
R1870 GNDA.n159 GNDA.n158 150
R1871 GNDA.n163 GNDA.n162 150
R1872 GNDA.n165 GNDA.n83 150
R1873 GNDA.n1202 GNDA.n1201 150
R1874 GNDA.n1198 GNDA.n1197 150
R1875 GNDA.n1194 GNDA.n1193 150
R1876 GNDA.n1190 GNDA.n1189 150
R1877 GNDA.n1186 GNDA.n1185 150
R1878 GNDA.n1182 GNDA.n1181 150
R1879 GNDA.n1178 GNDA.n1177 150
R1880 GNDA.n1174 GNDA.n1173 150
R1881 GNDA.n1225 GNDA.n1063 150
R1882 GNDA.n1147 GNDA.n1064 150
R1883 GNDA.n1155 GNDA.n1154 150
R1884 GNDA.n1162 GNDA.n1161 150
R1885 GNDA.n1210 GNDA.n1209 150
R1886 GNDA.n1214 GNDA.n1213 150
R1887 GNDA.n1218 GNDA.n1217 150
R1888 GNDA.n1222 GNDA.n1221 150
R1889 GNDA.n1782 GNDA.n1781 150
R1890 GNDA.n1778 GNDA.n1777 150
R1891 GNDA.n1774 GNDA.n1773 150
R1892 GNDA.n1770 GNDA.n1769 150
R1893 GNDA.n1766 GNDA.n1765 150
R1894 GNDA.n1762 GNDA.n1761 150
R1895 GNDA.n1758 GNDA.n1757 150
R1896 GNDA.n1754 GNDA.n1753 150
R1897 GNDA.n1807 GNDA.n847 150
R1898 GNDA.n1727 GNDA.n848 150
R1899 GNDA.n1735 GNDA.n1734 150
R1900 GNDA.n1742 GNDA.n1741 150
R1901 GNDA.n1790 GNDA.n1789 150
R1902 GNDA.n1794 GNDA.n1793 150
R1903 GNDA.n1798 GNDA.n1797 150
R1904 GNDA.n1804 GNDA.n865 150
R1905 GNDA.n1683 GNDA.n1682 150
R1906 GNDA.n1679 GNDA.n1678 150
R1907 GNDA.n1675 GNDA.n1674 150
R1908 GNDA.n1671 GNDA.n1670 150
R1909 GNDA.n1667 GNDA.n1666 150
R1910 GNDA.n1663 GNDA.n1662 150
R1911 GNDA.n1659 GNDA.n1658 150
R1912 GNDA.n1655 GNDA.n1654 150
R1913 GNDA.n1706 GNDA.n874 150
R1914 GNDA.n1628 GNDA.n875 150
R1915 GNDA.n1636 GNDA.n1635 150
R1916 GNDA.n1643 GNDA.n1642 150
R1917 GNDA.n1691 GNDA.n1690 150
R1918 GNDA.n1695 GNDA.n1694 150
R1919 GNDA.n1699 GNDA.n1698 150
R1920 GNDA.n1703 GNDA.n1702 150
R1921 GNDA.n999 GNDA.n998 150
R1922 GNDA.n995 GNDA.n994 150
R1923 GNDA.n991 GNDA.n990 150
R1924 GNDA.n987 GNDA.n986 150
R1925 GNDA.n983 GNDA.n982 150
R1926 GNDA.n979 GNDA.n978 150
R1927 GNDA.n975 GNDA.n974 150
R1928 GNDA.n971 GNDA.n970 150
R1929 GNDA.n1046 GNDA.n968 150
R1930 GNDA.n1036 GNDA.n1035 150
R1931 GNDA.n1029 GNDA.n1028 150
R1932 GNDA.n1049 GNDA.n948 150
R1933 GNDA.n1007 GNDA.n1006 150
R1934 GNDA.n1011 GNDA.n1010 150
R1935 GNDA.n1015 GNDA.n1014 150
R1936 GNDA.n1017 GNDA.n967 150
R1937 GNDA.n1967 GNDA.n1966 150
R1938 GNDA.n1963 GNDA.n1962 150
R1939 GNDA.n1959 GNDA.n1958 150
R1940 GNDA.n1955 GNDA.n1954 150
R1941 GNDA.n1951 GNDA.n1950 150
R1942 GNDA.n1947 GNDA.n1946 150
R1943 GNDA.n1943 GNDA.n1942 150
R1944 GNDA.n1939 GNDA.n1938 150
R1945 GNDA.n1996 GNDA.n1995 150
R1946 GNDA.n1988 GNDA.n1896 150
R1947 GNDA.n1920 GNDA.n1897 150
R1948 GNDA.n1927 GNDA.n1926 150
R1949 GNDA.n1985 GNDA.n1913 150
R1950 GNDA.n1981 GNDA.n1980 150
R1951 GNDA.n1977 GNDA.n1976 150
R1952 GNDA.n1973 GNDA.n1972 150
R1953 GNDA.n650 GNDA.n648 150
R1954 GNDA.n646 GNDA.n579 150
R1955 GNDA.n642 GNDA.n640 150
R1956 GNDA.n638 GNDA.n581 150
R1957 GNDA.n634 GNDA.n632 150
R1958 GNDA.n630 GNDA.n583 150
R1959 GNDA.n626 GNDA.n625 150
R1960 GNDA.n623 GNDA.n586 150
R1961 GNDA.n675 GNDA.n674 150
R1962 GNDA.n677 GNDA.n572 150
R1963 GNDA.n605 GNDA.n603 150
R1964 GNDA.n616 GNDA.n590 150
R1965 GNDA.n658 GNDA.n656 150
R1966 GNDA.n662 GNDA.n575 150
R1967 GNDA.n666 GNDA.n664 150
R1968 GNDA.n670 GNDA.n573 150
R1969 GNDA.n762 GNDA.n760 150
R1970 GNDA.n758 GNDA.n557 150
R1971 GNDA.n754 GNDA.n752 150
R1972 GNDA.n750 GNDA.n559 150
R1973 GNDA.n746 GNDA.n744 150
R1974 GNDA.n742 GNDA.n561 150
R1975 GNDA.n738 GNDA.n737 150
R1976 GNDA.n735 GNDA.n564 150
R1977 GNDA.n787 GNDA.n786 150
R1978 GNDA.n789 GNDA.n550 150
R1979 GNDA.n717 GNDA.n715 150
R1980 GNDA.n728 GNDA.n694 150
R1981 GNDA.n770 GNDA.n768 150
R1982 GNDA.n774 GNDA.n553 150
R1983 GNDA.n778 GNDA.n776 150
R1984 GNDA.n782 GNDA.n551 150
R1985 GNDA.n1585 GNDA.n1584 150
R1986 GNDA.n1581 GNDA.n1580 150
R1987 GNDA.n1577 GNDA.n1576 150
R1988 GNDA.n1573 GNDA.n1572 150
R1989 GNDA.n1569 GNDA.n1568 150
R1990 GNDA.n1565 GNDA.n1564 150
R1991 GNDA.n1561 GNDA.n1560 150
R1992 GNDA.n1557 GNDA.n1556 150
R1993 GNDA.n1608 GNDA.n1264 150
R1994 GNDA.n1530 GNDA.n1265 150
R1995 GNDA.n1538 GNDA.n1537 150
R1996 GNDA.n1545 GNDA.n1544 150
R1997 GNDA.n1593 GNDA.n1592 150
R1998 GNDA.n1597 GNDA.n1596 150
R1999 GNDA.n1601 GNDA.n1600 150
R2000 GNDA.n1605 GNDA.n1604 150
R2001 GNDA.t163 GNDA.t45 148.435
R2002 GNDA.n317 GNDA.n316 148.017
R2003 GNDA.n334 GNDA.n333 148.017
R2004 GNDA.n2277 GNDA.n2276 148.017
R2005 GNDA.n2294 GNDA.n2293 148.017
R2006 GNDA.t135 GNDA.t43 144.9
R2007 GNDA.t60 GNDA.t337 139.599
R2008 GNDA.n1887 GNDA.n1886 132.721
R2009 GNDA.n530 GNDA.n495 132.721
R2010 GNDA.n2191 GNDA.n2190 124.832
R2011 GNDA.n1235 GNDA.n1234 124.832
R2012 GNDA.n1619 GNDA.n893 124.832
R2013 GNDA.n1716 GNDA.n1715 124.832
R2014 GNDA.n1719 GNDA.n1718 124.832
R2015 GNDA.n1058 GNDA.n943 124.832
R2016 GNDA.n2006 GNDA.n458 124.832
R2017 GNDA.n466 GNDA.n463 124.832
R2018 GNDA.n2184 GNDA.n99 124.832
R2019 GNDA.n566 GNDA.n195 124.832
R2020 GNDA.n2154 GNDA.n2153 124.832
R2021 GNDA.n1617 GNDA.n1260 124.832
R2022 GNDA.n23 GNDA.n22 118.861
R2023 GNDA.n26 GNDA.n25 118.861
R2024 GNDA.n29 GNDA.n28 118.861
R2025 GNDA.n33 GNDA.n32 118.861
R2026 GNDA.n36 GNDA.n35 118.861
R2027 GNDA.n39 GNDA.n38 118.861
R2028 GNDA.n295 GNDA.n294 118.861
R2029 GNDA.n298 GNDA.n297 118.861
R2030 GNDA.n301 GNDA.n300 118.861
R2031 GNDA.n305 GNDA.n304 118.861
R2032 GNDA.n308 GNDA.n307 118.861
R2033 GNDA.n311 GNDA.n310 118.861
R2034 GNDA.n2206 GNDA.t277 118.281
R2035 GNDA.n544 GNDA.t220 116.501
R2036 GNDA.n2157 GNDA.t210 116.501
R2037 GNDA.n2181 GNDA.t193 116.501
R2038 GNDA.n2163 GNDA.t241 116.501
R2039 GNDA.n2211 GNDA.t265 116.501
R2040 GNDA.n2226 GNDA.t185 116.501
R2041 GNDA.n93 GNDA.t338 115.948
R2042 GNDA.n1314 GNDA.t137 115.105
R2043 GNDA.n93 GNDA.t44 114.635
R2044 GNDA.n1315 GNDA.t134 114.635
R2045 GNDA.t91 GNDA.t130 109.35
R2046 GNDA.t249 GNDA.n252 107.805
R2047 GNDA.t259 GNDA.n17 107.805
R2048 GNDA.n183 GNDA.t192 103.15
R2049 GNDA.n686 GNDA.n685 100.025
R2050 GNDA.t182 GNDA.n182 47.6748
R2051 GNDA.n188 GNDA.n187 97.1505
R2052 GNDA.n537 GNDA.n536 97.1505
R2053 GNDA.n540 GNDA.n539 97.1505
R2054 GNDA.n2177 GNDA.n2176 97.1505
R2055 GNDA.n2173 GNDA.n2172 97.1505
R2056 GNDA.n2170 GNDA.n2169 97.1505
R2057 GNDA.n2166 GNDA.n2165 97.1505
R2058 GNDA.n2214 GNDA.n2213 97.1505
R2059 GNDA.n2218 GNDA.n2217 97.1505
R2060 GNDA.n2221 GNDA.n2220 97.1505
R2061 GNDA.t20 GNDA.t92 95.8263
R2062 GNDA.t166 GNDA.t20 95.8263
R2063 GNDA.t136 GNDA.t166 95.8263
R2064 GNDA.t270 GNDA.t332 95.8263
R2065 GNDA.t219 GNDA.n793 91.6889
R2066 GNDA.n109 GNDA.t151 91.6889
R2067 GNDA.n795 GNDA.t9 90.647
R2068 GNDA.n2048 GNDA.t182 90.5399
R2069 GNDA.n1372 GNDA.n413 88.5317
R2070 GNDA.n1372 GNDA.n1370 88.5317
R2071 GNDA.n1378 GNDA.n1370 88.5317
R2072 GNDA.n1379 GNDA.n1378 88.5317
R2073 GNDA.n1380 GNDA.n1379 88.5317
R2074 GNDA.n1386 GNDA.n1366 88.5317
R2075 GNDA.n1387 GNDA.n1386 88.5317
R2076 GNDA.n1388 GNDA.n1387 88.5317
R2077 GNDA.n1388 GNDA.n1325 88.5317
R2078 GNDA.n1394 GNDA.n1325 88.5317
R2079 GNDA.n1396 GNDA.n1320 88.5317
R2080 GNDA.n1403 GNDA.n1320 88.5317
R2081 GNDA.n1404 GNDA.n1403 88.5317
R2082 GNDA.n1405 GNDA.n1404 88.5317
R2083 GNDA.n1405 GNDA.n1311 88.5317
R2084 GNDA.n1413 GNDA.n1412 88.5317
R2085 GNDA.n1413 GNDA.n1307 88.5317
R2086 GNDA.n1420 GNDA.n1307 88.5317
R2087 GNDA.n1421 GNDA.n1420 88.5317
R2088 GNDA.n1423 GNDA.n1421 88.5317
R2089 GNDA.n1475 GNDA.n1303 88.5317
R2090 GNDA.n1476 GNDA.n1475 88.5317
R2091 GNDA.n1477 GNDA.n1476 88.5317
R2092 GNDA.n1477 GNDA.n1299 88.5317
R2093 GNDA.n1483 GNDA.n1299 88.5317
R2094 GNDA.n1485 GNDA.n1484 88.5317
R2095 GNDA.n1485 GNDA.n1295 88.5317
R2096 GNDA.n1491 GNDA.n1295 88.5317
R2097 GNDA.n1492 GNDA.n1491 88.5317
R2098 GNDA.n1493 GNDA.n1492 88.5317
R2099 GNDA.t271 GNDA.t25 87.8408
R2100 GNDA.t2 GNDA.t140 87.8408
R2101 GNDA.t117 GNDA.t10 87.8408
R2102 GNDA.t328 GNDA.t283 87.8408
R2103 GNDA.t324 GNDA.t326 87.8408
R2104 GNDA.t164 GNDA.t249 87.8408
R2105 GNDA.t147 GNDA.t164 87.8408
R2106 GNDA.t40 GNDA.t147 87.8408
R2107 GNDA.t46 GNDA.t78 87.8408
R2108 GNDA.t78 GNDA.t6 87.8408
R2109 GNDA.t48 GNDA.t80 87.8408
R2110 GNDA.t113 GNDA.t131 87.8408
R2111 GNDA.t131 GNDA.t259 87.8408
R2112 GNDA.t0 GNDA.t305 87.8408
R2113 GNDA.t298 GNDA.t308 87.8408
R2114 GNDA.t294 GNDA.t314 87.8408
R2115 GNDA.t82 GNDA.t304 87.8408
R2116 GNDA.t225 GNDA.t311 87.8408
R2117 GNDA.n707 GNDA.t159 85.4374
R2118 GNDA.t339 GNDA.n596 85.4374
R2119 GNDA.n1313 GNDA.n1312 84.306
R2120 GNDA.t187 GNDA.t205 83.848
R2121 GNDA.t196 GNDA.t199 83.848
R2122 GNDA.n2306 GNDA.t85 83.848
R2123 GNDA.t243 GNDA.t317 83.848
R2124 GNDA.n1089 GNDA.t133 81.9681
R2125 GNDA.n610 GNDA.t268 81.2697
R2126 GNDA.n1395 GNDA.n1324 80.9821
R2127 GNDA.n2275 GNDA.t327 80.7106
R2128 GNDA.t22 GNDA.t124 78.144
R2129 GNDA.t182 GNDA.n232 76.3879
R2130 GNDA.n2099 GNDA.n2098 76.3222
R2131 GNDA.n2096 GNDA.n2071 76.3222
R2132 GNDA.n2092 GNDA.n2091 76.3222
R2133 GNDA.n2085 GNDA.n2077 76.3222
R2134 GNDA.n2084 GNDA.n2083 76.3222
R2135 GNDA.n2189 GNDA.n2188 76.3222
R2136 GNDA.n2069 GNDA.n2068 76.3222
R2137 GNDA.n2064 GNDA.n224 76.3222
R2138 GNDA.n2062 GNDA.n2061 76.3222
R2139 GNDA.n2057 GNDA.n227 76.3222
R2140 GNDA.n2055 GNDA.n2054 76.3222
R2141 GNDA.n2050 GNDA.n230 76.3222
R2142 GNDA.n1233 GNDA.n474 76.3222
R2143 GNDA.n1228 GNDA.n473 76.3222
R2144 GNDA.n1145 GNDA.n472 76.3222
R2145 GNDA.n1151 GNDA.n471 76.3222
R2146 GNDA.n1157 GNDA.n470 76.3222
R2147 GNDA.n1166 GNDA.n469 76.3222
R2148 GNDA.n1257 GNDA.n1256 76.3222
R2149 GNDA.n1254 GNDA.n1253 76.3222
R2150 GNDA.n1249 GNDA.n924 76.3222
R2151 GNDA.n1246 GNDA.n923 76.3222
R2152 GNDA.n1242 GNDA.n922 76.3222
R2153 GNDA.n1238 GNDA.n921 76.3222
R2154 GNDA.n1092 GNDA.n418 76.3222
R2155 GNDA.n1096 GNDA.n419 76.3222
R2156 GNDA.n1100 GNDA.n420 76.3222
R2157 GNDA.n1104 GNDA.n421 76.3222
R2158 GNDA.n1108 GNDA.n422 76.3222
R2159 GNDA.n1111 GNDA.n423 76.3222
R2160 GNDA.n1429 GNDA.n1428 76.3222
R2161 GNDA.n1432 GNDA.n1431 76.3222
R2162 GNDA.n1437 GNDA.n1436 76.3222
R2163 GNDA.n1440 GNDA.n1439 76.3222
R2164 GNDA.n1446 GNDA.n1445 76.3222
R2165 GNDA.n1447 GNDA.n893 76.3222
R2166 GNDA.n1714 GNDA.n839 76.3222
R2167 GNDA.n1709 GNDA.n838 76.3222
R2168 GNDA.n1626 GNDA.n837 76.3222
R2169 GNDA.n1632 GNDA.n836 76.3222
R2170 GNDA.n1638 GNDA.n835 76.3222
R2171 GNDA.n1647 GNDA.n834 76.3222
R2172 GNDA.n1838 GNDA.n1837 76.3222
R2173 GNDA.n1832 GNDA.n489 76.3222
R2174 GNDA.n1829 GNDA.n490 76.3222
R2175 GNDA.n1825 GNDA.n491 76.3222
R2176 GNDA.n1821 GNDA.n492 76.3222
R2177 GNDA.n1814 GNDA.n1813 76.3222
R2178 GNDA.n1811 GNDA.n1810 76.3222
R2179 GNDA.n1725 GNDA.n843 76.3222
R2180 GNDA.n1731 GNDA.n842 76.3222
R2181 GNDA.n1737 GNDA.n841 76.3222
R2182 GNDA.n1746 GNDA.n840 76.3222
R2183 GNDA.n936 GNDA.n935 76.3222
R2184 GNDA.n937 GNDA.n927 76.3222
R2185 GNDA.n938 GNDA.n929 76.3222
R2186 GNDA.n939 GNDA.n931 76.3222
R2187 GNDA.n940 GNDA.n933 76.3222
R2188 GNDA.n943 GNDA.n942 76.3222
R2189 GNDA.n896 GNDA.n424 76.3222
R2190 GNDA.n900 GNDA.n425 76.3222
R2191 GNDA.n904 GNDA.n426 76.3222
R2192 GNDA.n908 GNDA.n427 76.3222
R2193 GNDA.n912 GNDA.n428 76.3222
R2194 GNDA.n916 GNDA.n429 76.3222
R2195 GNDA.n2005 GNDA.n2004 76.3222
R2196 GNDA.n1043 GNDA.n479 76.3222
R2197 GNDA.n1039 GNDA.n478 76.3222
R2198 GNDA.n1032 GNDA.n477 76.3222
R2199 GNDA.n1025 GNDA.n476 76.3222
R2200 GNDA.n1053 GNDA.n475 76.3222
R2201 GNDA.n2030 GNDA.n2029 76.3222
R2202 GNDA.n2022 GNDA.n442 76.3222
R2203 GNDA.n2021 GNDA.n2020 76.3222
R2204 GNDA.n2014 GNDA.n450 76.3222
R2205 GNDA.n2013 GNDA.n2012 76.3222
R2206 GNDA.n1867 GNDA.n1866 76.3222
R2207 GNDA.n1870 GNDA.n1869 76.3222
R2208 GNDA.n1875 GNDA.n1874 76.3222
R2209 GNDA.n1878 GNDA.n1877 76.3222
R2210 GNDA.n1883 GNDA.n1882 76.3222
R2211 GNDA.n1886 GNDA.n1885 76.3222
R2212 GNDA.n1862 GNDA.n430 76.3222
R2213 GNDA.n1858 GNDA.n431 76.3222
R2214 GNDA.n1854 GNDA.n432 76.3222
R2215 GNDA.n1850 GNDA.n433 76.3222
R2216 GNDA.n1846 GNDA.n434 76.3222
R2217 GNDA.n2035 GNDA.n2034 76.3222
R2218 GNDA.n2002 GNDA.n2001 76.3222
R2219 GNDA.n1890 GNDA.n485 76.3222
R2220 GNDA.n1991 GNDA.n484 76.3222
R2221 GNDA.n1918 GNDA.n483 76.3222
R2222 GNDA.n1922 GNDA.n482 76.3222
R2223 GNDA.n1931 GNDA.n481 76.3222
R2224 GNDA.n443 GNDA.n436 76.3222
R2225 GNDA.n446 GNDA.n445 76.3222
R2226 GNDA.n451 GNDA.n448 76.3222
R2227 GNDA.n454 GNDA.n453 76.3222
R2228 GNDA.n459 GNDA.n456 76.3222
R2229 GNDA.n462 GNDA.n461 76.3222
R2230 GNDA.n2072 GNDA.n174 76.3222
R2231 GNDA.n2074 GNDA.n175 76.3222
R2232 GNDA.n2078 GNDA.n176 76.3222
R2233 GNDA.n2080 GNDA.n177 76.3222
R2234 GNDA.n178 GNDA.n173 76.3222
R2235 GNDA.n2185 GNDA.n2184 76.3222
R2236 GNDA.n2121 GNDA.n2120 76.3222
R2237 GNDA.n2116 GNDA.n213 76.3222
R2238 GNDA.n2114 GNDA.n2113 76.3222
R2239 GNDA.n2109 GNDA.n216 76.3222
R2240 GNDA.n2107 GNDA.n2106 76.3222
R2241 GNDA.n2102 GNDA.n219 76.3222
R2242 GNDA.n2124 GNDA.n2123 76.3222
R2243 GNDA.n2134 GNDA.n2133 76.3222
R2244 GNDA.n205 GNDA.n204 76.3222
R2245 GNDA.n2145 GNDA.n2144 76.3222
R2246 GNDA.n2148 GNDA.n2147 76.3222
R2247 GNDA.n821 GNDA.n820 76.3222
R2248 GNDA.n816 GNDA.n499 76.3222
R2249 GNDA.n813 GNDA.n498 76.3222
R2250 GNDA.n809 GNDA.n497 76.3222
R2251 GNDA.n805 GNDA.n496 76.3222
R2252 GNDA.n801 GNDA.n495 76.3222
R2253 GNDA.n527 GNDA.n503 76.3222
R2254 GNDA.n525 GNDA.n524 76.3222
R2255 GNDA.n520 GNDA.n506 76.3222
R2256 GNDA.n518 GNDA.n517 76.3222
R2257 GNDA.n513 GNDA.n510 76.3222
R2258 GNDA.n511 GNDA.n208 76.3222
R2259 GNDA.n2127 GNDA.n2126 76.3222
R2260 GNDA.n2130 GNDA.n2129 76.3222
R2261 GNDA.n2138 GNDA.n2137 76.3222
R2262 GNDA.n2141 GNDA.n2140 76.3222
R2263 GNDA.n200 GNDA.n199 76.3222
R2264 GNDA.n2152 GNDA.n2151 76.3222
R2265 GNDA.n2153 GNDA.n2152 76.3222
R2266 GNDA.n199 GNDA.n193 76.3222
R2267 GNDA.n2142 GNDA.n2141 76.3222
R2268 GNDA.n2139 GNDA.n2138 76.3222
R2269 GNDA.n2129 GNDA.n202 76.3222
R2270 GNDA.n2128 GNDA.n2127 76.3222
R2271 GNDA.n2123 GNDA.n206 76.3222
R2272 GNDA.n2135 GNDA.n2134 76.3222
R2273 GNDA.n204 GNDA.n197 76.3222
R2274 GNDA.n2146 GNDA.n2145 76.3222
R2275 GNDA.n2149 GNDA.n2148 76.3222
R2276 GNDA.n463 GNDA.n462 76.3222
R2277 GNDA.n460 GNDA.n459 76.3222
R2278 GNDA.n455 GNDA.n454 76.3222
R2279 GNDA.n452 GNDA.n451 76.3222
R2280 GNDA.n447 GNDA.n446 76.3222
R2281 GNDA.n444 GNDA.n443 76.3222
R2282 GNDA.n2029 GNDA.n2028 76.3222
R2283 GNDA.n2023 GNDA.n2022 76.3222
R2284 GNDA.n2020 GNDA.n2019 76.3222
R2285 GNDA.n2015 GNDA.n2014 76.3222
R2286 GNDA.n2012 GNDA.n2011 76.3222
R2287 GNDA.n2035 GNDA.n435 76.3222
R2288 GNDA.n1849 GNDA.n434 76.3222
R2289 GNDA.n1853 GNDA.n433 76.3222
R2290 GNDA.n1857 GNDA.n432 76.3222
R2291 GNDA.n1861 GNDA.n431 76.3222
R2292 GNDA.n1845 GNDA.n430 76.3222
R2293 GNDA.n913 GNDA.n429 76.3222
R2294 GNDA.n909 GNDA.n428 76.3222
R2295 GNDA.n905 GNDA.n427 76.3222
R2296 GNDA.n901 GNDA.n426 76.3222
R2297 GNDA.n897 GNDA.n425 76.3222
R2298 GNDA.n441 GNDA.n424 76.3222
R2299 GNDA.n1109 GNDA.n423 76.3222
R2300 GNDA.n1105 GNDA.n422 76.3222
R2301 GNDA.n1101 GNDA.n421 76.3222
R2302 GNDA.n1097 GNDA.n420 76.3222
R2303 GNDA.n1093 GNDA.n419 76.3222
R2304 GNDA.n919 GNDA.n418 76.3222
R2305 GNDA.n1813 GNDA.n827 76.3222
R2306 GNDA.n1811 GNDA.n844 76.3222
R2307 GNDA.n1730 GNDA.n843 76.3222
R2308 GNDA.n1738 GNDA.n842 76.3222
R2309 GNDA.n1745 GNDA.n841 76.3222
R2310 GNDA.n1720 GNDA.n840 76.3222
R2311 GNDA.n1710 GNDA.n839 76.3222
R2312 GNDA.n1625 GNDA.n838 76.3222
R2313 GNDA.n1631 GNDA.n837 76.3222
R2314 GNDA.n1639 GNDA.n836 76.3222
R2315 GNDA.n1646 GNDA.n835 76.3222
R2316 GNDA.n1620 GNDA.n834 76.3222
R2317 GNDA.n512 GNDA.n511 76.3222
R2318 GNDA.n510 GNDA.n507 76.3222
R2319 GNDA.n519 GNDA.n518 76.3222
R2320 GNDA.n506 GNDA.n504 76.3222
R2321 GNDA.n526 GNDA.n525 76.3222
R2322 GNDA.n503 GNDA.n501 76.3222
R2323 GNDA.n219 GNDA.n217 76.3222
R2324 GNDA.n2108 GNDA.n2107 76.3222
R2325 GNDA.n216 GNDA.n214 76.3222
R2326 GNDA.n2115 GNDA.n2114 76.3222
R2327 GNDA.n213 GNDA.n211 76.3222
R2328 GNDA.n2122 GNDA.n2121 76.3222
R2329 GNDA.n230 GNDA.n228 76.3222
R2330 GNDA.n2056 GNDA.n2055 76.3222
R2331 GNDA.n227 GNDA.n225 76.3222
R2332 GNDA.n2063 GNDA.n2062 76.3222
R2333 GNDA.n224 GNDA.n222 76.3222
R2334 GNDA.n2070 GNDA.n2069 76.3222
R2335 GNDA.n2002 GNDA.n486 76.3222
R2336 GNDA.n1992 GNDA.n485 76.3222
R2337 GNDA.n1917 GNDA.n484 76.3222
R2338 GNDA.n1923 GNDA.n483 76.3222
R2339 GNDA.n1930 GNDA.n482 76.3222
R2340 GNDA.n481 GNDA.n480 76.3222
R2341 GNDA.n2004 GNDA.n468 76.3222
R2342 GNDA.n1040 GNDA.n479 76.3222
R2343 GNDA.n1033 GNDA.n478 76.3222
R2344 GNDA.n1026 GNDA.n477 76.3222
R2345 GNDA.n1052 GNDA.n476 76.3222
R2346 GNDA.n1057 GNDA.n475 76.3222
R2347 GNDA.n1229 GNDA.n474 76.3222
R2348 GNDA.n1144 GNDA.n473 76.3222
R2349 GNDA.n1150 GNDA.n472 76.3222
R2350 GNDA.n1158 GNDA.n471 76.3222
R2351 GNDA.n1165 GNDA.n470 76.3222
R2352 GNDA.n1139 GNDA.n469 76.3222
R2353 GNDA.n821 GNDA.n500 76.3222
R2354 GNDA.n814 GNDA.n499 76.3222
R2355 GNDA.n810 GNDA.n498 76.3222
R2356 GNDA.n806 GNDA.n497 76.3222
R2357 GNDA.n802 GNDA.n496 76.3222
R2358 GNDA.n1868 GNDA.n1867 76.3222
R2359 GNDA.n1869 GNDA.n1843 76.3222
R2360 GNDA.n1876 GNDA.n1875 76.3222
R2361 GNDA.n1877 GNDA.n1841 76.3222
R2362 GNDA.n1884 GNDA.n1883 76.3222
R2363 GNDA.n1838 GNDA.n823 76.3222
R2364 GNDA.n1830 GNDA.n489 76.3222
R2365 GNDA.n1826 GNDA.n490 76.3222
R2366 GNDA.n1822 GNDA.n491 76.3222
R2367 GNDA.n1818 GNDA.n492 76.3222
R2368 GNDA.n1469 GNDA.n1468 76.3222
R2369 GNDA.n1466 GNDA.n1427 76.3222
R2370 GNDA.n1462 GNDA.n1461 76.3222
R2371 GNDA.n1455 GNDA.n1434 76.3222
R2372 GNDA.n1454 GNDA.n1453 76.3222
R2373 GNDA.n1443 GNDA.n1442 76.3222
R2374 GNDA.n1616 GNDA.n833 76.3222
R2375 GNDA.n1611 GNDA.n832 76.3222
R2376 GNDA.n1528 GNDA.n831 76.3222
R2377 GNDA.n1534 GNDA.n830 76.3222
R2378 GNDA.n1540 GNDA.n829 76.3222
R2379 GNDA.n1549 GNDA.n828 76.3222
R2380 GNDA.n1612 GNDA.n833 76.3222
R2381 GNDA.n1527 GNDA.n832 76.3222
R2382 GNDA.n1533 GNDA.n831 76.3222
R2383 GNDA.n1541 GNDA.n830 76.3222
R2384 GNDA.n1548 GNDA.n829 76.3222
R2385 GNDA.n1522 GNDA.n828 76.3222
R2386 GNDA.n1448 GNDA.n1447 76.3222
R2387 GNDA.n1445 GNDA.n1444 76.3222
R2388 GNDA.n1439 GNDA.n1438 76.3222
R2389 GNDA.n1436 GNDA.n1435 76.3222
R2390 GNDA.n1431 GNDA.n1430 76.3222
R2391 GNDA.n1428 GNDA.n1425 76.3222
R2392 GNDA.n1468 GNDA.n1467 76.3222
R2393 GNDA.n1463 GNDA.n1427 76.3222
R2394 GNDA.n1461 GNDA.n1460 76.3222
R2395 GNDA.n1456 GNDA.n1455 76.3222
R2396 GNDA.n1453 GNDA.n1452 76.3222
R2397 GNDA.n1442 GNDA.n1260 76.3222
R2398 GNDA.n942 GNDA.n934 76.3222
R2399 GNDA.n940 GNDA.n932 76.3222
R2400 GNDA.n939 GNDA.n930 76.3222
R2401 GNDA.n938 GNDA.n928 76.3222
R2402 GNDA.n937 GNDA.n926 76.3222
R2403 GNDA.n936 GNDA.n917 76.3222
R2404 GNDA.n1256 GNDA.n920 76.3222
R2405 GNDA.n1254 GNDA.n925 76.3222
R2406 GNDA.n1247 GNDA.n924 76.3222
R2407 GNDA.n1243 GNDA.n923 76.3222
R2408 GNDA.n1239 GNDA.n922 76.3222
R2409 GNDA.n1235 GNDA.n921 76.3222
R2410 GNDA.n2186 GNDA.n2185 76.3222
R2411 GNDA.n2081 GNDA.n178 76.3222
R2412 GNDA.n2079 GNDA.n177 76.3222
R2413 GNDA.n2075 GNDA.n176 76.3222
R2414 GNDA.n2073 GNDA.n175 76.3222
R2415 GNDA.n2101 GNDA.n174 76.3222
R2416 GNDA.n2098 GNDA.n2097 76.3222
R2417 GNDA.n2093 GNDA.n2071 76.3222
R2418 GNDA.n2091 GNDA.n2090 76.3222
R2419 GNDA.n2086 GNDA.n2085 76.3222
R2420 GNDA.n2083 GNDA.n171 76.3222
R2421 GNDA.n2190 GNDA.n2189 76.3222
R2422 GNDA.t254 GNDA.t212 75.8626
R2423 GNDA.t317 GNDA.t23 75.8626
R2424 GNDA.n612 GNDA.t330 75.0183
R2425 GNDA.n134 GNDA.n72 74.5978
R2426 GNDA.n131 GNDA.n72 74.5978
R2427 GNDA.n1189 GNDA.n1070 74.5978
R2428 GNDA.n1186 GNDA.n1070 74.5978
R2429 GNDA.n1769 GNDA.n854 74.5978
R2430 GNDA.n1766 GNDA.n854 74.5978
R2431 GNDA.n1670 GNDA.n881 74.5978
R2432 GNDA.n1667 GNDA.n881 74.5978
R2433 GNDA.n986 GNDA.n955 74.5978
R2434 GNDA.n983 GNDA.n955 74.5978
R2435 GNDA.n1954 GNDA.n1902 74.5978
R2436 GNDA.n1951 GNDA.n1902 74.5978
R2437 GNDA.n633 GNDA.n581 74.5978
R2438 GNDA.n634 GNDA.n633 74.5978
R2439 GNDA.n745 GNDA.n559 74.5978
R2440 GNDA.n746 GNDA.n745 74.5978
R2441 GNDA.n1572 GNDA.n1271 74.5978
R2442 GNDA.n1569 GNDA.n1271 74.5978
R2443 GNDA.n2273 GNDA.t276 74.4678
R2444 GNDA.n2156 GNDA.t291 72.9344
R2445 GNDA.t28 GNDA.n682 70.8506
R2446 GNDA.t264 GNDA.n108 70.8506
R2447 GNDA.t143 GNDA.n106 69.8087
R2448 GNDA.n2249 GNDA.n2248 69.3109
R2449 GNDA.n2249 GNDA.n83 69.3109
R2450 GNDA.n1223 GNDA.n1063 69.3109
R2451 GNDA.n1223 GNDA.n1222 69.3109
R2452 GNDA.n1805 GNDA.n847 69.3109
R2453 GNDA.n1805 GNDA.n1804 69.3109
R2454 GNDA.n1704 GNDA.n874 69.3109
R2455 GNDA.n1704 GNDA.n1703 69.3109
R2456 GNDA.n1047 GNDA.n1046 69.3109
R2457 GNDA.n1047 GNDA.n967 69.3109
R2458 GNDA.n1996 GNDA.n1892 69.3109
R2459 GNDA.n1972 GNDA.n1892 69.3109
R2460 GNDA.n674 GNDA.n671 69.3109
R2461 GNDA.n671 GNDA.n670 69.3109
R2462 GNDA.n786 GNDA.n783 69.3109
R2463 GNDA.n783 GNDA.n782 69.3109
R2464 GNDA.n1606 GNDA.n1264 69.3109
R2465 GNDA.n1606 GNDA.n1605 69.3109
R2466 GNDA.t25 GNDA.t286 67.8771
R2467 GNDA.t95 GNDA.t324 67.8771
R2468 GNDA.t38 GNDA.n286 67.8771
R2469 GNDA.n2305 GNDA.t98 67.8771
R2470 GNDA.n257 GNDA.t114 67.8771
R2471 GNDA.n2292 GNDA.t212 67.8771
R2472 GNDA.t58 GNDA.n2273 66.8849
R2473 GNDA.t227 GNDA.n82 65.8183
R2474 GNDA.t227 GNDA.n81 65.8183
R2475 GNDA.t227 GNDA.n80 65.8183
R2476 GNDA.t227 GNDA.n79 65.8183
R2477 GNDA.t227 GNDA.n70 65.8183
R2478 GNDA.t227 GNDA.n77 65.8183
R2479 GNDA.t227 GNDA.n68 65.8183
R2480 GNDA.t227 GNDA.n78 65.8183
R2481 GNDA.t227 GNDA.n76 65.8183
R2482 GNDA.t227 GNDA.n75 65.8183
R2483 GNDA.t227 GNDA.n74 65.8183
R2484 GNDA.t227 GNDA.n73 65.8183
R2485 GNDA.t227 GNDA.n71 65.8183
R2486 GNDA.n2250 GNDA.t227 65.8183
R2487 GNDA.t227 GNDA.n69 65.8183
R2488 GNDA.t227 GNDA.n67 65.8183
R2489 GNDA.t223 GNDA.n1080 65.8183
R2490 GNDA.t223 GNDA.n1079 65.8183
R2491 GNDA.t223 GNDA.n1078 65.8183
R2492 GNDA.t223 GNDA.n1077 65.8183
R2493 GNDA.t223 GNDA.n1068 65.8183
R2494 GNDA.t223 GNDA.n1075 65.8183
R2495 GNDA.t223 GNDA.n1065 65.8183
R2496 GNDA.t223 GNDA.n1076 65.8183
R2497 GNDA.t223 GNDA.n1074 65.8183
R2498 GNDA.t223 GNDA.n1073 65.8183
R2499 GNDA.t223 GNDA.n1072 65.8183
R2500 GNDA.t223 GNDA.n1071 65.8183
R2501 GNDA.t223 GNDA.n1069 65.8183
R2502 GNDA.t223 GNDA.n1067 65.8183
R2503 GNDA.t223 GNDA.n1066 65.8183
R2504 GNDA.n1224 GNDA.t223 65.8183
R2505 GNDA.t194 GNDA.n864 65.8183
R2506 GNDA.t194 GNDA.n863 65.8183
R2507 GNDA.t194 GNDA.n862 65.8183
R2508 GNDA.t194 GNDA.n861 65.8183
R2509 GNDA.t194 GNDA.n852 65.8183
R2510 GNDA.t194 GNDA.n859 65.8183
R2511 GNDA.t194 GNDA.n849 65.8183
R2512 GNDA.t194 GNDA.n860 65.8183
R2513 GNDA.t194 GNDA.n858 65.8183
R2514 GNDA.t194 GNDA.n857 65.8183
R2515 GNDA.t194 GNDA.n856 65.8183
R2516 GNDA.t194 GNDA.n855 65.8183
R2517 GNDA.t181 GNDA.n891 65.8183
R2518 GNDA.t181 GNDA.n890 65.8183
R2519 GNDA.t181 GNDA.n889 65.8183
R2520 GNDA.t181 GNDA.n888 65.8183
R2521 GNDA.t181 GNDA.n879 65.8183
R2522 GNDA.t181 GNDA.n886 65.8183
R2523 GNDA.t181 GNDA.n876 65.8183
R2524 GNDA.t181 GNDA.n887 65.8183
R2525 GNDA.t181 GNDA.n885 65.8183
R2526 GNDA.t181 GNDA.n884 65.8183
R2527 GNDA.t181 GNDA.n883 65.8183
R2528 GNDA.t181 GNDA.n882 65.8183
R2529 GNDA.t181 GNDA.n880 65.8183
R2530 GNDA.t181 GNDA.n878 65.8183
R2531 GNDA.t181 GNDA.n877 65.8183
R2532 GNDA.n1705 GNDA.t181 65.8183
R2533 GNDA.t194 GNDA.n853 65.8183
R2534 GNDA.t194 GNDA.n851 65.8183
R2535 GNDA.t194 GNDA.n850 65.8183
R2536 GNDA.n1806 GNDA.t194 65.8183
R2537 GNDA.t201 GNDA.n966 65.8183
R2538 GNDA.t201 GNDA.n965 65.8183
R2539 GNDA.t201 GNDA.n964 65.8183
R2540 GNDA.t201 GNDA.n963 65.8183
R2541 GNDA.t201 GNDA.n954 65.8183
R2542 GNDA.t201 GNDA.n961 65.8183
R2543 GNDA.t201 GNDA.n951 65.8183
R2544 GNDA.t201 GNDA.n962 65.8183
R2545 GNDA.t201 GNDA.n960 65.8183
R2546 GNDA.t201 GNDA.n958 65.8183
R2547 GNDA.t201 GNDA.n957 65.8183
R2548 GNDA.t201 GNDA.n956 65.8183
R2549 GNDA.n1048 GNDA.t201 65.8183
R2550 GNDA.t201 GNDA.n953 65.8183
R2551 GNDA.t201 GNDA.n952 65.8183
R2552 GNDA.t201 GNDA.n950 65.8183
R2553 GNDA.t221 GNDA.n1986 65.8183
R2554 GNDA.t221 GNDA.n1911 65.8183
R2555 GNDA.t221 GNDA.n1910 65.8183
R2556 GNDA.t221 GNDA.n1909 65.8183
R2557 GNDA.t221 GNDA.n1900 65.8183
R2558 GNDA.t221 GNDA.n1907 65.8183
R2559 GNDA.t221 GNDA.n1898 65.8183
R2560 GNDA.t221 GNDA.n1908 65.8183
R2561 GNDA.t221 GNDA.n1906 65.8183
R2562 GNDA.t221 GNDA.n1905 65.8183
R2563 GNDA.t221 GNDA.n1904 65.8183
R2564 GNDA.t221 GNDA.n1903 65.8183
R2565 GNDA.t221 GNDA.n1901 65.8183
R2566 GNDA.t221 GNDA.n1899 65.8183
R2567 GNDA.n1987 GNDA.t221 65.8183
R2568 GNDA.t221 GNDA.n1893 65.8183
R2569 GNDA.n655 GNDA.t202 65.8183
R2570 GNDA.n657 GNDA.t202 65.8183
R2571 GNDA.n663 GNDA.t202 65.8183
R2572 GNDA.n665 GNDA.t202 65.8183
R2573 GNDA.n639 GNDA.t202 65.8183
R2574 GNDA.n641 GNDA.t202 65.8183
R2575 GNDA.n647 GNDA.t202 65.8183
R2576 GNDA.n649 GNDA.t202 65.8183
R2577 GNDA.n587 GNDA.t202 65.8183
R2578 GNDA.n624 GNDA.t202 65.8183
R2579 GNDA.n585 GNDA.t202 65.8183
R2580 GNDA.n631 GNDA.t202 65.8183
R2581 GNDA.n617 GNDA.t202 65.8183
R2582 GNDA.n604 GNDA.t202 65.8183
R2583 GNDA.n602 GNDA.t202 65.8183
R2584 GNDA.n676 GNDA.t202 65.8183
R2585 GNDA.n767 GNDA.t222 65.8183
R2586 GNDA.n769 GNDA.t222 65.8183
R2587 GNDA.n775 GNDA.t222 65.8183
R2588 GNDA.n777 GNDA.t222 65.8183
R2589 GNDA.n751 GNDA.t222 65.8183
R2590 GNDA.n753 GNDA.t222 65.8183
R2591 GNDA.n759 GNDA.t222 65.8183
R2592 GNDA.n761 GNDA.t222 65.8183
R2593 GNDA.n692 GNDA.t222 65.8183
R2594 GNDA.n736 GNDA.t222 65.8183
R2595 GNDA.n563 GNDA.t222 65.8183
R2596 GNDA.n743 GNDA.t222 65.8183
R2597 GNDA.n729 GNDA.t222 65.8183
R2598 GNDA.n716 GNDA.t222 65.8183
R2599 GNDA.n714 GNDA.t222 65.8183
R2600 GNDA.n788 GNDA.t222 65.8183
R2601 GNDA.t207 GNDA.n1281 65.8183
R2602 GNDA.t207 GNDA.n1280 65.8183
R2603 GNDA.t207 GNDA.n1279 65.8183
R2604 GNDA.t207 GNDA.n1278 65.8183
R2605 GNDA.t207 GNDA.n1269 65.8183
R2606 GNDA.t207 GNDA.n1276 65.8183
R2607 GNDA.t207 GNDA.n1266 65.8183
R2608 GNDA.t207 GNDA.n1277 65.8183
R2609 GNDA.t207 GNDA.n1275 65.8183
R2610 GNDA.t207 GNDA.n1274 65.8183
R2611 GNDA.t207 GNDA.n1273 65.8183
R2612 GNDA.t207 GNDA.n1272 65.8183
R2613 GNDA.t207 GNDA.n1270 65.8183
R2614 GNDA.t207 GNDA.n1268 65.8183
R2615 GNDA.t207 GNDA.n1267 65.8183
R2616 GNDA.n1607 GNDA.t207 65.8183
R2617 GNDA.n546 GNDA.t3 65.641
R2618 GNDA.n723 GNDA.t148 65.641
R2619 GNDA.n681 GNDA.t41 64.5991
R2620 GNDA.t184 GNDA.n2228 64.5991
R2621 GNDA.n2277 GNDA.n2275 63.8843
R2622 GNDA.t327 GNDA.t91 62.4857
R2623 GNDA.t320 GNDA.t54 62.4857
R2624 GNDA.t54 GNDA.t19 62.4857
R2625 GNDA.n349 GNDA.t262 62.2505
R2626 GNDA.n351 GNDA.t250 62.2505
R2627 GNDA.n346 GNDA.t190 62.2505
R2628 GNDA.n287 GNDA.t174 62.2505
R2629 GNDA.n339 GNDA.t257 62.2505
R2630 GNDA.n2307 GNDA.t180 62.2505
R2631 GNDA.n255 GNDA.t233 62.2505
R2632 GNDA.n12 GNDA.t252 62.2505
R2633 GNDA.n9 GNDA.t238 62.2505
R2634 GNDA.n16 GNDA.t267 62.2505
R2635 GNDA.n2304 GNDA.t247 62.2505
R2636 GNDA.n4 GNDA.t260 62.2505
R2637 GNDA.n611 GNDA.t122 60.4315
R2638 GNDA.t312 GNDA.n2232 60.4315
R2639 GNDA.n318 GNDA.t187 59.8916
R2640 GNDA.n332 GNDA.t199 59.8916
R2641 GNDA.t321 GNDA.t0 59.8916
R2642 GNDA.t304 GNDA.t93 59.8916
R2643 GNDA.t182 GNDA.n406 59.4672
R2644 GNDA.n2279 GNDA.n2278 59.2425
R2645 GNDA.n2292 GNDA.n2291 59.2425
R2646 GNDA.n319 GNDA.n318 59.2425
R2647 GNDA.n332 GNDA.n331 59.2425
R2648 GNDA.t227 GNDA.n2249 57.8461
R2649 GNDA.t223 GNDA.n1223 57.8461
R2650 GNDA.t181 GNDA.n1704 57.8461
R2651 GNDA.t194 GNDA.n1805 57.8461
R2652 GNDA.t201 GNDA.n1047 57.8461
R2653 GNDA.t221 GNDA.n1892 57.8461
R2654 GNDA.n671 GNDA.t202 57.8461
R2655 GNDA.n783 GNDA.t222 57.8461
R2656 GNDA.t207 GNDA.n1606 57.8461
R2657 GNDA.t290 GNDA.t299 57.3057
R2658 GNDA.t240 GNDA.n96 57.3057
R2659 GNDA.t141 GNDA.t144 57.3057
R2660 GNDA.n1817 GNDA.n493 56.3995
R2661 GNDA.n1815 GNDA.n493 56.3995
R2662 GNDA.n54 GNDA.n51 56.3995
R2663 GNDA.n1137 GNDA.n1136 56.3995
R2664 GNDA.n530 GNDA.n494 56.3995
R2665 GNDA.n1887 GNDA.n487 56.3995
R2666 GNDA.n51 GNDA.n49 56.3995
R2667 GNDA.n1138 GNDA.n1137 56.3995
R2668 GNDA.n1520 GNDA.n1519 56.3995
R2669 GNDA.n1521 GNDA.n1520 56.3995
R2670 GNDA.n2278 GNDA.n2277 55.8989
R2671 GNDA.n2197 GNDA.n2196 55.2219
R2672 GNDA.t126 GNDA.n2243 55.2219
R2673 GNDA.t227 GNDA.n72 55.2026
R2674 GNDA.t223 GNDA.n1070 55.2026
R2675 GNDA.t194 GNDA.n854 55.2026
R2676 GNDA.t181 GNDA.n881 55.2026
R2677 GNDA.t201 GNDA.n955 55.2026
R2678 GNDA.t221 GNDA.n1902 55.2026
R2679 GNDA.n633 GNDA.t202 55.2026
R2680 GNDA.n745 GNDA.t222 55.2026
R2681 GNDA.t207 GNDA.n1271 55.2026
R2682 GNDA.n699 GNDA.t209 54.18
R2683 GNDA.t87 GNDA.n611 54.18
R2684 GNDA.n150 GNDA.n78 53.3664
R2685 GNDA.n146 GNDA.n68 53.3664
R2686 GNDA.n142 GNDA.n77 53.3664
R2687 GNDA.n138 GNDA.n70 53.3664
R2688 GNDA.n127 GNDA.n73 53.3664
R2689 GNDA.n123 GNDA.n74 53.3664
R2690 GNDA.n119 GNDA.n75 53.3664
R2691 GNDA.n115 GNDA.n76 53.3664
R2692 GNDA.n84 GNDA.n67 53.3664
R2693 GNDA.n2238 GNDA.n69 53.3664
R2694 GNDA.n2251 GNDA.n2250 53.3664
R2695 GNDA.n101 GNDA.n71 53.3664
R2696 GNDA.n154 GNDA.n82 53.3664
R2697 GNDA.n155 GNDA.n81 53.3664
R2698 GNDA.n159 GNDA.n80 53.3664
R2699 GNDA.n163 GNDA.n79 53.3664
R2700 GNDA.n151 GNDA.n82 53.3664
R2701 GNDA.n158 GNDA.n81 53.3664
R2702 GNDA.n162 GNDA.n80 53.3664
R2703 GNDA.n165 GNDA.n79 53.3664
R2704 GNDA.n135 GNDA.n70 53.3664
R2705 GNDA.n139 GNDA.n77 53.3664
R2706 GNDA.n143 GNDA.n68 53.3664
R2707 GNDA.n147 GNDA.n78 53.3664
R2708 GNDA.n118 GNDA.n76 53.3664
R2709 GNDA.n122 GNDA.n75 53.3664
R2710 GNDA.n126 GNDA.n74 53.3664
R2711 GNDA.n130 GNDA.n73 53.3664
R2712 GNDA.n114 GNDA.n71 53.3664
R2713 GNDA.n2250 GNDA.n66 53.3664
R2714 GNDA.n69 GNDA.n65 53.3664
R2715 GNDA.n2237 GNDA.n67 53.3664
R2716 GNDA.n1205 GNDA.n1076 53.3664
R2717 GNDA.n1201 GNDA.n1065 53.3664
R2718 GNDA.n1197 GNDA.n1075 53.3664
R2719 GNDA.n1193 GNDA.n1068 53.3664
R2720 GNDA.n1182 GNDA.n1071 53.3664
R2721 GNDA.n1178 GNDA.n1072 53.3664
R2722 GNDA.n1174 GNDA.n1073 53.3664
R2723 GNDA.n1170 GNDA.n1074 53.3664
R2724 GNDA.n1225 GNDA.n1224 53.3664
R2725 GNDA.n1147 GNDA.n1066 53.3664
R2726 GNDA.n1155 GNDA.n1067 53.3664
R2727 GNDA.n1162 GNDA.n1069 53.3664
R2728 GNDA.n1209 GNDA.n1080 53.3664
R2729 GNDA.n1210 GNDA.n1079 53.3664
R2730 GNDA.n1214 GNDA.n1078 53.3664
R2731 GNDA.n1218 GNDA.n1077 53.3664
R2732 GNDA.n1206 GNDA.n1080 53.3664
R2733 GNDA.n1213 GNDA.n1079 53.3664
R2734 GNDA.n1217 GNDA.n1078 53.3664
R2735 GNDA.n1221 GNDA.n1077 53.3664
R2736 GNDA.n1190 GNDA.n1068 53.3664
R2737 GNDA.n1194 GNDA.n1075 53.3664
R2738 GNDA.n1198 GNDA.n1065 53.3664
R2739 GNDA.n1202 GNDA.n1076 53.3664
R2740 GNDA.n1173 GNDA.n1074 53.3664
R2741 GNDA.n1177 GNDA.n1073 53.3664
R2742 GNDA.n1181 GNDA.n1072 53.3664
R2743 GNDA.n1185 GNDA.n1071 53.3664
R2744 GNDA.n1169 GNDA.n1069 53.3664
R2745 GNDA.n1161 GNDA.n1067 53.3664
R2746 GNDA.n1154 GNDA.n1066 53.3664
R2747 GNDA.n1224 GNDA.n1064 53.3664
R2748 GNDA.n1785 GNDA.n860 53.3664
R2749 GNDA.n1781 GNDA.n849 53.3664
R2750 GNDA.n1777 GNDA.n859 53.3664
R2751 GNDA.n1773 GNDA.n852 53.3664
R2752 GNDA.n1762 GNDA.n855 53.3664
R2753 GNDA.n1758 GNDA.n856 53.3664
R2754 GNDA.n1754 GNDA.n857 53.3664
R2755 GNDA.n1750 GNDA.n858 53.3664
R2756 GNDA.n1807 GNDA.n1806 53.3664
R2757 GNDA.n1727 GNDA.n850 53.3664
R2758 GNDA.n1735 GNDA.n851 53.3664
R2759 GNDA.n1742 GNDA.n853 53.3664
R2760 GNDA.n1789 GNDA.n864 53.3664
R2761 GNDA.n1790 GNDA.n863 53.3664
R2762 GNDA.n1794 GNDA.n862 53.3664
R2763 GNDA.n1798 GNDA.n861 53.3664
R2764 GNDA.n1786 GNDA.n864 53.3664
R2765 GNDA.n1793 GNDA.n863 53.3664
R2766 GNDA.n1797 GNDA.n862 53.3664
R2767 GNDA.n865 GNDA.n861 53.3664
R2768 GNDA.n1770 GNDA.n852 53.3664
R2769 GNDA.n1774 GNDA.n859 53.3664
R2770 GNDA.n1778 GNDA.n849 53.3664
R2771 GNDA.n1782 GNDA.n860 53.3664
R2772 GNDA.n1753 GNDA.n858 53.3664
R2773 GNDA.n1757 GNDA.n857 53.3664
R2774 GNDA.n1761 GNDA.n856 53.3664
R2775 GNDA.n1765 GNDA.n855 53.3664
R2776 GNDA.n1686 GNDA.n887 53.3664
R2777 GNDA.n1682 GNDA.n876 53.3664
R2778 GNDA.n1678 GNDA.n886 53.3664
R2779 GNDA.n1674 GNDA.n879 53.3664
R2780 GNDA.n1663 GNDA.n882 53.3664
R2781 GNDA.n1659 GNDA.n883 53.3664
R2782 GNDA.n1655 GNDA.n884 53.3664
R2783 GNDA.n1651 GNDA.n885 53.3664
R2784 GNDA.n1706 GNDA.n1705 53.3664
R2785 GNDA.n1628 GNDA.n877 53.3664
R2786 GNDA.n1636 GNDA.n878 53.3664
R2787 GNDA.n1643 GNDA.n880 53.3664
R2788 GNDA.n1690 GNDA.n891 53.3664
R2789 GNDA.n1691 GNDA.n890 53.3664
R2790 GNDA.n1695 GNDA.n889 53.3664
R2791 GNDA.n1699 GNDA.n888 53.3664
R2792 GNDA.n1687 GNDA.n891 53.3664
R2793 GNDA.n1694 GNDA.n890 53.3664
R2794 GNDA.n1698 GNDA.n889 53.3664
R2795 GNDA.n1702 GNDA.n888 53.3664
R2796 GNDA.n1671 GNDA.n879 53.3664
R2797 GNDA.n1675 GNDA.n886 53.3664
R2798 GNDA.n1679 GNDA.n876 53.3664
R2799 GNDA.n1683 GNDA.n887 53.3664
R2800 GNDA.n1654 GNDA.n885 53.3664
R2801 GNDA.n1658 GNDA.n884 53.3664
R2802 GNDA.n1662 GNDA.n883 53.3664
R2803 GNDA.n1666 GNDA.n882 53.3664
R2804 GNDA.n1650 GNDA.n880 53.3664
R2805 GNDA.n1642 GNDA.n878 53.3664
R2806 GNDA.n1635 GNDA.n877 53.3664
R2807 GNDA.n1705 GNDA.n875 53.3664
R2808 GNDA.n1749 GNDA.n853 53.3664
R2809 GNDA.n1741 GNDA.n851 53.3664
R2810 GNDA.n1734 GNDA.n850 53.3664
R2811 GNDA.n1806 GNDA.n848 53.3664
R2812 GNDA.n1002 GNDA.n962 53.3664
R2813 GNDA.n998 GNDA.n951 53.3664
R2814 GNDA.n994 GNDA.n961 53.3664
R2815 GNDA.n990 GNDA.n954 53.3664
R2816 GNDA.n979 GNDA.n956 53.3664
R2817 GNDA.n975 GNDA.n957 53.3664
R2818 GNDA.n971 GNDA.n958 53.3664
R2819 GNDA.n960 GNDA.n959 53.3664
R2820 GNDA.n968 GNDA.n950 53.3664
R2821 GNDA.n1036 GNDA.n952 53.3664
R2822 GNDA.n1029 GNDA.n953 53.3664
R2823 GNDA.n1049 GNDA.n1048 53.3664
R2824 GNDA.n1006 GNDA.n966 53.3664
R2825 GNDA.n1007 GNDA.n965 53.3664
R2826 GNDA.n1011 GNDA.n964 53.3664
R2827 GNDA.n1015 GNDA.n963 53.3664
R2828 GNDA.n1003 GNDA.n966 53.3664
R2829 GNDA.n1010 GNDA.n965 53.3664
R2830 GNDA.n1014 GNDA.n964 53.3664
R2831 GNDA.n1017 GNDA.n963 53.3664
R2832 GNDA.n987 GNDA.n954 53.3664
R2833 GNDA.n991 GNDA.n961 53.3664
R2834 GNDA.n995 GNDA.n951 53.3664
R2835 GNDA.n999 GNDA.n962 53.3664
R2836 GNDA.n970 GNDA.n960 53.3664
R2837 GNDA.n974 GNDA.n958 53.3664
R2838 GNDA.n978 GNDA.n957 53.3664
R2839 GNDA.n982 GNDA.n956 53.3664
R2840 GNDA.n1048 GNDA.n949 53.3664
R2841 GNDA.n953 GNDA.n948 53.3664
R2842 GNDA.n1028 GNDA.n952 53.3664
R2843 GNDA.n1035 GNDA.n950 53.3664
R2844 GNDA.n1969 GNDA.n1908 53.3664
R2845 GNDA.n1966 GNDA.n1898 53.3664
R2846 GNDA.n1962 GNDA.n1907 53.3664
R2847 GNDA.n1958 GNDA.n1900 53.3664
R2848 GNDA.n1947 GNDA.n1903 53.3664
R2849 GNDA.n1943 GNDA.n1904 53.3664
R2850 GNDA.n1939 GNDA.n1905 53.3664
R2851 GNDA.n1935 GNDA.n1906 53.3664
R2852 GNDA.n1995 GNDA.n1893 53.3664
R2853 GNDA.n1988 GNDA.n1987 53.3664
R2854 GNDA.n1920 GNDA.n1899 53.3664
R2855 GNDA.n1927 GNDA.n1901 53.3664
R2856 GNDA.n1986 GNDA.n1985 53.3664
R2857 GNDA.n1913 GNDA.n1911 53.3664
R2858 GNDA.n1980 GNDA.n1910 53.3664
R2859 GNDA.n1976 GNDA.n1909 53.3664
R2860 GNDA.n1986 GNDA.n1912 53.3664
R2861 GNDA.n1981 GNDA.n1911 53.3664
R2862 GNDA.n1977 GNDA.n1910 53.3664
R2863 GNDA.n1973 GNDA.n1909 53.3664
R2864 GNDA.n1955 GNDA.n1900 53.3664
R2865 GNDA.n1959 GNDA.n1907 53.3664
R2866 GNDA.n1963 GNDA.n1898 53.3664
R2867 GNDA.n1967 GNDA.n1908 53.3664
R2868 GNDA.n1938 GNDA.n1906 53.3664
R2869 GNDA.n1942 GNDA.n1905 53.3664
R2870 GNDA.n1946 GNDA.n1904 53.3664
R2871 GNDA.n1950 GNDA.n1903 53.3664
R2872 GNDA.n1934 GNDA.n1901 53.3664
R2873 GNDA.n1926 GNDA.n1899 53.3664
R2874 GNDA.n1987 GNDA.n1897 53.3664
R2875 GNDA.n1896 GNDA.n1893 53.3664
R2876 GNDA.n649 GNDA.n577 53.3664
R2877 GNDA.n648 GNDA.n647 53.3664
R2878 GNDA.n641 GNDA.n579 53.3664
R2879 GNDA.n640 GNDA.n639 53.3664
R2880 GNDA.n631 GNDA.n630 53.3664
R2881 GNDA.n626 GNDA.n585 53.3664
R2882 GNDA.n624 GNDA.n623 53.3664
R2883 GNDA.n619 GNDA.n587 53.3664
R2884 GNDA.n676 GNDA.n675 53.3664
R2885 GNDA.n602 GNDA.n572 53.3664
R2886 GNDA.n605 GNDA.n604 53.3664
R2887 GNDA.n617 GNDA.n616 53.3664
R2888 GNDA.n656 GNDA.n655 53.3664
R2889 GNDA.n658 GNDA.n657 53.3664
R2890 GNDA.n663 GNDA.n662 53.3664
R2891 GNDA.n666 GNDA.n665 53.3664
R2892 GNDA.n655 GNDA.n654 53.3664
R2893 GNDA.n657 GNDA.n575 53.3664
R2894 GNDA.n664 GNDA.n663 53.3664
R2895 GNDA.n665 GNDA.n573 53.3664
R2896 GNDA.n639 GNDA.n638 53.3664
R2897 GNDA.n642 GNDA.n641 53.3664
R2898 GNDA.n647 GNDA.n646 53.3664
R2899 GNDA.n650 GNDA.n649 53.3664
R2900 GNDA.n587 GNDA.n586 53.3664
R2901 GNDA.n625 GNDA.n624 53.3664
R2902 GNDA.n585 GNDA.n583 53.3664
R2903 GNDA.n632 GNDA.n631 53.3664
R2904 GNDA.n618 GNDA.n617 53.3664
R2905 GNDA.n604 GNDA.n590 53.3664
R2906 GNDA.n603 GNDA.n602 53.3664
R2907 GNDA.n677 GNDA.n676 53.3664
R2908 GNDA.n761 GNDA.n555 53.3664
R2909 GNDA.n760 GNDA.n759 53.3664
R2910 GNDA.n753 GNDA.n557 53.3664
R2911 GNDA.n752 GNDA.n751 53.3664
R2912 GNDA.n743 GNDA.n742 53.3664
R2913 GNDA.n738 GNDA.n563 53.3664
R2914 GNDA.n736 GNDA.n735 53.3664
R2915 GNDA.n731 GNDA.n692 53.3664
R2916 GNDA.n788 GNDA.n787 53.3664
R2917 GNDA.n714 GNDA.n550 53.3664
R2918 GNDA.n717 GNDA.n716 53.3664
R2919 GNDA.n729 GNDA.n728 53.3664
R2920 GNDA.n768 GNDA.n767 53.3664
R2921 GNDA.n770 GNDA.n769 53.3664
R2922 GNDA.n775 GNDA.n774 53.3664
R2923 GNDA.n778 GNDA.n777 53.3664
R2924 GNDA.n767 GNDA.n766 53.3664
R2925 GNDA.n769 GNDA.n553 53.3664
R2926 GNDA.n776 GNDA.n775 53.3664
R2927 GNDA.n777 GNDA.n551 53.3664
R2928 GNDA.n751 GNDA.n750 53.3664
R2929 GNDA.n754 GNDA.n753 53.3664
R2930 GNDA.n759 GNDA.n758 53.3664
R2931 GNDA.n762 GNDA.n761 53.3664
R2932 GNDA.n692 GNDA.n564 53.3664
R2933 GNDA.n737 GNDA.n736 53.3664
R2934 GNDA.n563 GNDA.n561 53.3664
R2935 GNDA.n744 GNDA.n743 53.3664
R2936 GNDA.n730 GNDA.n729 53.3664
R2937 GNDA.n716 GNDA.n694 53.3664
R2938 GNDA.n715 GNDA.n714 53.3664
R2939 GNDA.n789 GNDA.n788 53.3664
R2940 GNDA.n1588 GNDA.n1277 53.3664
R2941 GNDA.n1584 GNDA.n1266 53.3664
R2942 GNDA.n1580 GNDA.n1276 53.3664
R2943 GNDA.n1576 GNDA.n1269 53.3664
R2944 GNDA.n1565 GNDA.n1272 53.3664
R2945 GNDA.n1561 GNDA.n1273 53.3664
R2946 GNDA.n1557 GNDA.n1274 53.3664
R2947 GNDA.n1553 GNDA.n1275 53.3664
R2948 GNDA.n1608 GNDA.n1607 53.3664
R2949 GNDA.n1530 GNDA.n1267 53.3664
R2950 GNDA.n1538 GNDA.n1268 53.3664
R2951 GNDA.n1545 GNDA.n1270 53.3664
R2952 GNDA.n1592 GNDA.n1281 53.3664
R2953 GNDA.n1593 GNDA.n1280 53.3664
R2954 GNDA.n1597 GNDA.n1279 53.3664
R2955 GNDA.n1601 GNDA.n1278 53.3664
R2956 GNDA.n1589 GNDA.n1281 53.3664
R2957 GNDA.n1596 GNDA.n1280 53.3664
R2958 GNDA.n1600 GNDA.n1279 53.3664
R2959 GNDA.n1604 GNDA.n1278 53.3664
R2960 GNDA.n1573 GNDA.n1269 53.3664
R2961 GNDA.n1577 GNDA.n1276 53.3664
R2962 GNDA.n1581 GNDA.n1266 53.3664
R2963 GNDA.n1585 GNDA.n1277 53.3664
R2964 GNDA.n1556 GNDA.n1275 53.3664
R2965 GNDA.n1560 GNDA.n1274 53.3664
R2966 GNDA.n1564 GNDA.n1273 53.3664
R2967 GNDA.n1568 GNDA.n1272 53.3664
R2968 GNDA.n1552 GNDA.n1270 53.3664
R2969 GNDA.n1544 GNDA.n1268 53.3664
R2970 GNDA.n1537 GNDA.n1267 53.3664
R2971 GNDA.n1607 GNDA.n1265 53.3664
R2972 GNDA.t182 GNDA.n180 52.0962
R2973 GNDA.t182 GNDA.n2182 52.0962
R2974 GNDA.t275 GNDA.n2227 52.0962
R2975 GNDA.t140 GNDA.t7 51.9061
R2976 GNDA.t295 GNDA.t328 51.9061
R2977 GNDA.t146 GNDA.t64 51.9061
R2978 GNDA.n2278 GNDA.t225 51.9061
R2979 GNDA.t149 GNDA.n681 50.0123
R2980 GNDA.n545 GNDA.n236 48.9704
R2981 GNDA.t182 GNDA.n405 48.9704
R2982 GNDA.t14 GNDA.n88 48.9704
R2983 GNDA.n1499 GNDA.n1291 48.2167
R2984 GNDA.n1500 GNDA.n1499 48.2167
R2985 GNDA.n1502 GNDA.n1500 48.2167
R2986 GNDA.n1502 GNDA.n1501 48.2167
R2987 GNDA.n1501 GNDA.n412 48.2167
R2988 GNDA.n1509 GNDA.n411 48.2167
R2989 GNDA.n1509 GNDA.n1285 48.2167
R2990 GNDA.n1516 GNDA.n1285 48.2167
R2991 GNDA.n1517 GNDA.n1516 48.2167
R2992 GNDA.n1518 GNDA.n1517 48.2167
R2993 GNDA.n1518 GNDA.n1283 48.2167
R2994 GNDA.n1283 GNDA.t55 48.2167
R2995 GNDA.n1116 GNDA.n1089 48.2167
R2996 GNDA.n1117 GNDA.n1116 48.2167
R2997 GNDA.n1119 GNDA.n1117 48.2167
R2998 GNDA.n1119 GNDA.n1118 48.2167
R2999 GNDA.n1118 GNDA.n409 48.2167
R3000 GNDA.n1126 GNDA.n408 48.2167
R3001 GNDA.n1126 GNDA.n1083 48.2167
R3002 GNDA.n1133 GNDA.n1083 48.2167
R3003 GNDA.n1134 GNDA.n1133 48.2167
R3004 GNDA.n1135 GNDA.n1134 48.2167
R3005 GNDA.n1135 GNDA.n406 48.2167
R3006 GNDA.n2048 GNDA.n2047 48.2167
R3007 GNDA.n2047 GNDA.n2046 48.2167
R3008 GNDA.n2046 GNDA.n2037 48.2167
R3009 GNDA.n2040 GNDA.n2037 48.2167
R3010 GNDA.n2040 GNDA.n59 48.2167
R3011 GNDA.n2256 GNDA.n55 48.2167
R3012 GNDA.n2262 GNDA.n55 48.2167
R3013 GNDA.n2263 GNDA.n2262 48.2167
R3014 GNDA.n2266 GNDA.n2263 48.2167
R3015 GNDA.n2266 GNDA.n2265 48.2167
R3016 GNDA.n2265 GNDA.n2264 48.2167
R3017 GNDA.n374 GNDA.t279 48.0005
R3018 GNDA.n374 GNDA.t102 48.0005
R3019 GNDA.n371 GNDA.t139 48.0005
R3020 GNDA.n371 GNDA.t169 48.0005
R3021 GNDA.n367 GNDA.t128 48.0005
R3022 GNDA.n367 GNDA.t108 48.0005
R3023 GNDA.n364 GNDA.t104 48.0005
R3024 GNDA.n364 GNDA.t16 48.0005
R3025 GNDA.n360 GNDA.t51 48.0005
R3026 GNDA.n360 GNDA.t106 48.0005
R3027 GNDA.n2155 GNDA.t26 47.9285
R3028 GNDA.n318 GNDA.n317 47.9134
R3029 GNDA.n333 GNDA.n332 47.9134
R3030 GNDA.t167 GNDA.t176 47.9134
R3031 GNDA.t84 GNDA.t52 47.9134
R3032 GNDA.t86 GNDA.t118 47.9134
R3033 GNDA.t329 GNDA.t32 47.9134
R3034 GNDA.t5 GNDA.t70 47.9134
R3035 GNDA.t31 GNDA.t109 47.9134
R3036 GNDA.t173 GNDA.t153 47.9134
R3037 GNDA.t120 GNDA.t246 47.9134
R3038 GNDA.t111 GNDA.t72 47.9134
R3039 GNDA.t155 GNDA.t37 47.9134
R3040 GNDA.t66 GNDA.t157 47.9134
R3041 GNDA.t34 GNDA.t165 47.9134
R3042 GNDA.t272 GNDA.t17 47.9134
R3043 GNDA.t68 GNDA.t13 47.9134
R3044 GNDA.t215 GNDA.t12 47.9134
R3045 GNDA.t182 GNDA.n2036 47.6748
R3046 GNDA.t27 GNDA.t280 46.8866
R3047 GNDA.n1380 GNDA.t182 46.2335
R3048 GNDA.t182 GNDA.n1311 46.2335
R3049 GNDA.t182 GNDA.n1483 46.2335
R3050 GNDA.n593 GNDA.t182 44.8028
R3051 GNDA.n381 GNDA.t6 43.9206
R3052 GNDA.n381 GNDA.t85 43.9206
R3053 GNDA.t284 GNDA.t298 43.9206
R3054 GNDA.t314 GNDA.t284 43.9206
R3055 GNDA.n546 GNDA.t76 43.7609
R3056 GNDA.n682 GNDA.t149 43.7609
R3057 GNDA.n597 GNDA.t288 42.7189
R3058 GNDA.t100 GNDA.t163 42.4101
R3059 GNDA.t43 GNDA.t100 42.4101
R3060 GNDA.t319 GNDA.t135 42.4101
R3061 GNDA.t337 GNDA.t319 42.4101
R3062 GNDA.t182 GNDA.n1366 42.2987
R3063 GNDA.n1412 GNDA.t182 42.2987
R3064 GNDA.n1484 GNDA.t182 42.2987
R3065 GNDA.t182 GNDA.t26 41.677
R3066 GNDA.t182 GNDA.t14 41.677
R3067 GNDA.n2200 GNDA.t59 41.0662
R3068 GNDA.n2202 GNDA.t39 40.4338
R3069 GNDA.n258 GNDA.t217 40.4338
R3070 GNDA.n285 GNDA.t177 40.4338
R3071 GNDA.n399 GNDA.n240 40.1221
R3072 GNDA.t176 GNDA.t38 39.9279
R3073 GNDA.t52 GNDA.t167 39.9279
R3074 GNDA.t118 GNDA.t84 39.9279
R3075 GNDA.t32 GNDA.t86 39.9279
R3076 GNDA.t70 GNDA.t329 39.9279
R3077 GNDA.t109 GNDA.t5 39.9279
R3078 GNDA.t153 GNDA.t31 39.9279
R3079 GNDA.t64 GNDA.t173 39.9279
R3080 GNDA.t13 GNDA.t272 39.9279
R3081 GNDA.t12 GNDA.t68 39.9279
R3082 GNDA.t114 GNDA.t215 39.9279
R3083 GNDA.n2293 GNDA.n2292 39.9279
R3084 GNDA.t209 GNDA.n698 39.5932
R3085 GNDA.n612 GNDA.t87 39.5932
R3086 GNDA.t334 GNDA.n2255 39.5932
R3087 GNDA.n685 GNDA.n180 38.5513
R3088 GNDA.n2197 GNDA.n97 38.5513
R3089 GNDA.n2244 GNDA.t126 38.5513
R3090 GNDA.n2255 GNDA.t11 38.5513
R3091 GNDA.n108 GNDA.t171 38.5513
R3092 GNDA.t325 GNDA.t320 38.533
R3093 GNDA.n262 GNDA.n261 37.5297
R3094 GNDA.n264 GNDA.n263 37.5297
R3095 GNDA.n266 GNDA.n265 37.5297
R3096 GNDA.n268 GNDA.n267 37.5297
R3097 GNDA.n270 GNDA.n269 37.5297
R3098 GNDA.n272 GNDA.n271 37.5297
R3099 GNDA.n274 GNDA.n273 37.5297
R3100 GNDA.n276 GNDA.n275 37.5297
R3101 GNDA.n278 GNDA.n277 37.5297
R3102 GNDA.n280 GNDA.n279 37.5297
R3103 GNDA.n282 GNDA.n281 37.5297
R3104 GNDA.n2182 GNDA.n183 37.5094
R3105 GNDA.t315 GNDA.t11 36.4675
R3106 GNDA.t7 GNDA.t117 35.9352
R3107 GNDA.t10 GNDA.t295 35.9352
R3108 GNDA.n256 GNDA.t34 35.9352
R3109 GNDA.n795 GNDA.t292 34.3836
R3110 GNDA.t289 GNDA.n405 34.3836
R3111 GNDA.n724 GNDA.t27 34.3836
R3112 GNDA.n683 GNDA.n96 34.3836
R3113 GNDA.t122 GNDA.n610 33.3417
R3114 GNDA.n2242 GNDA.t312 33.3417
R3115 GNDA.t182 GNDA.n410 32.9056
R3116 GNDA.t182 GNDA.n407 32.9056
R3117 GNDA.t182 GNDA.n412 32.6804
R3118 GNDA.t182 GNDA.n409 32.6804
R3119 GNDA.t182 GNDA.n59 32.6804
R3120 GNDA.n702 GNDA.n701 31.4662
R3121 GNDA.t171 GNDA.n47 31.2579
R3122 GNDA.n41 GNDA.n40 31.1567
R3123 GNDA.n316 GNDA.t188 31.1255
R3124 GNDA.n334 GNDA.t200 31.1255
R3125 GNDA.n2276 GNDA.t226 31.1255
R3126 GNDA.n2294 GNDA.t213 31.1255
R3127 GNDA.n313 GNDA.n312 31.1255
R3128 GNDA.n704 GNDA.n703 30.8338
R3129 GNDA.n2311 GNDA.n0 30.4627
R3130 GNDA.n352 GNDA.n351 29.8672
R3131 GNDA.n340 GNDA.n339 29.8672
R3132 GNDA.n2300 GNDA.n4 29.8672
R3133 GNDA.n596 GNDA.t41 29.1741
R3134 GNDA.n2229 GNDA.t184 29.1741
R3135 GNDA.t148 GNDA.n722 28.1322
R3136 GNDA.n698 GNDA.t291 28.1322
R3137 GNDA.t308 GNDA.t321 27.9497
R3138 GNDA.t93 GNDA.t294 27.9497
R3139 GNDA.n152 GNDA.n149 27.5561
R3140 GNDA.n1207 GNDA.n1204 27.5561
R3141 GNDA.n1787 GNDA.n1784 27.5561
R3142 GNDA.n1688 GNDA.n1685 27.5561
R3143 GNDA.n1004 GNDA.n1001 27.5561
R3144 GNDA.n1971 GNDA.n1970 27.5561
R3145 GNDA.n653 GNDA.n652 27.5561
R3146 GNDA.n765 GNDA.n764 27.5561
R3147 GNDA.n1590 GNDA.n1587 27.5561
R3148 GNDA.n133 GNDA.n132 26.6672
R3149 GNDA.n1188 GNDA.n1187 26.6672
R3150 GNDA.n1768 GNDA.n1767 26.6672
R3151 GNDA.n1669 GNDA.n1668 26.6672
R3152 GNDA.n985 GNDA.n984 26.6672
R3153 GNDA.n1953 GNDA.n1952 26.6672
R3154 GNDA.n636 GNDA.n635 26.6672
R3155 GNDA.n748 GNDA.n747 26.6672
R3156 GNDA.n1571 GNDA.n1570 26.6672
R3157 GNDA.t299 GNDA.t21 26.0483
R3158 GNDA.n2273 GNDA.n2272 25.0064
R3159 GNDA.n187 GNDA.t281 24.0005
R3160 GNDA.n187 GNDA.t300 24.0005
R3161 GNDA.n536 GNDA.t162 24.0005
R3162 GNDA.n536 GNDA.t160 24.0005
R3163 GNDA.n539 GNDA.t90 24.0005
R3164 GNDA.n539 GNDA.t77 24.0005
R3165 GNDA.n2176 GNDA.t88 24.0005
R3166 GNDA.n2176 GNDA.t331 24.0005
R3167 GNDA.n2172 GNDA.t269 24.0005
R3168 GNDA.n2172 GNDA.t123 24.0005
R3169 GNDA.n2169 GNDA.t42 24.0005
R3170 GNDA.n2169 GNDA.t340 24.0005
R3171 GNDA.n2165 GNDA.t29 24.0005
R3172 GNDA.n2165 GNDA.t150 24.0005
R3173 GNDA.n2213 GNDA.t316 24.0005
R3174 GNDA.n2213 GNDA.t152 24.0005
R3175 GNDA.n2217 GNDA.t313 24.0005
R3176 GNDA.n2217 GNDA.t335 24.0005
R3177 GNDA.n2220 GNDA.t125 24.0005
R3178 GNDA.n2220 GNDA.t142 24.0005
R3179 GNDA.n2227 GNDA.n88 23.9645
R3180 GNDA.n2228 GNDA.t275 23.9645
R3181 GNDA.t144 GNDA.n2242 23.9645
R3182 GNDA.n107 GNDA.t143 23.9645
R3183 GNDA.n2272 GNDA.n47 23.9645
R3184 GNDA.t246 GNDA.t132 23.9569
R3185 GNDA.t72 GNDA.t336 23.9569
R3186 GNDA.t37 GNDA.t18 23.9569
R3187 GNDA.t157 GNDA.t333 23.9569
R3188 GNDA.t165 GNDA.t232 23.9569
R3189 GNDA.t130 GNDA.t325 23.9532
R3190 GNDA.n793 GNDA.t89 22.9226
R3191 GNDA.n683 GNDA.t28 22.9226
R3192 GNDA.n385 GNDA.n384 21.7827
R3193 GNDA.n242 GNDA.n43 21.7827
R3194 GNDA.n2311 GNDA.n2310 21.383
R3195 GNDA.n1316 GNDA.n1315 21.0192
R3196 GNDA.t182 GNDA.n236 20.8388
R3197 GNDA.t293 GNDA.n706 20.8388
R3198 GNDA.t4 GNDA.n61 20.8388
R3199 GNDA.t182 GNDA.n61 20.8388
R3200 GNDA.t182 GNDA.n404 20.0574
R3201 GNDA.t286 GNDA.t2 19.9642
R3202 GNDA.t283 GNDA.t95 19.9642
R3203 GNDA.n286 GNDA.t40 19.9642
R3204 GNDA.n348 GNDA.t46 19.9642
R3205 GNDA.n257 GNDA.t113 19.9642
R3206 GNDA.n22 GNDA.t170 19.7005
R3207 GNDA.n22 GNDA.t302 19.7005
R3208 GNDA.n25 GNDA.t310 19.7005
R3209 GNDA.n25 GNDA.t318 19.7005
R3210 GNDA.n28 GNDA.t303 19.7005
R3211 GNDA.n28 GNDA.t307 19.7005
R3212 GNDA.n32 GNDA.t301 19.7005
R3213 GNDA.n32 GNDA.t309 19.7005
R3214 GNDA.n35 GNDA.t297 19.7005
R3215 GNDA.n35 GNDA.t83 19.7005
R3216 GNDA.n38 GNDA.t306 19.7005
R3217 GNDA.n38 GNDA.t145 19.7005
R3218 GNDA.n294 GNDA.t56 19.7005
R3219 GNDA.n294 GNDA.t62 19.7005
R3220 GNDA.n297 GNDA.t30 19.7005
R3221 GNDA.n297 GNDA.t74 19.7005
R3222 GNDA.n300 GNDA.t158 19.7005
R3223 GNDA.n300 GNDA.t73 19.7005
R3224 GNDA.n304 GNDA.t282 19.7005
R3225 GNDA.n304 GNDA.t115 19.7005
R3226 GNDA.n307 GNDA.t323 19.7005
R3227 GNDA.n307 GNDA.t75 19.7005
R3228 GNDA.n310 GNDA.t63 19.7005
R3229 GNDA.n310 GNDA.t116 19.7005
R3230 GNDA.t182 GNDA.n413 19.6741
R3231 GNDA.t330 GNDA.n97 18.7549
R3232 GNDA.n106 GNDA.t315 18.7549
R3233 GNDA.n1410 GNDA.n1409 18.5605
R3234 GNDA GNDA.n94 18.1604
R3235 GNDA.n2051 GNDA.n229 17.5843
R3236 GNDA.n1113 GNDA.n1112 17.5843
R3237 GNDA.n1496 GNDA.n1495 17.5843
R3238 GNDA.n351 GNDA.n350 17.5172
R3239 GNDA.n2303 GNDA.n4 17.4755
R3240 GNDA.n1836 GNDA.n825 16.9379
R3241 GNDA.n1865 GNDA.n1864 16.9379
R3242 GNDA.n819 GNDA.n529 16.9379
R3243 GNDA.n2007 GNDA.n209 16.7709
R3244 GNDA.n2032 GNDA.n439 16.7709
R3245 GNDA.n1618 GNDA.n1259 16.7709
R3246 GNDA.n1059 GNDA.n218 16.7709
R3247 GNDA.n2207 GNDA.n2206 16.0112
R3248 GNDA.n153 GNDA.n152 16.0005
R3249 GNDA.n156 GNDA.n153 16.0005
R3250 GNDA.n157 GNDA.n156 16.0005
R3251 GNDA.n160 GNDA.n157 16.0005
R3252 GNDA.n161 GNDA.n160 16.0005
R3253 GNDA.n164 GNDA.n161 16.0005
R3254 GNDA.n166 GNDA.n164 16.0005
R3255 GNDA.n167 GNDA.n166 16.0005
R3256 GNDA.n149 GNDA.n148 16.0005
R3257 GNDA.n148 GNDA.n145 16.0005
R3258 GNDA.n145 GNDA.n144 16.0005
R3259 GNDA.n144 GNDA.n141 16.0005
R3260 GNDA.n141 GNDA.n140 16.0005
R3261 GNDA.n140 GNDA.n137 16.0005
R3262 GNDA.n137 GNDA.n136 16.0005
R3263 GNDA.n136 GNDA.n133 16.0005
R3264 GNDA.n132 GNDA.n129 16.0005
R3265 GNDA.n129 GNDA.n128 16.0005
R3266 GNDA.n128 GNDA.n125 16.0005
R3267 GNDA.n125 GNDA.n124 16.0005
R3268 GNDA.n124 GNDA.n121 16.0005
R3269 GNDA.n121 GNDA.n120 16.0005
R3270 GNDA.n120 GNDA.n117 16.0005
R3271 GNDA.n117 GNDA.n116 16.0005
R3272 GNDA.n1208 GNDA.n1207 16.0005
R3273 GNDA.n1211 GNDA.n1208 16.0005
R3274 GNDA.n1212 GNDA.n1211 16.0005
R3275 GNDA.n1215 GNDA.n1212 16.0005
R3276 GNDA.n1216 GNDA.n1215 16.0005
R3277 GNDA.n1219 GNDA.n1216 16.0005
R3278 GNDA.n1220 GNDA.n1219 16.0005
R3279 GNDA.n1220 GNDA.n1060 16.0005
R3280 GNDA.n1204 GNDA.n1203 16.0005
R3281 GNDA.n1203 GNDA.n1200 16.0005
R3282 GNDA.n1200 GNDA.n1199 16.0005
R3283 GNDA.n1199 GNDA.n1196 16.0005
R3284 GNDA.n1196 GNDA.n1195 16.0005
R3285 GNDA.n1195 GNDA.n1192 16.0005
R3286 GNDA.n1192 GNDA.n1191 16.0005
R3287 GNDA.n1191 GNDA.n1188 16.0005
R3288 GNDA.n1187 GNDA.n1184 16.0005
R3289 GNDA.n1184 GNDA.n1183 16.0005
R3290 GNDA.n1183 GNDA.n1180 16.0005
R3291 GNDA.n1180 GNDA.n1179 16.0005
R3292 GNDA.n1179 GNDA.n1176 16.0005
R3293 GNDA.n1176 GNDA.n1175 16.0005
R3294 GNDA.n1175 GNDA.n1172 16.0005
R3295 GNDA.n1172 GNDA.n1171 16.0005
R3296 GNDA.n1317 GNDA.n1316 16.0005
R3297 GNDA.n1410 GNDA.n1317 16.0005
R3298 GNDA.n1788 GNDA.n1787 16.0005
R3299 GNDA.n1791 GNDA.n1788 16.0005
R3300 GNDA.n1792 GNDA.n1791 16.0005
R3301 GNDA.n1795 GNDA.n1792 16.0005
R3302 GNDA.n1796 GNDA.n1795 16.0005
R3303 GNDA.n1799 GNDA.n1796 16.0005
R3304 GNDA.n1800 GNDA.n1799 16.0005
R3305 GNDA.n1803 GNDA.n1800 16.0005
R3306 GNDA.n1784 GNDA.n1783 16.0005
R3307 GNDA.n1783 GNDA.n1780 16.0005
R3308 GNDA.n1780 GNDA.n1779 16.0005
R3309 GNDA.n1779 GNDA.n1776 16.0005
R3310 GNDA.n1776 GNDA.n1775 16.0005
R3311 GNDA.n1775 GNDA.n1772 16.0005
R3312 GNDA.n1772 GNDA.n1771 16.0005
R3313 GNDA.n1771 GNDA.n1768 16.0005
R3314 GNDA.n1767 GNDA.n1764 16.0005
R3315 GNDA.n1764 GNDA.n1763 16.0005
R3316 GNDA.n1763 GNDA.n1760 16.0005
R3317 GNDA.n1760 GNDA.n1759 16.0005
R3318 GNDA.n1759 GNDA.n1756 16.0005
R3319 GNDA.n1756 GNDA.n1755 16.0005
R3320 GNDA.n1755 GNDA.n1752 16.0005
R3321 GNDA.n1752 GNDA.n1751 16.0005
R3322 GNDA.n1689 GNDA.n1688 16.0005
R3323 GNDA.n1692 GNDA.n1689 16.0005
R3324 GNDA.n1693 GNDA.n1692 16.0005
R3325 GNDA.n1696 GNDA.n1693 16.0005
R3326 GNDA.n1697 GNDA.n1696 16.0005
R3327 GNDA.n1700 GNDA.n1697 16.0005
R3328 GNDA.n1701 GNDA.n1700 16.0005
R3329 GNDA.n1701 GNDA.n871 16.0005
R3330 GNDA.n1685 GNDA.n1684 16.0005
R3331 GNDA.n1684 GNDA.n1681 16.0005
R3332 GNDA.n1681 GNDA.n1680 16.0005
R3333 GNDA.n1680 GNDA.n1677 16.0005
R3334 GNDA.n1677 GNDA.n1676 16.0005
R3335 GNDA.n1676 GNDA.n1673 16.0005
R3336 GNDA.n1673 GNDA.n1672 16.0005
R3337 GNDA.n1672 GNDA.n1669 16.0005
R3338 GNDA.n1668 GNDA.n1665 16.0005
R3339 GNDA.n1665 GNDA.n1664 16.0005
R3340 GNDA.n1664 GNDA.n1661 16.0005
R3341 GNDA.n1661 GNDA.n1660 16.0005
R3342 GNDA.n1660 GNDA.n1657 16.0005
R3343 GNDA.n1657 GNDA.n1656 16.0005
R3344 GNDA.n1656 GNDA.n1653 16.0005
R3345 GNDA.n1653 GNDA.n1652 16.0005
R3346 GNDA.n1005 GNDA.n1004 16.0005
R3347 GNDA.n1008 GNDA.n1005 16.0005
R3348 GNDA.n1009 GNDA.n1008 16.0005
R3349 GNDA.n1012 GNDA.n1009 16.0005
R3350 GNDA.n1013 GNDA.n1012 16.0005
R3351 GNDA.n1016 GNDA.n1013 16.0005
R3352 GNDA.n1018 GNDA.n1016 16.0005
R3353 GNDA.n1019 GNDA.n1018 16.0005
R3354 GNDA.n1001 GNDA.n1000 16.0005
R3355 GNDA.n1000 GNDA.n997 16.0005
R3356 GNDA.n997 GNDA.n996 16.0005
R3357 GNDA.n996 GNDA.n993 16.0005
R3358 GNDA.n993 GNDA.n992 16.0005
R3359 GNDA.n992 GNDA.n989 16.0005
R3360 GNDA.n989 GNDA.n988 16.0005
R3361 GNDA.n988 GNDA.n985 16.0005
R3362 GNDA.n984 GNDA.n981 16.0005
R3363 GNDA.n981 GNDA.n980 16.0005
R3364 GNDA.n980 GNDA.n977 16.0005
R3365 GNDA.n977 GNDA.n976 16.0005
R3366 GNDA.n976 GNDA.n973 16.0005
R3367 GNDA.n973 GNDA.n972 16.0005
R3368 GNDA.n972 GNDA.n969 16.0005
R3369 GNDA.n969 GNDA.n945 16.0005
R3370 GNDA.n1984 GNDA.n1971 16.0005
R3371 GNDA.n1984 GNDA.n1983 16.0005
R3372 GNDA.n1983 GNDA.n1982 16.0005
R3373 GNDA.n1982 GNDA.n1979 16.0005
R3374 GNDA.n1979 GNDA.n1978 16.0005
R3375 GNDA.n1978 GNDA.n1975 16.0005
R3376 GNDA.n1975 GNDA.n1974 16.0005
R3377 GNDA.n1974 GNDA.n1889 16.0005
R3378 GNDA.n1970 GNDA.n1968 16.0005
R3379 GNDA.n1968 GNDA.n1965 16.0005
R3380 GNDA.n1965 GNDA.n1964 16.0005
R3381 GNDA.n1964 GNDA.n1961 16.0005
R3382 GNDA.n1961 GNDA.n1960 16.0005
R3383 GNDA.n1960 GNDA.n1957 16.0005
R3384 GNDA.n1957 GNDA.n1956 16.0005
R3385 GNDA.n1956 GNDA.n1953 16.0005
R3386 GNDA.n1952 GNDA.n1949 16.0005
R3387 GNDA.n1949 GNDA.n1948 16.0005
R3388 GNDA.n1948 GNDA.n1945 16.0005
R3389 GNDA.n1945 GNDA.n1944 16.0005
R3390 GNDA.n1944 GNDA.n1941 16.0005
R3391 GNDA.n1941 GNDA.n1940 16.0005
R3392 GNDA.n1940 GNDA.n1937 16.0005
R3393 GNDA.n1937 GNDA.n1936 16.0005
R3394 GNDA.n653 GNDA.n576 16.0005
R3395 GNDA.n659 GNDA.n576 16.0005
R3396 GNDA.n660 GNDA.n659 16.0005
R3397 GNDA.n661 GNDA.n660 16.0005
R3398 GNDA.n661 GNDA.n574 16.0005
R3399 GNDA.n667 GNDA.n574 16.0005
R3400 GNDA.n668 GNDA.n667 16.0005
R3401 GNDA.n669 GNDA.n668 16.0005
R3402 GNDA.n652 GNDA.n651 16.0005
R3403 GNDA.n651 GNDA.n578 16.0005
R3404 GNDA.n645 GNDA.n578 16.0005
R3405 GNDA.n645 GNDA.n644 16.0005
R3406 GNDA.n644 GNDA.n643 16.0005
R3407 GNDA.n643 GNDA.n580 16.0005
R3408 GNDA.n637 GNDA.n580 16.0005
R3409 GNDA.n637 GNDA.n636 16.0005
R3410 GNDA.n635 GNDA.n582 16.0005
R3411 GNDA.n629 GNDA.n582 16.0005
R3412 GNDA.n629 GNDA.n628 16.0005
R3413 GNDA.n628 GNDA.n627 16.0005
R3414 GNDA.n627 GNDA.n584 16.0005
R3415 GNDA.n622 GNDA.n584 16.0005
R3416 GNDA.n622 GNDA.n621 16.0005
R3417 GNDA.n621 GNDA.n620 16.0005
R3418 GNDA.n765 GNDA.n554 16.0005
R3419 GNDA.n771 GNDA.n554 16.0005
R3420 GNDA.n772 GNDA.n771 16.0005
R3421 GNDA.n773 GNDA.n772 16.0005
R3422 GNDA.n773 GNDA.n552 16.0005
R3423 GNDA.n779 GNDA.n552 16.0005
R3424 GNDA.n780 GNDA.n779 16.0005
R3425 GNDA.n781 GNDA.n780 16.0005
R3426 GNDA.n764 GNDA.n763 16.0005
R3427 GNDA.n763 GNDA.n556 16.0005
R3428 GNDA.n757 GNDA.n556 16.0005
R3429 GNDA.n757 GNDA.n756 16.0005
R3430 GNDA.n756 GNDA.n755 16.0005
R3431 GNDA.n755 GNDA.n558 16.0005
R3432 GNDA.n749 GNDA.n558 16.0005
R3433 GNDA.n749 GNDA.n748 16.0005
R3434 GNDA.n747 GNDA.n560 16.0005
R3435 GNDA.n741 GNDA.n560 16.0005
R3436 GNDA.n741 GNDA.n740 16.0005
R3437 GNDA.n740 GNDA.n739 16.0005
R3438 GNDA.n739 GNDA.n562 16.0005
R3439 GNDA.n734 GNDA.n562 16.0005
R3440 GNDA.n734 GNDA.n733 16.0005
R3441 GNDA.n733 GNDA.n732 16.0005
R3442 GNDA.n1591 GNDA.n1590 16.0005
R3443 GNDA.n1594 GNDA.n1591 16.0005
R3444 GNDA.n1595 GNDA.n1594 16.0005
R3445 GNDA.n1598 GNDA.n1595 16.0005
R3446 GNDA.n1599 GNDA.n1598 16.0005
R3447 GNDA.n1602 GNDA.n1599 16.0005
R3448 GNDA.n1603 GNDA.n1602 16.0005
R3449 GNDA.n1603 GNDA.n1261 16.0005
R3450 GNDA.n1587 GNDA.n1586 16.0005
R3451 GNDA.n1586 GNDA.n1583 16.0005
R3452 GNDA.n1583 GNDA.n1582 16.0005
R3453 GNDA.n1582 GNDA.n1579 16.0005
R3454 GNDA.n1579 GNDA.n1578 16.0005
R3455 GNDA.n1578 GNDA.n1575 16.0005
R3456 GNDA.n1575 GNDA.n1574 16.0005
R3457 GNDA.n1574 GNDA.n1571 16.0005
R3458 GNDA.n1570 GNDA.n1567 16.0005
R3459 GNDA.n1567 GNDA.n1566 16.0005
R3460 GNDA.n1566 GNDA.n1563 16.0005
R3461 GNDA.n1563 GNDA.n1562 16.0005
R3462 GNDA.n1562 GNDA.n1559 16.0005
R3463 GNDA.n1559 GNDA.n1558 16.0005
R3464 GNDA.n1558 GNDA.n1555 16.0005
R3465 GNDA.n1555 GNDA.n1554 16.0005
R3466 GNDA.n348 GNDA.t146 15.9715
R3467 GNDA.t80 GNDA.t179 15.9715
R3468 GNDA.t132 GNDA.t98 15.9715
R3469 GNDA.t336 GNDA.t120 15.9715
R3470 GNDA.t18 GNDA.t111 15.9715
R3471 GNDA.t333 GNDA.t155 15.9715
R3472 GNDA.t232 GNDA.t66 15.9715
R3473 GNDA.t76 GNDA.t289 15.6292
R3474 GNDA.t182 GNDA.t161 15.6292
R3475 GNDA.t1 GNDA.t264 15.6292
R3476 GNDA.t182 GNDA.n411 15.5368
R3477 GNDA.t182 GNDA.n408 15.5368
R3478 GNDA.n2256 GNDA.t182 15.5368
R3479 GNDA.n335 GNDA.n290 15.1255
R3480 GNDA.n2295 GNDA.n8 15.1255
R3481 GNDA.n345 GNDA.n288 14.6634
R3482 GNDA.n15 GNDA.n13 14.6634
R3483 GNDA.n1812 GNDA.n410 14.555
R3484 GNDA.n2003 GNDA.n407 14.555
R3485 GNDA.n353 GNDA.n352 14.0922
R3486 GNDA.n2301 GNDA.n2300 14.0922
R3487 GNDA.n2205 GNDA.n2204 12.7542
R3488 GNDA.n2279 GNDA.t244 12.6791
R3489 GNDA.n2291 GNDA.t255 12.6791
R3490 GNDA.n319 GNDA.t206 12.6791
R3491 GNDA.n331 GNDA.t197 12.6791
R3492 GNDA.t280 GNDA.n723 12.5035
R3493 GNDA.n593 GNDA.t268 12.5035
R3494 GNDA.n2243 GNDA.t141 12.5035
R3495 GNDA.n359 GNDA.n354 12.2817
R3496 GNDA.n2199 GNDA.n2198 12.2193
R3497 GNDA.t305 GNDA.t254 11.9787
R3498 GNDA.t23 GNDA.t82 11.9787
R3499 GNDA.n2039 GNDA.n229 11.6369
R3500 GNDA.n2044 GNDA.n2039 11.6369
R3501 GNDA.n2044 GNDA.n2043 11.6369
R3502 GNDA.n2043 GNDA.n2042 11.6369
R3503 GNDA.n2042 GNDA.n57 11.6369
R3504 GNDA.n2258 GNDA.n57 11.6369
R3505 GNDA.n2259 GNDA.n2258 11.6369
R3506 GNDA.n2260 GNDA.n2259 11.6369
R3507 GNDA.n2260 GNDA.n52 11.6369
R3508 GNDA.n2268 GNDA.n52 11.6369
R3509 GNDA.n2067 GNDA.n221 11.6369
R3510 GNDA.n2067 GNDA.n2066 11.6369
R3511 GNDA.n2066 GNDA.n2065 11.6369
R3512 GNDA.n2065 GNDA.n223 11.6369
R3513 GNDA.n2060 GNDA.n223 11.6369
R3514 GNDA.n2060 GNDA.n2059 11.6369
R3515 GNDA.n2059 GNDA.n2058 11.6369
R3516 GNDA.n2058 GNDA.n226 11.6369
R3517 GNDA.n2053 GNDA.n226 11.6369
R3518 GNDA.n2053 GNDA.n2052 11.6369
R3519 GNDA.n2052 GNDA.n2051 11.6369
R3520 GNDA.n1114 GNDA.n1113 11.6369
R3521 GNDA.n1114 GNDA.n1087 11.6369
R3522 GNDA.n1121 GNDA.n1087 11.6369
R3523 GNDA.n1122 GNDA.n1121 11.6369
R3524 GNDA.n1123 GNDA.n1122 11.6369
R3525 GNDA.n1123 GNDA.n1085 11.6369
R3526 GNDA.n1128 GNDA.n1085 11.6369
R3527 GNDA.n1129 GNDA.n1128 11.6369
R3528 GNDA.n1131 GNDA.n1129 11.6369
R3529 GNDA.n1131 GNDA.n1130 11.6369
R3530 GNDA.n1091 GNDA.n894 11.6369
R3531 GNDA.n1094 GNDA.n1091 11.6369
R3532 GNDA.n1095 GNDA.n1094 11.6369
R3533 GNDA.n1098 GNDA.n1095 11.6369
R3534 GNDA.n1099 GNDA.n1098 11.6369
R3535 GNDA.n1102 GNDA.n1099 11.6369
R3536 GNDA.n1103 GNDA.n1102 11.6369
R3537 GNDA.n1106 GNDA.n1103 11.6369
R3538 GNDA.n1107 GNDA.n1106 11.6369
R3539 GNDA.n1110 GNDA.n1107 11.6369
R3540 GNDA.n1112 GNDA.n1110 11.6369
R3541 GNDA.n1374 GNDA.n825 11.6369
R3542 GNDA.n1375 GNDA.n1374 11.6369
R3543 GNDA.n1376 GNDA.n1375 11.6369
R3544 GNDA.n1376 GNDA.n1368 11.6369
R3545 GNDA.n1382 GNDA.n1368 11.6369
R3546 GNDA.n1383 GNDA.n1382 11.6369
R3547 GNDA.n1384 GNDA.n1383 11.6369
R3548 GNDA.n1384 GNDA.n1364 11.6369
R3549 GNDA.n1390 GNDA.n1364 11.6369
R3550 GNDA.n1391 GNDA.n1390 11.6369
R3551 GNDA.n1392 GNDA.n1391 11.6369
R3552 GNDA.n1836 GNDA.n1835 11.6369
R3553 GNDA.n1835 GNDA.n1834 11.6369
R3554 GNDA.n1834 GNDA.n1833 11.6369
R3555 GNDA.n1833 GNDA.n1831 11.6369
R3556 GNDA.n1831 GNDA.n1828 11.6369
R3557 GNDA.n1828 GNDA.n1827 11.6369
R3558 GNDA.n1827 GNDA.n1824 11.6369
R3559 GNDA.n1824 GNDA.n1823 11.6369
R3560 GNDA.n1823 GNDA.n1820 11.6369
R3561 GNDA.n1820 GNDA.n1819 11.6369
R3562 GNDA.n1865 GNDA.n1844 11.6369
R3563 GNDA.n1871 GNDA.n1844 11.6369
R3564 GNDA.n1872 GNDA.n1871 11.6369
R3565 GNDA.n1873 GNDA.n1872 11.6369
R3566 GNDA.n1873 GNDA.n1842 11.6369
R3567 GNDA.n1879 GNDA.n1842 11.6369
R3568 GNDA.n1880 GNDA.n1879 11.6369
R3569 GNDA.n1881 GNDA.n1880 11.6369
R3570 GNDA.n1881 GNDA.n1840 11.6369
R3571 GNDA.n1840 GNDA.n488 11.6369
R3572 GNDA.n895 GNDA.n438 11.6369
R3573 GNDA.n898 GNDA.n895 11.6369
R3574 GNDA.n899 GNDA.n898 11.6369
R3575 GNDA.n902 GNDA.n899 11.6369
R3576 GNDA.n903 GNDA.n902 11.6369
R3577 GNDA.n906 GNDA.n903 11.6369
R3578 GNDA.n907 GNDA.n906 11.6369
R3579 GNDA.n910 GNDA.n907 11.6369
R3580 GNDA.n911 GNDA.n910 11.6369
R3581 GNDA.n914 GNDA.n911 11.6369
R3582 GNDA.n915 GNDA.n914 11.6369
R3583 GNDA.n1864 GNDA.n1863 11.6369
R3584 GNDA.n1863 GNDA.n1860 11.6369
R3585 GNDA.n1860 GNDA.n1859 11.6369
R3586 GNDA.n1859 GNDA.n1856 11.6369
R3587 GNDA.n1856 GNDA.n1855 11.6369
R3588 GNDA.n1855 GNDA.n1852 11.6369
R3589 GNDA.n1852 GNDA.n1851 11.6369
R3590 GNDA.n1851 GNDA.n1848 11.6369
R3591 GNDA.n1848 GNDA.n1847 11.6369
R3592 GNDA.n1847 GNDA.n437 11.6369
R3593 GNDA.n2033 GNDA.n437 11.6369
R3594 GNDA.n819 GNDA.n818 11.6369
R3595 GNDA.n818 GNDA.n817 11.6369
R3596 GNDA.n817 GNDA.n815 11.6369
R3597 GNDA.n815 GNDA.n812 11.6369
R3598 GNDA.n812 GNDA.n811 11.6369
R3599 GNDA.n811 GNDA.n808 11.6369
R3600 GNDA.n808 GNDA.n807 11.6369
R3601 GNDA.n807 GNDA.n804 11.6369
R3602 GNDA.n804 GNDA.n803 11.6369
R3603 GNDA.n803 GNDA.n800 11.6369
R3604 GNDA.n2119 GNDA.n210 11.6369
R3605 GNDA.n2119 GNDA.n2118 11.6369
R3606 GNDA.n2118 GNDA.n2117 11.6369
R3607 GNDA.n2117 GNDA.n212 11.6369
R3608 GNDA.n2112 GNDA.n212 11.6369
R3609 GNDA.n2112 GNDA.n2111 11.6369
R3610 GNDA.n2111 GNDA.n2110 11.6369
R3611 GNDA.n2110 GNDA.n215 11.6369
R3612 GNDA.n2105 GNDA.n215 11.6369
R3613 GNDA.n2105 GNDA.n2104 11.6369
R3614 GNDA.n2104 GNDA.n2103 11.6369
R3615 GNDA.n529 GNDA.n528 11.6369
R3616 GNDA.n528 GNDA.n502 11.6369
R3617 GNDA.n523 GNDA.n502 11.6369
R3618 GNDA.n523 GNDA.n522 11.6369
R3619 GNDA.n522 GNDA.n521 11.6369
R3620 GNDA.n521 GNDA.n505 11.6369
R3621 GNDA.n516 GNDA.n505 11.6369
R3622 GNDA.n516 GNDA.n515 11.6369
R3623 GNDA.n515 GNDA.n514 11.6369
R3624 GNDA.n514 GNDA.n509 11.6369
R3625 GNDA.n509 GNDA.n508 11.6369
R3626 GNDA.n1497 GNDA.n1496 11.6369
R3627 GNDA.n1497 GNDA.n1289 11.6369
R3628 GNDA.n1504 GNDA.n1289 11.6369
R3629 GNDA.n1505 GNDA.n1504 11.6369
R3630 GNDA.n1506 GNDA.n1505 11.6369
R3631 GNDA.n1506 GNDA.n1287 11.6369
R3632 GNDA.n1511 GNDA.n1287 11.6369
R3633 GNDA.n1512 GNDA.n1511 11.6369
R3634 GNDA.n1514 GNDA.n1512 11.6369
R3635 GNDA.n1514 GNDA.n1513 11.6369
R3636 GNDA.n1473 GNDA.n1472 11.6369
R3637 GNDA.n1473 GNDA.n1301 11.6369
R3638 GNDA.n1479 GNDA.n1301 11.6369
R3639 GNDA.n1480 GNDA.n1479 11.6369
R3640 GNDA.n1481 GNDA.n1480 11.6369
R3641 GNDA.n1481 GNDA.n1297 11.6369
R3642 GNDA.n1487 GNDA.n1297 11.6369
R3643 GNDA.n1488 GNDA.n1487 11.6369
R3644 GNDA.n1489 GNDA.n1488 11.6369
R3645 GNDA.n1489 GNDA.n1293 11.6369
R3646 GNDA.n1495 GNDA.n1293 11.6369
R3647 GNDA.n1399 GNDA.n1398 11.6369
R3648 GNDA.n1401 GNDA.n1399 11.6369
R3649 GNDA.n1401 GNDA.n1400 11.6369
R3650 GNDA.n1400 GNDA.n1318 11.6369
R3651 GNDA.n1408 GNDA.n1318 11.6369
R3652 GNDA.n1415 GNDA.n1309 11.6369
R3653 GNDA.n1416 GNDA.n1415 11.6369
R3654 GNDA.n1418 GNDA.n1416 11.6369
R3655 GNDA.n1418 GNDA.n1417 11.6369
R3656 GNDA.n1417 GNDA.n1305 11.6369
R3657 GNDA.n2209 GNDA.n2208 11.473
R3658 GNDA.t55 GNDA.t36 10.7152
R3659 GNDA.t292 GNDA.n545 10.4196
R3660 GNDA.n92 GNDA.n0 9.75668
R3661 GNDA.n2283 GNDA.n2282 9.73997
R3662 GNDA.n2286 GNDA.n2285 9.73997
R3663 GNDA.n323 GNDA.n322 9.73997
R3664 GNDA.n326 GNDA.n325 9.73997
R3665 GNDA.n702 GNDA.t61 9.6005
R3666 GNDA.n703 GNDA.t57 9.6005
R3667 GNDA.n261 GNDA.t69 9.6005
R3668 GNDA.n261 GNDA.t216 9.6005
R3669 GNDA.n263 GNDA.t35 9.6005
R3670 GNDA.n263 GNDA.t273 9.6005
R3671 GNDA.n265 GNDA.t156 9.6005
R3672 GNDA.n265 GNDA.t67 9.6005
R3673 GNDA.n267 GNDA.t121 9.6005
R3674 GNDA.n267 GNDA.t112 9.6005
R3675 GNDA.n269 GNDA.t81 9.6005
R3676 GNDA.n269 GNDA.t99 9.6005
R3677 GNDA.n271 GNDA.t274 9.6005
R3678 GNDA.n271 GNDA.t49 9.6005
R3679 GNDA.n273 GNDA.t79 9.6005
R3680 GNDA.n273 GNDA.t97 9.6005
R3681 GNDA.n275 GNDA.t65 9.6005
R3682 GNDA.n275 GNDA.t47 9.6005
R3683 GNDA.n277 GNDA.t110 9.6005
R3684 GNDA.n277 GNDA.t154 9.6005
R3685 GNDA.n279 GNDA.t33 9.6005
R3686 GNDA.n279 GNDA.t71 9.6005
R3687 GNDA.n281 GNDA.t53 9.6005
R3688 GNDA.n281 GNDA.t119 9.6005
R3689 GNDA.n379 GNDA.n378 9.3005
R3690 GNDA.n341 GNDA.n340 9.3005
R3691 GNDA.n357 GNDA.n356 9.3005
R3692 GNDA.n344 GNDA.n342 9.04217
R3693 GNDA.n11 GNDA.n6 9.04217
R3694 GNDA.n2199 GNDA.n95 8.8452
R3695 GNDA.n353 GNDA.n251 8.79217
R3696 GNDA.n337 GNDA.n289 8.79217
R3697 GNDA.n2297 GNDA.n7 8.79217
R3698 GNDA.n2302 GNDA.n2301 8.79217
R3699 GNDA.n867 GNDA.n410 8.60107
R3700 GNDA.n467 GNDA.n407 8.60107
R3701 GNDA.t182 GNDA.t133 8.57228
R3702 GNDA.n2301 GNDA.n2299 8.34425
R3703 GNDA.n722 GNDA.t159 8.33581
R3704 GNDA.n597 GNDA.t339 8.33581
R3705 GNDA.n94 GNDA.n93 7.56675
R3706 GNDA.n1314 GNDA.n92 7.56675
R3707 GNDA.n19 GNDA.n5 7.46925
R3708 GNDA.n253 GNDA.n1 7.40675
R3709 GNDA.n2290 GNDA.n18 7.33383
R3710 GNDA.n2281 GNDA.n2280 7.33383
R3711 GNDA.n330 GNDA.n291 7.33383
R3712 GNDA.n321 GNDA.n320 7.33383
R3713 GNDA.n724 GNDA.t21 7.29389
R3714 GNDA.n2229 GNDA.t22 7.29389
R3715 GNDA.n2232 GNDA.t4 7.29389
R3716 GNDA.n109 GNDA.t1 7.29389
R3717 GNDA.n283 GNDA.n253 7.063
R3718 GNDA.n1392 GNDA.n1322 6.72373
R3719 GNDA.n1259 GNDA.n915 6.72373
R3720 GNDA.n2033 GNDA.n2032 6.72373
R3721 GNDA.n2103 GNDA.n218 6.72373
R3722 GNDA.n508 GNDA.n209 6.72373
R3723 GNDA.n1471 GNDA.n1305 6.72373
R3724 GNDA.n260 GNDA.n5 6.71925
R3725 GNDA.n2310 GNDA.n1 6.34425
R3726 GNDA.n2284 GNDA.n2283 6.313
R3727 GNDA.n2287 GNDA.n2286 6.313
R3728 GNDA.n324 GNDA.n323 6.313
R3729 GNDA.n327 GNDA.n326 6.313
R3730 GNDA.t288 GNDA.t182 6.25198
R3731 GNDA.n2283 GNDA.n2281 6.20883
R3732 GNDA.n2286 GNDA.n18 6.20883
R3733 GNDA.n323 GNDA.n321 6.20883
R3734 GNDA.n326 GNDA.n291 6.20883
R3735 GNDA.n221 GNDA.n218 6.20656
R3736 GNDA.n1259 GNDA.n894 6.20656
R3737 GNDA.n2032 GNDA.n438 6.20656
R3738 GNDA.n210 GNDA.n209 6.20656
R3739 GNDA.n1472 GNDA.n1471 6.20656
R3740 GNDA.n1398 GNDA.n1322 6.20656
R3741 GNDA.n1409 GNDA.n1408 6.07727
R3742 GNDA.n39 GNDA.n37 5.79217
R3743 GNDA.n24 GNDA.n23 5.79217
R3744 GNDA.n311 GNDA.n309 5.79217
R3745 GNDA.n296 GNDA.n295 5.79217
R3746 GNDA.n94 GNDA.n0 5.737
R3747 GNDA.n27 GNDA.n23 5.72967
R3748 GNDA.n299 GNDA.n295 5.72967
R3749 GNDA.n1409 GNDA.n1309 5.5601
R3750 GNDA.n354 GNDA.n353 5.53175
R3751 GNDA.n116 GNDA.n50 5.51161
R3752 GNDA.n1171 GNDA.n1141 5.51161
R3753 GNDA.n1751 GNDA.n1722 5.51161
R3754 GNDA.n1652 GNDA.n1622 5.51161
R3755 GNDA.n1055 GNDA.n945 5.51161
R3756 GNDA.n1936 GNDA.n1914 5.51161
R3757 GNDA.n620 GNDA.n100 5.51161
R3758 GNDA.n732 GNDA.n691 5.51161
R3759 GNDA.n1554 GNDA.n1524 5.51161
R3760 GNDA.n357 GNDA.n249 5.47967
R3761 GNDA.n378 GNDA.n247 5.47967
R3762 GNDA.n543 GNDA.n534 5.33383
R3763 GNDA.n2158 GNDA.n189 5.33383
R3764 GNDA.n2167 GNDA.n2164 5.33383
R3765 GNDA.n2180 GNDA.n2178 5.33383
R3766 GNDA.n2225 GNDA.n89 5.33383
R3767 GNDA.n2215 GNDA.n2212 5.33383
R3768 GNDA.n26 GNDA.n24 5.22967
R3769 GNDA.n29 GNDA.n21 5.22967
R3770 GNDA.n34 GNDA.n33 5.22967
R3771 GNDA.n37 GNDA.n36 5.22967
R3772 GNDA.n298 GNDA.n296 5.22967
R3773 GNDA.n301 GNDA.n293 5.22967
R3774 GNDA.n306 GNDA.n305 5.22967
R3775 GNDA.n309 GNDA.n308 5.22967
R3776 GNDA.t3 GNDA.t89 5.21007
R3777 GNDA.n706 GNDA.t161 5.21007
R3778 GNDA.t124 GNDA.t276 5.21007
R3779 GNDA.t182 GNDA.t334 5.21007
R3780 GNDA.n2270 GNDA.n2269 5.1717
R3781 GNDA.n1140 GNDA.n1081 5.1717
R3782 GNDA.n1523 GNDA.n1282 5.1717
R3783 GNDA.n27 GNDA.n26 5.16717
R3784 GNDA.n30 GNDA.n29 5.16717
R3785 GNDA.n33 GNDA.n31 5.16717
R3786 GNDA.n36 GNDA.n20 5.16717
R3787 GNDA.n40 GNDA.n39 5.16717
R3788 GNDA.n299 GNDA.n298 5.16717
R3789 GNDA.n302 GNDA.n301 5.16717
R3790 GNDA.n305 GNDA.n303 5.16717
R3791 GNDA.n308 GNDA.n292 5.16717
R3792 GNDA.n312 GNDA.n311 5.16717
R3793 GNDA.n542 GNDA.n541 5.063
R3794 GNDA.n377 GNDA.n376 5.063
R3795 GNDA.n2309 GNDA.n2308 5.02133
R3796 GNDA.n254 GNDA.n2 5.02133
R3797 GNDA.n375 GNDA.n247 4.91717
R3798 GNDA.n372 GNDA.n370 4.91717
R3799 GNDA.n369 GNDA.n368 4.91717
R3800 GNDA.n366 GNDA.n365 4.91717
R3801 GNDA.n361 GNDA.n249 4.91717
R3802 GNDA.n1816 GNDA.n826 4.9157
R3803 GNDA.n2000 GNDA.n1888 4.9157
R3804 GNDA.n799 GNDA.n798 4.9157
R3805 GNDA.n188 GNDA.n186 4.83383
R3806 GNDA.n538 GNDA.n537 4.83383
R3807 GNDA.n541 GNDA.n540 4.83383
R3808 GNDA.n2177 GNDA.n2175 4.83383
R3809 GNDA.n2174 GNDA.n2173 4.83383
R3810 GNDA.n2171 GNDA.n2170 4.83383
R3811 GNDA.n2166 GNDA.n185 4.83383
R3812 GNDA.n2214 GNDA.n91 4.83383
R3813 GNDA.n2219 GNDA.n2218 4.83383
R3814 GNDA.n2222 GNDA.n2221 4.83383
R3815 GNDA.n342 GNDA.n341 4.79217
R3816 GNDA.n337 GNDA.n336 4.79217
R3817 GNDA.n2297 GNDA.n2296 4.79217
R3818 GNDA.n14 GNDA.n6 4.79217
R3819 GNDA.n2204 GNDA.n2203 4.7827
R3820 GNDA.n189 GNDA.n188 4.77133
R3821 GNDA.n537 GNDA.n535 4.77133
R3822 GNDA.n540 GNDA.n534 4.77133
R3823 GNDA.n2178 GNDA.n2177 4.77133
R3824 GNDA.n2173 GNDA.n184 4.77133
R3825 GNDA.n2170 GNDA.n2168 4.77133
R3826 GNDA.n2167 GNDA.n2166 4.77133
R3827 GNDA.n2215 GNDA.n2214 4.77133
R3828 GNDA.n2218 GNDA.n2216 4.77133
R3829 GNDA.n2221 GNDA.n89 4.77133
R3830 GNDA.n376 GNDA.n375 4.72967
R3831 GNDA.n373 GNDA.n372 4.72967
R3832 GNDA.n368 GNDA.n248 4.72967
R3833 GNDA.n365 GNDA.n363 4.72967
R3834 GNDA.n362 GNDA.n361 4.72967
R3835 GNDA.n2289 GNDA.n2288 4.70883
R3836 GNDA.n42 GNDA.n41 4.70883
R3837 GNDA.n329 GNDA.n328 4.70883
R3838 GNDA.n314 GNDA.n313 4.70883
R3839 GNDA.n2158 GNDA.n2157 4.6505
R3840 GNDA.n2164 GNDA.n2163 4.6505
R3841 GNDA.n2181 GNDA.n2180 4.6505
R3842 GNDA.n2226 GNDA.n2225 4.6505
R3843 GNDA.n2212 GNDA.n2211 4.6505
R3844 GNDA.n544 GNDA.n543 4.6505
R3845 GNDA.n2210 GNDA.n2209 4.5005
R3846 GNDA.n2224 GNDA.n2223 4.5005
R3847 GNDA.n2179 GNDA.n90 4.5005
R3848 GNDA.n2162 GNDA.n2161 4.5005
R3849 GNDA.n2160 GNDA.n2159 4.5005
R3850 GNDA.n284 GNDA.n283 4.5005
R3851 GNDA.n260 GNDA.n259 4.5005
R3852 GNDA.n2299 GNDA.n2298 4.5005
R3853 GNDA.n338 GNDA.n250 4.5005
R3854 GNDA.n359 GNDA.n358 4.5005
R3855 GNDA.n2125 GNDA.n207 4.26717
R3856 GNDA.n2131 GNDA.n207 4.26717
R3857 GNDA.n2131 GNDA.n203 4.26717
R3858 GNDA.n2136 GNDA.n203 4.26717
R3859 GNDA.n2136 GNDA.n201 4.26717
R3860 GNDA.n201 GNDA.n198 4.26717
R3861 GNDA.n2143 GNDA.n198 4.26717
R3862 GNDA.n2143 GNDA.n196 4.26717
R3863 GNDA.n196 GNDA.n194 4.26717
R3864 GNDA.n2150 GNDA.n194 4.26717
R3865 GNDA.n2150 GNDA.n192 4.26717
R3866 GNDA.n2031 GNDA.n440 4.26717
R3867 GNDA.n2026 GNDA.n440 4.26717
R3868 GNDA.n2026 GNDA.n2025 4.26717
R3869 GNDA.n2025 GNDA.n2024 4.26717
R3870 GNDA.n2024 GNDA.n449 4.26717
R3871 GNDA.n2018 GNDA.n449 4.26717
R3872 GNDA.n2018 GNDA.n2017 4.26717
R3873 GNDA.n2017 GNDA.n2016 4.26717
R3874 GNDA.n2016 GNDA.n457 4.26717
R3875 GNDA.n2010 GNDA.n457 4.26717
R3876 GNDA.n2010 GNDA.n2009 4.26717
R3877 GNDA.n1362 GNDA.n1361 4.26717
R3878 GNDA.n1361 GNDA.n1328 4.26717
R3879 GNDA.n1355 GNDA.n1328 4.26717
R3880 GNDA.n1355 GNDA.n1354 4.26717
R3881 GNDA.n1354 GNDA.n1353 4.26717
R3882 GNDA.n1353 GNDA.n1336 4.26717
R3883 GNDA.n1338 GNDA.n1336 4.26717
R3884 GNDA.n1344 GNDA.n1338 4.26717
R3885 GNDA.n1345 GNDA.n1344 4.26717
R3886 GNDA.n1345 GNDA.n869 4.26717
R3887 GNDA.n1717 GNDA.n869 4.26717
R3888 GNDA.n1470 GNDA.n1426 4.26717
R3889 GNDA.n1465 GNDA.n1426 4.26717
R3890 GNDA.n1465 GNDA.n1464 4.26717
R3891 GNDA.n1464 GNDA.n1433 4.26717
R3892 GNDA.n1459 GNDA.n1433 4.26717
R3893 GNDA.n1459 GNDA.n1458 4.26717
R3894 GNDA.n1458 GNDA.n1457 4.26717
R3895 GNDA.n1457 GNDA.n1441 4.26717
R3896 GNDA.n1451 GNDA.n1441 4.26717
R3897 GNDA.n1451 GNDA.n1450 4.26717
R3898 GNDA.n1450 GNDA.n1449 4.26717
R3899 GNDA.n1258 GNDA.n918 4.26717
R3900 GNDA.n1252 GNDA.n918 4.26717
R3901 GNDA.n1252 GNDA.n1251 4.26717
R3902 GNDA.n1251 GNDA.n1250 4.26717
R3903 GNDA.n1250 GNDA.n1248 4.26717
R3904 GNDA.n1248 GNDA.n1245 4.26717
R3905 GNDA.n1245 GNDA.n1244 4.26717
R3906 GNDA.n1244 GNDA.n1241 4.26717
R3907 GNDA.n1241 GNDA.n1240 4.26717
R3908 GNDA.n1240 GNDA.n1237 4.26717
R3909 GNDA.n1237 GNDA.n1236 4.26717
R3910 GNDA.n2100 GNDA.n220 4.26717
R3911 GNDA.n2095 GNDA.n220 4.26717
R3912 GNDA.n2095 GNDA.n2094 4.26717
R3913 GNDA.n2094 GNDA.n2076 4.26717
R3914 GNDA.n2089 GNDA.n2076 4.26717
R3915 GNDA.n2089 GNDA.n2088 4.26717
R3916 GNDA.n2088 GNDA.n2087 4.26717
R3917 GNDA.n2087 GNDA.n2082 4.26717
R3918 GNDA.n2082 GNDA.n172 4.26717
R3919 GNDA.n2187 GNDA.n172 4.26717
R3920 GNDA.n2187 GNDA.n170 4.26717
R3921 GNDA GNDA.n2311 4.2117
R3922 GNDA.n2156 GNDA.n2155 4.16815
R3923 GNDA.n2204 GNDA.n2199 4.063
R3924 GNDA.t205 GNDA.t271 3.99324
R3925 GNDA.t326 GNDA.t196 3.99324
R3926 GNDA.n2306 GNDA.t48 3.99324
R3927 GNDA.t179 GNDA.n2305 3.99324
R3928 GNDA.t17 GNDA.n256 3.99324
R3929 GNDA.t311 GNDA.t243 3.99324
R3930 GNDA.n2125 GNDA.n209 3.93531
R3931 GNDA.n2032 GNDA.n2031 3.93531
R3932 GNDA.n1362 GNDA.n1322 3.93531
R3933 GNDA.n1471 GNDA.n1470 3.93531
R3934 GNDA.n1259 GNDA.n1258 3.93531
R3935 GNDA.n2100 GNDA.n218 3.93531
R3936 GNDA.n2247 GNDA.n85 3.7893
R3937 GNDA.n2246 GNDA.n86 3.7893
R3938 GNDA.n2234 GNDA.n2233 3.7893
R3939 GNDA.n2240 GNDA.n2239 3.7893
R3940 GNDA.n2236 GNDA.n2235 3.7893
R3941 GNDA.n103 GNDA.n64 3.7893
R3942 GNDA.n104 GNDA.n102 3.7893
R3943 GNDA.n113 GNDA.n111 3.7893
R3944 GNDA.n1230 GNDA.n1061 3.7893
R3945 GNDA.n1227 GNDA.n1226 3.7893
R3946 GNDA.n1143 GNDA.n1062 3.7893
R3947 GNDA.n1148 GNDA.n1146 3.7893
R3948 GNDA.n1153 GNDA.n1149 3.7893
R3949 GNDA.n1160 GNDA.n1159 3.7893
R3950 GNDA.n1163 GNDA.n1142 3.7893
R3951 GNDA.n1168 GNDA.n1164 3.7893
R3952 GNDA.n1711 GNDA.n872 3.7893
R3953 GNDA.n1708 GNDA.n1707 3.7893
R3954 GNDA.n1624 GNDA.n873 3.7893
R3955 GNDA.n1629 GNDA.n1627 3.7893
R3956 GNDA.n1634 GNDA.n1630 3.7893
R3957 GNDA.n1641 GNDA.n1640 3.7893
R3958 GNDA.n1644 GNDA.n1623 3.7893
R3959 GNDA.n1649 GNDA.n1645 3.7893
R3960 GNDA.n1801 GNDA.n845 3.7893
R3961 GNDA.n1809 GNDA.n1808 3.7893
R3962 GNDA.n1724 GNDA.n846 3.7893
R3963 GNDA.n1728 GNDA.n1726 3.7893
R3964 GNDA.n1733 GNDA.n1729 3.7893
R3965 GNDA.n1740 GNDA.n1739 3.7893
R3966 GNDA.n1743 GNDA.n1723 3.7893
R3967 GNDA.n1748 GNDA.n1744 3.7893
R3968 GNDA.n1045 GNDA.n1021 3.7893
R3969 GNDA.n1044 GNDA.n1042 3.7893
R3970 GNDA.n1041 GNDA.n1022 3.7893
R3971 GNDA.n1038 GNDA.n1037 3.7893
R3972 GNDA.n1034 GNDA.n1023 3.7893
R3973 GNDA.n1027 GNDA.n1024 3.7893
R3974 GNDA.n1050 GNDA.n947 3.7893
R3975 GNDA.n1051 GNDA.n946 3.7893
R3976 GNDA.n1998 GNDA.n1997 3.7893
R3977 GNDA.n1994 GNDA.n1891 3.7893
R3978 GNDA.n1993 GNDA.n1894 3.7893
R3979 GNDA.n1990 GNDA.n1989 3.7893
R3980 GNDA.n1916 GNDA.n1895 3.7893
R3981 GNDA.n1925 GNDA.n1924 3.7893
R3982 GNDA.n1928 GNDA.n1915 3.7893
R3983 GNDA.n1933 GNDA.n1929 3.7893
R3984 GNDA.n673 GNDA.n568 3.7893
R3985 GNDA.n672 GNDA.n570 3.7893
R3986 GNDA.n679 GNDA.n678 3.7893
R3987 GNDA.n595 GNDA.n571 3.7893
R3988 GNDA.n601 GNDA.n599 3.7893
R3989 GNDA.n608 GNDA.n607 3.7893
R3990 GNDA.n615 GNDA.n591 3.7893
R3991 GNDA.n614 GNDA.n589 3.7893
R3992 GNDA.n785 GNDA.n533 3.7893
R3993 GNDA.n784 GNDA.n548 3.7893
R3994 GNDA.n791 GNDA.n790 3.7893
R3995 GNDA.n709 GNDA.n549 3.7893
R3996 GNDA.n713 GNDA.n711 3.7893
R3997 GNDA.n720 GNDA.n719 3.7893
R3998 GNDA.n727 GNDA.n695 3.7893
R3999 GNDA.n726 GNDA.n693 3.7893
R4000 GNDA.n1613 GNDA.n1262 3.7893
R4001 GNDA.n1610 GNDA.n1609 3.7893
R4002 GNDA.n1526 GNDA.n1263 3.7893
R4003 GNDA.n1531 GNDA.n1529 3.7893
R4004 GNDA.n1536 GNDA.n1532 3.7893
R4005 GNDA.n1543 GNDA.n1542 3.7893
R4006 GNDA.n1546 GNDA.n1525 3.7893
R4007 GNDA.n1551 GNDA.n1547 3.7893
R4008 GNDA GNDA.n2252 3.7381
R4009 GNDA.n1156 GNDA 3.7381
R4010 GNDA.n1637 GNDA 3.7381
R4011 GNDA.n1736 GNDA 3.7381
R4012 GNDA GNDA.n1030 3.7381
R4013 GNDA.n1921 GNDA 3.7381
R4014 GNDA.n606 GNDA 3.7381
R4015 GNDA.n718 GNDA 3.7381
R4016 GNDA.n1539 GNDA 3.7381
R4017 GNDA.n347 GNDA.n287 3.65764
R4018 GNDA.n347 GNDA.n346 3.65764
R4019 GNDA.n9 GNDA.n3 3.65764
R4020 GNDA.n12 GNDA.n3 3.65764
R4021 GNDA.n19 GNDA.n2 3.53175
R4022 GNDA.n253 GNDA.n250 3.53175
R4023 GNDA.n2299 GNDA.n5 3.46925
R4024 GNDA.n2282 GNDA.t94 3.42907
R4025 GNDA.n2282 GNDA.t24 3.42907
R4026 GNDA.n2285 GNDA.t322 3.42907
R4027 GNDA.n2285 GNDA.t285 3.42907
R4028 GNDA.n322 GNDA.t287 3.42907
R4029 GNDA.n322 GNDA.t8 3.42907
R4030 GNDA.n325 GNDA.t296 3.42907
R4031 GNDA.n325 GNDA.t96 3.42907
R4032 GNDA.n2308 GNDA.n2307 3.39217
R4033 GNDA.n255 GNDA.n254 3.39217
R4034 GNDA.n2208 GNDA.n92 3.32575
R4035 GNDA.t9 GNDA.n794 3.12624
R4036 GNDA.n707 GNDA.t293 3.12624
R4037 GNDA.n699 GNDA.t290 3.12624
R4038 GNDA.n2244 GNDA.t276 3.12624
R4039 GNDA.n350 GNDA.n349 3.1005
R4040 GNDA.n339 GNDA.n288 3.1005
R4041 GNDA.n345 GNDA.n287 3.1005
R4042 GNDA.n346 GNDA.n345 3.1005
R4043 GNDA.n16 GNDA.n15 3.1005
R4044 GNDA.n13 GNDA.n9 3.1005
R4045 GNDA.n13 GNDA.n12 3.1005
R4046 GNDA.n2304 GNDA.n2303 3.1005
R4047 GNDA.n354 GNDA.n250 2.813
R4048 GNDA.n169 GNDA.n168 2.6629
R4049 GNDA.n1232 GNDA.n1231 2.6629
R4050 GNDA.n1713 GNDA.n1712 2.6629
R4051 GNDA.n1621 GNDA.n892 2.6629
R4052 GNDA.n1802 GNDA.n826 2.6629
R4053 GNDA.n1721 GNDA.n866 2.6629
R4054 GNDA.n1020 GNDA.n464 2.6629
R4055 GNDA.n1056 GNDA.n944 2.6629
R4056 GNDA.n2000 GNDA.n1999 2.6629
R4057 GNDA.n2008 GNDA.n465 2.6629
R4058 GNDA.n688 GNDA.n565 2.6629
R4059 GNDA.n2194 GNDA.n2193 2.6629
R4060 GNDA.n798 GNDA.n531 2.6629
R4061 GNDA.n690 GNDA.n689 2.6629
R4062 GNDA.n1615 GNDA.n1614 2.6629
R4063 GNDA.n2193 GNDA.n169 2.4581
R4064 GNDA.n2270 GNDA.n50 2.4581
R4065 GNDA.n1232 GNDA.n944 2.4581
R4066 GNDA.n1141 GNDA.n1140 2.4581
R4067 GNDA.n1713 GNDA.n866 2.4581
R4068 GNDA.n1622 GNDA.n1621 2.4581
R4069 GNDA.n1722 GNDA.n1721 2.4581
R4070 GNDA.n2008 GNDA.n464 2.4581
R4071 GNDA.n1056 GNDA.n1055 2.4581
R4072 GNDA.n1914 GNDA.n465 2.4581
R4073 GNDA.n689 GNDA.n688 2.4581
R4074 GNDA.n2194 GNDA.n100 2.4581
R4075 GNDA.n691 GNDA.n690 2.4581
R4076 GNDA.n1615 GNDA.n892 2.4581
R4077 GNDA.n1524 GNDA.n1523 2.4581
R4078 GNDA.n2205 GNDA 2.26825
R4079 GNDA.n285 GNDA.n284 2.19633
R4080 GNDA.n689 GNDA.n192 2.18124
R4081 GNDA.n2009 GNDA.n2008 2.18124
R4082 GNDA.n1717 GNDA.n866 2.18124
R4083 GNDA.n1449 GNDA.n892 2.18124
R4084 GNDA.n1236 GNDA.n944 2.18124
R4085 GNDA.n2193 GNDA.n170 2.18124
R4086 GNDA.n112 GNDA.n50 2.1509
R4087 GNDA.n1167 GNDA.n1141 2.1509
R4088 GNDA.n1648 GNDA.n1622 2.1509
R4089 GNDA.n1747 GNDA.n1722 2.1509
R4090 GNDA.n1055 GNDA.n1054 2.1509
R4091 GNDA.n1932 GNDA.n1914 2.1509
R4092 GNDA.n588 GNDA.n100 2.1509
R4093 GNDA.n697 GNDA.n691 2.1509
R4094 GNDA.n1550 GNDA.n1524 2.1509
R4095 GNDA.n2202 GNDA.n2201 2.13383
R4096 GNDA.n168 GNDA.n167 2.13383
R4097 GNDA.n1231 GNDA.n1060 2.13383
R4098 GNDA.n1803 GNDA.n1802 2.13383
R4099 GNDA.n1712 GNDA.n871 2.13383
R4100 GNDA.n1020 GNDA.n1019 2.13383
R4101 GNDA.n1999 GNDA.n1889 2.13383
R4102 GNDA.n669 GNDA.n565 2.13383
R4103 GNDA.n781 GNDA.n531 2.13383
R4104 GNDA.n1614 GNDA.n1261 2.13383
R4105 GNDA.n705 GNDA.n704 2.13383
R4106 GNDA.n689 GNDA.n191 2.08643
R4107 GNDA.n2008 GNDA.n2007 2.08643
R4108 GNDA.n866 GNDA.n439 2.08643
R4109 GNDA.n1618 GNDA.n892 2.08643
R4110 GNDA.n1059 GNDA.n944 2.08643
R4111 GNDA.n2193 GNDA.n2192 2.08643
R4112 GNDA.n794 GNDA.t219 2.08433
R4113 GNDA.n686 GNDA.t240 2.08433
R4114 GNDA.n2196 GNDA.t192 2.08433
R4115 GNDA.t151 GNDA.n107 2.08433
R4116 GNDA.n168 GNDA.n85 1.9461
R4117 GNDA.n1231 GNDA.n1230 1.9461
R4118 GNDA.n1712 GNDA.n1711 1.9461
R4119 GNDA.n1802 GNDA.n1801 1.9461
R4120 GNDA.n1021 GNDA.n1020 1.9461
R4121 GNDA.n1999 GNDA.n1998 1.9461
R4122 GNDA.n568 GNDA.n565 1.9461
R4123 GNDA.n533 GNDA.n531 1.9461
R4124 GNDA.n1614 GNDA.n1613 1.9461
R4125 GNDA.n2309 GNDA.n2 1.938
R4126 GNDA.n259 GNDA.n258 1.91062
R4127 GNDA.n1315 GNDA.n1314 1.90675
R4128 GNDA.n404 GNDA.t60 1.8483
R4129 GNDA.n2290 GNDA.n2289 1.60467
R4130 GNDA.n2280 GNDA.n42 1.60467
R4131 GNDA.n330 GNDA.n329 1.60467
R4132 GNDA.n320 GNDA.n314 1.60467
R4133 GNDA.n2203 GNDA.n2202 1.5505
R4134 GNDA.n704 GNDA.n95 1.5505
R4135 GNDA.n328 GNDA.n1 1.53175
R4136 GNDA.n2288 GNDA.n19 1.5005
R4137 GNDA.n2269 GNDA.n2268 1.47392
R4138 GNDA.n1130 GNDA.n1081 1.47392
R4139 GNDA.n1819 GNDA.n1816 1.47392
R4140 GNDA.n1888 GNDA.n488 1.47392
R4141 GNDA.n800 GNDA.n799 1.47392
R4142 GNDA.n1513 GNDA.n1282 1.47392
R4143 GNDA.n338 GNDA.n337 1.34425
R4144 GNDA.n2298 GNDA.n2297 1.34425
R4145 GNDA.n335 GNDA.n334 1.163
R4146 GNDA.n316 GNDA.n290 1.163
R4147 GNDA.n2295 GNDA.n2294 1.163
R4148 GNDA.n2276 GNDA.n8 1.163
R4149 GNDA.n2281 GNDA.n18 1.1255
R4150 GNDA.n2284 GNDA.n41 1.1255
R4151 GNDA.n2287 GNDA.n2284 1.1255
R4152 GNDA.n2288 GNDA.n2287 1.1255
R4153 GNDA.n321 GNDA.n291 1.1255
R4154 GNDA.n324 GNDA.n313 1.1255
R4155 GNDA.n327 GNDA.n324 1.1255
R4156 GNDA.n328 GNDA.n327 1.1255
R4157 GNDA.n342 GNDA.n338 1.03175
R4158 GNDA.n2298 GNDA.n6 1.03175
R4159 GNDA.n2223 GNDA.n90 0.8755
R4160 GNDA.n2247 GNDA.n2246 0.8197
R4161 GNDA.n2233 GNDA.n86 0.8197
R4162 GNDA.n2240 GNDA.n2234 0.8197
R4163 GNDA.n2239 GNDA.n2236 0.8197
R4164 GNDA.n2252 GNDA.n64 0.8197
R4165 GNDA.n104 GNDA.n103 0.8197
R4166 GNDA.n111 GNDA.n102 0.8197
R4167 GNDA.n113 GNDA.n112 0.8197
R4168 GNDA.n1227 GNDA.n1061 0.8197
R4169 GNDA.n1226 GNDA.n1062 0.8197
R4170 GNDA.n1146 GNDA.n1143 0.8197
R4171 GNDA.n1149 GNDA.n1148 0.8197
R4172 GNDA.n1159 GNDA.n1156 0.8197
R4173 GNDA.n1160 GNDA.n1142 0.8197
R4174 GNDA.n1164 GNDA.n1163 0.8197
R4175 GNDA.n1168 GNDA.n1167 0.8197
R4176 GNDA.n1708 GNDA.n872 0.8197
R4177 GNDA.n1707 GNDA.n873 0.8197
R4178 GNDA.n1627 GNDA.n1624 0.8197
R4179 GNDA.n1630 GNDA.n1629 0.8197
R4180 GNDA.n1640 GNDA.n1637 0.8197
R4181 GNDA.n1641 GNDA.n1623 0.8197
R4182 GNDA.n1645 GNDA.n1644 0.8197
R4183 GNDA.n1649 GNDA.n1648 0.8197
R4184 GNDA.n1809 GNDA.n845 0.8197
R4185 GNDA.n1808 GNDA.n846 0.8197
R4186 GNDA.n1726 GNDA.n1724 0.8197
R4187 GNDA.n1729 GNDA.n1728 0.8197
R4188 GNDA.n1739 GNDA.n1736 0.8197
R4189 GNDA.n1740 GNDA.n1723 0.8197
R4190 GNDA.n1744 GNDA.n1743 0.8197
R4191 GNDA.n1748 GNDA.n1747 0.8197
R4192 GNDA.n1045 GNDA.n1044 0.8197
R4193 GNDA.n1042 GNDA.n1041 0.8197
R4194 GNDA.n1038 GNDA.n1022 0.8197
R4195 GNDA.n1037 GNDA.n1034 0.8197
R4196 GNDA.n1030 GNDA.n1027 0.8197
R4197 GNDA.n1024 GNDA.n947 0.8197
R4198 GNDA.n1051 GNDA.n1050 0.8197
R4199 GNDA.n1054 GNDA.n946 0.8197
R4200 GNDA.n1997 GNDA.n1891 0.8197
R4201 GNDA.n1994 GNDA.n1993 0.8197
R4202 GNDA.n1990 GNDA.n1894 0.8197
R4203 GNDA.n1989 GNDA.n1895 0.8197
R4204 GNDA.n1924 GNDA.n1921 0.8197
R4205 GNDA.n1925 GNDA.n1915 0.8197
R4206 GNDA.n1929 GNDA.n1928 0.8197
R4207 GNDA.n1933 GNDA.n1932 0.8197
R4208 GNDA.n673 GNDA.n672 0.8197
R4209 GNDA.n679 GNDA.n570 0.8197
R4210 GNDA.n678 GNDA.n571 0.8197
R4211 GNDA.n599 GNDA.n595 0.8197
R4212 GNDA.n608 GNDA.n606 0.8197
R4213 GNDA.n607 GNDA.n591 0.8197
R4214 GNDA.n615 GNDA.n614 0.8197
R4215 GNDA.n589 GNDA.n588 0.8197
R4216 GNDA.n785 GNDA.n784 0.8197
R4217 GNDA.n791 GNDA.n548 0.8197
R4218 GNDA.n790 GNDA.n549 0.8197
R4219 GNDA.n711 GNDA.n709 0.8197
R4220 GNDA.n720 GNDA.n718 0.8197
R4221 GNDA.n719 GNDA.n695 0.8197
R4222 GNDA.n727 GNDA.n726 0.8197
R4223 GNDA.n697 GNDA.n693 0.8197
R4224 GNDA.n1610 GNDA.n1262 0.8197
R4225 GNDA.n1609 GNDA.n1263 0.8197
R4226 GNDA.n1529 GNDA.n1526 0.8197
R4227 GNDA.n1532 GNDA.n1531 0.8197
R4228 GNDA.n1542 GNDA.n1539 0.8197
R4229 GNDA.n1543 GNDA.n1525 0.8197
R4230 GNDA.n1547 GNDA.n1546 0.8197
R4231 GNDA.n1551 GNDA.n1550 0.8197
R4232 GNDA.n2161 GNDA.n2160 0.813
R4233 GNDA.n336 GNDA.n335 0.771333
R4234 GNDA.n290 GNDA.n289 0.771333
R4235 GNDA.n2296 GNDA.n2295 0.771333
R4236 GNDA.n8 GNDA.n7 0.771333
R4237 GNDA.n2201 GNDA.n2200 0.632847
R4238 GNDA.n705 GNDA.n701 0.632847
R4239 GNDA.n2310 GNDA.n2309 0.6255
R4240 GNDA.n1839 GNDA.n404 0.574752
R4241 GNDA.n2235 GNDA 0.5637
R4242 GNDA.n1153 GNDA 0.5637
R4243 GNDA.n1634 GNDA 0.5637
R4244 GNDA.n1733 GNDA 0.5637
R4245 GNDA GNDA.n1023 0.5637
R4246 GNDA GNDA.n1916 0.5637
R4247 GNDA.n601 GNDA 0.5637
R4248 GNDA.n713 GNDA 0.5637
R4249 GNDA.n1536 GNDA 0.5637
R4250 GNDA.n535 GNDA.n534 0.563
R4251 GNDA.n535 GNDA.n189 0.563
R4252 GNDA.n2168 GNDA.n2167 0.563
R4253 GNDA.n2168 GNDA.n184 0.563
R4254 GNDA.n2178 GNDA.n184 0.563
R4255 GNDA.n2216 GNDA.n89 0.563
R4256 GNDA.n2216 GNDA.n2215 0.563
R4257 GNDA.n2209 GNDA.n91 0.563
R4258 GNDA.n2219 GNDA.n91 0.563
R4259 GNDA.n2222 GNDA.n2219 0.563
R4260 GNDA.n2223 GNDA.n2222 0.563
R4261 GNDA.n2175 GNDA.n90 0.563
R4262 GNDA.n2175 GNDA.n2174 0.563
R4263 GNDA.n2174 GNDA.n2171 0.563
R4264 GNDA.n2171 GNDA.n185 0.563
R4265 GNDA.n2161 GNDA.n185 0.563
R4266 GNDA.n2160 GNDA.n186 0.563
R4267 GNDA.n538 GNDA.n186 0.563
R4268 GNDA.n541 GNDA.n538 0.563
R4269 GNDA.n366 GNDA.n249 0.563
R4270 GNDA.n369 GNDA.n366 0.563
R4271 GNDA.n370 GNDA.n369 0.563
R4272 GNDA.n370 GNDA.n247 0.563
R4273 GNDA.n376 GNDA.n373 0.563
R4274 GNDA.n373 GNDA.n248 0.563
R4275 GNDA.n363 GNDA.n248 0.563
R4276 GNDA.n363 GNDA.n362 0.563
R4277 GNDA.n362 GNDA.n359 0.563
R4278 GNDA.n283 GNDA.n282 0.563
R4279 GNDA.n282 GNDA.n280 0.563
R4280 GNDA.n280 GNDA.n278 0.563
R4281 GNDA.n278 GNDA.n276 0.563
R4282 GNDA.n276 GNDA.n274 0.563
R4283 GNDA.n274 GNDA.n272 0.563
R4284 GNDA.n272 GNDA.n270 0.563
R4285 GNDA.n270 GNDA.n268 0.563
R4286 GNDA.n268 GNDA.n266 0.563
R4287 GNDA.n266 GNDA.n264 0.563
R4288 GNDA.n264 GNDA.n262 0.563
R4289 GNDA.n37 GNDA.n34 0.563
R4290 GNDA.n34 GNDA.n21 0.563
R4291 GNDA.n24 GNDA.n21 0.563
R4292 GNDA.n30 GNDA.n27 0.563
R4293 GNDA.n31 GNDA.n30 0.563
R4294 GNDA.n31 GNDA.n20 0.563
R4295 GNDA.n40 GNDA.n20 0.563
R4296 GNDA.n309 GNDA.n306 0.563
R4297 GNDA.n306 GNDA.n293 0.563
R4298 GNDA.n296 GNDA.n293 0.563
R4299 GNDA.n302 GNDA.n299 0.563
R4300 GNDA.n303 GNDA.n302 0.563
R4301 GNDA.n303 GNDA.n292 0.563
R4302 GNDA.n312 GNDA.n292 0.563
R4303 GNDA.t182 GNDA.t36 0.536236
R4304 GNDA.n2291 GNDA.n2290 0.489974
R4305 GNDA.n2280 GNDA.n2279 0.489974
R4306 GNDA.n331 GNDA.n330 0.489974
R4307 GNDA.n320 GNDA.n319 0.489974
R4308 GNDA.n2203 GNDA.n2200 0.460076
R4309 GNDA.n701 GNDA.n95 0.460076
R4310 GNDA.n341 GNDA.n288 0.458833
R4311 GNDA.n15 GNDA.n14 0.458833
R4312 GNDA.n2159 GNDA.n2158 0.333833
R4313 GNDA.n2164 GNDA.n2162 0.333833
R4314 GNDA.n2180 GNDA.n2179 0.333833
R4315 GNDA.n2225 GNDA.n2224 0.333833
R4316 GNDA.n2212 GNDA.n2210 0.333833
R4317 GNDA.n543 GNDA.n542 0.333833
R4318 GNDA.n2208 GNDA.n2207 0.300125
R4319 GNDA.n350 GNDA.n251 0.292167
R4320 GNDA.n2303 GNDA.n2302 0.292167
R4321 GNDA.n2253 GNDA 0.2565
R4322 GNDA GNDA.n1152 0.2565
R4323 GNDA GNDA.n1633 0.2565
R4324 GNDA GNDA.n1732 0.2565
R4325 GNDA.n1031 GNDA 0.2565
R4326 GNDA.n1919 GNDA 0.2565
R4327 GNDA GNDA.n600 0.2565
R4328 GNDA GNDA.n712 0.2565
R4329 GNDA GNDA.n1535 0.2565
R4330 GNDA.n345 GNDA.n344 0.246712
R4331 GNDA.n13 GNDA.n11 0.246712
R4332 GNDA.n378 GNDA.n377 0.229667
R4333 GNDA.n358 GNDA.n357 0.229667
R4334 GNDA.n262 GNDA.n260 0.21925
R4335 GNDA.n2207 GNDA.n2205 0.217875
R4336 GNDA.n2253 GNDA 0.0517
R4337 GNDA.n1152 GNDA 0.0517
R4338 GNDA.n1633 GNDA 0.0517
R4339 GNDA.n1732 GNDA 0.0517
R4340 GNDA.n1031 GNDA 0.0517
R4341 GNDA GNDA.n1919 0.0517
R4342 GNDA.n600 GNDA 0.0517
R4343 GNDA.n712 GNDA 0.0517
R4344 GNDA.n1535 GNDA 0.0517
R4345 two_stage_opamp_dummy_magic_0.Y.n61 two_stage_opamp_dummy_magic_0.Y.t34 1172.87
R4346 two_stage_opamp_dummy_magic_0.Y.n64 two_stage_opamp_dummy_magic_0.Y.t26 1172.87
R4347 two_stage_opamp_dummy_magic_0.Y.n68 two_stage_opamp_dummy_magic_0.Y.t28 996.134
R4348 two_stage_opamp_dummy_magic_0.Y.n61 two_stage_opamp_dummy_magic_0.Y.t49 996.134
R4349 two_stage_opamp_dummy_magic_0.Y.n62 two_stage_opamp_dummy_magic_0.Y.t36 996.134
R4350 two_stage_opamp_dummy_magic_0.Y.n63 two_stage_opamp_dummy_magic_0.Y.t51 996.134
R4351 two_stage_opamp_dummy_magic_0.Y.n67 two_stage_opamp_dummy_magic_0.Y.t44 996.134
R4352 two_stage_opamp_dummy_magic_0.Y.n66 two_stage_opamp_dummy_magic_0.Y.t31 996.134
R4353 two_stage_opamp_dummy_magic_0.Y.n65 two_stage_opamp_dummy_magic_0.Y.t46 996.134
R4354 two_stage_opamp_dummy_magic_0.Y.n64 two_stage_opamp_dummy_magic_0.Y.t40 996.134
R4355 two_stage_opamp_dummy_magic_0.Y.n53 two_stage_opamp_dummy_magic_0.Y.t53 690.867
R4356 two_stage_opamp_dummy_magic_0.Y.n50 two_stage_opamp_dummy_magic_0.Y.t29 690.867
R4357 two_stage_opamp_dummy_magic_0.Y.n42 two_stage_opamp_dummy_magic_0.Y.t37 530.201
R4358 two_stage_opamp_dummy_magic_0.Y.n45 two_stage_opamp_dummy_magic_0.Y.t30 530.201
R4359 two_stage_opamp_dummy_magic_0.Y.n57 two_stage_opamp_dummy_magic_0.Y.t54 514.134
R4360 two_stage_opamp_dummy_magic_0.Y.n53 two_stage_opamp_dummy_magic_0.Y.t38 514.134
R4361 two_stage_opamp_dummy_magic_0.Y.n54 two_stage_opamp_dummy_magic_0.Y.t42 514.134
R4362 two_stage_opamp_dummy_magic_0.Y.n55 two_stage_opamp_dummy_magic_0.Y.t27 514.134
R4363 two_stage_opamp_dummy_magic_0.Y.n56 two_stage_opamp_dummy_magic_0.Y.t41 514.134
R4364 two_stage_opamp_dummy_magic_0.Y.n52 two_stage_opamp_dummy_magic_0.Y.t48 514.134
R4365 two_stage_opamp_dummy_magic_0.Y.n51 two_stage_opamp_dummy_magic_0.Y.t33 514.134
R4366 two_stage_opamp_dummy_magic_0.Y.n50 two_stage_opamp_dummy_magic_0.Y.t45 514.134
R4367 two_stage_opamp_dummy_magic_0.Y.n58 two_stage_opamp_dummy_magic_0.Y.n49 473.967
R4368 two_stage_opamp_dummy_magic_0.Y.n69 two_stage_opamp_dummy_magic_0.Y.n68 446.967
R4369 two_stage_opamp_dummy_magic_0.Y.n58 two_stage_opamp_dummy_magic_0.Y.n57 441.834
R4370 two_stage_opamp_dummy_magic_0.Y.n49 two_stage_opamp_dummy_magic_0.Y.t32 353.467
R4371 two_stage_opamp_dummy_magic_0.Y.n42 two_stage_opamp_dummy_magic_0.Y.t52 353.467
R4372 two_stage_opamp_dummy_magic_0.Y.n43 two_stage_opamp_dummy_magic_0.Y.t39 353.467
R4373 two_stage_opamp_dummy_magic_0.Y.n44 two_stage_opamp_dummy_magic_0.Y.t25 353.467
R4374 two_stage_opamp_dummy_magic_0.Y.n48 two_stage_opamp_dummy_magic_0.Y.t47 353.467
R4375 two_stage_opamp_dummy_magic_0.Y.n47 two_stage_opamp_dummy_magic_0.Y.t35 353.467
R4376 two_stage_opamp_dummy_magic_0.Y.n46 two_stage_opamp_dummy_magic_0.Y.t50 353.467
R4377 two_stage_opamp_dummy_magic_0.Y.n45 two_stage_opamp_dummy_magic_0.Y.t43 353.467
R4378 two_stage_opamp_dummy_magic_0.Y.n62 two_stage_opamp_dummy_magic_0.Y.n61 176.733
R4379 two_stage_opamp_dummy_magic_0.Y.n63 two_stage_opamp_dummy_magic_0.Y.n62 176.733
R4380 two_stage_opamp_dummy_magic_0.Y.n68 two_stage_opamp_dummy_magic_0.Y.n63 176.733
R4381 two_stage_opamp_dummy_magic_0.Y.n68 two_stage_opamp_dummy_magic_0.Y.n67 176.733
R4382 two_stage_opamp_dummy_magic_0.Y.n67 two_stage_opamp_dummy_magic_0.Y.n66 176.733
R4383 two_stage_opamp_dummy_magic_0.Y.n66 two_stage_opamp_dummy_magic_0.Y.n65 176.733
R4384 two_stage_opamp_dummy_magic_0.Y.n65 two_stage_opamp_dummy_magic_0.Y.n64 176.733
R4385 two_stage_opamp_dummy_magic_0.Y.n43 two_stage_opamp_dummy_magic_0.Y.n42 176.733
R4386 two_stage_opamp_dummy_magic_0.Y.n44 two_stage_opamp_dummy_magic_0.Y.n43 176.733
R4387 two_stage_opamp_dummy_magic_0.Y.n49 two_stage_opamp_dummy_magic_0.Y.n44 176.733
R4388 two_stage_opamp_dummy_magic_0.Y.n49 two_stage_opamp_dummy_magic_0.Y.n48 176.733
R4389 two_stage_opamp_dummy_magic_0.Y.n48 two_stage_opamp_dummy_magic_0.Y.n47 176.733
R4390 two_stage_opamp_dummy_magic_0.Y.n47 two_stage_opamp_dummy_magic_0.Y.n46 176.733
R4391 two_stage_opamp_dummy_magic_0.Y.n46 two_stage_opamp_dummy_magic_0.Y.n45 176.733
R4392 two_stage_opamp_dummy_magic_0.Y.n51 two_stage_opamp_dummy_magic_0.Y.n50 176.733
R4393 two_stage_opamp_dummy_magic_0.Y.n52 two_stage_opamp_dummy_magic_0.Y.n51 176.733
R4394 two_stage_opamp_dummy_magic_0.Y.n57 two_stage_opamp_dummy_magic_0.Y.n52 176.733
R4395 two_stage_opamp_dummy_magic_0.Y.n57 two_stage_opamp_dummy_magic_0.Y.n56 176.733
R4396 two_stage_opamp_dummy_magic_0.Y.n56 two_stage_opamp_dummy_magic_0.Y.n55 176.733
R4397 two_stage_opamp_dummy_magic_0.Y.n55 two_stage_opamp_dummy_magic_0.Y.n54 176.733
R4398 two_stage_opamp_dummy_magic_0.Y.n54 two_stage_opamp_dummy_magic_0.Y.n53 176.733
R4399 two_stage_opamp_dummy_magic_0.Y.n59 two_stage_opamp_dummy_magic_0.Y.n58 176.238
R4400 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.n23 66.0338
R4401 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.n26 66.0338
R4402 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.n29 66.0338
R4403 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.n33 66.0338
R4404 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.n36 66.0338
R4405 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n39 66.0338
R4406 two_stage_opamp_dummy_magic_0.Y.t23 two_stage_opamp_dummy_magic_0.Y.n69 49.9906
R4407 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.n0 49.3505
R4408 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.n5 49.3505
R4409 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.n8 49.3505
R4410 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.n11 49.3505
R4411 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.n3 49.3505
R4412 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.n16 49.3505
R4413 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t0 16.0005
R4414 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t24 16.0005
R4415 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.t20 16.0005
R4416 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.t9 16.0005
R4417 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.t4 16.0005
R4418 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.t15 16.0005
R4419 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t17 16.0005
R4420 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t1 16.0005
R4421 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.t12 16.0005
R4422 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.t21 16.0005
R4423 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.t11 16.0005
R4424 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.t10 16.0005
R4425 two_stage_opamp_dummy_magic_0.Y.n59 two_stage_opamp_dummy_magic_0.Y.n41 12.7193
R4426 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.t18 11.2576
R4427 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.t7 11.2576
R4428 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.t8 11.2576
R4429 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.t16 11.2576
R4430 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.t13 11.2576
R4431 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.t19 11.2576
R4432 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.t5 11.2576
R4433 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.t2 11.2576
R4434 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.t6 11.2576
R4435 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.t22 11.2576
R4436 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.t3 11.2576
R4437 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.t14 11.2576
R4438 two_stage_opamp_dummy_magic_0.Y.n60 two_stage_opamp_dummy_magic_0.Y.n20 10.6255
R4439 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.n24 6.10467
R4440 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n38 5.91717
R4441 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.n24 5.91717
R4442 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.n4 5.6255
R4443 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n6 5.6255
R4444 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.n27 5.47967
R4445 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.n30 5.47967
R4446 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.n32 5.47967
R4447 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.n21 5.47967
R4448 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.n40 5.47967
R4449 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.n4 5.438
R4450 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.n6 5.438
R4451 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.n25 5.29217
R4452 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.n22 5.29217
R4453 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.n34 5.29217
R4454 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.n37 5.29217
R4455 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n9 5.063
R4456 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.n12 5.063
R4457 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.n15 5.063
R4458 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.n1 5.063
R4459 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.n7 4.8755
R4460 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.n2 4.8755
R4461 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.n17 4.8755
R4462 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.n19 4.5005
R4463 two_stage_opamp_dummy_magic_0.Y.n60 two_stage_opamp_dummy_magic_0.Y.n59 4.5005
R4464 two_stage_opamp_dummy_magic_0.Y.n69 two_stage_opamp_dummy_magic_0.Y.n60 2.3755
R4465 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.n35 0.6255
R4466 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.n22 0.6255
R4467 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.n22 0.6255
R4468 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.n28 0.6255
R4469 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.n31 0.6255
R4470 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.n21 0.6255
R4471 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.n21 0.6255
R4472 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.n14 0.563
R4473 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.n18 0.563
R4474 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.n2 0.563
R4475 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.n2 0.563
R4476 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.n10 0.563
R4477 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.n13 0.563
R4478 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.n1 0.3755
R4479 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 297.151
R4480 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 297.151
R4481 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 297.151
R4482 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n26 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 123.067
R4483 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 118.861
R4484 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 118.861
R4485 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n18 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n17 118.861
R4486 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n21 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n20 118.861
R4487 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n24 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n23 118.861
R4488 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n26 42.063
R4489 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 39.4005
R4490 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 39.4005
R4491 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 39.4005
R4492 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 39.4005
R4493 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 39.4005
R4494 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 39.4005
R4495 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 19.7005
R4496 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 19.7005
R4497 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 19.7005
R4498 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 19.7005
R4499 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n17 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 19.7005
R4500 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n17 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 19.7005
R4501 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n20 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 19.7005
R4502 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n20 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 19.7005
R4503 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n23 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 19.7005
R4504 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n23 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 19.7005
R4505 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n26 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n25 6.2505
R4506 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 5.60467
R4507 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 5.588
R4508 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n24 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n22 5.54217
R4509 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 5.54217
R4510 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 5.32967
R4511 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 5.32967
R4512 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 5.063
R4513 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 5.04217
R4514 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n18 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n16 5.04217
R4515 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n21 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 5.04217
R4516 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n25 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n24 5.04217
R4517 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 5.0255
R4518 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 4.97967
R4519 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n19 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n18 4.97967
R4520 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n22 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n21 4.97967
R4521 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 4.76717
R4522 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 1.28175
R4523 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n22 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n19 0.563
R4524 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n19 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 0.563
R4525 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 0.563
R4526 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 0.563
R4527 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n25 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 0.563
R4528 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 0.5255
R4529 VDDA.n209 VDDA.t131 1231.74
R4530 VDDA.n230 VDDA.t110 1231.74
R4531 VDDA.n68 VDDA.t201 1231.74
R4532 VDDA.n89 VDDA.t92 1231.74
R4533 VDDA.t159 VDDA.n199 1095.3
R4534 VDDA.n200 VDDA.t174 1095.3
R4535 VDDA.n135 VDDA.t150 1095.3
R4536 VDDA.t138 VDDA.n134 1095.3
R4537 VDDA.n59 VDDA.t165 1095.3
R4538 VDDA.t177 VDDA.n58 1095.3
R4539 VDDA.n145 VDDA.t179 671.418
R4540 VDDA.n166 VDDA.t107 671.418
R4541 VDDA.n4 VDDA.t161 671.418
R4542 VDDA.n25 VDDA.t104 671.418
R4543 VDDA.t141 VDDA.n344 665.689
R4544 VDDA.n345 VDDA.t117 665.689
R4545 VDDA.t196 VDDA.n305 665.689
R4546 VDDA.n306 VDDA.t96 665.689
R4547 VDDA.n199 VDDA.t160 663.801
R4548 VDDA.n200 VDDA.t175 663.801
R4549 VDDA.n135 VDDA.t151 663.801
R4550 VDDA.n134 VDDA.t139 663.801
R4551 VDDA.n59 VDDA.t166 663.801
R4552 VDDA.n58 VDDA.t178 663.801
R4553 VDDA.n245 VDDA.t198 661.375
R4554 VDDA.n248 VDDA.t119 661.375
R4555 VDDA.t129 VDDA.n382 648.726
R4556 VDDA.n383 VDDA.t126 648.726
R4557 VDDA.t153 VDDA.n352 648.726
R4558 VDDA.n353 VDDA.t190 648.726
R4559 VDDA.t171 VDDA.n444 648.726
R4560 VDDA.n445 VDDA.t135 648.726
R4561 VDDA.t147 VDDA.n433 648.726
R4562 VDDA.n434 VDDA.t102 648.726
R4563 VDDA.t114 VDDA.n410 648.726
R4564 VDDA.n411 VDDA.t156 648.726
R4565 VDDA.n130 VDDA.n129 594.301
R4566 VDDA.n127 VDDA.n126 594.301
R4567 VDDA.n123 VDDA.n122 594.301
R4568 VDDA.n120 VDDA.n119 594.301
R4569 VDDA.n116 VDDA.n115 594.301
R4570 VDDA.n113 VDDA.n112 594.301
R4571 VDDA.n109 VDDA.n108 594.301
R4572 VDDA.n106 VDDA.n105 594.301
R4573 VDDA.n102 VDDA.n101 594.301
R4574 VDDA.n99 VDDA.n98 594.301
R4575 VDDA.n189 VDDA.t122 589.076
R4576 VDDA.n194 VDDA.t98 589.076
R4577 VDDA.n48 VDDA.t192 589.076
R4578 VDDA.n53 VDDA.t204 589.076
R4579 VDDA.t53 VDDA.t159 580.557
R4580 VDDA.t419 VDDA.t53 580.557
R4581 VDDA.t291 VDDA.t419 580.557
R4582 VDDA.t209 VDDA.t291 580.557
R4583 VDDA.t288 VDDA.t209 580.557
R4584 VDDA.t17 VDDA.t288 580.557
R4585 VDDA.t433 VDDA.t17 580.557
R4586 VDDA.t432 VDDA.t433 580.557
R4587 VDDA.t2 VDDA.t432 580.557
R4588 VDDA.t270 VDDA.t2 580.557
R4589 VDDA.t174 VDDA.t270 580.557
R4590 VDDA.t150 VDDA.t268 580.557
R4591 VDDA.t268 VDDA.t76 580.557
R4592 VDDA.t76 VDDA.t0 580.557
R4593 VDDA.t0 VDDA.t26 580.557
R4594 VDDA.t26 VDDA.t446 580.557
R4595 VDDA.t446 VDDA.t264 580.557
R4596 VDDA.t264 VDDA.t266 580.557
R4597 VDDA.t266 VDDA.t295 580.557
R4598 VDDA.t295 VDDA.t453 580.557
R4599 VDDA.t453 VDDA.t422 580.557
R4600 VDDA.t422 VDDA.t424 580.557
R4601 VDDA.t424 VDDA.t24 580.557
R4602 VDDA.t24 VDDA.t231 580.557
R4603 VDDA.t231 VDDA.t297 580.557
R4604 VDDA.t297 VDDA.t277 580.557
R4605 VDDA.t277 VDDA.t459 580.557
R4606 VDDA.t459 VDDA.t339 580.557
R4607 VDDA.t339 VDDA.t444 580.557
R4608 VDDA.t444 VDDA.t293 580.557
R4609 VDDA.t293 VDDA.t235 580.557
R4610 VDDA.t235 VDDA.t138 580.557
R4611 VDDA.t165 VDDA.t292 580.557
R4612 VDDA.t292 VDDA.t214 580.557
R4613 VDDA.t214 VDDA.t237 580.557
R4614 VDDA.t237 VDDA.t336 580.557
R4615 VDDA.t336 VDDA.t230 580.557
R4616 VDDA.t230 VDDA.t5 580.557
R4617 VDDA.t5 VDDA.t31 580.557
R4618 VDDA.t31 VDDA.t71 580.557
R4619 VDDA.t71 VDDA.t450 580.557
R4620 VDDA.t450 VDDA.t416 580.557
R4621 VDDA.t416 VDDA.t177 580.557
R4622 VDDA.n350 VDDA.t152 524.808
R4623 VDDA.n355 VDDA.t189 524.808
R4624 VDDA.n379 VDDA.t128 514.768
R4625 VDDA.n385 VDDA.t125 514.768
R4626 VDDA.n237 VDDA.t182 456.526
R4627 VDDA.n240 VDDA.t167 456.526
R4628 VDDA.n447 VDDA.t134 418.368
R4629 VDDA.n431 VDDA.t146 418.368
R4630 VDDA.n436 VDDA.t101 418.368
R4631 VDDA.n408 VDDA.t113 418.368
R4632 VDDA.t313 VDDA.t141 407.144
R4633 VDDA.t252 VDDA.t313 407.144
R4634 VDDA.t74 VDDA.t252 407.144
R4635 VDDA.t434 VDDA.t74 407.144
R4636 VDDA.t18 VDDA.t434 407.144
R4637 VDDA.t355 VDDA.t18 407.144
R4638 VDDA.t303 VDDA.t355 407.144
R4639 VDDA.t254 VDDA.t303 407.144
R4640 VDDA.t273 VDDA.t254 407.144
R4641 VDDA.t451 VDDA.t273 407.144
R4642 VDDA.t420 VDDA.t451 407.144
R4643 VDDA.t357 VDDA.t420 407.144
R4644 VDDA.t372 VDDA.t357 407.144
R4645 VDDA.t72 VDDA.t372 407.144
R4646 VDDA.t271 VDDA.t72 407.144
R4647 VDDA.t463 VDDA.t271 407.144
R4648 VDDA.t233 VDDA.t463 407.144
R4649 VDDA.t315 VDDA.t233 407.144
R4650 VDDA.t117 VDDA.t315 407.144
R4651 VDDA.t56 VDDA.t196 407.144
R4652 VDDA.t286 VDDA.t56 407.144
R4653 VDDA.t12 VDDA.t286 407.144
R4654 VDDA.t90 VDDA.t12 407.144
R4655 VDDA.t86 VDDA.t90 407.144
R4656 VDDA.t67 VDDA.t86 407.144
R4657 VDDA.t317 VDDA.t67 407.144
R4658 VDDA.t284 VDDA.t317 407.144
R4659 VDDA.t37 VDDA.t284 407.144
R4660 VDDA.t58 VDDA.t37 407.144
R4661 VDDA.t348 VDDA.t58 407.144
R4662 VDDA.t84 VDDA.t348 407.144
R4663 VDDA.t369 VDDA.t84 407.144
R4664 VDDA.t65 VDDA.t369 407.144
R4665 VDDA.t417 VDDA.t65 407.144
R4666 VDDA.t60 VDDA.t417 407.144
R4667 VDDA.t88 VDDA.t60 407.144
R4668 VDDA.t69 VDDA.t88 407.144
R4669 VDDA.t96 VDDA.t69 407.144
R4670 VDDA.n442 VDDA.t170 399.623
R4671 VDDA.n413 VDDA.t155 399.623
R4672 VDDA.n239 VDDA.t168 397.784
R4673 VDDA.t183 VDDA.n238 397.784
R4674 VDDA.n342 VDDA.t140 382.217
R4675 VDDA.n347 VDDA.t116 382.217
R4676 VDDA.n303 VDDA.t195 382.217
R4677 VDDA.n308 VDDA.t95 382.217
R4678 VDDA.n376 VDDA.t143 374.668
R4679 VDDA.t275 VDDA.t129 373.214
R4680 VDDA.t22 VDDA.t275 373.214
R4681 VDDA.t126 VDDA.t22 373.214
R4682 VDDA.t305 VDDA.t153 373.214
R4683 VDDA.t52 VDDA.t305 373.214
R4684 VDDA.t190 VDDA.t52 373.214
R4685 VDDA.t455 VDDA.t171 373.214
R4686 VDDA.t256 VDDA.t455 373.214
R4687 VDDA.t440 VDDA.t256 373.214
R4688 VDDA.t258 VDDA.t440 373.214
R4689 VDDA.t135 VDDA.t258 373.214
R4690 VDDA.t436 VDDA.t147 373.214
R4691 VDDA.t212 VDDA.t436 373.214
R4692 VDDA.t299 VDDA.t212 373.214
R4693 VDDA.t20 VDDA.t299 373.214
R4694 VDDA.t219 VDDA.t20 373.214
R4695 VDDA.t438 VDDA.t219 373.214
R4696 VDDA.t217 VDDA.t438 373.214
R4697 VDDA.t262 VDDA.t217 373.214
R4698 VDDA.t457 VDDA.t262 373.214
R4699 VDDA.t319 VDDA.t457 373.214
R4700 VDDA.t102 VDDA.t319 373.214
R4701 VDDA.t337 VDDA.t114 373.214
R4702 VDDA.t260 VDDA.t337 373.214
R4703 VDDA.t210 VDDA.t260 373.214
R4704 VDDA.t442 VDDA.t210 373.214
R4705 VDDA.t156 VDDA.t442 373.214
R4706 VDDA.t144 VDDA.t145 371.774
R4707 VDDA.n358 VDDA.t186 370.168
R4708 VDDA.n197 VDDA.t158 348.075
R4709 VDDA.n202 VDDA.t173 348.075
R4710 VDDA.n132 VDDA.t137 348.075
R4711 VDDA.n92 VDDA.t149 348.075
R4712 VDDA.n56 VDDA.t176 348.075
R4713 VDDA.n61 VDDA.t164 348.075
R4714 VDDA.n192 VDDA.t99 343.882
R4715 VDDA.t123 VDDA.n191 343.882
R4716 VDDA.t193 VDDA.n50 343.882
R4717 VDDA.n51 VDDA.t205 343.882
R4718 VDDA.n344 VDDA.t142 331.901
R4719 VDDA.n345 VDDA.t118 331.901
R4720 VDDA.n305 VDDA.t197 331.901
R4721 VDDA.n306 VDDA.t97 331.901
R4722 VDDA.n382 VDDA.t130 331.901
R4723 VDDA.n383 VDDA.t127 331.901
R4724 VDDA.n352 VDDA.t154 331.901
R4725 VDDA.n353 VDDA.t191 331.901
R4726 VDDA.n444 VDDA.t172 331.901
R4727 VDDA.n445 VDDA.t136 331.901
R4728 VDDA.n433 VDDA.t148 331.901
R4729 VDDA.n434 VDDA.t103 331.901
R4730 VDDA.n410 VDDA.t115 331.901
R4731 VDDA.n411 VDDA.t157 331.901
R4732 VDDA.n339 VDDA.n338 297.151
R4733 VDDA.n336 VDDA.n335 297.151
R4734 VDDA.n332 VDDA.n331 297.151
R4735 VDDA.n329 VDDA.n328 297.151
R4736 VDDA.n325 VDDA.n324 297.151
R4737 VDDA.n322 VDDA.n321 297.151
R4738 VDDA.n318 VDDA.n317 297.151
R4739 VDDA.n315 VDDA.n314 297.151
R4740 VDDA.n264 VDDA.n263 297.151
R4741 VDDA.n301 VDDA.n300 297.151
R4742 VDDA.n298 VDDA.n297 297.151
R4743 VDDA.n294 VDDA.n293 297.151
R4744 VDDA.n291 VDDA.n290 297.151
R4745 VDDA.n287 VDDA.n286 297.151
R4746 VDDA.n284 VDDA.n283 297.151
R4747 VDDA.n280 VDDA.n279 297.151
R4748 VDDA.n277 VDDA.n276 297.151
R4749 VDDA.n269 VDDA.n268 297.151
R4750 VDDA.n378 VDDA.n377 297.151
R4751 VDDA.n439 VDDA.n438 297.151
R4752 VDDA.n392 VDDA.n391 297.151
R4753 VDDA.n428 VDDA.n427 297.151
R4754 VDDA.n425 VDDA.n424 297.151
R4755 VDDA.n421 VDDA.n420 297.151
R4756 VDDA.n418 VDDA.n417 297.151
R4757 VDDA.n397 VDDA.n396 297.151
R4758 VDDA.n406 VDDA.n405 297.151
R4759 VDDA.n402 VDDA.n401 297.151
R4760 VDDA.n357 VDDA.t187 285.517
R4761 VDDA.t168 VDDA.t241 259.091
R4762 VDDA.t241 VDDA.t183 259.091
R4763 VDDA.t187 VDDA.t309 251.471
R4764 VDDA.t309 VDDA.t311 251.471
R4765 VDDA.t311 VDDA.t250 251.471
R4766 VDDA.t250 VDDA.t228 251.471
R4767 VDDA.t228 VDDA.t45 251.471
R4768 VDDA.t45 VDDA.t225 251.471
R4769 VDDA.t225 VDDA.t32 251.471
R4770 VDDA.t32 VDDA.t9 251.471
R4771 VDDA.t9 VDDA.t43 251.471
R4772 VDDA.t43 VDDA.t81 251.471
R4773 VDDA.t81 VDDA.t243 251.471
R4774 VDDA.t243 VDDA.t248 251.471
R4775 VDDA.t248 VDDA.t352 251.471
R4776 VDDA.t352 VDDA.t307 251.471
R4777 VDDA.t307 VDDA.t329 251.471
R4778 VDDA.t329 VDDA.t39 251.471
R4779 VDDA.t39 VDDA.t144 251.471
R4780 VDDA.t99 VDDA.t399 217.708
R4781 VDDA.t399 VDDA.t379 217.708
R4782 VDDA.t379 VDDA.t398 217.708
R4783 VDDA.t398 VDDA.t415 217.708
R4784 VDDA.t415 VDDA.t405 217.708
R4785 VDDA.t405 VDDA.t387 217.708
R4786 VDDA.t387 VDDA.t402 217.708
R4787 VDDA.t402 VDDA.t383 217.708
R4788 VDDA.t383 VDDA.t394 217.708
R4789 VDDA.t394 VDDA.t409 217.708
R4790 VDDA.t409 VDDA.t123 217.708
R4791 VDDA.t222 VDDA.t193 217.708
R4792 VDDA.t428 VDDA.t222 217.708
R4793 VDDA.t80 VDDA.t428 217.708
R4794 VDDA.t363 VDDA.t80 217.708
R4795 VDDA.t221 VDDA.t363 217.708
R4796 VDDA.t281 VDDA.t221 217.708
R4797 VDDA.t78 VDDA.t281 217.708
R4798 VDDA.t36 VDDA.t78 217.708
R4799 VDDA.t79 VDDA.t36 217.708
R4800 VDDA.t62 VDDA.t79 217.708
R4801 VDDA.t205 VDDA.t62 217.708
R4802 VDDA.t199 VDDA.n246 213.131
R4803 VDDA.n247 VDDA.t120 213.131
R4804 VDDA.n164 VDDA.t108 213.131
R4805 VDDA.t180 VDDA.n163 213.131
R4806 VDDA.t162 VDDA.n22 213.131
R4807 VDDA.n23 VDDA.t105 213.131
R4808 VDDA.n258 VDDA.t471 169.55
R4809 VDDA.n239 VDDA.t169 168.139
R4810 VDDA.n238 VDDA.t185 168.139
R4811 VDDA.n260 VDDA.t470 165.8
R4812 VDDA.n259 VDDA.t472 165.8
R4813 VDDA.n258 VDDA.t469 165.8
R4814 VDDA.n236 VDDA.n235 153.576
R4815 VDDA.t14 VDDA.t199 146.155
R4816 VDDA.t120 VDDA.t14 146.155
R4817 VDDA.t108 VDDA.t448 146.155
R4818 VDDA.t448 VDDA.t346 146.155
R4819 VDDA.t346 VDDA.t301 146.155
R4820 VDDA.t301 VDDA.t344 146.155
R4821 VDDA.t344 VDDA.t359 146.155
R4822 VDDA.t359 VDDA.t3 146.155
R4823 VDDA.t3 VDDA.t367 146.155
R4824 VDDA.t367 VDDA.t7 146.155
R4825 VDDA.t7 VDDA.t342 146.155
R4826 VDDA.t342 VDDA.t461 146.155
R4827 VDDA.t461 VDDA.t180 146.155
R4828 VDDA.t215 VDDA.t162 146.155
R4829 VDDA.t467 VDDA.t215 146.155
R4830 VDDA.t365 VDDA.t467 146.155
R4831 VDDA.t426 VDDA.t365 146.155
R4832 VDDA.t29 VDDA.t426 146.155
R4833 VDDA.t465 VDDA.t29 146.155
R4834 VDDA.t289 VDDA.t465 146.155
R4835 VDDA.t279 VDDA.t289 146.155
R4836 VDDA.t374 VDDA.t279 146.155
R4837 VDDA.t207 VDDA.t374 146.155
R4838 VDDA.t105 VDDA.t207 146.155
R4839 VDDA.n192 VDDA.t100 136.701
R4840 VDDA.n191 VDDA.t124 136.701
R4841 VDDA.n50 VDDA.t194 136.701
R4842 VDDA.n51 VDDA.t206 136.701
R4843 VDDA.n228 VDDA.t111 122.829
R4844 VDDA.t132 VDDA.n227 122.829
R4845 VDDA.t202 VDDA.n86 122.829
R4846 VDDA.n87 VDDA.t93 122.829
R4847 VDDA.n357 VDDA.t188 86.2588
R4848 VDDA.t111 VDDA.t403 81.6411
R4849 VDDA.t403 VDDA.t384 81.6411
R4850 VDDA.t384 VDDA.t400 81.6411
R4851 VDDA.t400 VDDA.t380 81.6411
R4852 VDDA.t380 VDDA.t410 81.6411
R4853 VDDA.t410 VDDA.t392 81.6411
R4854 VDDA.t392 VDDA.t406 81.6411
R4855 VDDA.t406 VDDA.t388 81.6411
R4856 VDDA.t388 VDDA.t395 81.6411
R4857 VDDA.t395 VDDA.t413 81.6411
R4858 VDDA.t413 VDDA.t132 81.6411
R4859 VDDA.t361 VDDA.t202 81.6411
R4860 VDDA.t238 VDDA.t361 81.6411
R4861 VDDA.t325 VDDA.t238 81.6411
R4862 VDDA.t50 VDDA.t325 81.6411
R4863 VDDA.t54 VDDA.t50 81.6411
R4864 VDDA.t48 VDDA.t54 81.6411
R4865 VDDA.t321 VDDA.t48 81.6411
R4866 VDDA.t282 VDDA.t321 81.6411
R4867 VDDA.t323 VDDA.t282 81.6411
R4868 VDDA.t63 VDDA.t323 81.6411
R4869 VDDA.t93 VDDA.t63 81.6411
R4870 VDDA.n375 VDDA.n374 79.538
R4871 VDDA.n373 VDDA.n372 79.538
R4872 VDDA.n371 VDDA.n370 79.538
R4873 VDDA.n369 VDDA.n368 79.538
R4874 VDDA.n367 VDDA.n366 79.538
R4875 VDDA.n365 VDDA.n364 79.538
R4876 VDDA.n363 VDDA.n362 79.538
R4877 VDDA.n361 VDDA.n360 79.538
R4878 VDDA.n129 VDDA.t294 78.8005
R4879 VDDA.n129 VDDA.t236 78.8005
R4880 VDDA.n126 VDDA.t340 78.8005
R4881 VDDA.n126 VDDA.t445 78.8005
R4882 VDDA.n122 VDDA.t278 78.8005
R4883 VDDA.n122 VDDA.t460 78.8005
R4884 VDDA.n119 VDDA.t232 78.8005
R4885 VDDA.n119 VDDA.t298 78.8005
R4886 VDDA.n115 VDDA.t425 78.8005
R4887 VDDA.n115 VDDA.t25 78.8005
R4888 VDDA.n112 VDDA.t454 78.8005
R4889 VDDA.n112 VDDA.t423 78.8005
R4890 VDDA.n108 VDDA.t267 78.8005
R4891 VDDA.n108 VDDA.t296 78.8005
R4892 VDDA.n105 VDDA.t447 78.8005
R4893 VDDA.n105 VDDA.t265 78.8005
R4894 VDDA.n101 VDDA.t1 78.8005
R4895 VDDA.n101 VDDA.t27 78.8005
R4896 VDDA.n98 VDDA.t269 78.8005
R4897 VDDA.n98 VDDA.t77 78.8005
R4898 VDDA.n246 VDDA.t200 76.2576
R4899 VDDA.n247 VDDA.t121 76.2576
R4900 VDDA.n164 VDDA.t109 76.2576
R4901 VDDA.n163 VDDA.t181 76.2576
R4902 VDDA.n22 VDDA.t163 76.2576
R4903 VDDA.n23 VDDA.t106 76.2576
R4904 VDDA.n244 VDDA.n243 71.388
R4905 VDDA.n160 VDDA.n159 66.0338
R4906 VDDA.n156 VDDA.n155 66.0338
R4907 VDDA.n153 VDDA.n152 66.0338
R4908 VDDA.n149 VDDA.n148 66.0338
R4909 VDDA.n143 VDDA.n142 66.0338
R4910 VDDA.n19 VDDA.n18 66.0338
R4911 VDDA.n15 VDDA.n14 66.0338
R4912 VDDA.n12 VDDA.n11 66.0338
R4913 VDDA.n8 VDDA.n7 66.0338
R4914 VDDA.n2 VDDA.n1 66.0338
R4915 VDDA.n228 VDDA.t112 40.9789
R4916 VDDA.n227 VDDA.t133 40.9789
R4917 VDDA.n86 VDDA.t203 40.9789
R4918 VDDA.n87 VDDA.t94 40.9789
R4919 VDDA.n338 VDDA.t314 39.4005
R4920 VDDA.n338 VDDA.t253 39.4005
R4921 VDDA.n335 VDDA.t75 39.4005
R4922 VDDA.n335 VDDA.t435 39.4005
R4923 VDDA.n331 VDDA.t19 39.4005
R4924 VDDA.n331 VDDA.t356 39.4005
R4925 VDDA.n328 VDDA.t304 39.4005
R4926 VDDA.n328 VDDA.t255 39.4005
R4927 VDDA.n324 VDDA.t274 39.4005
R4928 VDDA.n324 VDDA.t452 39.4005
R4929 VDDA.n321 VDDA.t421 39.4005
R4930 VDDA.n321 VDDA.t358 39.4005
R4931 VDDA.n317 VDDA.t373 39.4005
R4932 VDDA.n317 VDDA.t73 39.4005
R4933 VDDA.n314 VDDA.t272 39.4005
R4934 VDDA.n314 VDDA.t464 39.4005
R4935 VDDA.n263 VDDA.t234 39.4005
R4936 VDDA.n263 VDDA.t316 39.4005
R4937 VDDA.n300 VDDA.t57 39.4005
R4938 VDDA.n300 VDDA.t287 39.4005
R4939 VDDA.n297 VDDA.t13 39.4005
R4940 VDDA.n297 VDDA.t91 39.4005
R4941 VDDA.n293 VDDA.t87 39.4005
R4942 VDDA.n293 VDDA.t68 39.4005
R4943 VDDA.n290 VDDA.t318 39.4005
R4944 VDDA.n290 VDDA.t285 39.4005
R4945 VDDA.n286 VDDA.t38 39.4005
R4946 VDDA.n286 VDDA.t59 39.4005
R4947 VDDA.n283 VDDA.t349 39.4005
R4948 VDDA.n283 VDDA.t85 39.4005
R4949 VDDA.n279 VDDA.t370 39.4005
R4950 VDDA.n279 VDDA.t66 39.4005
R4951 VDDA.n276 VDDA.t418 39.4005
R4952 VDDA.n276 VDDA.t61 39.4005
R4953 VDDA.n268 VDDA.t89 39.4005
R4954 VDDA.n268 VDDA.t70 39.4005
R4955 VDDA.n377 VDDA.t276 39.4005
R4956 VDDA.n377 VDDA.t23 39.4005
R4957 VDDA.n438 VDDA.t456 39.4005
R4958 VDDA.n438 VDDA.t257 39.4005
R4959 VDDA.n391 VDDA.t441 39.4005
R4960 VDDA.n391 VDDA.t259 39.4005
R4961 VDDA.n427 VDDA.t437 39.4005
R4962 VDDA.n427 VDDA.t213 39.4005
R4963 VDDA.n424 VDDA.t300 39.4005
R4964 VDDA.n424 VDDA.t21 39.4005
R4965 VDDA.n420 VDDA.t220 39.4005
R4966 VDDA.n420 VDDA.t439 39.4005
R4967 VDDA.n417 VDDA.t218 39.4005
R4968 VDDA.n417 VDDA.t263 39.4005
R4969 VDDA.n396 VDDA.t458 39.4005
R4970 VDDA.n396 VDDA.t320 39.4005
R4971 VDDA.n405 VDDA.t338 39.4005
R4972 VDDA.n405 VDDA.t261 39.4005
R4973 VDDA.n401 VDDA.t211 39.4005
R4974 VDDA.n401 VDDA.t443 39.4005
R4975 VDDA.n224 VDDA.n223 34.9935
R4976 VDDA.n220 VDDA.n219 34.9935
R4977 VDDA.n217 VDDA.n216 34.9935
R4978 VDDA.n213 VDDA.n212 34.9935
R4979 VDDA.n207 VDDA.n206 34.9935
R4980 VDDA.n83 VDDA.n82 34.9935
R4981 VDDA.n79 VDDA.n78 34.9935
R4982 VDDA.n76 VDDA.n75 34.9935
R4983 VDDA.n72 VDDA.n71 34.9935
R4984 VDDA.n66 VDDA.n65 34.9935
R4985 VDDA.n257 VDDA.n251 27.9413
R4986 VDDA.n171 VDDA.n170 24.288
R4987 VDDA.n174 VDDA.n173 24.288
R4988 VDDA.n177 VDDA.n176 24.288
R4989 VDDA.n181 VDDA.n180 24.288
R4990 VDDA.n184 VDDA.n183 24.288
R4991 VDDA.n187 VDDA.n186 24.288
R4992 VDDA.n30 VDDA.n29 24.288
R4993 VDDA.n33 VDDA.n32 24.288
R4994 VDDA.n36 VDDA.n35 24.288
R4995 VDDA.n40 VDDA.n39 24.288
R4996 VDDA.n43 VDDA.n42 24.288
R4997 VDDA.n46 VDDA.n45 24.288
R4998 VDDA.n235 VDDA.t242 21.8894
R4999 VDDA.n235 VDDA.t184 21.8894
R5000 VDDA.n251 VDDA.n250 20.1017
R5001 VDDA.n257 VDDA.t224 19.9244
R5002 VDDA.n193 VDDA.n190 14.8338
R5003 VDDA.n52 VDDA.n49 14.8338
R5004 VDDA.n201 VDDA.n198 14.0838
R5005 VDDA.n60 VDDA.n57 14.0838
R5006 VDDA.n374 VDDA.t330 13.1338
R5007 VDDA.n374 VDDA.t40 13.1338
R5008 VDDA.n372 VDDA.t353 13.1338
R5009 VDDA.n372 VDDA.t308 13.1338
R5010 VDDA.n370 VDDA.t244 13.1338
R5011 VDDA.n370 VDDA.t249 13.1338
R5012 VDDA.n368 VDDA.t44 13.1338
R5013 VDDA.n368 VDDA.t82 13.1338
R5014 VDDA.n366 VDDA.t33 13.1338
R5015 VDDA.n366 VDDA.t10 13.1338
R5016 VDDA.n364 VDDA.t46 13.1338
R5017 VDDA.n364 VDDA.t226 13.1338
R5018 VDDA.n362 VDDA.t251 13.1338
R5019 VDDA.n362 VDDA.t229 13.1338
R5020 VDDA.n360 VDDA.t310 13.1338
R5021 VDDA.n360 VDDA.t312 13.1338
R5022 VDDA.n196 VDDA.n188 11.9693
R5023 VDDA.n55 VDDA.n47 11.9693
R5024 VDDA.n449 VDDA.n448 11.4105
R5025 VDDA.n261 VDDA.n260 11.348
R5026 VDDA.t200 VDDA.n244 11.2576
R5027 VDDA.n244 VDDA.t15 11.2576
R5028 VDDA.n159 VDDA.t343 11.2576
R5029 VDDA.n159 VDDA.t462 11.2576
R5030 VDDA.n155 VDDA.t368 11.2576
R5031 VDDA.n155 VDDA.t8 11.2576
R5032 VDDA.n152 VDDA.t360 11.2576
R5033 VDDA.n152 VDDA.t4 11.2576
R5034 VDDA.n148 VDDA.t302 11.2576
R5035 VDDA.n148 VDDA.t345 11.2576
R5036 VDDA.n142 VDDA.t449 11.2576
R5037 VDDA.n142 VDDA.t347 11.2576
R5038 VDDA.n18 VDDA.t216 11.2576
R5039 VDDA.n18 VDDA.t468 11.2576
R5040 VDDA.n14 VDDA.t366 11.2576
R5041 VDDA.n14 VDDA.t427 11.2576
R5042 VDDA.n11 VDDA.t30 11.2576
R5043 VDDA.n11 VDDA.t466 11.2576
R5044 VDDA.n7 VDDA.t290 11.2576
R5045 VDDA.n7 VDDA.t280 11.2576
R5046 VDDA.n1 VDDA.t375 11.2576
R5047 VDDA.n1 VDDA.t208 11.2576
R5048 VDDA.n354 VDDA.n351 11.1672
R5049 VDDA.n389 VDDA.n388 9.7855
R5050 VDDA.n201 VDDA.n200 9.3005
R5051 VDDA.n199 VDDA.n198 9.3005
R5052 VDDA.n136 VDDA.n135 9.3005
R5053 VDDA.n134 VDDA.n133 9.3005
R5054 VDDA.n60 VDDA.n59 9.3005
R5055 VDDA.n58 VDDA.n57 9.3005
R5056 VDDA.n203 VDDA.n197 9.02133
R5057 VDDA.n62 VDDA.n56 9.02133
R5058 VDDA.n349 VDDA.n348 8.973
R5059 VDDA.n233 VDDA.n232 8.8755
R5060 VDDA.n140 VDDA.n139 8.8755
R5061 VDDA.n195 VDDA.n189 8.79217
R5062 VDDA.n54 VDDA.n48 8.79217
R5063 VDDA.n170 VDDA.t377 8.0005
R5064 VDDA.n170 VDDA.t335 8.0005
R5065 VDDA.n173 VDDA.t390 8.0005
R5066 VDDA.n173 VDDA.t397 8.0005
R5067 VDDA.n176 VDDA.t382 8.0005
R5068 VDDA.n176 VDDA.t412 8.0005
R5069 VDDA.n180 VDDA.t386 8.0005
R5070 VDDA.n180 VDDA.t378 8.0005
R5071 VDDA.n183 VDDA.t391 8.0005
R5072 VDDA.n183 VDDA.t376 8.0005
R5073 VDDA.n186 VDDA.t334 8.0005
R5074 VDDA.n186 VDDA.t408 8.0005
R5075 VDDA.n29 VDDA.t332 8.0005
R5076 VDDA.n29 VDDA.t341 8.0005
R5077 VDDA.n32 VDDA.t28 8.0005
R5078 VDDA.n32 VDDA.t6 8.0005
R5079 VDDA.n35 VDDA.t240 8.0005
R5080 VDDA.n35 VDDA.t223 8.0005
R5081 VDDA.n39 VDDA.t16 8.0005
R5082 VDDA.n39 VDDA.t431 8.0005
R5083 VDDA.n42 VDDA.t364 8.0005
R5084 VDDA.n42 VDDA.t429 8.0005
R5085 VDDA.n45 VDDA.t430 8.0005
R5086 VDDA.n45 VDDA.t333 8.0005
R5087 VDDA.n234 VDDA.n233 6.90675
R5088 VDDA.n234 VDDA.n140 6.90675
R5089 VDDA.n242 VDDA.n234 6.813
R5090 VDDA.n223 VDDA.t396 6.56717
R5091 VDDA.n223 VDDA.t414 6.56717
R5092 VDDA.n219 VDDA.t407 6.56717
R5093 VDDA.n219 VDDA.t389 6.56717
R5094 VDDA.n216 VDDA.t411 6.56717
R5095 VDDA.n216 VDDA.t393 6.56717
R5096 VDDA.n212 VDDA.t401 6.56717
R5097 VDDA.n212 VDDA.t381 6.56717
R5098 VDDA.n206 VDDA.t404 6.56717
R5099 VDDA.n206 VDDA.t385 6.56717
R5100 VDDA.n82 VDDA.t362 6.56717
R5101 VDDA.n82 VDDA.t239 6.56717
R5102 VDDA.n78 VDDA.t326 6.56717
R5103 VDDA.n78 VDDA.t51 6.56717
R5104 VDDA.n75 VDDA.t55 6.56717
R5105 VDDA.n75 VDDA.t49 6.56717
R5106 VDDA.n71 VDDA.t322 6.56717
R5107 VDDA.n71 VDDA.t283 6.56717
R5108 VDDA.n65 VDDA.t324 6.56717
R5109 VDDA.n65 VDDA.t64 6.56717
R5110 VDDA.n229 VDDA.n208 6.563
R5111 VDDA.n226 VDDA.n225 6.563
R5112 VDDA.n88 VDDA.n67 6.563
R5113 VDDA.n85 VDDA.n84 6.563
R5114 VDDA.n224 VDDA.n222 6.20883
R5115 VDDA.n221 VDDA.n220 6.20883
R5116 VDDA.n218 VDDA.n217 6.20883
R5117 VDDA.n213 VDDA.n211 6.20883
R5118 VDDA.n207 VDDA.n205 6.20883
R5119 VDDA.n83 VDDA.n81 6.20883
R5120 VDDA.n80 VDDA.n79 6.20883
R5121 VDDA.n77 VDDA.n76 6.20883
R5122 VDDA.n72 VDDA.n70 6.20883
R5123 VDDA.n66 VDDA.n64 6.20883
R5124 VDDA.n165 VDDA.n144 6.10467
R5125 VDDA.n162 VDDA.n161 6.10467
R5126 VDDA.n24 VDDA.n3 6.10467
R5127 VDDA.n21 VDDA.n20 6.10467
R5128 VDDA.n204 VDDA.n203 6.09425
R5129 VDDA.n63 VDDA.n62 6.09425
R5130 VDDA.n225 VDDA.n224 6.0005
R5131 VDDA.n220 VDDA.n210 6.0005
R5132 VDDA.n217 VDDA.n215 6.0005
R5133 VDDA.n214 VDDA.n213 6.0005
R5134 VDDA.n208 VDDA.n207 6.0005
R5135 VDDA.n84 VDDA.n83 6.0005
R5136 VDDA.n79 VDDA.n69 6.0005
R5137 VDDA.n76 VDDA.n74 6.0005
R5138 VDDA.n73 VDDA.n72 6.0005
R5139 VDDA.n67 VDDA.n66 6.0005
R5140 VDDA.n356 VDDA.n350 5.97967
R5141 VDDA.n187 VDDA.n185 5.938
R5142 VDDA.n172 VDDA.n171 5.938
R5143 VDDA.n175 VDDA.n171 5.938
R5144 VDDA.n46 VDDA.n44 5.938
R5145 VDDA.n31 VDDA.n30 5.938
R5146 VDDA.n34 VDDA.n30 5.938
R5147 VDDA.n346 VDDA.n265 5.85467
R5148 VDDA.n343 VDDA.n266 5.85467
R5149 VDDA.n307 VDDA.n270 5.85467
R5150 VDDA.n304 VDDA.n271 5.85467
R5151 VDDA.n160 VDDA.n158 5.813
R5152 VDDA.n157 VDDA.n156 5.813
R5153 VDDA.n154 VDDA.n153 5.813
R5154 VDDA.n149 VDDA.n147 5.813
R5155 VDDA.n143 VDDA.n141 5.813
R5156 VDDA.n19 VDDA.n17 5.813
R5157 VDDA.n16 VDDA.n15 5.813
R5158 VDDA.n13 VDDA.n12 5.813
R5159 VDDA.n8 VDDA.n6 5.813
R5160 VDDA.n2 VDDA.n0 5.813
R5161 VDDA.n133 VDDA.n93 5.60467
R5162 VDDA.n303 VDDA.n302 5.60467
R5163 VDDA.n158 VDDA.n145 5.563
R5164 VDDA.n17 VDDA.n4 5.563
R5165 VDDA.n435 VDDA.n398 5.52133
R5166 VDDA.n432 VDDA.n399 5.52133
R5167 VDDA.n446 VDDA.n393 5.51717
R5168 VDDA.n443 VDDA.n394 5.51717
R5169 VDDA.n412 VDDA.n403 5.51717
R5170 VDDA.n409 VDDA.n404 5.51717
R5171 VDDA.n161 VDDA.n160 5.47967
R5172 VDDA.n156 VDDA.n146 5.47967
R5173 VDDA.n153 VDDA.n151 5.47967
R5174 VDDA.n150 VDDA.n149 5.47967
R5175 VDDA.n144 VDDA.n143 5.47967
R5176 VDDA.n20 VDDA.n19 5.47967
R5177 VDDA.n15 VDDA.n5 5.47967
R5178 VDDA.n12 VDDA.n10 5.47967
R5179 VDDA.n9 VDDA.n8 5.47967
R5180 VDDA.n3 VDDA.n2 5.47967
R5181 VDDA.n222 VDDA.n209 5.3755
R5182 VDDA.n175 VDDA.n174 5.3755
R5183 VDDA.n174 VDDA.n172 5.3755
R5184 VDDA.n178 VDDA.n177 5.3755
R5185 VDDA.n177 VDDA.n169 5.3755
R5186 VDDA.n181 VDDA.n179 5.3755
R5187 VDDA.n182 VDDA.n181 5.3755
R5188 VDDA.n184 VDDA.n168 5.3755
R5189 VDDA.n185 VDDA.n184 5.3755
R5190 VDDA.n188 VDDA.n187 5.3755
R5191 VDDA.n81 VDDA.n68 5.3755
R5192 VDDA.n34 VDDA.n33 5.3755
R5193 VDDA.n33 VDDA.n31 5.3755
R5194 VDDA.n37 VDDA.n36 5.3755
R5195 VDDA.n36 VDDA.n28 5.3755
R5196 VDDA.n40 VDDA.n38 5.3755
R5197 VDDA.n41 VDDA.n40 5.3755
R5198 VDDA.n43 VDDA.n27 5.3755
R5199 VDDA.n44 VDDA.n43 5.3755
R5200 VDDA.n47 VDDA.n46 5.3755
R5201 VDDA.n100 VDDA.n92 5.35467
R5202 VDDA.n132 VDDA.n131 5.35467
R5203 VDDA.n340 VDDA.n339 5.35467
R5204 VDDA.n337 VDDA.n336 5.35467
R5205 VDDA.n332 VDDA.n310 5.35467
R5206 VDDA.n329 VDDA.n327 5.35467
R5207 VDDA.n326 VDDA.n325 5.35467
R5208 VDDA.n323 VDDA.n322 5.35467
R5209 VDDA.n318 VDDA.n312 5.35467
R5210 VDDA.n315 VDDA.n313 5.35467
R5211 VDDA.n264 VDDA.n262 5.35467
R5212 VDDA.n302 VDDA.n301 5.35467
R5213 VDDA.n299 VDDA.n298 5.35467
R5214 VDDA.n294 VDDA.n272 5.35467
R5215 VDDA.n291 VDDA.n289 5.35467
R5216 VDDA.n288 VDDA.n287 5.35467
R5217 VDDA.n285 VDDA.n284 5.35467
R5218 VDDA.n280 VDDA.n274 5.35467
R5219 VDDA.n277 VDDA.n275 5.35467
R5220 VDDA.n269 VDDA.n267 5.35467
R5221 VDDA.n384 VDDA.n380 5.33383
R5222 VDDA.n381 VDDA.n380 5.33383
R5223 VDDA.n250 VDDA.n249 5.28175
R5224 VDDA.n242 VDDA.n241 5.28175
R5225 VDDA.n232 VDDA.n231 5.28175
R5226 VDDA.n196 VDDA.n195 5.28175
R5227 VDDA.n55 VDDA.n54 5.28175
R5228 VDDA.n339 VDDA.n266 5.22967
R5229 VDDA.n336 VDDA.n334 5.22967
R5230 VDDA.n333 VDDA.n332 5.22967
R5231 VDDA.n330 VDDA.n329 5.22967
R5232 VDDA.n325 VDDA.n311 5.22967
R5233 VDDA.n322 VDDA.n320 5.22967
R5234 VDDA.n319 VDDA.n318 5.22967
R5235 VDDA.n316 VDDA.n315 5.22967
R5236 VDDA.n265 VDDA.n264 5.22967
R5237 VDDA.n301 VDDA.n271 5.22967
R5238 VDDA.n298 VDDA.n296 5.22967
R5239 VDDA.n295 VDDA.n294 5.22967
R5240 VDDA.n292 VDDA.n291 5.22967
R5241 VDDA.n287 VDDA.n273 5.22967
R5242 VDDA.n284 VDDA.n282 5.22967
R5243 VDDA.n281 VDDA.n280 5.22967
R5244 VDDA.n278 VDDA.n277 5.22967
R5245 VDDA.n270 VDDA.n269 5.22967
R5246 VDDA.n386 VDDA.n385 5.063
R5247 VDDA.n386 VDDA.n379 5.063
R5248 VDDA.n408 VDDA.n407 5.063
R5249 VDDA.n130 VDDA.n93 5.04217
R5250 VDDA.n131 VDDA.n130 5.04217
R5251 VDDA.n127 VDDA.n125 5.04217
R5252 VDDA.n128 VDDA.n127 5.04217
R5253 VDDA.n124 VDDA.n123 5.04217
R5254 VDDA.n123 VDDA.n94 5.04217
R5255 VDDA.n121 VDDA.n120 5.04217
R5256 VDDA.n120 VDDA.n118 5.04217
R5257 VDDA.n116 VDDA.n95 5.04217
R5258 VDDA.n117 VDDA.n116 5.04217
R5259 VDDA.n113 VDDA.n111 5.04217
R5260 VDDA.n114 VDDA.n113 5.04217
R5261 VDDA.n110 VDDA.n109 5.04217
R5262 VDDA.n109 VDDA.n96 5.04217
R5263 VDDA.n107 VDDA.n106 5.04217
R5264 VDDA.n106 VDDA.n104 5.04217
R5265 VDDA.n102 VDDA.n97 5.04217
R5266 VDDA.n103 VDDA.n102 5.04217
R5267 VDDA.n99 VDDA.n91 5.04217
R5268 VDDA.n100 VDDA.n99 5.04217
R5269 VDDA.n137 VDDA.n136 5.04217
R5270 VDDA.n203 VDDA.n202 5.02133
R5271 VDDA.n62 VDDA.n61 5.02133
R5272 VDDA.n348 VDDA.n347 4.97967
R5273 VDDA.n342 VDDA.n341 4.97967
R5274 VDDA.n309 VDDA.n308 4.97967
R5275 VDDA.n428 VDDA.n399 4.95883
R5276 VDDA.n425 VDDA.n423 4.95883
R5277 VDDA.n422 VDDA.n421 4.95883
R5278 VDDA.n419 VDDA.n418 4.95883
R5279 VDDA.n398 VDDA.n397 4.95883
R5280 VDDA.n439 VDDA.n394 4.95467
R5281 VDDA.n393 VDDA.n392 4.95467
R5282 VDDA.n406 VDDA.n404 4.95467
R5283 VDDA.n403 VDDA.n402 4.95467
R5284 VDDA.n167 VDDA.n166 4.938
R5285 VDDA.n26 VDDA.n25 4.938
R5286 VDDA.n440 VDDA.n439 4.838
R5287 VDDA.n392 VDDA.n390 4.838
R5288 VDDA.n407 VDDA.n406 4.838
R5289 VDDA.n402 VDDA.n400 4.838
R5290 VDDA.n429 VDDA.n428 4.83383
R5291 VDDA.n426 VDDA.n425 4.83383
R5292 VDDA.n421 VDDA.n415 4.83383
R5293 VDDA.n418 VDDA.n416 4.83383
R5294 VDDA.n397 VDDA.n395 4.83383
R5295 VDDA.n231 VDDA.n230 4.813
R5296 VDDA.n90 VDDA.n89 4.813
R5297 VDDA.n195 VDDA.n194 4.79217
R5298 VDDA.n54 VDDA.n53 4.79217
R5299 VDDA.n380 VDDA.n378 4.77133
R5300 VDDA.n245 VDDA.n243 4.7505
R5301 VDDA.n237 VDDA.n236 4.7505
R5302 VDDA.n388 VDDA.n387 4.7505
R5303 VDDA.n356 VDDA.n355 4.72967
R5304 VDDA.n346 VDDA.n345 4.6505
R5305 VDDA.n344 VDDA.n343 4.6505
R5306 VDDA.n307 VDDA.n306 4.6505
R5307 VDDA.n305 VDDA.n304 4.6505
R5308 VDDA.n384 VDDA.n383 4.6505
R5309 VDDA.n382 VDDA.n381 4.6505
R5310 VDDA.n354 VDDA.n353 4.6505
R5311 VDDA.n352 VDDA.n351 4.6505
R5312 VDDA.n446 VDDA.n445 4.6505
R5313 VDDA.n444 VDDA.n443 4.6505
R5314 VDDA.n435 VDDA.n434 4.6505
R5315 VDDA.n433 VDDA.n432 4.6505
R5316 VDDA.n412 VDDA.n411 4.6505
R5317 VDDA.n410 VDDA.n409 4.6505
R5318 VDDA.n249 VDDA.n248 4.5005
R5319 VDDA.n241 VDDA.n240 4.5005
R5320 VDDA.n139 VDDA.n138 4.5005
R5321 VDDA.n387 VDDA.n386 4.5005
R5322 VDDA.n359 VDDA.n358 4.5005
R5323 VDDA.n414 VDDA.n413 4.5005
R5324 VDDA.n431 VDDA.n430 4.5005
R5325 VDDA.n437 VDDA.n436 4.5005
R5326 VDDA.n442 VDDA.n441 4.5005
R5327 VDDA.n448 VDDA.n447 4.5005
R5328 VDDA.n261 VDDA.n257 4.38325
R5329 VDDA.n259 VDDA.n258 4.3755
R5330 VDDA.n232 VDDA.n204 4.15675
R5331 VDDA.n139 VDDA.n63 4.15675
R5332 VDDA.n260 VDDA.n259 3.7505
R5333 VDDA.n450 VDDA.n449 3.62787
R5334 VDDA.n138 VDDA.n137 3.1255
R5335 VDDA.n240 VDDA.n239 2.8255
R5336 VDDA.n238 VDDA.n237 2.8255
R5337 VDDA.n388 VDDA.n376 2.5005
R5338 VDDA.n450 VDDA.n251 2.1343
R5339 VDDA VDDA.n450 2.0779
R5340 VDDA.n358 VDDA.n357 1.913
R5341 VDDA.n248 VDDA.n247 1.888
R5342 VDDA.n246 VDDA.n245 1.888
R5343 VDDA.n341 VDDA.n309 1.8755
R5344 VDDA.n193 VDDA.n192 1.8605
R5345 VDDA.n191 VDDA.n190 1.8605
R5346 VDDA.n52 VDDA.n51 1.8605
R5347 VDDA.n50 VDDA.n49 1.8605
R5348 VDDA.n359 VDDA.n356 1.84425
R5349 VDDA.n430 VDDA.n414 1.813
R5350 VDDA.n441 VDDA.n437 1.813
R5351 VDDA.n204 VDDA.n196 1.438
R5352 VDDA.n63 VDDA.n55 1.438
R5353 VDDA.n230 VDDA.n229 1.39633
R5354 VDDA.n226 VDDA.n209 1.39633
R5355 VDDA.n89 VDDA.n88 1.39633
R5356 VDDA.n85 VDDA.n68 1.39633
R5357 VDDA.n349 VDDA.n261 1.06387
R5358 VDDA.n165 VDDA.n164 1.03383
R5359 VDDA.n163 VDDA.n162 1.03383
R5360 VDDA.n24 VDDA.n23 1.03383
R5361 VDDA.n22 VDDA.n21 1.03383
R5362 VDDA.n361 VDDA.n359 1.0005
R5363 VDDA.n363 VDDA.n361 1.0005
R5364 VDDA.n365 VDDA.n363 1.0005
R5365 VDDA.n367 VDDA.n365 1.0005
R5366 VDDA.n369 VDDA.n367 1.0005
R5367 VDDA.n371 VDDA.n369 1.0005
R5368 VDDA.n373 VDDA.n371 1.0005
R5369 VDDA.n375 VDDA.n373 1.0005
R5370 VDDA.n376 VDDA.n375 1.0005
R5371 VDDA.n250 VDDA.n242 0.938
R5372 VDDA.n166 VDDA.n165 0.8755
R5373 VDDA.n162 VDDA.n145 0.8755
R5374 VDDA.n25 VDDA.n24 0.8755
R5375 VDDA.n21 VDDA.n4 0.8755
R5376 VDDA.n138 VDDA.n90 0.78175
R5377 VDDA.n389 VDDA.n349 0.723125
R5378 VDDA.n249 VDDA.n243 0.6255
R5379 VDDA.n241 VDDA.n236 0.6255
R5380 VDDA.n150 VDDA.n144 0.6255
R5381 VDDA.n151 VDDA.n150 0.6255
R5382 VDDA.n151 VDDA.n146 0.6255
R5383 VDDA.n161 VDDA.n146 0.6255
R5384 VDDA.n158 VDDA.n157 0.6255
R5385 VDDA.n157 VDDA.n154 0.6255
R5386 VDDA.n154 VDDA.n147 0.6255
R5387 VDDA.n147 VDDA.n141 0.6255
R5388 VDDA.n167 VDDA.n141 0.6255
R5389 VDDA.n9 VDDA.n3 0.6255
R5390 VDDA.n10 VDDA.n9 0.6255
R5391 VDDA.n10 VDDA.n5 0.6255
R5392 VDDA.n20 VDDA.n5 0.6255
R5393 VDDA.n17 VDDA.n16 0.6255
R5394 VDDA.n16 VDDA.n13 0.6255
R5395 VDDA.n13 VDDA.n6 0.6255
R5396 VDDA.n6 VDDA.n0 0.6255
R5397 VDDA.n26 VDDA.n0 0.6255
R5398 VDDA.n316 VDDA.n265 0.6255
R5399 VDDA.n319 VDDA.n316 0.6255
R5400 VDDA.n320 VDDA.n319 0.6255
R5401 VDDA.n320 VDDA.n311 0.6255
R5402 VDDA.n330 VDDA.n311 0.6255
R5403 VDDA.n333 VDDA.n330 0.6255
R5404 VDDA.n334 VDDA.n333 0.6255
R5405 VDDA.n334 VDDA.n266 0.6255
R5406 VDDA.n278 VDDA.n270 0.6255
R5407 VDDA.n281 VDDA.n278 0.6255
R5408 VDDA.n282 VDDA.n281 0.6255
R5409 VDDA.n282 VDDA.n273 0.6255
R5410 VDDA.n292 VDDA.n273 0.6255
R5411 VDDA.n295 VDDA.n292 0.6255
R5412 VDDA.n296 VDDA.n295 0.6255
R5413 VDDA.n296 VDDA.n271 0.6255
R5414 VDDA.n302 VDDA.n299 0.6255
R5415 VDDA.n299 VDDA.n272 0.6255
R5416 VDDA.n289 VDDA.n272 0.6255
R5417 VDDA.n289 VDDA.n288 0.6255
R5418 VDDA.n288 VDDA.n285 0.6255
R5419 VDDA.n285 VDDA.n274 0.6255
R5420 VDDA.n275 VDDA.n274 0.6255
R5421 VDDA.n275 VDDA.n267 0.6255
R5422 VDDA.n309 VDDA.n267 0.6255
R5423 VDDA.n341 VDDA.n340 0.6255
R5424 VDDA.n340 VDDA.n337 0.6255
R5425 VDDA.n337 VDDA.n310 0.6255
R5426 VDDA.n327 VDDA.n310 0.6255
R5427 VDDA.n327 VDDA.n326 0.6255
R5428 VDDA.n326 VDDA.n323 0.6255
R5429 VDDA.n323 VDDA.n312 0.6255
R5430 VDDA.n313 VDDA.n312 0.6255
R5431 VDDA.n313 VDDA.n262 0.6255
R5432 VDDA.n348 VDDA.n262 0.6255
R5433 VDDA.n140 VDDA.n26 0.59425
R5434 VDDA.n229 VDDA.n228 0.58175
R5435 VDDA.n227 VDDA.n226 0.58175
R5436 VDDA.n88 VDDA.n87 0.58175
R5437 VDDA.n86 VDDA.n85 0.58175
R5438 VDDA.n214 VDDA.n208 0.563
R5439 VDDA.n215 VDDA.n214 0.563
R5440 VDDA.n215 VDDA.n210 0.563
R5441 VDDA.n225 VDDA.n210 0.563
R5442 VDDA.n222 VDDA.n221 0.563
R5443 VDDA.n221 VDDA.n218 0.563
R5444 VDDA.n218 VDDA.n211 0.563
R5445 VDDA.n211 VDDA.n205 0.563
R5446 VDDA.n231 VDDA.n205 0.563
R5447 VDDA.n194 VDDA.n193 0.563
R5448 VDDA.n190 VDDA.n189 0.563
R5449 VDDA.n185 VDDA.n182 0.563
R5450 VDDA.n182 VDDA.n169 0.563
R5451 VDDA.n172 VDDA.n169 0.563
R5452 VDDA.n178 VDDA.n175 0.563
R5453 VDDA.n179 VDDA.n178 0.563
R5454 VDDA.n179 VDDA.n168 0.563
R5455 VDDA.n188 VDDA.n168 0.563
R5456 VDDA.n233 VDDA.n167 0.563
R5457 VDDA.n103 VDDA.n100 0.563
R5458 VDDA.n104 VDDA.n103 0.563
R5459 VDDA.n104 VDDA.n96 0.563
R5460 VDDA.n114 VDDA.n96 0.563
R5461 VDDA.n117 VDDA.n114 0.563
R5462 VDDA.n118 VDDA.n117 0.563
R5463 VDDA.n118 VDDA.n94 0.563
R5464 VDDA.n128 VDDA.n94 0.563
R5465 VDDA.n131 VDDA.n128 0.563
R5466 VDDA.n125 VDDA.n93 0.563
R5467 VDDA.n125 VDDA.n124 0.563
R5468 VDDA.n124 VDDA.n121 0.563
R5469 VDDA.n121 VDDA.n95 0.563
R5470 VDDA.n111 VDDA.n95 0.563
R5471 VDDA.n111 VDDA.n110 0.563
R5472 VDDA.n110 VDDA.n107 0.563
R5473 VDDA.n107 VDDA.n97 0.563
R5474 VDDA.n97 VDDA.n91 0.563
R5475 VDDA.n137 VDDA.n91 0.563
R5476 VDDA.n73 VDDA.n67 0.563
R5477 VDDA.n74 VDDA.n73 0.563
R5478 VDDA.n74 VDDA.n69 0.563
R5479 VDDA.n84 VDDA.n69 0.563
R5480 VDDA.n81 VDDA.n80 0.563
R5481 VDDA.n80 VDDA.n77 0.563
R5482 VDDA.n77 VDDA.n70 0.563
R5483 VDDA.n70 VDDA.n64 0.563
R5484 VDDA.n90 VDDA.n64 0.563
R5485 VDDA.n53 VDDA.n52 0.563
R5486 VDDA.n49 VDDA.n48 0.563
R5487 VDDA.n44 VDDA.n41 0.563
R5488 VDDA.n41 VDDA.n28 0.563
R5489 VDDA.n31 VDDA.n28 0.563
R5490 VDDA.n37 VDDA.n34 0.563
R5491 VDDA.n38 VDDA.n37 0.563
R5492 VDDA.n38 VDDA.n27 0.563
R5493 VDDA.n47 VDDA.n27 0.563
R5494 VDDA.n394 VDDA.n393 0.563
R5495 VDDA.n419 VDDA.n398 0.563
R5496 VDDA.n422 VDDA.n419 0.563
R5497 VDDA.n423 VDDA.n422 0.563
R5498 VDDA.n423 VDDA.n399 0.563
R5499 VDDA.n404 VDDA.n403 0.563
R5500 VDDA.n407 VDDA.n400 0.563
R5501 VDDA.n414 VDDA.n400 0.563
R5502 VDDA.n430 VDDA.n429 0.563
R5503 VDDA.n429 VDDA.n426 0.563
R5504 VDDA.n426 VDDA.n415 0.563
R5505 VDDA.n416 VDDA.n415 0.563
R5506 VDDA.n416 VDDA.n395 0.563
R5507 VDDA.n437 VDDA.n395 0.563
R5508 VDDA.n441 VDDA.n440 0.563
R5509 VDDA.n440 VDDA.n390 0.563
R5510 VDDA.n448 VDDA.n390 0.563
R5511 VDDA.n355 VDDA.n354 0.479667
R5512 VDDA.n351 VDDA.n350 0.479667
R5513 VDDA VDDA.n389 0.464625
R5514 VDDA.n385 VDDA.n384 0.458833
R5515 VDDA.n381 VDDA.n379 0.458833
R5516 VDDA.n387 VDDA.n378 0.458833
R5517 VDDA.n347 VDDA.n346 0.3755
R5518 VDDA.n343 VDDA.n342 0.3755
R5519 VDDA.n308 VDDA.n307 0.3755
R5520 VDDA.n304 VDDA.n303 0.3755
R5521 VDDA.n447 VDDA.n446 0.338
R5522 VDDA.n443 VDDA.n442 0.338
R5523 VDDA.n413 VDDA.n412 0.338
R5524 VDDA.n409 VDDA.n408 0.338
R5525 VDDA.n436 VDDA.n435 0.333833
R5526 VDDA.n432 VDDA.n431 0.333833
R5527 VDDA.n202 VDDA.n201 0.2505
R5528 VDDA.n198 VDDA.n197 0.2505
R5529 VDDA.n136 VDDA.n92 0.2505
R5530 VDDA.n133 VDDA.n132 0.2505
R5531 VDDA.n61 VDDA.n60 0.2505
R5532 VDDA.n57 VDDA.n56 0.2505
R5533 VDDA.t306 VDDA.t331 0.1603
R5534 VDDA.t350 VDDA.t35 0.1603
R5535 VDDA.t371 VDDA.t327 0.1603
R5536 VDDA.t351 VDDA.t247 0.1603
R5537 VDDA.t11 VDDA.t354 0.1603
R5538 VDDA.n253 VDDA.t227 0.159278
R5539 VDDA.n254 VDDA.t47 0.159278
R5540 VDDA.n255 VDDA.t34 0.159278
R5541 VDDA.n256 VDDA.t246 0.159278
R5542 VDDA.n256 VDDA.t41 0.1368
R5543 VDDA.n256 VDDA.t306 0.1368
R5544 VDDA.n255 VDDA.t328 0.1368
R5545 VDDA.n255 VDDA.t350 0.1368
R5546 VDDA.n254 VDDA.t245 0.1368
R5547 VDDA.n254 VDDA.t371 0.1368
R5548 VDDA.n253 VDDA.t83 0.1368
R5549 VDDA.n253 VDDA.t351 0.1368
R5550 VDDA.n252 VDDA.t42 0.1368
R5551 VDDA.n252 VDDA.t11 0.1368
R5552 VDDA.n449 VDDA 0.135625
R5553 VDDA.t227 VDDA.n252 0.00152174
R5554 VDDA.t47 VDDA.n253 0.00152174
R5555 VDDA.t34 VDDA.n254 0.00152174
R5556 VDDA.t246 VDDA.n255 0.00152174
R5557 VDDA.t224 VDDA.n256 0.00152174
R5558 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 594.301
R5559 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 594.301
R5560 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 594.301
R5561 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 289.2
R5562 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 289.2
R5563 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 194.3
R5564 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.n24 194.3
R5565 two_stage_opamp_dummy_magic_0.err_amp_mir.n26 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 194.3
R5566 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 176.733
R5567 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 176.733
R5568 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 176.733
R5569 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 176.733
R5570 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 176.733
R5571 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 161.3
R5572 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 161.3
R5573 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 112.468
R5574 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 112.468
R5575 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 112.468
R5576 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 112.468
R5577 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 112.468
R5578 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 112.468
R5579 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 112.468
R5580 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 112.468
R5581 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 78.8005
R5582 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 78.8005
R5583 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 78.8005
R5584 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 78.8005
R5585 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 78.8005
R5586 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 78.8005
R5587 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 48.0005
R5588 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 48.0005
R5589 two_stage_opamp_dummy_magic_0.err_amp_mir.n24 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 48.0005
R5590 two_stage_opamp_dummy_magic_0.err_amp_mir.n24 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 48.0005
R5591 two_stage_opamp_dummy_magic_0.err_amp_mir.n26 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 48.0005
R5592 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 two_stage_opamp_dummy_magic_0.err_amp_mir.n26 48.0005
R5593 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 45.5227
R5594 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 45.5227
R5595 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 45.5227
R5596 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 45.5227
R5597 two_stage_opamp_dummy_magic_0.err_amp_mir.n22 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 6.60467
R5598 two_stage_opamp_dummy_magic_0.err_amp_mir.n25 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 6.39633
R5599 two_stage_opamp_dummy_magic_0.err_amp_mir.n25 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 6.39633
R5600 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 6.10467
R5601 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 6.10467
R5602 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.n23 5.97967
R5603 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 5.91717
R5604 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 5.91717
R5605 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.n25 5.14633
R5606 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 4.85467
R5607 two_stage_opamp_dummy_magic_0.err_amp_mir.n22 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 4.72967
R5608 two_stage_opamp_dummy_magic_0.err_amp_mir.n23 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 4.72967
R5609 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 4.66717
R5610 two_stage_opamp_dummy_magic_0.err_amp_mir.n23 two_stage_opamp_dummy_magic_0.err_amp_mir.n22 1.2505
R5611 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.t12 840.657
R5612 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.n1 601.072
R5613 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.n4 599.822
R5614 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.n2 599.822
R5615 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.n7 194.3
R5616 two_stage_opamp_dummy_magic_0.err_amp_out.n11 two_stage_opamp_dummy_magic_0.err_amp_out.n10 194.3
R5617 two_stage_opamp_dummy_magic_0.err_amp_out.n14 two_stage_opamp_dummy_magic_0.err_amp_out.n13 194.3
R5618 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.t0 78.8005
R5619 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.t11 78.8005
R5620 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.t5 78.8005
R5621 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.t2 78.8005
R5622 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t1 78.8005
R5623 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t3 78.8005
R5624 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.t9 48.0005
R5625 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.t6 48.0005
R5626 two_stage_opamp_dummy_magic_0.err_amp_out.n10 two_stage_opamp_dummy_magic_0.err_amp_out.t7 48.0005
R5627 two_stage_opamp_dummy_magic_0.err_amp_out.n10 two_stage_opamp_dummy_magic_0.err_amp_out.t4 48.0005
R5628 two_stage_opamp_dummy_magic_0.err_amp_out.n14 two_stage_opamp_dummy_magic_0.err_amp_out.t8 48.0005
R5629 two_stage_opamp_dummy_magic_0.err_amp_out.t10 two_stage_opamp_dummy_magic_0.err_amp_out.n14 48.0005
R5630 two_stage_opamp_dummy_magic_0.err_amp_out.n11 two_stage_opamp_dummy_magic_0.err_amp_out.n0 6.39633
R5631 two_stage_opamp_dummy_magic_0.err_amp_out.n12 two_stage_opamp_dummy_magic_0.err_amp_out.n11 6.20883
R5632 two_stage_opamp_dummy_magic_0.err_amp_out.n13 two_stage_opamp_dummy_magic_0.err_amp_out.n0 5.14633
R5633 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.n6 5.14633
R5634 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n8 4.95883
R5635 two_stage_opamp_dummy_magic_0.err_amp_out.n13 two_stage_opamp_dummy_magic_0.err_amp_out.n12 4.95883
R5636 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.n0 1.2505
R5637 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.n3 1.2505
R5638 two_stage_opamp_dummy_magic_0.err_amp_out.n12 two_stage_opamp_dummy_magic_0.err_amp_out.n9 1.2505
R5639 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.n5 1.063
R5640 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 610.534
R5641 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 610.534
R5642 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 433.8
R5643 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 433.8
R5644 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 433.8
R5645 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 433.8
R5646 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 433.8
R5647 two_stage_opamp_dummy_magic_0.V_tail_gate.n30 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 433.8
R5648 two_stage_opamp_dummy_magic_0.V_tail_gate.n31 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 433.8
R5649 two_stage_opamp_dummy_magic_0.V_tail_gate.n32 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 433.8
R5650 two_stage_opamp_dummy_magic_0.V_tail_gate.n33 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 433.8
R5651 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 433.8
R5652 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 433.8
R5653 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 433.8
R5654 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 433.8
R5655 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 433.8
R5656 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 433.8
R5657 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 433.8
R5658 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 433.8
R5659 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 433.8
R5660 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 297.151
R5661 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 297.151
R5662 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 297.151
R5663 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 297.151
R5664 two_stage_opamp_dummy_magic_0.V_tail_gate.n33 two_stage_opamp_dummy_magic_0.V_tail_gate.n32 176.733
R5665 two_stage_opamp_dummy_magic_0.V_tail_gate.n32 two_stage_opamp_dummy_magic_0.V_tail_gate.n31 176.733
R5666 two_stage_opamp_dummy_magic_0.V_tail_gate.n31 two_stage_opamp_dummy_magic_0.V_tail_gate.n30 176.733
R5667 two_stage_opamp_dummy_magic_0.V_tail_gate.n30 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 176.733
R5668 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 176.733
R5669 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 176.733
R5670 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 176.733
R5671 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 176.733
R5672 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 176.733
R5673 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 176.733
R5674 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 176.733
R5675 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 176.733
R5676 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 176.733
R5677 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 176.733
R5678 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 176.733
R5679 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 176.733
R5680 two_stage_opamp_dummy_magic_0.V_tail_gate.n35 two_stage_opamp_dummy_magic_0.V_tail_gate.n34 162.508
R5681 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_0.V_tail_gate 61.8443
R5682 two_stage_opamp_dummy_magic_0.V_tail_gate.n34 two_stage_opamp_dummy_magic_0.V_tail_gate.n33 56.2338
R5683 two_stage_opamp_dummy_magic_0.V_tail_gate.n34 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 56.2338
R5684 two_stage_opamp_dummy_magic_0.V_tail_gate.n37 two_stage_opamp_dummy_magic_0.V_tail_gate.n36 49.3505
R5685 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 49.3505
R5686 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 39.4005
R5687 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 39.4005
R5688 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 39.4005
R5689 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 39.4005
R5690 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 39.4005
R5691 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 39.4005
R5692 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 39.4005
R5693 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 39.4005
R5694 two_stage_opamp_dummy_magic_0.V_tail_gate.n36 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 16.0005
R5695 two_stage_opamp_dummy_magic_0.V_tail_gate.n36 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 16.0005
R5696 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 16.0005
R5697 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 16.0005
R5698 two_stage_opamp_dummy_magic_0.V_tail_gate.n37 two_stage_opamp_dummy_magic_0.V_tail_gate.n35 10.7922
R5699 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 5.96925
R5700 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 5.58383
R5701 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 5.58383
R5702 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 5.33383
R5703 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 5.33383
R5704 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 5.02133
R5705 two_stage_opamp_dummy_magic_0.V_tail_gate two_stage_opamp_dummy_magic_0.V_tail_gate.n13 4.82862
R5706 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 4.77133
R5707 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 4.77133
R5708 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 4.5005
R5709 two_stage_opamp_dummy_magic_0.V_tail_gate two_stage_opamp_dummy_magic_0.V_tail_gate.n12 1.28175
R5710 two_stage_opamp_dummy_magic_0.V_tail_gate.n35 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 1.22967
R5711 two_stage_opamp_dummy_magic_0.V_tail_gate two_stage_opamp_dummy_magic_0.V_tail_gate.n37 1.14112
R5712 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 0.563
R5713 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 0.563
R5714 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 0.521333
R5715 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.n0 97.1193
R5716 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t0 16.0005
R5717 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t3 16.0005
R5718 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.t1 9.6005
R5719 two_stage_opamp_dummy_magic_0.V_p_mir.t2 two_stage_opamp_dummy_magic_0.V_p_mir.n1 9.6005
R5720 two_stage_opamp_dummy_magic_0.VD2.n20 two_stage_opamp_dummy_magic_0.VD2.n19 49.3505
R5721 two_stage_opamp_dummy_magic_0.VD2.n23 two_stage_opamp_dummy_magic_0.VD2.n22 49.3505
R5722 two_stage_opamp_dummy_magic_0.VD2.n26 two_stage_opamp_dummy_magic_0.VD2.n25 49.3505
R5723 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.n3 49.3505
R5724 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.n7 49.3505
R5725 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.n9 49.3505
R5726 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.n5 49.3505
R5727 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.n14 49.3505
R5728 two_stage_opamp_dummy_magic_0.VD2.n35 two_stage_opamp_dummy_magic_0.VD2.n34 49.3505
R5729 two_stage_opamp_dummy_magic_0.VD2.n31 two_stage_opamp_dummy_magic_0.VD2.n30 49.3505
R5730 two_stage_opamp_dummy_magic_0.VD2.n29 two_stage_opamp_dummy_magic_0.VD2.n28 49.3505
R5731 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.t15 16.0005
R5732 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.t17 16.0005
R5733 two_stage_opamp_dummy_magic_0.VD2.n22 two_stage_opamp_dummy_magic_0.VD2.t4 16.0005
R5734 two_stage_opamp_dummy_magic_0.VD2.n22 two_stage_opamp_dummy_magic_0.VD2.t21 16.0005
R5735 two_stage_opamp_dummy_magic_0.VD2.n25 two_stage_opamp_dummy_magic_0.VD2.t18 16.0005
R5736 two_stage_opamp_dummy_magic_0.VD2.n25 two_stage_opamp_dummy_magic_0.VD2.t9 16.0005
R5737 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t3 16.0005
R5738 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t2 16.0005
R5739 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.t6 16.0005
R5740 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.t5 16.0005
R5741 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.t12 16.0005
R5742 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.t13 16.0005
R5743 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t7 16.0005
R5744 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t11 16.0005
R5745 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t20 16.0005
R5746 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t8 16.0005
R5747 two_stage_opamp_dummy_magic_0.VD2.n34 two_stage_opamp_dummy_magic_0.VD2.t1 16.0005
R5748 two_stage_opamp_dummy_magic_0.VD2.n34 two_stage_opamp_dummy_magic_0.VD2.t0 16.0005
R5749 two_stage_opamp_dummy_magic_0.VD2.n30 two_stage_opamp_dummy_magic_0.VD2.t10 16.0005
R5750 two_stage_opamp_dummy_magic_0.VD2.n30 two_stage_opamp_dummy_magic_0.VD2.t14 16.0005
R5751 two_stage_opamp_dummy_magic_0.VD2.n28 two_stage_opamp_dummy_magic_0.VD2.t19 16.0005
R5752 two_stage_opamp_dummy_magic_0.VD2.n28 two_stage_opamp_dummy_magic_0.VD2.t16 16.0005
R5753 two_stage_opamp_dummy_magic_0.VD2.n29 two_stage_opamp_dummy_magic_0.VD2.n18 5.64633
R5754 two_stage_opamp_dummy_magic_0.VD2.n21 two_stage_opamp_dummy_magic_0.VD2.n20 5.64633
R5755 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n6 5.6255
R5756 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n8 5.6255
R5757 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n6 5.438
R5758 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.n4 5.438
R5759 two_stage_opamp_dummy_magic_0.VD2.n24 two_stage_opamp_dummy_magic_0.VD2.n20 5.438
R5760 two_stage_opamp_dummy_magic_0.VD2.n32 two_stage_opamp_dummy_magic_0.VD2.n29 5.438
R5761 two_stage_opamp_dummy_magic_0.VD2.n23 two_stage_opamp_dummy_magic_0.VD2.n21 5.08383
R5762 two_stage_opamp_dummy_magic_0.VD2.n26 two_stage_opamp_dummy_magic_0.VD2.n2 5.08383
R5763 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.n35 5.08383
R5764 two_stage_opamp_dummy_magic_0.VD2.n31 two_stage_opamp_dummy_magic_0.VD2.n18 5.08383
R5765 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n10 5.063
R5766 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.n13 5.063
R5767 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.n0 5.063
R5768 two_stage_opamp_dummy_magic_0.VD2 two_stage_opamp_dummy_magic_0.VD2.n2 5.02133
R5769 two_stage_opamp_dummy_magic_0.VD2.n24 two_stage_opamp_dummy_magic_0.VD2.n23 4.8755
R5770 two_stage_opamp_dummy_magic_0.VD2.n27 two_stage_opamp_dummy_magic_0.VD2.n26 4.8755
R5771 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.n4 4.8755
R5772 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n15 4.8755
R5773 two_stage_opamp_dummy_magic_0.VD2.n35 two_stage_opamp_dummy_magic_0.VD2.n33 4.8755
R5774 two_stage_opamp_dummy_magic_0.VD2.n32 two_stage_opamp_dummy_magic_0.VD2.n31 4.8755
R5775 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.n17 4.5005
R5776 two_stage_opamp_dummy_magic_0.VD2 two_stage_opamp_dummy_magic_0.VD2.n0 1.1255
R5777 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n12 0.563
R5778 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.n16 0.563
R5779 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.n4 0.563
R5780 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.n11 0.563
R5781 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.n18 0.563
R5782 two_stage_opamp_dummy_magic_0.VD2.n21 two_stage_opamp_dummy_magic_0.VD2.n2 0.563
R5783 two_stage_opamp_dummy_magic_0.VD2.n27 two_stage_opamp_dummy_magic_0.VD2.n24 0.563
R5784 two_stage_opamp_dummy_magic_0.VD2.n33 two_stage_opamp_dummy_magic_0.VD2.n27 0.563
R5785 two_stage_opamp_dummy_magic_0.VD2.n33 two_stage_opamp_dummy_magic_0.VD2.n32 0.563
R5786 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.n1 0.46925
R5787 VOUT+.n9 VOUT+.t18 113.16
R5788 VOUT+.n11 VOUT+.n10 34.9935
R5789 VOUT+.n13 VOUT+.n12 34.9935
R5790 VOUT+.n17 VOUT+.n16 34.9935
R5791 VOUT+.n20 VOUT+.n19 34.9935
R5792 VOUT+.n23 VOUT+.n22 34.9935
R5793 VOUT+.n27 VOUT+.n26 34.9935
R5794 VOUT+.n110 VOUT+.n30 21.0005
R5795 VOUT+.n110 VOUT+.n109 11.6871
R5796 VOUT+ VOUT+.n110 9.90675
R5797 VOUT+.n2 VOUT+.n1 9.73997
R5798 VOUT+.n4 VOUT+.n3 9.73997
R5799 VOUT+.n7 VOUT+.n6 9.73997
R5800 VOUT+.n7 VOUT+.n5 7.14633
R5801 VOUT+.n5 VOUT+.n2 7.14633
R5802 VOUT+.n2 VOUT+.n0 7.14633
R5803 VOUT+.n10 VOUT+.t8 6.56717
R5804 VOUT+.n10 VOUT+.t12 6.56717
R5805 VOUT+.n12 VOUT+.t1 6.56717
R5806 VOUT+.n12 VOUT+.t13 6.56717
R5807 VOUT+.n16 VOUT+.t16 6.56717
R5808 VOUT+.n16 VOUT+.t2 6.56717
R5809 VOUT+.n19 VOUT+.t9 6.56717
R5810 VOUT+.n19 VOUT+.t11 6.56717
R5811 VOUT+.n22 VOUT+.t10 6.56717
R5812 VOUT+.n22 VOUT+.t14 6.56717
R5813 VOUT+.n26 VOUT+.t7 6.56717
R5814 VOUT+.n26 VOUT+.t15 6.56717
R5815 VOUT+.n21 VOUT+.n17 6.3755
R5816 VOUT+.n18 VOUT+.n17 6.3755
R5817 VOUT+.n29 VOUT+.n13 6.3755
R5818 VOUT+.n15 VOUT+.n13 6.3755
R5819 VOUT+.n4 VOUT+.n0 6.02133
R5820 VOUT+.n5 VOUT+.n4 6.02133
R5821 VOUT+.n8 VOUT+.n7 6.02133
R5822 VOUT+.n20 VOUT+.n18 5.813
R5823 VOUT+.n21 VOUT+.n20 5.813
R5824 VOUT+.n23 VOUT+.n14 5.813
R5825 VOUT+.n24 VOUT+.n23 5.813
R5826 VOUT+.n28 VOUT+.n27 5.813
R5827 VOUT+.n27 VOUT+.n25 5.813
R5828 VOUT+.n15 VOUT+.n11 5.813
R5829 VOUT+.n57 VOUT+.t85 4.8295
R5830 VOUT+.n59 VOUT+.t131 4.8295
R5831 VOUT+.n61 VOUT+.t31 4.8295
R5832 VOUT+.n63 VOUT+.t62 4.8295
R5833 VOUT+.n65 VOUT+.t114 4.8295
R5834 VOUT+.n77 VOUT+.t40 4.8295
R5835 VOUT+.n79 VOUT+.t34 4.8295
R5836 VOUT+.n80 VOUT+.t136 4.8295
R5837 VOUT+.n82 VOUT+.t70 4.8295
R5838 VOUT+.n83 VOUT+.t36 4.8295
R5839 VOUT+.n85 VOUT+.t95 4.8295
R5840 VOUT+.n86 VOUT+.t66 4.8295
R5841 VOUT+.n88 VOUT+.t55 4.8295
R5842 VOUT+.n89 VOUT+.t29 4.8295
R5843 VOUT+.n91 VOUT+.t91 4.8295
R5844 VOUT+.n92 VOUT+.t58 4.8295
R5845 VOUT+.n94 VOUT+.t49 4.8295
R5846 VOUT+.n95 VOUT+.t20 4.8295
R5847 VOUT+.n97 VOUT+.t148 4.8295
R5848 VOUT+.n98 VOUT+.t122 4.8295
R5849 VOUT+.n100 VOUT+.t44 4.8295
R5850 VOUT+.n101 VOUT+.t152 4.8295
R5851 VOUT+.n103 VOUT+.t142 4.8295
R5852 VOUT+.n104 VOUT+.t116 4.8295
R5853 VOUT+.n31 VOUT+.t108 4.8295
R5854 VOUT+.n43 VOUT+.t28 4.8295
R5855 VOUT+.n45 VOUT+.t24 4.8295
R5856 VOUT+.n46 VOUT+.t129 4.8295
R5857 VOUT+.n48 VOUT+.t61 4.8295
R5858 VOUT+.n49 VOUT+.t32 4.8295
R5859 VOUT+.n51 VOUT+.t100 4.8295
R5860 VOUT+.n52 VOUT+.t71 4.8295
R5861 VOUT+.n54 VOUT+.t69 4.8295
R5862 VOUT+.n55 VOUT+.t35 4.8295
R5863 VOUT+.n106 VOUT+.t77 4.8295
R5864 VOUT+.n70 VOUT+.t26 4.8154
R5865 VOUT+.n69 VOUT+.t59 4.8154
R5866 VOUT+.n68 VOUT+.t37 4.8154
R5867 VOUT+.n67 VOUT+.t81 4.8154
R5868 VOUT+.n76 VOUT+.t132 4.806
R5869 VOUT+.n75 VOUT+.t115 4.806
R5870 VOUT+.n74 VOUT+.t146 4.806
R5871 VOUT+.n73 VOUT+.t46 4.806
R5872 VOUT+.n72 VOUT+.t87 4.806
R5873 VOUT+.n71 VOUT+.t65 4.806
R5874 VOUT+.n70 VOUT+.t102 4.806
R5875 VOUT+.n69 VOUT+.t134 4.806
R5876 VOUT+.n68 VOUT+.t120 4.806
R5877 VOUT+.n67 VOUT+.t155 4.806
R5878 VOUT+.n42 VOUT+.t48 4.806
R5879 VOUT+.n41 VOUT+.t92 4.806
R5880 VOUT+.n40 VOUT+.t42 4.806
R5881 VOUT+.n39 VOUT+.t130 4.806
R5882 VOUT+.n38 VOUT+.t84 4.806
R5883 VOUT+.n37 VOUT+.t125 4.806
R5884 VOUT+.n36 VOUT+.t74 4.806
R5885 VOUT+.n35 VOUT+.t23 4.806
R5886 VOUT+.n34 VOUT+.t64 4.806
R5887 VOUT+.n33 VOUT+.t150 4.806
R5888 VOUT+.n58 VOUT+.t96 4.5005
R5889 VOUT+.n57 VOUT+.t57 4.5005
R5890 VOUT+.n59 VOUT+.t104 4.5005
R5891 VOUT+.n60 VOUT+.t73 4.5005
R5892 VOUT+.n61 VOUT+.t138 4.5005
R5893 VOUT+.n62 VOUT+.t107 4.5005
R5894 VOUT+.n63 VOUT+.t41 4.5005
R5895 VOUT+.n64 VOUT+.t143 4.5005
R5896 VOUT+.n65 VOUT+.t21 4.5005
R5897 VOUT+.n66 VOUT+.t126 4.5005
R5898 VOUT+.n67 VOUT+.t119 4.5005
R5899 VOUT+.n68 VOUT+.t82 4.5005
R5900 VOUT+.n69 VOUT+.t97 4.5005
R5901 VOUT+.n70 VOUT+.t63 4.5005
R5902 VOUT+.n71 VOUT+.t27 4.5005
R5903 VOUT+.n72 VOUT+.t45 4.5005
R5904 VOUT+.n73 VOUT+.t144 4.5005
R5905 VOUT+.n74 VOUT+.t112 4.5005
R5906 VOUT+.n75 VOUT+.t76 4.5005
R5907 VOUT+.n76 VOUT+.t93 4.5005
R5908 VOUT+.n78 VOUT+.t56 4.5005
R5909 VOUT+.n77 VOUT+.t19 4.5005
R5910 VOUT+.n79 VOUT+.t52 4.5005
R5911 VOUT+.n81 VOUT+.t156 4.5005
R5912 VOUT+.n80 VOUT+.t121 4.5005
R5913 VOUT+.n82 VOUT+.t89 4.5005
R5914 VOUT+.n84 VOUT+.t50 4.5005
R5915 VOUT+.n83 VOUT+.t151 4.5005
R5916 VOUT+.n85 VOUT+.t43 4.5005
R5917 VOUT+.n87 VOUT+.t145 4.5005
R5918 VOUT+.n86 VOUT+.t118 4.5005
R5919 VOUT+.n88 VOUT+.t141 4.5005
R5920 VOUT+.n90 VOUT+.t111 4.5005
R5921 VOUT+.n89 VOUT+.t80 4.5005
R5922 VOUT+.n91 VOUT+.t39 4.5005
R5923 VOUT+.n93 VOUT+.t139 4.5005
R5924 VOUT+.n92 VOUT+.t109 4.5005
R5925 VOUT+.n94 VOUT+.t135 4.5005
R5926 VOUT+.n96 VOUT+.t103 4.5005
R5927 VOUT+.n95 VOUT+.t72 4.5005
R5928 VOUT+.n97 VOUT+.t99 4.5005
R5929 VOUT+.n99 VOUT+.t68 4.5005
R5930 VOUT+.n98 VOUT+.t33 4.5005
R5931 VOUT+.n100 VOUT+.t133 4.5005
R5932 VOUT+.n102 VOUT+.t98 4.5005
R5933 VOUT+.n101 VOUT+.t67 4.5005
R5934 VOUT+.n103 VOUT+.t94 4.5005
R5935 VOUT+.n105 VOUT+.t60 4.5005
R5936 VOUT+.n104 VOUT+.t30 4.5005
R5937 VOUT+.n32 VOUT+.t101 4.5005
R5938 VOUT+.n31 VOUT+.t149 4.5005
R5939 VOUT+.n33 VOUT+.t88 4.5005
R5940 VOUT+.n34 VOUT+.t51 4.5005
R5941 VOUT+.n35 VOUT+.t137 4.5005
R5942 VOUT+.n36 VOUT+.t106 4.5005
R5943 VOUT+.n37 VOUT+.t75 4.5005
R5944 VOUT+.n38 VOUT+.t25 4.5005
R5945 VOUT+.n39 VOUT+.t128 4.5005
R5946 VOUT+.n40 VOUT+.t90 4.5005
R5947 VOUT+.n41 VOUT+.t54 4.5005
R5948 VOUT+.n42 VOUT+.t140 4.5005
R5949 VOUT+.n44 VOUT+.t110 4.5005
R5950 VOUT+.n43 VOUT+.t79 4.5005
R5951 VOUT+.n45 VOUT+.t113 4.5005
R5952 VOUT+.n47 VOUT+.t78 4.5005
R5953 VOUT+.n46 VOUT+.t38 4.5005
R5954 VOUT+.n48 VOUT+.t147 4.5005
R5955 VOUT+.n50 VOUT+.t117 4.5005
R5956 VOUT+.n49 VOUT+.t83 4.5005
R5957 VOUT+.n51 VOUT+.t47 4.5005
R5958 VOUT+.n53 VOUT+.t153 4.5005
R5959 VOUT+.n52 VOUT+.t123 4.5005
R5960 VOUT+.n54 VOUT+.t154 4.5005
R5961 VOUT+.n56 VOUT+.t124 4.5005
R5962 VOUT+.n55 VOUT+.t86 4.5005
R5963 VOUT+.n109 VOUT+.t105 4.5005
R5964 VOUT+.n108 VOUT+.t53 4.5005
R5965 VOUT+.n107 VOUT+.t22 4.5005
R5966 VOUT+.n106 VOUT+.t127 4.5005
R5967 VOUT+.n30 VOUT+.n29 4.5005
R5968 VOUT+.n1 VOUT+.t5 3.42907
R5969 VOUT+.n1 VOUT+.t17 3.42907
R5970 VOUT+.n3 VOUT+.t6 3.42907
R5971 VOUT+.n3 VOUT+.t3 3.42907
R5972 VOUT+.n6 VOUT+.t0 3.42907
R5973 VOUT+.n6 VOUT+.t4 3.42907
R5974 VOUT+ VOUT+.n9 1.84425
R5975 VOUT+.n9 VOUT+.n8 1.688
R5976 VOUT+.n30 VOUT+.n11 1.313
R5977 VOUT+.n8 VOUT+.n0 1.1255
R5978 VOUT+.n25 VOUT+.n15 0.563
R5979 VOUT+.n25 VOUT+.n24 0.563
R5980 VOUT+.n24 VOUT+.n21 0.563
R5981 VOUT+.n18 VOUT+.n14 0.563
R5982 VOUT+.n28 VOUT+.n14 0.563
R5983 VOUT+.n29 VOUT+.n28 0.563
R5984 VOUT+.n58 VOUT+.n57 0.3295
R5985 VOUT+.n60 VOUT+.n59 0.3295
R5986 VOUT+.n62 VOUT+.n61 0.3295
R5987 VOUT+.n64 VOUT+.n63 0.3295
R5988 VOUT+.n66 VOUT+.n65 0.3295
R5989 VOUT+.n68 VOUT+.n67 0.3295
R5990 VOUT+.n69 VOUT+.n68 0.3295
R5991 VOUT+.n70 VOUT+.n69 0.3295
R5992 VOUT+.n71 VOUT+.n70 0.3295
R5993 VOUT+.n72 VOUT+.n71 0.3295
R5994 VOUT+.n73 VOUT+.n72 0.3295
R5995 VOUT+.n74 VOUT+.n73 0.3295
R5996 VOUT+.n75 VOUT+.n74 0.3295
R5997 VOUT+.n76 VOUT+.n75 0.3295
R5998 VOUT+.n78 VOUT+.n76 0.3295
R5999 VOUT+.n78 VOUT+.n77 0.3295
R6000 VOUT+.n81 VOUT+.n79 0.3295
R6001 VOUT+.n81 VOUT+.n80 0.3295
R6002 VOUT+.n84 VOUT+.n82 0.3295
R6003 VOUT+.n84 VOUT+.n83 0.3295
R6004 VOUT+.n87 VOUT+.n85 0.3295
R6005 VOUT+.n87 VOUT+.n86 0.3295
R6006 VOUT+.n90 VOUT+.n88 0.3295
R6007 VOUT+.n90 VOUT+.n89 0.3295
R6008 VOUT+.n93 VOUT+.n91 0.3295
R6009 VOUT+.n93 VOUT+.n92 0.3295
R6010 VOUT+.n96 VOUT+.n94 0.3295
R6011 VOUT+.n96 VOUT+.n95 0.3295
R6012 VOUT+.n99 VOUT+.n97 0.3295
R6013 VOUT+.n99 VOUT+.n98 0.3295
R6014 VOUT+.n102 VOUT+.n100 0.3295
R6015 VOUT+.n102 VOUT+.n101 0.3295
R6016 VOUT+.n105 VOUT+.n103 0.3295
R6017 VOUT+.n105 VOUT+.n104 0.3295
R6018 VOUT+.n32 VOUT+.n31 0.3295
R6019 VOUT+.n34 VOUT+.n33 0.3295
R6020 VOUT+.n35 VOUT+.n34 0.3295
R6021 VOUT+.n36 VOUT+.n35 0.3295
R6022 VOUT+.n37 VOUT+.n36 0.3295
R6023 VOUT+.n38 VOUT+.n37 0.3295
R6024 VOUT+.n39 VOUT+.n38 0.3295
R6025 VOUT+.n40 VOUT+.n39 0.3295
R6026 VOUT+.n41 VOUT+.n40 0.3295
R6027 VOUT+.n42 VOUT+.n41 0.3295
R6028 VOUT+.n44 VOUT+.n42 0.3295
R6029 VOUT+.n44 VOUT+.n43 0.3295
R6030 VOUT+.n47 VOUT+.n45 0.3295
R6031 VOUT+.n47 VOUT+.n46 0.3295
R6032 VOUT+.n50 VOUT+.n48 0.3295
R6033 VOUT+.n50 VOUT+.n49 0.3295
R6034 VOUT+.n53 VOUT+.n51 0.3295
R6035 VOUT+.n53 VOUT+.n52 0.3295
R6036 VOUT+.n56 VOUT+.n54 0.3295
R6037 VOUT+.n56 VOUT+.n55 0.3295
R6038 VOUT+.n109 VOUT+.n108 0.3295
R6039 VOUT+.n108 VOUT+.n107 0.3295
R6040 VOUT+.n107 VOUT+.n106 0.3295
R6041 VOUT+.n74 VOUT+.n60 0.306
R6042 VOUT+.n73 VOUT+.n62 0.306
R6043 VOUT+.n72 VOUT+.n64 0.306
R6044 VOUT+.n71 VOUT+.n66 0.306
R6045 VOUT+.n78 VOUT+.n58 0.2825
R6046 VOUT+.n81 VOUT+.n78 0.2825
R6047 VOUT+.n84 VOUT+.n81 0.2825
R6048 VOUT+.n87 VOUT+.n84 0.2825
R6049 VOUT+.n90 VOUT+.n87 0.2825
R6050 VOUT+.n93 VOUT+.n90 0.2825
R6051 VOUT+.n96 VOUT+.n93 0.2825
R6052 VOUT+.n99 VOUT+.n96 0.2825
R6053 VOUT+.n102 VOUT+.n99 0.2825
R6054 VOUT+.n105 VOUT+.n102 0.2825
R6055 VOUT+.n44 VOUT+.n32 0.2825
R6056 VOUT+.n47 VOUT+.n44 0.2825
R6057 VOUT+.n50 VOUT+.n47 0.2825
R6058 VOUT+.n53 VOUT+.n50 0.2825
R6059 VOUT+.n56 VOUT+.n53 0.2825
R6060 VOUT+.n107 VOUT+.n56 0.2825
R6061 VOUT+.n107 VOUT+.n105 0.2825
R6062 two_stage_opamp_dummy_magic_0.cap_res_Y two_stage_opamp_dummy_magic_0.cap_res_Y.t138 49.2388
R6063 two_stage_opamp_dummy_magic_0.cap_res_Y two_stage_opamp_dummy_magic_0.cap_res_Y.t125 0.922875
R6064 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 0.1603
R6065 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 0.1603
R6066 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 0.1603
R6067 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 0.1603
R6068 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 0.1603
R6069 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 0.1603
R6070 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 0.1603
R6071 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 0.1603
R6072 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 0.1603
R6073 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 0.1603
R6074 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 0.1603
R6075 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 0.1603
R6076 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 0.1603
R6077 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 0.1603
R6078 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 0.1603
R6079 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 0.1603
R6080 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 0.1603
R6081 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 0.1603
R6082 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 0.1603
R6083 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 0.1603
R6084 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 0.1603
R6085 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 0.1603
R6086 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 0.1603
R6087 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 0.1603
R6088 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 0.1603
R6089 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 0.1603
R6090 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 0.1603
R6091 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 0.1603
R6092 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 0.1603
R6093 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 0.1603
R6094 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 0.1603
R6095 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 0.1603
R6096 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 0.1603
R6097 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 0.1603
R6098 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 0.1603
R6099 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 0.1603
R6100 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 0.1603
R6101 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 0.1603
R6102 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 0.1603
R6103 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 0.1603
R6104 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 0.1603
R6105 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 0.1603
R6106 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 0.1603
R6107 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 0.1603
R6108 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 0.1603
R6109 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 0.1603
R6110 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 0.1603
R6111 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 0.1603
R6112 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 0.1603
R6113 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 0.1603
R6114 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 0.1603
R6115 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 0.1603
R6116 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 0.1603
R6117 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 0.1603
R6118 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 0.1603
R6119 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 0.1603
R6120 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 0.1603
R6121 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 0.1603
R6122 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 0.159278
R6123 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 0.159278
R6124 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 0.159278
R6125 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 0.159278
R6126 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 0.159278
R6127 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 0.159278
R6128 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 0.159278
R6129 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 0.159278
R6130 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 0.159278
R6131 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 0.159278
R6132 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 0.159278
R6133 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 0.159278
R6134 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 0.159278
R6135 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 0.159278
R6136 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 0.159278
R6137 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 0.159278
R6138 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 0.159278
R6139 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 0.159278
R6140 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 0.159278
R6141 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 0.159278
R6142 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 0.159278
R6143 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 0.159278
R6144 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 0.159278
R6145 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 0.159278
R6146 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 0.159278
R6147 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 0.159278
R6148 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 0.159278
R6149 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 0.137822
R6150 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 0.1368
R6151 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 0.1368
R6152 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 0.1368
R6153 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 0.1368
R6154 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 0.1368
R6155 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 0.1368
R6156 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 0.1368
R6157 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 0.1368
R6158 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 0.1368
R6159 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 0.1368
R6160 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 0.1368
R6161 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 0.1368
R6162 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 0.1368
R6163 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 0.1368
R6164 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 0.1368
R6165 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 0.1368
R6166 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 0.1368
R6167 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 0.1368
R6168 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 0.1368
R6169 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 0.1368
R6170 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 0.1368
R6171 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 0.1368
R6172 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 0.1368
R6173 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 0.1368
R6174 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 0.1368
R6175 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 0.1368
R6176 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 0.1368
R6177 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 0.1368
R6178 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 0.1368
R6179 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 0.1368
R6180 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 0.1368
R6181 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 0.114322
R6182 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 0.1133
R6183 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 0.1133
R6184 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 0.1133
R6185 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 0.1133
R6186 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 0.1133
R6187 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 0.1133
R6188 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 0.1133
R6189 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 0.1133
R6190 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 0.1133
R6191 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 0.1133
R6192 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 0.1133
R6193 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 0.1133
R6194 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 0.1133
R6195 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 0.1133
R6196 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 0.1133
R6197 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 0.1133
R6198 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 0.1133
R6199 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 0.1133
R6200 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 0.1133
R6201 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 0.00152174
R6202 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 0.00152174
R6203 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 0.00152174
R6204 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 0.00152174
R6205 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 0.00152174
R6206 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 0.00152174
R6207 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 0.00152174
R6208 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 0.00152174
R6209 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 0.00152174
R6210 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 0.00152174
R6211 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 0.00152174
R6212 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 0.00152174
R6213 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 0.00152174
R6214 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 0.00152174
R6215 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 0.00152174
R6216 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 0.00152174
R6217 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 0.00152174
R6218 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 0.00152174
R6219 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 0.00152174
R6220 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 0.00152174
R6221 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 0.00152174
R6222 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 0.00152174
R6223 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 0.00152174
R6224 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 0.00152174
R6225 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 0.00152174
R6226 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 0.00152174
R6227 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 0.00152174
R6228 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 0.00152174
R6229 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 0.00152174
R6230 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 0.00152174
R6231 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 0.00152174
R6232 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 0.00152174
R6233 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 0.00152174
R6234 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 0.00152174
R6235 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 0.00152174
R6236 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 0.00152174
R6237 bgr_0.V_mir1.n17 bgr_0.V_mir1.t20 310.488
R6238 bgr_0.V_mir1.n8 bgr_0.V_mir1.t22 310.488
R6239 bgr_0.V_mir1.n14 bgr_0.V_mir1.t21 310.488
R6240 bgr_0.V_mir1.n13 bgr_0.V_mir1.n12 297.151
R6241 bgr_0.V_mir1.n24 bgr_0.V_mir1.n23 297.151
R6242 bgr_0.V_mir1.n27 bgr_0.V_mir1.n26 297.151
R6243 bgr_0.V_mir1.n2 bgr_0.V_mir1.t2 242.3
R6244 bgr_0.V_mir1.n1 bgr_0.V_mir1.n0 194.3
R6245 bgr_0.V_mir1.n5 bgr_0.V_mir1.n4 194.3
R6246 bgr_0.V_mir1.n19 bgr_0.V_mir1.t6 184.097
R6247 bgr_0.V_mir1.n10 bgr_0.V_mir1.t14 184.097
R6248 bgr_0.V_mir1.n16 bgr_0.V_mir1.t12 184.097
R6249 bgr_0.V_mir1.n18 bgr_0.V_mir1.n17 167.094
R6250 bgr_0.V_mir1.n9 bgr_0.V_mir1.n8 167.094
R6251 bgr_0.V_mir1.n15 bgr_0.V_mir1.n14 167.094
R6252 bgr_0.V_mir1.n20 bgr_0.V_mir1.n19 161.3
R6253 bgr_0.V_mir1.n11 bgr_0.V_mir1.n10 161.3
R6254 bgr_0.V_mir1.n22 bgr_0.V_mir1.n16 161.3
R6255 bgr_0.V_mir1.n17 bgr_0.V_mir1.t17 120.501
R6256 bgr_0.V_mir1.n18 bgr_0.V_mir1.t10 120.501
R6257 bgr_0.V_mir1.n8 bgr_0.V_mir1.t18 120.501
R6258 bgr_0.V_mir1.n9 bgr_0.V_mir1.t8 120.501
R6259 bgr_0.V_mir1.n14 bgr_0.V_mir1.t19 120.501
R6260 bgr_0.V_mir1.n15 bgr_0.V_mir1.t4 120.501
R6261 bgr_0.V_mir1.n0 bgr_0.V_mir1.t1 48.0005
R6262 bgr_0.V_mir1.n0 bgr_0.V_mir1.t0 48.0005
R6263 bgr_0.V_mir1.n4 bgr_0.V_mir1.t16 48.0005
R6264 bgr_0.V_mir1.n4 bgr_0.V_mir1.t3 48.0005
R6265 bgr_0.V_mir1.n19 bgr_0.V_mir1.n18 40.7027
R6266 bgr_0.V_mir1.n10 bgr_0.V_mir1.n9 40.7027
R6267 bgr_0.V_mir1.n16 bgr_0.V_mir1.n15 40.7027
R6268 bgr_0.V_mir1.n12 bgr_0.V_mir1.t7 39.4005
R6269 bgr_0.V_mir1.n12 bgr_0.V_mir1.t11 39.4005
R6270 bgr_0.V_mir1.n23 bgr_0.V_mir1.t13 39.4005
R6271 bgr_0.V_mir1.n23 bgr_0.V_mir1.t5 39.4005
R6272 bgr_0.V_mir1.t15 bgr_0.V_mir1.n27 39.4005
R6273 bgr_0.V_mir1.n27 bgr_0.V_mir1.t9 39.4005
R6274 bgr_0.V_mir1.n25 bgr_0.V_mir1.n24 6.89633
R6275 bgr_0.V_mir1.n25 bgr_0.V_mir1.n13 6.89633
R6276 bgr_0.V_mir1.n22 bgr_0.V_mir1.n21 6.6255
R6277 bgr_0.V_mir1.n21 bgr_0.V_mir1.n20 6.6255
R6278 bgr_0.V_mir1.n6 bgr_0.V_mir1.n2 6.22967
R6279 bgr_0.V_mir1.n3 bgr_0.V_mir1.n2 6.04217
R6280 bgr_0.V_mir1.n3 bgr_0.V_mir1.n1 6.04217
R6281 bgr_0.V_mir1.n7 bgr_0.V_mir1.n6 5.8755
R6282 bgr_0.V_mir1.n6 bgr_0.V_mir1.n5 4.85467
R6283 bgr_0.V_mir1.n26 bgr_0.V_mir1.n25 4.77133
R6284 bgr_0.V_mir1.n5 bgr_0.V_mir1.n3 4.66717
R6285 bgr_0.V_mir1.n21 bgr_0.V_mir1.n11 4.5005
R6286 bgr_0.V_mir1.n11 bgr_0.V_mir1.n7 1.7505
R6287 bgr_0.V_mir1.n7 bgr_0.V_mir1.n1 0.354667
R6288 bgr_0.V_mir1.n26 bgr_0.V_mir1.n11 0.333833
R6289 bgr_0.V_mir1.n24 bgr_0.V_mir1.n22 0.333833
R6290 bgr_0.V_mir1.n20 bgr_0.V_mir1.n13 0.333833
R6291 bgr_0.1st_Vout_1.n18 bgr_0.1st_Vout_1.t17 703.528
R6292 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t27 703.231
R6293 bgr_0.1st_Vout_1.n20 bgr_0.1st_Vout_1.n19 540.556
R6294 bgr_0.1st_Vout_1.n17 bgr_0.1st_Vout_1.n16 540.556
R6295 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.n8 297.151
R6296 bgr_0.1st_Vout_1.n24 bgr_0.1st_Vout_1.n23 297.151
R6297 bgr_0.1st_Vout_1.n27 bgr_0.1st_Vout_1.n26 297.151
R6298 bgr_0.1st_Vout_1.n19 bgr_0.1st_Vout_1.t13 291.209
R6299 bgr_0.1st_Vout_1.n16 bgr_0.1st_Vout_1.t15 291.209
R6300 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t7 242.3
R6301 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.n10 194.3
R6302 bgr_0.1st_Vout_1.n14 bgr_0.1st_Vout_1.n13 194.3
R6303 bgr_0.1st_Vout_1.n19 bgr_0.1st_Vout_1.t29 162.675
R6304 bgr_0.1st_Vout_1.n16 bgr_0.1st_Vout_1.t24 162.675
R6305 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.n4 53.7603
R6306 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t6 48.0005
R6307 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t10 48.0005
R6308 bgr_0.1st_Vout_1.n13 bgr_0.1st_Vout_1.t9 48.0005
R6309 bgr_0.1st_Vout_1.n13 bgr_0.1st_Vout_1.t8 48.0005
R6310 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t3 39.4005
R6311 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t1 39.4005
R6312 bgr_0.1st_Vout_1.n23 bgr_0.1st_Vout_1.t4 39.4005
R6313 bgr_0.1st_Vout_1.n23 bgr_0.1st_Vout_1.t0 39.4005
R6314 bgr_0.1st_Vout_1.t5 bgr_0.1st_Vout_1.n27 39.4005
R6315 bgr_0.1st_Vout_1.n27 bgr_0.1st_Vout_1.t2 39.4005
R6316 bgr_0.1st_Vout_1.n25 bgr_0.1st_Vout_1.n9 7.08383
R6317 bgr_0.1st_Vout_1.n26 bgr_0.1st_Vout_1.n25 7.08383
R6318 bgr_0.1st_Vout_1.n14 bgr_0.1st_Vout_1.n12 6.22967
R6319 bgr_0.1st_Vout_1.n12 bgr_0.1st_Vout_1.n11 6.22967
R6320 bgr_0.1st_Vout_1.n15 bgr_0.1st_Vout_1.n14 6.04217
R6321 bgr_0.1st_Vout_1.n15 bgr_0.1st_Vout_1.n11 6.04217
R6322 bgr_0.1st_Vout_1.n26 bgr_0.1st_Vout_1.n7 5.45883
R6323 bgr_0.1st_Vout_1.n18 bgr_0.1st_Vout_1.n9 5.45883
R6324 bgr_0.1st_Vout_1.n25 bgr_0.1st_Vout_1.n24 4.95883
R6325 bgr_0.1st_Vout_1.n12 bgr_0.1st_Vout_1.n5 4.85467
R6326 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t11 4.8295
R6327 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t31 4.8295
R6328 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t33 4.8295
R6329 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t21 4.8295
R6330 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t23 4.8295
R6331 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t14 4.8295
R6332 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t32 4.8295
R6333 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t19 4.8295
R6334 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t22 4.8295
R6335 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.n15 4.5005
R6336 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t16 4.5005
R6337 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t36 4.5005
R6338 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t35 4.5005
R6339 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t30 4.5005
R6340 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t28 4.5005
R6341 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t20 4.5005
R6342 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t34 4.5005
R6343 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t26 4.5005
R6344 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t25 4.5005
R6345 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t18 4.5005
R6346 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t12 4.5005
R6347 bgr_0.1st_Vout_1.n22 bgr_0.1st_Vout_1.n21 4.5005
R6348 bgr_0.1st_Vout_1.n22 bgr_0.1st_Vout_1.n5 1.26092
R6349 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.n6 1.04738
R6350 bgr_0.1st_Vout_1.n21 bgr_0.1st_Vout_1.n17 1.04738
R6351 bgr_0.1st_Vout_1.n20 bgr_0.1st_Vout_1.n18 1.04738
R6352 bgr_0.1st_Vout_1.n17 bgr_0.1st_Vout_1.n7 0.984875
R6353 bgr_0.1st_Vout_1.n21 bgr_0.1st_Vout_1.n20 0.984875
R6354 bgr_0.1st_Vout_1.n24 bgr_0.1st_Vout_1.n22 0.958833
R6355 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n2 0.8935
R6356 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.n0 0.8935
R6357 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.n3 0.6585
R6358 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.n1 0.6585
R6359 VOUT-.n110 VOUT-.t15 113.16
R6360 VOUT-.n1 VOUT-.n0 34.9935
R6361 VOUT-.n5 VOUT-.n4 34.9935
R6362 VOUT-.n7 VOUT-.n6 34.9935
R6363 VOUT-.n11 VOUT-.n10 34.9935
R6364 VOUT-.n14 VOUT-.n13 34.9935
R6365 VOUT-.n18 VOUT-.n17 34.9935
R6366 VOUT-.n100 VOUT-.n20 21.0005
R6367 VOUT-.n100 VOUT-.n99 11.6871
R6368 VOUT- VOUT-.n100 10.188
R6369 VOUT-.n103 VOUT-.n102 9.73997
R6370 VOUT-.n105 VOUT-.n104 9.73997
R6371 VOUT-.n108 VOUT-.n107 9.73997
R6372 VOUT-.n108 VOUT-.n106 7.14633
R6373 VOUT-.n106 VOUT-.n103 7.14633
R6374 VOUT-.n103 VOUT-.n101 7.14633
R6375 VOUT-.n0 VOUT-.t9 6.56717
R6376 VOUT-.n0 VOUT-.t11 6.56717
R6377 VOUT-.n4 VOUT-.t6 6.56717
R6378 VOUT-.n4 VOUT-.t16 6.56717
R6379 VOUT-.n6 VOUT-.t8 6.56717
R6380 VOUT-.n6 VOUT-.t12 6.56717
R6381 VOUT-.n10 VOUT-.t2 6.56717
R6382 VOUT-.n10 VOUT-.t3 6.56717
R6383 VOUT-.n13 VOUT-.t1 6.56717
R6384 VOUT-.n13 VOUT-.t10 6.56717
R6385 VOUT-.n17 VOUT-.t4 6.56717
R6386 VOUT-.n17 VOUT-.t5 6.56717
R6387 VOUT-.n18 VOUT-.n16 6.3755
R6388 VOUT-.n19 VOUT-.n18 6.3755
R6389 VOUT-.n8 VOUT-.n5 6.3755
R6390 VOUT-.n5 VOUT-.n3 6.3755
R6391 VOUT-.n105 VOUT-.n101 6.02133
R6392 VOUT-.n106 VOUT-.n105 6.02133
R6393 VOUT-.n109 VOUT-.n108 6.02133
R6394 VOUT-.n7 VOUT-.n3 5.813
R6395 VOUT-.n8 VOUT-.n7 5.813
R6396 VOUT-.n12 VOUT-.n11 5.813
R6397 VOUT-.n11 VOUT-.n9 5.813
R6398 VOUT-.n15 VOUT-.n14 5.813
R6399 VOUT-.n14 VOUT-.n2 5.813
R6400 VOUT-.n16 VOUT-.n1 5.813
R6401 VOUT-.n47 VOUT-.t108 4.8295
R6402 VOUT-.n56 VOUT-.t65 4.8295
R6403 VOUT-.n54 VOUT-.t118 4.8295
R6404 VOUT-.n52 VOUT-.t151 4.8295
R6405 VOUT-.n50 VOUT-.t44 4.8295
R6406 VOUT-.n49 VOUT-.t67 4.8295
R6407 VOUT-.n69 VOUT-.t27 4.8295
R6408 VOUT-.n70 VOUT-.t76 4.8295
R6409 VOUT-.n72 VOUT-.t62 4.8295
R6410 VOUT-.n73 VOUT-.t112 4.8295
R6411 VOUT-.n75 VOUT-.t114 4.8295
R6412 VOUT-.n76 VOUT-.t99 4.8295
R6413 VOUT-.n78 VOUT-.t74 4.8295
R6414 VOUT-.n79 VOUT-.t55 4.8295
R6415 VOUT-.n81 VOUT-.t109 4.8295
R6416 VOUT-.n82 VOUT-.t91 4.8295
R6417 VOUT-.n84 VOUT-.t68 4.8295
R6418 VOUT-.n85 VOUT-.t52 4.8295
R6419 VOUT-.n87 VOUT-.t29 4.8295
R6420 VOUT-.n88 VOUT-.t153 4.8295
R6421 VOUT-.n90 VOUT-.t63 4.8295
R6422 VOUT-.n91 VOUT-.t46 4.8295
R6423 VOUT-.n93 VOUT-.t22 4.8295
R6424 VOUT-.n94 VOUT-.t146 4.8295
R6425 VOUT-.n21 VOUT-.t117 4.8295
R6426 VOUT-.n23 VOUT-.t72 4.8295
R6427 VOUT-.n35 VOUT-.t37 4.8295
R6428 VOUT-.n36 VOUT-.t20 4.8295
R6429 VOUT-.n38 VOUT-.t79 4.8295
R6430 VOUT-.n39 VOUT-.t60 4.8295
R6431 VOUT-.n41 VOUT-.t121 4.8295
R6432 VOUT-.n42 VOUT-.t104 4.8295
R6433 VOUT-.n44 VOUT-.t84 4.8295
R6434 VOUT-.n45 VOUT-.t66 4.8295
R6435 VOUT-.n96 VOUT-.t123 4.8295
R6436 VOUT-.n58 VOUT-.t95 4.8154
R6437 VOUT-.n59 VOUT-.t70 4.8154
R6438 VOUT-.n60 VOUT-.t110 4.8154
R6439 VOUT-.n61 VOUT-.t145 4.8154
R6440 VOUT-.n58 VOUT-.t32 4.806
R6441 VOUT-.n59 VOUT-.t150 4.806
R6442 VOUT-.n60 VOUT-.t50 4.806
R6443 VOUT-.n61 VOUT-.t87 4.806
R6444 VOUT-.n62 VOUT-.t125 4.806
R6445 VOUT-.n63 VOUT-.t105 4.806
R6446 VOUT-.n64 VOUT-.t140 4.806
R6447 VOUT-.n65 VOUT-.t36 4.806
R6448 VOUT-.n66 VOUT-.t156 4.806
R6449 VOUT-.n67 VOUT-.t53 4.806
R6450 VOUT-.n24 VOUT-.t73 4.806
R6451 VOUT-.n25 VOUT-.t116 4.806
R6452 VOUT-.n26 VOUT-.t64 4.806
R6453 VOUT-.n27 VOUT-.t154 4.806
R6454 VOUT-.n28 VOUT-.t106 4.806
R6455 VOUT-.n29 VOUT-.t143 4.806
R6456 VOUT-.n30 VOUT-.t96 4.806
R6457 VOUT-.n31 VOUT-.t42 4.806
R6458 VOUT-.n32 VOUT-.t86 4.806
R6459 VOUT-.n33 VOUT-.t34 4.806
R6460 VOUT-.n47 VOUT-.t69 4.5005
R6461 VOUT-.n48 VOUT-.t90 4.5005
R6462 VOUT-.n56 VOUT-.t80 4.5005
R6463 VOUT-.n57 VOUT-.t43 4.5005
R6464 VOUT-.n54 VOUT-.t56 4.5005
R6465 VOUT-.n55 VOUT-.t21 4.5005
R6466 VOUT-.n52 VOUT-.t98 4.5005
R6467 VOUT-.n53 VOUT-.t59 4.5005
R6468 VOUT-.n50 VOUT-.t136 4.5005
R6469 VOUT-.n51 VOUT-.t101 4.5005
R6470 VOUT-.n49 VOUT-.t30 4.5005
R6471 VOUT-.n68 VOUT-.t51 4.5005
R6472 VOUT-.n67 VOUT-.t155 4.5005
R6473 VOUT-.n66 VOUT-.t119 4.5005
R6474 VOUT-.n65 VOUT-.t139 4.5005
R6475 VOUT-.n64 VOUT-.t102 4.5005
R6476 VOUT-.n63 VOUT-.t61 4.5005
R6477 VOUT-.n62 VOUT-.t85 4.5005
R6478 VOUT-.n61 VOUT-.t45 4.5005
R6479 VOUT-.n60 VOUT-.t147 4.5005
R6480 VOUT-.n59 VOUT-.t111 4.5005
R6481 VOUT-.n58 VOUT-.t134 4.5005
R6482 VOUT-.n69 VOUT-.t130 4.5005
R6483 VOUT-.n71 VOUT-.t152 4.5005
R6484 VOUT-.n70 VOUT-.t115 4.5005
R6485 VOUT-.n72 VOUT-.t23 4.5005
R6486 VOUT-.n74 VOUT-.t47 4.5005
R6487 VOUT-.n73 VOUT-.t148 4.5005
R6488 VOUT-.n75 VOUT-.t78 4.5005
R6489 VOUT-.n77 VOUT-.t26 4.5005
R6490 VOUT-.n76 VOUT-.t132 4.5005
R6491 VOUT-.n78 VOUT-.t39 4.5005
R6492 VOUT-.n80 VOUT-.t128 4.5005
R6493 VOUT-.n79 VOUT-.t92 4.5005
R6494 VOUT-.n81 VOUT-.t71 4.5005
R6495 VOUT-.n83 VOUT-.t19 4.5005
R6496 VOUT-.n82 VOUT-.t126 4.5005
R6497 VOUT-.n84 VOUT-.t33 4.5005
R6498 VOUT-.n86 VOUT-.t122 4.5005
R6499 VOUT-.n85 VOUT-.t88 4.5005
R6500 VOUT-.n87 VOUT-.t135 4.5005
R6501 VOUT-.n89 VOUT-.t82 4.5005
R6502 VOUT-.n88 VOUT-.t48 4.5005
R6503 VOUT-.n90 VOUT-.t28 4.5005
R6504 VOUT-.n92 VOUT-.t120 4.5005
R6505 VOUT-.n91 VOUT-.t81 4.5005
R6506 VOUT-.n93 VOUT-.t129 4.5005
R6507 VOUT-.n95 VOUT-.t77 4.5005
R6508 VOUT-.n94 VOUT-.t40 4.5005
R6509 VOUT-.n21 VOUT-.t25 4.5005
R6510 VOUT-.n22 VOUT-.t124 4.5005
R6511 VOUT-.n23 VOUT-.t38 4.5005
R6512 VOUT-.n34 VOUT-.t127 4.5005
R6513 VOUT-.n33 VOUT-.t94 4.5005
R6514 VOUT-.n32 VOUT-.t54 4.5005
R6515 VOUT-.n31 VOUT-.t144 4.5005
R6516 VOUT-.n30 VOUT-.t113 4.5005
R6517 VOUT-.n29 VOUT-.t75 4.5005
R6518 VOUT-.n28 VOUT-.t24 4.5005
R6519 VOUT-.n27 VOUT-.t131 4.5005
R6520 VOUT-.n26 VOUT-.t97 4.5005
R6521 VOUT-.n25 VOUT-.t58 4.5005
R6522 VOUT-.n24 VOUT-.t149 4.5005
R6523 VOUT-.n35 VOUT-.t142 4.5005
R6524 VOUT-.n37 VOUT-.t93 4.5005
R6525 VOUT-.n36 VOUT-.t57 4.5005
R6526 VOUT-.n38 VOUT-.t41 4.5005
R6527 VOUT-.n40 VOUT-.t133 4.5005
R6528 VOUT-.n39 VOUT-.t100 4.5005
R6529 VOUT-.n41 VOUT-.t83 4.5005
R6530 VOUT-.n43 VOUT-.t31 4.5005
R6531 VOUT-.n42 VOUT-.t137 4.5005
R6532 VOUT-.n44 VOUT-.t49 4.5005
R6533 VOUT-.n46 VOUT-.t138 4.5005
R6534 VOUT-.n45 VOUT-.t103 4.5005
R6535 VOUT-.n96 VOUT-.t89 4.5005
R6536 VOUT-.n97 VOUT-.t35 4.5005
R6537 VOUT-.n98 VOUT-.t141 4.5005
R6538 VOUT-.n99 VOUT-.t107 4.5005
R6539 VOUT-.n20 VOUT-.n19 4.5005
R6540 VOUT-.n102 VOUT-.t7 3.42907
R6541 VOUT-.n102 VOUT-.t13 3.42907
R6542 VOUT-.n104 VOUT-.t0 3.42907
R6543 VOUT-.n104 VOUT-.t18 3.42907
R6544 VOUT-.n107 VOUT-.t14 3.42907
R6545 VOUT-.n107 VOUT-.t17 3.42907
R6546 VOUT-.n110 VOUT-.n109 1.688
R6547 VOUT- VOUT-.n110 1.53175
R6548 VOUT-.n20 VOUT-.n1 1.313
R6549 VOUT-.n109 VOUT-.n101 1.1255
R6550 VOUT-.n19 VOUT-.n2 0.563
R6551 VOUT-.n9 VOUT-.n2 0.563
R6552 VOUT-.n9 VOUT-.n8 0.563
R6553 VOUT-.n12 VOUT-.n3 0.563
R6554 VOUT-.n15 VOUT-.n12 0.563
R6555 VOUT-.n16 VOUT-.n15 0.563
R6556 VOUT-.n48 VOUT-.n47 0.3295
R6557 VOUT-.n57 VOUT-.n56 0.3295
R6558 VOUT-.n55 VOUT-.n54 0.3295
R6559 VOUT-.n53 VOUT-.n52 0.3295
R6560 VOUT-.n51 VOUT-.n50 0.3295
R6561 VOUT-.n68 VOUT-.n49 0.3295
R6562 VOUT-.n68 VOUT-.n67 0.3295
R6563 VOUT-.n67 VOUT-.n66 0.3295
R6564 VOUT-.n66 VOUT-.n65 0.3295
R6565 VOUT-.n65 VOUT-.n64 0.3295
R6566 VOUT-.n64 VOUT-.n63 0.3295
R6567 VOUT-.n63 VOUT-.n62 0.3295
R6568 VOUT-.n62 VOUT-.n61 0.3295
R6569 VOUT-.n61 VOUT-.n60 0.3295
R6570 VOUT-.n60 VOUT-.n59 0.3295
R6571 VOUT-.n59 VOUT-.n58 0.3295
R6572 VOUT-.n71 VOUT-.n69 0.3295
R6573 VOUT-.n71 VOUT-.n70 0.3295
R6574 VOUT-.n74 VOUT-.n72 0.3295
R6575 VOUT-.n74 VOUT-.n73 0.3295
R6576 VOUT-.n77 VOUT-.n75 0.3295
R6577 VOUT-.n77 VOUT-.n76 0.3295
R6578 VOUT-.n80 VOUT-.n78 0.3295
R6579 VOUT-.n80 VOUT-.n79 0.3295
R6580 VOUT-.n83 VOUT-.n81 0.3295
R6581 VOUT-.n83 VOUT-.n82 0.3295
R6582 VOUT-.n86 VOUT-.n84 0.3295
R6583 VOUT-.n86 VOUT-.n85 0.3295
R6584 VOUT-.n89 VOUT-.n87 0.3295
R6585 VOUT-.n89 VOUT-.n88 0.3295
R6586 VOUT-.n92 VOUT-.n90 0.3295
R6587 VOUT-.n92 VOUT-.n91 0.3295
R6588 VOUT-.n95 VOUT-.n93 0.3295
R6589 VOUT-.n95 VOUT-.n94 0.3295
R6590 VOUT-.n22 VOUT-.n21 0.3295
R6591 VOUT-.n34 VOUT-.n23 0.3295
R6592 VOUT-.n34 VOUT-.n33 0.3295
R6593 VOUT-.n33 VOUT-.n32 0.3295
R6594 VOUT-.n32 VOUT-.n31 0.3295
R6595 VOUT-.n31 VOUT-.n30 0.3295
R6596 VOUT-.n30 VOUT-.n29 0.3295
R6597 VOUT-.n29 VOUT-.n28 0.3295
R6598 VOUT-.n28 VOUT-.n27 0.3295
R6599 VOUT-.n27 VOUT-.n26 0.3295
R6600 VOUT-.n26 VOUT-.n25 0.3295
R6601 VOUT-.n25 VOUT-.n24 0.3295
R6602 VOUT-.n37 VOUT-.n35 0.3295
R6603 VOUT-.n37 VOUT-.n36 0.3295
R6604 VOUT-.n40 VOUT-.n38 0.3295
R6605 VOUT-.n40 VOUT-.n39 0.3295
R6606 VOUT-.n43 VOUT-.n41 0.3295
R6607 VOUT-.n43 VOUT-.n42 0.3295
R6608 VOUT-.n46 VOUT-.n44 0.3295
R6609 VOUT-.n46 VOUT-.n45 0.3295
R6610 VOUT-.n97 VOUT-.n96 0.3295
R6611 VOUT-.n98 VOUT-.n97 0.3295
R6612 VOUT-.n99 VOUT-.n98 0.3295
R6613 VOUT-.n62 VOUT-.n57 0.306
R6614 VOUT-.n63 VOUT-.n55 0.306
R6615 VOUT-.n64 VOUT-.n53 0.306
R6616 VOUT-.n65 VOUT-.n51 0.306
R6617 VOUT-.n68 VOUT-.n48 0.2825
R6618 VOUT-.n71 VOUT-.n68 0.2825
R6619 VOUT-.n74 VOUT-.n71 0.2825
R6620 VOUT-.n77 VOUT-.n74 0.2825
R6621 VOUT-.n80 VOUT-.n77 0.2825
R6622 VOUT-.n83 VOUT-.n80 0.2825
R6623 VOUT-.n86 VOUT-.n83 0.2825
R6624 VOUT-.n89 VOUT-.n86 0.2825
R6625 VOUT-.n92 VOUT-.n89 0.2825
R6626 VOUT-.n95 VOUT-.n92 0.2825
R6627 VOUT-.n34 VOUT-.n22 0.2825
R6628 VOUT-.n37 VOUT-.n34 0.2825
R6629 VOUT-.n40 VOUT-.n37 0.2825
R6630 VOUT-.n43 VOUT-.n40 0.2825
R6631 VOUT-.n46 VOUT-.n43 0.2825
R6632 VOUT-.n97 VOUT-.n46 0.2825
R6633 VOUT-.n97 VOUT-.n95 0.2825
R6634 bgr_0.V_TOP.n20 bgr_0.V_TOP.t27 369.534
R6635 bgr_0.V_TOP.n14 bgr_0.V_TOP.t45 369.534
R6636 bgr_0.V_TOP.n37 bgr_0.V_TOP.n35 299.866
R6637 bgr_0.V_TOP.n37 bgr_0.V_TOP.n36 299.579
R6638 bgr_0.V_TOP.n13 bgr_0.V_TOP.n12 297.151
R6639 bgr_0.V_TOP.n33 bgr_0.V_TOP.n32 297.151
R6640 bgr_0.V_TOP.n40 bgr_0.V_TOP.n39 297.151
R6641 bgr_0.V_TOP.n43 bgr_0.V_TOP.n42 297.151
R6642 bgr_0.V_TOP.n21 bgr_0.V_TOP.n20 224.934
R6643 bgr_0.V_TOP.n22 bgr_0.V_TOP.n21 224.934
R6644 bgr_0.V_TOP.n23 bgr_0.V_TOP.n22 224.934
R6645 bgr_0.V_TOP.n24 bgr_0.V_TOP.n23 224.934
R6646 bgr_0.V_TOP.n25 bgr_0.V_TOP.n24 224.934
R6647 bgr_0.V_TOP.n26 bgr_0.V_TOP.n25 224.934
R6648 bgr_0.V_TOP.n27 bgr_0.V_TOP.n26 224.934
R6649 bgr_0.V_TOP.n15 bgr_0.V_TOP.n14 224.934
R6650 bgr_0.V_TOP.n16 bgr_0.V_TOP.n15 224.934
R6651 bgr_0.V_TOP.n17 bgr_0.V_TOP.n16 224.934
R6652 bgr_0.V_TOP.n18 bgr_0.V_TOP.n17 224.934
R6653 bgr_0.V_TOP.n19 bgr_0.V_TOP.n18 224.934
R6654 bgr_0.V_TOP.n29 bgr_0.V_TOP.n28 162.977
R6655 bgr_0.V_TOP.n20 bgr_0.V_TOP.t35 144.601
R6656 bgr_0.V_TOP.n21 bgr_0.V_TOP.t48 144.601
R6657 bgr_0.V_TOP.n22 bgr_0.V_TOP.t23 144.601
R6658 bgr_0.V_TOP.n23 bgr_0.V_TOP.t33 144.601
R6659 bgr_0.V_TOP.n24 bgr_0.V_TOP.t31 144.601
R6660 bgr_0.V_TOP.n25 bgr_0.V_TOP.t43 144.601
R6661 bgr_0.V_TOP.n26 bgr_0.V_TOP.t20 144.601
R6662 bgr_0.V_TOP.n27 bgr_0.V_TOP.t29 144.601
R6663 bgr_0.V_TOP.n14 bgr_0.V_TOP.t46 144.601
R6664 bgr_0.V_TOP.n15 bgr_0.V_TOP.t34 144.601
R6665 bgr_0.V_TOP.n16 bgr_0.V_TOP.t26 144.601
R6666 bgr_0.V_TOP.n17 bgr_0.V_TOP.t17 144.601
R6667 bgr_0.V_TOP.n18 bgr_0.V_TOP.t38 144.601
R6668 bgr_0.V_TOP.n19 bgr_0.V_TOP.t41 144.601
R6669 bgr_0.V_TOP.t1 bgr_0.V_TOP.n45 108.424
R6670 bgr_0.V_TOP.n28 bgr_0.V_TOP.n27 77.4126
R6671 bgr_0.V_TOP.n28 bgr_0.V_TOP.n19 77.4126
R6672 bgr_0.V_TOP.n29 bgr_0.V_TOP.t6 47.9838
R6673 bgr_0.V_TOP.n12 bgr_0.V_TOP.t10 39.4005
R6674 bgr_0.V_TOP.n12 bgr_0.V_TOP.t2 39.4005
R6675 bgr_0.V_TOP.n32 bgr_0.V_TOP.t12 39.4005
R6676 bgr_0.V_TOP.n32 bgr_0.V_TOP.t7 39.4005
R6677 bgr_0.V_TOP.n39 bgr_0.V_TOP.t11 39.4005
R6678 bgr_0.V_TOP.n39 bgr_0.V_TOP.t9 39.4005
R6679 bgr_0.V_TOP.n35 bgr_0.V_TOP.t3 39.4005
R6680 bgr_0.V_TOP.n35 bgr_0.V_TOP.t13 39.4005
R6681 bgr_0.V_TOP.n36 bgr_0.V_TOP.t0 39.4005
R6682 bgr_0.V_TOP.n36 bgr_0.V_TOP.t4 39.4005
R6683 bgr_0.V_TOP.n42 bgr_0.V_TOP.t5 39.4005
R6684 bgr_0.V_TOP.n42 bgr_0.V_TOP.t8 39.4005
R6685 bgr_0.V_TOP.n45 bgr_0.V_TOP.n10 37.1479
R6686 bgr_0.V_TOP.n45 bgr_0.V_TOP.n44 28.1496
R6687 bgr_0.V_TOP.n38 bgr_0.V_TOP.n37 9.61217
R6688 bgr_0.V_TOP.n43 bgr_0.V_TOP.n41 7.14633
R6689 bgr_0.V_TOP.n34 bgr_0.V_TOP.n13 7.14633
R6690 bgr_0.V_TOP.n30 bgr_0.V_TOP.n29 5.188
R6691 bgr_0.V_TOP.n33 bgr_0.V_TOP.n31 5.14633
R6692 bgr_0.V_TOP.n44 bgr_0.V_TOP.n43 5.14633
R6693 bgr_0.V_TOP.n30 bgr_0.V_TOP.n13 5.14633
R6694 bgr_0.V_TOP.n34 bgr_0.V_TOP.n33 5.02133
R6695 bgr_0.V_TOP.n41 bgr_0.V_TOP.n40 5.02133
R6696 bgr_0.V_TOP.n0 bgr_0.V_TOP.t24 4.8295
R6697 bgr_0.V_TOP.n1 bgr_0.V_TOP.t19 4.8295
R6698 bgr_0.V_TOP.n2 bgr_0.V_TOP.t16 4.8295
R6699 bgr_0.V_TOP.n3 bgr_0.V_TOP.t44 4.8295
R6700 bgr_0.V_TOP.n4 bgr_0.V_TOP.t39 4.8295
R6701 bgr_0.V_TOP.n5 bgr_0.V_TOP.t32 4.8295
R6702 bgr_0.V_TOP.n6 bgr_0.V_TOP.t14 4.8295
R6703 bgr_0.V_TOP.n7 bgr_0.V_TOP.t40 4.8295
R6704 bgr_0.V_TOP.n8 bgr_0.V_TOP.t28 4.8295
R6705 bgr_0.V_TOP.n0 bgr_0.V_TOP.t30 4.5005
R6706 bgr_0.V_TOP.n1 bgr_0.V_TOP.t25 4.5005
R6707 bgr_0.V_TOP.n2 bgr_0.V_TOP.t22 4.5005
R6708 bgr_0.V_TOP.n3 bgr_0.V_TOP.t18 4.5005
R6709 bgr_0.V_TOP.n4 bgr_0.V_TOP.t49 4.5005
R6710 bgr_0.V_TOP.n5 bgr_0.V_TOP.t42 4.5005
R6711 bgr_0.V_TOP.n6 bgr_0.V_TOP.t21 4.5005
R6712 bgr_0.V_TOP.n7 bgr_0.V_TOP.t15 4.5005
R6713 bgr_0.V_TOP.n10 bgr_0.V_TOP.t36 4.5005
R6714 bgr_0.V_TOP.n9 bgr_0.V_TOP.t47 4.5005
R6715 bgr_0.V_TOP.n8 bgr_0.V_TOP.t37 4.5005
R6716 bgr_0.V_TOP.n38 bgr_0.V_TOP.n11 4.5005
R6717 bgr_0.V_TOP.n41 bgr_0.V_TOP.n34 2.1255
R6718 bgr_0.V_TOP.n31 bgr_0.V_TOP.n30 2.1255
R6719 bgr_0.V_TOP.n31 bgr_0.V_TOP.n11 2.1255
R6720 bgr_0.V_TOP.n44 bgr_0.V_TOP.n11 2.1255
R6721 bgr_0.V_TOP.n40 bgr_0.V_TOP.n38 0.646333
R6722 bgr_0.V_TOP.n1 bgr_0.V_TOP.n0 0.3295
R6723 bgr_0.V_TOP.n3 bgr_0.V_TOP.n2 0.3295
R6724 bgr_0.V_TOP.n5 bgr_0.V_TOP.n4 0.3295
R6725 bgr_0.V_TOP.n7 bgr_0.V_TOP.n6 0.3295
R6726 bgr_0.V_TOP.n10 bgr_0.V_TOP.n9 0.3295
R6727 bgr_0.V_TOP.n9 bgr_0.V_TOP.n8 0.3295
R6728 bgr_0.V_TOP.n3 bgr_0.V_TOP.n1 0.2825
R6729 bgr_0.V_TOP.n5 bgr_0.V_TOP.n3 0.2825
R6730 bgr_0.V_TOP.n7 bgr_0.V_TOP.n5 0.2825
R6731 bgr_0.V_TOP.n8 bgr_0.V_TOP.n7 0.2825
R6732 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t13 703.528
R6733 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t14 703.231
R6734 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n15 540.556
R6735 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n16 540.556
R6736 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n8 297.151
R6737 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.n17 297.151
R6738 bgr_0.1st_Vout_2.n20 bgr_0.1st_Vout_2.n19 297.151
R6739 bgr_0.1st_Vout_2.n15 bgr_0.1st_Vout_2.t20 291.209
R6740 bgr_0.1st_Vout_2.n16 bgr_0.1st_Vout_2.t25 291.209
R6741 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.t9 242.3
R6742 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.n9 194.3
R6743 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.n10 194.3
R6744 bgr_0.1st_Vout_2.n15 bgr_0.1st_Vout_2.t33 162.675
R6745 bgr_0.1st_Vout_2.n16 bgr_0.1st_Vout_2.t34 162.675
R6746 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.n7 52.4165
R6747 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.t0 48.0005
R6748 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.t1 48.0005
R6749 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t10 48.0005
R6750 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t2 48.0005
R6751 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t5 39.4005
R6752 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t4 39.4005
R6753 bgr_0.1st_Vout_2.n17 bgr_0.1st_Vout_2.t6 39.4005
R6754 bgr_0.1st_Vout_2.n17 bgr_0.1st_Vout_2.t8 39.4005
R6755 bgr_0.1st_Vout_2.t3 bgr_0.1st_Vout_2.n20 39.4005
R6756 bgr_0.1st_Vout_2.n20 bgr_0.1st_Vout_2.t7 39.4005
R6757 bgr_0.1st_Vout_2.n18 bgr_0.1st_Vout_2.n0 7.08383
R6758 bgr_0.1st_Vout_2.n19 bgr_0.1st_Vout_2.n18 7.08383
R6759 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.n12 6.22967
R6760 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.n11 6.22967
R6761 bgr_0.1st_Vout_2.n14 bgr_0.1st_Vout_2.n13 6.04217
R6762 bgr_0.1st_Vout_2.n14 bgr_0.1st_Vout_2.n11 6.04217
R6763 bgr_0.1st_Vout_2.n19 bgr_0.1st_Vout_2.n3 5.45883
R6764 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n0 5.45883
R6765 bgr_0.1st_Vout_2.n18 bgr_0.1st_Vout_2.n5 4.95883
R6766 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.n4 4.85467
R6767 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t17 4.8295
R6768 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t35 4.8295
R6769 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t11 4.8295
R6770 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t27 4.8295
R6771 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t30 4.8295
R6772 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t19 4.8295
R6773 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t36 4.8295
R6774 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t26 4.8295
R6775 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t18 4.8295
R6776 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.n14 4.5005
R6777 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t12 4.5005
R6778 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t32 4.5005
R6779 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t31 4.5005
R6780 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t24 4.5005
R6781 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t23 4.5005
R6782 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t16 4.5005
R6783 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t29 4.5005
R6784 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t22 4.5005
R6785 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t28 4.5005
R6786 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t21 4.5005
R6787 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t15 4.5005
R6788 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.n1 4.5005
R6789 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.n6 3.1025
R6790 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n3 3.07862
R6791 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.n4 2.21925
R6792 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n2 2.03175
R6793 bgr_0.cap_res2.t0 bgr_0.cap_res2.t18 121.245
R6794 bgr_0.cap_res2.t13 bgr_0.cap_res2.t7 0.1603
R6795 bgr_0.cap_res2.t6 bgr_0.cap_res2.t1 0.1603
R6796 bgr_0.cap_res2.t11 bgr_0.cap_res2.t5 0.1603
R6797 bgr_0.cap_res2.t4 bgr_0.cap_res2.t20 0.1603
R6798 bgr_0.cap_res2.t19 bgr_0.cap_res2.t16 0.1603
R6799 bgr_0.cap_res2.n1 bgr_0.cap_res2.t3 0.159278
R6800 bgr_0.cap_res2.n2 bgr_0.cap_res2.t10 0.159278
R6801 bgr_0.cap_res2.n3 bgr_0.cap_res2.t17 0.159278
R6802 bgr_0.cap_res2.n4 bgr_0.cap_res2.t12 0.159278
R6803 bgr_0.cap_res2.n4 bgr_0.cap_res2.t15 0.1368
R6804 bgr_0.cap_res2.n4 bgr_0.cap_res2.t13 0.1368
R6805 bgr_0.cap_res2.n3 bgr_0.cap_res2.t9 0.1368
R6806 bgr_0.cap_res2.n3 bgr_0.cap_res2.t6 0.1368
R6807 bgr_0.cap_res2.n2 bgr_0.cap_res2.t14 0.1368
R6808 bgr_0.cap_res2.n2 bgr_0.cap_res2.t11 0.1368
R6809 bgr_0.cap_res2.n1 bgr_0.cap_res2.t8 0.1368
R6810 bgr_0.cap_res2.n1 bgr_0.cap_res2.t4 0.1368
R6811 bgr_0.cap_res2.n0 bgr_0.cap_res2.t2 0.1368
R6812 bgr_0.cap_res2.n0 bgr_0.cap_res2.t19 0.1368
R6813 bgr_0.cap_res2.t3 bgr_0.cap_res2.n0 0.00152174
R6814 bgr_0.cap_res2.t10 bgr_0.cap_res2.n1 0.00152174
R6815 bgr_0.cap_res2.t17 bgr_0.cap_res2.n2 0.00152174
R6816 bgr_0.cap_res2.t12 bgr_0.cap_res2.n3 0.00152174
R6817 bgr_0.cap_res2.t18 bgr_0.cap_res2.n4 0.00152174
R6818 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 120.504
R6819 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 100.322
R6820 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 99.7078
R6821 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n21 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n20 35.7193
R6822 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n21 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 31.4376
R6823 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 24.288
R6824 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 24.288
R6825 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 24.288
R6826 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n14 24.288
R6827 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n17 24.288
R6828 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 24.0005
R6829 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 24.0005
R6830 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 24.0005
R6831 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 24.0005
R6832 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 8.0005
R6833 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 8.0005
R6834 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 8.0005
R6835 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 8.0005
R6836 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 8.0005
R6837 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 8.0005
R6838 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 8.0005
R6839 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 8.0005
R6840 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 8.0005
R6841 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 8.0005
R6842 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n19 5.96925
R6843 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n16 5.7505
R6844 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 5.7505
R6845 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 5.7505
R6846 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 5.188
R6847 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 5.188
R6848 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 5.188
R6849 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 5.188
R6850 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 5.188
R6851 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n15 5.188
R6852 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n18 5.188
R6853 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n13 0.563
R6854 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 0.563
R6855 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 0.563
R6856 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 0.563
R6857 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 0.563
R6858 bgr_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n21 0.047375
R6859 two_stage_opamp_dummy_magic_0.V_source.n70 two_stage_opamp_dummy_magic_0.V_source.t29 66.2047
R6860 two_stage_opamp_dummy_magic_0.V_source.n1 two_stage_opamp_dummy_magic_0.V_source.n0 49.3505
R6861 two_stage_opamp_dummy_magic_0.V_source.n4 two_stage_opamp_dummy_magic_0.V_source.n3 49.3505
R6862 two_stage_opamp_dummy_magic_0.V_source.n7 two_stage_opamp_dummy_magic_0.V_source.n6 49.3505
R6863 two_stage_opamp_dummy_magic_0.V_source.n10 two_stage_opamp_dummy_magic_0.V_source.n9 49.3505
R6864 two_stage_opamp_dummy_magic_0.V_source.n14 two_stage_opamp_dummy_magic_0.V_source.n13 49.3505
R6865 two_stage_opamp_dummy_magic_0.V_source.n19 two_stage_opamp_dummy_magic_0.V_source.n18 49.3505
R6866 two_stage_opamp_dummy_magic_0.V_source.n21 two_stage_opamp_dummy_magic_0.V_source.n20 49.3505
R6867 two_stage_opamp_dummy_magic_0.V_source.n25 two_stage_opamp_dummy_magic_0.V_source.n24 49.3505
R6868 two_stage_opamp_dummy_magic_0.V_source.n28 two_stage_opamp_dummy_magic_0.V_source.n27 49.3505
R6869 two_stage_opamp_dummy_magic_0.V_source.n31 two_stage_opamp_dummy_magic_0.V_source.n30 49.3505
R6870 two_stage_opamp_dummy_magic_0.V_source.n39 two_stage_opamp_dummy_magic_0.V_source.n38 32.3838
R6871 two_stage_opamp_dummy_magic_0.V_source.n41 two_stage_opamp_dummy_magic_0.V_source.n40 32.3838
R6872 two_stage_opamp_dummy_magic_0.V_source.n47 two_stage_opamp_dummy_magic_0.V_source.n46 32.3838
R6873 two_stage_opamp_dummy_magic_0.V_source.n49 two_stage_opamp_dummy_magic_0.V_source.n48 32.3838
R6874 two_stage_opamp_dummy_magic_0.V_source.n53 two_stage_opamp_dummy_magic_0.V_source.n52 32.3838
R6875 two_stage_opamp_dummy_magic_0.V_source.n56 two_stage_opamp_dummy_magic_0.V_source.n55 32.3838
R6876 two_stage_opamp_dummy_magic_0.V_source.n60 two_stage_opamp_dummy_magic_0.V_source.n59 32.3838
R6877 two_stage_opamp_dummy_magic_0.V_source.n63 two_stage_opamp_dummy_magic_0.V_source.n62 32.3838
R6878 two_stage_opamp_dummy_magic_0.V_source.n67 two_stage_opamp_dummy_magic_0.V_source.n66 32.3838
R6879 two_stage_opamp_dummy_magic_0.V_source.n72 two_stage_opamp_dummy_magic_0.V_source.n71 32.3838
R6880 two_stage_opamp_dummy_magic_0.V_source.n0 two_stage_opamp_dummy_magic_0.V_source.t0 16.0005
R6881 two_stage_opamp_dummy_magic_0.V_source.n0 two_stage_opamp_dummy_magic_0.V_source.t3 16.0005
R6882 two_stage_opamp_dummy_magic_0.V_source.n3 two_stage_opamp_dummy_magic_0.V_source.t31 16.0005
R6883 two_stage_opamp_dummy_magic_0.V_source.n3 two_stage_opamp_dummy_magic_0.V_source.t38 16.0005
R6884 two_stage_opamp_dummy_magic_0.V_source.n6 two_stage_opamp_dummy_magic_0.V_source.t6 16.0005
R6885 two_stage_opamp_dummy_magic_0.V_source.n6 two_stage_opamp_dummy_magic_0.V_source.t5 16.0005
R6886 two_stage_opamp_dummy_magic_0.V_source.n9 two_stage_opamp_dummy_magic_0.V_source.t33 16.0005
R6887 two_stage_opamp_dummy_magic_0.V_source.n9 two_stage_opamp_dummy_magic_0.V_source.t30 16.0005
R6888 two_stage_opamp_dummy_magic_0.V_source.n13 two_stage_opamp_dummy_magic_0.V_source.t25 16.0005
R6889 two_stage_opamp_dummy_magic_0.V_source.n13 two_stage_opamp_dummy_magic_0.V_source.t39 16.0005
R6890 two_stage_opamp_dummy_magic_0.V_source.n18 two_stage_opamp_dummy_magic_0.V_source.t32 16.0005
R6891 two_stage_opamp_dummy_magic_0.V_source.n18 two_stage_opamp_dummy_magic_0.V_source.t37 16.0005
R6892 two_stage_opamp_dummy_magic_0.V_source.n20 two_stage_opamp_dummy_magic_0.V_source.t1 16.0005
R6893 two_stage_opamp_dummy_magic_0.V_source.n20 two_stage_opamp_dummy_magic_0.V_source.t28 16.0005
R6894 two_stage_opamp_dummy_magic_0.V_source.n24 two_stage_opamp_dummy_magic_0.V_source.t26 16.0005
R6895 two_stage_opamp_dummy_magic_0.V_source.n24 two_stage_opamp_dummy_magic_0.V_source.t2 16.0005
R6896 two_stage_opamp_dummy_magic_0.V_source.n27 two_stage_opamp_dummy_magic_0.V_source.t40 16.0005
R6897 two_stage_opamp_dummy_magic_0.V_source.n27 two_stage_opamp_dummy_magic_0.V_source.t36 16.0005
R6898 two_stage_opamp_dummy_magic_0.V_source.n30 two_stage_opamp_dummy_magic_0.V_source.t35 16.0005
R6899 two_stage_opamp_dummy_magic_0.V_source.n30 two_stage_opamp_dummy_magic_0.V_source.t4 16.0005
R6900 two_stage_opamp_dummy_magic_0.V_source.n38 two_stage_opamp_dummy_magic_0.V_source.t34 9.6005
R6901 two_stage_opamp_dummy_magic_0.V_source.n38 two_stage_opamp_dummy_magic_0.V_source.t27 9.6005
R6902 two_stage_opamp_dummy_magic_0.V_source.n40 two_stage_opamp_dummy_magic_0.V_source.t23 9.6005
R6903 two_stage_opamp_dummy_magic_0.V_source.n40 two_stage_opamp_dummy_magic_0.V_source.t17 9.6005
R6904 two_stage_opamp_dummy_magic_0.V_source.n46 two_stage_opamp_dummy_magic_0.V_source.t10 9.6005
R6905 two_stage_opamp_dummy_magic_0.V_source.n46 two_stage_opamp_dummy_magic_0.V_source.t16 9.6005
R6906 two_stage_opamp_dummy_magic_0.V_source.n48 two_stage_opamp_dummy_magic_0.V_source.t12 9.6005
R6907 two_stage_opamp_dummy_magic_0.V_source.n48 two_stage_opamp_dummy_magic_0.V_source.t20 9.6005
R6908 two_stage_opamp_dummy_magic_0.V_source.n52 two_stage_opamp_dummy_magic_0.V_source.t14 9.6005
R6909 two_stage_opamp_dummy_magic_0.V_source.n52 two_stage_opamp_dummy_magic_0.V_source.t22 9.6005
R6910 two_stage_opamp_dummy_magic_0.V_source.n55 two_stage_opamp_dummy_magic_0.V_source.t18 9.6005
R6911 two_stage_opamp_dummy_magic_0.V_source.n55 two_stage_opamp_dummy_magic_0.V_source.t8 9.6005
R6912 two_stage_opamp_dummy_magic_0.V_source.n59 two_stage_opamp_dummy_magic_0.V_source.t15 9.6005
R6913 two_stage_opamp_dummy_magic_0.V_source.n59 two_stage_opamp_dummy_magic_0.V_source.t7 9.6005
R6914 two_stage_opamp_dummy_magic_0.V_source.n62 two_stage_opamp_dummy_magic_0.V_source.t19 9.6005
R6915 two_stage_opamp_dummy_magic_0.V_source.n62 two_stage_opamp_dummy_magic_0.V_source.t9 9.6005
R6916 two_stage_opamp_dummy_magic_0.V_source.n66 two_stage_opamp_dummy_magic_0.V_source.t21 9.6005
R6917 two_stage_opamp_dummy_magic_0.V_source.n66 two_stage_opamp_dummy_magic_0.V_source.t11 9.6005
R6918 two_stage_opamp_dummy_magic_0.V_source.t24 two_stage_opamp_dummy_magic_0.V_source.n72 9.6005
R6919 two_stage_opamp_dummy_magic_0.V_source.n72 two_stage_opamp_dummy_magic_0.V_source.t13 9.6005
R6920 two_stage_opamp_dummy_magic_0.V_source.n47 two_stage_opamp_dummy_magic_0.V_source.n45 5.89633
R6921 two_stage_opamp_dummy_magic_0.V_source.n39 two_stage_opamp_dummy_magic_0.V_source.n36 5.89633
R6922 two_stage_opamp_dummy_magic_0.V_source.n50 two_stage_opamp_dummy_magic_0.V_source.n47 5.70883
R6923 two_stage_opamp_dummy_magic_0.V_source.n42 two_stage_opamp_dummy_magic_0.V_source.n39 5.70883
R6924 two_stage_opamp_dummy_magic_0.V_source.n22 two_stage_opamp_dummy_magic_0.V_source.n19 5.6255
R6925 two_stage_opamp_dummy_magic_0.V_source.n5 two_stage_opamp_dummy_magic_0.V_source.n4 5.6255
R6926 two_stage_opamp_dummy_magic_0.V_source.n31 two_stage_opamp_dummy_magic_0.V_source.n29 5.45883
R6927 two_stage_opamp_dummy_magic_0.V_source.n19 two_stage_opamp_dummy_magic_0.V_source.n17 5.45883
R6928 two_stage_opamp_dummy_magic_0.V_source.n8 two_stage_opamp_dummy_magic_0.V_source.n4 5.45883
R6929 two_stage_opamp_dummy_magic_0.V_source.n12 two_stage_opamp_dummy_magic_0.V_source.n1 5.45883
R6930 two_stage_opamp_dummy_magic_0.V_source.n41 two_stage_opamp_dummy_magic_0.V_source.n36 5.33383
R6931 two_stage_opamp_dummy_magic_0.V_source.n49 two_stage_opamp_dummy_magic_0.V_source.n45 5.33383
R6932 two_stage_opamp_dummy_magic_0.V_source.n54 two_stage_opamp_dummy_magic_0.V_source.n53 5.33383
R6933 two_stage_opamp_dummy_magic_0.V_source.n57 two_stage_opamp_dummy_magic_0.V_source.n56 5.33383
R6934 two_stage_opamp_dummy_magic_0.V_source.n60 two_stage_opamp_dummy_magic_0.V_source.n58 5.33383
R6935 two_stage_opamp_dummy_magic_0.V_source.n63 two_stage_opamp_dummy_magic_0.V_source.n37 5.33383
R6936 two_stage_opamp_dummy_magic_0.V_source.n68 two_stage_opamp_dummy_magic_0.V_source.n67 5.33383
R6937 two_stage_opamp_dummy_magic_0.V_source.n42 two_stage_opamp_dummy_magic_0.V_source.n41 5.14633
R6938 two_stage_opamp_dummy_magic_0.V_source.n50 two_stage_opamp_dummy_magic_0.V_source.n49 5.14633
R6939 two_stage_opamp_dummy_magic_0.V_source.n53 two_stage_opamp_dummy_magic_0.V_source.n51 5.14633
R6940 two_stage_opamp_dummy_magic_0.V_source.n56 two_stage_opamp_dummy_magic_0.V_source.n44 5.14633
R6941 two_stage_opamp_dummy_magic_0.V_source.n61 two_stage_opamp_dummy_magic_0.V_source.n60 5.14633
R6942 two_stage_opamp_dummy_magic_0.V_source.n64 two_stage_opamp_dummy_magic_0.V_source.n63 5.14633
R6943 two_stage_opamp_dummy_magic_0.V_source.n67 two_stage_opamp_dummy_magic_0.V_source.n65 5.14633
R6944 two_stage_opamp_dummy_magic_0.V_source.n7 two_stage_opamp_dummy_magic_0.V_source.n5 5.063
R6945 two_stage_opamp_dummy_magic_0.V_source.n10 two_stage_opamp_dummy_magic_0.V_source.n2 5.063
R6946 two_stage_opamp_dummy_magic_0.V_source.n15 two_stage_opamp_dummy_magic_0.V_source.n14 5.063
R6947 two_stage_opamp_dummy_magic_0.V_source.n22 two_stage_opamp_dummy_magic_0.V_source.n21 5.063
R6948 two_stage_opamp_dummy_magic_0.V_source.n25 two_stage_opamp_dummy_magic_0.V_source.n23 5.063
R6949 two_stage_opamp_dummy_magic_0.V_source.n28 two_stage_opamp_dummy_magic_0.V_source.n16 5.063
R6950 two_stage_opamp_dummy_magic_0.V_source.n32 two_stage_opamp_dummy_magic_0.V_source.n31 5.063
R6951 two_stage_opamp_dummy_magic_0.V_source.n8 two_stage_opamp_dummy_magic_0.V_source.n7 4.89633
R6952 two_stage_opamp_dummy_magic_0.V_source.n11 two_stage_opamp_dummy_magic_0.V_source.n10 4.89633
R6953 two_stage_opamp_dummy_magic_0.V_source.n14 two_stage_opamp_dummy_magic_0.V_source.n12 4.89633
R6954 two_stage_opamp_dummy_magic_0.V_source.n21 two_stage_opamp_dummy_magic_0.V_source.n17 4.89633
R6955 two_stage_opamp_dummy_magic_0.V_source.n26 two_stage_opamp_dummy_magic_0.V_source.n25 4.89633
R6956 two_stage_opamp_dummy_magic_0.V_source.n29 two_stage_opamp_dummy_magic_0.V_source.n28 4.89633
R6957 two_stage_opamp_dummy_magic_0.V_source.n34 two_stage_opamp_dummy_magic_0.V_source.n33 4.5005
R6958 two_stage_opamp_dummy_magic_0.V_source.n43 two_stage_opamp_dummy_magic_0.V_source.n35 4.5005
R6959 two_stage_opamp_dummy_magic_0.V_source.n70 two_stage_opamp_dummy_magic_0.V_source.n69 4.5005
R6960 two_stage_opamp_dummy_magic_0.V_source.n33 two_stage_opamp_dummy_magic_0.V_source.n32 3.6255
R6961 two_stage_opamp_dummy_magic_0.V_source.n35 two_stage_opamp_dummy_magic_0.V_source.n34 1.738
R6962 two_stage_opamp_dummy_magic_0.V_source.n71 two_stage_opamp_dummy_magic_0.V_source.n70 0.833833
R6963 two_stage_opamp_dummy_magic_0.V_source.n71 two_stage_opamp_dummy_magic_0.V_source.n35 0.633833
R6964 two_stage_opamp_dummy_magic_0.V_source.n29 two_stage_opamp_dummy_magic_0.V_source.n26 0.563
R6965 two_stage_opamp_dummy_magic_0.V_source.n26 two_stage_opamp_dummy_magic_0.V_source.n17 0.563
R6966 two_stage_opamp_dummy_magic_0.V_source.n23 two_stage_opamp_dummy_magic_0.V_source.n22 0.563
R6967 two_stage_opamp_dummy_magic_0.V_source.n23 two_stage_opamp_dummy_magic_0.V_source.n16 0.563
R6968 two_stage_opamp_dummy_magic_0.V_source.n32 two_stage_opamp_dummy_magic_0.V_source.n16 0.563
R6969 two_stage_opamp_dummy_magic_0.V_source.n33 two_stage_opamp_dummy_magic_0.V_source.n15 0.563
R6970 two_stage_opamp_dummy_magic_0.V_source.n15 two_stage_opamp_dummy_magic_0.V_source.n2 0.563
R6971 two_stage_opamp_dummy_magic_0.V_source.n5 two_stage_opamp_dummy_magic_0.V_source.n2 0.563
R6972 two_stage_opamp_dummy_magic_0.V_source.n11 two_stage_opamp_dummy_magic_0.V_source.n8 0.563
R6973 two_stage_opamp_dummy_magic_0.V_source.n12 two_stage_opamp_dummy_magic_0.V_source.n11 0.563
R6974 two_stage_opamp_dummy_magic_0.V_source.n34 two_stage_opamp_dummy_magic_0.V_source.n1 0.563
R6975 two_stage_opamp_dummy_magic_0.V_source.n69 two_stage_opamp_dummy_magic_0.V_source.n68 0.563
R6976 two_stage_opamp_dummy_magic_0.V_source.n68 two_stage_opamp_dummy_magic_0.V_source.n37 0.563
R6977 two_stage_opamp_dummy_magic_0.V_source.n58 two_stage_opamp_dummy_magic_0.V_source.n37 0.563
R6978 two_stage_opamp_dummy_magic_0.V_source.n58 two_stage_opamp_dummy_magic_0.V_source.n57 0.563
R6979 two_stage_opamp_dummy_magic_0.V_source.n57 two_stage_opamp_dummy_magic_0.V_source.n54 0.563
R6980 two_stage_opamp_dummy_magic_0.V_source.n54 two_stage_opamp_dummy_magic_0.V_source.n45 0.563
R6981 two_stage_opamp_dummy_magic_0.V_source.n51 two_stage_opamp_dummy_magic_0.V_source.n50 0.563
R6982 two_stage_opamp_dummy_magic_0.V_source.n51 two_stage_opamp_dummy_magic_0.V_source.n44 0.563
R6983 two_stage_opamp_dummy_magic_0.V_source.n61 two_stage_opamp_dummy_magic_0.V_source.n44 0.563
R6984 two_stage_opamp_dummy_magic_0.V_source.n64 two_stage_opamp_dummy_magic_0.V_source.n61 0.563
R6985 two_stage_opamp_dummy_magic_0.V_source.n65 two_stage_opamp_dummy_magic_0.V_source.n64 0.563
R6986 two_stage_opamp_dummy_magic_0.V_source.n65 two_stage_opamp_dummy_magic_0.V_source.n43 0.563
R6987 two_stage_opamp_dummy_magic_0.V_source.n43 two_stage_opamp_dummy_magic_0.V_source.n42 0.563
R6988 two_stage_opamp_dummy_magic_0.V_source.n69 two_stage_opamp_dummy_magic_0.V_source.n36 0.563
R6989 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.t1 530.833
R6990 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n13 490.228
R6991 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n8 490.166
R6992 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n14 420.858
R6993 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t13 385.601
R6994 bgr_0.NFET_GATE_10uA.t1 bgr_0.NFET_GATE_10uA.n18 385.601
R6995 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t17 369.534
R6996 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t20 369.534
R6997 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n20 330.276
R6998 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.t23 208.868
R6999 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.t6 208.868
R7000 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t14 208.868
R7001 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.t22 208.868
R7002 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.t10 208.868
R7003 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.t16 208.868
R7004 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.t11 192.8
R7005 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.t18 192.8
R7006 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.t5 192.8
R7007 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t12 192.8
R7008 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t19 192.8
R7009 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.t7 192.8
R7010 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t8 192.8
R7011 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.t15 192.8
R7012 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.t21 192.8
R7013 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t9 192.8
R7014 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.n2 176.733
R7015 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.n1 176.733
R7016 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n12 176.733
R7017 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.n11 176.733
R7018 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.n10 176.733
R7019 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.n9 176.733
R7020 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.n4 176.733
R7021 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.n5 176.733
R7022 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.n6 176.733
R7023 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n7 176.733
R7024 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.n17 176.733
R7025 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.n16 176.733
R7026 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.n0 97.638
R7027 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n3 56.2338
R7028 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.n15 56.2338
R7029 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t0 39.4005
R7030 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t4 39.4005
R7031 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t3 24.0005
R7032 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t2 24.0005
R7033 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n19 21.0505
R7034 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.t27 746.673
R7035 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.t1 721.625
R7036 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.t17 611.739
R7037 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.t29 611.739
R7038 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.t32 611.739
R7039 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.t22 611.739
R7040 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.t13 563.451
R7041 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.t24 463.925
R7042 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.t18 463.925
R7043 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.t15 421.75
R7044 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.t12 421.75
R7045 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.t30 421.75
R7046 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.t11 421.75
R7047 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.t14 421.75
R7048 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.t16 421.75
R7049 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.t19 421.75
R7050 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.t26 421.75
R7051 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.t21 421.75
R7052 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.t23 421.75
R7053 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.t20 421.75
R7054 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.t28 421.75
R7055 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.t25 421.75
R7056 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.t31 421.75
R7057 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.n14 391.913
R7058 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.n22 391.351
R7059 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.n19 167.094
R7060 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.n20 167.094
R7061 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.n15 167.094
R7062 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.n16 167.094
R7063 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.n17 167.094
R7064 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.n10 167.094
R7065 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.n11 167.094
R7066 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.n12 167.094
R7067 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.n7 167.094
R7068 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.n8 167.094
R7069 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.n21 147.814
R7070 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.n18 147.814
R7071 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.n13 147.814
R7072 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.n9 147.814
R7073 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.n0 100.323
R7074 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.n1 99.707
R7075 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n27 97.1505
R7076 two_stage_opamp_dummy_magic_0.Vb2.n30 two_stage_opamp_dummy_magic_0.Vb2.n29 97.1505
R7077 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.n4 67.013
R7078 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.n25 62.4786
R7079 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.t7 24.0005
R7080 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.t4 24.0005
R7081 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t5 24.0005
R7082 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t3 24.0005
R7083 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.t9 24.0005
R7084 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.t6 24.0005
R7085 two_stage_opamp_dummy_magic_0.Vb2.t8 two_stage_opamp_dummy_magic_0.Vb2.n30 24.0005
R7086 two_stage_opamp_dummy_magic_0.Vb2.n30 two_stage_opamp_dummy_magic_0.Vb2.t10 24.0005
R7087 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.n23 13.4067
R7088 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n28 11.2922
R7089 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.t2 11.2576
R7090 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.t0 11.2576
R7091 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.n2 7.39572
R7092 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.n5 7.35988
R7093 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n3 5.188
R7094 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n26 5.188
R7095 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.n24 4.55362
R7096 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.n3 1.2505
R7097 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.n6 1.14112
R7098 two_stage_opamp_dummy_magic_0.VD4.n24 two_stage_opamp_dummy_magic_0.VD4.t27 671.418
R7099 two_stage_opamp_dummy_magic_0.VD4.n23 two_stage_opamp_dummy_magic_0.VD4.t24 671.418
R7100 two_stage_opamp_dummy_magic_0.VD4.t28 two_stage_opamp_dummy_magic_0.VD4.n41 213.131
R7101 two_stage_opamp_dummy_magic_0.VD4.n42 two_stage_opamp_dummy_magic_0.VD4.t25 213.131
R7102 two_stage_opamp_dummy_magic_0.VD4.t10 two_stage_opamp_dummy_magic_0.VD4.t28 146.155
R7103 two_stage_opamp_dummy_magic_0.VD4.t14 two_stage_opamp_dummy_magic_0.VD4.t10 146.155
R7104 two_stage_opamp_dummy_magic_0.VD4.t18 two_stage_opamp_dummy_magic_0.VD4.t14 146.155
R7105 two_stage_opamp_dummy_magic_0.VD4.t2 two_stage_opamp_dummy_magic_0.VD4.t18 146.155
R7106 two_stage_opamp_dummy_magic_0.VD4.t6 two_stage_opamp_dummy_magic_0.VD4.t2 146.155
R7107 two_stage_opamp_dummy_magic_0.VD4.t8 two_stage_opamp_dummy_magic_0.VD4.t6 146.155
R7108 two_stage_opamp_dummy_magic_0.VD4.t12 two_stage_opamp_dummy_magic_0.VD4.t8 146.155
R7109 two_stage_opamp_dummy_magic_0.VD4.t16 two_stage_opamp_dummy_magic_0.VD4.t12 146.155
R7110 two_stage_opamp_dummy_magic_0.VD4.t20 two_stage_opamp_dummy_magic_0.VD4.t16 146.155
R7111 two_stage_opamp_dummy_magic_0.VD4.t4 two_stage_opamp_dummy_magic_0.VD4.t20 146.155
R7112 two_stage_opamp_dummy_magic_0.VD4.t25 two_stage_opamp_dummy_magic_0.VD4.t4 146.155
R7113 two_stage_opamp_dummy_magic_0.VD4.n41 two_stage_opamp_dummy_magic_0.VD4.t29 76.2576
R7114 two_stage_opamp_dummy_magic_0.VD4.n42 two_stage_opamp_dummy_magic_0.VD4.t26 76.2576
R7115 two_stage_opamp_dummy_magic_0.VD4.n38 two_stage_opamp_dummy_magic_0.VD4.n37 66.0338
R7116 two_stage_opamp_dummy_magic_0.VD4.n34 two_stage_opamp_dummy_magic_0.VD4.n33 66.0338
R7117 two_stage_opamp_dummy_magic_0.VD4.n31 two_stage_opamp_dummy_magic_0.VD4.n30 66.0338
R7118 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n26 66.0338
R7119 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.n4 66.0338
R7120 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n7 66.0338
R7121 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n10 66.0338
R7122 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.n14 66.0338
R7123 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.n17 66.0338
R7124 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.n20 66.0338
R7125 two_stage_opamp_dummy_magic_0.VD4.n47 two_stage_opamp_dummy_magic_0.VD4.n46 66.0338
R7126 two_stage_opamp_dummy_magic_0.VD4.n37 two_stage_opamp_dummy_magic_0.VD4.t11 11.2576
R7127 two_stage_opamp_dummy_magic_0.VD4.n37 two_stage_opamp_dummy_magic_0.VD4.t15 11.2576
R7128 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.t19 11.2576
R7129 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.t3 11.2576
R7130 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.t7 11.2576
R7131 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.t9 11.2576
R7132 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.t13 11.2576
R7133 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.t17 11.2576
R7134 two_stage_opamp_dummy_magic_0.VD4.n4 two_stage_opamp_dummy_magic_0.VD4.t37 11.2576
R7135 two_stage_opamp_dummy_magic_0.VD4.n4 two_stage_opamp_dummy_magic_0.VD4.t23 11.2576
R7136 two_stage_opamp_dummy_magic_0.VD4.n7 two_stage_opamp_dummy_magic_0.VD4.t1 11.2576
R7137 two_stage_opamp_dummy_magic_0.VD4.n7 two_stage_opamp_dummy_magic_0.VD4.t31 11.2576
R7138 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.t0 11.2576
R7139 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.t35 11.2576
R7140 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.t32 11.2576
R7141 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.t34 11.2576
R7142 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.t33 11.2576
R7143 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.t30 11.2576
R7144 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.t22 11.2576
R7145 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.t36 11.2576
R7146 two_stage_opamp_dummy_magic_0.VD4.t21 two_stage_opamp_dummy_magic_0.VD4.n47 11.2576
R7147 two_stage_opamp_dummy_magic_0.VD4.n47 two_stage_opamp_dummy_magic_0.VD4.t5 11.2576
R7148 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.n19 5.91717
R7149 two_stage_opamp_dummy_magic_0.VD4.n6 two_stage_opamp_dummy_magic_0.VD4.n5 5.91717
R7150 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.n5 5.91717
R7151 two_stage_opamp_dummy_magic_0.VD4.n40 two_stage_opamp_dummy_magic_0.VD4.n39 5.91717
R7152 two_stage_opamp_dummy_magic_0.VD4.n38 two_stage_opamp_dummy_magic_0.VD4.n36 5.563
R7153 two_stage_opamp_dummy_magic_0.VD4.n35 two_stage_opamp_dummy_magic_0.VD4.n34 5.563
R7154 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.n31 5.563
R7155 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.n27 5.563
R7156 two_stage_opamp_dummy_magic_0.VD4.n46 two_stage_opamp_dummy_magic_0.VD4.n0 5.563
R7157 two_stage_opamp_dummy_magic_0.VD4.n23 two_stage_opamp_dummy_magic_0.VD4.n0 5.313
R7158 two_stage_opamp_dummy_magic_0.VD4.n36 two_stage_opamp_dummy_magic_0.VD4.n24 5.313
R7159 two_stage_opamp_dummy_magic_0.VD4.n39 two_stage_opamp_dummy_magic_0.VD4.n38 5.29217
R7160 two_stage_opamp_dummy_magic_0.VD4.n34 two_stage_opamp_dummy_magic_0.VD4.n25 5.29217
R7161 two_stage_opamp_dummy_magic_0.VD4.n31 two_stage_opamp_dummy_magic_0.VD4.n29 5.29217
R7162 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n1 5.29217
R7163 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.n8 5.29217
R7164 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n6 5.29217
R7165 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n11 5.29217
R7166 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n3 5.29217
R7167 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.n13 5.29217
R7168 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.n15 5.29217
R7169 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.n2 5.29217
R7170 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.n18 5.29217
R7171 two_stage_opamp_dummy_magic_0.VD4.n22 two_stage_opamp_dummy_magic_0.VD4.n21 5.29217
R7172 two_stage_opamp_dummy_magic_0.VD4.n44 two_stage_opamp_dummy_magic_0.VD4.n43 5.29217
R7173 two_stage_opamp_dummy_magic_0.VD4.n46 two_stage_opamp_dummy_magic_0.VD4.n45 5.29217
R7174 two_stage_opamp_dummy_magic_0.VD4.n44 two_stage_opamp_dummy_magic_0.VD4.n22 2.5005
R7175 two_stage_opamp_dummy_magic_0.VD4.n43 two_stage_opamp_dummy_magic_0.VD4.n42 1.03383
R7176 two_stage_opamp_dummy_magic_0.VD4.n41 two_stage_opamp_dummy_magic_0.VD4.n40 1.03383
R7177 two_stage_opamp_dummy_magic_0.VD4.n43 two_stage_opamp_dummy_magic_0.VD4.n23 0.8755
R7178 two_stage_opamp_dummy_magic_0.VD4.n40 two_stage_opamp_dummy_magic_0.VD4.n24 0.8755
R7179 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.n16 0.6255
R7180 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.n3 0.6255
R7181 two_stage_opamp_dummy_magic_0.VD4.n6 two_stage_opamp_dummy_magic_0.VD4.n3 0.6255
R7182 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n9 0.6255
R7183 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.n12 0.6255
R7184 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.n2 0.6255
R7185 two_stage_opamp_dummy_magic_0.VD4.n22 two_stage_opamp_dummy_magic_0.VD4.n2 0.6255
R7186 two_stage_opamp_dummy_magic_0.VD4.n45 two_stage_opamp_dummy_magic_0.VD4.n44 0.6255
R7187 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.n0 0.6255
R7188 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.n28 0.6255
R7189 two_stage_opamp_dummy_magic_0.VD4.n35 two_stage_opamp_dummy_magic_0.VD4.n32 0.6255
R7190 two_stage_opamp_dummy_magic_0.VD4.n36 two_stage_opamp_dummy_magic_0.VD4.n35 0.6255
R7191 two_stage_opamp_dummy_magic_0.VD4.n39 two_stage_opamp_dummy_magic_0.VD4.n25 0.6255
R7192 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.n25 0.6255
R7193 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.n1 0.6255
R7194 two_stage_opamp_dummy_magic_0.VD4.n45 two_stage_opamp_dummy_magic_0.VD4.n1 0.6255
R7195 a_7460_23988.t0 a_7460_23988.t1 178.133
R7196 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 739.067
R7197 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 724.936
R7198 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 688.859
R7199 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 577.866
R7200 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 530.201
R7201 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 530.201
R7202 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 530.201
R7203 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 514.134
R7204 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 361.531
R7205 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 208.868
R7206 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 208.868
R7207 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 208.868
R7208 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 208.868
R7209 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 208.868
R7210 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 208.868
R7211 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 208.868
R7212 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 208.868
R7213 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 208.868
R7214 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 176.733
R7215 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 176.733
R7216 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 176.733
R7217 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 176.733
R7218 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 174.726
R7219 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 174.726
R7220 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 174.726
R7221 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 174.726
R7222 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 128.534
R7223 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 128.534
R7224 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 124.579
R7225 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 74.288
R7226 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 74.288
R7227 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n21 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n20 74.288
R7228 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n23 45.6567
R7229 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 13.1338
R7230 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 13.1338
R7231 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 13.1338
R7232 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 13.1338
R7233 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n20 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 13.1338
R7234 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n20 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 13.1338
R7235 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 10.1672
R7236 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n23 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n22 10.0317
R7237 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n21 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 9.813
R7238 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 9.813
R7239 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 5.79217
R7240 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n22 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n21 5.79217
R7241 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 5.438
R7242 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n23 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 4.438
R7243 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n22 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 4.3755
R7244 bgr_0.V_p_2.n3 bgr_0.V_p_2.n4 194.3
R7245 bgr_0.V_p_2.n6 bgr_0.V_p_2.n5 194.3
R7246 bgr_0.V_p_2.n2 bgr_0.V_p_2.n7 194.3
R7247 bgr_0.V_p_2.n9 bgr_0.V_p_2.n8 194.3
R7248 bgr_0.V_p_2.n11 bgr_0.V_p_2.n10 194.3
R7249 bgr_0.V_p_2.n0 bgr_0.V_p_2.t8 49.713
R7250 bgr_0.V_p_2.n4 bgr_0.V_p_2.t3 48.0005
R7251 bgr_0.V_p_2.n4 bgr_0.V_p_2.t10 48.0005
R7252 bgr_0.V_p_2.n5 bgr_0.V_p_2.t2 48.0005
R7253 bgr_0.V_p_2.n5 bgr_0.V_p_2.t5 48.0005
R7254 bgr_0.V_p_2.n7 bgr_0.V_p_2.t7 48.0005
R7255 bgr_0.V_p_2.n7 bgr_0.V_p_2.t9 48.0005
R7256 bgr_0.V_p_2.n8 bgr_0.V_p_2.t1 48.0005
R7257 bgr_0.V_p_2.n8 bgr_0.V_p_2.t4 48.0005
R7258 bgr_0.V_p_2.n11 bgr_0.V_p_2.t6 48.0005
R7259 bgr_0.V_p_2.t0 bgr_0.V_p_2.n11 48.0005
R7260 bgr_0.V_p_2.n0 bgr_0.V_p_2.n2 6.91717
R7261 bgr_0.V_p_2.n1 bgr_0.V_p_2.n6 6.29217
R7262 bgr_0.V_p_2.n1 bgr_0.V_p_2.n2 5.66717
R7263 bgr_0.V_p_2.n0 bgr_0.V_p_2.n3 5.66717
R7264 bgr_0.V_p_2.n1 bgr_0.V_p_2.n3 5.66717
R7265 bgr_0.V_p_2.n6 bgr_0.V_p_2.n0 5.04217
R7266 bgr_0.V_p_2.n10 bgr_0.V_p_2.n0 5.04217
R7267 bgr_0.V_p_2.n9 bgr_0.V_p_2.n0 5.04217
R7268 bgr_0.V_p_2.n1 bgr_0.V_p_2.n9 5.04217
R7269 bgr_0.V_p_2.n10 bgr_0.V_p_2.n1 5.04217
R7270 bgr_0.V_mir2.n17 bgr_0.V_mir2.t17 310.488
R7271 bgr_0.V_mir2.n14 bgr_0.V_mir2.t22 310.488
R7272 bgr_0.V_mir2.n0 bgr_0.V_mir2.t21 310.488
R7273 bgr_0.V_mir2.n5 bgr_0.V_mir2.n4 297.151
R7274 bgr_0.V_mir2.n24 bgr_0.V_mir2.n23 297.151
R7275 bgr_0.V_mir2.n27 bgr_0.V_mir2.n26 297.151
R7276 bgr_0.V_mir2.n8 bgr_0.V_mir2.t1 242.3
R7277 bgr_0.V_mir2.n7 bgr_0.V_mir2.n6 194.3
R7278 bgr_0.V_mir2.n11 bgr_0.V_mir2.n10 194.3
R7279 bgr_0.V_mir2.n19 bgr_0.V_mir2.t11 184.097
R7280 bgr_0.V_mir2.n16 bgr_0.V_mir2.t13 184.097
R7281 bgr_0.V_mir2.n2 bgr_0.V_mir2.t15 184.097
R7282 bgr_0.V_mir2.n18 bgr_0.V_mir2.n17 167.094
R7283 bgr_0.V_mir2.n15 bgr_0.V_mir2.n14 167.094
R7284 bgr_0.V_mir2.n1 bgr_0.V_mir2.n0 167.094
R7285 bgr_0.V_mir2.n20 bgr_0.V_mir2.n19 161.3
R7286 bgr_0.V_mir2.n22 bgr_0.V_mir2.n16 161.3
R7287 bgr_0.V_mir2.n3 bgr_0.V_mir2.n2 161.3
R7288 bgr_0.V_mir2.n17 bgr_0.V_mir2.t19 120.501
R7289 bgr_0.V_mir2.n18 bgr_0.V_mir2.t5 120.501
R7290 bgr_0.V_mir2.n14 bgr_0.V_mir2.t20 120.501
R7291 bgr_0.V_mir2.n15 bgr_0.V_mir2.t9 120.501
R7292 bgr_0.V_mir2.n0 bgr_0.V_mir2.t18 120.501
R7293 bgr_0.V_mir2.n1 bgr_0.V_mir2.t7 120.501
R7294 bgr_0.V_mir2.n6 bgr_0.V_mir2.t2 48.0005
R7295 bgr_0.V_mir2.n6 bgr_0.V_mir2.t0 48.0005
R7296 bgr_0.V_mir2.n10 bgr_0.V_mir2.t3 48.0005
R7297 bgr_0.V_mir2.n10 bgr_0.V_mir2.t4 48.0005
R7298 bgr_0.V_mir2.n19 bgr_0.V_mir2.n18 40.7027
R7299 bgr_0.V_mir2.n16 bgr_0.V_mir2.n15 40.7027
R7300 bgr_0.V_mir2.n2 bgr_0.V_mir2.n1 40.7027
R7301 bgr_0.V_mir2.n4 bgr_0.V_mir2.t6 39.4005
R7302 bgr_0.V_mir2.n4 bgr_0.V_mir2.t12 39.4005
R7303 bgr_0.V_mir2.n23 bgr_0.V_mir2.t10 39.4005
R7304 bgr_0.V_mir2.n23 bgr_0.V_mir2.t14 39.4005
R7305 bgr_0.V_mir2.n27 bgr_0.V_mir2.t8 39.4005
R7306 bgr_0.V_mir2.t16 bgr_0.V_mir2.n27 39.4005
R7307 bgr_0.V_mir2.n25 bgr_0.V_mir2.n5 6.89633
R7308 bgr_0.V_mir2.n26 bgr_0.V_mir2.n25 6.89633
R7309 bgr_0.V_mir2.n21 bgr_0.V_mir2.n3 6.6255
R7310 bgr_0.V_mir2.n21 bgr_0.V_mir2.n20 6.6255
R7311 bgr_0.V_mir2.n12 bgr_0.V_mir2.n8 6.22967
R7312 bgr_0.V_mir2.n9 bgr_0.V_mir2.n8 6.04217
R7313 bgr_0.V_mir2.n9 bgr_0.V_mir2.n7 6.04217
R7314 bgr_0.V_mir2.n13 bgr_0.V_mir2.n12 5.8755
R7315 bgr_0.V_mir2.n12 bgr_0.V_mir2.n11 4.85467
R7316 bgr_0.V_mir2.n25 bgr_0.V_mir2.n24 4.77133
R7317 bgr_0.V_mir2.n11 bgr_0.V_mir2.n9 4.66717
R7318 bgr_0.V_mir2.n22 bgr_0.V_mir2.n21 4.5005
R7319 bgr_0.V_mir2.n22 bgr_0.V_mir2.n13 1.7505
R7320 bgr_0.V_mir2.n13 bgr_0.V_mir2.n7 0.354667
R7321 bgr_0.V_mir2.n24 bgr_0.V_mir2.n22 0.333833
R7322 bgr_0.V_mir2.n26 bgr_0.V_mir2.n3 0.333833
R7323 bgr_0.V_mir2.n20 bgr_0.V_mir2.n5 0.333833
R7324 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.n2 443.433
R7325 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.n14 438.933
R7326 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.n10 438.933
R7327 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t24 369.534
R7328 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t20 369.534
R7329 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t27 369.534
R7330 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t11 369.534
R7331 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n16 297.151
R7332 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.n20 297.151
R7333 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.n22 297.151
R7334 bgr_0.PFET_GATE_10uA.n27 bgr_0.PFET_GATE_10uA.n26 297.151
R7335 bgr_0.PFET_GATE_10uA.n31 bgr_0.PFET_GATE_10uA.n30 289.829
R7336 bgr_0.PFET_GATE_10uA.n30 bgr_0.PFET_GATE_10uA.t10 249.034
R7337 bgr_0.PFET_GATE_10uA.n30 bgr_0.PFET_GATE_10uA.t18 249.034
R7338 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.t23 192.8
R7339 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t17 192.8
R7340 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.t29 192.8
R7341 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.t22 192.8
R7342 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t13 192.8
R7343 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.t14 192.8
R7344 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t26 192.8
R7345 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t16 192.8
R7346 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.t28 192.8
R7347 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t21 192.8
R7348 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t15 192.8
R7349 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.t12 192.8
R7350 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t25 192.8
R7351 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t19 192.8
R7352 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.n13 176.733
R7353 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n12 176.733
R7354 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.n3 176.733
R7355 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n4 176.733
R7356 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.n5 176.733
R7357 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n6 176.733
R7358 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n9 176.733
R7359 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.n8 176.733
R7360 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n7 176.733
R7361 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.n0 176.733
R7362 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n1 176.733
R7363 bgr_0.PFET_GATE_10uA.n31 bgr_0.PFET_GATE_10uA.t0 137.667
R7364 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.t3 53.1713
R7365 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.t4 39.4005
R7366 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.t6 39.4005
R7367 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.t2 39.4005
R7368 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.t9 39.4005
R7369 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.t5 39.4005
R7370 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.t7 39.4005
R7371 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.t8 39.4005
R7372 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.t1 39.4005
R7373 bgr_0.PFET_GATE_10uA.n28 bgr_0.PFET_GATE_10uA.n27 7.27133
R7374 bgr_0.PFET_GATE_10uA.n27 bgr_0.PFET_GATE_10uA.n25 7.14633
R7375 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.n21 7.14633
R7376 bgr_0.PFET_GATE_10uA.n32 bgr_0.PFET_GATE_10uA.n31 6.188
R7377 bgr_0.PFET_GATE_10uA.n33 bgr_0.PFET_GATE_10uA.n15 5.79738
R7378 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.n18 5.14633
R7379 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.n19 5.14633
R7380 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.n23 5.02133
R7381 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.n17 5.02133
R7382 bgr_0.PFET_GATE_10uA.n33 bgr_0.PFET_GATE_10uA.n32 4.90675
R7383 bgr_0.PFET_GATE_10uA.n29 bgr_0.PFET_GATE_10uA.n28 4.5005
R7384 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.n11 4.2505
R7385 bgr_0.PFET_GATE_10uA.n28 bgr_0.PFET_GATE_10uA.n18 2.1255
R7386 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.n18 2.1255
R7387 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.n24 2.1255
R7388 bgr_0.PFET_GATE_10uA.n29 bgr_0.PFET_GATE_10uA.n17 0.646333
R7389 bgr_0.PFET_GATE_10uA.n32 bgr_0.PFET_GATE_10uA.n29 0.53175
R7390 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n33 0.063
R7391 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.n15 634.533
R7392 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.t8 449.868
R7393 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.t2 449.868
R7394 two_stage_opamp_dummy_magic_0.Vb1.n26 two_stage_opamp_dummy_magic_0.Vb1.t24 449.868
R7395 two_stage_opamp_dummy_magic_0.Vb1.n35 two_stage_opamp_dummy_magic_0.Vb1.n25 306.173
R7396 two_stage_opamp_dummy_magic_0.Vb1.n35 two_stage_opamp_dummy_magic_0.Vb1.n34 305.485
R7397 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.n2 299.861
R7398 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.n3 299.586
R7399 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.t4 273.134
R7400 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.t6 273.134
R7401 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.t27 273.134
R7402 two_stage_opamp_dummy_magic_0.Vb1.n25 two_stage_opamp_dummy_magic_0.Vb1.t23 273.134
R7403 two_stage_opamp_dummy_magic_0.Vb1.n34 two_stage_opamp_dummy_magic_0.Vb1.t28 273.134
R7404 two_stage_opamp_dummy_magic_0.Vb1.n26 two_stage_opamp_dummy_magic_0.Vb1.t34 273.134
R7405 two_stage_opamp_dummy_magic_0.Vb1.n27 two_stage_opamp_dummy_magic_0.Vb1.t22 273.134
R7406 two_stage_opamp_dummy_magic_0.Vb1.n28 two_stage_opamp_dummy_magic_0.Vb1.t31 273.134
R7407 two_stage_opamp_dummy_magic_0.Vb1.n29 two_stage_opamp_dummy_magic_0.Vb1.t19 273.134
R7408 two_stage_opamp_dummy_magic_0.Vb1.n30 two_stage_opamp_dummy_magic_0.Vb1.t16 273.134
R7409 two_stage_opamp_dummy_magic_0.Vb1.n31 two_stage_opamp_dummy_magic_0.Vb1.t20 273.134
R7410 two_stage_opamp_dummy_magic_0.Vb1.n32 two_stage_opamp_dummy_magic_0.Vb1.t29 273.134
R7411 two_stage_opamp_dummy_magic_0.Vb1.n33 two_stage_opamp_dummy_magic_0.Vb1.t18 273.134
R7412 two_stage_opamp_dummy_magic_0.Vb1.n24 two_stage_opamp_dummy_magic_0.Vb1.t32 273.134
R7413 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.t21 273.134
R7414 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.t30 273.134
R7415 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.t26 273.134
R7416 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.t15 273.134
R7417 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.t25 273.134
R7418 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.t14 273.134
R7419 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.t17 273.134
R7420 two_stage_opamp_dummy_magic_0.Vb1.n34 two_stage_opamp_dummy_magic_0.Vb1.n33 176.733
R7421 two_stage_opamp_dummy_magic_0.Vb1.n33 two_stage_opamp_dummy_magic_0.Vb1.n32 176.733
R7422 two_stage_opamp_dummy_magic_0.Vb1.n32 two_stage_opamp_dummy_magic_0.Vb1.n31 176.733
R7423 two_stage_opamp_dummy_magic_0.Vb1.n31 two_stage_opamp_dummy_magic_0.Vb1.n30 176.733
R7424 two_stage_opamp_dummy_magic_0.Vb1.n30 two_stage_opamp_dummy_magic_0.Vb1.n29 176.733
R7425 two_stage_opamp_dummy_magic_0.Vb1.n29 two_stage_opamp_dummy_magic_0.Vb1.n28 176.733
R7426 two_stage_opamp_dummy_magic_0.Vb1.n28 two_stage_opamp_dummy_magic_0.Vb1.n27 176.733
R7427 two_stage_opamp_dummy_magic_0.Vb1.n27 two_stage_opamp_dummy_magic_0.Vb1.n26 176.733
R7428 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.n16 176.733
R7429 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.n17 176.733
R7430 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.n18 176.733
R7431 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.n19 176.733
R7432 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.n20 176.733
R7433 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.n21 176.733
R7434 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.n22 176.733
R7435 two_stage_opamp_dummy_magic_0.Vb1.n24 two_stage_opamp_dummy_magic_0.Vb1.n23 176.733
R7436 two_stage_opamp_dummy_magic_0.Vb1.n25 two_stage_opamp_dummy_magic_0.Vb1.n24 176.733
R7437 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.t33 165.8
R7438 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.n9 161.3
R7439 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb1.n35 54.8755
R7440 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.n12 49.3505
R7441 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.n10 49.3505
R7442 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.n5 49.3505
R7443 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.n8 45.5227
R7444 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.n7 45.5227
R7445 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.t1 39.4005
R7446 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.t13 39.4005
R7447 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t12 39.4005
R7448 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t0 39.4005
R7449 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.t10 16.0005
R7450 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.t3 16.0005
R7451 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.t7 16.0005
R7452 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.t5 16.0005
R7453 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.t9 16.0005
R7454 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.t11 16.0005
R7455 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb1.n4 13.4872
R7456 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.n11 5.6255
R7457 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.n6 5.6255
R7458 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.n0 5.5005
R7459 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.n1 5.063
R7460 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.n13 4.938
R7461 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.n0 4.938
R7462 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.n14 1.96925
R7463 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.n0 0.563
R7464 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.n25 594.301
R7465 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.n26 594.301
R7466 two_stage_opamp_dummy_magic_0.V_err_gate.n29 two_stage_opamp_dummy_magic_0.V_err_gate.n28 594.301
R7467 two_stage_opamp_dummy_magic_0.V_err_gate.n31 two_stage_opamp_dummy_magic_0.V_err_gate.n30 594.301
R7468 two_stage_opamp_dummy_magic_0.V_err_gate.n33 two_stage_opamp_dummy_magic_0.V_err_gate.n32 594.301
R7469 two_stage_opamp_dummy_magic_0.V_err_gate.n35 two_stage_opamp_dummy_magic_0.V_err_gate.n34 594.301
R7470 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n24 571
R7471 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.t14 289.2
R7472 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.t22 289.2
R7473 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.n7 176.733
R7474 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.n8 176.733
R7475 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.n9 176.733
R7476 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.n10 176.733
R7477 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.n11 176.733
R7478 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.n12 176.733
R7479 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.n13 176.733
R7480 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.n14 176.733
R7481 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.n15 176.733
R7482 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.n16 176.733
R7483 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.n23 176.733
R7484 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.n22 176.733
R7485 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.n21 176.733
R7486 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.n20 176.733
R7487 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.n19 176.733
R7488 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.n18 176.733
R7489 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.n17 176.733
R7490 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n6 138.577
R7491 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.t30 112.468
R7492 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.t25 112.468
R7493 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.t31 112.468
R7494 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.t24 112.468
R7495 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.t16 112.468
R7496 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.t27 112.468
R7497 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.t18 112.468
R7498 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.t29 112.468
R7499 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.t20 112.468
R7500 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.t33 112.468
R7501 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.t23 112.468
R7502 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.t21 112.468
R7503 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.t15 112.468
R7504 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.t26 112.468
R7505 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.t17 112.468
R7506 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.t28 112.468
R7507 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.t19 112.468
R7508 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.t32 112.468
R7509 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate.t4 78.8005
R7510 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate.t8 78.8005
R7511 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate.t13 78.8005
R7512 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate.t0 78.8005
R7513 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.t5 78.8005
R7514 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.t3 78.8005
R7515 two_stage_opamp_dummy_magic_0.V_err_gate.n30 two_stage_opamp_dummy_magic_0.V_err_gate.t11 78.8005
R7516 two_stage_opamp_dummy_magic_0.V_err_gate.n30 two_stage_opamp_dummy_magic_0.V_err_gate.t12 78.8005
R7517 two_stage_opamp_dummy_magic_0.V_err_gate.n32 two_stage_opamp_dummy_magic_0.V_err_gate.t6 78.8005
R7518 two_stage_opamp_dummy_magic_0.V_err_gate.n32 two_stage_opamp_dummy_magic_0.V_err_gate.t2 78.8005
R7519 two_stage_opamp_dummy_magic_0.V_err_gate.n34 two_stage_opamp_dummy_magic_0.V_err_gate.t7 78.8005
R7520 two_stage_opamp_dummy_magic_0.V_err_gate.n34 two_stage_opamp_dummy_magic_0.V_err_gate.t1 78.8005
R7521 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.t9 24.0005
R7522 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.t10 24.0005
R7523 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n3 6.8755
R7524 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.n2 5.41717
R7525 two_stage_opamp_dummy_magic_0.V_err_gate.n35 two_stage_opamp_dummy_magic_0.V_err_gate.n1 5.22967
R7526 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n2 5.22967
R7527 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.n27 4.85467
R7528 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.n29 4.85467
R7529 two_stage_opamp_dummy_magic_0.V_err_gate.n31 two_stage_opamp_dummy_magic_0.V_err_gate.n5 4.85467
R7530 two_stage_opamp_dummy_magic_0.V_err_gate.n33 two_stage_opamp_dummy_magic_0.V_err_gate.n3 4.85467
R7531 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.n35 4.85467
R7532 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.n0 4.66717
R7533 two_stage_opamp_dummy_magic_0.V_err_gate.n29 two_stage_opamp_dummy_magic_0.V_err_gate.n0 4.66717
R7534 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n31 4.66717
R7535 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n33 4.66717
R7536 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n0 1.688
R7537 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.n3 1.1255
R7538 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.n4 1.1255
R7539 two_stage_opamp_dummy_magic_0.V_err_p.n20 two_stage_opamp_dummy_magic_0.V_err_p.n19 594.301
R7540 two_stage_opamp_dummy_magic_0.V_err_p.n23 two_stage_opamp_dummy_magic_0.V_err_p.n22 594.301
R7541 two_stage_opamp_dummy_magic_0.V_err_p.n26 two_stage_opamp_dummy_magic_0.V_err_p.n25 594.301
R7542 two_stage_opamp_dummy_magic_0.V_err_p.n30 two_stage_opamp_dummy_magic_0.V_err_p.n29 594.301
R7543 two_stage_opamp_dummy_magic_0.V_err_p.n33 two_stage_opamp_dummy_magic_0.V_err_p.n32 594.301
R7544 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.n1 594.301
R7545 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n4 594.301
R7546 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.n7 594.301
R7547 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n10 594.301
R7548 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n14 594.301
R7549 two_stage_opamp_dummy_magic_0.V_err_p.n37 two_stage_opamp_dummy_magic_0.V_err_p.n36 594.301
R7550 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.t15 78.8005
R7551 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.t7 78.8005
R7552 two_stage_opamp_dummy_magic_0.V_err_p.n22 two_stage_opamp_dummy_magic_0.V_err_p.t18 78.8005
R7553 two_stage_opamp_dummy_magic_0.V_err_p.n22 two_stage_opamp_dummy_magic_0.V_err_p.t13 78.8005
R7554 two_stage_opamp_dummy_magic_0.V_err_p.n25 two_stage_opamp_dummy_magic_0.V_err_p.t11 78.8005
R7555 two_stage_opamp_dummy_magic_0.V_err_p.n25 two_stage_opamp_dummy_magic_0.V_err_p.t16 78.8005
R7556 two_stage_opamp_dummy_magic_0.V_err_p.n29 two_stage_opamp_dummy_magic_0.V_err_p.t12 78.8005
R7557 two_stage_opamp_dummy_magic_0.V_err_p.n29 two_stage_opamp_dummy_magic_0.V_err_p.t17 78.8005
R7558 two_stage_opamp_dummy_magic_0.V_err_p.n32 two_stage_opamp_dummy_magic_0.V_err_p.t14 78.8005
R7559 two_stage_opamp_dummy_magic_0.V_err_p.n32 two_stage_opamp_dummy_magic_0.V_err_p.t19 78.8005
R7560 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t2 78.8005
R7561 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t9 78.8005
R7562 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t6 78.8005
R7563 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t21 78.8005
R7564 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.t1 78.8005
R7565 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.t4 78.8005
R7566 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.t5 78.8005
R7567 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.t0 78.8005
R7568 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t10 78.8005
R7569 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t3 78.8005
R7570 two_stage_opamp_dummy_magic_0.V_err_p.n37 two_stage_opamp_dummy_magic_0.V_err_p.t8 78.8005
R7571 two_stage_opamp_dummy_magic_0.V_err_p.t20 two_stage_opamp_dummy_magic_0.V_err_p.n37 78.8005
R7572 two_stage_opamp_dummy_magic_0.V_err_p.n35 two_stage_opamp_dummy_magic_0.V_err_p.n17 7.188
R7573 two_stage_opamp_dummy_magic_0.V_err_p.n36 two_stage_opamp_dummy_magic_0.V_err_p.n0 6.10467
R7574 two_stage_opamp_dummy_magic_0.V_err_p.n24 two_stage_opamp_dummy_magic_0.V_err_p.n20 6.10467
R7575 two_stage_opamp_dummy_magic_0.V_err_p.n21 two_stage_opamp_dummy_magic_0.V_err_p.n20 5.91717
R7576 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.n5 5.41717
R7577 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n5 5.22967
R7578 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.n2 5.22967
R7579 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n16 5.063
R7580 two_stage_opamp_dummy_magic_0.V_err_p.n24 two_stage_opamp_dummy_magic_0.V_err_p.n23 4.85467
R7581 two_stage_opamp_dummy_magic_0.V_err_p.n27 two_stage_opamp_dummy_magic_0.V_err_p.n26 4.85467
R7582 two_stage_opamp_dummy_magic_0.V_err_p.n30 two_stage_opamp_dummy_magic_0.V_err_p.n28 4.85467
R7583 two_stage_opamp_dummy_magic_0.V_err_p.n33 two_stage_opamp_dummy_magic_0.V_err_p.n0 4.85467
R7584 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.n6 4.85467
R7585 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n3 4.85467
R7586 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.n15 4.85467
R7587 two_stage_opamp_dummy_magic_0.V_err_p.n23 two_stage_opamp_dummy_magic_0.V_err_p.n21 4.66717
R7588 two_stage_opamp_dummy_magic_0.V_err_p.n26 two_stage_opamp_dummy_magic_0.V_err_p.n18 4.66717
R7589 two_stage_opamp_dummy_magic_0.V_err_p.n31 two_stage_opamp_dummy_magic_0.V_err_p.n30 4.66717
R7590 two_stage_opamp_dummy_magic_0.V_err_p.n34 two_stage_opamp_dummy_magic_0.V_err_p.n33 4.66717
R7591 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n8 4.66717
R7592 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n11 4.66717
R7593 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n13 4.66717
R7594 two_stage_opamp_dummy_magic_0.V_err_p.n36 two_stage_opamp_dummy_magic_0.V_err_p.n35 4.66717
R7595 two_stage_opamp_dummy_magic_0.V_err_p.n28 two_stage_opamp_dummy_magic_0.V_err_p.n0 1.2505
R7596 two_stage_opamp_dummy_magic_0.V_err_p.n28 two_stage_opamp_dummy_magic_0.V_err_p.n27 1.2505
R7597 two_stage_opamp_dummy_magic_0.V_err_p.n27 two_stage_opamp_dummy_magic_0.V_err_p.n24 1.2505
R7598 two_stage_opamp_dummy_magic_0.V_err_p.n21 two_stage_opamp_dummy_magic_0.V_err_p.n18 1.2505
R7599 two_stage_opamp_dummy_magic_0.V_err_p.n31 two_stage_opamp_dummy_magic_0.V_err_p.n18 1.2505
R7600 two_stage_opamp_dummy_magic_0.V_err_p.n34 two_stage_opamp_dummy_magic_0.V_err_p.n31 1.2505
R7601 two_stage_opamp_dummy_magic_0.V_err_p.n35 two_stage_opamp_dummy_magic_0.V_err_p.n34 1.2505
R7602 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.n3 0.563
R7603 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.n3 0.563
R7604 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n9 0.563
R7605 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.n12 0.563
R7606 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n2 0.354667
R7607 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.t41 1172.87
R7608 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.t34 1172.87
R7609 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.t32 996.134
R7610 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.t26 996.134
R7611 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.t43 996.134
R7612 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.t28 996.134
R7613 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.t47 996.134
R7614 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.t50 996.134
R7615 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.t35 996.134
R7616 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.t49 996.134
R7617 two_stage_opamp_dummy_magic_0.X.n63 two_stage_opamp_dummy_magic_0.X.t30 690.867
R7618 two_stage_opamp_dummy_magic_0.X.n59 two_stage_opamp_dummy_magic_0.X.t37 690.867
R7619 two_stage_opamp_dummy_magic_0.X.n51 two_stage_opamp_dummy_magic_0.X.t44 530.201
R7620 two_stage_opamp_dummy_magic_0.X.n55 two_stage_opamp_dummy_magic_0.X.t38 530.201
R7621 two_stage_opamp_dummy_magic_0.X.n66 two_stage_opamp_dummy_magic_0.X.t27 514.134
R7622 two_stage_opamp_dummy_magic_0.X.n63 two_stage_opamp_dummy_magic_0.X.t45 514.134
R7623 two_stage_opamp_dummy_magic_0.X.n64 two_stage_opamp_dummy_magic_0.X.t31 514.134
R7624 two_stage_opamp_dummy_magic_0.X.n65 two_stage_opamp_dummy_magic_0.X.t46 514.134
R7625 two_stage_opamp_dummy_magic_0.X.n62 two_stage_opamp_dummy_magic_0.X.t42 514.134
R7626 two_stage_opamp_dummy_magic_0.X.n61 two_stage_opamp_dummy_magic_0.X.t25 514.134
R7627 two_stage_opamp_dummy_magic_0.X.n60 two_stage_opamp_dummy_magic_0.X.t40 514.134
R7628 two_stage_opamp_dummy_magic_0.X.n59 two_stage_opamp_dummy_magic_0.X.t54 514.134
R7629 two_stage_opamp_dummy_magic_0.X.n67 two_stage_opamp_dummy_magic_0.X.n58 473.967
R7630 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.n28 446.967
R7631 two_stage_opamp_dummy_magic_0.X.n67 two_stage_opamp_dummy_magic_0.X.n66 441.834
R7632 two_stage_opamp_dummy_magic_0.X.n58 two_stage_opamp_dummy_magic_0.X.t36 353.467
R7633 two_stage_opamp_dummy_magic_0.X.n51 two_stage_opamp_dummy_magic_0.X.t29 353.467
R7634 two_stage_opamp_dummy_magic_0.X.n52 two_stage_opamp_dummy_magic_0.X.t48 353.467
R7635 two_stage_opamp_dummy_magic_0.X.n53 two_stage_opamp_dummy_magic_0.X.t33 353.467
R7636 two_stage_opamp_dummy_magic_0.X.n54 two_stage_opamp_dummy_magic_0.X.t51 353.467
R7637 two_stage_opamp_dummy_magic_0.X.n57 two_stage_opamp_dummy_magic_0.X.t53 353.467
R7638 two_stage_opamp_dummy_magic_0.X.n56 two_stage_opamp_dummy_magic_0.X.t39 353.467
R7639 two_stage_opamp_dummy_magic_0.X.n55 two_stage_opamp_dummy_magic_0.X.t52 353.467
R7640 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.n21 176.733
R7641 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.n22 176.733
R7642 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.n23 176.733
R7643 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.n24 176.733
R7644 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.n27 176.733
R7645 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.n26 176.733
R7646 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.n25 176.733
R7647 two_stage_opamp_dummy_magic_0.X.n52 two_stage_opamp_dummy_magic_0.X.n51 176.733
R7648 two_stage_opamp_dummy_magic_0.X.n53 two_stage_opamp_dummy_magic_0.X.n52 176.733
R7649 two_stage_opamp_dummy_magic_0.X.n54 two_stage_opamp_dummy_magic_0.X.n53 176.733
R7650 two_stage_opamp_dummy_magic_0.X.n58 two_stage_opamp_dummy_magic_0.X.n54 176.733
R7651 two_stage_opamp_dummy_magic_0.X.n58 two_stage_opamp_dummy_magic_0.X.n57 176.733
R7652 two_stage_opamp_dummy_magic_0.X.n57 two_stage_opamp_dummy_magic_0.X.n56 176.733
R7653 two_stage_opamp_dummy_magic_0.X.n56 two_stage_opamp_dummy_magic_0.X.n55 176.733
R7654 two_stage_opamp_dummy_magic_0.X.n60 two_stage_opamp_dummy_magic_0.X.n59 176.733
R7655 two_stage_opamp_dummy_magic_0.X.n61 two_stage_opamp_dummy_magic_0.X.n60 176.733
R7656 two_stage_opamp_dummy_magic_0.X.n62 two_stage_opamp_dummy_magic_0.X.n61 176.733
R7657 two_stage_opamp_dummy_magic_0.X.n66 two_stage_opamp_dummy_magic_0.X.n62 176.733
R7658 two_stage_opamp_dummy_magic_0.X.n66 two_stage_opamp_dummy_magic_0.X.n65 176.733
R7659 two_stage_opamp_dummy_magic_0.X.n65 two_stage_opamp_dummy_magic_0.X.n64 176.733
R7660 two_stage_opamp_dummy_magic_0.X.n64 two_stage_opamp_dummy_magic_0.X.n63 176.733
R7661 two_stage_opamp_dummy_magic_0.X.n68 two_stage_opamp_dummy_magic_0.X.n67 176.238
R7662 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.n32 66.0338
R7663 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.n35 66.0338
R7664 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.n38 66.0338
R7665 two_stage_opamp_dummy_magic_0.X.n43 two_stage_opamp_dummy_magic_0.X.n42 66.0338
R7666 two_stage_opamp_dummy_magic_0.X.n46 two_stage_opamp_dummy_magic_0.X.n45 66.0338
R7667 two_stage_opamp_dummy_magic_0.X.n49 two_stage_opamp_dummy_magic_0.X.n48 66.0338
R7668 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.t11 49.9898
R7669 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.n0 49.3505
R7670 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.n4 49.3505
R7671 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.n6 49.3505
R7672 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.n10 49.3505
R7673 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.n12 49.3505
R7674 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.n16 49.3505
R7675 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t16 16.0005
R7676 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t17 16.0005
R7677 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.t22 16.0005
R7678 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.t20 16.0005
R7679 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.t13 16.0005
R7680 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.t14 16.0005
R7681 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.t15 16.0005
R7682 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.t23 16.0005
R7683 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.t18 16.0005
R7684 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.t12 16.0005
R7685 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.t19 16.0005
R7686 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.t21 16.0005
R7687 two_stage_opamp_dummy_magic_0.X.n68 two_stage_opamp_dummy_magic_0.X.n50 12.7193
R7688 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.t4 11.2576
R7689 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.t24 11.2576
R7690 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.t3 11.2576
R7691 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.t2 11.2576
R7692 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.t6 11.2576
R7693 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.t1 11.2576
R7694 two_stage_opamp_dummy_magic_0.X.n42 two_stage_opamp_dummy_magic_0.X.t9 11.2576
R7695 two_stage_opamp_dummy_magic_0.X.n42 two_stage_opamp_dummy_magic_0.X.t0 11.2576
R7696 two_stage_opamp_dummy_magic_0.X.n45 two_stage_opamp_dummy_magic_0.X.t7 11.2576
R7697 two_stage_opamp_dummy_magic_0.X.n45 two_stage_opamp_dummy_magic_0.X.t8 11.2576
R7698 two_stage_opamp_dummy_magic_0.X.n48 two_stage_opamp_dummy_magic_0.X.t10 11.2576
R7699 two_stage_opamp_dummy_magic_0.X.n48 two_stage_opamp_dummy_magic_0.X.t5 11.2576
R7700 two_stage_opamp_dummy_magic_0.X.n70 two_stage_opamp_dummy_magic_0.X.n69 8.09425
R7701 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.n33 6.10467
R7702 two_stage_opamp_dummy_magic_0.X.n49 two_stage_opamp_dummy_magic_0.X.n47 5.91717
R7703 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.n33 5.91717
R7704 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.n11 5.6255
R7705 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.n5 5.6255
R7706 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.n36 5.47967
R7707 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n39 5.47967
R7708 two_stage_opamp_dummy_magic_0.X.n43 two_stage_opamp_dummy_magic_0.X.n41 5.47967
R7709 two_stage_opamp_dummy_magic_0.X.n46 two_stage_opamp_dummy_magic_0.X.n30 5.47967
R7710 two_stage_opamp_dummy_magic_0.X.n50 two_stage_opamp_dummy_magic_0.X.n49 5.47967
R7711 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.n3 5.438
R7712 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.n2 5.438
R7713 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.n34 5.29217
R7714 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.n31 5.29217
R7715 two_stage_opamp_dummy_magic_0.X.n44 two_stage_opamp_dummy_magic_0.X.n43 5.29217
R7716 two_stage_opamp_dummy_magic_0.X.n47 two_stage_opamp_dummy_magic_0.X.n46 5.29217
R7717 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.n7 5.063
R7718 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.n13 5.063
R7719 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.n15 5.063
R7720 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.n1 5.063
R7721 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.n2 4.8755
R7722 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.n3 4.8755
R7723 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.n17 4.8755
R7724 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.n19 4.5005
R7725 two_stage_opamp_dummy_magic_0.X.n69 two_stage_opamp_dummy_magic_0.X.n68 4.5005
R7726 two_stage_opamp_dummy_magic_0.X.n70 two_stage_opamp_dummy_magic_0.X.n20 2.46925
R7727 two_stage_opamp_dummy_magic_0.X.n69 two_stage_opamp_dummy_magic_0.X.n29 2.3755
R7728 two_stage_opamp_dummy_magic_0.X.n47 two_stage_opamp_dummy_magic_0.X.n44 0.6255
R7729 two_stage_opamp_dummy_magic_0.X.n44 two_stage_opamp_dummy_magic_0.X.n31 0.6255
R7730 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.n31 0.6255
R7731 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n37 0.6255
R7732 two_stage_opamp_dummy_magic_0.X.n41 two_stage_opamp_dummy_magic_0.X.n40 0.6255
R7733 two_stage_opamp_dummy_magic_0.X.n41 two_stage_opamp_dummy_magic_0.X.n30 0.6255
R7734 two_stage_opamp_dummy_magic_0.X.n50 two_stage_opamp_dummy_magic_0.X.n30 0.6255
R7735 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.n9 0.563
R7736 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.n14 0.563
R7737 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.n3 0.563
R7738 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n18 0.563
R7739 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n2 0.563
R7740 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.n8 0.563
R7741 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.n1 0.3755
R7742 two_stage_opamp_dummy_magic_0.X two_stage_opamp_dummy_magic_0.X.n70 0.063
R7743 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n1 49.3505
R7744 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.n4 49.3505
R7745 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.n6 49.3505
R7746 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n10 49.3505
R7747 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.n14 49.3505
R7748 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n17 49.3505
R7749 two_stage_opamp_dummy_magic_0.VD1.n21 two_stage_opamp_dummy_magic_0.VD1.n20 49.3505
R7750 two_stage_opamp_dummy_magic_0.VD1.n24 two_stage_opamp_dummy_magic_0.VD1.n23 49.3505
R7751 two_stage_opamp_dummy_magic_0.VD1.n26 two_stage_opamp_dummy_magic_0.VD1.n25 49.3505
R7752 two_stage_opamp_dummy_magic_0.VD1.n30 two_stage_opamp_dummy_magic_0.VD1.n29 49.3505
R7753 two_stage_opamp_dummy_magic_0.VD1.n37 two_stage_opamp_dummy_magic_0.VD1.n36 49.3505
R7754 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t7 16.0005
R7755 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t12 16.0005
R7756 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t5 16.0005
R7757 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t10 16.0005
R7758 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.t6 16.0005
R7759 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.t11 16.0005
R7760 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.t13 16.0005
R7761 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.t8 16.0005
R7762 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.t19 16.0005
R7763 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.t16 16.0005
R7764 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t20 16.0005
R7765 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t3 16.0005
R7766 two_stage_opamp_dummy_magic_0.VD1.n20 two_stage_opamp_dummy_magic_0.VD1.t2 16.0005
R7767 two_stage_opamp_dummy_magic_0.VD1.n20 two_stage_opamp_dummy_magic_0.VD1.t17 16.0005
R7768 two_stage_opamp_dummy_magic_0.VD1.n23 two_stage_opamp_dummy_magic_0.VD1.t1 16.0005
R7769 two_stage_opamp_dummy_magic_0.VD1.n23 two_stage_opamp_dummy_magic_0.VD1.t18 16.0005
R7770 two_stage_opamp_dummy_magic_0.VD1.n25 two_stage_opamp_dummy_magic_0.VD1.t21 16.0005
R7771 two_stage_opamp_dummy_magic_0.VD1.n25 two_stage_opamp_dummy_magic_0.VD1.t0 16.0005
R7772 two_stage_opamp_dummy_magic_0.VD1.n29 two_stage_opamp_dummy_magic_0.VD1.t15 16.0005
R7773 two_stage_opamp_dummy_magic_0.VD1.n29 two_stage_opamp_dummy_magic_0.VD1.t4 16.0005
R7774 two_stage_opamp_dummy_magic_0.VD1.t14 two_stage_opamp_dummy_magic_0.VD1.n37 16.0005
R7775 two_stage_opamp_dummy_magic_0.VD1.n37 two_stage_opamp_dummy_magic_0.VD1.t9 16.0005
R7776 two_stage_opamp_dummy_magic_0.VD1.n33 two_stage_opamp_dummy_magic_0.VD1.n32 5.77133
R7777 two_stage_opamp_dummy_magic_0.VD1.n24 two_stage_opamp_dummy_magic_0.VD1.n13 5.64633
R7778 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n15 5.64633
R7779 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.n5 5.6255
R7780 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n0 5.6255
R7781 two_stage_opamp_dummy_magic_0.VD1.n27 two_stage_opamp_dummy_magic_0.VD1.n24 5.438
R7782 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.n15 5.438
R7783 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.n3 5.438
R7784 two_stage_opamp_dummy_magic_0.VD1.n35 two_stage_opamp_dummy_magic_0.VD1.n2 5.438
R7785 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n16 5.08383
R7786 two_stage_opamp_dummy_magic_0.VD1.n21 two_stage_opamp_dummy_magic_0.VD1.n12 5.08383
R7787 two_stage_opamp_dummy_magic_0.VD1.n26 two_stage_opamp_dummy_magic_0.VD1.n13 5.08383
R7788 two_stage_opamp_dummy_magic_0.VD1.n31 two_stage_opamp_dummy_magic_0.VD1.n30 5.08383
R7789 two_stage_opamp_dummy_magic_0.VD1.n36 two_stage_opamp_dummy_magic_0.VD1.n0 5.063
R7790 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.n7 5.063
R7791 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n9 5.063
R7792 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.n3 4.8755
R7793 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.n18 4.8755
R7794 two_stage_opamp_dummy_magic_0.VD1.n22 two_stage_opamp_dummy_magic_0.VD1.n21 4.8755
R7795 two_stage_opamp_dummy_magic_0.VD1.n27 two_stage_opamp_dummy_magic_0.VD1.n26 4.8755
R7796 two_stage_opamp_dummy_magic_0.VD1.n30 two_stage_opamp_dummy_magic_0.VD1.n28 4.8755
R7797 two_stage_opamp_dummy_magic_0.VD1.n36 two_stage_opamp_dummy_magic_0.VD1.n35 4.8755
R7798 two_stage_opamp_dummy_magic_0.VD1.n34 two_stage_opamp_dummy_magic_0.VD1.n33 4.5005
R7799 two_stage_opamp_dummy_magic_0.VD1.n31 two_stage_opamp_dummy_magic_0.VD1.n13 0.563
R7800 two_stage_opamp_dummy_magic_0.VD1.n28 two_stage_opamp_dummy_magic_0.VD1.n27 0.563
R7801 two_stage_opamp_dummy_magic_0.VD1.n28 two_stage_opamp_dummy_magic_0.VD1.n22 0.563
R7802 two_stage_opamp_dummy_magic_0.VD1.n22 two_stage_opamp_dummy_magic_0.VD1.n19 0.563
R7803 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n12 0.563
R7804 two_stage_opamp_dummy_magic_0.VD1.n35 two_stage_opamp_dummy_magic_0.VD1.n34 0.563
R7805 two_stage_opamp_dummy_magic_0.VD1.n34 two_stage_opamp_dummy_magic_0.VD1.n3 0.563
R7806 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.n8 0.563
R7807 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.n0 0.563
R7808 two_stage_opamp_dummy_magic_0.VD1.n33 two_stage_opamp_dummy_magic_0.VD1.n11 0.3755
R7809 two_stage_opamp_dummy_magic_0.VD1.n32 two_stage_opamp_dummy_magic_0.VD1.n31 0.234875
R7810 two_stage_opamp_dummy_magic_0.VD1.n32 two_stage_opamp_dummy_magic_0.VD1.n12 0.234875
R7811 a_6930_22564.t0 a_6930_22564.t1 178.133
R7812 two_stage_opamp_dummy_magic_0.cap_res_X.t0 two_stage_opamp_dummy_magic_0.cap_res_X.t6 50.1603
R7813 two_stage_opamp_dummy_magic_0.cap_res_X.t23 two_stage_opamp_dummy_magic_0.cap_res_X.t62 0.1603
R7814 two_stage_opamp_dummy_magic_0.cap_res_X.t46 two_stage_opamp_dummy_magic_0.cap_res_X.t87 0.1603
R7815 two_stage_opamp_dummy_magic_0.cap_res_X.t10 two_stage_opamp_dummy_magic_0.cap_res_X.t47 0.1603
R7816 two_stage_opamp_dummy_magic_0.cap_res_X.t112 two_stage_opamp_dummy_magic_0.cap_res_X.t12 0.1603
R7817 two_stage_opamp_dummy_magic_0.cap_res_X.t77 two_stage_opamp_dummy_magic_0.cap_res_X.t92 0.1603
R7818 two_stage_opamp_dummy_magic_0.cap_res_X.t114 two_stage_opamp_dummy_magic_0.cap_res_X.t77 0.1603
R7819 two_stage_opamp_dummy_magic_0.cap_res_X.t72 two_stage_opamp_dummy_magic_0.cap_res_X.t114 0.1603
R7820 two_stage_opamp_dummy_magic_0.cap_res_X.t101 two_stage_opamp_dummy_magic_0.cap_res_X.t39 0.1603
R7821 two_stage_opamp_dummy_magic_0.cap_res_X.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t101 0.1603
R7822 two_stage_opamp_dummy_magic_0.cap_res_X.t96 two_stage_opamp_dummy_magic_0.cap_res_X.t136 0.1603
R7823 two_stage_opamp_dummy_magic_0.cap_res_X.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t90 0.1603
R7824 two_stage_opamp_dummy_magic_0.cap_res_X.t88 two_stage_opamp_dummy_magic_0.cap_res_X.t49 0.1603
R7825 two_stage_opamp_dummy_magic_0.cap_res_X.t42 two_stage_opamp_dummy_magic_0.cap_res_X.t81 0.1603
R7826 two_stage_opamp_dummy_magic_0.cap_res_X.t27 two_stage_opamp_dummy_magic_0.cap_res_X.t130 0.1603
R7827 two_stage_opamp_dummy_magic_0.cap_res_X.t9 two_stage_opamp_dummy_magic_0.cap_res_X.t45 0.1603
R7828 two_stage_opamp_dummy_magic_0.cap_res_X.t134 two_stage_opamp_dummy_magic_0.cap_res_X.t95 0.1603
R7829 two_stage_opamp_dummy_magic_0.cap_res_X.t25 two_stage_opamp_dummy_magic_0.cap_res_X.t58 0.1603
R7830 two_stage_opamp_dummy_magic_0.cap_res_X.t79 two_stage_opamp_dummy_magic_0.cap_res_X.t43 0.1603
R7831 two_stage_opamp_dummy_magic_0.cap_res_X.t65 two_stage_opamp_dummy_magic_0.cap_res_X.t102 0.1603
R7832 two_stage_opamp_dummy_magic_0.cap_res_X.t118 two_stage_opamp_dummy_magic_0.cap_res_X.t83 0.1603
R7833 two_stage_opamp_dummy_magic_0.cap_res_X.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t66 0.1603
R7834 two_stage_opamp_dummy_magic_0.cap_res_X.t86 two_stage_opamp_dummy_magic_0.cap_res_X.t48 0.1603
R7835 two_stage_opamp_dummy_magic_0.cap_res_X.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t105 0.1603
R7836 two_stage_opamp_dummy_magic_0.cap_res_X.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t89 0.1603
R7837 two_stage_opamp_dummy_magic_0.cap_res_X.t109 two_stage_opamp_dummy_magic_0.cap_res_X.t4 0.1603
R7838 two_stage_opamp_dummy_magic_0.cap_res_X.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t128 0.1603
R7839 two_stage_opamp_dummy_magic_0.cap_res_X.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t111 0.1603
R7840 two_stage_opamp_dummy_magic_0.cap_res_X.t129 two_stage_opamp_dummy_magic_0.cap_res_X.t94 0.1603
R7841 two_stage_opamp_dummy_magic_0.cap_res_X.t117 two_stage_opamp_dummy_magic_0.cap_res_X.t11 0.1603
R7842 two_stage_opamp_dummy_magic_0.cap_res_X.t28 two_stage_opamp_dummy_magic_0.cap_res_X.t135 0.1603
R7843 two_stage_opamp_dummy_magic_0.cap_res_X.t16 two_stage_opamp_dummy_magic_0.cap_res_X.t50 0.1603
R7844 two_stage_opamp_dummy_magic_0.cap_res_X.t68 two_stage_opamp_dummy_magic_0.cap_res_X.t34 0.1603
R7845 two_stage_opamp_dummy_magic_0.cap_res_X.t54 two_stage_opamp_dummy_magic_0.cap_res_X.t91 0.1603
R7846 two_stage_opamp_dummy_magic_0.cap_res_X.t108 two_stage_opamp_dummy_magic_0.cap_res_X.t73 0.1603
R7847 two_stage_opamp_dummy_magic_0.cap_res_X.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t53 0.1603
R7848 two_stage_opamp_dummy_magic_0.cap_res_X.t74 two_stage_opamp_dummy_magic_0.cap_res_X.t36 0.1603
R7849 two_stage_opamp_dummy_magic_0.cap_res_X.t57 two_stage_opamp_dummy_magic_0.cap_res_X.t97 0.1603
R7850 two_stage_opamp_dummy_magic_0.cap_res_X.t116 two_stage_opamp_dummy_magic_0.cap_res_X.t78 0.1603
R7851 two_stage_opamp_dummy_magic_0.cap_res_X.t100 two_stage_opamp_dummy_magic_0.cap_res_X.t137 0.1603
R7852 two_stage_opamp_dummy_magic_0.cap_res_X.t15 two_stage_opamp_dummy_magic_0.cap_res_X.t120 0.1603
R7853 two_stage_opamp_dummy_magic_0.cap_res_X.t8 two_stage_opamp_dummy_magic_0.cap_res_X.t84 0.1603
R7854 two_stage_opamp_dummy_magic_0.cap_res_X.t99 two_stage_opamp_dummy_magic_0.cap_res_X.t41 0.1603
R7855 two_stage_opamp_dummy_magic_0.cap_res_X.t60 two_stage_opamp_dummy_magic_0.cap_res_X.t93 0.1603
R7856 two_stage_opamp_dummy_magic_0.cap_res_X.t26 two_stage_opamp_dummy_magic_0.cap_res_X.t3 0.1603
R7857 two_stage_opamp_dummy_magic_0.cap_res_X.t133 two_stage_opamp_dummy_magic_0.cap_res_X.t51 0.1603
R7858 two_stage_opamp_dummy_magic_0.cap_res_X.t82 two_stage_opamp_dummy_magic_0.cap_res_X.t14 0.1603
R7859 two_stage_opamp_dummy_magic_0.cap_res_X.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t61 0.1603
R7860 two_stage_opamp_dummy_magic_0.cap_res_X.t13 two_stage_opamp_dummy_magic_0.cap_res_X.t115 0.1603
R7861 two_stage_opamp_dummy_magic_0.cap_res_X.t103 two_stage_opamp_dummy_magic_0.cap_res_X.t71 0.1603
R7862 two_stage_opamp_dummy_magic_0.cap_res_X.t63 two_stage_opamp_dummy_magic_0.cap_res_X.t123 0.1603
R7863 two_stage_opamp_dummy_magic_0.cap_res_X.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t85 0.1603
R7864 two_stage_opamp_dummy_magic_0.cap_res_X.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t40 0.1603
R7865 two_stage_opamp_dummy_magic_0.cap_res_X.t21 two_stage_opamp_dummy_magic_0.cap_res_X.t113 0.1603
R7866 two_stage_opamp_dummy_magic_0.cap_res_X.t56 two_stage_opamp_dummy_magic_0.cap_res_X.t21 0.1603
R7867 two_stage_opamp_dummy_magic_0.cap_res_X.t18 two_stage_opamp_dummy_magic_0.cap_res_X.t56 0.1603
R7868 two_stage_opamp_dummy_magic_0.cap_res_X.t98 two_stage_opamp_dummy_magic_0.cap_res_X.t55 0.1603
R7869 two_stage_opamp_dummy_magic_0.cap_res_X.t59 two_stage_opamp_dummy_magic_0.cap_res_X.t98 0.1603
R7870 two_stage_opamp_dummy_magic_0.cap_res_X.t6 two_stage_opamp_dummy_magic_0.cap_res_X.t59 0.1603
R7871 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t125 0.159278
R7872 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t7 0.159278
R7873 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t107 0.159278
R7874 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t70 0.159278
R7875 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t32 0.159278
R7876 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t52 0.159278
R7877 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t67 0.159278
R7878 two_stage_opamp_dummy_magic_0.cap_res_X.t30 two_stage_opamp_dummy_magic_0.cap_res_X.n9 0.159278
R7879 two_stage_opamp_dummy_magic_0.cap_res_X.t64 two_stage_opamp_dummy_magic_0.cap_res_X.n10 0.159278
R7880 two_stage_opamp_dummy_magic_0.cap_res_X.t24 two_stage_opamp_dummy_magic_0.cap_res_X.n11 0.159278
R7881 two_stage_opamp_dummy_magic_0.cap_res_X.t126 two_stage_opamp_dummy_magic_0.cap_res_X.n12 0.159278
R7882 two_stage_opamp_dummy_magic_0.cap_res_X.t19 two_stage_opamp_dummy_magic_0.cap_res_X.n13 0.159278
R7883 two_stage_opamp_dummy_magic_0.cap_res_X.t122 two_stage_opamp_dummy_magic_0.cap_res_X.n14 0.159278
R7884 two_stage_opamp_dummy_magic_0.cap_res_X.t80 two_stage_opamp_dummy_magic_0.cap_res_X.n15 0.159278
R7885 two_stage_opamp_dummy_magic_0.cap_res_X.t37 two_stage_opamp_dummy_magic_0.cap_res_X.n16 0.159278
R7886 two_stage_opamp_dummy_magic_0.cap_res_X.t75 two_stage_opamp_dummy_magic_0.cap_res_X.n17 0.159278
R7887 two_stage_opamp_dummy_magic_0.cap_res_X.t35 two_stage_opamp_dummy_magic_0.cap_res_X.n18 0.159278
R7888 two_stage_opamp_dummy_magic_0.cap_res_X.t138 two_stage_opamp_dummy_magic_0.cap_res_X.n19 0.159278
R7889 two_stage_opamp_dummy_magic_0.cap_res_X.t29 two_stage_opamp_dummy_magic_0.cap_res_X.n20 0.159278
R7890 two_stage_opamp_dummy_magic_0.cap_res_X.t131 two_stage_opamp_dummy_magic_0.cap_res_X.n21 0.159278
R7891 two_stage_opamp_dummy_magic_0.cap_res_X.t110 two_stage_opamp_dummy_magic_0.cap_res_X.n22 0.159278
R7892 two_stage_opamp_dummy_magic_0.cap_res_X.t5 two_stage_opamp_dummy_magic_0.cap_res_X.n23 0.159278
R7893 two_stage_opamp_dummy_magic_0.cap_res_X.t106 two_stage_opamp_dummy_magic_0.cap_res_X.n24 0.159278
R7894 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t104 0.159278
R7895 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t1 0.159278
R7896 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t121 0.159278
R7897 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.t17 0.159278
R7898 two_stage_opamp_dummy_magic_0.cap_res_X.t67 two_stage_opamp_dummy_magic_0.cap_res_X.t88 0.137822
R7899 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t127 0.1368
R7900 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t42 0.1368
R7901 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t27 0.1368
R7902 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t9 0.1368
R7903 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t134 0.1368
R7904 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t25 0.1368
R7905 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t79 0.1368
R7906 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t65 0.1368
R7907 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t118 0.1368
R7908 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t31 0.1368
R7909 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t86 0.1368
R7910 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t69 0.1368
R7911 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t124 0.1368
R7912 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t109 0.1368
R7913 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t22 0.1368
R7914 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t76 0.1368
R7915 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t129 0.1368
R7916 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t117 0.1368
R7917 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t28 0.1368
R7918 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t16 0.1368
R7919 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t68 0.1368
R7920 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t54 0.1368
R7921 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t108 0.1368
R7922 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t20 0.1368
R7923 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t74 0.1368
R7924 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t57 0.1368
R7925 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t116 0.1368
R7926 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t100 0.1368
R7927 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t15 0.1368
R7928 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.t119 0.1368
R7929 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.t132 0.1368
R7930 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t8 0.114322
R7931 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.n29 0.1133
R7932 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.n30 0.1133
R7933 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.n31 0.1133
R7934 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.n32 0.1133
R7935 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.n33 0.1133
R7936 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.n0 0.1133
R7937 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.n1 0.1133
R7938 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.n2 0.1133
R7939 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.n3 0.1133
R7940 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.n4 0.1133
R7941 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.n5 0.1133
R7942 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.n6 0.1133
R7943 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.n7 0.1133
R7944 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.n8 0.1133
R7945 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.n25 0.1133
R7946 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.n26 0.1133
R7947 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.n27 0.1133
R7948 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n28 0.1133
R7949 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n34 0.1133
R7950 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t23 0.00152174
R7951 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t46 0.00152174
R7952 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t10 0.00152174
R7953 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t112 0.00152174
R7954 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t72 0.00152174
R7955 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t96 0.00152174
R7956 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t99 0.00152174
R7957 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.t60 0.00152174
R7958 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.t26 0.00152174
R7959 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.t133 0.00152174
R7960 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.t82 0.00152174
R7961 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.t44 0.00152174
R7962 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.t13 0.00152174
R7963 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.t103 0.00152174
R7964 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.t63 0.00152174
R7965 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.t33 0.00152174
R7966 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.t30 0.00152174
R7967 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t64 0.00152174
R7968 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t24 0.00152174
R7969 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t126 0.00152174
R7970 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t19 0.00152174
R7971 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t122 0.00152174
R7972 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t80 0.00152174
R7973 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t37 0.00152174
R7974 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t75 0.00152174
R7975 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t35 0.00152174
R7976 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t138 0.00152174
R7977 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t29 0.00152174
R7978 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t131 0.00152174
R7979 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t110 0.00152174
R7980 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t5 0.00152174
R7981 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t106 0.00152174
R7982 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t2 0.00152174
R7983 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t38 0.00152174
R7984 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t18 0.00152174
R7985 two_stage_opamp_dummy_magic_0.cap_res_X.t55 two_stage_opamp_dummy_magic_0.cap_res_X.n35 0.00152174
R7986 bgr_0.cap_res1.t0 bgr_0.cap_res1.t10 121.245
R7987 bgr_0.cap_res1.t16 bgr_0.cap_res1.t19 0.1603
R7988 bgr_0.cap_res1.t9 bgr_0.cap_res1.t15 0.1603
R7989 bgr_0.cap_res1.t14 bgr_0.cap_res1.t18 0.1603
R7990 bgr_0.cap_res1.t7 bgr_0.cap_res1.t13 0.1603
R7991 bgr_0.cap_res1.t1 bgr_0.cap_res1.t6 0.1603
R7992 bgr_0.cap_res1.n1 bgr_0.cap_res1.t17 0.159278
R7993 bgr_0.cap_res1.n2 bgr_0.cap_res1.t2 0.159278
R7994 bgr_0.cap_res1.n3 bgr_0.cap_res1.t8 0.159278
R7995 bgr_0.cap_res1.n4 bgr_0.cap_res1.t3 0.159278
R7996 bgr_0.cap_res1.n4 bgr_0.cap_res1.t16 0.1368
R7997 bgr_0.cap_res1.n4 bgr_0.cap_res1.t12 0.1368
R7998 bgr_0.cap_res1.n3 bgr_0.cap_res1.t9 0.1368
R7999 bgr_0.cap_res1.n3 bgr_0.cap_res1.t5 0.1368
R8000 bgr_0.cap_res1.n2 bgr_0.cap_res1.t14 0.1368
R8001 bgr_0.cap_res1.n2 bgr_0.cap_res1.t11 0.1368
R8002 bgr_0.cap_res1.n1 bgr_0.cap_res1.t7 0.1368
R8003 bgr_0.cap_res1.n1 bgr_0.cap_res1.t4 0.1368
R8004 bgr_0.cap_res1.n0 bgr_0.cap_res1.t1 0.1368
R8005 bgr_0.cap_res1.n0 bgr_0.cap_res1.t20 0.1368
R8006 bgr_0.cap_res1.t17 bgr_0.cap_res1.n0 0.00152174
R8007 bgr_0.cap_res1.t2 bgr_0.cap_res1.n1 0.00152174
R8008 bgr_0.cap_res1.t8 bgr_0.cap_res1.n2 0.00152174
R8009 bgr_0.cap_res1.t3 bgr_0.cap_res1.n3 0.00152174
R8010 bgr_0.cap_res1.t10 bgr_0.cap_res1.n4 0.00152174
R8011 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 297.151
R8012 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 297.151
R8013 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 297.151
R8014 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n26 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 123.067
R8015 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 118.861
R8016 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 118.861
R8017 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n18 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n17 118.861
R8018 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n21 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n20 118.861
R8019 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n24 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n23 118.861
R8020 bgr_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n26 42.063
R8021 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 39.4005
R8022 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 39.4005
R8023 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 39.4005
R8024 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 39.4005
R8025 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 39.4005
R8026 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 39.4005
R8027 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 19.7005
R8028 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 19.7005
R8029 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 19.7005
R8030 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 19.7005
R8031 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n17 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 19.7005
R8032 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n17 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 19.7005
R8033 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n20 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 19.7005
R8034 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n20 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 19.7005
R8035 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n23 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 19.7005
R8036 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n23 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 19.7005
R8037 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n26 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n25 6.2505
R8038 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 5.60467
R8039 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 5.588
R8040 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n24 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n22 5.54217
R8041 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 5.54217
R8042 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 5.32967
R8043 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 5.32967
R8044 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 5.063
R8045 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 5.04217
R8046 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n18 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n16 5.04217
R8047 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n21 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 5.04217
R8048 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n25 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n24 5.04217
R8049 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 5.0255
R8050 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 4.97967
R8051 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n19 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n18 4.97967
R8052 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n22 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n21 4.97967
R8053 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 4.76717
R8054 bgr_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 1.28175
R8055 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n22 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n19 0.563
R8056 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n19 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 0.563
R8057 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 0.563
R8058 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 0.563
R8059 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n25 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 0.563
R8060 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 0.5255
R8061 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.n5 1092.47
R8062 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.n0 755.798
R8063 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.n10 755.798
R8064 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.n2 530.201
R8065 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.n4 530.201
R8066 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.n6 530.201
R8067 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.n8 530.201
R8068 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t11 208.868
R8069 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.t4 208.868
R8070 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.t12 208.868
R8071 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.t6 208.868
R8072 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.t8 208.868
R8073 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.t5 208.868
R8074 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.t10 208.868
R8075 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.t7 208.868
R8076 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.t9 208.868
R8077 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.t13 208.868
R8078 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.n1 176.733
R8079 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.n3 176.733
R8080 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.n7 176.733
R8081 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n9 176.733
R8082 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.t2 117.591
R8083 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t1 117.591
R8084 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t3 108.424
R8085 two_stage_opamp_dummy_magic_0.V_tot.t0 two_stage_opamp_dummy_magic_0.V_tot.n11 108.424
R8086 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 120.504
R8087 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 100.322
R8088 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 99.7078
R8089 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n21 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n20 35.7193
R8090 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n21 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 31.5001
R8091 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 24.288
R8092 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 24.288
R8093 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 24.288
R8094 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n14 24.288
R8095 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n17 24.288
R8096 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 24.0005
R8097 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 24.0005
R8098 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 24.0005
R8099 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 24.0005
R8100 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 8.0005
R8101 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 8.0005
R8102 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 8.0005
R8103 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 8.0005
R8104 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 8.0005
R8105 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 8.0005
R8106 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 8.0005
R8107 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 8.0005
R8108 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 8.0005
R8109 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 8.0005
R8110 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n19 5.96925
R8111 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n16 5.7505
R8112 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 5.7505
R8113 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 5.7505
R8114 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 5.188
R8115 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 5.188
R8116 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 5.188
R8117 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 5.188
R8118 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 5.188
R8119 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n15 5.188
R8120 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n18 5.188
R8121 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n13 0.563
R8122 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 0.563
R8123 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 0.563
R8124 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 0.563
R8125 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 0.563
R8126 bgr_0.V_CMFB_S2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n21 0.047375
R8127 bgr_0.START_UP.n4 bgr_0.START_UP.t6 246.113
R8128 bgr_0.START_UP.n4 bgr_0.START_UP.t7 246.113
R8129 bgr_0.START_UP.n0 bgr_0.START_UP.t0 168.925
R8130 bgr_0.START_UP.n5 bgr_0.START_UP.n4 166.852
R8131 bgr_0.START_UP.n0 bgr_0.START_UP.t1 125.984
R8132 bgr_0.START_UP.n3 bgr_0.START_UP.n1 80.4102
R8133 bgr_0.START_UP.n3 bgr_0.START_UP.n2 77.0939
R8134 bgr_0.START_UP bgr_0.START_UP.n5 14.6567
R8135 bgr_0.START_UP.n1 bgr_0.START_UP.t2 13.1338
R8136 bgr_0.START_UP.n1 bgr_0.START_UP.t4 13.1338
R8137 bgr_0.START_UP.n2 bgr_0.START_UP.t3 13.1338
R8138 bgr_0.START_UP.n2 bgr_0.START_UP.t5 13.1338
R8139 bgr_0.START_UP bgr_0.START_UP.n0 8.688
R8140 bgr_0.START_UP.n5 bgr_0.START_UP.n3 6.13903
R8141 bgr_0.START_UP_NFET1 bgr_0.START_UP_NFET1.t1 161.3
R8142 bgr_0.START_UP_NFET1 bgr_0.START_UP_NFET1.t0 109.609
R8143 two_stage_opamp_dummy_magic_0.V_er_mir_p.n20 two_stage_opamp_dummy_magic_0.V_er_mir_p.n19 594.301
R8144 two_stage_opamp_dummy_magic_0.V_er_mir_p.n32 two_stage_opamp_dummy_magic_0.V_er_mir_p.n31 594.301
R8145 two_stage_opamp_dummy_magic_0.V_er_mir_p.n1 two_stage_opamp_dummy_magic_0.V_er_mir_p.n0 594.301
R8146 two_stage_opamp_dummy_magic_0.V_er_mir_p.n4 two_stage_opamp_dummy_magic_0.V_er_mir_p.n3 594.301
R8147 two_stage_opamp_dummy_magic_0.V_er_mir_p.n7 two_stage_opamp_dummy_magic_0.V_er_mir_p.n6 594.301
R8148 two_stage_opamp_dummy_magic_0.V_er_mir_p.n10 two_stage_opamp_dummy_magic_0.V_er_mir_p.n9 594.301
R8149 two_stage_opamp_dummy_magic_0.V_er_mir_p.n14 two_stage_opamp_dummy_magic_0.V_er_mir_p.n13 594.301
R8150 two_stage_opamp_dummy_magic_0.V_er_mir_p.n29 two_stage_opamp_dummy_magic_0.V_er_mir_p.n28 594.301
R8151 two_stage_opamp_dummy_magic_0.V_er_mir_p.n26 two_stage_opamp_dummy_magic_0.V_er_mir_p.n25 594.301
R8152 two_stage_opamp_dummy_magic_0.V_er_mir_p.n22 two_stage_opamp_dummy_magic_0.V_er_mir_p.n21 594.301
R8153 two_stage_opamp_dummy_magic_0.V_er_mir_p.n19 two_stage_opamp_dummy_magic_0.V_er_mir_p.t15 78.8005
R8154 two_stage_opamp_dummy_magic_0.V_er_mir_p.n19 two_stage_opamp_dummy_magic_0.V_er_mir_p.t12 78.8005
R8155 two_stage_opamp_dummy_magic_0.V_er_mir_p.n31 two_stage_opamp_dummy_magic_0.V_er_mir_p.t17 78.8005
R8156 two_stage_opamp_dummy_magic_0.V_er_mir_p.n31 two_stage_opamp_dummy_magic_0.V_er_mir_p.t11 78.8005
R8157 two_stage_opamp_dummy_magic_0.V_er_mir_p.n0 two_stage_opamp_dummy_magic_0.V_er_mir_p.t9 78.8005
R8158 two_stage_opamp_dummy_magic_0.V_er_mir_p.n0 two_stage_opamp_dummy_magic_0.V_er_mir_p.t1 78.8005
R8159 two_stage_opamp_dummy_magic_0.V_er_mir_p.n3 two_stage_opamp_dummy_magic_0.V_er_mir_p.t5 78.8005
R8160 two_stage_opamp_dummy_magic_0.V_er_mir_p.n3 two_stage_opamp_dummy_magic_0.V_er_mir_p.t3 78.8005
R8161 two_stage_opamp_dummy_magic_0.V_er_mir_p.n6 two_stage_opamp_dummy_magic_0.V_er_mir_p.t0 78.8005
R8162 two_stage_opamp_dummy_magic_0.V_er_mir_p.n6 two_stage_opamp_dummy_magic_0.V_er_mir_p.t7 78.8005
R8163 two_stage_opamp_dummy_magic_0.V_er_mir_p.n9 two_stage_opamp_dummy_magic_0.V_er_mir_p.t8 78.8005
R8164 two_stage_opamp_dummy_magic_0.V_er_mir_p.n9 two_stage_opamp_dummy_magic_0.V_er_mir_p.t2 78.8005
R8165 two_stage_opamp_dummy_magic_0.V_er_mir_p.n13 two_stage_opamp_dummy_magic_0.V_er_mir_p.t4 78.8005
R8166 two_stage_opamp_dummy_magic_0.V_er_mir_p.n13 two_stage_opamp_dummy_magic_0.V_er_mir_p.t6 78.8005
R8167 two_stage_opamp_dummy_magic_0.V_er_mir_p.n28 two_stage_opamp_dummy_magic_0.V_er_mir_p.t19 78.8005
R8168 two_stage_opamp_dummy_magic_0.V_er_mir_p.n28 two_stage_opamp_dummy_magic_0.V_er_mir_p.t14 78.8005
R8169 two_stage_opamp_dummy_magic_0.V_er_mir_p.n25 two_stage_opamp_dummy_magic_0.V_er_mir_p.t10 78.8005
R8170 two_stage_opamp_dummy_magic_0.V_er_mir_p.n25 two_stage_opamp_dummy_magic_0.V_er_mir_p.t16 78.8005
R8171 two_stage_opamp_dummy_magic_0.V_er_mir_p.n21 two_stage_opamp_dummy_magic_0.V_er_mir_p.t13 78.8005
R8172 two_stage_opamp_dummy_magic_0.V_er_mir_p.n21 two_stage_opamp_dummy_magic_0.V_er_mir_p.t18 78.8005
R8173 two_stage_opamp_dummy_magic_0.V_er_mir_p two_stage_opamp_dummy_magic_0.V_er_mir_p.n33 6.2505
R8174 two_stage_opamp_dummy_magic_0.V_er_mir_p.n23 two_stage_opamp_dummy_magic_0.V_er_mir_p.n20 6.10467
R8175 two_stage_opamp_dummy_magic_0.V_er_mir_p.n32 two_stage_opamp_dummy_magic_0.V_er_mir_p.n30 5.91717
R8176 two_stage_opamp_dummy_magic_0.V_er_mir_p.n20 two_stage_opamp_dummy_magic_0.V_er_mir_p.n18 5.91717
R8177 two_stage_opamp_dummy_magic_0.V_er_mir_p.n5 two_stage_opamp_dummy_magic_0.V_er_mir_p.n4 5.41717
R8178 two_stage_opamp_dummy_magic_0.V_er_mir_p.n8 two_stage_opamp_dummy_magic_0.V_er_mir_p.n4 5.22967
R8179 two_stage_opamp_dummy_magic_0.V_er_mir_p.n12 two_stage_opamp_dummy_magic_0.V_er_mir_p.n1 5.22967
R8180 two_stage_opamp_dummy_magic_0.V_er_mir_p.n16 two_stage_opamp_dummy_magic_0.V_er_mir_p.n15 5.063
R8181 two_stage_opamp_dummy_magic_0.V_er_mir_p.n7 two_stage_opamp_dummy_magic_0.V_er_mir_p.n5 4.85467
R8182 two_stage_opamp_dummy_magic_0.V_er_mir_p.n10 two_stage_opamp_dummy_magic_0.V_er_mir_p.n2 4.85467
R8183 two_stage_opamp_dummy_magic_0.V_er_mir_p.n15 two_stage_opamp_dummy_magic_0.V_er_mir_p.n14 4.85467
R8184 two_stage_opamp_dummy_magic_0.V_er_mir_p.n29 two_stage_opamp_dummy_magic_0.V_er_mir_p.n17 4.85467
R8185 two_stage_opamp_dummy_magic_0.V_er_mir_p.n26 two_stage_opamp_dummy_magic_0.V_er_mir_p.n24 4.85467
R8186 two_stage_opamp_dummy_magic_0.V_er_mir_p.n33 two_stage_opamp_dummy_magic_0.V_er_mir_p.n32 4.85467
R8187 two_stage_opamp_dummy_magic_0.V_er_mir_p.n23 two_stage_opamp_dummy_magic_0.V_er_mir_p.n22 4.85467
R8188 two_stage_opamp_dummy_magic_0.V_er_mir_p.n22 two_stage_opamp_dummy_magic_0.V_er_mir_p.n18 4.66717
R8189 two_stage_opamp_dummy_magic_0.V_er_mir_p.n8 two_stage_opamp_dummy_magic_0.V_er_mir_p.n7 4.66717
R8190 two_stage_opamp_dummy_magic_0.V_er_mir_p.n11 two_stage_opamp_dummy_magic_0.V_er_mir_p.n10 4.66717
R8191 two_stage_opamp_dummy_magic_0.V_er_mir_p.n14 two_stage_opamp_dummy_magic_0.V_er_mir_p.n12 4.66717
R8192 two_stage_opamp_dummy_magic_0.V_er_mir_p.n30 two_stage_opamp_dummy_magic_0.V_er_mir_p.n29 4.66717
R8193 two_stage_opamp_dummy_magic_0.V_er_mir_p.n27 two_stage_opamp_dummy_magic_0.V_er_mir_p.n26 4.66717
R8194 two_stage_opamp_dummy_magic_0.V_er_mir_p.n24 two_stage_opamp_dummy_magic_0.V_er_mir_p.n23 1.2505
R8195 two_stage_opamp_dummy_magic_0.V_er_mir_p.n24 two_stage_opamp_dummy_magic_0.V_er_mir_p.n17 1.2505
R8196 two_stage_opamp_dummy_magic_0.V_er_mir_p.n33 two_stage_opamp_dummy_magic_0.V_er_mir_p.n17 1.2505
R8197 two_stage_opamp_dummy_magic_0.V_er_mir_p.n30 two_stage_opamp_dummy_magic_0.V_er_mir_p.n27 1.2505
R8198 two_stage_opamp_dummy_magic_0.V_er_mir_p.n27 two_stage_opamp_dummy_magic_0.V_er_mir_p.n18 1.2505
R8199 two_stage_opamp_dummy_magic_0.V_er_mir_p two_stage_opamp_dummy_magic_0.V_er_mir_p.n16 0.938
R8200 two_stage_opamp_dummy_magic_0.V_er_mir_p.n15 two_stage_opamp_dummy_magic_0.V_er_mir_p.n2 0.563
R8201 two_stage_opamp_dummy_magic_0.V_er_mir_p.n5 two_stage_opamp_dummy_magic_0.V_er_mir_p.n2 0.563
R8202 two_stage_opamp_dummy_magic_0.V_er_mir_p.n11 two_stage_opamp_dummy_magic_0.V_er_mir_p.n8 0.563
R8203 two_stage_opamp_dummy_magic_0.V_er_mir_p.n12 two_stage_opamp_dummy_magic_0.V_er_mir_p.n11 0.563
R8204 two_stage_opamp_dummy_magic_0.V_er_mir_p.n16 two_stage_opamp_dummy_magic_0.V_er_mir_p.n1 0.354667
R8205 VIN-.n0 VIN-.t2 1001.34
R8206 VIN- VIN-.n9 593.684
R8207 VIN-.n9 VIN-.t7 273.134
R8208 VIN-.n0 VIN-.t4 273.134
R8209 VIN-.n1 VIN-.t9 273.134
R8210 VIN-.n2 VIN-.t3 273.134
R8211 VIN-.n3 VIN-.t8 273.134
R8212 VIN-.n4 VIN-.t6 273.134
R8213 VIN-.n5 VIN-.t0 273.134
R8214 VIN-.n6 VIN-.t5 273.134
R8215 VIN-.n7 VIN-.t10 273.134
R8216 VIN-.n8 VIN-.t1 273.134
R8217 VIN-.n9 VIN-.n8 176.733
R8218 VIN-.n8 VIN-.n7 176.733
R8219 VIN-.n7 VIN-.n6 176.733
R8220 VIN-.n6 VIN-.n5 176.733
R8221 VIN-.n5 VIN-.n4 176.733
R8222 VIN-.n4 VIN-.n3 176.733
R8223 VIN-.n3 VIN-.n2 176.733
R8224 VIN-.n2 VIN-.n1 176.733
R8225 VIN-.n1 VIN-.n0 176.733
R8226 two_stage_opamp_dummy_magic_0.Vb3.n27 two_stage_opamp_dummy_magic_0.Vb3.t25 768.551
R8227 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.t19 611.739
R8228 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.t13 611.739
R8229 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.t10 611.739
R8230 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.t27 611.739
R8231 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.n25 507.113
R8232 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.n17 506.582
R8233 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.t26 463.925
R8234 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.t20 463.925
R8235 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.t15 421.75
R8236 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.t17 421.75
R8237 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.t14 421.75
R8238 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.t16 421.75
R8239 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.t21 421.75
R8240 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.t18 421.75
R8241 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.t22 421.75
R8242 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.t12 421.75
R8243 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.t9 421.75
R8244 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.t28 421.75
R8245 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.t24 421.75
R8246 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.t8 421.75
R8247 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.t11 421.75
R8248 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.t23 421.75
R8249 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.n22 167.094
R8250 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.n23 167.094
R8251 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.n18 167.094
R8252 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.n19 167.094
R8253 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.n20 167.094
R8254 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.n13 167.094
R8255 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.n14 167.094
R8256 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.n15 167.094
R8257 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.n10 167.094
R8258 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.n11 167.094
R8259 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.n24 147.814
R8260 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.n21 147.814
R8261 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.n16 147.814
R8262 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.n12 147.814
R8263 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.n2 97.1505
R8264 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.n5 97.1505
R8265 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.n0 97.1505
R8266 two_stage_opamp_dummy_magic_0.Vb3.n28 two_stage_opamp_dummy_magic_0.Vb3.n9 73.3151
R8267 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb3.n28 47.563
R8268 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb3.n8 40.9693
R8269 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.t2 24.0005
R8270 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.t1 24.0005
R8271 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t4 24.0005
R8272 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t7 24.0005
R8273 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t5 24.0005
R8274 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t3 24.0005
R8275 two_stage_opamp_dummy_magic_0.Vb3.n27 two_stage_opamp_dummy_magic_0.Vb3.n26 14.4693
R8276 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.t6 11.2576
R8277 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.t0 11.2576
R8278 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.n4 5.58383
R8279 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.n3 5.58383
R8280 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.n6 5.52133
R8281 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.n3 5.52133
R8282 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.n1 5.02133
R8283 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.n7 4.5005
R8284 two_stage_opamp_dummy_magic_0.Vb3.n28 two_stage_opamp_dummy_magic_0.Vb3.n27 1.21925
R8285 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.n1 0.458833
R8286 two_stage_opamp_dummy_magic_0.VD3.n3 two_stage_opamp_dummy_magic_0.VD3.t35 671.418
R8287 two_stage_opamp_dummy_magic_0.VD3.n37 two_stage_opamp_dummy_magic_0.VD3.t32 671.418
R8288 two_stage_opamp_dummy_magic_0.VD3.t36 two_stage_opamp_dummy_magic_0.VD3.n34 213.131
R8289 two_stage_opamp_dummy_magic_0.VD3.n35 two_stage_opamp_dummy_magic_0.VD3.t33 213.131
R8290 two_stage_opamp_dummy_magic_0.VD3.t0 two_stage_opamp_dummy_magic_0.VD3.t36 146.155
R8291 two_stage_opamp_dummy_magic_0.VD3.t6 two_stage_opamp_dummy_magic_0.VD3.t0 146.155
R8292 two_stage_opamp_dummy_magic_0.VD3.t14 two_stage_opamp_dummy_magic_0.VD3.t6 146.155
R8293 two_stage_opamp_dummy_magic_0.VD3.t10 two_stage_opamp_dummy_magic_0.VD3.t14 146.155
R8294 two_stage_opamp_dummy_magic_0.VD3.t16 two_stage_opamp_dummy_magic_0.VD3.t10 146.155
R8295 two_stage_opamp_dummy_magic_0.VD3.t18 two_stage_opamp_dummy_magic_0.VD3.t16 146.155
R8296 two_stage_opamp_dummy_magic_0.VD3.t2 two_stage_opamp_dummy_magic_0.VD3.t18 146.155
R8297 two_stage_opamp_dummy_magic_0.VD3.t8 two_stage_opamp_dummy_magic_0.VD3.t2 146.155
R8298 two_stage_opamp_dummy_magic_0.VD3.t4 two_stage_opamp_dummy_magic_0.VD3.t8 146.155
R8299 two_stage_opamp_dummy_magic_0.VD3.t12 two_stage_opamp_dummy_magic_0.VD3.t4 146.155
R8300 two_stage_opamp_dummy_magic_0.VD3.t33 two_stage_opamp_dummy_magic_0.VD3.t12 146.155
R8301 two_stage_opamp_dummy_magic_0.VD3.n34 two_stage_opamp_dummy_magic_0.VD3.t37 76.2576
R8302 two_stage_opamp_dummy_magic_0.VD3.n35 two_stage_opamp_dummy_magic_0.VD3.t34 76.2576
R8303 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.n29 66.0338
R8304 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.n25 66.0338
R8305 two_stage_opamp_dummy_magic_0.VD3.n39 two_stage_opamp_dummy_magic_0.VD3.n38 66.0338
R8306 two_stage_opamp_dummy_magic_0.VD3.n43 two_stage_opamp_dummy_magic_0.VD3.n42 66.0338
R8307 two_stage_opamp_dummy_magic_0.VD3.n7 two_stage_opamp_dummy_magic_0.VD3.n6 66.0338
R8308 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.n9 66.0338
R8309 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.n12 66.0338
R8310 two_stage_opamp_dummy_magic_0.VD3.n17 two_stage_opamp_dummy_magic_0.VD3.n16 66.0338
R8311 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.n19 66.0338
R8312 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n22 66.0338
R8313 two_stage_opamp_dummy_magic_0.VD3.n47 two_stage_opamp_dummy_magic_0.VD3.n46 66.0338
R8314 two_stage_opamp_dummy_magic_0.VD3.n29 two_stage_opamp_dummy_magic_0.VD3.t1 11.2576
R8315 two_stage_opamp_dummy_magic_0.VD3.n29 two_stage_opamp_dummy_magic_0.VD3.t7 11.2576
R8316 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.t15 11.2576
R8317 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.t11 11.2576
R8318 two_stage_opamp_dummy_magic_0.VD3.n38 two_stage_opamp_dummy_magic_0.VD3.t5 11.2576
R8319 two_stage_opamp_dummy_magic_0.VD3.n38 two_stage_opamp_dummy_magic_0.VD3.t13 11.2576
R8320 two_stage_opamp_dummy_magic_0.VD3.n42 two_stage_opamp_dummy_magic_0.VD3.t3 11.2576
R8321 two_stage_opamp_dummy_magic_0.VD3.n42 two_stage_opamp_dummy_magic_0.VD3.t9 11.2576
R8322 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.t21 11.2576
R8323 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.t29 11.2576
R8324 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.t27 11.2576
R8325 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.t30 11.2576
R8326 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.t22 11.2576
R8327 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.t24 11.2576
R8328 two_stage_opamp_dummy_magic_0.VD3.n16 two_stage_opamp_dummy_magic_0.VD3.t26 11.2576
R8329 two_stage_opamp_dummy_magic_0.VD3.n16 two_stage_opamp_dummy_magic_0.VD3.t25 11.2576
R8330 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.t28 11.2576
R8331 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.t31 11.2576
R8332 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.t23 11.2576
R8333 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.t20 11.2576
R8334 two_stage_opamp_dummy_magic_0.VD3.n47 two_stage_opamp_dummy_magic_0.VD3.t17 11.2576
R8335 two_stage_opamp_dummy_magic_0.VD3.t19 two_stage_opamp_dummy_magic_0.VD3.n47 11.2576
R8336 two_stage_opamp_dummy_magic_0.VD3.n36 two_stage_opamp_dummy_magic_0.VD3.n2 5.91717
R8337 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n21 5.91717
R8338 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n7 5.91717
R8339 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.n7 5.91717
R8340 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.n28 5.563
R8341 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.n26 5.563
R8342 two_stage_opamp_dummy_magic_0.VD3.n46 two_stage_opamp_dummy_magic_0.VD3.n0 5.563
R8343 two_stage_opamp_dummy_magic_0.VD3.n40 two_stage_opamp_dummy_magic_0.VD3.n39 5.563
R8344 two_stage_opamp_dummy_magic_0.VD3.n43 two_stage_opamp_dummy_magic_0.VD3.n41 5.563
R8345 two_stage_opamp_dummy_magic_0.VD3.n40 two_stage_opamp_dummy_magic_0.VD3.n37 5.313
R8346 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.n3 5.313
R8347 two_stage_opamp_dummy_magic_0.VD3.n31 two_stage_opamp_dummy_magic_0.VD3.n30 5.29217
R8348 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.n1 5.29217
R8349 two_stage_opamp_dummy_magic_0.VD3.n39 two_stage_opamp_dummy_magic_0.VD3.n2 5.29217
R8350 two_stage_opamp_dummy_magic_0.VD3.n44 two_stage_opamp_dummy_magic_0.VD3.n43 5.29217
R8351 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.n32 5.29217
R8352 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.n10 5.29217
R8353 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.n8 5.29217
R8354 two_stage_opamp_dummy_magic_0.VD3.n14 two_stage_opamp_dummy_magic_0.VD3.n13 5.29217
R8355 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.n5 5.29217
R8356 two_stage_opamp_dummy_magic_0.VD3.n17 two_stage_opamp_dummy_magic_0.VD3.n15 5.29217
R8357 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.n17 5.29217
R8358 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.n4 5.29217
R8359 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.n20 5.29217
R8360 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.n23 5.29217
R8361 two_stage_opamp_dummy_magic_0.VD3.n46 two_stage_opamp_dummy_magic_0.VD3.n45 5.29217
R8362 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.n24 2.53175
R8363 two_stage_opamp_dummy_magic_0.VD3.n36 two_stage_opamp_dummy_magic_0.VD3.n35 1.03383
R8364 two_stage_opamp_dummy_magic_0.VD3.n34 two_stage_opamp_dummy_magic_0.VD3.n33 1.03383
R8365 two_stage_opamp_dummy_magic_0.VD3.n37 two_stage_opamp_dummy_magic_0.VD3.n36 0.8755
R8366 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.n3 0.8755
R8367 two_stage_opamp_dummy_magic_0.VD3.n45 two_stage_opamp_dummy_magic_0.VD3.n44 0.6255
R8368 two_stage_opamp_dummy_magic_0.VD3.n44 two_stage_opamp_dummy_magic_0.VD3.n2 0.6255
R8369 two_stage_opamp_dummy_magic_0.VD3.n41 two_stage_opamp_dummy_magic_0.VD3.n40 0.6255
R8370 two_stage_opamp_dummy_magic_0.VD3.n41 two_stage_opamp_dummy_magic_0.VD3.n0 0.6255
R8371 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.n0 0.6255
R8372 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.n27 0.6255
R8373 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.n18 0.6255
R8374 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.n5 0.6255
R8375 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n5 0.6255
R8376 two_stage_opamp_dummy_magic_0.VD3.n14 two_stage_opamp_dummy_magic_0.VD3.n11 0.6255
R8377 two_stage_opamp_dummy_magic_0.VD3.n15 two_stage_opamp_dummy_magic_0.VD3.n14 0.6255
R8378 two_stage_opamp_dummy_magic_0.VD3.n15 two_stage_opamp_dummy_magic_0.VD3.n4 0.6255
R8379 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.n4 0.6255
R8380 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.n31 0.6255
R8381 two_stage_opamp_dummy_magic_0.VD3.n31 two_stage_opamp_dummy_magic_0.VD3.n1 0.6255
R8382 two_stage_opamp_dummy_magic_0.VD3.n45 two_stage_opamp_dummy_magic_0.VD3.n1 0.6255
R8383 VIN+.n0 VIN+.t9 1001.34
R8384 VIN+ VIN+.n9 593.684
R8385 VIN+.n9 VIN+.t5 273.134
R8386 VIN+.n0 VIN+.t6 273.134
R8387 VIN+.n8 VIN+.t10 273.134
R8388 VIN+.n7 VIN+.t4 273.134
R8389 VIN+.n6 VIN+.t8 273.134
R8390 VIN+.n5 VIN+.t2 273.134
R8391 VIN+.n4 VIN+.t0 273.134
R8392 VIN+.n3 VIN+.t3 273.134
R8393 VIN+.n2 VIN+.t7 273.134
R8394 VIN+.n1 VIN+.t1 273.134
R8395 VIN+.n1 VIN+.n0 176.733
R8396 VIN+.n2 VIN+.n1 176.733
R8397 VIN+.n3 VIN+.n2 176.733
R8398 VIN+.n4 VIN+.n3 176.733
R8399 VIN+.n5 VIN+.n4 176.733
R8400 VIN+.n6 VIN+.n5 176.733
R8401 VIN+.n7 VIN+.n6 176.733
R8402 VIN+.n8 VIN+.n7 176.733
R8403 VIN+.n9 VIN+.n8 176.733
R8404 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.n1 514.134
R8405 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.n3 514.134
R8406 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n4 384.567
R8407 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n0 324.587
R8408 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t5 303.259
R8409 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t3 174.726
R8410 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.t7 174.726
R8411 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.t4 174.726
R8412 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t6 174.726
R8413 bgr_0.V_CUR_REF_REG.t1 bgr_0.V_CUR_REF_REG.n5 152.474
R8414 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.n2 128.534
R8415 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t2 39.4005
R8416 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t0 39.4005
R8417 two_stage_opamp_dummy_magic_0.Vb2_2.n2 two_stage_opamp_dummy_magic_0.Vb2_2.t4 661.375
R8418 two_stage_opamp_dummy_magic_0.Vb2_2.n4 two_stage_opamp_dummy_magic_0.Vb2_2.t7 661.375
R8419 two_stage_opamp_dummy_magic_0.Vb2_2.t5 two_stage_opamp_dummy_magic_0.Vb2_2.n0 213.131
R8420 two_stage_opamp_dummy_magic_0.Vb2_2.n3 two_stage_opamp_dummy_magic_0.Vb2_2.t8 213.131
R8421 two_stage_opamp_dummy_magic_0.Vb2_2.n6 two_stage_opamp_dummy_magic_0.Vb2_2.n1 154.983
R8422 two_stage_opamp_dummy_magic_0.Vb2_2.t0 two_stage_opamp_dummy_magic_0.Vb2_2.t5 146.155
R8423 two_stage_opamp_dummy_magic_0.Vb2_2.t8 two_stage_opamp_dummy_magic_0.Vb2_2.t0 146.155
R8424 two_stage_opamp_dummy_magic_0.Vb2_2.t6 two_stage_opamp_dummy_magic_0.Vb2_2.n0 76.2576
R8425 two_stage_opamp_dummy_magic_0.Vb2_2.n3 two_stage_opamp_dummy_magic_0.Vb2_2.t9 76.2576
R8426 two_stage_opamp_dummy_magic_0.Vb2_2.n7 two_stage_opamp_dummy_magic_0.Vb2_2.n6 66.4421
R8427 two_stage_opamp_dummy_magic_0.Vb2_2.n1 two_stage_opamp_dummy_magic_0.Vb2_2.t3 21.8894
R8428 two_stage_opamp_dummy_magic_0.Vb2_2.n1 two_stage_opamp_dummy_magic_0.Vb2_2.t2 21.8894
R8429 two_stage_opamp_dummy_magic_0.Vb2_2.t6 two_stage_opamp_dummy_magic_0.Vb2_2.n7 11.2576
R8430 two_stage_opamp_dummy_magic_0.Vb2_2.n7 two_stage_opamp_dummy_magic_0.Vb2_2.t1 11.2576
R8431 two_stage_opamp_dummy_magic_0.Vb2_2.n5 two_stage_opamp_dummy_magic_0.Vb2_2.n4 5.1255
R8432 two_stage_opamp_dummy_magic_0.Vb2_2.n6 two_stage_opamp_dummy_magic_0.Vb2_2.n5 4.92067
R8433 two_stage_opamp_dummy_magic_0.Vb2_2.n5 two_stage_opamp_dummy_magic_0.Vb2_2.n2 4.7505
R8434 two_stage_opamp_dummy_magic_0.Vb2_2.n4 two_stage_opamp_dummy_magic_0.Vb2_2.n3 1.888
R8435 two_stage_opamp_dummy_magic_0.Vb2_2.n2 two_stage_opamp_dummy_magic_0.Vb2_2.n0 1.888
R8436 bgr_0.Vin-.n7 bgr_0.Vin-.t12 688.859
R8437 bgr_0.Vin-.n11 bgr_0.Vin-.n10 577.21
R8438 bgr_0.Vin-.n9 bgr_0.Vin-.n8 514.134
R8439 bgr_0.Vin-.n6 bgr_0.Vin-.n5 314.046
R8440 bgr_0.Vin-.n7 bgr_0.Vin-.t8 174.726
R8441 bgr_0.Vin-.n8 bgr_0.Vin-.t10 174.726
R8442 bgr_0.Vin-.n9 bgr_0.Vin-.t9 174.726
R8443 bgr_0.Vin-.n10 bgr_0.Vin-.t11 174.726
R8444 bgr_0.Vin-.n8 bgr_0.Vin-.n7 128.534
R8445 bgr_0.Vin-.n10 bgr_0.Vin-.n9 128.534
R8446 bgr_0.Vin-.n12 bgr_0.Vin-.t6 118.785
R8447 bgr_0.Vin-.n16 bgr_0.Vin-.n15 83.5719
R8448 bgr_0.Vin-.n1 bgr_0.Vin-.n0 83.5719
R8449 bgr_0.Vin-.n4 bgr_0.Vin-.n2 79.3085
R8450 bgr_0.Vin-.n4 bgr_0.Vin-.n3 77.0655
R8451 bgr_0.Vin-.n19 bgr_0.Vin-.n1 73.8495
R8452 bgr_0.Vin-.t7 bgr_0.Vin-.n14 65.0341
R8453 bgr_0.Vin-.n5 bgr_0.Vin-.t0 39.4005
R8454 bgr_0.Vin-.n5 bgr_0.Vin-.t1 39.4005
R8455 bgr_0.Vin-.n13 bgr_0.Vin-.n12 28.5005
R8456 bgr_0.Vin-.n15 bgr_0.Vin-.n1 26.074
R8457 bgr_0.Vin-.n12 bgr_0.Vin-.n11 15.3443
R8458 bgr_0.Vin-.n2 bgr_0.Vin-.t2 13.1338
R8459 bgr_0.Vin-.n2 bgr_0.Vin-.t4 13.1338
R8460 bgr_0.Vin-.n3 bgr_0.Vin-.t3 13.1338
R8461 bgr_0.Vin-.n3 bgr_0.Vin-.t5 13.1338
R8462 bgr_0.Vin-.n11 bgr_0.Vin-.n6 12.6255
R8463 bgr_0.Vin-.n6 bgr_0.Vin-.n4 5.57549
R8464 bgr_0.Vin-.n16 bgr_0.Vin-.n14 1.56483
R8465 bgr_0.Vin-.n18 bgr_0.Vin-.n17 1.5505
R8466 bgr_0.Vin-.n17 bgr_0.Vin-.n0 0.885803
R8467 bgr_0.Vin-.n17 bgr_0.Vin-.n16 0.77514
R8468 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_0.Vin-.n0 0.756696
R8469 bgr_0.Vin-.n19 bgr_0.Vin-.n18 0.711459
R8470 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_0.Vin-.n19 0.576566
R8471 bgr_0.Vin-.n14 bgr_0.Vin-.n13 0.531499
R8472 bgr_0.Vin-.n15 bgr_0.Vin-.t7 0.290206
R8473 bgr_0.Vin-.n18 bgr_0.Vin-.n13 0.00817857
R8474 bgr_0.V_p_1.n5 bgr_0.V_p_1.n4 194.3
R8475 bgr_0.V_p_1.n7 bgr_0.V_p_1.n6 194.3
R8476 bgr_0.V_p_1.n9 bgr_0.V_p_1.n8 194.3
R8477 bgr_0.V_p_1.n11 bgr_0.V_p_1.n10 194.3
R8478 bgr_0.V_p_1.n13 bgr_0.V_p_1.n12 194.3
R8479 bgr_0.V_p_1.n0 bgr_0.V_p_1.t5 49.713
R8480 bgr_0.V_p_1.n4 bgr_0.V_p_1.t9 48.0005
R8481 bgr_0.V_p_1.n4 bgr_0.V_p_1.t1 48.0005
R8482 bgr_0.V_p_1.n6 bgr_0.V_p_1.t3 48.0005
R8483 bgr_0.V_p_1.n6 bgr_0.V_p_1.t6 48.0005
R8484 bgr_0.V_p_1.n8 bgr_0.V_p_1.t10 48.0005
R8485 bgr_0.V_p_1.n8 bgr_0.V_p_1.t2 48.0005
R8486 bgr_0.V_p_1.n10 bgr_0.V_p_1.t8 48.0005
R8487 bgr_0.V_p_1.n10 bgr_0.V_p_1.t0 48.0005
R8488 bgr_0.V_p_1.t4 bgr_0.V_p_1.n13 48.0005
R8489 bgr_0.V_p_1.n13 bgr_0.V_p_1.t7 48.0005
R8490 bgr_0.V_p_1.n3 bgr_0.V_p_1.n11 5.66717
R8491 bgr_0.V_p_1.n11 bgr_0.V_p_1.n1 5.66717
R8492 bgr_0.V_p_1.n5 bgr_0.V_p_1.n2 5.66717
R8493 bgr_0.V_p_1.n7 bgr_0.V_p_1.n2 5.04217
R8494 bgr_0.V_p_1.n0 bgr_0.V_p_1.n7 5.04217
R8495 bgr_0.V_p_1.n3 bgr_0.V_p_1.n9 5.04217
R8496 bgr_0.V_p_1.n9 bgr_0.V_p_1.n1 5.04217
R8497 bgr_0.V_p_1.n12 bgr_0.V_p_1.n1 5.04217
R8498 bgr_0.V_p_1.n0 bgr_0.V_p_1.n5 5.04217
R8499 bgr_0.V_p_1.n12 bgr_0.V_p_1.n3 5.04217
R8500 bgr_0.V_p_1.n1 bgr_0.V_p_1.n0 1.8755
R8501 bgr_0.V_p_1.n3 bgr_0.V_p_1.n2 1.2505
R8502 a_5310_4968.t0 a_5310_4968.t1 169.905
R8503 a_14560_4968.t0 a_14560_4968.t1 294.339
R8504 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 525.38
R8505 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 525.38
R8506 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 483.608
R8507 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 483.608
R8508 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 291.209
R8509 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 291.209
R8510 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 281.168
R8511 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 281.168
R8512 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 202.502
R8513 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 202.502
R8514 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 202.44
R8515 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 202.44
R8516 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 117.567
R8517 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 117.567
R8518 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 19.2193
R8519 a_12530_23988.t0 a_12530_23988.t1 178.133
R8520 a_14680_4968.t0 a_14680_4968.t1 169.905
R8521 a_7580_22380.t0 a_7580_22380.t1 178.133
R8522 two_stage_opamp_dummy_magic_0.Vb1_2.n1 two_stage_opamp_dummy_magic_0.Vb1_2.t0 65.3505
R8523 two_stage_opamp_dummy_magic_0.Vb1_2.n3 two_stage_opamp_dummy_magic_0.Vb1_2.n2 49.3505
R8524 two_stage_opamp_dummy_magic_0.Vb1_2.n6 two_stage_opamp_dummy_magic_0.Vb1_2.n5 49.3505
R8525 two_stage_opamp_dummy_magic_0.Vb1_2.n2 two_stage_opamp_dummy_magic_0.Vb1_2.t4 16.0005
R8526 two_stage_opamp_dummy_magic_0.Vb1_2.n2 two_stage_opamp_dummy_magic_0.Vb1_2.t2 16.0005
R8527 two_stage_opamp_dummy_magic_0.Vb1_2.t3 two_stage_opamp_dummy_magic_0.Vb1_2.n6 16.0005
R8528 two_stage_opamp_dummy_magic_0.Vb1_2.n6 two_stage_opamp_dummy_magic_0.Vb1_2.t1 16.0005
R8529 two_stage_opamp_dummy_magic_0.Vb1_2.n1 two_stage_opamp_dummy_magic_0.Vb1_2.n0 6.3755
R8530 two_stage_opamp_dummy_magic_0.Vb1_2.n4 two_stage_opamp_dummy_magic_0.Vb1_2.n1 6.1255
R8531 two_stage_opamp_dummy_magic_0.Vb1_2.n5 two_stage_opamp_dummy_magic_0.Vb1_2.n0 5.688
R8532 two_stage_opamp_dummy_magic_0.Vb1_2.n5 two_stage_opamp_dummy_magic_0.Vb1_2.n4 5.438
R8533 two_stage_opamp_dummy_magic_0.Vb1_2.n3 two_stage_opamp_dummy_magic_0.Vb1_2.n0 5.1255
R8534 two_stage_opamp_dummy_magic_0.Vb1_2.n4 two_stage_opamp_dummy_magic_0.Vb1_2.n3 4.8755
R8535 a_5190_4968.t0 a_5190_4968.t1 294.339
R8536 a_14240_1956.t0 a_14240_1956.t1 169.905
R8537 a_6810_23838.t0 a_6810_23838.t1 178.133
R8538 a_12410_22380.t0 a_12410_22380.t1 178.133
R8539 a_13060_22630.t0 a_13060_22630.t1 178.133
R8540 a_5760_1956.t0 a_5760_1956.t1 169.905
R8541 a_13180_23838.t0 a_13180_23838.t1 178.133
R8542 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 661.375
R8543 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 661.375
R8544 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 213.131
R8545 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 213.131
R8546 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 146.155
R8547 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 146.155
R8548 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 76.2576
R8549 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 76.2576
R8550 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 72.4424
R8551 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 66.4532
R8552 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 11.2576
R8553 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 11.2576
R8554 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 11.2576
R8555 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 11.2576
R8556 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 5.1255
R8557 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 4.9096
R8558 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 4.7505
R8559 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 1.888
R8560 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 1.888
C0 bgr_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_tail_gate 0.194271f
C1 bgr_0.START_UP_NFET1 bgr_0.START_UP 0.107665f
C2 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_er_mir_p 0.121861f
C3 bgr_0.NFET_GATE_10uA VDDA 0.896596f
C4 two_stage_opamp_dummy_magic_0.V_err_gate VDDA 3.79413f
C5 VOUT+ VOUT- 0.305434f
C6 two_stage_opamp_dummy_magic_0.V_err_amp_ref VOUT+ 0.039377f
C7 VIN+ two_stage_opamp_dummy_magic_0.VD2 0.44526f
C8 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.X 0.048253f
C9 bgr_0.START_UP VDDA 1.96085f
C10 m2_9370_16340# VDDA 0.010037f
C11 bgr_0.NFET_GATE_10uA bgr_0.PFET_GATE_10uA 0.517701f
C12 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_tail_gate 1.26251f
C13 VDDA two_stage_opamp_dummy_magic_0.V_er_mir_p 4.61308f
C14 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter VDDA 0.046803f
C15 two_stage_opamp_dummy_magic_0.X two_stage_opamp_dummy_magic_0.V_er_mir_p 0.015553f
C16 bgr_0.PFET_GATE_10uA m2_9370_16340# 0.010495f
C17 VDDA VOUT+ 15.2453f
C18 VOUT+ two_stage_opamp_dummy_magic_0.cap_res_Y 50.857998f
C19 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_gate 3.68994f
C20 two_stage_opamp_dummy_magic_0.V_tail_gate two_stage_opamp_dummy_magic_0.VD2 0.010726f
C21 VIN+ VIN- 0.155333f
C22 bgr_0.NFET_GATE_10uA bgr_0.START_UP 1.57006f
C23 VDDA VOUT- 15.2493f
C24 two_stage_opamp_dummy_magic_0.V_err_amp_ref VDDA 7.200779f
C25 VOUT- two_stage_opamp_dummy_magic_0.cap_res_Y 0.028842f
C26 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.cap_res_Y 0.244277f
C27 VOUT+ two_stage_opamp_dummy_magic_0.V_tail_gate 0.010419f
C28 VOUT- two_stage_opamp_dummy_magic_0.X 1.89641f
C29 VOUT- two_stage_opamp_dummy_magic_0.V_tail_gate 0.02548f
C30 bgr_0.NFET_GATE_10uA bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.016355f
C31 bgr_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.98661f
C32 bgr_0.START_UP_NFET1 VDDA 0.108124f
C33 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_er_mir_p 3.41966f
C34 VIN+ two_stage_opamp_dummy_magic_0.V_tail_gate 0.204972f
C35 m2_10730_16340# VDDA 0.010036f
C36 VIN- two_stage_opamp_dummy_magic_0.V_tail_gate 0.201317f
C37 VDDA two_stage_opamp_dummy_magic_0.cap_res_Y 0.685156f
C38 VDDA two_stage_opamp_dummy_magic_0.X 5.94769f
C39 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.053168f
C40 two_stage_opamp_dummy_magic_0.V_err_gate VOUT- 0.038284f
C41 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.466539f
C42 two_stage_opamp_dummy_magic_0.V_er_mir_p two_stage_opamp_dummy_magic_0.VD2 0.014803f
C43 bgr_0.START_UP two_stage_opamp_dummy_magic_0.V_err_amp_ref 2.52476f
C44 VDDA two_stage_opamp_dummy_magic_0.V_tail_gate 6.28625f
C45 bgr_0.PFET_GATE_10uA VDDA 10.1904f
C46 two_stage_opamp_dummy_magic_0.V_tail_gate two_stage_opamp_dummy_magic_0.cap_res_Y 0.034719f
C47 two_stage_opamp_dummy_magic_0.V_tail_gate two_stage_opamp_dummy_magic_0.X 0.128694f
C48 bgr_0.NFET_GATE_10uA bgr_0.START_UP_NFET1 0.253883f
C49 VIN- GNDA 2.10578f
C50 VIN+ GNDA 2.1107f
C51 VOUT- GNDA 20.803532f
C52 VOUT+ GNDA 20.84126f
C53 VDDA GNDA 0.133268p
C54 two_stage_opamp_dummy_magic_0.VD2 GNDA 2.810206f
C55 two_stage_opamp_dummy_magic_0.V_er_mir_p GNDA 1.054479f
C56 two_stage_opamp_dummy_magic_0.cap_res_Y GNDA 33.56648f
C57 two_stage_opamp_dummy_magic_0.X GNDA 7.658068f
C58 two_stage_opamp_dummy_magic_0.V_tail_gate GNDA 9.219989f
C59 bgr_0.START_UP GNDA 5.095123f
C60 bgr_0.START_UP_NFET1 GNDA 3.23382f
C61 two_stage_opamp_dummy_magic_0.V_err_gate GNDA 13.44459f
C62 bgr_0.NFET_GATE_10uA GNDA 7.81663f
C63 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA 17.7038f
C64 two_stage_opamp_dummy_magic_0.V_err_amp_ref GNDA 9.73803f
C65 bgr_0.PFET_GATE_10uA GNDA 5.972853f
C66 two_stage_opamp_dummy_magic_0.Vb1_2.t1 GNDA 0.047649f
C67 two_stage_opamp_dummy_magic_0.Vb1_2.n0 GNDA 0.318351f
C68 two_stage_opamp_dummy_magic_0.Vb1_2.t0 GNDA 0.161927f
C69 two_stage_opamp_dummy_magic_0.Vb1_2.n1 GNDA 0.491746f
C70 two_stage_opamp_dummy_magic_0.Vb1_2.t4 GNDA 0.047649f
C71 two_stage_opamp_dummy_magic_0.Vb1_2.t2 GNDA 0.047649f
C72 two_stage_opamp_dummy_magic_0.Vb1_2.n2 GNDA 0.103679f
C73 two_stage_opamp_dummy_magic_0.Vb1_2.n3 GNDA 0.407675f
C74 two_stage_opamp_dummy_magic_0.Vb1_2.n4 GNDA 0.297965f
C75 two_stage_opamp_dummy_magic_0.Vb1_2.n5 GNDA 0.42438f
C76 two_stage_opamp_dummy_magic_0.Vb1_2.n6 GNDA 0.103679f
C77 two_stage_opamp_dummy_magic_0.Vb1_2.t3 GNDA 0.047649f
C78 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 GNDA 0.104967f
C79 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 GNDA 0.306198f
C80 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 GNDA 0.26258f
C81 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 GNDA 0.311642f
C82 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 GNDA 0.163258f
C83 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 GNDA 0.265798f
C84 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 GNDA 0.176022f
C85 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 GNDA 0.509533f
C86 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 GNDA 0.26258f
C87 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 GNDA 0.311642f
C88 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 GNDA 0.163258f
C89 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 GNDA 0.306198f
C90 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 GNDA 0.265798f
C91 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 GNDA 0.176022f
C92 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 GNDA 0.509533f
C93 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 GNDA 0.104967f
C94 bgr_0.V_p_1.n0 GNDA 0.527156f
C95 bgr_0.V_p_1.n1 GNDA 0.157357f
C96 bgr_0.V_p_1.n2 GNDA 0.098819f
C97 bgr_0.V_p_1.n3 GNDA 0.157357f
C98 bgr_0.V_p_1.t5 GNDA 0.196701f
C99 bgr_0.V_p_1.n4 GNDA 0.017531f
C100 bgr_0.V_p_1.n5 GNDA 0.18041f
C101 bgr_0.V_p_1.n6 GNDA 0.017531f
C102 bgr_0.V_p_1.n7 GNDA 0.175416f
C103 bgr_0.V_p_1.n8 GNDA 0.017531f
C104 bgr_0.V_p_1.n9 GNDA 0.175416f
C105 bgr_0.V_p_1.n10 GNDA 0.017531f
C106 bgr_0.V_p_1.n11 GNDA 0.185403f
C107 bgr_0.V_p_1.n12 GNDA 0.175416f
C108 bgr_0.V_p_1.n13 GNDA 0.017531f
C109 bgr_0.Vin-.n0 GNDA 0.08443f
C110 bgr_0.Vin-.n1 GNDA 0.382704f
C111 bgr_0.Vin-.t2 GNDA 0.032806f
C112 bgr_0.Vin-.t4 GNDA 0.032806f
C113 bgr_0.Vin-.n2 GNDA 0.093858f
C114 bgr_0.Vin-.t3 GNDA 0.032806f
C115 bgr_0.Vin-.t5 GNDA 0.032806f
C116 bgr_0.Vin-.n3 GNDA 0.080724f
C117 bgr_0.Vin-.n4 GNDA 0.91389f
C118 bgr_0.Vin-.t0 GNDA 0.010935f
C119 bgr_0.Vin-.t1 GNDA 0.010935f
C120 bgr_0.Vin-.n5 GNDA 0.030922f
C121 bgr_0.Vin-.n6 GNDA 0.536105f
C122 bgr_0.Vin-.t12 GNDA 0.027051f
C123 bgr_0.Vin-.t8 GNDA 0.010115f
C124 bgr_0.Vin-.n7 GNDA 0.031727f
C125 bgr_0.Vin-.t10 GNDA 0.010115f
C126 bgr_0.Vin-.n8 GNDA 0.025972f
C127 bgr_0.Vin-.t9 GNDA 0.010115f
C128 bgr_0.Vin-.n9 GNDA 0.025972f
C129 bgr_0.Vin-.t11 GNDA 0.010115f
C130 bgr_0.Vin-.n10 GNDA 0.032247f
C131 bgr_0.Vin-.n11 GNDA 0.599168f
C132 bgr_0.Vin-.t6 GNDA 0.141676f
C133 bgr_0.Vin-.n12 GNDA 0.764746f
C134 bgr_0.Vin-.n13 GNDA 1.29395f
C135 bgr_0.Vin-.n14 GNDA 0.570547f
C136 bgr_0.Vin-.t7 GNDA 0.31671f
C137 bgr_0.Vin-.n15 GNDA 0.084586f
C138 bgr_0.Vin-.n16 GNDA 0.14477f
C139 bgr_0.Vin-.n17 GNDA 0.085378f
C140 bgr_0.Vin-.n18 GNDA 0.700926f
C141 bgr_0.Vin-.n19 GNDA 0.433629f
C142 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter GNDA 0.104756f
C143 bgr_0.V_CUR_REF_REG.n0 GNDA 0.045597f
C144 bgr_0.V_CUR_REF_REG.t5 GNDA 0.012811f
C145 bgr_0.V_CUR_REF_REG.n1 GNDA 0.027476f
C146 bgr_0.V_CUR_REF_REG.n2 GNDA 0.021381f
C147 bgr_0.V_CUR_REF_REG.n3 GNDA 0.021381f
C148 bgr_0.V_CUR_REF_REG.n4 GNDA 0.03263f
C149 bgr_0.V_CUR_REF_REG.n5 GNDA 1.7198f
C150 bgr_0.V_CUR_REF_REG.t1 GNDA 0.267612f
C151 two_stage_opamp_dummy_magic_0.VD3.t17 GNDA 0.067958f
C152 two_stage_opamp_dummy_magic_0.VD3.n0 GNDA 0.080546f
C153 two_stage_opamp_dummy_magic_0.VD3.n1 GNDA 0.073712f
C154 two_stage_opamp_dummy_magic_0.VD3.n2 GNDA 0.125745f
C155 two_stage_opamp_dummy_magic_0.VD3.t34 GNDA 0.241734f
C156 two_stage_opamp_dummy_magic_0.VD3.t37 GNDA 0.241734f
C157 two_stage_opamp_dummy_magic_0.VD3.t35 GNDA 0.118974f
C158 two_stage_opamp_dummy_magic_0.VD3.n3 GNDA 0.184796f
C159 two_stage_opamp_dummy_magic_0.VD3.n4 GNDA 0.073712f
C160 two_stage_opamp_dummy_magic_0.VD3.n5 GNDA 0.073712f
C161 two_stage_opamp_dummy_magic_0.VD3.t21 GNDA 0.067958f
C162 two_stage_opamp_dummy_magic_0.VD3.t29 GNDA 0.067958f
C163 two_stage_opamp_dummy_magic_0.VD3.n6 GNDA 0.139014f
C164 two_stage_opamp_dummy_magic_0.VD3.n7 GNDA 0.450087f
C165 two_stage_opamp_dummy_magic_0.VD3.n8 GNDA 0.125745f
C166 two_stage_opamp_dummy_magic_0.VD3.t27 GNDA 0.067958f
C167 two_stage_opamp_dummy_magic_0.VD3.t30 GNDA 0.067958f
C168 two_stage_opamp_dummy_magic_0.VD3.n9 GNDA 0.139014f
C169 two_stage_opamp_dummy_magic_0.VD3.n10 GNDA 0.437796f
C170 two_stage_opamp_dummy_magic_0.VD3.n11 GNDA 0.125745f
C171 two_stage_opamp_dummy_magic_0.VD3.t22 GNDA 0.067958f
C172 two_stage_opamp_dummy_magic_0.VD3.t24 GNDA 0.067958f
C173 two_stage_opamp_dummy_magic_0.VD3.n12 GNDA 0.139014f
C174 two_stage_opamp_dummy_magic_0.VD3.n13 GNDA 0.437796f
C175 two_stage_opamp_dummy_magic_0.VD3.n14 GNDA 0.073712f
C176 two_stage_opamp_dummy_magic_0.VD3.n15 GNDA 0.073712f
C177 two_stage_opamp_dummy_magic_0.VD3.t26 GNDA 0.067958f
C178 two_stage_opamp_dummy_magic_0.VD3.t25 GNDA 0.067958f
C179 two_stage_opamp_dummy_magic_0.VD3.n16 GNDA 0.139014f
C180 two_stage_opamp_dummy_magic_0.VD3.n17 GNDA 0.437796f
C181 two_stage_opamp_dummy_magic_0.VD3.n18 GNDA 0.073712f
C182 two_stage_opamp_dummy_magic_0.VD3.t28 GNDA 0.067958f
C183 two_stage_opamp_dummy_magic_0.VD3.t31 GNDA 0.067958f
C184 two_stage_opamp_dummy_magic_0.VD3.n19 GNDA 0.139014f
C185 two_stage_opamp_dummy_magic_0.VD3.n20 GNDA 0.437796f
C186 two_stage_opamp_dummy_magic_0.VD3.n21 GNDA 0.125745f
C187 two_stage_opamp_dummy_magic_0.VD3.t23 GNDA 0.067958f
C188 two_stage_opamp_dummy_magic_0.VD3.t20 GNDA 0.067958f
C189 two_stage_opamp_dummy_magic_0.VD3.n22 GNDA 0.139014f
C190 two_stage_opamp_dummy_magic_0.VD3.n23 GNDA 0.443941f
C191 two_stage_opamp_dummy_magic_0.VD3.n24 GNDA 0.132932f
C192 two_stage_opamp_dummy_magic_0.VD3.t15 GNDA 0.067958f
C193 two_stage_opamp_dummy_magic_0.VD3.t11 GNDA 0.067958f
C194 two_stage_opamp_dummy_magic_0.VD3.n25 GNDA 0.139014f
C195 two_stage_opamp_dummy_magic_0.VD3.n26 GNDA 0.468824f
C196 two_stage_opamp_dummy_magic_0.VD3.n27 GNDA 0.080546f
C197 two_stage_opamp_dummy_magic_0.VD3.n28 GNDA 0.122873f
C198 two_stage_opamp_dummy_magic_0.VD3.t1 GNDA 0.067958f
C199 two_stage_opamp_dummy_magic_0.VD3.t7 GNDA 0.067958f
C200 two_stage_opamp_dummy_magic_0.VD3.n29 GNDA 0.139014f
C201 two_stage_opamp_dummy_magic_0.VD3.n30 GNDA 0.468824f
C202 two_stage_opamp_dummy_magic_0.VD3.n31 GNDA 0.073712f
C203 two_stage_opamp_dummy_magic_0.VD3.n32 GNDA 0.132932f
C204 two_stage_opamp_dummy_magic_0.VD3.n33 GNDA 0.182585f
C205 two_stage_opamp_dummy_magic_0.VD3.n34 GNDA 0.701251f
C206 two_stage_opamp_dummy_magic_0.VD3.t36 GNDA 0.579264f
C207 two_stage_opamp_dummy_magic_0.VD3.t0 GNDA 0.454345f
C208 two_stage_opamp_dummy_magic_0.VD3.t6 GNDA 0.454345f
C209 two_stage_opamp_dummy_magic_0.VD3.t14 GNDA 0.454345f
C210 two_stage_opamp_dummy_magic_0.VD3.t10 GNDA 0.454345f
C211 two_stage_opamp_dummy_magic_0.VD3.t16 GNDA 0.454345f
C212 two_stage_opamp_dummy_magic_0.VD3.t18 GNDA 0.454345f
C213 two_stage_opamp_dummy_magic_0.VD3.t2 GNDA 0.454345f
C214 two_stage_opamp_dummy_magic_0.VD3.t8 GNDA 0.454345f
C215 two_stage_opamp_dummy_magic_0.VD3.t4 GNDA 0.454345f
C216 two_stage_opamp_dummy_magic_0.VD3.t12 GNDA 0.454345f
C217 two_stage_opamp_dummy_magic_0.VD3.t33 GNDA 0.579264f
C218 two_stage_opamp_dummy_magic_0.VD3.n35 GNDA 0.701251f
C219 two_stage_opamp_dummy_magic_0.VD3.n36 GNDA 0.188731f
C220 two_stage_opamp_dummy_magic_0.VD3.t32 GNDA 0.118974f
C221 two_stage_opamp_dummy_magic_0.VD3.n37 GNDA 0.184796f
C222 two_stage_opamp_dummy_magic_0.VD3.t5 GNDA 0.067958f
C223 two_stage_opamp_dummy_magic_0.VD3.t13 GNDA 0.067958f
C224 two_stage_opamp_dummy_magic_0.VD3.n38 GNDA 0.139014f
C225 two_stage_opamp_dummy_magic_0.VD3.n39 GNDA 0.468824f
C226 two_stage_opamp_dummy_magic_0.VD3.n40 GNDA 0.122873f
C227 two_stage_opamp_dummy_magic_0.VD3.n41 GNDA 0.080546f
C228 two_stage_opamp_dummy_magic_0.VD3.t3 GNDA 0.067958f
C229 two_stage_opamp_dummy_magic_0.VD3.t9 GNDA 0.067958f
C230 two_stage_opamp_dummy_magic_0.VD3.n42 GNDA 0.139014f
C231 two_stage_opamp_dummy_magic_0.VD3.n43 GNDA 0.468824f
C232 two_stage_opamp_dummy_magic_0.VD3.n44 GNDA 0.073712f
C233 two_stage_opamp_dummy_magic_0.VD3.n45 GNDA 0.073712f
C234 two_stage_opamp_dummy_magic_0.VD3.n46 GNDA 0.468824f
C235 two_stage_opamp_dummy_magic_0.VD3.n47 GNDA 0.139014f
C236 two_stage_opamp_dummy_magic_0.VD3.t19 GNDA 0.067958f
C237 two_stage_opamp_dummy_magic_0.Vb3.t5 GNDA 0.015858f
C238 two_stage_opamp_dummy_magic_0.Vb3.t3 GNDA 0.015858f
C239 two_stage_opamp_dummy_magic_0.Vb3.n0 GNDA 0.033764f
C240 two_stage_opamp_dummy_magic_0.Vb3.n1 GNDA 0.140069f
C241 two_stage_opamp_dummy_magic_0.Vb3.t2 GNDA 0.015858f
C242 two_stage_opamp_dummy_magic_0.Vb3.t1 GNDA 0.015858f
C243 two_stage_opamp_dummy_magic_0.Vb3.n2 GNDA 0.033764f
C244 two_stage_opamp_dummy_magic_0.Vb3.n3 GNDA 0.188325f
C245 two_stage_opamp_dummy_magic_0.Vb3.n4 GNDA 0.126997f
C246 two_stage_opamp_dummy_magic_0.Vb3.t4 GNDA 0.015858f
C247 two_stage_opamp_dummy_magic_0.Vb3.t7 GNDA 0.015858f
C248 two_stage_opamp_dummy_magic_0.Vb3.n5 GNDA 0.033764f
C249 two_stage_opamp_dummy_magic_0.Vb3.n6 GNDA 0.188325f
C250 two_stage_opamp_dummy_magic_0.Vb3.n7 GNDA 0.120394f
C251 two_stage_opamp_dummy_magic_0.Vb3.n8 GNDA 0.805152f
C252 two_stage_opamp_dummy_magic_0.Vb3.t6 GNDA 0.055501f
C253 two_stage_opamp_dummy_magic_0.Vb3.t0 GNDA 0.055501f
C254 two_stage_opamp_dummy_magic_0.Vb3.n9 GNDA 0.153113f
C255 two_stage_opamp_dummy_magic_0.Vb3.t23 GNDA 0.078494f
C256 two_stage_opamp_dummy_magic_0.Vb3.t11 GNDA 0.078494f
C257 two_stage_opamp_dummy_magic_0.Vb3.t8 GNDA 0.078494f
C258 two_stage_opamp_dummy_magic_0.Vb3.t27 GNDA 0.090582f
C259 two_stage_opamp_dummy_magic_0.Vb3.n10 GNDA 0.073543f
C260 two_stage_opamp_dummy_magic_0.Vb3.n11 GNDA 0.045194f
C261 two_stage_opamp_dummy_magic_0.Vb3.n12 GNDA 0.044315f
C262 two_stage_opamp_dummy_magic_0.Vb3.t24 GNDA 0.078494f
C263 two_stage_opamp_dummy_magic_0.Vb3.t28 GNDA 0.078494f
C264 two_stage_opamp_dummy_magic_0.Vb3.t9 GNDA 0.078494f
C265 two_stage_opamp_dummy_magic_0.Vb3.t12 GNDA 0.078494f
C266 two_stage_opamp_dummy_magic_0.Vb3.t10 GNDA 0.090582f
C267 two_stage_opamp_dummy_magic_0.Vb3.n13 GNDA 0.073543f
C268 two_stage_opamp_dummy_magic_0.Vb3.n14 GNDA 0.045194f
C269 two_stage_opamp_dummy_magic_0.Vb3.n15 GNDA 0.045194f
C270 two_stage_opamp_dummy_magic_0.Vb3.n16 GNDA 0.044315f
C271 two_stage_opamp_dummy_magic_0.Vb3.t20 GNDA 0.081269f
C272 two_stage_opamp_dummy_magic_0.Vb3.n17 GNDA 0.08575f
C273 two_stage_opamp_dummy_magic_0.Vb3.t22 GNDA 0.078494f
C274 two_stage_opamp_dummy_magic_0.Vb3.t18 GNDA 0.078494f
C275 two_stage_opamp_dummy_magic_0.Vb3.t21 GNDA 0.078494f
C276 two_stage_opamp_dummy_magic_0.Vb3.t16 GNDA 0.078494f
C277 two_stage_opamp_dummy_magic_0.Vb3.t13 GNDA 0.090582f
C278 two_stage_opamp_dummy_magic_0.Vb3.n18 GNDA 0.073543f
C279 two_stage_opamp_dummy_magic_0.Vb3.n19 GNDA 0.045194f
C280 two_stage_opamp_dummy_magic_0.Vb3.n20 GNDA 0.045194f
C281 two_stage_opamp_dummy_magic_0.Vb3.n21 GNDA 0.044315f
C282 two_stage_opamp_dummy_magic_0.Vb3.t14 GNDA 0.078494f
C283 two_stage_opamp_dummy_magic_0.Vb3.t17 GNDA 0.078494f
C284 two_stage_opamp_dummy_magic_0.Vb3.t15 GNDA 0.078494f
C285 two_stage_opamp_dummy_magic_0.Vb3.t19 GNDA 0.090582f
C286 two_stage_opamp_dummy_magic_0.Vb3.n22 GNDA 0.073543f
C287 two_stage_opamp_dummy_magic_0.Vb3.n23 GNDA 0.045194f
C288 two_stage_opamp_dummy_magic_0.Vb3.n24 GNDA 0.044315f
C289 two_stage_opamp_dummy_magic_0.Vb3.t26 GNDA 0.081269f
C290 two_stage_opamp_dummy_magic_0.Vb3.n25 GNDA 0.086364f
C291 two_stage_opamp_dummy_magic_0.Vb3.n26 GNDA 1.33624f
C292 two_stage_opamp_dummy_magic_0.Vb3.t25 GNDA 0.102539f
C293 two_stage_opamp_dummy_magic_0.Vb3.n27 GNDA 0.363304f
C294 two_stage_opamp_dummy_magic_0.Vb3.n28 GNDA 1.1613f
C295 bgr_0.VB3_CUR_BIAS GNDA 1.7683f
C296 two_stage_opamp_dummy_magic_0.V_er_mir_p.t9 GNDA 0.030734f
C297 two_stage_opamp_dummy_magic_0.V_er_mir_p.t1 GNDA 0.030734f
C298 two_stage_opamp_dummy_magic_0.V_er_mir_p.n0 GNDA 0.062623f
C299 two_stage_opamp_dummy_magic_0.V_er_mir_p.n1 GNDA 0.309237f
C300 two_stage_opamp_dummy_magic_0.V_er_mir_p.n2 GNDA 0.195142f
C301 two_stage_opamp_dummy_magic_0.V_er_mir_p.t5 GNDA 0.030734f
C302 two_stage_opamp_dummy_magic_0.V_er_mir_p.t3 GNDA 0.030734f
C303 two_stage_opamp_dummy_magic_0.V_er_mir_p.n3 GNDA 0.062623f
C304 two_stage_opamp_dummy_magic_0.V_er_mir_p.n4 GNDA 0.461459f
C305 two_stage_opamp_dummy_magic_0.V_er_mir_p.n5 GNDA 0.33146f
C306 two_stage_opamp_dummy_magic_0.V_er_mir_p.t0 GNDA 0.030734f
C307 two_stage_opamp_dummy_magic_0.V_er_mir_p.t7 GNDA 0.030734f
C308 two_stage_opamp_dummy_magic_0.V_er_mir_p.n6 GNDA 0.062623f
C309 two_stage_opamp_dummy_magic_0.V_er_mir_p.n7 GNDA 0.430057f
C310 two_stage_opamp_dummy_magic_0.V_er_mir_p.n8 GNDA 0.317572f
C311 two_stage_opamp_dummy_magic_0.V_er_mir_p.t8 GNDA 0.030734f
C312 two_stage_opamp_dummy_magic_0.V_er_mir_p.t2 GNDA 0.030734f
C313 two_stage_opamp_dummy_magic_0.V_er_mir_p.n9 GNDA 0.062623f
C314 two_stage_opamp_dummy_magic_0.V_er_mir_p.n10 GNDA 0.430057f
C315 two_stage_opamp_dummy_magic_0.V_er_mir_p.n11 GNDA 0.188103f
C316 two_stage_opamp_dummy_magic_0.V_er_mir_p.n12 GNDA 0.317572f
C317 two_stage_opamp_dummy_magic_0.V_er_mir_p.t4 GNDA 0.030734f
C318 two_stage_opamp_dummy_magic_0.V_er_mir_p.t6 GNDA 0.030734f
C319 two_stage_opamp_dummy_magic_0.V_er_mir_p.n13 GNDA 0.062623f
C320 two_stage_opamp_dummy_magic_0.V_er_mir_p.n14 GNDA 0.430057f
C321 two_stage_opamp_dummy_magic_0.V_er_mir_p.n15 GNDA 0.320811f
C322 two_stage_opamp_dummy_magic_0.V_er_mir_p.n16 GNDA 0.241551f
C323 two_stage_opamp_dummy_magic_0.V_er_mir_p.n17 GNDA 0.330373f
C324 two_stage_opamp_dummy_magic_0.V_er_mir_p.n18 GNDA 0.491089f
C325 two_stage_opamp_dummy_magic_0.V_er_mir_p.t15 GNDA 0.030734f
C326 two_stage_opamp_dummy_magic_0.V_er_mir_p.t12 GNDA 0.030734f
C327 two_stage_opamp_dummy_magic_0.V_er_mir_p.n19 GNDA 0.062623f
C328 two_stage_opamp_dummy_magic_0.V_er_mir_p.n20 GNDA 0.519987f
C329 two_stage_opamp_dummy_magic_0.V_er_mir_p.t13 GNDA 0.030734f
C330 two_stage_opamp_dummy_magic_0.V_er_mir_p.t18 GNDA 0.030734f
C331 two_stage_opamp_dummy_magic_0.V_er_mir_p.n21 GNDA 0.062623f
C332 two_stage_opamp_dummy_magic_0.V_er_mir_p.n22 GNDA 0.430057f
C333 two_stage_opamp_dummy_magic_0.V_er_mir_p.n23 GNDA 0.505107f
C334 two_stage_opamp_dummy_magic_0.V_er_mir_p.n24 GNDA 0.330373f
C335 two_stage_opamp_dummy_magic_0.V_er_mir_p.t10 GNDA 0.030734f
C336 two_stage_opamp_dummy_magic_0.V_er_mir_p.t16 GNDA 0.030734f
C337 two_stage_opamp_dummy_magic_0.V_er_mir_p.n25 GNDA 0.062623f
C338 two_stage_opamp_dummy_magic_0.V_er_mir_p.n26 GNDA 0.430057f
C339 two_stage_opamp_dummy_magic_0.V_er_mir_p.n27 GNDA 0.323333f
C340 two_stage_opamp_dummy_magic_0.V_er_mir_p.t19 GNDA 0.030734f
C341 two_stage_opamp_dummy_magic_0.V_er_mir_p.t14 GNDA 0.030734f
C342 two_stage_opamp_dummy_magic_0.V_er_mir_p.n28 GNDA 0.062623f
C343 two_stage_opamp_dummy_magic_0.V_er_mir_p.n29 GNDA 0.430057f
C344 two_stage_opamp_dummy_magic_0.V_er_mir_p.n30 GNDA 0.491089f
C345 two_stage_opamp_dummy_magic_0.V_er_mir_p.t17 GNDA 0.030734f
C346 two_stage_opamp_dummy_magic_0.V_er_mir_p.t11 GNDA 0.030734f
C347 two_stage_opamp_dummy_magic_0.V_er_mir_p.n31 GNDA 0.062623f
C348 two_stage_opamp_dummy_magic_0.V_er_mir_p.n32 GNDA 0.474991f
C349 two_stage_opamp_dummy_magic_0.V_er_mir_p.n33 GNDA 0.565428f
C350 bgr_0.START_UP.t0 GNDA 2.02004f
C351 bgr_0.START_UP.t1 GNDA 0.075562f
C352 bgr_0.START_UP.n0 GNDA 0.650598f
C353 bgr_0.START_UP.t2 GNDA 0.059442f
C354 bgr_0.START_UP.t4 GNDA 0.059442f
C355 bgr_0.START_UP.n1 GNDA 0.189396f
C356 bgr_0.START_UP.t3 GNDA 0.059442f
C357 bgr_0.START_UP.t5 GNDA 0.059442f
C358 bgr_0.START_UP.n2 GNDA 0.148916f
C359 bgr_0.START_UP.n3 GNDA 1.8941f
C360 bgr_0.START_UP.t7 GNDA 0.022671f
C361 bgr_0.START_UP.t6 GNDA 0.022671f
C362 bgr_0.START_UP.n4 GNDA 0.061199f
C363 bgr_0.START_UP.n5 GNDA 0.748295f
C364 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 GNDA 0.027874f
C365 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 GNDA 0.027874f
C366 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 GNDA 0.074525f
C367 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 GNDA 0.027874f
C368 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 GNDA 0.027874f
C369 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 GNDA 0.071124f
C370 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 GNDA 2.16068f
C371 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 GNDA 0.346139f
C372 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 GNDA 0.096954f
C373 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 GNDA 0.16682f
C374 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA 0.083621f
C375 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 GNDA 0.083621f
C376 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 GNDA 0.17885f
C377 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 GNDA 0.559442f
C378 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 GNDA 0.083621f
C379 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 GNDA 0.083621f
C380 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 GNDA 0.17885f
C381 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 GNDA 0.54429f
C382 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 GNDA 0.16682f
C383 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 GNDA 0.096954f
C384 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA 0.083621f
C385 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 GNDA 0.083621f
C386 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 GNDA 0.17885f
C387 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 GNDA 0.54429f
C388 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n13 GNDA 0.096954f
C389 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 GNDA 0.083621f
C390 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 GNDA 0.083621f
C391 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n14 GNDA 0.17885f
C392 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n15 GNDA 0.54429f
C393 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n16 GNDA 0.16682f
C394 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 GNDA 0.083621f
C395 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 GNDA 0.083621f
C396 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n17 GNDA 0.17885f
C397 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n18 GNDA 0.551866f
C398 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n19 GNDA 0.216176f
C399 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n20 GNDA 2.12983f
C400 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n21 GNDA 2.31013f
C401 bgr_0.V_CMFB_S2 GNDA 0.013937f
C402 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 GNDA 0.021174f
C403 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 GNDA 0.021174f
C404 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 GNDA 0.043243f
C405 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 GNDA 0.16469f
C406 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 GNDA 0.021174f
C407 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 GNDA 0.021174f
C408 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 GNDA 0.043243f
C409 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 GNDA 0.227515f
C410 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 GNDA 0.157479f
C411 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 GNDA 0.021174f
C412 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 GNDA 0.021174f
C413 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 GNDA 0.043243f
C414 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 GNDA 0.216541f
C415 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 GNDA 0.163297f
C416 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 GNDA 0.108203f
C417 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 GNDA 0.273637f
C418 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 GNDA 0.06689f
C419 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 GNDA 0.118314f
C420 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 GNDA 0.042349f
C421 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 GNDA 0.042349f
C422 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 GNDA 0.086586f
C423 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 GNDA 0.290839f
C424 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 GNDA 0.042349f
C425 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 GNDA 0.042349f
C426 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 GNDA 0.086586f
C427 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 GNDA 0.28008f
C428 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 GNDA 0.113731f
C429 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n16 GNDA 0.06689f
C430 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 GNDA 0.042349f
C431 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 GNDA 0.042349f
C432 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n17 GNDA 0.086586f
C433 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n18 GNDA 0.28008f
C434 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n19 GNDA 0.069335f
C435 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 GNDA 0.042349f
C436 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 GNDA 0.042349f
C437 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n20 GNDA 0.086586f
C438 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n21 GNDA 0.28008f
C439 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n22 GNDA 0.118314f
C440 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 GNDA 0.042349f
C441 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 GNDA 0.042349f
C442 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n23 GNDA 0.086586f
C443 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n24 GNDA 0.285613f
C444 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n25 GNDA 0.171152f
C445 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n26 GNDA 1.94694f
C446 bgr_0.V_CMFB_S1 GNDA 1.08719f
C447 bgr_0.cap_res1.t12 GNDA 0.331712f
C448 bgr_0.cap_res1.t19 GNDA 0.349187f
C449 bgr_0.cap_res1.t16 GNDA 0.350452f
C450 bgr_0.cap_res1.t5 GNDA 0.331712f
C451 bgr_0.cap_res1.t15 GNDA 0.349187f
C452 bgr_0.cap_res1.t9 GNDA 0.350452f
C453 bgr_0.cap_res1.t11 GNDA 0.331712f
C454 bgr_0.cap_res1.t18 GNDA 0.349187f
C455 bgr_0.cap_res1.t14 GNDA 0.350452f
C456 bgr_0.cap_res1.t4 GNDA 0.331712f
C457 bgr_0.cap_res1.t13 GNDA 0.349187f
C458 bgr_0.cap_res1.t7 GNDA 0.350452f
C459 bgr_0.cap_res1.t20 GNDA 0.331712f
C460 bgr_0.cap_res1.t6 GNDA 0.349187f
C461 bgr_0.cap_res1.t1 GNDA 0.350452f
C462 bgr_0.cap_res1.n0 GNDA 0.23406f
C463 bgr_0.cap_res1.t17 GNDA 0.186395f
C464 bgr_0.cap_res1.n1 GNDA 0.253961f
C465 bgr_0.cap_res1.t2 GNDA 0.186395f
C466 bgr_0.cap_res1.n2 GNDA 0.253961f
C467 bgr_0.cap_res1.t8 GNDA 0.186395f
C468 bgr_0.cap_res1.n3 GNDA 0.253961f
C469 bgr_0.cap_res1.t3 GNDA 0.186395f
C470 bgr_0.cap_res1.n4 GNDA 0.253961f
C471 bgr_0.cap_res1.t10 GNDA 0.363549f
C472 bgr_0.cap_res1.t0 GNDA 0.08421f
C473 two_stage_opamp_dummy_magic_0.cap_res_X.t90 GNDA 0.34556f
C474 two_stage_opamp_dummy_magic_0.cap_res_X.t127 GNDA 0.346812f
C475 two_stage_opamp_dummy_magic_0.cap_res_X.t49 GNDA 0.34556f
C476 two_stage_opamp_dummy_magic_0.cap_res_X.t88 GNDA 0.348269f
C477 two_stage_opamp_dummy_magic_0.cap_res_X.t67 GNDA 0.378793f
C478 two_stage_opamp_dummy_magic_0.cap_res_X.t130 GNDA 0.34556f
C479 two_stage_opamp_dummy_magic_0.cap_res_X.t27 GNDA 0.346812f
C480 two_stage_opamp_dummy_magic_0.cap_res_X.t81 GNDA 0.34556f
C481 two_stage_opamp_dummy_magic_0.cap_res_X.t42 GNDA 0.346812f
C482 two_stage_opamp_dummy_magic_0.cap_res_X.t95 GNDA 0.34556f
C483 two_stage_opamp_dummy_magic_0.cap_res_X.t134 GNDA 0.346812f
C484 two_stage_opamp_dummy_magic_0.cap_res_X.t45 GNDA 0.34556f
C485 two_stage_opamp_dummy_magic_0.cap_res_X.t9 GNDA 0.346812f
C486 two_stage_opamp_dummy_magic_0.cap_res_X.t43 GNDA 0.34556f
C487 two_stage_opamp_dummy_magic_0.cap_res_X.t79 GNDA 0.346812f
C488 two_stage_opamp_dummy_magic_0.cap_res_X.t58 GNDA 0.34556f
C489 two_stage_opamp_dummy_magic_0.cap_res_X.t25 GNDA 0.346812f
C490 two_stage_opamp_dummy_magic_0.cap_res_X.t83 GNDA 0.34556f
C491 two_stage_opamp_dummy_magic_0.cap_res_X.t118 GNDA 0.346812f
C492 two_stage_opamp_dummy_magic_0.cap_res_X.t102 GNDA 0.34556f
C493 two_stage_opamp_dummy_magic_0.cap_res_X.t65 GNDA 0.346812f
C494 two_stage_opamp_dummy_magic_0.cap_res_X.t48 GNDA 0.34556f
C495 two_stage_opamp_dummy_magic_0.cap_res_X.t86 GNDA 0.346812f
C496 two_stage_opamp_dummy_magic_0.cap_res_X.t66 GNDA 0.34556f
C497 two_stage_opamp_dummy_magic_0.cap_res_X.t31 GNDA 0.346812f
C498 two_stage_opamp_dummy_magic_0.cap_res_X.t89 GNDA 0.34556f
C499 two_stage_opamp_dummy_magic_0.cap_res_X.t124 GNDA 0.346812f
C500 two_stage_opamp_dummy_magic_0.cap_res_X.t105 GNDA 0.34556f
C501 two_stage_opamp_dummy_magic_0.cap_res_X.t69 GNDA 0.346812f
C502 two_stage_opamp_dummy_magic_0.cap_res_X.t128 GNDA 0.34556f
C503 two_stage_opamp_dummy_magic_0.cap_res_X.t22 GNDA 0.346812f
C504 two_stage_opamp_dummy_magic_0.cap_res_X.t4 GNDA 0.34556f
C505 two_stage_opamp_dummy_magic_0.cap_res_X.t109 GNDA 0.346812f
C506 two_stage_opamp_dummy_magic_0.cap_res_X.t94 GNDA 0.34556f
C507 two_stage_opamp_dummy_magic_0.cap_res_X.t129 GNDA 0.346812f
C508 two_stage_opamp_dummy_magic_0.cap_res_X.t111 GNDA 0.34556f
C509 two_stage_opamp_dummy_magic_0.cap_res_X.t76 GNDA 0.346812f
C510 two_stage_opamp_dummy_magic_0.cap_res_X.t135 GNDA 0.34556f
C511 two_stage_opamp_dummy_magic_0.cap_res_X.t28 GNDA 0.346812f
C512 two_stage_opamp_dummy_magic_0.cap_res_X.t11 GNDA 0.34556f
C513 two_stage_opamp_dummy_magic_0.cap_res_X.t117 GNDA 0.346812f
C514 two_stage_opamp_dummy_magic_0.cap_res_X.t34 GNDA 0.34556f
C515 two_stage_opamp_dummy_magic_0.cap_res_X.t68 GNDA 0.346812f
C516 two_stage_opamp_dummy_magic_0.cap_res_X.t50 GNDA 0.34556f
C517 two_stage_opamp_dummy_magic_0.cap_res_X.t16 GNDA 0.346812f
C518 two_stage_opamp_dummy_magic_0.cap_res_X.t73 GNDA 0.34556f
C519 two_stage_opamp_dummy_magic_0.cap_res_X.t108 GNDA 0.346812f
C520 two_stage_opamp_dummy_magic_0.cap_res_X.t91 GNDA 0.34556f
C521 two_stage_opamp_dummy_magic_0.cap_res_X.t54 GNDA 0.346812f
C522 two_stage_opamp_dummy_magic_0.cap_res_X.t36 GNDA 0.34556f
C523 two_stage_opamp_dummy_magic_0.cap_res_X.t74 GNDA 0.346812f
C524 two_stage_opamp_dummy_magic_0.cap_res_X.t53 GNDA 0.34556f
C525 two_stage_opamp_dummy_magic_0.cap_res_X.t20 GNDA 0.346812f
C526 two_stage_opamp_dummy_magic_0.cap_res_X.t78 GNDA 0.34556f
C527 two_stage_opamp_dummy_magic_0.cap_res_X.t116 GNDA 0.346812f
C528 two_stage_opamp_dummy_magic_0.cap_res_X.t97 GNDA 0.34556f
C529 two_stage_opamp_dummy_magic_0.cap_res_X.t57 GNDA 0.346812f
C530 two_stage_opamp_dummy_magic_0.cap_res_X.t120 GNDA 0.34556f
C531 two_stage_opamp_dummy_magic_0.cap_res_X.t15 GNDA 0.346812f
C532 two_stage_opamp_dummy_magic_0.cap_res_X.t137 GNDA 0.34556f
C533 two_stage_opamp_dummy_magic_0.cap_res_X.t100 GNDA 0.346812f
C534 two_stage_opamp_dummy_magic_0.cap_res_X.t85 GNDA 0.34556f
C535 two_stage_opamp_dummy_magic_0.cap_res_X.t119 GNDA 0.346812f
C536 two_stage_opamp_dummy_magic_0.cap_res_X.t84 GNDA 0.34556f
C537 two_stage_opamp_dummy_magic_0.cap_res_X.t8 GNDA 0.362503f
C538 two_stage_opamp_dummy_magic_0.cap_res_X.t41 GNDA 0.34556f
C539 two_stage_opamp_dummy_magic_0.cap_res_X.t99 GNDA 0.185607f
C540 two_stage_opamp_dummy_magic_0.cap_res_X.n0 GNDA 0.198646f
C541 two_stage_opamp_dummy_magic_0.cap_res_X.t93 GNDA 0.34556f
C542 two_stage_opamp_dummy_magic_0.cap_res_X.t60 GNDA 0.185607f
C543 two_stage_opamp_dummy_magic_0.cap_res_X.n1 GNDA 0.197043f
C544 two_stage_opamp_dummy_magic_0.cap_res_X.t3 GNDA 0.34556f
C545 two_stage_opamp_dummy_magic_0.cap_res_X.t26 GNDA 0.185607f
C546 two_stage_opamp_dummy_magic_0.cap_res_X.n2 GNDA 0.197043f
C547 two_stage_opamp_dummy_magic_0.cap_res_X.t51 GNDA 0.34556f
C548 two_stage_opamp_dummy_magic_0.cap_res_X.t133 GNDA 0.185607f
C549 two_stage_opamp_dummy_magic_0.cap_res_X.n3 GNDA 0.197043f
C550 two_stage_opamp_dummy_magic_0.cap_res_X.t14 GNDA 0.34556f
C551 two_stage_opamp_dummy_magic_0.cap_res_X.t82 GNDA 0.185607f
C552 two_stage_opamp_dummy_magic_0.cap_res_X.n4 GNDA 0.197043f
C553 two_stage_opamp_dummy_magic_0.cap_res_X.t61 GNDA 0.34556f
C554 two_stage_opamp_dummy_magic_0.cap_res_X.t44 GNDA 0.185607f
C555 two_stage_opamp_dummy_magic_0.cap_res_X.n5 GNDA 0.197043f
C556 two_stage_opamp_dummy_magic_0.cap_res_X.t115 GNDA 0.34556f
C557 two_stage_opamp_dummy_magic_0.cap_res_X.t13 GNDA 0.185607f
C558 two_stage_opamp_dummy_magic_0.cap_res_X.n6 GNDA 0.197043f
C559 two_stage_opamp_dummy_magic_0.cap_res_X.t71 GNDA 0.34556f
C560 two_stage_opamp_dummy_magic_0.cap_res_X.t103 GNDA 0.185607f
C561 two_stage_opamp_dummy_magic_0.cap_res_X.n7 GNDA 0.197043f
C562 two_stage_opamp_dummy_magic_0.cap_res_X.t123 GNDA 0.34556f
C563 two_stage_opamp_dummy_magic_0.cap_res_X.t63 GNDA 0.185607f
C564 two_stage_opamp_dummy_magic_0.cap_res_X.n8 GNDA 0.197043f
C565 two_stage_opamp_dummy_magic_0.cap_res_X.t40 GNDA 0.34556f
C566 two_stage_opamp_dummy_magic_0.cap_res_X.t132 GNDA 0.346812f
C567 two_stage_opamp_dummy_magic_0.cap_res_X.t33 GNDA 0.167062f
C568 two_stage_opamp_dummy_magic_0.cap_res_X.n9 GNDA 0.215485f
C569 two_stage_opamp_dummy_magic_0.cap_res_X.t30 GNDA 0.184458f
C570 two_stage_opamp_dummy_magic_0.cap_res_X.n10 GNDA 0.23403f
C571 two_stage_opamp_dummy_magic_0.cap_res_X.t64 GNDA 0.184458f
C572 two_stage_opamp_dummy_magic_0.cap_res_X.n11 GNDA 0.251323f
C573 two_stage_opamp_dummy_magic_0.cap_res_X.t24 GNDA 0.184458f
C574 two_stage_opamp_dummy_magic_0.cap_res_X.n12 GNDA 0.251323f
C575 two_stage_opamp_dummy_magic_0.cap_res_X.t126 GNDA 0.184458f
C576 two_stage_opamp_dummy_magic_0.cap_res_X.n13 GNDA 0.251323f
C577 two_stage_opamp_dummy_magic_0.cap_res_X.t19 GNDA 0.184458f
C578 two_stage_opamp_dummy_magic_0.cap_res_X.n14 GNDA 0.251323f
C579 two_stage_opamp_dummy_magic_0.cap_res_X.t122 GNDA 0.184458f
C580 two_stage_opamp_dummy_magic_0.cap_res_X.n15 GNDA 0.251323f
C581 two_stage_opamp_dummy_magic_0.cap_res_X.t80 GNDA 0.184458f
C582 two_stage_opamp_dummy_magic_0.cap_res_X.n16 GNDA 0.251323f
C583 two_stage_opamp_dummy_magic_0.cap_res_X.t37 GNDA 0.184458f
C584 two_stage_opamp_dummy_magic_0.cap_res_X.n17 GNDA 0.251323f
C585 two_stage_opamp_dummy_magic_0.cap_res_X.t75 GNDA 0.184458f
C586 two_stage_opamp_dummy_magic_0.cap_res_X.n18 GNDA 0.251323f
C587 two_stage_opamp_dummy_magic_0.cap_res_X.t35 GNDA 0.184458f
C588 two_stage_opamp_dummy_magic_0.cap_res_X.n19 GNDA 0.251323f
C589 two_stage_opamp_dummy_magic_0.cap_res_X.t138 GNDA 0.184458f
C590 two_stage_opamp_dummy_magic_0.cap_res_X.n20 GNDA 0.251323f
C591 two_stage_opamp_dummy_magic_0.cap_res_X.t29 GNDA 0.184458f
C592 two_stage_opamp_dummy_magic_0.cap_res_X.n21 GNDA 0.251323f
C593 two_stage_opamp_dummy_magic_0.cap_res_X.t131 GNDA 0.184458f
C594 two_stage_opamp_dummy_magic_0.cap_res_X.n22 GNDA 0.251323f
C595 two_stage_opamp_dummy_magic_0.cap_res_X.t110 GNDA 0.184458f
C596 two_stage_opamp_dummy_magic_0.cap_res_X.n23 GNDA 0.251323f
C597 two_stage_opamp_dummy_magic_0.cap_res_X.t5 GNDA 0.184458f
C598 two_stage_opamp_dummy_magic_0.cap_res_X.n24 GNDA 0.251323f
C599 two_stage_opamp_dummy_magic_0.cap_res_X.t106 GNDA 0.184458f
C600 two_stage_opamp_dummy_magic_0.cap_res_X.n25 GNDA 0.23403f
C601 two_stage_opamp_dummy_magic_0.cap_res_X.t104 GNDA 0.344411f
C602 two_stage_opamp_dummy_magic_0.cap_res_X.t2 GNDA 0.167062f
C603 two_stage_opamp_dummy_magic_0.cap_res_X.n26 GNDA 0.216737f
C604 two_stage_opamp_dummy_magic_0.cap_res_X.t1 GNDA 0.344411f
C605 two_stage_opamp_dummy_magic_0.cap_res_X.t38 GNDA 0.167062f
C606 two_stage_opamp_dummy_magic_0.cap_res_X.n27 GNDA 0.216737f
C607 two_stage_opamp_dummy_magic_0.cap_res_X.t121 GNDA 0.344411f
C608 two_stage_opamp_dummy_magic_0.cap_res_X.t113 GNDA 0.34556f
C609 two_stage_opamp_dummy_magic_0.cap_res_X.t21 GNDA 0.364105f
C610 two_stage_opamp_dummy_magic_0.cap_res_X.t56 GNDA 0.364105f
C611 two_stage_opamp_dummy_magic_0.cap_res_X.t18 GNDA 0.185607f
C612 two_stage_opamp_dummy_magic_0.cap_res_X.n28 GNDA 0.216737f
C613 two_stage_opamp_dummy_magic_0.cap_res_X.t125 GNDA 0.344411f
C614 two_stage_opamp_dummy_magic_0.cap_res_X.t62 GNDA 0.34556f
C615 two_stage_opamp_dummy_magic_0.cap_res_X.t23 GNDA 0.185607f
C616 two_stage_opamp_dummy_magic_0.cap_res_X.n29 GNDA 0.198192f
C617 two_stage_opamp_dummy_magic_0.cap_res_X.t7 GNDA 0.344411f
C618 two_stage_opamp_dummy_magic_0.cap_res_X.t87 GNDA 0.34556f
C619 two_stage_opamp_dummy_magic_0.cap_res_X.t46 GNDA 0.185607f
C620 two_stage_opamp_dummy_magic_0.cap_res_X.n30 GNDA 0.216737f
C621 two_stage_opamp_dummy_magic_0.cap_res_X.t107 GNDA 0.344411f
C622 two_stage_opamp_dummy_magic_0.cap_res_X.t47 GNDA 0.34556f
C623 two_stage_opamp_dummy_magic_0.cap_res_X.t10 GNDA 0.185607f
C624 two_stage_opamp_dummy_magic_0.cap_res_X.n31 GNDA 0.216737f
C625 two_stage_opamp_dummy_magic_0.cap_res_X.t70 GNDA 0.344411f
C626 two_stage_opamp_dummy_magic_0.cap_res_X.t12 GNDA 0.34556f
C627 two_stage_opamp_dummy_magic_0.cap_res_X.t112 GNDA 0.185607f
C628 two_stage_opamp_dummy_magic_0.cap_res_X.n32 GNDA 0.216737f
C629 two_stage_opamp_dummy_magic_0.cap_res_X.t32 GNDA 0.344411f
C630 two_stage_opamp_dummy_magic_0.cap_res_X.t92 GNDA 0.34556f
C631 two_stage_opamp_dummy_magic_0.cap_res_X.t77 GNDA 0.364105f
C632 two_stage_opamp_dummy_magic_0.cap_res_X.t114 GNDA 0.364105f
C633 two_stage_opamp_dummy_magic_0.cap_res_X.t72 GNDA 0.185607f
C634 two_stage_opamp_dummy_magic_0.cap_res_X.n33 GNDA 0.216737f
C635 two_stage_opamp_dummy_magic_0.cap_res_X.t52 GNDA 0.344411f
C636 two_stage_opamp_dummy_magic_0.cap_res_X.t39 GNDA 0.34556f
C637 two_stage_opamp_dummy_magic_0.cap_res_X.t101 GNDA 0.364105f
C638 two_stage_opamp_dummy_magic_0.cap_res_X.t136 GNDA 0.364105f
C639 two_stage_opamp_dummy_magic_0.cap_res_X.t96 GNDA 0.185607f
C640 two_stage_opamp_dummy_magic_0.cap_res_X.n34 GNDA 0.216737f
C641 two_stage_opamp_dummy_magic_0.cap_res_X.t17 GNDA 0.344411f
C642 two_stage_opamp_dummy_magic_0.cap_res_X.n35 GNDA 0.216737f
C643 two_stage_opamp_dummy_magic_0.cap_res_X.t55 GNDA 0.185607f
C644 two_stage_opamp_dummy_magic_0.cap_res_X.t98 GNDA 0.364105f
C645 two_stage_opamp_dummy_magic_0.cap_res_X.t59 GNDA 0.364105f
C646 two_stage_opamp_dummy_magic_0.cap_res_X.t6 GNDA 0.738067f
C647 two_stage_opamp_dummy_magic_0.cap_res_X.t0 GNDA 0.298118f
C648 two_stage_opamp_dummy_magic_0.VD1.t9 GNDA 0.053331f
C649 two_stage_opamp_dummy_magic_0.VD1.n0 GNDA 0.203944f
C650 two_stage_opamp_dummy_magic_0.VD1.t7 GNDA 0.053331f
C651 two_stage_opamp_dummy_magic_0.VD1.t12 GNDA 0.053331f
C652 two_stage_opamp_dummy_magic_0.VD1.n1 GNDA 0.116042f
C653 two_stage_opamp_dummy_magic_0.VD1.n2 GNDA 0.461069f
C654 two_stage_opamp_dummy_magic_0.VD1.n3 GNDA 0.192793f
C655 two_stage_opamp_dummy_magic_0.VD1.t5 GNDA 0.053331f
C656 two_stage_opamp_dummy_magic_0.VD1.t10 GNDA 0.053331f
C657 two_stage_opamp_dummy_magic_0.VD1.n4 GNDA 0.116042f
C658 two_stage_opamp_dummy_magic_0.VD1.n5 GNDA 0.461069f
C659 two_stage_opamp_dummy_magic_0.VD1.t6 GNDA 0.053331f
C660 two_stage_opamp_dummy_magic_0.VD1.t11 GNDA 0.053331f
C661 two_stage_opamp_dummy_magic_0.VD1.n6 GNDA 0.116042f
C662 two_stage_opamp_dummy_magic_0.VD1.n7 GNDA 0.442486f
C663 two_stage_opamp_dummy_magic_0.VD1.n8 GNDA 0.203944f
C664 two_stage_opamp_dummy_magic_0.VD1.n9 GNDA 0.119128f
C665 two_stage_opamp_dummy_magic_0.VD1.t13 GNDA 0.053331f
C666 two_stage_opamp_dummy_magic_0.VD1.t8 GNDA 0.053331f
C667 two_stage_opamp_dummy_magic_0.VD1.n10 GNDA 0.116042f
C668 two_stage_opamp_dummy_magic_0.VD1.n11 GNDA 0.361396f
C669 two_stage_opamp_dummy_magic_0.VD1.n12 GNDA 0.099935f
C670 two_stage_opamp_dummy_magic_0.VD1.n13 GNDA 0.205342f
C671 two_stage_opamp_dummy_magic_0.VD1.t19 GNDA 0.053331f
C672 two_stage_opamp_dummy_magic_0.VD1.t16 GNDA 0.053331f
C673 two_stage_opamp_dummy_magic_0.VD1.n14 GNDA 0.116042f
C674 two_stage_opamp_dummy_magic_0.VD1.n15 GNDA 0.465721f
C675 two_stage_opamp_dummy_magic_0.VD1.n16 GNDA 0.205342f
C676 two_stage_opamp_dummy_magic_0.VD1.t20 GNDA 0.053331f
C677 two_stage_opamp_dummy_magic_0.VD1.t3 GNDA 0.053331f
C678 two_stage_opamp_dummy_magic_0.VD1.n17 GNDA 0.116042f
C679 two_stage_opamp_dummy_magic_0.VD1.n18 GNDA 0.447102f
C680 two_stage_opamp_dummy_magic_0.VD1.n19 GNDA 0.192793f
C681 two_stage_opamp_dummy_magic_0.VD1.t2 GNDA 0.053331f
C682 two_stage_opamp_dummy_magic_0.VD1.t17 GNDA 0.053331f
C683 two_stage_opamp_dummy_magic_0.VD1.n20 GNDA 0.116042f
C684 two_stage_opamp_dummy_magic_0.VD1.n21 GNDA 0.447102f
C685 two_stage_opamp_dummy_magic_0.VD1.n22 GNDA 0.113419f
C686 two_stage_opamp_dummy_magic_0.VD1.t1 GNDA 0.053331f
C687 two_stage_opamp_dummy_magic_0.VD1.t18 GNDA 0.053331f
C688 two_stage_opamp_dummy_magic_0.VD1.n23 GNDA 0.116042f
C689 two_stage_opamp_dummy_magic_0.VD1.n24 GNDA 0.465721f
C690 two_stage_opamp_dummy_magic_0.VD1.t21 GNDA 0.053331f
C691 two_stage_opamp_dummy_magic_0.VD1.t0 GNDA 0.053331f
C692 two_stage_opamp_dummy_magic_0.VD1.n25 GNDA 0.116042f
C693 two_stage_opamp_dummy_magic_0.VD1.n26 GNDA 0.447102f
C694 two_stage_opamp_dummy_magic_0.VD1.n27 GNDA 0.192793f
C695 two_stage_opamp_dummy_magic_0.VD1.n28 GNDA 0.113419f
C696 two_stage_opamp_dummy_magic_0.VD1.t15 GNDA 0.053331f
C697 two_stage_opamp_dummy_magic_0.VD1.t4 GNDA 0.053331f
C698 two_stage_opamp_dummy_magic_0.VD1.n29 GNDA 0.116042f
C699 two_stage_opamp_dummy_magic_0.VD1.n30 GNDA 0.447102f
C700 two_stage_opamp_dummy_magic_0.VD1.n31 GNDA 0.099935f
C701 two_stage_opamp_dummy_magic_0.VD1.n32 GNDA 0.08441f
C702 two_stage_opamp_dummy_magic_0.VD1.n33 GNDA 0.235249f
C703 two_stage_opamp_dummy_magic_0.VD1.n34 GNDA 0.106662f
C704 two_stage_opamp_dummy_magic_0.VD1.n35 GNDA 0.192793f
C705 two_stage_opamp_dummy_magic_0.VD1.n36 GNDA 0.442486f
C706 two_stage_opamp_dummy_magic_0.VD1.n37 GNDA 0.116042f
C707 two_stage_opamp_dummy_magic_0.VD1.t14 GNDA 0.053331f
C708 two_stage_opamp_dummy_magic_0.X.t16 GNDA 0.03768f
C709 two_stage_opamp_dummy_magic_0.X.t17 GNDA 0.03768f
C710 two_stage_opamp_dummy_magic_0.X.n0 GNDA 0.081988f
C711 two_stage_opamp_dummy_magic_0.X.n1 GNDA 0.25534f
C712 two_stage_opamp_dummy_magic_0.X.n2 GNDA 0.136216f
C713 two_stage_opamp_dummy_magic_0.X.n3 GNDA 0.136215f
C714 two_stage_opamp_dummy_magic_0.X.t22 GNDA 0.03768f
C715 two_stage_opamp_dummy_magic_0.X.t20 GNDA 0.03768f
C716 two_stage_opamp_dummy_magic_0.X.n4 GNDA 0.081988f
C717 two_stage_opamp_dummy_magic_0.X.n5 GNDA 0.325763f
C718 two_stage_opamp_dummy_magic_0.X.t13 GNDA 0.03768f
C719 two_stage_opamp_dummy_magic_0.X.t14 GNDA 0.03768f
C720 two_stage_opamp_dummy_magic_0.X.n6 GNDA 0.081988f
C721 two_stage_opamp_dummy_magic_0.X.n7 GNDA 0.312634f
C722 two_stage_opamp_dummy_magic_0.X.n8 GNDA 0.144094f
C723 two_stage_opamp_dummy_magic_0.X.n9 GNDA 0.084168f
C724 two_stage_opamp_dummy_magic_0.X.t15 GNDA 0.03768f
C725 two_stage_opamp_dummy_magic_0.X.t23 GNDA 0.03768f
C726 two_stage_opamp_dummy_magic_0.X.n10 GNDA 0.081988f
C727 two_stage_opamp_dummy_magic_0.X.n11 GNDA 0.325763f
C728 two_stage_opamp_dummy_magic_0.X.t18 GNDA 0.03768f
C729 two_stage_opamp_dummy_magic_0.X.t12 GNDA 0.03768f
C730 two_stage_opamp_dummy_magic_0.X.n12 GNDA 0.081988f
C731 two_stage_opamp_dummy_magic_0.X.n13 GNDA 0.312634f
C732 two_stage_opamp_dummy_magic_0.X.n14 GNDA 0.144094f
C733 two_stage_opamp_dummy_magic_0.X.n15 GNDA 0.084168f
C734 two_stage_opamp_dummy_magic_0.X.t19 GNDA 0.03768f
C735 two_stage_opamp_dummy_magic_0.X.t21 GNDA 0.03768f
C736 two_stage_opamp_dummy_magic_0.X.n16 GNDA 0.081988f
C737 two_stage_opamp_dummy_magic_0.X.n17 GNDA 0.312634f
C738 two_stage_opamp_dummy_magic_0.X.n18 GNDA 0.080135f
C739 two_stage_opamp_dummy_magic_0.X.n19 GNDA 0.075361f
C740 two_stage_opamp_dummy_magic_0.X.n20 GNDA 0.156078f
C741 two_stage_opamp_dummy_magic_0.X.t11 GNDA 1.21356f
C742 two_stage_opamp_dummy_magic_0.X.t32 GNDA 0.165794f
C743 two_stage_opamp_dummy_magic_0.X.t47 GNDA 0.165794f
C744 two_stage_opamp_dummy_magic_0.X.t28 GNDA 0.165794f
C745 two_stage_opamp_dummy_magic_0.X.t43 GNDA 0.165794f
C746 two_stage_opamp_dummy_magic_0.X.t26 GNDA 0.165794f
C747 two_stage_opamp_dummy_magic_0.X.t41 GNDA 0.176582f
C748 two_stage_opamp_dummy_magic_0.X.n21 GNDA 0.139934f
C749 two_stage_opamp_dummy_magic_0.X.n22 GNDA 0.079129f
C750 two_stage_opamp_dummy_magic_0.X.n23 GNDA 0.079129f
C751 two_stage_opamp_dummy_magic_0.X.n24 GNDA 0.079129f
C752 two_stage_opamp_dummy_magic_0.X.t50 GNDA 0.165794f
C753 two_stage_opamp_dummy_magic_0.X.t35 GNDA 0.165794f
C754 two_stage_opamp_dummy_magic_0.X.t49 GNDA 0.165794f
C755 two_stage_opamp_dummy_magic_0.X.t34 GNDA 0.176582f
C756 two_stage_opamp_dummy_magic_0.X.n25 GNDA 0.139934f
C757 two_stage_opamp_dummy_magic_0.X.n26 GNDA 0.079129f
C758 two_stage_opamp_dummy_magic_0.X.n27 GNDA 0.079129f
C759 two_stage_opamp_dummy_magic_0.X.n28 GNDA 0.117701f
C760 two_stage_opamp_dummy_magic_0.X.n29 GNDA 1.3031f
C761 two_stage_opamp_dummy_magic_0.X.n30 GNDA 0.101322f
C762 two_stage_opamp_dummy_magic_0.X.n31 GNDA 0.095366f
C763 two_stage_opamp_dummy_magic_0.X.t4 GNDA 0.087921f
C764 two_stage_opamp_dummy_magic_0.X.t24 GNDA 0.087921f
C765 two_stage_opamp_dummy_magic_0.X.n32 GNDA 0.179851f
C766 two_stage_opamp_dummy_magic_0.X.n33 GNDA 0.610627f
C767 two_stage_opamp_dummy_magic_0.X.n34 GNDA 0.162684f
C768 two_stage_opamp_dummy_magic_0.X.t3 GNDA 0.087921f
C769 two_stage_opamp_dummy_magic_0.X.t2 GNDA 0.087921f
C770 two_stage_opamp_dummy_magic_0.X.n35 GNDA 0.179851f
C771 two_stage_opamp_dummy_magic_0.X.n36 GNDA 0.59436f
C772 two_stage_opamp_dummy_magic_0.X.n37 GNDA 0.17423f
C773 two_stage_opamp_dummy_magic_0.X.t6 GNDA 0.087921f
C774 two_stage_opamp_dummy_magic_0.X.t1 GNDA 0.087921f
C775 two_stage_opamp_dummy_magic_0.X.n38 GNDA 0.179851f
C776 two_stage_opamp_dummy_magic_0.X.n39 GNDA 0.59436f
C777 two_stage_opamp_dummy_magic_0.X.n40 GNDA 0.101322f
C778 two_stage_opamp_dummy_magic_0.X.n41 GNDA 0.101322f
C779 two_stage_opamp_dummy_magic_0.X.t9 GNDA 0.087921f
C780 two_stage_opamp_dummy_magic_0.X.t0 GNDA 0.087921f
C781 two_stage_opamp_dummy_magic_0.X.n42 GNDA 0.179851f
C782 two_stage_opamp_dummy_magic_0.X.n43 GNDA 0.59436f
C783 two_stage_opamp_dummy_magic_0.X.n44 GNDA 0.095366f
C784 two_stage_opamp_dummy_magic_0.X.t7 GNDA 0.087921f
C785 two_stage_opamp_dummy_magic_0.X.t8 GNDA 0.087921f
C786 two_stage_opamp_dummy_magic_0.X.n45 GNDA 0.179851f
C787 two_stage_opamp_dummy_magic_0.X.n46 GNDA 0.59436f
C788 two_stage_opamp_dummy_magic_0.X.n47 GNDA 0.162684f
C789 two_stage_opamp_dummy_magic_0.X.t10 GNDA 0.087921f
C790 two_stage_opamp_dummy_magic_0.X.t5 GNDA 0.087921f
C791 two_stage_opamp_dummy_magic_0.X.n48 GNDA 0.179851f
C792 two_stage_opamp_dummy_magic_0.X.n49 GNDA 0.602311f
C793 two_stage_opamp_dummy_magic_0.X.n50 GNDA 0.395522f
C794 two_stage_opamp_dummy_magic_0.X.t36 GNDA 0.052753f
C795 two_stage_opamp_dummy_magic_0.X.t51 GNDA 0.052753f
C796 two_stage_opamp_dummy_magic_0.X.t33 GNDA 0.052753f
C797 two_stage_opamp_dummy_magic_0.X.t48 GNDA 0.052753f
C798 two_stage_opamp_dummy_magic_0.X.t29 GNDA 0.052753f
C799 two_stage_opamp_dummy_magic_0.X.t44 GNDA 0.064057f
C800 two_stage_opamp_dummy_magic_0.X.n51 GNDA 0.064057f
C801 two_stage_opamp_dummy_magic_0.X.n52 GNDA 0.041448f
C802 two_stage_opamp_dummy_magic_0.X.n53 GNDA 0.041448f
C803 two_stage_opamp_dummy_magic_0.X.n54 GNDA 0.041448f
C804 two_stage_opamp_dummy_magic_0.X.t53 GNDA 0.052753f
C805 two_stage_opamp_dummy_magic_0.X.t39 GNDA 0.052753f
C806 two_stage_opamp_dummy_magic_0.X.t52 GNDA 0.052753f
C807 two_stage_opamp_dummy_magic_0.X.t38 GNDA 0.064057f
C808 two_stage_opamp_dummy_magic_0.X.n55 GNDA 0.064057f
C809 two_stage_opamp_dummy_magic_0.X.n56 GNDA 0.041448f
C810 two_stage_opamp_dummy_magic_0.X.n57 GNDA 0.041448f
C811 two_stage_opamp_dummy_magic_0.X.n58 GNDA 0.069677f
C812 two_stage_opamp_dummy_magic_0.X.t27 GNDA 0.081013f
C813 two_stage_opamp_dummy_magic_0.X.t42 GNDA 0.081013f
C814 two_stage_opamp_dummy_magic_0.X.t25 GNDA 0.081013f
C815 two_stage_opamp_dummy_magic_0.X.t40 GNDA 0.081013f
C816 two_stage_opamp_dummy_magic_0.X.t54 GNDA 0.081013f
C817 two_stage_opamp_dummy_magic_0.X.t37 GNDA 0.092098f
C818 two_stage_opamp_dummy_magic_0.X.n59 GNDA 0.083116f
C819 two_stage_opamp_dummy_magic_0.X.n60 GNDA 0.050869f
C820 two_stage_opamp_dummy_magic_0.X.n61 GNDA 0.050869f
C821 two_stage_opamp_dummy_magic_0.X.n62 GNDA 0.050869f
C822 two_stage_opamp_dummy_magic_0.X.t46 GNDA 0.081013f
C823 two_stage_opamp_dummy_magic_0.X.t31 GNDA 0.081013f
C824 two_stage_opamp_dummy_magic_0.X.t45 GNDA 0.081013f
C825 two_stage_opamp_dummy_magic_0.X.t30 GNDA 0.092098f
C826 two_stage_opamp_dummy_magic_0.X.n63 GNDA 0.083116f
C827 two_stage_opamp_dummy_magic_0.X.n64 GNDA 0.050869f
C828 two_stage_opamp_dummy_magic_0.X.n65 GNDA 0.050869f
C829 two_stage_opamp_dummy_magic_0.X.n66 GNDA 0.077245f
C830 two_stage_opamp_dummy_magic_0.X.n67 GNDA 0.113576f
C831 two_stage_opamp_dummy_magic_0.X.n68 GNDA 1.07875f
C832 two_stage_opamp_dummy_magic_0.X.n69 GNDA 0.369903f
C833 two_stage_opamp_dummy_magic_0.X.n70 GNDA 0.20931f
C834 two_stage_opamp_dummy_magic_0.V_err_p.t8 GNDA 0.026629f
C835 two_stage_opamp_dummy_magic_0.V_err_p.n0 GNDA 0.437635f
C836 two_stage_opamp_dummy_magic_0.V_err_p.t2 GNDA 0.026629f
C837 two_stage_opamp_dummy_magic_0.V_err_p.t9 GNDA 0.026629f
C838 two_stage_opamp_dummy_magic_0.V_err_p.n1 GNDA 0.054258f
C839 two_stage_opamp_dummy_magic_0.V_err_p.n2 GNDA 0.267929f
C840 two_stage_opamp_dummy_magic_0.V_err_p.n3 GNDA 0.169075f
C841 two_stage_opamp_dummy_magic_0.V_err_p.t6 GNDA 0.026629f
C842 two_stage_opamp_dummy_magic_0.V_err_p.t21 GNDA 0.026629f
C843 two_stage_opamp_dummy_magic_0.V_err_p.n4 GNDA 0.054258f
C844 two_stage_opamp_dummy_magic_0.V_err_p.n5 GNDA 0.399818f
C845 two_stage_opamp_dummy_magic_0.V_err_p.n6 GNDA 0.287184f
C846 two_stage_opamp_dummy_magic_0.V_err_p.t1 GNDA 0.026629f
C847 two_stage_opamp_dummy_magic_0.V_err_p.t4 GNDA 0.026629f
C848 two_stage_opamp_dummy_magic_0.V_err_p.n7 GNDA 0.054258f
C849 two_stage_opamp_dummy_magic_0.V_err_p.n8 GNDA 0.37261f
C850 two_stage_opamp_dummy_magic_0.V_err_p.n9 GNDA 0.275151f
C851 two_stage_opamp_dummy_magic_0.V_err_p.t5 GNDA 0.026629f
C852 two_stage_opamp_dummy_magic_0.V_err_p.t0 GNDA 0.026629f
C853 two_stage_opamp_dummy_magic_0.V_err_p.n10 GNDA 0.054258f
C854 two_stage_opamp_dummy_magic_0.V_err_p.n11 GNDA 0.37261f
C855 two_stage_opamp_dummy_magic_0.V_err_p.n12 GNDA 0.162976f
C856 two_stage_opamp_dummy_magic_0.V_err_p.n13 GNDA 0.275151f
C857 two_stage_opamp_dummy_magic_0.V_err_p.t10 GNDA 0.026629f
C858 two_stage_opamp_dummy_magic_0.V_err_p.t3 GNDA 0.026629f
C859 two_stage_opamp_dummy_magic_0.V_err_p.n14 GNDA 0.054258f
C860 two_stage_opamp_dummy_magic_0.V_err_p.n15 GNDA 0.37261f
C861 two_stage_opamp_dummy_magic_0.V_err_p.n16 GNDA 0.277957f
C862 two_stage_opamp_dummy_magic_0.V_err_p.n17 GNDA 0.42243f
C863 two_stage_opamp_dummy_magic_0.V_err_p.n18 GNDA 0.280143f
C864 two_stage_opamp_dummy_magic_0.V_err_p.t15 GNDA 0.026629f
C865 two_stage_opamp_dummy_magic_0.V_err_p.t7 GNDA 0.026629f
C866 two_stage_opamp_dummy_magic_0.V_err_p.n19 GNDA 0.054258f
C867 two_stage_opamp_dummy_magic_0.V_err_p.n20 GNDA 0.450528f
C868 two_stage_opamp_dummy_magic_0.V_err_p.n21 GNDA 0.42549f
C869 two_stage_opamp_dummy_magic_0.V_err_p.t18 GNDA 0.026629f
C870 two_stage_opamp_dummy_magic_0.V_err_p.t13 GNDA 0.026629f
C871 two_stage_opamp_dummy_magic_0.V_err_p.n22 GNDA 0.054258f
C872 two_stage_opamp_dummy_magic_0.V_err_p.n23 GNDA 0.37261f
C873 two_stage_opamp_dummy_magic_0.V_err_p.n24 GNDA 0.437635f
C874 two_stage_opamp_dummy_magic_0.V_err_p.t11 GNDA 0.026629f
C875 two_stage_opamp_dummy_magic_0.V_err_p.t16 GNDA 0.026629f
C876 two_stage_opamp_dummy_magic_0.V_err_p.n25 GNDA 0.054258f
C877 two_stage_opamp_dummy_magic_0.V_err_p.n26 GNDA 0.37261f
C878 two_stage_opamp_dummy_magic_0.V_err_p.n27 GNDA 0.286242f
C879 two_stage_opamp_dummy_magic_0.V_err_p.n28 GNDA 0.286242f
C880 two_stage_opamp_dummy_magic_0.V_err_p.t12 GNDA 0.026629f
C881 two_stage_opamp_dummy_magic_0.V_err_p.t17 GNDA 0.026629f
C882 two_stage_opamp_dummy_magic_0.V_err_p.n29 GNDA 0.054258f
C883 two_stage_opamp_dummy_magic_0.V_err_p.n30 GNDA 0.37261f
C884 two_stage_opamp_dummy_magic_0.V_err_p.n31 GNDA 0.280143f
C885 two_stage_opamp_dummy_magic_0.V_err_p.t14 GNDA 0.026629f
C886 two_stage_opamp_dummy_magic_0.V_err_p.t19 GNDA 0.026629f
C887 two_stage_opamp_dummy_magic_0.V_err_p.n32 GNDA 0.054258f
C888 two_stage_opamp_dummy_magic_0.V_err_p.n33 GNDA 0.37261f
C889 two_stage_opamp_dummy_magic_0.V_err_p.n34 GNDA 0.280143f
C890 two_stage_opamp_dummy_magic_0.V_err_p.n35 GNDA 0.395596f
C891 two_stage_opamp_dummy_magic_0.V_err_p.n36 GNDA 0.411595f
C892 two_stage_opamp_dummy_magic_0.V_err_p.n37 GNDA 0.054258f
C893 two_stage_opamp_dummy_magic_0.V_err_p.t20 GNDA 0.026629f
C894 two_stage_opamp_dummy_magic_0.V_err_gate.n0 GNDA 0.302465f
C895 two_stage_opamp_dummy_magic_0.V_err_gate.n1 GNDA 0.302465f
C896 two_stage_opamp_dummy_magic_0.V_err_gate.n2 GNDA 0.276018f
C897 two_stage_opamp_dummy_magic_0.V_err_gate.n3 GNDA 0.372156f
C898 two_stage_opamp_dummy_magic_0.V_err_gate.n4 GNDA 0.19826f
C899 two_stage_opamp_dummy_magic_0.V_err_gate.n5 GNDA 0.233445f
C900 two_stage_opamp_dummy_magic_0.V_err_gate.t9 GNDA 0.036767f
C901 two_stage_opamp_dummy_magic_0.V_err_gate.t10 GNDA 0.036767f
C902 two_stage_opamp_dummy_magic_0.V_err_gate.n6 GNDA 0.674676f
C903 two_stage_opamp_dummy_magic_0.V_err_gate.t30 GNDA 0.015166f
C904 two_stage_opamp_dummy_magic_0.V_err_gate.t23 GNDA 0.015166f
C905 two_stage_opamp_dummy_magic_0.V_err_gate.t33 GNDA 0.015166f
C906 two_stage_opamp_dummy_magic_0.V_err_gate.t20 GNDA 0.015166f
C907 two_stage_opamp_dummy_magic_0.V_err_gate.t29 GNDA 0.015166f
C908 two_stage_opamp_dummy_magic_0.V_err_gate.t18 GNDA 0.015166f
C909 two_stage_opamp_dummy_magic_0.V_err_gate.t27 GNDA 0.015166f
C910 two_stage_opamp_dummy_magic_0.V_err_gate.t16 GNDA 0.015166f
C911 two_stage_opamp_dummy_magic_0.V_err_gate.t24 GNDA 0.015166f
C912 two_stage_opamp_dummy_magic_0.V_err_gate.t31 GNDA 0.015166f
C913 two_stage_opamp_dummy_magic_0.V_err_gate.t25 GNDA 0.015166f
C914 two_stage_opamp_dummy_magic_0.V_err_gate.t14 GNDA 0.03286f
C915 two_stage_opamp_dummy_magic_0.V_err_gate.n7 GNDA 0.051244f
C916 two_stage_opamp_dummy_magic_0.V_err_gate.n8 GNDA 0.039984f
C917 two_stage_opamp_dummy_magic_0.V_err_gate.n9 GNDA 0.039984f
C918 two_stage_opamp_dummy_magic_0.V_err_gate.n10 GNDA 0.039984f
C919 two_stage_opamp_dummy_magic_0.V_err_gate.n11 GNDA 0.039984f
C920 two_stage_opamp_dummy_magic_0.V_err_gate.n12 GNDA 0.039984f
C921 two_stage_opamp_dummy_magic_0.V_err_gate.n13 GNDA 0.039984f
C922 two_stage_opamp_dummy_magic_0.V_err_gate.n14 GNDA 0.039984f
C923 two_stage_opamp_dummy_magic_0.V_err_gate.n15 GNDA 0.039984f
C924 two_stage_opamp_dummy_magic_0.V_err_gate.n16 GNDA 0.039984f
C925 two_stage_opamp_dummy_magic_0.V_err_gate.t21 GNDA 0.015166f
C926 two_stage_opamp_dummy_magic_0.V_err_gate.t15 GNDA 0.015166f
C927 two_stage_opamp_dummy_magic_0.V_err_gate.t26 GNDA 0.015166f
C928 two_stage_opamp_dummy_magic_0.V_err_gate.t17 GNDA 0.015166f
C929 two_stage_opamp_dummy_magic_0.V_err_gate.t28 GNDA 0.015166f
C930 two_stage_opamp_dummy_magic_0.V_err_gate.t19 GNDA 0.015166f
C931 two_stage_opamp_dummy_magic_0.V_err_gate.t32 GNDA 0.015166f
C932 two_stage_opamp_dummy_magic_0.V_err_gate.t22 GNDA 0.03286f
C933 two_stage_opamp_dummy_magic_0.V_err_gate.n17 GNDA 0.051244f
C934 two_stage_opamp_dummy_magic_0.V_err_gate.n18 GNDA 0.039984f
C935 two_stage_opamp_dummy_magic_0.V_err_gate.n19 GNDA 0.039984f
C936 two_stage_opamp_dummy_magic_0.V_err_gate.n20 GNDA 0.039984f
C937 two_stage_opamp_dummy_magic_0.V_err_gate.n21 GNDA 0.039984f
C938 two_stage_opamp_dummy_magic_0.V_err_gate.n22 GNDA 0.039984f
C939 two_stage_opamp_dummy_magic_0.V_err_gate.n23 GNDA 0.039984f
C940 two_stage_opamp_dummy_magic_0.V_err_gate.n24 GNDA 0.102015f
C941 two_stage_opamp_dummy_magic_0.V_err_gate.t4 GNDA 0.018383f
C942 two_stage_opamp_dummy_magic_0.V_err_gate.t8 GNDA 0.018383f
C943 two_stage_opamp_dummy_magic_0.V_err_gate.n25 GNDA 0.037457f
C944 two_stage_opamp_dummy_magic_0.V_err_gate.t13 GNDA 0.018383f
C945 two_stage_opamp_dummy_magic_0.V_err_gate.t0 GNDA 0.018383f
C946 two_stage_opamp_dummy_magic_0.V_err_gate.n26 GNDA 0.037457f
C947 two_stage_opamp_dummy_magic_0.V_err_gate.n27 GNDA 0.257235f
C948 two_stage_opamp_dummy_magic_0.V_err_gate.t5 GNDA 0.018383f
C949 two_stage_opamp_dummy_magic_0.V_err_gate.t3 GNDA 0.018383f
C950 two_stage_opamp_dummy_magic_0.V_err_gate.n28 GNDA 0.037457f
C951 two_stage_opamp_dummy_magic_0.V_err_gate.n29 GNDA 0.257235f
C952 two_stage_opamp_dummy_magic_0.V_err_gate.t11 GNDA 0.018383f
C953 two_stage_opamp_dummy_magic_0.V_err_gate.t12 GNDA 0.018383f
C954 two_stage_opamp_dummy_magic_0.V_err_gate.n30 GNDA 0.037457f
C955 two_stage_opamp_dummy_magic_0.V_err_gate.n31 GNDA 0.257235f
C956 two_stage_opamp_dummy_magic_0.V_err_gate.t6 GNDA 0.018383f
C957 two_stage_opamp_dummy_magic_0.V_err_gate.t2 GNDA 0.018383f
C958 two_stage_opamp_dummy_magic_0.V_err_gate.n32 GNDA 0.037457f
C959 two_stage_opamp_dummy_magic_0.V_err_gate.n33 GNDA 0.257235f
C960 two_stage_opamp_dummy_magic_0.V_err_gate.t7 GNDA 0.018383f
C961 two_stage_opamp_dummy_magic_0.V_err_gate.t1 GNDA 0.018383f
C962 two_stage_opamp_dummy_magic_0.V_err_gate.n34 GNDA 0.037457f
C963 two_stage_opamp_dummy_magic_0.V_err_gate.n35 GNDA 0.266569f
C964 two_stage_opamp_dummy_magic_0.Vb1.n0 GNDA 0.085417f
C965 two_stage_opamp_dummy_magic_0.Vb1.n1 GNDA 0.236102f
C966 two_stage_opamp_dummy_magic_0.Vb1.t1 GNDA 0.016179f
C967 two_stage_opamp_dummy_magic_0.Vb1.t13 GNDA 0.016179f
C968 two_stage_opamp_dummy_magic_0.Vb1.n2 GNDA 0.034871f
C969 two_stage_opamp_dummy_magic_0.Vb1.t12 GNDA 0.016179f
C970 two_stage_opamp_dummy_magic_0.Vb1.t0 GNDA 0.016179f
C971 two_stage_opamp_dummy_magic_0.Vb1.n3 GNDA 0.034652f
C972 two_stage_opamp_dummy_magic_0.Vb1.n4 GNDA 0.626025f
C973 two_stage_opamp_dummy_magic_0.Vb1.t23 GNDA 0.024875f
C974 two_stage_opamp_dummy_magic_0.Vb1.t32 GNDA 0.024875f
C975 two_stage_opamp_dummy_magic_0.Vb1.t21 GNDA 0.024875f
C976 two_stage_opamp_dummy_magic_0.Vb1.t30 GNDA 0.024875f
C977 two_stage_opamp_dummy_magic_0.Vb1.t26 GNDA 0.024875f
C978 two_stage_opamp_dummy_magic_0.Vb1.t15 GNDA 0.024875f
C979 two_stage_opamp_dummy_magic_0.Vb1.t25 GNDA 0.024875f
C980 two_stage_opamp_dummy_magic_0.Vb1.t14 GNDA 0.024875f
C981 two_stage_opamp_dummy_magic_0.Vb1.t17 GNDA 0.024875f
C982 two_stage_opamp_dummy_magic_0.Vb1.t27 GNDA 0.024875f
C983 two_stage_opamp_dummy_magic_0.Vb1.t9 GNDA 0.024268f
C984 two_stage_opamp_dummy_magic_0.Vb1.t11 GNDA 0.024268f
C985 two_stage_opamp_dummy_magic_0.Vb1.n5 GNDA 0.052805f
C986 two_stage_opamp_dummy_magic_0.Vb1.n6 GNDA 0.216328f
C987 two_stage_opamp_dummy_magic_0.Vb1.t6 GNDA 0.024875f
C988 two_stage_opamp_dummy_magic_0.Vb1.t2 GNDA 0.032264f
C989 two_stage_opamp_dummy_magic_0.Vb1.n7 GNDA 0.033171f
C990 two_stage_opamp_dummy_magic_0.Vb1.t4 GNDA 0.024875f
C991 two_stage_opamp_dummy_magic_0.Vb1.t8 GNDA 0.032264f
C992 two_stage_opamp_dummy_magic_0.Vb1.n8 GNDA 0.033171f
C993 two_stage_opamp_dummy_magic_0.Vb1.n9 GNDA 0.024726f
C994 two_stage_opamp_dummy_magic_0.Vb1.t7 GNDA 0.024268f
C995 two_stage_opamp_dummy_magic_0.Vb1.t5 GNDA 0.024268f
C996 two_stage_opamp_dummy_magic_0.Vb1.n10 GNDA 0.052805f
C997 two_stage_opamp_dummy_magic_0.Vb1.n11 GNDA 0.1314f
C998 two_stage_opamp_dummy_magic_0.Vb1.t10 GNDA 0.024268f
C999 two_stage_opamp_dummy_magic_0.Vb1.t3 GNDA 0.024268f
C1000 two_stage_opamp_dummy_magic_0.Vb1.n12 GNDA 0.052805f
C1001 two_stage_opamp_dummy_magic_0.Vb1.n13 GNDA 0.212127f
C1002 two_stage_opamp_dummy_magic_0.Vb1.n14 GNDA 0.088809f
C1003 two_stage_opamp_dummy_magic_0.Vb1.t33 GNDA 0.75679f
C1004 two_stage_opamp_dummy_magic_0.Vb1.n15 GNDA 1.09347f
C1005 two_stage_opamp_dummy_magic_0.Vb1.n16 GNDA 0.067129f
C1006 two_stage_opamp_dummy_magic_0.Vb1.n17 GNDA 0.023662f
C1007 two_stage_opamp_dummy_magic_0.Vb1.n18 GNDA 0.023662f
C1008 two_stage_opamp_dummy_magic_0.Vb1.n19 GNDA 0.023662f
C1009 two_stage_opamp_dummy_magic_0.Vb1.n20 GNDA 0.023662f
C1010 two_stage_opamp_dummy_magic_0.Vb1.n21 GNDA 0.023662f
C1011 two_stage_opamp_dummy_magic_0.Vb1.n22 GNDA 0.023662f
C1012 two_stage_opamp_dummy_magic_0.Vb1.n23 GNDA 0.023662f
C1013 two_stage_opamp_dummy_magic_0.Vb1.n24 GNDA 0.023662f
C1014 two_stage_opamp_dummy_magic_0.Vb1.n25 GNDA 0.039897f
C1015 two_stage_opamp_dummy_magic_0.Vb1.t28 GNDA 0.024875f
C1016 two_stage_opamp_dummy_magic_0.Vb1.t18 GNDA 0.024875f
C1017 two_stage_opamp_dummy_magic_0.Vb1.t29 GNDA 0.024875f
C1018 two_stage_opamp_dummy_magic_0.Vb1.t20 GNDA 0.024875f
C1019 two_stage_opamp_dummy_magic_0.Vb1.t16 GNDA 0.024875f
C1020 two_stage_opamp_dummy_magic_0.Vb1.t19 GNDA 0.024875f
C1021 two_stage_opamp_dummy_magic_0.Vb1.t31 GNDA 0.024875f
C1022 two_stage_opamp_dummy_magic_0.Vb1.t22 GNDA 0.024875f
C1023 two_stage_opamp_dummy_magic_0.Vb1.t34 GNDA 0.024875f
C1024 two_stage_opamp_dummy_magic_0.Vb1.t24 GNDA 0.032264f
C1025 two_stage_opamp_dummy_magic_0.Vb1.n26 GNDA 0.035081f
C1026 two_stage_opamp_dummy_magic_0.Vb1.n27 GNDA 0.023662f
C1027 two_stage_opamp_dummy_magic_0.Vb1.n28 GNDA 0.023662f
C1028 two_stage_opamp_dummy_magic_0.Vb1.n29 GNDA 0.023662f
C1029 two_stage_opamp_dummy_magic_0.Vb1.n30 GNDA 0.023662f
C1030 two_stage_opamp_dummy_magic_0.Vb1.n31 GNDA 0.023662f
C1031 two_stage_opamp_dummy_magic_0.Vb1.n32 GNDA 0.023662f
C1032 two_stage_opamp_dummy_magic_0.Vb1.n33 GNDA 0.023662f
C1033 two_stage_opamp_dummy_magic_0.Vb1.n34 GNDA 0.039581f
C1034 two_stage_opamp_dummy_magic_0.Vb1.n35 GNDA 1.17864f
C1035 bgr_0.VB1_CUR_BIAS GNDA 1.28978f
C1036 bgr_0.PFET_GATE_10uA.t12 GNDA 0.030647f
C1037 bgr_0.PFET_GATE_10uA.t25 GNDA 0.030647f
C1038 bgr_0.PFET_GATE_10uA.t19 GNDA 0.030647f
C1039 bgr_0.PFET_GATE_10uA.t11 GNDA 0.045305f
C1040 bgr_0.PFET_GATE_10uA.n0 GNDA 0.056067f
C1041 bgr_0.PFET_GATE_10uA.n1 GNDA 0.040077f
C1042 bgr_0.PFET_GATE_10uA.n2 GNDA 0.076523f
C1043 bgr_0.PFET_GATE_10uA.t22 GNDA 0.030647f
C1044 bgr_0.PFET_GATE_10uA.t16 GNDA 0.030647f
C1045 bgr_0.PFET_GATE_10uA.t28 GNDA 0.030647f
C1046 bgr_0.PFET_GATE_10uA.t21 GNDA 0.030647f
C1047 bgr_0.PFET_GATE_10uA.t15 GNDA 0.030647f
C1048 bgr_0.PFET_GATE_10uA.t27 GNDA 0.045305f
C1049 bgr_0.PFET_GATE_10uA.n3 GNDA 0.056067f
C1050 bgr_0.PFET_GATE_10uA.n4 GNDA 0.040077f
C1051 bgr_0.PFET_GATE_10uA.n5 GNDA 0.040077f
C1052 bgr_0.PFET_GATE_10uA.n6 GNDA 0.040077f
C1053 bgr_0.PFET_GATE_10uA.t26 GNDA 0.030647f
C1054 bgr_0.PFET_GATE_10uA.t14 GNDA 0.030647f
C1055 bgr_0.PFET_GATE_10uA.t13 GNDA 0.030647f
C1056 bgr_0.PFET_GATE_10uA.t20 GNDA 0.045305f
C1057 bgr_0.PFET_GATE_10uA.n7 GNDA 0.056067f
C1058 bgr_0.PFET_GATE_10uA.n8 GNDA 0.040077f
C1059 bgr_0.PFET_GATE_10uA.n9 GNDA 0.040077f
C1060 bgr_0.PFET_GATE_10uA.n10 GNDA 0.082242f
C1061 bgr_0.PFET_GATE_10uA.n11 GNDA 0.936677f
C1062 bgr_0.PFET_GATE_10uA.t23 GNDA 0.030647f
C1063 bgr_0.PFET_GATE_10uA.t29 GNDA 0.030647f
C1064 bgr_0.PFET_GATE_10uA.t17 GNDA 0.030647f
C1065 bgr_0.PFET_GATE_10uA.t24 GNDA 0.045305f
C1066 bgr_0.PFET_GATE_10uA.n12 GNDA 0.056067f
C1067 bgr_0.PFET_GATE_10uA.n13 GNDA 0.040077f
C1068 bgr_0.PFET_GATE_10uA.n14 GNDA 0.072812f
C1069 bgr_0.PFET_GATE_10uA.n15 GNDA 0.498452f
C1070 bgr_0.PFET_GATE_10uA.t4 GNDA 0.031433f
C1071 bgr_0.PFET_GATE_10uA.t6 GNDA 0.031433f
C1072 bgr_0.PFET_GATE_10uA.n16 GNDA 0.064194f
C1073 bgr_0.PFET_GATE_10uA.n17 GNDA 0.301383f
C1074 bgr_0.PFET_GATE_10uA.n18 GNDA 0.265107f
C1075 bgr_0.PFET_GATE_10uA.t3 GNDA 0.460977f
C1076 bgr_0.PFET_GATE_10uA.n19 GNDA 1.17461f
C1077 bgr_0.PFET_GATE_10uA.t2 GNDA 0.031433f
C1078 bgr_0.PFET_GATE_10uA.t9 GNDA 0.031433f
C1079 bgr_0.PFET_GATE_10uA.n20 GNDA 0.064194f
C1080 bgr_0.PFET_GATE_10uA.n21 GNDA 0.444219f
C1081 bgr_0.PFET_GATE_10uA.t5 GNDA 0.031433f
C1082 bgr_0.PFET_GATE_10uA.t7 GNDA 0.031433f
C1083 bgr_0.PFET_GATE_10uA.n22 GNDA 0.064194f
C1084 bgr_0.PFET_GATE_10uA.n23 GNDA 0.396438f
C1085 bgr_0.PFET_GATE_10uA.n24 GNDA 0.374153f
C1086 bgr_0.PFET_GATE_10uA.n25 GNDA 0.374153f
C1087 bgr_0.PFET_GATE_10uA.t8 GNDA 0.031433f
C1088 bgr_0.PFET_GATE_10uA.t1 GNDA 0.031433f
C1089 bgr_0.PFET_GATE_10uA.n26 GNDA 0.064194f
C1090 bgr_0.PFET_GATE_10uA.n27 GNDA 0.492302f
C1091 bgr_0.PFET_GATE_10uA.n28 GNDA 0.367902f
C1092 bgr_0.PFET_GATE_10uA.n29 GNDA 0.129129f
C1093 bgr_0.PFET_GATE_10uA.t0 GNDA 0.687037f
C1094 bgr_0.PFET_GATE_10uA.t18 GNDA 0.035571f
C1095 bgr_0.PFET_GATE_10uA.t10 GNDA 0.035571f
C1096 bgr_0.PFET_GATE_10uA.n30 GNDA 0.095516f
C1097 bgr_0.PFET_GATE_10uA.n31 GNDA 2.90812f
C1098 bgr_0.PFET_GATE_10uA.n32 GNDA 0.346215f
C1099 bgr_0.PFET_GATE_10uA.n33 GNDA 0.308982f
C1100 bgr_0.V_mir2.t8 GNDA 0.031034f
C1101 bgr_0.V_mir2.t7 GNDA 0.037241f
C1102 bgr_0.V_mir2.t18 GNDA 0.037241f
C1103 bgr_0.V_mir2.t21 GNDA 0.060113f
C1104 bgr_0.V_mir2.n0 GNDA 0.067129f
C1105 bgr_0.V_mir2.n1 GNDA 0.045857f
C1106 bgr_0.V_mir2.t15 GNDA 0.047277f
C1107 bgr_0.V_mir2.n2 GNDA 0.074211f
C1108 bgr_0.V_mir2.n3 GNDA 0.166486f
C1109 bgr_0.V_mir2.t6 GNDA 0.031034f
C1110 bgr_0.V_mir2.t12 GNDA 0.031034f
C1111 bgr_0.V_mir2.n4 GNDA 0.06338f
C1112 bgr_0.V_mir2.n5 GNDA 0.260312f
C1113 bgr_0.V_mir2.t2 GNDA 0.015517f
C1114 bgr_0.V_mir2.t0 GNDA 0.015517f
C1115 bgr_0.V_mir2.n6 GNDA 0.032817f
C1116 bgr_0.V_mir2.n7 GNDA 0.172902f
C1117 bgr_0.V_mir2.t1 GNDA 0.054276f
C1118 bgr_0.V_mir2.n8 GNDA 0.277215f
C1119 bgr_0.V_mir2.n9 GNDA 0.351139f
C1120 bgr_0.V_mir2.t3 GNDA 0.015517f
C1121 bgr_0.V_mir2.t4 GNDA 0.015517f
C1122 bgr_0.V_mir2.n10 GNDA 0.032817f
C1123 bgr_0.V_mir2.n11 GNDA 0.21593f
C1124 bgr_0.V_mir2.n12 GNDA 0.356077f
C1125 bgr_0.V_mir2.n13 GNDA 0.181138f
C1126 bgr_0.V_mir2.t9 GNDA 0.037241f
C1127 bgr_0.V_mir2.t20 GNDA 0.037241f
C1128 bgr_0.V_mir2.t22 GNDA 0.060113f
C1129 bgr_0.V_mir2.n14 GNDA 0.067129f
C1130 bgr_0.V_mir2.n15 GNDA 0.045857f
C1131 bgr_0.V_mir2.t13 GNDA 0.047277f
C1132 bgr_0.V_mir2.n16 GNDA 0.074211f
C1133 bgr_0.V_mir2.t5 GNDA 0.037241f
C1134 bgr_0.V_mir2.t19 GNDA 0.037241f
C1135 bgr_0.V_mir2.t17 GNDA 0.060113f
C1136 bgr_0.V_mir2.n17 GNDA 0.067129f
C1137 bgr_0.V_mir2.n18 GNDA 0.045857f
C1138 bgr_0.V_mir2.t11 GNDA 0.047277f
C1139 bgr_0.V_mir2.n19 GNDA 0.074211f
C1140 bgr_0.V_mir2.n20 GNDA 0.166486f
C1141 bgr_0.V_mir2.n21 GNDA 0.450644f
C1142 bgr_0.V_mir2.n22 GNDA 0.199395f
C1143 bgr_0.V_mir2.t10 GNDA 0.031034f
C1144 bgr_0.V_mir2.t14 GNDA 0.031034f
C1145 bgr_0.V_mir2.n23 GNDA 0.06338f
C1146 bgr_0.V_mir2.n24 GNDA 0.213276f
C1147 bgr_0.V_mir2.n25 GNDA 0.463152f
C1148 bgr_0.V_mir2.n26 GNDA 0.260312f
C1149 bgr_0.V_mir2.n27 GNDA 0.06338f
C1150 bgr_0.V_mir2.t16 GNDA 0.031034f
C1151 bgr_0.V_p_2.n0 GNDA 0.684513f
C1152 bgr_0.V_p_2.n1 GNDA 0.256175f
C1153 bgr_0.V_p_2.n2 GNDA 0.18041f
C1154 bgr_0.V_p_2.n3 GNDA 0.185403f
C1155 bgr_0.V_p_2.n4 GNDA 0.017531f
C1156 bgr_0.V_p_2.n5 GNDA 0.017531f
C1157 bgr_0.V_p_2.n6 GNDA 0.175416f
C1158 bgr_0.V_p_2.n7 GNDA 0.017531f
C1159 bgr_0.V_p_2.t8 GNDA 0.196701f
C1160 bgr_0.V_p_2.n8 GNDA 0.017531f
C1161 bgr_0.V_p_2.n9 GNDA 0.175416f
C1162 bgr_0.V_p_2.n10 GNDA 0.175416f
C1163 bgr_0.V_p_2.n11 GNDA 0.017531f
C1164 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 GNDA 0.021934f
C1165 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 GNDA 0.021934f
C1166 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 GNDA 0.021934f
C1167 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 GNDA 0.021934f
C1168 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 GNDA 0.021934f
C1169 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 GNDA 0.021934f
C1170 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 GNDA 0.021934f
C1171 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 GNDA 0.021934f
C1172 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 GNDA 0.021934f
C1173 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 GNDA 0.067288f
C1174 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 GNDA 0.091409f
C1175 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 GNDA 0.073542f
C1176 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 GNDA 0.073542f
C1177 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 GNDA 0.433083f
C1178 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 GNDA 0.433083f
C1179 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 GNDA 0.073542f
C1180 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 GNDA 0.073542f
C1181 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 GNDA 0.073542f
C1182 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 GNDA 0.109382f
C1183 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 GNDA 0.526865f
C1184 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 GNDA 0.085109f
C1185 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 GNDA 0.031825f
C1186 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 GNDA 0.099822f
C1187 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 GNDA 0.031825f
C1188 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 GNDA 0.081714f
C1189 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 GNDA 0.031825f
C1190 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 GNDA 0.081714f
C1191 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 GNDA 0.031825f
C1192 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 GNDA 0.102647f
C1193 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 GNDA 2.74879f
C1194 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 GNDA 0.757364f
C1195 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 GNDA 0.103217f
C1196 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 GNDA 0.103217f
C1197 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 GNDA 0.211119f
C1198 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 GNDA 1.13907f
C1199 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 GNDA 0.103217f
C1200 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 GNDA 0.103217f
C1201 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 GNDA 0.211119f
C1202 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 GNDA 0.854779f
C1203 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 GNDA 0.899716f
C1204 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 GNDA 0.103217f
C1205 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 GNDA 0.103217f
C1206 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n20 GNDA 0.211119f
C1207 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n21 GNDA 0.995574f
C1208 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n22 GNDA 0.789261f
C1209 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n23 GNDA 2.41641f
C1210 two_stage_opamp_dummy_magic_0.VD4.t5 GNDA 0.067965f
C1211 two_stage_opamp_dummy_magic_0.VD4.n0 GNDA 0.122886f
C1212 two_stage_opamp_dummy_magic_0.VD4.n1 GNDA 0.07372f
C1213 two_stage_opamp_dummy_magic_0.VD4.n2 GNDA 0.07372f
C1214 two_stage_opamp_dummy_magic_0.VD4.n3 GNDA 0.07372f
C1215 two_stage_opamp_dummy_magic_0.VD4.t37 GNDA 0.067965f
C1216 two_stage_opamp_dummy_magic_0.VD4.t23 GNDA 0.067965f
C1217 two_stage_opamp_dummy_magic_0.VD4.n4 GNDA 0.139029f
C1218 two_stage_opamp_dummy_magic_0.VD4.n5 GNDA 0.450134f
C1219 two_stage_opamp_dummy_magic_0.VD4.n6 GNDA 0.125758f
C1220 two_stage_opamp_dummy_magic_0.VD4.t1 GNDA 0.067965f
C1221 two_stage_opamp_dummy_magic_0.VD4.t31 GNDA 0.067965f
C1222 two_stage_opamp_dummy_magic_0.VD4.n7 GNDA 0.139029f
C1223 two_stage_opamp_dummy_magic_0.VD4.n8 GNDA 0.437842f
C1224 two_stage_opamp_dummy_magic_0.VD4.n9 GNDA 0.125758f
C1225 two_stage_opamp_dummy_magic_0.VD4.t0 GNDA 0.067965f
C1226 two_stage_opamp_dummy_magic_0.VD4.t35 GNDA 0.067965f
C1227 two_stage_opamp_dummy_magic_0.VD4.n10 GNDA 0.139029f
C1228 two_stage_opamp_dummy_magic_0.VD4.n11 GNDA 0.437842f
C1229 two_stage_opamp_dummy_magic_0.VD4.n12 GNDA 0.07372f
C1230 two_stage_opamp_dummy_magic_0.VD4.n13 GNDA 0.07372f
C1231 two_stage_opamp_dummy_magic_0.VD4.t32 GNDA 0.067965f
C1232 two_stage_opamp_dummy_magic_0.VD4.t34 GNDA 0.067965f
C1233 two_stage_opamp_dummy_magic_0.VD4.n14 GNDA 0.139029f
C1234 two_stage_opamp_dummy_magic_0.VD4.n15 GNDA 0.437842f
C1235 two_stage_opamp_dummy_magic_0.VD4.n16 GNDA 0.07372f
C1236 two_stage_opamp_dummy_magic_0.VD4.t33 GNDA 0.067965f
C1237 two_stage_opamp_dummy_magic_0.VD4.t30 GNDA 0.067965f
C1238 two_stage_opamp_dummy_magic_0.VD4.n17 GNDA 0.139029f
C1239 two_stage_opamp_dummy_magic_0.VD4.n18 GNDA 0.437842f
C1240 two_stage_opamp_dummy_magic_0.VD4.n19 GNDA 0.125758f
C1241 two_stage_opamp_dummy_magic_0.VD4.t22 GNDA 0.067965f
C1242 two_stage_opamp_dummy_magic_0.VD4.t36 GNDA 0.067965f
C1243 two_stage_opamp_dummy_magic_0.VD4.n20 GNDA 0.139029f
C1244 two_stage_opamp_dummy_magic_0.VD4.n21 GNDA 0.443988f
C1245 two_stage_opamp_dummy_magic_0.VD4.n22 GNDA 0.131975f
C1246 two_stage_opamp_dummy_magic_0.VD4.t24 GNDA 0.118986f
C1247 two_stage_opamp_dummy_magic_0.VD4.n23 GNDA 0.184816f
C1248 two_stage_opamp_dummy_magic_0.VD4.t26 GNDA 0.24176f
C1249 two_stage_opamp_dummy_magic_0.VD4.t29 GNDA 0.24176f
C1250 two_stage_opamp_dummy_magic_0.VD4.t27 GNDA 0.118986f
C1251 two_stage_opamp_dummy_magic_0.VD4.n24 GNDA 0.184816f
C1252 two_stage_opamp_dummy_magic_0.VD4.n25 GNDA 0.07372f
C1253 two_stage_opamp_dummy_magic_0.VD4.t13 GNDA 0.067965f
C1254 two_stage_opamp_dummy_magic_0.VD4.t17 GNDA 0.067965f
C1255 two_stage_opamp_dummy_magic_0.VD4.n26 GNDA 0.139029f
C1256 two_stage_opamp_dummy_magic_0.VD4.n27 GNDA 0.468873f
C1257 two_stage_opamp_dummy_magic_0.VD4.n28 GNDA 0.080554f
C1258 two_stage_opamp_dummy_magic_0.VD4.n29 GNDA 0.07372f
C1259 two_stage_opamp_dummy_magic_0.VD4.t7 GNDA 0.067965f
C1260 two_stage_opamp_dummy_magic_0.VD4.t9 GNDA 0.067965f
C1261 two_stage_opamp_dummy_magic_0.VD4.n30 GNDA 0.139029f
C1262 two_stage_opamp_dummy_magic_0.VD4.n31 GNDA 0.468873f
C1263 two_stage_opamp_dummy_magic_0.VD4.n32 GNDA 0.080554f
C1264 two_stage_opamp_dummy_magic_0.VD4.t19 GNDA 0.067965f
C1265 two_stage_opamp_dummy_magic_0.VD4.t3 GNDA 0.067965f
C1266 two_stage_opamp_dummy_magic_0.VD4.n33 GNDA 0.139029f
C1267 two_stage_opamp_dummy_magic_0.VD4.n34 GNDA 0.468873f
C1268 two_stage_opamp_dummy_magic_0.VD4.n35 GNDA 0.080554f
C1269 two_stage_opamp_dummy_magic_0.VD4.n36 GNDA 0.122886f
C1270 two_stage_opamp_dummy_magic_0.VD4.t11 GNDA 0.067965f
C1271 two_stage_opamp_dummy_magic_0.VD4.t15 GNDA 0.067965f
C1272 two_stage_opamp_dummy_magic_0.VD4.n37 GNDA 0.139029f
C1273 two_stage_opamp_dummy_magic_0.VD4.n38 GNDA 0.468873f
C1274 two_stage_opamp_dummy_magic_0.VD4.n39 GNDA 0.125758f
C1275 two_stage_opamp_dummy_magic_0.VD4.n40 GNDA 0.188751f
C1276 two_stage_opamp_dummy_magic_0.VD4.n41 GNDA 0.701325f
C1277 two_stage_opamp_dummy_magic_0.VD4.t28 GNDA 0.579325f
C1278 two_stage_opamp_dummy_magic_0.VD4.t10 GNDA 0.454393f
C1279 two_stage_opamp_dummy_magic_0.VD4.t14 GNDA 0.454393f
C1280 two_stage_opamp_dummy_magic_0.VD4.t18 GNDA 0.454393f
C1281 two_stage_opamp_dummy_magic_0.VD4.t2 GNDA 0.454393f
C1282 two_stage_opamp_dummy_magic_0.VD4.t6 GNDA 0.454393f
C1283 two_stage_opamp_dummy_magic_0.VD4.t8 GNDA 0.454393f
C1284 two_stage_opamp_dummy_magic_0.VD4.t12 GNDA 0.454393f
C1285 two_stage_opamp_dummy_magic_0.VD4.t16 GNDA 0.454393f
C1286 two_stage_opamp_dummy_magic_0.VD4.t20 GNDA 0.454393f
C1287 two_stage_opamp_dummy_magic_0.VD4.t4 GNDA 0.454393f
C1288 two_stage_opamp_dummy_magic_0.VD4.t25 GNDA 0.579325f
C1289 two_stage_opamp_dummy_magic_0.VD4.n42 GNDA 0.701325f
C1290 two_stage_opamp_dummy_magic_0.VD4.n43 GNDA 0.182605f
C1291 two_stage_opamp_dummy_magic_0.VD4.n44 GNDA 0.131975f
C1292 two_stage_opamp_dummy_magic_0.VD4.n45 GNDA 0.07372f
C1293 two_stage_opamp_dummy_magic_0.VD4.n46 GNDA 0.468873f
C1294 two_stage_opamp_dummy_magic_0.VD4.n47 GNDA 0.139029f
C1295 two_stage_opamp_dummy_magic_0.VD4.t21 GNDA 0.067965f
C1296 two_stage_opamp_dummy_magic_0.Vb2.n0 GNDA 0.023174f
C1297 two_stage_opamp_dummy_magic_0.Vb2.n1 GNDA 0.022113f
C1298 two_stage_opamp_dummy_magic_0.Vb2.n2 GNDA 0.397356f
C1299 two_stage_opamp_dummy_magic_0.Vb2.n3 GNDA 0.14203f
C1300 two_stage_opamp_dummy_magic_0.Vb2.t2 GNDA 0.030326f
C1301 two_stage_opamp_dummy_magic_0.Vb2.t0 GNDA 0.030326f
C1302 two_stage_opamp_dummy_magic_0.Vb2.n4 GNDA 0.0644f
C1303 two_stage_opamp_dummy_magic_0.Vb2.t1 GNDA 0.056611f
C1304 two_stage_opamp_dummy_magic_0.Vb2.n5 GNDA 0.262142f
C1305 two_stage_opamp_dummy_magic_0.Vb2.t13 GNDA 0.033997f
C1306 two_stage_opamp_dummy_magic_0.Vb2.n6 GNDA 0.130516f
C1307 two_stage_opamp_dummy_magic_0.Vb2.t31 GNDA 0.04289f
C1308 two_stage_opamp_dummy_magic_0.Vb2.t25 GNDA 0.04289f
C1309 two_stage_opamp_dummy_magic_0.Vb2.t28 GNDA 0.04289f
C1310 two_stage_opamp_dummy_magic_0.Vb2.t22 GNDA 0.049495f
C1311 two_stage_opamp_dummy_magic_0.Vb2.n7 GNDA 0.040184f
C1312 two_stage_opamp_dummy_magic_0.Vb2.n8 GNDA 0.024694f
C1313 two_stage_opamp_dummy_magic_0.Vb2.n9 GNDA 0.024214f
C1314 two_stage_opamp_dummy_magic_0.Vb2.t20 GNDA 0.04289f
C1315 two_stage_opamp_dummy_magic_0.Vb2.t23 GNDA 0.04289f
C1316 two_stage_opamp_dummy_magic_0.Vb2.t21 GNDA 0.04289f
C1317 two_stage_opamp_dummy_magic_0.Vb2.t26 GNDA 0.04289f
C1318 two_stage_opamp_dummy_magic_0.Vb2.t32 GNDA 0.049495f
C1319 two_stage_opamp_dummy_magic_0.Vb2.n10 GNDA 0.040184f
C1320 two_stage_opamp_dummy_magic_0.Vb2.n11 GNDA 0.024694f
C1321 two_stage_opamp_dummy_magic_0.Vb2.n12 GNDA 0.024694f
C1322 two_stage_opamp_dummy_magic_0.Vb2.n13 GNDA 0.024214f
C1323 two_stage_opamp_dummy_magic_0.Vb2.t18 GNDA 0.044406f
C1324 two_stage_opamp_dummy_magic_0.Vb2.n14 GNDA 0.041031f
C1325 two_stage_opamp_dummy_magic_0.Vb2.t19 GNDA 0.04289f
C1326 two_stage_opamp_dummy_magic_0.Vb2.t16 GNDA 0.04289f
C1327 two_stage_opamp_dummy_magic_0.Vb2.t14 GNDA 0.04289f
C1328 two_stage_opamp_dummy_magic_0.Vb2.t11 GNDA 0.04289f
C1329 two_stage_opamp_dummy_magic_0.Vb2.t29 GNDA 0.049495f
C1330 two_stage_opamp_dummy_magic_0.Vb2.n15 GNDA 0.040184f
C1331 two_stage_opamp_dummy_magic_0.Vb2.n16 GNDA 0.024694f
C1332 two_stage_opamp_dummy_magic_0.Vb2.n17 GNDA 0.024694f
C1333 two_stage_opamp_dummy_magic_0.Vb2.n18 GNDA 0.024214f
C1334 two_stage_opamp_dummy_magic_0.Vb2.t30 GNDA 0.04289f
C1335 two_stage_opamp_dummy_magic_0.Vb2.t12 GNDA 0.04289f
C1336 two_stage_opamp_dummy_magic_0.Vb2.t15 GNDA 0.04289f
C1337 two_stage_opamp_dummy_magic_0.Vb2.t17 GNDA 0.049495f
C1338 two_stage_opamp_dummy_magic_0.Vb2.n19 GNDA 0.040184f
C1339 two_stage_opamp_dummy_magic_0.Vb2.n20 GNDA 0.024694f
C1340 two_stage_opamp_dummy_magic_0.Vb2.n21 GNDA 0.024214f
C1341 two_stage_opamp_dummy_magic_0.Vb2.t24 GNDA 0.044406f
C1342 two_stage_opamp_dummy_magic_0.Vb2.n22 GNDA 0.040843f
C1343 two_stage_opamp_dummy_magic_0.Vb2.n23 GNDA 0.344613f
C1344 two_stage_opamp_dummy_magic_0.Vb2.n24 GNDA 0.16247f
C1345 two_stage_opamp_dummy_magic_0.Vb2.t27 GNDA 0.055738f
C1346 two_stage_opamp_dummy_magic_0.Vb2.n25 GNDA 0.733611f
C1347 two_stage_opamp_dummy_magic_0.Vb2.n26 GNDA 0.743682f
C1348 two_stage_opamp_dummy_magic_0.Vb2.n27 GNDA 0.018449f
C1349 two_stage_opamp_dummy_magic_0.Vb2.n28 GNDA 0.142901f
C1350 two_stage_opamp_dummy_magic_0.Vb2.n29 GNDA 0.142901f
C1351 two_stage_opamp_dummy_magic_0.Vb2.n30 GNDA 0.018449f
C1352 bgr_0.NFET_GATE_10uA.t3 GNDA 0.015735f
C1353 bgr_0.NFET_GATE_10uA.t2 GNDA 0.015735f
C1354 bgr_0.NFET_GATE_10uA.n0 GNDA 0.033951f
C1355 bgr_0.NFET_GATE_10uA.t22 GNDA 0.015931f
C1356 bgr_0.NFET_GATE_10uA.t10 GNDA 0.015931f
C1357 bgr_0.NFET_GATE_10uA.t16 GNDA 0.015931f
C1358 bgr_0.NFET_GATE_10uA.t23 GNDA 0.015931f
C1359 bgr_0.NFET_GATE_10uA.t6 GNDA 0.015931f
C1360 bgr_0.NFET_GATE_10uA.t14 GNDA 0.015931f
C1361 bgr_0.NFET_GATE_10uA.t13 GNDA 0.023233f
C1362 bgr_0.NFET_GATE_10uA.n1 GNDA 0.029281f
C1363 bgr_0.NFET_GATE_10uA.n2 GNDA 0.020652f
C1364 bgr_0.NFET_GATE_10uA.n3 GNDA 0.016226f
C1365 bgr_0.NFET_GATE_10uA.t7 GNDA 0.015341f
C1366 bgr_0.NFET_GATE_10uA.t9 GNDA 0.015341f
C1367 bgr_0.NFET_GATE_10uA.t21 GNDA 0.015341f
C1368 bgr_0.NFET_GATE_10uA.t15 GNDA 0.015341f
C1369 bgr_0.NFET_GATE_10uA.t8 GNDA 0.015341f
C1370 bgr_0.NFET_GATE_10uA.t20 GNDA 0.022678f
C1371 bgr_0.NFET_GATE_10uA.n4 GNDA 0.028066f
C1372 bgr_0.NFET_GATE_10uA.n5 GNDA 0.020062f
C1373 bgr_0.NFET_GATE_10uA.n6 GNDA 0.020062f
C1374 bgr_0.NFET_GATE_10uA.n7 GNDA 0.020062f
C1375 bgr_0.NFET_GATE_10uA.n8 GNDA 0.038642f
C1376 bgr_0.NFET_GATE_10uA.t11 GNDA 0.015341f
C1377 bgr_0.NFET_GATE_10uA.t18 GNDA 0.015341f
C1378 bgr_0.NFET_GATE_10uA.t5 GNDA 0.015341f
C1379 bgr_0.NFET_GATE_10uA.t12 GNDA 0.015341f
C1380 bgr_0.NFET_GATE_10uA.t19 GNDA 0.015341f
C1381 bgr_0.NFET_GATE_10uA.t17 GNDA 0.022678f
C1382 bgr_0.NFET_GATE_10uA.n9 GNDA 0.028066f
C1383 bgr_0.NFET_GATE_10uA.n10 GNDA 0.020062f
C1384 bgr_0.NFET_GATE_10uA.n11 GNDA 0.020062f
C1385 bgr_0.NFET_GATE_10uA.n12 GNDA 0.020062f
C1386 bgr_0.NFET_GATE_10uA.n13 GNDA 0.038671f
C1387 bgr_0.NFET_GATE_10uA.n14 GNDA 0.520479f
C1388 bgr_0.NFET_GATE_10uA.n15 GNDA 0.03651f
C1389 bgr_0.NFET_GATE_10uA.n16 GNDA 0.016226f
C1390 bgr_0.NFET_GATE_10uA.n17 GNDA 0.020652f
C1391 bgr_0.NFET_GATE_10uA.n18 GNDA 0.029281f
C1392 bgr_0.NFET_GATE_10uA.t1 GNDA 0.038233f
C1393 bgr_0.NFET_GATE_10uA.n19 GNDA 0.491201f
C1394 bgr_0.NFET_GATE_10uA.t0 GNDA 0.015735f
C1395 bgr_0.NFET_GATE_10uA.t4 GNDA 0.015735f
C1396 bgr_0.NFET_GATE_10uA.n20 GNDA 0.10107f
C1397 two_stage_opamp_dummy_magic_0.V_source.t13 GNDA 0.038168f
C1398 two_stage_opamp_dummy_magic_0.V_source.t0 GNDA 0.022901f
C1399 two_stage_opamp_dummy_magic_0.V_source.t3 GNDA 0.022901f
C1400 two_stage_opamp_dummy_magic_0.V_source.n0 GNDA 0.049829f
C1401 two_stage_opamp_dummy_magic_0.V_source.n1 GNDA 0.153174f
C1402 two_stage_opamp_dummy_magic_0.V_source.n2 GNDA 0.051155f
C1403 two_stage_opamp_dummy_magic_0.V_source.t31 GNDA 0.022901f
C1404 two_stage_opamp_dummy_magic_0.V_source.t38 GNDA 0.022901f
C1405 two_stage_opamp_dummy_magic_0.V_source.n3 GNDA 0.049829f
C1406 two_stage_opamp_dummy_magic_0.V_source.n4 GNDA 0.200044f
C1407 two_stage_opamp_dummy_magic_0.V_source.n5 GNDA 0.087575f
C1408 two_stage_opamp_dummy_magic_0.V_source.t6 GNDA 0.022901f
C1409 two_stage_opamp_dummy_magic_0.V_source.t5 GNDA 0.022901f
C1410 two_stage_opamp_dummy_magic_0.V_source.n6 GNDA 0.049829f
C1411 two_stage_opamp_dummy_magic_0.V_source.n7 GNDA 0.192055f
C1412 two_stage_opamp_dummy_magic_0.V_source.n8 GNDA 0.083262f
C1413 two_stage_opamp_dummy_magic_0.V_source.t33 GNDA 0.022901f
C1414 two_stage_opamp_dummy_magic_0.V_source.t30 GNDA 0.022901f
C1415 two_stage_opamp_dummy_magic_0.V_source.n9 GNDA 0.049829f
C1416 two_stage_opamp_dummy_magic_0.V_source.n10 GNDA 0.192055f
C1417 two_stage_opamp_dummy_magic_0.V_source.n11 GNDA 0.048946f
C1418 two_stage_opamp_dummy_magic_0.V_source.n12 GNDA 0.083262f
C1419 two_stage_opamp_dummy_magic_0.V_source.t25 GNDA 0.022901f
C1420 two_stage_opamp_dummy_magic_0.V_source.t39 GNDA 0.022901f
C1421 two_stage_opamp_dummy_magic_0.V_source.n13 GNDA 0.049829f
C1422 two_stage_opamp_dummy_magic_0.V_source.n14 GNDA 0.192055f
C1423 two_stage_opamp_dummy_magic_0.V_source.n15 GNDA 0.051155f
C1424 two_stage_opamp_dummy_magic_0.V_source.n16 GNDA 0.051155f
C1425 two_stage_opamp_dummy_magic_0.V_source.n17 GNDA 0.083262f
C1426 two_stage_opamp_dummy_magic_0.V_source.t32 GNDA 0.022901f
C1427 two_stage_opamp_dummy_magic_0.V_source.t37 GNDA 0.022901f
C1428 two_stage_opamp_dummy_magic_0.V_source.n18 GNDA 0.049829f
C1429 two_stage_opamp_dummy_magic_0.V_source.n19 GNDA 0.200044f
C1430 two_stage_opamp_dummy_magic_0.V_source.t1 GNDA 0.022901f
C1431 two_stage_opamp_dummy_magic_0.V_source.t28 GNDA 0.022901f
C1432 two_stage_opamp_dummy_magic_0.V_source.n20 GNDA 0.049829f
C1433 two_stage_opamp_dummy_magic_0.V_source.n21 GNDA 0.192055f
C1434 two_stage_opamp_dummy_magic_0.V_source.n22 GNDA 0.087575f
C1435 two_stage_opamp_dummy_magic_0.V_source.n23 GNDA 0.051155f
C1436 two_stage_opamp_dummy_magic_0.V_source.t26 GNDA 0.022901f
C1437 two_stage_opamp_dummy_magic_0.V_source.t2 GNDA 0.022901f
C1438 two_stage_opamp_dummy_magic_0.V_source.n24 GNDA 0.049829f
C1439 two_stage_opamp_dummy_magic_0.V_source.n25 GNDA 0.192055f
C1440 two_stage_opamp_dummy_magic_0.V_source.n26 GNDA 0.048946f
C1441 two_stage_opamp_dummy_magic_0.V_source.t40 GNDA 0.022901f
C1442 two_stage_opamp_dummy_magic_0.V_source.t36 GNDA 0.022901f
C1443 two_stage_opamp_dummy_magic_0.V_source.n27 GNDA 0.049829f
C1444 two_stage_opamp_dummy_magic_0.V_source.n28 GNDA 0.192055f
C1445 two_stage_opamp_dummy_magic_0.V_source.n29 GNDA 0.083262f
C1446 two_stage_opamp_dummy_magic_0.V_source.t35 GNDA 0.022901f
C1447 two_stage_opamp_dummy_magic_0.V_source.t4 GNDA 0.022901f
C1448 two_stage_opamp_dummy_magic_0.V_source.n30 GNDA 0.049829f
C1449 two_stage_opamp_dummy_magic_0.V_source.n31 GNDA 0.195998f
C1450 two_stage_opamp_dummy_magic_0.V_source.n32 GNDA 0.125964f
C1451 two_stage_opamp_dummy_magic_0.V_source.n33 GNDA 0.120611f
C1452 two_stage_opamp_dummy_magic_0.V_source.n34 GNDA 0.087586f
C1453 two_stage_opamp_dummy_magic_0.V_source.n35 GNDA 0.099442f
C1454 two_stage_opamp_dummy_magic_0.V_source.t29 GNDA 0.079851f
C1455 two_stage_opamp_dummy_magic_0.V_source.n36 GNDA 0.096361f
C1456 two_stage_opamp_dummy_magic_0.V_source.n37 GNDA 0.05567f
C1457 two_stage_opamp_dummy_magic_0.V_source.t34 GNDA 0.038168f
C1458 two_stage_opamp_dummy_magic_0.V_source.t27 GNDA 0.038168f
C1459 two_stage_opamp_dummy_magic_0.V_source.n38 GNDA 0.081597f
C1460 two_stage_opamp_dummy_magic_0.V_source.n39 GNDA 0.294282f
C1461 two_stage_opamp_dummy_magic_0.V_source.t23 GNDA 0.038168f
C1462 two_stage_opamp_dummy_magic_0.V_source.t17 GNDA 0.038168f
C1463 two_stage_opamp_dummy_magic_0.V_source.n40 GNDA 0.081597f
C1464 two_stage_opamp_dummy_magic_0.V_source.n41 GNDA 0.285878f
C1465 two_stage_opamp_dummy_magic_0.V_source.n42 GNDA 0.090055f
C1466 two_stage_opamp_dummy_magic_0.V_source.n43 GNDA 0.045802f
C1467 two_stage_opamp_dummy_magic_0.V_source.n44 GNDA 0.052428f
C1468 two_stage_opamp_dummy_magic_0.V_source.n45 GNDA 0.096361f
C1469 two_stage_opamp_dummy_magic_0.V_source.t10 GNDA 0.038168f
C1470 two_stage_opamp_dummy_magic_0.V_source.t16 GNDA 0.038168f
C1471 two_stage_opamp_dummy_magic_0.V_source.n46 GNDA 0.081597f
C1472 two_stage_opamp_dummy_magic_0.V_source.n47 GNDA 0.294282f
C1473 two_stage_opamp_dummy_magic_0.V_source.t12 GNDA 0.038168f
C1474 two_stage_opamp_dummy_magic_0.V_source.t20 GNDA 0.038168f
C1475 two_stage_opamp_dummy_magic_0.V_source.n48 GNDA 0.081597f
C1476 two_stage_opamp_dummy_magic_0.V_source.n49 GNDA 0.285878f
C1477 two_stage_opamp_dummy_magic_0.V_source.n50 GNDA 0.090055f
C1478 two_stage_opamp_dummy_magic_0.V_source.n51 GNDA 0.052428f
C1479 two_stage_opamp_dummy_magic_0.V_source.t14 GNDA 0.038168f
C1480 two_stage_opamp_dummy_magic_0.V_source.t22 GNDA 0.038168f
C1481 two_stage_opamp_dummy_magic_0.V_source.n52 GNDA 0.081597f
C1482 two_stage_opamp_dummy_magic_0.V_source.n53 GNDA 0.285878f
C1483 two_stage_opamp_dummy_magic_0.V_source.n54 GNDA 0.05567f
C1484 two_stage_opamp_dummy_magic_0.V_source.t18 GNDA 0.038168f
C1485 two_stage_opamp_dummy_magic_0.V_source.t8 GNDA 0.038168f
C1486 two_stage_opamp_dummy_magic_0.V_source.n55 GNDA 0.081597f
C1487 two_stage_opamp_dummy_magic_0.V_source.n56 GNDA 0.285878f
C1488 two_stage_opamp_dummy_magic_0.V_source.n57 GNDA 0.05567f
C1489 two_stage_opamp_dummy_magic_0.V_source.n58 GNDA 0.05567f
C1490 two_stage_opamp_dummy_magic_0.V_source.t15 GNDA 0.038168f
C1491 two_stage_opamp_dummy_magic_0.V_source.t7 GNDA 0.038168f
C1492 two_stage_opamp_dummy_magic_0.V_source.n59 GNDA 0.081597f
C1493 two_stage_opamp_dummy_magic_0.V_source.n60 GNDA 0.285878f
C1494 two_stage_opamp_dummy_magic_0.V_source.n61 GNDA 0.052428f
C1495 two_stage_opamp_dummy_magic_0.V_source.t19 GNDA 0.038168f
C1496 two_stage_opamp_dummy_magic_0.V_source.t9 GNDA 0.038168f
C1497 two_stage_opamp_dummy_magic_0.V_source.n62 GNDA 0.081597f
C1498 two_stage_opamp_dummy_magic_0.V_source.n63 GNDA 0.285878f
C1499 two_stage_opamp_dummy_magic_0.V_source.n64 GNDA 0.052428f
C1500 two_stage_opamp_dummy_magic_0.V_source.n65 GNDA 0.052428f
C1501 two_stage_opamp_dummy_magic_0.V_source.t21 GNDA 0.038168f
C1502 two_stage_opamp_dummy_magic_0.V_source.t11 GNDA 0.038168f
C1503 two_stage_opamp_dummy_magic_0.V_source.n66 GNDA 0.081597f
C1504 two_stage_opamp_dummy_magic_0.V_source.n67 GNDA 0.285878f
C1505 two_stage_opamp_dummy_magic_0.V_source.n68 GNDA 0.05567f
C1506 two_stage_opamp_dummy_magic_0.V_source.n69 GNDA 0.045802f
C1507 two_stage_opamp_dummy_magic_0.V_source.n70 GNDA 0.258117f
C1508 two_stage_opamp_dummy_magic_0.V_source.n71 GNDA 0.185859f
C1509 two_stage_opamp_dummy_magic_0.V_source.n72 GNDA 0.081597f
C1510 two_stage_opamp_dummy_magic_0.V_source.t24 GNDA 0.038168f
C1511 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 GNDA 0.028313f
C1512 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 GNDA 0.028313f
C1513 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 GNDA 0.075699f
C1514 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 GNDA 0.028313f
C1515 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 GNDA 0.028313f
C1516 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 GNDA 0.072244f
C1517 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 GNDA 2.19144f
C1518 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 GNDA 0.35159f
C1519 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 GNDA 0.098481f
C1520 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 GNDA 0.169447f
C1521 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 GNDA 0.084938f
C1522 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 GNDA 0.084938f
C1523 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 GNDA 0.181667f
C1524 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 GNDA 0.568252f
C1525 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 GNDA 0.084938f
C1526 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 GNDA 0.084938f
C1527 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 GNDA 0.181667f
C1528 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 GNDA 0.552862f
C1529 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 GNDA 0.169447f
C1530 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 GNDA 0.098481f
C1531 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 GNDA 0.084938f
C1532 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 GNDA 0.084938f
C1533 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 GNDA 0.181667f
C1534 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 GNDA 0.552862f
C1535 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n13 GNDA 0.098481f
C1536 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 GNDA 0.084938f
C1537 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 GNDA 0.084938f
C1538 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n14 GNDA 0.181667f
C1539 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n15 GNDA 0.552862f
C1540 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n16 GNDA 0.169447f
C1541 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 GNDA 0.084938f
C1542 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 GNDA 0.084938f
C1543 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n17 GNDA 0.181667f
C1544 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n18 GNDA 0.560557f
C1545 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n19 GNDA 0.219581f
C1546 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n20 GNDA 2.16409f
C1547 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n21 GNDA 2.34906f
C1548 bgr_0.V_CMFB_S4 GNDA 0.014156f
C1549 bgr_0.cap_res2.t7 GNDA 0.358376f
C1550 bgr_0.cap_res2.t13 GNDA 0.359675f
C1551 bgr_0.cap_res2.t15 GNDA 0.340442f
C1552 bgr_0.cap_res2.t1 GNDA 0.358376f
C1553 bgr_0.cap_res2.t6 GNDA 0.359675f
C1554 bgr_0.cap_res2.t9 GNDA 0.340442f
C1555 bgr_0.cap_res2.t5 GNDA 0.358376f
C1556 bgr_0.cap_res2.t11 GNDA 0.359675f
C1557 bgr_0.cap_res2.t14 GNDA 0.340442f
C1558 bgr_0.cap_res2.t20 GNDA 0.358376f
C1559 bgr_0.cap_res2.t4 GNDA 0.359675f
C1560 bgr_0.cap_res2.t8 GNDA 0.340442f
C1561 bgr_0.cap_res2.t16 GNDA 0.358376f
C1562 bgr_0.cap_res2.t19 GNDA 0.359675f
C1563 bgr_0.cap_res2.t2 GNDA 0.340442f
C1564 bgr_0.cap_res2.n0 GNDA 0.24022f
C1565 bgr_0.cap_res2.t3 GNDA 0.1913f
C1566 bgr_0.cap_res2.n1 GNDA 0.260644f
C1567 bgr_0.cap_res2.t10 GNDA 0.1913f
C1568 bgr_0.cap_res2.n2 GNDA 0.260644f
C1569 bgr_0.cap_res2.t17 GNDA 0.1913f
C1570 bgr_0.cap_res2.n3 GNDA 0.260644f
C1571 bgr_0.cap_res2.t12 GNDA 0.1913f
C1572 bgr_0.cap_res2.n4 GNDA 0.260644f
C1573 bgr_0.cap_res2.t18 GNDA 0.373116f
C1574 bgr_0.cap_res2.t0 GNDA 0.086426f
C1575 bgr_0.1st_Vout_2.n0 GNDA 0.205909f
C1576 bgr_0.1st_Vout_2.n1 GNDA 0.3069f
C1577 bgr_0.1st_Vout_2.n2 GNDA 1.00621f
C1578 bgr_0.1st_Vout_2.n3 GNDA 0.178696f
C1579 bgr_0.1st_Vout_2.n4 GNDA 0.113f
C1580 bgr_0.1st_Vout_2.n5 GNDA 0.21697f
C1581 bgr_0.1st_Vout_2.n6 GNDA 2.61681f
C1582 bgr_0.1st_Vout_2.n7 GNDA 2.65427f
C1583 bgr_0.1st_Vout_2.t7 GNDA 0.013189f
C1584 bgr_0.1st_Vout_2.t28 GNDA 0.52755f
C1585 bgr_0.1st_Vout_2.t17 GNDA 0.536536f
C1586 bgr_0.1st_Vout_2.t12 GNDA 0.52755f
C1587 bgr_0.1st_Vout_2.t32 GNDA 0.52755f
C1588 bgr_0.1st_Vout_2.t35 GNDA 0.536536f
C1589 bgr_0.1st_Vout_2.t11 GNDA 0.536536f
C1590 bgr_0.1st_Vout_2.t31 GNDA 0.52755f
C1591 bgr_0.1st_Vout_2.t24 GNDA 0.52755f
C1592 bgr_0.1st_Vout_2.t27 GNDA 0.536536f
C1593 bgr_0.1st_Vout_2.t30 GNDA 0.536536f
C1594 bgr_0.1st_Vout_2.t23 GNDA 0.52755f
C1595 bgr_0.1st_Vout_2.t16 GNDA 0.52755f
C1596 bgr_0.1st_Vout_2.t19 GNDA 0.536536f
C1597 bgr_0.1st_Vout_2.t36 GNDA 0.536536f
C1598 bgr_0.1st_Vout_2.t29 GNDA 0.52755f
C1599 bgr_0.1st_Vout_2.t22 GNDA 0.52755f
C1600 bgr_0.1st_Vout_2.t26 GNDA 0.536536f
C1601 bgr_0.1st_Vout_2.t18 GNDA 0.536536f
C1602 bgr_0.1st_Vout_2.t15 GNDA 0.52755f
C1603 bgr_0.1st_Vout_2.t21 GNDA 0.52755f
C1604 bgr_0.1st_Vout_2.t14 GNDA 0.049375f
C1605 bgr_0.1st_Vout_2.t5 GNDA 0.013189f
C1606 bgr_0.1st_Vout_2.t4 GNDA 0.013189f
C1607 bgr_0.1st_Vout_2.n8 GNDA 0.026935f
C1608 bgr_0.1st_Vout_2.n9 GNDA 0.013946f
C1609 bgr_0.1st_Vout_2.n10 GNDA 0.013946f
C1610 bgr_0.1st_Vout_2.n11 GNDA 0.113739f
C1611 bgr_0.1st_Vout_2.n12 GNDA 0.15375f
C1612 bgr_0.1st_Vout_2.t9 GNDA 0.023066f
C1613 bgr_0.1st_Vout_2.n13 GNDA 0.117808f
C1614 bgr_0.1st_Vout_2.n14 GNDA 0.14843f
C1615 bgr_0.1st_Vout_2.t13 GNDA 0.04941f
C1616 bgr_0.1st_Vout_2.t20 GNDA 0.024683f
C1617 bgr_0.1st_Vout_2.t33 GNDA 0.018135f
C1618 bgr_0.1st_Vout_2.n15 GNDA 0.052887f
C1619 bgr_0.1st_Vout_2.t25 GNDA 0.024683f
C1620 bgr_0.1st_Vout_2.t34 GNDA 0.018135f
C1621 bgr_0.1st_Vout_2.n16 GNDA 0.052887f
C1622 bgr_0.1st_Vout_2.t6 GNDA 0.013189f
C1623 bgr_0.1st_Vout_2.t8 GNDA 0.013189f
C1624 bgr_0.1st_Vout_2.n17 GNDA 0.026935f
C1625 bgr_0.1st_Vout_2.n18 GNDA 0.202261f
C1626 bgr_0.1st_Vout_2.n19 GNDA 0.205909f
C1627 bgr_0.1st_Vout_2.n20 GNDA 0.026935f
C1628 bgr_0.1st_Vout_2.t3 GNDA 0.013189f
C1629 bgr_0.V_TOP.t36 GNDA 0.474011f
C1630 bgr_0.V_TOP.t24 GNDA 0.482085f
C1631 bgr_0.V_TOP.t30 GNDA 0.474011f
C1632 bgr_0.V_TOP.n0 GNDA 0.317809f
C1633 bgr_0.V_TOP.t25 GNDA 0.474011f
C1634 bgr_0.V_TOP.t19 GNDA 0.482085f
C1635 bgr_0.V_TOP.n1 GNDA 0.406686f
C1636 bgr_0.V_TOP.t16 GNDA 0.482085f
C1637 bgr_0.V_TOP.t22 GNDA 0.474011f
C1638 bgr_0.V_TOP.n2 GNDA 0.317809f
C1639 bgr_0.V_TOP.t18 GNDA 0.474011f
C1640 bgr_0.V_TOP.t44 GNDA 0.482085f
C1641 bgr_0.V_TOP.n3 GNDA 0.495564f
C1642 bgr_0.V_TOP.t39 GNDA 0.482085f
C1643 bgr_0.V_TOP.t49 GNDA 0.474011f
C1644 bgr_0.V_TOP.n4 GNDA 0.317809f
C1645 bgr_0.V_TOP.t42 GNDA 0.474011f
C1646 bgr_0.V_TOP.t32 GNDA 0.482085f
C1647 bgr_0.V_TOP.n5 GNDA 0.495564f
C1648 bgr_0.V_TOP.t14 GNDA 0.482085f
C1649 bgr_0.V_TOP.t21 GNDA 0.474011f
C1650 bgr_0.V_TOP.n6 GNDA 0.317809f
C1651 bgr_0.V_TOP.t15 GNDA 0.474011f
C1652 bgr_0.V_TOP.t40 GNDA 0.482085f
C1653 bgr_0.V_TOP.n7 GNDA 0.495564f
C1654 bgr_0.V_TOP.t28 GNDA 0.482085f
C1655 bgr_0.V_TOP.t37 GNDA 0.474011f
C1656 bgr_0.V_TOP.n8 GNDA 0.406686f
C1657 bgr_0.V_TOP.t47 GNDA 0.474011f
C1658 bgr_0.V_TOP.n9 GNDA 0.20738f
C1659 bgr_0.V_TOP.n10 GNDA 0.709704f
C1660 bgr_0.V_TOP.n11 GNDA 0.094802f
C1661 bgr_0.V_TOP.t10 GNDA 0.01185f
C1662 bgr_0.V_TOP.t2 GNDA 0.01185f
C1663 bgr_0.V_TOP.n12 GNDA 0.024201f
C1664 bgr_0.V_TOP.n13 GNDA 0.167471f
C1665 bgr_0.V_TOP.t6 GNDA 0.136551f
C1666 bgr_0.V_TOP.t41 GNDA 0.124428f
C1667 bgr_0.V_TOP.t38 GNDA 0.124428f
C1668 bgr_0.V_TOP.t17 GNDA 0.124428f
C1669 bgr_0.V_TOP.t26 GNDA 0.124428f
C1670 bgr_0.V_TOP.t34 GNDA 0.124428f
C1671 bgr_0.V_TOP.t46 GNDA 0.124428f
C1672 bgr_0.V_TOP.t45 GNDA 0.162658f
C1673 bgr_0.V_TOP.n14 GNDA 0.090938f
C1674 bgr_0.V_TOP.n15 GNDA 0.066362f
C1675 bgr_0.V_TOP.n16 GNDA 0.066362f
C1676 bgr_0.V_TOP.n17 GNDA 0.066362f
C1677 bgr_0.V_TOP.n18 GNDA 0.066362f
C1678 bgr_0.V_TOP.n19 GNDA 0.061574f
C1679 bgr_0.V_TOP.t29 GNDA 0.124428f
C1680 bgr_0.V_TOP.t20 GNDA 0.124428f
C1681 bgr_0.V_TOP.t43 GNDA 0.124428f
C1682 bgr_0.V_TOP.t31 GNDA 0.124428f
C1683 bgr_0.V_TOP.t33 GNDA 0.124428f
C1684 bgr_0.V_TOP.t23 GNDA 0.124428f
C1685 bgr_0.V_TOP.t48 GNDA 0.124428f
C1686 bgr_0.V_TOP.t35 GNDA 0.124428f
C1687 bgr_0.V_TOP.t27 GNDA 0.162658f
C1688 bgr_0.V_TOP.n20 GNDA 0.090938f
C1689 bgr_0.V_TOP.n21 GNDA 0.066362f
C1690 bgr_0.V_TOP.n22 GNDA 0.066362f
C1691 bgr_0.V_TOP.n23 GNDA 0.066362f
C1692 bgr_0.V_TOP.n24 GNDA 0.066362f
C1693 bgr_0.V_TOP.n25 GNDA 0.066362f
C1694 bgr_0.V_TOP.n26 GNDA 0.066362f
C1695 bgr_0.V_TOP.n27 GNDA 0.061574f
C1696 bgr_0.V_TOP.n28 GNDA 0.025195f
C1697 bgr_0.V_TOP.n29 GNDA 0.466786f
C1698 bgr_0.V_TOP.n30 GNDA 0.098389f
C1699 bgr_0.V_TOP.n31 GNDA 0.099945f
C1700 bgr_0.V_TOP.t12 GNDA 0.01185f
C1701 bgr_0.V_TOP.t7 GNDA 0.01185f
C1702 bgr_0.V_TOP.n32 GNDA 0.024201f
C1703 bgr_0.V_TOP.n33 GNDA 0.149457f
C1704 bgr_0.V_TOP.n34 GNDA 0.141056f
C1705 bgr_0.V_TOP.t3 GNDA 0.01185f
C1706 bgr_0.V_TOP.t13 GNDA 0.01185f
C1707 bgr_0.V_TOP.n35 GNDA 0.025558f
C1708 bgr_0.V_TOP.t0 GNDA 0.01185f
C1709 bgr_0.V_TOP.t4 GNDA 0.01185f
C1710 bgr_0.V_TOP.n36 GNDA 0.025392f
C1711 bgr_0.V_TOP.n37 GNDA 0.409784f
C1712 bgr_0.V_TOP.n38 GNDA 0.154984f
C1713 bgr_0.V_TOP.t11 GNDA 0.01185f
C1714 bgr_0.V_TOP.t9 GNDA 0.01185f
C1715 bgr_0.V_TOP.n39 GNDA 0.024201f
C1716 bgr_0.V_TOP.n40 GNDA 0.113621f
C1717 bgr_0.V_TOP.n41 GNDA 0.141056f
C1718 bgr_0.V_TOP.t5 GNDA 0.01185f
C1719 bgr_0.V_TOP.t8 GNDA 0.01185f
C1720 bgr_0.V_TOP.n42 GNDA 0.024201f
C1721 bgr_0.V_TOP.n43 GNDA 0.167471f
C1722 bgr_0.V_TOP.n44 GNDA 0.482466f
C1723 bgr_0.V_TOP.n45 GNDA 0.950439f
C1724 bgr_0.V_TOP.t1 GNDA 0.133346f
C1725 VOUT-.t9 GNDA 0.04706f
C1726 VOUT-.t11 GNDA 0.04706f
C1727 VOUT-.n0 GNDA 0.096426f
C1728 VOUT-.n1 GNDA 0.246395f
C1729 VOUT-.n2 GNDA 0.03392f
C1730 VOUT-.n3 GNDA 0.059842f
C1731 VOUT-.t6 GNDA 0.04706f
C1732 VOUT-.t16 GNDA 0.04706f
C1733 VOUT-.n4 GNDA 0.096426f
C1734 VOUT-.n5 GNDA 0.287036f
C1735 VOUT-.t8 GNDA 0.04706f
C1736 VOUT-.t12 GNDA 0.04706f
C1737 VOUT-.n6 GNDA 0.096426f
C1738 VOUT-.n7 GNDA 0.282019f
C1739 VOUT-.n8 GNDA 0.059842f
C1740 VOUT-.n9 GNDA 0.03392f
C1741 VOUT-.t2 GNDA 0.04706f
C1742 VOUT-.t3 GNDA 0.04706f
C1743 VOUT-.n10 GNDA 0.096426f
C1744 VOUT-.n11 GNDA 0.282019f
C1745 VOUT-.n12 GNDA 0.03392f
C1746 VOUT-.t1 GNDA 0.04706f
C1747 VOUT-.t10 GNDA 0.04706f
C1748 VOUT-.n13 GNDA 0.096426f
C1749 VOUT-.n14 GNDA 0.282019f
C1750 VOUT-.n15 GNDA 0.03392f
C1751 VOUT-.n16 GNDA 0.059842f
C1752 VOUT-.t4 GNDA 0.04706f
C1753 VOUT-.t5 GNDA 0.04706f
C1754 VOUT-.n17 GNDA 0.096426f
C1755 VOUT-.n18 GNDA 0.287036f
C1756 VOUT-.n19 GNDA 0.049452f
C1757 VOUT-.n20 GNDA 0.202653f
C1758 VOUT-.t117 GNDA 0.319077f
C1759 VOUT-.t25 GNDA 0.313734f
C1760 VOUT-.n21 GNDA 0.210348f
C1761 VOUT-.t124 GNDA 0.313734f
C1762 VOUT-.n22 GNDA 0.137258f
C1763 VOUT-.t72 GNDA 0.319077f
C1764 VOUT-.t38 GNDA 0.313734f
C1765 VOUT-.n23 GNDA 0.210348f
C1766 VOUT-.t127 GNDA 0.313734f
C1767 VOUT-.t34 GNDA 0.318408f
C1768 VOUT-.t86 GNDA 0.318408f
C1769 VOUT-.t42 GNDA 0.318408f
C1770 VOUT-.t96 GNDA 0.318408f
C1771 VOUT-.t143 GNDA 0.318408f
C1772 VOUT-.t106 GNDA 0.318408f
C1773 VOUT-.t154 GNDA 0.318408f
C1774 VOUT-.t64 GNDA 0.318408f
C1775 VOUT-.t116 GNDA 0.318408f
C1776 VOUT-.t73 GNDA 0.318408f
C1777 VOUT-.t149 GNDA 0.313734f
C1778 VOUT-.n24 GNDA 0.211017f
C1779 VOUT-.t58 GNDA 0.313734f
C1780 VOUT-.n25 GNDA 0.269842f
C1781 VOUT-.t97 GNDA 0.313734f
C1782 VOUT-.n26 GNDA 0.269842f
C1783 VOUT-.t131 GNDA 0.313734f
C1784 VOUT-.n27 GNDA 0.269842f
C1785 VOUT-.t24 GNDA 0.313734f
C1786 VOUT-.n28 GNDA 0.269842f
C1787 VOUT-.t75 GNDA 0.313734f
C1788 VOUT-.n29 GNDA 0.269842f
C1789 VOUT-.t113 GNDA 0.313734f
C1790 VOUT-.n30 GNDA 0.269842f
C1791 VOUT-.t144 GNDA 0.313734f
C1792 VOUT-.n31 GNDA 0.269842f
C1793 VOUT-.t54 GNDA 0.313734f
C1794 VOUT-.n32 GNDA 0.269842f
C1795 VOUT-.t94 GNDA 0.313734f
C1796 VOUT-.n33 GNDA 0.269842f
C1797 VOUT-.n34 GNDA 0.254908f
C1798 VOUT-.t37 GNDA 0.319077f
C1799 VOUT-.t142 GNDA 0.313734f
C1800 VOUT-.n35 GNDA 0.210348f
C1801 VOUT-.t93 GNDA 0.313734f
C1802 VOUT-.t20 GNDA 0.319077f
C1803 VOUT-.t57 GNDA 0.313734f
C1804 VOUT-.n36 GNDA 0.210348f
C1805 VOUT-.n37 GNDA 0.254908f
C1806 VOUT-.t79 GNDA 0.319077f
C1807 VOUT-.t41 GNDA 0.313734f
C1808 VOUT-.n38 GNDA 0.210348f
C1809 VOUT-.t133 GNDA 0.313734f
C1810 VOUT-.t60 GNDA 0.319077f
C1811 VOUT-.t100 GNDA 0.313734f
C1812 VOUT-.n39 GNDA 0.210348f
C1813 VOUT-.n40 GNDA 0.254908f
C1814 VOUT-.t121 GNDA 0.319077f
C1815 VOUT-.t83 GNDA 0.313734f
C1816 VOUT-.n41 GNDA 0.210348f
C1817 VOUT-.t31 GNDA 0.313734f
C1818 VOUT-.t104 GNDA 0.319077f
C1819 VOUT-.t137 GNDA 0.313734f
C1820 VOUT-.n42 GNDA 0.210348f
C1821 VOUT-.n43 GNDA 0.254908f
C1822 VOUT-.t84 GNDA 0.319077f
C1823 VOUT-.t49 GNDA 0.313734f
C1824 VOUT-.n44 GNDA 0.210348f
C1825 VOUT-.t138 GNDA 0.313734f
C1826 VOUT-.t66 GNDA 0.319077f
C1827 VOUT-.t103 GNDA 0.313734f
C1828 VOUT-.n45 GNDA 0.210348f
C1829 VOUT-.n46 GNDA 0.254908f
C1830 VOUT-.t108 GNDA 0.319077f
C1831 VOUT-.t69 GNDA 0.313734f
C1832 VOUT-.n47 GNDA 0.210348f
C1833 VOUT-.t90 GNDA 0.313734f
C1834 VOUT-.n48 GNDA 0.137258f
C1835 VOUT-.t67 GNDA 0.319077f
C1836 VOUT-.t30 GNDA 0.313734f
C1837 VOUT-.n49 GNDA 0.210348f
C1838 VOUT-.t51 GNDA 0.313734f
C1839 VOUT-.t53 GNDA 0.318408f
C1840 VOUT-.t156 GNDA 0.318408f
C1841 VOUT-.t44 GNDA 0.319077f
C1842 VOUT-.t136 GNDA 0.313734f
C1843 VOUT-.n50 GNDA 0.210348f
C1844 VOUT-.t101 GNDA 0.313734f
C1845 VOUT-.n51 GNDA 0.132356f
C1846 VOUT-.t36 GNDA 0.318408f
C1847 VOUT-.t151 GNDA 0.319077f
C1848 VOUT-.t98 GNDA 0.313734f
C1849 VOUT-.n52 GNDA 0.210348f
C1850 VOUT-.t59 GNDA 0.313734f
C1851 VOUT-.n53 GNDA 0.132356f
C1852 VOUT-.t140 GNDA 0.318408f
C1853 VOUT-.t118 GNDA 0.319077f
C1854 VOUT-.t56 GNDA 0.313734f
C1855 VOUT-.n54 GNDA 0.210348f
C1856 VOUT-.t21 GNDA 0.313734f
C1857 VOUT-.n55 GNDA 0.132356f
C1858 VOUT-.t105 GNDA 0.318408f
C1859 VOUT-.t65 GNDA 0.319077f
C1860 VOUT-.t80 GNDA 0.313734f
C1861 VOUT-.n56 GNDA 0.210348f
C1862 VOUT-.t43 GNDA 0.313734f
C1863 VOUT-.n57 GNDA 0.132356f
C1864 VOUT-.t125 GNDA 0.318408f
C1865 VOUT-.t145 GNDA 0.318671f
C1866 VOUT-.t87 GNDA 0.318408f
C1867 VOUT-.t110 GNDA 0.318671f
C1868 VOUT-.t50 GNDA 0.318408f
C1869 VOUT-.t70 GNDA 0.318671f
C1870 VOUT-.t150 GNDA 0.318408f
C1871 VOUT-.t95 GNDA 0.318671f
C1872 VOUT-.t32 GNDA 0.318408f
C1873 VOUT-.t134 GNDA 0.313734f
C1874 VOUT-.n58 GNDA 0.34726f
C1875 VOUT-.t111 GNDA 0.313734f
C1876 VOUT-.n59 GNDA 0.406085f
C1877 VOUT-.t147 GNDA 0.313734f
C1878 VOUT-.n60 GNDA 0.406085f
C1879 VOUT-.t45 GNDA 0.313734f
C1880 VOUT-.n61 GNDA 0.406085f
C1881 VOUT-.t85 GNDA 0.313734f
C1882 VOUT-.n62 GNDA 0.333569f
C1883 VOUT-.t61 GNDA 0.313734f
C1884 VOUT-.n63 GNDA 0.333569f
C1885 VOUT-.t102 GNDA 0.313734f
C1886 VOUT-.n64 GNDA 0.333569f
C1887 VOUT-.t139 GNDA 0.313734f
C1888 VOUT-.n65 GNDA 0.333569f
C1889 VOUT-.t119 GNDA 0.313734f
C1890 VOUT-.n66 GNDA 0.269842f
C1891 VOUT-.t155 GNDA 0.313734f
C1892 VOUT-.n67 GNDA 0.269842f
C1893 VOUT-.n68 GNDA 0.254908f
C1894 VOUT-.t27 GNDA 0.319077f
C1895 VOUT-.t130 GNDA 0.313734f
C1896 VOUT-.n69 GNDA 0.210348f
C1897 VOUT-.t152 GNDA 0.313734f
C1898 VOUT-.t76 GNDA 0.319077f
C1899 VOUT-.t115 GNDA 0.313734f
C1900 VOUT-.n70 GNDA 0.210348f
C1901 VOUT-.n71 GNDA 0.254908f
C1902 VOUT-.t62 GNDA 0.319077f
C1903 VOUT-.t23 GNDA 0.313734f
C1904 VOUT-.n72 GNDA 0.210348f
C1905 VOUT-.t47 GNDA 0.313734f
C1906 VOUT-.t112 GNDA 0.319077f
C1907 VOUT-.t148 GNDA 0.313734f
C1908 VOUT-.n73 GNDA 0.210348f
C1909 VOUT-.n74 GNDA 0.254908f
C1910 VOUT-.t114 GNDA 0.319077f
C1911 VOUT-.t78 GNDA 0.313734f
C1912 VOUT-.n75 GNDA 0.210348f
C1913 VOUT-.t26 GNDA 0.313734f
C1914 VOUT-.t99 GNDA 0.319077f
C1915 VOUT-.t132 GNDA 0.313734f
C1916 VOUT-.n76 GNDA 0.210348f
C1917 VOUT-.n77 GNDA 0.254908f
C1918 VOUT-.t74 GNDA 0.319077f
C1919 VOUT-.t39 GNDA 0.313734f
C1920 VOUT-.n78 GNDA 0.210348f
C1921 VOUT-.t128 GNDA 0.313734f
C1922 VOUT-.t55 GNDA 0.319077f
C1923 VOUT-.t92 GNDA 0.313734f
C1924 VOUT-.n79 GNDA 0.210348f
C1925 VOUT-.n80 GNDA 0.254908f
C1926 VOUT-.t109 GNDA 0.319077f
C1927 VOUT-.t71 GNDA 0.313734f
C1928 VOUT-.n81 GNDA 0.210348f
C1929 VOUT-.t19 GNDA 0.313734f
C1930 VOUT-.t91 GNDA 0.319077f
C1931 VOUT-.t126 GNDA 0.313734f
C1932 VOUT-.n82 GNDA 0.210348f
C1933 VOUT-.n83 GNDA 0.254908f
C1934 VOUT-.t68 GNDA 0.319077f
C1935 VOUT-.t33 GNDA 0.313734f
C1936 VOUT-.n84 GNDA 0.210348f
C1937 VOUT-.t122 GNDA 0.313734f
C1938 VOUT-.t52 GNDA 0.319077f
C1939 VOUT-.t88 GNDA 0.313734f
C1940 VOUT-.n85 GNDA 0.210348f
C1941 VOUT-.n86 GNDA 0.254908f
C1942 VOUT-.t29 GNDA 0.319077f
C1943 VOUT-.t135 GNDA 0.313734f
C1944 VOUT-.n87 GNDA 0.210348f
C1945 VOUT-.t82 GNDA 0.313734f
C1946 VOUT-.t153 GNDA 0.319077f
C1947 VOUT-.t48 GNDA 0.313734f
C1948 VOUT-.n88 GNDA 0.210348f
C1949 VOUT-.n89 GNDA 0.254908f
C1950 VOUT-.t63 GNDA 0.319077f
C1951 VOUT-.t28 GNDA 0.313734f
C1952 VOUT-.n90 GNDA 0.210348f
C1953 VOUT-.t120 GNDA 0.313734f
C1954 VOUT-.t46 GNDA 0.319077f
C1955 VOUT-.t81 GNDA 0.313734f
C1956 VOUT-.n91 GNDA 0.210348f
C1957 VOUT-.n92 GNDA 0.254908f
C1958 VOUT-.t22 GNDA 0.319077f
C1959 VOUT-.t129 GNDA 0.313734f
C1960 VOUT-.n93 GNDA 0.210348f
C1961 VOUT-.t77 GNDA 0.313734f
C1962 VOUT-.t146 GNDA 0.319077f
C1963 VOUT-.t40 GNDA 0.313734f
C1964 VOUT-.n94 GNDA 0.210348f
C1965 VOUT-.n95 GNDA 0.254908f
C1966 VOUT-.t123 GNDA 0.319077f
C1967 VOUT-.t89 GNDA 0.313734f
C1968 VOUT-.n96 GNDA 0.210348f
C1969 VOUT-.t35 GNDA 0.313734f
C1970 VOUT-.n97 GNDA 0.254908f
C1971 VOUT-.t141 GNDA 0.313734f
C1972 VOUT-.n98 GNDA 0.137258f
C1973 VOUT-.t107 GNDA 0.313734f
C1974 VOUT-.n99 GNDA 0.249494f
C1975 VOUT-.n100 GNDA 0.31936f
C1976 VOUT-.n101 GNDA 0.082953f
C1977 VOUT-.t7 GNDA 0.054903f
C1978 VOUT-.t13 GNDA 0.054903f
C1979 VOUT-.n102 GNDA 0.117966f
C1980 VOUT-.n103 GNDA 0.329815f
C1981 VOUT-.t0 GNDA 0.054903f
C1982 VOUT-.t18 GNDA 0.054903f
C1983 VOUT-.n104 GNDA 0.117966f
C1984 VOUT-.n105 GNDA 0.317784f
C1985 VOUT-.n106 GNDA 0.115148f
C1986 VOUT-.t14 GNDA 0.054903f
C1987 VOUT-.t17 GNDA 0.054903f
C1988 VOUT-.n107 GNDA 0.117966f
C1989 VOUT-.n108 GNDA 0.3238f
C1990 VOUT-.n109 GNDA 0.057818f
C1991 VOUT-.t15 GNDA 0.09073f
C1992 VOUT-.n110 GNDA 0.107022f
C1993 bgr_0.1st_Vout_1.n0 GNDA 0.816409f
C1994 bgr_0.1st_Vout_1.n1 GNDA 0.358128f
C1995 bgr_0.1st_Vout_1.n2 GNDA 1.47499f
C1996 bgr_0.1st_Vout_1.n3 GNDA 1.37484f
C1997 bgr_0.1st_Vout_1.n4 GNDA 1.34019f
C1998 bgr_0.1st_Vout_1.n5 GNDA 0.114413f
C1999 bgr_0.1st_Vout_1.t2 GNDA 0.013354f
C2000 bgr_0.1st_Vout_1.t11 GNDA 0.543245f
C2001 bgr_0.1st_Vout_1.t16 GNDA 0.534147f
C2002 bgr_0.1st_Vout_1.t31 GNDA 0.543245f
C2003 bgr_0.1st_Vout_1.t36 GNDA 0.534147f
C2004 bgr_0.1st_Vout_1.t33 GNDA 0.543245f
C2005 bgr_0.1st_Vout_1.t35 GNDA 0.534147f
C2006 bgr_0.1st_Vout_1.t21 GNDA 0.543245f
C2007 bgr_0.1st_Vout_1.t30 GNDA 0.534147f
C2008 bgr_0.1st_Vout_1.t23 GNDA 0.543245f
C2009 bgr_0.1st_Vout_1.t28 GNDA 0.534147f
C2010 bgr_0.1st_Vout_1.t14 GNDA 0.543245f
C2011 bgr_0.1st_Vout_1.t20 GNDA 0.534147f
C2012 bgr_0.1st_Vout_1.t32 GNDA 0.543245f
C2013 bgr_0.1st_Vout_1.t34 GNDA 0.534147f
C2014 bgr_0.1st_Vout_1.t19 GNDA 0.543245f
C2015 bgr_0.1st_Vout_1.t26 GNDA 0.534147f
C2016 bgr_0.1st_Vout_1.t22 GNDA 0.543245f
C2017 bgr_0.1st_Vout_1.t25 GNDA 0.534147f
C2018 bgr_0.1st_Vout_1.t18 GNDA 0.534147f
C2019 bgr_0.1st_Vout_1.t12 GNDA 0.534147f
C2020 bgr_0.1st_Vout_1.t27 GNDA 0.049992f
C2021 bgr_0.1st_Vout_1.n6 GNDA 1.04864f
C2022 bgr_0.1st_Vout_1.n7 GNDA 0.069966f
C2023 bgr_0.1st_Vout_1.t3 GNDA 0.013354f
C2024 bgr_0.1st_Vout_1.t1 GNDA 0.013354f
C2025 bgr_0.1st_Vout_1.n8 GNDA 0.027271f
C2026 bgr_0.1st_Vout_1.n9 GNDA 0.208484f
C2027 bgr_0.1st_Vout_1.n10 GNDA 0.014121f
C2028 bgr_0.1st_Vout_1.t7 GNDA 0.023354f
C2029 bgr_0.1st_Vout_1.n11 GNDA 0.119281f
C2030 bgr_0.1st_Vout_1.n12 GNDA 0.155672f
C2031 bgr_0.1st_Vout_1.n13 GNDA 0.014121f
C2032 bgr_0.1st_Vout_1.n14 GNDA 0.115161f
C2033 bgr_0.1st_Vout_1.n15 GNDA 0.150286f
C2034 bgr_0.1st_Vout_1.t15 GNDA 0.024992f
C2035 bgr_0.1st_Vout_1.t24 GNDA 0.018361f
C2036 bgr_0.1st_Vout_1.n16 GNDA 0.053548f
C2037 bgr_0.1st_Vout_1.n17 GNDA 0.110964f
C2038 bgr_0.1st_Vout_1.t17 GNDA 0.050028f
C2039 bgr_0.1st_Vout_1.n18 GNDA 0.140566f
C2040 bgr_0.1st_Vout_1.t13 GNDA 0.024992f
C2041 bgr_0.1st_Vout_1.t29 GNDA 0.018361f
C2042 bgr_0.1st_Vout_1.n19 GNDA 0.053548f
C2043 bgr_0.1st_Vout_1.n20 GNDA 0.110964f
C2044 bgr_0.1st_Vout_1.n21 GNDA 0.059208f
C2045 bgr_0.1st_Vout_1.n22 GNDA 0.081973f
C2046 bgr_0.1st_Vout_1.t4 GNDA 0.013354f
C2047 bgr_0.1st_Vout_1.t0 GNDA 0.013354f
C2048 bgr_0.1st_Vout_1.n23 GNDA 0.027271f
C2049 bgr_0.1st_Vout_1.n24 GNDA 0.13771f
C2050 bgr_0.1st_Vout_1.n25 GNDA 0.20479f
C2051 bgr_0.1st_Vout_1.n26 GNDA 0.208484f
C2052 bgr_0.1st_Vout_1.n27 GNDA 0.027271f
C2053 bgr_0.1st_Vout_1.t5 GNDA 0.013354f
C2054 bgr_0.V_mir1.t9 GNDA 0.031034f
C2055 bgr_0.V_mir1.t1 GNDA 0.015517f
C2056 bgr_0.V_mir1.t0 GNDA 0.015517f
C2057 bgr_0.V_mir1.n0 GNDA 0.032817f
C2058 bgr_0.V_mir1.n1 GNDA 0.172902f
C2059 bgr_0.V_mir1.t2 GNDA 0.054276f
C2060 bgr_0.V_mir1.n2 GNDA 0.277214f
C2061 bgr_0.V_mir1.n3 GNDA 0.351139f
C2062 bgr_0.V_mir1.t16 GNDA 0.015517f
C2063 bgr_0.V_mir1.t3 GNDA 0.015517f
C2064 bgr_0.V_mir1.n4 GNDA 0.032817f
C2065 bgr_0.V_mir1.n5 GNDA 0.21593f
C2066 bgr_0.V_mir1.n6 GNDA 0.356077f
C2067 bgr_0.V_mir1.n7 GNDA 0.181138f
C2068 bgr_0.V_mir1.t14 GNDA 0.047277f
C2069 bgr_0.V_mir1.t8 GNDA 0.037241f
C2070 bgr_0.V_mir1.t18 GNDA 0.037241f
C2071 bgr_0.V_mir1.t22 GNDA 0.060113f
C2072 bgr_0.V_mir1.n8 GNDA 0.067129f
C2073 bgr_0.V_mir1.n9 GNDA 0.045857f
C2074 bgr_0.V_mir1.n10 GNDA 0.074211f
C2075 bgr_0.V_mir1.n11 GNDA 0.199395f
C2076 bgr_0.V_mir1.t7 GNDA 0.031034f
C2077 bgr_0.V_mir1.t11 GNDA 0.031034f
C2078 bgr_0.V_mir1.n12 GNDA 0.06338f
C2079 bgr_0.V_mir1.n13 GNDA 0.260312f
C2080 bgr_0.V_mir1.t12 GNDA 0.047277f
C2081 bgr_0.V_mir1.t4 GNDA 0.037241f
C2082 bgr_0.V_mir1.t19 GNDA 0.037241f
C2083 bgr_0.V_mir1.t21 GNDA 0.060113f
C2084 bgr_0.V_mir1.n14 GNDA 0.067129f
C2085 bgr_0.V_mir1.n15 GNDA 0.045857f
C2086 bgr_0.V_mir1.n16 GNDA 0.074211f
C2087 bgr_0.V_mir1.t6 GNDA 0.047277f
C2088 bgr_0.V_mir1.t10 GNDA 0.037241f
C2089 bgr_0.V_mir1.t17 GNDA 0.037241f
C2090 bgr_0.V_mir1.t20 GNDA 0.060113f
C2091 bgr_0.V_mir1.n17 GNDA 0.067129f
C2092 bgr_0.V_mir1.n18 GNDA 0.045857f
C2093 bgr_0.V_mir1.n19 GNDA 0.074211f
C2094 bgr_0.V_mir1.n20 GNDA 0.166486f
C2095 bgr_0.V_mir1.n21 GNDA 0.450644f
C2096 bgr_0.V_mir1.n22 GNDA 0.166486f
C2097 bgr_0.V_mir1.t13 GNDA 0.031034f
C2098 bgr_0.V_mir1.t5 GNDA 0.031034f
C2099 bgr_0.V_mir1.n23 GNDA 0.06338f
C2100 bgr_0.V_mir1.n24 GNDA 0.260312f
C2101 bgr_0.V_mir1.n25 GNDA 0.463152f
C2102 bgr_0.V_mir1.n26 GNDA 0.213276f
C2103 bgr_0.V_mir1.n27 GNDA 0.06338f
C2104 bgr_0.V_mir1.t15 GNDA 0.031034f
C2105 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 GNDA 0.344411f
C2106 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 GNDA 0.34556f
C2107 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 GNDA 0.185607f
C2108 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 GNDA 0.198192f
C2109 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 GNDA 0.344411f
C2110 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 GNDA 0.34556f
C2111 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 GNDA 0.185607f
C2112 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 GNDA 0.216737f
C2113 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 GNDA 0.344411f
C2114 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 GNDA 0.34556f
C2115 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 GNDA 0.185607f
C2116 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 GNDA 0.216737f
C2117 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 GNDA 0.344411f
C2118 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 GNDA 0.34556f
C2119 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 GNDA 0.185607f
C2120 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 GNDA 0.216737f
C2121 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 GNDA 0.344411f
C2122 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 GNDA 0.34556f
C2123 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 GNDA 0.364105f
C2124 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 GNDA 0.364105f
C2125 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 GNDA 0.185607f
C2126 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 GNDA 0.216737f
C2127 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 GNDA 0.344411f
C2128 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 GNDA 0.34556f
C2129 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 GNDA 0.364105f
C2130 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 GNDA 0.364105f
C2131 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 GNDA 0.185607f
C2132 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 GNDA 0.216737f
C2133 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 GNDA 0.34556f
C2134 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 GNDA 0.346812f
C2135 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 GNDA 0.34556f
C2136 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 GNDA 0.348269f
C2137 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 GNDA 0.378792f
C2138 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 GNDA 0.34556f
C2139 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 GNDA 0.346812f
C2140 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 GNDA 0.34556f
C2141 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 GNDA 0.346812f
C2142 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 GNDA 0.34556f
C2143 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 GNDA 0.346812f
C2144 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 GNDA 0.34556f
C2145 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 GNDA 0.346812f
C2146 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 GNDA 0.34556f
C2147 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 GNDA 0.346812f
C2148 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 GNDA 0.34556f
C2149 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 GNDA 0.346812f
C2150 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 GNDA 0.34556f
C2151 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 GNDA 0.346812f
C2152 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 GNDA 0.34556f
C2153 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 GNDA 0.346812f
C2154 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 GNDA 0.34556f
C2155 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 GNDA 0.346812f
C2156 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 GNDA 0.34556f
C2157 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 GNDA 0.346812f
C2158 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 GNDA 0.34556f
C2159 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 GNDA 0.346812f
C2160 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 GNDA 0.34556f
C2161 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 GNDA 0.346812f
C2162 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 GNDA 0.34556f
C2163 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 GNDA 0.346812f
C2164 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 GNDA 0.34556f
C2165 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 GNDA 0.346812f
C2166 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 GNDA 0.34556f
C2167 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 GNDA 0.346812f
C2168 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 GNDA 0.34556f
C2169 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 GNDA 0.346812f
C2170 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 GNDA 0.34556f
C2171 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 GNDA 0.346812f
C2172 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 GNDA 0.34556f
C2173 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 GNDA 0.346812f
C2174 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 GNDA 0.34556f
C2175 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 GNDA 0.346812f
C2176 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 GNDA 0.34556f
C2177 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 GNDA 0.346812f
C2178 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 GNDA 0.34556f
C2179 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 GNDA 0.346812f
C2180 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 GNDA 0.34556f
C2181 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 GNDA 0.346812f
C2182 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 GNDA 0.34556f
C2183 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 GNDA 0.346812f
C2184 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 GNDA 0.34556f
C2185 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 GNDA 0.346812f
C2186 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 GNDA 0.34556f
C2187 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 GNDA 0.346812f
C2188 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 GNDA 0.34556f
C2189 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 GNDA 0.346812f
C2190 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 GNDA 0.34556f
C2191 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 GNDA 0.346812f
C2192 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 GNDA 0.34556f
C2193 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 GNDA 0.346812f
C2194 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 GNDA 0.34556f
C2195 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 GNDA 0.362503f
C2196 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 GNDA 0.34556f
C2197 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 GNDA 0.185607f
C2198 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 GNDA 0.198646f
C2199 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 GNDA 0.34556f
C2200 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 GNDA 0.185607f
C2201 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 GNDA 0.197043f
C2202 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 GNDA 0.34556f
C2203 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 GNDA 0.185607f
C2204 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 GNDA 0.197043f
C2205 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 GNDA 0.34556f
C2206 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 GNDA 0.185607f
C2207 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 GNDA 0.197043f
C2208 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 GNDA 0.34556f
C2209 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 GNDA 0.185607f
C2210 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 GNDA 0.197043f
C2211 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 GNDA 0.34556f
C2212 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 GNDA 0.185607f
C2213 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 GNDA 0.197043f
C2214 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 GNDA 0.34556f
C2215 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 GNDA 0.185607f
C2216 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 GNDA 0.197043f
C2217 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 GNDA 0.34556f
C2218 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 GNDA 0.185607f
C2219 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 GNDA 0.197043f
C2220 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 GNDA 0.34556f
C2221 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 GNDA 0.185607f
C2222 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 GNDA 0.197043f
C2223 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 GNDA 0.34556f
C2224 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 GNDA 0.346812f
C2225 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 GNDA 0.34556f
C2226 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 GNDA 0.346812f
C2227 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 GNDA 0.167062f
C2228 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 GNDA 0.215485f
C2229 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 GNDA 0.184458f
C2230 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 GNDA 0.23403f
C2231 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 GNDA 0.184458f
C2232 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 GNDA 0.251323f
C2233 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 GNDA 0.184458f
C2234 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 GNDA 0.251323f
C2235 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 GNDA 0.184458f
C2236 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 GNDA 0.251323f
C2237 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 GNDA 0.184458f
C2238 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 GNDA 0.251323f
C2239 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 GNDA 0.184458f
C2240 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 GNDA 0.251323f
C2241 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 GNDA 0.184458f
C2242 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 GNDA 0.251323f
C2243 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 GNDA 0.184458f
C2244 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 GNDA 0.251323f
C2245 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 GNDA 0.184458f
C2246 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 GNDA 0.251323f
C2247 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 GNDA 0.184458f
C2248 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 GNDA 0.251323f
C2249 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 GNDA 0.184458f
C2250 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 GNDA 0.251323f
C2251 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 GNDA 0.184458f
C2252 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 GNDA 0.251323f
C2253 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 GNDA 0.184458f
C2254 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 GNDA 0.251323f
C2255 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 GNDA 0.184458f
C2256 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 GNDA 0.251323f
C2257 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 GNDA 0.184458f
C2258 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 GNDA 0.251323f
C2259 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 GNDA 0.184458f
C2260 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 GNDA 0.23403f
C2261 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 GNDA 0.344411f
C2262 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 GNDA 0.167062f
C2263 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 GNDA 0.216737f
C2264 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 GNDA 0.344411f
C2265 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 GNDA 0.167062f
C2266 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 GNDA 0.216737f
C2267 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 GNDA 0.344411f
C2268 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 GNDA 0.34556f
C2269 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 GNDA 0.364105f
C2270 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 GNDA 0.364105f
C2271 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 GNDA 0.185607f
C2272 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 GNDA 0.216737f
C2273 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 GNDA 0.344411f
C2274 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 GNDA 0.216737f
C2275 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 GNDA 0.185607f
C2276 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 GNDA 0.364105f
C2277 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 GNDA 0.364105f
C2278 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 GNDA 0.435648f
C2279 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 GNDA 0.292454f
C2280 VOUT+.n0 GNDA 0.082952f
C2281 VOUT+.t5 GNDA 0.054903f
C2282 VOUT+.t17 GNDA 0.054903f
C2283 VOUT+.n1 GNDA 0.117965f
C2284 VOUT+.n2 GNDA 0.329812f
C2285 VOUT+.t6 GNDA 0.054903f
C2286 VOUT+.t3 GNDA 0.054903f
C2287 VOUT+.n3 GNDA 0.117965f
C2288 VOUT+.n4 GNDA 0.317781f
C2289 VOUT+.n5 GNDA 0.115146f
C2290 VOUT+.t0 GNDA 0.054903f
C2291 VOUT+.t4 GNDA 0.054903f
C2292 VOUT+.n6 GNDA 0.117965f
C2293 VOUT+.n7 GNDA 0.323796f
C2294 VOUT+.n8 GNDA 0.057818f
C2295 VOUT+.t18 GNDA 0.090729f
C2296 VOUT+.n9 GNDA 0.110958f
C2297 VOUT+.t8 GNDA 0.04706f
C2298 VOUT+.t12 GNDA 0.04706f
C2299 VOUT+.n10 GNDA 0.096425f
C2300 VOUT+.n11 GNDA 0.246393f
C2301 VOUT+.t1 GNDA 0.04706f
C2302 VOUT+.t13 GNDA 0.04706f
C2303 VOUT+.n12 GNDA 0.096425f
C2304 VOUT+.n13 GNDA 0.287033f
C2305 VOUT+.n14 GNDA 0.03392f
C2306 VOUT+.n15 GNDA 0.059841f
C2307 VOUT+.t16 GNDA 0.04706f
C2308 VOUT+.t2 GNDA 0.04706f
C2309 VOUT+.n16 GNDA 0.096425f
C2310 VOUT+.n17 GNDA 0.287033f
C2311 VOUT+.n18 GNDA 0.059841f
C2312 VOUT+.t9 GNDA 0.04706f
C2313 VOUT+.t11 GNDA 0.04706f
C2314 VOUT+.n19 GNDA 0.096425f
C2315 VOUT+.n20 GNDA 0.282016f
C2316 VOUT+.n21 GNDA 0.059841f
C2317 VOUT+.t10 GNDA 0.04706f
C2318 VOUT+.t14 GNDA 0.04706f
C2319 VOUT+.n22 GNDA 0.096425f
C2320 VOUT+.n23 GNDA 0.282016f
C2321 VOUT+.n24 GNDA 0.03392f
C2322 VOUT+.n25 GNDA 0.03392f
C2323 VOUT+.t7 GNDA 0.04706f
C2324 VOUT+.t15 GNDA 0.04706f
C2325 VOUT+.n26 GNDA 0.096425f
C2326 VOUT+.n27 GNDA 0.282016f
C2327 VOUT+.n28 GNDA 0.03392f
C2328 VOUT+.n29 GNDA 0.049451f
C2329 VOUT+.n30 GNDA 0.202651f
C2330 VOUT+.t101 GNDA 0.31373f
C2331 VOUT+.t108 GNDA 0.319074f
C2332 VOUT+.t149 GNDA 0.31373f
C2333 VOUT+.n31 GNDA 0.210346f
C2334 VOUT+.n32 GNDA 0.137257f
C2335 VOUT+.t48 GNDA 0.318405f
C2336 VOUT+.t92 GNDA 0.318405f
C2337 VOUT+.t42 GNDA 0.318405f
C2338 VOUT+.t130 GNDA 0.318405f
C2339 VOUT+.t84 GNDA 0.318405f
C2340 VOUT+.t125 GNDA 0.318405f
C2341 VOUT+.t74 GNDA 0.318405f
C2342 VOUT+.t23 GNDA 0.318405f
C2343 VOUT+.t64 GNDA 0.318405f
C2344 VOUT+.t150 GNDA 0.318405f
C2345 VOUT+.t88 GNDA 0.31373f
C2346 VOUT+.n33 GNDA 0.211015f
C2347 VOUT+.t51 GNDA 0.31373f
C2348 VOUT+.n34 GNDA 0.269839f
C2349 VOUT+.t137 GNDA 0.31373f
C2350 VOUT+.n35 GNDA 0.269839f
C2351 VOUT+.t106 GNDA 0.31373f
C2352 VOUT+.n36 GNDA 0.269839f
C2353 VOUT+.t75 GNDA 0.31373f
C2354 VOUT+.n37 GNDA 0.269839f
C2355 VOUT+.t25 GNDA 0.31373f
C2356 VOUT+.n38 GNDA 0.269839f
C2357 VOUT+.t128 GNDA 0.31373f
C2358 VOUT+.n39 GNDA 0.269839f
C2359 VOUT+.t90 GNDA 0.31373f
C2360 VOUT+.n40 GNDA 0.269839f
C2361 VOUT+.t54 GNDA 0.31373f
C2362 VOUT+.n41 GNDA 0.269839f
C2363 VOUT+.t140 GNDA 0.31373f
C2364 VOUT+.n42 GNDA 0.269839f
C2365 VOUT+.t110 GNDA 0.31373f
C2366 VOUT+.t28 GNDA 0.319074f
C2367 VOUT+.t79 GNDA 0.31373f
C2368 VOUT+.n43 GNDA 0.210346f
C2369 VOUT+.n44 GNDA 0.254906f
C2370 VOUT+.t24 GNDA 0.319074f
C2371 VOUT+.t113 GNDA 0.31373f
C2372 VOUT+.n45 GNDA 0.210346f
C2373 VOUT+.t78 GNDA 0.31373f
C2374 VOUT+.t129 GNDA 0.319074f
C2375 VOUT+.t38 GNDA 0.31373f
C2376 VOUT+.n46 GNDA 0.210346f
C2377 VOUT+.n47 GNDA 0.254906f
C2378 VOUT+.t61 GNDA 0.319074f
C2379 VOUT+.t147 GNDA 0.31373f
C2380 VOUT+.n48 GNDA 0.210346f
C2381 VOUT+.t117 GNDA 0.31373f
C2382 VOUT+.t32 GNDA 0.319074f
C2383 VOUT+.t83 GNDA 0.31373f
C2384 VOUT+.n49 GNDA 0.210346f
C2385 VOUT+.n50 GNDA 0.254906f
C2386 VOUT+.t100 GNDA 0.319074f
C2387 VOUT+.t47 GNDA 0.31373f
C2388 VOUT+.n51 GNDA 0.210346f
C2389 VOUT+.t153 GNDA 0.31373f
C2390 VOUT+.t71 GNDA 0.319074f
C2391 VOUT+.t123 GNDA 0.31373f
C2392 VOUT+.n52 GNDA 0.210346f
C2393 VOUT+.n53 GNDA 0.254906f
C2394 VOUT+.t69 GNDA 0.319074f
C2395 VOUT+.t154 GNDA 0.31373f
C2396 VOUT+.n54 GNDA 0.210346f
C2397 VOUT+.t124 GNDA 0.31373f
C2398 VOUT+.t35 GNDA 0.319074f
C2399 VOUT+.t86 GNDA 0.31373f
C2400 VOUT+.n55 GNDA 0.210346f
C2401 VOUT+.n56 GNDA 0.254906f
C2402 VOUT+.t96 GNDA 0.31373f
C2403 VOUT+.t85 GNDA 0.319074f
C2404 VOUT+.t57 GNDA 0.31373f
C2405 VOUT+.n57 GNDA 0.210346f
C2406 VOUT+.n58 GNDA 0.137257f
C2407 VOUT+.t132 GNDA 0.318405f
C2408 VOUT+.t115 GNDA 0.318405f
C2409 VOUT+.t131 GNDA 0.319074f
C2410 VOUT+.t104 GNDA 0.31373f
C2411 VOUT+.n59 GNDA 0.210346f
C2412 VOUT+.t73 GNDA 0.31373f
C2413 VOUT+.n60 GNDA 0.132355f
C2414 VOUT+.t146 GNDA 0.318405f
C2415 VOUT+.t31 GNDA 0.319074f
C2416 VOUT+.t138 GNDA 0.31373f
C2417 VOUT+.n61 GNDA 0.210346f
C2418 VOUT+.t107 GNDA 0.31373f
C2419 VOUT+.n62 GNDA 0.132355f
C2420 VOUT+.t46 GNDA 0.318405f
C2421 VOUT+.t62 GNDA 0.319074f
C2422 VOUT+.t41 GNDA 0.31373f
C2423 VOUT+.n63 GNDA 0.210346f
C2424 VOUT+.t143 GNDA 0.31373f
C2425 VOUT+.n64 GNDA 0.132355f
C2426 VOUT+.t87 GNDA 0.318405f
C2427 VOUT+.t114 GNDA 0.319074f
C2428 VOUT+.t21 GNDA 0.31373f
C2429 VOUT+.n65 GNDA 0.210346f
C2430 VOUT+.t126 GNDA 0.31373f
C2431 VOUT+.n66 GNDA 0.132355f
C2432 VOUT+.t65 GNDA 0.318405f
C2433 VOUT+.t26 GNDA 0.318667f
C2434 VOUT+.t102 GNDA 0.318405f
C2435 VOUT+.t59 GNDA 0.318667f
C2436 VOUT+.t134 GNDA 0.318405f
C2437 VOUT+.t37 GNDA 0.318667f
C2438 VOUT+.t120 GNDA 0.318405f
C2439 VOUT+.t81 GNDA 0.318667f
C2440 VOUT+.t155 GNDA 0.318405f
C2441 VOUT+.t119 GNDA 0.31373f
C2442 VOUT+.n67 GNDA 0.347256f
C2443 VOUT+.t82 GNDA 0.31373f
C2444 VOUT+.n68 GNDA 0.406081f
C2445 VOUT+.t97 GNDA 0.31373f
C2446 VOUT+.n69 GNDA 0.406081f
C2447 VOUT+.t63 GNDA 0.31373f
C2448 VOUT+.n70 GNDA 0.406081f
C2449 VOUT+.t27 GNDA 0.31373f
C2450 VOUT+.n71 GNDA 0.333566f
C2451 VOUT+.t45 GNDA 0.31373f
C2452 VOUT+.n72 GNDA 0.333566f
C2453 VOUT+.t144 GNDA 0.31373f
C2454 VOUT+.n73 GNDA 0.333566f
C2455 VOUT+.t112 GNDA 0.31373f
C2456 VOUT+.n74 GNDA 0.333566f
C2457 VOUT+.t76 GNDA 0.31373f
C2458 VOUT+.n75 GNDA 0.269839f
C2459 VOUT+.t93 GNDA 0.31373f
C2460 VOUT+.n76 GNDA 0.269839f
C2461 VOUT+.t56 GNDA 0.31373f
C2462 VOUT+.t40 GNDA 0.319074f
C2463 VOUT+.t19 GNDA 0.31373f
C2464 VOUT+.n77 GNDA 0.210346f
C2465 VOUT+.n78 GNDA 0.254906f
C2466 VOUT+.t34 GNDA 0.319074f
C2467 VOUT+.t52 GNDA 0.31373f
C2468 VOUT+.n79 GNDA 0.210346f
C2469 VOUT+.t156 GNDA 0.31373f
C2470 VOUT+.t136 GNDA 0.319074f
C2471 VOUT+.t121 GNDA 0.31373f
C2472 VOUT+.n80 GNDA 0.210346f
C2473 VOUT+.n81 GNDA 0.254906f
C2474 VOUT+.t70 GNDA 0.319074f
C2475 VOUT+.t89 GNDA 0.31373f
C2476 VOUT+.n82 GNDA 0.210346f
C2477 VOUT+.t50 GNDA 0.31373f
C2478 VOUT+.t36 GNDA 0.319074f
C2479 VOUT+.t151 GNDA 0.31373f
C2480 VOUT+.n83 GNDA 0.210346f
C2481 VOUT+.n84 GNDA 0.254906f
C2482 VOUT+.t95 GNDA 0.319074f
C2483 VOUT+.t43 GNDA 0.31373f
C2484 VOUT+.n85 GNDA 0.210346f
C2485 VOUT+.t145 GNDA 0.31373f
C2486 VOUT+.t66 GNDA 0.319074f
C2487 VOUT+.t118 GNDA 0.31373f
C2488 VOUT+.n86 GNDA 0.210346f
C2489 VOUT+.n87 GNDA 0.254906f
C2490 VOUT+.t55 GNDA 0.319074f
C2491 VOUT+.t141 GNDA 0.31373f
C2492 VOUT+.n88 GNDA 0.210346f
C2493 VOUT+.t111 GNDA 0.31373f
C2494 VOUT+.t29 GNDA 0.319074f
C2495 VOUT+.t80 GNDA 0.31373f
C2496 VOUT+.n89 GNDA 0.210346f
C2497 VOUT+.n90 GNDA 0.254906f
C2498 VOUT+.t91 GNDA 0.319074f
C2499 VOUT+.t39 GNDA 0.31373f
C2500 VOUT+.n91 GNDA 0.210346f
C2501 VOUT+.t139 GNDA 0.31373f
C2502 VOUT+.t58 GNDA 0.319074f
C2503 VOUT+.t109 GNDA 0.31373f
C2504 VOUT+.n92 GNDA 0.210346f
C2505 VOUT+.n93 GNDA 0.254906f
C2506 VOUT+.t49 GNDA 0.319074f
C2507 VOUT+.t135 GNDA 0.31373f
C2508 VOUT+.n94 GNDA 0.210346f
C2509 VOUT+.t103 GNDA 0.31373f
C2510 VOUT+.t20 GNDA 0.319074f
C2511 VOUT+.t72 GNDA 0.31373f
C2512 VOUT+.n95 GNDA 0.210346f
C2513 VOUT+.n96 GNDA 0.254906f
C2514 VOUT+.t148 GNDA 0.319074f
C2515 VOUT+.t99 GNDA 0.31373f
C2516 VOUT+.n97 GNDA 0.210346f
C2517 VOUT+.t68 GNDA 0.31373f
C2518 VOUT+.t122 GNDA 0.319074f
C2519 VOUT+.t33 GNDA 0.31373f
C2520 VOUT+.n98 GNDA 0.210346f
C2521 VOUT+.n99 GNDA 0.254906f
C2522 VOUT+.t44 GNDA 0.319074f
C2523 VOUT+.t133 GNDA 0.31373f
C2524 VOUT+.n100 GNDA 0.210346f
C2525 VOUT+.t98 GNDA 0.31373f
C2526 VOUT+.t152 GNDA 0.319074f
C2527 VOUT+.t67 GNDA 0.31373f
C2528 VOUT+.n101 GNDA 0.210346f
C2529 VOUT+.n102 GNDA 0.254906f
C2530 VOUT+.t142 GNDA 0.319074f
C2531 VOUT+.t94 GNDA 0.31373f
C2532 VOUT+.n103 GNDA 0.210346f
C2533 VOUT+.t60 GNDA 0.31373f
C2534 VOUT+.t116 GNDA 0.319074f
C2535 VOUT+.t30 GNDA 0.31373f
C2536 VOUT+.n104 GNDA 0.210346f
C2537 VOUT+.n105 GNDA 0.254906f
C2538 VOUT+.t77 GNDA 0.319074f
C2539 VOUT+.t127 GNDA 0.31373f
C2540 VOUT+.n106 GNDA 0.210346f
C2541 VOUT+.t22 GNDA 0.31373f
C2542 VOUT+.n107 GNDA 0.254906f
C2543 VOUT+.t53 GNDA 0.31373f
C2544 VOUT+.n108 GNDA 0.137257f
C2545 VOUT+.t105 GNDA 0.31373f
C2546 VOUT+.n109 GNDA 0.249491f
C2547 VOUT+.n110 GNDA 0.317475f
C2548 two_stage_opamp_dummy_magic_0.VD2.n0 GNDA 0.483909f
C2549 two_stage_opamp_dummy_magic_0.VD2.n1 GNDA 0.099935f
C2550 two_stage_opamp_dummy_magic_0.VD2.n2 GNDA 0.167505f
C2551 two_stage_opamp_dummy_magic_0.VD2.t3 GNDA 0.053331f
C2552 two_stage_opamp_dummy_magic_0.VD2.t2 GNDA 0.053331f
C2553 two_stage_opamp_dummy_magic_0.VD2.n3 GNDA 0.116042f
C2554 two_stage_opamp_dummy_magic_0.VD2.n4 GNDA 0.192793f
C2555 two_stage_opamp_dummy_magic_0.VD2.t7 GNDA 0.053331f
C2556 two_stage_opamp_dummy_magic_0.VD2.t11 GNDA 0.053331f
C2557 two_stage_opamp_dummy_magic_0.VD2.n5 GNDA 0.116042f
C2558 two_stage_opamp_dummy_magic_0.VD2.n6 GNDA 0.461069f
C2559 two_stage_opamp_dummy_magic_0.VD2.t6 GNDA 0.053331f
C2560 two_stage_opamp_dummy_magic_0.VD2.t5 GNDA 0.053331f
C2561 two_stage_opamp_dummy_magic_0.VD2.n7 GNDA 0.116042f
C2562 two_stage_opamp_dummy_magic_0.VD2.n8 GNDA 0.461069f
C2563 two_stage_opamp_dummy_magic_0.VD2.t12 GNDA 0.053331f
C2564 two_stage_opamp_dummy_magic_0.VD2.t13 GNDA 0.053331f
C2565 two_stage_opamp_dummy_magic_0.VD2.n9 GNDA 0.116042f
C2566 two_stage_opamp_dummy_magic_0.VD2.n10 GNDA 0.442486f
C2567 two_stage_opamp_dummy_magic_0.VD2.n11 GNDA 0.203944f
C2568 two_stage_opamp_dummy_magic_0.VD2.n12 GNDA 0.119128f
C2569 two_stage_opamp_dummy_magic_0.VD2.n13 GNDA 0.203944f
C2570 two_stage_opamp_dummy_magic_0.VD2.t20 GNDA 0.053331f
C2571 two_stage_opamp_dummy_magic_0.VD2.t8 GNDA 0.053331f
C2572 two_stage_opamp_dummy_magic_0.VD2.n14 GNDA 0.116042f
C2573 two_stage_opamp_dummy_magic_0.VD2.n15 GNDA 0.442486f
C2574 two_stage_opamp_dummy_magic_0.VD2.n16 GNDA 0.192793f
C2575 two_stage_opamp_dummy_magic_0.VD2.n17 GNDA 0.106662f
C2576 two_stage_opamp_dummy_magic_0.VD2.n18 GNDA 0.205342f
C2577 two_stage_opamp_dummy_magic_0.VD2.t15 GNDA 0.053331f
C2578 two_stage_opamp_dummy_magic_0.VD2.t17 GNDA 0.053331f
C2579 two_stage_opamp_dummy_magic_0.VD2.n19 GNDA 0.116042f
C2580 two_stage_opamp_dummy_magic_0.VD2.n20 GNDA 0.465721f
C2581 two_stage_opamp_dummy_magic_0.VD2.n21 GNDA 0.205342f
C2582 two_stage_opamp_dummy_magic_0.VD2.t4 GNDA 0.053331f
C2583 two_stage_opamp_dummy_magic_0.VD2.t21 GNDA 0.053331f
C2584 two_stage_opamp_dummy_magic_0.VD2.n22 GNDA 0.116042f
C2585 two_stage_opamp_dummy_magic_0.VD2.n23 GNDA 0.447102f
C2586 two_stage_opamp_dummy_magic_0.VD2.n24 GNDA 0.192793f
C2587 two_stage_opamp_dummy_magic_0.VD2.t18 GNDA 0.053331f
C2588 two_stage_opamp_dummy_magic_0.VD2.t9 GNDA 0.053331f
C2589 two_stage_opamp_dummy_magic_0.VD2.n25 GNDA 0.116042f
C2590 two_stage_opamp_dummy_magic_0.VD2.n26 GNDA 0.447102f
C2591 two_stage_opamp_dummy_magic_0.VD2.n27 GNDA 0.113419f
C2592 two_stage_opamp_dummy_magic_0.VD2.t19 GNDA 0.053331f
C2593 two_stage_opamp_dummy_magic_0.VD2.t16 GNDA 0.053331f
C2594 two_stage_opamp_dummy_magic_0.VD2.n28 GNDA 0.116042f
C2595 two_stage_opamp_dummy_magic_0.VD2.n29 GNDA 0.465721f
C2596 two_stage_opamp_dummy_magic_0.VD2.t10 GNDA 0.053331f
C2597 two_stage_opamp_dummy_magic_0.VD2.t14 GNDA 0.053331f
C2598 two_stage_opamp_dummy_magic_0.VD2.n30 GNDA 0.116042f
C2599 two_stage_opamp_dummy_magic_0.VD2.n31 GNDA 0.447102f
C2600 two_stage_opamp_dummy_magic_0.VD2.n32 GNDA 0.192793f
C2601 two_stage_opamp_dummy_magic_0.VD2.n33 GNDA 0.113419f
C2602 two_stage_opamp_dummy_magic_0.VD2.t1 GNDA 0.053331f
C2603 two_stage_opamp_dummy_magic_0.VD2.t0 GNDA 0.053331f
C2604 two_stage_opamp_dummy_magic_0.VD2.n34 GNDA 0.116042f
C2605 two_stage_opamp_dummy_magic_0.VD2.n35 GNDA 0.447102f
C2606 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 GNDA 0.016904f
C2607 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 GNDA 0.016904f
C2608 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 GNDA 0.034522f
C2609 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 GNDA 0.127376f
C2610 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 GNDA 0.016904f
C2611 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 GNDA 0.016904f
C2612 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 GNDA 0.034522f
C2613 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 GNDA 0.181646f
C2614 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 GNDA 0.016904f
C2615 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 GNDA 0.016904f
C2616 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 GNDA 0.034522f
C2617 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 GNDA 0.181646f
C2618 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 GNDA 0.089279f
C2619 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 GNDA 0.089279f
C2620 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 GNDA 0.016904f
C2621 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 GNDA 0.016904f
C2622 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 GNDA 0.034522f
C2623 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 GNDA 0.172887f
C2624 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 GNDA 0.095677f
C2625 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 GNDA 0.090409f
C2626 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 GNDA 0.081803f
C2627 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 GNDA 1.17373f
C2628 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 GNDA 0.025355f
C2629 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 GNDA 0.025355f
C2630 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 GNDA 0.055171f
C2631 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 GNDA 0.197605f
C2632 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 GNDA 0.045006f
C2633 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 GNDA 0.045006f
C2634 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 GNDA 0.045006f
C2635 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 GNDA 0.045006f
C2636 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 GNDA 0.045006f
C2637 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 GNDA 0.045006f
C2638 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 GNDA 0.045006f
C2639 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 GNDA 0.045006f
C2640 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 GNDA 0.045006f
C2641 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 GNDA 0.052529f
C2642 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 GNDA 0.049527f
C2643 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 GNDA 0.031061f
C2644 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 GNDA 0.031061f
C2645 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 GNDA 0.031061f
C2646 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 GNDA 0.031061f
C2647 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 GNDA 0.031061f
C2648 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 GNDA 0.031061f
C2649 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 GNDA 0.031061f
C2650 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 GNDA 0.027755f
C2651 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 GNDA 0.045006f
C2652 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 GNDA 0.045006f
C2653 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 GNDA 0.045006f
C2654 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 GNDA 0.045006f
C2655 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 GNDA 0.045006f
C2656 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 GNDA 0.045006f
C2657 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 GNDA 0.045006f
C2658 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 GNDA 0.045006f
C2659 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 GNDA 0.045006f
C2660 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 GNDA 0.052529f
C2661 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 GNDA 0.049527f
C2662 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 GNDA 0.031061f
C2663 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 GNDA 0.031061f
C2664 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 GNDA 0.031061f
C2665 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 GNDA 0.031061f
C2666 two_stage_opamp_dummy_magic_0.V_tail_gate.n30 GNDA 0.031061f
C2667 two_stage_opamp_dummy_magic_0.V_tail_gate.n31 GNDA 0.031061f
C2668 two_stage_opamp_dummy_magic_0.V_tail_gate.n32 GNDA 0.031061f
C2669 two_stage_opamp_dummy_magic_0.V_tail_gate.n33 GNDA 0.027755f
C2670 two_stage_opamp_dummy_magic_0.V_tail_gate.n34 GNDA 0.023496f
C2671 two_stage_opamp_dummy_magic_0.V_tail_gate.n35 GNDA 0.205386f
C2672 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 GNDA 0.025355f
C2673 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 GNDA 0.025355f
C2674 two_stage_opamp_dummy_magic_0.V_tail_gate.n36 GNDA 0.055171f
C2675 two_stage_opamp_dummy_magic_0.V_tail_gate.n37 GNDA 0.244733f
C2676 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 GNDA 0.22024f
C2677 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 GNDA 0.157793f
C2678 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 GNDA 0.179507f
C2679 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 GNDA 0.015426f
C2680 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 GNDA 0.145366f
C2681 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 GNDA 0.013038f
C2682 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 GNDA 0.020333f
C2683 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 GNDA 0.015865f
C2684 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 GNDA 0.014143f
C2685 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 GNDA 0.022295f
C2686 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 GNDA 0.014143f
C2687 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 GNDA 0.015865f
C2688 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 GNDA 0.015865f
C2689 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 GNDA 0.014143f
C2690 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 GNDA 0.013038f
C2691 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 GNDA 0.018611f
C2692 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 GNDA 0.022295f
C2693 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 GNDA 0.014862f
C2694 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 GNDA 0.014862f
C2695 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 GNDA 0.123409f
C2696 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 GNDA 0.156365f
C2697 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 GNDA 0.014862f
C2698 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 GNDA 0.123409f
C2699 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 GNDA 0.158799f
C2700 two_stage_opamp_dummy_magic_0.err_amp_mir.n22 GNDA 0.122069f
C2701 two_stage_opamp_dummy_magic_0.err_amp_mir.n23 GNDA 0.114677f
C2702 two_stage_opamp_dummy_magic_0.err_amp_mir.n24 GNDA 0.015426f
C2703 two_stage_opamp_dummy_magic_0.err_amp_mir.n25 GNDA 0.172193f
C2704 two_stage_opamp_dummy_magic_0.err_amp_mir.n26 GNDA 0.015426f
C2705 VDDA.n0 GNDA 0.062237f
C2706 VDDA.t375 GNDA 0.048142f
C2707 VDDA.t208 GNDA 0.048142f
C2708 VDDA.n1 GNDA 0.098479f
C2709 VDDA.n2 GNDA 0.36701f
C2710 VDDA.n3 GNDA 0.095402f
C2711 VDDA.t106 GNDA 0.171248f
C2712 VDDA.t163 GNDA 0.171248f
C2713 VDDA.t161 GNDA 0.084283f
C2714 VDDA.n4 GNDA 0.153433f
C2715 VDDA.n5 GNDA 0.05548f
C2716 VDDA.n6 GNDA 0.062237f
C2717 VDDA.t290 GNDA 0.048142f
C2718 VDDA.t280 GNDA 0.048142f
C2719 VDDA.n7 GNDA 0.098479f
C2720 VDDA.n8 GNDA 0.36701f
C2721 VDDA.n9 GNDA 0.05548f
C2722 VDDA.n10 GNDA 0.05548f
C2723 VDDA.t30 GNDA 0.048142f
C2724 VDDA.t466 GNDA 0.048142f
C2725 VDDA.n11 GNDA 0.098479f
C2726 VDDA.n12 GNDA 0.36701f
C2727 VDDA.n13 GNDA 0.062237f
C2728 VDDA.t366 GNDA 0.048142f
C2729 VDDA.t427 GNDA 0.048142f
C2730 VDDA.n14 GNDA 0.098479f
C2731 VDDA.n15 GNDA 0.36701f
C2732 VDDA.n16 GNDA 0.062237f
C2733 VDDA.n17 GNDA 0.094461f
C2734 VDDA.t216 GNDA 0.048142f
C2735 VDDA.t468 GNDA 0.048142f
C2736 VDDA.n18 GNDA 0.098479f
C2737 VDDA.n19 GNDA 0.36701f
C2738 VDDA.n20 GNDA 0.095402f
C2739 VDDA.n21 GNDA 0.149207f
C2740 VDDA.n22 GNDA 0.496775f
C2741 VDDA.t162 GNDA 0.410358f
C2742 VDDA.t215 GNDA 0.321864f
C2743 VDDA.t467 GNDA 0.321864f
C2744 VDDA.t365 GNDA 0.321864f
C2745 VDDA.t426 GNDA 0.321864f
C2746 VDDA.t29 GNDA 0.321864f
C2747 VDDA.t465 GNDA 0.321864f
C2748 VDDA.t289 GNDA 0.321864f
C2749 VDDA.t279 GNDA 0.321864f
C2750 VDDA.t374 GNDA 0.321864f
C2751 VDDA.t207 GNDA 0.321864f
C2752 VDDA.t105 GNDA 0.410358f
C2753 VDDA.n23 GNDA 0.496775f
C2754 VDDA.n24 GNDA 0.149207f
C2755 VDDA.t104 GNDA 0.080156f
C2756 VDDA.n25 GNDA 0.149354f
C2757 VDDA.n26 GNDA 0.046618f
C2758 VDDA.n27 GNDA 0.050865f
C2759 VDDA.n28 GNDA 0.050865f
C2760 VDDA.t332 GNDA 0.041265f
C2761 VDDA.t341 GNDA 0.041265f
C2762 VDDA.n29 GNDA 0.088257f
C2763 VDDA.n30 GNDA 0.307499f
C2764 VDDA.n31 GNDA 0.088195f
C2765 VDDA.t28 GNDA 0.041265f
C2766 VDDA.t6 GNDA 0.041265f
C2767 VDDA.n32 GNDA 0.088257f
C2768 VDDA.n33 GNDA 0.299686f
C2769 VDDA.n34 GNDA 0.088195f
C2770 VDDA.t240 GNDA 0.041265f
C2771 VDDA.t223 GNDA 0.041265f
C2772 VDDA.n35 GNDA 0.088257f
C2773 VDDA.n36 GNDA 0.299686f
C2774 VDDA.n37 GNDA 0.050865f
C2775 VDDA.n38 GNDA 0.050865f
C2776 VDDA.t16 GNDA 0.041265f
C2777 VDDA.t431 GNDA 0.041265f
C2778 VDDA.n39 GNDA 0.088257f
C2779 VDDA.n40 GNDA 0.299686f
C2780 VDDA.n41 GNDA 0.050865f
C2781 VDDA.t364 GNDA 0.041265f
C2782 VDDA.t429 GNDA 0.041265f
C2783 VDDA.n42 GNDA 0.088257f
C2784 VDDA.n43 GNDA 0.299686f
C2785 VDDA.n44 GNDA 0.088195f
C2786 VDDA.t430 GNDA 0.041265f
C2787 VDDA.t333 GNDA 0.041265f
C2788 VDDA.n45 GNDA 0.088257f
C2789 VDDA.n46 GNDA 0.303593f
C2790 VDDA.n47 GNDA 0.187327f
C2791 VDDA.t192 GNDA 0.040179f
C2792 VDDA.n48 GNDA 0.158607f
C2793 VDDA.n49 GNDA 0.241742f
C2794 VDDA.t206 GNDA 0.098145f
C2795 VDDA.t194 GNDA 0.098145f
C2796 VDDA.n50 GNDA 0.285942f
C2797 VDDA.t193 GNDA 0.244509f
C2798 VDDA.t222 GNDA 0.181564f
C2799 VDDA.t428 GNDA 0.181564f
C2800 VDDA.t80 GNDA 0.181564f
C2801 VDDA.t363 GNDA 0.181564f
C2802 VDDA.t221 GNDA 0.181564f
C2803 VDDA.t281 GNDA 0.181564f
C2804 VDDA.t78 GNDA 0.181564f
C2805 VDDA.t36 GNDA 0.181564f
C2806 VDDA.t79 GNDA 0.181564f
C2807 VDDA.t62 GNDA 0.181564f
C2808 VDDA.t205 GNDA 0.244509f
C2809 VDDA.n51 GNDA 0.285942f
C2810 VDDA.n52 GNDA 0.241742f
C2811 VDDA.t204 GNDA 0.040179f
C2812 VDDA.n53 GNDA 0.10897f
C2813 VDDA.n54 GNDA 0.214061f
C2814 VDDA.n55 GNDA 0.271947f
C2815 VDDA.t176 GNDA 0.01955f
C2816 VDDA.n56 GNDA 0.15287f
C2817 VDDA.n57 GNDA 0.189129f
C2818 VDDA.t178 GNDA 0.02506f
C2819 VDDA.n58 GNDA 0.077586f
C2820 VDDA.t177 GNDA 0.102989f
C2821 VDDA.t416 GNDA 0.068086f
C2822 VDDA.t450 GNDA 0.068086f
C2823 VDDA.t71 GNDA 0.068086f
C2824 VDDA.t31 GNDA 0.068086f
C2825 VDDA.t5 GNDA 0.068086f
C2826 VDDA.t230 GNDA 0.068086f
C2827 VDDA.t336 GNDA 0.068086f
C2828 VDDA.t237 GNDA 0.068086f
C2829 VDDA.t214 GNDA 0.068086f
C2830 VDDA.t292 GNDA 0.068086f
C2831 VDDA.t165 GNDA 0.102989f
C2832 VDDA.t166 GNDA 0.02506f
C2833 VDDA.n59 GNDA 0.077586f
C2834 VDDA.n60 GNDA 0.189129f
C2835 VDDA.t164 GNDA 0.01955f
C2836 VDDA.n61 GNDA 0.103396f
C2837 VDDA.n62 GNDA 0.24612f
C2838 VDDA.n63 GNDA 0.153822f
C2839 VDDA.n64 GNDA 0.06887f
C2840 VDDA.t324 GNDA 0.082529f
C2841 VDDA.t64 GNDA 0.082529f
C2842 VDDA.n65 GNDA 0.169102f
C2843 VDDA.n66 GNDA 0.538686f
C2844 VDDA.n67 GNDA 0.113258f
C2845 VDDA.t94 GNDA 0.290441f
C2846 VDDA.t203 GNDA 0.290441f
C2847 VDDA.t201 GNDA 0.10013f
C2848 VDDA.n68 GNDA 0.178206f
C2849 VDDA.n69 GNDA 0.063763f
C2850 VDDA.n70 GNDA 0.06887f
C2851 VDDA.t322 GNDA 0.082529f
C2852 VDDA.t283 GNDA 0.082529f
C2853 VDDA.n71 GNDA 0.169102f
C2854 VDDA.n72 GNDA 0.538686f
C2855 VDDA.n73 GNDA 0.063763f
C2856 VDDA.n74 GNDA 0.063763f
C2857 VDDA.t55 GNDA 0.082529f
C2858 VDDA.t49 GNDA 0.082529f
C2859 VDDA.n75 GNDA 0.169102f
C2860 VDDA.n76 GNDA 0.538686f
C2861 VDDA.n77 GNDA 0.06887f
C2862 VDDA.t326 GNDA 0.082529f
C2863 VDDA.t51 GNDA 0.082529f
C2864 VDDA.n78 GNDA 0.169102f
C2865 VDDA.n79 GNDA 0.538686f
C2866 VDDA.n80 GNDA 0.06887f
C2867 VDDA.n81 GNDA 0.098987f
C2868 VDDA.t362 GNDA 0.082529f
C2869 VDDA.t239 GNDA 0.082529f
C2870 VDDA.n82 GNDA 0.169102f
C2871 VDDA.n83 GNDA 0.538686f
C2872 VDDA.n84 GNDA 0.113258f
C2873 VDDA.n85 GNDA 0.21563f
C2874 VDDA.n86 GNDA 0.836808f
C2875 VDDA.t202 GNDA 0.629245f
C2876 VDDA.t361 GNDA 0.484171f
C2877 VDDA.t238 GNDA 0.484171f
C2878 VDDA.t325 GNDA 0.484171f
C2879 VDDA.t50 GNDA 0.484171f
C2880 VDDA.t54 GNDA 0.484171f
C2881 VDDA.t48 GNDA 0.484171f
C2882 VDDA.t321 GNDA 0.484171f
C2883 VDDA.t282 GNDA 0.484171f
C2884 VDDA.t323 GNDA 0.484171f
C2885 VDDA.t63 GNDA 0.484171f
C2886 VDDA.t93 GNDA 0.629245f
C2887 VDDA.n87 GNDA 0.836808f
C2888 VDDA.n88 GNDA 0.21563f
C2889 VDDA.t92 GNDA 0.10013f
C2890 VDDA.n89 GNDA 0.174686f
C2891 VDDA.n90 GNDA 0.048079f
C2892 VDDA.n91 GNDA 0.045816f
C2893 VDDA.t149 GNDA 0.01955f
C2894 VDDA.n92 GNDA 0.08669f
C2895 VDDA.t139 GNDA 0.02506f
C2896 VDDA.n93 GNDA 0.078371f
C2897 VDDA.n94 GNDA 0.045816f
C2898 VDDA.n95 GNDA 0.045816f
C2899 VDDA.n96 GNDA 0.045816f
C2900 VDDA.n97 GNDA 0.045816f
C2901 VDDA.n98 GNDA 0.014013f
C2902 VDDA.n99 GNDA 0.146069f
C2903 VDDA.n100 GNDA 0.075749f
C2904 VDDA.n101 GNDA 0.014013f
C2905 VDDA.n102 GNDA 0.146069f
C2906 VDDA.n103 GNDA 0.045816f
C2907 VDDA.n104 GNDA 0.045816f
C2908 VDDA.n105 GNDA 0.014013f
C2909 VDDA.n106 GNDA 0.146069f
C2910 VDDA.n107 GNDA 0.045816f
C2911 VDDA.n108 GNDA 0.014013f
C2912 VDDA.n109 GNDA 0.146069f
C2913 VDDA.n110 GNDA 0.045816f
C2914 VDDA.n111 GNDA 0.045816f
C2915 VDDA.n112 GNDA 0.014013f
C2916 VDDA.n113 GNDA 0.146069f
C2917 VDDA.n114 GNDA 0.045816f
C2918 VDDA.n115 GNDA 0.014013f
C2919 VDDA.n116 GNDA 0.146069f
C2920 VDDA.n117 GNDA 0.045816f
C2921 VDDA.n118 GNDA 0.045816f
C2922 VDDA.n119 GNDA 0.014013f
C2923 VDDA.n120 GNDA 0.146069f
C2924 VDDA.n121 GNDA 0.045816f
C2925 VDDA.n122 GNDA 0.014013f
C2926 VDDA.n123 GNDA 0.146069f
C2927 VDDA.n124 GNDA 0.045816f
C2928 VDDA.n125 GNDA 0.045816f
C2929 VDDA.n126 GNDA 0.014013f
C2930 VDDA.n127 GNDA 0.146069f
C2931 VDDA.n128 GNDA 0.045816f
C2932 VDDA.n129 GNDA 0.014013f
C2933 VDDA.n130 GNDA 0.146069f
C2934 VDDA.n131 GNDA 0.075749f
C2935 VDDA.t137 GNDA 0.01955f
C2936 VDDA.n132 GNDA 0.08669f
C2937 VDDA.n133 GNDA 0.080922f
C2938 VDDA.n134 GNDA 0.077586f
C2939 VDDA.t138 GNDA 0.102989f
C2940 VDDA.t235 GNDA 0.068086f
C2941 VDDA.t293 GNDA 0.068086f
C2942 VDDA.t444 GNDA 0.068086f
C2943 VDDA.t339 GNDA 0.068086f
C2944 VDDA.t459 GNDA 0.068086f
C2945 VDDA.t277 GNDA 0.068086f
C2946 VDDA.t297 GNDA 0.068086f
C2947 VDDA.t231 GNDA 0.068086f
C2948 VDDA.t24 GNDA 0.068086f
C2949 VDDA.t424 GNDA 0.068086f
C2950 VDDA.t422 GNDA 0.068086f
C2951 VDDA.t453 GNDA 0.068086f
C2952 VDDA.t295 GNDA 0.068086f
C2953 VDDA.t266 GNDA 0.068086f
C2954 VDDA.t264 GNDA 0.068086f
C2955 VDDA.t446 GNDA 0.068086f
C2956 VDDA.t26 GNDA 0.068086f
C2957 VDDA.t0 GNDA 0.068086f
C2958 VDDA.t76 GNDA 0.068086f
C2959 VDDA.t268 GNDA 0.068086f
C2960 VDDA.t150 GNDA 0.102989f
C2961 VDDA.t151 GNDA 0.02506f
C2962 VDDA.n135 GNDA 0.077586f
C2963 VDDA.n136 GNDA 0.07729f
C2964 VDDA.n137 GNDA 0.102211f
C2965 VDDA.n138 GNDA 0.102474f
C2966 VDDA.n139 GNDA 0.262844f
C2967 VDDA.n140 GNDA 0.238521f
C2968 VDDA.n141 GNDA 0.062237f
C2969 VDDA.t449 GNDA 0.048142f
C2970 VDDA.t347 GNDA 0.048142f
C2971 VDDA.n142 GNDA 0.098479f
C2972 VDDA.n143 GNDA 0.36701f
C2973 VDDA.n144 GNDA 0.095402f
C2974 VDDA.t181 GNDA 0.171248f
C2975 VDDA.t179 GNDA 0.084283f
C2976 VDDA.n145 GNDA 0.153433f
C2977 VDDA.n146 GNDA 0.05548f
C2978 VDDA.n147 GNDA 0.062237f
C2979 VDDA.t302 GNDA 0.048142f
C2980 VDDA.t345 GNDA 0.048142f
C2981 VDDA.n148 GNDA 0.098479f
C2982 VDDA.n149 GNDA 0.36701f
C2983 VDDA.n150 GNDA 0.05548f
C2984 VDDA.n151 GNDA 0.05548f
C2985 VDDA.t360 GNDA 0.048142f
C2986 VDDA.t4 GNDA 0.048142f
C2987 VDDA.n152 GNDA 0.098479f
C2988 VDDA.n153 GNDA 0.36701f
C2989 VDDA.n154 GNDA 0.062237f
C2990 VDDA.t368 GNDA 0.048142f
C2991 VDDA.t8 GNDA 0.048142f
C2992 VDDA.n155 GNDA 0.098479f
C2993 VDDA.n156 GNDA 0.36701f
C2994 VDDA.n157 GNDA 0.062237f
C2995 VDDA.n158 GNDA 0.094461f
C2996 VDDA.t343 GNDA 0.048142f
C2997 VDDA.t462 GNDA 0.048142f
C2998 VDDA.n159 GNDA 0.098479f
C2999 VDDA.n160 GNDA 0.36701f
C3000 VDDA.n161 GNDA 0.095402f
C3001 VDDA.n162 GNDA 0.149207f
C3002 VDDA.n163 GNDA 0.496775f
C3003 VDDA.t180 GNDA 0.410358f
C3004 VDDA.t461 GNDA 0.321864f
C3005 VDDA.t342 GNDA 0.321864f
C3006 VDDA.t7 GNDA 0.321864f
C3007 VDDA.t367 GNDA 0.321864f
C3008 VDDA.t3 GNDA 0.321864f
C3009 VDDA.t359 GNDA 0.321864f
C3010 VDDA.t344 GNDA 0.321864f
C3011 VDDA.t301 GNDA 0.321864f
C3012 VDDA.t346 GNDA 0.321864f
C3013 VDDA.t448 GNDA 0.321864f
C3014 VDDA.t108 GNDA 0.410358f
C3015 VDDA.t109 GNDA 0.171248f
C3016 VDDA.n164 GNDA 0.496775f
C3017 VDDA.n165 GNDA 0.149207f
C3018 VDDA.t107 GNDA 0.080156f
C3019 VDDA.n166 GNDA 0.149354f
C3020 VDDA.n167 GNDA 0.045931f
C3021 VDDA.n168 GNDA 0.050865f
C3022 VDDA.n169 GNDA 0.050865f
C3023 VDDA.t377 GNDA 0.041265f
C3024 VDDA.t335 GNDA 0.041265f
C3025 VDDA.n170 GNDA 0.088257f
C3026 VDDA.n171 GNDA 0.307499f
C3027 VDDA.n172 GNDA 0.088195f
C3028 VDDA.t390 GNDA 0.041265f
C3029 VDDA.t397 GNDA 0.041265f
C3030 VDDA.n173 GNDA 0.088257f
C3031 VDDA.n174 GNDA 0.299686f
C3032 VDDA.n175 GNDA 0.088195f
C3033 VDDA.t382 GNDA 0.041265f
C3034 VDDA.t412 GNDA 0.041265f
C3035 VDDA.n176 GNDA 0.088257f
C3036 VDDA.n177 GNDA 0.299686f
C3037 VDDA.n178 GNDA 0.050865f
C3038 VDDA.n179 GNDA 0.050865f
C3039 VDDA.t386 GNDA 0.041265f
C3040 VDDA.t378 GNDA 0.041265f
C3041 VDDA.n180 GNDA 0.088257f
C3042 VDDA.n181 GNDA 0.299686f
C3043 VDDA.n182 GNDA 0.050865f
C3044 VDDA.t391 GNDA 0.041265f
C3045 VDDA.t376 GNDA 0.041265f
C3046 VDDA.n183 GNDA 0.088257f
C3047 VDDA.n184 GNDA 0.299686f
C3048 VDDA.n185 GNDA 0.088195f
C3049 VDDA.t334 GNDA 0.041265f
C3050 VDDA.t408 GNDA 0.041265f
C3051 VDDA.n186 GNDA 0.088257f
C3052 VDDA.n187 GNDA 0.303593f
C3053 VDDA.n188 GNDA 0.187327f
C3054 VDDA.t122 GNDA 0.040179f
C3055 VDDA.n189 GNDA 0.158607f
C3056 VDDA.n190 GNDA 0.241742f
C3057 VDDA.t124 GNDA 0.098145f
C3058 VDDA.n191 GNDA 0.285942f
C3059 VDDA.t123 GNDA 0.244509f
C3060 VDDA.t409 GNDA 0.181564f
C3061 VDDA.t394 GNDA 0.181564f
C3062 VDDA.t383 GNDA 0.181564f
C3063 VDDA.t402 GNDA 0.181564f
C3064 VDDA.t387 GNDA 0.181564f
C3065 VDDA.t405 GNDA 0.181564f
C3066 VDDA.t415 GNDA 0.181564f
C3067 VDDA.t398 GNDA 0.181564f
C3068 VDDA.t379 GNDA 0.181564f
C3069 VDDA.t399 GNDA 0.181564f
C3070 VDDA.t99 GNDA 0.244509f
C3071 VDDA.t100 GNDA 0.098145f
C3072 VDDA.n192 GNDA 0.285942f
C3073 VDDA.n193 GNDA 0.241742f
C3074 VDDA.t98 GNDA 0.040179f
C3075 VDDA.n194 GNDA 0.10897f
C3076 VDDA.n195 GNDA 0.214061f
C3077 VDDA.n196 GNDA 0.271947f
C3078 VDDA.t158 GNDA 0.01955f
C3079 VDDA.n197 GNDA 0.15287f
C3080 VDDA.n198 GNDA 0.189129f
C3081 VDDA.t175 GNDA 0.02506f
C3082 VDDA.t160 GNDA 0.02506f
C3083 VDDA.n199 GNDA 0.077586f
C3084 VDDA.t159 GNDA 0.102989f
C3085 VDDA.t53 GNDA 0.068086f
C3086 VDDA.t419 GNDA 0.068086f
C3087 VDDA.t291 GNDA 0.068086f
C3088 VDDA.t209 GNDA 0.068086f
C3089 VDDA.t288 GNDA 0.068086f
C3090 VDDA.t17 GNDA 0.068086f
C3091 VDDA.t433 GNDA 0.068086f
C3092 VDDA.t432 GNDA 0.068086f
C3093 VDDA.t2 GNDA 0.068086f
C3094 VDDA.t270 GNDA 0.068086f
C3095 VDDA.t174 GNDA 0.102989f
C3096 VDDA.n200 GNDA 0.077586f
C3097 VDDA.n201 GNDA 0.189129f
C3098 VDDA.t173 GNDA 0.01955f
C3099 VDDA.n202 GNDA 0.103396f
C3100 VDDA.n203 GNDA 0.24612f
C3101 VDDA.n204 GNDA 0.153822f
C3102 VDDA.n205 GNDA 0.06887f
C3103 VDDA.t404 GNDA 0.082529f
C3104 VDDA.t385 GNDA 0.082529f
C3105 VDDA.n206 GNDA 0.169102f
C3106 VDDA.n207 GNDA 0.538686f
C3107 VDDA.n208 GNDA 0.113258f
C3108 VDDA.t133 GNDA 0.290441f
C3109 VDDA.t131 GNDA 0.10013f
C3110 VDDA.n209 GNDA 0.178206f
C3111 VDDA.n210 GNDA 0.063763f
C3112 VDDA.n211 GNDA 0.06887f
C3113 VDDA.t401 GNDA 0.082529f
C3114 VDDA.t381 GNDA 0.082529f
C3115 VDDA.n212 GNDA 0.169102f
C3116 VDDA.n213 GNDA 0.538686f
C3117 VDDA.n214 GNDA 0.063763f
C3118 VDDA.n215 GNDA 0.063763f
C3119 VDDA.t411 GNDA 0.082529f
C3120 VDDA.t393 GNDA 0.082529f
C3121 VDDA.n216 GNDA 0.169102f
C3122 VDDA.n217 GNDA 0.538686f
C3123 VDDA.n218 GNDA 0.06887f
C3124 VDDA.t407 GNDA 0.082529f
C3125 VDDA.t389 GNDA 0.082529f
C3126 VDDA.n219 GNDA 0.169102f
C3127 VDDA.n220 GNDA 0.538686f
C3128 VDDA.n221 GNDA 0.06887f
C3129 VDDA.n222 GNDA 0.098987f
C3130 VDDA.t396 GNDA 0.082529f
C3131 VDDA.t414 GNDA 0.082529f
C3132 VDDA.n223 GNDA 0.169102f
C3133 VDDA.n224 GNDA 0.538686f
C3134 VDDA.n225 GNDA 0.113258f
C3135 VDDA.n226 GNDA 0.21563f
C3136 VDDA.n227 GNDA 0.836808f
C3137 VDDA.t132 GNDA 0.629245f
C3138 VDDA.t413 GNDA 0.484171f
C3139 VDDA.t395 GNDA 0.484171f
C3140 VDDA.t388 GNDA 0.484171f
C3141 VDDA.t406 GNDA 0.484171f
C3142 VDDA.t392 GNDA 0.484171f
C3143 VDDA.t410 GNDA 0.484171f
C3144 VDDA.t380 GNDA 0.484171f
C3145 VDDA.t400 GNDA 0.484171f
C3146 VDDA.t384 GNDA 0.484171f
C3147 VDDA.t403 GNDA 0.484171f
C3148 VDDA.t111 GNDA 0.629245f
C3149 VDDA.t112 GNDA 0.290441f
C3150 VDDA.n228 GNDA 0.836808f
C3151 VDDA.n229 GNDA 0.21563f
C3152 VDDA.t110 GNDA 0.10013f
C3153 VDDA.n230 GNDA 0.174686f
C3154 VDDA.n231 GNDA 0.079138f
C3155 VDDA.n232 GNDA 0.268236f
C3156 VDDA.n233 GNDA 0.237833f
C3157 VDDA.n234 GNDA 0.3443f
C3158 VDDA.t242 GNDA 0.024759f
C3159 VDDA.t184 GNDA 0.024759f
C3160 VDDA.n235 GNDA 0.056001f
C3161 VDDA.n236 GNDA 0.223295f
C3162 VDDA.t167 GNDA 0.051743f
C3163 VDDA.t185 GNDA 0.089365f
C3164 VDDA.t182 GNDA 0.051743f
C3165 VDDA.n237 GNDA 0.136986f
C3166 VDDA.n238 GNDA 0.269067f
C3167 VDDA.t183 GNDA 0.239544f
C3168 VDDA.t241 GNDA 0.181564f
C3169 VDDA.t168 GNDA 0.239544f
C3170 VDDA.t169 GNDA 0.089365f
C3171 VDDA.n239 GNDA 0.269067f
C3172 VDDA.n240 GNDA 0.135683f
C3173 VDDA.n241 GNDA 0.078512f
C3174 VDDA.n242 GNDA 0.139761f
C3175 VDDA.n243 GNDA 0.345425f
C3176 VDDA.t119 GNDA 0.085252f
C3177 VDDA.t15 GNDA 0.048142f
C3178 VDDA.n244 GNDA 0.120937f
C3179 VDDA.t200 GNDA 0.21939f
C3180 VDDA.t198 GNDA 0.085252f
C3181 VDDA.n245 GNDA 0.180071f
C3182 VDDA.n246 GNDA 0.547741f
C3183 VDDA.t199 GNDA 0.410358f
C3184 VDDA.t14 GNDA 0.321864f
C3185 VDDA.t120 GNDA 0.410358f
C3186 VDDA.t121 GNDA 0.171248f
C3187 VDDA.n247 GNDA 0.547741f
C3188 VDDA.n248 GNDA 0.178768f
C3189 VDDA.n249 GNDA 0.078512f
C3190 VDDA.n250 GNDA 0.368762f
C3191 VDDA.n251 GNDA 7.60041f
C3192 VDDA.t331 GNDA 0.768896f
C3193 VDDA.t306 GNDA 0.771683f
C3194 VDDA.t41 GNDA 0.730418f
C3195 VDDA.t35 GNDA 0.768896f
C3196 VDDA.t350 GNDA 0.771683f
C3197 VDDA.t328 GNDA 0.730418f
C3198 VDDA.t327 GNDA 0.768896f
C3199 VDDA.t371 GNDA 0.771683f
C3200 VDDA.t245 GNDA 0.730418f
C3201 VDDA.t247 GNDA 0.768896f
C3202 VDDA.t351 GNDA 0.771683f
C3203 VDDA.t83 GNDA 0.730418f
C3204 VDDA.t354 GNDA 0.768896f
C3205 VDDA.t11 GNDA 0.771683f
C3206 VDDA.t42 GNDA 0.730418f
C3207 VDDA.n252 GNDA 0.515392f
C3208 VDDA.t227 GNDA 0.410434f
C3209 VDDA.n253 GNDA 0.559212f
C3210 VDDA.t47 GNDA 0.410434f
C3211 VDDA.n254 GNDA 0.559212f
C3212 VDDA.t34 GNDA 0.410434f
C3213 VDDA.n255 GNDA 0.559212f
C3214 VDDA.t246 GNDA 0.410434f
C3215 VDDA.n256 GNDA 0.559212f
C3216 VDDA.t224 GNDA 0.719012f
C3217 VDDA.n257 GNDA 6.36261f
C3218 VDDA.t471 GNDA 1.74393f
C3219 VDDA.t469 GNDA 1.74081f
C3220 VDDA.n258 GNDA 0.372118f
C3221 VDDA.t472 GNDA 1.74104f
C3222 VDDA.n259 GNDA 0.236905f
C3223 VDDA.t470 GNDA 1.74104f
C3224 VDDA.n260 GNDA 0.373589f
C3225 VDDA.n261 GNDA 1.41074f
C3226 VDDA.n262 GNDA 0.053259f
C3227 VDDA.t234 GNDA 0.013755f
C3228 VDDA.t316 GNDA 0.013755f
C3229 VDDA.n263 GNDA 0.028091f
C3230 VDDA.n264 GNDA 0.208544f
C3231 VDDA.n265 GNDA 0.087156f
C3232 VDDA.t118 GNDA 0.050121f
C3233 VDDA.t142 GNDA 0.050121f
C3234 VDDA.n266 GNDA 0.087156f
C3235 VDDA.n267 GNDA 0.053259f
C3236 VDDA.t89 GNDA 0.013755f
C3237 VDDA.t70 GNDA 0.013755f
C3238 VDDA.n268 GNDA 0.028091f
C3239 VDDA.n269 GNDA 0.208544f
C3240 VDDA.n270 GNDA 0.087156f
C3241 VDDA.t97 GNDA 0.050121f
C3242 VDDA.t197 GNDA 0.050121f
C3243 VDDA.n271 GNDA 0.087156f
C3244 VDDA.n272 GNDA 0.053259f
C3245 VDDA.n273 GNDA 0.051227f
C3246 VDDA.n274 GNDA 0.053259f
C3247 VDDA.n275 GNDA 0.053259f
C3248 VDDA.t418 GNDA 0.013755f
C3249 VDDA.t61 GNDA 0.013755f
C3250 VDDA.n276 GNDA 0.028091f
C3251 VDDA.n277 GNDA 0.208544f
C3252 VDDA.n278 GNDA 0.051227f
C3253 VDDA.t370 GNDA 0.013755f
C3254 VDDA.t66 GNDA 0.013755f
C3255 VDDA.n279 GNDA 0.028091f
C3256 VDDA.n280 GNDA 0.208544f
C3257 VDDA.n281 GNDA 0.051227f
C3258 VDDA.n282 GNDA 0.051227f
C3259 VDDA.t349 GNDA 0.013755f
C3260 VDDA.t85 GNDA 0.013755f
C3261 VDDA.n283 GNDA 0.028091f
C3262 VDDA.n284 GNDA 0.208544f
C3263 VDDA.n285 GNDA 0.053259f
C3264 VDDA.t38 GNDA 0.013755f
C3265 VDDA.t59 GNDA 0.013755f
C3266 VDDA.n286 GNDA 0.028091f
C3267 VDDA.n287 GNDA 0.208544f
C3268 VDDA.n288 GNDA 0.053259f
C3269 VDDA.n289 GNDA 0.053259f
C3270 VDDA.t318 GNDA 0.013755f
C3271 VDDA.t285 GNDA 0.013755f
C3272 VDDA.n290 GNDA 0.028091f
C3273 VDDA.n291 GNDA 0.208544f
C3274 VDDA.n292 GNDA 0.051227f
C3275 VDDA.t87 GNDA 0.013755f
C3276 VDDA.t68 GNDA 0.013755f
C3277 VDDA.n293 GNDA 0.028091f
C3278 VDDA.n294 GNDA 0.208544f
C3279 VDDA.n295 GNDA 0.051227f
C3280 VDDA.n296 GNDA 0.051227f
C3281 VDDA.t13 GNDA 0.013755f
C3282 VDDA.t91 GNDA 0.013755f
C3283 VDDA.n297 GNDA 0.028091f
C3284 VDDA.n298 GNDA 0.208544f
C3285 VDDA.n299 GNDA 0.053259f
C3286 VDDA.t57 GNDA 0.013755f
C3287 VDDA.t287 GNDA 0.013755f
C3288 VDDA.n300 GNDA 0.028091f
C3289 VDDA.n301 GNDA 0.208544f
C3290 VDDA.n302 GNDA 0.085943f
C3291 VDDA.t195 GNDA 0.034862f
C3292 VDDA.n303 GNDA 0.114361f
C3293 VDDA.n304 GNDA 0.103683f
C3294 VDDA.n305 GNDA 0.147334f
C3295 VDDA.t196 GNDA 0.158795f
C3296 VDDA.t56 GNDA 0.115541f
C3297 VDDA.t286 GNDA 0.115541f
C3298 VDDA.t12 GNDA 0.115541f
C3299 VDDA.t90 GNDA 0.115541f
C3300 VDDA.t86 GNDA 0.115541f
C3301 VDDA.t67 GNDA 0.115541f
C3302 VDDA.t317 GNDA 0.115541f
C3303 VDDA.t284 GNDA 0.115541f
C3304 VDDA.t37 GNDA 0.115541f
C3305 VDDA.t58 GNDA 0.115541f
C3306 VDDA.t348 GNDA 0.115541f
C3307 VDDA.t84 GNDA 0.115541f
C3308 VDDA.t369 GNDA 0.115541f
C3309 VDDA.t65 GNDA 0.115541f
C3310 VDDA.t417 GNDA 0.115541f
C3311 VDDA.t60 GNDA 0.115541f
C3312 VDDA.t88 GNDA 0.115541f
C3313 VDDA.t69 GNDA 0.115541f
C3314 VDDA.t96 GNDA 0.161553f
C3315 VDDA.n306 GNDA 0.154205f
C3316 VDDA.n307 GNDA 0.103683f
C3317 VDDA.t95 GNDA 0.034862f
C3318 VDDA.n308 GNDA 0.110258f
C3319 VDDA.n309 GNDA 0.075301f
C3320 VDDA.n310 GNDA 0.053259f
C3321 VDDA.n311 GNDA 0.051227f
C3322 VDDA.n312 GNDA 0.053259f
C3323 VDDA.n313 GNDA 0.053259f
C3324 VDDA.t272 GNDA 0.013755f
C3325 VDDA.t464 GNDA 0.013755f
C3326 VDDA.n314 GNDA 0.028091f
C3327 VDDA.n315 GNDA 0.208544f
C3328 VDDA.n316 GNDA 0.051227f
C3329 VDDA.t373 GNDA 0.013755f
C3330 VDDA.t73 GNDA 0.013755f
C3331 VDDA.n317 GNDA 0.028091f
C3332 VDDA.n318 GNDA 0.208544f
C3333 VDDA.n319 GNDA 0.051227f
C3334 VDDA.n320 GNDA 0.051227f
C3335 VDDA.t421 GNDA 0.013755f
C3336 VDDA.t358 GNDA 0.013755f
C3337 VDDA.n321 GNDA 0.028091f
C3338 VDDA.n322 GNDA 0.208544f
C3339 VDDA.n323 GNDA 0.053259f
C3340 VDDA.t274 GNDA 0.013755f
C3341 VDDA.t452 GNDA 0.013755f
C3342 VDDA.n324 GNDA 0.028091f
C3343 VDDA.n325 GNDA 0.208544f
C3344 VDDA.n326 GNDA 0.053259f
C3345 VDDA.n327 GNDA 0.053259f
C3346 VDDA.t304 GNDA 0.013755f
C3347 VDDA.t255 GNDA 0.013755f
C3348 VDDA.n328 GNDA 0.028091f
C3349 VDDA.n329 GNDA 0.208544f
C3350 VDDA.n330 GNDA 0.051227f
C3351 VDDA.t19 GNDA 0.013755f
C3352 VDDA.t356 GNDA 0.013755f
C3353 VDDA.n331 GNDA 0.028091f
C3354 VDDA.n332 GNDA 0.208544f
C3355 VDDA.n333 GNDA 0.051227f
C3356 VDDA.n334 GNDA 0.051227f
C3357 VDDA.t75 GNDA 0.013755f
C3358 VDDA.t435 GNDA 0.013755f
C3359 VDDA.n335 GNDA 0.028091f
C3360 VDDA.n336 GNDA 0.208544f
C3361 VDDA.n337 GNDA 0.053259f
C3362 VDDA.t314 GNDA 0.013755f
C3363 VDDA.t253 GNDA 0.013755f
C3364 VDDA.n338 GNDA 0.028091f
C3365 VDDA.n339 GNDA 0.208544f
C3366 VDDA.n340 GNDA 0.053259f
C3367 VDDA.n341 GNDA 0.075301f
C3368 VDDA.t140 GNDA 0.034862f
C3369 VDDA.n342 GNDA 0.110258f
C3370 VDDA.n343 GNDA 0.103683f
C3371 VDDA.n344 GNDA 0.154205f
C3372 VDDA.t141 GNDA 0.161553f
C3373 VDDA.t313 GNDA 0.115541f
C3374 VDDA.t252 GNDA 0.115541f
C3375 VDDA.t74 GNDA 0.115541f
C3376 VDDA.t434 GNDA 0.115541f
C3377 VDDA.t18 GNDA 0.115541f
C3378 VDDA.t355 GNDA 0.115541f
C3379 VDDA.t303 GNDA 0.115541f
C3380 VDDA.t254 GNDA 0.115541f
C3381 VDDA.t273 GNDA 0.115541f
C3382 VDDA.t451 GNDA 0.115541f
C3383 VDDA.t420 GNDA 0.115541f
C3384 VDDA.t357 GNDA 0.115541f
C3385 VDDA.t372 GNDA 0.115541f
C3386 VDDA.t72 GNDA 0.115541f
C3387 VDDA.t271 GNDA 0.115541f
C3388 VDDA.t463 GNDA 0.115541f
C3389 VDDA.t233 GNDA 0.115541f
C3390 VDDA.t315 GNDA 0.115541f
C3391 VDDA.t117 GNDA 0.158795f
C3392 VDDA.n345 GNDA 0.147334f
C3393 VDDA.n346 GNDA 0.103683f
C3394 VDDA.t116 GNDA 0.034862f
C3395 VDDA.n347 GNDA 0.110258f
C3396 VDDA.n348 GNDA 0.210298f
C3397 VDDA.n349 GNDA 0.505979f
C3398 VDDA.t152 GNDA 0.028257f
C3399 VDDA.n350 GNDA 0.090199f
C3400 VDDA.n351 GNDA 0.131703f
C3401 VDDA.t191 GNDA 0.050121f
C3402 VDDA.t154 GNDA 0.050121f
C3403 VDDA.n352 GNDA 0.144756f
C3404 VDDA.t153 GNDA 0.151746f
C3405 VDDA.t305 GNDA 0.105912f
C3406 VDDA.t52 GNDA 0.105912f
C3407 VDDA.t190 GNDA 0.151746f
C3408 VDDA.n353 GNDA 0.144756f
C3409 VDDA.n354 GNDA 0.131703f
C3410 VDDA.t189 GNDA 0.028257f
C3411 VDDA.n355 GNDA 0.080154f
C3412 VDDA.n356 GNDA 0.123882f
C3413 VDDA.t145 GNDA 0.413323f
C3414 VDDA.t144 GNDA 0.541264f
C3415 VDDA.t39 GNDA 0.420899f
C3416 VDDA.t329 GNDA 0.420899f
C3417 VDDA.t307 GNDA 0.420899f
C3418 VDDA.t352 GNDA 0.420899f
C3419 VDDA.t248 GNDA 0.420899f
C3420 VDDA.t243 GNDA 0.420899f
C3421 VDDA.t81 GNDA 0.420899f
C3422 VDDA.t43 GNDA 0.420899f
C3423 VDDA.t9 GNDA 0.420899f
C3424 VDDA.t32 GNDA 0.420899f
C3425 VDDA.t225 GNDA 0.420899f
C3426 VDDA.t45 GNDA 0.420899f
C3427 VDDA.t228 GNDA 0.420899f
C3428 VDDA.t250 GNDA 0.420899f
C3429 VDDA.t311 GNDA 0.420899f
C3430 VDDA.t309 GNDA 0.420899f
C3431 VDDA.t187 GNDA 0.460565f
C3432 VDDA.t188 GNDA 0.14621f
C3433 VDDA.n357 GNDA 0.505586f
C3434 VDDA.t186 GNDA 0.198371f
C3435 VDDA.n358 GNDA 0.174104f
C3436 VDDA.n359 GNDA 0.07909f
C3437 VDDA.t310 GNDA 0.041265f
C3438 VDDA.t312 GNDA 0.041265f
C3439 VDDA.n360 GNDA 0.101576f
C3440 VDDA.n361 GNDA 0.31107f
C3441 VDDA.t251 GNDA 0.041265f
C3442 VDDA.t229 GNDA 0.041265f
C3443 VDDA.n362 GNDA 0.101576f
C3444 VDDA.n363 GNDA 0.31107f
C3445 VDDA.t46 GNDA 0.041265f
C3446 VDDA.t226 GNDA 0.041265f
C3447 VDDA.n364 GNDA 0.101576f
C3448 VDDA.n365 GNDA 0.31107f
C3449 VDDA.t33 GNDA 0.041265f
C3450 VDDA.t10 GNDA 0.041265f
C3451 VDDA.n366 GNDA 0.101576f
C3452 VDDA.n367 GNDA 0.31107f
C3453 VDDA.t44 GNDA 0.041265f
C3454 VDDA.t82 GNDA 0.041265f
C3455 VDDA.n368 GNDA 0.101576f
C3456 VDDA.n369 GNDA 0.31107f
C3457 VDDA.t244 GNDA 0.041265f
C3458 VDDA.t249 GNDA 0.041265f
C3459 VDDA.n370 GNDA 0.101576f
C3460 VDDA.n371 GNDA 0.31107f
C3461 VDDA.t353 GNDA 0.041265f
C3462 VDDA.t308 GNDA 0.041265f
C3463 VDDA.n372 GNDA 0.101576f
C3464 VDDA.n373 GNDA 0.31107f
C3465 VDDA.t330 GNDA 0.041265f
C3466 VDDA.t40 GNDA 0.041265f
C3467 VDDA.n374 GNDA 0.101576f
C3468 VDDA.n375 GNDA 0.31107f
C3469 VDDA.t143 GNDA 0.199384f
C3470 VDDA.n376 GNDA 0.176812f
C3471 VDDA.t276 GNDA 0.013755f
C3472 VDDA.t23 GNDA 0.013755f
C3473 VDDA.n377 GNDA 0.028091f
C3474 VDDA.n378 GNDA 0.100593f
C3475 VDDA.t128 GNDA 0.029712f
C3476 VDDA.n379 GNDA 0.08592f
C3477 VDDA.n380 GNDA 0.102404f
C3478 VDDA.t127 GNDA 0.050121f
C3479 VDDA.t130 GNDA 0.050121f
C3480 VDDA.n381 GNDA 0.067544f
C3481 VDDA.n382 GNDA 0.144756f
C3482 VDDA.t129 GNDA 0.151746f
C3483 VDDA.t275 GNDA 0.105912f
C3484 VDDA.t22 GNDA 0.105912f
C3485 VDDA.t126 GNDA 0.151746f
C3486 VDDA.n383 GNDA 0.144756f
C3487 VDDA.n384 GNDA 0.067544f
C3488 VDDA.t125 GNDA 0.029712f
C3489 VDDA.n385 GNDA 0.08592f
C3490 VDDA.n386 GNDA 0.097507f
C3491 VDDA.n387 GNDA 0.064392f
C3492 VDDA.n388 GNDA 0.268732f
C3493 VDDA.n389 GNDA 0.3818f
C3494 VDDA.n390 GNDA 0.043503f
C3495 VDDA.t441 GNDA 0.013755f
C3496 VDDA.t259 GNDA 0.013755f
C3497 VDDA.n391 GNDA 0.028091f
C3498 VDDA.n392 GNDA 0.140876f
C3499 VDDA.n393 GNDA 0.076283f
C3500 VDDA.t136 GNDA 0.050121f
C3501 VDDA.t172 GNDA 0.050121f
C3502 VDDA.n394 GNDA 0.076283f
C3503 VDDA.t170 GNDA 0.028913f
C3504 VDDA.n395 GNDA 0.043463f
C3505 VDDA.t458 GNDA 0.013755f
C3506 VDDA.t320 GNDA 0.013755f
C3507 VDDA.n396 GNDA 0.028091f
C3508 VDDA.n397 GNDA 0.140868f
C3509 VDDA.n398 GNDA 0.076377f
C3510 VDDA.t103 GNDA 0.050121f
C3511 VDDA.t148 GNDA 0.050121f
C3512 VDDA.n399 GNDA 0.076377f
C3513 VDDA.t146 GNDA 0.027992f
C3514 VDDA.n400 GNDA 0.043503f
C3515 VDDA.t211 GNDA 0.013755f
C3516 VDDA.t443 GNDA 0.013755f
C3517 VDDA.n401 GNDA 0.028091f
C3518 VDDA.n402 GNDA 0.140876f
C3519 VDDA.n403 GNDA 0.076283f
C3520 VDDA.t157 GNDA 0.050121f
C3521 VDDA.t115 GNDA 0.050121f
C3522 VDDA.n404 GNDA 0.076283f
C3523 VDDA.t113 GNDA 0.027992f
C3524 VDDA.t338 GNDA 0.013755f
C3525 VDDA.t261 GNDA 0.013755f
C3526 VDDA.n405 GNDA 0.028091f
C3527 VDDA.n406 GNDA 0.140876f
C3528 VDDA.n407 GNDA 0.071624f
C3529 VDDA.n408 GNDA 0.07535f
C3530 VDDA.n409 GNDA 0.078054f
C3531 VDDA.n410 GNDA 0.144756f
C3532 VDDA.t114 GNDA 0.151746f
C3533 VDDA.t337 GNDA 0.105912f
C3534 VDDA.t260 GNDA 0.105912f
C3535 VDDA.t210 GNDA 0.105912f
C3536 VDDA.t442 GNDA 0.105912f
C3537 VDDA.t156 GNDA 0.151746f
C3538 VDDA.n411 GNDA 0.144756f
C3539 VDDA.n412 GNDA 0.078054f
C3540 VDDA.t155 GNDA 0.028913f
C3541 VDDA.n413 GNDA 0.072633f
C3542 VDDA.n414 GNDA 0.068774f
C3543 VDDA.n415 GNDA 0.043463f
C3544 VDDA.n416 GNDA 0.043463f
C3545 VDDA.t218 GNDA 0.013755f
C3546 VDDA.t263 GNDA 0.013755f
C3547 VDDA.n417 GNDA 0.028091f
C3548 VDDA.n418 GNDA 0.140868f
C3549 VDDA.n419 GNDA 0.044794f
C3550 VDDA.t220 GNDA 0.013755f
C3551 VDDA.t439 GNDA 0.013755f
C3552 VDDA.n420 GNDA 0.028091f
C3553 VDDA.n421 GNDA 0.140868f
C3554 VDDA.n422 GNDA 0.044794f
C3555 VDDA.n423 GNDA 0.044794f
C3556 VDDA.t300 GNDA 0.013755f
C3557 VDDA.t21 GNDA 0.013755f
C3558 VDDA.n424 GNDA 0.028091f
C3559 VDDA.n425 GNDA 0.140868f
C3560 VDDA.n426 GNDA 0.043463f
C3561 VDDA.t437 GNDA 0.013755f
C3562 VDDA.t213 GNDA 0.013755f
C3563 VDDA.n427 GNDA 0.028091f
C3564 VDDA.n428 GNDA 0.140868f
C3565 VDDA.n429 GNDA 0.043463f
C3566 VDDA.n430 GNDA 0.068774f
C3567 VDDA.n431 GNDA 0.071623f
C3568 VDDA.n432 GNDA 0.078219f
C3569 VDDA.n433 GNDA 0.144756f
C3570 VDDA.t147 GNDA 0.151746f
C3571 VDDA.t436 GNDA 0.105912f
C3572 VDDA.t212 GNDA 0.105912f
C3573 VDDA.t299 GNDA 0.105912f
C3574 VDDA.t20 GNDA 0.105912f
C3575 VDDA.t219 GNDA 0.105912f
C3576 VDDA.t438 GNDA 0.105912f
C3577 VDDA.t217 GNDA 0.105912f
C3578 VDDA.t262 GNDA 0.105912f
C3579 VDDA.t457 GNDA 0.105912f
C3580 VDDA.t319 GNDA 0.105912f
C3581 VDDA.t102 GNDA 0.151746f
C3582 VDDA.n434 GNDA 0.144756f
C3583 VDDA.n435 GNDA 0.078219f
C3584 VDDA.t101 GNDA 0.027992f
C3585 VDDA.n436 GNDA 0.071623f
C3586 VDDA.n437 GNDA 0.068774f
C3587 VDDA.t456 GNDA 0.013755f
C3588 VDDA.t257 GNDA 0.013755f
C3589 VDDA.n438 GNDA 0.028091f
C3590 VDDA.n439 GNDA 0.140876f
C3591 VDDA.n440 GNDA 0.043503f
C3592 VDDA.n441 GNDA 0.068774f
C3593 VDDA.n442 GNDA 0.072633f
C3594 VDDA.n443 GNDA 0.078054f
C3595 VDDA.n444 GNDA 0.144756f
C3596 VDDA.t171 GNDA 0.151746f
C3597 VDDA.t455 GNDA 0.105912f
C3598 VDDA.t256 GNDA 0.105912f
C3599 VDDA.t440 GNDA 0.105912f
C3600 VDDA.t258 GNDA 0.105912f
C3601 VDDA.t135 GNDA 0.151746f
C3602 VDDA.n445 GNDA 0.144756f
C3603 VDDA.n446 GNDA 0.078054f
C3604 VDDA.t134 GNDA 0.027992f
C3605 VDDA.n447 GNDA 0.071835f
C3606 VDDA.n448 GNDA 0.26332f
C3607 VDDA.n449 GNDA 0.28932f
C3608 VDDA.n450 GNDA 1.54497f
C3609 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 GNDA 0.021174f
C3610 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 GNDA 0.021174f
C3611 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 GNDA 0.043243f
C3612 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 GNDA 0.16469f
C3613 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 GNDA 0.021174f
C3614 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 GNDA 0.021174f
C3615 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 GNDA 0.043243f
C3616 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 GNDA 0.227515f
C3617 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 GNDA 0.157479f
C3618 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 GNDA 0.021174f
C3619 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 GNDA 0.021174f
C3620 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 GNDA 0.043243f
C3621 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 GNDA 0.216541f
C3622 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 GNDA 0.163297f
C3623 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 GNDA 0.108203f
C3624 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 GNDA 0.273637f
C3625 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 GNDA 0.06689f
C3626 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 GNDA 0.118314f
C3627 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 GNDA 0.042349f
C3628 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 GNDA 0.042349f
C3629 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 GNDA 0.086586f
C3630 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 GNDA 0.290839f
C3631 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 GNDA 0.042349f
C3632 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 GNDA 0.042349f
C3633 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 GNDA 0.086586f
C3634 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 GNDA 0.28008f
C3635 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 GNDA 0.113731f
C3636 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n16 GNDA 0.06689f
C3637 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 GNDA 0.042349f
C3638 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 GNDA 0.042349f
C3639 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n17 GNDA 0.086586f
C3640 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n18 GNDA 0.28008f
C3641 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n19 GNDA 0.069335f
C3642 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 GNDA 0.042349f
C3643 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 GNDA 0.042349f
C3644 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n20 GNDA 0.086586f
C3645 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n21 GNDA 0.28008f
C3646 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n22 GNDA 0.118314f
C3647 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 GNDA 0.042349f
C3648 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 GNDA 0.042349f
C3649 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n23 GNDA 0.086586f
C3650 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n24 GNDA 0.285613f
C3651 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n25 GNDA 0.171152f
C3652 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n26 GNDA 1.94694f
C3653 bgr_0.V_CMFB_S3 GNDA 1.08719f
C3654 two_stage_opamp_dummy_magic_0.Y.t0 GNDA 0.037869f
C3655 two_stage_opamp_dummy_magic_0.Y.t24 GNDA 0.037869f
C3656 two_stage_opamp_dummy_magic_0.Y.n0 GNDA 0.082398f
C3657 two_stage_opamp_dummy_magic_0.Y.n1 GNDA 0.256617f
C3658 two_stage_opamp_dummy_magic_0.Y.n2 GNDA 0.080536f
C3659 two_stage_opamp_dummy_magic_0.Y.t12 GNDA 0.037869f
C3660 two_stage_opamp_dummy_magic_0.Y.t21 GNDA 0.037869f
C3661 two_stage_opamp_dummy_magic_0.Y.n3 GNDA 0.082398f
C3662 two_stage_opamp_dummy_magic_0.Y.n4 GNDA 0.327392f
C3663 two_stage_opamp_dummy_magic_0.Y.t20 GNDA 0.037869f
C3664 two_stage_opamp_dummy_magic_0.Y.t9 GNDA 0.037869f
C3665 two_stage_opamp_dummy_magic_0.Y.n5 GNDA 0.082398f
C3666 two_stage_opamp_dummy_magic_0.Y.n6 GNDA 0.327392f
C3667 two_stage_opamp_dummy_magic_0.Y.n7 GNDA 0.136897f
C3668 two_stage_opamp_dummy_magic_0.Y.t4 GNDA 0.037869f
C3669 two_stage_opamp_dummy_magic_0.Y.t15 GNDA 0.037869f
C3670 two_stage_opamp_dummy_magic_0.Y.n8 GNDA 0.082398f
C3671 two_stage_opamp_dummy_magic_0.Y.n9 GNDA 0.314197f
C3672 two_stage_opamp_dummy_magic_0.Y.n10 GNDA 0.144815f
C3673 two_stage_opamp_dummy_magic_0.Y.t17 GNDA 0.037869f
C3674 two_stage_opamp_dummy_magic_0.Y.t1 GNDA 0.037869f
C3675 two_stage_opamp_dummy_magic_0.Y.n11 GNDA 0.082398f
C3676 two_stage_opamp_dummy_magic_0.Y.n12 GNDA 0.314197f
C3677 two_stage_opamp_dummy_magic_0.Y.n13 GNDA 0.084589f
C3678 two_stage_opamp_dummy_magic_0.Y.n14 GNDA 0.084589f
C3679 two_stage_opamp_dummy_magic_0.Y.n15 GNDA 0.144815f
C3680 two_stage_opamp_dummy_magic_0.Y.t11 GNDA 0.037869f
C3681 two_stage_opamp_dummy_magic_0.Y.t10 GNDA 0.037869f
C3682 two_stage_opamp_dummy_magic_0.Y.n16 GNDA 0.082398f
C3683 two_stage_opamp_dummy_magic_0.Y.n17 GNDA 0.314197f
C3684 two_stage_opamp_dummy_magic_0.Y.n18 GNDA 0.136897f
C3685 two_stage_opamp_dummy_magic_0.Y.n19 GNDA 0.075738f
C3686 two_stage_opamp_dummy_magic_0.Y.n20 GNDA 0.32544f
C3687 two_stage_opamp_dummy_magic_0.Y.n21 GNDA 0.101828f
C3688 two_stage_opamp_dummy_magic_0.Y.n22 GNDA 0.095842f
C3689 two_stage_opamp_dummy_magic_0.Y.t18 GNDA 0.08836f
C3690 two_stage_opamp_dummy_magic_0.Y.t7 GNDA 0.08836f
C3691 two_stage_opamp_dummy_magic_0.Y.n23 GNDA 0.180751f
C3692 two_stage_opamp_dummy_magic_0.Y.n24 GNDA 0.61368f
C3693 two_stage_opamp_dummy_magic_0.Y.n25 GNDA 0.163497f
C3694 two_stage_opamp_dummy_magic_0.Y.t8 GNDA 0.08836f
C3695 two_stage_opamp_dummy_magic_0.Y.t16 GNDA 0.08836f
C3696 two_stage_opamp_dummy_magic_0.Y.n26 GNDA 0.180751f
C3697 two_stage_opamp_dummy_magic_0.Y.n27 GNDA 0.597331f
C3698 two_stage_opamp_dummy_magic_0.Y.n28 GNDA 0.175101f
C3699 two_stage_opamp_dummy_magic_0.Y.t13 GNDA 0.08836f
C3700 two_stage_opamp_dummy_magic_0.Y.t19 GNDA 0.08836f
C3701 two_stage_opamp_dummy_magic_0.Y.n29 GNDA 0.180751f
C3702 two_stage_opamp_dummy_magic_0.Y.n30 GNDA 0.597331f
C3703 two_stage_opamp_dummy_magic_0.Y.n31 GNDA 0.101828f
C3704 two_stage_opamp_dummy_magic_0.Y.n32 GNDA 0.101828f
C3705 two_stage_opamp_dummy_magic_0.Y.t5 GNDA 0.08836f
C3706 two_stage_opamp_dummy_magic_0.Y.t2 GNDA 0.08836f
C3707 two_stage_opamp_dummy_magic_0.Y.n33 GNDA 0.180751f
C3708 two_stage_opamp_dummy_magic_0.Y.n34 GNDA 0.597331f
C3709 two_stage_opamp_dummy_magic_0.Y.n35 GNDA 0.095842f
C3710 two_stage_opamp_dummy_magic_0.Y.t6 GNDA 0.08836f
C3711 two_stage_opamp_dummy_magic_0.Y.t22 GNDA 0.08836f
C3712 two_stage_opamp_dummy_magic_0.Y.n36 GNDA 0.180751f
C3713 two_stage_opamp_dummy_magic_0.Y.n37 GNDA 0.597331f
C3714 two_stage_opamp_dummy_magic_0.Y.n38 GNDA 0.163497f
C3715 two_stage_opamp_dummy_magic_0.Y.t3 GNDA 0.08836f
C3716 two_stage_opamp_dummy_magic_0.Y.t14 GNDA 0.08836f
C3717 two_stage_opamp_dummy_magic_0.Y.n39 GNDA 0.180751f
C3718 two_stage_opamp_dummy_magic_0.Y.n40 GNDA 0.605322f
C3719 two_stage_opamp_dummy_magic_0.Y.n41 GNDA 0.397499f
C3720 two_stage_opamp_dummy_magic_0.Y.t32 GNDA 0.053016f
C3721 two_stage_opamp_dummy_magic_0.Y.t25 GNDA 0.053016f
C3722 two_stage_opamp_dummy_magic_0.Y.t39 GNDA 0.053016f
C3723 two_stage_opamp_dummy_magic_0.Y.t52 GNDA 0.053016f
C3724 two_stage_opamp_dummy_magic_0.Y.t37 GNDA 0.064377f
C3725 two_stage_opamp_dummy_magic_0.Y.n42 GNDA 0.064377f
C3726 two_stage_opamp_dummy_magic_0.Y.n43 GNDA 0.041656f
C3727 two_stage_opamp_dummy_magic_0.Y.n44 GNDA 0.041656f
C3728 two_stage_opamp_dummy_magic_0.Y.t47 GNDA 0.053016f
C3729 two_stage_opamp_dummy_magic_0.Y.t35 GNDA 0.053016f
C3730 two_stage_opamp_dummy_magic_0.Y.t50 GNDA 0.053016f
C3731 two_stage_opamp_dummy_magic_0.Y.t43 GNDA 0.053016f
C3732 two_stage_opamp_dummy_magic_0.Y.t30 GNDA 0.064377f
C3733 two_stage_opamp_dummy_magic_0.Y.n45 GNDA 0.064377f
C3734 two_stage_opamp_dummy_magic_0.Y.n46 GNDA 0.041656f
C3735 two_stage_opamp_dummy_magic_0.Y.n47 GNDA 0.041656f
C3736 two_stage_opamp_dummy_magic_0.Y.n48 GNDA 0.041656f
C3737 two_stage_opamp_dummy_magic_0.Y.n49 GNDA 0.070025f
C3738 two_stage_opamp_dummy_magic_0.Y.t54 GNDA 0.081418f
C3739 two_stage_opamp_dummy_magic_0.Y.t48 GNDA 0.081418f
C3740 two_stage_opamp_dummy_magic_0.Y.t33 GNDA 0.081418f
C3741 two_stage_opamp_dummy_magic_0.Y.t45 GNDA 0.081418f
C3742 two_stage_opamp_dummy_magic_0.Y.t29 GNDA 0.092558f
C3743 two_stage_opamp_dummy_magic_0.Y.n50 GNDA 0.083532f
C3744 two_stage_opamp_dummy_magic_0.Y.n51 GNDA 0.051123f
C3745 two_stage_opamp_dummy_magic_0.Y.n52 GNDA 0.051123f
C3746 two_stage_opamp_dummy_magic_0.Y.t41 GNDA 0.081418f
C3747 two_stage_opamp_dummy_magic_0.Y.t27 GNDA 0.081418f
C3748 two_stage_opamp_dummy_magic_0.Y.t42 GNDA 0.081418f
C3749 two_stage_opamp_dummy_magic_0.Y.t38 GNDA 0.081418f
C3750 two_stage_opamp_dummy_magic_0.Y.t53 GNDA 0.092558f
C3751 two_stage_opamp_dummy_magic_0.Y.n53 GNDA 0.083532f
C3752 two_stage_opamp_dummy_magic_0.Y.n54 GNDA 0.051123f
C3753 two_stage_opamp_dummy_magic_0.Y.n55 GNDA 0.051123f
C3754 two_stage_opamp_dummy_magic_0.Y.n56 GNDA 0.051123f
C3755 two_stage_opamp_dummy_magic_0.Y.n57 GNDA 0.077631f
C3756 two_stage_opamp_dummy_magic_0.Y.n58 GNDA 0.114144f
C3757 two_stage_opamp_dummy_magic_0.Y.n59 GNDA 1.08414f
C3758 two_stage_opamp_dummy_magic_0.Y.n60 GNDA 0.423626f
C3759 two_stage_opamp_dummy_magic_0.Y.t28 GNDA 0.166623f
C3760 two_stage_opamp_dummy_magic_0.Y.t51 GNDA 0.166623f
C3761 two_stage_opamp_dummy_magic_0.Y.t36 GNDA 0.166623f
C3762 two_stage_opamp_dummy_magic_0.Y.t49 GNDA 0.166623f
C3763 two_stage_opamp_dummy_magic_0.Y.t34 GNDA 0.177465f
C3764 two_stage_opamp_dummy_magic_0.Y.n61 GNDA 0.140633f
C3765 two_stage_opamp_dummy_magic_0.Y.n62 GNDA 0.079524f
C3766 two_stage_opamp_dummy_magic_0.Y.n63 GNDA 0.079524f
C3767 two_stage_opamp_dummy_magic_0.Y.t44 GNDA 0.166623f
C3768 two_stage_opamp_dummy_magic_0.Y.t31 GNDA 0.166623f
C3769 two_stage_opamp_dummy_magic_0.Y.t46 GNDA 0.166623f
C3770 two_stage_opamp_dummy_magic_0.Y.t40 GNDA 0.166623f
C3771 two_stage_opamp_dummy_magic_0.Y.t26 GNDA 0.177465f
C3772 two_stage_opamp_dummy_magic_0.Y.n64 GNDA 0.140633f
C3773 two_stage_opamp_dummy_magic_0.Y.n65 GNDA 0.079524f
C3774 two_stage_opamp_dummy_magic_0.Y.n66 GNDA 0.079524f
C3775 two_stage_opamp_dummy_magic_0.Y.n67 GNDA 0.079524f
C3776 two_stage_opamp_dummy_magic_0.Y.n68 GNDA 0.11829f
C3777 two_stage_opamp_dummy_magic_0.Y.n69 GNDA 1.30961f
C3778 two_stage_opamp_dummy_magic_0.Y.t23 GNDA 1.21964f
C3779 bgr_0.Vin+.t5 GNDA 0.249247f
C3780 bgr_0.Vin+.t8 GNDA 0.036348f
C3781 bgr_0.Vin+.t9 GNDA 0.023627f
C3782 bgr_0.Vin+.n0 GNDA 0.077956f
C3783 bgr_0.Vin+.t6 GNDA 0.023627f
C3784 bgr_0.Vin+.n1 GNDA 0.060664f
C3785 bgr_0.Vin+.t10 GNDA 0.023627f
C3786 bgr_0.Vin+.n2 GNDA 0.060664f
C3787 bgr_0.Vin+.t7 GNDA 0.023627f
C3788 bgr_0.Vin+.n3 GNDA 0.138961f
C3789 bgr_0.Vin+.n4 GNDA 1.72958f
C3790 bgr_0.Vin+.t2 GNDA 0.076628f
C3791 bgr_0.Vin+.t0 GNDA 0.076628f
C3792 bgr_0.Vin+.n5 GNDA 0.156734f
C3793 bgr_0.Vin+.n6 GNDA 0.79018f
C3794 bgr_0.Vin+.t1 GNDA 0.076628f
C3795 bgr_0.Vin+.t3 GNDA 0.076628f
C3796 bgr_0.Vin+.n7 GNDA 0.156734f
C3797 bgr_0.Vin+.n8 GNDA 0.79018f
C3798 bgr_0.Vin+.n9 GNDA 1.34635f
C3799 bgr_0.Vin+.n10 GNDA 2.47471f
C3800 bgr_0.Vin+.t4 GNDA 0.330676f
.ends

