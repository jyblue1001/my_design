magic
tech sky130A
timestamp 1754396681
<< nwell >>
rect 16315 1310 16695 1450
rect 16825 1310 17315 1450
rect 17445 1310 18155 1450
rect 18285 1310 18775 1450
rect 16375 745 16760 885
rect 16910 645 18690 985
rect 18845 745 19170 985
rect 16360 5 17725 145
rect 17880 5 19240 145
<< pwell >>
rect 17780 -4300 17820 -4120
<< nmos >>
rect 17000 -410 17020 -160
rect 17060 -410 17080 -160
rect 18520 -410 18540 -160
rect 18580 -410 18600 -160
rect 16570 -945 17070 -695
rect 17190 -945 17690 -695
rect 17910 -945 18410 -695
rect 18530 -945 19030 -695
rect 16780 -1250 17780 -1150
rect 17820 -1250 18820 -1150
rect 16640 -1640 16655 -1540
rect 16695 -1640 16710 -1540
rect 16750 -1640 16765 -1540
rect 16805 -1640 16820 -1540
rect 16860 -1640 16875 -1540
rect 17065 -1640 17080 -1540
rect 17120 -1640 17135 -1540
rect 17175 -1640 17190 -1540
rect 17230 -1640 17245 -1540
rect 17285 -1640 17300 -1540
rect 17340 -1640 17355 -1540
rect 17395 -1640 17410 -1540
rect 17450 -1640 17465 -1540
rect 17655 -1640 17670 -1540
rect 17710 -1640 17725 -1540
rect 17765 -1640 17780 -1540
rect 17820 -1640 17835 -1540
rect 17875 -1640 17890 -1540
rect 17930 -1640 17945 -1540
rect 18135 -1640 18150 -1540
rect 18190 -1640 18205 -1540
rect 18245 -1640 18260 -1540
rect 18300 -1640 18315 -1540
rect 18355 -1640 18370 -1540
rect 18410 -1640 18425 -1540
rect 18465 -1640 18480 -1540
rect 18520 -1640 18535 -1540
<< pmos >>
rect 16415 1330 16430 1430
rect 16470 1330 16485 1430
rect 16525 1330 16540 1430
rect 16580 1330 16595 1430
rect 16925 1330 16940 1430
rect 16980 1330 16995 1430
rect 17035 1330 17050 1430
rect 17090 1330 17105 1430
rect 17145 1330 17160 1430
rect 17200 1330 17215 1430
rect 17545 1330 17560 1430
rect 17600 1330 17615 1430
rect 17655 1330 17670 1430
rect 17710 1330 17725 1430
rect 17765 1330 17780 1430
rect 17820 1330 17835 1430
rect 17875 1330 17890 1430
rect 17930 1330 17945 1430
rect 17985 1330 18000 1430
rect 18040 1330 18055 1430
rect 18385 1330 18400 1430
rect 18440 1330 18455 1430
rect 18495 1330 18510 1430
rect 18550 1330 18565 1430
rect 18605 1330 18620 1430
rect 18660 1330 18675 1430
rect 16475 765 16490 865
rect 16530 765 16545 865
rect 16585 765 16600 865
rect 16640 765 16655 865
rect 17010 665 17060 965
rect 17100 665 17150 965
rect 17190 665 17240 965
rect 17280 665 17330 965
rect 17370 665 17420 965
rect 17460 665 17510 965
rect 17550 665 17600 965
rect 17640 665 17690 965
rect 17730 665 17780 965
rect 17820 665 17870 965
rect 17910 665 17960 965
rect 18000 665 18050 965
rect 18090 665 18140 965
rect 18180 665 18230 965
rect 18270 665 18320 965
rect 18360 665 18410 965
rect 18450 665 18500 965
rect 18540 665 18590 965
rect 18945 765 18960 965
rect 19000 765 19015 965
rect 19055 765 19070 965
rect 16460 25 16480 125
rect 16520 25 16540 125
rect 16580 25 16600 125
rect 16640 25 16660 125
rect 16700 25 16720 125
rect 16760 25 16780 125
rect 16820 25 16840 125
rect 16880 25 16900 125
rect 16940 25 16960 125
rect 17000 25 17020 125
rect 17060 25 17080 125
rect 17120 25 17140 125
rect 17180 25 17200 125
rect 17240 25 17260 125
rect 17300 25 17320 125
rect 17360 25 17380 125
rect 17420 25 17440 125
rect 17480 25 17500 125
rect 17540 25 17560 125
rect 17600 25 17620 125
rect 17980 25 18000 125
rect 18040 25 18060 125
rect 18100 25 18120 125
rect 18160 25 18180 125
rect 18220 25 18240 125
rect 18280 25 18300 125
rect 18340 25 18360 125
rect 18400 25 18420 125
rect 18460 25 18480 125
rect 18520 25 18540 125
rect 18580 25 18600 125
rect 18640 25 18660 125
rect 18700 25 18720 125
rect 18760 25 18780 125
rect 18820 25 18840 125
rect 18880 25 18900 125
rect 18940 25 18960 125
rect 19000 25 19020 125
rect 19060 25 19080 125
rect 19120 25 19140 125
<< ndiff >>
rect 16960 -175 17000 -160
rect 16960 -195 16970 -175
rect 16990 -195 17000 -175
rect 16960 -225 17000 -195
rect 16960 -245 16970 -225
rect 16990 -245 17000 -225
rect 16960 -275 17000 -245
rect 16960 -295 16970 -275
rect 16990 -295 17000 -275
rect 16960 -325 17000 -295
rect 16960 -345 16970 -325
rect 16990 -345 17000 -325
rect 16960 -375 17000 -345
rect 16960 -395 16970 -375
rect 16990 -395 17000 -375
rect 16960 -410 17000 -395
rect 17020 -175 17060 -160
rect 17020 -195 17030 -175
rect 17050 -195 17060 -175
rect 17020 -225 17060 -195
rect 17020 -245 17030 -225
rect 17050 -245 17060 -225
rect 17020 -275 17060 -245
rect 17020 -295 17030 -275
rect 17050 -295 17060 -275
rect 17020 -325 17060 -295
rect 17020 -345 17030 -325
rect 17050 -345 17060 -325
rect 17020 -375 17060 -345
rect 17020 -395 17030 -375
rect 17050 -395 17060 -375
rect 17020 -410 17060 -395
rect 17080 -175 17120 -160
rect 17080 -195 17090 -175
rect 17110 -195 17120 -175
rect 17080 -225 17120 -195
rect 17080 -245 17090 -225
rect 17110 -245 17120 -225
rect 17080 -275 17120 -245
rect 17080 -295 17090 -275
rect 17110 -295 17120 -275
rect 18480 -175 18520 -160
rect 18480 -195 18490 -175
rect 18510 -195 18520 -175
rect 18480 -225 18520 -195
rect 18480 -245 18490 -225
rect 18510 -245 18520 -225
rect 18480 -275 18520 -245
rect 17080 -325 17120 -295
rect 17080 -345 17090 -325
rect 17110 -345 17120 -325
rect 17080 -375 17120 -345
rect 17080 -395 17090 -375
rect 17110 -395 17120 -375
rect 17080 -410 17120 -395
rect 18480 -295 18490 -275
rect 18510 -295 18520 -275
rect 18480 -325 18520 -295
rect 18480 -345 18490 -325
rect 18510 -345 18520 -325
rect 18480 -375 18520 -345
rect 18480 -395 18490 -375
rect 18510 -395 18520 -375
rect 18480 -410 18520 -395
rect 18540 -175 18580 -160
rect 18540 -195 18550 -175
rect 18570 -195 18580 -175
rect 18540 -225 18580 -195
rect 18540 -245 18550 -225
rect 18570 -245 18580 -225
rect 18540 -275 18580 -245
rect 18540 -295 18550 -275
rect 18570 -295 18580 -275
rect 18540 -325 18580 -295
rect 18540 -345 18550 -325
rect 18570 -345 18580 -325
rect 18540 -375 18580 -345
rect 18540 -395 18550 -375
rect 18570 -395 18580 -375
rect 18540 -410 18580 -395
rect 18600 -175 18640 -160
rect 18600 -195 18610 -175
rect 18630 -195 18640 -175
rect 18600 -225 18640 -195
rect 18600 -245 18610 -225
rect 18630 -245 18640 -225
rect 18600 -275 18640 -245
rect 18600 -295 18610 -275
rect 18630 -295 18640 -275
rect 18600 -325 18640 -295
rect 18600 -345 18610 -325
rect 18630 -345 18640 -325
rect 18600 -375 18640 -345
rect 18600 -395 18610 -375
rect 18630 -395 18640 -375
rect 18600 -410 18640 -395
rect 16530 -710 16570 -695
rect 16530 -730 16540 -710
rect 16560 -730 16570 -710
rect 16530 -760 16570 -730
rect 16530 -780 16540 -760
rect 16560 -780 16570 -760
rect 16530 -810 16570 -780
rect 16530 -830 16540 -810
rect 16560 -830 16570 -810
rect 16530 -860 16570 -830
rect 16530 -880 16540 -860
rect 16560 -880 16570 -860
rect 16530 -910 16570 -880
rect 16530 -930 16540 -910
rect 16560 -930 16570 -910
rect 16530 -945 16570 -930
rect 17070 -710 17110 -695
rect 17150 -710 17190 -695
rect 17070 -730 17080 -710
rect 17100 -730 17110 -710
rect 17150 -730 17160 -710
rect 17180 -730 17190 -710
rect 17070 -760 17110 -730
rect 17150 -760 17190 -730
rect 17070 -780 17080 -760
rect 17100 -780 17110 -760
rect 17150 -780 17160 -760
rect 17180 -780 17190 -760
rect 17070 -810 17110 -780
rect 17150 -810 17190 -780
rect 17070 -830 17080 -810
rect 17100 -830 17110 -810
rect 17150 -830 17160 -810
rect 17180 -830 17190 -810
rect 17070 -860 17110 -830
rect 17150 -860 17190 -830
rect 17070 -880 17080 -860
rect 17100 -880 17110 -860
rect 17150 -880 17160 -860
rect 17180 -880 17190 -860
rect 17070 -910 17110 -880
rect 17150 -910 17190 -880
rect 17070 -930 17080 -910
rect 17100 -930 17110 -910
rect 17150 -930 17160 -910
rect 17180 -930 17190 -910
rect 17070 -940 17110 -930
rect 17150 -940 17190 -930
rect 17070 -945 17190 -940
rect 17690 -710 17730 -695
rect 17690 -730 17700 -710
rect 17720 -730 17730 -710
rect 17690 -760 17730 -730
rect 17690 -780 17700 -760
rect 17720 -780 17730 -760
rect 17690 -810 17730 -780
rect 17690 -830 17700 -810
rect 17720 -830 17730 -810
rect 17690 -860 17730 -830
rect 17690 -880 17700 -860
rect 17720 -880 17730 -860
rect 17690 -910 17730 -880
rect 17690 -930 17700 -910
rect 17720 -930 17730 -910
rect 17690 -945 17730 -930
rect 17870 -710 17910 -695
rect 17870 -730 17880 -710
rect 17900 -730 17910 -710
rect 17870 -760 17910 -730
rect 17870 -780 17880 -760
rect 17900 -780 17910 -760
rect 17870 -810 17910 -780
rect 17870 -830 17880 -810
rect 17900 -830 17910 -810
rect 17870 -860 17910 -830
rect 17870 -880 17880 -860
rect 17900 -880 17910 -860
rect 17870 -910 17910 -880
rect 17870 -930 17880 -910
rect 17900 -930 17910 -910
rect 17870 -945 17910 -930
rect 18410 -710 18450 -695
rect 18490 -710 18530 -695
rect 18410 -730 18420 -710
rect 18440 -730 18450 -710
rect 18490 -730 18500 -710
rect 18520 -730 18530 -710
rect 18410 -760 18450 -730
rect 18490 -760 18530 -730
rect 18410 -780 18420 -760
rect 18440 -780 18450 -760
rect 18490 -780 18500 -760
rect 18520 -780 18530 -760
rect 18410 -810 18450 -780
rect 18490 -810 18530 -780
rect 18410 -830 18420 -810
rect 18440 -830 18450 -810
rect 18490 -830 18500 -810
rect 18520 -830 18530 -810
rect 18410 -860 18450 -830
rect 18490 -860 18530 -830
rect 18410 -880 18420 -860
rect 18440 -880 18450 -860
rect 18490 -880 18500 -860
rect 18520 -880 18530 -860
rect 18410 -910 18450 -880
rect 18490 -910 18530 -880
rect 18410 -930 18420 -910
rect 18440 -930 18450 -910
rect 18490 -930 18500 -910
rect 18520 -930 18530 -910
rect 18410 -945 18450 -930
rect 18490 -945 18530 -930
rect 19030 -710 19070 -695
rect 19030 -730 19040 -710
rect 19060 -730 19070 -710
rect 19030 -760 19070 -730
rect 19030 -780 19040 -760
rect 19060 -780 19070 -760
rect 19030 -810 19070 -780
rect 19030 -830 19040 -810
rect 19060 -830 19070 -810
rect 19030 -860 19070 -830
rect 19030 -880 19040 -860
rect 19060 -880 19070 -860
rect 19030 -910 19070 -880
rect 19030 -930 19040 -910
rect 19060 -930 19070 -910
rect 19030 -945 19070 -930
rect 16740 -1165 16780 -1150
rect 16740 -1185 16750 -1165
rect 16770 -1185 16780 -1165
rect 16740 -1215 16780 -1185
rect 16740 -1235 16750 -1215
rect 16770 -1235 16780 -1215
rect 16740 -1250 16780 -1235
rect 17780 -1165 17820 -1150
rect 17780 -1185 17790 -1165
rect 17810 -1185 17820 -1165
rect 17780 -1215 17820 -1185
rect 17780 -1235 17790 -1215
rect 17810 -1235 17820 -1215
rect 17780 -1250 17820 -1235
rect 18820 -1165 18860 -1150
rect 18820 -1185 18830 -1165
rect 18850 -1185 18860 -1165
rect 18820 -1215 18860 -1185
rect 18820 -1235 18830 -1215
rect 18850 -1235 18860 -1215
rect 18820 -1250 18860 -1235
rect 16600 -1555 16640 -1540
rect 16600 -1575 16610 -1555
rect 16630 -1575 16640 -1555
rect 16600 -1605 16640 -1575
rect 16600 -1625 16610 -1605
rect 16630 -1625 16640 -1605
rect 16600 -1640 16640 -1625
rect 16655 -1555 16695 -1540
rect 16655 -1575 16665 -1555
rect 16685 -1575 16695 -1555
rect 16655 -1605 16695 -1575
rect 16655 -1625 16665 -1605
rect 16685 -1625 16695 -1605
rect 16655 -1640 16695 -1625
rect 16710 -1555 16750 -1540
rect 16710 -1575 16720 -1555
rect 16740 -1575 16750 -1555
rect 16710 -1605 16750 -1575
rect 16710 -1625 16720 -1605
rect 16740 -1625 16750 -1605
rect 16710 -1640 16750 -1625
rect 16765 -1555 16805 -1540
rect 16765 -1575 16775 -1555
rect 16795 -1575 16805 -1555
rect 16765 -1605 16805 -1575
rect 16765 -1625 16775 -1605
rect 16795 -1625 16805 -1605
rect 16765 -1640 16805 -1625
rect 16820 -1555 16860 -1540
rect 16820 -1575 16830 -1555
rect 16850 -1575 16860 -1555
rect 16820 -1605 16860 -1575
rect 16820 -1625 16830 -1605
rect 16850 -1625 16860 -1605
rect 16820 -1640 16860 -1625
rect 16875 -1555 16915 -1540
rect 16875 -1575 16885 -1555
rect 16905 -1575 16915 -1555
rect 16875 -1605 16915 -1575
rect 16875 -1625 16885 -1605
rect 16905 -1625 16915 -1605
rect 16875 -1640 16915 -1625
rect 17025 -1555 17065 -1540
rect 17025 -1575 17035 -1555
rect 17055 -1575 17065 -1555
rect 17025 -1605 17065 -1575
rect 17025 -1625 17035 -1605
rect 17055 -1625 17065 -1605
rect 17025 -1640 17065 -1625
rect 17080 -1555 17120 -1540
rect 17080 -1575 17090 -1555
rect 17110 -1575 17120 -1555
rect 17080 -1605 17120 -1575
rect 17080 -1625 17090 -1605
rect 17110 -1625 17120 -1605
rect 17080 -1640 17120 -1625
rect 17135 -1555 17175 -1540
rect 17135 -1575 17145 -1555
rect 17165 -1575 17175 -1555
rect 17135 -1605 17175 -1575
rect 17135 -1625 17145 -1605
rect 17165 -1625 17175 -1605
rect 17135 -1640 17175 -1625
rect 17190 -1555 17230 -1540
rect 17190 -1575 17200 -1555
rect 17220 -1575 17230 -1555
rect 17190 -1605 17230 -1575
rect 17190 -1625 17200 -1605
rect 17220 -1625 17230 -1605
rect 17190 -1640 17230 -1625
rect 17245 -1555 17285 -1540
rect 17245 -1575 17255 -1555
rect 17275 -1575 17285 -1555
rect 17245 -1605 17285 -1575
rect 17245 -1625 17255 -1605
rect 17275 -1625 17285 -1605
rect 17245 -1640 17285 -1625
rect 17300 -1555 17340 -1540
rect 17300 -1575 17310 -1555
rect 17330 -1575 17340 -1555
rect 17300 -1605 17340 -1575
rect 17300 -1625 17310 -1605
rect 17330 -1625 17340 -1605
rect 17300 -1640 17340 -1625
rect 17355 -1555 17395 -1540
rect 17355 -1575 17365 -1555
rect 17385 -1575 17395 -1555
rect 17355 -1605 17395 -1575
rect 17355 -1625 17365 -1605
rect 17385 -1625 17395 -1605
rect 17355 -1640 17395 -1625
rect 17410 -1555 17450 -1540
rect 17410 -1575 17420 -1555
rect 17440 -1575 17450 -1555
rect 17410 -1605 17450 -1575
rect 17410 -1625 17420 -1605
rect 17440 -1625 17450 -1605
rect 17410 -1640 17450 -1625
rect 17465 -1555 17505 -1540
rect 17465 -1575 17475 -1555
rect 17495 -1575 17505 -1555
rect 17465 -1605 17505 -1575
rect 17465 -1625 17475 -1605
rect 17495 -1625 17505 -1605
rect 17465 -1640 17505 -1625
rect 17615 -1555 17655 -1540
rect 17615 -1575 17625 -1555
rect 17645 -1575 17655 -1555
rect 17615 -1605 17655 -1575
rect 17615 -1625 17625 -1605
rect 17645 -1625 17655 -1605
rect 17615 -1640 17655 -1625
rect 17670 -1555 17710 -1540
rect 17670 -1575 17680 -1555
rect 17700 -1575 17710 -1555
rect 17670 -1605 17710 -1575
rect 17670 -1625 17680 -1605
rect 17700 -1625 17710 -1605
rect 17670 -1640 17710 -1625
rect 17725 -1555 17765 -1540
rect 17725 -1575 17735 -1555
rect 17755 -1575 17765 -1555
rect 17725 -1605 17765 -1575
rect 17725 -1625 17735 -1605
rect 17755 -1625 17765 -1605
rect 17725 -1640 17765 -1625
rect 17780 -1555 17820 -1540
rect 17780 -1575 17790 -1555
rect 17810 -1575 17820 -1555
rect 17780 -1605 17820 -1575
rect 17780 -1625 17790 -1605
rect 17810 -1625 17820 -1605
rect 17780 -1640 17820 -1625
rect 17835 -1555 17875 -1540
rect 17835 -1575 17845 -1555
rect 17865 -1575 17875 -1555
rect 17835 -1605 17875 -1575
rect 17835 -1625 17845 -1605
rect 17865 -1625 17875 -1605
rect 17835 -1640 17875 -1625
rect 17890 -1555 17930 -1540
rect 17890 -1575 17900 -1555
rect 17920 -1575 17930 -1555
rect 17890 -1605 17930 -1575
rect 17890 -1625 17900 -1605
rect 17920 -1625 17930 -1605
rect 17890 -1640 17930 -1625
rect 17945 -1555 17985 -1540
rect 17945 -1575 17955 -1555
rect 17975 -1575 17985 -1555
rect 17945 -1605 17985 -1575
rect 17945 -1625 17955 -1605
rect 17975 -1625 17985 -1605
rect 17945 -1640 17985 -1625
rect 18095 -1555 18135 -1540
rect 18095 -1575 18105 -1555
rect 18125 -1575 18135 -1555
rect 18095 -1605 18135 -1575
rect 18095 -1625 18105 -1605
rect 18125 -1625 18135 -1605
rect 18095 -1640 18135 -1625
rect 18150 -1555 18190 -1540
rect 18150 -1575 18160 -1555
rect 18180 -1575 18190 -1555
rect 18150 -1605 18190 -1575
rect 18150 -1625 18160 -1605
rect 18180 -1625 18190 -1605
rect 18150 -1640 18190 -1625
rect 18205 -1555 18245 -1540
rect 18205 -1575 18215 -1555
rect 18235 -1575 18245 -1555
rect 18205 -1605 18245 -1575
rect 18205 -1625 18215 -1605
rect 18235 -1625 18245 -1605
rect 18205 -1640 18245 -1625
rect 18260 -1555 18300 -1540
rect 18260 -1575 18270 -1555
rect 18290 -1575 18300 -1555
rect 18260 -1605 18300 -1575
rect 18260 -1625 18270 -1605
rect 18290 -1625 18300 -1605
rect 18260 -1640 18300 -1625
rect 18315 -1555 18355 -1540
rect 18315 -1575 18325 -1555
rect 18345 -1575 18355 -1555
rect 18315 -1605 18355 -1575
rect 18315 -1625 18325 -1605
rect 18345 -1625 18355 -1605
rect 18315 -1640 18355 -1625
rect 18370 -1555 18410 -1540
rect 18370 -1575 18380 -1555
rect 18400 -1575 18410 -1555
rect 18370 -1605 18410 -1575
rect 18370 -1625 18380 -1605
rect 18400 -1625 18410 -1605
rect 18370 -1640 18410 -1625
rect 18425 -1555 18465 -1540
rect 18425 -1575 18435 -1555
rect 18455 -1575 18465 -1555
rect 18425 -1605 18465 -1575
rect 18425 -1625 18435 -1605
rect 18455 -1625 18465 -1605
rect 18425 -1640 18465 -1625
rect 18480 -1555 18520 -1540
rect 18480 -1575 18490 -1555
rect 18510 -1575 18520 -1555
rect 18480 -1605 18520 -1575
rect 18480 -1625 18490 -1605
rect 18510 -1625 18520 -1605
rect 18480 -1640 18520 -1625
rect 18535 -1555 18575 -1540
rect 18535 -1575 18545 -1555
rect 18565 -1575 18575 -1555
rect 18535 -1605 18575 -1575
rect 18535 -1625 18545 -1605
rect 18565 -1625 18575 -1605
rect 18535 -1640 18575 -1625
<< pdiff >>
rect 16375 1415 16415 1430
rect 16375 1395 16385 1415
rect 16405 1395 16415 1415
rect 16375 1365 16415 1395
rect 16375 1345 16385 1365
rect 16405 1345 16415 1365
rect 16375 1330 16415 1345
rect 16430 1415 16470 1430
rect 16430 1395 16440 1415
rect 16460 1395 16470 1415
rect 16430 1365 16470 1395
rect 16430 1345 16440 1365
rect 16460 1345 16470 1365
rect 16430 1330 16470 1345
rect 16485 1415 16525 1430
rect 16485 1395 16495 1415
rect 16515 1395 16525 1415
rect 16485 1365 16525 1395
rect 16485 1345 16495 1365
rect 16515 1345 16525 1365
rect 16485 1330 16525 1345
rect 16540 1415 16580 1430
rect 16540 1395 16550 1415
rect 16570 1395 16580 1415
rect 16540 1365 16580 1395
rect 16540 1345 16550 1365
rect 16570 1345 16580 1365
rect 16540 1330 16580 1345
rect 16595 1415 16635 1430
rect 16595 1395 16605 1415
rect 16625 1395 16635 1415
rect 16595 1365 16635 1395
rect 16595 1345 16605 1365
rect 16625 1345 16635 1365
rect 16595 1330 16635 1345
rect 16885 1415 16925 1430
rect 16885 1343 16895 1415
rect 16915 1343 16925 1415
rect 16885 1330 16925 1343
rect 16940 1415 16980 1430
rect 16940 1343 16950 1415
rect 16970 1343 16980 1415
rect 16940 1330 16980 1343
rect 16995 1415 17035 1430
rect 16995 1343 17005 1415
rect 17025 1343 17035 1415
rect 16995 1330 17035 1343
rect 17050 1415 17090 1430
rect 17050 1343 17060 1415
rect 17080 1343 17090 1415
rect 17050 1330 17090 1343
rect 17105 1415 17145 1430
rect 17105 1343 17115 1415
rect 17135 1343 17145 1415
rect 17105 1330 17145 1343
rect 17160 1415 17200 1430
rect 17160 1343 17170 1415
rect 17190 1343 17200 1415
rect 17160 1330 17200 1343
rect 17215 1415 17255 1430
rect 17215 1343 17225 1415
rect 17245 1343 17255 1415
rect 17215 1330 17255 1343
rect 17505 1415 17545 1430
rect 17505 1395 17515 1415
rect 17535 1395 17545 1415
rect 17505 1365 17545 1395
rect 17505 1345 17515 1365
rect 17535 1345 17545 1365
rect 17505 1330 17545 1345
rect 17560 1415 17600 1430
rect 17560 1395 17570 1415
rect 17590 1395 17600 1415
rect 17560 1365 17600 1395
rect 17560 1345 17570 1365
rect 17590 1345 17600 1365
rect 17560 1330 17600 1345
rect 17615 1415 17655 1430
rect 17615 1395 17625 1415
rect 17645 1395 17655 1415
rect 17615 1365 17655 1395
rect 17615 1345 17625 1365
rect 17645 1345 17655 1365
rect 17615 1330 17655 1345
rect 17670 1415 17710 1430
rect 17670 1395 17680 1415
rect 17700 1395 17710 1415
rect 17670 1365 17710 1395
rect 17670 1345 17680 1365
rect 17700 1345 17710 1365
rect 17670 1330 17710 1345
rect 17725 1415 17765 1430
rect 17725 1395 17735 1415
rect 17755 1395 17765 1415
rect 17725 1365 17765 1395
rect 17725 1345 17735 1365
rect 17755 1345 17765 1365
rect 17725 1330 17765 1345
rect 17780 1415 17820 1430
rect 17780 1395 17790 1415
rect 17810 1395 17820 1415
rect 17780 1365 17820 1395
rect 17780 1345 17790 1365
rect 17810 1345 17820 1365
rect 17780 1330 17820 1345
rect 17835 1415 17875 1430
rect 17835 1395 17845 1415
rect 17865 1395 17875 1415
rect 17835 1365 17875 1395
rect 17835 1345 17845 1365
rect 17865 1345 17875 1365
rect 17835 1330 17875 1345
rect 17890 1415 17930 1430
rect 17890 1395 17900 1415
rect 17920 1395 17930 1415
rect 17890 1365 17930 1395
rect 17890 1345 17900 1365
rect 17920 1345 17930 1365
rect 17890 1330 17930 1345
rect 17945 1415 17985 1430
rect 17945 1395 17955 1415
rect 17975 1395 17985 1415
rect 17945 1365 17985 1395
rect 17945 1345 17955 1365
rect 17975 1345 17985 1365
rect 17945 1330 17985 1345
rect 18000 1415 18040 1430
rect 18000 1395 18010 1415
rect 18030 1395 18040 1415
rect 18000 1365 18040 1395
rect 18000 1345 18010 1365
rect 18030 1345 18040 1365
rect 18000 1330 18040 1345
rect 18055 1415 18095 1430
rect 18055 1395 18065 1415
rect 18085 1395 18095 1415
rect 18055 1365 18095 1395
rect 18055 1345 18065 1365
rect 18085 1345 18095 1365
rect 18055 1330 18095 1345
rect 18345 1415 18385 1430
rect 18345 1345 18355 1415
rect 18375 1345 18385 1415
rect 18345 1330 18385 1345
rect 18400 1415 18440 1430
rect 18400 1345 18410 1415
rect 18430 1345 18440 1415
rect 18400 1330 18440 1345
rect 18455 1415 18495 1430
rect 18455 1345 18465 1415
rect 18485 1345 18495 1415
rect 18455 1330 18495 1345
rect 18510 1415 18550 1430
rect 18510 1345 18520 1415
rect 18540 1345 18550 1415
rect 18510 1330 18550 1345
rect 18565 1415 18605 1430
rect 18565 1345 18575 1415
rect 18595 1345 18605 1415
rect 18565 1330 18605 1345
rect 18620 1415 18660 1430
rect 18620 1345 18630 1415
rect 18650 1345 18660 1415
rect 18620 1330 18660 1345
rect 18675 1415 18715 1430
rect 18675 1345 18685 1415
rect 18705 1345 18715 1415
rect 18675 1330 18715 1345
rect 16970 950 17010 965
rect 16970 930 16980 950
rect 17000 930 17010 950
rect 16970 900 17010 930
rect 16970 880 16980 900
rect 17000 880 17010 900
rect 16435 850 16475 865
rect 16435 830 16445 850
rect 16465 830 16475 850
rect 16435 800 16475 830
rect 16435 780 16445 800
rect 16465 780 16475 800
rect 16435 765 16475 780
rect 16490 850 16530 865
rect 16490 830 16500 850
rect 16520 830 16530 850
rect 16490 800 16530 830
rect 16490 780 16500 800
rect 16520 780 16530 800
rect 16490 765 16530 780
rect 16545 850 16585 865
rect 16545 830 16555 850
rect 16575 830 16585 850
rect 16545 800 16585 830
rect 16545 780 16555 800
rect 16575 780 16585 800
rect 16545 765 16585 780
rect 16600 850 16640 865
rect 16600 830 16610 850
rect 16630 830 16640 850
rect 16600 800 16640 830
rect 16600 780 16610 800
rect 16630 780 16640 800
rect 16600 765 16640 780
rect 16655 850 16700 865
rect 16655 830 16665 850
rect 16685 830 16700 850
rect 16655 800 16700 830
rect 16655 780 16665 800
rect 16685 780 16700 800
rect 16655 765 16700 780
rect 16970 850 17010 880
rect 16970 830 16980 850
rect 17000 830 17010 850
rect 16970 800 17010 830
rect 16970 780 16980 800
rect 17000 780 17010 800
rect 16970 750 17010 780
rect 16970 730 16980 750
rect 17000 730 17010 750
rect 16970 700 17010 730
rect 16970 680 16980 700
rect 17000 680 17010 700
rect 16970 665 17010 680
rect 17060 950 17100 965
rect 17060 930 17070 950
rect 17090 930 17100 950
rect 17060 900 17100 930
rect 17060 880 17070 900
rect 17090 880 17100 900
rect 17060 850 17100 880
rect 17060 830 17070 850
rect 17090 830 17100 850
rect 17060 800 17100 830
rect 17060 780 17070 800
rect 17090 780 17100 800
rect 17060 750 17100 780
rect 17060 730 17070 750
rect 17090 730 17100 750
rect 17060 700 17100 730
rect 17060 680 17070 700
rect 17090 680 17100 700
rect 17060 665 17100 680
rect 17150 950 17190 965
rect 17150 930 17160 950
rect 17180 930 17190 950
rect 17150 900 17190 930
rect 17150 880 17160 900
rect 17180 880 17190 900
rect 17150 850 17190 880
rect 17150 830 17160 850
rect 17180 830 17190 850
rect 17150 800 17190 830
rect 17150 780 17160 800
rect 17180 780 17190 800
rect 17150 750 17190 780
rect 17150 730 17160 750
rect 17180 730 17190 750
rect 17150 700 17190 730
rect 17150 680 17160 700
rect 17180 680 17190 700
rect 17150 665 17190 680
rect 17240 950 17280 965
rect 17240 930 17250 950
rect 17270 930 17280 950
rect 17240 900 17280 930
rect 17240 880 17250 900
rect 17270 880 17280 900
rect 17240 850 17280 880
rect 17240 830 17250 850
rect 17270 830 17280 850
rect 17240 800 17280 830
rect 17240 780 17250 800
rect 17270 780 17280 800
rect 17240 750 17280 780
rect 17240 730 17250 750
rect 17270 730 17280 750
rect 17240 700 17280 730
rect 17240 680 17250 700
rect 17270 680 17280 700
rect 17240 665 17280 680
rect 17330 950 17370 965
rect 17330 930 17340 950
rect 17360 930 17370 950
rect 17330 900 17370 930
rect 17330 880 17340 900
rect 17360 880 17370 900
rect 17330 850 17370 880
rect 17330 830 17340 850
rect 17360 830 17370 850
rect 17330 800 17370 830
rect 17330 780 17340 800
rect 17360 780 17370 800
rect 17330 750 17370 780
rect 17330 730 17340 750
rect 17360 730 17370 750
rect 17330 700 17370 730
rect 17330 680 17340 700
rect 17360 680 17370 700
rect 17330 665 17370 680
rect 17420 950 17460 965
rect 17420 930 17430 950
rect 17450 930 17460 950
rect 17420 900 17460 930
rect 17420 880 17430 900
rect 17450 880 17460 900
rect 17420 850 17460 880
rect 17420 830 17430 850
rect 17450 830 17460 850
rect 17420 800 17460 830
rect 17420 780 17430 800
rect 17450 780 17460 800
rect 17420 750 17460 780
rect 17420 730 17430 750
rect 17450 730 17460 750
rect 17420 700 17460 730
rect 17420 680 17430 700
rect 17450 680 17460 700
rect 17420 665 17460 680
rect 17510 950 17550 965
rect 17510 930 17520 950
rect 17540 930 17550 950
rect 17510 900 17550 930
rect 17510 880 17520 900
rect 17540 880 17550 900
rect 17510 850 17550 880
rect 17510 830 17520 850
rect 17540 830 17550 850
rect 17510 800 17550 830
rect 17510 780 17520 800
rect 17540 780 17550 800
rect 17510 750 17550 780
rect 17510 730 17520 750
rect 17540 730 17550 750
rect 17510 700 17550 730
rect 17510 680 17520 700
rect 17540 680 17550 700
rect 17510 665 17550 680
rect 17600 950 17640 965
rect 17600 930 17610 950
rect 17630 930 17640 950
rect 17600 900 17640 930
rect 17600 880 17610 900
rect 17630 880 17640 900
rect 17600 850 17640 880
rect 17600 830 17610 850
rect 17630 830 17640 850
rect 17600 800 17640 830
rect 17600 780 17610 800
rect 17630 780 17640 800
rect 17600 750 17640 780
rect 17600 730 17610 750
rect 17630 730 17640 750
rect 17600 700 17640 730
rect 17600 680 17610 700
rect 17630 680 17640 700
rect 17600 665 17640 680
rect 17690 950 17730 965
rect 17690 930 17700 950
rect 17720 930 17730 950
rect 17690 900 17730 930
rect 17690 880 17700 900
rect 17720 880 17730 900
rect 17690 850 17730 880
rect 17690 830 17700 850
rect 17720 830 17730 850
rect 17690 800 17730 830
rect 17690 780 17700 800
rect 17720 780 17730 800
rect 17690 750 17730 780
rect 17690 730 17700 750
rect 17720 730 17730 750
rect 17690 700 17730 730
rect 17690 680 17700 700
rect 17720 680 17730 700
rect 17690 665 17730 680
rect 17780 950 17820 965
rect 17780 930 17790 950
rect 17810 930 17820 950
rect 17780 900 17820 930
rect 17780 880 17790 900
rect 17810 880 17820 900
rect 17780 850 17820 880
rect 17780 830 17790 850
rect 17810 830 17820 850
rect 17780 800 17820 830
rect 17780 780 17790 800
rect 17810 780 17820 800
rect 17780 750 17820 780
rect 17780 730 17790 750
rect 17810 730 17820 750
rect 17780 700 17820 730
rect 17780 680 17790 700
rect 17810 680 17820 700
rect 17780 665 17820 680
rect 17870 950 17910 965
rect 17870 930 17880 950
rect 17900 930 17910 950
rect 17870 900 17910 930
rect 17870 880 17880 900
rect 17900 880 17910 900
rect 17870 850 17910 880
rect 17870 830 17880 850
rect 17900 830 17910 850
rect 17870 800 17910 830
rect 17870 780 17880 800
rect 17900 780 17910 800
rect 17870 750 17910 780
rect 17870 730 17880 750
rect 17900 730 17910 750
rect 17870 700 17910 730
rect 17870 680 17880 700
rect 17900 680 17910 700
rect 17870 665 17910 680
rect 17960 950 18000 965
rect 17960 930 17970 950
rect 17990 930 18000 950
rect 17960 900 18000 930
rect 17960 880 17970 900
rect 17990 880 18000 900
rect 17960 850 18000 880
rect 17960 830 17970 850
rect 17990 830 18000 850
rect 17960 800 18000 830
rect 17960 780 17970 800
rect 17990 780 18000 800
rect 17960 750 18000 780
rect 17960 730 17970 750
rect 17990 730 18000 750
rect 17960 700 18000 730
rect 17960 680 17970 700
rect 17990 680 18000 700
rect 17960 665 18000 680
rect 18050 950 18090 965
rect 18050 930 18060 950
rect 18080 930 18090 950
rect 18050 900 18090 930
rect 18050 880 18060 900
rect 18080 880 18090 900
rect 18050 850 18090 880
rect 18050 830 18060 850
rect 18080 830 18090 850
rect 18050 800 18090 830
rect 18050 780 18060 800
rect 18080 780 18090 800
rect 18050 750 18090 780
rect 18050 730 18060 750
rect 18080 730 18090 750
rect 18050 700 18090 730
rect 18050 680 18060 700
rect 18080 680 18090 700
rect 18050 665 18090 680
rect 18140 950 18180 965
rect 18140 930 18150 950
rect 18170 930 18180 950
rect 18140 900 18180 930
rect 18140 880 18150 900
rect 18170 880 18180 900
rect 18140 850 18180 880
rect 18140 830 18150 850
rect 18170 830 18180 850
rect 18140 800 18180 830
rect 18140 780 18150 800
rect 18170 780 18180 800
rect 18140 750 18180 780
rect 18140 730 18150 750
rect 18170 730 18180 750
rect 18140 700 18180 730
rect 18140 680 18150 700
rect 18170 680 18180 700
rect 18140 665 18180 680
rect 18230 950 18270 965
rect 18230 930 18240 950
rect 18260 930 18270 950
rect 18230 900 18270 930
rect 18230 880 18240 900
rect 18260 880 18270 900
rect 18230 850 18270 880
rect 18230 830 18240 850
rect 18260 830 18270 850
rect 18230 800 18270 830
rect 18230 780 18240 800
rect 18260 780 18270 800
rect 18230 750 18270 780
rect 18230 730 18240 750
rect 18260 730 18270 750
rect 18230 700 18270 730
rect 18230 680 18240 700
rect 18260 680 18270 700
rect 18230 665 18270 680
rect 18320 950 18360 965
rect 18320 930 18330 950
rect 18350 930 18360 950
rect 18320 900 18360 930
rect 18320 880 18330 900
rect 18350 880 18360 900
rect 18320 850 18360 880
rect 18320 830 18330 850
rect 18350 830 18360 850
rect 18320 800 18360 830
rect 18320 780 18330 800
rect 18350 780 18360 800
rect 18320 750 18360 780
rect 18320 730 18330 750
rect 18350 730 18360 750
rect 18320 700 18360 730
rect 18320 680 18330 700
rect 18350 680 18360 700
rect 18320 665 18360 680
rect 18410 950 18450 965
rect 18410 930 18420 950
rect 18440 930 18450 950
rect 18410 900 18450 930
rect 18410 880 18420 900
rect 18440 880 18450 900
rect 18410 850 18450 880
rect 18410 830 18420 850
rect 18440 830 18450 850
rect 18410 800 18450 830
rect 18410 780 18420 800
rect 18440 780 18450 800
rect 18410 750 18450 780
rect 18410 730 18420 750
rect 18440 730 18450 750
rect 18410 700 18450 730
rect 18410 680 18420 700
rect 18440 680 18450 700
rect 18410 665 18450 680
rect 18500 950 18540 965
rect 18500 930 18510 950
rect 18530 930 18540 950
rect 18500 900 18540 930
rect 18500 880 18510 900
rect 18530 880 18540 900
rect 18500 850 18540 880
rect 18500 830 18510 850
rect 18530 830 18540 850
rect 18500 800 18540 830
rect 18500 780 18510 800
rect 18530 780 18540 800
rect 18500 750 18540 780
rect 18500 730 18510 750
rect 18530 730 18540 750
rect 18500 700 18540 730
rect 18500 680 18510 700
rect 18530 680 18540 700
rect 18500 665 18540 680
rect 18590 950 18630 965
rect 18590 930 18600 950
rect 18620 930 18630 950
rect 18590 900 18630 930
rect 18590 880 18600 900
rect 18620 880 18630 900
rect 18590 850 18630 880
rect 18590 830 18600 850
rect 18620 830 18630 850
rect 18590 800 18630 830
rect 18590 780 18600 800
rect 18620 780 18630 800
rect 18590 750 18630 780
rect 18905 950 18945 965
rect 18905 930 18915 950
rect 18935 930 18945 950
rect 18905 900 18945 930
rect 18905 880 18915 900
rect 18935 880 18945 900
rect 18905 850 18945 880
rect 18905 830 18915 850
rect 18935 830 18945 850
rect 18905 800 18945 830
rect 18905 780 18915 800
rect 18935 780 18945 800
rect 18905 765 18945 780
rect 18960 950 19000 965
rect 18960 930 18970 950
rect 18990 930 19000 950
rect 18960 900 19000 930
rect 18960 880 18970 900
rect 18990 880 19000 900
rect 18960 850 19000 880
rect 18960 830 18970 850
rect 18990 830 19000 850
rect 18960 800 19000 830
rect 18960 780 18970 800
rect 18990 780 19000 800
rect 18960 765 19000 780
rect 19015 950 19055 965
rect 19015 930 19025 950
rect 19045 930 19055 950
rect 19015 900 19055 930
rect 19015 880 19025 900
rect 19045 880 19055 900
rect 19015 850 19055 880
rect 19015 830 19025 850
rect 19045 830 19055 850
rect 19015 800 19055 830
rect 19015 780 19025 800
rect 19045 780 19055 800
rect 19015 765 19055 780
rect 19070 950 19110 965
rect 19070 930 19080 950
rect 19100 930 19110 950
rect 19070 900 19110 930
rect 19070 880 19080 900
rect 19100 880 19110 900
rect 19070 850 19110 880
rect 19070 830 19080 850
rect 19100 830 19110 850
rect 19070 800 19110 830
rect 19070 780 19080 800
rect 19100 780 19110 800
rect 19070 765 19110 780
rect 18590 730 18600 750
rect 18620 730 18630 750
rect 18590 700 18630 730
rect 18590 680 18600 700
rect 18620 680 18630 700
rect 18590 665 18630 680
rect 16420 110 16460 125
rect 16420 90 16430 110
rect 16450 90 16460 110
rect 16420 60 16460 90
rect 16420 40 16430 60
rect 16450 40 16460 60
rect 16420 25 16460 40
rect 16480 110 16520 125
rect 16480 90 16490 110
rect 16510 90 16520 110
rect 16480 60 16520 90
rect 16480 40 16490 60
rect 16510 40 16520 60
rect 16480 25 16520 40
rect 16540 110 16580 125
rect 16540 90 16550 110
rect 16570 90 16580 110
rect 16540 60 16580 90
rect 16540 40 16550 60
rect 16570 40 16580 60
rect 16540 25 16580 40
rect 16600 110 16640 125
rect 16600 90 16610 110
rect 16630 90 16640 110
rect 16600 60 16640 90
rect 16600 40 16610 60
rect 16630 40 16640 60
rect 16600 25 16640 40
rect 16660 110 16700 125
rect 16660 90 16670 110
rect 16690 90 16700 110
rect 16660 60 16700 90
rect 16660 40 16670 60
rect 16690 40 16700 60
rect 16660 25 16700 40
rect 16720 110 16760 125
rect 16720 90 16730 110
rect 16750 90 16760 110
rect 16720 60 16760 90
rect 16720 40 16730 60
rect 16750 40 16760 60
rect 16720 25 16760 40
rect 16780 110 16820 125
rect 16780 90 16790 110
rect 16810 90 16820 110
rect 16780 60 16820 90
rect 16780 40 16790 60
rect 16810 40 16820 60
rect 16780 25 16820 40
rect 16840 110 16880 125
rect 16840 90 16850 110
rect 16870 90 16880 110
rect 16840 60 16880 90
rect 16840 40 16850 60
rect 16870 40 16880 60
rect 16840 25 16880 40
rect 16900 110 16940 125
rect 16900 90 16910 110
rect 16930 90 16940 110
rect 16900 60 16940 90
rect 16900 40 16910 60
rect 16930 40 16940 60
rect 16900 25 16940 40
rect 16960 110 17000 125
rect 16960 90 16970 110
rect 16990 90 17000 110
rect 16960 60 17000 90
rect 16960 40 16970 60
rect 16990 40 17000 60
rect 16960 25 17000 40
rect 17020 110 17060 125
rect 17020 90 17030 110
rect 17050 90 17060 110
rect 17020 60 17060 90
rect 17020 40 17030 60
rect 17050 40 17060 60
rect 17020 25 17060 40
rect 17080 110 17120 125
rect 17080 90 17090 110
rect 17110 90 17120 110
rect 17080 60 17120 90
rect 17080 40 17090 60
rect 17110 40 17120 60
rect 17080 25 17120 40
rect 17140 110 17180 125
rect 17140 90 17150 110
rect 17170 90 17180 110
rect 17140 60 17180 90
rect 17140 40 17150 60
rect 17170 40 17180 60
rect 17140 25 17180 40
rect 17200 110 17240 125
rect 17200 90 17210 110
rect 17230 90 17240 110
rect 17200 60 17240 90
rect 17200 40 17210 60
rect 17230 40 17240 60
rect 17200 25 17240 40
rect 17260 110 17300 125
rect 17260 90 17270 110
rect 17290 90 17300 110
rect 17260 60 17300 90
rect 17260 40 17270 60
rect 17290 40 17300 60
rect 17260 25 17300 40
rect 17320 110 17360 125
rect 17320 90 17330 110
rect 17350 90 17360 110
rect 17320 60 17360 90
rect 17320 40 17330 60
rect 17350 40 17360 60
rect 17320 25 17360 40
rect 17380 110 17420 125
rect 17380 90 17390 110
rect 17410 90 17420 110
rect 17380 60 17420 90
rect 17380 40 17390 60
rect 17410 40 17420 60
rect 17380 25 17420 40
rect 17440 110 17480 125
rect 17440 90 17450 110
rect 17470 90 17480 110
rect 17440 60 17480 90
rect 17440 40 17450 60
rect 17470 40 17480 60
rect 17440 25 17480 40
rect 17500 110 17540 125
rect 17500 90 17510 110
rect 17530 90 17540 110
rect 17500 60 17540 90
rect 17500 40 17510 60
rect 17530 40 17540 60
rect 17500 25 17540 40
rect 17560 110 17600 125
rect 17560 90 17570 110
rect 17590 90 17600 110
rect 17560 60 17600 90
rect 17560 40 17570 60
rect 17590 40 17600 60
rect 17560 25 17600 40
rect 17620 110 17660 125
rect 17620 90 17630 110
rect 17650 90 17660 110
rect 17620 60 17660 90
rect 17620 40 17630 60
rect 17650 40 17660 60
rect 17620 25 17660 40
rect 17940 110 17980 125
rect 17940 90 17950 110
rect 17970 90 17980 110
rect 17940 60 17980 90
rect 17940 40 17950 60
rect 17970 40 17980 60
rect 17940 25 17980 40
rect 18000 110 18040 125
rect 18000 90 18010 110
rect 18030 90 18040 110
rect 18000 60 18040 90
rect 18000 40 18010 60
rect 18030 40 18040 60
rect 18000 25 18040 40
rect 18060 110 18100 125
rect 18060 90 18070 110
rect 18090 90 18100 110
rect 18060 60 18100 90
rect 18060 40 18070 60
rect 18090 40 18100 60
rect 18060 25 18100 40
rect 18120 110 18160 125
rect 18120 90 18130 110
rect 18150 90 18160 110
rect 18120 60 18160 90
rect 18120 40 18130 60
rect 18150 40 18160 60
rect 18120 25 18160 40
rect 18180 110 18220 125
rect 18180 90 18190 110
rect 18210 90 18220 110
rect 18180 60 18220 90
rect 18180 40 18190 60
rect 18210 40 18220 60
rect 18180 25 18220 40
rect 18240 110 18280 125
rect 18240 90 18250 110
rect 18270 90 18280 110
rect 18240 60 18280 90
rect 18240 40 18250 60
rect 18270 40 18280 60
rect 18240 25 18280 40
rect 18300 110 18340 125
rect 18300 90 18310 110
rect 18330 90 18340 110
rect 18300 60 18340 90
rect 18300 40 18310 60
rect 18330 40 18340 60
rect 18300 25 18340 40
rect 18360 110 18400 125
rect 18360 90 18370 110
rect 18390 90 18400 110
rect 18360 60 18400 90
rect 18360 40 18370 60
rect 18390 40 18400 60
rect 18360 25 18400 40
rect 18420 110 18460 125
rect 18420 90 18430 110
rect 18450 90 18460 110
rect 18420 60 18460 90
rect 18420 40 18430 60
rect 18450 40 18460 60
rect 18420 25 18460 40
rect 18480 110 18520 125
rect 18480 90 18490 110
rect 18510 90 18520 110
rect 18480 60 18520 90
rect 18480 40 18490 60
rect 18510 40 18520 60
rect 18480 25 18520 40
rect 18540 110 18580 125
rect 18540 90 18550 110
rect 18570 90 18580 110
rect 18540 60 18580 90
rect 18540 40 18550 60
rect 18570 40 18580 60
rect 18540 25 18580 40
rect 18600 110 18640 125
rect 18600 90 18610 110
rect 18630 90 18640 110
rect 18600 60 18640 90
rect 18600 40 18610 60
rect 18630 40 18640 60
rect 18600 25 18640 40
rect 18660 110 18700 125
rect 18660 90 18670 110
rect 18690 90 18700 110
rect 18660 60 18700 90
rect 18660 40 18670 60
rect 18690 40 18700 60
rect 18660 25 18700 40
rect 18720 110 18760 125
rect 18720 90 18730 110
rect 18750 90 18760 110
rect 18720 60 18760 90
rect 18720 40 18730 60
rect 18750 40 18760 60
rect 18720 25 18760 40
rect 18780 110 18820 125
rect 18780 90 18790 110
rect 18810 90 18820 110
rect 18780 60 18820 90
rect 18780 40 18790 60
rect 18810 40 18820 60
rect 18780 25 18820 40
rect 18840 110 18880 125
rect 18840 90 18850 110
rect 18870 90 18880 110
rect 18840 60 18880 90
rect 18840 40 18850 60
rect 18870 40 18880 60
rect 18840 25 18880 40
rect 18900 110 18940 125
rect 18900 90 18910 110
rect 18930 90 18940 110
rect 18900 60 18940 90
rect 18900 40 18910 60
rect 18930 40 18940 60
rect 18900 25 18940 40
rect 18960 110 19000 125
rect 18960 90 18970 110
rect 18990 90 19000 110
rect 18960 60 19000 90
rect 18960 40 18970 60
rect 18990 40 19000 60
rect 18960 25 19000 40
rect 19020 110 19060 125
rect 19020 90 19030 110
rect 19050 90 19060 110
rect 19020 60 19060 90
rect 19020 40 19030 60
rect 19050 40 19060 60
rect 19020 25 19060 40
rect 19080 110 19120 125
rect 19080 90 19090 110
rect 19110 90 19120 110
rect 19080 60 19120 90
rect 19080 40 19090 60
rect 19110 40 19120 60
rect 19080 25 19120 40
rect 19140 110 19180 125
rect 19140 90 19150 110
rect 19170 90 19180 110
rect 19140 60 19180 90
rect 19140 40 19150 60
rect 19170 40 19180 60
rect 19140 25 19180 40
<< ndiffc >>
rect 16970 -195 16990 -175
rect 16970 -245 16990 -225
rect 16970 -295 16990 -275
rect 16970 -345 16990 -325
rect 16970 -395 16990 -375
rect 17030 -195 17050 -175
rect 17030 -245 17050 -225
rect 17030 -295 17050 -275
rect 17030 -345 17050 -325
rect 17030 -395 17050 -375
rect 17090 -195 17110 -175
rect 17090 -245 17110 -225
rect 17090 -295 17110 -275
rect 18490 -195 18510 -175
rect 18490 -245 18510 -225
rect 17090 -345 17110 -325
rect 17090 -395 17110 -375
rect 18490 -295 18510 -275
rect 18490 -345 18510 -325
rect 18490 -395 18510 -375
rect 18550 -195 18570 -175
rect 18550 -245 18570 -225
rect 18550 -295 18570 -275
rect 18550 -345 18570 -325
rect 18550 -395 18570 -375
rect 18610 -195 18630 -175
rect 18610 -245 18630 -225
rect 18610 -295 18630 -275
rect 18610 -345 18630 -325
rect 18610 -395 18630 -375
rect 16540 -730 16560 -710
rect 16540 -780 16560 -760
rect 16540 -830 16560 -810
rect 16540 -880 16560 -860
rect 16540 -930 16560 -910
rect 17080 -730 17100 -710
rect 17160 -730 17180 -710
rect 17080 -780 17100 -760
rect 17160 -780 17180 -760
rect 17080 -830 17100 -810
rect 17160 -830 17180 -810
rect 17080 -880 17100 -860
rect 17160 -880 17180 -860
rect 17080 -930 17100 -910
rect 17160 -930 17180 -910
rect 17700 -730 17720 -710
rect 17700 -780 17720 -760
rect 17700 -830 17720 -810
rect 17700 -880 17720 -860
rect 17700 -930 17720 -910
rect 17880 -730 17900 -710
rect 17880 -780 17900 -760
rect 17880 -830 17900 -810
rect 17880 -880 17900 -860
rect 17880 -930 17900 -910
rect 18420 -730 18440 -710
rect 18500 -730 18520 -710
rect 18420 -780 18440 -760
rect 18500 -780 18520 -760
rect 18420 -830 18440 -810
rect 18500 -830 18520 -810
rect 18420 -880 18440 -860
rect 18500 -880 18520 -860
rect 18420 -930 18440 -910
rect 18500 -930 18520 -910
rect 19040 -730 19060 -710
rect 19040 -780 19060 -760
rect 19040 -830 19060 -810
rect 19040 -880 19060 -860
rect 19040 -930 19060 -910
rect 16750 -1185 16770 -1165
rect 16750 -1235 16770 -1215
rect 17790 -1185 17810 -1165
rect 17790 -1235 17810 -1215
rect 18830 -1185 18850 -1165
rect 18830 -1235 18850 -1215
rect 16610 -1575 16630 -1555
rect 16610 -1625 16630 -1605
rect 16665 -1575 16685 -1555
rect 16665 -1625 16685 -1605
rect 16720 -1575 16740 -1555
rect 16720 -1625 16740 -1605
rect 16775 -1575 16795 -1555
rect 16775 -1625 16795 -1605
rect 16830 -1575 16850 -1555
rect 16830 -1625 16850 -1605
rect 16885 -1575 16905 -1555
rect 16885 -1625 16905 -1605
rect 17035 -1575 17055 -1555
rect 17035 -1625 17055 -1605
rect 17090 -1575 17110 -1555
rect 17090 -1625 17110 -1605
rect 17145 -1575 17165 -1555
rect 17145 -1625 17165 -1605
rect 17200 -1575 17220 -1555
rect 17200 -1625 17220 -1605
rect 17255 -1575 17275 -1555
rect 17255 -1625 17275 -1605
rect 17310 -1575 17330 -1555
rect 17310 -1625 17330 -1605
rect 17365 -1575 17385 -1555
rect 17365 -1625 17385 -1605
rect 17420 -1575 17440 -1555
rect 17420 -1625 17440 -1605
rect 17475 -1575 17495 -1555
rect 17475 -1625 17495 -1605
rect 17625 -1575 17645 -1555
rect 17625 -1625 17645 -1605
rect 17680 -1575 17700 -1555
rect 17680 -1625 17700 -1605
rect 17735 -1575 17755 -1555
rect 17735 -1625 17755 -1605
rect 17790 -1575 17810 -1555
rect 17790 -1625 17810 -1605
rect 17845 -1575 17865 -1555
rect 17845 -1625 17865 -1605
rect 17900 -1575 17920 -1555
rect 17900 -1625 17920 -1605
rect 17955 -1575 17975 -1555
rect 17955 -1625 17975 -1605
rect 18105 -1575 18125 -1555
rect 18105 -1625 18125 -1605
rect 18160 -1575 18180 -1555
rect 18160 -1625 18180 -1605
rect 18215 -1575 18235 -1555
rect 18215 -1625 18235 -1605
rect 18270 -1575 18290 -1555
rect 18270 -1625 18290 -1605
rect 18325 -1575 18345 -1555
rect 18325 -1625 18345 -1605
rect 18380 -1575 18400 -1555
rect 18380 -1625 18400 -1605
rect 18435 -1575 18455 -1555
rect 18435 -1625 18455 -1605
rect 18490 -1575 18510 -1555
rect 18490 -1625 18510 -1605
rect 18545 -1575 18565 -1555
rect 18545 -1625 18565 -1605
<< pdiffc >>
rect 16385 1395 16405 1415
rect 16385 1345 16405 1365
rect 16440 1395 16460 1415
rect 16440 1345 16460 1365
rect 16495 1395 16515 1415
rect 16495 1345 16515 1365
rect 16550 1395 16570 1415
rect 16550 1345 16570 1365
rect 16605 1395 16625 1415
rect 16605 1345 16625 1365
rect 16895 1343 16915 1415
rect 16950 1343 16970 1415
rect 17005 1343 17025 1415
rect 17060 1343 17080 1415
rect 17115 1343 17135 1415
rect 17170 1343 17190 1415
rect 17225 1343 17245 1415
rect 17515 1395 17535 1415
rect 17515 1345 17535 1365
rect 17570 1395 17590 1415
rect 17570 1345 17590 1365
rect 17625 1395 17645 1415
rect 17625 1345 17645 1365
rect 17680 1395 17700 1415
rect 17680 1345 17700 1365
rect 17735 1395 17755 1415
rect 17735 1345 17755 1365
rect 17790 1395 17810 1415
rect 17790 1345 17810 1365
rect 17845 1395 17865 1415
rect 17845 1345 17865 1365
rect 17900 1395 17920 1415
rect 17900 1345 17920 1365
rect 17955 1395 17975 1415
rect 17955 1345 17975 1365
rect 18010 1395 18030 1415
rect 18010 1345 18030 1365
rect 18065 1395 18085 1415
rect 18065 1345 18085 1365
rect 18355 1345 18375 1415
rect 18410 1345 18430 1415
rect 18465 1345 18485 1415
rect 18520 1345 18540 1415
rect 18575 1345 18595 1415
rect 18630 1345 18650 1415
rect 18685 1345 18705 1415
rect 16980 930 17000 950
rect 16980 880 17000 900
rect 16445 830 16465 850
rect 16445 780 16465 800
rect 16500 830 16520 850
rect 16500 780 16520 800
rect 16555 830 16575 850
rect 16555 780 16575 800
rect 16610 830 16630 850
rect 16610 780 16630 800
rect 16665 830 16685 850
rect 16665 780 16685 800
rect 16980 830 17000 850
rect 16980 780 17000 800
rect 16980 730 17000 750
rect 16980 680 17000 700
rect 17070 930 17090 950
rect 17070 880 17090 900
rect 17070 830 17090 850
rect 17070 780 17090 800
rect 17070 730 17090 750
rect 17070 680 17090 700
rect 17160 930 17180 950
rect 17160 880 17180 900
rect 17160 830 17180 850
rect 17160 780 17180 800
rect 17160 730 17180 750
rect 17160 680 17180 700
rect 17250 930 17270 950
rect 17250 880 17270 900
rect 17250 830 17270 850
rect 17250 780 17270 800
rect 17250 730 17270 750
rect 17250 680 17270 700
rect 17340 930 17360 950
rect 17340 880 17360 900
rect 17340 830 17360 850
rect 17340 780 17360 800
rect 17340 730 17360 750
rect 17340 680 17360 700
rect 17430 930 17450 950
rect 17430 880 17450 900
rect 17430 830 17450 850
rect 17430 780 17450 800
rect 17430 730 17450 750
rect 17430 680 17450 700
rect 17520 930 17540 950
rect 17520 880 17540 900
rect 17520 830 17540 850
rect 17520 780 17540 800
rect 17520 730 17540 750
rect 17520 680 17540 700
rect 17610 930 17630 950
rect 17610 880 17630 900
rect 17610 830 17630 850
rect 17610 780 17630 800
rect 17610 730 17630 750
rect 17610 680 17630 700
rect 17700 930 17720 950
rect 17700 880 17720 900
rect 17700 830 17720 850
rect 17700 780 17720 800
rect 17700 730 17720 750
rect 17700 680 17720 700
rect 17790 930 17810 950
rect 17790 880 17810 900
rect 17790 830 17810 850
rect 17790 780 17810 800
rect 17790 730 17810 750
rect 17790 680 17810 700
rect 17880 930 17900 950
rect 17880 880 17900 900
rect 17880 830 17900 850
rect 17880 780 17900 800
rect 17880 730 17900 750
rect 17880 680 17900 700
rect 17970 930 17990 950
rect 17970 880 17990 900
rect 17970 830 17990 850
rect 17970 780 17990 800
rect 17970 730 17990 750
rect 17970 680 17990 700
rect 18060 930 18080 950
rect 18060 880 18080 900
rect 18060 830 18080 850
rect 18060 780 18080 800
rect 18060 730 18080 750
rect 18060 680 18080 700
rect 18150 930 18170 950
rect 18150 880 18170 900
rect 18150 830 18170 850
rect 18150 780 18170 800
rect 18150 730 18170 750
rect 18150 680 18170 700
rect 18240 930 18260 950
rect 18240 880 18260 900
rect 18240 830 18260 850
rect 18240 780 18260 800
rect 18240 730 18260 750
rect 18240 680 18260 700
rect 18330 930 18350 950
rect 18330 880 18350 900
rect 18330 830 18350 850
rect 18330 780 18350 800
rect 18330 730 18350 750
rect 18330 680 18350 700
rect 18420 930 18440 950
rect 18420 880 18440 900
rect 18420 830 18440 850
rect 18420 780 18440 800
rect 18420 730 18440 750
rect 18420 680 18440 700
rect 18510 930 18530 950
rect 18510 880 18530 900
rect 18510 830 18530 850
rect 18510 780 18530 800
rect 18510 730 18530 750
rect 18510 680 18530 700
rect 18600 930 18620 950
rect 18600 880 18620 900
rect 18600 830 18620 850
rect 18600 780 18620 800
rect 18915 930 18935 950
rect 18915 880 18935 900
rect 18915 830 18935 850
rect 18915 780 18935 800
rect 18970 930 18990 950
rect 18970 880 18990 900
rect 18970 830 18990 850
rect 18970 780 18990 800
rect 19025 930 19045 950
rect 19025 880 19045 900
rect 19025 830 19045 850
rect 19025 780 19045 800
rect 19080 930 19100 950
rect 19080 880 19100 900
rect 19080 830 19100 850
rect 19080 780 19100 800
rect 18600 730 18620 750
rect 18600 680 18620 700
rect 16430 90 16450 110
rect 16430 40 16450 60
rect 16490 90 16510 110
rect 16490 40 16510 60
rect 16550 90 16570 110
rect 16550 40 16570 60
rect 16610 90 16630 110
rect 16610 40 16630 60
rect 16670 90 16690 110
rect 16670 40 16690 60
rect 16730 90 16750 110
rect 16730 40 16750 60
rect 16790 90 16810 110
rect 16790 40 16810 60
rect 16850 90 16870 110
rect 16850 40 16870 60
rect 16910 90 16930 110
rect 16910 40 16930 60
rect 16970 90 16990 110
rect 16970 40 16990 60
rect 17030 90 17050 110
rect 17030 40 17050 60
rect 17090 90 17110 110
rect 17090 40 17110 60
rect 17150 90 17170 110
rect 17150 40 17170 60
rect 17210 90 17230 110
rect 17210 40 17230 60
rect 17270 90 17290 110
rect 17270 40 17290 60
rect 17330 90 17350 110
rect 17330 40 17350 60
rect 17390 90 17410 110
rect 17390 40 17410 60
rect 17450 90 17470 110
rect 17450 40 17470 60
rect 17510 90 17530 110
rect 17510 40 17530 60
rect 17570 90 17590 110
rect 17570 40 17590 60
rect 17630 90 17650 110
rect 17630 40 17650 60
rect 17950 90 17970 110
rect 17950 40 17970 60
rect 18010 90 18030 110
rect 18010 40 18030 60
rect 18070 90 18090 110
rect 18070 40 18090 60
rect 18130 90 18150 110
rect 18130 40 18150 60
rect 18190 90 18210 110
rect 18190 40 18210 60
rect 18250 90 18270 110
rect 18250 40 18270 60
rect 18310 90 18330 110
rect 18310 40 18330 60
rect 18370 90 18390 110
rect 18370 40 18390 60
rect 18430 90 18450 110
rect 18430 40 18450 60
rect 18490 90 18510 110
rect 18490 40 18510 60
rect 18550 90 18570 110
rect 18550 40 18570 60
rect 18610 90 18630 110
rect 18610 40 18630 60
rect 18670 90 18690 110
rect 18670 40 18690 60
rect 18730 90 18750 110
rect 18730 40 18750 60
rect 18790 90 18810 110
rect 18790 40 18810 60
rect 18850 90 18870 110
rect 18850 40 18870 60
rect 18910 90 18930 110
rect 18910 40 18930 60
rect 18970 90 18990 110
rect 18970 40 18990 60
rect 19030 90 19050 110
rect 19030 40 19050 60
rect 19090 90 19110 110
rect 19090 40 19110 60
rect 19150 90 19170 110
rect 19150 40 19170 60
<< psubdiff >>
rect 17560 -175 17600 -160
rect 17560 -195 17570 -175
rect 17590 -195 17600 -175
rect 17560 -215 17600 -195
rect 17560 -235 17570 -215
rect 17590 -235 17600 -215
rect 17560 -255 17600 -235
rect 17560 -275 17570 -255
rect 17590 -275 17600 -255
rect 17560 -290 17600 -275
rect 18000 -175 18040 -160
rect 18000 -195 18010 -175
rect 18030 -195 18040 -175
rect 18000 -215 18040 -195
rect 18000 -235 18010 -215
rect 18030 -235 18040 -215
rect 18000 -255 18040 -235
rect 18000 -275 18010 -255
rect 18030 -275 18040 -255
rect 18000 -290 18040 -275
rect 17110 -710 17150 -695
rect 17110 -730 17120 -710
rect 17140 -730 17150 -710
rect 17110 -760 17150 -730
rect 17110 -780 17120 -760
rect 17140 -780 17150 -760
rect 17110 -810 17150 -780
rect 17110 -830 17120 -810
rect 17140 -830 17150 -810
rect 17110 -860 17150 -830
rect 17110 -880 17120 -860
rect 17140 -880 17150 -860
rect 17110 -910 17150 -880
rect 17110 -930 17120 -910
rect 17140 -930 17150 -910
rect 17110 -940 17150 -930
rect 18450 -710 18490 -695
rect 18450 -730 18460 -710
rect 18480 -730 18490 -710
rect 18450 -760 18490 -730
rect 18450 -780 18460 -760
rect 18480 -780 18490 -760
rect 18450 -810 18490 -780
rect 18450 -830 18460 -810
rect 18480 -830 18490 -810
rect 18450 -860 18490 -830
rect 18450 -880 18460 -860
rect 18480 -880 18490 -860
rect 18450 -910 18490 -880
rect 18450 -930 18460 -910
rect 18480 -930 18490 -910
rect 18450 -945 18490 -930
rect 18860 -1165 18900 -1150
rect 18860 -1185 18870 -1165
rect 18890 -1185 18900 -1165
rect 18860 -1215 18900 -1185
rect 18860 -1235 18870 -1215
rect 18890 -1235 18900 -1215
rect 18860 -1250 18900 -1235
rect 16560 -1555 16600 -1540
rect 16560 -1575 16570 -1555
rect 16590 -1575 16600 -1555
rect 16560 -1605 16600 -1575
rect 16560 -1625 16570 -1605
rect 16590 -1625 16600 -1605
rect 16560 -1640 16600 -1625
rect 16915 -1555 16955 -1540
rect 16915 -1575 16925 -1555
rect 16945 -1575 16955 -1555
rect 16915 -1605 16955 -1575
rect 16915 -1625 16925 -1605
rect 16945 -1625 16955 -1605
rect 16915 -1640 16955 -1625
rect 16985 -1555 17025 -1540
rect 16985 -1575 16995 -1555
rect 17015 -1575 17025 -1555
rect 16985 -1605 17025 -1575
rect 16985 -1625 16995 -1605
rect 17015 -1625 17025 -1605
rect 16985 -1640 17025 -1625
rect 17505 -1555 17545 -1540
rect 17505 -1575 17515 -1555
rect 17535 -1575 17545 -1555
rect 17505 -1605 17545 -1575
rect 17505 -1625 17515 -1605
rect 17535 -1625 17545 -1605
rect 17505 -1640 17545 -1625
rect 17575 -1555 17615 -1540
rect 17575 -1575 17585 -1555
rect 17605 -1575 17615 -1555
rect 17575 -1605 17615 -1575
rect 17575 -1625 17585 -1605
rect 17605 -1625 17615 -1605
rect 17575 -1640 17615 -1625
rect 17985 -1555 18025 -1540
rect 17985 -1575 17995 -1555
rect 18015 -1575 18025 -1555
rect 17985 -1605 18025 -1575
rect 17985 -1625 17995 -1605
rect 18015 -1625 18025 -1605
rect 17985 -1640 18025 -1625
rect 18055 -1555 18095 -1540
rect 18055 -1575 18065 -1555
rect 18085 -1575 18095 -1555
rect 18055 -1605 18095 -1575
rect 18055 -1625 18065 -1605
rect 18085 -1625 18095 -1605
rect 18055 -1640 18095 -1625
rect 18575 -1555 18615 -1540
rect 18575 -1575 18585 -1555
rect 18605 -1575 18615 -1555
rect 18575 -1605 18615 -1575
rect 18575 -1625 18585 -1605
rect 18605 -1625 18615 -1605
rect 18575 -1640 18615 -1625
rect 17775 -4170 17825 -4155
rect 17775 -4190 17790 -4170
rect 17810 -4190 17825 -4170
rect 17775 -4220 17825 -4190
rect 17775 -4240 17790 -4220
rect 17810 -4240 17825 -4220
rect 17775 -4270 17825 -4240
rect 17775 -4290 17790 -4270
rect 17810 -4290 17825 -4270
rect 17775 -4305 17825 -4290
<< nsubdiff >>
rect 16335 1417 16375 1430
rect 16335 1395 16345 1417
rect 16365 1395 16375 1417
rect 16335 1365 16375 1395
rect 16335 1345 16345 1365
rect 16365 1345 16375 1365
rect 16335 1330 16375 1345
rect 16635 1417 16675 1430
rect 16635 1395 16645 1417
rect 16665 1395 16675 1417
rect 16635 1365 16675 1395
rect 16635 1345 16645 1365
rect 16665 1345 16675 1365
rect 16635 1330 16675 1345
rect 16845 1417 16885 1430
rect 16845 1345 16855 1417
rect 16875 1345 16885 1417
rect 16845 1330 16885 1345
rect 17255 1417 17295 1430
rect 17255 1345 17265 1417
rect 17285 1345 17295 1417
rect 17255 1330 17295 1345
rect 17465 1417 17505 1430
rect 17465 1395 17475 1417
rect 17495 1395 17505 1417
rect 17465 1365 17505 1395
rect 17465 1345 17475 1365
rect 17495 1345 17505 1365
rect 17465 1330 17505 1345
rect 18095 1417 18135 1430
rect 18095 1395 18105 1417
rect 18125 1395 18135 1417
rect 18095 1365 18135 1395
rect 18095 1345 18105 1365
rect 18125 1345 18135 1365
rect 18095 1330 18135 1345
rect 18305 1417 18345 1430
rect 18305 1345 18315 1417
rect 18335 1345 18345 1417
rect 18305 1330 18345 1345
rect 18715 1417 18755 1430
rect 18715 1345 18725 1417
rect 18745 1345 18755 1417
rect 18715 1330 18755 1345
rect 16930 950 16970 965
rect 16930 930 16940 950
rect 16960 930 16970 950
rect 16930 900 16970 930
rect 16930 880 16940 900
rect 16960 880 16970 900
rect 16395 850 16435 865
rect 16395 830 16405 850
rect 16425 830 16435 850
rect 16395 800 16435 830
rect 16395 780 16405 800
rect 16425 780 16435 800
rect 16395 765 16435 780
rect 16700 850 16740 865
rect 16700 830 16710 850
rect 16730 830 16740 850
rect 16700 800 16740 830
rect 16700 780 16710 800
rect 16730 780 16740 800
rect 16700 765 16740 780
rect 16930 850 16970 880
rect 16930 830 16940 850
rect 16960 830 16970 850
rect 16930 800 16970 830
rect 16930 780 16940 800
rect 16960 780 16970 800
rect 16930 750 16970 780
rect 16930 730 16940 750
rect 16960 730 16970 750
rect 16930 700 16970 730
rect 16930 680 16940 700
rect 16960 680 16970 700
rect 16930 665 16970 680
rect 18630 950 18670 965
rect 18630 930 18640 950
rect 18660 930 18670 950
rect 18630 900 18670 930
rect 18630 880 18640 900
rect 18660 880 18670 900
rect 18630 850 18670 880
rect 18630 830 18640 850
rect 18660 830 18670 850
rect 18630 800 18670 830
rect 18630 780 18640 800
rect 18660 780 18670 800
rect 18630 750 18670 780
rect 18865 950 18905 965
rect 18865 930 18875 950
rect 18895 930 18905 950
rect 18865 900 18905 930
rect 18865 880 18875 900
rect 18895 880 18905 900
rect 18865 850 18905 880
rect 18865 830 18875 850
rect 18895 830 18905 850
rect 18865 800 18905 830
rect 18865 780 18875 800
rect 18895 780 18905 800
rect 18865 765 18905 780
rect 19110 950 19150 965
rect 19110 930 19120 950
rect 19140 930 19150 950
rect 19110 900 19150 930
rect 19110 880 19120 900
rect 19140 880 19150 900
rect 19110 850 19150 880
rect 19110 830 19120 850
rect 19140 830 19150 850
rect 19110 800 19150 830
rect 19110 780 19120 800
rect 19140 780 19150 800
rect 19110 765 19150 780
rect 18630 730 18640 750
rect 18660 730 18670 750
rect 18630 700 18670 730
rect 18630 680 18640 700
rect 18660 680 18670 700
rect 18630 665 18670 680
rect 16380 110 16420 125
rect 16380 90 16390 110
rect 16410 90 16420 110
rect 16380 60 16420 90
rect 16380 40 16390 60
rect 16410 40 16420 60
rect 16380 25 16420 40
rect 17660 110 17700 125
rect 17660 90 17670 110
rect 17690 90 17700 110
rect 17660 60 17700 90
rect 17660 40 17670 60
rect 17690 40 17700 60
rect 17660 25 17700 40
rect 17900 110 17940 125
rect 17900 90 17910 110
rect 17930 90 17940 110
rect 17900 60 17940 90
rect 17900 40 17910 60
rect 17930 40 17940 60
rect 17900 25 17940 40
rect 19180 110 19220 125
rect 19180 90 19190 110
rect 19210 90 19220 110
rect 19180 60 19220 90
rect 19180 40 19190 60
rect 19210 40 19220 60
rect 19180 25 19220 40
<< psubdiffcont >>
rect 17570 -195 17590 -175
rect 17570 -235 17590 -215
rect 17570 -275 17590 -255
rect 18010 -195 18030 -175
rect 18010 -235 18030 -215
rect 18010 -275 18030 -255
rect 17120 -730 17140 -710
rect 17120 -780 17140 -760
rect 17120 -830 17140 -810
rect 17120 -880 17140 -860
rect 17120 -930 17140 -910
rect 18460 -730 18480 -710
rect 18460 -780 18480 -760
rect 18460 -830 18480 -810
rect 18460 -880 18480 -860
rect 18460 -930 18480 -910
rect 18870 -1185 18890 -1165
rect 18870 -1235 18890 -1215
rect 16570 -1575 16590 -1555
rect 16570 -1625 16590 -1605
rect 16925 -1575 16945 -1555
rect 16925 -1625 16945 -1605
rect 16995 -1575 17015 -1555
rect 16995 -1625 17015 -1605
rect 17515 -1575 17535 -1555
rect 17515 -1625 17535 -1605
rect 17585 -1575 17605 -1555
rect 17585 -1625 17605 -1605
rect 17995 -1575 18015 -1555
rect 17995 -1625 18015 -1605
rect 18065 -1575 18085 -1555
rect 18065 -1625 18085 -1605
rect 18585 -1575 18605 -1555
rect 18585 -1625 18605 -1605
rect 17790 -4190 17810 -4170
rect 17790 -4240 17810 -4220
rect 17790 -4290 17810 -4270
<< nsubdiffcont >>
rect 16345 1395 16365 1417
rect 16345 1345 16365 1365
rect 16645 1395 16665 1417
rect 16645 1345 16665 1365
rect 16855 1345 16875 1417
rect 17265 1345 17285 1417
rect 17475 1395 17495 1417
rect 17475 1345 17495 1365
rect 18105 1395 18125 1417
rect 18105 1345 18125 1365
rect 18315 1345 18335 1417
rect 18725 1345 18745 1417
rect 16940 930 16960 950
rect 16940 880 16960 900
rect 16405 830 16425 850
rect 16405 780 16425 800
rect 16710 830 16730 850
rect 16710 780 16730 800
rect 16940 830 16960 850
rect 16940 780 16960 800
rect 16940 730 16960 750
rect 16940 680 16960 700
rect 18640 930 18660 950
rect 18640 880 18660 900
rect 18640 830 18660 850
rect 18640 780 18660 800
rect 18875 930 18895 950
rect 18875 880 18895 900
rect 18875 830 18895 850
rect 18875 780 18895 800
rect 19120 930 19140 950
rect 19120 880 19140 900
rect 19120 830 19140 850
rect 19120 780 19140 800
rect 18640 730 18660 750
rect 18640 680 18660 700
rect 16390 90 16410 110
rect 16390 40 16410 60
rect 17670 90 17690 110
rect 17670 40 17690 60
rect 17910 90 17930 110
rect 17910 40 17930 60
rect 19190 90 19210 110
rect 19190 40 19210 60
<< poly >>
rect 16485 1610 16525 1620
rect 16485 1590 16495 1610
rect 16515 1590 16525 1610
rect 16485 1580 16525 1590
rect 17780 1610 17820 1620
rect 17780 1590 17790 1610
rect 17810 1590 17820 1610
rect 17780 1580 17820 1590
rect 16365 1475 16405 1485
rect 16365 1455 16375 1475
rect 16395 1460 16405 1475
rect 16395 1455 16430 1460
rect 16495 1455 16515 1580
rect 16605 1475 16645 1485
rect 16605 1460 16615 1475
rect 16580 1455 16615 1460
rect 16635 1455 16645 1475
rect 16365 1445 16430 1455
rect 16415 1430 16430 1445
rect 16470 1440 16540 1455
rect 16470 1430 16485 1440
rect 16525 1430 16540 1440
rect 16580 1445 16645 1455
rect 16885 1475 16925 1485
rect 16885 1455 16895 1475
rect 16915 1455 16925 1475
rect 17055 1475 17085 1485
rect 17055 1455 17060 1475
rect 17080 1455 17085 1475
rect 17215 1475 17255 1485
rect 17215 1455 17225 1475
rect 17245 1455 17255 1475
rect 16580 1430 16595 1445
rect 16885 1440 16940 1455
rect 16925 1430 16940 1440
rect 16980 1440 17160 1455
rect 16980 1430 16995 1440
rect 17035 1430 17050 1440
rect 17090 1430 17105 1440
rect 17145 1430 17160 1440
rect 17200 1440 17255 1455
rect 17495 1475 17535 1485
rect 17495 1455 17505 1475
rect 17525 1460 17535 1475
rect 17525 1455 17560 1460
rect 17790 1455 17810 1580
rect 18065 1475 18105 1485
rect 18065 1460 18075 1475
rect 18040 1455 18075 1460
rect 18095 1455 18105 1475
rect 17495 1445 17560 1455
rect 17200 1430 17215 1440
rect 17545 1430 17560 1445
rect 17600 1440 18000 1455
rect 17600 1430 17615 1440
rect 17655 1430 17670 1440
rect 17710 1430 17725 1440
rect 17765 1430 17780 1440
rect 17820 1430 17835 1440
rect 17875 1430 17890 1440
rect 17930 1430 17945 1440
rect 17985 1430 18000 1440
rect 18040 1445 18105 1455
rect 18345 1475 18385 1485
rect 18345 1455 18355 1475
rect 18375 1460 18385 1475
rect 18515 1475 18545 1485
rect 18375 1455 18400 1460
rect 18515 1455 18520 1475
rect 18540 1455 18545 1475
rect 18675 1475 18715 1485
rect 18675 1460 18685 1475
rect 18660 1455 18685 1460
rect 18705 1455 18715 1475
rect 18345 1445 18400 1455
rect 18040 1430 18055 1445
rect 18385 1430 18400 1445
rect 18440 1440 18620 1455
rect 18440 1430 18455 1440
rect 18495 1430 18510 1440
rect 18550 1430 18565 1440
rect 18605 1430 18620 1440
rect 18660 1445 18715 1455
rect 18660 1430 18675 1445
rect 16415 1315 16430 1330
rect 16470 1315 16485 1330
rect 16525 1315 16540 1330
rect 16580 1315 16595 1330
rect 16925 1315 16940 1330
rect 16980 1315 16995 1330
rect 17035 1315 17050 1330
rect 17090 1315 17105 1330
rect 17145 1315 17160 1330
rect 17200 1315 17215 1330
rect 17545 1315 17560 1330
rect 17600 1315 17615 1330
rect 17655 1315 17670 1330
rect 17710 1315 17725 1330
rect 17765 1315 17780 1330
rect 17820 1315 17835 1330
rect 17875 1315 17890 1330
rect 17930 1315 17945 1330
rect 17985 1315 18000 1330
rect 18040 1315 18055 1330
rect 18385 1315 18400 1330
rect 18440 1315 18455 1330
rect 18495 1315 18510 1330
rect 18550 1315 18565 1330
rect 18605 1315 18620 1330
rect 18660 1315 18675 1330
rect 16970 1010 17010 1020
rect 16970 990 16980 1010
rect 17000 995 17010 1010
rect 18590 1010 18630 1020
rect 18590 995 18600 1010
rect 17000 990 17060 995
rect 16970 980 17060 990
rect 18540 990 18600 995
rect 18620 990 18630 1010
rect 18540 980 18630 990
rect 18910 1010 18940 1020
rect 18910 990 18915 1010
rect 18935 995 18940 1010
rect 19080 1010 19110 1020
rect 19080 995 19085 1010
rect 18935 990 18960 995
rect 18910 980 18960 990
rect 19055 990 19085 995
rect 19105 990 19110 1010
rect 19055 980 19110 990
rect 17010 965 17060 980
rect 17100 965 17150 980
rect 17190 965 17240 980
rect 17280 965 17330 980
rect 17370 965 17420 980
rect 17460 965 17510 980
rect 17550 965 17600 980
rect 17640 965 17690 980
rect 17730 965 17780 980
rect 17820 965 17870 980
rect 17910 965 17960 980
rect 18000 965 18050 980
rect 18090 965 18140 980
rect 18180 965 18230 980
rect 18270 965 18320 980
rect 18360 965 18410 980
rect 18450 965 18500 980
rect 18540 965 18590 980
rect 18945 965 18960 980
rect 19000 965 19015 980
rect 19055 965 19070 980
rect 16440 910 16470 920
rect 16440 890 16445 910
rect 16465 890 16470 910
rect 16660 910 16690 920
rect 16660 890 16665 910
rect 16685 890 16690 910
rect 16440 875 16490 890
rect 16475 865 16490 875
rect 16530 865 16545 880
rect 16585 865 16600 880
rect 16640 875 16690 890
rect 16640 865 16655 875
rect 16475 750 16490 765
rect 16530 755 16545 765
rect 16585 755 16600 765
rect 16530 740 16600 755
rect 16640 750 16655 765
rect 16545 720 16555 740
rect 16575 720 16585 740
rect 16545 710 16585 720
rect 18945 750 18960 765
rect 19000 690 19015 765
rect 19055 750 19070 765
rect 19000 680 19040 690
rect 17010 650 17060 665
rect 17100 655 17150 665
rect 17190 655 17240 665
rect 17280 655 17330 665
rect 17370 655 17420 665
rect 17460 655 17510 665
rect 17550 655 17600 665
rect 17640 655 17690 665
rect 17730 655 17780 665
rect 17820 655 17870 665
rect 17910 655 17960 665
rect 18000 655 18050 665
rect 18090 655 18140 665
rect 18180 655 18230 665
rect 18270 655 18320 665
rect 18360 655 18410 665
rect 18450 655 18500 665
rect 17100 640 18500 655
rect 18540 650 18590 665
rect 19000 660 19010 680
rect 19030 660 19040 680
rect 19000 650 19040 660
rect 17690 620 17700 640
rect 17720 620 17730 640
rect 17690 610 17730 620
rect 16425 170 16455 180
rect 16425 150 16430 170
rect 16450 150 16455 170
rect 17625 170 17655 180
rect 17625 150 17630 170
rect 17650 150 17655 170
rect 16425 135 16480 150
rect 16460 125 16480 135
rect 16520 125 16540 140
rect 16580 125 16600 140
rect 16640 125 16660 140
rect 16700 125 16720 140
rect 16760 125 16780 140
rect 16820 125 16840 140
rect 16880 125 16900 140
rect 16940 125 16960 140
rect 17000 125 17020 140
rect 17060 125 17080 140
rect 17120 125 17140 140
rect 17180 125 17200 140
rect 17240 125 17260 140
rect 17300 125 17320 140
rect 17360 125 17380 140
rect 17420 125 17440 140
rect 17480 125 17500 140
rect 17540 125 17560 140
rect 17600 135 17655 150
rect 17945 170 17975 180
rect 17945 150 17950 170
rect 17970 150 17975 170
rect 19145 170 19175 180
rect 19145 150 19150 170
rect 19170 150 19175 170
rect 17945 135 18000 150
rect 17600 125 17620 135
rect 17980 125 18000 135
rect 18040 125 18060 140
rect 18100 125 18120 140
rect 18160 125 18180 140
rect 18220 125 18240 140
rect 18280 125 18300 140
rect 18340 125 18360 140
rect 18400 125 18420 140
rect 18460 125 18480 140
rect 18520 125 18540 140
rect 18580 125 18600 140
rect 18640 125 18660 140
rect 18700 125 18720 140
rect 18760 125 18780 140
rect 18820 125 18840 140
rect 18880 125 18900 140
rect 18940 125 18960 140
rect 19000 125 19020 140
rect 19060 125 19080 140
rect 19120 135 19175 150
rect 19120 125 19140 135
rect 16460 15 16480 25
rect 16425 0 16480 15
rect 16520 10 16540 25
rect 16580 15 16600 25
rect 16640 15 16660 25
rect 16700 15 16720 25
rect 16760 15 16780 25
rect 16510 0 16550 10
rect 16580 0 16780 15
rect 16820 15 16840 25
rect 16880 15 16900 25
rect 16820 0 16900 15
rect 16940 15 16960 25
rect 17000 15 17020 25
rect 17060 15 17080 25
rect 17120 15 17140 25
rect 16940 0 17140 15
rect 17180 15 17200 25
rect 17240 15 17260 25
rect 17180 0 17260 15
rect 17300 15 17320 25
rect 17360 15 17380 25
rect 17420 15 17440 25
rect 17480 15 17500 25
rect 17300 0 17500 15
rect 17540 10 17560 25
rect 17600 10 17620 25
rect 17980 15 18000 25
rect 17535 0 17565 10
rect 16425 -20 16430 0
rect 16450 -20 16455 0
rect 16425 -30 16455 -20
rect 16510 -20 16520 0
rect 16540 -20 16550 0
rect 16510 -30 16550 -20
rect 16600 -20 16610 0
rect 16630 -20 16640 0
rect 16600 -30 16640 -20
rect 16840 -20 16850 0
rect 16870 -20 16880 0
rect 16840 -30 16880 -20
rect 16960 -20 16970 0
rect 16990 -20 17000 0
rect 16960 -30 17000 -20
rect 17200 -20 17210 0
rect 17230 -20 17240 0
rect 17200 -30 17240 -20
rect 17320 -20 17330 0
rect 17350 -20 17360 0
rect 17320 -30 17360 -20
rect 17535 -20 17540 0
rect 17560 -20 17565 0
rect 17535 -30 17565 -20
rect 17945 0 18000 15
rect 18040 10 18060 25
rect 18100 15 18120 25
rect 18160 15 18180 25
rect 18220 15 18240 25
rect 18280 15 18300 25
rect 18035 0 18065 10
rect 18100 0 18300 15
rect 18340 15 18360 25
rect 18400 15 18420 25
rect 18340 0 18420 15
rect 18460 15 18480 25
rect 18520 15 18540 25
rect 18580 15 18600 25
rect 18640 15 18660 25
rect 18460 0 18660 15
rect 18700 15 18720 25
rect 18760 15 18780 25
rect 18700 0 18780 15
rect 18820 15 18840 25
rect 18880 15 18900 25
rect 18940 15 18960 25
rect 19000 15 19020 25
rect 18820 0 19020 15
rect 19060 10 19080 25
rect 19120 15 19140 25
rect 19050 0 19090 10
rect 19120 0 19175 15
rect 17945 -20 17950 0
rect 17970 -20 17975 0
rect 17945 -30 17975 -20
rect 18035 -20 18040 0
rect 18060 -20 18065 0
rect 18035 -30 18065 -20
rect 18240 -20 18250 0
rect 18270 -20 18280 0
rect 18240 -30 18280 -20
rect 18360 -20 18370 0
rect 18390 -20 18400 0
rect 18360 -30 18400 -20
rect 18600 -20 18610 0
rect 18630 -20 18640 0
rect 18600 -30 18640 -20
rect 18720 -20 18730 0
rect 18750 -20 18760 0
rect 18720 -30 18760 -20
rect 18960 -20 18970 0
rect 18990 -20 19000 0
rect 18960 -30 19000 -20
rect 19050 -20 19060 0
rect 19080 -20 19090 0
rect 19050 -30 19090 -20
rect 19145 -20 19150 0
rect 19170 -20 19175 0
rect 19145 -30 19175 -20
rect 17007 -115 17037 -105
rect 17007 -130 17012 -115
rect 17000 -135 17012 -130
rect 17032 -135 17037 -115
rect 17000 -145 17037 -135
rect 18563 -115 18593 -105
rect 18563 -135 18568 -115
rect 18588 -130 18593 -115
rect 18588 -135 18600 -130
rect 18563 -145 18600 -135
rect 17000 -160 17020 -145
rect 17060 -160 17080 -145
rect 18520 -160 18540 -145
rect 18580 -160 18600 -145
rect 17000 -425 17020 -410
rect 17060 -425 17080 -410
rect 18520 -425 18540 -410
rect 18580 -425 18600 -410
rect 17060 -435 17105 -425
rect 17060 -455 17080 -435
rect 17100 -455 17105 -435
rect 17060 -465 17105 -455
rect 18495 -435 18540 -425
rect 18495 -455 18500 -435
rect 18520 -455 18540 -435
rect 18495 -465 18540 -455
rect 16620 -650 16660 -640
rect 16620 -670 16630 -650
rect 16650 -670 16660 -650
rect 16620 -680 16660 -670
rect 16740 -650 16780 -640
rect 16740 -670 16750 -650
rect 16770 -670 16780 -650
rect 16740 -680 16780 -670
rect 16860 -650 16900 -640
rect 16860 -670 16870 -650
rect 16890 -670 16900 -650
rect 16860 -680 16900 -670
rect 16980 -650 17020 -640
rect 16980 -670 16990 -650
rect 17010 -670 17020 -650
rect 16980 -680 17020 -670
rect 17300 -650 17340 -640
rect 17300 -670 17310 -650
rect 17330 -670 17340 -650
rect 17300 -680 17340 -670
rect 17420 -650 17460 -640
rect 17420 -670 17430 -650
rect 17450 -670 17460 -650
rect 17420 -680 17460 -670
rect 17540 -650 17580 -640
rect 17540 -670 17550 -650
rect 17570 -670 17580 -650
rect 17540 -680 17580 -670
rect 18020 -650 18060 -640
rect 18020 -670 18030 -650
rect 18050 -670 18060 -650
rect 18020 -680 18060 -670
rect 18140 -650 18180 -640
rect 18140 -670 18150 -650
rect 18170 -670 18180 -650
rect 18140 -680 18180 -670
rect 18260 -650 18300 -640
rect 18260 -670 18270 -650
rect 18290 -670 18300 -650
rect 18260 -680 18300 -670
rect 18580 -650 18620 -640
rect 18580 -670 18590 -650
rect 18610 -670 18620 -650
rect 18580 -680 18620 -670
rect 18700 -650 18740 -640
rect 18700 -670 18710 -650
rect 18730 -670 18740 -650
rect 18700 -680 18740 -670
rect 18820 -650 18860 -640
rect 18820 -670 18830 -650
rect 18850 -670 18860 -650
rect 18820 -680 18860 -670
rect 18940 -650 18980 -640
rect 18940 -670 18950 -650
rect 18970 -670 18980 -650
rect 18940 -680 18980 -670
rect 16570 -695 17070 -680
rect 17190 -695 17690 -680
rect 17910 -695 18410 -680
rect 18530 -695 19030 -680
rect 16570 -960 17070 -945
rect 17190 -960 17690 -945
rect 17910 -960 18410 -945
rect 18530 -960 19030 -945
rect 16820 -1105 16860 -1095
rect 16820 -1125 16830 -1105
rect 16850 -1125 16860 -1105
rect 16820 -1135 16860 -1125
rect 16900 -1105 16940 -1095
rect 16900 -1125 16910 -1105
rect 16930 -1125 16940 -1105
rect 16900 -1135 16940 -1125
rect 16980 -1105 17020 -1095
rect 16980 -1125 16990 -1105
rect 17010 -1125 17020 -1105
rect 16980 -1135 17020 -1125
rect 17060 -1105 17100 -1095
rect 17060 -1125 17070 -1105
rect 17090 -1125 17100 -1105
rect 17060 -1135 17100 -1125
rect 17140 -1105 17180 -1095
rect 17140 -1125 17150 -1105
rect 17170 -1125 17180 -1105
rect 17140 -1135 17180 -1125
rect 17220 -1105 17260 -1095
rect 17220 -1125 17230 -1105
rect 17250 -1125 17260 -1105
rect 17220 -1135 17260 -1125
rect 17300 -1105 17340 -1095
rect 17300 -1125 17310 -1105
rect 17330 -1125 17340 -1105
rect 17300 -1135 17340 -1125
rect 17380 -1105 17420 -1095
rect 17380 -1125 17390 -1105
rect 17410 -1125 17420 -1105
rect 17380 -1135 17420 -1125
rect 17460 -1105 17500 -1095
rect 17460 -1125 17470 -1105
rect 17490 -1125 17500 -1105
rect 17460 -1135 17500 -1125
rect 17540 -1105 17580 -1095
rect 17540 -1125 17550 -1105
rect 17570 -1125 17580 -1105
rect 17540 -1135 17580 -1125
rect 17620 -1105 17660 -1095
rect 17620 -1125 17630 -1105
rect 17650 -1125 17660 -1105
rect 17620 -1135 17660 -1125
rect 17700 -1105 17740 -1095
rect 17700 -1125 17710 -1105
rect 17730 -1125 17740 -1105
rect 17700 -1135 17740 -1125
rect 17860 -1105 17900 -1095
rect 17860 -1125 17870 -1105
rect 17890 -1125 17900 -1105
rect 17860 -1135 17900 -1125
rect 17940 -1105 17980 -1095
rect 17940 -1125 17950 -1105
rect 17970 -1125 17980 -1105
rect 17940 -1135 17980 -1125
rect 18020 -1105 18060 -1095
rect 18020 -1125 18030 -1105
rect 18050 -1125 18060 -1105
rect 18020 -1135 18060 -1125
rect 18100 -1105 18140 -1095
rect 18100 -1125 18110 -1105
rect 18130 -1125 18140 -1105
rect 18100 -1135 18140 -1125
rect 18180 -1105 18220 -1095
rect 18180 -1125 18190 -1105
rect 18210 -1125 18220 -1105
rect 18180 -1135 18220 -1125
rect 18260 -1105 18300 -1095
rect 18260 -1125 18270 -1105
rect 18290 -1125 18300 -1105
rect 18260 -1135 18300 -1125
rect 18340 -1105 18380 -1095
rect 18340 -1125 18350 -1105
rect 18370 -1125 18380 -1105
rect 18340 -1135 18380 -1125
rect 18420 -1105 18460 -1095
rect 18420 -1125 18430 -1105
rect 18450 -1125 18460 -1105
rect 18420 -1135 18460 -1125
rect 18500 -1105 18540 -1095
rect 18500 -1125 18510 -1105
rect 18530 -1125 18540 -1105
rect 18500 -1135 18540 -1125
rect 18580 -1105 18620 -1095
rect 18580 -1125 18590 -1105
rect 18610 -1125 18620 -1105
rect 18580 -1135 18620 -1125
rect 18660 -1105 18700 -1095
rect 18660 -1125 18670 -1105
rect 18690 -1125 18700 -1105
rect 18660 -1135 18700 -1125
rect 18740 -1105 18780 -1095
rect 18740 -1125 18750 -1105
rect 18770 -1125 18780 -1105
rect 18740 -1135 18780 -1125
rect 16780 -1150 17780 -1135
rect 17820 -1150 18820 -1135
rect 16780 -1265 17780 -1250
rect 17820 -1265 18820 -1250
rect 16600 -1495 16640 -1485
rect 16600 -1515 16610 -1495
rect 16630 -1510 16640 -1495
rect 16770 -1495 16800 -1485
rect 16630 -1515 16655 -1510
rect 16770 -1515 16775 -1495
rect 16795 -1515 16800 -1495
rect 16880 -1495 16920 -1485
rect 16880 -1510 16890 -1495
rect 16860 -1515 16890 -1510
rect 16910 -1515 16920 -1495
rect 16600 -1525 16655 -1515
rect 16640 -1540 16655 -1525
rect 16695 -1530 16820 -1515
rect 16695 -1540 16710 -1530
rect 16750 -1540 16765 -1530
rect 16805 -1540 16820 -1530
rect 16860 -1525 16920 -1515
rect 17025 -1495 17065 -1485
rect 17025 -1515 17035 -1495
rect 17055 -1510 17065 -1495
rect 17305 -1495 17335 -1485
rect 17055 -1515 17080 -1510
rect 17305 -1515 17310 -1495
rect 17330 -1515 17335 -1495
rect 17465 -1495 17505 -1485
rect 17465 -1510 17475 -1495
rect 17450 -1515 17475 -1510
rect 17495 -1515 17505 -1495
rect 17025 -1525 17080 -1515
rect 16860 -1540 16875 -1525
rect 17065 -1540 17080 -1525
rect 17120 -1530 17410 -1515
rect 17120 -1540 17135 -1530
rect 17175 -1540 17190 -1530
rect 17230 -1540 17245 -1530
rect 17285 -1540 17300 -1530
rect 17340 -1540 17355 -1530
rect 17395 -1540 17410 -1530
rect 17450 -1525 17505 -1515
rect 17615 -1495 17655 -1485
rect 17615 -1515 17625 -1495
rect 17645 -1510 17655 -1495
rect 17785 -1495 17815 -1485
rect 17645 -1515 17670 -1510
rect 17785 -1515 17790 -1495
rect 17810 -1515 17815 -1495
rect 17945 -1495 17985 -1485
rect 17945 -1510 17955 -1495
rect 17930 -1515 17955 -1510
rect 17975 -1515 17985 -1495
rect 17615 -1525 17670 -1515
rect 17450 -1540 17465 -1525
rect 17655 -1540 17670 -1525
rect 17710 -1530 17890 -1515
rect 17710 -1540 17725 -1530
rect 17765 -1540 17780 -1530
rect 17820 -1540 17835 -1530
rect 17875 -1540 17890 -1530
rect 17930 -1525 17985 -1515
rect 18095 -1495 18135 -1485
rect 18095 -1515 18105 -1495
rect 18125 -1510 18135 -1495
rect 18265 -1495 18295 -1485
rect 18125 -1515 18150 -1510
rect 18265 -1515 18270 -1495
rect 18290 -1515 18295 -1495
rect 18535 -1495 18575 -1485
rect 18535 -1510 18545 -1495
rect 18520 -1515 18545 -1510
rect 18565 -1515 18575 -1495
rect 18095 -1525 18150 -1515
rect 17930 -1540 17945 -1525
rect 18135 -1540 18150 -1525
rect 18190 -1530 18480 -1515
rect 18190 -1540 18205 -1530
rect 18245 -1540 18260 -1530
rect 18300 -1540 18315 -1530
rect 18355 -1540 18370 -1530
rect 18410 -1540 18425 -1530
rect 18465 -1540 18480 -1530
rect 18520 -1525 18575 -1515
rect 18520 -1540 18535 -1525
rect 16640 -1655 16655 -1640
rect 16695 -1655 16710 -1640
rect 16750 -1655 16765 -1640
rect 16805 -1655 16820 -1640
rect 16860 -1655 16875 -1640
rect 17065 -1655 17080 -1640
rect 17120 -1655 17135 -1640
rect 17175 -1655 17190 -1640
rect 17230 -1655 17245 -1640
rect 17285 -1655 17300 -1640
rect 17340 -1655 17355 -1640
rect 17395 -1655 17410 -1640
rect 17450 -1655 17465 -1640
rect 17655 -1655 17670 -1640
rect 17710 -1655 17725 -1640
rect 17765 -1655 17780 -1640
rect 17820 -1655 17835 -1640
rect 17875 -1655 17890 -1640
rect 17930 -1655 17945 -1640
rect 18135 -1655 18150 -1640
rect 18190 -1655 18205 -1640
rect 18245 -1655 18260 -1640
rect 18300 -1655 18315 -1640
rect 18355 -1655 18370 -1640
rect 18410 -1655 18425 -1640
rect 18465 -1655 18480 -1640
rect 18520 -1655 18535 -1640
<< polycont >>
rect 16495 1590 16515 1610
rect 17790 1590 17810 1610
rect 16375 1455 16395 1475
rect 16615 1455 16635 1475
rect 16895 1455 16915 1475
rect 17060 1455 17080 1475
rect 17225 1455 17245 1475
rect 17505 1455 17525 1475
rect 18075 1455 18095 1475
rect 18355 1455 18375 1475
rect 18520 1455 18540 1475
rect 18685 1455 18705 1475
rect 16980 990 17000 1010
rect 18600 990 18620 1010
rect 18915 990 18935 1010
rect 19085 990 19105 1010
rect 16445 890 16465 910
rect 16665 890 16685 910
rect 16555 720 16575 740
rect 19010 660 19030 680
rect 17700 620 17720 640
rect 16430 150 16450 170
rect 17630 150 17650 170
rect 17950 150 17970 170
rect 19150 150 19170 170
rect 16430 -20 16450 0
rect 16520 -20 16540 0
rect 16610 -20 16630 0
rect 16850 -20 16870 0
rect 16970 -20 16990 0
rect 17210 -20 17230 0
rect 17330 -20 17350 0
rect 17540 -20 17560 0
rect 17950 -20 17970 0
rect 18040 -20 18060 0
rect 18250 -20 18270 0
rect 18370 -20 18390 0
rect 18610 -20 18630 0
rect 18730 -20 18750 0
rect 18970 -20 18990 0
rect 19060 -20 19080 0
rect 19150 -20 19170 0
rect 17012 -135 17032 -115
rect 18568 -135 18588 -115
rect 17080 -455 17100 -435
rect 18500 -455 18520 -435
rect 16630 -670 16650 -650
rect 16750 -670 16770 -650
rect 16870 -670 16890 -650
rect 16990 -670 17010 -650
rect 17310 -670 17330 -650
rect 17430 -670 17450 -650
rect 17550 -670 17570 -650
rect 18030 -670 18050 -650
rect 18150 -670 18170 -650
rect 18270 -670 18290 -650
rect 18590 -670 18610 -650
rect 18710 -670 18730 -650
rect 18830 -670 18850 -650
rect 18950 -670 18970 -650
rect 16830 -1125 16850 -1105
rect 16910 -1125 16930 -1105
rect 16990 -1125 17010 -1105
rect 17070 -1125 17090 -1105
rect 17150 -1125 17170 -1105
rect 17230 -1125 17250 -1105
rect 17310 -1125 17330 -1105
rect 17390 -1125 17410 -1105
rect 17470 -1125 17490 -1105
rect 17550 -1125 17570 -1105
rect 17630 -1125 17650 -1105
rect 17710 -1125 17730 -1105
rect 17870 -1125 17890 -1105
rect 17950 -1125 17970 -1105
rect 18030 -1125 18050 -1105
rect 18110 -1125 18130 -1105
rect 18190 -1125 18210 -1105
rect 18270 -1125 18290 -1105
rect 18350 -1125 18370 -1105
rect 18430 -1125 18450 -1105
rect 18510 -1125 18530 -1105
rect 18590 -1125 18610 -1105
rect 18670 -1125 18690 -1105
rect 18750 -1125 18770 -1105
rect 16610 -1515 16630 -1495
rect 16775 -1515 16795 -1495
rect 16890 -1515 16910 -1495
rect 17035 -1515 17055 -1495
rect 17310 -1515 17330 -1495
rect 17475 -1515 17495 -1495
rect 17625 -1515 17645 -1495
rect 17790 -1515 17810 -1495
rect 17955 -1515 17975 -1495
rect 18105 -1515 18125 -1495
rect 18270 -1515 18290 -1495
rect 18545 -1515 18565 -1495
<< xpolycontact >>
rect 17470 -2035 17690 -2000
rect 17904 -2035 18124 -2000
rect 15950 -3376 15985 -3156
rect 15950 -3784 15985 -3565
rect 16160 -3285 16195 -3065
rect 16160 -3889 16195 -3669
rect 16220 -3285 16255 -3065
rect 16220 -3889 16255 -3669
rect 16280 -3285 16315 -3065
rect 16280 -3889 16315 -3669
rect 16485 -3160 16520 -2940
rect 16485 -3964 16520 -3744
rect 16545 -3160 16580 -2940
rect 16545 -3964 16580 -3744
rect 16605 -3160 16640 -2940
rect 16605 -3964 16640 -3744
rect 18960 -3160 18995 -2940
rect 18960 -3964 18995 -3744
rect 19020 -3160 19055 -2940
rect 19020 -3964 19055 -3744
rect 19080 -3160 19115 -2940
rect 19080 -3964 19115 -3744
rect 19285 -3257 19320 -3037
rect 19285 -3889 19320 -3669
rect 19345 -3257 19380 -3037
rect 19345 -3889 19380 -3669
rect 19405 -3257 19440 -3037
rect 19405 -3889 19440 -3669
rect 19610 -3376 19645 -3156
rect 19610 -3784 19645 -3565
<< ppolyres >>
rect 15950 -3565 15985 -3376
rect 19610 -3565 19645 -3376
<< xpolyres >>
rect 17690 -2035 17904 -2000
rect 16160 -3669 16195 -3285
rect 16220 -3669 16255 -3285
rect 16280 -3669 16315 -3285
rect 16485 -3744 16520 -3160
rect 16545 -3744 16580 -3160
rect 16605 -3744 16640 -3160
rect 18960 -3744 18995 -3160
rect 19020 -3744 19055 -3160
rect 19080 -3744 19115 -3160
rect 19285 -3669 19320 -3257
rect 19345 -3669 19380 -3257
rect 19405 -3669 19440 -3257
<< locali >>
rect 16485 1610 16525 1620
rect 16485 1590 16495 1610
rect 16515 1590 16525 1610
rect 16485 1580 16525 1590
rect 17780 1610 17820 1620
rect 17780 1590 17790 1610
rect 17810 1590 17820 1610
rect 17780 1580 17820 1590
rect 16365 1475 16405 1485
rect 16365 1455 16375 1475
rect 16395 1455 16405 1475
rect 16365 1445 16405 1455
rect 16485 1475 16525 1485
rect 16485 1455 16495 1475
rect 16515 1455 16525 1475
rect 16485 1445 16525 1455
rect 16605 1475 16645 1485
rect 16605 1455 16615 1475
rect 16635 1455 16645 1475
rect 16605 1445 16645 1455
rect 16885 1475 16925 1485
rect 16885 1455 16895 1475
rect 16915 1455 16925 1475
rect 16885 1445 16925 1455
rect 16945 1475 16975 1485
rect 16945 1455 16950 1475
rect 16970 1455 16975 1475
rect 16945 1445 16975 1455
rect 16995 1475 17035 1485
rect 16995 1455 17005 1475
rect 17025 1455 17035 1475
rect 16995 1445 17035 1455
rect 17055 1475 17085 1485
rect 17055 1455 17060 1475
rect 17080 1455 17085 1475
rect 17055 1445 17085 1455
rect 17105 1475 17145 1485
rect 17105 1455 17115 1475
rect 17135 1455 17145 1475
rect 17105 1445 17145 1455
rect 17215 1475 17255 1485
rect 17215 1455 17225 1475
rect 17245 1455 17255 1475
rect 17215 1445 17255 1455
rect 17495 1475 17535 1485
rect 17495 1455 17505 1475
rect 17525 1455 17535 1475
rect 17495 1445 17535 1455
rect 17560 1475 17600 1485
rect 17560 1455 17570 1475
rect 17590 1455 17600 1475
rect 17560 1445 17600 1455
rect 17620 1475 17650 1485
rect 17620 1455 17625 1475
rect 17645 1455 17650 1475
rect 16385 1425 16405 1445
rect 16495 1425 16515 1445
rect 16605 1425 16625 1445
rect 16895 1425 16915 1445
rect 16950 1425 16970 1445
rect 17005 1425 17025 1445
rect 17115 1425 17135 1445
rect 17225 1425 17245 1445
rect 17515 1425 17535 1445
rect 17570 1425 17590 1445
rect 16340 1417 16410 1425
rect 16340 1395 16345 1417
rect 16365 1415 16410 1417
rect 16365 1395 16385 1415
rect 16405 1395 16410 1415
rect 16340 1365 16410 1395
rect 16340 1345 16345 1365
rect 16365 1345 16385 1365
rect 16405 1345 16410 1365
rect 16340 1335 16410 1345
rect 16435 1415 16465 1425
rect 16435 1395 16440 1415
rect 16460 1395 16465 1415
rect 16435 1365 16465 1395
rect 16435 1345 16440 1365
rect 16460 1345 16465 1365
rect 16435 1335 16465 1345
rect 16490 1415 16520 1425
rect 16490 1395 16495 1415
rect 16515 1395 16520 1415
rect 16490 1365 16520 1395
rect 16490 1345 16495 1365
rect 16515 1345 16520 1365
rect 16490 1335 16520 1345
rect 16545 1415 16575 1425
rect 16545 1395 16550 1415
rect 16570 1395 16575 1415
rect 16545 1365 16575 1395
rect 16545 1345 16550 1365
rect 16570 1345 16575 1365
rect 16545 1335 16575 1345
rect 16600 1417 16670 1425
rect 16600 1415 16645 1417
rect 16600 1395 16605 1415
rect 16625 1395 16645 1415
rect 16665 1395 16670 1417
rect 16600 1365 16670 1395
rect 16600 1345 16605 1365
rect 16625 1345 16645 1365
rect 16665 1345 16670 1365
rect 16600 1335 16670 1345
rect 16850 1417 16920 1425
rect 16850 1345 16855 1417
rect 16875 1415 16920 1417
rect 16875 1345 16895 1415
rect 16850 1343 16895 1345
rect 16915 1343 16920 1415
rect 16850 1335 16920 1343
rect 16945 1415 16975 1425
rect 16945 1343 16950 1415
rect 16970 1343 16975 1415
rect 16945 1335 16975 1343
rect 17000 1415 17030 1425
rect 17000 1343 17005 1415
rect 17025 1343 17030 1415
rect 17000 1335 17030 1343
rect 17055 1415 17085 1425
rect 17055 1343 17060 1415
rect 17080 1343 17085 1415
rect 17055 1335 17085 1343
rect 17110 1415 17140 1425
rect 17110 1343 17115 1415
rect 17135 1343 17140 1415
rect 17110 1335 17140 1343
rect 17165 1415 17195 1425
rect 17165 1343 17170 1415
rect 17190 1343 17195 1415
rect 17165 1335 17195 1343
rect 17220 1417 17290 1425
rect 17220 1415 17265 1417
rect 17220 1343 17225 1415
rect 17245 1345 17265 1415
rect 17285 1345 17290 1417
rect 17245 1343 17290 1345
rect 17220 1335 17290 1343
rect 17470 1417 17540 1425
rect 17470 1395 17475 1417
rect 17495 1415 17540 1417
rect 17495 1395 17515 1415
rect 17535 1395 17540 1415
rect 17470 1365 17540 1395
rect 17470 1345 17475 1365
rect 17495 1345 17515 1365
rect 17535 1345 17540 1365
rect 17470 1335 17540 1345
rect 17565 1415 17595 1425
rect 17565 1395 17570 1415
rect 17590 1395 17595 1415
rect 17565 1365 17595 1395
rect 17565 1345 17570 1365
rect 17590 1345 17595 1365
rect 17565 1335 17595 1345
rect 17620 1415 17650 1455
rect 17670 1475 17710 1485
rect 17670 1455 17680 1475
rect 17700 1455 17710 1475
rect 17670 1445 17710 1455
rect 17730 1475 17760 1485
rect 17730 1455 17735 1475
rect 17755 1455 17760 1475
rect 17680 1425 17700 1445
rect 17620 1395 17625 1415
rect 17645 1395 17650 1415
rect 17620 1365 17650 1395
rect 17620 1345 17625 1365
rect 17645 1345 17650 1365
rect 17620 1335 17650 1345
rect 17675 1415 17705 1425
rect 17675 1395 17680 1415
rect 17700 1395 17705 1415
rect 17675 1365 17705 1395
rect 17675 1345 17680 1365
rect 17700 1345 17705 1365
rect 17675 1335 17705 1345
rect 17730 1415 17760 1455
rect 17780 1475 17820 1485
rect 17780 1455 17790 1475
rect 17810 1455 17820 1475
rect 17780 1445 17820 1455
rect 17840 1475 17870 1485
rect 17840 1455 17845 1475
rect 17865 1455 17870 1475
rect 17790 1425 17810 1445
rect 17730 1395 17735 1415
rect 17755 1395 17760 1415
rect 17730 1365 17760 1395
rect 17730 1345 17735 1365
rect 17755 1345 17760 1365
rect 17730 1335 17760 1345
rect 17785 1415 17815 1425
rect 17785 1395 17790 1415
rect 17810 1395 17815 1415
rect 17785 1365 17815 1395
rect 17785 1345 17790 1365
rect 17810 1345 17815 1365
rect 17785 1335 17815 1345
rect 17840 1415 17870 1455
rect 17890 1475 17930 1485
rect 17890 1455 17900 1475
rect 17920 1455 17930 1475
rect 17890 1445 17930 1455
rect 17950 1475 17980 1485
rect 17950 1455 17955 1475
rect 17975 1455 17980 1475
rect 17900 1425 17920 1445
rect 17840 1395 17845 1415
rect 17865 1395 17870 1415
rect 17840 1365 17870 1395
rect 17840 1345 17845 1365
rect 17865 1345 17870 1365
rect 17840 1335 17870 1345
rect 17895 1415 17925 1425
rect 17895 1395 17900 1415
rect 17920 1395 17925 1415
rect 17895 1365 17925 1395
rect 17895 1345 17900 1365
rect 17920 1345 17925 1365
rect 17895 1335 17925 1345
rect 17950 1415 17980 1455
rect 18000 1475 18040 1485
rect 18000 1455 18010 1475
rect 18030 1455 18040 1475
rect 18000 1445 18040 1455
rect 18065 1475 18105 1485
rect 18065 1455 18075 1475
rect 18095 1455 18105 1475
rect 18065 1445 18105 1455
rect 18345 1475 18385 1485
rect 18345 1455 18355 1475
rect 18375 1455 18385 1475
rect 18345 1445 18385 1455
rect 18455 1475 18495 1485
rect 18455 1455 18465 1475
rect 18485 1455 18495 1475
rect 18455 1445 18495 1455
rect 18515 1475 18545 1485
rect 18515 1455 18520 1475
rect 18540 1455 18545 1475
rect 18515 1445 18545 1455
rect 18565 1475 18605 1485
rect 18565 1455 18575 1475
rect 18595 1455 18605 1475
rect 18565 1445 18605 1455
rect 18625 1475 18655 1485
rect 18625 1455 18630 1475
rect 18650 1455 18655 1475
rect 18625 1445 18655 1455
rect 18675 1475 18715 1485
rect 18675 1455 18685 1475
rect 18705 1455 18715 1475
rect 18675 1445 18715 1455
rect 18010 1425 18030 1445
rect 18065 1425 18085 1445
rect 18355 1425 18375 1445
rect 18465 1425 18485 1445
rect 18575 1425 18595 1445
rect 18630 1425 18650 1445
rect 18685 1425 18705 1445
rect 17950 1395 17955 1415
rect 17975 1395 17980 1415
rect 17950 1365 17980 1395
rect 17950 1345 17955 1365
rect 17975 1345 17980 1365
rect 17950 1335 17980 1345
rect 18005 1415 18035 1425
rect 18005 1395 18010 1415
rect 18030 1395 18035 1415
rect 18005 1365 18035 1395
rect 18005 1345 18010 1365
rect 18030 1345 18035 1365
rect 18005 1335 18035 1345
rect 18060 1417 18130 1425
rect 18060 1415 18105 1417
rect 18060 1395 18065 1415
rect 18085 1395 18105 1415
rect 18125 1395 18130 1417
rect 18060 1365 18130 1395
rect 18060 1345 18065 1365
rect 18085 1345 18105 1365
rect 18125 1345 18130 1365
rect 18060 1335 18130 1345
rect 18310 1417 18380 1425
rect 18310 1345 18315 1417
rect 18335 1415 18380 1417
rect 18335 1345 18355 1415
rect 18375 1345 18380 1415
rect 18310 1335 18380 1345
rect 18405 1415 18435 1425
rect 18405 1345 18410 1415
rect 18430 1345 18435 1415
rect 18405 1335 18435 1345
rect 18460 1415 18490 1425
rect 18460 1345 18465 1415
rect 18485 1345 18490 1415
rect 18460 1335 18490 1345
rect 18515 1415 18545 1425
rect 18515 1345 18520 1415
rect 18540 1345 18545 1415
rect 18515 1335 18545 1345
rect 18570 1415 18600 1425
rect 18570 1345 18575 1415
rect 18595 1345 18600 1415
rect 18570 1335 18600 1345
rect 18625 1415 18655 1425
rect 18625 1345 18630 1415
rect 18650 1345 18655 1415
rect 18625 1335 18655 1345
rect 18680 1417 18750 1425
rect 18680 1415 18725 1417
rect 18680 1345 18685 1415
rect 18705 1345 18725 1415
rect 18745 1345 18750 1417
rect 18680 1335 18750 1345
rect 16440 1315 16460 1335
rect 16550 1315 16570 1335
rect 16950 1315 16970 1335
rect 17060 1315 17080 1335
rect 17170 1315 17190 1335
rect 17625 1315 17645 1335
rect 17735 1315 17755 1335
rect 17845 1315 17865 1335
rect 17955 1315 17975 1335
rect 18410 1315 18430 1335
rect 18520 1315 18540 1335
rect 18630 1315 18650 1335
rect 16430 1305 16470 1315
rect 16430 1285 16440 1305
rect 16460 1285 16470 1305
rect 16430 1275 16470 1285
rect 16540 1305 16580 1315
rect 16540 1285 16550 1305
rect 16570 1285 16580 1305
rect 16540 1275 16580 1285
rect 16940 1305 16980 1315
rect 16940 1285 16950 1305
rect 16970 1285 16980 1305
rect 16940 1275 16980 1285
rect 17050 1305 17090 1315
rect 17050 1285 17060 1305
rect 17080 1285 17090 1305
rect 17050 1275 17090 1285
rect 17160 1305 17200 1315
rect 17160 1285 17170 1305
rect 17190 1285 17200 1305
rect 17160 1275 17200 1285
rect 17615 1305 17655 1315
rect 17615 1285 17625 1305
rect 17645 1285 17655 1305
rect 17615 1275 17655 1285
rect 17725 1305 17765 1315
rect 17725 1285 17735 1305
rect 17755 1285 17765 1305
rect 17725 1275 17765 1285
rect 17835 1305 17875 1315
rect 17835 1285 17845 1305
rect 17865 1285 17875 1305
rect 17835 1275 17875 1285
rect 17945 1305 17985 1315
rect 17945 1285 17955 1305
rect 17975 1285 17985 1305
rect 17945 1275 17985 1285
rect 18400 1305 18440 1315
rect 18400 1285 18410 1305
rect 18430 1285 18440 1305
rect 18400 1275 18440 1285
rect 18510 1305 18550 1315
rect 18510 1285 18520 1305
rect 18540 1285 18550 1305
rect 18510 1275 18550 1285
rect 18620 1305 18660 1315
rect 18620 1285 18630 1305
rect 18650 1285 18660 1305
rect 18620 1275 18660 1285
rect 16970 1010 17010 1020
rect 16970 990 16980 1010
rect 17000 990 17010 1010
rect 16970 980 17010 990
rect 17150 1010 17190 1020
rect 17150 990 17160 1010
rect 17180 990 17190 1010
rect 17150 980 17190 990
rect 17330 1010 17370 1020
rect 17330 990 17340 1010
rect 17360 990 17370 1010
rect 17330 980 17370 990
rect 17510 1010 17550 1020
rect 17510 990 17520 1010
rect 17540 990 17550 1010
rect 17510 980 17550 990
rect 17690 1010 17730 1020
rect 17690 990 17700 1010
rect 17720 990 17730 1010
rect 17690 980 17730 990
rect 17870 1010 17910 1020
rect 17870 990 17880 1010
rect 17900 990 17910 1010
rect 17870 980 17910 990
rect 18050 1010 18090 1020
rect 18050 990 18060 1010
rect 18080 990 18090 1010
rect 18050 980 18090 990
rect 18230 1010 18270 1020
rect 18230 990 18240 1010
rect 18260 990 18270 1010
rect 18230 980 18270 990
rect 18410 1010 18450 1020
rect 18410 990 18420 1010
rect 18440 990 18450 1010
rect 18410 980 18450 990
rect 18590 1010 18630 1020
rect 18590 990 18600 1010
rect 18620 990 18630 1010
rect 18590 980 18630 990
rect 18905 1010 18945 1020
rect 18905 990 18915 1010
rect 18935 990 18945 1010
rect 18905 980 18945 990
rect 19015 1010 19055 1020
rect 19015 990 19025 1010
rect 19045 990 19055 1010
rect 19015 980 19055 990
rect 19075 1010 19115 1020
rect 19075 990 19085 1010
rect 19105 990 19115 1010
rect 19075 980 19115 990
rect 16980 960 17000 980
rect 17160 960 17180 980
rect 17340 960 17360 980
rect 17520 960 17540 980
rect 17700 960 17720 980
rect 17880 960 17900 980
rect 18060 960 18080 980
rect 18240 960 18260 980
rect 18420 960 18440 980
rect 18600 960 18620 980
rect 18915 960 18935 980
rect 19025 960 19045 980
rect 19080 960 19100 980
rect 16935 950 17005 960
rect 16935 930 16940 950
rect 16960 930 16980 950
rect 17000 930 17005 950
rect 16440 910 16470 920
rect 16440 890 16445 910
rect 16465 890 16470 910
rect 16440 860 16470 890
rect 16545 910 16585 920
rect 16545 890 16555 910
rect 16575 890 16585 910
rect 16545 880 16585 890
rect 16655 910 16695 920
rect 16655 890 16665 910
rect 16685 890 16695 910
rect 16655 880 16695 890
rect 16935 900 17005 930
rect 16935 880 16940 900
rect 16960 880 16980 900
rect 17000 880 17005 900
rect 16555 860 16575 880
rect 16660 860 16690 880
rect 16400 850 16470 860
rect 16400 830 16405 850
rect 16425 830 16445 850
rect 16465 830 16470 850
rect 16400 800 16470 830
rect 16400 780 16405 800
rect 16425 780 16445 800
rect 16465 780 16470 800
rect 16400 770 16470 780
rect 16495 850 16525 860
rect 16495 830 16500 850
rect 16520 830 16525 850
rect 16495 800 16525 830
rect 16495 780 16500 800
rect 16520 780 16525 800
rect 16495 770 16525 780
rect 16550 850 16580 860
rect 16550 830 16555 850
rect 16575 830 16580 850
rect 16550 800 16580 830
rect 16550 780 16555 800
rect 16575 780 16580 800
rect 16550 770 16580 780
rect 16605 850 16635 860
rect 16605 830 16610 850
rect 16630 830 16635 850
rect 16605 800 16635 830
rect 16605 780 16610 800
rect 16630 780 16635 800
rect 16605 770 16635 780
rect 16660 850 16735 860
rect 16660 830 16665 850
rect 16685 830 16710 850
rect 16730 830 16735 850
rect 16660 800 16735 830
rect 16660 780 16665 800
rect 16685 780 16710 800
rect 16730 780 16735 800
rect 16660 770 16735 780
rect 16935 850 17005 880
rect 16935 830 16940 850
rect 16960 830 16980 850
rect 17000 830 17005 850
rect 16935 800 17005 830
rect 16935 780 16940 800
rect 16960 780 16980 800
rect 17000 780 17005 800
rect 16500 750 16520 770
rect 16610 750 16630 770
rect 16935 750 17005 780
rect 16480 740 16520 750
rect 16480 720 16490 740
rect 16510 720 16520 740
rect 16480 710 16520 720
rect 16545 740 16585 750
rect 16545 720 16555 740
rect 16575 720 16585 740
rect 16545 710 16585 720
rect 16610 740 16650 750
rect 16610 720 16620 740
rect 16640 720 16650 740
rect 16610 710 16650 720
rect 16935 730 16940 750
rect 16960 730 16980 750
rect 17000 730 17005 750
rect 16935 700 17005 730
rect 16935 680 16940 700
rect 16960 680 16980 700
rect 17000 680 17005 700
rect 16935 670 17005 680
rect 17065 950 17095 960
rect 17065 930 17070 950
rect 17090 930 17095 950
rect 17065 900 17095 930
rect 17065 880 17070 900
rect 17090 880 17095 900
rect 17065 850 17095 880
rect 17065 830 17070 850
rect 17090 830 17095 850
rect 17065 800 17095 830
rect 17065 780 17070 800
rect 17090 780 17095 800
rect 17065 750 17095 780
rect 17065 730 17070 750
rect 17090 730 17095 750
rect 17065 700 17095 730
rect 17065 680 17070 700
rect 17090 680 17095 700
rect 17065 670 17095 680
rect 17155 950 17185 960
rect 17155 930 17160 950
rect 17180 930 17185 950
rect 17155 900 17185 930
rect 17155 880 17160 900
rect 17180 880 17185 900
rect 17155 850 17185 880
rect 17155 830 17160 850
rect 17180 830 17185 850
rect 17155 800 17185 830
rect 17155 780 17160 800
rect 17180 780 17185 800
rect 17155 750 17185 780
rect 17155 730 17160 750
rect 17180 730 17185 750
rect 17155 700 17185 730
rect 17155 680 17160 700
rect 17180 680 17185 700
rect 17155 670 17185 680
rect 17245 950 17275 960
rect 17245 930 17250 950
rect 17270 930 17275 950
rect 17245 900 17275 930
rect 17245 880 17250 900
rect 17270 880 17275 900
rect 17245 850 17275 880
rect 17245 830 17250 850
rect 17270 830 17275 850
rect 17245 800 17275 830
rect 17245 780 17250 800
rect 17270 780 17275 800
rect 17245 750 17275 780
rect 17245 730 17250 750
rect 17270 730 17275 750
rect 17245 700 17275 730
rect 17245 680 17250 700
rect 17270 680 17275 700
rect 17245 670 17275 680
rect 17335 950 17365 960
rect 17335 930 17340 950
rect 17360 930 17365 950
rect 17335 900 17365 930
rect 17335 880 17340 900
rect 17360 880 17365 900
rect 17335 850 17365 880
rect 17335 830 17340 850
rect 17360 830 17365 850
rect 17335 800 17365 830
rect 17335 780 17340 800
rect 17360 780 17365 800
rect 17335 750 17365 780
rect 17335 730 17340 750
rect 17360 730 17365 750
rect 17335 700 17365 730
rect 17335 680 17340 700
rect 17360 680 17365 700
rect 17335 670 17365 680
rect 17425 950 17455 960
rect 17425 930 17430 950
rect 17450 930 17455 950
rect 17425 900 17455 930
rect 17425 880 17430 900
rect 17450 880 17455 900
rect 17425 850 17455 880
rect 17425 830 17430 850
rect 17450 830 17455 850
rect 17425 800 17455 830
rect 17425 780 17430 800
rect 17450 780 17455 800
rect 17425 750 17455 780
rect 17425 730 17430 750
rect 17450 730 17455 750
rect 17425 700 17455 730
rect 17425 680 17430 700
rect 17450 680 17455 700
rect 17425 670 17455 680
rect 17515 950 17545 960
rect 17515 930 17520 950
rect 17540 930 17545 950
rect 17515 900 17545 930
rect 17515 880 17520 900
rect 17540 880 17545 900
rect 17515 850 17545 880
rect 17515 830 17520 850
rect 17540 830 17545 850
rect 17515 800 17545 830
rect 17515 780 17520 800
rect 17540 780 17545 800
rect 17515 750 17545 780
rect 17515 730 17520 750
rect 17540 730 17545 750
rect 17515 700 17545 730
rect 17515 680 17520 700
rect 17540 680 17545 700
rect 17515 670 17545 680
rect 17605 950 17635 960
rect 17605 930 17610 950
rect 17630 930 17635 950
rect 17605 900 17635 930
rect 17605 880 17610 900
rect 17630 880 17635 900
rect 17605 850 17635 880
rect 17605 830 17610 850
rect 17630 830 17635 850
rect 17605 800 17635 830
rect 17605 780 17610 800
rect 17630 780 17635 800
rect 17605 750 17635 780
rect 17605 730 17610 750
rect 17630 730 17635 750
rect 17605 700 17635 730
rect 17605 680 17610 700
rect 17630 680 17635 700
rect 17605 670 17635 680
rect 17695 950 17725 960
rect 17695 930 17700 950
rect 17720 930 17725 950
rect 17695 900 17725 930
rect 17695 880 17700 900
rect 17720 880 17725 900
rect 17695 850 17725 880
rect 17695 830 17700 850
rect 17720 830 17725 850
rect 17695 800 17725 830
rect 17695 780 17700 800
rect 17720 780 17725 800
rect 17695 750 17725 780
rect 17695 730 17700 750
rect 17720 730 17725 750
rect 17695 700 17725 730
rect 17695 680 17700 700
rect 17720 680 17725 700
rect 17695 670 17725 680
rect 17785 950 17815 960
rect 17785 930 17790 950
rect 17810 930 17815 950
rect 17785 900 17815 930
rect 17785 880 17790 900
rect 17810 880 17815 900
rect 17785 850 17815 880
rect 17785 830 17790 850
rect 17810 830 17815 850
rect 17785 800 17815 830
rect 17785 780 17790 800
rect 17810 780 17815 800
rect 17785 750 17815 780
rect 17785 730 17790 750
rect 17810 730 17815 750
rect 17785 700 17815 730
rect 17785 680 17790 700
rect 17810 680 17815 700
rect 17785 670 17815 680
rect 17875 950 17905 960
rect 17875 930 17880 950
rect 17900 930 17905 950
rect 17875 900 17905 930
rect 17875 880 17880 900
rect 17900 880 17905 900
rect 17875 850 17905 880
rect 17875 830 17880 850
rect 17900 830 17905 850
rect 17875 800 17905 830
rect 17875 780 17880 800
rect 17900 780 17905 800
rect 17875 750 17905 780
rect 17875 730 17880 750
rect 17900 730 17905 750
rect 17875 700 17905 730
rect 17875 680 17880 700
rect 17900 680 17905 700
rect 17875 670 17905 680
rect 17965 950 17995 960
rect 17965 930 17970 950
rect 17990 930 17995 950
rect 17965 900 17995 930
rect 17965 880 17970 900
rect 17990 880 17995 900
rect 17965 850 17995 880
rect 17965 830 17970 850
rect 17990 830 17995 850
rect 17965 800 17995 830
rect 17965 780 17970 800
rect 17990 780 17995 800
rect 17965 750 17995 780
rect 17965 730 17970 750
rect 17990 730 17995 750
rect 17965 700 17995 730
rect 17965 680 17970 700
rect 17990 680 17995 700
rect 17965 670 17995 680
rect 18055 950 18085 960
rect 18055 930 18060 950
rect 18080 930 18085 950
rect 18055 900 18085 930
rect 18055 880 18060 900
rect 18080 880 18085 900
rect 18055 850 18085 880
rect 18055 830 18060 850
rect 18080 830 18085 850
rect 18055 800 18085 830
rect 18055 780 18060 800
rect 18080 780 18085 800
rect 18055 750 18085 780
rect 18055 730 18060 750
rect 18080 730 18085 750
rect 18055 700 18085 730
rect 18055 680 18060 700
rect 18080 680 18085 700
rect 18055 670 18085 680
rect 18145 950 18175 960
rect 18145 930 18150 950
rect 18170 930 18175 950
rect 18145 900 18175 930
rect 18145 880 18150 900
rect 18170 880 18175 900
rect 18145 850 18175 880
rect 18145 830 18150 850
rect 18170 830 18175 850
rect 18145 800 18175 830
rect 18145 780 18150 800
rect 18170 780 18175 800
rect 18145 750 18175 780
rect 18145 730 18150 750
rect 18170 730 18175 750
rect 18145 700 18175 730
rect 18145 680 18150 700
rect 18170 680 18175 700
rect 18145 670 18175 680
rect 18235 950 18265 960
rect 18235 930 18240 950
rect 18260 930 18265 950
rect 18235 900 18265 930
rect 18235 880 18240 900
rect 18260 880 18265 900
rect 18235 850 18265 880
rect 18235 830 18240 850
rect 18260 830 18265 850
rect 18235 800 18265 830
rect 18235 780 18240 800
rect 18260 780 18265 800
rect 18235 750 18265 780
rect 18235 730 18240 750
rect 18260 730 18265 750
rect 18235 700 18265 730
rect 18235 680 18240 700
rect 18260 680 18265 700
rect 18235 670 18265 680
rect 18325 950 18355 960
rect 18325 930 18330 950
rect 18350 930 18355 950
rect 18325 900 18355 930
rect 18325 880 18330 900
rect 18350 880 18355 900
rect 18325 850 18355 880
rect 18325 830 18330 850
rect 18350 830 18355 850
rect 18325 800 18355 830
rect 18325 780 18330 800
rect 18350 780 18355 800
rect 18325 750 18355 780
rect 18325 730 18330 750
rect 18350 730 18355 750
rect 18325 700 18355 730
rect 18325 680 18330 700
rect 18350 680 18355 700
rect 18325 670 18355 680
rect 18415 950 18445 960
rect 18415 930 18420 950
rect 18440 930 18445 950
rect 18415 900 18445 930
rect 18415 880 18420 900
rect 18440 880 18445 900
rect 18415 850 18445 880
rect 18415 830 18420 850
rect 18440 830 18445 850
rect 18415 800 18445 830
rect 18415 780 18420 800
rect 18440 780 18445 800
rect 18415 750 18445 780
rect 18415 730 18420 750
rect 18440 730 18445 750
rect 18415 700 18445 730
rect 18415 680 18420 700
rect 18440 680 18445 700
rect 18415 670 18445 680
rect 18505 950 18535 960
rect 18505 930 18510 950
rect 18530 930 18535 950
rect 18505 900 18535 930
rect 18505 880 18510 900
rect 18530 880 18535 900
rect 18505 850 18535 880
rect 18505 830 18510 850
rect 18530 830 18535 850
rect 18505 800 18535 830
rect 18505 780 18510 800
rect 18530 780 18535 800
rect 18505 750 18535 780
rect 18505 730 18510 750
rect 18530 730 18535 750
rect 18505 700 18535 730
rect 18505 680 18510 700
rect 18530 680 18535 700
rect 18505 670 18535 680
rect 18595 950 18665 960
rect 18595 930 18600 950
rect 18620 930 18640 950
rect 18660 930 18665 950
rect 18595 900 18665 930
rect 18595 880 18600 900
rect 18620 880 18640 900
rect 18660 880 18665 900
rect 18595 850 18665 880
rect 18595 830 18600 850
rect 18620 830 18640 850
rect 18660 830 18665 850
rect 18595 800 18665 830
rect 18595 780 18600 800
rect 18620 780 18640 800
rect 18660 780 18665 800
rect 18595 750 18665 780
rect 18870 950 18940 960
rect 18870 930 18875 950
rect 18895 930 18915 950
rect 18935 930 18940 950
rect 18870 900 18940 930
rect 18870 880 18875 900
rect 18895 880 18915 900
rect 18935 880 18940 900
rect 18870 850 18940 880
rect 18870 830 18875 850
rect 18895 830 18915 850
rect 18935 830 18940 850
rect 18870 800 18940 830
rect 18870 780 18875 800
rect 18895 780 18915 800
rect 18935 780 18940 800
rect 18870 770 18940 780
rect 18965 950 18995 960
rect 18965 930 18970 950
rect 18990 930 18995 950
rect 18965 900 18995 930
rect 18965 880 18970 900
rect 18990 880 18995 900
rect 18965 850 18995 880
rect 18965 830 18970 850
rect 18990 830 18995 850
rect 18965 800 18995 830
rect 18965 780 18970 800
rect 18990 780 18995 800
rect 18965 770 18995 780
rect 19020 950 19050 960
rect 19020 930 19025 950
rect 19045 930 19050 950
rect 19020 900 19050 930
rect 19020 880 19025 900
rect 19045 880 19050 900
rect 19020 850 19050 880
rect 19020 830 19025 850
rect 19045 830 19050 850
rect 19020 800 19050 830
rect 19020 780 19025 800
rect 19045 780 19050 800
rect 19020 770 19050 780
rect 19075 950 19145 960
rect 19075 930 19080 950
rect 19100 930 19120 950
rect 19140 930 19145 950
rect 19075 900 19145 930
rect 19075 880 19080 900
rect 19100 880 19120 900
rect 19140 880 19145 900
rect 19075 850 19145 880
rect 19075 830 19080 850
rect 19100 830 19120 850
rect 19140 830 19145 850
rect 19075 800 19145 830
rect 19075 780 19080 800
rect 19100 780 19120 800
rect 19140 780 19145 800
rect 19075 770 19145 780
rect 18970 750 18990 770
rect 18595 730 18600 750
rect 18620 730 18640 750
rect 18660 730 18665 750
rect 18595 700 18665 730
rect 18950 740 18990 750
rect 18950 720 18960 740
rect 18980 720 18990 740
rect 18950 710 18990 720
rect 18595 680 18600 700
rect 18620 680 18640 700
rect 18660 680 18665 700
rect 18595 670 18665 680
rect 19000 680 19040 690
rect 17070 650 17090 670
rect 17250 650 17270 670
rect 17430 650 17450 670
rect 17610 650 17630 670
rect 17790 650 17810 670
rect 17970 650 17990 670
rect 18150 650 18170 670
rect 18330 650 18350 670
rect 18510 650 18530 670
rect 19000 660 19010 680
rect 19030 660 19040 680
rect 19000 650 19040 660
rect 17060 640 17100 650
rect 17060 620 17070 640
rect 17090 620 17100 640
rect 17060 610 17100 620
rect 17240 640 17280 650
rect 17240 620 17250 640
rect 17270 620 17280 640
rect 17240 610 17280 620
rect 17420 640 17460 650
rect 17420 620 17430 640
rect 17450 620 17460 640
rect 17420 610 17460 620
rect 17600 640 17640 650
rect 17600 620 17610 640
rect 17630 620 17640 640
rect 17600 610 17640 620
rect 17690 640 17730 650
rect 17690 620 17700 640
rect 17720 620 17730 640
rect 17690 610 17730 620
rect 17780 640 17820 650
rect 17780 620 17790 640
rect 17810 620 17820 640
rect 17780 610 17820 620
rect 17960 640 18000 650
rect 17960 620 17970 640
rect 17990 620 18000 640
rect 17960 610 18000 620
rect 18140 640 18180 650
rect 18140 620 18150 640
rect 18170 620 18180 640
rect 18140 610 18180 620
rect 18320 640 18360 650
rect 18320 620 18330 640
rect 18350 620 18360 640
rect 18320 610 18360 620
rect 18500 640 18540 650
rect 18500 620 18510 640
rect 18530 620 18540 640
rect 18500 610 18540 620
rect 16425 170 16455 180
rect 16425 150 16430 170
rect 16450 150 16455 170
rect 16425 120 16455 150
rect 16480 170 16520 180
rect 16480 150 16490 170
rect 16510 150 16520 170
rect 16480 140 16520 150
rect 16545 170 16575 180
rect 16545 150 16550 170
rect 16570 150 16575 170
rect 16545 140 16575 150
rect 16665 170 16695 180
rect 16665 150 16670 170
rect 16690 150 16695 170
rect 16665 140 16695 150
rect 16785 170 16815 180
rect 16785 150 16790 170
rect 16810 150 16815 170
rect 16785 140 16815 150
rect 16840 170 16880 180
rect 16840 150 16850 170
rect 16870 150 16880 170
rect 16840 140 16880 150
rect 16905 170 16935 180
rect 16905 150 16910 170
rect 16930 150 16935 170
rect 16905 140 16935 150
rect 17025 170 17055 180
rect 17025 150 17030 170
rect 17050 150 17055 170
rect 17025 140 17055 150
rect 17145 170 17175 180
rect 17145 150 17150 170
rect 17170 150 17175 170
rect 17145 140 17175 150
rect 17200 170 17240 180
rect 17200 150 17210 170
rect 17230 150 17240 170
rect 17200 140 17240 150
rect 17265 170 17295 180
rect 17265 150 17270 170
rect 17290 150 17295 170
rect 17265 140 17295 150
rect 17385 170 17415 180
rect 17385 150 17390 170
rect 17410 150 17415 170
rect 17385 140 17415 150
rect 17505 170 17535 180
rect 17505 150 17510 170
rect 17530 150 17535 170
rect 17505 140 17535 150
rect 17560 170 17600 180
rect 17560 150 17570 170
rect 17590 150 17600 170
rect 17560 140 17600 150
rect 17625 170 17655 180
rect 17625 150 17630 170
rect 17650 150 17655 170
rect 16490 120 16510 140
rect 16550 120 16570 140
rect 16670 120 16690 140
rect 16790 120 16810 140
rect 16850 120 16870 140
rect 16910 120 16930 140
rect 17030 120 17050 140
rect 17150 120 17170 140
rect 17210 120 17230 140
rect 17270 120 17290 140
rect 17390 120 17410 140
rect 17510 120 17530 140
rect 17570 120 17590 140
rect 17625 120 17655 150
rect 17945 170 17975 180
rect 17945 150 17950 170
rect 17970 150 17975 170
rect 17945 120 17975 150
rect 18000 170 18040 180
rect 18000 150 18010 170
rect 18030 150 18040 170
rect 18000 140 18040 150
rect 18065 170 18095 180
rect 18065 150 18070 170
rect 18090 150 18095 170
rect 18065 140 18095 150
rect 18185 170 18215 180
rect 18185 150 18190 170
rect 18210 150 18215 170
rect 18185 140 18215 150
rect 18305 170 18335 180
rect 18305 150 18310 170
rect 18330 150 18335 170
rect 18305 140 18335 150
rect 18360 170 18400 180
rect 18360 150 18370 170
rect 18390 150 18400 170
rect 18360 140 18400 150
rect 18425 170 18455 180
rect 18425 150 18430 170
rect 18450 150 18455 170
rect 18425 140 18455 150
rect 18545 170 18575 180
rect 18545 150 18550 170
rect 18570 150 18575 170
rect 18545 140 18575 150
rect 18665 170 18695 180
rect 18665 150 18670 170
rect 18690 150 18695 170
rect 18665 140 18695 150
rect 18720 170 18760 180
rect 18720 150 18730 170
rect 18750 150 18760 170
rect 18720 140 18760 150
rect 18785 170 18815 180
rect 18785 150 18790 170
rect 18810 150 18815 170
rect 18785 140 18815 150
rect 18905 170 18935 180
rect 18905 150 18910 170
rect 18930 150 18935 170
rect 18905 140 18935 150
rect 19025 170 19055 180
rect 19025 150 19030 170
rect 19050 150 19055 170
rect 19025 140 19055 150
rect 19080 170 19120 180
rect 19080 150 19090 170
rect 19110 150 19120 170
rect 19080 140 19120 150
rect 19145 170 19175 180
rect 19145 150 19150 170
rect 19170 150 19175 170
rect 18010 120 18030 140
rect 18070 120 18090 140
rect 18190 120 18210 140
rect 18310 120 18330 140
rect 18370 120 18390 140
rect 18430 120 18450 140
rect 18550 120 18570 140
rect 18670 120 18690 140
rect 18730 120 18750 140
rect 18790 120 18810 140
rect 18910 120 18930 140
rect 19030 120 19050 140
rect 19090 120 19110 140
rect 19145 120 19175 150
rect 16385 110 16455 120
rect 16385 90 16390 110
rect 16410 90 16430 110
rect 16450 90 16455 110
rect 16385 60 16455 90
rect 16385 40 16390 60
rect 16410 40 16430 60
rect 16450 40 16455 60
rect 16385 30 16455 40
rect 16485 110 16515 120
rect 16485 90 16490 110
rect 16510 90 16515 110
rect 16485 60 16515 90
rect 16485 40 16490 60
rect 16510 40 16515 60
rect 16485 30 16515 40
rect 16545 110 16575 120
rect 16545 90 16550 110
rect 16570 90 16575 110
rect 16545 60 16575 90
rect 16545 40 16550 60
rect 16570 40 16575 60
rect 16545 30 16575 40
rect 16605 110 16635 120
rect 16605 90 16610 110
rect 16630 90 16635 110
rect 16605 60 16635 90
rect 16605 40 16610 60
rect 16630 40 16635 60
rect 16605 30 16635 40
rect 16665 110 16695 120
rect 16665 90 16670 110
rect 16690 90 16695 110
rect 16665 60 16695 90
rect 16665 40 16670 60
rect 16690 40 16695 60
rect 16665 30 16695 40
rect 16725 110 16755 120
rect 16725 90 16730 110
rect 16750 90 16755 110
rect 16725 60 16755 90
rect 16725 40 16730 60
rect 16750 40 16755 60
rect 16725 30 16755 40
rect 16785 110 16815 120
rect 16785 90 16790 110
rect 16810 90 16815 110
rect 16785 60 16815 90
rect 16785 40 16790 60
rect 16810 40 16815 60
rect 16785 30 16815 40
rect 16845 110 16875 120
rect 16845 90 16850 110
rect 16870 90 16875 110
rect 16845 60 16875 90
rect 16845 40 16850 60
rect 16870 40 16875 60
rect 16845 30 16875 40
rect 16905 110 16935 120
rect 16905 90 16910 110
rect 16930 90 16935 110
rect 16905 60 16935 90
rect 16905 40 16910 60
rect 16930 40 16935 60
rect 16905 30 16935 40
rect 16965 110 16995 120
rect 16965 90 16970 110
rect 16990 90 16995 110
rect 16965 60 16995 90
rect 16965 40 16970 60
rect 16990 40 16995 60
rect 16965 30 16995 40
rect 17025 110 17055 120
rect 17025 90 17030 110
rect 17050 90 17055 110
rect 17025 60 17055 90
rect 17025 40 17030 60
rect 17050 40 17055 60
rect 17025 30 17055 40
rect 17085 110 17115 120
rect 17085 90 17090 110
rect 17110 90 17115 110
rect 17085 60 17115 90
rect 17085 40 17090 60
rect 17110 40 17115 60
rect 17085 30 17115 40
rect 17145 110 17175 120
rect 17145 90 17150 110
rect 17170 90 17175 110
rect 17145 60 17175 90
rect 17145 40 17150 60
rect 17170 40 17175 60
rect 17145 30 17175 40
rect 17205 110 17235 120
rect 17205 90 17210 110
rect 17230 90 17235 110
rect 17205 60 17235 90
rect 17205 40 17210 60
rect 17230 40 17235 60
rect 17205 30 17235 40
rect 17265 110 17295 120
rect 17265 90 17270 110
rect 17290 90 17295 110
rect 17265 60 17295 90
rect 17265 40 17270 60
rect 17290 40 17295 60
rect 17265 30 17295 40
rect 17325 110 17355 120
rect 17325 90 17330 110
rect 17350 90 17355 110
rect 17325 60 17355 90
rect 17325 40 17330 60
rect 17350 40 17355 60
rect 17325 30 17355 40
rect 17385 110 17415 120
rect 17385 90 17390 110
rect 17410 90 17415 110
rect 17385 60 17415 90
rect 17385 40 17390 60
rect 17410 40 17415 60
rect 17385 30 17415 40
rect 17445 110 17475 120
rect 17445 90 17450 110
rect 17470 90 17475 110
rect 17445 60 17475 90
rect 17445 40 17450 60
rect 17470 40 17475 60
rect 17445 30 17475 40
rect 17505 110 17535 120
rect 17505 90 17510 110
rect 17530 90 17535 110
rect 17505 60 17535 90
rect 17505 40 17510 60
rect 17530 40 17535 60
rect 17505 30 17535 40
rect 17565 110 17595 120
rect 17565 90 17570 110
rect 17590 90 17595 110
rect 17565 60 17595 90
rect 17565 40 17570 60
rect 17590 40 17595 60
rect 17565 30 17595 40
rect 17625 110 17695 120
rect 17625 90 17630 110
rect 17650 90 17670 110
rect 17690 90 17695 110
rect 17625 60 17695 90
rect 17625 40 17630 60
rect 17650 40 17670 60
rect 17690 40 17695 60
rect 17625 30 17695 40
rect 17905 110 17975 120
rect 17905 90 17910 110
rect 17930 90 17950 110
rect 17970 90 17975 110
rect 17905 60 17975 90
rect 17905 40 17910 60
rect 17930 40 17950 60
rect 17970 40 17975 60
rect 17905 30 17975 40
rect 18005 110 18035 120
rect 18005 90 18010 110
rect 18030 90 18035 110
rect 18005 60 18035 90
rect 18005 40 18010 60
rect 18030 40 18035 60
rect 18005 30 18035 40
rect 18065 110 18095 120
rect 18065 90 18070 110
rect 18090 90 18095 110
rect 18065 60 18095 90
rect 18065 40 18070 60
rect 18090 40 18095 60
rect 18065 30 18095 40
rect 18125 110 18155 120
rect 18125 90 18130 110
rect 18150 90 18155 110
rect 18125 60 18155 90
rect 18125 40 18130 60
rect 18150 40 18155 60
rect 18125 30 18155 40
rect 18185 110 18215 120
rect 18185 90 18190 110
rect 18210 90 18215 110
rect 18185 60 18215 90
rect 18185 40 18190 60
rect 18210 40 18215 60
rect 18185 30 18215 40
rect 18245 110 18275 120
rect 18245 90 18250 110
rect 18270 90 18275 110
rect 18245 60 18275 90
rect 18245 40 18250 60
rect 18270 40 18275 60
rect 18245 30 18275 40
rect 18305 110 18335 120
rect 18305 90 18310 110
rect 18330 90 18335 110
rect 18305 60 18335 90
rect 18305 40 18310 60
rect 18330 40 18335 60
rect 18305 30 18335 40
rect 18365 110 18395 120
rect 18365 90 18370 110
rect 18390 90 18395 110
rect 18365 60 18395 90
rect 18365 40 18370 60
rect 18390 40 18395 60
rect 18365 30 18395 40
rect 18425 110 18455 120
rect 18425 90 18430 110
rect 18450 90 18455 110
rect 18425 60 18455 90
rect 18425 40 18430 60
rect 18450 40 18455 60
rect 18425 30 18455 40
rect 18485 110 18515 120
rect 18485 90 18490 110
rect 18510 90 18515 110
rect 18485 60 18515 90
rect 18485 40 18490 60
rect 18510 40 18515 60
rect 18485 30 18515 40
rect 18545 110 18575 120
rect 18545 90 18550 110
rect 18570 90 18575 110
rect 18545 60 18575 90
rect 18545 40 18550 60
rect 18570 40 18575 60
rect 18545 30 18575 40
rect 18605 110 18635 120
rect 18605 90 18610 110
rect 18630 90 18635 110
rect 18605 60 18635 90
rect 18605 40 18610 60
rect 18630 40 18635 60
rect 18605 30 18635 40
rect 18665 110 18695 120
rect 18665 90 18670 110
rect 18690 90 18695 110
rect 18665 60 18695 90
rect 18665 40 18670 60
rect 18690 40 18695 60
rect 18665 30 18695 40
rect 18725 110 18755 120
rect 18725 90 18730 110
rect 18750 90 18755 110
rect 18725 60 18755 90
rect 18725 40 18730 60
rect 18750 40 18755 60
rect 18725 30 18755 40
rect 18785 110 18815 120
rect 18785 90 18790 110
rect 18810 90 18815 110
rect 18785 60 18815 90
rect 18785 40 18790 60
rect 18810 40 18815 60
rect 18785 30 18815 40
rect 18845 110 18875 120
rect 18845 90 18850 110
rect 18870 90 18875 110
rect 18845 60 18875 90
rect 18845 40 18850 60
rect 18870 40 18875 60
rect 18845 30 18875 40
rect 18905 110 18935 120
rect 18905 90 18910 110
rect 18930 90 18935 110
rect 18905 60 18935 90
rect 18905 40 18910 60
rect 18930 40 18935 60
rect 18905 30 18935 40
rect 18965 110 18995 120
rect 18965 90 18970 110
rect 18990 90 18995 110
rect 18965 60 18995 90
rect 18965 40 18970 60
rect 18990 40 18995 60
rect 18965 30 18995 40
rect 19025 110 19055 120
rect 19025 90 19030 110
rect 19050 90 19055 110
rect 19025 60 19055 90
rect 19025 40 19030 60
rect 19050 40 19055 60
rect 19025 30 19055 40
rect 19085 110 19115 120
rect 19085 90 19090 110
rect 19110 90 19115 110
rect 19085 60 19115 90
rect 19085 40 19090 60
rect 19110 40 19115 60
rect 19085 30 19115 40
rect 19145 110 19215 120
rect 19145 90 19150 110
rect 19170 90 19190 110
rect 19210 90 19215 110
rect 19145 60 19215 90
rect 19145 40 19150 60
rect 19170 40 19190 60
rect 19210 40 19215 60
rect 19145 30 19215 40
rect 16425 0 16455 30
rect 16610 10 16630 30
rect 16730 10 16750 30
rect 16970 10 16990 30
rect 17090 10 17110 30
rect 17330 10 17350 30
rect 17450 10 17470 30
rect 16425 -20 16430 0
rect 16450 -20 16455 0
rect 16425 -30 16455 -20
rect 16510 0 16550 10
rect 16510 -20 16520 0
rect 16540 -20 16550 0
rect 16510 -30 16550 -20
rect 16600 0 16640 10
rect 16600 -20 16610 0
rect 16630 -20 16640 0
rect 16600 -30 16640 -20
rect 16720 0 16760 10
rect 16720 -20 16730 0
rect 16750 -20 16760 0
rect 16720 -30 16760 -20
rect 16840 0 16880 10
rect 16840 -20 16850 0
rect 16870 -20 16880 0
rect 16840 -30 16880 -20
rect 16960 0 17000 10
rect 16960 -20 16970 0
rect 16990 -20 17000 0
rect 16960 -30 17000 -20
rect 17080 0 17120 10
rect 17080 -20 17090 0
rect 17110 -20 17120 0
rect 17080 -30 17120 -20
rect 17200 0 17240 10
rect 17200 -20 17210 0
rect 17230 -20 17240 0
rect 17200 -30 17240 -20
rect 17320 0 17360 10
rect 17320 -20 17330 0
rect 17350 -20 17360 0
rect 17320 -30 17360 -20
rect 17440 0 17480 10
rect 17440 -20 17450 0
rect 17470 -20 17480 0
rect 17440 -30 17480 -20
rect 17535 0 17565 10
rect 17535 -20 17540 0
rect 17560 -20 17565 0
rect 17535 -30 17565 -20
rect 17945 0 17975 30
rect 18130 10 18150 30
rect 18250 10 18270 30
rect 18490 10 18510 30
rect 18610 10 18630 30
rect 18850 10 18870 30
rect 18970 10 18990 30
rect 19145 25 19180 30
rect 17945 -20 17950 0
rect 17970 -20 17975 0
rect 17945 -30 17975 -20
rect 18035 0 18065 10
rect 18035 -20 18040 0
rect 18060 -20 18065 0
rect 18035 -30 18065 -20
rect 18120 0 18160 10
rect 18120 -20 18130 0
rect 18150 -20 18160 0
rect 18120 -30 18160 -20
rect 18240 0 18280 10
rect 18240 -20 18250 0
rect 18270 -20 18280 0
rect 18240 -30 18280 -20
rect 18360 0 18400 10
rect 18360 -20 18370 0
rect 18390 -20 18400 0
rect 18360 -30 18400 -20
rect 18480 0 18520 10
rect 18480 -20 18490 0
rect 18510 -20 18520 0
rect 18480 -30 18520 -20
rect 18600 0 18640 10
rect 18600 -20 18610 0
rect 18630 -20 18640 0
rect 18600 -30 18640 -20
rect 18720 0 18760 10
rect 18720 -20 18730 0
rect 18750 -20 18760 0
rect 18720 -30 18760 -20
rect 18840 0 18880 10
rect 18840 -20 18850 0
rect 18870 -20 18880 0
rect 18840 -30 18880 -20
rect 18960 0 19000 10
rect 18960 -20 18970 0
rect 18990 -20 19000 0
rect 18960 -30 19000 -20
rect 19050 0 19090 10
rect 19050 -20 19060 0
rect 19080 -20 19090 0
rect 19050 -30 19090 -20
rect 19145 0 19175 25
rect 19145 -20 19150 0
rect 19170 -20 19175 0
rect 19145 -30 19175 -20
rect 16960 -115 16990 -105
rect 16960 -135 16965 -115
rect 16985 -135 16990 -115
rect 16960 -145 16990 -135
rect 17007 -115 17037 -105
rect 17007 -135 17012 -115
rect 17032 -135 17037 -115
rect 17007 -145 17037 -135
rect 17090 -115 17120 -105
rect 17090 -135 17095 -115
rect 17115 -135 17120 -115
rect 17090 -145 17120 -135
rect 18480 -115 18510 -105
rect 18480 -135 18485 -115
rect 18505 -135 18510 -115
rect 18480 -145 18510 -135
rect 18563 -115 18593 -105
rect 18563 -135 18568 -115
rect 18588 -135 18593 -115
rect 18563 -145 18593 -135
rect 18610 -115 18640 -105
rect 18610 -135 18615 -115
rect 18635 -135 18640 -115
rect 18610 -145 18640 -135
rect 16970 -165 16990 -145
rect 17090 -165 17110 -145
rect 18490 -165 18510 -145
rect 18610 -165 18630 -145
rect 16965 -175 16995 -165
rect 16965 -195 16970 -175
rect 16990 -195 16995 -175
rect 16965 -225 16995 -195
rect 16965 -245 16970 -225
rect 16990 -245 16995 -225
rect 16965 -275 16995 -245
rect 16965 -295 16970 -275
rect 16990 -295 16995 -275
rect 16965 -325 16995 -295
rect 16965 -345 16970 -325
rect 16990 -345 16995 -325
rect 16965 -375 16995 -345
rect 16965 -395 16970 -375
rect 16990 -395 16995 -375
rect 16965 -405 16995 -395
rect 17025 -175 17055 -165
rect 17025 -195 17030 -175
rect 17050 -195 17055 -175
rect 17025 -225 17055 -195
rect 17025 -245 17030 -225
rect 17050 -245 17055 -225
rect 17025 -275 17055 -245
rect 17025 -295 17030 -275
rect 17050 -295 17055 -275
rect 17025 -325 17055 -295
rect 17025 -345 17030 -325
rect 17050 -345 17055 -325
rect 17025 -375 17055 -345
rect 17025 -395 17030 -375
rect 17050 -395 17055 -375
rect 17025 -405 17055 -395
rect 17085 -175 17115 -165
rect 17085 -195 17090 -175
rect 17110 -195 17115 -175
rect 17085 -225 17115 -195
rect 17085 -245 17090 -225
rect 17110 -245 17115 -225
rect 17085 -275 17115 -245
rect 17085 -295 17090 -275
rect 17110 -295 17115 -275
rect 17560 -175 17600 -165
rect 17560 -195 17570 -175
rect 17590 -195 17600 -175
rect 17560 -215 17600 -195
rect 17560 -235 17570 -215
rect 17590 -235 17600 -215
rect 17560 -255 17600 -235
rect 17560 -275 17570 -255
rect 17590 -275 17600 -255
rect 17560 -285 17600 -275
rect 18000 -175 18040 -165
rect 18000 -195 18010 -175
rect 18030 -195 18040 -175
rect 18000 -215 18040 -195
rect 18000 -235 18010 -215
rect 18030 -235 18040 -215
rect 18000 -255 18040 -235
rect 18000 -275 18010 -255
rect 18030 -275 18040 -255
rect 18000 -285 18040 -275
rect 18485 -175 18515 -165
rect 18485 -195 18490 -175
rect 18510 -195 18515 -175
rect 18485 -225 18515 -195
rect 18485 -245 18490 -225
rect 18510 -245 18515 -225
rect 18485 -275 18515 -245
rect 17085 -325 17115 -295
rect 17085 -345 17090 -325
rect 17110 -345 17115 -325
rect 17085 -375 17115 -345
rect 17085 -395 17090 -375
rect 17110 -395 17115 -375
rect 17085 -405 17115 -395
rect 18485 -295 18490 -275
rect 18510 -295 18515 -275
rect 18485 -325 18515 -295
rect 18485 -345 18490 -325
rect 18510 -345 18515 -325
rect 18485 -375 18515 -345
rect 18485 -395 18490 -375
rect 18510 -395 18515 -375
rect 18485 -405 18515 -395
rect 18545 -175 18575 -165
rect 18545 -195 18550 -175
rect 18570 -195 18575 -175
rect 18545 -225 18575 -195
rect 18545 -245 18550 -225
rect 18570 -245 18575 -225
rect 18545 -275 18575 -245
rect 18545 -295 18550 -275
rect 18570 -295 18575 -275
rect 18545 -325 18575 -295
rect 18545 -345 18550 -325
rect 18570 -345 18575 -325
rect 18545 -375 18575 -345
rect 18545 -395 18550 -375
rect 18570 -395 18575 -375
rect 18545 -405 18575 -395
rect 18605 -175 18635 -165
rect 18605 -195 18610 -175
rect 18630 -195 18635 -175
rect 18605 -225 18635 -195
rect 18605 -245 18610 -225
rect 18630 -245 18635 -225
rect 18605 -275 18635 -245
rect 18605 -295 18610 -275
rect 18630 -295 18635 -275
rect 18605 -325 18635 -295
rect 18605 -345 18610 -325
rect 18630 -345 18635 -325
rect 18605 -375 18635 -345
rect 18605 -395 18610 -375
rect 18630 -395 18635 -375
rect 18605 -405 18635 -395
rect 18550 -425 18570 -405
rect 17075 -435 17105 -425
rect 17075 -455 17080 -435
rect 17100 -455 17105 -435
rect 17075 -465 17105 -455
rect 18495 -435 18525 -425
rect 18495 -455 18500 -435
rect 18520 -455 18525 -435
rect 18495 -465 18525 -455
rect 18545 -435 18575 -425
rect 18545 -455 18550 -435
rect 18570 -455 18575 -435
rect 18545 -465 18575 -455
rect 16620 -650 16660 -640
rect 16620 -670 16630 -650
rect 16650 -670 16660 -650
rect 16620 -680 16660 -670
rect 16740 -650 16780 -640
rect 16740 -670 16750 -650
rect 16770 -670 16780 -650
rect 16740 -680 16780 -670
rect 16860 -650 16900 -640
rect 16860 -670 16870 -650
rect 16890 -670 16900 -650
rect 16860 -680 16900 -670
rect 16980 -650 17020 -640
rect 16980 -670 16990 -650
rect 17010 -670 17020 -650
rect 16980 -680 17020 -670
rect 17300 -650 17340 -640
rect 17300 -670 17310 -650
rect 17330 -670 17340 -650
rect 17300 -680 17340 -670
rect 17420 -650 17460 -640
rect 17420 -670 17430 -650
rect 17450 -670 17460 -650
rect 17420 -680 17460 -670
rect 17540 -650 17580 -640
rect 17540 -670 17550 -650
rect 17570 -670 17580 -650
rect 18020 -650 18060 -640
rect 17540 -680 17580 -670
rect 17695 -665 17725 -655
rect 17695 -685 17700 -665
rect 17720 -685 17725 -665
rect 16535 -710 16565 -700
rect 16535 -730 16540 -710
rect 16560 -730 16565 -710
rect 16535 -760 16565 -730
rect 16535 -780 16540 -760
rect 16560 -780 16565 -760
rect 16535 -810 16565 -780
rect 16535 -830 16540 -810
rect 16560 -830 16565 -810
rect 16535 -860 16565 -830
rect 16535 -880 16540 -860
rect 16560 -880 16565 -860
rect 16535 -910 16565 -880
rect 16535 -930 16540 -910
rect 16560 -930 16565 -910
rect 16535 -940 16565 -930
rect 17075 -710 17185 -700
rect 17075 -730 17080 -710
rect 17100 -730 17120 -710
rect 17140 -730 17160 -710
rect 17180 -730 17185 -710
rect 17075 -760 17185 -730
rect 17075 -780 17080 -760
rect 17100 -780 17120 -760
rect 17140 -780 17160 -760
rect 17180 -780 17185 -760
rect 17075 -810 17185 -780
rect 17075 -830 17080 -810
rect 17100 -830 17120 -810
rect 17140 -830 17160 -810
rect 17180 -830 17185 -810
rect 17075 -860 17185 -830
rect 17075 -880 17080 -860
rect 17100 -880 17120 -860
rect 17140 -880 17160 -860
rect 17180 -880 17185 -860
rect 17075 -910 17185 -880
rect 17075 -930 17080 -910
rect 17100 -930 17120 -910
rect 17140 -930 17160 -910
rect 17180 -930 17185 -910
rect 17075 -940 17185 -930
rect 17695 -710 17725 -685
rect 17695 -730 17700 -710
rect 17720 -730 17725 -710
rect 17695 -760 17725 -730
rect 17695 -780 17700 -760
rect 17720 -780 17725 -760
rect 17695 -810 17725 -780
rect 17695 -830 17700 -810
rect 17720 -830 17725 -810
rect 17695 -860 17725 -830
rect 17695 -880 17700 -860
rect 17720 -880 17725 -860
rect 17695 -910 17725 -880
rect 17695 -930 17700 -910
rect 17720 -930 17725 -910
rect 17695 -940 17725 -930
rect 17875 -665 17905 -655
rect 17875 -685 17880 -665
rect 17900 -685 17905 -665
rect 18020 -670 18030 -650
rect 18050 -670 18060 -650
rect 18020 -680 18060 -670
rect 18140 -650 18180 -640
rect 18140 -670 18150 -650
rect 18170 -670 18180 -650
rect 18140 -680 18180 -670
rect 18260 -650 18300 -640
rect 18260 -670 18270 -650
rect 18290 -670 18300 -650
rect 18260 -680 18300 -670
rect 18580 -650 18620 -640
rect 18580 -670 18590 -650
rect 18610 -670 18620 -650
rect 18580 -680 18620 -670
rect 18700 -650 18740 -640
rect 18700 -670 18710 -650
rect 18730 -670 18740 -650
rect 18700 -680 18740 -670
rect 18820 -650 18860 -640
rect 18820 -670 18830 -650
rect 18850 -670 18860 -650
rect 18820 -680 18860 -670
rect 18940 -650 18980 -640
rect 18940 -670 18950 -650
rect 18970 -670 18980 -650
rect 18940 -680 18980 -670
rect 19030 -670 19070 -660
rect 17875 -710 17905 -685
rect 19030 -690 19040 -670
rect 19060 -690 19070 -670
rect 19030 -700 19070 -690
rect 17875 -730 17880 -710
rect 17900 -730 17905 -710
rect 17875 -760 17905 -730
rect 17875 -780 17880 -760
rect 17900 -780 17905 -760
rect 17875 -810 17905 -780
rect 17875 -830 17880 -810
rect 17900 -830 17905 -810
rect 17875 -860 17905 -830
rect 17875 -880 17880 -860
rect 17900 -880 17905 -860
rect 17875 -910 17905 -880
rect 17875 -930 17880 -910
rect 17900 -930 17905 -910
rect 17875 -940 17905 -930
rect 18415 -710 18525 -700
rect 18415 -730 18420 -710
rect 18440 -730 18460 -710
rect 18480 -730 18500 -710
rect 18520 -730 18525 -710
rect 18415 -760 18525 -730
rect 18415 -780 18420 -760
rect 18440 -780 18460 -760
rect 18480 -780 18500 -760
rect 18520 -780 18525 -760
rect 18415 -810 18525 -780
rect 18415 -830 18420 -810
rect 18440 -830 18460 -810
rect 18480 -830 18500 -810
rect 18520 -830 18525 -810
rect 18415 -860 18525 -830
rect 18415 -880 18420 -860
rect 18440 -880 18460 -860
rect 18480 -880 18500 -860
rect 18520 -880 18525 -860
rect 18415 -910 18525 -880
rect 18415 -930 18420 -910
rect 18440 -930 18460 -910
rect 18480 -930 18500 -910
rect 18520 -930 18525 -910
rect 18415 -940 18525 -930
rect 19035 -710 19065 -700
rect 19035 -730 19040 -710
rect 19060 -730 19065 -710
rect 19035 -760 19065 -730
rect 19035 -780 19040 -760
rect 19060 -780 19065 -760
rect 19035 -810 19065 -780
rect 19035 -830 19040 -810
rect 19060 -830 19065 -810
rect 19035 -860 19065 -830
rect 19035 -880 19040 -860
rect 19060 -880 19065 -860
rect 19035 -910 19065 -880
rect 19035 -930 19040 -910
rect 19060 -930 19065 -910
rect 19035 -940 19065 -930
rect 17120 -960 17140 -940
rect 18460 -960 18480 -940
rect 17110 -970 17150 -960
rect 17110 -990 17120 -970
rect 17140 -990 17150 -970
rect 17110 -1000 17150 -990
rect 18450 -970 18490 -960
rect 18450 -990 18460 -970
rect 18480 -990 18490 -970
rect 18450 -1000 18490 -990
rect 16740 -1105 16780 -1095
rect 16740 -1125 16750 -1105
rect 16770 -1125 16780 -1105
rect 16740 -1135 16780 -1125
rect 16820 -1105 16860 -1095
rect 16820 -1125 16830 -1105
rect 16850 -1125 16860 -1105
rect 16820 -1135 16860 -1125
rect 16900 -1105 16940 -1095
rect 16900 -1125 16910 -1105
rect 16930 -1125 16940 -1105
rect 16900 -1135 16940 -1125
rect 16980 -1105 17020 -1095
rect 16980 -1125 16990 -1105
rect 17010 -1125 17020 -1105
rect 16980 -1135 17020 -1125
rect 17060 -1105 17100 -1095
rect 17060 -1125 17070 -1105
rect 17090 -1125 17100 -1105
rect 17060 -1135 17100 -1125
rect 17140 -1105 17180 -1095
rect 17140 -1125 17150 -1105
rect 17170 -1125 17180 -1105
rect 17140 -1135 17180 -1125
rect 17220 -1105 17260 -1095
rect 17220 -1125 17230 -1105
rect 17250 -1125 17260 -1105
rect 17220 -1135 17260 -1125
rect 17300 -1105 17340 -1095
rect 17300 -1125 17310 -1105
rect 17330 -1125 17340 -1105
rect 17300 -1135 17340 -1125
rect 17380 -1105 17420 -1095
rect 17380 -1125 17390 -1105
rect 17410 -1125 17420 -1105
rect 17380 -1135 17420 -1125
rect 17460 -1105 17500 -1095
rect 17460 -1125 17470 -1105
rect 17490 -1125 17500 -1105
rect 17460 -1135 17500 -1125
rect 17540 -1105 17580 -1095
rect 17540 -1125 17550 -1105
rect 17570 -1125 17580 -1105
rect 17540 -1135 17580 -1125
rect 17620 -1105 17660 -1095
rect 17620 -1125 17630 -1105
rect 17650 -1125 17660 -1105
rect 17620 -1135 17660 -1125
rect 17700 -1105 17740 -1095
rect 17700 -1125 17710 -1105
rect 17730 -1125 17740 -1105
rect 17700 -1135 17740 -1125
rect 17780 -1105 17820 -1095
rect 17780 -1125 17790 -1105
rect 17810 -1125 17820 -1105
rect 17780 -1135 17820 -1125
rect 17860 -1105 17900 -1095
rect 17860 -1125 17870 -1105
rect 17890 -1125 17900 -1105
rect 17860 -1135 17900 -1125
rect 17940 -1105 17980 -1095
rect 17940 -1125 17950 -1105
rect 17970 -1125 17980 -1105
rect 17940 -1135 17980 -1125
rect 18020 -1105 18060 -1095
rect 18020 -1125 18030 -1105
rect 18050 -1125 18060 -1105
rect 18020 -1135 18060 -1125
rect 18100 -1105 18140 -1095
rect 18100 -1125 18110 -1105
rect 18130 -1125 18140 -1105
rect 18100 -1135 18140 -1125
rect 18180 -1105 18220 -1095
rect 18180 -1125 18190 -1105
rect 18210 -1125 18220 -1105
rect 18180 -1135 18220 -1125
rect 18260 -1105 18300 -1095
rect 18260 -1125 18270 -1105
rect 18290 -1125 18300 -1105
rect 18260 -1135 18300 -1125
rect 18340 -1105 18380 -1095
rect 18340 -1125 18350 -1105
rect 18370 -1125 18380 -1105
rect 18340 -1135 18380 -1125
rect 18420 -1105 18460 -1095
rect 18420 -1125 18430 -1105
rect 18450 -1125 18460 -1105
rect 18420 -1135 18460 -1125
rect 18500 -1105 18540 -1095
rect 18500 -1125 18510 -1105
rect 18530 -1125 18540 -1105
rect 18500 -1135 18540 -1125
rect 18580 -1105 18620 -1095
rect 18580 -1125 18590 -1105
rect 18610 -1125 18620 -1105
rect 18580 -1135 18620 -1125
rect 18660 -1105 18700 -1095
rect 18660 -1125 18670 -1105
rect 18690 -1125 18700 -1105
rect 18660 -1135 18700 -1125
rect 18740 -1105 18780 -1095
rect 18740 -1125 18750 -1105
rect 18770 -1125 18780 -1105
rect 18740 -1135 18780 -1125
rect 16750 -1155 16770 -1135
rect 17790 -1155 17810 -1135
rect 16745 -1165 16775 -1155
rect 16745 -1180 16750 -1165
rect 16700 -1185 16750 -1180
rect 16770 -1185 16775 -1165
rect 16700 -1190 16775 -1185
rect 16700 -1210 16710 -1190
rect 16730 -1210 16775 -1190
rect 16700 -1215 16775 -1210
rect 16700 -1220 16750 -1215
rect 16745 -1235 16750 -1220
rect 16770 -1235 16775 -1215
rect 16745 -1245 16775 -1235
rect 17785 -1165 17815 -1155
rect 17785 -1185 17790 -1165
rect 17810 -1185 17815 -1165
rect 17785 -1215 17815 -1185
rect 17785 -1235 17790 -1215
rect 17810 -1235 17815 -1215
rect 17785 -1245 17815 -1235
rect 18825 -1160 18895 -1155
rect 18825 -1165 18935 -1160
rect 18825 -1185 18830 -1165
rect 18850 -1185 18870 -1165
rect 18890 -1170 18935 -1165
rect 18890 -1185 18905 -1170
rect 18825 -1190 18905 -1185
rect 18925 -1190 18935 -1170
rect 18825 -1210 18935 -1190
rect 18825 -1215 18905 -1210
rect 18825 -1235 18830 -1215
rect 18850 -1235 18870 -1215
rect 18890 -1230 18905 -1215
rect 18925 -1230 18935 -1210
rect 18890 -1235 18935 -1230
rect 18825 -1240 18935 -1235
rect 18825 -1245 18895 -1240
rect 16600 -1495 16640 -1485
rect 16600 -1515 16610 -1495
rect 16630 -1515 16640 -1495
rect 16600 -1525 16640 -1515
rect 16660 -1495 16690 -1485
rect 16660 -1515 16665 -1495
rect 16685 -1515 16690 -1495
rect 16660 -1525 16690 -1515
rect 16710 -1495 16750 -1485
rect 16710 -1515 16720 -1495
rect 16740 -1515 16750 -1495
rect 16710 -1525 16750 -1515
rect 16770 -1495 16800 -1485
rect 16770 -1515 16775 -1495
rect 16795 -1515 16800 -1495
rect 16770 -1525 16800 -1515
rect 16820 -1495 16860 -1485
rect 16820 -1515 16830 -1495
rect 16850 -1515 16860 -1495
rect 16820 -1525 16860 -1515
rect 16880 -1495 16920 -1485
rect 16880 -1515 16890 -1495
rect 16910 -1515 16920 -1495
rect 16880 -1525 16920 -1515
rect 17025 -1495 17065 -1485
rect 17025 -1515 17035 -1495
rect 17055 -1515 17065 -1495
rect 17025 -1525 17065 -1515
rect 17135 -1495 17175 -1485
rect 17135 -1515 17145 -1495
rect 17165 -1515 17175 -1495
rect 17135 -1525 17175 -1515
rect 17245 -1495 17285 -1485
rect 17245 -1515 17255 -1495
rect 17275 -1515 17285 -1495
rect 17245 -1525 17285 -1515
rect 17305 -1495 17335 -1485
rect 17305 -1515 17310 -1495
rect 17330 -1515 17335 -1495
rect 17305 -1525 17335 -1515
rect 17355 -1495 17395 -1485
rect 17355 -1515 17365 -1495
rect 17385 -1515 17395 -1495
rect 17355 -1525 17395 -1515
rect 17465 -1495 17505 -1485
rect 17465 -1515 17475 -1495
rect 17495 -1515 17505 -1495
rect 17465 -1525 17505 -1515
rect 17615 -1495 17655 -1485
rect 17615 -1515 17625 -1495
rect 17645 -1515 17655 -1495
rect 17615 -1525 17655 -1515
rect 17725 -1495 17765 -1485
rect 17725 -1515 17735 -1495
rect 17755 -1515 17765 -1495
rect 17725 -1525 17765 -1515
rect 17785 -1495 17815 -1485
rect 17785 -1515 17790 -1495
rect 17810 -1515 17815 -1495
rect 17785 -1525 17815 -1515
rect 17835 -1495 17875 -1485
rect 17835 -1515 17845 -1495
rect 17865 -1515 17875 -1495
rect 17835 -1525 17875 -1515
rect 17945 -1495 17985 -1485
rect 17945 -1515 17955 -1495
rect 17975 -1515 17985 -1495
rect 17945 -1525 17985 -1515
rect 18095 -1495 18135 -1485
rect 18095 -1515 18105 -1495
rect 18125 -1515 18135 -1495
rect 18095 -1525 18135 -1515
rect 18205 -1495 18245 -1485
rect 18205 -1515 18215 -1495
rect 18235 -1515 18245 -1495
rect 18205 -1525 18245 -1515
rect 18265 -1495 18295 -1485
rect 18265 -1515 18270 -1495
rect 18290 -1515 18295 -1495
rect 18265 -1525 18295 -1515
rect 18315 -1495 18355 -1485
rect 18315 -1515 18325 -1495
rect 18345 -1515 18355 -1495
rect 18315 -1525 18355 -1515
rect 18425 -1495 18465 -1485
rect 18425 -1515 18435 -1495
rect 18455 -1515 18465 -1495
rect 18425 -1525 18465 -1515
rect 18535 -1495 18575 -1485
rect 18535 -1515 18545 -1495
rect 18565 -1515 18575 -1495
rect 18535 -1525 18575 -1515
rect 16605 -1545 16635 -1525
rect 16665 -1545 16685 -1525
rect 16720 -1545 16740 -1525
rect 16830 -1545 16850 -1525
rect 16880 -1545 16910 -1525
rect 17030 -1545 17060 -1525
rect 17145 -1545 17165 -1525
rect 17255 -1545 17275 -1525
rect 17365 -1545 17385 -1525
rect 17470 -1545 17500 -1525
rect 17620 -1545 17650 -1525
rect 17735 -1545 17755 -1525
rect 17845 -1545 17865 -1525
rect 17950 -1545 17980 -1525
rect 18100 -1545 18130 -1525
rect 18215 -1545 18235 -1525
rect 18325 -1545 18345 -1525
rect 18435 -1545 18455 -1525
rect 18540 -1545 18570 -1525
rect 16565 -1555 16635 -1545
rect 16565 -1575 16570 -1555
rect 16590 -1575 16610 -1555
rect 16630 -1575 16635 -1555
rect 16565 -1605 16635 -1575
rect 16565 -1625 16570 -1605
rect 16590 -1625 16610 -1605
rect 16630 -1625 16635 -1605
rect 16565 -1635 16635 -1625
rect 16660 -1555 16690 -1545
rect 16660 -1575 16665 -1555
rect 16685 -1575 16690 -1555
rect 16660 -1605 16690 -1575
rect 16660 -1625 16665 -1605
rect 16685 -1625 16690 -1605
rect 16660 -1635 16690 -1625
rect 16715 -1555 16745 -1545
rect 16715 -1575 16720 -1555
rect 16740 -1575 16745 -1555
rect 16715 -1605 16745 -1575
rect 16715 -1625 16720 -1605
rect 16740 -1625 16745 -1605
rect 16715 -1635 16745 -1625
rect 16770 -1555 16800 -1545
rect 16770 -1575 16775 -1555
rect 16795 -1575 16800 -1555
rect 16770 -1605 16800 -1575
rect 16770 -1625 16775 -1605
rect 16795 -1625 16800 -1605
rect 16770 -1635 16800 -1625
rect 16825 -1555 16855 -1545
rect 16825 -1575 16830 -1555
rect 16850 -1575 16855 -1555
rect 16825 -1605 16855 -1575
rect 16825 -1625 16830 -1605
rect 16850 -1625 16855 -1605
rect 16825 -1635 16855 -1625
rect 16880 -1555 16950 -1545
rect 16880 -1575 16885 -1555
rect 16905 -1575 16925 -1555
rect 16945 -1575 16950 -1555
rect 16880 -1605 16950 -1575
rect 16880 -1625 16885 -1605
rect 16905 -1625 16925 -1605
rect 16945 -1625 16950 -1605
rect 16880 -1635 16950 -1625
rect 16990 -1555 17060 -1545
rect 16990 -1575 16995 -1555
rect 17015 -1575 17035 -1555
rect 17055 -1575 17060 -1555
rect 16990 -1605 17060 -1575
rect 16990 -1625 16995 -1605
rect 17015 -1625 17035 -1605
rect 17055 -1625 17060 -1605
rect 16990 -1635 17060 -1625
rect 17085 -1555 17115 -1545
rect 17085 -1575 17090 -1555
rect 17110 -1575 17115 -1555
rect 17085 -1605 17115 -1575
rect 17085 -1625 17090 -1605
rect 17110 -1625 17115 -1605
rect 17085 -1635 17115 -1625
rect 17140 -1555 17170 -1545
rect 17140 -1575 17145 -1555
rect 17165 -1575 17170 -1555
rect 17140 -1605 17170 -1575
rect 17140 -1625 17145 -1605
rect 17165 -1625 17170 -1605
rect 17140 -1635 17170 -1625
rect 17195 -1555 17225 -1545
rect 17195 -1575 17200 -1555
rect 17220 -1575 17225 -1555
rect 17195 -1605 17225 -1575
rect 17195 -1625 17200 -1605
rect 17220 -1625 17225 -1605
rect 17195 -1635 17225 -1625
rect 17250 -1555 17280 -1545
rect 17250 -1575 17255 -1555
rect 17275 -1575 17280 -1555
rect 17250 -1605 17280 -1575
rect 17250 -1625 17255 -1605
rect 17275 -1625 17280 -1605
rect 17250 -1635 17280 -1625
rect 17305 -1555 17335 -1545
rect 17305 -1575 17310 -1555
rect 17330 -1575 17335 -1555
rect 17305 -1605 17335 -1575
rect 17305 -1625 17310 -1605
rect 17330 -1625 17335 -1605
rect 17305 -1635 17335 -1625
rect 17360 -1555 17390 -1545
rect 17360 -1575 17365 -1555
rect 17385 -1575 17390 -1555
rect 17360 -1605 17390 -1575
rect 17360 -1625 17365 -1605
rect 17385 -1625 17390 -1605
rect 17360 -1635 17390 -1625
rect 17415 -1555 17445 -1545
rect 17415 -1575 17420 -1555
rect 17440 -1575 17445 -1555
rect 17415 -1605 17445 -1575
rect 17415 -1625 17420 -1605
rect 17440 -1625 17445 -1605
rect 17415 -1635 17445 -1625
rect 17470 -1555 17540 -1545
rect 17470 -1575 17475 -1555
rect 17495 -1575 17515 -1555
rect 17535 -1575 17540 -1555
rect 17470 -1605 17540 -1575
rect 17470 -1625 17475 -1605
rect 17495 -1625 17515 -1605
rect 17535 -1625 17540 -1605
rect 17470 -1635 17540 -1625
rect 17580 -1555 17650 -1545
rect 17580 -1575 17585 -1555
rect 17605 -1575 17625 -1555
rect 17645 -1575 17650 -1555
rect 17580 -1605 17650 -1575
rect 17580 -1625 17585 -1605
rect 17605 -1625 17625 -1605
rect 17645 -1625 17650 -1605
rect 17580 -1635 17650 -1625
rect 17675 -1555 17705 -1545
rect 17675 -1575 17680 -1555
rect 17700 -1575 17705 -1555
rect 17675 -1605 17705 -1575
rect 17675 -1625 17680 -1605
rect 17700 -1625 17705 -1605
rect 17675 -1635 17705 -1625
rect 17730 -1555 17760 -1545
rect 17730 -1575 17735 -1555
rect 17755 -1575 17760 -1555
rect 17730 -1605 17760 -1575
rect 17730 -1625 17735 -1605
rect 17755 -1625 17760 -1605
rect 17730 -1635 17760 -1625
rect 17785 -1555 17815 -1545
rect 17785 -1575 17790 -1555
rect 17810 -1575 17815 -1555
rect 17785 -1605 17815 -1575
rect 17785 -1625 17790 -1605
rect 17810 -1625 17815 -1605
rect 17785 -1635 17815 -1625
rect 17840 -1555 17870 -1545
rect 17840 -1575 17845 -1555
rect 17865 -1575 17870 -1555
rect 17840 -1605 17870 -1575
rect 17840 -1625 17845 -1605
rect 17865 -1625 17870 -1605
rect 17840 -1635 17870 -1625
rect 17895 -1555 17925 -1545
rect 17895 -1575 17900 -1555
rect 17920 -1575 17925 -1555
rect 17895 -1605 17925 -1575
rect 17895 -1625 17900 -1605
rect 17920 -1625 17925 -1605
rect 17895 -1635 17925 -1625
rect 17950 -1555 18020 -1545
rect 17950 -1575 17955 -1555
rect 17975 -1575 17995 -1555
rect 18015 -1575 18020 -1555
rect 17950 -1605 18020 -1575
rect 17950 -1625 17955 -1605
rect 17975 -1625 17995 -1605
rect 18015 -1625 18020 -1605
rect 17950 -1635 18020 -1625
rect 18060 -1555 18130 -1545
rect 18060 -1575 18065 -1555
rect 18085 -1575 18105 -1555
rect 18125 -1575 18130 -1555
rect 18060 -1605 18130 -1575
rect 18060 -1625 18065 -1605
rect 18085 -1625 18105 -1605
rect 18125 -1625 18130 -1605
rect 18060 -1635 18130 -1625
rect 18155 -1555 18185 -1545
rect 18155 -1575 18160 -1555
rect 18180 -1575 18185 -1555
rect 18155 -1605 18185 -1575
rect 18155 -1625 18160 -1605
rect 18180 -1625 18185 -1605
rect 18155 -1635 18185 -1625
rect 18210 -1555 18240 -1545
rect 18210 -1575 18215 -1555
rect 18235 -1575 18240 -1555
rect 18210 -1605 18240 -1575
rect 18210 -1625 18215 -1605
rect 18235 -1625 18240 -1605
rect 18210 -1635 18240 -1625
rect 18265 -1555 18295 -1545
rect 18265 -1575 18270 -1555
rect 18290 -1575 18295 -1555
rect 18265 -1605 18295 -1575
rect 18265 -1625 18270 -1605
rect 18290 -1625 18295 -1605
rect 18265 -1635 18295 -1625
rect 18320 -1555 18350 -1545
rect 18320 -1575 18325 -1555
rect 18345 -1575 18350 -1555
rect 18320 -1605 18350 -1575
rect 18320 -1625 18325 -1605
rect 18345 -1625 18350 -1605
rect 18320 -1635 18350 -1625
rect 18375 -1555 18405 -1545
rect 18375 -1575 18380 -1555
rect 18400 -1575 18405 -1555
rect 18375 -1605 18405 -1575
rect 18375 -1625 18380 -1605
rect 18400 -1625 18405 -1605
rect 18375 -1635 18405 -1625
rect 18430 -1555 18460 -1545
rect 18430 -1575 18435 -1555
rect 18455 -1575 18460 -1555
rect 18430 -1605 18460 -1575
rect 18430 -1625 18435 -1605
rect 18455 -1625 18460 -1605
rect 18430 -1635 18460 -1625
rect 18485 -1555 18515 -1545
rect 18485 -1575 18490 -1555
rect 18510 -1575 18515 -1555
rect 18485 -1605 18515 -1575
rect 18485 -1625 18490 -1605
rect 18510 -1625 18515 -1605
rect 18485 -1635 18515 -1625
rect 18540 -1555 18610 -1545
rect 18540 -1575 18545 -1555
rect 18565 -1575 18585 -1555
rect 18605 -1575 18610 -1555
rect 18540 -1605 18610 -1575
rect 18540 -1625 18545 -1605
rect 18565 -1625 18585 -1605
rect 18605 -1625 18610 -1605
rect 18540 -1635 18610 -1625
rect 16775 -1655 16795 -1635
rect 17090 -1655 17110 -1635
rect 17310 -1655 17330 -1635
rect 17680 -1655 17700 -1635
rect 17790 -1655 17810 -1635
rect 17900 -1655 17920 -1635
rect 18270 -1655 18290 -1635
rect 18490 -1655 18510 -1635
rect 16765 -1665 16805 -1655
rect 16765 -1685 16775 -1665
rect 16795 -1685 16805 -1665
rect 16765 -1695 16805 -1685
rect 17080 -1665 17120 -1655
rect 17080 -1685 17090 -1665
rect 17110 -1685 17120 -1665
rect 17080 -1695 17120 -1685
rect 17190 -1665 17230 -1655
rect 17190 -1685 17200 -1665
rect 17220 -1685 17230 -1665
rect 17190 -1695 17230 -1685
rect 17300 -1665 17340 -1655
rect 17300 -1685 17310 -1665
rect 17330 -1685 17340 -1665
rect 17300 -1695 17340 -1685
rect 17410 -1665 17450 -1655
rect 17410 -1685 17420 -1665
rect 17440 -1685 17450 -1665
rect 17410 -1695 17450 -1685
rect 17670 -1665 17710 -1655
rect 17670 -1685 17680 -1665
rect 17700 -1685 17710 -1665
rect 17670 -1695 17710 -1685
rect 17780 -1665 17820 -1655
rect 17780 -1685 17790 -1665
rect 17810 -1685 17820 -1665
rect 17780 -1695 17820 -1685
rect 17890 -1665 17930 -1655
rect 17890 -1685 17900 -1665
rect 17920 -1685 17930 -1665
rect 17890 -1695 17930 -1685
rect 18150 -1665 18190 -1655
rect 18150 -1685 18160 -1665
rect 18180 -1685 18190 -1665
rect 18150 -1695 18190 -1685
rect 18260 -1665 18300 -1655
rect 18260 -1685 18270 -1665
rect 18290 -1685 18300 -1665
rect 18260 -1695 18300 -1685
rect 18370 -1665 18410 -1655
rect 18370 -1685 18380 -1665
rect 18400 -1685 18410 -1665
rect 18370 -1695 18410 -1685
rect 18480 -1665 18520 -1655
rect 18480 -1685 18490 -1665
rect 18510 -1685 18520 -1665
rect 18480 -1695 18520 -1685
rect 17425 -2005 17470 -2000
rect 17425 -2030 17435 -2005
rect 17460 -2030 17470 -2005
rect 17425 -2035 17470 -2030
rect 18124 -2005 18169 -2000
rect 18124 -2030 18134 -2005
rect 18159 -2030 18169 -2005
rect 18124 -2035 18169 -2030
rect 16795 -2240 18805 -2115
rect 17440 -2795 17480 -2240
rect 18120 -2795 18160 -2240
rect 16485 -2905 16520 -2895
rect 16485 -2930 16490 -2905
rect 16515 -2930 16520 -2905
rect 16795 -2920 18805 -2795
rect 19080 -2905 19115 -2895
rect 16485 -2940 16520 -2930
rect 16160 -3030 16195 -3020
rect 16160 -3055 16165 -3030
rect 16190 -3055 16195 -3030
rect 16160 -3065 16195 -3055
rect 15950 -3121 15985 -3110
rect 15950 -3146 15955 -3121
rect 15980 -3146 15985 -3121
rect 15950 -3156 15985 -3146
rect 16255 -3100 16280 -3065
rect 16580 -2975 16605 -2940
rect 17440 -3475 17480 -2920
rect 18120 -3475 18160 -2920
rect 19080 -2930 19085 -2905
rect 19110 -2930 19115 -2905
rect 19080 -2940 19115 -2930
rect 18995 -2975 19020 -2940
rect 19405 -3002 19440 -2992
rect 19405 -3027 19410 -3002
rect 19435 -3027 19440 -3002
rect 19405 -3037 19440 -3027
rect 19320 -3072 19345 -3037
rect 19610 -3120 19645 -3110
rect 19610 -3145 19615 -3120
rect 19640 -3145 19645 -3120
rect 19610 -3156 19645 -3145
rect 16795 -3600 18805 -3475
rect 15950 -3794 15985 -3784
rect 15950 -3819 15955 -3794
rect 15980 -3819 15985 -3794
rect 15950 -3829 15985 -3819
rect 16195 -3889 16220 -3854
rect 16280 -3899 16315 -3889
rect 16280 -3924 16285 -3899
rect 16310 -3924 16315 -3899
rect 16280 -3934 16315 -3924
rect 16520 -3964 16545 -3929
rect 16605 -3974 16640 -3964
rect 16605 -3999 16610 -3974
rect 16635 -3999 16640 -3974
rect 16605 -4009 16640 -3999
rect 17440 -4125 17480 -3600
rect 17780 -4170 17820 -4120
rect 18120 -4125 18160 -3600
rect 19055 -3964 19080 -3929
rect 19380 -3889 19405 -3854
rect 19610 -3794 19645 -3784
rect 19610 -3819 19615 -3794
rect 19640 -3819 19645 -3794
rect 19610 -3829 19645 -3819
rect 19285 -3899 19320 -3889
rect 19285 -3924 19290 -3899
rect 19315 -3924 19320 -3899
rect 19285 -3934 19320 -3924
rect 18960 -3974 18995 -3964
rect 18960 -3999 18965 -3974
rect 18990 -3999 18995 -3974
rect 18960 -4009 18995 -3999
rect 17780 -4190 17790 -4170
rect 17810 -4190 17820 -4170
rect 17780 -4220 17820 -4190
rect 17780 -4240 17790 -4220
rect 17810 -4240 17820 -4220
rect 17780 -4270 17820 -4240
rect 17780 -4290 17790 -4270
rect 17810 -4290 17820 -4270
rect 17780 -4300 17820 -4290
<< viali >>
rect 16495 1590 16515 1610
rect 17790 1590 17810 1610
rect 16375 1455 16395 1475
rect 16495 1455 16515 1475
rect 16615 1455 16635 1475
rect 16895 1455 16915 1475
rect 16950 1455 16970 1475
rect 17005 1455 17025 1475
rect 17060 1455 17080 1475
rect 17115 1455 17135 1475
rect 17225 1455 17245 1475
rect 17505 1455 17525 1475
rect 17570 1455 17590 1475
rect 17625 1455 17645 1475
rect 17680 1455 17700 1475
rect 17735 1455 17755 1475
rect 17790 1455 17810 1475
rect 17845 1455 17865 1475
rect 17900 1455 17920 1475
rect 17955 1455 17975 1475
rect 18010 1455 18030 1475
rect 18075 1455 18095 1475
rect 18355 1455 18375 1475
rect 18465 1455 18485 1475
rect 18520 1455 18540 1475
rect 18575 1455 18595 1475
rect 18630 1455 18650 1475
rect 18685 1455 18705 1475
rect 16440 1285 16460 1305
rect 16550 1285 16570 1305
rect 16950 1285 16970 1305
rect 17060 1285 17080 1305
rect 17170 1285 17190 1305
rect 17625 1285 17645 1305
rect 17735 1285 17755 1305
rect 17845 1285 17865 1305
rect 17955 1285 17975 1305
rect 18410 1285 18430 1305
rect 18520 1285 18540 1305
rect 18630 1285 18650 1305
rect 16980 990 17000 1010
rect 17160 990 17180 1010
rect 17340 990 17360 1010
rect 17520 990 17540 1010
rect 17700 990 17720 1010
rect 17880 990 17900 1010
rect 18060 990 18080 1010
rect 18240 990 18260 1010
rect 18420 990 18440 1010
rect 18600 990 18620 1010
rect 18915 990 18935 1010
rect 19025 990 19045 1010
rect 19085 990 19105 1010
rect 16445 890 16465 910
rect 16555 890 16575 910
rect 16665 890 16685 910
rect 16490 720 16510 740
rect 16555 720 16575 740
rect 16620 720 16640 740
rect 18960 720 18980 740
rect 19010 660 19030 680
rect 17070 620 17090 640
rect 17250 620 17270 640
rect 17430 620 17450 640
rect 17610 620 17630 640
rect 17700 620 17720 640
rect 17790 620 17810 640
rect 17970 620 17990 640
rect 18150 620 18170 640
rect 18330 620 18350 640
rect 18510 620 18530 640
rect 16430 150 16450 170
rect 16490 150 16510 170
rect 16550 150 16570 170
rect 16670 150 16690 170
rect 16790 150 16810 170
rect 16850 150 16870 170
rect 16910 150 16930 170
rect 17030 150 17050 170
rect 17150 150 17170 170
rect 17210 150 17230 170
rect 17270 150 17290 170
rect 17390 150 17410 170
rect 17510 150 17530 170
rect 17570 150 17590 170
rect 17630 150 17650 170
rect 17950 150 17970 170
rect 18010 150 18030 170
rect 18070 150 18090 170
rect 18190 150 18210 170
rect 18310 150 18330 170
rect 18370 150 18390 170
rect 18430 150 18450 170
rect 18550 150 18570 170
rect 18670 150 18690 170
rect 18730 150 18750 170
rect 18790 150 18810 170
rect 18910 150 18930 170
rect 19030 150 19050 170
rect 19090 150 19110 170
rect 19150 150 19170 170
rect 16520 -20 16540 0
rect 16610 -20 16630 0
rect 16730 -20 16750 0
rect 16850 -20 16870 0
rect 16970 -20 16990 0
rect 17090 -20 17110 0
rect 17210 -20 17230 0
rect 17330 -20 17350 0
rect 17450 -20 17470 0
rect 17540 -20 17560 0
rect 18040 -20 18060 0
rect 18130 -20 18150 0
rect 18250 -20 18270 0
rect 18370 -20 18390 0
rect 18490 -20 18510 0
rect 18610 -20 18630 0
rect 18730 -20 18750 0
rect 18850 -20 18870 0
rect 18970 -20 18990 0
rect 19060 -20 19080 0
rect 16965 -135 16985 -115
rect 17012 -135 17032 -115
rect 17095 -135 17115 -115
rect 18485 -135 18505 -115
rect 18568 -135 18588 -115
rect 18615 -135 18635 -115
rect 17030 -195 17050 -175
rect 17030 -245 17050 -225
rect 17030 -295 17050 -275
rect 17030 -345 17050 -325
rect 17030 -395 17050 -375
rect 17570 -195 17590 -175
rect 17570 -235 17590 -215
rect 17570 -275 17590 -255
rect 18010 -195 18030 -175
rect 18010 -235 18030 -215
rect 18010 -275 18030 -255
rect 17080 -455 17100 -435
rect 18500 -455 18520 -435
rect 18550 -455 18570 -435
rect 16630 -670 16650 -650
rect 16750 -670 16770 -650
rect 16870 -670 16890 -650
rect 16990 -670 17010 -650
rect 17310 -670 17330 -650
rect 17430 -670 17450 -650
rect 17550 -670 17570 -650
rect 17700 -685 17720 -665
rect 16540 -730 16560 -710
rect 16540 -780 16560 -760
rect 16540 -830 16560 -810
rect 16540 -880 16560 -860
rect 16540 -930 16560 -910
rect 17880 -685 17900 -665
rect 18030 -670 18050 -650
rect 18150 -670 18170 -650
rect 18270 -670 18290 -650
rect 18590 -670 18610 -650
rect 18710 -670 18730 -650
rect 18830 -670 18850 -650
rect 18950 -670 18970 -650
rect 19040 -690 19060 -670
rect 17120 -990 17140 -970
rect 18460 -990 18480 -970
rect 16750 -1125 16770 -1105
rect 16830 -1125 16850 -1105
rect 16910 -1125 16930 -1105
rect 16990 -1125 17010 -1105
rect 17070 -1125 17090 -1105
rect 17150 -1125 17170 -1105
rect 17230 -1125 17250 -1105
rect 17310 -1125 17330 -1105
rect 17390 -1125 17410 -1105
rect 17470 -1125 17490 -1105
rect 17550 -1125 17570 -1105
rect 17630 -1125 17650 -1105
rect 17710 -1125 17730 -1105
rect 17790 -1125 17810 -1105
rect 17870 -1125 17890 -1105
rect 17950 -1125 17970 -1105
rect 18030 -1125 18050 -1105
rect 18110 -1125 18130 -1105
rect 18190 -1125 18210 -1105
rect 18270 -1125 18290 -1105
rect 18350 -1125 18370 -1105
rect 18430 -1125 18450 -1105
rect 18510 -1125 18530 -1105
rect 18590 -1125 18610 -1105
rect 18670 -1125 18690 -1105
rect 18750 -1125 18770 -1105
rect 16710 -1210 16730 -1190
rect 18905 -1190 18925 -1170
rect 18905 -1230 18925 -1210
rect 16610 -1515 16630 -1495
rect 16665 -1515 16685 -1495
rect 16720 -1515 16740 -1495
rect 16775 -1515 16795 -1495
rect 16830 -1515 16850 -1495
rect 16890 -1515 16910 -1495
rect 17035 -1515 17055 -1495
rect 17145 -1515 17165 -1495
rect 17255 -1515 17275 -1495
rect 17310 -1515 17330 -1495
rect 17365 -1515 17385 -1495
rect 17475 -1515 17495 -1495
rect 17625 -1515 17645 -1495
rect 17735 -1515 17755 -1495
rect 17790 -1515 17810 -1495
rect 17845 -1515 17865 -1495
rect 17955 -1515 17975 -1495
rect 18105 -1515 18125 -1495
rect 18215 -1515 18235 -1495
rect 18270 -1515 18290 -1495
rect 18325 -1515 18345 -1495
rect 18435 -1515 18455 -1495
rect 18545 -1515 18565 -1495
rect 17200 -1575 17220 -1555
rect 17200 -1625 17220 -1605
rect 17420 -1575 17440 -1555
rect 17420 -1625 17440 -1605
rect 18160 -1575 18180 -1555
rect 18160 -1625 18180 -1605
rect 18380 -1575 18400 -1555
rect 18380 -1625 18400 -1605
rect 16775 -1685 16795 -1665
rect 17090 -1685 17110 -1665
rect 17200 -1685 17220 -1665
rect 17310 -1685 17330 -1665
rect 17420 -1685 17440 -1665
rect 17680 -1685 17700 -1665
rect 17790 -1685 17810 -1665
rect 17900 -1685 17920 -1665
rect 18160 -1685 18180 -1665
rect 18270 -1685 18290 -1665
rect 18380 -1685 18400 -1665
rect 18490 -1685 18510 -1665
rect 17435 -2030 17460 -2005
rect 18134 -2030 18159 -2005
rect 16490 -2930 16515 -2905
rect 16165 -3055 16190 -3030
rect 15955 -3146 15980 -3121
rect 19085 -2930 19110 -2905
rect 19410 -3027 19435 -3002
rect 19615 -3145 19640 -3120
rect 15955 -3819 15980 -3794
rect 16285 -3924 16310 -3899
rect 16610 -3999 16635 -3974
rect 19615 -3819 19640 -3794
rect 19290 -3924 19315 -3899
rect 18965 -3999 18990 -3974
rect 17790 -4290 17810 -4270
<< metal1 >>
rect 15725 -55 15765 -50
rect 15725 -85 15730 -55
rect 15760 -85 15765 -55
rect 15725 -90 15765 -85
rect 15735 -4310 15755 -90
rect 15790 -1765 15815 1795
rect 15890 1310 15930 1315
rect 15890 1280 15895 1310
rect 15925 1280 15930 1310
rect 15890 -1355 15930 1280
rect 15945 175 15985 180
rect 15945 145 15950 175
rect 15980 145 15985 175
rect 15945 140 15985 145
rect 15890 -1385 15895 -1355
rect 15925 -1385 15930 -1355
rect 15890 -1390 15930 -1385
rect 15785 -1770 15825 -1765
rect 15785 -1800 15790 -1770
rect 15820 -1800 15825 -1770
rect 15785 -1805 15825 -1800
rect 15955 -3110 15975 140
rect 16040 -1710 16060 1795
rect 16030 -1715 16070 -1710
rect 16030 -1745 16035 -1715
rect 16065 -1745 16070 -1715
rect 16030 -1750 16070 -1745
rect 16115 -1860 16135 1795
rect 16485 1615 16525 1620
rect 16485 1585 16490 1615
rect 16520 1585 16525 1615
rect 16485 1580 16525 1585
rect 16365 1560 16405 1565
rect 16365 1530 16370 1560
rect 16400 1530 16405 1560
rect 16365 1520 16405 1530
rect 16365 1490 16370 1520
rect 16400 1490 16405 1520
rect 16365 1480 16405 1490
rect 16365 1450 16370 1480
rect 16400 1450 16405 1480
rect 16365 1445 16405 1450
rect 16485 1560 16525 1565
rect 16485 1530 16490 1560
rect 16520 1530 16525 1560
rect 16485 1520 16525 1530
rect 16485 1490 16490 1520
rect 16520 1490 16525 1520
rect 16485 1480 16525 1490
rect 16485 1450 16490 1480
rect 16520 1450 16525 1480
rect 16485 1445 16525 1450
rect 16605 1560 16645 1565
rect 16605 1530 16610 1560
rect 16640 1530 16645 1560
rect 16605 1520 16645 1530
rect 16605 1490 16610 1520
rect 16640 1490 16645 1520
rect 16605 1480 16645 1490
rect 16605 1450 16610 1480
rect 16640 1450 16645 1480
rect 16605 1445 16645 1450
rect 16885 1560 16925 1565
rect 16885 1530 16890 1560
rect 16920 1530 16925 1560
rect 16885 1520 16925 1530
rect 16885 1490 16890 1520
rect 16920 1490 16925 1520
rect 16885 1480 16925 1490
rect 16950 1485 16970 1795
rect 17050 1615 17090 1620
rect 17050 1585 17055 1615
rect 17085 1585 17090 1615
rect 17050 1580 17090 1585
rect 16995 1560 17035 1565
rect 16995 1530 17000 1560
rect 17030 1530 17035 1560
rect 16995 1520 17035 1530
rect 16995 1490 17000 1520
rect 17030 1490 17035 1520
rect 16885 1450 16890 1480
rect 16920 1450 16925 1480
rect 16885 1445 16925 1450
rect 16945 1475 16975 1485
rect 16945 1455 16950 1475
rect 16970 1455 16975 1475
rect 16945 1445 16975 1455
rect 16995 1480 17035 1490
rect 16995 1450 17000 1480
rect 17030 1450 17035 1480
rect 16995 1445 17035 1450
rect 17055 1475 17085 1580
rect 17055 1455 17060 1475
rect 17080 1455 17085 1475
rect 17055 1445 17085 1455
rect 17105 1560 17145 1565
rect 17105 1530 17110 1560
rect 17140 1530 17145 1560
rect 17105 1520 17145 1530
rect 17105 1490 17110 1520
rect 17140 1490 17145 1520
rect 17105 1480 17145 1490
rect 17105 1450 17110 1480
rect 17140 1450 17145 1480
rect 17105 1445 17145 1450
rect 17215 1560 17255 1565
rect 17215 1530 17220 1560
rect 17250 1530 17255 1560
rect 17215 1520 17255 1530
rect 17215 1490 17220 1520
rect 17250 1490 17255 1520
rect 17215 1480 17255 1490
rect 17215 1450 17220 1480
rect 17250 1450 17255 1480
rect 17215 1445 17255 1450
rect 17495 1560 17535 1565
rect 17495 1530 17500 1560
rect 17530 1530 17535 1560
rect 17495 1520 17535 1530
rect 17495 1490 17500 1520
rect 17530 1490 17535 1520
rect 17495 1480 17535 1490
rect 17495 1450 17500 1480
rect 17530 1450 17535 1480
rect 17495 1445 17535 1450
rect 17560 1560 17600 1565
rect 17560 1530 17565 1560
rect 17595 1530 17600 1560
rect 17560 1520 17600 1530
rect 17560 1490 17565 1520
rect 17595 1490 17600 1520
rect 17560 1480 17600 1490
rect 17560 1450 17565 1480
rect 17595 1450 17600 1480
rect 17560 1445 17600 1450
rect 17620 1475 17650 1795
rect 17620 1455 17625 1475
rect 17645 1455 17650 1475
rect 17620 1445 17650 1455
rect 17670 1560 17710 1565
rect 17670 1530 17675 1560
rect 17705 1530 17710 1560
rect 17670 1520 17710 1530
rect 17670 1490 17675 1520
rect 17705 1490 17710 1520
rect 17670 1480 17710 1490
rect 17670 1450 17675 1480
rect 17705 1450 17710 1480
rect 17670 1445 17710 1450
rect 17730 1475 17760 1795
rect 17780 1615 17820 1620
rect 17780 1585 17785 1615
rect 17815 1585 17820 1615
rect 17780 1580 17820 1585
rect 17730 1455 17735 1475
rect 17755 1455 17760 1475
rect 17730 1445 17760 1455
rect 17780 1560 17820 1565
rect 17780 1530 17785 1560
rect 17815 1530 17820 1560
rect 17780 1520 17820 1530
rect 17780 1490 17785 1520
rect 17815 1490 17820 1520
rect 17780 1480 17820 1490
rect 17780 1450 17785 1480
rect 17815 1450 17820 1480
rect 17780 1445 17820 1450
rect 17840 1475 17870 1795
rect 17840 1455 17845 1475
rect 17865 1455 17870 1475
rect 17840 1445 17870 1455
rect 17890 1560 17930 1565
rect 17890 1530 17895 1560
rect 17925 1530 17930 1560
rect 17890 1520 17930 1530
rect 17890 1490 17895 1520
rect 17925 1490 17930 1520
rect 17890 1480 17930 1490
rect 17890 1450 17895 1480
rect 17925 1450 17930 1480
rect 17890 1445 17930 1450
rect 17950 1475 17980 1795
rect 18510 1585 18515 1615
rect 18545 1585 18550 1615
rect 18510 1580 18550 1585
rect 17950 1455 17955 1475
rect 17975 1455 17980 1475
rect 17950 1445 17980 1455
rect 18000 1560 18040 1565
rect 18000 1530 18005 1560
rect 18035 1530 18040 1560
rect 18000 1520 18040 1530
rect 18000 1490 18005 1520
rect 18035 1490 18040 1520
rect 18000 1480 18040 1490
rect 18000 1450 18005 1480
rect 18035 1450 18040 1480
rect 18000 1445 18040 1450
rect 18065 1560 18105 1565
rect 18065 1530 18070 1560
rect 18100 1530 18105 1560
rect 18065 1520 18105 1530
rect 18065 1490 18070 1520
rect 18100 1490 18105 1520
rect 18065 1480 18105 1490
rect 18065 1450 18070 1480
rect 18100 1450 18105 1480
rect 18065 1445 18105 1450
rect 18345 1560 18385 1565
rect 18345 1530 18350 1560
rect 18380 1530 18385 1560
rect 18345 1520 18385 1530
rect 18345 1490 18350 1520
rect 18380 1490 18385 1520
rect 18345 1480 18385 1490
rect 18345 1450 18350 1480
rect 18380 1450 18385 1480
rect 18345 1445 18385 1450
rect 18455 1560 18495 1565
rect 18455 1530 18460 1560
rect 18490 1530 18495 1560
rect 18455 1520 18495 1530
rect 18455 1490 18460 1520
rect 18490 1490 18495 1520
rect 18455 1480 18495 1490
rect 18520 1485 18540 1580
rect 18565 1560 18605 1565
rect 18565 1530 18570 1560
rect 18600 1530 18605 1560
rect 18565 1520 18605 1530
rect 18565 1490 18570 1520
rect 18600 1490 18605 1520
rect 18455 1450 18460 1480
rect 18490 1450 18495 1480
rect 18455 1445 18495 1450
rect 18515 1475 18545 1485
rect 18515 1455 18520 1475
rect 18540 1455 18545 1475
rect 18515 1445 18545 1455
rect 18565 1480 18605 1490
rect 18630 1485 18650 1795
rect 18675 1560 18715 1565
rect 18675 1530 18680 1560
rect 18710 1530 18715 1560
rect 18675 1520 18715 1530
rect 18675 1490 18680 1520
rect 18710 1490 18715 1520
rect 18565 1450 18570 1480
rect 18600 1450 18605 1480
rect 18565 1445 18605 1450
rect 18625 1475 18655 1485
rect 18625 1455 18630 1475
rect 18650 1455 18655 1475
rect 18625 1445 18655 1455
rect 18675 1480 18715 1490
rect 18675 1450 18680 1480
rect 18710 1450 18715 1480
rect 18675 1445 18715 1450
rect 16430 1310 16470 1315
rect 16430 1280 16435 1310
rect 16465 1280 16470 1310
rect 16430 1275 16470 1280
rect 16540 1310 16580 1315
rect 16540 1280 16545 1310
rect 16575 1280 16580 1310
rect 16540 1275 16580 1280
rect 16940 1310 16980 1315
rect 16940 1280 16945 1310
rect 16975 1280 16980 1310
rect 16940 1275 16980 1280
rect 17050 1310 17090 1315
rect 17050 1280 17055 1310
rect 17085 1280 17090 1310
rect 17050 1275 17090 1280
rect 17160 1310 17200 1315
rect 17160 1280 17165 1310
rect 17195 1280 17200 1310
rect 17160 1275 17200 1280
rect 17615 1310 17655 1315
rect 17615 1280 17620 1310
rect 17650 1280 17655 1310
rect 17615 1275 17655 1280
rect 17725 1310 17765 1315
rect 17725 1280 17730 1310
rect 17760 1280 17765 1310
rect 17725 1275 17765 1280
rect 17835 1310 17875 1315
rect 17835 1280 17840 1310
rect 17870 1280 17875 1310
rect 17835 1275 17875 1280
rect 17945 1310 17985 1315
rect 17945 1280 17950 1310
rect 17980 1280 17985 1310
rect 17945 1275 17985 1280
rect 18400 1310 18440 1315
rect 18400 1280 18405 1310
rect 18435 1280 18440 1310
rect 18400 1275 18440 1280
rect 18510 1310 18550 1315
rect 18510 1280 18515 1310
rect 18545 1280 18550 1310
rect 18510 1275 18550 1280
rect 18620 1310 18660 1315
rect 18620 1280 18625 1310
rect 18655 1280 18660 1310
rect 18620 1275 18660 1280
rect 16550 1215 16570 1275
rect 16540 1210 16580 1215
rect 16540 1180 16545 1210
rect 16575 1180 16580 1210
rect 16540 1175 16580 1180
rect 16435 1095 16475 1100
rect 16435 1065 16440 1095
rect 16470 1065 16475 1095
rect 16435 1055 16475 1065
rect 16435 1025 16440 1055
rect 16470 1025 16475 1055
rect 16435 1015 16475 1025
rect 16435 985 16440 1015
rect 16470 985 16475 1015
rect 16435 980 16475 985
rect 16655 1095 16695 1100
rect 16655 1065 16660 1095
rect 16690 1065 16695 1095
rect 16655 1055 16695 1065
rect 16655 1025 16660 1055
rect 16690 1025 16695 1055
rect 16655 1015 16695 1025
rect 16655 985 16660 1015
rect 16690 985 16695 1015
rect 16655 980 16695 985
rect 16970 1095 17010 1100
rect 16970 1065 16975 1095
rect 17005 1065 17010 1095
rect 16970 1055 17010 1065
rect 16970 1025 16975 1055
rect 17005 1025 17010 1055
rect 16970 1015 17010 1025
rect 16970 985 16975 1015
rect 17005 985 17010 1015
rect 16970 980 17010 985
rect 17150 1095 17190 1100
rect 17150 1065 17155 1095
rect 17185 1065 17190 1095
rect 17150 1055 17190 1065
rect 17150 1025 17155 1055
rect 17185 1025 17190 1055
rect 17150 1015 17190 1025
rect 17150 985 17155 1015
rect 17185 985 17190 1015
rect 17150 980 17190 985
rect 17330 1095 17370 1100
rect 17330 1065 17335 1095
rect 17365 1065 17370 1095
rect 17330 1055 17370 1065
rect 17330 1025 17335 1055
rect 17365 1025 17370 1055
rect 17330 1015 17370 1025
rect 17330 985 17335 1015
rect 17365 985 17370 1015
rect 17330 980 17370 985
rect 17510 1095 17550 1100
rect 17510 1065 17515 1095
rect 17545 1065 17550 1095
rect 17510 1055 17550 1065
rect 17510 1025 17515 1055
rect 17545 1025 17550 1055
rect 17510 1015 17550 1025
rect 17510 985 17515 1015
rect 17545 985 17550 1015
rect 17510 980 17550 985
rect 17690 1095 17730 1100
rect 17690 1065 17695 1095
rect 17725 1065 17730 1095
rect 17690 1055 17730 1065
rect 17690 1025 17695 1055
rect 17725 1025 17730 1055
rect 17690 1015 17730 1025
rect 17690 985 17695 1015
rect 17725 985 17730 1015
rect 17690 980 17730 985
rect 17870 1095 17910 1100
rect 17870 1065 17875 1095
rect 17905 1065 17910 1095
rect 17870 1055 17910 1065
rect 17870 1025 17875 1055
rect 17905 1025 17910 1055
rect 17870 1015 17910 1025
rect 17870 985 17875 1015
rect 17905 985 17910 1015
rect 17870 980 17910 985
rect 18050 1095 18090 1100
rect 18050 1065 18055 1095
rect 18085 1065 18090 1095
rect 18050 1055 18090 1065
rect 18050 1025 18055 1055
rect 18085 1025 18090 1055
rect 18050 1015 18090 1025
rect 18050 985 18055 1015
rect 18085 985 18090 1015
rect 18050 980 18090 985
rect 18230 1095 18270 1100
rect 18230 1065 18235 1095
rect 18265 1065 18270 1095
rect 18230 1055 18270 1065
rect 18230 1025 18235 1055
rect 18265 1025 18270 1055
rect 18230 1015 18270 1025
rect 18230 985 18235 1015
rect 18265 985 18270 1015
rect 18230 980 18270 985
rect 18410 1095 18450 1100
rect 18410 1065 18415 1095
rect 18445 1065 18450 1095
rect 18410 1055 18450 1065
rect 18410 1025 18415 1055
rect 18445 1025 18450 1055
rect 18410 1015 18450 1025
rect 18410 985 18415 1015
rect 18445 985 18450 1015
rect 18410 980 18450 985
rect 18590 1095 18630 1100
rect 18590 1065 18595 1095
rect 18625 1065 18630 1095
rect 18590 1055 18630 1065
rect 18590 1025 18595 1055
rect 18625 1025 18630 1055
rect 18590 1015 18630 1025
rect 18590 985 18595 1015
rect 18625 985 18630 1015
rect 18590 980 18630 985
rect 18905 1095 18945 1100
rect 18905 1065 18910 1095
rect 18940 1065 18945 1095
rect 18905 1055 18945 1065
rect 18905 1025 18910 1055
rect 18940 1025 18945 1055
rect 18905 1015 18945 1025
rect 18905 985 18910 1015
rect 18940 985 18945 1015
rect 18905 980 18945 985
rect 19015 1095 19055 1100
rect 19015 1065 19020 1095
rect 19050 1065 19055 1095
rect 19015 1055 19055 1065
rect 19015 1025 19020 1055
rect 19050 1025 19055 1055
rect 19015 1015 19055 1025
rect 19015 985 19020 1015
rect 19050 985 19055 1015
rect 19015 980 19055 985
rect 19075 1095 19115 1100
rect 19075 1065 19080 1095
rect 19110 1065 19115 1095
rect 19075 1055 19115 1065
rect 19075 1025 19080 1055
rect 19110 1025 19115 1055
rect 19075 1015 19115 1025
rect 19075 985 19080 1015
rect 19110 985 19115 1015
rect 19075 980 19115 985
rect 16445 920 16465 980
rect 16665 920 16685 980
rect 16435 910 16475 920
rect 16435 890 16445 910
rect 16465 890 16475 910
rect 16435 880 16475 890
rect 16545 915 16585 920
rect 16545 885 16550 915
rect 16580 885 16585 915
rect 16545 880 16585 885
rect 16655 910 16695 920
rect 16655 890 16665 910
rect 16685 890 16695 910
rect 16655 880 16695 890
rect 16780 915 16820 920
rect 16780 885 16785 915
rect 16815 885 16820 915
rect 16780 880 16820 885
rect 16480 745 16520 750
rect 16480 715 16485 745
rect 16515 715 16520 745
rect 16480 710 16520 715
rect 16545 740 16585 750
rect 16545 720 16555 740
rect 16575 720 16585 740
rect 16545 710 16585 720
rect 16610 745 16650 750
rect 16610 715 16615 745
rect 16645 715 16650 745
rect 16610 710 16650 715
rect 16315 645 16355 650
rect 16315 615 16320 645
rect 16350 615 16355 645
rect 16260 590 16300 595
rect 16260 560 16265 590
rect 16295 560 16300 590
rect 16205 535 16245 540
rect 16205 505 16210 535
rect 16240 505 16245 535
rect 16205 500 16245 505
rect 16215 -1180 16235 500
rect 16260 -110 16300 560
rect 16260 -140 16265 -110
rect 16295 -140 16300 -110
rect 16205 -1185 16245 -1180
rect 16205 -1215 16210 -1185
rect 16240 -1215 16245 -1185
rect 16205 -1220 16245 -1215
rect 16105 -1865 16145 -1860
rect 16105 -1895 16110 -1865
rect 16140 -1895 16145 -1865
rect 16105 -1900 16145 -1895
rect 16155 -1950 16195 -1945
rect 16155 -1980 16160 -1950
rect 16190 -1980 16195 -1950
rect 16155 -1985 16195 -1980
rect 16165 -3020 16185 -1985
rect 16260 -2100 16300 -140
rect 16315 -430 16355 615
rect 16420 390 16460 395
rect 16420 360 16425 390
rect 16455 360 16460 390
rect 16420 350 16460 360
rect 16420 320 16425 350
rect 16455 320 16460 350
rect 16420 310 16460 320
rect 16420 280 16425 310
rect 16455 280 16460 310
rect 16420 275 16460 280
rect 16430 180 16450 275
rect 16490 180 16510 710
rect 16555 540 16575 710
rect 16790 595 16810 880
rect 19270 750 19290 1795
rect 19325 1210 19365 1215
rect 19325 1180 19330 1210
rect 19360 1180 19365 1210
rect 19325 1175 19365 1180
rect 18950 745 18990 750
rect 18950 715 18955 745
rect 18985 715 18990 745
rect 18950 710 18990 715
rect 19260 745 19300 750
rect 19260 715 19265 745
rect 19295 715 19300 745
rect 19260 710 19300 715
rect 19000 685 19040 690
rect 19000 655 19005 685
rect 19035 655 19040 685
rect 19000 650 19040 655
rect 17060 640 17100 650
rect 17060 620 17070 640
rect 17090 620 17100 640
rect 17060 610 17100 620
rect 17240 640 17280 650
rect 17240 620 17250 640
rect 17270 620 17280 640
rect 17240 610 17280 620
rect 17420 640 17460 650
rect 17420 620 17430 640
rect 17450 620 17460 640
rect 17420 610 17460 620
rect 17600 645 17640 650
rect 17600 615 17605 645
rect 17635 615 17640 645
rect 17600 610 17640 615
rect 17690 640 17730 650
rect 17690 620 17700 640
rect 17720 620 17730 640
rect 17690 610 17730 620
rect 17780 640 17820 650
rect 17780 620 17790 640
rect 17810 620 17820 640
rect 17780 610 17820 620
rect 17960 645 18000 650
rect 17960 615 17965 645
rect 17995 615 18000 645
rect 17960 610 18000 615
rect 18140 640 18180 650
rect 18140 620 18150 640
rect 18170 620 18180 640
rect 18140 610 18180 620
rect 18320 640 18360 650
rect 18320 620 18330 640
rect 18350 620 18360 640
rect 18320 610 18360 620
rect 18500 640 18540 650
rect 18500 620 18510 640
rect 18530 620 18540 640
rect 18500 610 18540 620
rect 16780 590 16820 595
rect 16780 560 16785 590
rect 16815 560 16820 590
rect 16780 555 16820 560
rect 16545 535 16585 540
rect 16545 505 16550 535
rect 16580 505 16585 535
rect 16545 500 16585 505
rect 17070 495 17090 610
rect 17250 540 17270 610
rect 17430 595 17450 610
rect 17420 590 17460 595
rect 17420 560 17425 590
rect 17455 560 17460 590
rect 17420 555 17460 560
rect 17240 535 17280 540
rect 17240 505 17245 535
rect 17275 505 17280 535
rect 17240 500 17280 505
rect 17060 490 17100 495
rect 17060 460 17065 490
rect 17095 460 17100 490
rect 17060 455 17100 460
rect 16540 390 16580 395
rect 16540 360 16545 390
rect 16575 360 16580 390
rect 16540 350 16580 360
rect 16540 320 16545 350
rect 16575 320 16580 350
rect 16540 310 16580 320
rect 16540 280 16545 310
rect 16575 280 16580 310
rect 16540 275 16580 280
rect 16660 390 16700 395
rect 16660 360 16665 390
rect 16695 360 16700 390
rect 16660 350 16700 360
rect 16660 320 16665 350
rect 16695 320 16700 350
rect 16660 310 16700 320
rect 16660 280 16665 310
rect 16695 280 16700 310
rect 16660 275 16700 280
rect 16780 390 16820 395
rect 16780 360 16785 390
rect 16815 360 16820 390
rect 16780 350 16820 360
rect 16780 320 16785 350
rect 16815 320 16820 350
rect 16780 310 16820 320
rect 16780 280 16785 310
rect 16815 280 16820 310
rect 16780 275 16820 280
rect 16900 390 16940 395
rect 16900 360 16905 390
rect 16935 360 16940 390
rect 16900 350 16940 360
rect 16900 320 16905 350
rect 16935 320 16940 350
rect 16900 310 16940 320
rect 16900 280 16905 310
rect 16935 280 16940 310
rect 16900 275 16940 280
rect 17020 390 17060 395
rect 17020 360 17025 390
rect 17055 360 17060 390
rect 17020 350 17060 360
rect 17020 320 17025 350
rect 17055 320 17060 350
rect 17020 310 17060 320
rect 17020 280 17025 310
rect 17055 280 17060 310
rect 17020 275 17060 280
rect 17140 390 17180 395
rect 17140 360 17145 390
rect 17175 360 17180 390
rect 17140 350 17180 360
rect 17140 320 17145 350
rect 17175 320 17180 350
rect 17140 310 17180 320
rect 17140 280 17145 310
rect 17175 280 17180 310
rect 17140 275 17180 280
rect 17260 390 17300 395
rect 17260 360 17265 390
rect 17295 360 17300 390
rect 17260 350 17300 360
rect 17260 320 17265 350
rect 17295 320 17300 350
rect 17260 310 17300 320
rect 17260 280 17265 310
rect 17295 280 17300 310
rect 17260 275 17300 280
rect 17380 390 17420 395
rect 17380 360 17385 390
rect 17415 360 17420 390
rect 17380 350 17420 360
rect 17380 320 17385 350
rect 17415 320 17420 350
rect 17380 310 17420 320
rect 17380 280 17385 310
rect 17415 280 17420 310
rect 17380 275 17420 280
rect 17500 390 17540 395
rect 17500 360 17505 390
rect 17535 360 17540 390
rect 17500 350 17540 360
rect 17500 320 17505 350
rect 17535 320 17540 350
rect 17500 310 17540 320
rect 17500 280 17505 310
rect 17535 280 17540 310
rect 17500 275 17540 280
rect 17620 390 17660 395
rect 17620 360 17625 390
rect 17655 360 17660 390
rect 17620 350 17660 360
rect 17620 320 17625 350
rect 17655 320 17660 350
rect 17620 310 17660 320
rect 17620 280 17625 310
rect 17655 280 17660 310
rect 17620 275 17660 280
rect 16550 180 16570 275
rect 16670 180 16690 275
rect 16790 180 16810 275
rect 16910 180 16930 275
rect 17030 180 17050 275
rect 17150 180 17170 275
rect 17270 180 17290 275
rect 17390 180 17410 275
rect 17510 180 17530 275
rect 17630 180 17650 275
rect 17700 180 17720 610
rect 17790 495 17810 610
rect 18150 595 18170 610
rect 18140 590 18180 595
rect 18140 560 18145 590
rect 18175 560 18180 590
rect 18140 555 18180 560
rect 18330 540 18350 610
rect 18320 535 18360 540
rect 18320 505 18325 535
rect 18355 505 18360 535
rect 18320 500 18360 505
rect 18510 495 18530 610
rect 17780 490 17820 495
rect 17780 460 17785 490
rect 17815 460 17820 490
rect 17780 455 17820 460
rect 18500 490 18540 495
rect 18500 460 18505 490
rect 18535 460 18540 490
rect 18500 455 18540 460
rect 17940 390 17980 395
rect 17940 360 17945 390
rect 17975 360 17980 390
rect 17940 350 17980 360
rect 17940 320 17945 350
rect 17975 320 17980 350
rect 17940 310 17980 320
rect 17940 280 17945 310
rect 17975 280 17980 310
rect 17940 275 17980 280
rect 18060 390 18100 395
rect 18060 360 18065 390
rect 18095 360 18100 390
rect 18060 350 18100 360
rect 18060 320 18065 350
rect 18095 320 18100 350
rect 18060 310 18100 320
rect 18060 280 18065 310
rect 18095 280 18100 310
rect 18060 275 18100 280
rect 18180 390 18220 395
rect 18180 360 18185 390
rect 18215 360 18220 390
rect 18180 350 18220 360
rect 18180 320 18185 350
rect 18215 320 18220 350
rect 18180 310 18220 320
rect 18180 280 18185 310
rect 18215 280 18220 310
rect 18180 275 18220 280
rect 18300 390 18340 395
rect 18300 360 18305 390
rect 18335 360 18340 390
rect 18300 350 18340 360
rect 18300 320 18305 350
rect 18335 320 18340 350
rect 18300 310 18340 320
rect 18300 280 18305 310
rect 18335 280 18340 310
rect 18300 275 18340 280
rect 18420 390 18460 395
rect 18420 360 18425 390
rect 18455 360 18460 390
rect 18420 350 18460 360
rect 18420 320 18425 350
rect 18455 320 18460 350
rect 18420 310 18460 320
rect 18420 280 18425 310
rect 18455 280 18460 310
rect 18420 275 18460 280
rect 18540 390 18580 395
rect 18540 360 18545 390
rect 18575 360 18580 390
rect 18540 350 18580 360
rect 18540 320 18545 350
rect 18575 320 18580 350
rect 18540 310 18580 320
rect 18540 280 18545 310
rect 18575 280 18580 310
rect 18540 275 18580 280
rect 18660 390 18700 395
rect 18660 360 18665 390
rect 18695 360 18700 390
rect 18660 350 18700 360
rect 18660 320 18665 350
rect 18695 320 18700 350
rect 18660 310 18700 320
rect 18660 280 18665 310
rect 18695 280 18700 310
rect 18660 275 18700 280
rect 18780 390 18820 395
rect 18780 360 18785 390
rect 18815 360 18820 390
rect 18780 350 18820 360
rect 18780 320 18785 350
rect 18815 320 18820 350
rect 18780 310 18820 320
rect 18780 280 18785 310
rect 18815 280 18820 310
rect 18780 275 18820 280
rect 18900 390 18940 395
rect 18900 360 18905 390
rect 18935 360 18940 390
rect 18900 350 18940 360
rect 18900 320 18905 350
rect 18935 320 18940 350
rect 18900 310 18940 320
rect 18900 280 18905 310
rect 18935 280 18940 310
rect 18900 275 18940 280
rect 19020 390 19060 395
rect 19020 360 19025 390
rect 19055 360 19060 390
rect 19020 350 19060 360
rect 19020 320 19025 350
rect 19055 320 19060 350
rect 19020 310 19060 320
rect 19020 280 19025 310
rect 19055 280 19060 310
rect 19020 275 19060 280
rect 19140 390 19180 395
rect 19140 360 19145 390
rect 19175 360 19180 390
rect 19140 350 19180 360
rect 19140 320 19145 350
rect 19175 320 19180 350
rect 19140 310 19180 320
rect 19140 280 19145 310
rect 19175 280 19180 310
rect 19140 275 19180 280
rect 17950 180 17970 275
rect 18070 180 18090 275
rect 18190 180 18210 275
rect 18310 180 18330 275
rect 18430 180 18450 275
rect 18550 180 18570 275
rect 18670 180 18690 275
rect 18790 180 18810 275
rect 18910 180 18930 275
rect 19030 180 19050 275
rect 19150 180 19170 275
rect 16425 170 16455 180
rect 16425 150 16430 170
rect 16450 150 16455 170
rect 16425 135 16455 150
rect 16480 175 16520 180
rect 16480 145 16485 175
rect 16515 145 16520 175
rect 16480 140 16520 145
rect 16545 170 16575 180
rect 16545 150 16550 170
rect 16570 150 16575 170
rect 16545 140 16575 150
rect 16665 170 16695 180
rect 16665 150 16670 170
rect 16690 150 16695 170
rect 16665 140 16695 150
rect 16785 170 16815 180
rect 16785 150 16790 170
rect 16810 150 16815 170
rect 16785 140 16815 150
rect 16840 175 16880 180
rect 16840 145 16845 175
rect 16875 145 16880 175
rect 16840 140 16880 145
rect 16905 170 16935 180
rect 16905 150 16910 170
rect 16930 150 16935 170
rect 16905 140 16935 150
rect 17025 170 17055 180
rect 17025 150 17030 170
rect 17050 150 17055 170
rect 17025 140 17055 150
rect 17145 170 17175 180
rect 17145 150 17150 170
rect 17170 150 17175 170
rect 17145 140 17175 150
rect 17200 175 17240 180
rect 17200 145 17205 175
rect 17235 145 17240 175
rect 17200 140 17240 145
rect 17265 170 17295 180
rect 17265 150 17270 170
rect 17290 150 17295 170
rect 17265 140 17295 150
rect 17385 170 17415 180
rect 17385 150 17390 170
rect 17410 150 17415 170
rect 17385 140 17415 150
rect 17505 170 17535 180
rect 17505 150 17510 170
rect 17530 150 17535 170
rect 17505 140 17535 150
rect 17560 175 17600 180
rect 17560 145 17565 175
rect 17595 145 17600 175
rect 17560 140 17600 145
rect 17625 170 17655 180
rect 17625 150 17630 170
rect 17650 150 17655 170
rect 17625 135 17655 150
rect 17690 175 17730 180
rect 17690 145 17695 175
rect 17725 145 17730 175
rect 17690 140 17730 145
rect 17870 175 17910 180
rect 17870 145 17875 175
rect 17905 145 17910 175
rect 17870 140 17910 145
rect 17945 170 17975 180
rect 17945 150 17950 170
rect 17970 150 17975 170
rect 16510 0 16550 10
rect 16510 -20 16520 0
rect 16540 -20 16550 0
rect 16510 -30 16550 -20
rect 16600 5 16640 10
rect 16600 -25 16605 5
rect 16635 -25 16640 5
rect 16600 -30 16640 -25
rect 16720 0 16760 10
rect 16720 -20 16730 0
rect 16750 -20 16760 0
rect 16720 -30 16760 -20
rect 16840 0 16880 10
rect 16840 -20 16850 0
rect 16870 -20 16880 0
rect 16840 -30 16880 -20
rect 16960 5 17000 10
rect 16960 -25 16965 5
rect 16995 -25 17000 5
rect 16960 -30 17000 -25
rect 17080 0 17120 10
rect 17080 -20 17090 0
rect 17110 -20 17120 0
rect 17080 -30 17120 -20
rect 17200 0 17240 10
rect 17200 -20 17210 0
rect 17230 -20 17240 0
rect 17200 -30 17240 -20
rect 17320 5 17360 10
rect 17320 -25 17325 5
rect 17355 -25 17360 5
rect 17320 -30 17360 -25
rect 17440 0 17480 10
rect 17440 -20 17450 0
rect 17470 -20 17480 0
rect 17440 -30 17480 -20
rect 17535 0 17565 10
rect 17535 -20 17540 0
rect 17560 -20 17565 0
rect 17535 -30 17565 -20
rect 16520 -50 16540 -30
rect 16730 -50 16750 -30
rect 16850 -50 16870 -30
rect 16510 -55 16550 -50
rect 16510 -85 16515 -55
rect 16545 -85 16550 -55
rect 16510 -90 16550 -85
rect 16720 -55 16760 -50
rect 16720 -85 16725 -55
rect 16755 -85 16760 -55
rect 16720 -90 16760 -85
rect 16840 -55 16880 -50
rect 16840 -85 16845 -55
rect 16875 -85 16880 -55
rect 16840 -90 16880 -85
rect 16970 -105 16990 -30
rect 17090 -50 17110 -30
rect 17210 -50 17230 -30
rect 17450 -50 17470 -30
rect 17540 -50 17560 -30
rect 17080 -55 17120 -50
rect 17080 -85 17085 -55
rect 17115 -85 17120 -55
rect 17080 -90 17120 -85
rect 17200 -55 17240 -50
rect 17200 -85 17205 -55
rect 17235 -85 17240 -55
rect 17200 -90 17240 -85
rect 17440 -55 17480 -50
rect 17440 -85 17445 -55
rect 17475 -85 17480 -55
rect 17440 -90 17480 -85
rect 17530 -55 17570 -50
rect 17530 -85 17535 -55
rect 17565 -85 17570 -55
rect 17530 -90 17570 -85
rect 17090 -105 17110 -90
rect 16960 -115 16990 -105
rect 16960 -135 16965 -115
rect 16985 -135 16990 -115
rect 16960 -145 16990 -135
rect 17007 -110 17037 -105
rect 17007 -145 17037 -140
rect 17090 -115 17120 -105
rect 17090 -135 17095 -115
rect 17115 -135 17120 -115
rect 17090 -145 17120 -135
rect 16315 -460 16320 -430
rect 16350 -460 16355 -430
rect 16315 -2000 16355 -460
rect 17025 -175 17055 -165
rect 17025 -195 17030 -175
rect 17050 -195 17055 -175
rect 17025 -225 17055 -195
rect 17025 -245 17030 -225
rect 17050 -245 17055 -225
rect 17025 -275 17055 -245
rect 17025 -295 17030 -275
rect 17050 -295 17055 -275
rect 17560 -170 17600 -165
rect 17560 -200 17565 -170
rect 17595 -200 17600 -170
rect 17560 -210 17600 -200
rect 17560 -240 17565 -210
rect 17595 -240 17600 -210
rect 17560 -250 17600 -240
rect 17560 -280 17565 -250
rect 17595 -280 17600 -250
rect 17560 -285 17600 -280
rect 17025 -325 17055 -295
rect 17025 -345 17030 -325
rect 17050 -345 17055 -325
rect 17025 -375 17055 -345
rect 17025 -395 17030 -375
rect 17050 -395 17055 -375
rect 17025 -505 17055 -395
rect 17075 -430 17105 -425
rect 17075 -465 17105 -460
rect 16530 -510 16570 -505
rect 16530 -540 16535 -510
rect 16565 -540 16570 -510
rect 16530 -545 16570 -540
rect 17020 -510 17060 -505
rect 17020 -540 17025 -510
rect 17055 -540 17060 -510
rect 17020 -545 17060 -540
rect 16535 -710 16565 -545
rect 16620 -565 16660 -560
rect 16620 -595 16625 -565
rect 16655 -595 16660 -565
rect 16620 -605 16660 -595
rect 16620 -635 16625 -605
rect 16655 -635 16660 -605
rect 16620 -645 16660 -635
rect 16620 -675 16625 -645
rect 16655 -675 16660 -645
rect 16620 -680 16660 -675
rect 16740 -565 16780 -560
rect 16740 -595 16745 -565
rect 16775 -595 16780 -565
rect 16740 -605 16780 -595
rect 16740 -635 16745 -605
rect 16775 -635 16780 -605
rect 16740 -645 16780 -635
rect 16740 -675 16745 -645
rect 16775 -675 16780 -645
rect 16740 -680 16780 -675
rect 16860 -565 16900 -560
rect 16860 -595 16865 -565
rect 16895 -595 16900 -565
rect 16860 -605 16900 -595
rect 16860 -635 16865 -605
rect 16895 -635 16900 -605
rect 16860 -645 16900 -635
rect 16860 -675 16865 -645
rect 16895 -675 16900 -645
rect 16860 -680 16900 -675
rect 16980 -565 17020 -560
rect 16980 -595 16985 -565
rect 17015 -595 17020 -565
rect 16980 -605 17020 -595
rect 16980 -635 16985 -605
rect 17015 -635 17020 -605
rect 16980 -645 17020 -635
rect 16980 -675 16985 -645
rect 17015 -675 17020 -645
rect 16980 -680 17020 -675
rect 17300 -565 17340 -560
rect 17300 -595 17305 -565
rect 17335 -595 17340 -565
rect 17300 -605 17340 -595
rect 17300 -635 17305 -605
rect 17335 -635 17340 -605
rect 17300 -645 17340 -635
rect 17300 -675 17305 -645
rect 17335 -675 17340 -645
rect 17300 -680 17340 -675
rect 17420 -565 17460 -560
rect 17420 -595 17425 -565
rect 17455 -595 17460 -565
rect 17420 -605 17460 -595
rect 17420 -635 17425 -605
rect 17455 -635 17460 -605
rect 17420 -645 17460 -635
rect 17420 -675 17425 -645
rect 17455 -675 17460 -645
rect 17420 -680 17460 -675
rect 17540 -565 17580 -560
rect 17540 -595 17545 -565
rect 17575 -595 17580 -565
rect 17540 -605 17580 -595
rect 17540 -635 17545 -605
rect 17575 -635 17580 -605
rect 17540 -645 17580 -635
rect 17540 -675 17545 -645
rect 17575 -675 17580 -645
rect 17700 -655 17720 140
rect 17740 -170 17860 -165
rect 17740 -200 17745 -170
rect 17775 -200 17785 -170
rect 17815 -200 17825 -170
rect 17855 -200 17860 -170
rect 17740 -210 17860 -200
rect 17740 -240 17745 -210
rect 17775 -240 17785 -210
rect 17815 -240 17825 -210
rect 17855 -240 17860 -210
rect 17740 -250 17860 -240
rect 17740 -280 17745 -250
rect 17775 -280 17785 -250
rect 17815 -280 17825 -250
rect 17855 -280 17860 -250
rect 17540 -680 17580 -675
rect 17695 -665 17725 -655
rect 17695 -685 17700 -665
rect 17720 -685 17725 -665
rect 17695 -695 17725 -685
rect 16535 -730 16540 -710
rect 16560 -730 16565 -710
rect 16535 -760 16565 -730
rect 16535 -780 16540 -760
rect 16560 -780 16565 -760
rect 16535 -810 16565 -780
rect 16535 -830 16540 -810
rect 16560 -830 16565 -810
rect 16535 -860 16565 -830
rect 16535 -880 16540 -860
rect 16560 -880 16565 -860
rect 16535 -910 16565 -880
rect 16535 -930 16540 -910
rect 16560 -930 16565 -910
rect 16535 -940 16565 -930
rect 17110 -965 17150 -960
rect 17110 -995 17115 -965
rect 17145 -995 17150 -965
rect 17110 -1005 17150 -995
rect 17110 -1035 17115 -1005
rect 17145 -1035 17150 -1005
rect 17110 -1045 17150 -1035
rect 17110 -1075 17115 -1045
rect 17145 -1075 17150 -1045
rect 17110 -1080 17150 -1075
rect 17740 -965 17860 -280
rect 17880 -655 17900 140
rect 17945 135 17975 150
rect 18000 175 18040 180
rect 18000 145 18005 175
rect 18035 145 18040 175
rect 18000 140 18040 145
rect 18065 170 18095 180
rect 18065 150 18070 170
rect 18090 150 18095 170
rect 18065 140 18095 150
rect 18185 170 18215 180
rect 18185 150 18190 170
rect 18210 150 18215 170
rect 18185 140 18215 150
rect 18305 170 18335 180
rect 18305 150 18310 170
rect 18330 150 18335 170
rect 18305 140 18335 150
rect 18360 175 18400 180
rect 18360 145 18365 175
rect 18395 145 18400 175
rect 18360 140 18400 145
rect 18425 170 18455 180
rect 18425 150 18430 170
rect 18450 150 18455 170
rect 18425 140 18455 150
rect 18545 170 18575 180
rect 18545 150 18550 170
rect 18570 150 18575 170
rect 18545 140 18575 150
rect 18665 170 18695 180
rect 18665 150 18670 170
rect 18690 150 18695 170
rect 18665 140 18695 150
rect 18720 175 18760 180
rect 18720 145 18725 175
rect 18755 145 18760 175
rect 18720 140 18760 145
rect 18785 170 18815 180
rect 18785 150 18790 170
rect 18810 150 18815 170
rect 18785 140 18815 150
rect 18905 170 18935 180
rect 18905 150 18910 170
rect 18930 150 18935 170
rect 18905 140 18935 150
rect 19025 170 19055 180
rect 19025 150 19030 170
rect 19050 150 19055 170
rect 19025 140 19055 150
rect 19080 175 19120 180
rect 19080 145 19085 175
rect 19115 145 19120 175
rect 19080 140 19120 145
rect 19145 170 19175 180
rect 19145 150 19150 170
rect 19170 150 19175 170
rect 19145 135 19175 150
rect 18035 0 18065 10
rect 18035 -20 18040 0
rect 18060 -20 18065 0
rect 18035 -30 18065 -20
rect 18120 0 18160 10
rect 18120 -20 18130 0
rect 18150 -20 18160 0
rect 18120 -30 18160 -20
rect 18240 5 18280 10
rect 18240 -25 18245 5
rect 18275 -25 18280 5
rect 18240 -30 18280 -25
rect 18360 0 18400 10
rect 18360 -20 18370 0
rect 18390 -20 18400 0
rect 18360 -30 18400 -20
rect 18480 0 18520 10
rect 18480 -20 18490 0
rect 18510 -20 18520 0
rect 18480 -30 18520 -20
rect 18600 5 18640 10
rect 18600 -25 18605 5
rect 18635 -25 18640 5
rect 18600 -30 18640 -25
rect 18720 0 18760 10
rect 18720 -20 18730 0
rect 18750 -20 18760 0
rect 18720 -30 18760 -20
rect 18840 0 18880 10
rect 18840 -20 18850 0
rect 18870 -20 18880 0
rect 18840 -30 18880 -20
rect 18960 5 19000 10
rect 18960 -25 18965 5
rect 18995 -25 19000 5
rect 18960 -30 19000 -25
rect 19050 0 19090 10
rect 19050 -20 19060 0
rect 19080 -20 19090 0
rect 19050 -30 19090 -20
rect 18040 -50 18060 -30
rect 18130 -50 18150 -30
rect 18370 -50 18390 -30
rect 18490 -50 18510 -30
rect 18030 -55 18070 -50
rect 18030 -85 18035 -55
rect 18065 -85 18070 -55
rect 18030 -90 18070 -85
rect 18120 -55 18160 -50
rect 18120 -85 18125 -55
rect 18155 -85 18160 -55
rect 18120 -90 18160 -85
rect 18360 -55 18400 -50
rect 18360 -85 18365 -55
rect 18395 -85 18400 -55
rect 18360 -90 18400 -85
rect 18480 -55 18520 -50
rect 18480 -85 18485 -55
rect 18515 -85 18520 -55
rect 18480 -90 18520 -85
rect 18490 -105 18510 -90
rect 18610 -105 18630 -30
rect 18730 -50 18750 -30
rect 18850 -50 18870 -30
rect 19060 -50 19080 -30
rect 18720 -55 18760 -50
rect 18720 -85 18725 -55
rect 18755 -85 18760 -55
rect 18720 -90 18760 -85
rect 18840 -55 18880 -50
rect 18840 -85 18845 -55
rect 18875 -85 18880 -55
rect 18840 -90 18880 -85
rect 19050 -55 19090 -50
rect 19050 -85 19055 -55
rect 19085 -85 19090 -55
rect 19050 -90 19090 -85
rect 18480 -115 18510 -105
rect 18480 -135 18485 -115
rect 18505 -135 18510 -115
rect 18480 -145 18510 -135
rect 18563 -110 18593 -105
rect 18563 -145 18593 -140
rect 18610 -115 18640 -105
rect 18610 -135 18615 -115
rect 18635 -135 18640 -115
rect 18610 -145 18640 -135
rect 18000 -170 18040 -165
rect 18000 -200 18005 -170
rect 18035 -200 18040 -170
rect 18000 -210 18040 -200
rect 18000 -240 18005 -210
rect 18035 -240 18040 -210
rect 18000 -250 18040 -240
rect 18000 -280 18005 -250
rect 18035 -280 18040 -250
rect 18000 -285 18040 -280
rect 19335 -425 19355 1175
rect 19415 495 19435 1795
rect 19405 490 19445 495
rect 19405 460 19410 490
rect 19440 460 19445 490
rect 19405 455 19445 460
rect 19415 -105 19435 455
rect 19405 -110 19445 -105
rect 19405 -140 19410 -110
rect 19440 -140 19445 -110
rect 19405 -145 19445 -140
rect 18495 -430 18525 -425
rect 18495 -465 18525 -460
rect 18545 -435 18575 -425
rect 18545 -455 18550 -435
rect 18570 -455 18575 -435
rect 18545 -465 18575 -455
rect 19325 -430 19365 -425
rect 19325 -460 19330 -430
rect 19360 -460 19365 -430
rect 19325 -465 19365 -460
rect 18550 -505 18570 -465
rect 18540 -510 18580 -505
rect 18540 -540 18545 -510
rect 18575 -540 18580 -510
rect 18540 -545 18580 -540
rect 19030 -510 19070 -505
rect 19030 -540 19035 -510
rect 19065 -540 19070 -510
rect 19030 -545 19070 -540
rect 18020 -565 18060 -560
rect 18020 -595 18025 -565
rect 18055 -595 18060 -565
rect 18020 -605 18060 -595
rect 18020 -635 18025 -605
rect 18055 -635 18060 -605
rect 18020 -645 18060 -635
rect 17875 -665 17905 -655
rect 17875 -685 17880 -665
rect 17900 -685 17905 -665
rect 18020 -675 18025 -645
rect 18055 -675 18060 -645
rect 18020 -680 18060 -675
rect 18140 -565 18180 -560
rect 18140 -595 18145 -565
rect 18175 -595 18180 -565
rect 18140 -605 18180 -595
rect 18140 -635 18145 -605
rect 18175 -635 18180 -605
rect 18140 -645 18180 -635
rect 18140 -675 18145 -645
rect 18175 -675 18180 -645
rect 18140 -680 18180 -675
rect 18260 -565 18300 -560
rect 18260 -595 18265 -565
rect 18295 -595 18300 -565
rect 18260 -605 18300 -595
rect 18260 -635 18265 -605
rect 18295 -635 18300 -605
rect 18260 -645 18300 -635
rect 18260 -675 18265 -645
rect 18295 -675 18300 -645
rect 18260 -680 18300 -675
rect 18580 -565 18620 -560
rect 18580 -595 18585 -565
rect 18615 -595 18620 -565
rect 18580 -605 18620 -595
rect 18580 -635 18585 -605
rect 18615 -635 18620 -605
rect 18580 -645 18620 -635
rect 18580 -675 18585 -645
rect 18615 -675 18620 -645
rect 18580 -680 18620 -675
rect 18700 -565 18740 -560
rect 18700 -595 18705 -565
rect 18735 -595 18740 -565
rect 18700 -605 18740 -595
rect 18700 -635 18705 -605
rect 18735 -635 18740 -605
rect 18700 -645 18740 -635
rect 18700 -675 18705 -645
rect 18735 -675 18740 -645
rect 18700 -680 18740 -675
rect 18820 -565 18860 -560
rect 18820 -595 18825 -565
rect 18855 -595 18860 -565
rect 18820 -605 18860 -595
rect 18820 -635 18825 -605
rect 18855 -635 18860 -605
rect 18820 -645 18860 -635
rect 18820 -675 18825 -645
rect 18855 -675 18860 -645
rect 18820 -680 18860 -675
rect 18940 -565 18980 -560
rect 18940 -595 18945 -565
rect 18975 -595 18980 -565
rect 18940 -605 18980 -595
rect 18940 -635 18945 -605
rect 18975 -635 18980 -605
rect 18940 -645 18980 -635
rect 18940 -675 18945 -645
rect 18975 -675 18980 -645
rect 19040 -660 19060 -545
rect 18940 -680 18980 -675
rect 19030 -670 19070 -660
rect 17875 -695 17905 -685
rect 19030 -690 19040 -670
rect 19060 -690 19070 -670
rect 19030 -700 19070 -690
rect 17740 -995 17745 -965
rect 17775 -995 17785 -965
rect 17815 -995 17825 -965
rect 17855 -995 17860 -965
rect 17740 -1005 17860 -995
rect 17740 -1035 17745 -1005
rect 17775 -1035 17785 -1005
rect 17815 -1035 17825 -1005
rect 17855 -1035 17860 -1005
rect 17740 -1045 17860 -1035
rect 17740 -1075 17745 -1045
rect 17775 -1075 17785 -1045
rect 17815 -1075 17825 -1045
rect 17855 -1075 17860 -1045
rect 17740 -1080 17860 -1075
rect 18450 -965 18490 -960
rect 18450 -995 18455 -965
rect 18485 -995 18490 -965
rect 18450 -1005 18490 -995
rect 18450 -1035 18455 -1005
rect 18485 -1035 18490 -1005
rect 18450 -1045 18490 -1035
rect 18450 -1075 18455 -1045
rect 18485 -1075 18490 -1045
rect 18450 -1080 18490 -1075
rect 16740 -1100 16780 -1095
rect 16740 -1130 16745 -1100
rect 16775 -1130 16780 -1100
rect 16740 -1135 16780 -1130
rect 16820 -1100 16860 -1095
rect 16820 -1130 16825 -1100
rect 16855 -1130 16860 -1100
rect 16820 -1135 16860 -1130
rect 16900 -1100 16940 -1095
rect 16900 -1130 16905 -1100
rect 16935 -1130 16940 -1100
rect 16900 -1135 16940 -1130
rect 16980 -1100 17020 -1095
rect 16980 -1130 16985 -1100
rect 17015 -1130 17020 -1100
rect 16980 -1135 17020 -1130
rect 17060 -1100 17100 -1095
rect 17060 -1130 17065 -1100
rect 17095 -1130 17100 -1100
rect 17060 -1135 17100 -1130
rect 17140 -1100 17180 -1095
rect 17140 -1130 17145 -1100
rect 17175 -1130 17180 -1100
rect 17140 -1135 17180 -1130
rect 17220 -1100 17260 -1095
rect 17220 -1130 17225 -1100
rect 17255 -1130 17260 -1100
rect 17220 -1135 17260 -1130
rect 17300 -1100 17340 -1095
rect 17300 -1130 17305 -1100
rect 17335 -1130 17340 -1100
rect 17300 -1135 17340 -1130
rect 17380 -1100 17420 -1095
rect 17380 -1130 17385 -1100
rect 17415 -1130 17420 -1100
rect 17380 -1135 17420 -1130
rect 17460 -1100 17500 -1095
rect 17460 -1130 17465 -1100
rect 17495 -1130 17500 -1100
rect 17460 -1135 17500 -1130
rect 17540 -1100 17580 -1095
rect 17540 -1130 17545 -1100
rect 17575 -1130 17580 -1100
rect 17540 -1135 17580 -1130
rect 17620 -1100 17660 -1095
rect 17620 -1130 17625 -1100
rect 17655 -1130 17660 -1100
rect 17620 -1135 17660 -1130
rect 17700 -1100 17740 -1095
rect 17700 -1130 17705 -1100
rect 17735 -1130 17740 -1100
rect 17700 -1135 17740 -1130
rect 17780 -1100 17820 -1095
rect 17780 -1130 17785 -1100
rect 17815 -1130 17820 -1100
rect 17780 -1135 17820 -1130
rect 17860 -1100 17900 -1095
rect 17860 -1130 17865 -1100
rect 17895 -1130 17900 -1100
rect 17860 -1135 17900 -1130
rect 17940 -1100 17980 -1095
rect 17940 -1130 17945 -1100
rect 17975 -1130 17980 -1100
rect 17940 -1135 17980 -1130
rect 18020 -1100 18060 -1095
rect 18020 -1130 18025 -1100
rect 18055 -1130 18060 -1100
rect 18020 -1135 18060 -1130
rect 18100 -1100 18140 -1095
rect 18100 -1130 18105 -1100
rect 18135 -1130 18140 -1100
rect 18100 -1135 18140 -1130
rect 18180 -1100 18220 -1095
rect 18180 -1130 18185 -1100
rect 18215 -1130 18220 -1100
rect 18180 -1135 18220 -1130
rect 18260 -1100 18300 -1095
rect 18260 -1130 18265 -1100
rect 18295 -1130 18300 -1100
rect 18260 -1135 18300 -1130
rect 18340 -1100 18380 -1095
rect 18340 -1130 18345 -1100
rect 18375 -1130 18380 -1100
rect 18340 -1135 18380 -1130
rect 18420 -1100 18460 -1095
rect 18420 -1130 18425 -1100
rect 18455 -1130 18460 -1100
rect 18420 -1135 18460 -1130
rect 18500 -1100 18540 -1095
rect 18500 -1130 18505 -1100
rect 18535 -1130 18540 -1100
rect 18500 -1135 18540 -1130
rect 18580 -1100 18620 -1095
rect 18580 -1130 18585 -1100
rect 18615 -1130 18620 -1100
rect 18580 -1135 18620 -1130
rect 18660 -1100 18700 -1095
rect 18660 -1130 18665 -1100
rect 18695 -1130 18700 -1100
rect 18660 -1135 18700 -1130
rect 18740 -1100 18780 -1095
rect 18740 -1130 18745 -1100
rect 18775 -1130 18780 -1100
rect 18740 -1135 18780 -1130
rect 18895 -1165 18935 -1160
rect 16700 -1185 16740 -1180
rect 16700 -1215 16705 -1185
rect 16735 -1215 16740 -1185
rect 16700 -1220 16740 -1215
rect 18895 -1195 18900 -1165
rect 18930 -1195 18935 -1165
rect 18895 -1205 18935 -1195
rect 18895 -1235 18900 -1205
rect 18930 -1235 18935 -1205
rect 18895 -1240 18935 -1235
rect 16655 -1355 16695 -1350
rect 16655 -1385 16660 -1355
rect 16690 -1385 16695 -1355
rect 16655 -1390 16695 -1385
rect 16765 -1355 16805 -1350
rect 16765 -1385 16770 -1355
rect 16800 -1385 16805 -1355
rect 16765 -1390 16805 -1385
rect 17300 -1355 17340 -1350
rect 17300 -1385 17305 -1355
rect 17335 -1385 17340 -1355
rect 17300 -1390 17340 -1385
rect 17780 -1355 17820 -1350
rect 17780 -1385 17785 -1355
rect 17815 -1385 17820 -1355
rect 17780 -1390 17820 -1385
rect 18260 -1355 18300 -1350
rect 18260 -1385 18265 -1355
rect 18295 -1385 18300 -1355
rect 18260 -1390 18300 -1385
rect 16600 -1410 16640 -1405
rect 16600 -1440 16605 -1410
rect 16635 -1440 16640 -1410
rect 16600 -1450 16640 -1440
rect 16600 -1480 16605 -1450
rect 16635 -1480 16640 -1450
rect 16600 -1490 16640 -1480
rect 16600 -1520 16605 -1490
rect 16635 -1520 16640 -1490
rect 16600 -1525 16640 -1520
rect 16660 -1495 16690 -1390
rect 16660 -1515 16665 -1495
rect 16685 -1515 16690 -1495
rect 16660 -1525 16690 -1515
rect 16710 -1410 16750 -1405
rect 16710 -1440 16715 -1410
rect 16745 -1440 16750 -1410
rect 16710 -1450 16750 -1440
rect 16710 -1480 16715 -1450
rect 16745 -1480 16750 -1450
rect 16710 -1490 16750 -1480
rect 16710 -1520 16715 -1490
rect 16745 -1520 16750 -1490
rect 16710 -1525 16750 -1520
rect 16770 -1495 16800 -1390
rect 16770 -1515 16775 -1495
rect 16795 -1515 16800 -1495
rect 16770 -1525 16800 -1515
rect 16820 -1410 16860 -1405
rect 16820 -1440 16825 -1410
rect 16855 -1440 16860 -1410
rect 16820 -1450 16860 -1440
rect 16820 -1480 16825 -1450
rect 16855 -1480 16860 -1450
rect 16820 -1490 16860 -1480
rect 16820 -1520 16825 -1490
rect 16855 -1520 16860 -1490
rect 16820 -1525 16860 -1520
rect 16880 -1410 16920 -1405
rect 16880 -1440 16885 -1410
rect 16915 -1440 16920 -1410
rect 16880 -1450 16920 -1440
rect 16880 -1480 16885 -1450
rect 16915 -1480 16920 -1450
rect 16880 -1490 16920 -1480
rect 16880 -1520 16885 -1490
rect 16915 -1520 16920 -1490
rect 16880 -1525 16920 -1520
rect 17025 -1410 17065 -1405
rect 17025 -1440 17030 -1410
rect 17060 -1440 17065 -1410
rect 17025 -1450 17065 -1440
rect 17025 -1480 17030 -1450
rect 17060 -1480 17065 -1450
rect 17025 -1490 17065 -1480
rect 17025 -1520 17030 -1490
rect 17060 -1520 17065 -1490
rect 17025 -1525 17065 -1520
rect 17135 -1410 17175 -1405
rect 17135 -1440 17140 -1410
rect 17170 -1440 17175 -1410
rect 17135 -1450 17175 -1440
rect 17135 -1480 17140 -1450
rect 17170 -1480 17175 -1450
rect 17135 -1490 17175 -1480
rect 17135 -1520 17140 -1490
rect 17170 -1520 17175 -1490
rect 17135 -1525 17175 -1520
rect 17245 -1410 17285 -1405
rect 17245 -1440 17250 -1410
rect 17280 -1440 17285 -1410
rect 17245 -1450 17285 -1440
rect 17245 -1480 17250 -1450
rect 17280 -1480 17285 -1450
rect 17245 -1490 17285 -1480
rect 17245 -1520 17250 -1490
rect 17280 -1520 17285 -1490
rect 17245 -1525 17285 -1520
rect 17305 -1495 17335 -1390
rect 17305 -1515 17310 -1495
rect 17330 -1515 17335 -1495
rect 17305 -1525 17335 -1515
rect 17355 -1410 17395 -1405
rect 17355 -1440 17360 -1410
rect 17390 -1440 17395 -1410
rect 17355 -1450 17395 -1440
rect 17355 -1480 17360 -1450
rect 17390 -1480 17395 -1450
rect 17355 -1490 17395 -1480
rect 17355 -1520 17360 -1490
rect 17390 -1520 17395 -1490
rect 17355 -1525 17395 -1520
rect 17465 -1410 17505 -1405
rect 17465 -1440 17470 -1410
rect 17500 -1440 17505 -1410
rect 17465 -1450 17505 -1440
rect 17465 -1480 17470 -1450
rect 17500 -1480 17505 -1450
rect 17465 -1490 17505 -1480
rect 17465 -1520 17470 -1490
rect 17500 -1520 17505 -1490
rect 17465 -1525 17505 -1520
rect 17615 -1410 17655 -1405
rect 17615 -1440 17620 -1410
rect 17650 -1440 17655 -1410
rect 17615 -1450 17655 -1440
rect 17615 -1480 17620 -1450
rect 17650 -1480 17655 -1450
rect 17615 -1490 17655 -1480
rect 17615 -1520 17620 -1490
rect 17650 -1520 17655 -1490
rect 17615 -1525 17655 -1520
rect 17725 -1410 17765 -1405
rect 17725 -1440 17730 -1410
rect 17760 -1440 17765 -1410
rect 17725 -1450 17765 -1440
rect 17725 -1480 17730 -1450
rect 17760 -1480 17765 -1450
rect 17725 -1490 17765 -1480
rect 17725 -1520 17730 -1490
rect 17760 -1520 17765 -1490
rect 17725 -1525 17765 -1520
rect 17785 -1495 17815 -1390
rect 17785 -1515 17790 -1495
rect 17810 -1515 17815 -1495
rect 17785 -1525 17815 -1515
rect 17835 -1410 17875 -1405
rect 17835 -1440 17840 -1410
rect 17870 -1440 17875 -1410
rect 17835 -1450 17875 -1440
rect 17835 -1480 17840 -1450
rect 17870 -1480 17875 -1450
rect 17835 -1490 17875 -1480
rect 17835 -1520 17840 -1490
rect 17870 -1520 17875 -1490
rect 17835 -1525 17875 -1520
rect 17945 -1410 17985 -1405
rect 17945 -1440 17950 -1410
rect 17980 -1440 17985 -1410
rect 17945 -1450 17985 -1440
rect 17945 -1480 17950 -1450
rect 17980 -1480 17985 -1450
rect 17945 -1490 17985 -1480
rect 17945 -1520 17950 -1490
rect 17980 -1520 17985 -1490
rect 17945 -1525 17985 -1520
rect 18095 -1410 18135 -1405
rect 18095 -1440 18100 -1410
rect 18130 -1440 18135 -1410
rect 18095 -1450 18135 -1440
rect 18095 -1480 18100 -1450
rect 18130 -1480 18135 -1450
rect 18095 -1490 18135 -1480
rect 18095 -1520 18100 -1490
rect 18130 -1520 18135 -1490
rect 18095 -1525 18135 -1520
rect 18205 -1410 18245 -1405
rect 18205 -1440 18210 -1410
rect 18240 -1440 18245 -1410
rect 18205 -1450 18245 -1440
rect 18205 -1480 18210 -1450
rect 18240 -1480 18245 -1450
rect 18205 -1490 18245 -1480
rect 18205 -1520 18210 -1490
rect 18240 -1520 18245 -1490
rect 18205 -1525 18245 -1520
rect 18265 -1495 18295 -1390
rect 18265 -1515 18270 -1495
rect 18290 -1515 18295 -1495
rect 18265 -1525 18295 -1515
rect 18315 -1410 18355 -1405
rect 18315 -1440 18320 -1410
rect 18350 -1440 18355 -1410
rect 18315 -1450 18355 -1440
rect 18315 -1480 18320 -1450
rect 18350 -1480 18355 -1450
rect 18315 -1490 18355 -1480
rect 18315 -1520 18320 -1490
rect 18350 -1520 18355 -1490
rect 18315 -1525 18355 -1520
rect 18425 -1410 18465 -1405
rect 18425 -1440 18430 -1410
rect 18460 -1440 18465 -1410
rect 18425 -1450 18465 -1440
rect 18425 -1480 18430 -1450
rect 18460 -1480 18465 -1450
rect 18425 -1490 18465 -1480
rect 18425 -1520 18430 -1490
rect 18460 -1520 18465 -1490
rect 18425 -1525 18465 -1520
rect 18535 -1410 18575 -1405
rect 18535 -1440 18540 -1410
rect 18570 -1440 18575 -1410
rect 18535 -1450 18575 -1440
rect 18535 -1480 18540 -1450
rect 18570 -1480 18575 -1450
rect 18535 -1490 18575 -1480
rect 18535 -1520 18540 -1490
rect 18570 -1520 18575 -1490
rect 18535 -1525 18575 -1520
rect 17195 -1555 17225 -1545
rect 17195 -1575 17200 -1555
rect 17220 -1575 17225 -1555
rect 17195 -1605 17225 -1575
rect 17195 -1625 17200 -1605
rect 17220 -1625 17225 -1605
rect 17195 -1655 17225 -1625
rect 17415 -1555 17445 -1545
rect 17415 -1575 17420 -1555
rect 17440 -1575 17445 -1555
rect 17415 -1605 17445 -1575
rect 17415 -1625 17420 -1605
rect 17440 -1625 17445 -1605
rect 17415 -1655 17445 -1625
rect 18155 -1555 18185 -1545
rect 18155 -1575 18160 -1555
rect 18180 -1575 18185 -1555
rect 18155 -1605 18185 -1575
rect 18155 -1625 18160 -1605
rect 18180 -1625 18185 -1605
rect 18155 -1655 18185 -1625
rect 18375 -1555 18405 -1545
rect 18375 -1575 18380 -1555
rect 18400 -1575 18405 -1555
rect 18375 -1605 18405 -1575
rect 18375 -1625 18380 -1605
rect 18400 -1625 18405 -1605
rect 18375 -1655 18405 -1625
rect 16765 -1665 16805 -1655
rect 16765 -1685 16775 -1665
rect 16795 -1685 16805 -1665
rect 16765 -1695 16805 -1685
rect 17080 -1665 17120 -1655
rect 17080 -1685 17090 -1665
rect 17110 -1685 17120 -1665
rect 17080 -1695 17120 -1685
rect 17190 -1660 17230 -1655
rect 17190 -1690 17195 -1660
rect 17225 -1690 17230 -1660
rect 16775 -1860 16795 -1695
rect 17090 -1710 17110 -1695
rect 17080 -1715 17120 -1710
rect 17080 -1745 17085 -1715
rect 17115 -1745 17120 -1715
rect 17080 -1750 17120 -1745
rect 17190 -1770 17230 -1690
rect 17300 -1665 17340 -1655
rect 17300 -1685 17310 -1665
rect 17330 -1685 17340 -1665
rect 17300 -1695 17340 -1685
rect 17410 -1660 17450 -1655
rect 17410 -1690 17415 -1660
rect 17445 -1690 17450 -1660
rect 17410 -1695 17450 -1690
rect 17670 -1660 17710 -1655
rect 17670 -1690 17675 -1660
rect 17705 -1690 17710 -1660
rect 17670 -1695 17710 -1690
rect 17780 -1660 17820 -1655
rect 17780 -1690 17785 -1660
rect 17815 -1690 17820 -1660
rect 17780 -1695 17820 -1690
rect 17890 -1660 17930 -1655
rect 17890 -1690 17895 -1660
rect 17925 -1690 17930 -1660
rect 17890 -1695 17930 -1690
rect 18150 -1660 18190 -1655
rect 18150 -1690 18155 -1660
rect 18185 -1690 18190 -1660
rect 18150 -1695 18190 -1690
rect 18260 -1665 18300 -1655
rect 18260 -1685 18270 -1665
rect 18290 -1685 18300 -1665
rect 18260 -1695 18300 -1685
rect 18370 -1660 18410 -1655
rect 18370 -1690 18375 -1660
rect 18405 -1690 18410 -1660
rect 18370 -1695 18410 -1690
rect 18480 -1665 18520 -1655
rect 18480 -1685 18490 -1665
rect 18510 -1685 18520 -1665
rect 18480 -1695 18520 -1685
rect 17310 -1710 17330 -1695
rect 17300 -1715 17340 -1710
rect 17300 -1745 17305 -1715
rect 17335 -1745 17340 -1715
rect 17300 -1750 17340 -1745
rect 17190 -1800 17195 -1770
rect 17225 -1800 17230 -1770
rect 17190 -1805 17230 -1800
rect 16765 -1865 16805 -1860
rect 16765 -1895 16770 -1865
rect 16800 -1895 16805 -1865
rect 17790 -1895 17810 -1695
rect 18270 -1710 18290 -1695
rect 18260 -1715 18300 -1710
rect 18260 -1745 18265 -1715
rect 18295 -1745 18300 -1715
rect 18260 -1750 18300 -1745
rect 18380 -1765 18400 -1695
rect 18490 -1710 18510 -1695
rect 18480 -1715 18520 -1710
rect 18480 -1745 18485 -1715
rect 18515 -1745 18520 -1715
rect 18480 -1750 18520 -1745
rect 18370 -1770 18410 -1765
rect 18370 -1800 18375 -1770
rect 18405 -1800 18410 -1770
rect 18370 -1805 18410 -1800
rect 16765 -1900 16805 -1895
rect 17780 -1900 17820 -1895
rect 17780 -1930 17785 -1900
rect 17815 -1930 17820 -1900
rect 17780 -1935 17820 -1930
rect 19335 -1945 19355 -465
rect 19325 -1950 19365 -1945
rect 19325 -1980 19330 -1950
rect 19360 -1980 19365 -1950
rect 19325 -1985 19365 -1980
rect 16315 -2030 16320 -2000
rect 16350 -2030 16355 -2000
rect 16315 -2035 16355 -2030
rect 17425 -2035 17430 -2000
rect 17465 -2035 17470 -2000
rect 18124 -2035 18129 -2000
rect 18164 -2035 18169 -2000
rect 18830 -2005 18870 -2000
rect 18830 -2035 18835 -2005
rect 18865 -2035 18870 -2005
rect 17425 -2060 17465 -2035
rect 17425 -2090 17430 -2060
rect 17460 -2090 17465 -2060
rect 17425 -2095 17465 -2090
rect 16260 -2130 16265 -2100
rect 16295 -2130 16300 -2100
rect 16260 -2135 16300 -2130
rect 16480 -2100 16520 -2095
rect 16480 -2130 16485 -2100
rect 16515 -2130 16520 -2100
rect 16480 -2895 16520 -2130
rect 16485 -2900 16520 -2895
rect 16485 -2940 16520 -2935
rect 16730 -2100 16770 -2095
rect 16730 -2130 16735 -2100
rect 16765 -2130 16770 -2100
rect 16160 -3025 16195 -3020
rect 16160 -3065 16195 -3060
rect 16730 -3105 16770 -2130
rect 15820 -3115 15860 -3110
rect 15820 -3145 15825 -3115
rect 15855 -3145 15860 -3115
rect 15820 -3150 15860 -3145
rect 15950 -3116 15985 -3110
rect 16730 -3135 16735 -3105
rect 16765 -3135 16770 -3105
rect 16730 -3140 16770 -3135
rect 16945 -2615 18655 -2265
rect 15830 -4260 15850 -3150
rect 15950 -3156 15985 -3151
rect 16945 -3625 17295 -2615
rect 17625 -3105 17975 -2945
rect 17625 -3135 17785 -3105
rect 17815 -3135 17975 -3105
rect 17625 -3295 17975 -3135
rect 18305 -3105 18655 -2615
rect 18305 -3135 18620 -3105
rect 18650 -3135 18655 -3105
rect 18305 -3625 18655 -3135
rect 18830 -3105 18870 -2035
rect 19080 -2060 19120 -2055
rect 19080 -2090 19085 -2060
rect 19115 -2090 19120 -2060
rect 19080 -2895 19120 -2090
rect 19080 -2900 19115 -2895
rect 19080 -2940 19115 -2935
rect 19415 -2992 19435 -145
rect 19545 -1895 19565 1795
rect 19610 1615 19650 1620
rect 19610 1585 19615 1615
rect 19645 1585 19650 1615
rect 19610 685 19650 1585
rect 19610 655 19615 685
rect 19645 655 19650 685
rect 19610 175 19650 655
rect 19610 145 19615 175
rect 19645 145 19650 175
rect 19535 -1900 19575 -1895
rect 19535 -1930 19540 -1900
rect 19570 -1930 19575 -1900
rect 19535 -1935 19575 -1930
rect 19405 -2997 19440 -2992
rect 19405 -3037 19440 -3032
rect 18830 -3135 18835 -3105
rect 18865 -3135 18870 -3105
rect 18830 -3140 18870 -3135
rect 19610 -3115 19650 145
rect 19785 -1765 19805 1795
rect 19830 -55 19870 -50
rect 19830 -85 19835 -55
rect 19865 -85 19870 -55
rect 19830 -90 19870 -85
rect 19775 -1770 19815 -1765
rect 19775 -1800 19780 -1770
rect 19810 -1800 19815 -1770
rect 19775 -1805 19815 -1800
rect 19610 -3160 19645 -3150
rect 15950 -3789 15985 -3784
rect 15950 -3829 15985 -3824
rect 15820 -4265 15860 -4260
rect 15820 -4295 15825 -4265
rect 15855 -4295 15860 -4265
rect 15820 -4300 15860 -4295
rect 15725 -4315 15765 -4310
rect 15725 -4345 15730 -4315
rect 15760 -4345 15765 -4315
rect 15725 -4350 15765 -4345
rect 15960 -4355 15980 -3829
rect 16280 -3894 16315 -3889
rect 16280 -3934 16315 -3929
rect 16290 -4185 16310 -3934
rect 16605 -3969 16640 -3964
rect 16945 -3975 18655 -3625
rect 19610 -3789 19645 -3784
rect 19610 -3829 19645 -3824
rect 19285 -3894 19320 -3889
rect 19285 -3934 19320 -3929
rect 18960 -3969 18995 -3964
rect 16605 -4009 16640 -4004
rect 18960 -4009 18995 -4004
rect 16615 -4185 16635 -4009
rect 16280 -4190 16320 -4185
rect 16280 -4220 16285 -4190
rect 16315 -4220 16320 -4190
rect 16280 -4225 16320 -4220
rect 16605 -4190 16645 -4185
rect 16605 -4220 16610 -4190
rect 16640 -4220 16645 -4190
rect 16605 -4225 16645 -4220
rect 17250 -4265 17300 -4255
rect 18965 -4260 18985 -4009
rect 19290 -4260 19310 -3934
rect 17250 -4295 17260 -4265
rect 17290 -4295 17300 -4265
rect 17250 -4305 17300 -4295
rect 17780 -4265 17820 -4260
rect 17780 -4295 17785 -4265
rect 17815 -4295 17820 -4265
rect 17780 -4300 17820 -4295
rect 18955 -4265 18995 -4260
rect 18955 -4295 18960 -4265
rect 18990 -4295 18995 -4265
rect 18955 -4300 18995 -4295
rect 19280 -4265 19320 -4260
rect 19280 -4295 19285 -4265
rect 19315 -4295 19320 -4265
rect 19280 -4300 19320 -4295
rect 16900 -4315 16950 -4305
rect 16900 -4345 16910 -4315
rect 16940 -4345 16950 -4315
rect 16900 -4355 16950 -4345
rect 18650 -4315 18700 -4305
rect 18650 -4345 18660 -4315
rect 18690 -4345 18700 -4315
rect 18650 -4355 18700 -4345
rect 19620 -4355 19640 -3829
rect 19840 -4310 19860 -90
rect 19830 -4315 19870 -4310
rect 19830 -4345 19835 -4315
rect 19865 -4345 19870 -4315
rect 19830 -4350 19870 -4345
rect 15950 -4360 15990 -4355
rect 15950 -4390 15955 -4360
rect 15985 -4390 15990 -4360
rect 15950 -4395 15990 -4390
rect 16205 -4360 16245 -4355
rect 16205 -4390 16210 -4360
rect 16240 -4390 16245 -4360
rect 16205 -4395 16245 -4390
rect 19355 -4360 19395 -4355
rect 19355 -4390 19360 -4360
rect 19390 -4390 19395 -4360
rect 19355 -4395 19395 -4390
rect 19610 -4360 19650 -4355
rect 19610 -4390 19615 -4360
rect 19645 -4390 19650 -4360
rect 19610 -4395 19650 -4390
rect 17955 -4410 17995 -4405
rect 17955 -4440 17960 -4410
rect 17990 -4440 17995 -4410
rect 17955 -4445 17995 -4440
<< via1 >>
rect 15730 -85 15760 -55
rect 15895 1280 15925 1310
rect 15950 145 15980 175
rect 15895 -1385 15925 -1355
rect 15790 -1800 15820 -1770
rect 16035 -1745 16065 -1715
rect 16490 1610 16520 1615
rect 16490 1590 16495 1610
rect 16495 1590 16515 1610
rect 16515 1590 16520 1610
rect 16490 1585 16520 1590
rect 16370 1530 16400 1560
rect 16370 1490 16400 1520
rect 16370 1475 16400 1480
rect 16370 1455 16375 1475
rect 16375 1455 16395 1475
rect 16395 1455 16400 1475
rect 16370 1450 16400 1455
rect 16490 1530 16520 1560
rect 16490 1490 16520 1520
rect 16490 1475 16520 1480
rect 16490 1455 16495 1475
rect 16495 1455 16515 1475
rect 16515 1455 16520 1475
rect 16490 1450 16520 1455
rect 16610 1530 16640 1560
rect 16610 1490 16640 1520
rect 16610 1475 16640 1480
rect 16610 1455 16615 1475
rect 16615 1455 16635 1475
rect 16635 1455 16640 1475
rect 16610 1450 16640 1455
rect 16890 1530 16920 1560
rect 16890 1490 16920 1520
rect 17055 1585 17085 1615
rect 17000 1530 17030 1560
rect 17000 1490 17030 1520
rect 16890 1475 16920 1480
rect 16890 1455 16895 1475
rect 16895 1455 16915 1475
rect 16915 1455 16920 1475
rect 16890 1450 16920 1455
rect 17000 1475 17030 1480
rect 17000 1455 17005 1475
rect 17005 1455 17025 1475
rect 17025 1455 17030 1475
rect 17000 1450 17030 1455
rect 17110 1530 17140 1560
rect 17110 1490 17140 1520
rect 17110 1475 17140 1480
rect 17110 1455 17115 1475
rect 17115 1455 17135 1475
rect 17135 1455 17140 1475
rect 17110 1450 17140 1455
rect 17220 1530 17250 1560
rect 17220 1490 17250 1520
rect 17220 1475 17250 1480
rect 17220 1455 17225 1475
rect 17225 1455 17245 1475
rect 17245 1455 17250 1475
rect 17220 1450 17250 1455
rect 17500 1530 17530 1560
rect 17500 1490 17530 1520
rect 17500 1475 17530 1480
rect 17500 1455 17505 1475
rect 17505 1455 17525 1475
rect 17525 1455 17530 1475
rect 17500 1450 17530 1455
rect 17565 1530 17595 1560
rect 17565 1490 17595 1520
rect 17565 1475 17595 1480
rect 17565 1455 17570 1475
rect 17570 1455 17590 1475
rect 17590 1455 17595 1475
rect 17565 1450 17595 1455
rect 17675 1530 17705 1560
rect 17675 1490 17705 1520
rect 17675 1475 17705 1480
rect 17675 1455 17680 1475
rect 17680 1455 17700 1475
rect 17700 1455 17705 1475
rect 17675 1450 17705 1455
rect 17785 1610 17815 1615
rect 17785 1590 17790 1610
rect 17790 1590 17810 1610
rect 17810 1590 17815 1610
rect 17785 1585 17815 1590
rect 17785 1530 17815 1560
rect 17785 1490 17815 1520
rect 17785 1475 17815 1480
rect 17785 1455 17790 1475
rect 17790 1455 17810 1475
rect 17810 1455 17815 1475
rect 17785 1450 17815 1455
rect 17895 1530 17925 1560
rect 17895 1490 17925 1520
rect 17895 1475 17925 1480
rect 17895 1455 17900 1475
rect 17900 1455 17920 1475
rect 17920 1455 17925 1475
rect 17895 1450 17925 1455
rect 18515 1585 18545 1615
rect 18005 1530 18035 1560
rect 18005 1490 18035 1520
rect 18005 1475 18035 1480
rect 18005 1455 18010 1475
rect 18010 1455 18030 1475
rect 18030 1455 18035 1475
rect 18005 1450 18035 1455
rect 18070 1530 18100 1560
rect 18070 1490 18100 1520
rect 18070 1475 18100 1480
rect 18070 1455 18075 1475
rect 18075 1455 18095 1475
rect 18095 1455 18100 1475
rect 18070 1450 18100 1455
rect 18350 1530 18380 1560
rect 18350 1490 18380 1520
rect 18350 1475 18380 1480
rect 18350 1455 18355 1475
rect 18355 1455 18375 1475
rect 18375 1455 18380 1475
rect 18350 1450 18380 1455
rect 18460 1530 18490 1560
rect 18460 1490 18490 1520
rect 18570 1530 18600 1560
rect 18570 1490 18600 1520
rect 18460 1475 18490 1480
rect 18460 1455 18465 1475
rect 18465 1455 18485 1475
rect 18485 1455 18490 1475
rect 18460 1450 18490 1455
rect 18680 1530 18710 1560
rect 18680 1490 18710 1520
rect 18570 1475 18600 1480
rect 18570 1455 18575 1475
rect 18575 1455 18595 1475
rect 18595 1455 18600 1475
rect 18570 1450 18600 1455
rect 18680 1475 18710 1480
rect 18680 1455 18685 1475
rect 18685 1455 18705 1475
rect 18705 1455 18710 1475
rect 18680 1450 18710 1455
rect 16435 1305 16465 1310
rect 16435 1285 16440 1305
rect 16440 1285 16460 1305
rect 16460 1285 16465 1305
rect 16435 1280 16465 1285
rect 16545 1305 16575 1310
rect 16545 1285 16550 1305
rect 16550 1285 16570 1305
rect 16570 1285 16575 1305
rect 16545 1280 16575 1285
rect 16945 1305 16975 1310
rect 16945 1285 16950 1305
rect 16950 1285 16970 1305
rect 16970 1285 16975 1305
rect 16945 1280 16975 1285
rect 17055 1305 17085 1310
rect 17055 1285 17060 1305
rect 17060 1285 17080 1305
rect 17080 1285 17085 1305
rect 17055 1280 17085 1285
rect 17165 1305 17195 1310
rect 17165 1285 17170 1305
rect 17170 1285 17190 1305
rect 17190 1285 17195 1305
rect 17165 1280 17195 1285
rect 17620 1305 17650 1310
rect 17620 1285 17625 1305
rect 17625 1285 17645 1305
rect 17645 1285 17650 1305
rect 17620 1280 17650 1285
rect 17730 1305 17760 1310
rect 17730 1285 17735 1305
rect 17735 1285 17755 1305
rect 17755 1285 17760 1305
rect 17730 1280 17760 1285
rect 17840 1305 17870 1310
rect 17840 1285 17845 1305
rect 17845 1285 17865 1305
rect 17865 1285 17870 1305
rect 17840 1280 17870 1285
rect 17950 1305 17980 1310
rect 17950 1285 17955 1305
rect 17955 1285 17975 1305
rect 17975 1285 17980 1305
rect 17950 1280 17980 1285
rect 18405 1305 18435 1310
rect 18405 1285 18410 1305
rect 18410 1285 18430 1305
rect 18430 1285 18435 1305
rect 18405 1280 18435 1285
rect 18515 1305 18545 1310
rect 18515 1285 18520 1305
rect 18520 1285 18540 1305
rect 18540 1285 18545 1305
rect 18515 1280 18545 1285
rect 18625 1305 18655 1310
rect 18625 1285 18630 1305
rect 18630 1285 18650 1305
rect 18650 1285 18655 1305
rect 18625 1280 18655 1285
rect 16545 1180 16575 1210
rect 16440 1065 16470 1095
rect 16440 1025 16470 1055
rect 16440 985 16470 1015
rect 16660 1065 16690 1095
rect 16660 1025 16690 1055
rect 16660 985 16690 1015
rect 16975 1065 17005 1095
rect 16975 1025 17005 1055
rect 16975 1010 17005 1015
rect 16975 990 16980 1010
rect 16980 990 17000 1010
rect 17000 990 17005 1010
rect 16975 985 17005 990
rect 17155 1065 17185 1095
rect 17155 1025 17185 1055
rect 17155 1010 17185 1015
rect 17155 990 17160 1010
rect 17160 990 17180 1010
rect 17180 990 17185 1010
rect 17155 985 17185 990
rect 17335 1065 17365 1095
rect 17335 1025 17365 1055
rect 17335 1010 17365 1015
rect 17335 990 17340 1010
rect 17340 990 17360 1010
rect 17360 990 17365 1010
rect 17335 985 17365 990
rect 17515 1065 17545 1095
rect 17515 1025 17545 1055
rect 17515 1010 17545 1015
rect 17515 990 17520 1010
rect 17520 990 17540 1010
rect 17540 990 17545 1010
rect 17515 985 17545 990
rect 17695 1065 17725 1095
rect 17695 1025 17725 1055
rect 17695 1010 17725 1015
rect 17695 990 17700 1010
rect 17700 990 17720 1010
rect 17720 990 17725 1010
rect 17695 985 17725 990
rect 17875 1065 17905 1095
rect 17875 1025 17905 1055
rect 17875 1010 17905 1015
rect 17875 990 17880 1010
rect 17880 990 17900 1010
rect 17900 990 17905 1010
rect 17875 985 17905 990
rect 18055 1065 18085 1095
rect 18055 1025 18085 1055
rect 18055 1010 18085 1015
rect 18055 990 18060 1010
rect 18060 990 18080 1010
rect 18080 990 18085 1010
rect 18055 985 18085 990
rect 18235 1065 18265 1095
rect 18235 1025 18265 1055
rect 18235 1010 18265 1015
rect 18235 990 18240 1010
rect 18240 990 18260 1010
rect 18260 990 18265 1010
rect 18235 985 18265 990
rect 18415 1065 18445 1095
rect 18415 1025 18445 1055
rect 18415 1010 18445 1015
rect 18415 990 18420 1010
rect 18420 990 18440 1010
rect 18440 990 18445 1010
rect 18415 985 18445 990
rect 18595 1065 18625 1095
rect 18595 1025 18625 1055
rect 18595 1010 18625 1015
rect 18595 990 18600 1010
rect 18600 990 18620 1010
rect 18620 990 18625 1010
rect 18595 985 18625 990
rect 18910 1065 18940 1095
rect 18910 1025 18940 1055
rect 18910 1010 18940 1015
rect 18910 990 18915 1010
rect 18915 990 18935 1010
rect 18935 990 18940 1010
rect 18910 985 18940 990
rect 19020 1065 19050 1095
rect 19020 1025 19050 1055
rect 19020 1010 19050 1015
rect 19020 990 19025 1010
rect 19025 990 19045 1010
rect 19045 990 19050 1010
rect 19020 985 19050 990
rect 19080 1065 19110 1095
rect 19080 1025 19110 1055
rect 19080 1010 19110 1015
rect 19080 990 19085 1010
rect 19085 990 19105 1010
rect 19105 990 19110 1010
rect 19080 985 19110 990
rect 16550 910 16580 915
rect 16550 890 16555 910
rect 16555 890 16575 910
rect 16575 890 16580 910
rect 16550 885 16580 890
rect 16785 885 16815 915
rect 16485 740 16515 745
rect 16485 720 16490 740
rect 16490 720 16510 740
rect 16510 720 16515 740
rect 16485 715 16515 720
rect 16615 740 16645 745
rect 16615 720 16620 740
rect 16620 720 16640 740
rect 16640 720 16645 740
rect 16615 715 16645 720
rect 16320 615 16350 645
rect 16265 560 16295 590
rect 16210 505 16240 535
rect 16265 -140 16295 -110
rect 16210 -1215 16240 -1185
rect 16110 -1895 16140 -1865
rect 16160 -1980 16190 -1950
rect 16425 360 16455 390
rect 16425 320 16455 350
rect 16425 280 16455 310
rect 19330 1180 19360 1210
rect 18955 740 18985 745
rect 18955 720 18960 740
rect 18960 720 18980 740
rect 18980 720 18985 740
rect 18955 715 18985 720
rect 19265 715 19295 745
rect 19005 680 19035 685
rect 19005 660 19010 680
rect 19010 660 19030 680
rect 19030 660 19035 680
rect 19005 655 19035 660
rect 17605 640 17635 645
rect 17605 620 17610 640
rect 17610 620 17630 640
rect 17630 620 17635 640
rect 17605 615 17635 620
rect 17965 640 17995 645
rect 17965 620 17970 640
rect 17970 620 17990 640
rect 17990 620 17995 640
rect 17965 615 17995 620
rect 16785 560 16815 590
rect 16550 505 16580 535
rect 17425 560 17455 590
rect 17245 505 17275 535
rect 17065 460 17095 490
rect 16545 360 16575 390
rect 16545 320 16575 350
rect 16545 280 16575 310
rect 16665 360 16695 390
rect 16665 320 16695 350
rect 16665 280 16695 310
rect 16785 360 16815 390
rect 16785 320 16815 350
rect 16785 280 16815 310
rect 16905 360 16935 390
rect 16905 320 16935 350
rect 16905 280 16935 310
rect 17025 360 17055 390
rect 17025 320 17055 350
rect 17025 280 17055 310
rect 17145 360 17175 390
rect 17145 320 17175 350
rect 17145 280 17175 310
rect 17265 360 17295 390
rect 17265 320 17295 350
rect 17265 280 17295 310
rect 17385 360 17415 390
rect 17385 320 17415 350
rect 17385 280 17415 310
rect 17505 360 17535 390
rect 17505 320 17535 350
rect 17505 280 17535 310
rect 17625 360 17655 390
rect 17625 320 17655 350
rect 17625 280 17655 310
rect 18145 560 18175 590
rect 18325 505 18355 535
rect 17785 460 17815 490
rect 18505 460 18535 490
rect 17945 360 17975 390
rect 17945 320 17975 350
rect 17945 280 17975 310
rect 18065 360 18095 390
rect 18065 320 18095 350
rect 18065 280 18095 310
rect 18185 360 18215 390
rect 18185 320 18215 350
rect 18185 280 18215 310
rect 18305 360 18335 390
rect 18305 320 18335 350
rect 18305 280 18335 310
rect 18425 360 18455 390
rect 18425 320 18455 350
rect 18425 280 18455 310
rect 18545 360 18575 390
rect 18545 320 18575 350
rect 18545 280 18575 310
rect 18665 360 18695 390
rect 18665 320 18695 350
rect 18665 280 18695 310
rect 18785 360 18815 390
rect 18785 320 18815 350
rect 18785 280 18815 310
rect 18905 360 18935 390
rect 18905 320 18935 350
rect 18905 280 18935 310
rect 19025 360 19055 390
rect 19025 320 19055 350
rect 19025 280 19055 310
rect 19145 360 19175 390
rect 19145 320 19175 350
rect 19145 280 19175 310
rect 16485 170 16515 175
rect 16485 150 16490 170
rect 16490 150 16510 170
rect 16510 150 16515 170
rect 16485 145 16515 150
rect 16845 170 16875 175
rect 16845 150 16850 170
rect 16850 150 16870 170
rect 16870 150 16875 170
rect 16845 145 16875 150
rect 17205 170 17235 175
rect 17205 150 17210 170
rect 17210 150 17230 170
rect 17230 150 17235 170
rect 17205 145 17235 150
rect 17565 170 17595 175
rect 17565 150 17570 170
rect 17570 150 17590 170
rect 17590 150 17595 170
rect 17565 145 17595 150
rect 17695 145 17725 175
rect 17875 145 17905 175
rect 16605 0 16635 5
rect 16605 -20 16610 0
rect 16610 -20 16630 0
rect 16630 -20 16635 0
rect 16605 -25 16635 -20
rect 16965 0 16995 5
rect 16965 -20 16970 0
rect 16970 -20 16990 0
rect 16990 -20 16995 0
rect 16965 -25 16995 -20
rect 17325 0 17355 5
rect 17325 -20 17330 0
rect 17330 -20 17350 0
rect 17350 -20 17355 0
rect 17325 -25 17355 -20
rect 16515 -85 16545 -55
rect 16725 -85 16755 -55
rect 16845 -85 16875 -55
rect 17085 -85 17115 -55
rect 17205 -85 17235 -55
rect 17445 -85 17475 -55
rect 17535 -85 17565 -55
rect 17007 -115 17037 -110
rect 17007 -135 17012 -115
rect 17012 -135 17032 -115
rect 17032 -135 17037 -115
rect 17007 -140 17037 -135
rect 16320 -460 16350 -430
rect 17565 -175 17595 -170
rect 17565 -195 17570 -175
rect 17570 -195 17590 -175
rect 17590 -195 17595 -175
rect 17565 -200 17595 -195
rect 17565 -215 17595 -210
rect 17565 -235 17570 -215
rect 17570 -235 17590 -215
rect 17590 -235 17595 -215
rect 17565 -240 17595 -235
rect 17565 -255 17595 -250
rect 17565 -275 17570 -255
rect 17570 -275 17590 -255
rect 17590 -275 17595 -255
rect 17565 -280 17595 -275
rect 17075 -435 17105 -430
rect 17075 -455 17080 -435
rect 17080 -455 17100 -435
rect 17100 -455 17105 -435
rect 17075 -460 17105 -455
rect 16535 -540 16565 -510
rect 17025 -540 17055 -510
rect 16625 -595 16655 -565
rect 16625 -635 16655 -605
rect 16625 -650 16655 -645
rect 16625 -670 16630 -650
rect 16630 -670 16650 -650
rect 16650 -670 16655 -650
rect 16625 -675 16655 -670
rect 16745 -595 16775 -565
rect 16745 -635 16775 -605
rect 16745 -650 16775 -645
rect 16745 -670 16750 -650
rect 16750 -670 16770 -650
rect 16770 -670 16775 -650
rect 16745 -675 16775 -670
rect 16865 -595 16895 -565
rect 16865 -635 16895 -605
rect 16865 -650 16895 -645
rect 16865 -670 16870 -650
rect 16870 -670 16890 -650
rect 16890 -670 16895 -650
rect 16865 -675 16895 -670
rect 16985 -595 17015 -565
rect 16985 -635 17015 -605
rect 16985 -650 17015 -645
rect 16985 -670 16990 -650
rect 16990 -670 17010 -650
rect 17010 -670 17015 -650
rect 16985 -675 17015 -670
rect 17305 -595 17335 -565
rect 17305 -635 17335 -605
rect 17305 -650 17335 -645
rect 17305 -670 17310 -650
rect 17310 -670 17330 -650
rect 17330 -670 17335 -650
rect 17305 -675 17335 -670
rect 17425 -595 17455 -565
rect 17425 -635 17455 -605
rect 17425 -650 17455 -645
rect 17425 -670 17430 -650
rect 17430 -670 17450 -650
rect 17450 -670 17455 -650
rect 17425 -675 17455 -670
rect 17545 -595 17575 -565
rect 17545 -635 17575 -605
rect 17545 -650 17575 -645
rect 17545 -670 17550 -650
rect 17550 -670 17570 -650
rect 17570 -670 17575 -650
rect 17545 -675 17575 -670
rect 17745 -200 17775 -170
rect 17785 -200 17815 -170
rect 17825 -200 17855 -170
rect 17745 -240 17775 -210
rect 17785 -240 17815 -210
rect 17825 -240 17855 -210
rect 17745 -280 17775 -250
rect 17785 -280 17815 -250
rect 17825 -280 17855 -250
rect 17115 -970 17145 -965
rect 17115 -990 17120 -970
rect 17120 -990 17140 -970
rect 17140 -990 17145 -970
rect 17115 -995 17145 -990
rect 17115 -1035 17145 -1005
rect 17115 -1075 17145 -1045
rect 18005 170 18035 175
rect 18005 150 18010 170
rect 18010 150 18030 170
rect 18030 150 18035 170
rect 18005 145 18035 150
rect 18365 170 18395 175
rect 18365 150 18370 170
rect 18370 150 18390 170
rect 18390 150 18395 170
rect 18365 145 18395 150
rect 18725 170 18755 175
rect 18725 150 18730 170
rect 18730 150 18750 170
rect 18750 150 18755 170
rect 18725 145 18755 150
rect 19085 170 19115 175
rect 19085 150 19090 170
rect 19090 150 19110 170
rect 19110 150 19115 170
rect 19085 145 19115 150
rect 18245 0 18275 5
rect 18245 -20 18250 0
rect 18250 -20 18270 0
rect 18270 -20 18275 0
rect 18245 -25 18275 -20
rect 18605 0 18635 5
rect 18605 -20 18610 0
rect 18610 -20 18630 0
rect 18630 -20 18635 0
rect 18605 -25 18635 -20
rect 18965 0 18995 5
rect 18965 -20 18970 0
rect 18970 -20 18990 0
rect 18990 -20 18995 0
rect 18965 -25 18995 -20
rect 18035 -85 18065 -55
rect 18125 -85 18155 -55
rect 18365 -85 18395 -55
rect 18485 -85 18515 -55
rect 18725 -85 18755 -55
rect 18845 -85 18875 -55
rect 19055 -85 19085 -55
rect 18563 -115 18593 -110
rect 18563 -135 18568 -115
rect 18568 -135 18588 -115
rect 18588 -135 18593 -115
rect 18563 -140 18593 -135
rect 18005 -175 18035 -170
rect 18005 -195 18010 -175
rect 18010 -195 18030 -175
rect 18030 -195 18035 -175
rect 18005 -200 18035 -195
rect 18005 -215 18035 -210
rect 18005 -235 18010 -215
rect 18010 -235 18030 -215
rect 18030 -235 18035 -215
rect 18005 -240 18035 -235
rect 18005 -255 18035 -250
rect 18005 -275 18010 -255
rect 18010 -275 18030 -255
rect 18030 -275 18035 -255
rect 18005 -280 18035 -275
rect 19410 460 19440 490
rect 19410 -140 19440 -110
rect 18495 -435 18525 -430
rect 18495 -455 18500 -435
rect 18500 -455 18520 -435
rect 18520 -455 18525 -435
rect 18495 -460 18525 -455
rect 19330 -460 19360 -430
rect 18545 -540 18575 -510
rect 19035 -540 19065 -510
rect 18025 -595 18055 -565
rect 18025 -635 18055 -605
rect 18025 -650 18055 -645
rect 18025 -670 18030 -650
rect 18030 -670 18050 -650
rect 18050 -670 18055 -650
rect 18025 -675 18055 -670
rect 18145 -595 18175 -565
rect 18145 -635 18175 -605
rect 18145 -650 18175 -645
rect 18145 -670 18150 -650
rect 18150 -670 18170 -650
rect 18170 -670 18175 -650
rect 18145 -675 18175 -670
rect 18265 -595 18295 -565
rect 18265 -635 18295 -605
rect 18265 -650 18295 -645
rect 18265 -670 18270 -650
rect 18270 -670 18290 -650
rect 18290 -670 18295 -650
rect 18265 -675 18295 -670
rect 18585 -595 18615 -565
rect 18585 -635 18615 -605
rect 18585 -650 18615 -645
rect 18585 -670 18590 -650
rect 18590 -670 18610 -650
rect 18610 -670 18615 -650
rect 18585 -675 18615 -670
rect 18705 -595 18735 -565
rect 18705 -635 18735 -605
rect 18705 -650 18735 -645
rect 18705 -670 18710 -650
rect 18710 -670 18730 -650
rect 18730 -670 18735 -650
rect 18705 -675 18735 -670
rect 18825 -595 18855 -565
rect 18825 -635 18855 -605
rect 18825 -650 18855 -645
rect 18825 -670 18830 -650
rect 18830 -670 18850 -650
rect 18850 -670 18855 -650
rect 18825 -675 18855 -670
rect 18945 -595 18975 -565
rect 18945 -635 18975 -605
rect 18945 -650 18975 -645
rect 18945 -670 18950 -650
rect 18950 -670 18970 -650
rect 18970 -670 18975 -650
rect 18945 -675 18975 -670
rect 17745 -995 17775 -965
rect 17785 -995 17815 -965
rect 17825 -995 17855 -965
rect 17745 -1035 17775 -1005
rect 17785 -1035 17815 -1005
rect 17825 -1035 17855 -1005
rect 17745 -1075 17775 -1045
rect 17785 -1075 17815 -1045
rect 17825 -1075 17855 -1045
rect 18455 -970 18485 -965
rect 18455 -990 18460 -970
rect 18460 -990 18480 -970
rect 18480 -990 18485 -970
rect 18455 -995 18485 -990
rect 18455 -1035 18485 -1005
rect 18455 -1075 18485 -1045
rect 16745 -1105 16775 -1100
rect 16745 -1125 16750 -1105
rect 16750 -1125 16770 -1105
rect 16770 -1125 16775 -1105
rect 16745 -1130 16775 -1125
rect 16825 -1105 16855 -1100
rect 16825 -1125 16830 -1105
rect 16830 -1125 16850 -1105
rect 16850 -1125 16855 -1105
rect 16825 -1130 16855 -1125
rect 16905 -1105 16935 -1100
rect 16905 -1125 16910 -1105
rect 16910 -1125 16930 -1105
rect 16930 -1125 16935 -1105
rect 16905 -1130 16935 -1125
rect 16985 -1105 17015 -1100
rect 16985 -1125 16990 -1105
rect 16990 -1125 17010 -1105
rect 17010 -1125 17015 -1105
rect 16985 -1130 17015 -1125
rect 17065 -1105 17095 -1100
rect 17065 -1125 17070 -1105
rect 17070 -1125 17090 -1105
rect 17090 -1125 17095 -1105
rect 17065 -1130 17095 -1125
rect 17145 -1105 17175 -1100
rect 17145 -1125 17150 -1105
rect 17150 -1125 17170 -1105
rect 17170 -1125 17175 -1105
rect 17145 -1130 17175 -1125
rect 17225 -1105 17255 -1100
rect 17225 -1125 17230 -1105
rect 17230 -1125 17250 -1105
rect 17250 -1125 17255 -1105
rect 17225 -1130 17255 -1125
rect 17305 -1105 17335 -1100
rect 17305 -1125 17310 -1105
rect 17310 -1125 17330 -1105
rect 17330 -1125 17335 -1105
rect 17305 -1130 17335 -1125
rect 17385 -1105 17415 -1100
rect 17385 -1125 17390 -1105
rect 17390 -1125 17410 -1105
rect 17410 -1125 17415 -1105
rect 17385 -1130 17415 -1125
rect 17465 -1105 17495 -1100
rect 17465 -1125 17470 -1105
rect 17470 -1125 17490 -1105
rect 17490 -1125 17495 -1105
rect 17465 -1130 17495 -1125
rect 17545 -1105 17575 -1100
rect 17545 -1125 17550 -1105
rect 17550 -1125 17570 -1105
rect 17570 -1125 17575 -1105
rect 17545 -1130 17575 -1125
rect 17625 -1105 17655 -1100
rect 17625 -1125 17630 -1105
rect 17630 -1125 17650 -1105
rect 17650 -1125 17655 -1105
rect 17625 -1130 17655 -1125
rect 17705 -1105 17735 -1100
rect 17705 -1125 17710 -1105
rect 17710 -1125 17730 -1105
rect 17730 -1125 17735 -1105
rect 17705 -1130 17735 -1125
rect 17785 -1105 17815 -1100
rect 17785 -1125 17790 -1105
rect 17790 -1125 17810 -1105
rect 17810 -1125 17815 -1105
rect 17785 -1130 17815 -1125
rect 17865 -1105 17895 -1100
rect 17865 -1125 17870 -1105
rect 17870 -1125 17890 -1105
rect 17890 -1125 17895 -1105
rect 17865 -1130 17895 -1125
rect 17945 -1105 17975 -1100
rect 17945 -1125 17950 -1105
rect 17950 -1125 17970 -1105
rect 17970 -1125 17975 -1105
rect 17945 -1130 17975 -1125
rect 18025 -1105 18055 -1100
rect 18025 -1125 18030 -1105
rect 18030 -1125 18050 -1105
rect 18050 -1125 18055 -1105
rect 18025 -1130 18055 -1125
rect 18105 -1105 18135 -1100
rect 18105 -1125 18110 -1105
rect 18110 -1125 18130 -1105
rect 18130 -1125 18135 -1105
rect 18105 -1130 18135 -1125
rect 18185 -1105 18215 -1100
rect 18185 -1125 18190 -1105
rect 18190 -1125 18210 -1105
rect 18210 -1125 18215 -1105
rect 18185 -1130 18215 -1125
rect 18265 -1105 18295 -1100
rect 18265 -1125 18270 -1105
rect 18270 -1125 18290 -1105
rect 18290 -1125 18295 -1105
rect 18265 -1130 18295 -1125
rect 18345 -1105 18375 -1100
rect 18345 -1125 18350 -1105
rect 18350 -1125 18370 -1105
rect 18370 -1125 18375 -1105
rect 18345 -1130 18375 -1125
rect 18425 -1105 18455 -1100
rect 18425 -1125 18430 -1105
rect 18430 -1125 18450 -1105
rect 18450 -1125 18455 -1105
rect 18425 -1130 18455 -1125
rect 18505 -1105 18535 -1100
rect 18505 -1125 18510 -1105
rect 18510 -1125 18530 -1105
rect 18530 -1125 18535 -1105
rect 18505 -1130 18535 -1125
rect 18585 -1105 18615 -1100
rect 18585 -1125 18590 -1105
rect 18590 -1125 18610 -1105
rect 18610 -1125 18615 -1105
rect 18585 -1130 18615 -1125
rect 18665 -1105 18695 -1100
rect 18665 -1125 18670 -1105
rect 18670 -1125 18690 -1105
rect 18690 -1125 18695 -1105
rect 18665 -1130 18695 -1125
rect 18745 -1105 18775 -1100
rect 18745 -1125 18750 -1105
rect 18750 -1125 18770 -1105
rect 18770 -1125 18775 -1105
rect 18745 -1130 18775 -1125
rect 16705 -1190 16735 -1185
rect 16705 -1210 16710 -1190
rect 16710 -1210 16730 -1190
rect 16730 -1210 16735 -1190
rect 16705 -1215 16735 -1210
rect 18900 -1170 18930 -1165
rect 18900 -1190 18905 -1170
rect 18905 -1190 18925 -1170
rect 18925 -1190 18930 -1170
rect 18900 -1195 18930 -1190
rect 18900 -1210 18930 -1205
rect 18900 -1230 18905 -1210
rect 18905 -1230 18925 -1210
rect 18925 -1230 18930 -1210
rect 18900 -1235 18930 -1230
rect 16660 -1385 16690 -1355
rect 16770 -1385 16800 -1355
rect 17305 -1385 17335 -1355
rect 17785 -1385 17815 -1355
rect 18265 -1385 18295 -1355
rect 16605 -1440 16635 -1410
rect 16605 -1480 16635 -1450
rect 16605 -1495 16635 -1490
rect 16605 -1515 16610 -1495
rect 16610 -1515 16630 -1495
rect 16630 -1515 16635 -1495
rect 16605 -1520 16635 -1515
rect 16715 -1440 16745 -1410
rect 16715 -1480 16745 -1450
rect 16715 -1495 16745 -1490
rect 16715 -1515 16720 -1495
rect 16720 -1515 16740 -1495
rect 16740 -1515 16745 -1495
rect 16715 -1520 16745 -1515
rect 16825 -1440 16855 -1410
rect 16825 -1480 16855 -1450
rect 16825 -1495 16855 -1490
rect 16825 -1515 16830 -1495
rect 16830 -1515 16850 -1495
rect 16850 -1515 16855 -1495
rect 16825 -1520 16855 -1515
rect 16885 -1440 16915 -1410
rect 16885 -1480 16915 -1450
rect 16885 -1495 16915 -1490
rect 16885 -1515 16890 -1495
rect 16890 -1515 16910 -1495
rect 16910 -1515 16915 -1495
rect 16885 -1520 16915 -1515
rect 17030 -1440 17060 -1410
rect 17030 -1480 17060 -1450
rect 17030 -1495 17060 -1490
rect 17030 -1515 17035 -1495
rect 17035 -1515 17055 -1495
rect 17055 -1515 17060 -1495
rect 17030 -1520 17060 -1515
rect 17140 -1440 17170 -1410
rect 17140 -1480 17170 -1450
rect 17140 -1495 17170 -1490
rect 17140 -1515 17145 -1495
rect 17145 -1515 17165 -1495
rect 17165 -1515 17170 -1495
rect 17140 -1520 17170 -1515
rect 17250 -1440 17280 -1410
rect 17250 -1480 17280 -1450
rect 17250 -1495 17280 -1490
rect 17250 -1515 17255 -1495
rect 17255 -1515 17275 -1495
rect 17275 -1515 17280 -1495
rect 17250 -1520 17280 -1515
rect 17360 -1440 17390 -1410
rect 17360 -1480 17390 -1450
rect 17360 -1495 17390 -1490
rect 17360 -1515 17365 -1495
rect 17365 -1515 17385 -1495
rect 17385 -1515 17390 -1495
rect 17360 -1520 17390 -1515
rect 17470 -1440 17500 -1410
rect 17470 -1480 17500 -1450
rect 17470 -1495 17500 -1490
rect 17470 -1515 17475 -1495
rect 17475 -1515 17495 -1495
rect 17495 -1515 17500 -1495
rect 17470 -1520 17500 -1515
rect 17620 -1440 17650 -1410
rect 17620 -1480 17650 -1450
rect 17620 -1495 17650 -1490
rect 17620 -1515 17625 -1495
rect 17625 -1515 17645 -1495
rect 17645 -1515 17650 -1495
rect 17620 -1520 17650 -1515
rect 17730 -1440 17760 -1410
rect 17730 -1480 17760 -1450
rect 17730 -1495 17760 -1490
rect 17730 -1515 17735 -1495
rect 17735 -1515 17755 -1495
rect 17755 -1515 17760 -1495
rect 17730 -1520 17760 -1515
rect 17840 -1440 17870 -1410
rect 17840 -1480 17870 -1450
rect 17840 -1495 17870 -1490
rect 17840 -1515 17845 -1495
rect 17845 -1515 17865 -1495
rect 17865 -1515 17870 -1495
rect 17840 -1520 17870 -1515
rect 17950 -1440 17980 -1410
rect 17950 -1480 17980 -1450
rect 17950 -1495 17980 -1490
rect 17950 -1515 17955 -1495
rect 17955 -1515 17975 -1495
rect 17975 -1515 17980 -1495
rect 17950 -1520 17980 -1515
rect 18100 -1440 18130 -1410
rect 18100 -1480 18130 -1450
rect 18100 -1495 18130 -1490
rect 18100 -1515 18105 -1495
rect 18105 -1515 18125 -1495
rect 18125 -1515 18130 -1495
rect 18100 -1520 18130 -1515
rect 18210 -1440 18240 -1410
rect 18210 -1480 18240 -1450
rect 18210 -1495 18240 -1490
rect 18210 -1515 18215 -1495
rect 18215 -1515 18235 -1495
rect 18235 -1515 18240 -1495
rect 18210 -1520 18240 -1515
rect 18320 -1440 18350 -1410
rect 18320 -1480 18350 -1450
rect 18320 -1495 18350 -1490
rect 18320 -1515 18325 -1495
rect 18325 -1515 18345 -1495
rect 18345 -1515 18350 -1495
rect 18320 -1520 18350 -1515
rect 18430 -1440 18460 -1410
rect 18430 -1480 18460 -1450
rect 18430 -1495 18460 -1490
rect 18430 -1515 18435 -1495
rect 18435 -1515 18455 -1495
rect 18455 -1515 18460 -1495
rect 18430 -1520 18460 -1515
rect 18540 -1440 18570 -1410
rect 18540 -1480 18570 -1450
rect 18540 -1495 18570 -1490
rect 18540 -1515 18545 -1495
rect 18545 -1515 18565 -1495
rect 18565 -1515 18570 -1495
rect 18540 -1520 18570 -1515
rect 17195 -1665 17225 -1660
rect 17195 -1685 17200 -1665
rect 17200 -1685 17220 -1665
rect 17220 -1685 17225 -1665
rect 17195 -1690 17225 -1685
rect 17085 -1745 17115 -1715
rect 17415 -1665 17445 -1660
rect 17415 -1685 17420 -1665
rect 17420 -1685 17440 -1665
rect 17440 -1685 17445 -1665
rect 17415 -1690 17445 -1685
rect 17675 -1665 17705 -1660
rect 17675 -1685 17680 -1665
rect 17680 -1685 17700 -1665
rect 17700 -1685 17705 -1665
rect 17675 -1690 17705 -1685
rect 17785 -1665 17815 -1660
rect 17785 -1685 17790 -1665
rect 17790 -1685 17810 -1665
rect 17810 -1685 17815 -1665
rect 17785 -1690 17815 -1685
rect 17895 -1665 17925 -1660
rect 17895 -1685 17900 -1665
rect 17900 -1685 17920 -1665
rect 17920 -1685 17925 -1665
rect 17895 -1690 17925 -1685
rect 18155 -1665 18185 -1660
rect 18155 -1685 18160 -1665
rect 18160 -1685 18180 -1665
rect 18180 -1685 18185 -1665
rect 18155 -1690 18185 -1685
rect 18375 -1665 18405 -1660
rect 18375 -1685 18380 -1665
rect 18380 -1685 18400 -1665
rect 18400 -1685 18405 -1665
rect 18375 -1690 18405 -1685
rect 17305 -1745 17335 -1715
rect 17195 -1800 17225 -1770
rect 16770 -1895 16800 -1865
rect 18265 -1745 18295 -1715
rect 18485 -1745 18515 -1715
rect 18375 -1800 18405 -1770
rect 17785 -1930 17815 -1900
rect 19330 -1980 19360 -1950
rect 16320 -2030 16350 -2000
rect 17430 -2005 17465 -2000
rect 17430 -2030 17435 -2005
rect 17435 -2030 17460 -2005
rect 17460 -2030 17465 -2005
rect 17430 -2035 17465 -2030
rect 18129 -2005 18164 -2000
rect 18129 -2030 18134 -2005
rect 18134 -2030 18159 -2005
rect 18159 -2030 18164 -2005
rect 18129 -2035 18164 -2030
rect 18835 -2035 18865 -2005
rect 17430 -2090 17460 -2060
rect 16265 -2130 16295 -2100
rect 16485 -2130 16515 -2100
rect 16485 -2905 16520 -2900
rect 16485 -2930 16490 -2905
rect 16490 -2930 16515 -2905
rect 16515 -2930 16520 -2905
rect 16485 -2935 16520 -2930
rect 16735 -2130 16765 -2100
rect 16160 -3030 16195 -3025
rect 16160 -3055 16165 -3030
rect 16165 -3055 16190 -3030
rect 16190 -3055 16195 -3030
rect 16160 -3060 16195 -3055
rect 15825 -3145 15855 -3115
rect 15950 -3121 15985 -3116
rect 15950 -3146 15955 -3121
rect 15955 -3146 15980 -3121
rect 15980 -3146 15985 -3121
rect 16735 -3135 16765 -3105
rect 15950 -3151 15985 -3146
rect 17785 -3135 17815 -3105
rect 18620 -3135 18650 -3105
rect 19085 -2090 19115 -2060
rect 19080 -2905 19115 -2900
rect 19080 -2930 19085 -2905
rect 19085 -2930 19110 -2905
rect 19110 -2930 19115 -2905
rect 19080 -2935 19115 -2930
rect 19615 1585 19645 1615
rect 19615 655 19645 685
rect 19615 145 19645 175
rect 19540 -1930 19570 -1900
rect 19405 -3002 19440 -2997
rect 19405 -3027 19410 -3002
rect 19410 -3027 19435 -3002
rect 19435 -3027 19440 -3002
rect 19405 -3032 19440 -3027
rect 18835 -3135 18865 -3105
rect 19835 -85 19865 -55
rect 19780 -1800 19810 -1770
rect 19610 -3120 19645 -3115
rect 19610 -3145 19615 -3120
rect 19615 -3145 19640 -3120
rect 19640 -3145 19645 -3120
rect 19610 -3150 19645 -3145
rect 15950 -3794 15985 -3789
rect 15950 -3819 15955 -3794
rect 15955 -3819 15980 -3794
rect 15980 -3819 15985 -3794
rect 15950 -3824 15985 -3819
rect 15825 -4295 15855 -4265
rect 15730 -4345 15760 -4315
rect 16280 -3899 16315 -3894
rect 16280 -3924 16285 -3899
rect 16285 -3924 16310 -3899
rect 16310 -3924 16315 -3899
rect 16280 -3929 16315 -3924
rect 16605 -3974 16640 -3969
rect 16605 -3999 16610 -3974
rect 16610 -3999 16635 -3974
rect 16635 -3999 16640 -3974
rect 19610 -3794 19645 -3789
rect 19610 -3819 19615 -3794
rect 19615 -3819 19640 -3794
rect 19640 -3819 19645 -3794
rect 19610 -3824 19645 -3819
rect 19285 -3899 19320 -3894
rect 19285 -3924 19290 -3899
rect 19290 -3924 19315 -3899
rect 19315 -3924 19320 -3899
rect 19285 -3929 19320 -3924
rect 18960 -3974 18995 -3969
rect 16605 -4004 16640 -3999
rect 18960 -3999 18965 -3974
rect 18965 -3999 18990 -3974
rect 18990 -3999 18995 -3974
rect 18960 -4004 18995 -3999
rect 16285 -4220 16315 -4190
rect 16610 -4220 16640 -4190
rect 17260 -4295 17290 -4265
rect 17785 -4270 17815 -4265
rect 17785 -4290 17790 -4270
rect 17790 -4290 17810 -4270
rect 17810 -4290 17815 -4270
rect 17785 -4295 17815 -4290
rect 18960 -4295 18990 -4265
rect 19285 -4295 19315 -4265
rect 16910 -4345 16940 -4315
rect 18660 -4345 18690 -4315
rect 19835 -4345 19865 -4315
rect 15955 -4390 15985 -4360
rect 16210 -4390 16240 -4360
rect 19360 -4390 19390 -4360
rect 19615 -4390 19645 -4360
rect 17960 -4440 17990 -4410
<< metal2 >>
rect 16485 1615 18500 1620
rect 18590 1615 19650 1620
rect 16485 1585 16490 1615
rect 16520 1585 17055 1615
rect 17085 1585 17785 1615
rect 17815 1585 18515 1615
rect 18545 1585 19615 1615
rect 19645 1585 19650 1615
rect 16485 1580 19650 1585
rect 16365 1560 18715 1565
rect 16365 1530 16370 1560
rect 16400 1530 16490 1560
rect 16520 1530 16610 1560
rect 16640 1530 16890 1560
rect 16920 1530 17000 1560
rect 17030 1530 17110 1560
rect 17140 1530 17220 1560
rect 17250 1530 17500 1560
rect 17530 1530 17565 1560
rect 17595 1530 17675 1560
rect 17705 1530 17785 1560
rect 17815 1530 17895 1560
rect 17925 1530 18005 1560
rect 18035 1530 18070 1560
rect 18100 1530 18350 1560
rect 18380 1530 18460 1560
rect 18490 1530 18570 1560
rect 18600 1530 18680 1560
rect 18710 1530 18715 1560
rect 16365 1520 18715 1530
rect 16365 1490 16370 1520
rect 16400 1490 16490 1520
rect 16520 1490 16610 1520
rect 16640 1490 16890 1520
rect 16920 1490 17000 1520
rect 17030 1490 17110 1520
rect 17140 1490 17220 1520
rect 17250 1490 17500 1520
rect 17530 1490 17565 1520
rect 17595 1490 17675 1520
rect 17705 1490 17785 1520
rect 17815 1490 17895 1520
rect 17925 1490 18005 1520
rect 18035 1490 18070 1520
rect 18100 1490 18350 1520
rect 18380 1490 18460 1520
rect 18490 1490 18570 1520
rect 18600 1490 18680 1520
rect 18710 1490 18715 1520
rect 16365 1480 18715 1490
rect 16365 1450 16370 1480
rect 16400 1450 16490 1480
rect 16520 1450 16610 1480
rect 16640 1450 16890 1480
rect 16920 1450 17000 1480
rect 17030 1450 17110 1480
rect 17140 1450 17220 1480
rect 17250 1450 17500 1480
rect 17530 1450 17565 1480
rect 17595 1450 17675 1480
rect 17705 1450 17785 1480
rect 17815 1450 17895 1480
rect 17925 1450 18005 1480
rect 18035 1450 18070 1480
rect 18100 1450 18350 1480
rect 18380 1450 18460 1480
rect 18490 1450 18570 1480
rect 18600 1450 18680 1480
rect 18710 1450 18715 1480
rect 16365 1445 18715 1450
rect 15890 1310 16470 1315
rect 15890 1280 15895 1310
rect 15925 1280 16435 1310
rect 16465 1280 16470 1310
rect 15890 1275 16470 1280
rect 16540 1310 16580 1315
rect 16540 1280 16545 1310
rect 16575 1280 16580 1310
rect 16540 1275 16580 1280
rect 16940 1310 16980 1315
rect 16940 1280 16945 1310
rect 16975 1305 16980 1310
rect 17050 1310 17090 1315
rect 17050 1305 17055 1310
rect 16975 1285 17055 1305
rect 16975 1280 16980 1285
rect 16940 1275 16980 1280
rect 17050 1280 17055 1285
rect 17085 1305 17090 1310
rect 17160 1310 17200 1315
rect 17160 1305 17165 1310
rect 17085 1285 17165 1305
rect 17085 1280 17090 1285
rect 17050 1275 17090 1280
rect 17160 1280 17165 1285
rect 17195 1280 17200 1310
rect 17160 1275 17200 1280
rect 17615 1310 17655 1315
rect 17615 1280 17620 1310
rect 17650 1305 17655 1310
rect 17725 1310 17765 1315
rect 17725 1305 17730 1310
rect 17650 1285 17730 1305
rect 17650 1280 17655 1285
rect 17615 1275 17655 1280
rect 17725 1280 17730 1285
rect 17760 1305 17765 1310
rect 17835 1310 17875 1315
rect 17835 1305 17840 1310
rect 17760 1285 17840 1305
rect 17760 1280 17765 1285
rect 17725 1275 17765 1280
rect 17835 1280 17840 1285
rect 17870 1305 17875 1310
rect 17945 1310 17985 1315
rect 17945 1305 17950 1310
rect 17870 1285 17950 1305
rect 17870 1280 17875 1285
rect 17835 1275 17875 1280
rect 17945 1280 17950 1285
rect 17980 1280 17985 1310
rect 17945 1275 17985 1280
rect 18400 1310 18440 1315
rect 18400 1280 18405 1310
rect 18435 1305 18440 1310
rect 18510 1310 18550 1315
rect 18510 1305 18515 1310
rect 18435 1285 18515 1305
rect 18435 1280 18440 1285
rect 18400 1275 18440 1280
rect 18510 1280 18515 1285
rect 18545 1305 18550 1310
rect 18620 1310 18660 1315
rect 18620 1305 18625 1310
rect 18545 1285 18625 1305
rect 18545 1280 18550 1285
rect 18510 1275 18550 1280
rect 18620 1280 18625 1285
rect 18655 1280 18660 1310
rect 18620 1275 18660 1280
rect 16540 1210 16580 1215
rect 16540 1180 16545 1210
rect 16575 1205 16580 1210
rect 19325 1210 19365 1215
rect 19325 1205 19330 1210
rect 16575 1185 19330 1205
rect 16575 1180 16580 1185
rect 16540 1175 16580 1180
rect 19325 1180 19330 1185
rect 19360 1180 19365 1210
rect 19325 1175 19365 1180
rect 16435 1095 18630 1100
rect 16435 1065 16440 1095
rect 16470 1065 16660 1095
rect 16690 1065 16975 1095
rect 17005 1065 17155 1095
rect 17185 1065 17335 1095
rect 17365 1065 17515 1095
rect 17545 1065 17695 1095
rect 17725 1065 17875 1095
rect 17905 1065 18055 1095
rect 18085 1065 18235 1095
rect 18265 1065 18415 1095
rect 18445 1065 18595 1095
rect 18625 1065 18630 1095
rect 16435 1055 18630 1065
rect 16435 1025 16440 1055
rect 16470 1025 16660 1055
rect 16690 1025 16975 1055
rect 17005 1025 17155 1055
rect 17185 1025 17335 1055
rect 17365 1025 17515 1055
rect 17545 1025 17695 1055
rect 17725 1025 17875 1055
rect 17905 1025 18055 1055
rect 18085 1025 18235 1055
rect 18265 1025 18415 1055
rect 18445 1025 18595 1055
rect 18625 1025 18630 1055
rect 16435 1015 18630 1025
rect 16435 985 16440 1015
rect 16470 985 16660 1015
rect 16690 985 16975 1015
rect 17005 985 17155 1015
rect 17185 985 17335 1015
rect 17365 985 17515 1015
rect 17545 985 17695 1015
rect 17725 985 17875 1015
rect 17905 985 18055 1015
rect 18085 985 18235 1015
rect 18265 985 18415 1015
rect 18445 985 18595 1015
rect 18625 985 18630 1015
rect 16435 980 18630 985
rect 18905 1095 19115 1100
rect 18905 1065 18910 1095
rect 18940 1065 19020 1095
rect 19050 1065 19080 1095
rect 19110 1065 19115 1095
rect 18905 1055 19115 1065
rect 18905 1025 18910 1055
rect 18940 1025 19020 1055
rect 19050 1025 19080 1055
rect 19110 1025 19115 1055
rect 18905 1015 19115 1025
rect 18905 985 18910 1015
rect 18940 985 19020 1015
rect 19050 985 19080 1015
rect 19110 985 19115 1015
rect 18905 980 19115 985
rect 16545 915 16585 920
rect 16545 885 16550 915
rect 16580 910 16585 915
rect 16780 915 16820 920
rect 16780 910 16785 915
rect 16580 890 16785 910
rect 16580 885 16585 890
rect 16545 880 16585 885
rect 16780 885 16785 890
rect 16815 885 16820 915
rect 16780 880 16820 885
rect 16480 745 16520 750
rect 16480 715 16485 745
rect 16515 740 16520 745
rect 16610 745 16650 750
rect 16610 740 16615 745
rect 16515 720 16615 740
rect 16515 715 16520 720
rect 16480 710 16520 715
rect 16610 715 16615 720
rect 16645 715 16650 745
rect 16610 710 16650 715
rect 18950 745 18990 750
rect 18950 715 18955 745
rect 18985 740 18990 745
rect 19260 745 19300 750
rect 19260 740 19265 745
rect 18985 720 19265 740
rect 18985 715 18990 720
rect 18950 710 18990 715
rect 19260 715 19265 720
rect 19295 715 19300 745
rect 19260 710 19300 715
rect 19000 685 19650 690
rect 19000 655 19005 685
rect 19035 655 19615 685
rect 19645 655 19650 685
rect 19000 650 19650 655
rect 16315 645 18000 650
rect 16315 615 16320 645
rect 16350 615 17605 645
rect 17635 615 17965 645
rect 17995 615 18000 645
rect 16315 610 18000 615
rect 16260 590 18180 595
rect 16260 560 16265 590
rect 16295 560 16785 590
rect 16815 560 17425 590
rect 17455 560 18145 590
rect 18175 560 18180 590
rect 16260 555 18180 560
rect 16205 535 16245 540
rect 16205 505 16210 535
rect 16240 530 16245 535
rect 16545 535 16585 540
rect 16545 530 16550 535
rect 16240 510 16550 530
rect 16240 505 16245 510
rect 16205 500 16245 505
rect 16545 505 16550 510
rect 16580 530 16585 535
rect 17240 535 17280 540
rect 17240 530 17245 535
rect 16580 510 17245 530
rect 16580 505 16585 510
rect 16545 500 16585 505
rect 17240 505 17245 510
rect 17275 530 17280 535
rect 18320 535 18360 540
rect 18320 530 18325 535
rect 17275 510 18325 530
rect 17275 505 17280 510
rect 17240 500 17280 505
rect 18320 505 18325 510
rect 18355 505 18360 535
rect 18320 500 18360 505
rect 17060 490 17100 495
rect 17060 460 17065 490
rect 17095 485 17100 490
rect 17780 490 17820 495
rect 17780 485 17785 490
rect 17095 465 17785 485
rect 17095 460 17100 465
rect 17060 455 17100 460
rect 17780 460 17785 465
rect 17815 485 17820 490
rect 18500 490 18540 495
rect 18500 485 18505 490
rect 17815 465 18505 485
rect 17815 460 17820 465
rect 17780 455 17820 460
rect 18500 460 18505 465
rect 18535 485 18540 490
rect 19405 490 19445 495
rect 19405 485 19410 490
rect 18535 465 19410 485
rect 18535 460 18540 465
rect 18500 455 18540 460
rect 19405 460 19410 465
rect 19440 460 19445 490
rect 19405 455 19445 460
rect 16420 390 19180 395
rect 16420 360 16425 390
rect 16455 360 16545 390
rect 16575 360 16665 390
rect 16695 360 16785 390
rect 16815 360 16905 390
rect 16935 360 17025 390
rect 17055 360 17145 390
rect 17175 360 17265 390
rect 17295 360 17385 390
rect 17415 360 17505 390
rect 17535 360 17625 390
rect 17655 360 17945 390
rect 17975 360 18065 390
rect 18095 360 18185 390
rect 18215 360 18305 390
rect 18335 360 18425 390
rect 18455 360 18545 390
rect 18575 360 18665 390
rect 18695 360 18785 390
rect 18815 360 18905 390
rect 18935 360 19025 390
rect 19055 360 19145 390
rect 19175 360 19180 390
rect 16420 350 19180 360
rect 16420 320 16425 350
rect 16455 320 16545 350
rect 16575 320 16665 350
rect 16695 320 16785 350
rect 16815 320 16905 350
rect 16935 320 17025 350
rect 17055 320 17145 350
rect 17175 320 17265 350
rect 17295 320 17385 350
rect 17415 320 17505 350
rect 17535 320 17625 350
rect 17655 320 17945 350
rect 17975 320 18065 350
rect 18095 320 18185 350
rect 18215 320 18305 350
rect 18335 320 18425 350
rect 18455 320 18545 350
rect 18575 320 18665 350
rect 18695 320 18785 350
rect 18815 320 18905 350
rect 18935 320 19025 350
rect 19055 320 19145 350
rect 19175 320 19180 350
rect 16420 310 19180 320
rect 16420 280 16425 310
rect 16455 280 16545 310
rect 16575 280 16665 310
rect 16695 280 16785 310
rect 16815 280 16905 310
rect 16935 280 17025 310
rect 17055 280 17145 310
rect 17175 280 17265 310
rect 17295 280 17385 310
rect 17415 280 17505 310
rect 17535 280 17625 310
rect 17655 280 17945 310
rect 17975 280 18065 310
rect 18095 280 18185 310
rect 18215 280 18305 310
rect 18335 280 18425 310
rect 18455 280 18545 310
rect 18575 280 18665 310
rect 18695 280 18785 310
rect 18815 280 18905 310
rect 18935 280 19025 310
rect 19055 280 19145 310
rect 19175 280 19180 310
rect 16420 275 19180 280
rect 15945 175 15985 180
rect 15945 145 15950 175
rect 15980 170 15985 175
rect 16480 175 16520 180
rect 16480 170 16485 175
rect 15980 150 16485 170
rect 15980 145 15985 150
rect 15945 140 15985 145
rect 16480 145 16485 150
rect 16515 170 16520 175
rect 16840 175 16880 180
rect 16840 170 16845 175
rect 16515 150 16845 170
rect 16515 145 16520 150
rect 16480 140 16520 145
rect 16840 145 16845 150
rect 16875 170 16880 175
rect 17200 175 17240 180
rect 17200 170 17205 175
rect 16875 150 17205 170
rect 16875 145 16880 150
rect 16840 140 16880 145
rect 17200 145 17205 150
rect 17235 170 17240 175
rect 17560 175 17600 180
rect 17560 170 17565 175
rect 17235 150 17565 170
rect 17235 145 17240 150
rect 17200 140 17240 145
rect 17560 145 17565 150
rect 17595 170 17600 175
rect 17690 175 17730 180
rect 17690 170 17695 175
rect 17595 150 17695 170
rect 17595 145 17600 150
rect 17560 140 17600 145
rect 17690 145 17695 150
rect 17725 145 17730 175
rect 17690 140 17730 145
rect 17870 175 19650 180
rect 17870 145 17875 175
rect 17905 145 18005 175
rect 18035 145 18365 175
rect 18395 145 18725 175
rect 18755 145 19085 175
rect 19115 145 19615 175
rect 19645 145 19650 175
rect 17870 140 19650 145
rect 16600 5 16640 10
rect 16600 -25 16605 5
rect 16635 0 16640 5
rect 16960 5 17000 10
rect 16960 0 16965 5
rect 16635 -20 16965 0
rect 16635 -25 16640 -20
rect 16600 -30 16640 -25
rect 16960 -25 16965 -20
rect 16995 0 17000 5
rect 17320 5 17360 10
rect 17320 0 17325 5
rect 16995 -20 17325 0
rect 16995 -25 17000 -20
rect 16960 -30 17000 -25
rect 17320 -25 17325 -20
rect 17355 -25 17360 5
rect 17320 -30 17360 -25
rect 18240 5 18280 10
rect 18240 -25 18245 5
rect 18275 0 18280 5
rect 18600 5 18640 10
rect 18600 0 18605 5
rect 18275 -20 18605 0
rect 18275 -25 18280 -20
rect 18240 -30 18280 -25
rect 18600 -25 18605 -20
rect 18635 0 18640 5
rect 18960 5 19000 10
rect 18960 0 18965 5
rect 18635 -20 18965 0
rect 18635 -25 18640 -20
rect 18600 -30 18640 -25
rect 18960 -25 18965 -20
rect 18995 -25 19000 5
rect 18960 -30 19000 -25
rect 15725 -55 15765 -50
rect 15725 -85 15730 -55
rect 15760 -60 15765 -55
rect 16510 -55 16550 -50
rect 16510 -60 16515 -55
rect 15760 -80 16515 -60
rect 15760 -85 15765 -80
rect 15725 -90 15765 -85
rect 16510 -85 16515 -80
rect 16545 -60 16550 -55
rect 16720 -55 16760 -50
rect 16720 -60 16725 -55
rect 16545 -80 16725 -60
rect 16545 -85 16550 -80
rect 16510 -90 16550 -85
rect 16720 -85 16725 -80
rect 16755 -60 16760 -55
rect 16840 -55 16880 -50
rect 16840 -60 16845 -55
rect 16755 -80 16845 -60
rect 16755 -85 16760 -80
rect 16720 -90 16760 -85
rect 16840 -85 16845 -80
rect 16875 -60 16880 -55
rect 17080 -55 17120 -50
rect 17080 -60 17085 -55
rect 16875 -80 17085 -60
rect 16875 -85 16880 -80
rect 16840 -90 16880 -85
rect 17080 -85 17085 -80
rect 17115 -60 17120 -55
rect 17200 -55 17240 -50
rect 17200 -60 17205 -55
rect 17115 -80 17205 -60
rect 17115 -85 17120 -80
rect 17080 -90 17120 -85
rect 17200 -85 17205 -80
rect 17235 -60 17240 -55
rect 17440 -55 17480 -50
rect 17440 -60 17445 -55
rect 17235 -80 17445 -60
rect 17235 -85 17240 -80
rect 17200 -90 17240 -85
rect 17440 -85 17445 -80
rect 17475 -60 17480 -55
rect 17530 -55 17570 -50
rect 17530 -60 17535 -55
rect 17475 -80 17535 -60
rect 17475 -85 17480 -80
rect 17440 -90 17480 -85
rect 17530 -85 17535 -80
rect 17565 -85 17570 -55
rect 17530 -90 17570 -85
rect 18030 -55 18070 -50
rect 18030 -85 18035 -55
rect 18065 -60 18070 -55
rect 18120 -55 18160 -50
rect 18120 -60 18125 -55
rect 18065 -80 18125 -60
rect 18065 -85 18070 -80
rect 18030 -90 18070 -85
rect 18120 -85 18125 -80
rect 18155 -60 18160 -55
rect 18360 -55 18400 -50
rect 18360 -60 18365 -55
rect 18155 -80 18365 -60
rect 18155 -85 18160 -80
rect 18120 -90 18160 -85
rect 18360 -85 18365 -80
rect 18395 -60 18400 -55
rect 18480 -55 18520 -50
rect 18480 -60 18485 -55
rect 18395 -80 18485 -60
rect 18395 -85 18400 -80
rect 18360 -90 18400 -85
rect 18480 -85 18485 -80
rect 18515 -60 18520 -55
rect 18720 -55 18760 -50
rect 18720 -60 18725 -55
rect 18515 -80 18725 -60
rect 18515 -85 18520 -80
rect 18480 -90 18520 -85
rect 18720 -85 18725 -80
rect 18755 -60 18760 -55
rect 18840 -55 18880 -50
rect 18840 -60 18845 -55
rect 18755 -80 18845 -60
rect 18755 -85 18760 -80
rect 18720 -90 18760 -85
rect 18840 -85 18845 -80
rect 18875 -60 18880 -55
rect 19050 -55 19090 -50
rect 19050 -60 19055 -55
rect 18875 -80 19055 -60
rect 18875 -85 18880 -80
rect 18840 -90 18880 -85
rect 19050 -85 19055 -80
rect 19085 -60 19090 -55
rect 19830 -55 19870 -50
rect 19830 -60 19835 -55
rect 19085 -80 19835 -60
rect 19085 -85 19090 -80
rect 19050 -90 19090 -85
rect 19830 -85 19835 -80
rect 19865 -85 19870 -55
rect 19830 -90 19870 -85
rect 16260 -110 17037 -105
rect 16260 -140 16265 -110
rect 16295 -140 17007 -110
rect 18563 -110 18593 -105
rect 18562 -135 18563 -115
rect 16260 -145 17037 -140
rect 19405 -110 19445 -105
rect 19405 -115 19410 -110
rect 18593 -135 19410 -115
rect 18563 -145 18593 -140
rect 19405 -140 19410 -135
rect 19440 -140 19445 -110
rect 19405 -145 19445 -140
rect 17560 -170 18040 -165
rect 17560 -200 17565 -170
rect 17595 -200 17745 -170
rect 17775 -200 17785 -170
rect 17815 -200 17825 -170
rect 17855 -200 18005 -170
rect 18035 -200 18040 -170
rect 17560 -210 18040 -200
rect 17560 -240 17565 -210
rect 17595 -240 17745 -210
rect 17775 -240 17785 -210
rect 17815 -240 17825 -210
rect 17855 -240 18005 -210
rect 18035 -240 18040 -210
rect 17560 -250 18040 -240
rect 17560 -280 17565 -250
rect 17595 -280 17745 -250
rect 17775 -280 17785 -250
rect 17815 -280 17825 -250
rect 17855 -280 18005 -250
rect 18035 -280 18040 -250
rect 17560 -285 18040 -280
rect 16315 -430 17105 -425
rect 16315 -460 16320 -430
rect 16350 -460 17075 -430
rect 16315 -465 17105 -460
rect 18495 -430 18525 -425
rect 19325 -430 19365 -425
rect 19325 -435 19330 -430
rect 18525 -455 19330 -435
rect 18495 -465 18525 -460
rect 19325 -460 19330 -455
rect 19360 -460 19365 -430
rect 19325 -465 19365 -460
rect 16530 -510 17060 -505
rect 16530 -540 16535 -510
rect 16565 -540 17025 -510
rect 17055 -540 17060 -510
rect 16530 -545 17060 -540
rect 18540 -510 18580 -505
rect 18540 -540 18545 -510
rect 18575 -515 18580 -510
rect 19030 -510 19070 -505
rect 19030 -515 19035 -510
rect 18575 -535 19035 -515
rect 18575 -540 18580 -535
rect 18540 -545 18580 -540
rect 19030 -540 19035 -535
rect 19065 -540 19070 -510
rect 19030 -545 19070 -540
rect 16620 -565 18980 -560
rect 16620 -595 16625 -565
rect 16655 -595 16745 -565
rect 16775 -595 16865 -565
rect 16895 -595 16985 -565
rect 17015 -595 17305 -565
rect 17335 -595 17425 -565
rect 17455 -595 17545 -565
rect 17575 -595 18025 -565
rect 18055 -595 18145 -565
rect 18175 -595 18265 -565
rect 18295 -595 18585 -565
rect 18615 -595 18705 -565
rect 18735 -595 18825 -565
rect 18855 -595 18945 -565
rect 18975 -595 18980 -565
rect 16620 -605 18980 -595
rect 16620 -635 16625 -605
rect 16655 -635 16745 -605
rect 16775 -635 16865 -605
rect 16895 -635 16985 -605
rect 17015 -635 17305 -605
rect 17335 -635 17425 -605
rect 17455 -635 17545 -605
rect 17575 -635 18025 -605
rect 18055 -635 18145 -605
rect 18175 -635 18265 -605
rect 18295 -635 18585 -605
rect 18615 -635 18705 -605
rect 18735 -635 18825 -605
rect 18855 -635 18945 -605
rect 18975 -635 18980 -605
rect 16620 -645 18980 -635
rect 16620 -675 16625 -645
rect 16655 -675 16745 -645
rect 16775 -675 16865 -645
rect 16895 -675 16985 -645
rect 17015 -675 17305 -645
rect 17335 -675 17425 -645
rect 17455 -675 17545 -645
rect 17575 -675 18025 -645
rect 18055 -675 18145 -645
rect 18175 -675 18265 -645
rect 18295 -675 18585 -645
rect 18615 -675 18705 -645
rect 18735 -675 18825 -645
rect 18855 -675 18945 -645
rect 18975 -675 18980 -645
rect 16620 -680 18980 -675
rect 17110 -965 18490 -960
rect 17110 -995 17115 -965
rect 17145 -995 17745 -965
rect 17775 -995 17785 -965
rect 17815 -995 17825 -965
rect 17855 -995 18455 -965
rect 18485 -995 18490 -965
rect 17110 -1005 18490 -995
rect 17110 -1035 17115 -1005
rect 17145 -1035 17745 -1005
rect 17775 -1035 17785 -1005
rect 17815 -1035 17825 -1005
rect 17855 -1035 18455 -1005
rect 18485 -1035 18490 -1005
rect 17110 -1045 18490 -1035
rect 17110 -1075 17115 -1045
rect 17145 -1075 17745 -1045
rect 17775 -1075 17785 -1045
rect 17815 -1075 17825 -1045
rect 17855 -1075 18455 -1045
rect 18485 -1075 18490 -1045
rect 17110 -1080 18490 -1075
rect 16740 -1100 16780 -1095
rect 16740 -1130 16745 -1100
rect 16775 -1105 16780 -1100
rect 16820 -1100 16860 -1095
rect 16820 -1105 16825 -1100
rect 16775 -1125 16825 -1105
rect 16775 -1130 16780 -1125
rect 16740 -1135 16780 -1130
rect 16820 -1130 16825 -1125
rect 16855 -1105 16860 -1100
rect 16900 -1100 16940 -1095
rect 16900 -1105 16905 -1100
rect 16855 -1125 16905 -1105
rect 16855 -1130 16860 -1125
rect 16820 -1135 16860 -1130
rect 16900 -1130 16905 -1125
rect 16935 -1105 16940 -1100
rect 16980 -1100 17020 -1095
rect 16980 -1105 16985 -1100
rect 16935 -1125 16985 -1105
rect 16935 -1130 16940 -1125
rect 16900 -1135 16940 -1130
rect 16980 -1130 16985 -1125
rect 17015 -1105 17020 -1100
rect 17060 -1100 17100 -1095
rect 17060 -1105 17065 -1100
rect 17015 -1125 17065 -1105
rect 17015 -1130 17020 -1125
rect 16980 -1135 17020 -1130
rect 17060 -1130 17065 -1125
rect 17095 -1105 17100 -1100
rect 17140 -1100 17180 -1095
rect 17140 -1105 17145 -1100
rect 17095 -1125 17145 -1105
rect 17095 -1130 17100 -1125
rect 17060 -1135 17100 -1130
rect 17140 -1130 17145 -1125
rect 17175 -1105 17180 -1100
rect 17220 -1100 17260 -1095
rect 17220 -1105 17225 -1100
rect 17175 -1125 17225 -1105
rect 17175 -1130 17180 -1125
rect 17140 -1135 17180 -1130
rect 17220 -1130 17225 -1125
rect 17255 -1105 17260 -1100
rect 17300 -1100 17340 -1095
rect 17300 -1105 17305 -1100
rect 17255 -1125 17305 -1105
rect 17255 -1130 17260 -1125
rect 17220 -1135 17260 -1130
rect 17300 -1130 17305 -1125
rect 17335 -1105 17340 -1100
rect 17380 -1100 17420 -1095
rect 17380 -1105 17385 -1100
rect 17335 -1125 17385 -1105
rect 17335 -1130 17340 -1125
rect 17300 -1135 17340 -1130
rect 17380 -1130 17385 -1125
rect 17415 -1105 17420 -1100
rect 17460 -1100 17500 -1095
rect 17460 -1105 17465 -1100
rect 17415 -1125 17465 -1105
rect 17415 -1130 17420 -1125
rect 17380 -1135 17420 -1130
rect 17460 -1130 17465 -1125
rect 17495 -1105 17500 -1100
rect 17540 -1100 17580 -1095
rect 17540 -1105 17545 -1100
rect 17495 -1125 17545 -1105
rect 17495 -1130 17500 -1125
rect 17460 -1135 17500 -1130
rect 17540 -1130 17545 -1125
rect 17575 -1105 17580 -1100
rect 17620 -1100 17660 -1095
rect 17620 -1105 17625 -1100
rect 17575 -1125 17625 -1105
rect 17575 -1130 17580 -1125
rect 17540 -1135 17580 -1130
rect 17620 -1130 17625 -1125
rect 17655 -1105 17660 -1100
rect 17700 -1100 17740 -1095
rect 17700 -1105 17705 -1100
rect 17655 -1125 17705 -1105
rect 17655 -1130 17660 -1125
rect 17620 -1135 17660 -1130
rect 17700 -1130 17705 -1125
rect 17735 -1130 17740 -1100
rect 17700 -1135 17740 -1130
rect 17780 -1100 17820 -1095
rect 17780 -1130 17785 -1100
rect 17815 -1105 17820 -1100
rect 17860 -1100 17900 -1095
rect 17860 -1105 17865 -1100
rect 17815 -1125 17865 -1105
rect 17815 -1130 17820 -1125
rect 17780 -1135 17820 -1130
rect 17860 -1130 17865 -1125
rect 17895 -1105 17900 -1100
rect 17940 -1100 17980 -1095
rect 17940 -1105 17945 -1100
rect 17895 -1125 17945 -1105
rect 17895 -1130 17900 -1125
rect 17860 -1135 17900 -1130
rect 17940 -1130 17945 -1125
rect 17975 -1105 17980 -1100
rect 18020 -1100 18060 -1095
rect 18020 -1105 18025 -1100
rect 17975 -1125 18025 -1105
rect 17975 -1130 17980 -1125
rect 17940 -1135 17980 -1130
rect 18020 -1130 18025 -1125
rect 18055 -1105 18060 -1100
rect 18100 -1100 18140 -1095
rect 18100 -1105 18105 -1100
rect 18055 -1125 18105 -1105
rect 18055 -1130 18060 -1125
rect 18020 -1135 18060 -1130
rect 18100 -1130 18105 -1125
rect 18135 -1105 18140 -1100
rect 18180 -1100 18220 -1095
rect 18180 -1105 18185 -1100
rect 18135 -1125 18185 -1105
rect 18135 -1130 18140 -1125
rect 18100 -1135 18140 -1130
rect 18180 -1130 18185 -1125
rect 18215 -1105 18220 -1100
rect 18260 -1100 18300 -1095
rect 18260 -1105 18265 -1100
rect 18215 -1125 18265 -1105
rect 18215 -1130 18220 -1125
rect 18180 -1135 18220 -1130
rect 18260 -1130 18265 -1125
rect 18295 -1105 18300 -1100
rect 18340 -1100 18380 -1095
rect 18340 -1105 18345 -1100
rect 18295 -1125 18345 -1105
rect 18295 -1130 18300 -1125
rect 18260 -1135 18300 -1130
rect 18340 -1130 18345 -1125
rect 18375 -1105 18380 -1100
rect 18420 -1100 18460 -1095
rect 18420 -1105 18425 -1100
rect 18375 -1125 18425 -1105
rect 18375 -1130 18380 -1125
rect 18340 -1135 18380 -1130
rect 18420 -1130 18425 -1125
rect 18455 -1105 18460 -1100
rect 18500 -1100 18540 -1095
rect 18500 -1105 18505 -1100
rect 18455 -1125 18505 -1105
rect 18455 -1130 18460 -1125
rect 18420 -1135 18460 -1130
rect 18500 -1130 18505 -1125
rect 18535 -1105 18540 -1100
rect 18580 -1100 18620 -1095
rect 18580 -1105 18585 -1100
rect 18535 -1125 18585 -1105
rect 18535 -1130 18540 -1125
rect 18500 -1135 18540 -1130
rect 18580 -1130 18585 -1125
rect 18615 -1105 18620 -1100
rect 18660 -1100 18700 -1095
rect 18660 -1105 18665 -1100
rect 18615 -1125 18665 -1105
rect 18615 -1130 18620 -1125
rect 18580 -1135 18620 -1130
rect 18660 -1130 18665 -1125
rect 18695 -1105 18700 -1100
rect 18740 -1100 18780 -1095
rect 18740 -1105 18745 -1100
rect 18695 -1125 18745 -1105
rect 18695 -1130 18700 -1125
rect 18660 -1135 18700 -1130
rect 18740 -1130 18745 -1125
rect 18775 -1130 18780 -1100
rect 18740 -1135 18780 -1130
rect 18895 -1165 18935 -1160
rect 16205 -1185 16245 -1180
rect 16205 -1215 16210 -1185
rect 16240 -1190 16245 -1185
rect 16700 -1185 16740 -1180
rect 16700 -1190 16705 -1185
rect 16240 -1210 16705 -1190
rect 16240 -1215 16245 -1210
rect 16205 -1220 16245 -1215
rect 16700 -1215 16705 -1210
rect 16735 -1215 16740 -1185
rect 16700 -1220 16740 -1215
rect 18895 -1195 18900 -1165
rect 18930 -1195 18935 -1165
rect 18895 -1205 18935 -1195
rect 18895 -1235 18900 -1205
rect 18930 -1235 18935 -1205
rect 18895 -1240 18935 -1235
rect 15890 -1355 18300 -1350
rect 15890 -1385 15895 -1355
rect 15925 -1385 16660 -1355
rect 16690 -1385 16770 -1355
rect 16800 -1385 17305 -1355
rect 17335 -1385 17785 -1355
rect 17815 -1385 18265 -1355
rect 18295 -1385 18300 -1355
rect 15890 -1390 18300 -1385
rect 16600 -1410 18575 -1405
rect 16600 -1440 16605 -1410
rect 16635 -1440 16715 -1410
rect 16745 -1440 16825 -1410
rect 16855 -1440 16885 -1410
rect 16915 -1440 17030 -1410
rect 17060 -1440 17140 -1410
rect 17170 -1440 17250 -1410
rect 17280 -1440 17360 -1410
rect 17390 -1440 17470 -1410
rect 17500 -1440 17620 -1410
rect 17650 -1440 17730 -1410
rect 17760 -1440 17840 -1410
rect 17870 -1440 17950 -1410
rect 17980 -1440 18100 -1410
rect 18130 -1440 18210 -1410
rect 18240 -1440 18320 -1410
rect 18350 -1440 18430 -1410
rect 18460 -1440 18540 -1410
rect 18570 -1440 18575 -1410
rect 16600 -1450 18575 -1440
rect 16600 -1480 16605 -1450
rect 16635 -1480 16715 -1450
rect 16745 -1480 16825 -1450
rect 16855 -1480 16885 -1450
rect 16915 -1480 17030 -1450
rect 17060 -1480 17140 -1450
rect 17170 -1480 17250 -1450
rect 17280 -1480 17360 -1450
rect 17390 -1480 17470 -1450
rect 17500 -1480 17620 -1450
rect 17650 -1480 17730 -1450
rect 17760 -1480 17840 -1450
rect 17870 -1480 17950 -1450
rect 17980 -1480 18100 -1450
rect 18130 -1480 18210 -1450
rect 18240 -1480 18320 -1450
rect 18350 -1480 18430 -1450
rect 18460 -1480 18540 -1450
rect 18570 -1480 18575 -1450
rect 16600 -1490 18575 -1480
rect 16600 -1520 16605 -1490
rect 16635 -1520 16715 -1490
rect 16745 -1520 16825 -1490
rect 16855 -1520 16885 -1490
rect 16915 -1520 17030 -1490
rect 17060 -1520 17140 -1490
rect 17170 -1520 17250 -1490
rect 17280 -1520 17360 -1490
rect 17390 -1520 17470 -1490
rect 17500 -1520 17620 -1490
rect 17650 -1520 17730 -1490
rect 17760 -1520 17840 -1490
rect 17870 -1520 17950 -1490
rect 17980 -1520 18100 -1490
rect 18130 -1520 18210 -1490
rect 18240 -1520 18320 -1490
rect 18350 -1520 18430 -1490
rect 18460 -1520 18540 -1490
rect 18570 -1520 18575 -1490
rect 16600 -1525 18575 -1520
rect 17190 -1660 17450 -1655
rect 17190 -1690 17195 -1660
rect 17225 -1690 17415 -1660
rect 17445 -1690 17450 -1660
rect 17190 -1695 17450 -1690
rect 17670 -1660 17710 -1655
rect 17670 -1690 17675 -1660
rect 17705 -1665 17710 -1660
rect 17780 -1660 17820 -1655
rect 17780 -1665 17785 -1660
rect 17705 -1685 17785 -1665
rect 17705 -1690 17710 -1685
rect 17670 -1695 17710 -1690
rect 17780 -1690 17785 -1685
rect 17815 -1665 17820 -1660
rect 17890 -1660 17930 -1655
rect 17890 -1665 17895 -1660
rect 17815 -1685 17895 -1665
rect 17815 -1690 17820 -1685
rect 17780 -1695 17820 -1690
rect 17890 -1690 17895 -1685
rect 17925 -1690 17930 -1660
rect 17890 -1695 17930 -1690
rect 18150 -1660 18410 -1655
rect 18150 -1690 18155 -1660
rect 18185 -1690 18375 -1660
rect 18405 -1690 18410 -1660
rect 18150 -1695 18410 -1690
rect 16030 -1715 16070 -1710
rect 16030 -1745 16035 -1715
rect 16065 -1720 16070 -1715
rect 17080 -1715 17120 -1710
rect 17080 -1720 17085 -1715
rect 16065 -1740 17085 -1720
rect 16065 -1745 16070 -1740
rect 16030 -1750 16070 -1745
rect 17080 -1745 17085 -1740
rect 17115 -1720 17120 -1715
rect 17300 -1715 17340 -1710
rect 17300 -1720 17305 -1715
rect 17115 -1740 17305 -1720
rect 17115 -1745 17120 -1740
rect 17080 -1750 17120 -1745
rect 17300 -1745 17305 -1740
rect 17335 -1720 17340 -1715
rect 18260 -1715 18300 -1710
rect 18260 -1720 18265 -1715
rect 17335 -1740 18265 -1720
rect 17335 -1745 17340 -1740
rect 17300 -1750 17340 -1745
rect 18260 -1745 18265 -1740
rect 18295 -1720 18300 -1715
rect 18480 -1715 18520 -1710
rect 18480 -1720 18485 -1715
rect 18295 -1740 18485 -1720
rect 18295 -1745 18300 -1740
rect 18260 -1750 18300 -1745
rect 18480 -1745 18485 -1740
rect 18515 -1745 18520 -1715
rect 18480 -1750 18520 -1745
rect 15785 -1770 17230 -1765
rect 15785 -1800 15790 -1770
rect 15820 -1800 17195 -1770
rect 17225 -1800 17230 -1770
rect 15785 -1805 17230 -1800
rect 18370 -1770 18410 -1765
rect 18370 -1800 18375 -1770
rect 18405 -1775 18410 -1770
rect 19775 -1770 19815 -1765
rect 19775 -1775 19780 -1770
rect 18405 -1795 19780 -1775
rect 18405 -1800 18410 -1795
rect 18370 -1805 18410 -1800
rect 19775 -1800 19780 -1795
rect 19810 -1800 19815 -1770
rect 19775 -1805 19815 -1800
rect 16105 -1865 16145 -1860
rect 16105 -1895 16110 -1865
rect 16140 -1870 16145 -1865
rect 16765 -1865 16805 -1860
rect 16765 -1870 16770 -1865
rect 16140 -1890 16770 -1870
rect 16140 -1895 16145 -1890
rect 16105 -1900 16145 -1895
rect 16765 -1895 16770 -1890
rect 16800 -1895 16805 -1865
rect 16765 -1900 16805 -1895
rect 17780 -1900 17820 -1895
rect 17780 -1930 17785 -1900
rect 17815 -1905 17820 -1900
rect 19535 -1900 19575 -1895
rect 19535 -1905 19540 -1900
rect 17815 -1925 19540 -1905
rect 17815 -1930 17820 -1925
rect 17780 -1935 17820 -1930
rect 19535 -1930 19540 -1925
rect 19570 -1930 19575 -1900
rect 19535 -1935 19575 -1930
rect 16155 -1950 16195 -1945
rect 16155 -1980 16160 -1950
rect 16190 -1955 16195 -1950
rect 19325 -1950 19365 -1945
rect 19325 -1955 19330 -1950
rect 16190 -1975 19330 -1955
rect 16190 -1980 16195 -1975
rect 16155 -1985 16195 -1980
rect 19325 -1980 19330 -1975
rect 19360 -1980 19365 -1950
rect 19325 -1985 19365 -1980
rect 16315 -2000 16355 -1995
rect 16315 -2030 16320 -2000
rect 16350 -2030 17430 -2000
rect 16315 -2035 17430 -2030
rect 17465 -2035 17470 -2000
rect 18124 -2035 18129 -2000
rect 18164 -2005 18870 -2000
rect 18164 -2035 18835 -2005
rect 18865 -2035 18870 -2005
rect 18165 -2040 18870 -2035
rect 17425 -2060 19120 -2055
rect 17425 -2090 17430 -2060
rect 17460 -2090 19085 -2060
rect 19115 -2090 19120 -2060
rect 17425 -2095 19120 -2090
rect 16260 -2100 16770 -2095
rect 16260 -2130 16265 -2100
rect 16295 -2130 16485 -2100
rect 16515 -2130 16735 -2100
rect 16765 -2130 16770 -2100
rect 16260 -2135 16770 -2130
rect 16485 -2900 16520 -2895
rect 16485 -2940 16520 -2935
rect 19080 -2900 19115 -2895
rect 19080 -2940 19115 -2935
rect 19405 -2997 19440 -2992
rect 16160 -3025 16195 -3020
rect 19405 -3037 19440 -3032
rect 16160 -3065 16195 -3060
rect 16730 -3105 17820 -3100
rect 15820 -3115 15860 -3110
rect 15820 -3145 15825 -3115
rect 15855 -3120 15860 -3115
rect 15950 -3116 15985 -3110
rect 15855 -3140 15950 -3120
rect 15855 -3145 15860 -3140
rect 15820 -3150 15860 -3145
rect 16730 -3135 16735 -3105
rect 16765 -3135 17785 -3105
rect 17815 -3135 17820 -3105
rect 16730 -3140 17820 -3135
rect 18615 -3105 18870 -3100
rect 18615 -3135 18620 -3105
rect 18650 -3135 18835 -3105
rect 18865 -3135 18870 -3105
rect 18615 -3140 18870 -3135
rect 19610 -3115 19645 -3110
rect 15950 -3156 15985 -3151
rect 19610 -3160 19645 -3150
rect 15950 -3789 15985 -3784
rect 15950 -3829 15985 -3824
rect 19610 -3789 19645 -3784
rect 19610 -3829 19645 -3824
rect 15960 -3830 15980 -3829
rect 19620 -3830 19640 -3829
rect 16280 -3894 16315 -3889
rect 16280 -3934 16315 -3929
rect 19285 -3894 19320 -3889
rect 19285 -3934 19320 -3929
rect 16290 -3935 16310 -3934
rect 19290 -3935 19310 -3934
rect 16605 -3969 16640 -3964
rect 16605 -4009 16640 -4004
rect 18960 -3969 18995 -3964
rect 18960 -4009 18995 -4004
rect 16615 -4010 16635 -4009
rect 18965 -4010 18985 -4009
rect 16280 -4190 16320 -4185
rect 16280 -4195 16285 -4190
rect 15665 -4215 16285 -4195
rect 16280 -4220 16285 -4215
rect 16315 -4195 16320 -4190
rect 16605 -4190 16645 -4185
rect 16605 -4195 16610 -4190
rect 16315 -4215 16610 -4195
rect 16315 -4220 16320 -4215
rect 16280 -4225 16320 -4220
rect 16605 -4220 16610 -4215
rect 16640 -4220 16645 -4190
rect 16605 -4225 16645 -4220
rect 15820 -4265 15860 -4260
rect 15820 -4295 15825 -4265
rect 15855 -4270 15860 -4265
rect 17250 -4265 17300 -4255
rect 17250 -4270 17260 -4265
rect 15855 -4290 17260 -4270
rect 15855 -4295 15860 -4290
rect 15820 -4300 15860 -4295
rect 17250 -4295 17260 -4290
rect 17290 -4295 17300 -4265
rect 17250 -4305 17300 -4295
rect 17780 -4265 17820 -4260
rect 17780 -4295 17785 -4265
rect 17815 -4270 17820 -4265
rect 18955 -4265 18995 -4260
rect 18955 -4270 18960 -4265
rect 17815 -4290 18960 -4270
rect 17815 -4295 17820 -4290
rect 17780 -4300 17820 -4295
rect 18955 -4295 18960 -4290
rect 18990 -4270 18995 -4265
rect 19280 -4265 19320 -4260
rect 19280 -4270 19285 -4265
rect 18990 -4290 19285 -4270
rect 18990 -4295 18995 -4290
rect 18955 -4300 18995 -4295
rect 19280 -4295 19285 -4290
rect 19315 -4295 19320 -4265
rect 19280 -4300 19320 -4295
rect 15725 -4315 15765 -4310
rect 15725 -4345 15730 -4315
rect 15760 -4320 15765 -4315
rect 16900 -4315 16950 -4305
rect 16900 -4320 16910 -4315
rect 15760 -4340 16910 -4320
rect 15760 -4345 15765 -4340
rect 15725 -4350 15765 -4345
rect 16900 -4345 16910 -4340
rect 16940 -4345 16950 -4315
rect 16900 -4355 16950 -4345
rect 18650 -4315 18700 -4305
rect 18650 -4345 18660 -4315
rect 18690 -4320 18700 -4315
rect 19830 -4315 19870 -4310
rect 19830 -4320 19835 -4315
rect 18690 -4340 19835 -4320
rect 18690 -4345 18700 -4340
rect 18650 -4355 18700 -4345
rect 19830 -4345 19835 -4340
rect 19865 -4345 19870 -4315
rect 19830 -4350 19870 -4345
rect 15950 -4360 15990 -4355
rect 15950 -4390 15955 -4360
rect 15985 -4365 15990 -4360
rect 16205 -4360 16245 -4355
rect 16205 -4365 16210 -4360
rect 15985 -4385 16210 -4365
rect 15985 -4390 15990 -4385
rect 15950 -4395 15990 -4390
rect 16205 -4390 16210 -4385
rect 16240 -4390 16245 -4360
rect 16205 -4395 16245 -4390
rect 19355 -4360 19395 -4355
rect 19355 -4390 19360 -4360
rect 19390 -4365 19395 -4360
rect 19610 -4360 19650 -4355
rect 19610 -4365 19615 -4360
rect 19390 -4385 19615 -4365
rect 19390 -4390 19395 -4385
rect 19355 -4395 19395 -4390
rect 19610 -4390 19615 -4385
rect 19645 -4390 19650 -4360
rect 19610 -4395 19650 -4390
rect 17955 -4410 17995 -4405
rect 17955 -4440 17960 -4410
rect 17990 -4415 17995 -4410
rect 17990 -4435 19905 -4415
rect 17990 -4440 17995 -4435
rect 17955 -4445 17995 -4440
<< via2 >>
rect 17260 -4295 17290 -4265
rect 16910 -4345 16940 -4315
rect 18660 -4345 18690 -4315
rect 16210 -4390 16240 -4360
rect 19360 -4390 19390 -4360
rect 17960 -4440 17990 -4410
<< metal3 >>
rect 17250 -4260 17300 -4255
rect 17250 -4300 17255 -4260
rect 17295 -4300 17300 -4260
rect 17250 -4305 17300 -4300
rect 16900 -4310 16950 -4305
rect 16900 -4350 16905 -4310
rect 16945 -4350 16950 -4310
rect 16900 -4355 16950 -4350
rect 18650 -4310 18700 -4305
rect 18650 -4350 18655 -4310
rect 18695 -4350 18700 -4310
rect 18650 -4355 18700 -4350
rect 16205 -4360 16245 -4355
rect 16205 -4390 16210 -4360
rect 16240 -4390 16245 -4360
rect 16205 -4520 16245 -4390
rect 19355 -4360 19395 -4355
rect 19355 -4390 19360 -4360
rect 19390 -4390 19395 -4360
rect 17955 -4410 17995 -4405
rect 17955 -4440 17960 -4410
rect 17990 -4440 17995 -4410
rect 17955 -4520 17995 -4440
rect 19355 -4520 19395 -4390
rect 15760 -4615 15990 -4520
rect 16110 -4615 16340 -4520
rect 16460 -4615 16690 -4520
rect 16810 -4615 17040 -4520
rect 15760 -4665 17040 -4615
rect 15760 -4750 15990 -4665
rect 16110 -4750 16340 -4665
rect 16460 -4750 16690 -4665
rect 16810 -4750 17040 -4665
rect 17160 -4615 17390 -4520
rect 17510 -4615 17740 -4520
rect 17860 -4615 18090 -4520
rect 18210 -4615 18440 -4520
rect 17160 -4665 18440 -4615
rect 17160 -4750 17390 -4665
rect 17510 -4750 17740 -4665
rect 17860 -4750 18090 -4665
rect 18210 -4750 18440 -4665
rect 18560 -4615 18790 -4520
rect 18910 -4615 19140 -4520
rect 19260 -4615 19490 -4520
rect 19610 -4615 19840 -4520
rect 18560 -4665 19840 -4615
rect 18560 -4750 18790 -4665
rect 18910 -4750 19140 -4665
rect 19260 -4750 19490 -4665
rect 19610 -4750 19840 -4665
rect 16200 -4870 16250 -4750
rect 17950 -4870 18000 -4750
rect 19350 -4870 19400 -4750
rect 15760 -4965 15990 -4870
rect 16110 -4965 16340 -4870
rect 16460 -4965 16690 -4870
rect 16810 -4965 17040 -4870
rect 15760 -5015 17040 -4965
rect 15760 -5100 15990 -5015
rect 16110 -5100 16340 -5015
rect 16460 -5100 16690 -5015
rect 16810 -5100 17040 -5015
rect 17160 -4965 17390 -4870
rect 17510 -4965 17740 -4870
rect 17860 -4965 18090 -4870
rect 18210 -4965 18440 -4870
rect 17160 -5015 18440 -4965
rect 17160 -5100 17390 -5015
rect 17510 -5100 17740 -5015
rect 17860 -5100 18090 -5015
rect 18210 -5100 18440 -5015
rect 18560 -4965 18790 -4870
rect 18910 -4965 19140 -4870
rect 19260 -4965 19490 -4870
rect 19610 -4965 19840 -4870
rect 18560 -5015 19840 -4965
rect 18560 -5100 18790 -5015
rect 18910 -5100 19140 -5015
rect 19260 -5100 19490 -5015
rect 19610 -5100 19840 -5015
rect 16200 -5220 16250 -5100
rect 17950 -5220 18000 -5100
rect 19350 -5220 19400 -5100
rect 15760 -5315 15990 -5220
rect 16110 -5315 16340 -5220
rect 16460 -5315 16690 -5220
rect 16810 -5315 17040 -5220
rect 15760 -5365 17040 -5315
rect 15760 -5450 15990 -5365
rect 16110 -5450 16340 -5365
rect 16460 -5450 16690 -5365
rect 16810 -5450 17040 -5365
rect 17160 -5315 17390 -5220
rect 17510 -5315 17740 -5220
rect 17860 -5315 18090 -5220
rect 18210 -5315 18440 -5220
rect 17160 -5365 18440 -5315
rect 17160 -5450 17390 -5365
rect 17510 -5450 17740 -5365
rect 17860 -5450 18090 -5365
rect 18210 -5450 18440 -5365
rect 18560 -5315 18790 -5220
rect 18910 -5315 19140 -5220
rect 19260 -5315 19490 -5220
rect 19610 -5315 19840 -5220
rect 18560 -5365 19840 -5315
rect 18560 -5450 18790 -5365
rect 18910 -5450 19140 -5365
rect 19260 -5450 19490 -5365
rect 19610 -5450 19840 -5365
rect 16200 -5570 16250 -5450
rect 17950 -5570 18000 -5450
rect 19350 -5570 19400 -5450
rect 15760 -5665 15990 -5570
rect 16110 -5665 16340 -5570
rect 16460 -5665 16690 -5570
rect 16810 -5665 17040 -5570
rect 15760 -5715 17040 -5665
rect 15760 -5800 15990 -5715
rect 16110 -5800 16340 -5715
rect 16460 -5800 16690 -5715
rect 16810 -5800 17040 -5715
rect 17160 -5665 17390 -5570
rect 17510 -5665 17740 -5570
rect 17860 -5665 18090 -5570
rect 18210 -5665 18440 -5570
rect 17160 -5715 18440 -5665
rect 17160 -5800 17390 -5715
rect 17510 -5800 17740 -5715
rect 17860 -5800 18090 -5715
rect 18210 -5800 18440 -5715
rect 18560 -5665 18790 -5570
rect 18910 -5665 19140 -5570
rect 19260 -5665 19490 -5570
rect 19610 -5665 19840 -5570
rect 18560 -5715 19840 -5665
rect 18560 -5800 18790 -5715
rect 18910 -5800 19140 -5715
rect 19260 -5800 19490 -5715
rect 19610 -5800 19840 -5715
rect 16200 -5920 16250 -5800
rect 17950 -5920 18000 -5800
rect 19350 -5920 19400 -5800
rect 15760 -6015 15990 -5920
rect 16110 -6015 16340 -5920
rect 16460 -6015 16690 -5920
rect 16810 -6015 17040 -5920
rect 15760 -6065 17040 -6015
rect 15760 -6150 15990 -6065
rect 16110 -6150 16340 -6065
rect 16460 -6150 16690 -6065
rect 16810 -6150 17040 -6065
rect 17160 -6015 17390 -5920
rect 17510 -6015 17740 -5920
rect 17860 -6015 18090 -5920
rect 18210 -6015 18440 -5920
rect 17160 -6065 18440 -6015
rect 17160 -6150 17390 -6065
rect 17510 -6150 17740 -6065
rect 17860 -6150 18090 -6065
rect 18210 -6150 18440 -6065
rect 18560 -6015 18790 -5920
rect 18910 -6015 19140 -5920
rect 19260 -6015 19490 -5920
rect 19610 -6015 19840 -5920
rect 18560 -6065 19840 -6015
rect 18560 -6150 18790 -6065
rect 18910 -6150 19140 -6065
rect 19260 -6150 19490 -6065
rect 19610 -6150 19840 -6065
<< via3 >>
rect 17255 -4265 17295 -4260
rect 17255 -4295 17260 -4265
rect 17260 -4295 17290 -4265
rect 17290 -4295 17295 -4265
rect 17255 -4300 17295 -4295
rect 16905 -4315 16945 -4310
rect 16905 -4345 16910 -4315
rect 16910 -4345 16940 -4315
rect 16940 -4345 16945 -4315
rect 16905 -4350 16945 -4345
rect 18655 -4315 18695 -4310
rect 18655 -4345 18660 -4315
rect 18660 -4345 18690 -4315
rect 18690 -4345 18695 -4315
rect 18655 -4350 18695 -4345
<< mimcap >>
rect 15775 -4620 15975 -4535
rect 15775 -4660 15855 -4620
rect 15895 -4660 15975 -4620
rect 15775 -4735 15975 -4660
rect 16125 -4620 16325 -4535
rect 16125 -4660 16205 -4620
rect 16245 -4660 16325 -4620
rect 16125 -4735 16325 -4660
rect 16475 -4620 16675 -4535
rect 16475 -4660 16555 -4620
rect 16595 -4660 16675 -4620
rect 16475 -4735 16675 -4660
rect 16825 -4620 17025 -4535
rect 16825 -4660 16905 -4620
rect 16945 -4660 17025 -4620
rect 16825 -4735 17025 -4660
rect 17175 -4620 17375 -4535
rect 17175 -4660 17255 -4620
rect 17295 -4660 17375 -4620
rect 17175 -4735 17375 -4660
rect 17525 -4620 17725 -4535
rect 17525 -4660 17605 -4620
rect 17645 -4660 17725 -4620
rect 17525 -4735 17725 -4660
rect 17875 -4620 18075 -4535
rect 17875 -4660 17955 -4620
rect 17995 -4660 18075 -4620
rect 17875 -4735 18075 -4660
rect 18225 -4620 18425 -4535
rect 18225 -4660 18305 -4620
rect 18345 -4660 18425 -4620
rect 18225 -4735 18425 -4660
rect 18575 -4620 18775 -4535
rect 18575 -4660 18655 -4620
rect 18695 -4660 18775 -4620
rect 18575 -4735 18775 -4660
rect 18925 -4620 19125 -4535
rect 18925 -4660 19005 -4620
rect 19045 -4660 19125 -4620
rect 18925 -4735 19125 -4660
rect 19275 -4620 19475 -4535
rect 19275 -4660 19355 -4620
rect 19395 -4660 19475 -4620
rect 19275 -4735 19475 -4660
rect 19625 -4620 19825 -4535
rect 19625 -4660 19705 -4620
rect 19745 -4660 19825 -4620
rect 19625 -4735 19825 -4660
rect 15775 -4970 15975 -4885
rect 15775 -5010 15855 -4970
rect 15895 -5010 15975 -4970
rect 15775 -5085 15975 -5010
rect 16125 -4970 16325 -4885
rect 16125 -5010 16205 -4970
rect 16245 -5010 16325 -4970
rect 16125 -5085 16325 -5010
rect 16475 -4970 16675 -4885
rect 16475 -5010 16555 -4970
rect 16595 -5010 16675 -4970
rect 16475 -5085 16675 -5010
rect 16825 -4970 17025 -4885
rect 16825 -5010 16905 -4970
rect 16945 -5010 17025 -4970
rect 16825 -5085 17025 -5010
rect 17175 -4970 17375 -4885
rect 17175 -5010 17255 -4970
rect 17295 -5010 17375 -4970
rect 17175 -5085 17375 -5010
rect 17525 -4970 17725 -4885
rect 17525 -5010 17605 -4970
rect 17645 -5010 17725 -4970
rect 17525 -5085 17725 -5010
rect 17875 -4970 18075 -4885
rect 17875 -5010 17955 -4970
rect 17995 -5010 18075 -4970
rect 17875 -5085 18075 -5010
rect 18225 -4970 18425 -4885
rect 18225 -5010 18305 -4970
rect 18345 -5010 18425 -4970
rect 18225 -5085 18425 -5010
rect 18575 -4970 18775 -4885
rect 18575 -5010 18655 -4970
rect 18695 -5010 18775 -4970
rect 18575 -5085 18775 -5010
rect 18925 -4970 19125 -4885
rect 18925 -5010 19005 -4970
rect 19045 -5010 19125 -4970
rect 18925 -5085 19125 -5010
rect 19275 -4970 19475 -4885
rect 19275 -5010 19355 -4970
rect 19395 -5010 19475 -4970
rect 19275 -5085 19475 -5010
rect 19625 -4970 19825 -4885
rect 19625 -5010 19705 -4970
rect 19745 -5010 19825 -4970
rect 19625 -5085 19825 -5010
rect 15775 -5320 15975 -5235
rect 15775 -5360 15855 -5320
rect 15895 -5360 15975 -5320
rect 15775 -5435 15975 -5360
rect 16125 -5320 16325 -5235
rect 16125 -5360 16205 -5320
rect 16245 -5360 16325 -5320
rect 16125 -5435 16325 -5360
rect 16475 -5320 16675 -5235
rect 16475 -5360 16555 -5320
rect 16595 -5360 16675 -5320
rect 16475 -5435 16675 -5360
rect 16825 -5320 17025 -5235
rect 16825 -5360 16905 -5320
rect 16945 -5360 17025 -5320
rect 16825 -5435 17025 -5360
rect 17175 -5320 17375 -5235
rect 17175 -5360 17255 -5320
rect 17295 -5360 17375 -5320
rect 17175 -5435 17375 -5360
rect 17525 -5320 17725 -5235
rect 17525 -5360 17605 -5320
rect 17645 -5360 17725 -5320
rect 17525 -5435 17725 -5360
rect 17875 -5320 18075 -5235
rect 17875 -5360 17955 -5320
rect 17995 -5360 18075 -5320
rect 17875 -5435 18075 -5360
rect 18225 -5320 18425 -5235
rect 18225 -5360 18305 -5320
rect 18345 -5360 18425 -5320
rect 18225 -5435 18425 -5360
rect 18575 -5320 18775 -5235
rect 18575 -5360 18655 -5320
rect 18695 -5360 18775 -5320
rect 18575 -5435 18775 -5360
rect 18925 -5320 19125 -5235
rect 18925 -5360 19005 -5320
rect 19045 -5360 19125 -5320
rect 18925 -5435 19125 -5360
rect 19275 -5320 19475 -5235
rect 19275 -5360 19355 -5320
rect 19395 -5360 19475 -5320
rect 19275 -5435 19475 -5360
rect 19625 -5320 19825 -5235
rect 19625 -5360 19705 -5320
rect 19745 -5360 19825 -5320
rect 19625 -5435 19825 -5360
rect 15775 -5670 15975 -5585
rect 15775 -5710 15855 -5670
rect 15895 -5710 15975 -5670
rect 15775 -5785 15975 -5710
rect 16125 -5670 16325 -5585
rect 16125 -5710 16205 -5670
rect 16245 -5710 16325 -5670
rect 16125 -5785 16325 -5710
rect 16475 -5670 16675 -5585
rect 16475 -5710 16555 -5670
rect 16595 -5710 16675 -5670
rect 16475 -5785 16675 -5710
rect 16825 -5670 17025 -5585
rect 16825 -5710 16905 -5670
rect 16945 -5710 17025 -5670
rect 16825 -5785 17025 -5710
rect 17175 -5670 17375 -5585
rect 17175 -5710 17255 -5670
rect 17295 -5710 17375 -5670
rect 17175 -5785 17375 -5710
rect 17525 -5670 17725 -5585
rect 17525 -5710 17605 -5670
rect 17645 -5710 17725 -5670
rect 17525 -5785 17725 -5710
rect 17875 -5670 18075 -5585
rect 17875 -5710 17955 -5670
rect 17995 -5710 18075 -5670
rect 17875 -5785 18075 -5710
rect 18225 -5670 18425 -5585
rect 18225 -5710 18305 -5670
rect 18345 -5710 18425 -5670
rect 18225 -5785 18425 -5710
rect 18575 -5670 18775 -5585
rect 18575 -5710 18655 -5670
rect 18695 -5710 18775 -5670
rect 18575 -5785 18775 -5710
rect 18925 -5670 19125 -5585
rect 18925 -5710 19005 -5670
rect 19045 -5710 19125 -5670
rect 18925 -5785 19125 -5710
rect 19275 -5670 19475 -5585
rect 19275 -5710 19355 -5670
rect 19395 -5710 19475 -5670
rect 19275 -5785 19475 -5710
rect 19625 -5670 19825 -5585
rect 19625 -5710 19705 -5670
rect 19745 -5710 19825 -5670
rect 19625 -5785 19825 -5710
rect 15775 -6020 15975 -5935
rect 15775 -6060 15855 -6020
rect 15895 -6060 15975 -6020
rect 15775 -6135 15975 -6060
rect 16125 -6020 16325 -5935
rect 16125 -6060 16205 -6020
rect 16245 -6060 16325 -6020
rect 16125 -6135 16325 -6060
rect 16475 -6020 16675 -5935
rect 16475 -6060 16555 -6020
rect 16595 -6060 16675 -6020
rect 16475 -6135 16675 -6060
rect 16825 -6020 17025 -5935
rect 16825 -6060 16905 -6020
rect 16945 -6060 17025 -6020
rect 16825 -6135 17025 -6060
rect 17175 -6020 17375 -5935
rect 17175 -6060 17255 -6020
rect 17295 -6060 17375 -6020
rect 17175 -6135 17375 -6060
rect 17525 -6020 17725 -5935
rect 17525 -6060 17605 -6020
rect 17645 -6060 17725 -6020
rect 17525 -6135 17725 -6060
rect 17875 -6020 18075 -5935
rect 17875 -6060 17955 -6020
rect 17995 -6060 18075 -6020
rect 17875 -6135 18075 -6060
rect 18225 -6020 18425 -5935
rect 18225 -6060 18305 -6020
rect 18345 -6060 18425 -6020
rect 18225 -6135 18425 -6060
rect 18575 -6020 18775 -5935
rect 18575 -6060 18655 -6020
rect 18695 -6060 18775 -6020
rect 18575 -6135 18775 -6060
rect 18925 -6020 19125 -5935
rect 18925 -6060 19005 -6020
rect 19045 -6060 19125 -6020
rect 18925 -6135 19125 -6060
rect 19275 -6020 19475 -5935
rect 19275 -6060 19355 -6020
rect 19395 -6060 19475 -6020
rect 19275 -6135 19475 -6060
rect 19625 -6020 19825 -5935
rect 19625 -6060 19705 -6020
rect 19745 -6060 19825 -6020
rect 19625 -6135 19825 -6060
<< mimcapcontact >>
rect 15855 -4660 15895 -4620
rect 16205 -4660 16245 -4620
rect 16555 -4660 16595 -4620
rect 16905 -4660 16945 -4620
rect 17255 -4660 17295 -4620
rect 17605 -4660 17645 -4620
rect 17955 -4660 17995 -4620
rect 18305 -4660 18345 -4620
rect 18655 -4660 18695 -4620
rect 19005 -4660 19045 -4620
rect 19355 -4660 19395 -4620
rect 19705 -4660 19745 -4620
rect 15855 -5010 15895 -4970
rect 16205 -5010 16245 -4970
rect 16555 -5010 16595 -4970
rect 16905 -5010 16945 -4970
rect 17255 -5010 17295 -4970
rect 17605 -5010 17645 -4970
rect 17955 -5010 17995 -4970
rect 18305 -5010 18345 -4970
rect 18655 -5010 18695 -4970
rect 19005 -5010 19045 -4970
rect 19355 -5010 19395 -4970
rect 19705 -5010 19745 -4970
rect 15855 -5360 15895 -5320
rect 16205 -5360 16245 -5320
rect 16555 -5360 16595 -5320
rect 16905 -5360 16945 -5320
rect 17255 -5360 17295 -5320
rect 17605 -5360 17645 -5320
rect 17955 -5360 17995 -5320
rect 18305 -5360 18345 -5320
rect 18655 -5360 18695 -5320
rect 19005 -5360 19045 -5320
rect 19355 -5360 19395 -5320
rect 19705 -5360 19745 -5320
rect 15855 -5710 15895 -5670
rect 16205 -5710 16245 -5670
rect 16555 -5710 16595 -5670
rect 16905 -5710 16945 -5670
rect 17255 -5710 17295 -5670
rect 17605 -5710 17645 -5670
rect 17955 -5710 17995 -5670
rect 18305 -5710 18345 -5670
rect 18655 -5710 18695 -5670
rect 19005 -5710 19045 -5670
rect 19355 -5710 19395 -5670
rect 19705 -5710 19745 -5670
rect 15855 -6060 15895 -6020
rect 16205 -6060 16245 -6020
rect 16555 -6060 16595 -6020
rect 16905 -6060 16945 -6020
rect 17255 -6060 17295 -6020
rect 17605 -6060 17645 -6020
rect 17955 -6060 17995 -6020
rect 18305 -6060 18345 -6020
rect 18655 -6060 18695 -6020
rect 19005 -6060 19045 -6020
rect 19355 -6060 19395 -6020
rect 19705 -6060 19745 -6020
<< metal4 >>
rect 17250 -4260 17300 -4255
rect 17250 -4300 17255 -4260
rect 17295 -4300 17300 -4260
rect 16900 -4310 16950 -4305
rect 16900 -4350 16905 -4310
rect 16945 -4350 16950 -4310
rect 16900 -4615 16950 -4350
rect 15850 -4620 16950 -4615
rect 15850 -4660 15855 -4620
rect 15895 -4660 16205 -4620
rect 16245 -4660 16555 -4620
rect 16595 -4660 16905 -4620
rect 16945 -4660 16950 -4620
rect 15850 -4665 16950 -4660
rect 17250 -4615 17300 -4300
rect 18650 -4310 18700 -4305
rect 18650 -4350 18655 -4310
rect 18695 -4350 18700 -4310
rect 18650 -4615 18700 -4350
rect 17250 -4620 18350 -4615
rect 17250 -4660 17255 -4620
rect 17295 -4660 17605 -4620
rect 17645 -4660 17955 -4620
rect 17995 -4660 18305 -4620
rect 18345 -4660 18350 -4620
rect 17250 -4665 18350 -4660
rect 18650 -4620 19750 -4615
rect 18650 -4660 18655 -4620
rect 18695 -4660 19005 -4620
rect 19045 -4660 19355 -4620
rect 19395 -4660 19705 -4620
rect 19745 -4660 19750 -4620
rect 18650 -4665 19750 -4660
rect 16200 -4965 16250 -4665
rect 17950 -4965 18000 -4665
rect 19350 -4965 19400 -4665
rect 15850 -4970 16950 -4965
rect 15850 -5010 15855 -4970
rect 15895 -5010 16205 -4970
rect 16245 -5010 16555 -4970
rect 16595 -5010 16905 -4970
rect 16945 -5010 16950 -4970
rect 15850 -5015 16950 -5010
rect 17250 -4970 18350 -4965
rect 17250 -5010 17255 -4970
rect 17295 -5010 17605 -4970
rect 17645 -5010 17955 -4970
rect 17995 -5010 18305 -4970
rect 18345 -5010 18350 -4970
rect 17250 -5015 18350 -5010
rect 18650 -4970 19750 -4965
rect 18650 -5010 18655 -4970
rect 18695 -5010 19005 -4970
rect 19045 -5010 19355 -4970
rect 19395 -5010 19705 -4970
rect 19745 -5010 19750 -4970
rect 18650 -5015 19750 -5010
rect 16200 -5315 16250 -5015
rect 17950 -5315 18000 -5015
rect 19350 -5315 19400 -5015
rect 15850 -5320 16950 -5315
rect 15850 -5360 15855 -5320
rect 15895 -5360 16205 -5320
rect 16245 -5360 16555 -5320
rect 16595 -5360 16905 -5320
rect 16945 -5360 16950 -5320
rect 15850 -5365 16950 -5360
rect 17250 -5320 18350 -5315
rect 17250 -5360 17255 -5320
rect 17295 -5360 17605 -5320
rect 17645 -5360 17955 -5320
rect 17995 -5360 18305 -5320
rect 18345 -5360 18350 -5320
rect 17250 -5365 18350 -5360
rect 18650 -5320 19750 -5315
rect 18650 -5360 18655 -5320
rect 18695 -5360 19005 -5320
rect 19045 -5360 19355 -5320
rect 19395 -5360 19705 -5320
rect 19745 -5360 19750 -5320
rect 18650 -5365 19750 -5360
rect 16200 -5665 16250 -5365
rect 17950 -5665 18000 -5365
rect 19350 -5665 19400 -5365
rect 15850 -5670 16950 -5665
rect 15850 -5710 15855 -5670
rect 15895 -5710 16205 -5670
rect 16245 -5710 16555 -5670
rect 16595 -5710 16905 -5670
rect 16945 -5710 16950 -5670
rect 15850 -5715 16950 -5710
rect 17250 -5670 18350 -5665
rect 17250 -5710 17255 -5670
rect 17295 -5710 17605 -5670
rect 17645 -5710 17955 -5670
rect 17995 -5710 18305 -5670
rect 18345 -5710 18350 -5670
rect 17250 -5715 18350 -5710
rect 18650 -5670 19750 -5665
rect 18650 -5710 18655 -5670
rect 18695 -5710 19005 -5670
rect 19045 -5710 19355 -5670
rect 19395 -5710 19705 -5670
rect 19745 -5710 19750 -5670
rect 18650 -5715 19750 -5710
rect 16200 -6015 16250 -5715
rect 17950 -6015 18000 -5715
rect 19350 -6015 19400 -5715
rect 15850 -6020 16950 -6015
rect 15850 -6060 15855 -6020
rect 15895 -6060 16205 -6020
rect 16245 -6060 16555 -6020
rect 16595 -6060 16905 -6020
rect 16945 -6060 16950 -6020
rect 15850 -6065 16950 -6060
rect 17250 -6020 18350 -6015
rect 17250 -6060 17255 -6020
rect 17295 -6060 17605 -6020
rect 17645 -6060 17955 -6020
rect 17995 -6060 18305 -6020
rect 18345 -6060 18350 -6020
rect 17250 -6065 18350 -6060
rect 18650 -6020 19750 -6015
rect 18650 -6060 18655 -6020
rect 18695 -6060 19005 -6020
rect 19045 -6060 19355 -6020
rect 19395 -6060 19705 -6020
rect 19745 -6060 19750 -6020
rect 18650 -6065 19750 -6060
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 18145 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_18
timestamp 1723858470
transform 1 0 16785 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_19
timestamp 1723858470
transform 1 0 17465 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_20
timestamp 1723858470
transform 1 0 18145 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_21
timestamp 1723858470
transform 1 0 18145 0 1 -3455
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_22
timestamp 1723858470
transform 1 0 17465 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23
timestamp 1723858470
transform 1 0 17465 0 1 -3455
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_24
timestamp 1723858470
transform 1 0 16785 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25
timestamp 1723858470
transform 1 0 16785 0 1 -3455
box 0 0 670 670
<< labels >>
flabel metal2 15995 -4385 15995 -4385 5 FreeSans 400 0 0 -40 cap_res1
flabel metal3 19355 -4375 19355 -4375 7 FreeSans 400 180 -40 0 cap_res2
flabel via1 17800 1610 17800 1610 1 FreeSans 400 0 0 200 PFET_GATE_10uA
flabel metal2 16670 -435 16670 -435 1 FreeSans 400 0 0 80 Vin+
flabel metal1 19795 1795 19795 1795 1 FreeSans 240 0 0 80 V_CMFB_S4
port 9 n
flabel metal1 16960 1795 16960 1795 1 FreeSans 240 0 0 80 V_CMFB_S1
port 6 n
flabel metal1 18640 1795 18640 1795 1 FreeSans 240 0 0 80 V_CMFB_S3
port 3 n
flabel metal1 19280 1790 19280 1790 1 FreeSans 240 0 0 80 VB1_CUR_BIAS
port 4 n
flabel metal1 16125 1795 16125 1795 1 FreeSans 240 0 0 80 ERR_AMP_CUR_BIAS
port 7 n
flabel metal1 17750 1795 17750 1795 1 FreeSans 240 0 0 80 TAIL_CUR_MIR_BIAS
port 5 n
flabel metal1 15805 1795 15805 1795 1 FreeSans 240 0 0 80 V_CMFB_S2
port 10 n
flabel metal2 18980 -30 18980 -30 5 FreeSans 400 0 0 -40 V_mir2
flabel metal2 18030 -70 18030 -70 7 FreeSans 240 0 -120 0 1st_Vout_2
flabel metal2 16620 -30 16620 -30 5 FreeSans 400 0 0 -40 V_mir1
flabel metal2 17570 -70 17570 -70 3 FreeSans 240 0 120 0 1st_Vout_1
flabel metal2 18930 -435 18930 -435 1 FreeSans 400 0 0 80 V_CUR_REF_REG
flabel metal2 16665 -135 16665 -135 5 FreeSans 400 0 0 -80 Vin-
flabel metal2 17060 -545 17060 -545 3 FreeSans 400 0 200 0 V_p_1
flabel metal2 18580 -545 18580 -545 3 FreeSans 400 180 200 0 V_p_2
flabel metal1 19415 1790 19415 1790 7 FreeSans 240 0 -160 0 ERR_AMP_REF
port 2 w
flabel metal1 16040 1785 16040 1785 7 FreeSans 240 0 -160 0 VB2_CUR_BIAS
port 11 w
flabel metal1 16235 -915 16235 -915 3 FreeSans 400 0 200 0 START_UP
flabel metal1 18780 -1115 18780 -1115 3 FreeSans 400 0 200 0 START_UP_NFET1
flabel metal1 19560 1790 19560 1790 3 FreeSans 240 0 160 0 VB3_CUR_BIAS
port 8 e
flabel metal1 15890 -1300 15890 -1300 7 FreeSans 400 0 -200 0 NFET_GATE_10uA
flabel poly 18430 645 18430 645 5 FreeSans 400 0 0 -40 V_TOP
<< end >>
