v {xschem version=3.4.5 file_version=1.2
}
G {}
K {}
V {}
S {}
E {}
B 2 940 -2260 1700 -1780 {flags=graph
y1=-4e-05
y2=0.00017
ypos1=0
ypos2=2
divy=5
subdivy=1
unity=1
x1=0
x2=1e-06
divx=5
subdivx=1
xlabmag=1.0
ylabmag=1.0


dataset=0
unitx=1
logx=0
logy=0






color="11 6 5 9"
node="i(vmeas1)
i(vmeas2)
i(vmeas3)
\\"-i(vmeas4)\\""
linewidth_mult=4
}
B 2 2120 -2200 3480 -1540 {flags=graph
y1=0
y2=1.8
ypos1=0
ypos2=2
divy=5
subdivy=1
unity=1
x1=0
x2=1e-06
divx=5
subdivx=1
xlabmag=1.0
ylabmag=1.0


dataset=0
unitx=1
logx=0
logy=0








linewidth_mult=3







autoload=0
sim_type=tran
color="6 7"
node="f_ref
f_vco"}
B 2 2120 -810 3500 -130 {flags=graph
y1=0.15202008
y2=2.8885817
ypos1=0
ypos2=2
divy=5
subdivy=1
unity=1
x1=0
x2=1e-06
divx=5
subdivx=1
xlabmag=1.0
ylabmag=1.0


dataset=0
unitx=1
logx=0
logy=0








linewidth_mult=5





color="6 5"
node="up_pfd_b
down_pfd"}
B 2 2120 -1520 3500 -820 {flags=graph
y1=-0.028
y2=1.9
ypos1=0
ypos2=2
divy=5
subdivy=1
unity=1
x1=0
x2=1e-06
divx=5
subdivx=1
xlabmag=1.0
ylabmag=1.0


dataset=0
unitx=1
logx=0
logy=0








linewidth_mult=5

color="6 5"
node="up_pfd
down_pfd"}
B 2 2050 670 2820 1030 {flags=graph
y1=-0.093
y2=1.9
ypos1=0
ypos2=2
divy=5
subdivy=1
unity=1
x1=0
x2=1e-06
divx=5
subdivx=1
xlabmag=1.0
ylabmag=1.0


dataset=0
unitx=1
logx=0
logy=0








linewidth_mult=2




color="6 5"
node="up_input
down_input"}
B 2 2120 -2870 2970 -2210 {flags=graph
y1=-8.1e-05
y2=0.58
ypos1=0
ypos2=2
divy=5
subdivy=1
unity=1
x1=0
x2=1e-06
divx=5
subdivx=1
xlabmag=1.0
ylabmag=1.0


dataset=0
unitx=1
logx=0
logy=0








linewidth_mult=5



color=6
node=vout}
B 2 2050 0 2810 380 {flags=graph
y1=-0.029
y2=1.9
ypos1=0
ypos2=2
divy=5
subdivy=1
unity=1
x1=0
x2=1e-06
divx=5
subdivx=1
xlabmag=1.0
ylabmag=1.0


dataset=0
unitx=1
logx=0
logy=0








linewidth_mult=3



color="18 6 11 5 12"
node="opamp_out
up_input


down_gate
down_input


x"}
B 2 2050 400 2690 660 {flags=graph
y1=-0.038
y2=1.9
ypos1=0
ypos2=2
divy=5
subdivy=1
unity=1
x1=0
x2=1e-06
divx=5
subdivx=1
xlabmag=1.0
ylabmag=1.0


dataset=0
unitx=1
logx=0
logy=0








linewidth_mult=2


color="6 5"
node="up_b
down"}
B 2 940 -2760 1700 -2280 {flags=graph
y1=7.9969411e-05
y2=0.00018372516
ypos1=0
ypos2=2
divy=5
subdivy=1
unity=1
x1=0
x2=1e-06
divx=5
subdivx=1
xlabmag=1.0
ylabmag=1.0


dataset=0
unitx=1
logx=0
logy=0








linewidth_mult=4



color="5 6 11"
node="i(@m.xm1.msky130_fd_pr__nfet_01v8[id])
i(@m.xm2.msky130_fd_pr__nfet_01v8[id])
x"}
N 770 -220 900 -220 {
lab=DOWN_gate}
N 730 -190 730 -110 {
lab=GND}
N 730 -110 990 -110 {
lab=GND}
N 690 -220 730 -220 {
lab=GND}
N 690 -220 690 -110 {
lab=GND}
N 690 -110 730 -110 {
lab=GND}
N 940 -220 980 -220 {
lab=GND}
N 900 -1340 940 -1340 {
lab=VDD}
N 990 -110 1030 -110 {
lab=GND}
N 940 -1530 940 -1370 {
lab=VDD}
N 900 -1530 900 -1340 {
lab=VDD}
N 1590 -1530 1590 -1370 {
lab=VDD}
N 1410 -1530 1410 -1470 {
lab=VDD}
N 1410 -1440 1430 -1440 {
lab=VDD}
N 1430 -1530 1430 -1440 {
lab=VDD}
N 1610 -1530 1610 -1340 {
lab=VDD}
N 1590 -1340 1610 -1340 {
lab=VDD}
N 1590 -1310 1590 -1040 {
lab=Vout}
N 1440 -270 1550 -270 {
lab=DOWN_input}
N 1030 -110 1140 -110 {
lab=GND}
N 1140 -160 1140 -110 {
lab=GND}
N 1590 -390 1590 -300 {
lab=Vout}
N 1590 -240 1590 -110 {
lab=GND}
N 1140 -110 1590 -110 {
lab=GND}
N 1140 -190 1340 -190 {
lab=GND}
N 1340 -190 1340 -110 {
lab=GND}
N 1590 -270 1610 -270 {
lab=GND}
N 1610 -270 1610 -110 {
lab=GND}
N 1590 -110 1610 -110 {
lab=GND}
N 350 -1020 450 -1020 {
lab=UP_PFD_b}
N 390 -550 500 -550 {
lab=#net1}
N 90 -1020 130 -1020 {
lab=UP_PFD}
N 130 -550 170 -550 {
lab=DOWN_PFD}
N 1590 -980 1590 -450 {
lab=Vout}
N 940 -1310 940 -990 {
lab=x}
N 940 -870 1040 -870 {
lab=x}
N 1080 -870 1590 -870 {
lab=Vout}
N 1060 -1340 1060 -1000 {
lab=opamp_out}
N 1850 -490 1850 -440 {
lab=#net2}
N 1850 -870 1850 -550 {
lab=Vout}
N 1850 -380 1850 -320 {
lab=GND}
N 1800 -520 1830 -520 {
lab=GND}
N 1800 -520 1800 -350 {
lab=GND}
N 1800 -350 1850 -350 {
lab=GND}
N 1700 -870 1700 -550 {
lab=Vout}
N 1700 -490 1700 -430 {
lab=GND}
N 1420 140 1420 180 {
lab=F_REF}
N 1750 140 1750 180 {
lab=F_VCO}
N 880 -270 880 -220 {
lab=DOWN_gate}
N 1590 -870 1630 -870 {
lab=Vout}
N 1690 -870 1930 -870 {
lab=Vout}
N 810 -290 810 -220 {
lab=DOWN_gate}
N 730 -290 810 -290 {
lab=DOWN_gate}
N 980 -220 980 -110 {
lab=GND}
N 940 -190 940 -110 {
lab=GND}
N 880 -270 1380 -270 {
lab=DOWN_gate}
N 1460 -1530 1460 -1340 {
lab=VDD}
N 560 -550 1090 -550 {
lab=DOWN_b}
N 1460 -1300 1460 -1020 {
lab=UP_b}
N 1140 -1440 1370 -1440 {
lab=UP}
N 1140 -1440 1140 -1020 {
lab=UP}
N 1500 -1410 1500 -1340 {
lab=UP_input}
N 1410 -1410 1500 -1410 {
lab=UP_input}
N 1490 -1340 1550 -1340 {
lab=UP_input}
N 900 -1530 1610 -1530 {
lab=VDD}
N 1350 -550 1410 -550 {
lab=DOWN}
N 1410 -550 1410 -310 {
lab=DOWN}
N 1140 -220 1500 -220 {
lab=DOWN_input}
N 1500 -270 1500 -220 {
lab=DOWN_input}
N 1050 -550 1050 -190 {
lab=DOWN_b}
N 1050 -190 1100 -190 {
lab=DOWN_b}
N 1410 -270 1410 -110 {
lab=GND}
N 730 -1190 730 -250 {
lab=DOWN_gate}
N 940 -930 940 -250 {
lab=x}
N 1020 -1420 1020 -1340 {
lab=opamp_out}
N 1020 -1530 1020 -1480 {
lab=VDD}
N 1460 -1020 1520 -1020 {
lab=UP_b}
N 1500 -310 1500 -270 {
lab=DOWN_input}
N 1410 -370 1500 -370 {
lab=DOWN}
N 980 -1340 1430 -1340 {
lab=opamp_out}
N 500 -590 500 -510 {
lab=#net1}
N 560 -590 560 -510 {
lab=DOWN_b}
N 530 -670 530 -630 {
lab=VDD}
N 530 -520 530 -510 {
lab=VDD}
N 530 -520 570 -520 {
lab=VDD}
N 570 -640 570 -520 {
lab=VDD}
N 530 -640 570 -640 {
lab=VDD}
N 530 -590 530 -580 {
lab=GND}
N 490 -580 530 -580 {
lab=GND}
N 490 -580 490 -460 {
lab=GND}
N 490 -460 530 -460 {
lab=GND}
N 530 -470 530 -420 {
lab=GND}
N 290 -570 290 -530 {
lab=#net1}
N 220 -600 250 -600 {
lab=DOWN_PFD}
N 220 -600 220 -500 {
lab=DOWN_PFD}
N 220 -500 250 -500 {
lab=DOWN_PFD}
N 290 -550 390 -550 {
lab=#net1}
N 170 -550 220 -550 {
lab=DOWN_PFD}
N 290 -470 290 -430 {
lab=GND}
N 290 -670 290 -630 {
lab=VDD}
N 290 -600 320 -600 {
lab=VDD}
N 320 -650 320 -600 {
lab=VDD}
N 290 -650 320 -650 {
lab=VDD}
N 290 -500 320 -500 {
lab=GND}
N 320 -500 320 -450 {
lab=GND}
N 290 -450 320 -450 {
lab=GND}
N 250 -1040 250 -1000 {
lab=UP_PFD_b}
N 180 -1070 210 -1070 {
lab=UP_PFD}
N 180 -1070 180 -970 {
lab=UP_PFD}
N 180 -970 210 -970 {
lab=UP_PFD}
N 250 -1020 350 -1020 {
lab=UP_PFD_b}
N 130 -1020 180 -1020 {
lab=UP_PFD}
N 250 -940 250 -900 {
lab=GND}
N 250 -1140 250 -1100 {
lab=VDD}
N 250 -1070 280 -1070 {
lab=VDD}
N 280 -1120 280 -1070 {
lab=VDD}
N 250 -1120 280 -1120 {
lab=VDD}
N 250 -970 280 -970 {
lab=GND}
N 280 -970 280 -920 {
lab=GND}
N 250 -920 280 -920 {
lab=GND}
N 570 -1040 570 -1000 {
lab=UP}
N 500 -1070 530 -1070 {
lab=UP_PFD_b}
N 500 -1070 500 -970 {
lab=UP_PFD_b}
N 500 -970 530 -970 {
lab=UP_PFD_b}
N 450 -1020 500 -1020 {
lab=UP_PFD_b}
N 570 -940 570 -900 {
lab=GND}
N 570 -1140 570 -1100 {
lab=VDD}
N 570 -1070 600 -1070 {
lab=VDD}
N 600 -1120 600 -1070 {
lab=VDD}
N 570 -1120 600 -1120 {
lab=VDD}
N 570 -970 600 -970 {
lab=GND}
N 600 -970 600 -920 {
lab=GND}
N 570 -920 600 -920 {
lab=GND}
N 1210 -570 1210 -530 {
lab=DOWN}
N 1140 -600 1170 -600 {
lab=DOWN_b}
N 1140 -600 1140 -500 {
lab=DOWN_b}
N 1140 -500 1170 -500 {
lab=DOWN_b}
N 1090 -550 1140 -550 {
lab=DOWN_b}
N 1210 -470 1210 -430 {
lab=GND}
N 1210 -670 1210 -630 {
lab=VDD}
N 1210 -600 1240 -600 {
lab=VDD}
N 1240 -650 1240 -600 {
lab=VDD}
N 1210 -650 1240 -650 {
lab=VDD}
N 1210 -500 1240 -500 {
lab=GND}
N 1240 -500 1240 -450 {
lab=GND}
N 1210 -450 1240 -450 {
lab=GND}
N 1210 -550 1350 -550 {
lab=DOWN}
N 1260 -1040 1260 -1000 {
lab=UP_b}
N 1190 -1070 1220 -1070 {
lab=UP}
N 1190 -1070 1190 -970 {
lab=UP}
N 1190 -970 1220 -970 {
lab=UP}
N 1140 -1020 1190 -1020 {
lab=UP}
N 1260 -940 1260 -900 {
lab=GND}
N 1260 -1140 1260 -1100 {
lab=VDD}
N 1260 -1070 1290 -1070 {
lab=VDD}
N 1290 -1120 1290 -1070 {
lab=VDD}
N 1260 -1120 1290 -1120 {
lab=VDD}
N 1260 -970 1290 -970 {
lab=GND}
N 1290 -970 1290 -920 {
lab=GND}
N 1260 -920 1290 -920 {
lab=GND}
N 1260 -1020 1400 -1020 {
lab=UP_b}
N 1400 -1020 1460 -1020 {
lab=UP_b}
N 570 -1020 1140 -1020 {
lab=UP}
N 1520 -1080 1520 -1020 {
lab=UP_b}
N 1520 -1340 1520 -1140 {
lab=UP_input}
N 1750 310 1750 350 {
lab=DOWN_gate}
N 1590 -450 1590 -390 {
lab=Vout}
N 1630 -870 1690 -870 {
lab=Vout}
N 1590 -1040 1590 -980 {
lab=Vout}
N 940 -990 940 -930 {
lab=x}
C {sky130_fd_pr/nfet_01v8.sym} 750 -220 0 1 {name=M1
L=0.15
W=5
nf=5 
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=nfet_01v8
spiceprefix=X
}
C {sky130_fd_pr/nfet_01v8.sym} 920 -220 0 0 {name=M2
L=0.15
W=5
nf=5 
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=nfet_01v8
spiceprefix=X
}
C {sky130_fd_pr/pfet_01v8.sym} 960 -1340 2 0 {name=M3
L=0.15
W=10
nf=10
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=pfet_01v8
spiceprefix=X
}
C {devices/vdd.sym} 1060 -1530 0 0 {name=l13 lab=VDD}
C {devices/gnd.sym} 910 -110 0 0 {name=l14 lab=GND}
C {sky130_fd_pr/corner.sym} 730 130 0 0 {name=CORNER only_toplevel=false corner=tt}
C {devices/code.sym} 960 128.75 0 0 {name=STIMULI only_toplevel=false value="

.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

.option method=gear trtol1
.option wnflag=1
.option savecurrents

* .temp = 75

.ic v(vout) = 1.0

.save 
+v(up_pfd)
+v(down_pfd)
+v(up_pfd_b)
+v(down_pfd_b)
+v(up)
+v(up_b)
+v(down)
+v(down_b)
+v(v2)
+v(x)
+v(y)
+v(z)
+v(vout)
+v(up_input)
+v(down_input)
+v(down_gate)
+v(opamp_out)
+v(x2.p_bias)
+v(x2.n_bias)
+v(x2.v_common_p)
+v(x2.v_common_n)
+v(x2.p_left)
+v(x2.p_right)
+v(x2.n_left)
+v(x2.n_right)
+v(f_ref)
+v(f_vco)
+v(x4.qa)
+v(x4.qa_b)
+v(x4.qb)
+v(x4.qb_b)
+v(x4.qa)
+v(x4.e)
+v(x4.e_b)
+v(x4.f)
+v(x4.f_b)
+v(x4.before_reset)
+v(x4.reset)
+@m.xm6.msky130_fd_pr__pfet_01v8[id]
+@m.xm9.msky130_fd_pr__nfet_01v8[id]

.control
  let start_delay = 0ns
  let stop_delay = 24ns
  let index = -12
  dowhile start_delay <= stop_delay
    alter @V3[pulse] = [ 0 1.8 $&start_delay 1ns 1ns 24ns 50ns ]
    save @m.xm6.msky130_fd_pr__pfet_01v8[id] @m.xm9.msky130_fd_pr__nfet_01v8[id] v(F_REF) v(F_VCO) v(vout)
    tran 0.01ns 1us
    remzerovec
    linearize @m.xm6.msky130_fd_pr__pfet_01v8[id] @m.xm9.msky130_fd_pr__nfet_01v8[id] v(F_REF) v(F_VCO) v(vout)
    echo $&start_delay
    write pfd_charge_pump_dead_zone_check_2_\{$&index\}.raw
    wrdata /foss/designs/my_design/projects/pll/charge_pump/xschem_ngspice/pfd_charge_pump_dead_zone_check_2_\{$&index\}.txt @m.xm6.msky130_fd_pr__pfet_01v8[id] @m.xm9.msky130_fd_pr__nfet_01v8[id]
    set appendwrite
    reset
    let index = index + 1
    let start_delay = start_delay + 1ns
  end
.endc




"}
C {devices/vsource.sym} 1240 210 0 0 {name=V1 value=1.8 savecurrent=false}
C {devices/gnd.sym} 1240 240 0 0 {name=l2 lab=GND}
C {devices/lab_wire.sym} 940 -830 0 0 {name=p1 sig_type=std_logic lab=x}
C {devices/vdd.sym} 1240 180 0 1 {name=l3 lab=VDD}
C {sky130_fd_pr/pfet_01v8.sym} 1460 -1320 3 0 {name=M4
L=0.15
W=4
nf=4
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=pfet_01v8
spiceprefix=X
}
C {sky130_fd_pr/pfet_01v8.sym} 1390 -1440 0 0 {name=M5
L=0.15
W=5
nf=5
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=pfet_01v8
spiceprefix=X
}
C {sky130_fd_pr/pfet_01v8.sym} 1570 -1340 0 0 {name=M6
L=0.15
W=10
nf=10
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=pfet_01v8
spiceprefix=X
}
C {devices/lab_wire.sym} 1140 -1440 0 0 {name=p4 sig_type=std_logic lab=UP}
C {devices/lab_wire.sym} 1460 -1060 0 1 {name=p5 sig_type=std_logic lab=UP_b}
C {sky130_fd_pr/nfet_01v8.sym} 1410 -290 1 0 {name=M7
L=0.15
W=2
nf=2 
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=nfet_01v8
spiceprefix=X
}
C {sky130_fd_pr/nfet_01v8.sym} 1120 -190 0 0 {name=M8
L=0.15
W=2
nf=2 
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=nfet_01v8
spiceprefix=X
}
C {devices/lab_wire.sym} 1410 -500 0 1 {name=p6 sig_type=std_logic lab=DOWN}
C {devices/lab_wire.sym} 1050 -190 2 1 {name=p8 sig_type=std_logic lab=DOWN_b}
C {sky130_fd_pr/nfet_01v8.sym} 1570 -270 0 0 {name=M9
L=0.15
W=5
nf=5 
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=nfet_01v8
spiceprefix=X
}
C {devices/lab_wire.sym} 350 -1020 0 1 {name=p15 sig_type=std_logic lab=UP_PFD_b}
C {devices/lab_wire.sym} 1520 -1340 2 0 {name=p13 sig_type=std_logic lab=UP_input}
C {devices/lab_wire.sym} 1520 -270 0 0 {name=p14 sig_type=std_logic lab=DOWN_input}
C {devices/gnd.sym} 990 -930 0 1 {name=l7 lab=GND}
C {devices/lab_wire.sym} 1010 -1340 0 1 {name=p17 sig_type=std_logic lab=opamp_out}
C {devices/lab_wire.sym} 1930 -870 0 1 {name=p9 sig_type=std_logic lab=Vout}
C {devices/lab_wire.sym} 90 -1020 0 0 {name=p2 sig_type=std_logic lab=UP_PFD}
C {devices/lab_wire.sym} 130 -550 2 1 {name=p7 sig_type=std_logic lab=DOWN_PFD}
C {sky130_fd_pr/cap_mim_m3_1.sym} 1700 -520 0 0 {name=C2 model=cap_mim_m3_1 W=45 L=100 MF=1 spiceprefix=X}
C {sky130_fd_pr/cap_mim_m3_1.sym} 1850 -410 0 0 {name=C1 model=cap_mim_m3_1 W=230 L=100 MF=1 spiceprefix=X}
C {devices/gnd.sym} 1850 -320 0 0 {name=l4 lab=GND}
C {devices/gnd.sym} 1700 -430 0 0 {name=l9 lab=GND}
C {devices/vsource.sym} 1420 210 0 0 {name=V2 value="pulse(0 1.8 12ns 1ns 1ns 24ns 50ns)" savecurrent=false
}
C {devices/gnd.sym} 1420 240 0 0 {name=l10 lab=GND}
C {devices/lab_pin.sym} 1420 140 0 1 {name=p11 sig_type=std_logic lab=F_REF}
C {devices/vsource.sym} 1750 210 0 0 {name=V3 value="pulse(0 1.8 22ns 1ns 1ns 24ns 50ns)" savecurrent=false
* "sin(0.9 0.9 20.1MEG)" pulse(0 1.8 1ns 0.25ns 0.25ns 24.875ns 49.75ns)}
C {devices/gnd.sym} 1750 240 0 0 {name=l15 lab=GND}
C {devices/lab_pin.sym} 1750 140 0 1 {name=p12 sig_type=std_logic lab=F_VCO}
C {/foss/designs/my_design/projects/pll/pfd/xschem_ngspice/phase_frequency_detector.sym} 930 440 0 0 {name=x4}
C {devices/lab_pin.sym} 780 420 0 0 {name=p19 lab=F_REF}
C {devices/lab_pin.sym} 780 460 0 0 {name=p20 lab=F_VCO}
C {devices/lab_wire.sym} 1080 420 0 1 {name=p22 sig_type=std_logic lab=UP_PFD}
C {devices/lab_wire.sym} 1080 460 2 0 {name=p23 sig_type=std_logic lab=DOWN_PFD}
C {devices/vdd.sym} 930 380 0 1 {name=l1 lab=VDD}
C {devices/gnd.sym} 930 500 0 0 {name=l8 lab=GND}
C {devices/lab_wire.sym} 895 -270 0 0 {name=p10 sig_type=std_logic lab=DOWN_gate}
C {/foss/designs/my_design/projects/pll/charge_pump/xschem_ngspice/rail_to_rail_opamp3.sym} 1060 -930 1 1 {name=x2}
C {devices/vdd.sym} 1130 -930 0 0 {name=l6 lab=VDD}
C {sky130_fd_pr/res_xhigh_po_0p35.sym} 1850 -520 0 0 {name=R1
L=4
model=res_xhigh_po_0p35
spiceprefix=X
mult=1}
C {sky130_fd_pr/pfet_01v8.sym} 530 -490 3 0 {name=M12
L=0.15
W=2
nf=2
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=pfet_01v8
spiceprefix=X
}
C {sky130_fd_pr/nfet_01v8.sym} 530 -610 1 0 {name=M13
L=0.15
W=1
nf=1 
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=nfet_01v8
spiceprefix=X
}
C {devices/vdd.sym} 530 -670 0 0 {name=l11 lab=VDD}
C {devices/gnd.sym} 530 -420 0 0 {name=l12 lab=GND}
C {sky130_fd_pr/cap_mim_m3_1.sym} 1500 -340 0 0 {name=C3 model=cap_mim_m3_1 W=1 L=1 MF=1 spiceprefix=X}
C {sky130_fd_pr/cap_mim_m3_1.sym} 1520 -1110 0 0 {name=C4 model=cap_mim_m3_1 W=6 L=1 MF=1 spiceprefix=X}
C {sky130_fd_pr/cap_mim_m3_1.sym} 1020 -1450 0 0 {name=C5 model=cap_mim_m3_1 W=15 L=15 MF=1 spiceprefix=X}
C {sky130_fd_pr/pfet_01v8.sym} 270 -600 0 0 {name=M10
L=0.15
W=2
nf=2
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=pfet_01v8
spiceprefix=X
}
C {sky130_fd_pr/nfet_01v8.sym} 270 -500 2 1 {name=M11
L=0.15
W=1
nf=1 
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=nfet_01v8
spiceprefix=X
}
C {devices/gnd.sym} 290 -430 0 0 {name=l16 lab=GND}
C {devices/vdd.sym} 290 -670 0 0 {name=l17 lab=VDD}
C {sky130_fd_pr/pfet_01v8.sym} 230 -1070 0 0 {name=M14
L=0.15
W=2
nf=2
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=pfet_01v8
spiceprefix=X
}
C {sky130_fd_pr/nfet_01v8.sym} 230 -970 2 1 {name=M15
L=0.15
W=1
nf=1 
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=nfet_01v8
spiceprefix=X
}
C {devices/gnd.sym} 250 -900 0 0 {name=l18 lab=GND}
C {devices/vdd.sym} 250 -1140 0 0 {name=l19 lab=VDD}
C {sky130_fd_pr/pfet_01v8.sym} 550 -1070 0 0 {name=M16
L=0.15
W=2
nf=2
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=pfet_01v8
spiceprefix=X
}
C {sky130_fd_pr/nfet_01v8.sym} 550 -970 2 1 {name=M17
L=0.15
W=1
nf=1 
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=nfet_01v8
spiceprefix=X
}
C {devices/gnd.sym} 570 -900 0 0 {name=l20 lab=GND}
C {devices/vdd.sym} 570 -1140 0 0 {name=l21 lab=VDD}
C {sky130_fd_pr/pfet_01v8.sym} 1190 -600 0 0 {name=M18
L=0.15
W=2
nf=2
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=pfet_01v8
spiceprefix=X
}
C {sky130_fd_pr/nfet_01v8.sym} 1190 -500 2 1 {name=M19
L=0.15
W=1
nf=1 
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=nfet_01v8
spiceprefix=X
}
C {devices/gnd.sym} 1210 -430 0 0 {name=l22 lab=GND}
C {devices/vdd.sym} 1210 -670 0 0 {name=l23 lab=VDD}
C {sky130_fd_pr/pfet_01v8.sym} 1240 -1070 0 0 {name=M20
L=0.15
W=2
nf=2
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=pfet_01v8
spiceprefix=X
}
C {sky130_fd_pr/nfet_01v8.sym} 1240 -970 2 1 {name=M21
L=0.15
W=1
nf=1 
mult=1
ad="'int((nf+1)/2) * W/nf * 0.29'" 
pd="'2*int((nf+1)/2) * (W/nf + 0.29)'"
as="'int((nf+2)/2) * W/nf * 0.29'" 
ps="'2*int((nf+2)/2) * (W/nf + 0.29)'"
nrd="'0.29 / W'" nrs="'0.29 / W'"
sa=0 sb=0 sd=0
model=nfet_01v8
spiceprefix=X
}
C {devices/gnd.sym} 1260 -900 0 0 {name=l24 lab=GND}
C {devices/vdd.sym} 1260 -1140 0 0 {name=l25 lab=VDD}
C {devices/isource.sym} 1750 380 2 0 {name=I1 value=100u}
C {devices/gnd.sym} 1750 410 0 0 {name=l26 lab=GND}
C {devices/lab_pin.sym} 1750 310 2 1 {name=p3 sig_type=std_logic lab=DOWN_gate}
C {devices/lab_wire.sym} 730 -1190 0 1 {name=p16 sig_type=std_logic lab=DOWN_gate}
