* PEX produced on Sat Feb  1 12:18:14 PM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from TSPC_FF_ratioed_divide2_magic.ext - technology: sky130A

.subckt TSPC_FF_ratioed_divide2_magic
X0 VOUT.t1 C.t4 GNDA.t6 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X1 VOUT.t0 a_1250_n70.t3 VDDA.t5 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X2 C.t3 a_1250_n70.t4 GNDA.t10 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X3 C.t0 a_1580_n70.t2 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X4 a_1580_n70.t1 a_1250_n70.t5 a_1470_n70.t1 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X5 a_1250_n70.t1 VIN VDDA.t9 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X6 GNDA.t12 VIN a_1250_n70.t2 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X7 VDDA.t1 VOUT.t2 a_1580_n70.t0 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X8 GNDA.t8 a_1250_n70.t6 C.t2 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X9 GNDA.t4 a_1250_n70.t7 C.t1 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X10 a_1470_n70.t0 VOUT.t3 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X11 VDDA.t7 VIN a_1250_n70.t0 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
R0 C.n2 C.t0 721.4
R1 C.n1 C.t4 349.433
R2 C.t1 C.n2 276.733
R3 C.n1 C.n0 206.333
R4 C.n0 C.t2 48.0005
R5 C.n0 C.t3 48.0005
R6 C.n2 C.n1 48.0005
R7 GNDA.t3 GNDA.t2 4683.87
R8 GNDA GNDA.t5 3947.35
R9 GNDA.t5 GNDA.t7 1561.29
R10 GNDA.t7 GNDA.t9 1561.29
R11 GNDA.t9 GNDA.t3 1561.29
R12 GNDA.t2 GNDA.t0 1561.29
R13 GNDA.t0 GNDA.t11 1561.29
R14 GNDA GNDA.n2 195.262
R15 GNDA GNDA.n1 194.3
R16 GNDA GNDA.n0 194.3
R17 GNDA.n1 GNDA.t10 48.0005
R18 GNDA.n1 GNDA.t4 48.0005
R19 GNDA.n0 GNDA.t6 48.0005
R20 GNDA.n0 GNDA.t8 48.0005
R21 GNDA.n2 GNDA.t1 48.0005
R22 GNDA.n2 GNDA.t12 48.0005
R23 VOUT.t2 VOUT.t3 819.4
R24 VOUT.n0 VOUT.t0 663.801
R25 VOUT.n0 VOUT.t2 489.168
R26 VOUT.t1 VOUT.n0 340.733
R27 a_1250_n70.n5 a_1250_n70.t0 723.534
R28 a_1250_n70.n4 a_1250_n70.t1 723.534
R29 a_1250_n70.n0 a_1250_n70.t3 369.534
R30 a_1250_n70.n3 a_1250_n70.n2 366.856
R31 a_1250_n70.t2 a_1250_n70.n5 254.333
R32 a_1250_n70.n3 a_1250_n70.t5 190.123
R33 a_1250_n70.n4 a_1250_n70.n3 187.201
R34 a_1250_n70.n1 a_1250_n70.n0 176.733
R35 a_1250_n70.n2 a_1250_n70.n1 176.733
R36 a_1250_n70.n0 a_1250_n70.t6 112.468
R37 a_1250_n70.n2 a_1250_n70.t7 112.468
R38 a_1250_n70.n1 a_1250_n70.t4 112.468
R39 a_1250_n70.n5 a_1250_n70.n4 70.4005
R40 VDDA.t0 VDDA.t8 1130.95
R41 VDDA.n0 VDDA.t2 927.381
R42 VDDA.n1 VDDA.t5 667.62
R43 VDDA.n0 VDDA.t4 610.715
R44 VDDA VDDA.n2 594.301
R45 VDDA VDDA.n3 594.301
R46 VDDA.t2 VDDA.t0 497.62
R47 VDDA.t8 VDDA.t6 497.62
R48 VDDA.n1 VDDA.n0 373.781
R49 VDDA.n2 VDDA.t3 78.8005
R50 VDDA.n2 VDDA.t1 78.8005
R51 VDDA.n3 VDDA.t9 78.8005
R52 VDDA.n3 VDDA.t7 78.8005
R53 VDDA VDDA.n1 3.55124
R54 a_1580_n70.n0 a_1580_n70.t0 713.933
R55 a_1580_n70.n0 a_1580_n70.t2 314.233
R56 a_1580_n70.t1 a_1580_n70.n0 308.2
R57 a_1470_n70.t0 a_1470_n70.t1 96.0005
C0 VIN VDDA 0.125153f
C1 VIN GNDA 0.291288f
C2 VDDA GNDA 1.11299f
.ends

