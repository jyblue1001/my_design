* NGSPICE file created from opamp_6_6.ext - technology: sky130A

**.subckt opamp_6_6
X0 a_3420_n350# a_3000_310# w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X1 w_1980_260# a_3000_310# a_3420_n350# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X2 a_3420_n350# a_2280_n350# a_2150_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X3 a_3420_n350# a_4140_1066# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X4 a_2020_310# a_1980_n1180# w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X5 a_3420_n350# a_3000_310# w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X6 a_2280_n350# a_2020_n350# a_2150_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X7 w_1980_260# a_1980_n1180# a_2020_310# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X8 a_4140_1066# a_3000_310# a_2150_n350# sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X9 a_2150_n350# a_2280_n350# a_3420_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X10 a_2150_n350# a_2020_n350# a_2020_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X11 w_1980_260# a_1980_n1180# a_1980_n1180# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=1.25 ps=6 w=2.5 l=0.5
X12 a_2280_n350# a_1630_200# a_2020_310# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X13 a_2020_310# a_1470_530# a_2020_n350# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X14 a_2490_n1180# a_2490_n1180# a_2150_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=1.25 pd=6 as=0.625 ps=3 w=2.5 l=0.5
X15 w_1980_260# a_1980_n1180# a_2020_310# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X16 a_2020_n350# a_1470_530# a_2020_310# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X17 a_3420_n350# a_2280_n350# a_2150_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X18 a_1980_n1180# a_1980_n1180# w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X19 a_2020_310# a_1630_200# a_2280_n350# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X20 a_2020_n350# a_2020_n350# a_2150_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X21 a_2150_n350# a_2490_n1180# a_2740_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X22 a_2280_n350# a_4140_n1860# a_2150_n350# sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X23 a_2740_n350# a_1630_200# a_3000_310# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X24 a_2740_310# a_2740_310# w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X25 a_2020_310# a_1980_n1180# w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X26 a_3000_310# a_1630_200# a_2740_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X27 w_1980_260# a_2740_310# a_3000_310# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X28 a_2740_n350# a_2490_n1180# a_2150_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X29 a_2740_n350# a_1470_530# a_2740_310# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X30 a_3000_310# a_2740_310# w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X31 a_3420_n350# a_4140_n1860# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X32 a_1980_n1180# a_1980_n1180# w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0.625 ps=3 w=2.5 l=0.5
X33 w_1980_260# a_2740_310# a_2740_310# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X34 a_2150_n350# a_2280_n350# a_3420_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X35 a_1980_n1180# a_2490_n1180# a_2150_n350# sky130_fd_pr__res_xhigh_po_2p85 l=0.51
X36 w_1980_260# a_3000_310# a_3420_n350# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X37 w_1980_260# a_1980_n1180# a_1980_n1180# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X38 a_2150_n350# a_2020_n350# a_2280_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X39 a_2740_310# a_1470_530# a_2740_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X40 a_2150_n350# a_2490_n1180# a_2490_n1180# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=1.25 ps=6 w=2.5 l=0.5
.ends

