magic
tech sky130A
timestamp 1738350291
<< nwell >>
rect 605 195 1530 210
rect 1780 195 2095 210
rect 605 105 2095 195
<< nmos >>
rect 665 -35 680 15
rect 845 -35 860 15
rect 900 -35 915 15
rect 1025 -35 1040 15
rect 1080 -35 1095 15
rect 1135 -35 1150 15
rect 1190 -35 1205 15
rect 1425 -35 1440 15
rect 1480 -35 1495 15
rect 1535 -35 1550 15
rect 1660 -35 1675 15
rect 1715 -35 1730 15
rect 1770 -35 1785 15
rect 1825 -35 1840 15
rect 1965 -35 1980 15
<< pmos >>
rect 665 125 680 175
rect 720 125 735 175
rect 845 125 860 175
rect 900 125 915 175
rect 1125 125 1140 175
rect 1425 125 1440 175
rect 1480 125 1495 175
rect 1670 125 1685 175
rect 1725 125 1740 175
rect 1965 125 1980 175
rect 2020 125 2035 175
<< ndiff >>
rect 625 0 665 15
rect 625 -20 635 0
rect 655 -20 665 0
rect 625 -35 665 -20
rect 680 0 720 15
rect 680 -20 690 0
rect 710 -20 720 0
rect 680 -35 720 -20
rect 805 0 845 15
rect 805 -20 815 0
rect 835 -20 845 0
rect 805 -35 845 -20
rect 860 0 900 15
rect 860 -20 870 0
rect 890 -20 900 0
rect 860 -35 900 -20
rect 915 0 955 15
rect 915 -20 925 0
rect 945 -20 955 0
rect 915 -35 955 -20
rect 985 0 1025 15
rect 985 -20 995 0
rect 1015 -20 1025 0
rect 985 -35 1025 -20
rect 1040 0 1080 15
rect 1040 -20 1050 0
rect 1070 -20 1080 0
rect 1040 -35 1080 -20
rect 1095 0 1135 15
rect 1095 -20 1105 0
rect 1125 -20 1135 0
rect 1095 -35 1135 -20
rect 1150 0 1190 15
rect 1150 -20 1160 0
rect 1180 -20 1190 0
rect 1150 -35 1190 -20
rect 1205 0 1245 15
rect 1205 -20 1215 0
rect 1235 -20 1245 0
rect 1205 -35 1245 -20
rect 1385 0 1425 15
rect 1385 -20 1395 0
rect 1415 -20 1425 0
rect 1385 -35 1425 -20
rect 1440 0 1480 15
rect 1440 -20 1450 0
rect 1470 -20 1480 0
rect 1440 -35 1480 -20
rect 1495 0 1535 15
rect 1495 -20 1505 0
rect 1525 -20 1535 0
rect 1495 -35 1535 -20
rect 1550 0 1590 15
rect 1550 -20 1560 0
rect 1580 -20 1590 0
rect 1550 -35 1590 -20
rect 1620 0 1660 15
rect 1620 -20 1630 0
rect 1650 -20 1660 0
rect 1620 -35 1660 -20
rect 1675 0 1715 15
rect 1675 -20 1685 0
rect 1705 -20 1715 0
rect 1675 -35 1715 -20
rect 1730 0 1770 15
rect 1730 -20 1740 0
rect 1760 -20 1770 0
rect 1730 -35 1770 -20
rect 1785 0 1825 15
rect 1785 -20 1795 0
rect 1815 -20 1825 0
rect 1785 -35 1825 -20
rect 1840 0 1880 15
rect 1840 -20 1850 0
rect 1870 -20 1880 0
rect 1840 -35 1880 -20
rect 1925 0 1965 15
rect 1925 -20 1935 0
rect 1955 -20 1965 0
rect 1925 -35 1965 -20
rect 1980 0 2020 15
rect 1980 -20 1990 0
rect 2010 -20 2020 0
rect 1980 -35 2020 -20
<< pdiff >>
rect 625 160 665 175
rect 625 140 635 160
rect 655 140 665 160
rect 625 125 665 140
rect 680 160 720 175
rect 680 140 690 160
rect 710 140 720 160
rect 680 125 720 140
rect 735 160 775 175
rect 735 140 745 160
rect 765 140 775 160
rect 735 125 775 140
rect 805 160 845 175
rect 805 140 815 160
rect 835 140 845 160
rect 805 125 845 140
rect 860 160 900 175
rect 860 140 870 160
rect 890 140 900 160
rect 860 125 900 140
rect 915 160 955 175
rect 915 140 925 160
rect 945 140 955 160
rect 915 125 955 140
rect 1085 160 1125 175
rect 1085 140 1095 160
rect 1115 140 1125 160
rect 1085 125 1125 140
rect 1140 160 1180 175
rect 1140 140 1150 160
rect 1170 140 1180 160
rect 1140 125 1180 140
rect 1385 160 1425 175
rect 1385 140 1395 160
rect 1415 140 1425 160
rect 1385 125 1425 140
rect 1440 160 1480 175
rect 1440 140 1450 160
rect 1470 140 1480 160
rect 1440 125 1480 140
rect 1495 160 1535 175
rect 1495 140 1505 160
rect 1525 140 1535 160
rect 1495 125 1535 140
rect 1630 160 1670 175
rect 1630 140 1640 160
rect 1660 140 1670 160
rect 1630 125 1670 140
rect 1685 160 1725 175
rect 1685 140 1695 160
rect 1715 140 1725 160
rect 1685 125 1725 140
rect 1740 160 1780 175
rect 1740 140 1750 160
rect 1770 140 1780 160
rect 1740 125 1780 140
rect 1925 160 1965 175
rect 1925 140 1935 160
rect 1955 140 1965 160
rect 1925 125 1965 140
rect 1980 160 2020 175
rect 1980 140 1990 160
rect 2010 140 2020 160
rect 1980 125 2020 140
rect 2035 160 2075 175
rect 2035 140 2045 160
rect 2065 140 2075 160
rect 2035 125 2075 140
<< ndiffc >>
rect 635 -20 655 0
rect 690 -20 710 0
rect 815 -20 835 0
rect 870 -20 890 0
rect 925 -20 945 0
rect 995 -20 1015 0
rect 1050 -20 1070 0
rect 1105 -20 1125 0
rect 1160 -20 1180 0
rect 1215 -20 1235 0
rect 1395 -20 1415 0
rect 1450 -20 1470 0
rect 1505 -20 1525 0
rect 1560 -20 1580 0
rect 1630 -20 1650 0
rect 1685 -20 1705 0
rect 1740 -20 1760 0
rect 1795 -20 1815 0
rect 1850 -20 1870 0
rect 1935 -20 1955 0
rect 1990 -20 2010 0
<< pdiffc >>
rect 635 140 655 160
rect 690 140 710 160
rect 745 140 765 160
rect 815 140 835 160
rect 870 140 890 160
rect 925 140 945 160
rect 1095 140 1115 160
rect 1150 140 1170 160
rect 1395 140 1415 160
rect 1450 140 1470 160
rect 1505 140 1525 160
rect 1640 140 1660 160
rect 1695 140 1715 160
rect 1750 140 1770 160
rect 1935 140 1955 160
rect 1990 140 2010 160
rect 2045 140 2065 160
<< psubdiff >>
rect 765 0 805 15
rect 765 -20 775 0
rect 795 -20 805 0
rect 765 -35 805 -20
<< nsubdiff >>
rect 1045 160 1085 175
rect 1045 140 1055 160
rect 1075 140 1085 160
rect 1045 125 1085 140
<< psubdiffcont >>
rect 775 -20 795 0
<< nsubdiffcont >>
rect 1055 140 1075 160
<< poly >>
rect 1520 225 1560 235
rect 1520 210 1530 225
rect 1480 205 1530 210
rect 1550 205 1560 225
rect 665 185 735 200
rect 1480 195 1560 205
rect 665 175 680 185
rect 720 175 735 185
rect 845 175 860 190
rect 900 175 915 190
rect 1125 175 1140 190
rect 1425 175 1440 190
rect 1480 175 1495 195
rect 1670 175 1685 190
rect 1725 175 1740 190
rect 1965 175 1980 190
rect 2020 175 2035 190
rect 1230 160 1270 170
rect 1230 140 1240 160
rect 1260 145 1270 160
rect 1260 140 1375 145
rect 1230 130 1375 140
rect 665 70 680 125
rect 720 110 735 125
rect 605 55 680 70
rect 665 15 680 55
rect 705 60 745 70
rect 705 40 715 60
rect 735 40 745 60
rect 705 30 745 40
rect 845 15 860 125
rect 900 110 915 125
rect 900 100 990 110
rect 900 95 960 100
rect 950 80 960 95
rect 980 80 990 100
rect 950 70 990 80
rect 1125 105 1140 125
rect 1360 105 1375 130
rect 1425 105 1440 125
rect 1480 115 1495 125
rect 1575 120 1615 130
rect 1125 90 1295 105
rect 1360 90 1455 105
rect 1480 100 1550 115
rect 885 60 925 70
rect 885 40 895 60
rect 915 40 925 60
rect 1125 40 1140 90
rect 1175 60 1215 65
rect 1175 40 1185 60
rect 1205 40 1215 60
rect 885 30 1150 40
rect 1175 30 1215 40
rect 1280 45 1295 90
rect 1440 76 1455 90
rect 1370 60 1410 65
rect 1440 61 1495 76
rect 1370 45 1380 60
rect 1280 40 1380 45
rect 1400 40 1410 60
rect 1280 30 1440 40
rect 900 25 1150 30
rect 900 15 915 25
rect 1025 15 1040 25
rect 1080 15 1095 25
rect 1135 15 1150 25
rect 1190 15 1205 30
rect 1370 25 1440 30
rect 1425 15 1440 25
rect 1480 15 1495 61
rect 1535 15 1550 100
rect 1575 100 1585 120
rect 1605 110 1615 120
rect 1670 110 1685 125
rect 1605 100 1685 110
rect 1725 100 1740 125
rect 1965 115 1980 125
rect 2020 115 2035 125
rect 1575 95 1685 100
rect 1575 90 1615 95
rect 1715 80 1740 100
rect 1765 100 1805 110
rect 1765 80 1775 100
rect 1795 85 1805 100
rect 1965 100 2035 115
rect 1875 85 1915 95
rect 1795 80 1840 85
rect 1575 60 1615 65
rect 1575 40 1585 60
rect 1605 45 1615 60
rect 1715 45 1730 80
rect 1765 70 1840 80
rect 1605 40 1785 45
rect 1575 30 1785 40
rect 1660 15 1675 30
rect 1715 15 1730 30
rect 1770 15 1785 30
rect 1825 15 1840 70
rect 1875 65 1885 85
rect 1905 80 1915 85
rect 1965 80 1980 100
rect 1905 65 1980 80
rect 1875 55 1915 65
rect 1965 15 1980 65
rect 2010 65 2125 75
rect 2010 45 2020 65
rect 2040 60 2125 65
rect 2040 45 2050 60
rect 2010 35 2050 45
rect 665 -50 680 -35
rect 845 -75 860 -35
rect 900 -50 915 -35
rect 1025 -50 1040 -35
rect 1080 -50 1095 -35
rect 1135 -50 1150 -35
rect 1190 -50 1205 -35
rect 1425 -50 1440 -35
rect 1480 -50 1495 -35
rect 1535 -50 1550 -35
rect 1660 -50 1675 -35
rect 1715 -50 1730 -35
rect 1770 -50 1785 -35
rect 1825 -50 1840 -35
rect 1965 -50 1980 -35
rect 2035 -75 2050 35
rect 845 -90 2050 -75
<< polycont >>
rect 1530 205 1550 225
rect 1240 140 1260 160
rect 715 40 735 60
rect 960 80 980 100
rect 895 40 915 60
rect 1185 40 1205 60
rect 1380 40 1400 60
rect 1585 100 1605 120
rect 1775 80 1795 100
rect 1585 40 1605 60
rect 1885 65 1905 85
rect 2020 45 2040 65
<< locali >>
rect 1520 225 1560 235
rect 1520 205 1530 225
rect 1550 215 1560 225
rect 1550 205 1770 215
rect 1520 195 1770 205
rect 1750 170 1770 195
rect 630 160 660 170
rect 630 140 635 160
rect 655 140 660 160
rect 630 130 660 140
rect 685 160 715 170
rect 685 140 690 160
rect 710 140 715 160
rect 685 130 715 140
rect 740 160 770 170
rect 740 140 745 160
rect 765 140 770 160
rect 740 130 770 140
rect 810 160 840 170
rect 810 140 815 160
rect 835 140 840 160
rect 810 130 840 140
rect 865 160 895 170
rect 865 140 870 160
rect 890 140 895 160
rect 865 130 895 140
rect 920 160 1030 170
rect 920 140 925 160
rect 945 150 1030 160
rect 945 140 950 150
rect 920 130 950 140
rect 695 70 715 130
rect 815 110 835 130
rect 815 100 990 110
rect 815 90 960 100
rect 950 80 960 90
rect 980 80 990 100
rect 950 70 990 80
rect 695 60 745 70
rect 695 40 715 60
rect 735 50 745 60
rect 885 60 925 70
rect 885 50 895 60
rect 735 40 895 50
rect 915 40 925 60
rect 695 30 925 40
rect 695 10 715 30
rect 950 10 970 70
rect 1010 50 1030 150
rect 1050 160 1120 170
rect 1050 140 1055 160
rect 1075 140 1095 160
rect 1115 140 1120 160
rect 1050 130 1120 140
rect 1145 160 1175 170
rect 1230 160 1270 170
rect 1390 160 1420 170
rect 1145 140 1150 160
rect 1170 140 1240 160
rect 1260 140 1270 160
rect 1145 130 1175 140
rect 1230 130 1270 140
rect 1330 140 1395 160
rect 1415 140 1420 160
rect 1175 60 1215 65
rect 1175 50 1185 60
rect 995 40 1185 50
rect 1205 40 1215 60
rect 995 30 1215 40
rect 995 10 1015 30
rect 1105 10 1125 30
rect 1240 10 1260 130
rect 630 0 660 10
rect 630 -20 635 0
rect 655 -20 660 0
rect 630 -30 660 -20
rect 685 0 715 10
rect 685 -20 690 0
rect 710 -20 715 0
rect 685 -30 715 -20
rect 770 0 840 10
rect 770 -20 775 0
rect 795 -20 815 0
rect 835 -20 840 0
rect 770 -30 840 -20
rect 865 0 895 10
rect 865 -20 870 0
rect 890 -20 895 0
rect 865 -30 895 -20
rect 920 0 970 10
rect 920 -20 925 0
rect 945 -10 970 0
rect 990 0 1020 10
rect 945 -20 950 -10
rect 920 -30 950 -20
rect 990 -20 995 0
rect 1015 -20 1020 0
rect 990 -30 1020 -20
rect 1045 0 1075 10
rect 1045 -20 1050 0
rect 1070 -20 1075 0
rect 1045 -30 1075 -20
rect 1100 0 1130 10
rect 1100 -20 1105 0
rect 1125 -20 1130 0
rect 1100 -30 1130 -20
rect 1155 0 1185 10
rect 1155 -20 1160 0
rect 1180 -20 1185 0
rect 1155 -30 1185 -20
rect 1210 0 1260 10
rect 1210 -20 1215 0
rect 1235 -20 1260 0
rect 1330 0 1350 140
rect 1390 130 1420 140
rect 1445 160 1475 170
rect 1445 140 1450 160
rect 1470 140 1475 160
rect 1445 130 1475 140
rect 1500 160 1530 170
rect 1500 140 1505 160
rect 1525 140 1530 160
rect 1500 130 1530 140
rect 1635 160 1665 170
rect 1635 140 1640 160
rect 1660 140 1665 160
rect 1635 130 1665 140
rect 1690 160 1720 170
rect 1690 140 1695 160
rect 1715 140 1720 160
rect 1690 130 1720 140
rect 1745 160 1775 170
rect 1930 160 1960 170
rect 1745 140 1750 160
rect 1770 140 1875 160
rect 1745 130 1775 140
rect 1395 110 1415 130
rect 1505 110 1525 130
rect 1575 120 1615 130
rect 1575 110 1585 120
rect 1395 100 1585 110
rect 1605 100 1615 120
rect 1395 90 1615 100
rect 1370 60 1410 65
rect 1575 60 1615 65
rect 1370 40 1380 60
rect 1400 40 1585 60
rect 1605 40 1615 60
rect 1645 50 1665 130
rect 1765 100 1805 110
rect 1765 80 1775 100
rect 1795 80 1805 100
rect 1765 70 1805 80
rect 1855 95 1875 140
rect 1930 140 1935 160
rect 1955 140 1960 160
rect 1930 130 1960 140
rect 1985 160 2015 170
rect 1985 140 1990 160
rect 2010 140 2015 160
rect 1985 130 2015 140
rect 2040 160 2070 170
rect 2040 140 2045 160
rect 2065 140 2070 160
rect 2040 130 2070 140
rect 1855 85 1915 95
rect 1765 50 1785 70
rect 1370 30 1410 40
rect 1575 30 1615 40
rect 1635 30 1785 50
rect 1855 65 1885 85
rect 1905 65 1915 85
rect 1855 55 1915 65
rect 1990 75 2010 130
rect 1990 65 2050 75
rect 1635 10 1655 30
rect 1745 10 1765 30
rect 1855 10 1875 55
rect 1990 45 2020 65
rect 2040 45 2050 65
rect 1990 35 2050 45
rect 1990 10 2010 35
rect 1390 0 1420 10
rect 1330 -20 1395 0
rect 1415 -20 1420 0
rect 1210 -30 1240 -20
rect 1390 -30 1420 -20
rect 1445 0 1475 10
rect 1445 -20 1450 0
rect 1470 -20 1475 0
rect 1445 -30 1475 -20
rect 1500 0 1530 10
rect 1500 -20 1505 0
rect 1525 -20 1530 0
rect 1500 -30 1530 -20
rect 1555 0 1585 10
rect 1555 -20 1560 0
rect 1580 -20 1585 0
rect 1555 -30 1585 -20
rect 1625 0 1655 10
rect 1625 -20 1630 0
rect 1650 -20 1655 0
rect 1625 -30 1655 -20
rect 1680 0 1710 10
rect 1680 -20 1685 0
rect 1705 -20 1710 0
rect 1680 -30 1710 -20
rect 1735 0 1765 10
rect 1735 -20 1740 0
rect 1760 -20 1765 0
rect 1735 -30 1765 -20
rect 1790 0 1820 10
rect 1790 -20 1795 0
rect 1815 -20 1820 0
rect 1790 -30 1820 -20
rect 1845 0 1875 10
rect 1845 -20 1850 0
rect 1870 -20 1875 0
rect 1845 -30 1875 -20
rect 1930 0 1960 10
rect 1930 -20 1935 0
rect 1955 -20 1960 0
rect 1930 -30 1960 -20
rect 1985 0 2015 10
rect 1985 -20 1990 0
rect 2010 -20 2015 0
rect 1985 -30 2015 -20
<< viali >>
rect 635 140 655 160
rect 745 140 765 160
rect 870 140 890 160
rect 1055 140 1075 160
rect 1095 140 1115 160
rect 635 -20 655 0
rect 775 -20 795 0
rect 815 -20 835 0
rect 1050 -20 1070 0
rect 1160 -20 1180 0
rect 1450 140 1470 160
rect 1695 140 1715 160
rect 1935 140 1955 160
rect 2045 140 2065 160
rect 1560 -20 1580 0
rect 1685 -20 1705 0
rect 1795 -20 1815 0
rect 1935 -20 1955 0
<< metal1 >>
rect 605 160 2095 175
rect 605 140 635 160
rect 655 140 745 160
rect 765 140 870 160
rect 890 140 1055 160
rect 1075 140 1095 160
rect 1115 140 1450 160
rect 1470 140 1695 160
rect 1715 140 1935 160
rect 1955 140 2045 160
rect 2065 140 2095 160
rect 605 125 2095 140
rect 605 0 2095 15
rect 605 -20 635 0
rect 655 -20 775 0
rect 795 -20 815 0
rect 835 -20 1050 0
rect 1070 -20 1160 0
rect 1180 -20 1560 0
rect 1580 -20 1685 0
rect 1705 -20 1795 0
rect 1815 -20 1935 0
rect 1955 -20 2095 0
rect 605 -35 2095 -20
<< labels >>
flabel locali 1030 80 1030 80 3 FreeSans 160 0 80 0 C
flabel locali 815 90 815 90 5 FreeSans 160 0 0 0 A
flabel locali 760 50 760 50 1 FreeSans 160 0 0 80 CLK
flabel poly 605 60 605 60 7 FreeSans 160 0 -80 0 VIN
flabel metal1 605 -10 605 -10 7 FreeSans 160 0 -80 0 GNDA
flabel metal1 605 150 605 150 7 FreeSans 160 0 -80 0 VDDA
flabel ndiff 880 -35 880 -35 5 FreeSans 160 0 0 -80 B
flabel locali 1330 160 1330 160 7 FreeSans 160 0 -80 0 E
flabel locali 1460 -30 1460 -30 5 FreeSans 160 0 0 -80 F
flabel locali 1515 -30 1515 -30 5 FreeSans 160 0 0 -80 G
flabel locali 1665 70 1665 70 3 FreeSans 160 0 80 0 H
flabel locali 1875 160 1875 160 3 FreeSans 160 0 80 0 I
flabel poly 2125 70 2125 70 3 FreeSans 160 0 80 0 VOUT
<< end >>
