magic
tech sky130A
timestamp 1753013163
<< nwell >>
rect 16750 1180 17240 1320
rect 17390 1180 18210 1320
rect 18360 1180 18850 1320
rect 16375 580 16755 720
rect 16910 470 18690 810
rect 18840 580 19220 720
rect 16360 -70 17725 70
rect 17875 -70 19240 70
<< pwell >>
rect 17780 -4300 17820 -4120
<< nmos >>
rect 16890 -500 16910 -450
rect 16950 -500 16970 -450
rect 17010 -500 17030 -450
rect 17070 -500 17090 -450
rect 17130 -500 17150 -450
rect 17190 -500 17210 -450
rect 17250 -500 17270 -450
rect 17310 -500 17330 -450
rect 17370 -500 17390 -450
rect 17430 -500 17450 -450
rect 18150 -500 18170 -450
rect 18210 -500 18230 -450
rect 18270 -500 18290 -450
rect 18330 -500 18350 -450
rect 18390 -500 18410 -450
rect 18450 -500 18470 -450
rect 18510 -500 18530 -450
rect 18570 -500 18590 -450
rect 18630 -500 18650 -450
rect 18690 -500 18710 -450
rect 16570 -975 17070 -725
rect 17190 -975 17690 -725
rect 17910 -975 18410 -725
rect 18530 -975 19030 -725
rect 16780 -1245 17780 -1145
rect 17820 -1245 18820 -1145
rect 16955 -1585 16970 -1485
rect 17010 -1585 17025 -1485
rect 17065 -1585 17080 -1485
rect 17120 -1585 17135 -1485
rect 17175 -1585 17190 -1485
rect 17230 -1585 17245 -1485
rect 17285 -1585 17300 -1485
rect 17340 -1585 17355 -1485
rect 17545 -1585 17560 -1485
rect 17600 -1585 17615 -1485
rect 17655 -1585 17670 -1485
rect 17710 -1585 17725 -1485
rect 17765 -1585 17780 -1485
rect 17820 -1585 17835 -1485
rect 17875 -1585 17890 -1485
rect 17930 -1585 17945 -1485
rect 17985 -1585 18000 -1485
rect 18040 -1585 18055 -1485
rect 18255 -1585 18270 -1485
rect 18310 -1585 18325 -1485
rect 18365 -1585 18380 -1485
rect 18420 -1585 18435 -1485
rect 18475 -1585 18490 -1485
rect 18530 -1585 18545 -1485
rect 18585 -1585 18600 -1485
rect 18640 -1585 18655 -1485
<< pmos >>
rect 16850 1200 16865 1300
rect 16905 1200 16920 1300
rect 16960 1200 16975 1300
rect 17015 1200 17030 1300
rect 17070 1200 17085 1300
rect 17125 1200 17140 1300
rect 17490 1200 17505 1300
rect 17545 1200 17560 1300
rect 17600 1200 17615 1300
rect 17655 1200 17670 1300
rect 17710 1200 17725 1300
rect 17765 1200 17780 1300
rect 17820 1200 17835 1300
rect 17875 1200 17890 1300
rect 17930 1200 17945 1300
rect 17985 1200 18000 1300
rect 18040 1200 18055 1300
rect 18095 1200 18110 1300
rect 18460 1200 18475 1300
rect 18515 1200 18530 1300
rect 18570 1200 18585 1300
rect 18625 1200 18640 1300
rect 18680 1200 18695 1300
rect 18735 1200 18750 1300
rect 16475 600 16490 700
rect 16530 600 16545 700
rect 16585 600 16600 700
rect 16640 600 16655 700
rect 17010 490 17060 790
rect 17100 490 17150 790
rect 17190 490 17240 790
rect 17280 490 17330 790
rect 17370 490 17420 790
rect 17460 490 17510 790
rect 17550 490 17600 790
rect 17640 490 17690 790
rect 17730 490 17780 790
rect 17820 490 17870 790
rect 17910 490 17960 790
rect 18000 490 18050 790
rect 18090 490 18140 790
rect 18180 490 18230 790
rect 18270 490 18320 790
rect 18360 490 18410 790
rect 18450 490 18500 790
rect 18540 490 18590 790
rect 18940 600 18955 700
rect 18995 600 19010 700
rect 19050 600 19065 700
rect 19105 600 19120 700
rect 16460 -50 16480 50
rect 16520 -50 16540 50
rect 16580 -50 16600 50
rect 16640 -50 16660 50
rect 16700 -50 16720 50
rect 16760 -50 16780 50
rect 16820 -50 16840 50
rect 16880 -50 16900 50
rect 16940 -50 16960 50
rect 17000 -50 17020 50
rect 17060 -50 17080 50
rect 17120 -50 17140 50
rect 17180 -50 17200 50
rect 17240 -50 17260 50
rect 17300 -50 17320 50
rect 17360 -50 17380 50
rect 17420 -50 17440 50
rect 17480 -50 17500 50
rect 17540 -50 17560 50
rect 17600 -50 17620 50
rect 17980 -50 18000 50
rect 18040 -50 18060 50
rect 18100 -50 18120 50
rect 18160 -50 18180 50
rect 18220 -50 18240 50
rect 18280 -50 18300 50
rect 18340 -50 18360 50
rect 18400 -50 18420 50
rect 18460 -50 18480 50
rect 18520 -50 18540 50
rect 18580 -50 18600 50
rect 18640 -50 18660 50
rect 18700 -50 18720 50
rect 18760 -50 18780 50
rect 18820 -50 18840 50
rect 18880 -50 18900 50
rect 18940 -50 18960 50
rect 19000 -50 19020 50
rect 19060 -50 19080 50
rect 19120 -50 19140 50
<< ndiff >>
rect 16850 -465 16890 -450
rect 16850 -485 16860 -465
rect 16880 -485 16890 -465
rect 16850 -500 16890 -485
rect 16910 -465 16950 -450
rect 16910 -485 16920 -465
rect 16940 -485 16950 -465
rect 16910 -500 16950 -485
rect 16970 -465 17010 -450
rect 16970 -485 16980 -465
rect 17000 -485 17010 -465
rect 16970 -500 17010 -485
rect 17030 -465 17070 -450
rect 17030 -485 17040 -465
rect 17060 -485 17070 -465
rect 17030 -500 17070 -485
rect 17090 -465 17130 -450
rect 17090 -485 17100 -465
rect 17120 -485 17130 -465
rect 17090 -500 17130 -485
rect 17150 -465 17190 -450
rect 17150 -485 17160 -465
rect 17180 -485 17190 -465
rect 17150 -500 17190 -485
rect 17210 -465 17250 -450
rect 17210 -485 17220 -465
rect 17240 -485 17250 -465
rect 17210 -500 17250 -485
rect 17270 -465 17310 -450
rect 17270 -485 17280 -465
rect 17300 -485 17310 -465
rect 17270 -500 17310 -485
rect 17330 -465 17370 -450
rect 17330 -485 17340 -465
rect 17360 -485 17370 -465
rect 17330 -500 17370 -485
rect 17390 -465 17430 -450
rect 17390 -485 17400 -465
rect 17420 -485 17430 -465
rect 17390 -500 17430 -485
rect 17450 -465 17490 -450
rect 17450 -485 17460 -465
rect 17480 -485 17490 -465
rect 17450 -500 17490 -485
rect 18110 -465 18150 -450
rect 18110 -485 18120 -465
rect 18140 -485 18150 -465
rect 18110 -500 18150 -485
rect 18170 -465 18210 -450
rect 18170 -485 18180 -465
rect 18200 -485 18210 -465
rect 18170 -500 18210 -485
rect 18230 -465 18270 -450
rect 18230 -485 18240 -465
rect 18260 -485 18270 -465
rect 18230 -500 18270 -485
rect 18290 -465 18330 -450
rect 18290 -485 18300 -465
rect 18320 -485 18330 -465
rect 18290 -500 18330 -485
rect 18350 -465 18390 -450
rect 18350 -485 18360 -465
rect 18380 -485 18390 -465
rect 18350 -500 18390 -485
rect 18410 -465 18450 -450
rect 18410 -485 18420 -465
rect 18440 -485 18450 -465
rect 18410 -500 18450 -485
rect 18470 -465 18510 -450
rect 18470 -485 18480 -465
rect 18500 -485 18510 -465
rect 18470 -500 18510 -485
rect 18530 -465 18570 -450
rect 18530 -485 18540 -465
rect 18560 -485 18570 -465
rect 18530 -500 18570 -485
rect 18590 -465 18630 -450
rect 18590 -485 18600 -465
rect 18620 -485 18630 -465
rect 18590 -500 18630 -485
rect 18650 -465 18690 -450
rect 18650 -485 18660 -465
rect 18680 -485 18690 -465
rect 18650 -500 18690 -485
rect 18710 -465 18750 -450
rect 18710 -485 18720 -465
rect 18740 -485 18750 -465
rect 18710 -500 18750 -485
rect 16530 -740 16570 -725
rect 16530 -960 16540 -740
rect 16560 -960 16570 -740
rect 16530 -975 16570 -960
rect 17070 -740 17110 -725
rect 17150 -740 17190 -725
rect 17070 -960 17080 -740
rect 17100 -960 17110 -740
rect 17150 -960 17160 -740
rect 17180 -960 17190 -740
rect 17070 -970 17110 -960
rect 17150 -970 17190 -960
rect 17070 -975 17190 -970
rect 17690 -740 17730 -725
rect 17690 -960 17700 -740
rect 17720 -960 17730 -740
rect 17690 -975 17730 -960
rect 17870 -740 17910 -725
rect 17870 -960 17880 -740
rect 17900 -960 17910 -740
rect 17870 -975 17910 -960
rect 18410 -740 18450 -725
rect 18490 -740 18530 -725
rect 18410 -960 18420 -740
rect 18440 -960 18450 -740
rect 18490 -960 18500 -740
rect 18520 -960 18530 -740
rect 18410 -975 18450 -960
rect 18490 -975 18530 -960
rect 19030 -740 19070 -725
rect 19030 -960 19040 -740
rect 19060 -960 19070 -740
rect 19030 -975 19070 -960
rect 16740 -1160 16780 -1145
rect 16740 -1230 16750 -1160
rect 16770 -1230 16780 -1160
rect 16740 -1245 16780 -1230
rect 17780 -1160 17820 -1145
rect 17780 -1230 17790 -1160
rect 17810 -1230 17820 -1160
rect 17780 -1245 17820 -1230
rect 18820 -1160 18860 -1145
rect 18820 -1230 18830 -1160
rect 18850 -1230 18860 -1160
rect 18820 -1245 18860 -1230
rect 16915 -1500 16955 -1485
rect 16915 -1570 16925 -1500
rect 16945 -1570 16955 -1500
rect 16915 -1585 16955 -1570
rect 16970 -1500 17010 -1485
rect 16970 -1570 16980 -1500
rect 17000 -1570 17010 -1500
rect 16970 -1585 17010 -1570
rect 17025 -1500 17065 -1485
rect 17025 -1570 17035 -1500
rect 17055 -1570 17065 -1500
rect 17025 -1585 17065 -1570
rect 17080 -1500 17120 -1485
rect 17080 -1570 17090 -1500
rect 17110 -1570 17120 -1500
rect 17080 -1585 17120 -1570
rect 17135 -1500 17175 -1485
rect 17135 -1570 17145 -1500
rect 17165 -1570 17175 -1500
rect 17135 -1585 17175 -1570
rect 17190 -1500 17230 -1485
rect 17190 -1570 17200 -1500
rect 17220 -1570 17230 -1500
rect 17190 -1585 17230 -1570
rect 17245 -1500 17285 -1485
rect 17245 -1570 17255 -1500
rect 17275 -1570 17285 -1500
rect 17245 -1585 17285 -1570
rect 17300 -1500 17340 -1485
rect 17300 -1570 17310 -1500
rect 17330 -1570 17340 -1500
rect 17300 -1585 17340 -1570
rect 17355 -1500 17395 -1485
rect 17355 -1570 17365 -1500
rect 17385 -1570 17395 -1500
rect 17355 -1585 17395 -1570
rect 17505 -1500 17545 -1485
rect 17505 -1570 17515 -1500
rect 17535 -1570 17545 -1500
rect 17505 -1585 17545 -1570
rect 17560 -1500 17600 -1485
rect 17560 -1570 17570 -1500
rect 17590 -1570 17600 -1500
rect 17560 -1585 17600 -1570
rect 17615 -1500 17655 -1485
rect 17615 -1570 17625 -1500
rect 17645 -1570 17655 -1500
rect 17615 -1585 17655 -1570
rect 17670 -1500 17710 -1485
rect 17670 -1570 17680 -1500
rect 17700 -1570 17710 -1500
rect 17670 -1585 17710 -1570
rect 17725 -1500 17765 -1485
rect 17725 -1570 17735 -1500
rect 17755 -1570 17765 -1500
rect 17725 -1585 17765 -1570
rect 17780 -1500 17820 -1485
rect 17780 -1570 17790 -1500
rect 17810 -1570 17820 -1500
rect 17780 -1585 17820 -1570
rect 17835 -1500 17875 -1485
rect 17835 -1570 17845 -1500
rect 17865 -1570 17875 -1500
rect 17835 -1585 17875 -1570
rect 17890 -1500 17930 -1485
rect 17890 -1570 17900 -1500
rect 17920 -1570 17930 -1500
rect 17890 -1585 17930 -1570
rect 17945 -1500 17985 -1485
rect 17945 -1570 17955 -1500
rect 17975 -1570 17985 -1500
rect 17945 -1585 17985 -1570
rect 18000 -1500 18040 -1485
rect 18000 -1570 18010 -1500
rect 18030 -1570 18040 -1500
rect 18000 -1585 18040 -1570
rect 18055 -1500 18095 -1485
rect 18055 -1570 18065 -1500
rect 18085 -1570 18095 -1500
rect 18055 -1585 18095 -1570
rect 18215 -1500 18255 -1485
rect 18215 -1570 18225 -1500
rect 18245 -1570 18255 -1500
rect 18215 -1585 18255 -1570
rect 18270 -1500 18310 -1485
rect 18270 -1570 18280 -1500
rect 18300 -1570 18310 -1500
rect 18270 -1585 18310 -1570
rect 18325 -1500 18365 -1485
rect 18325 -1570 18335 -1500
rect 18355 -1570 18365 -1500
rect 18325 -1585 18365 -1570
rect 18380 -1500 18420 -1485
rect 18380 -1570 18390 -1500
rect 18410 -1570 18420 -1500
rect 18380 -1585 18420 -1570
rect 18435 -1500 18475 -1485
rect 18435 -1570 18445 -1500
rect 18465 -1570 18475 -1500
rect 18435 -1585 18475 -1570
rect 18490 -1500 18530 -1485
rect 18490 -1570 18500 -1500
rect 18520 -1570 18530 -1500
rect 18490 -1585 18530 -1570
rect 18545 -1500 18585 -1485
rect 18545 -1570 18555 -1500
rect 18575 -1570 18585 -1500
rect 18545 -1585 18585 -1570
rect 18600 -1500 18640 -1485
rect 18600 -1570 18610 -1500
rect 18630 -1570 18640 -1500
rect 18600 -1585 18640 -1570
rect 18655 -1500 18695 -1485
rect 18655 -1570 18665 -1500
rect 18685 -1570 18695 -1500
rect 18655 -1585 18695 -1570
<< pdiff >>
rect 16810 1285 16850 1300
rect 16810 1213 16820 1285
rect 16840 1213 16850 1285
rect 16810 1200 16850 1213
rect 16865 1285 16905 1300
rect 16865 1213 16875 1285
rect 16895 1213 16905 1285
rect 16865 1200 16905 1213
rect 16920 1285 16960 1300
rect 16920 1213 16930 1285
rect 16950 1213 16960 1285
rect 16920 1200 16960 1213
rect 16975 1285 17015 1300
rect 16975 1213 16985 1285
rect 17005 1213 17015 1285
rect 16975 1200 17015 1213
rect 17030 1285 17070 1300
rect 17030 1213 17040 1285
rect 17060 1213 17070 1285
rect 17030 1200 17070 1213
rect 17085 1285 17125 1300
rect 17085 1213 17095 1285
rect 17115 1213 17125 1285
rect 17085 1200 17125 1213
rect 17140 1285 17180 1300
rect 17140 1213 17150 1285
rect 17170 1213 17180 1285
rect 17140 1200 17180 1213
rect 17450 1285 17490 1300
rect 17450 1215 17460 1285
rect 17480 1215 17490 1285
rect 17450 1200 17490 1215
rect 17505 1285 17545 1300
rect 17505 1215 17515 1285
rect 17535 1215 17545 1285
rect 17505 1200 17545 1215
rect 17560 1285 17600 1300
rect 17560 1215 17570 1285
rect 17590 1215 17600 1285
rect 17560 1200 17600 1215
rect 17615 1285 17655 1300
rect 17615 1215 17625 1285
rect 17645 1215 17655 1285
rect 17615 1200 17655 1215
rect 17670 1285 17710 1300
rect 17670 1215 17680 1285
rect 17700 1215 17710 1285
rect 17670 1200 17710 1215
rect 17725 1285 17765 1300
rect 17725 1215 17735 1285
rect 17755 1215 17765 1285
rect 17725 1200 17765 1215
rect 17780 1285 17820 1300
rect 17780 1215 17790 1285
rect 17810 1215 17820 1285
rect 17780 1200 17820 1215
rect 17835 1285 17875 1300
rect 17835 1215 17845 1285
rect 17865 1215 17875 1285
rect 17835 1200 17875 1215
rect 17890 1285 17930 1300
rect 17890 1215 17900 1285
rect 17920 1215 17930 1285
rect 17890 1200 17930 1215
rect 17945 1285 17985 1300
rect 17945 1215 17955 1285
rect 17975 1215 17985 1285
rect 17945 1200 17985 1215
rect 18000 1285 18040 1300
rect 18000 1215 18010 1285
rect 18030 1215 18040 1285
rect 18000 1200 18040 1215
rect 18055 1285 18095 1300
rect 18055 1215 18065 1285
rect 18085 1215 18095 1285
rect 18055 1200 18095 1215
rect 18110 1285 18150 1300
rect 18110 1215 18120 1285
rect 18140 1215 18150 1285
rect 18110 1200 18150 1215
rect 18420 1285 18460 1300
rect 18420 1213 18430 1285
rect 18450 1213 18460 1285
rect 18420 1200 18460 1213
rect 18475 1285 18515 1300
rect 18475 1213 18485 1285
rect 18505 1213 18515 1285
rect 18475 1200 18515 1213
rect 18530 1285 18570 1300
rect 18530 1213 18540 1285
rect 18560 1213 18570 1285
rect 18530 1200 18570 1213
rect 18585 1285 18625 1300
rect 18585 1213 18595 1285
rect 18615 1213 18625 1285
rect 18585 1200 18625 1213
rect 18640 1285 18680 1300
rect 18640 1213 18650 1285
rect 18670 1213 18680 1285
rect 18640 1200 18680 1213
rect 18695 1285 18735 1300
rect 18695 1213 18705 1285
rect 18725 1213 18735 1285
rect 18695 1200 18735 1213
rect 18750 1285 18790 1300
rect 18750 1213 18760 1285
rect 18780 1213 18790 1285
rect 18750 1200 18790 1213
rect 16970 775 17010 790
rect 16435 685 16475 700
rect 16435 615 16445 685
rect 16465 615 16475 685
rect 16435 600 16475 615
rect 16490 685 16530 700
rect 16490 615 16500 685
rect 16520 615 16530 685
rect 16490 600 16530 615
rect 16545 685 16585 700
rect 16545 615 16555 685
rect 16575 615 16585 685
rect 16545 600 16585 615
rect 16600 685 16640 700
rect 16600 615 16610 685
rect 16630 615 16640 685
rect 16600 600 16640 615
rect 16655 685 16695 700
rect 16655 615 16665 685
rect 16685 615 16695 685
rect 16655 600 16695 615
rect 16970 505 16980 775
rect 17000 505 17010 775
rect 16970 490 17010 505
rect 17060 775 17100 790
rect 17060 505 17070 775
rect 17090 505 17100 775
rect 17060 490 17100 505
rect 17150 775 17190 790
rect 17150 505 17160 775
rect 17180 505 17190 775
rect 17150 490 17190 505
rect 17240 775 17280 790
rect 17240 505 17250 775
rect 17270 505 17280 775
rect 17240 490 17280 505
rect 17330 775 17370 790
rect 17330 505 17340 775
rect 17360 505 17370 775
rect 17330 490 17370 505
rect 17420 775 17460 790
rect 17420 505 17430 775
rect 17450 505 17460 775
rect 17420 490 17460 505
rect 17510 775 17550 790
rect 17510 505 17520 775
rect 17540 505 17550 775
rect 17510 490 17550 505
rect 17600 775 17640 790
rect 17600 505 17610 775
rect 17630 505 17640 775
rect 17600 490 17640 505
rect 17690 775 17730 790
rect 17690 505 17700 775
rect 17720 505 17730 775
rect 17690 490 17730 505
rect 17780 775 17820 790
rect 17780 505 17790 775
rect 17810 505 17820 775
rect 17780 490 17820 505
rect 17870 775 17910 790
rect 17870 505 17880 775
rect 17900 505 17910 775
rect 17870 490 17910 505
rect 17960 775 18000 790
rect 17960 505 17970 775
rect 17990 505 18000 775
rect 17960 490 18000 505
rect 18050 775 18090 790
rect 18050 505 18060 775
rect 18080 505 18090 775
rect 18050 490 18090 505
rect 18140 775 18180 790
rect 18140 505 18150 775
rect 18170 505 18180 775
rect 18140 490 18180 505
rect 18230 775 18270 790
rect 18230 505 18240 775
rect 18260 505 18270 775
rect 18230 490 18270 505
rect 18320 775 18360 790
rect 18320 505 18330 775
rect 18350 505 18360 775
rect 18320 490 18360 505
rect 18410 775 18450 790
rect 18410 505 18420 775
rect 18440 505 18450 775
rect 18410 490 18450 505
rect 18500 775 18540 790
rect 18500 505 18510 775
rect 18530 505 18540 775
rect 18500 490 18540 505
rect 18590 775 18630 790
rect 18590 505 18600 775
rect 18620 505 18630 775
rect 18900 685 18940 700
rect 18900 615 18910 685
rect 18930 615 18940 685
rect 18900 600 18940 615
rect 18955 685 18995 700
rect 18955 615 18965 685
rect 18985 615 18995 685
rect 18955 600 18995 615
rect 19010 685 19050 700
rect 19010 615 19020 685
rect 19040 615 19050 685
rect 19010 600 19050 615
rect 19065 685 19105 700
rect 19065 615 19075 685
rect 19095 615 19105 685
rect 19065 600 19105 615
rect 19120 685 19160 700
rect 19120 615 19130 685
rect 19150 615 19160 685
rect 19120 600 19160 615
rect 18590 490 18630 505
rect 16420 35 16460 50
rect 16420 -35 16430 35
rect 16450 -35 16460 35
rect 16420 -50 16460 -35
rect 16480 35 16520 50
rect 16480 -35 16490 35
rect 16510 -35 16520 35
rect 16480 -50 16520 -35
rect 16540 35 16580 50
rect 16540 -35 16550 35
rect 16570 -35 16580 35
rect 16540 -50 16580 -35
rect 16600 35 16640 50
rect 16600 -35 16610 35
rect 16630 -35 16640 35
rect 16600 -50 16640 -35
rect 16660 35 16700 50
rect 16660 -35 16670 35
rect 16690 -35 16700 35
rect 16660 -50 16700 -35
rect 16720 35 16760 50
rect 16720 -35 16730 35
rect 16750 -35 16760 35
rect 16720 -50 16760 -35
rect 16780 35 16820 50
rect 16780 -35 16790 35
rect 16810 -35 16820 35
rect 16780 -50 16820 -35
rect 16840 35 16880 50
rect 16840 -35 16850 35
rect 16870 -35 16880 35
rect 16840 -50 16880 -35
rect 16900 35 16940 50
rect 16900 -35 16910 35
rect 16930 -35 16940 35
rect 16900 -50 16940 -35
rect 16960 35 17000 50
rect 16960 -35 16970 35
rect 16990 -35 17000 35
rect 16960 -50 17000 -35
rect 17020 35 17060 50
rect 17020 -35 17030 35
rect 17050 -35 17060 35
rect 17020 -50 17060 -35
rect 17080 35 17120 50
rect 17080 -35 17090 35
rect 17110 -35 17120 35
rect 17080 -50 17120 -35
rect 17140 35 17180 50
rect 17140 -35 17150 35
rect 17170 -35 17180 35
rect 17140 -50 17180 -35
rect 17200 35 17240 50
rect 17200 -35 17210 35
rect 17230 -35 17240 35
rect 17200 -50 17240 -35
rect 17260 35 17300 50
rect 17260 -35 17270 35
rect 17290 -35 17300 35
rect 17260 -50 17300 -35
rect 17320 35 17360 50
rect 17320 -35 17330 35
rect 17350 -35 17360 35
rect 17320 -50 17360 -35
rect 17380 35 17420 50
rect 17380 -35 17390 35
rect 17410 -35 17420 35
rect 17380 -50 17420 -35
rect 17440 35 17480 50
rect 17440 -35 17450 35
rect 17470 -35 17480 35
rect 17440 -50 17480 -35
rect 17500 35 17540 50
rect 17500 -35 17510 35
rect 17530 -35 17540 35
rect 17500 -50 17540 -35
rect 17560 35 17600 50
rect 17560 -35 17570 35
rect 17590 -35 17600 35
rect 17560 -50 17600 -35
rect 17620 35 17660 50
rect 17620 -35 17630 35
rect 17650 -35 17660 35
rect 17620 -50 17660 -35
rect 17940 35 17980 50
rect 17940 -35 17950 35
rect 17970 -35 17980 35
rect 17940 -50 17980 -35
rect 18000 35 18040 50
rect 18000 -35 18010 35
rect 18030 -35 18040 35
rect 18000 -50 18040 -35
rect 18060 35 18100 50
rect 18060 -35 18070 35
rect 18090 -35 18100 35
rect 18060 -50 18100 -35
rect 18120 35 18160 50
rect 18120 -35 18130 35
rect 18150 -35 18160 35
rect 18120 -50 18160 -35
rect 18180 35 18220 50
rect 18180 -35 18190 35
rect 18210 -35 18220 35
rect 18180 -50 18220 -35
rect 18240 35 18280 50
rect 18240 -35 18250 35
rect 18270 -35 18280 35
rect 18240 -50 18280 -35
rect 18300 35 18340 50
rect 18300 -35 18310 35
rect 18330 -35 18340 35
rect 18300 -50 18340 -35
rect 18360 35 18400 50
rect 18360 -35 18370 35
rect 18390 -35 18400 35
rect 18360 -50 18400 -35
rect 18420 35 18460 50
rect 18420 -35 18430 35
rect 18450 -35 18460 35
rect 18420 -50 18460 -35
rect 18480 35 18520 50
rect 18480 -35 18490 35
rect 18510 -35 18520 35
rect 18480 -50 18520 -35
rect 18540 35 18580 50
rect 18540 -35 18550 35
rect 18570 -35 18580 35
rect 18540 -50 18580 -35
rect 18600 35 18640 50
rect 18600 -35 18610 35
rect 18630 -35 18640 35
rect 18600 -50 18640 -35
rect 18660 35 18700 50
rect 18660 -35 18670 35
rect 18690 -35 18700 35
rect 18660 -50 18700 -35
rect 18720 35 18760 50
rect 18720 -35 18730 35
rect 18750 -35 18760 35
rect 18720 -50 18760 -35
rect 18780 35 18820 50
rect 18780 -35 18790 35
rect 18810 -35 18820 35
rect 18780 -50 18820 -35
rect 18840 35 18880 50
rect 18840 -35 18850 35
rect 18870 -35 18880 35
rect 18840 -50 18880 -35
rect 18900 35 18940 50
rect 18900 -35 18910 35
rect 18930 -35 18940 35
rect 18900 -50 18940 -35
rect 18960 35 19000 50
rect 18960 -35 18970 35
rect 18990 -35 19000 35
rect 18960 -50 19000 -35
rect 19020 35 19060 50
rect 19020 -35 19030 35
rect 19050 -35 19060 35
rect 19020 -50 19060 -35
rect 19080 35 19120 50
rect 19080 -35 19090 35
rect 19110 -35 19120 35
rect 19080 -50 19120 -35
rect 19140 35 19180 50
rect 19140 -35 19150 35
rect 19170 -35 19180 35
rect 19140 -50 19180 -35
<< ndiffc >>
rect 16860 -485 16880 -465
rect 16920 -485 16940 -465
rect 16980 -485 17000 -465
rect 17040 -485 17060 -465
rect 17100 -485 17120 -465
rect 17160 -485 17180 -465
rect 17220 -485 17240 -465
rect 17280 -485 17300 -465
rect 17340 -485 17360 -465
rect 17400 -485 17420 -465
rect 17460 -485 17480 -465
rect 18120 -485 18140 -465
rect 18180 -485 18200 -465
rect 18240 -485 18260 -465
rect 18300 -485 18320 -465
rect 18360 -485 18380 -465
rect 18420 -485 18440 -465
rect 18480 -485 18500 -465
rect 18540 -485 18560 -465
rect 18600 -485 18620 -465
rect 18660 -485 18680 -465
rect 18720 -485 18740 -465
rect 16540 -960 16560 -740
rect 17080 -960 17100 -740
rect 17160 -960 17180 -740
rect 17700 -960 17720 -740
rect 17880 -960 17900 -740
rect 18420 -960 18440 -740
rect 18500 -960 18520 -740
rect 19040 -960 19060 -740
rect 16750 -1230 16770 -1160
rect 17790 -1230 17810 -1160
rect 18830 -1230 18850 -1160
rect 16925 -1570 16945 -1500
rect 16980 -1570 17000 -1500
rect 17035 -1570 17055 -1500
rect 17090 -1570 17110 -1500
rect 17145 -1570 17165 -1500
rect 17200 -1570 17220 -1500
rect 17255 -1570 17275 -1500
rect 17310 -1570 17330 -1500
rect 17365 -1570 17385 -1500
rect 17515 -1570 17535 -1500
rect 17570 -1570 17590 -1500
rect 17625 -1570 17645 -1500
rect 17680 -1570 17700 -1500
rect 17735 -1570 17755 -1500
rect 17790 -1570 17810 -1500
rect 17845 -1570 17865 -1500
rect 17900 -1570 17920 -1500
rect 17955 -1570 17975 -1500
rect 18010 -1570 18030 -1500
rect 18065 -1570 18085 -1500
rect 18225 -1570 18245 -1500
rect 18280 -1570 18300 -1500
rect 18335 -1570 18355 -1500
rect 18390 -1570 18410 -1500
rect 18445 -1570 18465 -1500
rect 18500 -1570 18520 -1500
rect 18555 -1570 18575 -1500
rect 18610 -1570 18630 -1500
rect 18665 -1570 18685 -1500
<< pdiffc >>
rect 16820 1213 16840 1285
rect 16875 1213 16895 1285
rect 16930 1213 16950 1285
rect 16985 1213 17005 1285
rect 17040 1213 17060 1285
rect 17095 1213 17115 1285
rect 17150 1213 17170 1285
rect 17460 1215 17480 1285
rect 17515 1215 17535 1285
rect 17570 1215 17590 1285
rect 17625 1215 17645 1285
rect 17680 1215 17700 1285
rect 17735 1215 17755 1285
rect 17790 1215 17810 1285
rect 17845 1215 17865 1285
rect 17900 1215 17920 1285
rect 17955 1215 17975 1285
rect 18010 1215 18030 1285
rect 18065 1215 18085 1285
rect 18120 1215 18140 1285
rect 18430 1213 18450 1285
rect 18485 1213 18505 1285
rect 18540 1213 18560 1285
rect 18595 1213 18615 1285
rect 18650 1213 18670 1285
rect 18705 1213 18725 1285
rect 18760 1213 18780 1285
rect 16445 615 16465 685
rect 16500 615 16520 685
rect 16555 615 16575 685
rect 16610 615 16630 685
rect 16665 615 16685 685
rect 16980 505 17000 775
rect 17070 505 17090 775
rect 17160 505 17180 775
rect 17250 505 17270 775
rect 17340 505 17360 775
rect 17430 505 17450 775
rect 17520 505 17540 775
rect 17610 505 17630 775
rect 17700 505 17720 775
rect 17790 505 17810 775
rect 17880 505 17900 775
rect 17970 505 17990 775
rect 18060 505 18080 775
rect 18150 505 18170 775
rect 18240 505 18260 775
rect 18330 505 18350 775
rect 18420 505 18440 775
rect 18510 505 18530 775
rect 18600 505 18620 775
rect 18910 615 18930 685
rect 18965 615 18985 685
rect 19020 615 19040 685
rect 19075 615 19095 685
rect 19130 615 19150 685
rect 16430 -35 16450 35
rect 16490 -35 16510 35
rect 16550 -35 16570 35
rect 16610 -35 16630 35
rect 16670 -35 16690 35
rect 16730 -35 16750 35
rect 16790 -35 16810 35
rect 16850 -35 16870 35
rect 16910 -35 16930 35
rect 16970 -35 16990 35
rect 17030 -35 17050 35
rect 17090 -35 17110 35
rect 17150 -35 17170 35
rect 17210 -35 17230 35
rect 17270 -35 17290 35
rect 17330 -35 17350 35
rect 17390 -35 17410 35
rect 17450 -35 17470 35
rect 17510 -35 17530 35
rect 17570 -35 17590 35
rect 17630 -35 17650 35
rect 17950 -35 17970 35
rect 18010 -35 18030 35
rect 18070 -35 18090 35
rect 18130 -35 18150 35
rect 18190 -35 18210 35
rect 18250 -35 18270 35
rect 18310 -35 18330 35
rect 18370 -35 18390 35
rect 18430 -35 18450 35
rect 18490 -35 18510 35
rect 18550 -35 18570 35
rect 18610 -35 18630 35
rect 18670 -35 18690 35
rect 18730 -35 18750 35
rect 18790 -35 18810 35
rect 18850 -35 18870 35
rect 18910 -35 18930 35
rect 18970 -35 18990 35
rect 19030 -35 19050 35
rect 19090 -35 19110 35
rect 19150 -35 19170 35
<< psubdiff >>
rect 17560 -465 17600 -450
rect 17560 -485 17570 -465
rect 17590 -485 17600 -465
rect 17560 -500 17600 -485
rect 18000 -465 18040 -450
rect 18000 -485 18010 -465
rect 18030 -485 18040 -465
rect 18000 -500 18040 -485
rect 17110 -740 17150 -725
rect 17110 -960 17120 -740
rect 17140 -960 17150 -740
rect 17110 -970 17150 -960
rect 18450 -740 18490 -725
rect 18450 -960 18460 -740
rect 18480 -960 18490 -740
rect 18450 -975 18490 -960
rect 18860 -1160 18900 -1145
rect 18860 -1230 18870 -1160
rect 18890 -1230 18900 -1160
rect 18860 -1245 18900 -1230
rect 16875 -1500 16915 -1485
rect 16875 -1570 16885 -1500
rect 16905 -1570 16915 -1500
rect 16875 -1585 16915 -1570
rect 17395 -1500 17435 -1485
rect 17395 -1570 17405 -1500
rect 17425 -1570 17435 -1500
rect 17395 -1585 17435 -1570
rect 17465 -1500 17505 -1485
rect 17465 -1570 17475 -1500
rect 17495 -1570 17505 -1500
rect 17465 -1585 17505 -1570
rect 18095 -1500 18135 -1485
rect 18095 -1570 18105 -1500
rect 18125 -1570 18135 -1500
rect 18095 -1585 18135 -1570
rect 18175 -1500 18215 -1485
rect 18175 -1570 18185 -1500
rect 18205 -1570 18215 -1500
rect 18175 -1585 18215 -1570
rect 18695 -1500 18735 -1485
rect 18695 -1570 18705 -1500
rect 18725 -1570 18735 -1500
rect 18695 -1585 18735 -1570
rect 17775 -4170 17825 -4155
rect 17775 -4190 17790 -4170
rect 17810 -4190 17825 -4170
rect 17775 -4220 17825 -4190
rect 17775 -4240 17790 -4220
rect 17810 -4240 17825 -4220
rect 17775 -4270 17825 -4240
rect 17775 -4290 17790 -4270
rect 17810 -4290 17825 -4270
rect 17775 -4305 17825 -4290
<< nsubdiff >>
rect 16770 1287 16810 1300
rect 16770 1215 16780 1287
rect 16800 1215 16810 1287
rect 16770 1200 16810 1215
rect 17180 1287 17220 1300
rect 17180 1215 17190 1287
rect 17210 1215 17220 1287
rect 17180 1200 17220 1215
rect 17410 1287 17450 1300
rect 17410 1215 17420 1287
rect 17440 1215 17450 1287
rect 17410 1200 17450 1215
rect 18150 1287 18190 1300
rect 18150 1215 18160 1287
rect 18180 1215 18190 1287
rect 18150 1200 18190 1215
rect 18380 1287 18420 1300
rect 18380 1215 18390 1287
rect 18410 1215 18420 1287
rect 18380 1200 18420 1215
rect 18790 1287 18830 1300
rect 18790 1215 18800 1287
rect 18820 1215 18830 1287
rect 18790 1200 18830 1215
rect 16930 775 16970 790
rect 16395 685 16435 700
rect 16395 615 16405 685
rect 16425 615 16435 685
rect 16395 600 16435 615
rect 16695 685 16735 700
rect 16695 615 16705 685
rect 16725 615 16735 685
rect 16695 600 16735 615
rect 16930 505 16940 775
rect 16960 505 16970 775
rect 16930 490 16970 505
rect 18630 775 18670 790
rect 18630 505 18640 775
rect 18660 505 18670 775
rect 18860 685 18900 700
rect 18860 615 18870 685
rect 18890 615 18900 685
rect 18860 600 18900 615
rect 19160 685 19200 700
rect 19160 615 19170 685
rect 19190 615 19200 685
rect 19160 600 19200 615
rect 18630 490 18670 505
rect 16380 35 16420 50
rect 16380 -35 16390 35
rect 16410 -35 16420 35
rect 16380 -50 16420 -35
rect 17660 35 17700 50
rect 17660 -35 17670 35
rect 17690 -35 17700 35
rect 17660 -50 17700 -35
rect 17900 35 17940 50
rect 17900 -35 17910 35
rect 17930 -35 17940 35
rect 17900 -50 17940 -35
rect 19180 35 19220 50
rect 19180 -35 19190 35
rect 19210 -35 19220 35
rect 19180 -50 19220 -35
<< psubdiffcont >>
rect 17570 -485 17590 -465
rect 18010 -485 18030 -465
rect 17120 -960 17140 -740
rect 18460 -960 18480 -740
rect 18870 -1230 18890 -1160
rect 16885 -1570 16905 -1500
rect 17405 -1570 17425 -1500
rect 17475 -1570 17495 -1500
rect 18105 -1570 18125 -1500
rect 18185 -1570 18205 -1500
rect 18705 -1570 18725 -1500
rect 17790 -4190 17810 -4170
rect 17790 -4240 17810 -4220
rect 17790 -4290 17810 -4270
<< nsubdiffcont >>
rect 16780 1215 16800 1287
rect 17190 1215 17210 1287
rect 17420 1215 17440 1287
rect 18160 1215 18180 1287
rect 18390 1215 18410 1287
rect 18800 1215 18820 1287
rect 16405 615 16425 685
rect 16705 615 16725 685
rect 16940 505 16960 775
rect 18640 505 18660 775
rect 18870 615 18890 685
rect 19170 615 19190 685
rect 16390 -35 16410 35
rect 17670 -35 17690 35
rect 17910 -35 17930 35
rect 19190 -35 19210 35
<< poly >>
rect 16810 1345 16850 1355
rect 16810 1325 16820 1345
rect 16840 1330 16850 1345
rect 17140 1345 17180 1355
rect 16840 1325 16865 1330
rect 17140 1325 17150 1345
rect 17170 1325 17180 1345
rect 16810 1315 16865 1325
rect 16850 1300 16865 1315
rect 16905 1300 16920 1315
rect 16960 1300 16975 1315
rect 17015 1300 17030 1315
rect 17070 1300 17085 1315
rect 17125 1310 17180 1325
rect 17450 1345 17490 1355
rect 17450 1325 17460 1345
rect 17480 1330 17490 1345
rect 18110 1345 18150 1355
rect 18110 1330 18120 1345
rect 17480 1325 17505 1330
rect 17450 1315 17505 1325
rect 18095 1325 18120 1330
rect 18140 1325 18150 1345
rect 18095 1315 18150 1325
rect 18420 1345 18460 1355
rect 18420 1325 18430 1345
rect 18450 1325 18460 1345
rect 18750 1345 18790 1355
rect 18750 1330 18760 1345
rect 18735 1325 18760 1330
rect 18780 1325 18790 1345
rect 17125 1300 17140 1310
rect 17490 1300 17505 1315
rect 17545 1300 17560 1315
rect 17600 1300 17615 1315
rect 17655 1300 17670 1315
rect 17710 1300 17725 1315
rect 17765 1300 17780 1315
rect 17820 1300 17835 1315
rect 17875 1300 17890 1315
rect 17930 1300 17945 1315
rect 17985 1300 18000 1315
rect 18040 1300 18055 1315
rect 18095 1300 18110 1315
rect 18420 1310 18475 1325
rect 18735 1315 18790 1325
rect 18460 1300 18475 1310
rect 18515 1300 18530 1315
rect 18570 1300 18585 1315
rect 18625 1300 18640 1315
rect 18680 1300 18695 1315
rect 18735 1300 18750 1315
rect 16850 1185 16865 1200
rect 16905 1190 16920 1200
rect 16960 1190 16975 1200
rect 17015 1190 17030 1200
rect 17070 1190 17085 1200
rect 16905 1175 17085 1190
rect 17125 1185 17140 1200
rect 17490 1185 17505 1200
rect 17545 1190 17560 1200
rect 17600 1190 17615 1200
rect 17655 1190 17670 1200
rect 17710 1190 17725 1200
rect 17765 1190 17780 1200
rect 17820 1190 17835 1200
rect 17875 1190 17890 1200
rect 17930 1190 17945 1200
rect 17985 1190 18000 1200
rect 18040 1190 18055 1200
rect 17545 1175 18055 1190
rect 18095 1185 18110 1200
rect 18460 1185 18475 1200
rect 18515 1190 18530 1200
rect 18570 1190 18585 1200
rect 18625 1190 18640 1200
rect 18680 1190 18695 1200
rect 18515 1175 18695 1190
rect 18735 1185 18750 1200
rect 17070 1100 17085 1175
rect 17820 1100 17835 1175
rect 18515 1100 18530 1175
rect 17070 1090 17100 1100
rect 17070 1070 17075 1090
rect 17095 1070 17100 1090
rect 17070 1060 17100 1070
rect 17805 1090 17835 1100
rect 17805 1070 17810 1090
rect 17830 1070 17835 1090
rect 17805 1060 17835 1070
rect 18500 1090 18530 1100
rect 18500 1070 18505 1090
rect 18525 1070 18530 1090
rect 18500 1060 18530 1070
rect 16970 835 17010 845
rect 16970 815 16980 835
rect 17000 820 17010 835
rect 18590 835 18630 845
rect 18590 820 18600 835
rect 17000 815 17060 820
rect 16970 805 17060 815
rect 18540 815 18600 820
rect 18620 815 18630 835
rect 18540 805 18630 815
rect 17010 790 17060 805
rect 17100 790 17150 805
rect 17190 790 17240 805
rect 17280 790 17330 805
rect 17370 790 17420 805
rect 17460 790 17510 805
rect 17550 790 17600 805
rect 17640 790 17690 805
rect 17730 790 17780 805
rect 17820 790 17870 805
rect 17910 790 17960 805
rect 18000 790 18050 805
rect 18090 790 18140 805
rect 18180 790 18230 805
rect 18270 790 18320 805
rect 18360 790 18410 805
rect 18450 790 18500 805
rect 18540 790 18590 805
rect 16440 775 16470 785
rect 16440 755 16445 775
rect 16465 760 16470 775
rect 16660 775 16690 785
rect 16660 760 16665 775
rect 16465 755 16490 760
rect 16440 745 16490 755
rect 16475 700 16490 745
rect 16640 755 16665 760
rect 16685 755 16690 775
rect 16640 745 16690 755
rect 16530 700 16545 715
rect 16585 700 16600 715
rect 16640 700 16655 745
rect 16475 585 16490 600
rect 16530 590 16545 600
rect 16585 590 16600 600
rect 16530 575 16600 590
rect 16640 585 16655 600
rect 16550 565 16580 575
rect 16550 545 16555 565
rect 16575 545 16580 565
rect 16550 535 16580 545
rect 18900 775 18940 785
rect 18900 755 18910 775
rect 18930 760 18940 775
rect 19120 775 19160 785
rect 19120 760 19130 775
rect 18930 755 18955 760
rect 18900 745 18955 755
rect 18940 700 18955 745
rect 19105 755 19130 760
rect 19150 755 19160 775
rect 19105 745 19160 755
rect 18995 700 19010 715
rect 19050 700 19065 715
rect 19105 700 19120 745
rect 18940 585 18955 600
rect 18995 590 19010 600
rect 19050 590 19065 600
rect 18995 575 19065 590
rect 19105 585 19120 600
rect 19020 545 19040 575
rect 19015 535 19045 545
rect 19015 515 19020 535
rect 19040 515 19045 535
rect 19015 505 19045 515
rect 17010 475 17060 490
rect 17100 480 17150 490
rect 17190 480 17240 490
rect 17280 480 17330 490
rect 17370 480 17420 490
rect 17460 480 17510 490
rect 17550 480 17600 490
rect 17640 480 17690 490
rect 17730 480 17780 490
rect 17820 480 17870 490
rect 17910 480 17960 490
rect 18000 480 18050 490
rect 18090 480 18140 490
rect 18180 480 18230 490
rect 18270 480 18320 490
rect 18360 480 18410 490
rect 18450 480 18500 490
rect 17100 465 18500 480
rect 18540 475 18590 490
rect 17695 455 17725 465
rect 17695 435 17700 455
rect 17720 435 17725 455
rect 17695 425 17725 435
rect 16425 100 16455 110
rect 16425 80 16430 100
rect 16450 85 16455 100
rect 17625 100 17655 110
rect 17625 85 17630 100
rect 16450 80 16480 85
rect 16425 70 16480 80
rect 16460 50 16480 70
rect 17600 80 17630 85
rect 17650 80 17655 100
rect 17600 70 17655 80
rect 17945 100 17975 110
rect 17945 80 17950 100
rect 17970 85 17975 100
rect 19145 100 19175 110
rect 19145 85 19150 100
rect 17970 80 18000 85
rect 17945 70 18000 80
rect 16520 50 16540 65
rect 16580 50 16600 65
rect 16640 50 16660 65
rect 16700 50 16720 65
rect 16760 50 16780 65
rect 16820 50 16840 65
rect 16880 50 16900 65
rect 16940 50 16960 65
rect 17000 50 17020 65
rect 17060 50 17080 65
rect 17120 50 17140 65
rect 17180 50 17200 65
rect 17240 50 17260 65
rect 17300 50 17320 65
rect 17360 50 17380 65
rect 17420 50 17440 65
rect 17480 50 17500 65
rect 17540 50 17560 65
rect 17600 50 17620 70
rect 17980 50 18000 70
rect 19120 80 19150 85
rect 19170 80 19175 100
rect 19120 70 19175 80
rect 18040 50 18060 65
rect 18100 50 18120 65
rect 18160 50 18180 65
rect 18220 50 18240 65
rect 18280 50 18300 65
rect 18340 50 18360 65
rect 18400 50 18420 65
rect 18460 50 18480 65
rect 18520 50 18540 65
rect 18580 50 18600 65
rect 18640 50 18660 65
rect 18700 50 18720 65
rect 18760 50 18780 65
rect 18820 50 18840 65
rect 18880 50 18900 65
rect 18940 50 18960 65
rect 19000 50 19020 65
rect 19060 50 19080 65
rect 19120 50 19140 70
rect 16460 -65 16480 -50
rect 16520 -215 16540 -50
rect 16580 -60 16600 -50
rect 16640 -60 16660 -50
rect 16700 -60 16720 -50
rect 16760 -60 16780 -50
rect 16580 -75 16780 -60
rect 16820 -60 16840 -50
rect 16880 -60 16900 -50
rect 16820 -75 16900 -60
rect 16940 -60 16960 -50
rect 17000 -60 17020 -50
rect 17060 -60 17080 -50
rect 17120 -60 17140 -50
rect 16940 -75 17140 -60
rect 17180 -60 17200 -50
rect 17240 -60 17260 -50
rect 17180 -75 17260 -60
rect 17300 -60 17320 -50
rect 17360 -60 17380 -50
rect 17420 -60 17440 -50
rect 17480 -60 17500 -50
rect 17300 -75 17500 -60
rect 16600 -95 16610 -75
rect 16630 -95 16640 -75
rect 16600 -105 16640 -95
rect 16880 -215 16900 -75
rect 16960 -95 16970 -75
rect 16990 -95 17000 -75
rect 16960 -105 17000 -95
rect 17240 -215 17260 -75
rect 17320 -95 17330 -75
rect 17350 -95 17360 -75
rect 17320 -105 17360 -95
rect 17540 -215 17560 -50
rect 17600 -65 17620 -50
rect 17980 -65 18000 -50
rect 16520 -225 16570 -215
rect 16520 -245 16545 -225
rect 16565 -245 16570 -225
rect 16880 -225 16930 -215
rect 16880 -245 16905 -225
rect 16925 -245 16930 -225
rect 17240 -225 17290 -215
rect 17240 -245 17265 -225
rect 17285 -245 17290 -225
rect 16540 -255 16570 -245
rect 16900 -255 16930 -245
rect 17260 -255 17290 -245
rect 17510 -225 17560 -215
rect 17510 -245 17515 -225
rect 17535 -245 17560 -225
rect 18040 -215 18060 -50
rect 18100 -60 18120 -50
rect 18160 -60 18180 -50
rect 18220 -60 18240 -50
rect 18280 -60 18300 -50
rect 18100 -75 18300 -60
rect 18340 -60 18360 -50
rect 18400 -60 18420 -50
rect 18340 -75 18420 -60
rect 18460 -60 18480 -50
rect 18520 -60 18540 -50
rect 18580 -60 18600 -50
rect 18640 -60 18660 -50
rect 18460 -75 18660 -60
rect 18700 -60 18720 -50
rect 18760 -60 18780 -50
rect 18700 -75 18780 -60
rect 18820 -60 18840 -50
rect 18880 -60 18900 -50
rect 18940 -60 18960 -50
rect 19000 -60 19020 -50
rect 18820 -75 19020 -60
rect 18240 -95 18250 -75
rect 18270 -95 18280 -75
rect 18240 -105 18280 -95
rect 18340 -215 18360 -75
rect 18600 -95 18610 -75
rect 18630 -95 18640 -75
rect 18600 -105 18640 -95
rect 18700 -215 18720 -75
rect 18960 -95 18970 -75
rect 18990 -95 19000 -75
rect 18960 -105 19000 -95
rect 19060 -215 19080 -50
rect 19120 -65 19140 -50
rect 18040 -225 18090 -215
rect 18040 -245 18065 -225
rect 18085 -245 18090 -225
rect 17510 -255 17540 -245
rect 18060 -255 18090 -245
rect 18310 -225 18360 -215
rect 18310 -245 18315 -225
rect 18335 -245 18360 -225
rect 18670 -225 18720 -215
rect 18670 -245 18675 -225
rect 18695 -245 18720 -225
rect 19030 -225 19080 -215
rect 19030 -245 19035 -225
rect 19055 -245 19080 -225
rect 18310 -255 18340 -245
rect 18670 -255 18700 -245
rect 19030 -255 19060 -245
rect 16800 -395 16830 -385
rect 18770 -395 18800 -385
rect 16800 -415 16805 -395
rect 16825 -410 17450 -395
rect 16825 -415 16830 -410
rect 16800 -425 16830 -415
rect 16890 -450 16910 -435
rect 16950 -450 16970 -410
rect 17010 -450 17030 -410
rect 17070 -450 17090 -435
rect 17130 -450 17150 -435
rect 17190 -450 17210 -410
rect 17250 -450 17270 -410
rect 17310 -450 17330 -435
rect 17370 -450 17390 -435
rect 17430 -450 17450 -410
rect 18150 -410 18775 -395
rect 18150 -450 18170 -410
rect 18210 -450 18230 -435
rect 18270 -450 18290 -435
rect 18330 -450 18350 -410
rect 18390 -450 18410 -410
rect 18450 -450 18470 -435
rect 18510 -450 18530 -435
rect 18570 -450 18590 -410
rect 18630 -450 18650 -410
rect 18770 -415 18775 -410
rect 18795 -415 18800 -395
rect 18770 -425 18800 -415
rect 18690 -450 18710 -435
rect 16800 -535 16830 -525
rect 16800 -555 16805 -535
rect 16825 -540 16830 -535
rect 16890 -540 16910 -500
rect 16950 -515 16970 -500
rect 17010 -515 17030 -500
rect 17070 -540 17090 -500
rect 17130 -540 17150 -500
rect 17190 -515 17210 -500
rect 17250 -515 17270 -500
rect 17310 -540 17330 -500
rect 17370 -540 17390 -500
rect 17430 -515 17450 -500
rect 18150 -515 18170 -500
rect 16825 -555 17390 -540
rect 18210 -540 18230 -500
rect 18270 -540 18290 -500
rect 18330 -515 18350 -500
rect 18390 -515 18410 -500
rect 18450 -540 18470 -500
rect 18510 -540 18530 -500
rect 18570 -515 18590 -500
rect 18630 -515 18650 -500
rect 18690 -540 18710 -500
rect 18770 -535 18800 -525
rect 18770 -540 18775 -535
rect 18210 -555 18775 -540
rect 18795 -555 18800 -535
rect 16800 -565 16830 -555
rect 18770 -565 18800 -555
rect 16800 -685 16840 -675
rect 16800 -705 16810 -685
rect 16830 -705 16840 -685
rect 16800 -710 16840 -705
rect 17420 -685 17460 -675
rect 17420 -705 17430 -685
rect 17450 -705 17460 -685
rect 17420 -710 17460 -705
rect 18140 -685 18180 -675
rect 18140 -705 18150 -685
rect 18170 -705 18180 -685
rect 18140 -710 18180 -705
rect 18760 -685 18800 -675
rect 18760 -705 18770 -685
rect 18790 -705 18800 -685
rect 18760 -710 18800 -705
rect 16570 -725 17070 -710
rect 17190 -725 17690 -710
rect 17910 -725 18410 -710
rect 18530 -725 19030 -710
rect 16570 -990 17070 -975
rect 17190 -990 17690 -975
rect 17910 -990 18410 -975
rect 18530 -990 19030 -975
rect 17260 -1100 17300 -1090
rect 17260 -1120 17270 -1100
rect 17290 -1120 17300 -1100
rect 17260 -1130 17300 -1120
rect 18300 -1100 18340 -1090
rect 18300 -1120 18310 -1100
rect 18330 -1120 18340 -1100
rect 18300 -1130 18340 -1120
rect 16780 -1145 17780 -1130
rect 17820 -1145 18820 -1130
rect 16780 -1260 17780 -1245
rect 17820 -1260 18820 -1245
rect 17285 -1340 17315 -1330
rect 17285 -1360 17290 -1340
rect 17310 -1360 17315 -1340
rect 17285 -1370 17315 -1360
rect 17785 -1340 17815 -1330
rect 17785 -1360 17790 -1340
rect 17810 -1360 17815 -1340
rect 17785 -1370 17815 -1360
rect 18295 -1340 18325 -1330
rect 18295 -1360 18300 -1340
rect 18320 -1360 18325 -1340
rect 18295 -1370 18325 -1360
rect 16915 -1440 16955 -1430
rect 16915 -1460 16925 -1440
rect 16945 -1455 16955 -1440
rect 16945 -1460 16970 -1455
rect 17285 -1460 17300 -1370
rect 17355 -1440 17395 -1430
rect 17355 -1455 17365 -1440
rect 16915 -1470 16970 -1460
rect 16955 -1485 16970 -1470
rect 17010 -1475 17300 -1460
rect 17010 -1485 17025 -1475
rect 17065 -1485 17080 -1475
rect 17120 -1485 17135 -1475
rect 17175 -1485 17190 -1475
rect 17230 -1485 17245 -1475
rect 17285 -1485 17300 -1475
rect 17340 -1460 17365 -1455
rect 17385 -1460 17395 -1440
rect 17340 -1470 17395 -1460
rect 17505 -1440 17545 -1430
rect 17505 -1460 17515 -1440
rect 17535 -1455 17545 -1440
rect 17790 -1455 17810 -1370
rect 18055 -1440 18095 -1430
rect 18055 -1455 18065 -1440
rect 17535 -1460 17560 -1455
rect 17505 -1470 17560 -1460
rect 17340 -1485 17355 -1470
rect 17545 -1485 17560 -1470
rect 17600 -1470 18000 -1455
rect 17600 -1485 17615 -1470
rect 17655 -1485 17670 -1470
rect 17710 -1485 17725 -1470
rect 17765 -1485 17780 -1470
rect 17820 -1485 17835 -1470
rect 17875 -1485 17890 -1470
rect 17930 -1485 17945 -1470
rect 17985 -1485 18000 -1470
rect 18040 -1460 18065 -1455
rect 18085 -1460 18095 -1440
rect 18040 -1470 18095 -1460
rect 18215 -1440 18255 -1430
rect 18215 -1460 18225 -1440
rect 18245 -1455 18255 -1440
rect 18245 -1460 18270 -1455
rect 18215 -1470 18270 -1460
rect 18040 -1485 18055 -1470
rect 18255 -1485 18270 -1470
rect 18310 -1460 18325 -1370
rect 18655 -1440 18695 -1430
rect 18655 -1455 18665 -1440
rect 18640 -1460 18665 -1455
rect 18685 -1460 18695 -1440
rect 18310 -1475 18600 -1460
rect 18310 -1485 18325 -1475
rect 18365 -1485 18380 -1475
rect 18420 -1485 18435 -1475
rect 18475 -1485 18490 -1475
rect 18530 -1485 18545 -1475
rect 18585 -1485 18600 -1475
rect 18640 -1470 18695 -1460
rect 18640 -1485 18655 -1470
rect 16955 -1600 16970 -1585
rect 17010 -1600 17025 -1585
rect 17065 -1600 17080 -1585
rect 17120 -1600 17135 -1585
rect 17175 -1600 17190 -1585
rect 17230 -1600 17245 -1585
rect 17285 -1600 17300 -1585
rect 17340 -1600 17355 -1585
rect 17545 -1600 17560 -1585
rect 17600 -1640 17615 -1585
rect 17655 -1600 17670 -1585
rect 17710 -1600 17725 -1585
rect 17765 -1600 17780 -1585
rect 17820 -1600 17835 -1585
rect 17875 -1600 17890 -1585
rect 17930 -1600 17945 -1585
rect 17985 -1600 18000 -1585
rect 18040 -1600 18055 -1585
rect 18255 -1600 18270 -1585
rect 18310 -1600 18325 -1585
rect 18365 -1600 18380 -1585
rect 18420 -1600 18435 -1585
rect 18475 -1600 18490 -1585
rect 18530 -1600 18545 -1585
rect 18585 -1600 18600 -1585
rect 18640 -1600 18655 -1585
rect 17585 -1650 17615 -1640
rect 17585 -1670 17590 -1650
rect 17610 -1670 17615 -1650
rect 17585 -1680 17615 -1670
<< polycont >>
rect 16820 1325 16840 1345
rect 17150 1325 17170 1345
rect 17460 1325 17480 1345
rect 18120 1325 18140 1345
rect 18430 1325 18450 1345
rect 18760 1325 18780 1345
rect 17075 1070 17095 1090
rect 17810 1070 17830 1090
rect 18505 1070 18525 1090
rect 16980 815 17000 835
rect 18600 815 18620 835
rect 16445 755 16465 775
rect 16665 755 16685 775
rect 16555 545 16575 565
rect 18910 755 18930 775
rect 19130 755 19150 775
rect 19020 515 19040 535
rect 17700 435 17720 455
rect 16430 80 16450 100
rect 17630 80 17650 100
rect 17950 80 17970 100
rect 19150 80 19170 100
rect 16610 -95 16630 -75
rect 16970 -95 16990 -75
rect 17330 -95 17350 -75
rect 16545 -245 16565 -225
rect 16905 -245 16925 -225
rect 17265 -245 17285 -225
rect 17515 -245 17535 -225
rect 18250 -95 18270 -75
rect 18610 -95 18630 -75
rect 18970 -95 18990 -75
rect 18065 -245 18085 -225
rect 18315 -245 18335 -225
rect 18675 -245 18695 -225
rect 19035 -245 19055 -225
rect 16805 -415 16825 -395
rect 18775 -415 18795 -395
rect 16805 -555 16825 -535
rect 18775 -555 18795 -535
rect 16810 -705 16830 -685
rect 17430 -705 17450 -685
rect 18150 -705 18170 -685
rect 18770 -705 18790 -685
rect 17270 -1120 17290 -1100
rect 18310 -1120 18330 -1100
rect 17290 -1360 17310 -1340
rect 17790 -1360 17810 -1340
rect 18300 -1360 18320 -1340
rect 16925 -1460 16945 -1440
rect 17365 -1460 17385 -1440
rect 17515 -1460 17535 -1440
rect 18065 -1460 18085 -1440
rect 18225 -1460 18245 -1440
rect 18665 -1460 18685 -1440
rect 17590 -1670 17610 -1650
<< xpolycontact >>
rect 17470 -1980 17690 -1945
rect 17904 -1980 18124 -1945
rect 15950 -3376 15985 -3156
rect 15950 -3784 15985 -3565
rect 16160 -3285 16195 -3065
rect 16160 -3889 16195 -3669
rect 16220 -3285 16255 -3065
rect 16220 -3889 16255 -3669
rect 16280 -3285 16315 -3065
rect 16280 -3889 16315 -3669
rect 16485 -3160 16520 -2940
rect 16485 -3964 16520 -3744
rect 16545 -3160 16580 -2940
rect 16545 -3964 16580 -3744
rect 16605 -3160 16640 -2940
rect 16605 -3964 16640 -3744
rect 18960 -3160 18995 -2940
rect 18960 -3964 18995 -3744
rect 19020 -3160 19055 -2940
rect 19020 -3964 19055 -3744
rect 19080 -3160 19115 -2940
rect 19080 -3964 19115 -3744
rect 19285 -3252 19320 -3032
rect 19285 -3889 19320 -3669
rect 19345 -3252 19380 -3032
rect 19345 -3889 19380 -3669
rect 19405 -3252 19440 -3032
rect 19405 -3889 19440 -3669
rect 19610 -3376 19645 -3156
rect 19610 -3784 19645 -3565
<< ppolyres >>
rect 15950 -3565 15985 -3376
rect 19610 -3565 19645 -3376
<< xpolyres >>
rect 17690 -1980 17904 -1945
rect 16160 -3669 16195 -3285
rect 16220 -3669 16255 -3285
rect 16280 -3669 16315 -3285
rect 16485 -3744 16520 -3160
rect 16545 -3744 16580 -3160
rect 16605 -3744 16640 -3160
rect 18960 -3744 18995 -3160
rect 19020 -3744 19055 -3160
rect 19080 -3744 19115 -3160
rect 19285 -3669 19320 -3252
rect 19345 -3669 19380 -3252
rect 19405 -3669 19440 -3252
<< locali >>
rect 16810 1345 16850 1355
rect 16810 1325 16820 1345
rect 16840 1325 16850 1345
rect 16810 1315 16850 1325
rect 17140 1345 17180 1355
rect 17140 1325 17150 1345
rect 17170 1325 17180 1345
rect 17140 1315 17180 1325
rect 17450 1345 17490 1355
rect 17450 1325 17460 1345
rect 17480 1325 17490 1345
rect 17450 1315 17490 1325
rect 18110 1345 18150 1355
rect 18110 1325 18120 1345
rect 18140 1325 18150 1345
rect 18110 1315 18150 1325
rect 18420 1345 18460 1355
rect 18420 1325 18430 1345
rect 18450 1325 18460 1345
rect 18420 1315 18460 1325
rect 18750 1345 18790 1355
rect 18750 1325 18760 1345
rect 18780 1325 18790 1345
rect 18750 1315 18790 1325
rect 16775 1287 16845 1295
rect 16775 1215 16780 1287
rect 16800 1285 16845 1287
rect 16800 1215 16820 1285
rect 16775 1213 16820 1215
rect 16840 1213 16845 1285
rect 16775 1205 16845 1213
rect 16870 1285 16900 1295
rect 16870 1213 16875 1285
rect 16895 1213 16900 1285
rect 16870 1205 16900 1213
rect 16925 1285 16955 1295
rect 16925 1213 16930 1285
rect 16950 1213 16955 1285
rect 16925 1205 16955 1213
rect 16980 1285 17010 1295
rect 16980 1213 16985 1285
rect 17005 1213 17010 1285
rect 16980 1205 17010 1213
rect 17035 1285 17065 1295
rect 17035 1213 17040 1285
rect 17060 1213 17065 1285
rect 17035 1205 17065 1213
rect 17090 1285 17120 1295
rect 17090 1213 17095 1285
rect 17115 1213 17120 1285
rect 17090 1205 17120 1213
rect 17145 1287 17215 1295
rect 17145 1285 17190 1287
rect 17145 1213 17150 1285
rect 17170 1215 17190 1285
rect 17210 1215 17215 1287
rect 17170 1213 17215 1215
rect 17145 1205 17215 1213
rect 17415 1287 17485 1295
rect 17415 1215 17420 1287
rect 17440 1285 17485 1287
rect 17440 1215 17460 1285
rect 17480 1215 17485 1285
rect 17415 1205 17485 1215
rect 17510 1285 17540 1295
rect 17510 1215 17515 1285
rect 17535 1215 17540 1285
rect 17510 1205 17540 1215
rect 17565 1285 17595 1295
rect 17565 1215 17570 1285
rect 17590 1215 17595 1285
rect 17565 1205 17595 1215
rect 17620 1285 17650 1295
rect 17620 1215 17625 1285
rect 17645 1215 17650 1285
rect 17620 1205 17650 1215
rect 17675 1285 17705 1295
rect 17675 1215 17680 1285
rect 17700 1215 17705 1285
rect 17675 1205 17705 1215
rect 17730 1285 17760 1295
rect 17730 1215 17735 1285
rect 17755 1215 17760 1285
rect 17730 1205 17760 1215
rect 17785 1285 17815 1295
rect 17785 1215 17790 1285
rect 17810 1215 17815 1285
rect 17785 1205 17815 1215
rect 17840 1285 17870 1295
rect 17840 1215 17845 1285
rect 17865 1215 17870 1285
rect 17840 1205 17870 1215
rect 17895 1285 17925 1295
rect 17895 1215 17900 1285
rect 17920 1215 17925 1285
rect 17895 1205 17925 1215
rect 17950 1285 17980 1295
rect 17950 1215 17955 1285
rect 17975 1215 17980 1285
rect 17950 1205 17980 1215
rect 18005 1285 18035 1295
rect 18005 1215 18010 1285
rect 18030 1215 18035 1285
rect 18005 1205 18035 1215
rect 18060 1285 18090 1295
rect 18060 1215 18065 1285
rect 18085 1215 18090 1285
rect 18060 1205 18090 1215
rect 18115 1287 18185 1295
rect 18115 1285 18160 1287
rect 18115 1215 18120 1285
rect 18140 1215 18160 1285
rect 18180 1215 18185 1287
rect 18115 1205 18185 1215
rect 18385 1287 18455 1295
rect 18385 1215 18390 1287
rect 18410 1285 18455 1287
rect 18410 1215 18430 1285
rect 18385 1213 18430 1215
rect 18450 1213 18455 1285
rect 18385 1205 18455 1213
rect 18480 1285 18510 1295
rect 18480 1213 18485 1285
rect 18505 1213 18510 1285
rect 18480 1205 18510 1213
rect 18535 1285 18565 1295
rect 18535 1213 18540 1285
rect 18560 1213 18565 1285
rect 18535 1205 18565 1213
rect 18590 1285 18620 1295
rect 18590 1213 18595 1285
rect 18615 1213 18620 1285
rect 18590 1205 18620 1213
rect 18645 1285 18675 1295
rect 18645 1213 18650 1285
rect 18670 1213 18675 1285
rect 18645 1205 18675 1213
rect 18700 1285 18730 1295
rect 18700 1213 18705 1285
rect 18725 1213 18730 1285
rect 18700 1205 18730 1213
rect 18755 1287 18825 1295
rect 18755 1285 18800 1287
rect 18755 1213 18760 1285
rect 18780 1215 18800 1285
rect 18820 1215 18825 1287
rect 18780 1213 18825 1215
rect 18755 1205 18825 1213
rect 17070 1090 17100 1100
rect 17070 1070 17075 1090
rect 17095 1070 17100 1090
rect 17070 1060 17100 1070
rect 17805 1090 17835 1100
rect 17805 1070 17810 1090
rect 17830 1070 17835 1090
rect 17805 1060 17835 1070
rect 18500 1090 18530 1100
rect 18500 1070 18505 1090
rect 18525 1070 18530 1090
rect 18500 1060 18530 1070
rect 16970 835 17010 845
rect 16970 815 16980 835
rect 17000 815 17010 835
rect 16970 805 17010 815
rect 18590 835 18630 845
rect 18590 815 18600 835
rect 18620 815 18630 835
rect 18590 805 18630 815
rect 16440 775 16470 785
rect 16440 755 16445 775
rect 16465 755 16470 775
rect 16440 745 16470 755
rect 16660 775 16690 785
rect 16660 755 16665 775
rect 16685 755 16690 775
rect 16660 745 16690 755
rect 16935 775 17005 785
rect 16400 685 16470 695
rect 16400 615 16405 685
rect 16425 615 16445 685
rect 16465 615 16470 685
rect 16400 605 16470 615
rect 16495 685 16525 695
rect 16495 615 16500 685
rect 16520 615 16525 685
rect 16495 605 16525 615
rect 16550 685 16580 695
rect 16550 615 16555 685
rect 16575 615 16580 685
rect 16550 605 16580 615
rect 16605 685 16635 695
rect 16605 615 16610 685
rect 16630 615 16635 685
rect 16605 605 16635 615
rect 16660 685 16730 695
rect 16660 615 16665 685
rect 16685 615 16705 685
rect 16725 615 16730 685
rect 16660 605 16730 615
rect 16550 565 16580 575
rect 16550 545 16555 565
rect 16575 545 16580 565
rect 16550 535 16580 545
rect 16935 505 16940 775
rect 16960 505 16980 775
rect 17000 505 17005 775
rect 16935 495 17005 505
rect 17065 775 17095 785
rect 17065 505 17070 775
rect 17090 505 17095 775
rect 17065 495 17095 505
rect 17155 775 17185 785
rect 17155 505 17160 775
rect 17180 505 17185 775
rect 17155 495 17185 505
rect 17245 775 17275 785
rect 17245 505 17250 775
rect 17270 505 17275 775
rect 17245 495 17275 505
rect 17335 775 17365 785
rect 17335 505 17340 775
rect 17360 505 17365 775
rect 17335 495 17365 505
rect 17425 775 17455 785
rect 17425 505 17430 775
rect 17450 505 17455 775
rect 17425 495 17455 505
rect 17515 775 17545 785
rect 17515 505 17520 775
rect 17540 505 17545 775
rect 17515 495 17545 505
rect 17605 775 17635 785
rect 17605 505 17610 775
rect 17630 505 17635 775
rect 17605 495 17635 505
rect 17695 775 17725 785
rect 17695 505 17700 775
rect 17720 505 17725 775
rect 17695 495 17725 505
rect 17785 775 17815 785
rect 17785 505 17790 775
rect 17810 505 17815 775
rect 17785 495 17815 505
rect 17875 775 17905 785
rect 17875 505 17880 775
rect 17900 505 17905 775
rect 17875 495 17905 505
rect 17965 775 17995 785
rect 17965 505 17970 775
rect 17990 505 17995 775
rect 17965 495 17995 505
rect 18055 775 18085 785
rect 18055 505 18060 775
rect 18080 505 18085 775
rect 18055 495 18085 505
rect 18145 775 18175 785
rect 18145 505 18150 775
rect 18170 505 18175 775
rect 18145 495 18175 505
rect 18235 775 18265 785
rect 18235 505 18240 775
rect 18260 505 18265 775
rect 18235 495 18265 505
rect 18325 775 18355 785
rect 18325 505 18330 775
rect 18350 505 18355 775
rect 18325 495 18355 505
rect 18415 775 18445 785
rect 18415 505 18420 775
rect 18440 505 18445 775
rect 18415 495 18445 505
rect 18505 775 18535 785
rect 18505 505 18510 775
rect 18530 505 18535 775
rect 18505 495 18535 505
rect 18595 775 18665 785
rect 18595 505 18600 775
rect 18620 505 18640 775
rect 18660 505 18665 775
rect 18900 775 18940 785
rect 18900 755 18910 775
rect 18930 755 18940 775
rect 18900 745 18940 755
rect 19120 775 19160 785
rect 19120 755 19130 775
rect 19150 755 19160 775
rect 19120 745 19160 755
rect 18865 685 18935 695
rect 18865 615 18870 685
rect 18890 615 18910 685
rect 18930 615 18935 685
rect 18865 605 18935 615
rect 18960 685 18990 695
rect 18960 615 18965 685
rect 18985 615 18990 685
rect 18960 605 18990 615
rect 19015 685 19045 695
rect 19015 615 19020 685
rect 19040 615 19045 685
rect 19015 605 19045 615
rect 19070 685 19100 695
rect 19070 615 19075 685
rect 19095 615 19100 685
rect 19070 605 19100 615
rect 19125 685 19195 695
rect 19125 615 19130 685
rect 19150 615 19170 685
rect 19190 615 19195 685
rect 19125 605 19195 615
rect 19015 535 19045 545
rect 19015 515 19020 535
rect 19040 515 19045 535
rect 19015 505 19045 515
rect 18595 495 18665 505
rect 17695 455 17725 465
rect 17695 435 17700 455
rect 17720 435 17725 455
rect 17695 425 17725 435
rect 16425 100 16455 110
rect 16425 80 16430 100
rect 16450 80 16455 100
rect 16425 70 16455 80
rect 17625 100 17655 110
rect 17625 80 17630 100
rect 17650 80 17655 100
rect 17625 70 17655 80
rect 17945 100 17975 110
rect 17945 80 17950 100
rect 17970 80 17975 100
rect 17945 70 17975 80
rect 19145 100 19175 110
rect 19145 80 19150 100
rect 19170 80 19175 100
rect 19145 70 19175 80
rect 16385 35 16455 45
rect 16385 -35 16390 35
rect 16410 -35 16430 35
rect 16450 -35 16455 35
rect 16385 -45 16455 -35
rect 16485 35 16515 45
rect 16485 -35 16490 35
rect 16510 -35 16515 35
rect 16485 -45 16515 -35
rect 16545 35 16575 45
rect 16545 -35 16550 35
rect 16570 -35 16575 35
rect 16545 -45 16575 -35
rect 16605 35 16635 45
rect 16605 -35 16610 35
rect 16630 -35 16635 35
rect 16605 -45 16635 -35
rect 16665 35 16695 45
rect 16665 -35 16670 35
rect 16690 -35 16695 35
rect 16665 -45 16695 -35
rect 16725 35 16755 45
rect 16725 -35 16730 35
rect 16750 -35 16755 35
rect 16725 -45 16755 -35
rect 16785 35 16815 45
rect 16785 -35 16790 35
rect 16810 -35 16815 35
rect 16785 -45 16815 -35
rect 16845 35 16875 45
rect 16845 -35 16850 35
rect 16870 -35 16875 35
rect 16845 -45 16875 -35
rect 16905 35 16935 45
rect 16905 -35 16910 35
rect 16930 -35 16935 35
rect 16905 -45 16935 -35
rect 16965 35 16995 45
rect 16965 -35 16970 35
rect 16990 -35 16995 35
rect 16965 -45 16995 -35
rect 17025 35 17055 45
rect 17025 -35 17030 35
rect 17050 -35 17055 35
rect 17025 -45 17055 -35
rect 17085 35 17115 45
rect 17085 -35 17090 35
rect 17110 -35 17115 35
rect 17085 -45 17115 -35
rect 17145 35 17175 45
rect 17145 -35 17150 35
rect 17170 -35 17175 35
rect 17145 -45 17175 -35
rect 17205 35 17235 45
rect 17205 -35 17210 35
rect 17230 -35 17235 35
rect 17205 -45 17235 -35
rect 17265 35 17295 45
rect 17265 -35 17270 35
rect 17290 -35 17295 35
rect 17265 -45 17295 -35
rect 17325 35 17355 45
rect 17325 -35 17330 35
rect 17350 -35 17355 35
rect 17325 -45 17355 -35
rect 17385 35 17415 45
rect 17385 -35 17390 35
rect 17410 -35 17415 35
rect 17385 -45 17415 -35
rect 17445 35 17475 45
rect 17445 -35 17450 35
rect 17470 -35 17475 35
rect 17445 -45 17475 -35
rect 17505 35 17535 45
rect 17505 -35 17510 35
rect 17530 -35 17535 35
rect 17505 -45 17535 -35
rect 17565 35 17595 45
rect 17565 -35 17570 35
rect 17590 -35 17595 35
rect 17565 -45 17595 -35
rect 17625 35 17695 45
rect 17625 -35 17630 35
rect 17650 -35 17670 35
rect 17690 -35 17695 35
rect 17625 -45 17695 -35
rect 17905 35 17975 45
rect 17905 -35 17910 35
rect 17930 -35 17950 35
rect 17970 -35 17975 35
rect 17905 -45 17975 -35
rect 18005 35 18035 45
rect 18005 -35 18010 35
rect 18030 -35 18035 35
rect 18005 -45 18035 -35
rect 18065 35 18095 45
rect 18065 -35 18070 35
rect 18090 -35 18095 35
rect 18065 -45 18095 -35
rect 18125 35 18155 45
rect 18125 -35 18130 35
rect 18150 -35 18155 35
rect 18125 -45 18155 -35
rect 18185 35 18215 45
rect 18185 -35 18190 35
rect 18210 -35 18215 35
rect 18185 -45 18215 -35
rect 18245 35 18275 45
rect 18245 -35 18250 35
rect 18270 -35 18275 35
rect 18245 -45 18275 -35
rect 18305 35 18335 45
rect 18305 -35 18310 35
rect 18330 -35 18335 35
rect 18305 -45 18335 -35
rect 18365 35 18395 45
rect 18365 -35 18370 35
rect 18390 -35 18395 35
rect 18365 -45 18395 -35
rect 18425 35 18455 45
rect 18425 -35 18430 35
rect 18450 -35 18455 35
rect 18425 -45 18455 -35
rect 18485 35 18515 45
rect 18485 -35 18490 35
rect 18510 -35 18515 35
rect 18485 -45 18515 -35
rect 18545 35 18575 45
rect 18545 -35 18550 35
rect 18570 -35 18575 35
rect 18545 -45 18575 -35
rect 18605 35 18635 45
rect 18605 -35 18610 35
rect 18630 -35 18635 35
rect 18605 -45 18635 -35
rect 18665 35 18695 45
rect 18665 -35 18670 35
rect 18690 -35 18695 35
rect 18665 -45 18695 -35
rect 18725 35 18755 45
rect 18725 -35 18730 35
rect 18750 -35 18755 35
rect 18725 -45 18755 -35
rect 18785 35 18815 45
rect 18785 -35 18790 35
rect 18810 -35 18815 35
rect 18785 -45 18815 -35
rect 18845 35 18875 45
rect 18845 -35 18850 35
rect 18870 -35 18875 35
rect 18845 -45 18875 -35
rect 18905 35 18935 45
rect 18905 -35 18910 35
rect 18930 -35 18935 35
rect 18905 -45 18935 -35
rect 18965 35 18995 45
rect 18965 -35 18970 35
rect 18990 -35 18995 35
rect 18965 -45 18995 -35
rect 19025 35 19055 45
rect 19025 -35 19030 35
rect 19050 -35 19055 35
rect 19025 -45 19055 -35
rect 19085 35 19115 45
rect 19085 -35 19090 35
rect 19110 -35 19115 35
rect 19085 -45 19115 -35
rect 19145 35 19215 45
rect 19145 -35 19150 35
rect 19170 -35 19190 35
rect 19210 -35 19215 35
rect 19145 -45 19215 -35
rect 16600 -75 16640 -65
rect 16600 -95 16610 -75
rect 16630 -95 16640 -75
rect 16600 -105 16640 -95
rect 16960 -75 17000 -65
rect 16960 -95 16970 -75
rect 16990 -95 17000 -75
rect 16960 -105 17000 -95
rect 17320 -75 17360 -65
rect 17320 -95 17330 -75
rect 17350 -95 17360 -75
rect 17320 -105 17360 -95
rect 18240 -75 18280 -65
rect 18240 -95 18250 -75
rect 18270 -95 18280 -75
rect 18240 -105 18280 -95
rect 18600 -75 18640 -65
rect 18600 -95 18610 -75
rect 18630 -95 18640 -75
rect 18600 -105 18640 -95
rect 18960 -75 19000 -65
rect 18960 -95 18970 -75
rect 18990 -95 19000 -75
rect 18960 -105 19000 -95
rect 16540 -225 16570 -215
rect 16540 -245 16545 -225
rect 16565 -245 16570 -225
rect 16540 -255 16570 -245
rect 16900 -225 16930 -215
rect 16900 -245 16905 -225
rect 16925 -245 16930 -225
rect 16900 -255 16930 -245
rect 17260 -225 17290 -215
rect 17260 -245 17265 -225
rect 17285 -245 17290 -225
rect 17260 -255 17290 -245
rect 17510 -225 17540 -215
rect 17510 -245 17515 -225
rect 17535 -245 17540 -225
rect 17510 -255 17540 -245
rect 18060 -225 18090 -215
rect 18060 -245 18065 -225
rect 18085 -245 18090 -225
rect 18060 -255 18090 -245
rect 18310 -225 18340 -215
rect 18310 -245 18315 -225
rect 18335 -245 18340 -225
rect 18310 -255 18340 -245
rect 18670 -225 18700 -215
rect 18670 -245 18675 -225
rect 18695 -245 18700 -225
rect 18670 -255 18700 -245
rect 19030 -225 19060 -215
rect 19030 -245 19035 -225
rect 19055 -245 19060 -225
rect 19030 -255 19060 -245
rect 16800 -395 16830 -385
rect 16800 -415 16805 -395
rect 16825 -415 16830 -395
rect 16800 -425 16830 -415
rect 18770 -395 18800 -385
rect 18770 -415 18775 -395
rect 18795 -415 18800 -395
rect 18770 -425 18800 -415
rect 16855 -465 16885 -455
rect 16855 -485 16860 -465
rect 16880 -485 16885 -465
rect 16855 -495 16885 -485
rect 16915 -465 16945 -455
rect 16915 -485 16920 -465
rect 16940 -485 16945 -465
rect 16915 -495 16945 -485
rect 16975 -465 17005 -455
rect 16975 -485 16980 -465
rect 17000 -485 17005 -465
rect 16975 -495 17005 -485
rect 17035 -465 17065 -455
rect 17035 -485 17040 -465
rect 17060 -485 17065 -465
rect 17035 -495 17065 -485
rect 17095 -465 17125 -455
rect 17095 -485 17100 -465
rect 17120 -485 17125 -465
rect 17095 -495 17125 -485
rect 17155 -465 17185 -455
rect 17155 -485 17160 -465
rect 17180 -485 17185 -465
rect 17155 -495 17185 -485
rect 17215 -465 17245 -455
rect 17215 -485 17220 -465
rect 17240 -485 17245 -465
rect 17215 -495 17245 -485
rect 17275 -465 17305 -455
rect 17275 -485 17280 -465
rect 17300 -485 17305 -465
rect 17275 -495 17305 -485
rect 17335 -465 17365 -455
rect 17335 -485 17340 -465
rect 17360 -485 17365 -465
rect 17335 -495 17365 -485
rect 17395 -465 17425 -455
rect 17395 -485 17400 -465
rect 17420 -485 17425 -465
rect 17395 -495 17425 -485
rect 17455 -465 17485 -455
rect 17455 -485 17460 -465
rect 17480 -485 17485 -465
rect 17455 -495 17485 -485
rect 17565 -465 17595 -455
rect 17565 -485 17570 -465
rect 17590 -485 17595 -465
rect 17565 -495 17595 -485
rect 18005 -465 18035 -455
rect 18005 -485 18010 -465
rect 18030 -485 18035 -465
rect 18005 -495 18035 -485
rect 18115 -465 18145 -455
rect 18115 -485 18120 -465
rect 18140 -485 18145 -465
rect 18115 -495 18145 -485
rect 18175 -465 18205 -455
rect 18175 -485 18180 -465
rect 18200 -485 18205 -465
rect 18175 -495 18205 -485
rect 18235 -465 18265 -455
rect 18235 -485 18240 -465
rect 18260 -485 18265 -465
rect 18235 -495 18265 -485
rect 18295 -465 18325 -455
rect 18295 -485 18300 -465
rect 18320 -485 18325 -465
rect 18295 -495 18325 -485
rect 18355 -465 18385 -455
rect 18355 -485 18360 -465
rect 18380 -485 18385 -465
rect 18355 -495 18385 -485
rect 18415 -465 18445 -455
rect 18415 -485 18420 -465
rect 18440 -485 18445 -465
rect 18415 -495 18445 -485
rect 18475 -465 18505 -455
rect 18475 -485 18480 -465
rect 18500 -485 18505 -465
rect 18475 -495 18505 -485
rect 18535 -465 18565 -455
rect 18535 -485 18540 -465
rect 18560 -485 18565 -465
rect 18535 -495 18565 -485
rect 18595 -465 18625 -455
rect 18595 -485 18600 -465
rect 18620 -485 18625 -465
rect 18595 -495 18625 -485
rect 18655 -465 18685 -455
rect 18655 -485 18660 -465
rect 18680 -485 18685 -465
rect 18655 -495 18685 -485
rect 18715 -465 18745 -455
rect 18715 -485 18720 -465
rect 18740 -485 18745 -465
rect 18715 -495 18745 -485
rect 16800 -535 16830 -525
rect 16800 -555 16805 -535
rect 16825 -555 16830 -535
rect 16800 -565 16830 -555
rect 18770 -535 18800 -525
rect 18770 -555 18775 -535
rect 18795 -555 18800 -535
rect 18770 -565 18800 -555
rect 16800 -685 16840 -680
rect 16800 -705 16810 -685
rect 16830 -705 16840 -685
rect 16800 -715 16840 -705
rect 17420 -685 17460 -680
rect 17420 -705 17430 -685
rect 17450 -705 17460 -685
rect 17420 -715 17460 -705
rect 18140 -685 18180 -675
rect 18140 -705 18150 -685
rect 18170 -705 18180 -685
rect 18140 -715 18180 -705
rect 18760 -685 18800 -675
rect 18760 -705 18770 -685
rect 18790 -705 18800 -685
rect 18760 -715 18800 -705
rect 16535 -740 16565 -730
rect 16535 -960 16540 -740
rect 16560 -960 16565 -740
rect 16535 -970 16565 -960
rect 17075 -740 17185 -730
rect 17075 -960 17080 -740
rect 17100 -960 17120 -740
rect 17140 -960 17160 -740
rect 17180 -960 17185 -740
rect 17075 -970 17185 -960
rect 17695 -740 17725 -730
rect 17695 -960 17700 -740
rect 17720 -960 17725 -740
rect 17695 -970 17725 -960
rect 17875 -740 17905 -730
rect 17875 -960 17880 -740
rect 17900 -960 17905 -740
rect 17875 -970 17905 -960
rect 18415 -740 18525 -730
rect 18415 -960 18420 -740
rect 18440 -960 18460 -740
rect 18480 -960 18500 -740
rect 18520 -960 18525 -740
rect 18415 -970 18525 -960
rect 19035 -740 19065 -730
rect 19035 -960 19040 -740
rect 19060 -960 19065 -740
rect 19035 -970 19065 -960
rect 17260 -1100 17300 -1090
rect 17260 -1120 17270 -1100
rect 17290 -1120 17300 -1100
rect 17260 -1130 17300 -1120
rect 18300 -1100 18340 -1090
rect 18300 -1120 18310 -1100
rect 18330 -1120 18340 -1100
rect 18300 -1130 18340 -1120
rect 16745 -1160 16775 -1150
rect 16745 -1230 16750 -1160
rect 16770 -1230 16775 -1160
rect 16745 -1240 16775 -1230
rect 17785 -1160 17815 -1150
rect 17785 -1230 17790 -1160
rect 17810 -1230 17815 -1160
rect 17785 -1240 17815 -1230
rect 18825 -1160 18895 -1150
rect 18825 -1230 18830 -1160
rect 18850 -1230 18870 -1160
rect 18890 -1230 18895 -1160
rect 18825 -1240 18895 -1230
rect 17285 -1340 17315 -1330
rect 17285 -1360 17290 -1340
rect 17310 -1360 17315 -1340
rect 17285 -1370 17315 -1360
rect 17785 -1340 17815 -1330
rect 17785 -1360 17790 -1340
rect 17810 -1360 17815 -1340
rect 17785 -1370 17815 -1360
rect 18295 -1340 18325 -1330
rect 18295 -1360 18300 -1340
rect 18320 -1360 18325 -1340
rect 18295 -1370 18325 -1360
rect 16915 -1440 16955 -1430
rect 16915 -1460 16925 -1440
rect 16945 -1460 16955 -1440
rect 16915 -1470 16955 -1460
rect 17355 -1440 17395 -1430
rect 17355 -1460 17365 -1440
rect 17385 -1460 17395 -1440
rect 17355 -1470 17395 -1460
rect 17505 -1440 17545 -1430
rect 17505 -1460 17515 -1440
rect 17535 -1460 17545 -1440
rect 17505 -1470 17545 -1460
rect 18055 -1440 18095 -1430
rect 18055 -1460 18065 -1440
rect 18085 -1460 18095 -1440
rect 18055 -1470 18095 -1460
rect 18215 -1440 18255 -1430
rect 18215 -1460 18225 -1440
rect 18245 -1460 18255 -1440
rect 18215 -1470 18255 -1460
rect 18655 -1440 18695 -1430
rect 18655 -1460 18665 -1440
rect 18685 -1460 18695 -1440
rect 18655 -1470 18695 -1460
rect 16880 -1500 16950 -1490
rect 16880 -1570 16885 -1500
rect 16905 -1570 16925 -1500
rect 16945 -1570 16950 -1500
rect 16880 -1580 16950 -1570
rect 16975 -1500 17005 -1490
rect 16975 -1570 16980 -1500
rect 17000 -1570 17005 -1500
rect 16975 -1580 17005 -1570
rect 17030 -1500 17060 -1490
rect 17030 -1570 17035 -1500
rect 17055 -1570 17060 -1500
rect 17030 -1580 17060 -1570
rect 17085 -1500 17115 -1490
rect 17085 -1570 17090 -1500
rect 17110 -1570 17115 -1500
rect 17085 -1580 17115 -1570
rect 17140 -1500 17170 -1490
rect 17140 -1570 17145 -1500
rect 17165 -1570 17170 -1500
rect 17140 -1580 17170 -1570
rect 17195 -1500 17225 -1490
rect 17195 -1570 17200 -1500
rect 17220 -1570 17225 -1500
rect 17195 -1580 17225 -1570
rect 17250 -1500 17280 -1490
rect 17250 -1570 17255 -1500
rect 17275 -1570 17280 -1500
rect 17250 -1580 17280 -1570
rect 17305 -1500 17335 -1490
rect 17305 -1570 17310 -1500
rect 17330 -1570 17335 -1500
rect 17305 -1580 17335 -1570
rect 17360 -1500 17430 -1490
rect 17360 -1570 17365 -1500
rect 17385 -1570 17405 -1500
rect 17425 -1570 17430 -1500
rect 17360 -1580 17430 -1570
rect 17470 -1500 17540 -1490
rect 17470 -1570 17475 -1500
rect 17495 -1570 17515 -1500
rect 17535 -1570 17540 -1500
rect 17470 -1580 17540 -1570
rect 17565 -1500 17595 -1490
rect 17565 -1570 17570 -1500
rect 17590 -1570 17595 -1500
rect 17565 -1580 17595 -1570
rect 17620 -1500 17650 -1490
rect 17620 -1570 17625 -1500
rect 17645 -1570 17650 -1500
rect 17620 -1580 17650 -1570
rect 17675 -1500 17705 -1490
rect 17675 -1570 17680 -1500
rect 17700 -1570 17705 -1500
rect 17675 -1580 17705 -1570
rect 17730 -1500 17760 -1490
rect 17730 -1570 17735 -1500
rect 17755 -1570 17760 -1500
rect 17730 -1580 17760 -1570
rect 17785 -1500 17815 -1490
rect 17785 -1570 17790 -1500
rect 17810 -1570 17815 -1500
rect 17785 -1580 17815 -1570
rect 17840 -1500 17870 -1490
rect 17840 -1570 17845 -1500
rect 17865 -1570 17870 -1500
rect 17840 -1580 17870 -1570
rect 17895 -1500 17925 -1490
rect 17895 -1570 17900 -1500
rect 17920 -1570 17925 -1500
rect 17895 -1580 17925 -1570
rect 17950 -1500 17980 -1490
rect 17950 -1570 17955 -1500
rect 17975 -1570 17980 -1500
rect 17950 -1580 17980 -1570
rect 18005 -1500 18035 -1490
rect 18005 -1570 18010 -1500
rect 18030 -1570 18035 -1500
rect 18005 -1580 18035 -1570
rect 18060 -1500 18130 -1490
rect 18060 -1570 18065 -1500
rect 18085 -1570 18105 -1500
rect 18125 -1570 18130 -1500
rect 18060 -1580 18130 -1570
rect 18180 -1500 18250 -1490
rect 18180 -1570 18185 -1500
rect 18205 -1570 18225 -1500
rect 18245 -1570 18250 -1500
rect 18180 -1580 18250 -1570
rect 18275 -1500 18305 -1490
rect 18275 -1570 18280 -1500
rect 18300 -1570 18305 -1500
rect 18275 -1580 18305 -1570
rect 18330 -1500 18360 -1490
rect 18330 -1570 18335 -1500
rect 18355 -1570 18360 -1500
rect 18330 -1580 18360 -1570
rect 18385 -1500 18415 -1490
rect 18385 -1570 18390 -1500
rect 18410 -1570 18415 -1500
rect 18385 -1580 18415 -1570
rect 18440 -1500 18470 -1490
rect 18440 -1570 18445 -1500
rect 18465 -1570 18470 -1500
rect 18440 -1580 18470 -1570
rect 18495 -1500 18525 -1490
rect 18495 -1570 18500 -1500
rect 18520 -1570 18525 -1500
rect 18495 -1580 18525 -1570
rect 18550 -1500 18580 -1490
rect 18550 -1570 18555 -1500
rect 18575 -1570 18580 -1500
rect 18550 -1580 18580 -1570
rect 18605 -1500 18635 -1490
rect 18605 -1570 18610 -1500
rect 18630 -1570 18635 -1500
rect 18605 -1580 18635 -1570
rect 18660 -1500 18730 -1490
rect 18660 -1570 18665 -1500
rect 18685 -1570 18705 -1500
rect 18725 -1570 18730 -1500
rect 18660 -1580 18730 -1570
rect 17585 -1650 17615 -1640
rect 17585 -1670 17590 -1650
rect 17610 -1670 17615 -1650
rect 17585 -1680 17615 -1670
rect 17425 -1950 17470 -1945
rect 17425 -1975 17435 -1950
rect 17460 -1975 17470 -1950
rect 17425 -1980 17470 -1975
rect 18124 -1950 18169 -1945
rect 18124 -1975 18134 -1950
rect 18159 -1975 18169 -1950
rect 18124 -1980 18169 -1975
rect 16795 -2240 18805 -2115
rect 17440 -2795 17480 -2240
rect 18120 -2795 18160 -2240
rect 16485 -2905 16520 -2895
rect 16485 -2930 16490 -2905
rect 16515 -2930 16520 -2905
rect 16795 -2920 18805 -2795
rect 19080 -2905 19115 -2895
rect 16485 -2940 16520 -2930
rect 16160 -3030 16195 -3020
rect 16160 -3055 16165 -3030
rect 16190 -3055 16195 -3030
rect 16160 -3065 16195 -3055
rect 15950 -3121 15985 -3111
rect 15950 -3146 15955 -3121
rect 15980 -3146 15985 -3121
rect 15950 -3156 15985 -3146
rect 16255 -3100 16280 -3065
rect 16580 -2975 16605 -2940
rect 17440 -3475 17480 -2920
rect 18120 -3475 18160 -2920
rect 19080 -2930 19085 -2905
rect 19110 -2930 19115 -2905
rect 19080 -2940 19115 -2930
rect 18995 -2975 19020 -2940
rect 19405 -2997 19440 -2987
rect 19405 -3022 19410 -2997
rect 19435 -3022 19440 -2997
rect 19405 -3032 19440 -3022
rect 19320 -3067 19345 -3032
rect 19610 -3121 19645 -3111
rect 19610 -3146 19615 -3121
rect 19640 -3146 19645 -3121
rect 19610 -3156 19645 -3146
rect 16795 -3600 18805 -3475
rect 15950 -3794 15985 -3784
rect 15950 -3819 15955 -3794
rect 15980 -3819 15985 -3794
rect 15950 -3829 15985 -3819
rect 16195 -3889 16220 -3854
rect 16280 -3899 16315 -3889
rect 16280 -3924 16285 -3899
rect 16310 -3924 16315 -3899
rect 16280 -3934 16315 -3924
rect 16520 -3964 16545 -3929
rect 16605 -3974 16640 -3964
rect 16605 -3999 16610 -3974
rect 16635 -3999 16640 -3974
rect 16605 -4009 16640 -3999
rect 17440 -4125 17480 -3600
rect 17780 -4170 17820 -4120
rect 18120 -4125 18160 -3600
rect 19055 -3964 19080 -3929
rect 19380 -3889 19405 -3854
rect 19610 -3794 19645 -3784
rect 19610 -3819 19615 -3794
rect 19640 -3819 19645 -3794
rect 19610 -3829 19645 -3819
rect 19285 -3899 19320 -3889
rect 19285 -3924 19290 -3899
rect 19315 -3924 19320 -3899
rect 19285 -3934 19320 -3924
rect 18960 -3974 18995 -3964
rect 18960 -3999 18965 -3974
rect 18990 -3999 18995 -3974
rect 18960 -4009 18995 -3999
rect 17780 -4190 17790 -4170
rect 17810 -4190 17820 -4170
rect 17780 -4220 17820 -4190
rect 17780 -4240 17790 -4220
rect 17810 -4240 17820 -4220
rect 17780 -4270 17820 -4240
rect 17780 -4290 17790 -4270
rect 17810 -4290 17820 -4270
rect 17780 -4300 17820 -4290
<< viali >>
rect 16820 1325 16840 1345
rect 17150 1325 17170 1345
rect 17460 1325 17480 1345
rect 18120 1325 18140 1345
rect 18430 1325 18450 1345
rect 18760 1325 18780 1345
rect 16820 1213 16840 1285
rect 16875 1213 16895 1285
rect 16930 1213 16950 1285
rect 16985 1213 17005 1285
rect 17040 1213 17060 1285
rect 17095 1213 17115 1285
rect 17150 1213 17170 1285
rect 17460 1215 17480 1285
rect 17515 1215 17535 1285
rect 17570 1215 17590 1285
rect 17625 1215 17645 1285
rect 17680 1215 17700 1285
rect 17735 1215 17755 1285
rect 17790 1215 17810 1285
rect 17845 1215 17865 1285
rect 17900 1215 17920 1285
rect 17955 1215 17975 1285
rect 18010 1215 18030 1285
rect 18065 1215 18085 1285
rect 18120 1215 18140 1285
rect 18430 1213 18450 1285
rect 18485 1213 18505 1285
rect 18540 1213 18560 1285
rect 18595 1213 18615 1285
rect 18650 1213 18670 1285
rect 18705 1213 18725 1285
rect 18760 1213 18780 1285
rect 17075 1070 17095 1090
rect 17810 1070 17830 1090
rect 18505 1070 18525 1090
rect 16980 815 17000 835
rect 18600 815 18620 835
rect 16445 755 16465 775
rect 16665 755 16685 775
rect 16445 615 16465 685
rect 16500 615 16520 685
rect 16555 615 16575 685
rect 16610 615 16630 685
rect 16665 615 16685 685
rect 16555 545 16575 565
rect 16980 505 17000 775
rect 17070 505 17090 775
rect 17160 505 17180 775
rect 17250 505 17270 775
rect 17340 505 17360 775
rect 17430 505 17450 775
rect 17520 505 17540 775
rect 17610 505 17630 775
rect 17700 505 17720 775
rect 17790 505 17810 775
rect 17880 505 17900 775
rect 17970 505 17990 775
rect 18060 505 18080 775
rect 18150 505 18170 775
rect 18240 505 18260 775
rect 18330 505 18350 775
rect 18420 505 18440 775
rect 18510 505 18530 775
rect 18600 505 18620 775
rect 18910 755 18930 775
rect 19130 755 19150 775
rect 18910 615 18930 685
rect 18965 615 18985 685
rect 19020 615 19040 685
rect 19075 615 19095 685
rect 19130 615 19150 685
rect 19020 515 19040 535
rect 17700 435 17720 455
rect 16430 80 16450 100
rect 17630 80 17650 100
rect 17950 80 17970 100
rect 19150 80 19170 100
rect 16430 -35 16450 35
rect 16490 -35 16510 35
rect 16550 -35 16570 35
rect 16610 -35 16630 35
rect 16670 -35 16690 35
rect 16730 -35 16750 35
rect 16790 -35 16810 35
rect 16850 -35 16870 35
rect 16910 -35 16930 35
rect 16970 -35 16990 35
rect 17030 -35 17050 35
rect 17090 -35 17110 35
rect 17150 -35 17170 35
rect 17210 -35 17230 35
rect 17270 -35 17290 35
rect 17330 -35 17350 35
rect 17390 -35 17410 35
rect 17450 -35 17470 35
rect 17510 -35 17530 35
rect 17570 -35 17590 35
rect 17630 -35 17650 35
rect 17950 -35 17970 35
rect 18010 -35 18030 35
rect 18070 -35 18090 35
rect 18130 -35 18150 35
rect 18190 -35 18210 35
rect 18250 -35 18270 35
rect 18310 -35 18330 35
rect 18370 -35 18390 35
rect 18430 -35 18450 35
rect 18490 -35 18510 35
rect 18550 -35 18570 35
rect 18610 -35 18630 35
rect 18670 -35 18690 35
rect 18730 -35 18750 35
rect 18790 -35 18810 35
rect 18850 -35 18870 35
rect 18910 -35 18930 35
rect 18970 -35 18990 35
rect 19030 -35 19050 35
rect 19090 -35 19110 35
rect 19150 -35 19170 35
rect 16610 -95 16630 -75
rect 16970 -95 16990 -75
rect 17330 -95 17350 -75
rect 18250 -95 18270 -75
rect 18610 -95 18630 -75
rect 18970 -95 18990 -75
rect 16545 -245 16565 -225
rect 16905 -245 16925 -225
rect 17265 -245 17285 -225
rect 17515 -245 17535 -225
rect 18065 -245 18085 -225
rect 18315 -245 18335 -225
rect 18675 -245 18695 -225
rect 19035 -245 19055 -225
rect 16805 -415 16825 -395
rect 18775 -415 18795 -395
rect 16860 -485 16880 -465
rect 16920 -485 16940 -465
rect 16980 -485 17000 -465
rect 17040 -485 17060 -465
rect 17100 -485 17120 -465
rect 17160 -485 17180 -465
rect 17220 -485 17240 -465
rect 17280 -485 17300 -465
rect 17340 -485 17360 -465
rect 17400 -485 17420 -465
rect 17460 -485 17480 -465
rect 17570 -485 17590 -465
rect 18010 -485 18030 -465
rect 18120 -485 18140 -465
rect 18180 -485 18200 -465
rect 18240 -485 18260 -465
rect 18300 -485 18320 -465
rect 18360 -485 18380 -465
rect 18420 -485 18440 -465
rect 18480 -485 18500 -465
rect 18540 -485 18560 -465
rect 18600 -485 18620 -465
rect 18660 -485 18680 -465
rect 18720 -485 18740 -465
rect 16805 -555 16825 -535
rect 18775 -555 18795 -535
rect 16810 -705 16830 -685
rect 17430 -705 17450 -685
rect 18150 -705 18170 -685
rect 18770 -705 18790 -685
rect 16540 -960 16560 -740
rect 17080 -960 17100 -740
rect 17120 -960 17140 -740
rect 17160 -960 17180 -740
rect 17700 -960 17720 -740
rect 17880 -960 17900 -740
rect 18420 -960 18440 -740
rect 18460 -960 18480 -740
rect 18500 -960 18520 -740
rect 19040 -960 19060 -740
rect 17270 -1120 17290 -1100
rect 18310 -1120 18330 -1100
rect 16750 -1230 16770 -1160
rect 17790 -1230 17810 -1160
rect 18830 -1230 18850 -1160
rect 18870 -1230 18890 -1160
rect 17290 -1360 17310 -1340
rect 17790 -1360 17810 -1340
rect 18300 -1360 18320 -1340
rect 16925 -1460 16945 -1440
rect 17365 -1460 17385 -1440
rect 17515 -1460 17535 -1440
rect 18065 -1460 18085 -1440
rect 18225 -1460 18245 -1440
rect 18665 -1460 18685 -1440
rect 16925 -1570 16945 -1500
rect 16980 -1570 17000 -1500
rect 17035 -1570 17055 -1500
rect 17090 -1570 17110 -1500
rect 17145 -1570 17165 -1500
rect 17200 -1570 17220 -1500
rect 17255 -1570 17275 -1500
rect 17310 -1570 17330 -1500
rect 17365 -1570 17385 -1500
rect 17515 -1570 17535 -1500
rect 17570 -1570 17590 -1500
rect 17625 -1570 17645 -1500
rect 17680 -1570 17700 -1500
rect 17735 -1570 17755 -1500
rect 17790 -1570 17810 -1500
rect 17845 -1570 17865 -1500
rect 17900 -1570 17920 -1500
rect 17955 -1570 17975 -1500
rect 18010 -1570 18030 -1500
rect 18065 -1570 18085 -1500
rect 18225 -1570 18245 -1500
rect 18280 -1570 18300 -1500
rect 18335 -1570 18355 -1500
rect 18390 -1570 18410 -1500
rect 18445 -1570 18465 -1500
rect 18500 -1570 18520 -1500
rect 18555 -1570 18575 -1500
rect 18610 -1570 18630 -1500
rect 18665 -1570 18685 -1500
rect 17590 -1670 17610 -1650
rect 17435 -1975 17460 -1950
rect 18134 -1975 18159 -1950
rect 16490 -2930 16515 -2905
rect 16165 -3055 16190 -3030
rect 15955 -3146 15980 -3121
rect 19085 -2930 19110 -2905
rect 19410 -3022 19435 -2997
rect 19615 -3146 19640 -3121
rect 15955 -3819 15980 -3794
rect 16285 -3924 16310 -3899
rect 16610 -3999 16635 -3974
rect 19615 -3819 19640 -3794
rect 19290 -3924 19315 -3899
rect 18965 -3999 18990 -3974
rect 17790 -4290 17810 -4270
<< metal1 >>
rect 15725 -215 15765 -210
rect 15725 -245 15730 -215
rect 15760 -245 15765 -215
rect 15725 -250 15765 -245
rect 15735 -4310 15755 -250
rect 15795 -1340 15815 1595
rect 15950 175 15990 180
rect 15950 145 15955 175
rect 15985 145 15990 175
rect 15950 140 15990 145
rect 15785 -1345 15825 -1340
rect 15785 -1375 15790 -1345
rect 15820 -1375 15825 -1345
rect 15785 -1380 15825 -1375
rect 15820 -3115 15860 -3110
rect 15960 -3111 15980 140
rect 16040 -1685 16060 1595
rect 16030 -1690 16070 -1685
rect 16030 -1720 16035 -1690
rect 16065 -1720 16070 -1690
rect 16030 -1725 16070 -1720
rect 16115 -1820 16135 1595
rect 17095 1400 17115 1595
rect 17740 1400 17760 1595
rect 18485 1400 18505 1595
rect 16865 1395 16905 1400
rect 16865 1365 16870 1395
rect 16900 1365 16905 1395
rect 16865 1360 16905 1365
rect 16975 1395 17015 1400
rect 16975 1365 16980 1395
rect 17010 1365 17015 1395
rect 16975 1360 17015 1365
rect 17085 1395 17125 1400
rect 17085 1365 17090 1395
rect 17120 1365 17125 1395
rect 17085 1360 17125 1365
rect 17615 1395 17655 1400
rect 17615 1365 17620 1395
rect 17650 1365 17655 1395
rect 17615 1360 17655 1365
rect 17725 1395 17765 1400
rect 17725 1365 17730 1395
rect 17760 1365 17765 1395
rect 17725 1360 17765 1365
rect 17835 1395 17875 1400
rect 17835 1365 17840 1395
rect 17870 1365 17875 1395
rect 17835 1360 17875 1365
rect 17945 1395 17985 1400
rect 17945 1365 17950 1395
rect 17980 1365 17985 1395
rect 17945 1360 17985 1365
rect 18475 1395 18515 1400
rect 18475 1365 18480 1395
rect 18510 1365 18515 1395
rect 18475 1360 18515 1365
rect 18585 1395 18625 1400
rect 18585 1365 18590 1395
rect 18620 1365 18625 1395
rect 18585 1360 18625 1365
rect 18695 1395 18735 1400
rect 18695 1365 18700 1395
rect 18730 1365 18735 1395
rect 18695 1360 18735 1365
rect 16810 1350 16850 1355
rect 16810 1320 16815 1350
rect 16845 1320 16850 1350
rect 16810 1315 16850 1320
rect 16815 1285 16845 1315
rect 16815 1213 16820 1285
rect 16840 1213 16845 1285
rect 16815 1155 16845 1213
rect 16870 1285 16900 1360
rect 16920 1350 16960 1355
rect 16920 1320 16925 1350
rect 16955 1320 16960 1350
rect 16920 1315 16960 1320
rect 16870 1213 16875 1285
rect 16895 1213 16900 1285
rect 16870 1200 16900 1213
rect 16925 1285 16955 1315
rect 16925 1213 16930 1285
rect 16950 1213 16955 1285
rect 16865 1195 16905 1200
rect 16865 1165 16870 1195
rect 16900 1165 16905 1195
rect 16865 1160 16905 1165
rect 16925 1155 16955 1213
rect 16980 1285 17010 1360
rect 17030 1350 17070 1355
rect 17030 1320 17035 1350
rect 17065 1320 17070 1350
rect 17030 1315 17070 1320
rect 16980 1213 16985 1285
rect 17005 1213 17010 1285
rect 16980 1200 17010 1213
rect 17035 1285 17065 1315
rect 17035 1213 17040 1285
rect 17060 1213 17065 1285
rect 16975 1195 17015 1200
rect 16975 1165 16980 1195
rect 17010 1165 17015 1195
rect 16975 1160 17015 1165
rect 17035 1155 17065 1213
rect 17090 1285 17120 1360
rect 17140 1350 17180 1355
rect 17140 1320 17145 1350
rect 17175 1320 17180 1350
rect 17140 1315 17180 1320
rect 17450 1350 17490 1355
rect 17450 1320 17455 1350
rect 17485 1320 17490 1350
rect 17450 1315 17490 1320
rect 17560 1350 17600 1355
rect 17560 1320 17565 1350
rect 17595 1320 17600 1350
rect 17560 1315 17600 1320
rect 17090 1213 17095 1285
rect 17115 1213 17120 1285
rect 17090 1200 17120 1213
rect 17145 1285 17175 1315
rect 17145 1213 17150 1285
rect 17170 1213 17175 1285
rect 17085 1195 17125 1200
rect 17085 1165 17090 1195
rect 17120 1165 17125 1195
rect 17085 1160 17125 1165
rect 17145 1155 17175 1213
rect 17455 1285 17485 1315
rect 17455 1215 17460 1285
rect 17480 1215 17485 1285
rect 17455 1155 17485 1215
rect 17510 1285 17540 1295
rect 17510 1215 17515 1285
rect 17535 1215 17540 1285
rect 16810 1150 16850 1155
rect 16810 1120 16815 1150
rect 16845 1120 16850 1150
rect 16810 1115 16850 1120
rect 16920 1150 16960 1155
rect 16920 1120 16925 1150
rect 16955 1120 16960 1150
rect 16920 1115 16960 1120
rect 17030 1150 17070 1155
rect 17030 1120 17035 1150
rect 17065 1120 17070 1150
rect 17030 1115 17070 1120
rect 17140 1150 17180 1155
rect 17140 1120 17145 1150
rect 17175 1120 17180 1150
rect 17140 1115 17180 1120
rect 17450 1150 17490 1155
rect 17450 1120 17455 1150
rect 17485 1120 17490 1150
rect 17450 1115 17490 1120
rect 17070 1095 17100 1100
rect 17070 1060 17100 1065
rect 17510 1055 17540 1215
rect 17565 1285 17595 1315
rect 17565 1215 17570 1285
rect 17590 1215 17595 1285
rect 17565 1155 17595 1215
rect 17620 1285 17650 1360
rect 17670 1350 17710 1355
rect 17670 1320 17675 1350
rect 17705 1320 17710 1350
rect 17670 1315 17710 1320
rect 17620 1215 17625 1285
rect 17645 1215 17650 1285
rect 17620 1200 17650 1215
rect 17675 1285 17705 1315
rect 17675 1215 17680 1285
rect 17700 1215 17705 1285
rect 17615 1195 17655 1200
rect 17615 1165 17620 1195
rect 17650 1165 17655 1195
rect 17615 1160 17655 1165
rect 17675 1155 17705 1215
rect 17730 1285 17760 1360
rect 17780 1350 17820 1355
rect 17780 1320 17785 1350
rect 17815 1320 17820 1350
rect 17780 1315 17820 1320
rect 17730 1215 17735 1285
rect 17755 1215 17760 1285
rect 17730 1200 17760 1215
rect 17785 1285 17815 1315
rect 17785 1215 17790 1285
rect 17810 1215 17815 1285
rect 17725 1195 17765 1200
rect 17725 1165 17730 1195
rect 17760 1165 17765 1195
rect 17725 1160 17765 1165
rect 17785 1155 17815 1215
rect 17840 1285 17870 1360
rect 17890 1350 17930 1355
rect 17890 1320 17895 1350
rect 17925 1320 17930 1350
rect 17890 1315 17930 1320
rect 17840 1215 17845 1285
rect 17865 1215 17870 1285
rect 17840 1200 17870 1215
rect 17895 1285 17925 1315
rect 17895 1215 17900 1285
rect 17920 1215 17925 1285
rect 17835 1195 17875 1200
rect 17835 1165 17840 1195
rect 17870 1165 17875 1195
rect 17835 1160 17875 1165
rect 17895 1155 17925 1215
rect 17950 1285 17980 1360
rect 18000 1350 18040 1355
rect 18000 1320 18005 1350
rect 18035 1320 18040 1350
rect 18000 1315 18040 1320
rect 18110 1350 18150 1355
rect 18110 1320 18115 1350
rect 18145 1320 18150 1350
rect 18110 1315 18150 1320
rect 18420 1350 18460 1355
rect 18420 1320 18425 1350
rect 18455 1320 18460 1350
rect 18420 1315 18460 1320
rect 17950 1215 17955 1285
rect 17975 1215 17980 1285
rect 17950 1200 17980 1215
rect 18005 1285 18035 1315
rect 18005 1215 18010 1285
rect 18030 1215 18035 1285
rect 17945 1195 17985 1200
rect 17945 1165 17950 1195
rect 17980 1165 17985 1195
rect 17945 1160 17985 1165
rect 18005 1155 18035 1215
rect 18060 1285 18090 1295
rect 18060 1215 18065 1285
rect 18085 1215 18090 1285
rect 17560 1150 17600 1155
rect 17560 1120 17565 1150
rect 17595 1120 17600 1150
rect 17560 1115 17600 1120
rect 17670 1150 17710 1155
rect 17670 1120 17675 1150
rect 17705 1120 17710 1150
rect 17670 1115 17710 1120
rect 17780 1150 17820 1155
rect 17780 1120 17785 1150
rect 17815 1120 17820 1150
rect 17780 1115 17820 1120
rect 17890 1150 17930 1155
rect 17890 1120 17895 1150
rect 17925 1120 17930 1150
rect 17890 1115 17930 1120
rect 18000 1150 18040 1155
rect 18000 1120 18005 1150
rect 18035 1120 18040 1150
rect 18000 1115 18040 1120
rect 17805 1095 17835 1100
rect 17805 1060 17835 1065
rect 18060 1055 18090 1215
rect 18115 1285 18145 1315
rect 18115 1215 18120 1285
rect 18140 1215 18145 1285
rect 18115 1155 18145 1215
rect 18425 1285 18455 1315
rect 18425 1213 18430 1285
rect 18450 1213 18455 1285
rect 18425 1155 18455 1213
rect 18480 1285 18510 1360
rect 18530 1350 18570 1355
rect 18530 1320 18535 1350
rect 18565 1320 18570 1350
rect 18530 1315 18570 1320
rect 18480 1213 18485 1285
rect 18505 1213 18510 1285
rect 18480 1200 18510 1213
rect 18535 1285 18565 1315
rect 18535 1213 18540 1285
rect 18560 1213 18565 1285
rect 18475 1195 18515 1200
rect 18475 1165 18480 1195
rect 18510 1165 18515 1195
rect 18475 1160 18515 1165
rect 18535 1155 18565 1213
rect 18590 1285 18620 1360
rect 18640 1350 18680 1355
rect 18640 1320 18645 1350
rect 18675 1320 18680 1350
rect 18640 1315 18680 1320
rect 18590 1213 18595 1285
rect 18615 1213 18620 1285
rect 18590 1200 18620 1213
rect 18645 1285 18675 1315
rect 18645 1213 18650 1285
rect 18670 1213 18675 1285
rect 18585 1195 18625 1200
rect 18585 1165 18590 1195
rect 18620 1165 18625 1195
rect 18585 1160 18625 1165
rect 18645 1155 18675 1213
rect 18700 1285 18730 1360
rect 18750 1350 18790 1355
rect 18750 1320 18755 1350
rect 18785 1320 18790 1350
rect 18750 1315 18790 1320
rect 18700 1213 18705 1285
rect 18725 1213 18730 1285
rect 18700 1200 18730 1213
rect 18755 1285 18785 1315
rect 18755 1213 18760 1285
rect 18780 1213 18785 1285
rect 18695 1195 18735 1200
rect 18695 1165 18700 1195
rect 18730 1165 18735 1195
rect 18695 1160 18735 1165
rect 18755 1155 18785 1213
rect 18110 1150 18150 1155
rect 18110 1120 18115 1150
rect 18145 1120 18150 1150
rect 18110 1115 18150 1120
rect 18420 1150 18460 1155
rect 18420 1120 18425 1150
rect 18455 1120 18460 1150
rect 18420 1115 18460 1120
rect 18530 1150 18570 1155
rect 18530 1120 18535 1150
rect 18565 1120 18570 1150
rect 18530 1115 18570 1120
rect 18640 1150 18680 1155
rect 18640 1120 18645 1150
rect 18675 1120 18680 1150
rect 18640 1115 18680 1120
rect 18750 1150 18790 1155
rect 18750 1120 18755 1150
rect 18785 1120 18790 1150
rect 18750 1115 18790 1120
rect 18500 1095 18530 1100
rect 18500 1060 18530 1065
rect 18720 1095 18760 1100
rect 18720 1065 18725 1095
rect 18755 1065 18760 1095
rect 18720 1060 18760 1065
rect 16160 1050 16200 1055
rect 16160 1020 16165 1050
rect 16195 1020 16200 1050
rect 16160 1015 16200 1020
rect 17505 1050 17545 1055
rect 17505 1020 17510 1050
rect 17540 1020 17545 1050
rect 18055 1050 18095 1055
rect 17505 1015 17545 1020
rect 17600 1020 17640 1025
rect 16170 -1775 16190 1015
rect 17600 990 17605 1020
rect 17635 990 17640 1020
rect 17600 985 17640 990
rect 17960 1020 18000 1025
rect 17960 990 17965 1020
rect 17995 990 18000 1020
rect 18055 1020 18060 1050
rect 18090 1020 18095 1050
rect 18055 1015 18095 1020
rect 17960 985 18000 990
rect 17420 975 17460 980
rect 17420 945 17425 975
rect 17455 945 17460 975
rect 17420 940 17460 945
rect 17240 930 17280 935
rect 17240 900 17245 930
rect 17275 900 17280 930
rect 17240 895 17280 900
rect 17060 885 17100 890
rect 17060 855 17065 885
rect 17095 855 17100 885
rect 17060 850 17100 855
rect 16435 840 16475 845
rect 16435 810 16440 840
rect 16470 810 16475 840
rect 16435 805 16475 810
rect 16655 840 16695 845
rect 16655 810 16660 840
rect 16690 810 16695 840
rect 16655 805 16695 810
rect 16970 840 17010 845
rect 16970 810 16975 840
rect 17005 810 17010 840
rect 16970 805 17010 810
rect 16440 780 16470 805
rect 16440 685 16470 750
rect 16490 780 16530 785
rect 16490 750 16495 780
rect 16525 750 16530 780
rect 16490 745 16530 750
rect 16600 780 16640 785
rect 16600 750 16605 780
rect 16635 750 16640 780
rect 16600 745 16640 750
rect 16660 780 16690 805
rect 16440 615 16445 685
rect 16465 615 16470 685
rect 16440 555 16470 615
rect 16495 685 16525 745
rect 16545 735 16585 740
rect 16545 705 16550 735
rect 16580 705 16585 735
rect 16545 700 16585 705
rect 16495 615 16500 685
rect 16520 615 16525 685
rect 16495 600 16525 615
rect 16550 685 16580 700
rect 16550 615 16555 685
rect 16575 615 16580 685
rect 16550 605 16580 615
rect 16605 685 16635 745
rect 16605 615 16610 685
rect 16630 615 16635 685
rect 16605 600 16635 615
rect 16660 685 16690 750
rect 16975 775 17005 805
rect 16780 735 16820 740
rect 16780 705 16785 735
rect 16815 705 16820 735
rect 16780 700 16820 705
rect 16660 615 16665 685
rect 16685 615 16690 685
rect 16490 595 16530 600
rect 16490 565 16495 595
rect 16525 565 16530 595
rect 16600 595 16640 600
rect 16490 560 16530 565
rect 16550 565 16580 575
rect 16435 550 16475 555
rect 16435 520 16440 550
rect 16470 520 16475 550
rect 16550 545 16555 565
rect 16575 545 16580 565
rect 16600 565 16605 595
rect 16635 565 16640 595
rect 16600 560 16640 565
rect 16660 555 16690 615
rect 16550 535 16580 545
rect 16655 550 16695 555
rect 16435 515 16475 520
rect 16305 485 16345 490
rect 16305 455 16310 485
rect 16340 455 16345 485
rect 16305 450 16345 455
rect 16260 430 16300 435
rect 16260 400 16265 430
rect 16295 400 16300 430
rect 16260 395 16300 400
rect 16205 385 16245 390
rect 16205 355 16210 385
rect 16240 355 16245 385
rect 16205 350 16245 355
rect 16215 -1090 16235 350
rect 16270 -385 16290 395
rect 16260 -390 16300 -385
rect 16260 -420 16265 -390
rect 16295 -420 16300 -390
rect 16260 -425 16300 -420
rect 16205 -1095 16245 -1090
rect 16205 -1125 16210 -1095
rect 16240 -1125 16245 -1095
rect 16205 -1130 16245 -1125
rect 16160 -1780 16200 -1775
rect 16160 -1810 16165 -1780
rect 16195 -1810 16200 -1780
rect 16160 -1815 16200 -1810
rect 16105 -1825 16145 -1820
rect 16105 -1855 16110 -1825
rect 16140 -1855 16145 -1825
rect 16105 -1860 16145 -1855
rect 16155 -1900 16195 -1895
rect 16155 -1930 16160 -1900
rect 16190 -1930 16195 -1900
rect 16155 -1935 16195 -1930
rect 16165 -3020 16185 -1935
rect 16270 -1940 16290 -425
rect 16315 -525 16335 450
rect 16555 390 16575 535
rect 16655 520 16660 550
rect 16690 520 16695 550
rect 16655 515 16695 520
rect 16790 435 16810 700
rect 16840 595 16880 600
rect 16840 565 16845 595
rect 16875 565 16880 595
rect 16840 560 16880 565
rect 16780 430 16820 435
rect 16780 400 16785 430
rect 16815 400 16820 430
rect 16780 395 16820 400
rect 16545 385 16585 390
rect 16545 355 16550 385
rect 16580 355 16585 385
rect 16545 350 16585 355
rect 16420 225 16460 230
rect 16420 195 16425 225
rect 16455 195 16460 225
rect 16420 190 16460 195
rect 16540 225 16580 230
rect 16540 195 16545 225
rect 16575 195 16580 225
rect 16540 190 16580 195
rect 16660 225 16700 230
rect 16660 195 16665 225
rect 16695 195 16700 225
rect 16660 190 16700 195
rect 16780 225 16820 230
rect 16780 195 16785 225
rect 16815 195 16820 225
rect 16780 190 16820 195
rect 16425 100 16455 190
rect 16480 175 16520 180
rect 16480 145 16485 175
rect 16515 145 16520 175
rect 16480 140 16520 145
rect 16425 80 16430 100
rect 16450 80 16455 100
rect 16425 35 16455 80
rect 16425 -35 16430 35
rect 16450 -35 16455 35
rect 16425 -160 16455 -35
rect 16485 35 16515 140
rect 16485 -35 16490 35
rect 16510 -35 16515 35
rect 16485 -110 16515 -35
rect 16545 35 16575 190
rect 16600 85 16640 90
rect 16600 55 16605 85
rect 16635 55 16640 85
rect 16600 50 16640 55
rect 16545 -35 16550 35
rect 16570 -35 16575 35
rect 16480 -115 16520 -110
rect 16480 -145 16485 -115
rect 16515 -145 16520 -115
rect 16480 -150 16520 -145
rect 16545 -160 16575 -35
rect 16605 35 16635 50
rect 16605 -35 16610 35
rect 16630 -35 16635 35
rect 16605 -65 16635 -35
rect 16665 35 16695 190
rect 16720 130 16760 135
rect 16720 100 16725 130
rect 16755 100 16760 130
rect 16720 95 16760 100
rect 16665 -35 16670 35
rect 16690 -35 16695 35
rect 16600 -70 16640 -65
rect 16600 -100 16605 -70
rect 16635 -100 16640 -70
rect 16600 -105 16640 -100
rect 16665 -160 16695 -35
rect 16725 35 16755 95
rect 16725 -35 16730 35
rect 16750 -35 16755 35
rect 16420 -165 16460 -160
rect 16420 -195 16425 -165
rect 16455 -195 16460 -165
rect 16420 -200 16460 -195
rect 16540 -165 16580 -160
rect 16540 -195 16545 -165
rect 16575 -195 16580 -165
rect 16540 -200 16580 -195
rect 16660 -165 16700 -160
rect 16660 -195 16665 -165
rect 16695 -195 16700 -165
rect 16660 -200 16700 -195
rect 16725 -215 16755 -35
rect 16785 35 16815 190
rect 16850 180 16870 560
rect 16975 505 16980 775
rect 17000 505 17005 775
rect 16975 495 17005 505
rect 17065 775 17095 850
rect 17150 840 17190 845
rect 17150 810 17155 840
rect 17185 810 17190 840
rect 17150 805 17190 810
rect 17065 505 17070 775
rect 17090 505 17095 775
rect 17065 345 17095 505
rect 17155 775 17185 805
rect 17155 505 17160 775
rect 17180 505 17185 775
rect 17155 495 17185 505
rect 17245 775 17275 895
rect 17330 840 17370 845
rect 17330 810 17335 840
rect 17365 810 17370 840
rect 17330 805 17370 810
rect 17245 505 17250 775
rect 17270 505 17275 775
rect 17245 390 17275 505
rect 17335 775 17365 805
rect 17335 505 17340 775
rect 17360 505 17365 775
rect 17335 495 17365 505
rect 17425 775 17455 940
rect 17510 840 17550 845
rect 17510 810 17515 840
rect 17545 810 17550 840
rect 17510 805 17550 810
rect 17425 505 17430 775
rect 17450 505 17455 775
rect 17425 435 17455 505
rect 17515 775 17545 805
rect 17515 505 17520 775
rect 17540 505 17545 775
rect 17515 495 17545 505
rect 17605 775 17635 985
rect 17780 885 17820 890
rect 17780 855 17785 885
rect 17815 855 17820 885
rect 17780 850 17820 855
rect 17690 840 17730 845
rect 17690 810 17695 840
rect 17725 810 17730 840
rect 17690 805 17730 810
rect 17605 505 17610 775
rect 17630 505 17635 775
rect 17605 490 17635 505
rect 17695 775 17725 805
rect 17695 505 17700 775
rect 17720 505 17725 775
rect 17695 495 17725 505
rect 17785 775 17815 850
rect 17870 840 17910 845
rect 17870 810 17875 840
rect 17905 810 17910 840
rect 17870 805 17910 810
rect 17785 505 17790 775
rect 17810 505 17815 775
rect 17600 485 17640 490
rect 17600 455 17605 485
rect 17635 455 17640 485
rect 17600 450 17640 455
rect 17695 455 17725 465
rect 17695 435 17700 455
rect 17720 435 17725 455
rect 17420 430 17460 435
rect 17420 400 17425 430
rect 17455 400 17460 430
rect 17695 425 17725 435
rect 17420 395 17460 400
rect 17240 385 17280 390
rect 17240 355 17245 385
rect 17275 355 17280 385
rect 17240 350 17280 355
rect 17060 340 17100 345
rect 17060 310 17065 340
rect 17095 310 17100 340
rect 17060 305 17100 310
rect 16900 225 16940 230
rect 16900 195 16905 225
rect 16935 195 16940 225
rect 16900 190 16940 195
rect 17020 225 17060 230
rect 17020 195 17025 225
rect 17055 195 17060 225
rect 17020 190 17060 195
rect 17140 225 17180 230
rect 17140 195 17145 225
rect 17175 195 17180 225
rect 17140 190 17180 195
rect 17260 225 17300 230
rect 17260 195 17265 225
rect 17295 195 17300 225
rect 17260 190 17300 195
rect 17380 225 17420 230
rect 17380 195 17385 225
rect 17415 195 17420 225
rect 17380 190 17420 195
rect 17500 225 17540 230
rect 17500 195 17505 225
rect 17535 195 17540 225
rect 17500 190 17540 195
rect 17620 225 17660 230
rect 17620 195 17625 225
rect 17655 195 17660 225
rect 17620 190 17660 195
rect 16840 175 16880 180
rect 16840 145 16845 175
rect 16875 145 16880 175
rect 16840 140 16880 145
rect 16785 -35 16790 35
rect 16810 -35 16815 35
rect 16785 -160 16815 -35
rect 16845 35 16875 140
rect 16845 -35 16850 35
rect 16870 -35 16875 35
rect 16845 -110 16875 -35
rect 16905 35 16935 190
rect 16960 85 17000 90
rect 16960 55 16965 85
rect 16995 55 17000 85
rect 16960 50 17000 55
rect 16905 -35 16910 35
rect 16930 -35 16935 35
rect 16840 -115 16880 -110
rect 16840 -145 16845 -115
rect 16875 -145 16880 -115
rect 16840 -150 16880 -145
rect 16905 -160 16935 -35
rect 16965 35 16995 50
rect 16965 -35 16970 35
rect 16990 -35 16995 35
rect 16965 -65 16995 -35
rect 17025 35 17055 190
rect 17080 130 17120 135
rect 17080 100 17085 130
rect 17115 100 17120 130
rect 17080 95 17120 100
rect 17025 -35 17030 35
rect 17050 -35 17055 35
rect 16960 -70 17000 -65
rect 16960 -100 16965 -70
rect 16995 -100 17000 -70
rect 16960 -105 17000 -100
rect 16780 -165 16820 -160
rect 16780 -195 16785 -165
rect 16815 -195 16820 -165
rect 16780 -200 16820 -195
rect 16900 -165 16940 -160
rect 16900 -195 16905 -165
rect 16935 -195 16940 -165
rect 16900 -200 16940 -195
rect 16540 -220 16570 -215
rect 16540 -255 16570 -250
rect 16720 -220 16760 -215
rect 16720 -250 16725 -220
rect 16755 -250 16760 -220
rect 16720 -255 16760 -250
rect 16900 -220 16930 -215
rect 16900 -255 16930 -250
rect 16910 -325 16950 -320
rect 16910 -355 16915 -325
rect 16945 -355 16950 -325
rect 16910 -360 16950 -355
rect 16800 -390 16830 -385
rect 16800 -425 16830 -420
rect 16850 -415 16890 -410
rect 16850 -445 16855 -415
rect 16885 -445 16890 -415
rect 16850 -450 16890 -445
rect 16855 -465 16885 -450
rect 16855 -485 16860 -465
rect 16880 -485 16885 -465
rect 16305 -530 16345 -525
rect 16305 -560 16310 -530
rect 16340 -560 16345 -530
rect 16305 -565 16345 -560
rect 16800 -530 16830 -525
rect 16855 -545 16885 -485
rect 16915 -465 16945 -360
rect 16980 -365 17000 -105
rect 17025 -160 17055 -35
rect 17085 35 17115 95
rect 17085 -35 17090 35
rect 17110 -35 17115 35
rect 17020 -165 17060 -160
rect 17020 -195 17025 -165
rect 17055 -195 17060 -165
rect 17020 -200 17060 -195
rect 17085 -215 17115 -35
rect 17145 35 17175 190
rect 17200 175 17240 180
rect 17200 145 17205 175
rect 17235 145 17240 175
rect 17200 140 17240 145
rect 17145 -35 17150 35
rect 17170 -35 17175 35
rect 17145 -160 17175 -35
rect 17205 35 17235 140
rect 17205 -35 17210 35
rect 17230 -35 17235 35
rect 17205 -110 17235 -35
rect 17265 35 17295 190
rect 17320 85 17360 90
rect 17320 55 17325 85
rect 17355 55 17360 85
rect 17320 50 17360 55
rect 17265 -35 17270 35
rect 17290 -35 17295 35
rect 17200 -115 17240 -110
rect 17200 -145 17205 -115
rect 17235 -145 17240 -115
rect 17200 -150 17240 -145
rect 17265 -160 17295 -35
rect 17325 35 17355 50
rect 17325 -35 17330 35
rect 17350 -35 17355 35
rect 17325 -65 17355 -35
rect 17385 35 17415 190
rect 17440 130 17480 135
rect 17440 100 17445 130
rect 17475 100 17480 130
rect 17440 95 17480 100
rect 17385 -35 17390 35
rect 17410 -35 17415 35
rect 17320 -70 17360 -65
rect 17320 -100 17325 -70
rect 17355 -100 17360 -70
rect 17320 -105 17360 -100
rect 17385 -160 17415 -35
rect 17445 35 17475 95
rect 17445 -35 17450 35
rect 17470 -35 17475 35
rect 17140 -165 17180 -160
rect 17140 -195 17145 -165
rect 17175 -195 17180 -165
rect 17140 -200 17180 -195
rect 17260 -165 17300 -160
rect 17260 -195 17265 -165
rect 17295 -195 17300 -165
rect 17260 -200 17300 -195
rect 17380 -165 17420 -160
rect 17380 -195 17385 -165
rect 17415 -195 17420 -165
rect 17380 -200 17420 -195
rect 17445 -215 17475 -35
rect 17505 35 17535 190
rect 17560 175 17600 180
rect 17560 145 17565 175
rect 17595 145 17600 175
rect 17560 140 17600 145
rect 17505 -35 17510 35
rect 17530 -35 17535 35
rect 17505 -160 17535 -35
rect 17565 35 17595 140
rect 17565 -35 17570 35
rect 17590 -35 17595 35
rect 17565 -110 17595 -35
rect 17625 100 17655 190
rect 17700 180 17720 425
rect 17785 345 17815 505
rect 17875 775 17905 805
rect 17875 505 17880 775
rect 17900 505 17905 775
rect 17875 495 17905 505
rect 17965 775 17995 985
rect 18140 975 18180 980
rect 18140 945 18145 975
rect 18175 945 18180 975
rect 18140 940 18180 945
rect 18050 840 18090 845
rect 18050 810 18055 840
rect 18085 810 18090 840
rect 18050 805 18090 810
rect 17965 505 17970 775
rect 17990 505 17995 775
rect 17965 490 17995 505
rect 18055 775 18085 805
rect 18055 505 18060 775
rect 18080 505 18085 775
rect 18055 495 18085 505
rect 18145 775 18175 940
rect 18320 930 18360 935
rect 18320 900 18325 930
rect 18355 900 18360 930
rect 18320 895 18360 900
rect 18230 840 18270 845
rect 18230 810 18235 840
rect 18265 810 18270 840
rect 18230 805 18270 810
rect 18145 505 18150 775
rect 18170 505 18175 775
rect 17960 485 18000 490
rect 17960 455 17965 485
rect 17995 455 18000 485
rect 17960 450 18000 455
rect 18145 435 18175 505
rect 18235 775 18265 805
rect 18235 505 18240 775
rect 18260 505 18265 775
rect 18235 495 18265 505
rect 18325 775 18355 895
rect 18500 885 18540 890
rect 18500 855 18505 885
rect 18535 855 18540 885
rect 18500 850 18540 855
rect 18410 840 18450 845
rect 18410 810 18415 840
rect 18445 810 18450 840
rect 18410 805 18450 810
rect 18325 505 18330 775
rect 18350 505 18355 775
rect 18140 430 18180 435
rect 18140 400 18145 430
rect 18175 400 18180 430
rect 18140 395 18180 400
rect 18325 390 18355 505
rect 18415 775 18445 805
rect 18415 505 18420 775
rect 18440 505 18445 775
rect 18415 495 18445 505
rect 18505 775 18535 850
rect 18590 840 18630 845
rect 18590 810 18595 840
rect 18625 810 18630 840
rect 18590 805 18630 810
rect 18505 505 18510 775
rect 18530 505 18535 775
rect 18320 385 18360 390
rect 18320 355 18325 385
rect 18355 355 18360 385
rect 18320 350 18360 355
rect 18505 345 18535 505
rect 18595 775 18625 785
rect 18595 505 18600 775
rect 18620 505 18625 775
rect 18595 495 18625 505
rect 17780 340 17820 345
rect 17780 310 17785 340
rect 17815 310 17820 340
rect 17780 305 17820 310
rect 18500 340 18540 345
rect 18500 310 18505 340
rect 18535 310 18540 340
rect 18500 305 18540 310
rect 18730 285 18750 1060
rect 19010 840 19050 845
rect 19010 810 19015 840
rect 19045 810 19050 840
rect 19010 805 19050 810
rect 19020 785 19040 805
rect 18900 780 18940 785
rect 18900 750 18905 780
rect 18935 750 18940 780
rect 18900 745 18940 750
rect 19010 780 19050 785
rect 19010 750 19015 780
rect 19045 750 19050 780
rect 19010 745 19050 750
rect 19120 780 19160 785
rect 19120 750 19125 780
rect 19155 750 19160 780
rect 19120 745 19160 750
rect 18905 685 18935 745
rect 18955 735 18995 740
rect 18955 705 18960 735
rect 18990 705 18995 735
rect 18955 700 18995 705
rect 18905 615 18910 685
rect 18930 615 18935 685
rect 18905 600 18935 615
rect 18960 685 18990 700
rect 18960 615 18965 685
rect 18985 615 18990 685
rect 18900 595 18940 600
rect 18900 565 18905 595
rect 18935 565 18940 595
rect 18900 560 18940 565
rect 18960 555 18990 615
rect 19015 685 19045 745
rect 19065 735 19105 740
rect 19065 705 19070 735
rect 19100 705 19105 735
rect 19065 700 19105 705
rect 19015 615 19020 685
rect 19040 615 19045 685
rect 19015 600 19045 615
rect 19070 685 19100 700
rect 19070 615 19075 685
rect 19095 615 19100 685
rect 19010 595 19050 600
rect 19010 565 19015 595
rect 19045 565 19050 595
rect 19010 560 19050 565
rect 19070 555 19100 615
rect 19125 685 19155 745
rect 19125 615 19130 685
rect 19150 615 19155 685
rect 19125 600 19155 615
rect 19120 595 19160 600
rect 19120 565 19125 595
rect 19155 565 19160 595
rect 19120 560 19160 565
rect 19270 555 19290 1595
rect 19325 1050 19365 1055
rect 19325 1020 19330 1050
rect 19360 1020 19365 1050
rect 19325 1015 19365 1020
rect 18955 550 18995 555
rect 18955 520 18960 550
rect 18990 520 18995 550
rect 19065 550 19105 555
rect 18955 515 18995 520
rect 19015 535 19045 545
rect 19015 515 19020 535
rect 19040 515 19045 535
rect 19065 520 19070 550
rect 19100 520 19105 550
rect 19065 515 19105 520
rect 19260 550 19300 555
rect 19260 520 19265 550
rect 19295 520 19300 550
rect 19260 515 19300 520
rect 19015 505 19045 515
rect 19020 285 19040 505
rect 18720 280 18760 285
rect 18720 250 18725 280
rect 18755 250 18760 280
rect 18720 245 18760 250
rect 19010 280 19050 285
rect 19010 250 19015 280
rect 19045 250 19050 280
rect 19010 245 19050 250
rect 17940 225 17980 230
rect 17940 195 17945 225
rect 17975 195 17980 225
rect 17940 190 17980 195
rect 18060 225 18100 230
rect 18060 195 18065 225
rect 18095 195 18100 225
rect 18060 190 18100 195
rect 18180 225 18220 230
rect 18180 195 18185 225
rect 18215 195 18220 225
rect 18180 190 18220 195
rect 18300 225 18340 230
rect 18300 195 18305 225
rect 18335 195 18340 225
rect 18300 190 18340 195
rect 18420 225 18460 230
rect 18420 195 18425 225
rect 18455 195 18460 225
rect 18420 190 18460 195
rect 18540 225 18580 230
rect 18540 195 18545 225
rect 18575 195 18580 225
rect 18540 190 18580 195
rect 18660 225 18700 230
rect 18660 195 18665 225
rect 18695 195 18700 225
rect 18660 190 18700 195
rect 17690 175 17730 180
rect 17690 145 17695 175
rect 17725 145 17730 175
rect 17690 140 17730 145
rect 17870 175 17910 180
rect 17870 145 17875 175
rect 17905 145 17910 175
rect 17870 140 17910 145
rect 17625 80 17630 100
rect 17650 80 17655 100
rect 17625 35 17655 80
rect 17625 -35 17630 35
rect 17650 -35 17655 35
rect 17560 -115 17600 -110
rect 17560 -145 17565 -115
rect 17595 -145 17600 -115
rect 17560 -150 17600 -145
rect 17625 -160 17655 -35
rect 17500 -165 17540 -160
rect 17500 -195 17505 -165
rect 17535 -195 17540 -165
rect 17500 -200 17540 -195
rect 17620 -165 17660 -160
rect 17620 -195 17625 -165
rect 17655 -195 17660 -165
rect 17620 -200 17660 -195
rect 17080 -220 17120 -215
rect 17080 -250 17085 -220
rect 17115 -250 17120 -220
rect 17080 -255 17120 -250
rect 17260 -220 17290 -215
rect 17260 -255 17290 -250
rect 17440 -220 17480 -215
rect 17440 -250 17445 -220
rect 17475 -250 17480 -220
rect 17440 -255 17480 -250
rect 17510 -220 17540 -215
rect 17510 -255 17540 -250
rect 17030 -325 17070 -320
rect 17030 -355 17035 -325
rect 17065 -355 17070 -325
rect 17030 -360 17070 -355
rect 16970 -370 17010 -365
rect 16970 -400 16975 -370
rect 17005 -400 17010 -370
rect 16970 -405 17010 -400
rect 16915 -485 16920 -465
rect 16940 -485 16945 -465
rect 16800 -565 16830 -560
rect 16850 -550 16890 -545
rect 16850 -580 16855 -550
rect 16885 -580 16890 -550
rect 16850 -585 16890 -580
rect 16915 -590 16945 -485
rect 16975 -465 17005 -405
rect 16975 -485 16980 -465
rect 17000 -485 17005 -465
rect 16975 -500 17005 -485
rect 17035 -465 17065 -360
rect 17090 -410 17110 -255
rect 17150 -325 17190 -320
rect 17150 -355 17155 -325
rect 17185 -355 17190 -325
rect 17150 -360 17190 -355
rect 17270 -325 17310 -320
rect 17270 -355 17275 -325
rect 17305 -355 17310 -325
rect 17270 -360 17310 -355
rect 17390 -325 17430 -320
rect 17390 -355 17395 -325
rect 17425 -355 17430 -325
rect 17390 -360 17430 -355
rect 17090 -415 17130 -410
rect 17090 -445 17095 -415
rect 17125 -445 17130 -415
rect 17090 -450 17130 -445
rect 17035 -485 17040 -465
rect 17060 -485 17065 -465
rect 16970 -505 17010 -500
rect 16970 -535 16975 -505
rect 17005 -535 17010 -505
rect 16970 -540 17010 -535
rect 17035 -590 17065 -485
rect 17095 -465 17125 -450
rect 17095 -485 17100 -465
rect 17120 -485 17125 -465
rect 17095 -545 17125 -485
rect 17155 -465 17185 -360
rect 17210 -370 17250 -365
rect 17210 -400 17215 -370
rect 17245 -400 17250 -370
rect 17210 -405 17250 -400
rect 17155 -485 17160 -465
rect 17180 -485 17185 -465
rect 17090 -550 17130 -545
rect 17090 -580 17095 -550
rect 17125 -580 17130 -550
rect 17090 -585 17130 -580
rect 17155 -590 17185 -485
rect 17215 -465 17245 -405
rect 17215 -485 17220 -465
rect 17240 -485 17245 -465
rect 17215 -500 17245 -485
rect 17275 -465 17305 -360
rect 17330 -415 17370 -410
rect 17330 -445 17335 -415
rect 17365 -445 17370 -415
rect 17330 -450 17370 -445
rect 17275 -485 17280 -465
rect 17300 -485 17305 -465
rect 17210 -505 17250 -500
rect 17210 -535 17215 -505
rect 17245 -535 17250 -505
rect 17210 -540 17250 -535
rect 17275 -590 17305 -485
rect 17335 -465 17365 -450
rect 17335 -485 17340 -465
rect 17360 -485 17365 -465
rect 17335 -545 17365 -485
rect 17395 -465 17425 -360
rect 17450 -370 17490 -365
rect 17450 -400 17455 -370
rect 17485 -400 17490 -370
rect 17450 -405 17490 -400
rect 17395 -485 17400 -465
rect 17420 -485 17425 -465
rect 17330 -550 17370 -545
rect 17330 -580 17335 -550
rect 17365 -580 17370 -550
rect 17330 -585 17370 -580
rect 17395 -590 17425 -485
rect 17455 -465 17485 -405
rect 17455 -485 17460 -465
rect 17480 -485 17485 -465
rect 17455 -500 17485 -485
rect 17565 -460 17595 -455
rect 17565 -495 17595 -490
rect 17450 -505 17490 -500
rect 17450 -535 17455 -505
rect 17485 -535 17490 -505
rect 17450 -540 17490 -535
rect 16530 -595 16570 -590
rect 16530 -625 16535 -595
rect 16565 -625 16570 -595
rect 16530 -630 16570 -625
rect 16910 -595 16950 -590
rect 16910 -625 16915 -595
rect 16945 -625 16950 -595
rect 16910 -630 16950 -625
rect 17030 -595 17070 -590
rect 17030 -625 17035 -595
rect 17065 -625 17070 -595
rect 17030 -630 17070 -625
rect 17150 -595 17190 -590
rect 17150 -625 17155 -595
rect 17185 -625 17190 -595
rect 17150 -630 17190 -625
rect 17270 -595 17310 -590
rect 17270 -625 17275 -595
rect 17305 -625 17310 -595
rect 17270 -630 17310 -625
rect 17390 -595 17430 -590
rect 17390 -625 17395 -595
rect 17425 -625 17430 -595
rect 17390 -630 17430 -625
rect 16535 -740 16565 -630
rect 16800 -680 16840 -675
rect 16800 -710 16805 -680
rect 16835 -710 16840 -680
rect 16800 -715 16840 -710
rect 17420 -680 17460 -675
rect 17420 -710 17425 -680
rect 17455 -710 17460 -680
rect 17420 -715 17460 -710
rect 17700 -730 17720 140
rect 17780 -460 17820 -455
rect 17780 -490 17785 -460
rect 17815 -490 17820 -460
rect 17780 -495 17820 -490
rect 16535 -960 16540 -740
rect 16560 -960 16565 -740
rect 16535 -970 16565 -960
rect 17075 -740 17185 -730
rect 17075 -960 17080 -740
rect 17100 -960 17120 -740
rect 17140 -960 17160 -740
rect 17180 -960 17185 -740
rect 17075 -970 17185 -960
rect 17695 -740 17725 -730
rect 17695 -960 17700 -740
rect 17720 -960 17725 -740
rect 17695 -970 17725 -960
rect 17115 -990 17145 -970
rect 17790 -990 17810 -495
rect 17880 -730 17900 140
rect 17945 100 17975 190
rect 18000 175 18040 180
rect 18000 145 18005 175
rect 18035 145 18040 175
rect 18000 140 18040 145
rect 17945 80 17950 100
rect 17970 80 17975 100
rect 17945 35 17975 80
rect 17945 -35 17950 35
rect 17970 -35 17975 35
rect 17945 -160 17975 -35
rect 18005 35 18035 140
rect 18005 -35 18010 35
rect 18030 -35 18035 35
rect 18005 -110 18035 -35
rect 18065 35 18095 190
rect 18120 130 18160 135
rect 18120 100 18125 130
rect 18155 100 18160 130
rect 18120 95 18160 100
rect 18065 -35 18070 35
rect 18090 -35 18095 35
rect 18000 -115 18040 -110
rect 18000 -145 18005 -115
rect 18035 -145 18040 -115
rect 18000 -150 18040 -145
rect 18065 -160 18095 -35
rect 18125 35 18155 95
rect 18125 -35 18130 35
rect 18150 -35 18155 35
rect 17940 -165 17980 -160
rect 17940 -195 17945 -165
rect 17975 -195 17980 -165
rect 17940 -200 17980 -195
rect 18060 -165 18100 -160
rect 18060 -195 18065 -165
rect 18095 -195 18100 -165
rect 18060 -200 18100 -195
rect 18125 -215 18155 -35
rect 18185 35 18215 190
rect 18240 85 18280 90
rect 18240 55 18245 85
rect 18275 55 18280 85
rect 18240 50 18280 55
rect 18185 -35 18190 35
rect 18210 -35 18215 35
rect 18185 -160 18215 -35
rect 18245 35 18275 50
rect 18245 -35 18250 35
rect 18270 -35 18275 35
rect 18245 -65 18275 -35
rect 18305 35 18335 190
rect 18360 175 18400 180
rect 18360 145 18365 175
rect 18395 145 18400 175
rect 18360 140 18400 145
rect 18305 -35 18310 35
rect 18330 -35 18335 35
rect 18240 -70 18280 -65
rect 18240 -100 18245 -70
rect 18275 -100 18280 -70
rect 18240 -105 18280 -100
rect 18305 -160 18335 -35
rect 18365 35 18395 140
rect 18365 -35 18370 35
rect 18390 -35 18395 35
rect 18365 -110 18395 -35
rect 18425 35 18455 190
rect 18480 130 18520 135
rect 18480 100 18485 130
rect 18515 100 18520 130
rect 18480 95 18520 100
rect 18425 -35 18430 35
rect 18450 -35 18455 35
rect 18360 -115 18400 -110
rect 18360 -145 18365 -115
rect 18395 -145 18400 -115
rect 18360 -150 18400 -145
rect 18425 -160 18455 -35
rect 18485 35 18515 95
rect 18485 -35 18490 35
rect 18510 -35 18515 35
rect 18180 -165 18220 -160
rect 18180 -195 18185 -165
rect 18215 -195 18220 -165
rect 18180 -200 18220 -195
rect 18300 -165 18340 -160
rect 18300 -195 18305 -165
rect 18335 -195 18340 -165
rect 18300 -200 18340 -195
rect 18420 -165 18460 -160
rect 18420 -195 18425 -165
rect 18455 -195 18460 -165
rect 18420 -200 18460 -195
rect 18485 -215 18515 -35
rect 18545 35 18575 190
rect 18600 85 18640 90
rect 18600 55 18605 85
rect 18635 55 18640 85
rect 18600 50 18640 55
rect 18545 -35 18550 35
rect 18570 -35 18575 35
rect 18545 -160 18575 -35
rect 18605 35 18635 50
rect 18605 -35 18610 35
rect 18630 -35 18635 35
rect 18605 -65 18635 -35
rect 18665 35 18695 190
rect 18730 180 18750 245
rect 18780 225 18820 230
rect 18780 195 18785 225
rect 18815 195 18820 225
rect 18780 190 18820 195
rect 18900 225 18940 230
rect 18900 195 18905 225
rect 18935 195 18940 225
rect 18900 190 18940 195
rect 19020 225 19060 230
rect 19020 195 19025 225
rect 19055 195 19060 225
rect 19020 190 19060 195
rect 19140 225 19180 230
rect 19140 195 19145 225
rect 19175 195 19180 225
rect 19140 190 19180 195
rect 18720 175 18760 180
rect 18720 145 18725 175
rect 18755 145 18760 175
rect 18720 140 18760 145
rect 18665 -35 18670 35
rect 18690 -35 18695 35
rect 18600 -70 18640 -65
rect 18600 -100 18605 -70
rect 18635 -100 18640 -70
rect 18600 -105 18640 -100
rect 18540 -165 18580 -160
rect 18540 -195 18545 -165
rect 18575 -195 18580 -165
rect 18540 -200 18580 -195
rect 18060 -220 18090 -215
rect 18060 -255 18090 -250
rect 18120 -220 18160 -215
rect 18120 -250 18125 -220
rect 18155 -250 18160 -220
rect 18120 -255 18160 -250
rect 18310 -220 18340 -215
rect 18310 -255 18340 -250
rect 18480 -220 18520 -215
rect 18480 -250 18485 -220
rect 18515 -250 18520 -220
rect 18480 -255 18520 -250
rect 18170 -325 18210 -320
rect 18170 -355 18175 -325
rect 18205 -355 18210 -325
rect 18170 -360 18210 -355
rect 18290 -325 18330 -320
rect 18290 -355 18295 -325
rect 18325 -355 18330 -325
rect 18290 -360 18330 -355
rect 18410 -325 18450 -320
rect 18410 -355 18415 -325
rect 18445 -355 18450 -325
rect 18410 -360 18450 -355
rect 18110 -370 18150 -365
rect 18110 -400 18115 -370
rect 18145 -400 18150 -370
rect 18110 -405 18150 -400
rect 18005 -460 18035 -455
rect 18005 -495 18035 -490
rect 18115 -465 18145 -405
rect 18115 -485 18120 -465
rect 18140 -485 18145 -465
rect 18115 -500 18145 -485
rect 18175 -465 18205 -360
rect 18230 -415 18270 -410
rect 18230 -445 18235 -415
rect 18265 -445 18270 -415
rect 18230 -450 18270 -445
rect 18175 -485 18180 -465
rect 18200 -485 18205 -465
rect 18110 -505 18150 -500
rect 18110 -535 18115 -505
rect 18145 -535 18150 -505
rect 18110 -540 18150 -535
rect 18175 -590 18205 -485
rect 18235 -465 18265 -450
rect 18235 -485 18240 -465
rect 18260 -485 18265 -465
rect 18235 -545 18265 -485
rect 18295 -465 18325 -360
rect 18350 -370 18390 -365
rect 18350 -400 18355 -370
rect 18385 -400 18390 -370
rect 18350 -405 18390 -400
rect 18295 -485 18300 -465
rect 18320 -485 18325 -465
rect 18230 -550 18270 -545
rect 18230 -580 18235 -550
rect 18265 -580 18270 -550
rect 18230 -585 18270 -580
rect 18295 -590 18325 -485
rect 18355 -465 18385 -405
rect 18355 -485 18360 -465
rect 18380 -485 18385 -465
rect 18355 -500 18385 -485
rect 18415 -465 18445 -360
rect 18490 -410 18510 -255
rect 18530 -325 18570 -320
rect 18530 -355 18535 -325
rect 18565 -355 18570 -325
rect 18530 -360 18570 -355
rect 18470 -415 18510 -410
rect 18470 -445 18475 -415
rect 18505 -445 18510 -415
rect 18470 -450 18510 -445
rect 18415 -485 18420 -465
rect 18440 -485 18445 -465
rect 18350 -505 18390 -500
rect 18350 -535 18355 -505
rect 18385 -535 18390 -505
rect 18350 -540 18390 -535
rect 18415 -590 18445 -485
rect 18475 -465 18505 -450
rect 18475 -485 18480 -465
rect 18500 -485 18505 -465
rect 18475 -545 18505 -485
rect 18535 -465 18565 -360
rect 18600 -365 18620 -105
rect 18665 -160 18695 -35
rect 18725 35 18755 140
rect 18725 -35 18730 35
rect 18750 -35 18755 35
rect 18725 -110 18755 -35
rect 18785 35 18815 190
rect 18840 130 18880 135
rect 18840 100 18845 130
rect 18875 100 18880 130
rect 18840 95 18880 100
rect 18785 -35 18790 35
rect 18810 -35 18815 35
rect 18720 -115 18760 -110
rect 18720 -145 18725 -115
rect 18755 -145 18760 -115
rect 18720 -150 18760 -145
rect 18785 -160 18815 -35
rect 18845 35 18875 95
rect 18845 -35 18850 35
rect 18870 -35 18875 35
rect 18660 -165 18700 -160
rect 18660 -195 18665 -165
rect 18695 -195 18700 -165
rect 18660 -200 18700 -195
rect 18780 -165 18820 -160
rect 18780 -195 18785 -165
rect 18815 -195 18820 -165
rect 18780 -200 18820 -195
rect 18845 -215 18875 -35
rect 18905 35 18935 190
rect 18960 85 19000 90
rect 18960 55 18965 85
rect 18995 55 19000 85
rect 18960 50 19000 55
rect 18905 -35 18910 35
rect 18930 -35 18935 35
rect 18905 -160 18935 -35
rect 18965 35 18995 50
rect 18965 -35 18970 35
rect 18990 -35 18995 35
rect 18965 -65 18995 -35
rect 19025 35 19055 190
rect 19080 175 19120 180
rect 19080 145 19085 175
rect 19115 145 19120 175
rect 19080 140 19120 145
rect 19025 -35 19030 35
rect 19050 -35 19055 35
rect 18960 -70 19000 -65
rect 18960 -100 18965 -70
rect 18995 -100 19000 -70
rect 18960 -105 19000 -100
rect 19025 -160 19055 -35
rect 19085 35 19115 140
rect 19085 -35 19090 35
rect 19110 -35 19115 35
rect 19085 -110 19115 -35
rect 19145 100 19175 190
rect 19145 80 19150 100
rect 19170 80 19175 100
rect 19145 35 19175 80
rect 19145 -35 19150 35
rect 19170 -35 19175 35
rect 19080 -115 19120 -110
rect 19080 -145 19085 -115
rect 19115 -145 19120 -115
rect 19080 -150 19120 -145
rect 19145 -160 19175 -35
rect 18900 -165 18940 -160
rect 18900 -195 18905 -165
rect 18935 -195 18940 -165
rect 18900 -200 18940 -195
rect 19020 -165 19060 -160
rect 19020 -195 19025 -165
rect 19055 -195 19060 -165
rect 19020 -200 19060 -195
rect 19140 -165 19180 -160
rect 19140 -195 19145 -165
rect 19175 -195 19180 -165
rect 19140 -200 19180 -195
rect 18670 -220 18700 -215
rect 18670 -255 18700 -250
rect 18840 -220 18880 -215
rect 18840 -250 18845 -220
rect 18875 -250 18880 -220
rect 18840 -255 18880 -250
rect 19030 -220 19060 -215
rect 19030 -255 19060 -250
rect 18650 -325 18690 -320
rect 18650 -355 18655 -325
rect 18685 -355 18690 -325
rect 18650 -360 18690 -355
rect 18590 -370 18630 -365
rect 18590 -400 18595 -370
rect 18625 -400 18630 -370
rect 18590 -405 18630 -400
rect 18535 -485 18540 -465
rect 18560 -485 18565 -465
rect 18470 -550 18510 -545
rect 18470 -580 18475 -550
rect 18505 -580 18510 -550
rect 18470 -585 18510 -580
rect 18535 -590 18565 -485
rect 18595 -465 18625 -405
rect 18595 -485 18600 -465
rect 18620 -485 18625 -465
rect 18595 -500 18625 -485
rect 18655 -465 18685 -360
rect 18770 -390 18800 -385
rect 18710 -415 18750 -410
rect 18710 -445 18715 -415
rect 18745 -445 18750 -415
rect 18770 -425 18800 -420
rect 18710 -450 18750 -445
rect 18655 -485 18660 -465
rect 18680 -485 18685 -465
rect 18590 -505 18630 -500
rect 18590 -535 18595 -505
rect 18625 -535 18630 -505
rect 18590 -540 18630 -535
rect 18655 -590 18685 -485
rect 18715 -465 18745 -450
rect 18715 -485 18720 -465
rect 18740 -485 18745 -465
rect 18715 -545 18745 -485
rect 19335 -525 19355 1015
rect 19415 345 19435 1600
rect 19460 485 19500 490
rect 19460 455 19465 485
rect 19495 455 19500 485
rect 19460 450 19500 455
rect 19405 340 19445 345
rect 19405 310 19410 340
rect 19440 310 19445 340
rect 19405 305 19445 310
rect 19415 -385 19435 305
rect 19405 -390 19445 -385
rect 19405 -420 19410 -390
rect 19440 -420 19445 -390
rect 19405 -425 19445 -420
rect 18770 -530 18800 -525
rect 18710 -550 18750 -545
rect 18710 -580 18715 -550
rect 18745 -580 18750 -550
rect 18770 -565 18800 -560
rect 19325 -530 19365 -525
rect 19325 -560 19330 -530
rect 19360 -560 19365 -530
rect 19325 -565 19365 -560
rect 18710 -585 18750 -580
rect 18170 -595 18210 -590
rect 18170 -625 18175 -595
rect 18205 -625 18210 -595
rect 18170 -630 18210 -625
rect 18290 -595 18330 -590
rect 18290 -625 18295 -595
rect 18325 -625 18330 -595
rect 18290 -630 18330 -625
rect 18410 -595 18450 -590
rect 18410 -625 18415 -595
rect 18445 -625 18450 -595
rect 18410 -630 18450 -625
rect 18530 -595 18570 -590
rect 18530 -625 18535 -595
rect 18565 -625 18570 -595
rect 18530 -630 18570 -625
rect 18650 -595 18690 -590
rect 18650 -625 18655 -595
rect 18685 -625 18690 -595
rect 18650 -630 18690 -625
rect 19030 -595 19070 -590
rect 19030 -625 19035 -595
rect 19065 -625 19070 -595
rect 19030 -630 19070 -625
rect 18140 -680 18180 -675
rect 18140 -710 18145 -680
rect 18175 -710 18180 -680
rect 18140 -715 18180 -710
rect 18760 -680 18800 -675
rect 18760 -710 18765 -680
rect 18795 -710 18800 -680
rect 18760 -715 18800 -710
rect 17875 -740 17905 -730
rect 17875 -960 17880 -740
rect 17900 -960 17905 -740
rect 17875 -970 17905 -960
rect 18415 -740 18525 -730
rect 18415 -960 18420 -740
rect 18440 -960 18460 -740
rect 18480 -960 18500 -740
rect 18520 -960 18525 -740
rect 18415 -970 18525 -960
rect 19035 -740 19065 -630
rect 19035 -960 19040 -740
rect 19060 -960 19065 -740
rect 19035 -970 19065 -960
rect 18455 -990 18485 -970
rect 17110 -995 17150 -990
rect 17110 -1025 17115 -995
rect 17145 -1025 17150 -995
rect 17110 -1030 17150 -1025
rect 17780 -995 17820 -990
rect 17780 -1025 17785 -995
rect 17815 -1025 17820 -995
rect 17780 -1030 17820 -1025
rect 18450 -995 18490 -990
rect 18450 -1025 18455 -995
rect 18485 -1025 18490 -995
rect 18450 -1030 18490 -1025
rect 16740 -1095 16780 -1090
rect 16740 -1125 16745 -1095
rect 16775 -1125 16780 -1095
rect 16740 -1130 16780 -1125
rect 17260 -1095 17300 -1090
rect 17260 -1125 17265 -1095
rect 17295 -1125 17300 -1095
rect 17260 -1130 17300 -1125
rect 17780 -1095 17820 -1090
rect 17780 -1125 17785 -1095
rect 17815 -1125 17820 -1095
rect 17780 -1130 17820 -1125
rect 18300 -1095 18340 -1090
rect 18300 -1125 18305 -1095
rect 18335 -1125 18340 -1095
rect 18300 -1130 18340 -1125
rect 16745 -1160 16775 -1130
rect 16745 -1230 16750 -1160
rect 16770 -1230 16775 -1160
rect 16745 -1240 16775 -1230
rect 17785 -1160 17815 -1130
rect 17785 -1230 17790 -1160
rect 17810 -1230 17815 -1160
rect 17785 -1240 17815 -1230
rect 18825 -1160 18895 -1150
rect 18825 -1230 18830 -1160
rect 18850 -1230 18870 -1160
rect 18890 -1175 18895 -1160
rect 18890 -1180 18935 -1175
rect 18890 -1210 18900 -1180
rect 18930 -1210 18935 -1180
rect 18890 -1215 18935 -1210
rect 18890 -1230 18895 -1215
rect 18825 -1240 18895 -1230
rect 17285 -1335 17315 -1330
rect 16970 -1345 17010 -1340
rect 16970 -1375 16975 -1345
rect 17005 -1375 17010 -1345
rect 16970 -1380 17010 -1375
rect 17190 -1345 17230 -1340
rect 17190 -1375 17195 -1345
rect 17225 -1375 17230 -1345
rect 17285 -1370 17315 -1365
rect 17785 -1335 17815 -1330
rect 17785 -1370 17815 -1365
rect 18295 -1335 18325 -1330
rect 18295 -1370 18325 -1365
rect 18380 -1345 18420 -1340
rect 17190 -1380 17230 -1375
rect 18380 -1375 18385 -1345
rect 18415 -1375 18420 -1345
rect 18380 -1380 18420 -1375
rect 18600 -1345 18640 -1340
rect 18600 -1375 18605 -1345
rect 18635 -1375 18640 -1345
rect 18600 -1380 18640 -1375
rect 16915 -1435 16955 -1430
rect 16915 -1465 16920 -1435
rect 16950 -1465 16955 -1435
rect 16915 -1470 16955 -1465
rect 16920 -1500 16950 -1470
rect 16920 -1570 16925 -1500
rect 16945 -1570 16950 -1500
rect 16920 -1585 16950 -1570
rect 16975 -1500 17005 -1380
rect 17080 -1390 17120 -1385
rect 17080 -1420 17085 -1390
rect 17115 -1420 17120 -1390
rect 17080 -1425 17120 -1420
rect 17025 -1435 17065 -1430
rect 17025 -1465 17030 -1435
rect 17060 -1465 17065 -1435
rect 17025 -1470 17065 -1465
rect 16975 -1570 16980 -1500
rect 17000 -1570 17005 -1500
rect 16915 -1590 16955 -1585
rect 16915 -1620 16920 -1590
rect 16950 -1620 16955 -1590
rect 16915 -1625 16955 -1620
rect 16975 -1640 17005 -1570
rect 17030 -1500 17060 -1470
rect 17030 -1570 17035 -1500
rect 17055 -1570 17060 -1500
rect 17030 -1585 17060 -1570
rect 17085 -1500 17115 -1425
rect 17135 -1435 17175 -1430
rect 17135 -1465 17140 -1435
rect 17170 -1465 17175 -1435
rect 17135 -1470 17175 -1465
rect 17085 -1570 17090 -1500
rect 17110 -1570 17115 -1500
rect 17025 -1590 17065 -1585
rect 17025 -1620 17030 -1590
rect 17060 -1620 17065 -1590
rect 17025 -1625 17065 -1620
rect 16970 -1645 17010 -1640
rect 16970 -1675 16975 -1645
rect 17005 -1675 17010 -1645
rect 16970 -1680 17010 -1675
rect 17085 -1685 17115 -1570
rect 17140 -1500 17170 -1470
rect 17140 -1570 17145 -1500
rect 17165 -1570 17170 -1500
rect 17140 -1585 17170 -1570
rect 17195 -1500 17225 -1380
rect 17300 -1390 17340 -1385
rect 17300 -1420 17305 -1390
rect 17335 -1420 17340 -1390
rect 17300 -1425 17340 -1420
rect 17780 -1390 17820 -1385
rect 17780 -1420 17785 -1390
rect 17815 -1420 17820 -1390
rect 17780 -1425 17820 -1420
rect 17890 -1390 17930 -1385
rect 17890 -1420 17895 -1390
rect 17925 -1420 17930 -1390
rect 17890 -1425 17930 -1420
rect 18000 -1390 18040 -1385
rect 18000 -1420 18005 -1390
rect 18035 -1420 18040 -1390
rect 18000 -1425 18040 -1420
rect 18270 -1390 18310 -1385
rect 18270 -1420 18275 -1390
rect 18305 -1420 18310 -1390
rect 18270 -1425 18310 -1420
rect 17245 -1435 17285 -1430
rect 17245 -1465 17250 -1435
rect 17280 -1465 17285 -1435
rect 17245 -1470 17285 -1465
rect 17195 -1570 17200 -1500
rect 17220 -1570 17225 -1500
rect 17135 -1590 17175 -1585
rect 17135 -1620 17140 -1590
rect 17170 -1620 17175 -1590
rect 17135 -1625 17175 -1620
rect 17195 -1640 17225 -1570
rect 17250 -1500 17280 -1470
rect 17250 -1570 17255 -1500
rect 17275 -1570 17280 -1500
rect 17250 -1585 17280 -1570
rect 17305 -1500 17335 -1425
rect 17355 -1435 17395 -1430
rect 17355 -1465 17360 -1435
rect 17390 -1465 17395 -1435
rect 17355 -1470 17395 -1465
rect 17505 -1435 17545 -1430
rect 17505 -1465 17510 -1435
rect 17540 -1465 17545 -1435
rect 17505 -1470 17545 -1465
rect 17615 -1435 17655 -1430
rect 17615 -1465 17620 -1435
rect 17650 -1465 17655 -1435
rect 17615 -1470 17655 -1465
rect 17725 -1435 17765 -1430
rect 17725 -1465 17730 -1435
rect 17760 -1465 17765 -1435
rect 17725 -1470 17765 -1465
rect 17305 -1570 17310 -1500
rect 17330 -1570 17335 -1500
rect 17245 -1590 17285 -1585
rect 17245 -1620 17250 -1590
rect 17280 -1620 17285 -1590
rect 17245 -1625 17285 -1620
rect 17190 -1645 17230 -1640
rect 17190 -1675 17195 -1645
rect 17225 -1675 17230 -1645
rect 17190 -1680 17230 -1675
rect 17305 -1685 17335 -1570
rect 17360 -1500 17390 -1470
rect 17360 -1570 17365 -1500
rect 17385 -1570 17390 -1500
rect 17360 -1585 17390 -1570
rect 17510 -1500 17540 -1470
rect 17510 -1570 17515 -1500
rect 17535 -1570 17540 -1500
rect 17510 -1585 17540 -1570
rect 17565 -1500 17595 -1490
rect 17565 -1570 17570 -1500
rect 17590 -1570 17595 -1500
rect 17355 -1590 17395 -1585
rect 17355 -1620 17360 -1590
rect 17390 -1620 17395 -1590
rect 17355 -1625 17395 -1620
rect 17505 -1590 17545 -1585
rect 17505 -1620 17510 -1590
rect 17540 -1620 17545 -1590
rect 17505 -1625 17545 -1620
rect 17565 -1640 17595 -1570
rect 17620 -1500 17650 -1470
rect 17620 -1570 17625 -1500
rect 17645 -1570 17650 -1500
rect 17620 -1585 17650 -1570
rect 17675 -1500 17705 -1490
rect 17675 -1570 17680 -1500
rect 17700 -1570 17705 -1500
rect 17615 -1590 17655 -1585
rect 17615 -1620 17620 -1590
rect 17650 -1620 17655 -1590
rect 17615 -1625 17655 -1620
rect 17675 -1630 17705 -1570
rect 17730 -1500 17760 -1470
rect 17730 -1570 17735 -1500
rect 17755 -1570 17760 -1500
rect 17730 -1585 17760 -1570
rect 17785 -1500 17815 -1425
rect 17835 -1435 17875 -1430
rect 17835 -1465 17840 -1435
rect 17870 -1465 17875 -1435
rect 17835 -1470 17875 -1465
rect 17785 -1570 17790 -1500
rect 17810 -1570 17815 -1500
rect 17725 -1590 17765 -1585
rect 17725 -1620 17730 -1590
rect 17760 -1620 17765 -1590
rect 17725 -1625 17765 -1620
rect 17785 -1630 17815 -1570
rect 17840 -1500 17870 -1470
rect 17840 -1570 17845 -1500
rect 17865 -1570 17870 -1500
rect 17840 -1585 17870 -1570
rect 17895 -1500 17925 -1425
rect 17945 -1435 17985 -1430
rect 17945 -1465 17950 -1435
rect 17980 -1465 17985 -1435
rect 17945 -1470 17985 -1465
rect 17895 -1570 17900 -1500
rect 17920 -1570 17925 -1500
rect 17835 -1590 17875 -1585
rect 17835 -1620 17840 -1590
rect 17870 -1620 17875 -1590
rect 17835 -1625 17875 -1620
rect 17895 -1630 17925 -1570
rect 17950 -1500 17980 -1470
rect 17950 -1570 17955 -1500
rect 17975 -1570 17980 -1500
rect 17950 -1585 17980 -1570
rect 18005 -1500 18035 -1425
rect 18055 -1435 18095 -1430
rect 18055 -1465 18060 -1435
rect 18090 -1465 18095 -1435
rect 18055 -1470 18095 -1465
rect 18215 -1435 18255 -1430
rect 18215 -1465 18220 -1435
rect 18250 -1465 18255 -1435
rect 18215 -1470 18255 -1465
rect 18005 -1570 18010 -1500
rect 18030 -1570 18035 -1500
rect 17945 -1590 17985 -1585
rect 17945 -1620 17950 -1590
rect 17980 -1620 17985 -1590
rect 17945 -1625 17985 -1620
rect 18005 -1630 18035 -1570
rect 18060 -1500 18090 -1470
rect 18060 -1570 18065 -1500
rect 18085 -1570 18090 -1500
rect 18060 -1585 18090 -1570
rect 18220 -1500 18250 -1470
rect 18220 -1570 18225 -1500
rect 18245 -1570 18250 -1500
rect 18220 -1585 18250 -1570
rect 18275 -1500 18305 -1425
rect 18325 -1435 18365 -1430
rect 18325 -1465 18330 -1435
rect 18360 -1465 18365 -1435
rect 18325 -1470 18365 -1465
rect 18275 -1570 18280 -1500
rect 18300 -1570 18305 -1500
rect 18055 -1590 18095 -1585
rect 18055 -1620 18060 -1590
rect 18090 -1620 18095 -1590
rect 18055 -1625 18095 -1620
rect 18215 -1590 18255 -1585
rect 18215 -1620 18220 -1590
rect 18250 -1620 18255 -1590
rect 18215 -1625 18255 -1620
rect 17670 -1635 17710 -1630
rect 17565 -1645 17615 -1640
rect 17565 -1675 17585 -1645
rect 17670 -1665 17675 -1635
rect 17705 -1665 17710 -1635
rect 17670 -1670 17710 -1665
rect 17780 -1635 17820 -1630
rect 17780 -1665 17785 -1635
rect 17815 -1665 17820 -1635
rect 17780 -1670 17820 -1665
rect 17890 -1635 17930 -1630
rect 17890 -1665 17895 -1635
rect 17925 -1665 17930 -1635
rect 17890 -1670 17930 -1665
rect 18000 -1635 18040 -1630
rect 18000 -1665 18005 -1635
rect 18035 -1665 18040 -1635
rect 18000 -1670 18040 -1665
rect 17565 -1680 17615 -1675
rect 17080 -1690 17120 -1685
rect 17080 -1720 17085 -1690
rect 17115 -1720 17120 -1690
rect 17080 -1725 17120 -1720
rect 17300 -1690 17340 -1685
rect 17300 -1720 17305 -1690
rect 17335 -1720 17340 -1690
rect 17300 -1725 17340 -1720
rect 17590 -1775 17610 -1680
rect 17580 -1780 17620 -1775
rect 17580 -1810 17585 -1780
rect 17615 -1810 17620 -1780
rect 17580 -1815 17620 -1810
rect 17680 -1820 17700 -1670
rect 17900 -1770 17920 -1670
rect 18275 -1685 18305 -1570
rect 18330 -1500 18360 -1470
rect 18330 -1570 18335 -1500
rect 18355 -1570 18360 -1500
rect 18330 -1585 18360 -1570
rect 18385 -1500 18415 -1380
rect 18490 -1390 18530 -1385
rect 18490 -1420 18495 -1390
rect 18525 -1420 18530 -1390
rect 18490 -1425 18530 -1420
rect 18435 -1435 18475 -1430
rect 18435 -1465 18440 -1435
rect 18470 -1465 18475 -1435
rect 18435 -1470 18475 -1465
rect 18385 -1570 18390 -1500
rect 18410 -1570 18415 -1500
rect 18325 -1590 18365 -1585
rect 18325 -1620 18330 -1590
rect 18360 -1620 18365 -1590
rect 18325 -1625 18365 -1620
rect 18385 -1640 18415 -1570
rect 18440 -1500 18470 -1470
rect 18440 -1570 18445 -1500
rect 18465 -1570 18470 -1500
rect 18440 -1585 18470 -1570
rect 18495 -1500 18525 -1425
rect 18545 -1435 18585 -1430
rect 18545 -1465 18550 -1435
rect 18580 -1465 18585 -1435
rect 18545 -1470 18585 -1465
rect 18495 -1570 18500 -1500
rect 18520 -1570 18525 -1500
rect 18435 -1590 18475 -1585
rect 18435 -1620 18440 -1590
rect 18470 -1620 18475 -1590
rect 18435 -1625 18475 -1620
rect 18380 -1645 18420 -1640
rect 18380 -1675 18385 -1645
rect 18415 -1675 18420 -1645
rect 18380 -1680 18420 -1675
rect 18495 -1685 18525 -1570
rect 18550 -1500 18580 -1470
rect 18550 -1570 18555 -1500
rect 18575 -1570 18580 -1500
rect 18550 -1585 18580 -1570
rect 18605 -1500 18635 -1380
rect 18655 -1435 18695 -1430
rect 18655 -1465 18660 -1435
rect 18690 -1465 18695 -1435
rect 18655 -1470 18695 -1465
rect 18605 -1570 18610 -1500
rect 18630 -1570 18635 -1500
rect 18545 -1590 18585 -1585
rect 18545 -1620 18550 -1590
rect 18580 -1620 18585 -1590
rect 18545 -1625 18585 -1620
rect 18605 -1640 18635 -1570
rect 18660 -1500 18690 -1470
rect 18660 -1570 18665 -1500
rect 18685 -1570 18690 -1500
rect 18660 -1585 18690 -1570
rect 18655 -1590 18695 -1585
rect 18655 -1620 18660 -1590
rect 18690 -1620 18695 -1590
rect 18655 -1625 18695 -1620
rect 18600 -1645 18640 -1640
rect 18600 -1675 18605 -1645
rect 18635 -1675 18640 -1645
rect 18600 -1680 18640 -1675
rect 18270 -1690 18310 -1685
rect 18270 -1720 18275 -1690
rect 18305 -1720 18310 -1690
rect 18270 -1725 18310 -1720
rect 18490 -1690 18530 -1685
rect 18490 -1720 18495 -1690
rect 18525 -1720 18530 -1690
rect 18490 -1725 18530 -1720
rect 17890 -1775 17930 -1770
rect 17890 -1805 17895 -1775
rect 17925 -1805 17930 -1775
rect 17890 -1810 17930 -1805
rect 17670 -1825 17710 -1820
rect 17670 -1855 17675 -1825
rect 17705 -1855 17710 -1825
rect 17670 -1860 17710 -1855
rect 19335 -1895 19355 -565
rect 19325 -1900 19365 -1895
rect 19325 -1930 19330 -1900
rect 19360 -1930 19365 -1900
rect 19325 -1935 19365 -1930
rect 16260 -1945 16300 -1940
rect 16260 -1975 16265 -1945
rect 16295 -1975 16300 -1945
rect 16260 -1980 16300 -1975
rect 16480 -1945 16520 -1940
rect 16480 -1975 16485 -1945
rect 16515 -1975 16520 -1945
rect 16480 -1980 16520 -1975
rect 16730 -1945 16770 -1940
rect 16730 -1975 16735 -1945
rect 16765 -1975 16770 -1945
rect 16730 -1980 16770 -1975
rect 17195 -1945 17235 -1940
rect 17195 -1975 17200 -1945
rect 17230 -1975 17235 -1945
rect 17195 -1980 17235 -1975
rect 17425 -1980 17430 -1945
rect 17465 -1980 17470 -1945
rect 18124 -1980 18129 -1945
rect 18164 -1980 18169 -1945
rect 19080 -1950 19120 -1945
rect 19080 -1980 19085 -1950
rect 19115 -1980 19120 -1950
rect 16490 -2895 16510 -1980
rect 16485 -2900 16520 -2895
rect 16485 -2940 16520 -2935
rect 16160 -3025 16195 -3020
rect 16160 -3065 16195 -3060
rect 16740 -3100 16760 -1980
rect 17205 -2010 17225 -1980
rect 19080 -1985 19120 -1980
rect 17195 -2015 17235 -2010
rect 17195 -2045 17200 -2015
rect 17230 -2045 17235 -2015
rect 17195 -2050 17235 -2045
rect 18830 -2015 18870 -2010
rect 18830 -2045 18835 -2015
rect 18865 -2045 18870 -2015
rect 18830 -2050 18870 -2045
rect 16945 -2615 18655 -2265
rect 16730 -3105 16770 -3100
rect 15820 -3145 15825 -3115
rect 15855 -3145 15860 -3115
rect 15820 -3150 15860 -3145
rect 15950 -3116 15985 -3111
rect 16730 -3135 16735 -3105
rect 16765 -3135 16770 -3105
rect 16730 -3140 16770 -3135
rect 15830 -4260 15850 -3150
rect 15950 -3156 15985 -3151
rect 16945 -3625 17295 -2615
rect 17625 -3105 17975 -2945
rect 17625 -3135 17785 -3105
rect 17815 -3135 17975 -3105
rect 17625 -3295 17975 -3135
rect 18305 -3105 18655 -2615
rect 18840 -3100 18860 -2050
rect 19090 -2895 19110 -1985
rect 19080 -2900 19115 -2895
rect 19080 -2940 19115 -2935
rect 19415 -2987 19435 -425
rect 19470 -1945 19490 450
rect 19545 -1770 19565 1600
rect 19610 280 19650 285
rect 19610 250 19615 280
rect 19645 250 19650 280
rect 19610 245 19650 250
rect 19535 -1775 19575 -1770
rect 19535 -1805 19540 -1775
rect 19570 -1805 19575 -1775
rect 19535 -1810 19575 -1805
rect 19460 -1950 19500 -1945
rect 19460 -1980 19465 -1950
rect 19495 -1980 19500 -1950
rect 19460 -1985 19500 -1980
rect 19405 -2992 19440 -2987
rect 19405 -3032 19440 -3027
rect 18305 -3135 18620 -3105
rect 18650 -3135 18655 -3105
rect 18305 -3625 18655 -3135
rect 18830 -3105 18870 -3100
rect 18830 -3135 18835 -3105
rect 18865 -3135 18870 -3105
rect 19620 -3111 19640 245
rect 19730 -220 19770 -215
rect 19730 -250 19735 -220
rect 19765 -250 19770 -220
rect 19730 -255 19770 -250
rect 18830 -3140 18870 -3135
rect 19610 -3116 19645 -3111
rect 19610 -3156 19645 -3151
rect 15950 -3789 15985 -3784
rect 15950 -3829 15985 -3824
rect 15820 -4265 15860 -4260
rect 15820 -4295 15825 -4265
rect 15855 -4295 15860 -4265
rect 15820 -4300 15860 -4295
rect 15725 -4315 15765 -4310
rect 15725 -4345 15730 -4315
rect 15760 -4345 15765 -4315
rect 15725 -4350 15765 -4345
rect 15960 -4355 15980 -3829
rect 16280 -3894 16315 -3889
rect 16280 -3934 16315 -3929
rect 16290 -4185 16310 -3934
rect 16605 -3969 16640 -3964
rect 16945 -3975 18655 -3625
rect 19610 -3789 19645 -3784
rect 19610 -3829 19645 -3824
rect 19285 -3894 19320 -3889
rect 19285 -3934 19320 -3929
rect 18960 -3969 18995 -3964
rect 16605 -4009 16640 -4004
rect 18960 -4009 18995 -4004
rect 16540 -4035 16580 -4030
rect 16540 -4065 16545 -4035
rect 16575 -4065 16580 -4035
rect 16540 -4070 16580 -4065
rect 16550 -4185 16570 -4070
rect 16615 -4185 16635 -4009
rect 16280 -4190 16320 -4185
rect 16280 -4220 16285 -4190
rect 16315 -4220 16320 -4190
rect 16280 -4225 16320 -4220
rect 16540 -4190 16580 -4185
rect 16540 -4220 16545 -4190
rect 16575 -4220 16580 -4190
rect 16540 -4225 16580 -4220
rect 16605 -4190 16645 -4185
rect 16605 -4220 16610 -4190
rect 16640 -4220 16645 -4190
rect 16605 -4225 16645 -4220
rect 17250 -4265 17300 -4255
rect 18965 -4260 18985 -4009
rect 19290 -4260 19310 -3934
rect 17250 -4295 17260 -4265
rect 17290 -4295 17300 -4265
rect 17250 -4305 17300 -4295
rect 17780 -4265 17820 -4260
rect 17780 -4295 17785 -4265
rect 17815 -4295 17820 -4265
rect 17780 -4300 17820 -4295
rect 18955 -4265 18995 -4260
rect 18955 -4295 18960 -4265
rect 18990 -4295 18995 -4265
rect 18955 -4300 18995 -4295
rect 19280 -4265 19320 -4260
rect 19280 -4295 19285 -4265
rect 19315 -4295 19320 -4265
rect 19280 -4300 19320 -4295
rect 16900 -4315 16950 -4305
rect 16900 -4345 16910 -4315
rect 16940 -4345 16950 -4315
rect 16900 -4355 16950 -4345
rect 18650 -4315 18700 -4305
rect 18650 -4345 18660 -4315
rect 18690 -4345 18700 -4315
rect 18650 -4355 18700 -4345
rect 19620 -4355 19640 -3829
rect 19740 -4310 19760 -255
rect 19785 -1340 19805 1595
rect 19775 -1345 19815 -1340
rect 19775 -1375 19780 -1345
rect 19810 -1375 19815 -1345
rect 19775 -1380 19815 -1375
rect 19730 -4315 19770 -4310
rect 19730 -4345 19735 -4315
rect 19765 -4345 19770 -4315
rect 19730 -4350 19770 -4345
rect 15950 -4360 15990 -4355
rect 15950 -4390 15955 -4360
rect 15985 -4390 15990 -4360
rect 15950 -4395 15990 -4390
rect 16205 -4360 16245 -4355
rect 16205 -4390 16210 -4360
rect 16240 -4390 16245 -4360
rect 16205 -4395 16245 -4390
rect 19355 -4360 19395 -4355
rect 19355 -4390 19360 -4360
rect 19390 -4390 19395 -4360
rect 19355 -4395 19395 -4390
rect 19610 -4360 19650 -4355
rect 19610 -4390 19615 -4360
rect 19645 -4390 19650 -4360
rect 19610 -4395 19650 -4390
rect 17955 -4410 17995 -4405
rect 17955 -4440 17960 -4410
rect 17990 -4440 17995 -4410
rect 17955 -4445 17995 -4440
<< via1 >>
rect 15730 -245 15760 -215
rect 15955 145 15985 175
rect 15790 -1375 15820 -1345
rect 16035 -1720 16065 -1690
rect 16870 1365 16900 1395
rect 16980 1365 17010 1395
rect 17090 1365 17120 1395
rect 17620 1365 17650 1395
rect 17730 1365 17760 1395
rect 17840 1365 17870 1395
rect 17950 1365 17980 1395
rect 18480 1365 18510 1395
rect 18590 1365 18620 1395
rect 18700 1365 18730 1395
rect 16815 1345 16845 1350
rect 16815 1325 16820 1345
rect 16820 1325 16840 1345
rect 16840 1325 16845 1345
rect 16815 1320 16845 1325
rect 16925 1320 16955 1350
rect 16870 1165 16900 1195
rect 17035 1320 17065 1350
rect 16980 1165 17010 1195
rect 17145 1345 17175 1350
rect 17145 1325 17150 1345
rect 17150 1325 17170 1345
rect 17170 1325 17175 1345
rect 17145 1320 17175 1325
rect 17455 1345 17485 1350
rect 17455 1325 17460 1345
rect 17460 1325 17480 1345
rect 17480 1325 17485 1345
rect 17455 1320 17485 1325
rect 17565 1320 17595 1350
rect 17090 1165 17120 1195
rect 16815 1120 16845 1150
rect 16925 1120 16955 1150
rect 17035 1120 17065 1150
rect 17145 1120 17175 1150
rect 17455 1120 17485 1150
rect 17070 1090 17100 1095
rect 17070 1070 17075 1090
rect 17075 1070 17095 1090
rect 17095 1070 17100 1090
rect 17070 1065 17100 1070
rect 17675 1320 17705 1350
rect 17620 1165 17650 1195
rect 17785 1320 17815 1350
rect 17730 1165 17760 1195
rect 17895 1320 17925 1350
rect 17840 1165 17870 1195
rect 18005 1320 18035 1350
rect 18115 1345 18145 1350
rect 18115 1325 18120 1345
rect 18120 1325 18140 1345
rect 18140 1325 18145 1345
rect 18115 1320 18145 1325
rect 18425 1345 18455 1350
rect 18425 1325 18430 1345
rect 18430 1325 18450 1345
rect 18450 1325 18455 1345
rect 18425 1320 18455 1325
rect 17950 1165 17980 1195
rect 17565 1120 17595 1150
rect 17675 1120 17705 1150
rect 17785 1120 17815 1150
rect 17895 1120 17925 1150
rect 18005 1120 18035 1150
rect 17805 1090 17835 1095
rect 17805 1070 17810 1090
rect 17810 1070 17830 1090
rect 17830 1070 17835 1090
rect 17805 1065 17835 1070
rect 18535 1320 18565 1350
rect 18480 1165 18510 1195
rect 18645 1320 18675 1350
rect 18590 1165 18620 1195
rect 18755 1345 18785 1350
rect 18755 1325 18760 1345
rect 18760 1325 18780 1345
rect 18780 1325 18785 1345
rect 18755 1320 18785 1325
rect 18700 1165 18730 1195
rect 18115 1120 18145 1150
rect 18425 1120 18455 1150
rect 18535 1120 18565 1150
rect 18645 1120 18675 1150
rect 18755 1120 18785 1150
rect 18500 1090 18530 1095
rect 18500 1070 18505 1090
rect 18505 1070 18525 1090
rect 18525 1070 18530 1090
rect 18500 1065 18530 1070
rect 18725 1065 18755 1095
rect 16165 1020 16195 1050
rect 17510 1020 17540 1050
rect 17605 990 17635 1020
rect 17965 990 17995 1020
rect 18060 1020 18090 1050
rect 17425 945 17455 975
rect 17245 900 17275 930
rect 17065 855 17095 885
rect 16440 810 16470 840
rect 16660 810 16690 840
rect 16975 835 17005 840
rect 16975 815 16980 835
rect 16980 815 17000 835
rect 17000 815 17005 835
rect 16975 810 17005 815
rect 16440 775 16470 780
rect 16440 755 16445 775
rect 16445 755 16465 775
rect 16465 755 16470 775
rect 16440 750 16470 755
rect 16495 750 16525 780
rect 16605 750 16635 780
rect 16660 775 16690 780
rect 16660 755 16665 775
rect 16665 755 16685 775
rect 16685 755 16690 775
rect 16660 750 16690 755
rect 16550 705 16580 735
rect 16785 705 16815 735
rect 16495 565 16525 595
rect 16440 520 16470 550
rect 16605 565 16635 595
rect 16310 455 16340 485
rect 16265 400 16295 430
rect 16210 355 16240 385
rect 16265 -420 16295 -390
rect 16210 -1125 16240 -1095
rect 16165 -1810 16195 -1780
rect 16110 -1855 16140 -1825
rect 16160 -1930 16190 -1900
rect 16660 520 16690 550
rect 16845 565 16875 595
rect 16785 400 16815 430
rect 16550 355 16580 385
rect 16425 195 16455 225
rect 16545 195 16575 225
rect 16665 195 16695 225
rect 16785 195 16815 225
rect 16485 145 16515 175
rect 16605 55 16635 85
rect 16485 -145 16515 -115
rect 16725 100 16755 130
rect 16605 -75 16635 -70
rect 16605 -95 16610 -75
rect 16610 -95 16630 -75
rect 16630 -95 16635 -75
rect 16605 -100 16635 -95
rect 16425 -195 16455 -165
rect 16545 -195 16575 -165
rect 16665 -195 16695 -165
rect 17155 810 17185 840
rect 17335 810 17365 840
rect 17515 810 17545 840
rect 17785 855 17815 885
rect 17695 810 17725 840
rect 17875 810 17905 840
rect 17605 455 17635 485
rect 17425 400 17455 430
rect 17245 355 17275 385
rect 17065 310 17095 340
rect 16905 195 16935 225
rect 17025 195 17055 225
rect 17145 195 17175 225
rect 17265 195 17295 225
rect 17385 195 17415 225
rect 17505 195 17535 225
rect 17625 195 17655 225
rect 16845 145 16875 175
rect 16965 55 16995 85
rect 16845 -145 16875 -115
rect 17085 100 17115 130
rect 16965 -75 16995 -70
rect 16965 -95 16970 -75
rect 16970 -95 16990 -75
rect 16990 -95 16995 -75
rect 16965 -100 16995 -95
rect 16785 -195 16815 -165
rect 16905 -195 16935 -165
rect 16540 -225 16570 -220
rect 16540 -245 16545 -225
rect 16545 -245 16565 -225
rect 16565 -245 16570 -225
rect 16540 -250 16570 -245
rect 16725 -250 16755 -220
rect 16900 -225 16930 -220
rect 16900 -245 16905 -225
rect 16905 -245 16925 -225
rect 16925 -245 16930 -225
rect 16900 -250 16930 -245
rect 16915 -355 16945 -325
rect 16800 -395 16830 -390
rect 16800 -415 16805 -395
rect 16805 -415 16825 -395
rect 16825 -415 16830 -395
rect 16800 -420 16830 -415
rect 16855 -445 16885 -415
rect 16310 -560 16340 -530
rect 16800 -535 16830 -530
rect 16800 -555 16805 -535
rect 16805 -555 16825 -535
rect 16825 -555 16830 -535
rect 17025 -195 17055 -165
rect 17205 145 17235 175
rect 17325 55 17355 85
rect 17205 -145 17235 -115
rect 17445 100 17475 130
rect 17325 -75 17355 -70
rect 17325 -95 17330 -75
rect 17330 -95 17350 -75
rect 17350 -95 17355 -75
rect 17325 -100 17355 -95
rect 17145 -195 17175 -165
rect 17265 -195 17295 -165
rect 17385 -195 17415 -165
rect 17565 145 17595 175
rect 18145 945 18175 975
rect 18055 810 18085 840
rect 18325 900 18355 930
rect 18235 810 18265 840
rect 17965 455 17995 485
rect 18505 855 18535 885
rect 18415 810 18445 840
rect 18145 400 18175 430
rect 18595 835 18625 840
rect 18595 815 18600 835
rect 18600 815 18620 835
rect 18620 815 18625 835
rect 18595 810 18625 815
rect 18325 355 18355 385
rect 17785 310 17815 340
rect 18505 310 18535 340
rect 19015 810 19045 840
rect 18905 775 18935 780
rect 18905 755 18910 775
rect 18910 755 18930 775
rect 18930 755 18935 775
rect 18905 750 18935 755
rect 19015 750 19045 780
rect 19125 775 19155 780
rect 19125 755 19130 775
rect 19130 755 19150 775
rect 19150 755 19155 775
rect 19125 750 19155 755
rect 18960 705 18990 735
rect 18905 565 18935 595
rect 19070 705 19100 735
rect 19015 565 19045 595
rect 19125 565 19155 595
rect 19330 1020 19360 1050
rect 18960 520 18990 550
rect 19070 520 19100 550
rect 19265 520 19295 550
rect 18725 250 18755 280
rect 19015 250 19045 280
rect 17945 195 17975 225
rect 18065 195 18095 225
rect 18185 195 18215 225
rect 18305 195 18335 225
rect 18425 195 18455 225
rect 18545 195 18575 225
rect 18665 195 18695 225
rect 17695 145 17725 175
rect 17875 145 17905 175
rect 17565 -145 17595 -115
rect 17505 -195 17535 -165
rect 17625 -195 17655 -165
rect 17085 -250 17115 -220
rect 17260 -225 17290 -220
rect 17260 -245 17265 -225
rect 17265 -245 17285 -225
rect 17285 -245 17290 -225
rect 17260 -250 17290 -245
rect 17445 -250 17475 -220
rect 17510 -225 17540 -220
rect 17510 -245 17515 -225
rect 17515 -245 17535 -225
rect 17535 -245 17540 -225
rect 17510 -250 17540 -245
rect 17035 -355 17065 -325
rect 16975 -400 17005 -370
rect 16800 -560 16830 -555
rect 16855 -580 16885 -550
rect 17155 -355 17185 -325
rect 17275 -355 17305 -325
rect 17395 -355 17425 -325
rect 17095 -445 17125 -415
rect 16975 -535 17005 -505
rect 17215 -400 17245 -370
rect 17095 -580 17125 -550
rect 17335 -445 17365 -415
rect 17215 -535 17245 -505
rect 17455 -400 17485 -370
rect 17335 -580 17365 -550
rect 17565 -465 17595 -460
rect 17565 -485 17570 -465
rect 17570 -485 17590 -465
rect 17590 -485 17595 -465
rect 17565 -490 17595 -485
rect 17455 -535 17485 -505
rect 16535 -625 16565 -595
rect 16915 -625 16945 -595
rect 17035 -625 17065 -595
rect 17155 -625 17185 -595
rect 17275 -625 17305 -595
rect 17395 -625 17425 -595
rect 16805 -685 16835 -680
rect 16805 -705 16810 -685
rect 16810 -705 16830 -685
rect 16830 -705 16835 -685
rect 16805 -710 16835 -705
rect 17425 -685 17455 -680
rect 17425 -705 17430 -685
rect 17430 -705 17450 -685
rect 17450 -705 17455 -685
rect 17425 -710 17455 -705
rect 17785 -490 17815 -460
rect 18005 145 18035 175
rect 18125 100 18155 130
rect 18005 -145 18035 -115
rect 17945 -195 17975 -165
rect 18065 -195 18095 -165
rect 18245 55 18275 85
rect 18365 145 18395 175
rect 18245 -75 18275 -70
rect 18245 -95 18250 -75
rect 18250 -95 18270 -75
rect 18270 -95 18275 -75
rect 18245 -100 18275 -95
rect 18485 100 18515 130
rect 18365 -145 18395 -115
rect 18185 -195 18215 -165
rect 18305 -195 18335 -165
rect 18425 -195 18455 -165
rect 18605 55 18635 85
rect 18785 195 18815 225
rect 18905 195 18935 225
rect 19025 195 19055 225
rect 19145 195 19175 225
rect 18725 145 18755 175
rect 18605 -75 18635 -70
rect 18605 -95 18610 -75
rect 18610 -95 18630 -75
rect 18630 -95 18635 -75
rect 18605 -100 18635 -95
rect 18545 -195 18575 -165
rect 18060 -225 18090 -220
rect 18060 -245 18065 -225
rect 18065 -245 18085 -225
rect 18085 -245 18090 -225
rect 18060 -250 18090 -245
rect 18125 -250 18155 -220
rect 18310 -225 18340 -220
rect 18310 -245 18315 -225
rect 18315 -245 18335 -225
rect 18335 -245 18340 -225
rect 18310 -250 18340 -245
rect 18485 -250 18515 -220
rect 18175 -355 18205 -325
rect 18295 -355 18325 -325
rect 18415 -355 18445 -325
rect 18115 -400 18145 -370
rect 18005 -465 18035 -460
rect 18005 -485 18010 -465
rect 18010 -485 18030 -465
rect 18030 -485 18035 -465
rect 18005 -490 18035 -485
rect 18235 -445 18265 -415
rect 18115 -535 18145 -505
rect 18355 -400 18385 -370
rect 18235 -580 18265 -550
rect 18535 -355 18565 -325
rect 18475 -445 18505 -415
rect 18355 -535 18385 -505
rect 18845 100 18875 130
rect 18725 -145 18755 -115
rect 18665 -195 18695 -165
rect 18785 -195 18815 -165
rect 18965 55 18995 85
rect 19085 145 19115 175
rect 18965 -75 18995 -70
rect 18965 -95 18970 -75
rect 18970 -95 18990 -75
rect 18990 -95 18995 -75
rect 18965 -100 18995 -95
rect 19085 -145 19115 -115
rect 18905 -195 18935 -165
rect 19025 -195 19055 -165
rect 19145 -195 19175 -165
rect 18670 -225 18700 -220
rect 18670 -245 18675 -225
rect 18675 -245 18695 -225
rect 18695 -245 18700 -225
rect 18670 -250 18700 -245
rect 18845 -250 18875 -220
rect 19030 -225 19060 -220
rect 19030 -245 19035 -225
rect 19035 -245 19055 -225
rect 19055 -245 19060 -225
rect 19030 -250 19060 -245
rect 18655 -355 18685 -325
rect 18595 -400 18625 -370
rect 18475 -580 18505 -550
rect 18770 -395 18800 -390
rect 18715 -445 18745 -415
rect 18770 -415 18775 -395
rect 18775 -415 18795 -395
rect 18795 -415 18800 -395
rect 18770 -420 18800 -415
rect 18595 -535 18625 -505
rect 19465 455 19495 485
rect 19410 310 19440 340
rect 19410 -420 19440 -390
rect 18770 -535 18800 -530
rect 18715 -580 18745 -550
rect 18770 -555 18775 -535
rect 18775 -555 18795 -535
rect 18795 -555 18800 -535
rect 18770 -560 18800 -555
rect 19330 -560 19360 -530
rect 18175 -625 18205 -595
rect 18295 -625 18325 -595
rect 18415 -625 18445 -595
rect 18535 -625 18565 -595
rect 18655 -625 18685 -595
rect 19035 -625 19065 -595
rect 18145 -685 18175 -680
rect 18145 -705 18150 -685
rect 18150 -705 18170 -685
rect 18170 -705 18175 -685
rect 18145 -710 18175 -705
rect 18765 -685 18795 -680
rect 18765 -705 18770 -685
rect 18770 -705 18790 -685
rect 18790 -705 18795 -685
rect 18765 -710 18795 -705
rect 17115 -1025 17145 -995
rect 17785 -1025 17815 -995
rect 18455 -1025 18485 -995
rect 16745 -1125 16775 -1095
rect 17265 -1100 17295 -1095
rect 17265 -1120 17270 -1100
rect 17270 -1120 17290 -1100
rect 17290 -1120 17295 -1100
rect 17265 -1125 17295 -1120
rect 17785 -1125 17815 -1095
rect 18305 -1100 18335 -1095
rect 18305 -1120 18310 -1100
rect 18310 -1120 18330 -1100
rect 18330 -1120 18335 -1100
rect 18305 -1125 18335 -1120
rect 18900 -1210 18930 -1180
rect 17285 -1340 17315 -1335
rect 16975 -1375 17005 -1345
rect 17195 -1375 17225 -1345
rect 17285 -1360 17290 -1340
rect 17290 -1360 17310 -1340
rect 17310 -1360 17315 -1340
rect 17285 -1365 17315 -1360
rect 17785 -1340 17815 -1335
rect 17785 -1360 17790 -1340
rect 17790 -1360 17810 -1340
rect 17810 -1360 17815 -1340
rect 17785 -1365 17815 -1360
rect 18295 -1340 18325 -1335
rect 18295 -1360 18300 -1340
rect 18300 -1360 18320 -1340
rect 18320 -1360 18325 -1340
rect 18295 -1365 18325 -1360
rect 18385 -1375 18415 -1345
rect 18605 -1375 18635 -1345
rect 16920 -1440 16950 -1435
rect 16920 -1460 16925 -1440
rect 16925 -1460 16945 -1440
rect 16945 -1460 16950 -1440
rect 16920 -1465 16950 -1460
rect 17085 -1420 17115 -1390
rect 17030 -1465 17060 -1435
rect 16920 -1620 16950 -1590
rect 17140 -1465 17170 -1435
rect 17030 -1620 17060 -1590
rect 16975 -1675 17005 -1645
rect 17305 -1420 17335 -1390
rect 17785 -1420 17815 -1390
rect 17895 -1420 17925 -1390
rect 18005 -1420 18035 -1390
rect 18275 -1420 18305 -1390
rect 17250 -1465 17280 -1435
rect 17140 -1620 17170 -1590
rect 17360 -1440 17390 -1435
rect 17360 -1460 17365 -1440
rect 17365 -1460 17385 -1440
rect 17385 -1460 17390 -1440
rect 17360 -1465 17390 -1460
rect 17510 -1440 17540 -1435
rect 17510 -1460 17515 -1440
rect 17515 -1460 17535 -1440
rect 17535 -1460 17540 -1440
rect 17510 -1465 17540 -1460
rect 17620 -1465 17650 -1435
rect 17730 -1465 17760 -1435
rect 17250 -1620 17280 -1590
rect 17195 -1675 17225 -1645
rect 17360 -1620 17390 -1590
rect 17510 -1620 17540 -1590
rect 17620 -1620 17650 -1590
rect 17840 -1465 17870 -1435
rect 17730 -1620 17760 -1590
rect 17950 -1465 17980 -1435
rect 17840 -1620 17870 -1590
rect 18060 -1440 18090 -1435
rect 18060 -1460 18065 -1440
rect 18065 -1460 18085 -1440
rect 18085 -1460 18090 -1440
rect 18060 -1465 18090 -1460
rect 18220 -1440 18250 -1435
rect 18220 -1460 18225 -1440
rect 18225 -1460 18245 -1440
rect 18245 -1460 18250 -1440
rect 18220 -1465 18250 -1460
rect 17950 -1620 17980 -1590
rect 18330 -1465 18360 -1435
rect 18060 -1620 18090 -1590
rect 18220 -1620 18250 -1590
rect 17585 -1650 17615 -1645
rect 17585 -1670 17590 -1650
rect 17590 -1670 17610 -1650
rect 17610 -1670 17615 -1650
rect 17675 -1665 17705 -1635
rect 17785 -1665 17815 -1635
rect 17895 -1665 17925 -1635
rect 18005 -1665 18035 -1635
rect 17585 -1675 17615 -1670
rect 17085 -1720 17115 -1690
rect 17305 -1720 17335 -1690
rect 17585 -1810 17615 -1780
rect 18495 -1420 18525 -1390
rect 18440 -1465 18470 -1435
rect 18330 -1620 18360 -1590
rect 18550 -1465 18580 -1435
rect 18440 -1620 18470 -1590
rect 18385 -1675 18415 -1645
rect 18660 -1440 18690 -1435
rect 18660 -1460 18665 -1440
rect 18665 -1460 18685 -1440
rect 18685 -1460 18690 -1440
rect 18660 -1465 18690 -1460
rect 18550 -1620 18580 -1590
rect 18660 -1620 18690 -1590
rect 18605 -1675 18635 -1645
rect 18275 -1720 18305 -1690
rect 18495 -1720 18525 -1690
rect 17895 -1805 17925 -1775
rect 17675 -1855 17705 -1825
rect 19330 -1930 19360 -1900
rect 16265 -1975 16295 -1945
rect 16485 -1975 16515 -1945
rect 16735 -1975 16765 -1945
rect 17200 -1975 17230 -1945
rect 17430 -1950 17465 -1945
rect 17430 -1975 17435 -1950
rect 17435 -1975 17460 -1950
rect 17460 -1975 17465 -1950
rect 17430 -1980 17465 -1975
rect 18129 -1950 18164 -1945
rect 18129 -1975 18134 -1950
rect 18134 -1975 18159 -1950
rect 18159 -1975 18164 -1950
rect 18129 -1980 18164 -1975
rect 19085 -1980 19115 -1950
rect 16485 -2905 16520 -2900
rect 16485 -2930 16490 -2905
rect 16490 -2930 16515 -2905
rect 16515 -2930 16520 -2905
rect 16485 -2935 16520 -2930
rect 16160 -3030 16195 -3025
rect 16160 -3055 16165 -3030
rect 16165 -3055 16190 -3030
rect 16190 -3055 16195 -3030
rect 16160 -3060 16195 -3055
rect 17200 -2045 17230 -2015
rect 18835 -2045 18865 -2015
rect 15825 -3145 15855 -3115
rect 15950 -3121 15985 -3116
rect 15950 -3146 15955 -3121
rect 15955 -3146 15980 -3121
rect 15980 -3146 15985 -3121
rect 16735 -3135 16765 -3105
rect 15950 -3151 15985 -3146
rect 17785 -3135 17815 -3105
rect 19080 -2905 19115 -2900
rect 19080 -2930 19085 -2905
rect 19085 -2930 19110 -2905
rect 19110 -2930 19115 -2905
rect 19080 -2935 19115 -2930
rect 19615 250 19645 280
rect 19540 -1805 19570 -1775
rect 19465 -1980 19495 -1950
rect 19405 -2997 19440 -2992
rect 19405 -3022 19410 -2997
rect 19410 -3022 19435 -2997
rect 19435 -3022 19440 -2997
rect 19405 -3027 19440 -3022
rect 18620 -3135 18650 -3105
rect 18835 -3135 18865 -3105
rect 19735 -250 19765 -220
rect 19610 -3121 19645 -3116
rect 19610 -3146 19615 -3121
rect 19615 -3146 19640 -3121
rect 19640 -3146 19645 -3121
rect 19610 -3151 19645 -3146
rect 15950 -3794 15985 -3789
rect 15950 -3819 15955 -3794
rect 15955 -3819 15980 -3794
rect 15980 -3819 15985 -3794
rect 15950 -3824 15985 -3819
rect 15825 -4295 15855 -4265
rect 15730 -4345 15760 -4315
rect 16280 -3899 16315 -3894
rect 16280 -3924 16285 -3899
rect 16285 -3924 16310 -3899
rect 16310 -3924 16315 -3899
rect 16280 -3929 16315 -3924
rect 16605 -3974 16640 -3969
rect 16605 -3999 16610 -3974
rect 16610 -3999 16635 -3974
rect 16635 -3999 16640 -3974
rect 19610 -3794 19645 -3789
rect 19610 -3819 19615 -3794
rect 19615 -3819 19640 -3794
rect 19640 -3819 19645 -3794
rect 19610 -3824 19645 -3819
rect 19285 -3899 19320 -3894
rect 19285 -3924 19290 -3899
rect 19290 -3924 19315 -3899
rect 19315 -3924 19320 -3899
rect 19285 -3929 19320 -3924
rect 18960 -3974 18995 -3969
rect 16605 -4004 16640 -3999
rect 18960 -3999 18965 -3974
rect 18965 -3999 18990 -3974
rect 18990 -3999 18995 -3974
rect 18960 -4004 18995 -3999
rect 16545 -4065 16575 -4035
rect 16285 -4220 16315 -4190
rect 16545 -4220 16575 -4190
rect 16610 -4220 16640 -4190
rect 17260 -4295 17290 -4265
rect 17785 -4270 17815 -4265
rect 17785 -4290 17790 -4270
rect 17790 -4290 17810 -4270
rect 17810 -4290 17815 -4270
rect 17785 -4295 17815 -4290
rect 18960 -4295 18990 -4265
rect 19285 -4295 19315 -4265
rect 16910 -4345 16940 -4315
rect 18660 -4345 18690 -4315
rect 19780 -1375 19810 -1345
rect 19735 -4345 19765 -4315
rect 15955 -4390 15985 -4360
rect 16210 -4390 16240 -4360
rect 19360 -4390 19390 -4360
rect 19615 -4390 19645 -4360
rect 17960 -4440 17990 -4410
<< metal2 >>
rect 16865 1395 16905 1400
rect 16865 1365 16870 1395
rect 16900 1390 16905 1395
rect 16975 1395 17015 1400
rect 16975 1390 16980 1395
rect 16900 1370 16980 1390
rect 16900 1365 16905 1370
rect 16865 1360 16905 1365
rect 16975 1365 16980 1370
rect 17010 1390 17015 1395
rect 17085 1395 17125 1400
rect 17085 1390 17090 1395
rect 17010 1370 17090 1390
rect 17010 1365 17015 1370
rect 16975 1360 17015 1365
rect 17085 1365 17090 1370
rect 17120 1365 17125 1395
rect 17085 1360 17125 1365
rect 17615 1395 17655 1400
rect 17615 1365 17620 1395
rect 17650 1390 17655 1395
rect 17725 1395 17765 1400
rect 17725 1390 17730 1395
rect 17650 1370 17730 1390
rect 17650 1365 17655 1370
rect 17615 1360 17655 1365
rect 17725 1365 17730 1370
rect 17760 1390 17765 1395
rect 17835 1395 17875 1400
rect 17835 1390 17840 1395
rect 17760 1370 17840 1390
rect 17760 1365 17765 1370
rect 17725 1360 17765 1365
rect 17835 1365 17840 1370
rect 17870 1390 17875 1395
rect 17945 1395 17985 1400
rect 17945 1390 17950 1395
rect 17870 1370 17950 1390
rect 17870 1365 17875 1370
rect 17835 1360 17875 1365
rect 17945 1365 17950 1370
rect 17980 1365 17985 1395
rect 17945 1360 17985 1365
rect 18475 1395 18515 1400
rect 18475 1365 18480 1395
rect 18510 1390 18515 1395
rect 18585 1395 18625 1400
rect 18585 1390 18590 1395
rect 18510 1370 18590 1390
rect 18510 1365 18515 1370
rect 18475 1360 18515 1365
rect 18585 1365 18590 1370
rect 18620 1390 18625 1395
rect 18695 1395 18735 1400
rect 18695 1390 18700 1395
rect 18620 1370 18700 1390
rect 18620 1365 18625 1370
rect 18585 1360 18625 1365
rect 18695 1365 18700 1370
rect 18730 1365 18735 1395
rect 18695 1360 18735 1365
rect 16810 1350 16850 1355
rect 16810 1320 16815 1350
rect 16845 1345 16850 1350
rect 16920 1350 16960 1355
rect 16920 1345 16925 1350
rect 16845 1325 16925 1345
rect 16845 1320 16850 1325
rect 16810 1315 16850 1320
rect 16920 1320 16925 1325
rect 16955 1345 16960 1350
rect 17030 1350 17070 1355
rect 17030 1345 17035 1350
rect 16955 1325 17035 1345
rect 16955 1320 16960 1325
rect 16920 1315 16960 1320
rect 17030 1320 17035 1325
rect 17065 1345 17070 1350
rect 17140 1350 17180 1355
rect 17140 1345 17145 1350
rect 17065 1325 17145 1345
rect 17065 1320 17070 1325
rect 17030 1315 17070 1320
rect 17140 1320 17145 1325
rect 17175 1345 17180 1350
rect 17450 1350 17490 1355
rect 17450 1345 17455 1350
rect 17175 1325 17455 1345
rect 17175 1320 17180 1325
rect 17140 1315 17180 1320
rect 17450 1320 17455 1325
rect 17485 1345 17490 1350
rect 17560 1350 17600 1355
rect 17560 1345 17565 1350
rect 17485 1325 17565 1345
rect 17485 1320 17490 1325
rect 17450 1315 17490 1320
rect 17560 1320 17565 1325
rect 17595 1345 17600 1350
rect 17670 1350 17710 1355
rect 17670 1345 17675 1350
rect 17595 1325 17675 1345
rect 17595 1320 17600 1325
rect 17560 1315 17600 1320
rect 17670 1320 17675 1325
rect 17705 1345 17710 1350
rect 17780 1350 17820 1355
rect 17780 1345 17785 1350
rect 17705 1325 17785 1345
rect 17705 1320 17710 1325
rect 17670 1315 17710 1320
rect 17780 1320 17785 1325
rect 17815 1345 17820 1350
rect 17890 1350 17930 1355
rect 17890 1345 17895 1350
rect 17815 1325 17895 1345
rect 17815 1320 17820 1325
rect 17780 1315 17820 1320
rect 17890 1320 17895 1325
rect 17925 1345 17930 1350
rect 18000 1350 18040 1355
rect 18000 1345 18005 1350
rect 17925 1325 18005 1345
rect 17925 1320 17930 1325
rect 17890 1315 17930 1320
rect 18000 1320 18005 1325
rect 18035 1345 18040 1350
rect 18110 1350 18150 1355
rect 18110 1345 18115 1350
rect 18035 1325 18115 1345
rect 18035 1320 18040 1325
rect 18000 1315 18040 1320
rect 18110 1320 18115 1325
rect 18145 1345 18150 1350
rect 18420 1350 18460 1355
rect 18420 1345 18425 1350
rect 18145 1325 18425 1345
rect 18145 1320 18150 1325
rect 18110 1315 18150 1320
rect 18420 1320 18425 1325
rect 18455 1345 18460 1350
rect 18530 1350 18570 1355
rect 18530 1345 18535 1350
rect 18455 1325 18535 1345
rect 18455 1320 18460 1325
rect 18420 1315 18460 1320
rect 18530 1320 18535 1325
rect 18565 1345 18570 1350
rect 18640 1350 18680 1355
rect 18640 1345 18645 1350
rect 18565 1325 18645 1345
rect 18565 1320 18570 1325
rect 18530 1315 18570 1320
rect 18640 1320 18645 1325
rect 18675 1345 18680 1350
rect 18750 1350 18790 1355
rect 18750 1345 18755 1350
rect 18675 1325 18755 1345
rect 18675 1320 18680 1325
rect 18640 1315 18680 1320
rect 18750 1320 18755 1325
rect 18785 1345 18790 1350
rect 20050 1350 20090 1355
rect 20050 1345 20055 1350
rect 18785 1325 20055 1345
rect 18785 1320 18790 1325
rect 18750 1315 18790 1320
rect 20050 1320 20055 1325
rect 20085 1320 20090 1350
rect 20050 1315 20090 1320
rect 16865 1195 16905 1200
rect 16865 1165 16870 1195
rect 16900 1190 16905 1195
rect 16975 1195 17015 1200
rect 16975 1190 16980 1195
rect 16900 1170 16980 1190
rect 16900 1165 16905 1170
rect 16865 1160 16905 1165
rect 16975 1165 16980 1170
rect 17010 1190 17015 1195
rect 17085 1195 17125 1200
rect 17085 1190 17090 1195
rect 17010 1170 17090 1190
rect 17010 1165 17015 1170
rect 16975 1160 17015 1165
rect 17085 1165 17090 1170
rect 17120 1165 17125 1195
rect 17085 1160 17125 1165
rect 17615 1195 17655 1200
rect 17615 1165 17620 1195
rect 17650 1190 17655 1195
rect 17725 1195 17765 1200
rect 17725 1190 17730 1195
rect 17650 1170 17730 1190
rect 17650 1165 17655 1170
rect 17615 1160 17655 1165
rect 17725 1165 17730 1170
rect 17760 1190 17765 1195
rect 17835 1195 17875 1200
rect 17835 1190 17840 1195
rect 17760 1170 17840 1190
rect 17760 1165 17765 1170
rect 17725 1160 17765 1165
rect 17835 1165 17840 1170
rect 17870 1190 17875 1195
rect 17945 1195 17985 1200
rect 17945 1190 17950 1195
rect 17870 1170 17950 1190
rect 17870 1165 17875 1170
rect 17835 1160 17875 1165
rect 17945 1165 17950 1170
rect 17980 1165 17985 1195
rect 17945 1160 17985 1165
rect 18475 1195 18515 1200
rect 18475 1165 18480 1195
rect 18510 1190 18515 1195
rect 18585 1195 18625 1200
rect 18585 1190 18590 1195
rect 18510 1170 18590 1190
rect 18510 1165 18515 1170
rect 18475 1160 18515 1165
rect 18585 1165 18590 1170
rect 18620 1190 18625 1195
rect 18695 1195 18735 1200
rect 18695 1190 18700 1195
rect 18620 1170 18700 1190
rect 18620 1165 18625 1170
rect 18585 1160 18625 1165
rect 18695 1165 18700 1170
rect 18730 1165 18735 1195
rect 18695 1160 18735 1165
rect 16810 1150 16850 1155
rect 16810 1120 16815 1150
rect 16845 1145 16850 1150
rect 16920 1150 16960 1155
rect 16920 1145 16925 1150
rect 16845 1125 16925 1145
rect 16845 1120 16850 1125
rect 16810 1115 16850 1120
rect 16920 1120 16925 1125
rect 16955 1145 16960 1150
rect 17030 1150 17070 1155
rect 17030 1145 17035 1150
rect 16955 1125 17035 1145
rect 16955 1120 16960 1125
rect 16920 1115 16960 1120
rect 17030 1120 17035 1125
rect 17065 1145 17070 1150
rect 17140 1150 17180 1155
rect 17140 1145 17145 1150
rect 17065 1125 17145 1145
rect 17065 1120 17070 1125
rect 17030 1115 17070 1120
rect 17140 1120 17145 1125
rect 17175 1120 17180 1150
rect 17140 1115 17180 1120
rect 17450 1150 17490 1155
rect 17450 1120 17455 1150
rect 17485 1145 17490 1150
rect 17560 1150 17600 1155
rect 17560 1145 17565 1150
rect 17485 1125 17565 1145
rect 17485 1120 17490 1125
rect 17450 1115 17490 1120
rect 17560 1120 17565 1125
rect 17595 1145 17600 1150
rect 17670 1150 17710 1155
rect 17670 1145 17675 1150
rect 17595 1125 17675 1145
rect 17595 1120 17600 1125
rect 17560 1115 17600 1120
rect 17670 1120 17675 1125
rect 17705 1145 17710 1150
rect 17780 1150 17820 1155
rect 17780 1145 17785 1150
rect 17705 1125 17785 1145
rect 17705 1120 17710 1125
rect 17670 1115 17710 1120
rect 17780 1120 17785 1125
rect 17815 1145 17820 1150
rect 17890 1150 17930 1155
rect 17890 1145 17895 1150
rect 17815 1125 17895 1145
rect 17815 1120 17820 1125
rect 17780 1115 17820 1120
rect 17890 1120 17895 1125
rect 17925 1145 17930 1150
rect 18000 1150 18040 1155
rect 18000 1145 18005 1150
rect 17925 1125 18005 1145
rect 17925 1120 17930 1125
rect 17890 1115 17930 1120
rect 18000 1120 18005 1125
rect 18035 1145 18040 1150
rect 18110 1150 18150 1155
rect 18110 1145 18115 1150
rect 18035 1125 18115 1145
rect 18035 1120 18040 1125
rect 18000 1115 18040 1120
rect 18110 1120 18115 1125
rect 18145 1120 18150 1150
rect 18110 1115 18150 1120
rect 18420 1150 18460 1155
rect 18420 1120 18425 1150
rect 18455 1145 18460 1150
rect 18530 1150 18570 1155
rect 18530 1145 18535 1150
rect 18455 1125 18535 1145
rect 18455 1120 18460 1125
rect 18420 1115 18460 1120
rect 18530 1120 18535 1125
rect 18565 1145 18570 1150
rect 18640 1150 18680 1155
rect 18640 1145 18645 1150
rect 18565 1125 18645 1145
rect 18565 1120 18570 1125
rect 18530 1115 18570 1120
rect 18640 1120 18645 1125
rect 18675 1145 18680 1150
rect 18750 1150 18790 1155
rect 18750 1145 18755 1150
rect 18675 1125 18755 1145
rect 18675 1120 18680 1125
rect 18640 1115 18680 1120
rect 18750 1120 18755 1125
rect 18785 1120 18790 1150
rect 18750 1115 18790 1120
rect 17070 1095 17100 1100
rect 17805 1095 17835 1100
rect 17100 1070 17805 1090
rect 17070 1060 17100 1065
rect 18500 1095 18530 1100
rect 17835 1070 18500 1090
rect 17805 1060 17835 1065
rect 18720 1095 18760 1100
rect 18720 1090 18725 1095
rect 18530 1070 18725 1090
rect 18500 1060 18530 1065
rect 18720 1065 18725 1070
rect 18755 1065 18760 1095
rect 18720 1060 18760 1065
rect 16160 1050 16200 1055
rect 16160 1020 16165 1050
rect 16195 1045 16200 1050
rect 17505 1050 17545 1055
rect 17505 1045 17510 1050
rect 16195 1025 17510 1045
rect 16195 1020 16200 1025
rect 16160 1015 16200 1020
rect 17505 1020 17510 1025
rect 17540 1020 17545 1050
rect 18055 1050 18095 1055
rect 17505 1015 17545 1020
rect 17600 1020 17640 1025
rect 17600 990 17605 1020
rect 17635 1015 17640 1020
rect 17960 1020 18000 1025
rect 17960 1015 17965 1020
rect 17635 995 17965 1015
rect 17635 990 17640 995
rect 17600 985 17640 990
rect 17960 990 17965 995
rect 17995 990 18000 1020
rect 18055 1020 18060 1050
rect 18090 1045 18095 1050
rect 19325 1050 19365 1055
rect 19325 1045 19330 1050
rect 18090 1025 19330 1045
rect 18090 1020 18095 1025
rect 18055 1015 18095 1020
rect 19325 1020 19330 1025
rect 19360 1020 19365 1050
rect 19325 1015 19365 1020
rect 17960 985 18000 990
rect 17420 975 17460 980
rect 17420 945 17425 975
rect 17455 970 17460 975
rect 18140 975 18180 980
rect 18140 970 18145 975
rect 17455 950 18145 970
rect 17455 945 17460 950
rect 17420 940 17460 945
rect 18140 945 18145 950
rect 18175 945 18180 975
rect 18140 940 18180 945
rect 17240 930 17280 935
rect 17240 900 17245 930
rect 17275 925 17280 930
rect 18320 930 18360 935
rect 18320 925 18325 930
rect 17275 905 18325 925
rect 17275 900 17280 905
rect 17240 895 17280 900
rect 18320 900 18325 905
rect 18355 900 18360 930
rect 18320 895 18360 900
rect 17060 885 17100 890
rect 17060 855 17065 885
rect 17095 880 17100 885
rect 17780 885 17820 890
rect 17780 880 17785 885
rect 17095 860 17785 880
rect 17095 855 17100 860
rect 17060 850 17100 855
rect 17780 855 17785 860
rect 17815 880 17820 885
rect 18500 885 18540 890
rect 18500 880 18505 885
rect 17815 860 18505 880
rect 17815 855 17820 860
rect 17780 850 17820 855
rect 18500 855 18505 860
rect 18535 855 18540 885
rect 18500 850 18540 855
rect 16435 840 16475 845
rect 16435 810 16440 840
rect 16470 835 16475 840
rect 16655 840 16695 845
rect 16655 835 16660 840
rect 16470 815 16660 835
rect 16470 810 16475 815
rect 16435 805 16475 810
rect 16655 810 16660 815
rect 16690 835 16695 840
rect 16970 840 17010 845
rect 16970 835 16975 840
rect 16690 815 16975 835
rect 16690 810 16695 815
rect 16655 805 16695 810
rect 16970 810 16975 815
rect 17005 835 17010 840
rect 17150 840 17190 845
rect 17150 835 17155 840
rect 17005 815 17155 835
rect 17005 810 17010 815
rect 16970 805 17010 810
rect 17150 810 17155 815
rect 17185 835 17190 840
rect 17330 840 17370 845
rect 17330 835 17335 840
rect 17185 815 17335 835
rect 17185 810 17190 815
rect 17150 805 17190 810
rect 17330 810 17335 815
rect 17365 835 17370 840
rect 17510 840 17550 845
rect 17510 835 17515 840
rect 17365 815 17515 835
rect 17365 810 17370 815
rect 17330 805 17370 810
rect 17510 810 17515 815
rect 17545 835 17550 840
rect 17690 840 17730 845
rect 17690 835 17695 840
rect 17545 815 17695 835
rect 17545 810 17550 815
rect 17510 805 17550 810
rect 17690 810 17695 815
rect 17725 835 17730 840
rect 17870 840 17910 845
rect 17870 835 17875 840
rect 17725 815 17875 835
rect 17725 810 17730 815
rect 17690 805 17730 810
rect 17870 810 17875 815
rect 17905 835 17910 840
rect 18050 840 18090 845
rect 18050 835 18055 840
rect 17905 815 18055 835
rect 17905 810 17910 815
rect 17870 805 17910 810
rect 18050 810 18055 815
rect 18085 835 18090 840
rect 18230 840 18270 845
rect 18230 835 18235 840
rect 18085 815 18235 835
rect 18085 810 18090 815
rect 18050 805 18090 810
rect 18230 810 18235 815
rect 18265 835 18270 840
rect 18410 840 18450 845
rect 18410 835 18415 840
rect 18265 815 18415 835
rect 18265 810 18270 815
rect 18230 805 18270 810
rect 18410 810 18415 815
rect 18445 835 18450 840
rect 18590 840 18630 845
rect 18590 835 18595 840
rect 18445 815 18595 835
rect 18445 810 18450 815
rect 18410 805 18450 810
rect 18590 810 18595 815
rect 18625 835 18630 840
rect 19010 840 19050 845
rect 19010 835 19015 840
rect 18625 815 19015 835
rect 18625 810 18630 815
rect 18590 805 18630 810
rect 19010 810 19015 815
rect 19045 835 19050 840
rect 20050 840 20090 845
rect 20050 835 20055 840
rect 19045 815 20055 835
rect 19045 810 19050 815
rect 19010 805 19050 810
rect 20050 810 20055 815
rect 20085 810 20090 840
rect 20050 805 20090 810
rect 16440 780 16470 785
rect 16440 745 16470 750
rect 16490 780 16530 785
rect 16490 750 16495 780
rect 16525 775 16530 780
rect 16600 780 16640 785
rect 16600 775 16605 780
rect 16525 755 16605 775
rect 16525 750 16530 755
rect 16490 745 16530 750
rect 16600 750 16605 755
rect 16635 750 16640 780
rect 16600 745 16640 750
rect 16660 780 16690 785
rect 16660 745 16690 750
rect 18900 780 18940 785
rect 18900 750 18905 780
rect 18935 775 18940 780
rect 19010 780 19050 785
rect 19010 775 19015 780
rect 18935 755 19015 775
rect 18935 750 18940 755
rect 18900 745 18940 750
rect 19010 750 19015 755
rect 19045 775 19050 780
rect 19120 780 19160 785
rect 19120 775 19125 780
rect 19045 755 19125 775
rect 19045 750 19050 755
rect 19010 745 19050 750
rect 19120 750 19125 755
rect 19155 750 19160 780
rect 19120 745 19160 750
rect 16545 735 16585 740
rect 16545 705 16550 735
rect 16580 730 16585 735
rect 16780 735 16820 740
rect 16780 730 16785 735
rect 16580 710 16785 730
rect 16580 705 16585 710
rect 16545 700 16585 705
rect 16780 705 16785 710
rect 16815 705 16820 735
rect 16780 700 16820 705
rect 18955 735 18995 740
rect 18955 705 18960 735
rect 18990 730 18995 735
rect 19065 735 19105 740
rect 19065 730 19070 735
rect 18990 710 19070 730
rect 18990 705 18995 710
rect 18955 700 18995 705
rect 19065 705 19070 710
rect 19100 705 19105 735
rect 19065 700 19105 705
rect 16490 595 16530 600
rect 16490 565 16495 595
rect 16525 590 16530 595
rect 16600 595 16640 600
rect 16600 590 16605 595
rect 16525 570 16605 590
rect 16525 565 16530 570
rect 16490 560 16530 565
rect 16600 565 16605 570
rect 16635 590 16640 595
rect 16840 595 16880 600
rect 16840 590 16845 595
rect 16635 570 16845 590
rect 16635 565 16640 570
rect 16600 560 16640 565
rect 16840 565 16845 570
rect 16875 565 16880 595
rect 16840 560 16880 565
rect 18900 595 18940 600
rect 18900 565 18905 595
rect 18935 590 18940 595
rect 19010 595 19050 600
rect 19010 590 19015 595
rect 18935 570 19015 590
rect 18935 565 18940 570
rect 18900 560 18940 565
rect 19010 565 19015 570
rect 19045 590 19050 595
rect 19120 595 19160 600
rect 19120 590 19125 595
rect 19045 570 19125 590
rect 19045 565 19050 570
rect 19010 560 19050 565
rect 19120 565 19125 570
rect 19155 565 19160 595
rect 19120 560 19160 565
rect 16435 550 16475 555
rect 16435 520 16440 550
rect 16470 545 16475 550
rect 16655 550 16695 555
rect 16655 545 16660 550
rect 16470 525 16660 545
rect 16470 520 16475 525
rect 16435 515 16475 520
rect 16655 520 16660 525
rect 16690 520 16695 550
rect 16655 515 16695 520
rect 18955 550 18995 555
rect 18955 520 18960 550
rect 18990 545 18995 550
rect 19065 550 19105 555
rect 19065 545 19070 550
rect 18990 525 19070 545
rect 18990 520 18995 525
rect 18955 515 18995 520
rect 19065 520 19070 525
rect 19100 545 19105 550
rect 19260 550 19300 555
rect 19260 545 19265 550
rect 19100 525 19265 545
rect 19100 520 19105 525
rect 19065 515 19105 520
rect 19260 520 19265 525
rect 19295 520 19300 550
rect 19260 515 19300 520
rect 16305 485 16345 490
rect 16305 455 16310 485
rect 16340 480 16345 485
rect 17600 485 17640 490
rect 17600 480 17605 485
rect 16340 460 17605 480
rect 16340 455 16345 460
rect 16305 450 16345 455
rect 17600 455 17605 460
rect 17635 480 17640 485
rect 17960 485 18000 490
rect 17960 480 17965 485
rect 17635 460 17965 480
rect 17635 455 17640 460
rect 17600 450 17640 455
rect 17960 455 17965 460
rect 17995 480 18000 485
rect 19460 485 19500 490
rect 19460 480 19465 485
rect 17995 460 19465 480
rect 17995 455 18000 460
rect 17960 450 18000 455
rect 19460 455 19465 460
rect 19495 455 19500 485
rect 19460 450 19500 455
rect 16260 430 16300 435
rect 16260 400 16265 430
rect 16295 425 16300 430
rect 16780 430 16820 435
rect 16780 425 16785 430
rect 16295 405 16785 425
rect 16295 400 16300 405
rect 16260 395 16300 400
rect 16780 400 16785 405
rect 16815 425 16820 430
rect 17420 430 17460 435
rect 17420 425 17425 430
rect 16815 405 17425 425
rect 16815 400 16820 405
rect 16780 395 16820 400
rect 17420 400 17425 405
rect 17455 425 17460 430
rect 18140 430 18180 435
rect 18140 425 18145 430
rect 17455 405 18145 425
rect 17455 400 17460 405
rect 17420 395 17460 400
rect 18140 400 18145 405
rect 18175 400 18180 430
rect 18140 395 18180 400
rect 16205 385 16245 390
rect 16205 355 16210 385
rect 16240 380 16245 385
rect 16545 385 16585 390
rect 16545 380 16550 385
rect 16240 360 16550 380
rect 16240 355 16245 360
rect 16205 350 16245 355
rect 16545 355 16550 360
rect 16580 380 16585 385
rect 17240 385 17280 390
rect 17240 380 17245 385
rect 16580 360 17245 380
rect 16580 355 16585 360
rect 16545 350 16585 355
rect 17240 355 17245 360
rect 17275 380 17280 385
rect 18320 385 18360 390
rect 18320 380 18325 385
rect 17275 360 18325 380
rect 17275 355 17280 360
rect 17240 350 17280 355
rect 18320 355 18325 360
rect 18355 355 18360 385
rect 18320 350 18360 355
rect 17060 340 17100 345
rect 17060 310 17065 340
rect 17095 335 17100 340
rect 17780 340 17820 345
rect 17780 335 17785 340
rect 17095 315 17785 335
rect 17095 310 17100 315
rect 17060 305 17100 310
rect 17780 310 17785 315
rect 17815 335 17820 340
rect 18500 340 18540 345
rect 18500 335 18505 340
rect 17815 315 18505 335
rect 17815 310 17820 315
rect 17780 305 17820 310
rect 18500 310 18505 315
rect 18535 335 18540 340
rect 19405 340 19445 345
rect 19405 335 19410 340
rect 18535 315 19410 335
rect 18535 310 18540 315
rect 18500 305 18540 310
rect 19405 310 19410 315
rect 19440 310 19445 340
rect 19405 305 19445 310
rect 18720 280 18760 285
rect 18720 250 18725 280
rect 18755 275 18760 280
rect 19010 280 19050 285
rect 19010 275 19015 280
rect 18755 255 19015 275
rect 18755 250 18760 255
rect 18720 245 18760 250
rect 19010 250 19015 255
rect 19045 275 19050 280
rect 19610 280 19650 285
rect 19610 275 19615 280
rect 19045 255 19615 275
rect 19045 250 19050 255
rect 19010 245 19050 250
rect 19610 250 19615 255
rect 19645 250 19650 280
rect 19610 245 19650 250
rect 16420 225 16460 230
rect 16420 195 16425 225
rect 16455 220 16460 225
rect 16540 225 16580 230
rect 16540 220 16545 225
rect 16455 200 16545 220
rect 16455 195 16460 200
rect 16420 190 16460 195
rect 16540 195 16545 200
rect 16575 220 16580 225
rect 16660 225 16700 230
rect 16660 220 16665 225
rect 16575 200 16665 220
rect 16575 195 16580 200
rect 16540 190 16580 195
rect 16660 195 16665 200
rect 16695 220 16700 225
rect 16780 225 16820 230
rect 16780 220 16785 225
rect 16695 200 16785 220
rect 16695 195 16700 200
rect 16660 190 16700 195
rect 16780 195 16785 200
rect 16815 220 16820 225
rect 16900 225 16940 230
rect 16900 220 16905 225
rect 16815 200 16905 220
rect 16815 195 16820 200
rect 16780 190 16820 195
rect 16900 195 16905 200
rect 16935 220 16940 225
rect 17020 225 17060 230
rect 17020 220 17025 225
rect 16935 200 17025 220
rect 16935 195 16940 200
rect 16900 190 16940 195
rect 17020 195 17025 200
rect 17055 220 17060 225
rect 17140 225 17180 230
rect 17140 220 17145 225
rect 17055 200 17145 220
rect 17055 195 17060 200
rect 17020 190 17060 195
rect 17140 195 17145 200
rect 17175 220 17180 225
rect 17260 225 17300 230
rect 17260 220 17265 225
rect 17175 200 17265 220
rect 17175 195 17180 200
rect 17140 190 17180 195
rect 17260 195 17265 200
rect 17295 220 17300 225
rect 17380 225 17420 230
rect 17380 220 17385 225
rect 17295 200 17385 220
rect 17295 195 17300 200
rect 17260 190 17300 195
rect 17380 195 17385 200
rect 17415 220 17420 225
rect 17500 225 17540 230
rect 17500 220 17505 225
rect 17415 200 17505 220
rect 17415 195 17420 200
rect 17380 190 17420 195
rect 17500 195 17505 200
rect 17535 220 17540 225
rect 17620 225 17660 230
rect 17620 220 17625 225
rect 17535 200 17625 220
rect 17535 195 17540 200
rect 17500 190 17540 195
rect 17620 195 17625 200
rect 17655 220 17660 225
rect 17940 225 17980 230
rect 17940 220 17945 225
rect 17655 200 17945 220
rect 17655 195 17660 200
rect 17620 190 17660 195
rect 17940 195 17945 200
rect 17975 220 17980 225
rect 18060 225 18100 230
rect 18060 220 18065 225
rect 17975 200 18065 220
rect 17975 195 17980 200
rect 17940 190 17980 195
rect 18060 195 18065 200
rect 18095 220 18100 225
rect 18180 225 18220 230
rect 18180 220 18185 225
rect 18095 200 18185 220
rect 18095 195 18100 200
rect 18060 190 18100 195
rect 18180 195 18185 200
rect 18215 220 18220 225
rect 18300 225 18340 230
rect 18300 220 18305 225
rect 18215 200 18305 220
rect 18215 195 18220 200
rect 18180 190 18220 195
rect 18300 195 18305 200
rect 18335 220 18340 225
rect 18420 225 18460 230
rect 18420 220 18425 225
rect 18335 200 18425 220
rect 18335 195 18340 200
rect 18300 190 18340 195
rect 18420 195 18425 200
rect 18455 220 18460 225
rect 18540 225 18580 230
rect 18540 220 18545 225
rect 18455 200 18545 220
rect 18455 195 18460 200
rect 18420 190 18460 195
rect 18540 195 18545 200
rect 18575 220 18580 225
rect 18660 225 18700 230
rect 18660 220 18665 225
rect 18575 200 18665 220
rect 18575 195 18580 200
rect 18540 190 18580 195
rect 18660 195 18665 200
rect 18695 220 18700 225
rect 18780 225 18820 230
rect 18780 220 18785 225
rect 18695 200 18785 220
rect 18695 195 18700 200
rect 18660 190 18700 195
rect 18780 195 18785 200
rect 18815 220 18820 225
rect 18900 225 18940 230
rect 18900 220 18905 225
rect 18815 200 18905 220
rect 18815 195 18820 200
rect 18780 190 18820 195
rect 18900 195 18905 200
rect 18935 220 18940 225
rect 19020 225 19060 230
rect 19020 220 19025 225
rect 18935 200 19025 220
rect 18935 195 18940 200
rect 18900 190 18940 195
rect 19020 195 19025 200
rect 19055 220 19060 225
rect 19140 225 19180 230
rect 19140 220 19145 225
rect 19055 200 19145 220
rect 19055 195 19060 200
rect 19020 190 19060 195
rect 19140 195 19145 200
rect 19175 220 19180 225
rect 20050 225 20090 230
rect 20050 220 20055 225
rect 19175 200 20055 220
rect 19175 195 19180 200
rect 19140 190 19180 195
rect 20050 195 20055 200
rect 20085 195 20090 225
rect 20050 190 20090 195
rect 15950 175 15990 180
rect 15950 145 15955 175
rect 15985 170 15990 175
rect 16480 175 16520 180
rect 16480 170 16485 175
rect 15985 150 16485 170
rect 15985 145 15990 150
rect 15950 140 15990 145
rect 16480 145 16485 150
rect 16515 170 16520 175
rect 16840 175 16880 180
rect 16840 170 16845 175
rect 16515 150 16845 170
rect 16515 145 16520 150
rect 16480 140 16520 145
rect 16840 145 16845 150
rect 16875 170 16880 175
rect 17200 175 17240 180
rect 17200 170 17205 175
rect 16875 150 17205 170
rect 16875 145 16880 150
rect 16840 140 16880 145
rect 17200 145 17205 150
rect 17235 170 17240 175
rect 17560 175 17600 180
rect 17560 170 17565 175
rect 17235 150 17565 170
rect 17235 145 17240 150
rect 17200 140 17240 145
rect 17560 145 17565 150
rect 17595 170 17600 175
rect 17690 175 17730 180
rect 17690 170 17695 175
rect 17595 150 17695 170
rect 17595 145 17600 150
rect 17560 140 17600 145
rect 17690 145 17695 150
rect 17725 145 17730 175
rect 17690 140 17730 145
rect 17870 175 17910 180
rect 17870 145 17875 175
rect 17905 170 17910 175
rect 18000 175 18040 180
rect 18000 170 18005 175
rect 17905 150 18005 170
rect 17905 145 17910 150
rect 17870 140 17910 145
rect 18000 145 18005 150
rect 18035 170 18040 175
rect 18360 175 18400 180
rect 18360 170 18365 175
rect 18035 150 18365 170
rect 18035 145 18040 150
rect 18000 140 18040 145
rect 18360 145 18365 150
rect 18395 170 18400 175
rect 18720 175 18760 180
rect 18720 170 18725 175
rect 18395 150 18725 170
rect 18395 145 18400 150
rect 18360 140 18400 145
rect 18720 145 18725 150
rect 18755 170 18760 175
rect 19080 175 19120 180
rect 19080 170 19085 175
rect 18755 150 19085 170
rect 18755 145 18760 150
rect 18720 140 18760 145
rect 19080 145 19085 150
rect 19115 145 19120 175
rect 19080 140 19120 145
rect 16720 130 16760 135
rect 16720 100 16725 130
rect 16755 125 16760 130
rect 17080 130 17120 135
rect 17080 125 17085 130
rect 16755 105 17085 125
rect 16755 100 16760 105
rect 16720 95 16760 100
rect 17080 100 17085 105
rect 17115 125 17120 130
rect 17440 130 17480 135
rect 17440 125 17445 130
rect 17115 105 17445 125
rect 17115 100 17120 105
rect 17080 95 17120 100
rect 17440 100 17445 105
rect 17475 100 17480 130
rect 17440 95 17480 100
rect 18120 130 18160 135
rect 18120 100 18125 130
rect 18155 125 18160 130
rect 18480 130 18520 135
rect 18480 125 18485 130
rect 18155 105 18485 125
rect 18155 100 18160 105
rect 18120 95 18160 100
rect 18480 100 18485 105
rect 18515 125 18520 130
rect 18840 130 18880 135
rect 18840 125 18845 130
rect 18515 105 18845 125
rect 18515 100 18520 105
rect 18480 95 18520 100
rect 18840 100 18845 105
rect 18875 100 18880 130
rect 18840 95 18880 100
rect 16600 85 16640 90
rect 16600 55 16605 85
rect 16635 80 16640 85
rect 16960 85 17000 90
rect 16960 80 16965 85
rect 16635 60 16965 80
rect 16635 55 16640 60
rect 16600 50 16640 55
rect 16960 55 16965 60
rect 16995 80 17000 85
rect 17320 85 17360 90
rect 17320 80 17325 85
rect 16995 60 17325 80
rect 16995 55 17000 60
rect 16960 50 17000 55
rect 17320 55 17325 60
rect 17355 55 17360 85
rect 18240 85 18280 90
rect 17440 60 17480 80
rect 18120 60 18160 80
rect 17320 50 17360 55
rect 18240 55 18245 85
rect 18275 80 18280 85
rect 18600 85 18640 90
rect 18600 80 18605 85
rect 18275 60 18605 80
rect 18275 55 18280 60
rect 18240 50 18280 55
rect 18600 55 18605 60
rect 18635 80 18640 85
rect 18960 85 19000 90
rect 18960 80 18965 85
rect 18635 60 18965 80
rect 18635 55 18640 60
rect 18600 50 18640 55
rect 18960 55 18965 60
rect 18995 55 19000 85
rect 18960 50 19000 55
rect 16600 -70 16640 -65
rect 16600 -100 16605 -70
rect 16635 -75 16640 -70
rect 16960 -70 17000 -65
rect 16960 -75 16965 -70
rect 16635 -95 16965 -75
rect 16635 -100 16640 -95
rect 16600 -105 16640 -100
rect 16960 -100 16965 -95
rect 16995 -75 17000 -70
rect 17320 -70 17360 -65
rect 17320 -75 17325 -70
rect 16995 -95 17325 -75
rect 16995 -100 17000 -95
rect 16960 -105 17000 -100
rect 17320 -100 17325 -95
rect 17355 -100 17360 -70
rect 17320 -105 17360 -100
rect 18240 -70 18280 -65
rect 18240 -100 18245 -70
rect 18275 -75 18280 -70
rect 18600 -70 18640 -65
rect 18600 -75 18605 -70
rect 18275 -95 18605 -75
rect 18275 -100 18280 -95
rect 18240 -105 18280 -100
rect 18600 -100 18605 -95
rect 18635 -75 18640 -70
rect 18960 -70 19000 -65
rect 18960 -75 18965 -70
rect 18635 -95 18965 -75
rect 18635 -100 18640 -95
rect 18600 -105 18640 -100
rect 18960 -100 18965 -95
rect 18995 -100 19000 -70
rect 18960 -105 19000 -100
rect 16480 -115 16520 -110
rect 16480 -145 16485 -115
rect 16515 -120 16520 -115
rect 16840 -115 16880 -110
rect 16840 -120 16845 -115
rect 16515 -140 16845 -120
rect 16515 -145 16520 -140
rect 16480 -150 16520 -145
rect 16840 -145 16845 -140
rect 16875 -120 16880 -115
rect 17200 -115 17240 -110
rect 17200 -120 17205 -115
rect 16875 -140 17205 -120
rect 16875 -145 16880 -140
rect 16840 -150 16880 -145
rect 17200 -145 17205 -140
rect 17235 -120 17240 -115
rect 17560 -115 17600 -110
rect 17560 -120 17565 -115
rect 17235 -140 17565 -120
rect 17235 -145 17240 -140
rect 17200 -150 17240 -145
rect 17560 -145 17565 -140
rect 17595 -145 17600 -115
rect 17560 -150 17600 -145
rect 18000 -115 18040 -110
rect 18000 -145 18005 -115
rect 18035 -120 18040 -115
rect 18360 -115 18400 -110
rect 18360 -120 18365 -115
rect 18035 -140 18365 -120
rect 18035 -145 18040 -140
rect 18000 -150 18040 -145
rect 18360 -145 18365 -140
rect 18395 -120 18400 -115
rect 18720 -115 18760 -110
rect 18720 -120 18725 -115
rect 18395 -140 18725 -120
rect 18395 -145 18400 -140
rect 18360 -150 18400 -145
rect 18720 -145 18725 -140
rect 18755 -120 18760 -115
rect 19080 -115 19120 -110
rect 19080 -120 19085 -115
rect 18755 -140 19085 -120
rect 18755 -145 18760 -140
rect 18720 -150 18760 -145
rect 19080 -145 19085 -140
rect 19115 -145 19120 -115
rect 19080 -150 19120 -145
rect 16420 -165 16460 -160
rect 16420 -195 16425 -165
rect 16455 -170 16460 -165
rect 16540 -165 16580 -160
rect 16540 -170 16545 -165
rect 16455 -190 16545 -170
rect 16455 -195 16460 -190
rect 16420 -200 16460 -195
rect 16540 -195 16545 -190
rect 16575 -170 16580 -165
rect 16660 -165 16700 -160
rect 16660 -170 16665 -165
rect 16575 -190 16665 -170
rect 16575 -195 16580 -190
rect 16540 -200 16580 -195
rect 16660 -195 16665 -190
rect 16695 -170 16700 -165
rect 16780 -165 16820 -160
rect 16780 -170 16785 -165
rect 16695 -190 16785 -170
rect 16695 -195 16700 -190
rect 16660 -200 16700 -195
rect 16780 -195 16785 -190
rect 16815 -170 16820 -165
rect 16900 -165 16940 -160
rect 16900 -170 16905 -165
rect 16815 -190 16905 -170
rect 16815 -195 16820 -190
rect 16780 -200 16820 -195
rect 16900 -195 16905 -190
rect 16935 -170 16940 -165
rect 17020 -165 17060 -160
rect 17020 -170 17025 -165
rect 16935 -190 17025 -170
rect 16935 -195 16940 -190
rect 16900 -200 16940 -195
rect 17020 -195 17025 -190
rect 17055 -170 17060 -165
rect 17140 -165 17180 -160
rect 17140 -170 17145 -165
rect 17055 -190 17145 -170
rect 17055 -195 17060 -190
rect 17020 -200 17060 -195
rect 17140 -195 17145 -190
rect 17175 -170 17180 -165
rect 17260 -165 17300 -160
rect 17260 -170 17265 -165
rect 17175 -190 17265 -170
rect 17175 -195 17180 -190
rect 17140 -200 17180 -195
rect 17260 -195 17265 -190
rect 17295 -170 17300 -165
rect 17380 -165 17420 -160
rect 17380 -170 17385 -165
rect 17295 -190 17385 -170
rect 17295 -195 17300 -190
rect 17260 -200 17300 -195
rect 17380 -195 17385 -190
rect 17415 -170 17420 -165
rect 17500 -165 17540 -160
rect 17500 -170 17505 -165
rect 17415 -190 17505 -170
rect 17415 -195 17420 -190
rect 17380 -200 17420 -195
rect 17500 -195 17505 -190
rect 17535 -170 17540 -165
rect 17620 -165 17660 -160
rect 17620 -170 17625 -165
rect 17535 -190 17625 -170
rect 17535 -195 17540 -190
rect 17500 -200 17540 -195
rect 17620 -195 17625 -190
rect 17655 -195 17660 -165
rect 17620 -200 17660 -195
rect 17940 -165 17980 -160
rect 17940 -195 17945 -165
rect 17975 -170 17980 -165
rect 18060 -165 18100 -160
rect 18060 -170 18065 -165
rect 17975 -190 18065 -170
rect 17975 -195 17980 -190
rect 17940 -200 17980 -195
rect 18060 -195 18065 -190
rect 18095 -170 18100 -165
rect 18180 -165 18220 -160
rect 18180 -170 18185 -165
rect 18095 -190 18185 -170
rect 18095 -195 18100 -190
rect 18060 -200 18100 -195
rect 18180 -195 18185 -190
rect 18215 -170 18220 -165
rect 18300 -165 18340 -160
rect 18300 -170 18305 -165
rect 18215 -190 18305 -170
rect 18215 -195 18220 -190
rect 18180 -200 18220 -195
rect 18300 -195 18305 -190
rect 18335 -170 18340 -165
rect 18420 -165 18460 -160
rect 18420 -170 18425 -165
rect 18335 -190 18425 -170
rect 18335 -195 18340 -190
rect 18300 -200 18340 -195
rect 18420 -195 18425 -190
rect 18455 -170 18460 -165
rect 18540 -165 18580 -160
rect 18540 -170 18545 -165
rect 18455 -190 18545 -170
rect 18455 -195 18460 -190
rect 18420 -200 18460 -195
rect 18540 -195 18545 -190
rect 18575 -170 18580 -165
rect 18660 -165 18700 -160
rect 18660 -170 18665 -165
rect 18575 -190 18665 -170
rect 18575 -195 18580 -190
rect 18540 -200 18580 -195
rect 18660 -195 18665 -190
rect 18695 -170 18700 -165
rect 18780 -165 18820 -160
rect 18780 -170 18785 -165
rect 18695 -190 18785 -170
rect 18695 -195 18700 -190
rect 18660 -200 18700 -195
rect 18780 -195 18785 -190
rect 18815 -170 18820 -165
rect 18900 -165 18940 -160
rect 18900 -170 18905 -165
rect 18815 -190 18905 -170
rect 18815 -195 18820 -190
rect 18780 -200 18820 -195
rect 18900 -195 18905 -190
rect 18935 -170 18940 -165
rect 19020 -165 19060 -160
rect 19020 -170 19025 -165
rect 18935 -190 19025 -170
rect 18935 -195 18940 -190
rect 18900 -200 18940 -195
rect 19020 -195 19025 -190
rect 19055 -170 19060 -165
rect 19140 -165 19180 -160
rect 19140 -170 19145 -165
rect 19055 -190 19145 -170
rect 19055 -195 19060 -190
rect 19020 -200 19060 -195
rect 19140 -195 19145 -190
rect 19175 -195 19180 -165
rect 19140 -200 19180 -195
rect 15725 -215 15765 -210
rect 15725 -245 15730 -215
rect 15760 -225 15765 -215
rect 16540 -220 16570 -215
rect 15760 -245 16540 -225
rect 15725 -250 15765 -245
rect 16720 -220 16760 -215
rect 16720 -225 16725 -220
rect 16570 -245 16725 -225
rect 16540 -255 16570 -250
rect 16720 -250 16725 -245
rect 16755 -225 16760 -220
rect 16900 -220 16930 -215
rect 16755 -245 16900 -225
rect 16755 -250 16760 -245
rect 16720 -255 16760 -250
rect 17080 -220 17120 -215
rect 17080 -225 17085 -220
rect 16930 -245 17085 -225
rect 16900 -255 16930 -250
rect 17080 -250 17085 -245
rect 17115 -225 17120 -220
rect 17260 -220 17290 -215
rect 17115 -245 17260 -225
rect 17115 -250 17120 -245
rect 17080 -255 17120 -250
rect 17440 -220 17480 -215
rect 17440 -225 17445 -220
rect 17290 -245 17445 -225
rect 17260 -255 17290 -250
rect 17440 -250 17445 -245
rect 17475 -225 17480 -220
rect 17510 -220 17540 -215
rect 17475 -245 17510 -225
rect 17475 -250 17480 -245
rect 17440 -255 17480 -250
rect 17510 -255 17540 -250
rect 18060 -220 18090 -215
rect 18120 -220 18160 -215
rect 18120 -225 18125 -220
rect 18090 -245 18125 -225
rect 18060 -255 18090 -250
rect 18120 -250 18125 -245
rect 18155 -225 18160 -220
rect 18310 -220 18340 -215
rect 18155 -245 18310 -225
rect 18155 -250 18160 -245
rect 18120 -255 18160 -250
rect 18480 -220 18520 -215
rect 18480 -225 18485 -220
rect 18340 -245 18485 -225
rect 18310 -255 18340 -250
rect 18480 -250 18485 -245
rect 18515 -225 18520 -220
rect 18670 -220 18700 -215
rect 18515 -245 18670 -225
rect 18515 -250 18520 -245
rect 18480 -255 18520 -250
rect 18840 -220 18880 -215
rect 18840 -225 18845 -220
rect 18700 -245 18845 -225
rect 18670 -255 18700 -250
rect 18840 -250 18845 -245
rect 18875 -225 18880 -220
rect 19030 -220 19060 -215
rect 18875 -245 19030 -225
rect 18875 -250 18880 -245
rect 18840 -255 18880 -250
rect 19730 -220 19770 -215
rect 19730 -225 19735 -220
rect 19060 -245 19735 -225
rect 19030 -255 19060 -250
rect 19730 -250 19735 -245
rect 19765 -250 19770 -220
rect 19730 -255 19770 -250
rect 16910 -325 16950 -320
rect 16910 -355 16915 -325
rect 16945 -330 16950 -325
rect 17030 -325 17070 -320
rect 17030 -330 17035 -325
rect 16945 -350 17035 -330
rect 16945 -355 16950 -350
rect 16910 -360 16950 -355
rect 17030 -355 17035 -350
rect 17065 -330 17070 -325
rect 17150 -325 17190 -320
rect 17150 -330 17155 -325
rect 17065 -350 17155 -330
rect 17065 -355 17070 -350
rect 17030 -360 17070 -355
rect 17150 -355 17155 -350
rect 17185 -330 17190 -325
rect 17270 -325 17310 -320
rect 17270 -330 17275 -325
rect 17185 -350 17275 -330
rect 17185 -355 17190 -350
rect 17150 -360 17190 -355
rect 17270 -355 17275 -350
rect 17305 -330 17310 -325
rect 17390 -325 17430 -320
rect 17390 -330 17395 -325
rect 17305 -350 17395 -330
rect 17305 -355 17310 -350
rect 17270 -360 17310 -355
rect 17390 -355 17395 -350
rect 17425 -355 17430 -325
rect 17390 -360 17430 -355
rect 18170 -325 18210 -320
rect 18170 -355 18175 -325
rect 18205 -330 18210 -325
rect 18290 -325 18330 -320
rect 18290 -330 18295 -325
rect 18205 -350 18295 -330
rect 18205 -355 18210 -350
rect 18170 -360 18210 -355
rect 18290 -355 18295 -350
rect 18325 -330 18330 -325
rect 18410 -325 18450 -320
rect 18410 -330 18415 -325
rect 18325 -350 18415 -330
rect 18325 -355 18330 -350
rect 18290 -360 18330 -355
rect 18410 -355 18415 -350
rect 18445 -330 18450 -325
rect 18530 -325 18570 -320
rect 18530 -330 18535 -325
rect 18445 -350 18535 -330
rect 18445 -355 18450 -350
rect 18410 -360 18450 -355
rect 18530 -355 18535 -350
rect 18565 -330 18570 -325
rect 18650 -325 18690 -320
rect 18650 -330 18655 -325
rect 18565 -350 18655 -330
rect 18565 -355 18570 -350
rect 18530 -360 18570 -355
rect 18650 -355 18655 -350
rect 18685 -355 18690 -325
rect 18650 -360 18690 -355
rect 16970 -370 17010 -365
rect 16260 -390 16300 -385
rect 16260 -420 16265 -390
rect 16295 -395 16300 -390
rect 16800 -390 16830 -385
rect 16295 -415 16800 -395
rect 16295 -420 16300 -415
rect 16260 -425 16300 -420
rect 16970 -400 16975 -370
rect 17005 -375 17010 -370
rect 17210 -370 17250 -365
rect 17210 -375 17215 -370
rect 17005 -395 17215 -375
rect 17005 -400 17010 -395
rect 16970 -405 17010 -400
rect 17210 -400 17215 -395
rect 17245 -375 17250 -370
rect 17450 -370 17490 -365
rect 17450 -375 17455 -370
rect 17245 -395 17455 -375
rect 17245 -400 17250 -395
rect 17210 -405 17250 -400
rect 17450 -400 17455 -395
rect 17485 -400 17490 -370
rect 17450 -405 17490 -400
rect 18110 -370 18150 -365
rect 18110 -400 18115 -370
rect 18145 -375 18150 -370
rect 18350 -370 18390 -365
rect 18350 -375 18355 -370
rect 18145 -395 18355 -375
rect 18145 -400 18150 -395
rect 18110 -405 18150 -400
rect 18350 -400 18355 -395
rect 18385 -375 18390 -370
rect 18590 -370 18630 -365
rect 18590 -375 18595 -370
rect 18385 -395 18595 -375
rect 18385 -400 18390 -395
rect 18350 -405 18390 -400
rect 18590 -400 18595 -395
rect 18625 -400 18630 -370
rect 18590 -405 18630 -400
rect 18770 -390 18800 -385
rect 16800 -425 16830 -420
rect 16850 -415 16890 -410
rect 16850 -445 16855 -415
rect 16885 -420 16890 -415
rect 17090 -415 17130 -410
rect 17090 -420 17095 -415
rect 16885 -440 17095 -420
rect 16885 -445 16890 -440
rect 16850 -450 16890 -445
rect 17090 -445 17095 -440
rect 17125 -420 17130 -415
rect 17330 -415 17370 -410
rect 17330 -420 17335 -415
rect 17125 -440 17335 -420
rect 17125 -445 17130 -440
rect 17090 -450 17130 -445
rect 17330 -445 17335 -440
rect 17365 -445 17370 -415
rect 18230 -415 18270 -410
rect 17390 -440 17430 -420
rect 18170 -440 18210 -420
rect 17330 -450 17370 -445
rect 18230 -445 18235 -415
rect 18265 -420 18270 -415
rect 18470 -415 18510 -410
rect 18470 -420 18475 -415
rect 18265 -440 18475 -420
rect 18265 -445 18270 -440
rect 18230 -450 18270 -445
rect 18470 -445 18475 -440
rect 18505 -420 18510 -415
rect 18710 -415 18750 -410
rect 18710 -420 18715 -415
rect 18505 -440 18715 -420
rect 18505 -445 18510 -440
rect 18470 -450 18510 -445
rect 18710 -445 18715 -440
rect 18745 -445 18750 -415
rect 19405 -390 19445 -385
rect 19405 -395 19410 -390
rect 18800 -415 19410 -395
rect 18770 -425 18800 -420
rect 19405 -420 19410 -415
rect 19440 -420 19445 -390
rect 19405 -425 19445 -420
rect 18710 -450 18750 -445
rect 17565 -460 17595 -455
rect 17780 -460 17820 -455
rect 17780 -465 17785 -460
rect 17595 -485 17785 -465
rect 17565 -495 17595 -490
rect 17780 -490 17785 -485
rect 17815 -465 17820 -460
rect 18005 -460 18035 -455
rect 17815 -485 18005 -465
rect 17815 -490 17820 -485
rect 17780 -495 17820 -490
rect 18005 -495 18035 -490
rect 16970 -505 17010 -500
rect 16305 -530 16345 -525
rect 16305 -560 16310 -530
rect 16340 -535 16345 -530
rect 16800 -530 16830 -525
rect 16340 -555 16800 -535
rect 16340 -560 16345 -555
rect 16305 -565 16345 -560
rect 16970 -535 16975 -505
rect 17005 -510 17010 -505
rect 17210 -505 17250 -500
rect 17210 -510 17215 -505
rect 17005 -530 17215 -510
rect 17005 -535 17010 -530
rect 16970 -540 17010 -535
rect 17210 -535 17215 -530
rect 17245 -510 17250 -505
rect 17450 -505 17490 -500
rect 17450 -510 17455 -505
rect 17245 -530 17455 -510
rect 17245 -535 17250 -530
rect 17210 -540 17250 -535
rect 17450 -535 17455 -530
rect 17485 -535 17490 -505
rect 17450 -540 17490 -535
rect 18110 -505 18150 -500
rect 18110 -535 18115 -505
rect 18145 -510 18150 -505
rect 18350 -505 18390 -500
rect 18350 -510 18355 -505
rect 18145 -530 18355 -510
rect 18145 -535 18150 -530
rect 18110 -540 18150 -535
rect 18350 -535 18355 -530
rect 18385 -510 18390 -505
rect 18590 -505 18630 -500
rect 18590 -510 18595 -505
rect 18385 -530 18595 -510
rect 18385 -535 18390 -530
rect 18350 -540 18390 -535
rect 18590 -535 18595 -530
rect 18625 -535 18630 -505
rect 18590 -540 18630 -535
rect 18770 -530 18800 -525
rect 16800 -565 16830 -560
rect 16850 -550 16890 -545
rect 16850 -580 16855 -550
rect 16885 -555 16890 -550
rect 17090 -550 17130 -545
rect 17090 -555 17095 -550
rect 16885 -575 17095 -555
rect 16885 -580 16890 -575
rect 16850 -585 16890 -580
rect 17090 -580 17095 -575
rect 17125 -555 17130 -550
rect 17330 -550 17370 -545
rect 17330 -555 17335 -550
rect 17125 -575 17335 -555
rect 17125 -580 17130 -575
rect 17090 -585 17130 -580
rect 17330 -580 17335 -575
rect 17365 -580 17370 -550
rect 17330 -585 17370 -580
rect 18230 -550 18270 -545
rect 18230 -580 18235 -550
rect 18265 -555 18270 -550
rect 18470 -550 18510 -545
rect 18470 -555 18475 -550
rect 18265 -575 18475 -555
rect 18265 -580 18270 -575
rect 18230 -585 18270 -580
rect 18470 -580 18475 -575
rect 18505 -555 18510 -550
rect 18710 -550 18750 -545
rect 18710 -555 18715 -550
rect 18505 -575 18715 -555
rect 18505 -580 18510 -575
rect 18470 -585 18510 -580
rect 18710 -580 18715 -575
rect 18745 -580 18750 -550
rect 19325 -530 19365 -525
rect 19325 -535 19330 -530
rect 18800 -555 19330 -535
rect 18770 -565 18800 -560
rect 19325 -560 19330 -555
rect 19360 -560 19365 -530
rect 19325 -565 19365 -560
rect 18710 -585 18750 -580
rect 16530 -595 16570 -590
rect 16530 -625 16535 -595
rect 16565 -600 16570 -595
rect 16910 -595 16950 -590
rect 16910 -600 16915 -595
rect 16565 -620 16915 -600
rect 16565 -625 16570 -620
rect 16530 -630 16570 -625
rect 16910 -625 16915 -620
rect 16945 -600 16950 -595
rect 17030 -595 17070 -590
rect 17030 -600 17035 -595
rect 16945 -620 17035 -600
rect 16945 -625 16950 -620
rect 16910 -630 16950 -625
rect 17030 -625 17035 -620
rect 17065 -600 17070 -595
rect 17150 -595 17190 -590
rect 17150 -600 17155 -595
rect 17065 -620 17155 -600
rect 17065 -625 17070 -620
rect 17030 -630 17070 -625
rect 17150 -625 17155 -620
rect 17185 -600 17190 -595
rect 17270 -595 17310 -590
rect 17270 -600 17275 -595
rect 17185 -620 17275 -600
rect 17185 -625 17190 -620
rect 17150 -630 17190 -625
rect 17270 -625 17275 -620
rect 17305 -600 17310 -595
rect 17390 -595 17430 -590
rect 17390 -600 17395 -595
rect 17305 -620 17395 -600
rect 17305 -625 17310 -620
rect 17270 -630 17310 -625
rect 17390 -625 17395 -620
rect 17425 -625 17430 -595
rect 17390 -630 17430 -625
rect 18170 -595 18210 -590
rect 18170 -625 18175 -595
rect 18205 -600 18210 -595
rect 18290 -595 18330 -590
rect 18290 -600 18295 -595
rect 18205 -620 18295 -600
rect 18205 -625 18210 -620
rect 18170 -630 18210 -625
rect 18290 -625 18295 -620
rect 18325 -600 18330 -595
rect 18410 -595 18450 -590
rect 18410 -600 18415 -595
rect 18325 -620 18415 -600
rect 18325 -625 18330 -620
rect 18290 -630 18330 -625
rect 18410 -625 18415 -620
rect 18445 -600 18450 -595
rect 18530 -595 18570 -590
rect 18530 -600 18535 -595
rect 18445 -620 18535 -600
rect 18445 -625 18450 -620
rect 18410 -630 18450 -625
rect 18530 -625 18535 -620
rect 18565 -600 18570 -595
rect 18650 -595 18690 -590
rect 18650 -600 18655 -595
rect 18565 -620 18655 -600
rect 18565 -625 18570 -620
rect 18530 -630 18570 -625
rect 18650 -625 18655 -620
rect 18685 -600 18690 -595
rect 19030 -595 19070 -590
rect 19030 -600 19035 -595
rect 18685 -620 19035 -600
rect 18685 -625 18690 -620
rect 18650 -630 18690 -625
rect 19030 -625 19035 -620
rect 19065 -625 19070 -595
rect 19030 -630 19070 -625
rect 16800 -680 16840 -675
rect 16800 -710 16805 -680
rect 16835 -685 16840 -680
rect 17420 -680 17460 -675
rect 17420 -685 17425 -680
rect 16835 -705 17425 -685
rect 16835 -710 16840 -705
rect 16800 -715 16840 -710
rect 17420 -710 17425 -705
rect 17455 -685 17460 -680
rect 18140 -680 18180 -675
rect 18140 -685 18145 -680
rect 17455 -705 18145 -685
rect 17455 -710 17460 -705
rect 17420 -715 17460 -710
rect 18140 -710 18145 -705
rect 18175 -685 18180 -680
rect 18760 -680 18800 -675
rect 18760 -685 18765 -680
rect 18175 -705 18765 -685
rect 18175 -710 18180 -705
rect 18140 -715 18180 -710
rect 18760 -710 18765 -705
rect 18795 -685 18800 -680
rect 20050 -680 20090 -675
rect 20050 -685 20055 -680
rect 18795 -705 20055 -685
rect 18795 -710 18800 -705
rect 18760 -715 18800 -710
rect 20050 -710 20055 -705
rect 20085 -710 20090 -680
rect 20050 -715 20090 -710
rect 17110 -995 17150 -990
rect 17110 -1025 17115 -995
rect 17145 -1000 17150 -995
rect 17780 -995 17820 -990
rect 17780 -1000 17785 -995
rect 17145 -1020 17785 -1000
rect 17145 -1025 17150 -1020
rect 17110 -1030 17150 -1025
rect 17780 -1025 17785 -1020
rect 17815 -1000 17820 -995
rect 18450 -995 18490 -990
rect 18450 -1000 18455 -995
rect 17815 -1020 18455 -1000
rect 17815 -1025 17820 -1020
rect 17780 -1030 17820 -1025
rect 18450 -1025 18455 -1020
rect 18485 -1000 18490 -995
rect 19965 -995 20005 -990
rect 19965 -1000 19970 -995
rect 18485 -1020 19970 -1000
rect 18485 -1025 18490 -1020
rect 18450 -1030 18490 -1025
rect 19965 -1025 19970 -1020
rect 20000 -1025 20005 -995
rect 19965 -1030 20005 -1025
rect 16205 -1095 16245 -1090
rect 16205 -1125 16210 -1095
rect 16240 -1100 16245 -1095
rect 16740 -1095 16780 -1090
rect 16740 -1100 16745 -1095
rect 16240 -1120 16745 -1100
rect 16240 -1125 16245 -1120
rect 16205 -1130 16245 -1125
rect 16740 -1125 16745 -1120
rect 16775 -1100 16780 -1095
rect 17260 -1095 17300 -1090
rect 17260 -1100 17265 -1095
rect 16775 -1120 17265 -1100
rect 16775 -1125 16780 -1120
rect 16740 -1130 16780 -1125
rect 17260 -1125 17265 -1120
rect 17295 -1125 17300 -1095
rect 17260 -1130 17300 -1125
rect 17780 -1095 17820 -1090
rect 17780 -1125 17785 -1095
rect 17815 -1100 17820 -1095
rect 18300 -1095 18340 -1090
rect 18300 -1100 18305 -1095
rect 17815 -1120 18305 -1100
rect 17815 -1125 17820 -1120
rect 17780 -1130 17820 -1125
rect 18300 -1125 18305 -1120
rect 18335 -1125 18340 -1095
rect 18300 -1130 18340 -1125
rect 18895 -1180 18935 -1175
rect 18895 -1210 18900 -1180
rect 18930 -1185 18935 -1180
rect 19965 -1180 20005 -1175
rect 19965 -1185 19970 -1180
rect 18930 -1205 19970 -1185
rect 18930 -1210 18935 -1205
rect 18895 -1215 18935 -1210
rect 19965 -1210 19970 -1205
rect 20000 -1210 20005 -1180
rect 19965 -1215 20005 -1210
rect 17285 -1335 17315 -1330
rect 15785 -1345 15825 -1340
rect 15785 -1375 15790 -1345
rect 15820 -1350 15825 -1345
rect 16970 -1345 17010 -1340
rect 16970 -1350 16975 -1345
rect 15820 -1370 16975 -1350
rect 15820 -1375 15825 -1370
rect 15785 -1380 15825 -1375
rect 16970 -1375 16975 -1370
rect 17005 -1350 17010 -1345
rect 17190 -1345 17230 -1340
rect 17190 -1350 17195 -1345
rect 17005 -1370 17195 -1350
rect 17005 -1375 17010 -1370
rect 16970 -1380 17010 -1375
rect 17190 -1375 17195 -1370
rect 17225 -1375 17230 -1345
rect 17785 -1335 17815 -1330
rect 17315 -1360 17785 -1340
rect 17285 -1370 17315 -1365
rect 18295 -1335 18325 -1330
rect 17815 -1360 18295 -1340
rect 17785 -1370 17815 -1365
rect 18295 -1370 18325 -1365
rect 18380 -1345 18420 -1340
rect 17190 -1380 17230 -1375
rect 18380 -1375 18385 -1345
rect 18415 -1350 18420 -1345
rect 18600 -1345 18640 -1340
rect 18600 -1350 18605 -1345
rect 18415 -1370 18605 -1350
rect 18415 -1375 18420 -1370
rect 18380 -1380 18420 -1375
rect 18600 -1375 18605 -1370
rect 18635 -1350 18640 -1345
rect 19775 -1345 19815 -1340
rect 19775 -1350 19780 -1345
rect 18635 -1370 19780 -1350
rect 18635 -1375 18640 -1370
rect 18600 -1380 18640 -1375
rect 19775 -1375 19780 -1370
rect 19810 -1375 19815 -1345
rect 19775 -1380 19815 -1375
rect 17080 -1390 17120 -1385
rect 17080 -1420 17085 -1390
rect 17115 -1395 17120 -1390
rect 17300 -1390 17340 -1385
rect 17300 -1395 17305 -1390
rect 17115 -1415 17305 -1395
rect 17115 -1420 17120 -1415
rect 17080 -1425 17120 -1420
rect 17300 -1420 17305 -1415
rect 17335 -1420 17340 -1390
rect 17300 -1425 17340 -1420
rect 17780 -1390 17820 -1385
rect 17780 -1420 17785 -1390
rect 17815 -1395 17820 -1390
rect 17890 -1390 17930 -1385
rect 17890 -1395 17895 -1390
rect 17815 -1415 17895 -1395
rect 17815 -1420 17820 -1415
rect 17780 -1425 17820 -1420
rect 17890 -1420 17895 -1415
rect 17925 -1395 17930 -1390
rect 18000 -1390 18040 -1385
rect 18000 -1395 18005 -1390
rect 17925 -1415 18005 -1395
rect 17925 -1420 17930 -1415
rect 17890 -1425 17930 -1420
rect 18000 -1420 18005 -1415
rect 18035 -1420 18040 -1390
rect 18000 -1425 18040 -1420
rect 18270 -1390 18310 -1385
rect 18270 -1420 18275 -1390
rect 18305 -1395 18310 -1390
rect 18490 -1390 18530 -1385
rect 18490 -1395 18495 -1390
rect 18305 -1415 18495 -1395
rect 18305 -1420 18310 -1415
rect 18270 -1425 18310 -1420
rect 18490 -1420 18495 -1415
rect 18525 -1420 18530 -1390
rect 18490 -1425 18530 -1420
rect 16915 -1435 16955 -1430
rect 16915 -1465 16920 -1435
rect 16950 -1440 16955 -1435
rect 17025 -1435 17065 -1430
rect 17025 -1440 17030 -1435
rect 16950 -1460 17030 -1440
rect 16950 -1465 16955 -1460
rect 16915 -1470 16955 -1465
rect 17025 -1465 17030 -1460
rect 17060 -1440 17065 -1435
rect 17135 -1435 17175 -1430
rect 17135 -1440 17140 -1435
rect 17060 -1460 17140 -1440
rect 17060 -1465 17065 -1460
rect 17025 -1470 17065 -1465
rect 17135 -1465 17140 -1460
rect 17170 -1440 17175 -1435
rect 17245 -1435 17285 -1430
rect 17245 -1440 17250 -1435
rect 17170 -1460 17250 -1440
rect 17170 -1465 17175 -1460
rect 17135 -1470 17175 -1465
rect 17245 -1465 17250 -1460
rect 17280 -1440 17285 -1435
rect 17355 -1435 17395 -1430
rect 17355 -1440 17360 -1435
rect 17280 -1460 17360 -1440
rect 17280 -1465 17285 -1460
rect 17245 -1470 17285 -1465
rect 17355 -1465 17360 -1460
rect 17390 -1440 17395 -1435
rect 17505 -1435 17545 -1430
rect 17505 -1440 17510 -1435
rect 17390 -1460 17510 -1440
rect 17390 -1465 17395 -1460
rect 17355 -1470 17395 -1465
rect 17505 -1465 17510 -1460
rect 17540 -1440 17545 -1435
rect 17615 -1435 17655 -1430
rect 17615 -1440 17620 -1435
rect 17540 -1460 17620 -1440
rect 17540 -1465 17545 -1460
rect 17505 -1470 17545 -1465
rect 17615 -1465 17620 -1460
rect 17650 -1440 17655 -1435
rect 17725 -1435 17765 -1430
rect 17725 -1440 17730 -1435
rect 17650 -1460 17730 -1440
rect 17650 -1465 17655 -1460
rect 17615 -1470 17655 -1465
rect 17725 -1465 17730 -1460
rect 17760 -1440 17765 -1435
rect 17835 -1435 17875 -1430
rect 17835 -1440 17840 -1435
rect 17760 -1460 17840 -1440
rect 17760 -1465 17765 -1460
rect 17725 -1470 17765 -1465
rect 17835 -1465 17840 -1460
rect 17870 -1440 17875 -1435
rect 17945 -1435 17985 -1430
rect 17945 -1440 17950 -1435
rect 17870 -1460 17950 -1440
rect 17870 -1465 17875 -1460
rect 17835 -1470 17875 -1465
rect 17945 -1465 17950 -1460
rect 17980 -1440 17985 -1435
rect 18055 -1435 18095 -1430
rect 18055 -1440 18060 -1435
rect 17980 -1460 18060 -1440
rect 17980 -1465 17985 -1460
rect 17945 -1470 17985 -1465
rect 18055 -1465 18060 -1460
rect 18090 -1440 18095 -1435
rect 18215 -1435 18255 -1430
rect 18215 -1440 18220 -1435
rect 18090 -1460 18220 -1440
rect 18090 -1465 18095 -1460
rect 18055 -1470 18095 -1465
rect 18215 -1465 18220 -1460
rect 18250 -1440 18255 -1435
rect 18325 -1435 18365 -1430
rect 18325 -1440 18330 -1435
rect 18250 -1460 18330 -1440
rect 18250 -1465 18255 -1460
rect 18215 -1470 18255 -1465
rect 18325 -1465 18330 -1460
rect 18360 -1440 18365 -1435
rect 18435 -1435 18475 -1430
rect 18435 -1440 18440 -1435
rect 18360 -1460 18440 -1440
rect 18360 -1465 18365 -1460
rect 18325 -1470 18365 -1465
rect 18435 -1465 18440 -1460
rect 18470 -1440 18475 -1435
rect 18545 -1435 18585 -1430
rect 18545 -1440 18550 -1435
rect 18470 -1460 18550 -1440
rect 18470 -1465 18475 -1460
rect 18435 -1470 18475 -1465
rect 18545 -1465 18550 -1460
rect 18580 -1440 18585 -1435
rect 18655 -1435 18695 -1430
rect 18655 -1440 18660 -1435
rect 18580 -1460 18660 -1440
rect 18580 -1465 18585 -1460
rect 18545 -1470 18585 -1465
rect 18655 -1465 18660 -1460
rect 18690 -1440 18695 -1435
rect 19965 -1435 20005 -1430
rect 19965 -1440 19970 -1435
rect 18690 -1460 19970 -1440
rect 18690 -1465 18695 -1460
rect 18655 -1470 18695 -1465
rect 19965 -1465 19970 -1460
rect 20000 -1465 20005 -1435
rect 19965 -1470 20005 -1465
rect 16915 -1590 16955 -1585
rect 16915 -1620 16920 -1590
rect 16950 -1595 16955 -1590
rect 17025 -1590 17065 -1585
rect 17025 -1595 17030 -1590
rect 16950 -1615 17030 -1595
rect 16950 -1620 16955 -1615
rect 16915 -1625 16955 -1620
rect 17025 -1620 17030 -1615
rect 17060 -1595 17065 -1590
rect 17135 -1590 17175 -1585
rect 17135 -1595 17140 -1590
rect 17060 -1615 17140 -1595
rect 17060 -1620 17065 -1615
rect 17025 -1625 17065 -1620
rect 17135 -1620 17140 -1615
rect 17170 -1595 17175 -1590
rect 17245 -1590 17285 -1585
rect 17245 -1595 17250 -1590
rect 17170 -1615 17250 -1595
rect 17170 -1620 17175 -1615
rect 17135 -1625 17175 -1620
rect 17245 -1620 17250 -1615
rect 17280 -1595 17285 -1590
rect 17355 -1590 17395 -1585
rect 17355 -1595 17360 -1590
rect 17280 -1615 17360 -1595
rect 17280 -1620 17285 -1615
rect 17245 -1625 17285 -1620
rect 17355 -1620 17360 -1615
rect 17390 -1620 17395 -1590
rect 17355 -1625 17395 -1620
rect 17505 -1590 17545 -1585
rect 17505 -1620 17510 -1590
rect 17540 -1595 17545 -1590
rect 17615 -1590 17655 -1585
rect 17615 -1595 17620 -1590
rect 17540 -1615 17620 -1595
rect 17540 -1620 17545 -1615
rect 17505 -1625 17545 -1620
rect 17615 -1620 17620 -1615
rect 17650 -1595 17655 -1590
rect 17725 -1590 17765 -1585
rect 17725 -1595 17730 -1590
rect 17650 -1615 17730 -1595
rect 17650 -1620 17655 -1615
rect 17615 -1625 17655 -1620
rect 17725 -1620 17730 -1615
rect 17760 -1595 17765 -1590
rect 17835 -1590 17875 -1585
rect 17835 -1595 17840 -1590
rect 17760 -1615 17840 -1595
rect 17760 -1620 17765 -1615
rect 17725 -1625 17765 -1620
rect 17835 -1620 17840 -1615
rect 17870 -1595 17875 -1590
rect 17945 -1590 17985 -1585
rect 17945 -1595 17950 -1590
rect 17870 -1615 17950 -1595
rect 17870 -1620 17875 -1615
rect 17835 -1625 17875 -1620
rect 17945 -1620 17950 -1615
rect 17980 -1595 17985 -1590
rect 18055 -1590 18095 -1585
rect 18055 -1595 18060 -1590
rect 17980 -1615 18060 -1595
rect 17980 -1620 17985 -1615
rect 17945 -1625 17985 -1620
rect 18055 -1620 18060 -1615
rect 18090 -1620 18095 -1590
rect 18055 -1625 18095 -1620
rect 18215 -1590 18255 -1585
rect 18215 -1620 18220 -1590
rect 18250 -1595 18255 -1590
rect 18325 -1590 18365 -1585
rect 18325 -1595 18330 -1590
rect 18250 -1615 18330 -1595
rect 18250 -1620 18255 -1615
rect 18215 -1625 18255 -1620
rect 18325 -1620 18330 -1615
rect 18360 -1595 18365 -1590
rect 18435 -1590 18475 -1585
rect 18435 -1595 18440 -1590
rect 18360 -1615 18440 -1595
rect 18360 -1620 18365 -1615
rect 18325 -1625 18365 -1620
rect 18435 -1620 18440 -1615
rect 18470 -1595 18475 -1590
rect 18545 -1590 18585 -1585
rect 18545 -1595 18550 -1590
rect 18470 -1615 18550 -1595
rect 18470 -1620 18475 -1615
rect 18435 -1625 18475 -1620
rect 18545 -1620 18550 -1615
rect 18580 -1595 18585 -1590
rect 18655 -1590 18695 -1585
rect 18655 -1595 18660 -1590
rect 18580 -1615 18660 -1595
rect 18580 -1620 18585 -1615
rect 18545 -1625 18585 -1620
rect 18655 -1620 18660 -1615
rect 18690 -1620 18695 -1590
rect 18655 -1625 18695 -1620
rect 17670 -1635 17710 -1630
rect 16970 -1645 17010 -1640
rect 16970 -1675 16975 -1645
rect 17005 -1650 17010 -1645
rect 17190 -1645 17230 -1640
rect 17190 -1650 17195 -1645
rect 17005 -1670 17195 -1650
rect 17005 -1675 17010 -1670
rect 16970 -1680 17010 -1675
rect 17190 -1675 17195 -1670
rect 17225 -1675 17230 -1645
rect 17190 -1680 17230 -1675
rect 17585 -1645 17615 -1640
rect 17670 -1665 17675 -1635
rect 17705 -1665 17710 -1635
rect 17670 -1670 17710 -1665
rect 17780 -1635 17820 -1630
rect 17780 -1665 17785 -1635
rect 17815 -1640 17820 -1635
rect 17890 -1635 17930 -1630
rect 17890 -1640 17895 -1635
rect 17815 -1660 17895 -1640
rect 17815 -1665 17820 -1660
rect 17780 -1670 17820 -1665
rect 17890 -1665 17895 -1660
rect 17925 -1640 17930 -1635
rect 18000 -1635 18040 -1630
rect 18000 -1640 18005 -1635
rect 17925 -1660 18005 -1640
rect 17925 -1665 17930 -1660
rect 17890 -1670 17930 -1665
rect 18000 -1665 18005 -1660
rect 18035 -1665 18040 -1635
rect 18000 -1670 18040 -1665
rect 18380 -1645 18420 -1640
rect 17585 -1680 17615 -1675
rect 18380 -1675 18385 -1645
rect 18415 -1650 18420 -1645
rect 18600 -1645 18640 -1640
rect 18600 -1650 18605 -1645
rect 18415 -1670 18605 -1650
rect 18415 -1675 18420 -1670
rect 18380 -1680 18420 -1675
rect 18600 -1675 18605 -1670
rect 18635 -1675 18640 -1645
rect 18600 -1680 18640 -1675
rect 16030 -1690 16070 -1685
rect 16030 -1720 16035 -1690
rect 16065 -1695 16070 -1690
rect 17080 -1690 17120 -1685
rect 17080 -1695 17085 -1690
rect 16065 -1715 17085 -1695
rect 16065 -1720 16070 -1715
rect 16030 -1725 16070 -1720
rect 17080 -1720 17085 -1715
rect 17115 -1695 17120 -1690
rect 17300 -1690 17340 -1685
rect 17300 -1695 17305 -1690
rect 17115 -1715 17305 -1695
rect 17115 -1720 17120 -1715
rect 17080 -1725 17120 -1720
rect 17300 -1720 17305 -1715
rect 17335 -1695 17340 -1690
rect 18270 -1690 18310 -1685
rect 18270 -1695 18275 -1690
rect 17335 -1715 18275 -1695
rect 17335 -1720 17340 -1715
rect 17300 -1725 17340 -1720
rect 18270 -1720 18275 -1715
rect 18305 -1695 18310 -1690
rect 18490 -1690 18530 -1685
rect 18490 -1695 18495 -1690
rect 18305 -1715 18495 -1695
rect 18305 -1720 18310 -1715
rect 18270 -1725 18310 -1720
rect 18490 -1720 18495 -1715
rect 18525 -1720 18530 -1690
rect 18490 -1725 18530 -1720
rect 17890 -1775 17930 -1770
rect 16160 -1780 16200 -1775
rect 16160 -1810 16165 -1780
rect 16195 -1785 16200 -1780
rect 17580 -1780 17620 -1775
rect 17580 -1785 17585 -1780
rect 16195 -1805 17585 -1785
rect 16195 -1810 16200 -1805
rect 16160 -1815 16200 -1810
rect 17580 -1810 17585 -1805
rect 17615 -1810 17620 -1780
rect 17890 -1805 17895 -1775
rect 17925 -1780 17930 -1775
rect 19535 -1775 19575 -1770
rect 19535 -1780 19540 -1775
rect 17925 -1800 19540 -1780
rect 17925 -1805 17930 -1800
rect 17890 -1810 17930 -1805
rect 19535 -1805 19540 -1800
rect 19570 -1805 19575 -1775
rect 19535 -1810 19575 -1805
rect 17580 -1815 17620 -1810
rect 16105 -1825 16145 -1820
rect 16105 -1855 16110 -1825
rect 16140 -1830 16145 -1825
rect 17670 -1825 17710 -1820
rect 17670 -1830 17675 -1825
rect 16140 -1850 17675 -1830
rect 16140 -1855 16145 -1850
rect 16105 -1860 16145 -1855
rect 17670 -1855 17675 -1850
rect 17705 -1855 17710 -1825
rect 17670 -1860 17710 -1855
rect 16155 -1900 16195 -1895
rect 16155 -1930 16160 -1900
rect 16190 -1905 16195 -1900
rect 19325 -1900 19365 -1895
rect 19325 -1905 19330 -1900
rect 16190 -1925 19330 -1905
rect 16190 -1930 16195 -1925
rect 16155 -1935 16195 -1930
rect 19325 -1930 19330 -1925
rect 19360 -1930 19365 -1900
rect 19325 -1935 19365 -1930
rect 16260 -1945 16300 -1940
rect 16260 -1975 16265 -1945
rect 16295 -1950 16300 -1945
rect 16480 -1945 16520 -1940
rect 16480 -1950 16485 -1945
rect 16295 -1970 16485 -1950
rect 16295 -1975 16300 -1970
rect 16260 -1980 16300 -1975
rect 16480 -1975 16485 -1970
rect 16515 -1950 16520 -1945
rect 16730 -1945 16770 -1940
rect 16730 -1950 16735 -1945
rect 16515 -1970 16735 -1950
rect 16515 -1975 16520 -1970
rect 16480 -1980 16520 -1975
rect 16730 -1975 16735 -1970
rect 16765 -1975 16770 -1945
rect 16730 -1980 16770 -1975
rect 17195 -1945 17235 -1940
rect 17195 -1975 17200 -1945
rect 17230 -1950 17235 -1945
rect 17425 -1950 17430 -1945
rect 17230 -1970 17430 -1950
rect 17230 -1975 17235 -1970
rect 17195 -1980 17235 -1975
rect 17425 -1980 17430 -1970
rect 17465 -1980 17470 -1945
rect 18124 -1980 18129 -1945
rect 18164 -1955 18169 -1945
rect 19080 -1950 19120 -1945
rect 19080 -1955 19085 -1950
rect 18164 -1975 19085 -1955
rect 18164 -1980 18169 -1975
rect 19080 -1980 19085 -1975
rect 19115 -1955 19120 -1950
rect 19460 -1950 19500 -1945
rect 19460 -1955 19465 -1950
rect 19115 -1975 19465 -1955
rect 19115 -1980 19120 -1975
rect 19080 -1985 19120 -1980
rect 19460 -1980 19465 -1975
rect 19495 -1980 19500 -1950
rect 19460 -1985 19500 -1980
rect 17195 -2015 17235 -2010
rect 17195 -2045 17200 -2015
rect 17230 -2020 17235 -2015
rect 18830 -2015 18870 -2010
rect 18830 -2020 18835 -2015
rect 17230 -2040 18835 -2020
rect 17230 -2045 17235 -2040
rect 17195 -2050 17235 -2045
rect 18830 -2045 18835 -2040
rect 18865 -2045 18870 -2015
rect 18830 -2050 18870 -2045
rect 16485 -2900 16520 -2895
rect 16485 -2940 16520 -2935
rect 19080 -2900 19115 -2895
rect 19080 -2940 19115 -2935
rect 19405 -2992 19440 -2987
rect 16160 -3025 16195 -3020
rect 19405 -3032 19440 -3027
rect 16160 -3065 16195 -3060
rect 16730 -3105 16770 -3100
rect 15820 -3115 15860 -3110
rect 15960 -3111 15980 -3110
rect 15820 -3145 15825 -3115
rect 15855 -3120 15860 -3115
rect 15950 -3116 15985 -3111
rect 15855 -3140 15950 -3120
rect 15855 -3145 15860 -3140
rect 15820 -3150 15860 -3145
rect 16730 -3135 16735 -3105
rect 16765 -3110 16770 -3105
rect 17780 -3105 17820 -3100
rect 17780 -3110 17785 -3105
rect 16765 -3130 17785 -3110
rect 16765 -3135 16770 -3130
rect 16730 -3140 16770 -3135
rect 17780 -3135 17785 -3130
rect 17815 -3135 17820 -3105
rect 17780 -3140 17820 -3135
rect 18615 -3105 18655 -3100
rect 18615 -3135 18620 -3105
rect 18650 -3110 18655 -3105
rect 18830 -3105 18870 -3100
rect 18830 -3110 18835 -3105
rect 18650 -3130 18835 -3110
rect 18650 -3135 18655 -3130
rect 18615 -3140 18655 -3135
rect 18830 -3135 18835 -3130
rect 18865 -3135 18870 -3105
rect 18830 -3140 18870 -3135
rect 19610 -3116 19645 -3111
rect 15950 -3156 15985 -3151
rect 19610 -3156 19645 -3151
rect 15950 -3789 15985 -3784
rect 15950 -3829 15985 -3824
rect 19610 -3789 19645 -3784
rect 19610 -3829 19645 -3824
rect 15960 -3830 15980 -3829
rect 19620 -3830 19640 -3829
rect 16280 -3894 16315 -3889
rect 16280 -3934 16315 -3929
rect 19285 -3894 19320 -3889
rect 19285 -3934 19320 -3929
rect 16290 -3935 16310 -3934
rect 19290 -3935 19310 -3934
rect 16605 -3969 16640 -3964
rect 16605 -4009 16640 -4004
rect 18960 -3969 18995 -3964
rect 18960 -4009 18995 -4004
rect 16615 -4010 16635 -4009
rect 18965 -4010 18985 -4009
rect 16540 -4035 16580 -4030
rect 16540 -4065 16545 -4035
rect 16575 -4065 16580 -4035
rect 16540 -4070 16580 -4065
rect 15595 -4190 15635 -4185
rect 15595 -4220 15600 -4190
rect 15630 -4195 15635 -4190
rect 16280 -4190 16320 -4185
rect 16280 -4195 16285 -4190
rect 15630 -4215 16285 -4195
rect 15630 -4220 15635 -4215
rect 15595 -4225 15635 -4220
rect 16280 -4220 16285 -4215
rect 16315 -4195 16320 -4190
rect 16540 -4190 16580 -4185
rect 16540 -4195 16545 -4190
rect 16315 -4215 16545 -4195
rect 16315 -4220 16320 -4215
rect 16280 -4225 16320 -4220
rect 16540 -4220 16545 -4215
rect 16575 -4195 16580 -4190
rect 16605 -4190 16645 -4185
rect 16605 -4195 16610 -4190
rect 16575 -4215 16610 -4195
rect 16575 -4220 16580 -4215
rect 16540 -4225 16580 -4220
rect 16605 -4220 16610 -4215
rect 16640 -4220 16645 -4190
rect 16605 -4225 16645 -4220
rect 15820 -4265 15860 -4260
rect 15820 -4295 15825 -4265
rect 15855 -4270 15860 -4265
rect 17250 -4265 17300 -4255
rect 17250 -4270 17260 -4265
rect 15855 -4290 17260 -4270
rect 15855 -4295 15860 -4290
rect 15820 -4300 15860 -4295
rect 17250 -4295 17260 -4290
rect 17290 -4295 17300 -4265
rect 17250 -4305 17300 -4295
rect 17780 -4265 17820 -4260
rect 17780 -4295 17785 -4265
rect 17815 -4270 17820 -4265
rect 18955 -4265 18995 -4260
rect 18955 -4270 18960 -4265
rect 17815 -4290 18960 -4270
rect 17815 -4295 17820 -4290
rect 17780 -4300 17820 -4295
rect 18955 -4295 18960 -4290
rect 18990 -4270 18995 -4265
rect 19280 -4265 19320 -4260
rect 19280 -4270 19285 -4265
rect 18990 -4290 19285 -4270
rect 18990 -4295 18995 -4290
rect 18955 -4300 18995 -4295
rect 19280 -4295 19285 -4290
rect 19315 -4270 19320 -4265
rect 19965 -4265 20005 -4260
rect 19965 -4270 19970 -4265
rect 19315 -4290 19970 -4270
rect 19315 -4295 19320 -4290
rect 19280 -4300 19320 -4295
rect 19965 -4295 19970 -4290
rect 20000 -4295 20005 -4265
rect 19965 -4300 20005 -4295
rect 15725 -4315 15765 -4310
rect 15725 -4345 15730 -4315
rect 15760 -4320 15765 -4315
rect 16900 -4315 16950 -4305
rect 16900 -4320 16910 -4315
rect 15760 -4340 16910 -4320
rect 15760 -4345 15765 -4340
rect 15725 -4350 15765 -4345
rect 16900 -4345 16910 -4340
rect 16940 -4345 16950 -4315
rect 16900 -4355 16950 -4345
rect 18650 -4315 18700 -4305
rect 18650 -4345 18660 -4315
rect 18690 -4320 18700 -4315
rect 19730 -4315 19770 -4310
rect 19730 -4320 19735 -4315
rect 18690 -4340 19735 -4320
rect 18690 -4345 18700 -4340
rect 18650 -4355 18700 -4345
rect 19730 -4345 19735 -4340
rect 19765 -4345 19770 -4315
rect 19730 -4350 19770 -4345
rect 15950 -4360 15990 -4355
rect 15950 -4390 15955 -4360
rect 15985 -4365 15990 -4360
rect 16205 -4360 16245 -4355
rect 16205 -4365 16210 -4360
rect 15985 -4385 16210 -4365
rect 15985 -4390 15990 -4385
rect 15950 -4395 15990 -4390
rect 16205 -4390 16210 -4385
rect 16240 -4390 16245 -4360
rect 16205 -4395 16245 -4390
rect 19355 -4360 19395 -4355
rect 19355 -4390 19360 -4360
rect 19390 -4365 19395 -4360
rect 19610 -4360 19650 -4355
rect 19610 -4365 19615 -4360
rect 19390 -4385 19615 -4365
rect 19390 -4390 19395 -4385
rect 19355 -4395 19395 -4390
rect 19610 -4390 19615 -4385
rect 19645 -4390 19650 -4360
rect 19610 -4395 19650 -4390
rect 17955 -4410 17995 -4405
rect 17955 -4440 17960 -4410
rect 17990 -4415 17995 -4410
rect 20050 -4410 20090 -4405
rect 20050 -4415 20055 -4410
rect 17990 -4435 20055 -4415
rect 17990 -4440 17995 -4435
rect 17955 -4445 17995 -4440
rect 20050 -4440 20055 -4435
rect 20085 -4440 20090 -4410
rect 20050 -4445 20090 -4440
<< via2 >>
rect 20055 1320 20085 1350
rect 20055 810 20085 840
rect 20055 195 20085 225
rect 20055 -710 20085 -680
rect 19970 -1025 20000 -995
rect 19970 -1210 20000 -1180
rect 19970 -1465 20000 -1435
rect 15600 -4220 15630 -4190
rect 17260 -4295 17290 -4265
rect 19970 -4295 20000 -4265
rect 16910 -4345 16940 -4315
rect 18660 -4345 18690 -4315
rect 16210 -4390 16240 -4360
rect 19360 -4390 19390 -4360
rect 17960 -4440 17990 -4410
rect 20055 -4440 20085 -4410
<< metal3 >>
rect 15505 1545 15555 1550
rect 15505 1505 15510 1545
rect 15550 1505 15555 1545
rect 15505 1500 15555 1505
rect 20045 1545 20095 1550
rect 20045 1505 20050 1545
rect 20090 1505 20095 1545
rect 20045 1500 20095 1505
rect 15510 -6245 15550 1500
rect 15590 1460 15640 1465
rect 15590 1420 15595 1460
rect 15635 1420 15640 1460
rect 15590 1415 15640 1420
rect 19960 1460 20010 1465
rect 19960 1420 19965 1460
rect 20005 1420 20010 1460
rect 19960 1415 20010 1420
rect 15595 -4190 15635 1415
rect 15595 -4220 15600 -4190
rect 15630 -4220 15635 -4190
rect 15595 -6165 15635 -4220
rect 19965 -995 20005 1415
rect 19965 -1025 19970 -995
rect 20000 -1025 20005 -995
rect 19965 -1180 20005 -1025
rect 19965 -1210 19970 -1180
rect 20000 -1210 20005 -1180
rect 19965 -1435 20005 -1210
rect 19965 -1465 19970 -1435
rect 20000 -1465 20005 -1435
rect 17250 -4260 17300 -4255
rect 17250 -4300 17255 -4260
rect 17295 -4300 17300 -4260
rect 17250 -4305 17300 -4300
rect 19965 -4265 20005 -1465
rect 19965 -4295 19970 -4265
rect 20000 -4295 20005 -4265
rect 16900 -4310 16950 -4305
rect 16900 -4350 16905 -4310
rect 16945 -4350 16950 -4310
rect 16900 -4355 16950 -4350
rect 18650 -4310 18700 -4305
rect 18650 -4350 18655 -4310
rect 18695 -4350 18700 -4310
rect 18650 -4355 18700 -4350
rect 16205 -4360 16245 -4355
rect 16205 -4390 16210 -4360
rect 16240 -4390 16245 -4360
rect 16205 -4520 16245 -4390
rect 19355 -4360 19395 -4355
rect 19355 -4390 19360 -4360
rect 19390 -4390 19395 -4360
rect 17955 -4410 17995 -4405
rect 17955 -4440 17960 -4410
rect 17990 -4440 17995 -4410
rect 17955 -4520 17995 -4440
rect 19355 -4520 19395 -4390
rect 15760 -4615 15990 -4520
rect 16110 -4615 16340 -4520
rect 16460 -4615 16690 -4520
rect 16810 -4615 17040 -4520
rect 15760 -4665 17040 -4615
rect 15760 -4750 15990 -4665
rect 16110 -4750 16340 -4665
rect 16460 -4750 16690 -4665
rect 16810 -4750 17040 -4665
rect 17160 -4615 17390 -4520
rect 17510 -4615 17740 -4520
rect 17860 -4615 18090 -4520
rect 18210 -4615 18440 -4520
rect 17160 -4665 18440 -4615
rect 17160 -4750 17390 -4665
rect 17510 -4750 17740 -4665
rect 17860 -4750 18090 -4665
rect 18210 -4750 18440 -4665
rect 18560 -4615 18790 -4520
rect 18910 -4615 19140 -4520
rect 19260 -4615 19490 -4520
rect 19610 -4615 19840 -4520
rect 18560 -4665 19840 -4615
rect 18560 -4750 18790 -4665
rect 18910 -4750 19140 -4665
rect 19260 -4750 19490 -4665
rect 19610 -4750 19840 -4665
rect 16200 -4870 16250 -4750
rect 17950 -4870 18000 -4750
rect 19350 -4870 19400 -4750
rect 15760 -4965 15990 -4870
rect 16110 -4965 16340 -4870
rect 16460 -4965 16690 -4870
rect 16810 -4965 17040 -4870
rect 15760 -5015 17040 -4965
rect 15760 -5100 15990 -5015
rect 16110 -5100 16340 -5015
rect 16460 -5100 16690 -5015
rect 16810 -5100 17040 -5015
rect 17160 -4965 17390 -4870
rect 17510 -4965 17740 -4870
rect 17860 -4965 18090 -4870
rect 18210 -4965 18440 -4870
rect 17160 -5015 18440 -4965
rect 17160 -5100 17390 -5015
rect 17510 -5100 17740 -5015
rect 17860 -5100 18090 -5015
rect 18210 -5100 18440 -5015
rect 18560 -4965 18790 -4870
rect 18910 -4965 19140 -4870
rect 19260 -4965 19490 -4870
rect 19610 -4965 19840 -4870
rect 18560 -5015 19840 -4965
rect 18560 -5100 18790 -5015
rect 18910 -5100 19140 -5015
rect 19260 -5100 19490 -5015
rect 19610 -5100 19840 -5015
rect 16200 -5220 16250 -5100
rect 17950 -5220 18000 -5100
rect 19350 -5220 19400 -5100
rect 15760 -5315 15990 -5220
rect 16110 -5315 16340 -5220
rect 16460 -5315 16690 -5220
rect 16810 -5315 17040 -5220
rect 15760 -5365 17040 -5315
rect 15760 -5450 15990 -5365
rect 16110 -5450 16340 -5365
rect 16460 -5450 16690 -5365
rect 16810 -5450 17040 -5365
rect 17160 -5315 17390 -5220
rect 17510 -5315 17740 -5220
rect 17860 -5315 18090 -5220
rect 18210 -5315 18440 -5220
rect 17160 -5365 18440 -5315
rect 17160 -5450 17390 -5365
rect 17510 -5450 17740 -5365
rect 17860 -5450 18090 -5365
rect 18210 -5450 18440 -5365
rect 18560 -5315 18790 -5220
rect 18910 -5315 19140 -5220
rect 19260 -5315 19490 -5220
rect 19610 -5315 19840 -5220
rect 18560 -5365 19840 -5315
rect 18560 -5450 18790 -5365
rect 18910 -5450 19140 -5365
rect 19260 -5450 19490 -5365
rect 19610 -5450 19840 -5365
rect 16200 -5570 16250 -5450
rect 17950 -5570 18000 -5450
rect 19350 -5570 19400 -5450
rect 15760 -5665 15990 -5570
rect 16110 -5665 16340 -5570
rect 16460 -5665 16690 -5570
rect 16810 -5665 17040 -5570
rect 15760 -5715 17040 -5665
rect 15760 -5800 15990 -5715
rect 16110 -5800 16340 -5715
rect 16460 -5800 16690 -5715
rect 16810 -5800 17040 -5715
rect 17160 -5665 17390 -5570
rect 17510 -5665 17740 -5570
rect 17860 -5665 18090 -5570
rect 18210 -5665 18440 -5570
rect 17160 -5715 18440 -5665
rect 17160 -5800 17390 -5715
rect 17510 -5800 17740 -5715
rect 17860 -5800 18090 -5715
rect 18210 -5800 18440 -5715
rect 18560 -5665 18790 -5570
rect 18910 -5665 19140 -5570
rect 19260 -5665 19490 -5570
rect 19610 -5665 19840 -5570
rect 18560 -5715 19840 -5665
rect 18560 -5800 18790 -5715
rect 18910 -5800 19140 -5715
rect 19260 -5800 19490 -5715
rect 19610 -5800 19840 -5715
rect 16200 -5920 16250 -5800
rect 17950 -5920 18000 -5800
rect 19350 -5920 19400 -5800
rect 15760 -6015 15990 -5920
rect 16110 -6015 16340 -5920
rect 16460 -6015 16690 -5920
rect 16810 -6015 17040 -5920
rect 15760 -6065 17040 -6015
rect 15760 -6150 15990 -6065
rect 16110 -6150 16340 -6065
rect 16460 -6150 16690 -6065
rect 16810 -6150 17040 -6065
rect 17160 -6015 17390 -5920
rect 17510 -6015 17740 -5920
rect 17860 -6015 18090 -5920
rect 18210 -6015 18440 -5920
rect 17160 -6065 18440 -6015
rect 17160 -6150 17390 -6065
rect 17510 -6150 17740 -6065
rect 17860 -6150 18090 -6065
rect 18210 -6150 18440 -6065
rect 18560 -6015 18790 -5920
rect 18910 -6015 19140 -5920
rect 19260 -6015 19490 -5920
rect 19610 -6015 19840 -5920
rect 18560 -6065 19840 -6015
rect 18560 -6150 18790 -6065
rect 18910 -6150 19140 -6065
rect 19260 -6150 19490 -6065
rect 19610 -6150 19840 -6065
rect 19965 -6165 20005 -4295
rect 20050 1350 20090 1500
rect 20050 1320 20055 1350
rect 20085 1320 20090 1350
rect 20050 840 20090 1320
rect 20050 810 20055 840
rect 20085 810 20090 840
rect 20050 225 20090 810
rect 20050 195 20055 225
rect 20085 195 20090 225
rect 20050 -680 20090 195
rect 20050 -710 20055 -680
rect 20085 -710 20090 -680
rect 20050 -4410 20090 -710
rect 20050 -4440 20055 -4410
rect 20085 -4440 20090 -4410
rect 15590 -6170 15640 -6165
rect 15590 -6210 15595 -6170
rect 15635 -6210 15640 -6170
rect 15590 -6215 15640 -6210
rect 19960 -6170 20010 -6165
rect 19960 -6210 19965 -6170
rect 20005 -6210 20010 -6170
rect 19960 -6215 20010 -6210
rect 20050 -6245 20090 -4440
rect 15505 -6250 15555 -6245
rect 15505 -6290 15510 -6250
rect 15550 -6290 15555 -6250
rect 15505 -6295 15555 -6290
rect 20045 -6250 20095 -6245
rect 20045 -6290 20050 -6250
rect 20090 -6290 20095 -6250
rect 20045 -6295 20095 -6290
<< via3 >>
rect 15510 1505 15550 1545
rect 20050 1505 20090 1545
rect 15595 1420 15635 1460
rect 19965 1420 20005 1460
rect 17255 -4265 17295 -4260
rect 17255 -4295 17260 -4265
rect 17260 -4295 17290 -4265
rect 17290 -4295 17295 -4265
rect 17255 -4300 17295 -4295
rect 16905 -4315 16945 -4310
rect 16905 -4345 16910 -4315
rect 16910 -4345 16940 -4315
rect 16940 -4345 16945 -4315
rect 16905 -4350 16945 -4345
rect 18655 -4315 18695 -4310
rect 18655 -4345 18660 -4315
rect 18660 -4345 18690 -4315
rect 18690 -4345 18695 -4315
rect 18655 -4350 18695 -4345
rect 15595 -6210 15635 -6170
rect 19965 -6210 20005 -6170
rect 15510 -6290 15550 -6250
rect 20050 -6290 20090 -6250
<< mimcap >>
rect 15775 -4620 15975 -4535
rect 15775 -4660 15855 -4620
rect 15895 -4660 15975 -4620
rect 15775 -4735 15975 -4660
rect 16125 -4620 16325 -4535
rect 16125 -4660 16205 -4620
rect 16245 -4660 16325 -4620
rect 16125 -4735 16325 -4660
rect 16475 -4620 16675 -4535
rect 16475 -4660 16555 -4620
rect 16595 -4660 16675 -4620
rect 16475 -4735 16675 -4660
rect 16825 -4620 17025 -4535
rect 16825 -4660 16905 -4620
rect 16945 -4660 17025 -4620
rect 16825 -4735 17025 -4660
rect 17175 -4620 17375 -4535
rect 17175 -4660 17255 -4620
rect 17295 -4660 17375 -4620
rect 17175 -4735 17375 -4660
rect 17525 -4620 17725 -4535
rect 17525 -4660 17605 -4620
rect 17645 -4660 17725 -4620
rect 17525 -4735 17725 -4660
rect 17875 -4620 18075 -4535
rect 17875 -4660 17955 -4620
rect 17995 -4660 18075 -4620
rect 17875 -4735 18075 -4660
rect 18225 -4620 18425 -4535
rect 18225 -4660 18305 -4620
rect 18345 -4660 18425 -4620
rect 18225 -4735 18425 -4660
rect 18575 -4620 18775 -4535
rect 18575 -4660 18655 -4620
rect 18695 -4660 18775 -4620
rect 18575 -4735 18775 -4660
rect 18925 -4620 19125 -4535
rect 18925 -4660 19005 -4620
rect 19045 -4660 19125 -4620
rect 18925 -4735 19125 -4660
rect 19275 -4620 19475 -4535
rect 19275 -4660 19355 -4620
rect 19395 -4660 19475 -4620
rect 19275 -4735 19475 -4660
rect 19625 -4620 19825 -4535
rect 19625 -4660 19705 -4620
rect 19745 -4660 19825 -4620
rect 19625 -4735 19825 -4660
rect 15775 -4970 15975 -4885
rect 15775 -5010 15855 -4970
rect 15895 -5010 15975 -4970
rect 15775 -5085 15975 -5010
rect 16125 -4970 16325 -4885
rect 16125 -5010 16205 -4970
rect 16245 -5010 16325 -4970
rect 16125 -5085 16325 -5010
rect 16475 -4970 16675 -4885
rect 16475 -5010 16555 -4970
rect 16595 -5010 16675 -4970
rect 16475 -5085 16675 -5010
rect 16825 -4970 17025 -4885
rect 16825 -5010 16905 -4970
rect 16945 -5010 17025 -4970
rect 16825 -5085 17025 -5010
rect 17175 -4970 17375 -4885
rect 17175 -5010 17255 -4970
rect 17295 -5010 17375 -4970
rect 17175 -5085 17375 -5010
rect 17525 -4970 17725 -4885
rect 17525 -5010 17605 -4970
rect 17645 -5010 17725 -4970
rect 17525 -5085 17725 -5010
rect 17875 -4970 18075 -4885
rect 17875 -5010 17955 -4970
rect 17995 -5010 18075 -4970
rect 17875 -5085 18075 -5010
rect 18225 -4970 18425 -4885
rect 18225 -5010 18305 -4970
rect 18345 -5010 18425 -4970
rect 18225 -5085 18425 -5010
rect 18575 -4970 18775 -4885
rect 18575 -5010 18655 -4970
rect 18695 -5010 18775 -4970
rect 18575 -5085 18775 -5010
rect 18925 -4970 19125 -4885
rect 18925 -5010 19005 -4970
rect 19045 -5010 19125 -4970
rect 18925 -5085 19125 -5010
rect 19275 -4970 19475 -4885
rect 19275 -5010 19355 -4970
rect 19395 -5010 19475 -4970
rect 19275 -5085 19475 -5010
rect 19625 -4970 19825 -4885
rect 19625 -5010 19705 -4970
rect 19745 -5010 19825 -4970
rect 19625 -5085 19825 -5010
rect 15775 -5320 15975 -5235
rect 15775 -5360 15855 -5320
rect 15895 -5360 15975 -5320
rect 15775 -5435 15975 -5360
rect 16125 -5320 16325 -5235
rect 16125 -5360 16205 -5320
rect 16245 -5360 16325 -5320
rect 16125 -5435 16325 -5360
rect 16475 -5320 16675 -5235
rect 16475 -5360 16555 -5320
rect 16595 -5360 16675 -5320
rect 16475 -5435 16675 -5360
rect 16825 -5320 17025 -5235
rect 16825 -5360 16905 -5320
rect 16945 -5360 17025 -5320
rect 16825 -5435 17025 -5360
rect 17175 -5320 17375 -5235
rect 17175 -5360 17255 -5320
rect 17295 -5360 17375 -5320
rect 17175 -5435 17375 -5360
rect 17525 -5320 17725 -5235
rect 17525 -5360 17605 -5320
rect 17645 -5360 17725 -5320
rect 17525 -5435 17725 -5360
rect 17875 -5320 18075 -5235
rect 17875 -5360 17955 -5320
rect 17995 -5360 18075 -5320
rect 17875 -5435 18075 -5360
rect 18225 -5320 18425 -5235
rect 18225 -5360 18305 -5320
rect 18345 -5360 18425 -5320
rect 18225 -5435 18425 -5360
rect 18575 -5320 18775 -5235
rect 18575 -5360 18655 -5320
rect 18695 -5360 18775 -5320
rect 18575 -5435 18775 -5360
rect 18925 -5320 19125 -5235
rect 18925 -5360 19005 -5320
rect 19045 -5360 19125 -5320
rect 18925 -5435 19125 -5360
rect 19275 -5320 19475 -5235
rect 19275 -5360 19355 -5320
rect 19395 -5360 19475 -5320
rect 19275 -5435 19475 -5360
rect 19625 -5320 19825 -5235
rect 19625 -5360 19705 -5320
rect 19745 -5360 19825 -5320
rect 19625 -5435 19825 -5360
rect 15775 -5670 15975 -5585
rect 15775 -5710 15855 -5670
rect 15895 -5710 15975 -5670
rect 15775 -5785 15975 -5710
rect 16125 -5670 16325 -5585
rect 16125 -5710 16205 -5670
rect 16245 -5710 16325 -5670
rect 16125 -5785 16325 -5710
rect 16475 -5670 16675 -5585
rect 16475 -5710 16555 -5670
rect 16595 -5710 16675 -5670
rect 16475 -5785 16675 -5710
rect 16825 -5670 17025 -5585
rect 16825 -5710 16905 -5670
rect 16945 -5710 17025 -5670
rect 16825 -5785 17025 -5710
rect 17175 -5670 17375 -5585
rect 17175 -5710 17255 -5670
rect 17295 -5710 17375 -5670
rect 17175 -5785 17375 -5710
rect 17525 -5670 17725 -5585
rect 17525 -5710 17605 -5670
rect 17645 -5710 17725 -5670
rect 17525 -5785 17725 -5710
rect 17875 -5670 18075 -5585
rect 17875 -5710 17955 -5670
rect 17995 -5710 18075 -5670
rect 17875 -5785 18075 -5710
rect 18225 -5670 18425 -5585
rect 18225 -5710 18305 -5670
rect 18345 -5710 18425 -5670
rect 18225 -5785 18425 -5710
rect 18575 -5670 18775 -5585
rect 18575 -5710 18655 -5670
rect 18695 -5710 18775 -5670
rect 18575 -5785 18775 -5710
rect 18925 -5670 19125 -5585
rect 18925 -5710 19005 -5670
rect 19045 -5710 19125 -5670
rect 18925 -5785 19125 -5710
rect 19275 -5670 19475 -5585
rect 19275 -5710 19355 -5670
rect 19395 -5710 19475 -5670
rect 19275 -5785 19475 -5710
rect 19625 -5670 19825 -5585
rect 19625 -5710 19705 -5670
rect 19745 -5710 19825 -5670
rect 19625 -5785 19825 -5710
rect 15775 -6020 15975 -5935
rect 15775 -6060 15855 -6020
rect 15895 -6060 15975 -6020
rect 15775 -6135 15975 -6060
rect 16125 -6020 16325 -5935
rect 16125 -6060 16205 -6020
rect 16245 -6060 16325 -6020
rect 16125 -6135 16325 -6060
rect 16475 -6020 16675 -5935
rect 16475 -6060 16555 -6020
rect 16595 -6060 16675 -6020
rect 16475 -6135 16675 -6060
rect 16825 -6020 17025 -5935
rect 16825 -6060 16905 -6020
rect 16945 -6060 17025 -6020
rect 16825 -6135 17025 -6060
rect 17175 -6020 17375 -5935
rect 17175 -6060 17255 -6020
rect 17295 -6060 17375 -6020
rect 17175 -6135 17375 -6060
rect 17525 -6020 17725 -5935
rect 17525 -6060 17605 -6020
rect 17645 -6060 17725 -6020
rect 17525 -6135 17725 -6060
rect 17875 -6020 18075 -5935
rect 17875 -6060 17955 -6020
rect 17995 -6060 18075 -6020
rect 17875 -6135 18075 -6060
rect 18225 -6020 18425 -5935
rect 18225 -6060 18305 -6020
rect 18345 -6060 18425 -6020
rect 18225 -6135 18425 -6060
rect 18575 -6020 18775 -5935
rect 18575 -6060 18655 -6020
rect 18695 -6060 18775 -6020
rect 18575 -6135 18775 -6060
rect 18925 -6020 19125 -5935
rect 18925 -6060 19005 -6020
rect 19045 -6060 19125 -6020
rect 18925 -6135 19125 -6060
rect 19275 -6020 19475 -5935
rect 19275 -6060 19355 -6020
rect 19395 -6060 19475 -6020
rect 19275 -6135 19475 -6060
rect 19625 -6020 19825 -5935
rect 19625 -6060 19705 -6020
rect 19745 -6060 19825 -6020
rect 19625 -6135 19825 -6060
<< mimcapcontact >>
rect 15855 -4660 15895 -4620
rect 16205 -4660 16245 -4620
rect 16555 -4660 16595 -4620
rect 16905 -4660 16945 -4620
rect 17255 -4660 17295 -4620
rect 17605 -4660 17645 -4620
rect 17955 -4660 17995 -4620
rect 18305 -4660 18345 -4620
rect 18655 -4660 18695 -4620
rect 19005 -4660 19045 -4620
rect 19355 -4660 19395 -4620
rect 19705 -4660 19745 -4620
rect 15855 -5010 15895 -4970
rect 16205 -5010 16245 -4970
rect 16555 -5010 16595 -4970
rect 16905 -5010 16945 -4970
rect 17255 -5010 17295 -4970
rect 17605 -5010 17645 -4970
rect 17955 -5010 17995 -4970
rect 18305 -5010 18345 -4970
rect 18655 -5010 18695 -4970
rect 19005 -5010 19045 -4970
rect 19355 -5010 19395 -4970
rect 19705 -5010 19745 -4970
rect 15855 -5360 15895 -5320
rect 16205 -5360 16245 -5320
rect 16555 -5360 16595 -5320
rect 16905 -5360 16945 -5320
rect 17255 -5360 17295 -5320
rect 17605 -5360 17645 -5320
rect 17955 -5360 17995 -5320
rect 18305 -5360 18345 -5320
rect 18655 -5360 18695 -5320
rect 19005 -5360 19045 -5320
rect 19355 -5360 19395 -5320
rect 19705 -5360 19745 -5320
rect 15855 -5710 15895 -5670
rect 16205 -5710 16245 -5670
rect 16555 -5710 16595 -5670
rect 16905 -5710 16945 -5670
rect 17255 -5710 17295 -5670
rect 17605 -5710 17645 -5670
rect 17955 -5710 17995 -5670
rect 18305 -5710 18345 -5670
rect 18655 -5710 18695 -5670
rect 19005 -5710 19045 -5670
rect 19355 -5710 19395 -5670
rect 19705 -5710 19745 -5670
rect 15855 -6060 15895 -6020
rect 16205 -6060 16245 -6020
rect 16555 -6060 16595 -6020
rect 16905 -6060 16945 -6020
rect 17255 -6060 17295 -6020
rect 17605 -6060 17645 -6020
rect 17955 -6060 17995 -6020
rect 18305 -6060 18345 -6020
rect 18655 -6060 18695 -6020
rect 19005 -6060 19045 -6020
rect 19355 -6060 19395 -6020
rect 19705 -6060 19745 -6020
<< metal4 >>
rect 15505 1545 20095 1550
rect 15505 1505 15510 1545
rect 15550 1505 20050 1545
rect 20090 1505 20095 1545
rect 15505 1500 20095 1505
rect 15590 1460 20010 1465
rect 15590 1420 15595 1460
rect 15635 1420 19965 1460
rect 20005 1420 20010 1460
rect 15590 1415 20010 1420
rect 17250 -4260 17300 -4255
rect 17250 -4300 17255 -4260
rect 17295 -4300 17300 -4260
rect 16900 -4310 16950 -4305
rect 16900 -4350 16905 -4310
rect 16945 -4350 16950 -4310
rect 16900 -4615 16950 -4350
rect 15850 -4620 16950 -4615
rect 15850 -4660 15855 -4620
rect 15895 -4660 16205 -4620
rect 16245 -4660 16555 -4620
rect 16595 -4660 16905 -4620
rect 16945 -4660 16950 -4620
rect 15850 -4665 16950 -4660
rect 17250 -4615 17300 -4300
rect 18650 -4310 18700 -4305
rect 18650 -4350 18655 -4310
rect 18695 -4350 18700 -4310
rect 18650 -4615 18700 -4350
rect 17250 -4620 18350 -4615
rect 17250 -4660 17255 -4620
rect 17295 -4660 17605 -4620
rect 17645 -4660 17955 -4620
rect 17995 -4660 18305 -4620
rect 18345 -4660 18350 -4620
rect 17250 -4665 18350 -4660
rect 18650 -4620 19750 -4615
rect 18650 -4660 18655 -4620
rect 18695 -4660 19005 -4620
rect 19045 -4660 19355 -4620
rect 19395 -4660 19705 -4620
rect 19745 -4660 19750 -4620
rect 18650 -4665 19750 -4660
rect 16200 -4965 16250 -4665
rect 17950 -4965 18000 -4665
rect 19350 -4965 19400 -4665
rect 15850 -4970 16950 -4965
rect 15850 -5010 15855 -4970
rect 15895 -5010 16205 -4970
rect 16245 -5010 16555 -4970
rect 16595 -5010 16905 -4970
rect 16945 -5010 16950 -4970
rect 15850 -5015 16950 -5010
rect 17250 -4970 18350 -4965
rect 17250 -5010 17255 -4970
rect 17295 -5010 17605 -4970
rect 17645 -5010 17955 -4970
rect 17995 -5010 18305 -4970
rect 18345 -5010 18350 -4970
rect 17250 -5015 18350 -5010
rect 18650 -4970 19750 -4965
rect 18650 -5010 18655 -4970
rect 18695 -5010 19005 -4970
rect 19045 -5010 19355 -4970
rect 19395 -5010 19705 -4970
rect 19745 -5010 19750 -4970
rect 18650 -5015 19750 -5010
rect 16200 -5315 16250 -5015
rect 17950 -5315 18000 -5015
rect 19350 -5315 19400 -5015
rect 15850 -5320 16950 -5315
rect 15850 -5360 15855 -5320
rect 15895 -5360 16205 -5320
rect 16245 -5360 16555 -5320
rect 16595 -5360 16905 -5320
rect 16945 -5360 16950 -5320
rect 15850 -5365 16950 -5360
rect 17250 -5320 18350 -5315
rect 17250 -5360 17255 -5320
rect 17295 -5360 17605 -5320
rect 17645 -5360 17955 -5320
rect 17995 -5360 18305 -5320
rect 18345 -5360 18350 -5320
rect 17250 -5365 18350 -5360
rect 18650 -5320 19750 -5315
rect 18650 -5360 18655 -5320
rect 18695 -5360 19005 -5320
rect 19045 -5360 19355 -5320
rect 19395 -5360 19705 -5320
rect 19745 -5360 19750 -5320
rect 18650 -5365 19750 -5360
rect 16200 -5665 16250 -5365
rect 17950 -5665 18000 -5365
rect 19350 -5665 19400 -5365
rect 15850 -5670 16950 -5665
rect 15850 -5710 15855 -5670
rect 15895 -5710 16205 -5670
rect 16245 -5710 16555 -5670
rect 16595 -5710 16905 -5670
rect 16945 -5710 16950 -5670
rect 15850 -5715 16950 -5710
rect 17250 -5670 18350 -5665
rect 17250 -5710 17255 -5670
rect 17295 -5710 17605 -5670
rect 17645 -5710 17955 -5670
rect 17995 -5710 18305 -5670
rect 18345 -5710 18350 -5670
rect 17250 -5715 18350 -5710
rect 18650 -5670 19750 -5665
rect 18650 -5710 18655 -5670
rect 18695 -5710 19005 -5670
rect 19045 -5710 19355 -5670
rect 19395 -5710 19705 -5670
rect 19745 -5710 19750 -5670
rect 18650 -5715 19750 -5710
rect 16200 -6015 16250 -5715
rect 17950 -6015 18000 -5715
rect 19350 -6015 19400 -5715
rect 15850 -6020 16950 -6015
rect 15850 -6060 15855 -6020
rect 15895 -6060 16205 -6020
rect 16245 -6060 16555 -6020
rect 16595 -6060 16905 -6020
rect 16945 -6060 16950 -6020
rect 15850 -6065 16950 -6060
rect 17250 -6020 18350 -6015
rect 17250 -6060 17255 -6020
rect 17295 -6060 17605 -6020
rect 17645 -6060 17955 -6020
rect 17995 -6060 18305 -6020
rect 18345 -6060 18350 -6020
rect 17250 -6065 18350 -6060
rect 18650 -6020 19750 -6015
rect 18650 -6060 18655 -6020
rect 18695 -6060 19005 -6020
rect 19045 -6060 19355 -6020
rect 19395 -6060 19705 -6020
rect 19745 -6060 19750 -6020
rect 18650 -6065 19750 -6060
rect 15590 -6170 20010 -6165
rect 15590 -6210 15595 -6170
rect 15635 -6210 19965 -6170
rect 20005 -6210 20010 -6170
rect 15590 -6215 20010 -6210
rect 15505 -6250 20095 -6245
rect 15505 -6290 15510 -6250
rect 15550 -6290 20050 -6250
rect 20090 -6290 20095 -6250
rect 15505 -6295 20095 -6290
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 18145 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_18
timestamp 1723858470
transform 1 0 16785 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_19
timestamp 1723858470
transform 1 0 17465 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_20
timestamp 1723858470
transform 1 0 18145 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_21
timestamp 1723858470
transform 1 0 18145 0 1 -3455
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_22
timestamp 1723858470
transform 1 0 17465 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23
timestamp 1723858470
transform 1 0 17465 0 1 -3455
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_24
timestamp 1723858470
transform 1 0 16785 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25
timestamp 1723858470
transform 1 0 16785 0 1 -3455
box 0 0 670 670
<< labels >>
flabel metal2 15995 -4385 15995 -4385 5 FreeSans 400 0 0 -40 cap_res1
flabel metal3 19355 -4375 19355 -4375 7 FreeSans 400 180 -40 0 cap_res2
flabel metal1 16125 1595 16125 1595 1 FreeSans 240 0 0 80 ERR_AMP_CUR_BIAS
port 7 n
flabel metal1 19280 1595 19280 1595 1 FreeSans 240 0 0 80 VB1_CUR_BIAS
port 4 n
flabel metal1 19795 1595 19795 1595 1 FreeSans 240 0 0 80 V_CMFB_S4
port 9 n
flabel metal1 16040 1585 16040 1585 7 FreeSans 240 0 -160 0 VB2_CUR_BIAS
port 11 w
flabel metal1 19415 1590 19415 1590 7 FreeSans 240 0 -160 0 ERR_AMP_REF
port 2 w
flabel metal1 19565 1590 19565 1590 3 FreeSans 240 0 160 0 VB3_CUR_BIAS
port 8 e
flabel metal1 15805 1595 15805 1595 1 FreeSans 240 0 0 80 V_CMFB_S2
port 10 n
flabel metal1 17750 1595 17750 1595 1 FreeSans 240 0 0 80 TAIL_CUR_MIR_BIAS
port 5 n
flabel metal1 17105 1595 17105 1595 1 FreeSans 240 0 0 80 V_CMFB_S1
port 6 n
flabel metal1 18495 1595 18495 1595 1 FreeSans 240 0 0 80 V_CMFB_S3
port 3 n
flabel metal3 20090 1220 20090 1220 3 FreeSans 400 0 200 0 VDDA
port 1 e
flabel metal2 16620 -105 16620 -105 5 FreeSans 400 0 0 -40 V_mir1
flabel metal1 16190 -1370 16190 -1370 3 FreeSans 400 0 40 0 NFET_GATE_10uA
flabel metal3 20005 920 20005 920 3 FreeSans 400 0 200 0 GNDA
port 12 e
flabel poly 18430 480 18430 480 5 FreeSans 400 0 0 -40 V_TOP
flabel metal1 16235 -945 16235 -945 3 FreeSans 400 0 200 0 START_UP
flabel metal2 17430 -630 17430 -630 3 FreeSans 400 0 200 0 V_p_1
flabel metal2 16670 -535 16670 -535 1 FreeSans 400 0 0 80 Vin+
flabel metal2 16665 -415 16665 -415 5 FreeSans 400 0 0 -80 Vin-
flabel metal2 18930 -535 18930 -535 1 FreeSans 400 0 0 80 V_CUR_REF_REG
flabel metal1 18340 -1110 18340 -1110 3 FreeSans 400 0 200 0 START_UP_NFET1
flabel metal1 18170 -630 18170 -630 7 FreeSans 400 0 -160 0 V_p_2
flabel metal1 17525 -255 17525 -255 5 FreeSans 400 0 0 -160 1st_Vout_1
flabel metal1 18075 -255 18075 -255 5 FreeSans 400 0 0 -160 1st_Vout_2
flabel metal1 18980 -105 18980 -105 5 FreeSans 400 0 0 -160 V_mir2
flabel metal1 18760 1080 18760 1080 3 FreeSans 400 0 160 0 PFET_GATE_10uA
<< end >>
