magic
tech sky130A
timestamp 1740284885
<< nwell >>
rect 1140 635 1245 675
rect 1135 530 1245 635
<< poly >>
rect 1175 520 1240 535
rect 150 260 170 275
<< locali >>
rect 1185 1140 1235 1150
rect 0 1120 25 1140
rect 1170 1120 1195 1140
rect 1185 1110 1195 1120
rect 1225 1110 1235 1140
rect 1185 1100 1235 1110
rect 1185 750 1235 760
rect 1185 720 1195 750
rect 1225 720 1235 750
rect 1185 710 1235 720
rect 6460 530 6470 550
rect 1185 350 1235 360
rect 1185 320 1195 350
rect 1225 320 1235 350
rect 1185 310 1235 320
rect 1185 100 1235 110
rect 1185 90 1195 100
rect 0 70 20 90
rect 1170 70 1195 90
rect 1225 70 1235 100
rect 1185 60 1235 70
<< viali >>
rect 1195 1110 1225 1140
rect 1195 720 1225 750
rect 1195 320 1225 350
rect 1195 70 1225 100
<< metal1 >>
rect 0 1140 20 1150
rect 1170 1140 1235 1150
rect 0 1120 25 1140
rect 0 1110 20 1120
rect 1170 1110 1195 1140
rect 1225 1110 1235 1140
rect 1185 1100 1235 1110
rect 1185 750 1235 760
rect 1185 720 1195 750
rect 1225 720 1235 750
rect 1185 710 1235 720
rect 1185 350 1235 360
rect 1185 320 1195 350
rect 1225 320 1235 350
rect 1185 310 1235 320
rect 1185 100 1235 110
rect 0 60 20 100
rect 1175 90 1195 100
rect 1170 70 1195 90
rect 1225 70 1235 100
rect 1175 60 1235 70
<< via1 >>
rect 1195 1110 1225 1140
rect 1195 720 1225 750
rect 1195 320 1225 350
rect 1195 70 1225 100
<< metal2 >>
rect 1185 1140 1235 1150
rect 1185 1110 1195 1140
rect 1225 1110 1235 1140
rect 1185 1100 1235 1110
rect 1185 750 1235 760
rect 1185 720 1195 750
rect 1225 720 1235 750
rect 1185 710 1235 720
rect 1185 350 1235 360
rect 1185 320 1195 350
rect 1225 320 1235 350
rect 1185 310 1235 320
rect 1185 100 1235 110
rect 1185 70 1195 100
rect 1225 70 1235 100
rect 1185 60 1235 70
<< via2 >>
rect 1195 1110 1225 1140
rect 1195 720 1225 750
rect 1195 320 1225 350
rect 1195 70 1225 100
<< metal3 >>
rect 1185 1145 1235 1150
rect 1185 1105 1190 1145
rect 1230 1105 1235 1145
rect 1185 1100 1235 1105
rect 1185 755 1235 760
rect 1185 715 1190 755
rect 1230 715 1235 755
rect 1185 710 1235 715
rect 1185 355 1235 360
rect 1185 315 1190 355
rect 1230 315 1235 355
rect 1185 310 1235 315
rect 1185 105 1235 110
rect 1185 65 1190 105
rect 1230 65 1235 105
rect 1185 60 1235 65
<< via3 >>
rect 1190 1140 1230 1145
rect 1190 1110 1195 1140
rect 1195 1110 1225 1140
rect 1225 1110 1230 1140
rect 1190 1105 1230 1110
rect 1190 750 1230 755
rect 1190 720 1195 750
rect 1195 720 1225 750
rect 1225 720 1230 750
rect 1190 715 1230 720
rect 1190 350 1230 355
rect 1190 320 1195 350
rect 1195 320 1225 350
rect 1225 320 1230 350
rect 1190 315 1230 320
rect 1190 100 1230 105
rect 1190 70 1195 100
rect 1195 70 1225 100
rect 1225 70 1230 100
rect 1190 65 1230 70
<< metal4 >>
rect 1185 1145 1235 1150
rect 1185 1105 1190 1145
rect 1230 1105 1235 1145
rect 1185 755 1235 1105
rect 1185 715 1190 755
rect 1230 715 1235 755
rect 1185 710 1235 715
rect 1185 355 1235 360
rect 1185 315 1190 355
rect 1230 315 1235 355
rect 1185 105 1235 315
rect 1185 65 1190 105
rect 1230 65 1235 105
rect 1185 60 1235 65
use div120_2  div120_2_0
timestamp 1740045839
transform 1 0 1245 0 1 890
box -10 -570 5215 -140
use vco2_3  vco2_3_0
timestamp 1740284794
transform 1 0 -1175 0 1 525
box 1175 -465 2350 625
<< labels >>
flabel metal1 0 1130 0 1130 7 FreeSans 800 0 -400 0 VDDA
port 2 w
flabel metal1 0 80 0 80 7 FreeSans 800 0 -400 0 GNDA
port 3 w
flabel poly 1205 520 1205 520 5 FreeSans 800 0 0 -400 V_OSC
flabel locali 6470 540 6470 540 3 FreeSans 800 0 400 0 V_OUT_120
port 1 e
flabel poly 150 270 150 270 7 FreeSans 800 0 -400 0 V_CONT
port 4 w
<< end >>
