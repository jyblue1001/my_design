* NGSPICE file created from charge_pump_2.ext - technology: sky130A

.subckt charge_pump_8 w_n3090_1240# a_n2950_2110# a_n2790_310# a_n3050_2170# a_n1130_2170#
X0 a_n3050_2170# a_n2950_2110# w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X1 a_n1130_2170# a_n1700_820# w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X2 a_n2790_310# a_n540_820# a_n1130_2170# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X3 w_n3090_1240# a_n1700_820# a_n1130_2170# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X4 w_n3090_1240# a_n2950_2110# a_n3050_2170# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X5 a_n1120_820# w_n3090_1240# a_n1540_820# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X6 a_n540_820# a_n1120_820# a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X7 a_n1120_820# a_n2790_310# a_n1540_820# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X8 a_n3050_2170# a_n3010_310# a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X9 a_n3050_2170# a_n2950_2110# w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X10 a_n3050_2170# a_n2950_2110# w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X11 a_n1990_820# a_n2280_820# w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X12 a_n3010_310# a_n3010_310# a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X13 a_n1130_2170# a_n540_820# a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X14 w_n3090_1240# a_n2950_2110# a_n3050_2170# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X15 a_n1700_820# a_n1990_820# a_n2950_2110# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X16 a_n2280_820# a_n2570_820# a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X17 a_n2790_310# a_n3010_310# a_n3010_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X18 a_n2790_310# a_n3010_310# a_n3010_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X19 a_n1700_820# a_n2280_820# w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X20 a_n2570_820# a_n3330_1140# a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X21 a_n1130_2170# a_n1700_820# w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X22 a_n3010_310# a_n3010_310# a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X23 a_n2790_310# a_n3330_710# a_n1540_820# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X24 a_n540_820# a_n830_820# a_n3010_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X25 a_n1130_2170# a_n1700_820# w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X26 a_n830_820# a_n1120_820# w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X27 w_n3090_1240# a_n1700_820# a_n1130_2170# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X28 a_n1130_2170# a_n1700_820# w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X29 a_n2570_820# a_n3330_1140# w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X30 w_n3090_1240# a_n2950_2110# a_n3050_2170# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X31 w_n3090_1240# a_n3330_710# a_n1540_820# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X32 w_n3090_1240# a_n1700_820# a_n1130_2170# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X33 a_n2790_310# a_n3010_310# a_n3050_2170# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X34 a_n3050_2170# a_n2950_2110# w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X35 a_n2280_820# a_n2570_820# w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X36 a_n2790_310# a_n540_820# a_n1130_2170# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X37 a_n1700_820# a_n2280_820# a_n2950_2110# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X38 a_n830_820# a_n1120_820# a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X39 w_n3090_1240# a_n2950_2110# a_n3050_2170# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X40 a_n3050_2170# a_n3010_310# a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X41 w_n3090_1240# a_n1700_820# a_n1130_2170# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X42 a_n1990_820# a_n2280_820# a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X43 a_n1130_2170# a_n540_820# a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X44 a_n540_820# a_n1120_820# a_n3010_310# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X45 a_n2790_310# a_n3010_310# a_n3050_2170# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X46 a_n1700_820# a_n1990_820# sky130_fd_pr__cap_mim_m3_1 l=4.2 w=6
X47 a_n540_820# a_n830_820# sky130_fd_pr__cap_mim_m3_1 l=2.6 w=2.6
.ends

.subckt opamp_6_6 a_1630_200# a_3420_n350# a_1470_530# w_1980_260# a_2150_n350#
X0 a_3420_n350# a_3000_310# w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X1 w_1980_260# a_3000_310# a_3420_n350# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X2 a_3420_n350# a_2280_n350# a_2150_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X3 a_3420_n350# a_4140_1066# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X4 a_2020_310# a_1980_n1180# w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X5 a_3420_n350# a_3000_310# w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X6 a_2280_n350# a_2020_n350# a_2150_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X7 w_1980_260# a_1980_n1180# a_2020_310# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X8 a_4140_1066# a_3000_310# a_2150_n350# sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X9 a_2150_n350# a_2280_n350# a_3420_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X10 a_2150_n350# a_2020_n350# a_2020_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X11 w_1980_260# a_1980_n1180# a_1980_n1180# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=1.25 ps=6 w=2.5 l=0.5
X12 a_2280_n350# a_1630_200# a_2020_310# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X13 a_2020_310# a_1470_530# a_2020_n350# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X14 a_2490_n1180# a_2490_n1180# a_2150_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=1.25 pd=6 as=0.625 ps=3 w=2.5 l=0.5
X15 w_1980_260# a_1980_n1180# a_2020_310# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X16 a_2020_n350# a_1470_530# a_2020_310# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X17 a_3420_n350# a_2280_n350# a_2150_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X18 a_1980_n1180# a_1980_n1180# w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X19 a_2020_310# a_1630_200# a_2280_n350# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X20 a_2020_n350# a_2020_n350# a_2150_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X21 a_2150_n350# a_2490_n1180# a_2740_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X22 a_2280_n350# a_4140_n1860# a_2150_n350# sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X23 a_2740_n350# a_1630_200# a_3000_310# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X24 a_2740_310# a_2740_310# w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X25 a_2020_310# a_1980_n1180# w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X26 a_3000_310# a_1630_200# a_2740_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X27 w_1980_260# a_2740_310# a_3000_310# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X28 a_2740_n350# a_2490_n1180# a_2150_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X29 a_2740_n350# a_1470_530# a_2740_310# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X30 a_3000_310# a_2740_310# w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X31 a_3420_n350# a_4140_n1860# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X32 a_1980_n1180# a_1980_n1180# w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0.625 ps=3 w=2.5 l=0.5
X33 w_1980_260# a_2740_310# a_2740_310# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X34 a_2150_n350# a_2280_n350# a_3420_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X35 a_1980_n1180# a_2490_n1180# a_2150_n350# sky130_fd_pr__res_xhigh_po_2p85 l=0.51
X36 w_1980_260# a_3000_310# a_3420_n350# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X37 w_1980_260# a_1980_n1180# a_1980_n1180# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X38 a_2150_n350# a_2020_n350# a_2280_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X39 a_2740_310# a_1470_530# a_2740_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X40 a_2150_n350# a_2490_n1180# a_2490_n1180# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=1.25 ps=6 w=2.5 l=0.5
.ends

.subckt charge_pump_2
Xcharge_pump_8_0 VDDA li_1590_1640# GNDA a_n310_5360# VOUT charge_pump_8
Xopamp_6_6_0 VOUT li_1590_1640# a_n310_5360# VDDA GNDA opamp_6_6
.ends

