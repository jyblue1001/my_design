magic
tech sky130A
timestamp 1737692480
<< nwell >>
rect -428 73 726 612
<< nmos >>
rect -258 -276 -243 -176
rect 19 -16 41 27
rect 296 -16 318 27
rect 573 -16 595 27
rect 26 -125 41 -82
rect 303 -125 318 -82
rect 580 -125 595 -82
rect 26 -276 41 -176
rect 303 -276 318 -176
rect 580 -276 595 -176
<< pmos >>
rect -323 382 -173 582
rect -46 382 104 582
rect 231 382 381 582
rect 508 382 658 582
rect 26 245 41 331
rect 303 245 318 331
rect 580 245 595 331
rect 19 93 41 179
rect 296 93 318 179
rect 573 93 595 179
<< ndiff >>
rect -308 -186 -258 -176
rect -308 -266 -293 -186
rect -273 -266 -258 -186
rect -308 -276 -258 -266
rect -243 -186 -193 -176
rect -243 -266 -228 -186
rect -208 -266 -193 -186
rect -243 -276 -193 -266
rect -31 19 19 27
rect -31 -6 -16 19
rect 4 -6 19 19
rect -31 -16 19 -6
rect 41 19 91 27
rect 41 -6 56 19
rect 76 -6 91 19
rect 41 -16 91 -6
rect 246 19 296 27
rect 246 -6 261 19
rect 281 -6 296 19
rect 246 -16 296 -6
rect 318 19 368 27
rect 318 -6 333 19
rect 353 -6 368 19
rect 318 -16 368 -6
rect 523 19 573 27
rect 523 -6 538 19
rect 558 -6 573 19
rect 523 -16 573 -6
rect 595 19 645 27
rect 595 -6 610 19
rect 630 -6 645 19
rect 595 -16 645 -6
rect -24 -92 26 -82
rect -24 -115 -9 -92
rect 11 -115 26 -92
rect -24 -125 26 -115
rect 41 -92 91 -82
rect 41 -115 56 -92
rect 76 -115 91 -92
rect 41 -125 91 -115
rect 253 -92 303 -82
rect 253 -115 268 -92
rect 288 -115 303 -92
rect 253 -125 303 -115
rect 318 -92 368 -82
rect 318 -115 333 -92
rect 353 -115 368 -92
rect 318 -125 368 -115
rect 530 -92 580 -82
rect 530 -115 545 -92
rect 565 -115 580 -92
rect 530 -125 580 -115
rect 595 -92 645 -82
rect 595 -115 610 -92
rect 630 -115 645 -92
rect 595 -125 645 -115
rect -24 -186 26 -176
rect -24 -266 -9 -186
rect 11 -266 26 -186
rect -24 -276 26 -266
rect 41 -186 91 -176
rect 41 -266 56 -186
rect 76 -266 91 -186
rect 41 -276 91 -266
rect 253 -186 303 -176
rect 253 -266 268 -186
rect 288 -266 303 -186
rect 253 -276 303 -266
rect 318 -186 368 -176
rect 318 -266 333 -186
rect 353 -266 368 -186
rect 318 -276 368 -266
rect 530 -186 580 -176
rect 530 -266 545 -186
rect 565 -266 580 -186
rect 530 -276 580 -266
rect 595 -186 645 -176
rect 595 -266 610 -186
rect 630 -266 645 -186
rect 595 -276 645 -266
<< pdiff >>
rect -373 572 -323 582
rect -373 392 -358 572
rect -338 392 -323 572
rect -373 382 -323 392
rect -173 572 -123 582
rect -173 392 -158 572
rect -138 392 -123 572
rect -173 382 -123 392
rect -96 572 -46 582
rect -96 392 -81 572
rect -61 392 -46 572
rect -96 382 -46 392
rect 104 572 154 582
rect 104 392 119 572
rect 139 392 154 572
rect 104 382 154 392
rect 181 572 231 582
rect 181 392 196 572
rect 216 392 231 572
rect 181 382 231 392
rect 381 572 431 582
rect 381 392 396 572
rect 416 392 431 572
rect 381 382 431 392
rect 458 572 508 582
rect 458 392 473 572
rect 493 392 508 572
rect 458 382 508 392
rect 658 572 708 582
rect 658 392 673 572
rect 693 392 708 572
rect 658 382 708 392
rect -24 321 26 331
rect -24 255 -9 321
rect 11 255 26 321
rect -24 245 26 255
rect 41 321 91 331
rect 41 255 56 321
rect 76 255 91 321
rect 41 245 91 255
rect 253 321 303 331
rect 253 255 268 321
rect 288 255 303 321
rect 253 245 303 255
rect 318 321 368 331
rect 318 255 333 321
rect 353 255 368 321
rect 318 245 368 255
rect 530 321 580 331
rect 530 255 545 321
rect 565 255 580 321
rect 530 245 580 255
rect 595 321 645 331
rect 595 255 610 321
rect 630 255 645 321
rect 595 245 645 255
rect -31 171 19 179
rect -31 103 -16 171
rect 4 103 19 171
rect -31 93 19 103
rect 41 171 91 179
rect 41 103 56 171
rect 76 103 91 171
rect 41 93 91 103
rect 246 171 296 179
rect 246 103 261 171
rect 281 103 296 171
rect 246 93 296 103
rect 318 171 368 179
rect 318 103 333 171
rect 353 103 368 171
rect 318 93 368 103
rect 523 171 573 179
rect 523 103 538 171
rect 558 103 573 171
rect 523 93 573 103
rect 595 171 645 179
rect 595 103 610 171
rect 630 103 645 171
rect 595 93 645 103
<< ndiffc >>
rect -293 -266 -273 -186
rect -228 -266 -208 -186
rect -16 -6 4 19
rect 56 -6 76 19
rect 261 -6 281 19
rect 333 -6 353 19
rect 538 -6 558 19
rect 610 -6 630 19
rect -9 -115 11 -92
rect 56 -115 76 -92
rect 268 -115 288 -92
rect 333 -115 353 -92
rect 545 -115 565 -92
rect 610 -115 630 -92
rect -9 -266 11 -186
rect 56 -266 76 -186
rect 268 -266 288 -186
rect 333 -266 353 -186
rect 545 -266 565 -186
rect 610 -266 630 -186
<< pdiffc >>
rect -358 392 -338 572
rect -158 392 -138 572
rect -81 392 -61 572
rect 119 392 139 572
rect 196 392 216 572
rect 396 392 416 572
rect 473 392 493 572
rect 673 392 693 572
rect -9 255 11 321
rect 56 255 76 321
rect 268 255 288 321
rect 333 255 353 321
rect 545 255 565 321
rect 610 255 630 321
rect -16 103 4 171
rect 56 103 76 171
rect 261 103 281 171
rect 333 103 353 171
rect 538 103 558 171
rect 610 103 630 171
<< psubdiff >>
rect 480 -92 530 -82
rect 480 -115 495 -92
rect 515 -115 530 -92
rect 480 -125 530 -115
<< nsubdiff >>
rect 203 321 253 331
rect 203 255 217 321
rect 237 255 253 321
rect 203 245 253 255
<< psubdiffcont >>
rect 495 -115 515 -92
<< nsubdiffcont >>
rect 217 255 237 321
<< poly >>
rect -323 626 -173 633
rect -323 606 -313 626
rect -185 606 -173 626
rect -323 582 -173 606
rect -46 626 104 633
rect -46 606 -36 626
rect 92 606 104 626
rect -46 582 104 606
rect 231 626 381 633
rect 231 606 241 626
rect 369 606 381 626
rect 231 582 381 606
rect 508 626 658 633
rect 508 606 518 626
rect 646 606 658 626
rect 508 582 658 606
rect -323 367 -173 382
rect -46 367 104 382
rect 231 367 381 382
rect 508 367 658 382
rect -323 357 -283 367
rect -323 337 -313 357
rect -293 337 -283 357
rect -323 327 -283 337
rect 26 331 41 346
rect 303 331 318 346
rect 580 331 595 346
rect 26 230 41 245
rect 303 230 318 245
rect 580 230 595 245
rect 26 220 595 230
rect 26 215 470 220
rect 460 200 470 215
rect 490 215 595 220
rect 490 200 500 215
rect 19 179 41 194
rect 296 179 318 194
rect 460 190 500 200
rect 573 179 595 194
rect 19 74 41 93
rect 296 74 318 93
rect 573 74 595 93
rect 19 69 81 74
rect -196 59 -156 69
rect -196 39 -186 59
rect -166 39 -156 59
rect -196 29 -156 39
rect -363 -161 -243 -146
rect -258 -176 -243 -161
rect -258 -291 -243 -276
rect -268 -299 -233 -291
rect -268 -318 -260 -299
rect -241 -318 -233 -299
rect -268 -326 -233 -318
rect -176 -350 -156 29
rect 19 49 51 69
rect 71 66 81 69
rect 239 69 275 74
rect 239 66 247 69
rect 71 51 247 66
rect 71 49 81 51
rect 19 44 81 49
rect 239 49 247 51
rect 267 49 275 69
rect 239 44 275 49
rect 296 69 354 74
rect 296 49 326 69
rect 346 66 354 69
rect 516 69 552 74
rect 516 66 524 69
rect 346 51 524 66
rect 346 49 354 51
rect 296 44 354 49
rect 516 49 524 51
rect 544 49 552 69
rect 516 44 552 49
rect 573 69 635 74
rect 573 49 605 69
rect 625 49 635 69
rect 573 44 635 49
rect 19 27 41 44
rect 296 27 318 44
rect 573 27 595 44
rect 19 -31 41 -16
rect 182 -37 222 -27
rect 296 -31 318 -16
rect 573 -31 595 -16
rect 182 -52 192 -37
rect 26 -57 192 -52
rect 212 -52 222 -37
rect 212 -57 595 -52
rect 26 -67 595 -57
rect 26 -82 41 -67
rect 303 -82 318 -67
rect 580 -82 595 -67
rect 26 -140 41 -125
rect 303 -140 318 -125
rect 580 -140 595 -125
rect 26 -176 41 -161
rect 303 -176 318 -161
rect 580 -176 595 -161
rect 26 -291 41 -276
rect 303 -291 318 -276
rect 580 -291 595 -276
rect 16 -299 51 -291
rect 16 -318 24 -299
rect 43 -318 51 -299
rect 16 -326 51 -318
rect 293 -299 328 -291
rect 293 -318 301 -299
rect 320 -318 328 -299
rect 293 -326 328 -318
rect 570 -299 605 -291
rect 570 -318 578 -299
rect 597 -318 605 -299
rect 570 -326 605 -318
rect -196 -360 -156 -350
rect -196 -380 -186 -360
rect -166 -380 -156 -360
rect -196 -390 -156 -380
<< polycont >>
rect -313 606 -185 626
rect -36 606 92 626
rect 241 606 369 626
rect 518 606 646 626
rect -313 337 -293 357
rect 470 200 490 220
rect -186 39 -166 59
rect -260 -318 -241 -299
rect 51 49 71 69
rect 247 49 267 69
rect 326 49 346 69
rect 524 49 544 69
rect 605 49 625 69
rect 192 -57 212 -37
rect 24 -318 43 -299
rect 301 -318 320 -299
rect 578 -318 597 -299
rect -186 -380 -166 -360
<< locali >>
rect -323 626 658 633
rect -323 606 -313 626
rect -185 606 -36 626
rect 92 606 241 626
rect 369 606 518 626
rect 646 606 658 626
rect -323 600 658 606
rect -368 572 -328 582
rect -368 392 -358 572
rect -338 392 -328 572
rect -368 385 -328 392
rect -168 572 -128 582
rect -168 392 -158 572
rect -138 392 -128 572
rect -368 347 -348 385
rect -168 382 -128 392
rect -91 572 -51 582
rect -91 392 -81 572
rect -61 392 -51 572
rect -91 382 -51 392
rect 109 572 149 582
rect 109 392 119 572
rect 139 392 149 572
rect -323 357 -283 367
rect -323 347 -313 357
rect -368 337 -313 347
rect -293 337 -283 357
rect -368 327 -283 337
rect 109 331 149 392
rect 186 572 226 582
rect 186 392 196 572
rect 216 392 226 572
rect 186 382 226 392
rect 386 572 426 582
rect 386 392 396 572
rect 416 392 426 572
rect 386 331 426 392
rect 463 572 503 582
rect 463 392 473 572
rect 493 392 503 572
rect 463 382 503 392
rect 663 572 703 582
rect 663 392 673 572
rect 693 392 703 572
rect 663 331 703 392
rect -303 -186 -283 327
rect -19 321 21 331
rect -19 292 -9 321
rect -24 255 -9 292
rect 11 255 21 321
rect -24 252 21 255
rect 46 321 149 331
rect 46 255 56 321
rect 76 297 149 321
rect 203 321 254 330
rect 323 321 426 331
rect 76 255 86 297
rect 46 171 86 255
rect 203 255 217 321
rect 237 255 268 321
rect 288 255 298 321
rect 323 255 333 321
rect 353 297 426 321
rect 535 321 575 331
rect 353 255 363 297
rect 203 245 254 255
rect -26 103 -16 171
rect 4 103 14 171
rect -26 69 14 103
rect 46 103 56 171
rect 76 103 86 171
rect 46 93 86 103
rect -196 59 14 69
rect -196 39 -186 59
rect -166 49 14 59
rect -166 39 -156 49
rect -196 29 -156 39
rect -26 19 14 49
rect 41 69 81 74
rect 41 49 51 69
rect 71 49 81 69
rect 41 44 81 49
rect -26 -6 -16 19
rect 4 -6 14 19
rect -26 -16 14 -6
rect 46 19 86 27
rect 46 -6 56 19
rect 76 -6 86 19
rect -19 -92 21 -82
rect -19 -115 -9 -92
rect 11 -115 21 -92
rect -19 -125 21 -115
rect 46 -92 86 -6
rect 202 -27 222 245
rect 323 171 363 255
rect 535 255 545 321
rect 565 255 575 321
rect 535 245 575 255
rect 600 321 703 331
rect 600 255 610 321
rect 630 297 703 321
rect 630 255 640 297
rect 251 103 261 171
rect 281 103 291 171
rect 251 74 291 103
rect 323 103 333 171
rect 353 103 363 171
rect 323 93 363 103
rect 460 220 500 230
rect 460 200 470 220
rect 490 200 500 220
rect 460 190 500 200
rect 239 69 291 74
rect 239 49 247 69
rect 267 49 291 69
rect 239 44 291 49
rect 318 69 354 74
rect 318 49 326 69
rect 346 49 354 69
rect 318 44 354 49
rect 251 19 291 44
rect 251 -6 261 19
rect 281 -6 291 19
rect 251 -16 291 -6
rect 323 19 363 27
rect 323 -6 333 19
rect 353 -6 363 19
rect 182 -37 222 -27
rect 182 -57 192 -37
rect 212 -57 222 -37
rect 182 -67 222 -57
rect 46 -115 56 -92
rect 76 -115 86 -92
rect 46 -186 86 -115
rect 258 -92 298 -82
rect 258 -115 268 -92
rect 288 -115 298 -92
rect 258 -125 298 -115
rect 323 -92 363 -6
rect 323 -115 333 -92
rect 353 -115 363 -92
rect 460 -82 480 190
rect 600 171 640 255
rect 528 103 538 171
rect 558 103 568 171
rect 528 75 568 103
rect 600 103 610 171
rect 630 103 640 171
rect 600 93 640 103
rect 527 74 568 75
rect 516 69 568 74
rect 516 49 524 69
rect 544 49 568 69
rect 516 44 568 49
rect 595 69 635 74
rect 595 49 605 69
rect 625 49 737 69
rect 595 44 635 49
rect 527 43 568 44
rect 528 19 568 43
rect 528 -6 538 19
rect 558 -6 568 19
rect 528 -16 568 -6
rect 600 19 640 27
rect 600 -6 610 19
rect 630 -6 640 19
rect 460 -92 575 -82
rect 460 -102 495 -92
rect 323 -186 363 -115
rect 480 -115 495 -102
rect 515 -115 545 -92
rect 565 -115 575 -92
rect 480 -125 575 -115
rect 600 -92 640 -6
rect 600 -115 610 -92
rect 630 -115 640 -92
rect -303 -266 -293 -186
rect -273 -266 -263 -186
rect -238 -266 -228 -186
rect -208 -266 -198 -186
rect -19 -266 -9 -186
rect 11 -266 21 -186
rect 46 -266 56 -186
rect 76 -266 86 -186
rect 253 -266 268 -186
rect 288 -266 298 -186
rect 323 -266 333 -186
rect 353 -266 363 -186
rect 535 -186 575 -176
rect 535 -266 545 -186
rect 565 -266 575 -186
rect 600 -186 640 -115
rect 600 -266 610 -186
rect 630 -266 640 -186
rect -268 -299 605 -291
rect -268 -318 -260 -299
rect -241 -318 24 -299
rect 43 -318 301 -299
rect 320 -318 578 -299
rect 597 -318 605 -299
rect -268 -326 605 -318
rect -196 -360 -156 -350
rect -196 -380 -186 -360
rect -166 -370 -156 -360
rect 657 -370 677 49
rect -166 -380 677 -370
rect -196 -390 677 -380
<< viali >>
rect -158 392 -138 572
rect -81 392 -61 572
rect 196 392 216 572
rect 473 392 493 572
rect -9 255 11 321
rect 217 255 237 321
rect 268 255 288 321
rect -9 -115 11 -92
rect 545 255 565 321
rect 268 -115 288 -92
rect 495 -115 515 -92
rect 545 -115 565 -92
rect -228 -266 -208 -186
rect -9 -266 11 -186
rect 268 -266 288 -186
rect 545 -266 565 -186
<< metal1 >>
rect -373 572 708 575
rect -373 392 -158 572
rect -138 392 -81 572
rect -61 392 196 572
rect 216 392 473 572
rect 493 392 708 572
rect -373 321 708 392
rect -373 255 -9 321
rect 11 255 217 321
rect 237 255 268 321
rect 288 255 545 321
rect 565 255 708 321
rect -373 252 708 255
rect -308 -92 645 -89
rect -308 -115 -9 -92
rect 11 -115 268 -92
rect 288 -115 495 -92
rect 515 -115 545 -92
rect 565 -115 645 -92
rect -308 -186 645 -115
rect -308 -266 -228 -186
rect -208 -266 -9 -186
rect 11 -266 268 -186
rect 288 -266 545 -186
rect 565 -266 645 -186
rect -308 -269 645 -266
<< labels >>
flabel metal1 -373 482 -373 482 7 FreeSans 80 0 0 0 VDDA
flabel locali 737 59 737 59 3 FreeSans 80 0 0 0 V_OSC
flabel poly -363 -154 -363 -154 7 FreeSans 80 0 0 0 V_CONT
flabel metal1 -308 -226 -308 -226 7 FreeSans 80 0 0 0 GNDA
<< end >>
