* PEX produced on Wed Jul 16 04:55:32 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic_13.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic_13 VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 GNDA.t192 bgr_9_0.NFET_GATE_10uA.t5 two_stage_opamp_dummy_magic_19_0.Vb3.t6 GNDA.t191 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1 bgr_9_0.V_TOP.t11 VDDA.t354 VDDA.t356 VDDA.t355 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.45 ps=2.9 w=1 l=0.15
X2 VOUT-.t19 two_stage_opamp_dummy_magic_19_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 two_stage_opamp_dummy_magic_19_0.err_amp_mir.t3 GNDA.t287 GNDA.t288 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X4 GNDA.t115 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t8 two_stage_opamp_dummy_magic_19_0.V_source.t37 GNDA.t114 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X5 VOUT+.t19 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 VOUT+.t14 GNDA.t284 GNDA.t286 GNDA.t285 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X7 VDDA.t101 two_stage_opamp_dummy_magic_19_0.X.t25 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t9 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X8 VOUT+.t20 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 VDDA.t82 bgr_9_0.V_TOP.t14 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t6 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X10 VDDA.t353 VDDA.t351 two_stage_opamp_dummy_magic_19_0.err_amp_out.t3 VDDA.t352 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X11 VOUT+.t21 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 GNDA.t283 GNDA.t281 VDDA.t240 GNDA.t282 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X13 bgr_9_0.Vin+.t5 bgr_9_0.V_TOP.t15 VDDA.t84 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X14 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t12 two_stage_opamp_dummy_magic_19_0.X.t26 GNDA.t84 VDDA.t102 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X15 VDDA.t146 bgr_9_0.V_mir1.t17 bgr_9_0.1st_Vout_1.t5 VDDA.t145 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X16 VOUT+.t22 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 bgr_9_0.1st_Vout_2.t11 bgr_9_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 two_stage_opamp_dummy_magic_19_0.X.t3 two_stage_opamp_dummy_magic_19_0.Vb2.t11 two_stage_opamp_dummy_magic_19_0.VD3.t19 two_stage_opamp_dummy_magic_19_0.VD3.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X19 GNDA.t37 two_stage_opamp_dummy_magic_19_0.Y.t25 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t12 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X20 VOUT+.t23 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 bgr_9_0.1st_Vout_2.t4 bgr_9_0.V_CUR_REF_REG.t3 bgr_9_0.V_p_2.t9 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X22 VOUT+.t24 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X23 VOUT+.t25 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X24 a_7460_23988.t0 bgr_9_0.Vin+.t1 GNDA.t90 sky130_fd_pr__res_xhigh_po_0p35 l=6
X25 two_stage_opamp_dummy_magic_19_0.VD2.t18 GNDA.t279 GNDA.t280 GNDA.t201 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X26 VDDA.t104 two_stage_opamp_dummy_magic_19_0.V_err_gate.t6 two_stage_opamp_dummy_magic_19_0.V_err_mir_p.t2 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X27 two_stage_opamp_dummy_magic_19_0.VD1.t13 two_stage_opamp_dummy_magic_19_0.Vb1.t12 two_stage_opamp_dummy_magic_19_0.X.t0 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X28 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t2 GNDA.t277 GNDA.t278 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X29 VOUT+.t26 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 VOUT+.t11 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t2 GNDA.t135 GNDA.t134 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X31 two_stage_opamp_dummy_magic_19_0.VD1.t12 two_stage_opamp_dummy_magic_19_0.Vb1.t13 two_stage_opamp_dummy_magic_19_0.X.t5 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X32 bgr_9_0.1st_Vout_2.t12 bgr_9_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 two_stage_opamp_dummy_magic_19_0.VD2.t4 two_stage_opamp_dummy_magic_19_0.Vb1.t14 two_stage_opamp_dummy_magic_19_0.Y.t13 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X34 GNDA.t89 a_6930_22564.t1 GNDA.t75 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X35 VDDA.t350 VDDA.t348 VDDA.t350 VDDA.t349 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0 ps=0 w=2 l=0.15
X36 GNDA.t276 GNDA.t275 two_stage_opamp_dummy_magic_19_0.Y.t22 GNDA.t270 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X37 VDDA.t358 bgr_9_0.PFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t4 VDDA.t357 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X38 VOUT-.t20 two_stage_opamp_dummy_magic_19_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 VOUT-.t21 two_stage_opamp_dummy_magic_19_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 VOUT-.t22 two_stage_opamp_dummy_magic_19_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X41 VOUT+.t27 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 bgr_9_0.1st_Vout_1.t11 bgr_9_0.cap_res1.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 bgr_9_0.1st_Vout_2.t5 bgr_9_0.V_mir2.t17 VDDA.t91 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X44 VDDA.t86 bgr_9_0.V_TOP.t16 bgr_9_0.Vin-.t6 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X45 VOUT+.t10 a_5820_2720.t1 GNDA.t133 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X46 bgr_9_0.1st_Vout_1.t6 bgr_9_0.Vin+.t6 bgr_9_0.V_p_1.t9 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X47 GNDA.t150 VDDA.t412 bgr_9_0.V_p_2.t10 GNDA.t149 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X48 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t8 two_stage_opamp_dummy_magic_19_0.X.t27 VDDA.t171 GNDA.t123 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X49 VOUT+.t28 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 bgr_9_0.cap_res2.t20 bgr_9_0.PFET_GATE_10uA.t6 GNDA.t103 sky130_fd_pr__res_high_po_0p35 l=2.05
X51 bgr_9_0.1st_Vout_1.t12 bgr_9_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t7 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t6 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0 ps=0 w=3.5 l=0.2
X53 VOUT-.t16 two_stage_opamp_dummy_magic_19_0.X.t28 VDDA.t375 VDDA.t374 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X54 two_stage_opamp_dummy_magic_19_0.V_source.t14 VIN-.t0 two_stage_opamp_dummy_magic_19_0.VD1.t17 GNDA.t102 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X55 VOUT+.t29 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X56 VOUT-.t23 two_stage_opamp_dummy_magic_19_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X57 two_stage_opamp_dummy_magic_19_0.V_source.t19 two_stage_opamp_dummy_magic_19_0.Vb1.t15 two_stage_opamp_dummy_magic_19_0.Vb1_2.t0 GNDA.t148 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.6 ps=3.8 w=1.5 l=3
X58 two_stage_opamp_dummy_magic_19_0.VD4.t35 two_stage_opamp_dummy_magic_19_0.Vb3.t8 VDDA.t236 VDDA.t235 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X59 two_stage_opamp_dummy_magic_19_0.V_source.t9 VIN+.t0 two_stage_opamp_dummy_magic_19_0.VD2.t8 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X60 VOUT-.t24 two_stage_opamp_dummy_magic_19_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 VOUT-.t25 two_stage_opamp_dummy_magic_19_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X62 VDDA.t34 two_stage_opamp_dummy_magic_19_0.Y.t26 VOUT+.t4 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X63 two_stage_opamp_dummy_magic_19_0.err_amp_out.t1 two_stage_opamp_dummy_magic_19_0.err_amp_mir.t5 GNDA.t72 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X64 two_stage_opamp_dummy_magic_19_0.V_source.t36 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t9 GNDA.t117 GNDA.t116 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X65 VDDA.t397 bgr_9_0.1st_Vout_1.t13 bgr_9_0.V_TOP.t13 VDDA.t396 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X66 bgr_9_0.V_TOP.t17 VDDA.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 VOUT-.t26 two_stage_opamp_dummy_magic_19_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 GNDA.t274 GNDA.t272 bgr_9_0.NFET_GATE_10uA.t0 GNDA.t273 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X69 bgr_9_0.START_UP.t5 bgr_9_0.V_TOP.t18 VDDA.t62 VDDA.t61 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X70 VOUT-.t27 two_stage_opamp_dummy_magic_19_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X71 two_stage_opamp_dummy_magic_19_0.V_err_gate.t3 bgr_9_0.NFET_GATE_10uA.t6 GNDA.t190 GNDA.t189 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X72 VDDA.t234 two_stage_opamp_dummy_magic_19_0.Vb3.t9 two_stage_opamp_dummy_magic_19_0.VD3.t35 VDDA.t233 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X73 bgr_9_0.1st_Vout_1.t10 bgr_9_0.Vin+.t7 bgr_9_0.V_p_1.t8 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X74 VOUT-.t28 two_stage_opamp_dummy_magic_19_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 GNDA.t14 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t10 two_stage_opamp_dummy_magic_19_0.V_source.t35 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X76 VOUT+.t30 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X77 VOUT-.t7 a_14170_2720.t0 GNDA.t120 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X78 VDDA.t66 two_stage_opamp_dummy_magic_19_0.X.t29 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t7 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X79 bgr_9_0.1st_Vout_1.t14 bgr_9_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X80 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t10 two_stage_opamp_dummy_magic_19_0.Y.t27 VDDA.t54 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X81 two_stage_opamp_dummy_magic_19_0.V_err_p.t2 two_stage_opamp_dummy_magic_19_0.V_err_gate.t7 VDDA.t13 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X82 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t7 VIN-.t1 two_stage_opamp_dummy_magic_19_0.V_p_mir.t5 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X83 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t9 two_stage_opamp_dummy_magic_19_0.Y.t28 VDDA.t40 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X84 bgr_9_0.V_TOP.t19 VDDA.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 bgr_9_0.V_mir2.t11 bgr_9_0.V_mir2.t10 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X86 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t15 VDDA.t333 VDDA.t335 VDDA.t334 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X87 VOUT-.t29 two_stage_opamp_dummy_magic_19_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t2 bgr_9_0.PFET_GATE_10uA.t11 VDDA.t164 VDDA.t163 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X89 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t10 VDDA.t345 VDDA.t347 VDDA.t346 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X90 VDDA.t7 bgr_9_0.PFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t0 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X91 GNDA.t36 two_stage_opamp_dummy_magic_19_0.Y.t29 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t11 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X92 VOUT+.t31 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X93 bgr_9_0.V_TOP.t20 VDDA.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X94 GNDA.t16 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t11 two_stage_opamp_dummy_magic_19_0.V_source.t34 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X95 bgr_9_0.1st_Vout_2.t2 bgr_9_0.V_CUR_REF_REG.t4 bgr_9_0.V_p_2.t8 GNDA.t50 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X96 two_stage_opamp_dummy_magic_19_0.VD4.t19 two_stage_opamp_dummy_magic_19_0.Vb2.t12 two_stage_opamp_dummy_magic_19_0.Y.t2 two_stage_opamp_dummy_magic_19_0.VD4.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X97 VOUT-.t30 two_stage_opamp_dummy_magic_19_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X98 VOUT-.t31 two_stage_opamp_dummy_magic_19_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X99 VOUT-.t32 two_stage_opamp_dummy_magic_19_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_19_0.Vb3.t2 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t3 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X101 two_stage_opamp_dummy_magic_19_0.VD2.t19 two_stage_opamp_dummy_magic_19_0.Vb1.t16 two_stage_opamp_dummy_magic_19_0.Y.t23 GNDA.t304 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X102 two_stage_opamp_dummy_magic_19_0.V_source.t33 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t12 GNDA.t57 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X103 bgr_9_0.PFET_GATE_10uA.t5 bgr_9_0.1st_Vout_2.t13 VDDA.t403 VDDA.t402 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X104 VOUT-.t33 two_stage_opamp_dummy_magic_19_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 bgr_9_0.V_TOP.t21 VDDA.t181 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X106 bgr_9_0.START_UP_NFET1.t0 bgr_9_0.START_UP_NFET1 GNDA.t86 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X107 two_stage_opamp_dummy_magic_19_0.VD3.t17 two_stage_opamp_dummy_magic_19_0.Vb2.t13 two_stage_opamp_dummy_magic_19_0.X.t10 two_stage_opamp_dummy_magic_19_0.VD3.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X108 VOUT+.t32 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X109 two_stage_opamp_dummy_magic_19_0.V_source.t4 VIN-.t2 two_stage_opamp_dummy_magic_19_0.VD1.t1 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X110 bgr_9_0.V_CUR_REF_REG.t2 VDDA.t342 VDDA.t344 VDDA.t343 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X111 VOUT-.t12 VDDA.t339 VDDA.t341 VDDA.t340 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X112 two_stage_opamp_dummy_magic_19_0.V_source.t11 VIN-.t3 two_stage_opamp_dummy_magic_19_0.VD1.t14 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X113 VOUT+.t33 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 bgr_9_0.V_TOP.t22 VDDA.t182 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 GNDA.t188 bgr_9_0.NFET_GATE_10uA.t7 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t13 GNDA.t187 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X116 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t12 bgr_9_0.NFET_GATE_10uA.t8 GNDA.t186 GNDA.t185 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X117 two_stage_opamp_dummy_magic_19_0.VD4.t17 two_stage_opamp_dummy_magic_19_0.Vb2.t14 two_stage_opamp_dummy_magic_19_0.Y.t7 two_stage_opamp_dummy_magic_19_0.VD4.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X118 two_stage_opamp_dummy_magic_19_0.V_source.t15 VIN+.t1 two_stage_opamp_dummy_magic_19_0.VD2.t14 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X119 VDDA.t53 two_stage_opamp_dummy_magic_19_0.Y.t30 VOUT+.t5 VDDA.t52 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X120 GNDA.t271 GNDA.t269 two_stage_opamp_dummy_magic_19_0.VD2.t17 GNDA.t270 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X121 VOUT-.t34 two_stage_opamp_dummy_magic_19_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 two_stage_opamp_dummy_magic_19_0.V_source.t32 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t13 GNDA.t59 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X123 VOUT-.t35 two_stage_opamp_dummy_magic_19_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 VOUT-.t36 two_stage_opamp_dummy_magic_19_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 VOUT-.t37 two_stage_opamp_dummy_magic_19_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 bgr_9_0.1st_Vout_2.t14 bgr_9_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X127 VOUT+.t34 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 VOUT+.t35 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 two_stage_opamp_dummy_magic_19_0.Vb1.t2 two_stage_opamp_dummy_magic_19_0.Vb1.t1 two_stage_opamp_dummy_magic_19_0.Vb1_2.t4 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X130 VOUT+.t36 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 VOUT+.t37 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X132 VOUT+.t38 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 GNDA.t60 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t14 two_stage_opamp_dummy_magic_19_0.V_source.t31 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X134 a_12530_23988.t0 bgr_9_0.Vin-.t1 GNDA.t66 sky130_fd_pr__res_xhigh_po_0p35 l=6
X135 two_stage_opamp_dummy_magic_19_0.VD3.t15 two_stage_opamp_dummy_magic_19_0.Vb2.t15 two_stage_opamp_dummy_magic_19_0.X.t13 two_stage_opamp_dummy_magic_19_0.VD3.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X136 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t8 two_stage_opamp_dummy_magic_19_0.Y.t31 VDDA.t139 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X137 VOUT-.t38 two_stage_opamp_dummy_magic_19_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 VOUT-.t39 two_stage_opamp_dummy_magic_19_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 bgr_9_0.1st_Vout_2.t9 bgr_9_0.V_mir2.t18 VDDA.t192 VDDA.t191 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X140 two_stage_opamp_dummy_magic_19_0.V_err_p.t0 two_stage_opamp_dummy_magic_19_0.V_tot.t4 two_stage_opamp_dummy_magic_19_0.err_amp_mir.t0 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X141 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t11 two_stage_opamp_dummy_magic_19_0.X.t30 GNDA.t40 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X142 VOUT-.t40 two_stage_opamp_dummy_magic_19_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X143 GNDA.t47 two_stage_opamp_dummy_magic_19_0.Y.t32 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t10 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X144 VOUT-.t41 two_stage_opamp_dummy_magic_19_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 bgr_9_0.1st_Vout_2.t15 bgr_9_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X146 VDDA.t338 VDDA.t336 VDDA.t338 VDDA.t337 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0 ps=0 w=2 l=0.15
X147 VOUT-.t42 two_stage_opamp_dummy_magic_19_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 VOUT+.t39 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 VOUT-.t43 two_stage_opamp_dummy_magic_19_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 VOUT+.t40 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 VOUT+.t41 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 bgr_9_0.1st_Vout_1.t15 bgr_9_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X153 VOUT+.t42 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 bgr_9_0.V_mir1.t14 bgr_9_0.Vin-.t8 bgr_9_0.V_p_1.t4 GNDA.t131 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X155 bgr_9_0.V_mir1.t12 bgr_9_0.V_mir1.t11 VDDA.t10 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X156 two_stage_opamp_dummy_magic_19_0.VD2.t10 two_stage_opamp_dummy_magic_19_0.Vb1.t17 two_stage_opamp_dummy_magic_19_0.Y.t16 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X157 GNDA.t119 a_7580_22380.t0 GNDA.t90 sky130_fd_pr__res_xhigh_po_0p35 l=6
X158 VOUT-.t44 two_stage_opamp_dummy_magic_19_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 two_stage_opamp_dummy_magic_19_0.Vb3.t1 two_stage_opamp_dummy_magic_19_0.Vb2.t16 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X160 VOUT-.t45 two_stage_opamp_dummy_magic_19_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X161 VOUT+.t43 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 VOUT-.t46 two_stage_opamp_dummy_magic_19_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X163 VOUT-.t47 two_stage_opamp_dummy_magic_19_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 VOUT-.t48 two_stage_opamp_dummy_magic_19_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 VDDA.t232 two_stage_opamp_dummy_magic_19_0.Vb3.t10 two_stage_opamp_dummy_magic_19_0.VD4.t34 VDDA.t231 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X166 bgr_9_0.V_TOP.t23 VDDA.t183 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X167 VDDA.t332 VDDA.t330 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t14 VDDA.t331 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X168 VOUT-.t49 two_stage_opamp_dummy_magic_19_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X169 VOUT-.t50 two_stage_opamp_dummy_magic_19_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X170 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t16 bgr_9_0.PFET_GATE_10uA.t13 VDDA.t409 VDDA.t408 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X171 VOUT-.t13 two_stage_opamp_dummy_magic_19_0.X.t31 VDDA.t371 VDDA.t370 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X172 VOUT+.t44 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X173 VOUT+.t45 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 two_stage_opamp_dummy_magic_19_0.V_source.t39 VIN+.t2 two_stage_opamp_dummy_magic_19_0.VD2.t20 GNDA.t304 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X175 bgr_9_0.V_mir1.t16 bgr_9_0.Vin-.t9 bgr_9_0.V_p_1.t3 GNDA.t300 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X176 two_stage_opamp_dummy_magic_19_0.X.t4 two_stage_opamp_dummy_magic_19_0.Vb1.t18 two_stage_opamp_dummy_magic_19_0.VD1.t11 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X177 VOUT+.t46 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X178 two_stage_opamp_dummy_magic_19_0.VD3.t34 two_stage_opamp_dummy_magic_19_0.Vb3.t11 VDDA.t230 VDDA.t229 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X179 VOUT+.t47 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X180 two_stage_opamp_dummy_magic_19_0.VD3.t13 two_stage_opamp_dummy_magic_19_0.Vb2.t17 two_stage_opamp_dummy_magic_19_0.X.t2 two_stage_opamp_dummy_magic_19_0.VD3.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X181 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t1 a_14170_2720.t1 GNDA.t128 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X182 two_stage_opamp_dummy_magic_19_0.Vb1.t10 GNDA.t267 GNDA.t268 GNDA.t136 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X183 bgr_9_0.START_UP.t4 bgr_9_0.V_TOP.t24 VDDA.t177 VDDA.t176 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X184 VOUT-.t51 two_stage_opamp_dummy_magic_19_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 bgr_9_0.PFET_GATE_10uA.t4 bgr_9_0.1st_Vout_2.t16 VDDA.t391 VDDA.t390 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X186 VDDA.t381 bgr_9_0.V_mir1.t18 bgr_9_0.1st_Vout_1.t4 VDDA.t380 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X187 VOUT+.t48 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 VOUT+.t49 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 VOUT-.t52 two_stage_opamp_dummy_magic_19_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X190 VDDA.t67 two_stage_opamp_dummy_magic_19_0.X.t32 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t6 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X191 VOUT-.t53 two_stage_opamp_dummy_magic_19_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 two_stage_opamp_dummy_magic_19_0.Vb2.t8 bgr_9_0.NFET_GATE_10uA.t9 GNDA.t184 GNDA.t183 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X193 VDDA.t228 two_stage_opamp_dummy_magic_19_0.Vb3.t12 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t9 VDDA.t227 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X194 GNDA.t182 bgr_9_0.NFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_19_0.Vb2.t7 GNDA.t181 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X195 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t7 two_stage_opamp_dummy_magic_19_0.Y.t33 VDDA.t138 GNDA.t99 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X196 VOUT+.t50 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 bgr_9_0.V_TOP.t25 VDDA.t178 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 GNDA.t180 bgr_9_0.NFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_19_0.Vb2.t6 GNDA.t179 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X199 two_stage_opamp_dummy_magic_19_0.Y.t4 two_stage_opamp_dummy_magic_19_0.Vb2.t18 two_stage_opamp_dummy_magic_19_0.VD4.t15 two_stage_opamp_dummy_magic_19_0.VD4.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X200 VDDA.t329 VDDA.t327 VOUT-.t11 VDDA.t328 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X201 VOUT+.t51 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 VOUT-.t54 two_stage_opamp_dummy_magic_19_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X203 GNDA.t291 VDDA.t324 VDDA.t326 VDDA.t325 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X204 GNDA.t92 two_stage_opamp_dummy_magic_19_0.Y.t34 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t9 VDDA.t117 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X205 VOUT+.t52 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X206 VOUT+.t53 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 VOUT+.t54 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 VOUT+.t55 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 VDDA.t180 bgr_9_0.V_TOP.t26 bgr_9_0.Vin+.t4 VDDA.t179 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X210 bgr_9_0.1st_Vout_2.t3 bgr_9_0.V_mir2.t19 VDDA.t73 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X211 VOUT-.t55 two_stage_opamp_dummy_magic_19_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 bgr_9_0.V_TOP.t2 bgr_9_0.1st_Vout_1.t16 VDDA.t106 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X213 VOUT-.t56 two_stage_opamp_dummy_magic_19_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X214 VOUT-.t57 two_stage_opamp_dummy_magic_19_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X215 VOUT-.t58 two_stage_opamp_dummy_magic_19_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 VOUT+.t56 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t5 bgr_9_0.PFET_GATE_10uA.t14 VDDA.t360 VDDA.t359 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X218 VOUT-.t59 two_stage_opamp_dummy_magic_19_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X219 two_stage_opamp_dummy_magic_19_0.X.t11 two_stage_opamp_dummy_magic_19_0.Vb2.t19 two_stage_opamp_dummy_magic_19_0.VD3.t11 two_stage_opamp_dummy_magic_19_0.VD3.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X220 a_14330_5524.t0 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t10 GNDA.t127 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X221 VOUT+.t57 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 VOUT+.t58 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 bgr_9_0.1st_Vout_2.t17 bgr_9_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X224 a_6810_23838.t1 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t0 GNDA.t75 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X225 two_stage_opamp_dummy_magic_19_0.Y.t1 two_stage_opamp_dummy_magic_19_0.Vb2.t20 two_stage_opamp_dummy_magic_19_0.VD4.t13 two_stage_opamp_dummy_magic_19_0.VD4.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X226 bgr_9_0.Vin+.t0 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 GNDA.t26 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X227 VOUT+.t59 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X228 VOUT+.t60 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 VOUT-.t60 two_stage_opamp_dummy_magic_19_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 VOUT-.t61 two_stage_opamp_dummy_magic_19_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X231 bgr_9_0.1st_Vout_2.t18 bgr_9_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 bgr_9_0.Vin+.t3 bgr_9_0.V_TOP.t27 VDDA.t156 VDDA.t155 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X233 VOUT-.t3 two_stage_opamp_dummy_magic_19_0.X.t33 VDDA.t97 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X234 VOUT-.t62 two_stage_opamp_dummy_magic_19_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X235 VDDA.t323 VDDA.t321 bgr_9_0.PFET_GATE_10uA.t9 VDDA.t322 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X236 VOUT+.t61 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X237 VDDA.t158 bgr_9_0.V_TOP.t28 bgr_9_0.Vin+.t2 VDDA.t157 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X238 two_stage_opamp_dummy_magic_19_0.V_source.t7 VIN+.t3 two_stage_opamp_dummy_magic_19_0.VD2.t7 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X239 VOUT+.t62 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 two_stage_opamp_dummy_magic_19_0.X.t23 two_stage_opamp_dummy_magic_19_0.Vb1.t19 two_stage_opamp_dummy_magic_19_0.VD1.t10 GNDA.t309 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X241 bgr_9_0.1st_Vout_1.t17 bgr_9_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X242 GNDA.t308 a_12410_22380.t1 GNDA.t307 sky130_fd_pr__res_xhigh_po_0p35 l=6
X243 GNDA.t178 bgr_9_0.NFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_19_0.Vb3.t5 GNDA.t177 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X244 VOUT-.t63 two_stage_opamp_dummy_magic_19_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 VOUT-.t64 two_stage_opamp_dummy_magic_19_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_19_0.Y.t11 GNDA.t25 sky130_fd_pr__res_high_po_1p41 l=1.41
X247 VOUT+.t63 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X248 bgr_9_0.cap_res1.t0 bgr_9_0.V_TOP.t3 GNDA.t96 sky130_fd_pr__res_high_po_0p35 l=2.05
X249 two_stage_opamp_dummy_magic_19_0.Vb3.t4 bgr_9_0.NFET_GATE_10uA.t13 GNDA.t176 GNDA.t175 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X250 bgr_9_0.V_mir2.t9 bgr_9_0.V_mir2.t8 VDDA.t141 VDDA.t140 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X251 GNDA.t302 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t3 VOUT-.t18 GNDA.t301 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X252 VDDA.t320 VDDA.t318 bgr_9_0.V_TOP.t10 VDDA.t319 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X253 two_stage_opamp_dummy_magic_19_0.X.t22 two_stage_opamp_dummy_magic_19_0.Vb2.t21 two_stage_opamp_dummy_magic_19_0.VD3.t9 two_stage_opamp_dummy_magic_19_0.VD3.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X254 VOUT+.t64 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X255 VOUT+.t65 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 VDDA.t239 GNDA.t264 GNDA.t266 GNDA.t265 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X257 bgr_9_0.1st_Vout_1.t18 bgr_9_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 VOUT-.t65 two_stage_opamp_dummy_magic_19_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X259 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t6 two_stage_opamp_dummy_magic_19_0.Y.t35 VDDA.t116 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X260 VOUT+.t66 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X261 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t5 bgr_9_0.V_TOP.t29 VDDA.t160 VDDA.t159 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X262 bgr_9_0.1st_Vout_2.t19 bgr_9_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 two_stage_opamp_dummy_magic_19_0.VD1.t0 VIN-.t4 two_stage_opamp_dummy_magic_19_0.V_source.t0 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X264 VOUT-.t66 two_stage_opamp_dummy_magic_19_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 GNDA.t312 a_13060_22630.t1 GNDA.t311 sky130_fd_pr__res_xhigh_po_0p35 l=4
X266 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t10 two_stage_opamp_dummy_magic_19_0.X.t34 GNDA.t316 VDDA.t411 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X267 VDDA.t71 two_stage_opamp_dummy_magic_19_0.X.t35 VOUT-.t2 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X268 VOUT+.t67 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 bgr_9_0.1st_Vout_1.t3 bgr_9_0.V_mir1.t19 VDDA.t383 VDDA.t382 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X270 VOUT+.t7 two_stage_opamp_dummy_magic_19_0.Y.t36 VDDA.t113 VDDA.t112 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X271 a_5420_5524.t1 two_stage_opamp_dummy_magic_19_0.V_tot.t2 GNDA.t294 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X272 bgr_9_0.1st_Vout_1.t19 bgr_9_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X273 two_stage_opamp_dummy_magic_19_0.X.t8 two_stage_opamp_dummy_magic_19_0.Vb2.t22 two_stage_opamp_dummy_magic_19_0.VD3.t7 two_stage_opamp_dummy_magic_19_0.VD3.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X274 VOUT-.t67 two_stage_opamp_dummy_magic_19_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X275 GNDA.t195 GNDA.t193 VOUT-.t10 GNDA.t194 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X276 two_stage_opamp_dummy_magic_19_0.VD4.t37 VDDA.t300 VDDA.t302 VDDA.t301 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X277 two_stage_opamp_dummy_magic_19_0.V_err_gate.t5 VDDA.t303 VDDA.t305 VDDA.t304 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X278 VDDA.t308 VDDA.t306 bgr_9_0.NFET_GATE_10uA.t3 VDDA.t307 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X279 two_stage_opamp_dummy_magic_19_0.Vb1_2.t3 two_stage_opamp_dummy_magic_19_0.Vb1.t7 two_stage_opamp_dummy_magic_19_0.Vb1.t8 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X280 VDDA.t362 bgr_9_0.PFET_GATE_10uA.t15 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t6 VDDA.t361 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X281 two_stage_opamp_dummy_magic_19_0.Y.t10 two_stage_opamp_dummy_magic_19_0.Vb2.t23 two_stage_opamp_dummy_magic_19_0.VD4.t11 two_stage_opamp_dummy_magic_19_0.VD4.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X282 two_stage_opamp_dummy_magic_19_0.VD2.t1 two_stage_opamp_dummy_magic_19_0.Vb1.t20 two_stage_opamp_dummy_magic_19_0.Y.t0 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X283 VOUT+.t68 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 two_stage_opamp_dummy_magic_19_0.V_p_mir.t3 GNDA.t262 GNDA.t263 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X285 VOUT+.t69 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 bgr_9_0.1st_Vout_1.t20 bgr_9_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X287 bgr_9_0.V_p_2.t4 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t7 bgr_9_0.V_mir2.t16 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X288 two_stage_opamp_dummy_magic_19_0.V_source.t17 two_stage_opamp_dummy_magic_19_0.err_amp_out.t4 GNDA.t125 GNDA.t124 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X289 VDDA.t226 two_stage_opamp_dummy_magic_19_0.Vb3.t13 two_stage_opamp_dummy_magic_19_0.VD3.t33 VDDA.t225 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X290 VDDA.t393 bgr_9_0.V_TOP.t30 bgr_9_0.START_UP.t3 VDDA.t392 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X291 VOUT+.t70 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 VOUT-.t68 two_stage_opamp_dummy_magic_19_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X293 VOUT-.t69 two_stage_opamp_dummy_magic_19_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X294 VOUT+.t71 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 VOUT+.t72 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X296 bgr_9_0.V_TOP.t31 VDDA.t394 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X297 bgr_9_0.V_TOP.t4 bgr_9_0.1st_Vout_1.t21 VDDA.t134 VDDA.t133 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X298 GNDA.t82 two_stage_opamp_dummy_magic_19_0.X.t36 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t9 VDDA.t98 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X299 VOUT+.t73 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 VDDA.t311 VDDA.t309 GNDA.t290 VDDA.t310 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X301 VDDA.t317 VDDA.t315 two_stage_opamp_dummy_magic_19_0.VD3.t37 VDDA.t316 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X302 VOUT+.t1 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t4 GNDA.t19 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X303 two_stage_opamp_dummy_magic_19_0.X.t21 two_stage_opamp_dummy_magic_19_0.Vb2.t24 two_stage_opamp_dummy_magic_19_0.VD3.t5 two_stage_opamp_dummy_magic_19_0.VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X304 VDDA.t314 VDDA.t312 two_stage_opamp_dummy_magic_19_0.V_err_gate.t4 VDDA.t313 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X305 VOUT-.t70 two_stage_opamp_dummy_magic_19_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X306 two_stage_opamp_dummy_magic_19_0.X.t16 two_stage_opamp_dummy_magic_19_0.Vb1.t21 two_stage_opamp_dummy_magic_19_0.VD1.t9 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X307 VOUT-.t71 two_stage_opamp_dummy_magic_19_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X308 bgr_9_0.V_TOP.t6 bgr_9_0.1st_Vout_1.t22 VDDA.t175 VDDA.t174 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X309 two_stage_opamp_dummy_magic_19_0.Y.t20 two_stage_opamp_dummy_magic_19_0.Vb1.t22 two_stage_opamp_dummy_magic_19_0.VD2.t16 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X310 VOUT+.t74 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X311 VOUT+.t75 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X312 VOUT+.t76 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 bgr_9_0.NFET_GATE_10uA.t2 bgr_9_0.NFET_GATE_10uA.t1 GNDA.t174 GNDA.t173 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X314 GNDA.t172 bgr_9_0.NFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_19_0.Vb3.t3 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X315 VOUT+.t77 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 bgr_9_0.V_TOP.t32 VDDA.t395 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 VDDA.t299 VDDA.t297 VDDA.t299 VDDA.t298 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X318 two_stage_opamp_dummy_magic_19_0.VD4.t9 two_stage_opamp_dummy_magic_19_0.Vb2.t25 two_stage_opamp_dummy_magic_19_0.Y.t9 two_stage_opamp_dummy_magic_19_0.VD4.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X319 VDDA.t118 two_stage_opamp_dummy_magic_19_0.X.t37 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t5 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X320 bgr_9_0.1st_Vout_2.t20 bgr_9_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X321 VOUT-.t72 two_stage_opamp_dummy_magic_19_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X322 VOUT-.t73 two_stage_opamp_dummy_magic_19_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 VOUT-.t74 two_stage_opamp_dummy_magic_19_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X324 VOUT+.t78 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X325 two_stage_opamp_dummy_magic_19_0.VD1.t21 VIN-.t5 two_stage_opamp_dummy_magic_19_0.V_source.t40 GNDA.t309 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X326 GNDA.t261 GNDA.t260 two_stage_opamp_dummy_magic_19_0.Vb1.t9 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X327 VDDA.t364 bgr_9_0.PFET_GATE_10uA.t16 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t16 VDDA.t363 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X328 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t8 two_stage_opamp_dummy_magic_19_0.X.t38 GNDA.t297 VDDA.t369 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X329 VOUT-.t75 two_stage_opamp_dummy_magic_19_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 VDDA.t69 two_stage_opamp_dummy_magic_19_0.X.t39 VOUT-.t1 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X331 bgr_9_0.1st_Vout_1.t23 bgr_9_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X332 bgr_9_0.V_mir1.t10 bgr_9_0.V_mir1.t9 VDDA.t148 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X333 VOUT+.t6 two_stage_opamp_dummy_magic_19_0.Y.t37 VDDA.t111 VDDA.t110 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X334 GNDA.t62 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t15 two_stage_opamp_dummy_magic_19_0.V_source.t30 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X335 VDDA.t405 bgr_9_0.V_TOP.t33 bgr_9_0.START_UP.t2 VDDA.t404 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X336 two_stage_opamp_dummy_magic_19_0.V_p_mir.t1 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t16 GNDA.t3 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X337 VOUT-.t76 two_stage_opamp_dummy_magic_19_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X338 bgr_9_0.1st_Vout_2.t21 bgr_9_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X339 VOUT+.t79 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X340 VOUT+.t80 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X341 a_7460_23988.t1 a_7580_22380.t1 GNDA.t90 sky130_fd_pr__res_xhigh_po_0p35 l=6
X342 bgr_9_0.V_p_2.t7 bgr_9_0.V_CUR_REF_REG.t5 bgr_9_0.1st_Vout_2.t8 GNDA.t140 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X343 VOUT-.t77 two_stage_opamp_dummy_magic_19_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X344 VOUT+.t81 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 two_stage_opamp_dummy_magic_19_0.VD3.t3 two_stage_opamp_dummy_magic_19_0.Vb2.t26 two_stage_opamp_dummy_magic_19_0.X.t7 two_stage_opamp_dummy_magic_19_0.VD3.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X346 VOUT-.t9 GNDA.t257 GNDA.t259 GNDA.t258 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X347 a_14450_5524.t0 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t15 GNDA.t303 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X348 two_stage_opamp_dummy_magic_19_0.V_source.t29 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t17 GNDA.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X349 GNDA.t256 GNDA.t254 VDDA.t238 GNDA.t255 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X350 bgr_9_0.1st_Vout_2.t22 bgr_9_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 two_stage_opamp_dummy_magic_19_0.VD4.t7 two_stage_opamp_dummy_magic_19_0.Vb2.t27 two_stage_opamp_dummy_magic_19_0.Y.t8 two_stage_opamp_dummy_magic_19_0.VD4.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X352 bgr_9_0.1st_Vout_1.t9 bgr_9_0.Vin+.t8 bgr_9_0.V_p_1.t7 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X353 VDDA.t379 bgr_9_0.V_mir2.t20 bgr_9_0.1st_Vout_2.t10 VDDA.t378 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X354 two_stage_opamp_dummy_magic_19_0.VD4.t33 two_stage_opamp_dummy_magic_19_0.Vb3.t14 VDDA.t224 VDDA.t223 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X355 VOUT-.t78 two_stage_opamp_dummy_magic_19_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X356 VOUT-.t79 two_stage_opamp_dummy_magic_19_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X357 GNDA.t97 two_stage_opamp_dummy_magic_19_0.X.t40 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t7 VDDA.t130 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X358 bgr_9_0.1st_Vout_1.t24 bgr_9_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 GNDA.t197 GNDA.t196 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X360 bgr_9_0.NFET_GATE_10uA.t4 bgr_9_0.PFET_GATE_10uA.t17 VDDA.t366 VDDA.t365 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X361 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t8 two_stage_opamp_dummy_magic_19_0.Y.t38 GNDA.t17 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X362 VOUT-.t80 two_stage_opamp_dummy_magic_19_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 bgr_9_0.1st_Vout_2.t23 bgr_9_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 GNDA.t170 bgr_9_0.NFET_GATE_10uA.t15 two_stage_opamp_dummy_magic_19_0.Vb2.t5 GNDA.t169 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X365 two_stage_opamp_dummy_magic_19_0.Vb2.t4 bgr_9_0.NFET_GATE_10uA.t16 GNDA.t168 GNDA.t167 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X366 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t7 two_stage_opamp_dummy_magic_19_0.Y.t39 GNDA.t35 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X367 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t14 GNDA.t251 GNDA.t253 GNDA.t252 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X368 VOUT+.t82 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X369 GNDA.t199 GNDA.t250 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X370 GNDA.t249 GNDA.t247 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t14 GNDA.t248 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X371 GNDA.t246 GNDA.t244 two_stage_opamp_dummy_magic_19_0.Vb2.t10 GNDA.t245 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X372 two_stage_opamp_dummy_magic_19_0.V_source.t2 VIN+.t4 two_stage_opamp_dummy_magic_19_0.VD2.t2 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X373 VOUT-.t81 two_stage_opamp_dummy_magic_19_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X374 two_stage_opamp_dummy_magic_19_0.V_err_mir_p.t1 two_stage_opamp_dummy_magic_19_0.V_err_gate.t8 VDDA.t15 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X375 VOUT+.t83 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X376 bgr_9_0.PFET_GATE_10uA.t8 VDDA.t294 VDDA.t296 VDDA.t295 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X377 two_stage_opamp_dummy_magic_19_0.X.t14 two_stage_opamp_dummy_magic_19_0.Vb1.t23 two_stage_opamp_dummy_magic_19_0.VD1.t8 GNDA.t118 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X378 VOUT+.t84 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 bgr_9_0.1st_Vout_1.t2 bgr_9_0.V_mir1.t20 VDDA.t58 VDDA.t57 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X380 two_stage_opamp_dummy_magic_19_0.X.t1 two_stage_opamp_dummy_magic_19_0.Vb1.t24 two_stage_opamp_dummy_magic_19_0.VD1.t7 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X381 two_stage_opamp_dummy_magic_19_0.Vb2_2.t2 two_stage_opamp_dummy_magic_19_0.Vb2.t28 VDDA.t399 VDDA.t398 sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.36 ps=2.2 w=1.8 l=0.2
X382 VOUT-.t82 two_stage_opamp_dummy_magic_19_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 two_stage_opamp_dummy_magic_19_0.Y.t24 two_stage_opamp_dummy_magic_19_0.Vb1.t25 two_stage_opamp_dummy_magic_19_0.VD2.t21 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X384 bgr_9_0.V_p_2.t6 bgr_9_0.V_CUR_REF_REG.t6 bgr_9_0.1st_Vout_2.t0 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X385 VOUT-.t83 two_stage_opamp_dummy_magic_19_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X386 VOUT+.t85 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X387 GNDA.t199 GNDA.t243 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X388 VOUT-.t84 two_stage_opamp_dummy_magic_19_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X389 VDDA.t93 two_stage_opamp_dummy_magic_19_0.X.t41 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t4 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X390 VOUT+.t86 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X391 GNDA.t199 GNDA.t242 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X392 VOUT-.t85 two_stage_opamp_dummy_magic_19_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X393 two_stage_opamp_dummy_magic_19_0.VD1.t2 VIN-.t6 two_stage_opamp_dummy_magic_19_0.V_source.t5 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X394 GNDA.t29 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t5 VOUT+.t2 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X395 a_5540_5524.t1 two_stage_opamp_dummy_magic_19_0.V_tot.t0 GNDA.t88 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X396 VDDA.t368 bgr_9_0.V_mir2.t6 bgr_9_0.V_mir2.t7 VDDA.t367 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X397 two_stage_opamp_dummy_magic_19_0.VD2.t0 VIN+.t5 two_stage_opamp_dummy_magic_19_0.V_source.t1 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X398 VDDA.t222 two_stage_opamp_dummy_magic_19_0.Vb3.t15 two_stage_opamp_dummy_magic_19_0.VD4.t32 VDDA.t221 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X399 VOUT+.t18 two_stage_opamp_dummy_magic_19_0.Y.t40 VDDA.t385 VDDA.t384 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X400 VOUT+.t87 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 VOUT+.t88 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X402 VOUT+.t89 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 GNDA.t137 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t18 two_stage_opamp_dummy_magic_19_0.V_source.t28 GNDA.t136 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X404 GNDA.t241 GNDA.t240 two_stage_opamp_dummy_magic_19_0.err_amp_out.t2 GNDA.t143 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X405 VOUT+.t90 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 VDDA.t21 bgr_9_0.PFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_19_0.Vb1.t0 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X407 bgr_9_0.V_p_2.t5 bgr_9_0.V_CUR_REF_REG.t7 bgr_9_0.1st_Vout_2.t1 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X408 two_stage_opamp_dummy_magic_19_0.VD4.t25 two_stage_opamp_dummy_magic_19_0.VD4.t23 two_stage_opamp_dummy_magic_19_0.Y.t15 two_stage_opamp_dummy_magic_19_0.VD4.t24 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X409 VOUT+.t91 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 a_13180_23838.t0 bgr_9_0.V_CUR_REF_REG.t0 GNDA.t44 sky130_fd_pr__res_xhigh_po_0p35 l=4
X411 two_stage_opamp_dummy_magic_19_0.VD3.t32 two_stage_opamp_dummy_magic_19_0.Vb3.t16 VDDA.t220 VDDA.t219 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X412 VOUT-.t86 two_stage_opamp_dummy_magic_19_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X413 bgr_9_0.V_TOP.t34 VDDA.t406 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 VOUT-.t87 two_stage_opamp_dummy_magic_19_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X415 VOUT-.t88 two_stage_opamp_dummy_magic_19_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 VOUT-.t89 two_stage_opamp_dummy_magic_19_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 VOUT-.t90 two_stage_opamp_dummy_magic_19_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X418 two_stage_opamp_dummy_magic_19_0.V_source.t27 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t19 GNDA.t139 GNDA.t138 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X419 VOUT-.t91 two_stage_opamp_dummy_magic_19_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X420 GNDA.t296 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t6 VOUT+.t17 GNDA.t295 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X421 VOUT+.t92 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X422 bgr_9_0.V_TOP.t35 VDDA.t407 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t3 two_stage_opamp_dummy_magic_19_0.X.t42 VDDA.t169 GNDA.t121 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X424 VDDA.t120 bgr_9_0.1st_Vout_2.t24 bgr_9_0.PFET_GATE_10uA.t3 VDDA.t119 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X425 two_stage_opamp_dummy_magic_19_0.err_amp_out.t0 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t8 two_stage_opamp_dummy_magic_19_0.V_err_p.t3 VDDA.t48 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X426 GNDA.t239 GNDA.t238 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t1 GNDA.t143 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X427 VOUT+.t93 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 VDDA.t387 two_stage_opamp_dummy_magic_19_0.Y.t41 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t5 GNDA.t305 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X429 VOUT-.t92 two_stage_opamp_dummy_magic_19_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X430 VOUT+.t94 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t6 two_stage_opamp_dummy_magic_19_0.Y.t42 GNDA.t147 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X432 VOUT+.t95 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 VOUT+.t96 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t2 bgr_9_0.PFET_GATE_10uA.t19 VDDA.t100 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X435 two_stage_opamp_dummy_magic_19_0.VD3.t25 two_stage_opamp_dummy_magic_19_0.VD3.t23 two_stage_opamp_dummy_magic_19_0.X.t12 two_stage_opamp_dummy_magic_19_0.VD3.t24 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X436 VOUT-.t93 two_stage_opamp_dummy_magic_19_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 VOUT-.t94 two_stage_opamp_dummy_magic_19_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 VDDA.t42 bgr_9_0.PFET_GATE_10uA.t20 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t0 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X439 VOUT-.t95 two_stage_opamp_dummy_magic_19_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 VOUT-.t96 two_stage_opamp_dummy_magic_19_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 two_stage_opamp_dummy_magic_19_0.V_err_mir_p.t3 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t9 two_stage_opamp_dummy_magic_19_0.V_err_gate.t1 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X442 two_stage_opamp_dummy_magic_19_0.X.t19 GNDA.t236 GNDA.t237 GNDA.t228 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X443 two_stage_opamp_dummy_magic_19_0.cap_res_X.t138 two_stage_opamp_dummy_magic_19_0.X.t17 GNDA.t145 sky130_fd_pr__res_high_po_1p41 l=1.41
X444 VOUT-.t97 two_stage_opamp_dummy_magic_19_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 bgr_9_0.V_TOP.t36 VDDA.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X446 VOUT-.t98 two_stage_opamp_dummy_magic_19_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X447 two_stage_opamp_dummy_magic_19_0.Y.t19 two_stage_opamp_dummy_magic_19_0.Vb1.t26 two_stage_opamp_dummy_magic_19_0.VD2.t13 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X448 bgr_9_0.Vin-.t5 bgr_9_0.V_TOP.t37 VDDA.t123 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X449 two_stage_opamp_dummy_magic_19_0.Y.t3 two_stage_opamp_dummy_magic_19_0.Vb2.t29 two_stage_opamp_dummy_magic_19_0.VD4.t5 two_stage_opamp_dummy_magic_19_0.VD4.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X450 VOUT-.t99 two_stage_opamp_dummy_magic_19_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X451 VDDA.t293 VDDA.t290 VDDA.t292 VDDA.t291 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0 ps=0 w=1.8 l=0.2
X452 VOUT+.t97 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X453 VOUT+.t98 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X454 VDDA.t218 two_stage_opamp_dummy_magic_19_0.Vb3.t17 two_stage_opamp_dummy_magic_19_0.VD4.t31 VDDA.t217 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X455 VOUT+.t99 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 GNDA.t166 bgr_9_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t13 GNDA.t165 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X457 bgr_9_0.1st_Vout_1.t1 bgr_9_0.V_mir1.t21 VDDA.t60 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X458 two_stage_opamp_dummy_magic_19_0.Vb2.t9 GNDA.t233 GNDA.t235 GNDA.t234 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X459 VOUT+.t100 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 VOUT+.t101 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 VOUT+.t102 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 bgr_9_0.1st_Vout_1.t25 bgr_9_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 VOUT-.t100 two_stage_opamp_dummy_magic_19_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X464 bgr_9_0.1st_Vout_2.t25 bgr_9_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X465 two_stage_opamp_dummy_magic_19_0.VD1.t18 VIN-.t7 two_stage_opamp_dummy_magic_19_0.V_source.t16 GNDA.t118 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X466 VDDA.t168 two_stage_opamp_dummy_magic_19_0.X.t43 VOUT-.t8 VDDA.t167 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X467 VOUT+.t103 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X468 two_stage_opamp_dummy_magic_19_0.VD1.t3 VIN-.t8 two_stage_opamp_dummy_magic_19_0.V_source.t8 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X469 two_stage_opamp_dummy_magic_19_0.VD2.t3 VIN+.t6 two_stage_opamp_dummy_magic_19_0.V_source.t3 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X470 VOUT-.t101 two_stage_opamp_dummy_magic_19_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X471 VOUT+.t3 two_stage_opamp_dummy_magic_19_0.Y.t43 VDDA.t30 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X472 GNDA.t70 two_stage_opamp_dummy_magic_19_0.err_amp_mir.t1 two_stage_opamp_dummy_magic_19_0.err_amp_mir.t2 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X473 bgr_9_0.1st_Vout_1.t26 bgr_9_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 GNDA.t142 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t20 two_stage_opamp_dummy_magic_19_0.V_source.t26 GNDA.t141 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X475 VOUT-.t102 two_stage_opamp_dummy_magic_19_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X476 VOUT-.t103 two_stage_opamp_dummy_magic_19_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X477 VOUT-.t104 two_stage_opamp_dummy_magic_19_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X478 a_14450_5524.t1 two_stage_opamp_dummy_magic_19_0.V_tot.t3 GNDA.t310 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X479 VOUT-.t105 two_stage_opamp_dummy_magic_19_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X480 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t4 bgr_9_0.V_TOP.t38 VDDA.t125 VDDA.t124 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X481 VOUT+.t104 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 VDDA.t1 bgr_9_0.V_mir2.t4 bgr_9_0.V_mir2.t5 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X483 VOUT+.t105 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X484 VDDA.t173 bgr_9_0.V_mir1.t7 bgr_9_0.V_mir1.t8 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X485 VDDA.t289 VDDA.t286 VDDA.t288 VDDA.t287 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.15
X486 two_stage_opamp_dummy_magic_19_0.V_source.t25 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t21 GNDA.t144 GNDA.t143 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X487 bgr_9_0.V_p_1.t2 bgr_9_0.Vin-.t10 bgr_9_0.V_mir1.t0 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X488 VDDA.t216 two_stage_opamp_dummy_magic_19_0.Vb3.t18 two_stage_opamp_dummy_magic_19_0.VD4.t30 VDDA.t215 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X489 two_stage_opamp_dummy_magic_19_0.Vb2.t0 two_stage_opamp_dummy_magic_19_0.Vb2_2.t6 two_stage_opamp_dummy_magic_19_0.Vb2_2.t8 two_stage_opamp_dummy_magic_19_0.Vb2_2.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X490 VOUT+.t106 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X491 bgr_9_0.1st_Vout_1.t27 bgr_9_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X492 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t2 two_stage_opamp_dummy_magic_19_0.X.t44 VDDA.t144 GNDA.t101 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X493 bgr_9_0.1st_Vout_2.t26 bgr_9_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X494 VDDA.t189 two_stage_opamp_dummy_magic_19_0.Y.t44 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t4 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X495 VDDA.t56 two_stage_opamp_dummy_magic_19_0.V_err_gate.t9 two_stage_opamp_dummy_magic_19_0.V_err_p.t1 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X496 two_stage_opamp_dummy_magic_19_0.V_p_mir.t4 VIN+.t7 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t3 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X497 GNDA.t315 two_stage_opamp_dummy_magic_19_0.X.t45 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t6 VDDA.t410 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X498 VOUT+.t107 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X499 VOUT+.t108 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X500 bgr_9_0.V_TOP.t9 VDDA.t283 VDDA.t285 VDDA.t284 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X501 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t5 two_stage_opamp_dummy_magic_19_0.Y.t45 GNDA.t46 VDDA.t50 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X502 VOUT+.t109 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X503 bgr_9_0.1st_Vout_1.t28 bgr_9_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X504 two_stage_opamp_dummy_magic_19_0.V_source.t24 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t22 GNDA.t108 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X505 VOUT-.t106 two_stage_opamp_dummy_magic_19_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X506 VDDA.t282 VDDA.t280 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t2 VDDA.t281 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X507 VDDA.t279 VDDA.t277 two_stage_opamp_dummy_magic_19_0.Vb2_2.t9 VDDA.t278 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.36 ps=2.2 w=1.8 l=0.2
X508 bgr_9_0.V_p_1.t1 bgr_9_0.Vin-.t11 bgr_9_0.V_mir1.t13 GNDA.t130 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X509 VOUT+.t110 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 VOUT-.t107 two_stage_opamp_dummy_magic_19_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 VOUT+.t111 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X512 VOUT+.t112 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X513 VOUT+.t113 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X514 bgr_9_0.1st_Vout_1.t29 bgr_9_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X515 two_stage_opamp_dummy_magic_19_0.Vb3.t0 GNDA.t230 GNDA.t232 GNDA.t231 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X516 VOUT+.t114 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X517 bgr_9_0.Vin-.t7 bgr_9_0.START_UP.t6 bgr_9_0.V_TOP.t12 VDDA.t386 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X518 two_stage_opamp_dummy_magic_19_0.Y.t17 two_stage_opamp_dummy_magic_19_0.Vb1.t27 two_stage_opamp_dummy_magic_19_0.VD2.t11 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X519 bgr_9_0.V_TOP.t0 bgr_9_0.START_UP.t7 bgr_9_0.Vin-.t0 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X520 VOUT-.t108 two_stage_opamp_dummy_magic_19_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X521 VOUT+.t115 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X522 VOUT+.t116 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 VDDA.t154 bgr_9_0.1st_Vout_2.t27 bgr_9_0.PFET_GATE_10uA.t2 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X524 bgr_9_0.V_mir1.t6 bgr_9_0.V_mir1.t5 VDDA.t389 VDDA.t388 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X525 VOUT-.t109 two_stage_opamp_dummy_magic_19_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X526 a_5540_5524.t0 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t1 GNDA.t21 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X527 VOUT-.t110 two_stage_opamp_dummy_magic_19_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 VOUT-.t111 two_stage_opamp_dummy_magic_19_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X529 GNDA.t199 GNDA.t222 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X530 bgr_9_0.START_UP.t1 bgr_9_0.START_UP.t0 bgr_9_0.START_UP_NFET1.t0 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X531 two_stage_opamp_dummy_magic_19_0.VD4.t29 two_stage_opamp_dummy_magic_19_0.Vb3.t19 VDDA.t214 VDDA.t213 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X532 bgr_9_0.V_p_2.t3 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t10 bgr_9_0.V_mir2.t15 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X533 two_stage_opamp_dummy_magic_19_0.VD1.t20 GNDA.t227 GNDA.t229 GNDA.t228 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X534 VOUT+.t16 VDDA.t274 VDDA.t276 VDDA.t275 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X535 VOUT+.t8 two_stage_opamp_dummy_magic_19_0.Y.t46 VDDA.t137 VDDA.t136 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X536 two_stage_opamp_dummy_magic_19_0.VD2.t6 VIN+.t8 two_stage_opamp_dummy_magic_19_0.V_source.t6 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X537 GNDA.t226 GNDA.t223 GNDA.t225 GNDA.t224 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X538 GNDA.t221 GNDA.t220 two_stage_opamp_dummy_magic_19_0.X.t18 GNDA.t218 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X539 VOUT+.t117 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X540 VOUT+.t118 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X541 VDDA.t212 two_stage_opamp_dummy_magic_19_0.Vb3.t20 two_stage_opamp_dummy_magic_19_0.VD3.t31 VDDA.t211 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X542 VOUT-.t112 two_stage_opamp_dummy_magic_19_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X543 bgr_9_0.1st_Vout_2.t28 bgr_9_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X544 VOUT-.t113 two_stage_opamp_dummy_magic_19_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X545 VOUT+.t119 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X546 two_stage_opamp_dummy_magic_19_0.Vb1_2.t2 two_stage_opamp_dummy_magic_19_0.Vb1.t5 two_stage_opamp_dummy_magic_19_0.Vb1.t6 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X547 VDDA.t162 bgr_9_0.V_mir2.t21 bgr_9_0.1st_Vout_2.t6 VDDA.t161 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X548 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t0 bgr_9_0.PFET_GATE_10uA.t21 VDDA.t143 VDDA.t142 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X549 VOUT-.t114 two_stage_opamp_dummy_magic_19_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X550 bgr_9_0.V_p_1.t0 bgr_9_0.Vin-.t12 bgr_9_0.V_mir1.t15 GNDA.t289 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X551 GNDA.t199 GNDA.t214 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X552 bgr_9_0.1st_Vout_2.t29 bgr_9_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X553 VOUT-.t115 two_stage_opamp_dummy_magic_19_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X554 VOUT-.t116 two_stage_opamp_dummy_magic_19_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X555 two_stage_opamp_dummy_magic_19_0.V_source.t23 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t23 GNDA.t109 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X556 VOUT+.t120 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X557 VDDA.t135 two_stage_opamp_dummy_magic_19_0.Y.t47 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t3 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X558 two_stage_opamp_dummy_magic_19_0.err_amp_mir.t4 VDDA.t271 VDDA.t273 VDDA.t272 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X559 VOUT-.t117 two_stage_opamp_dummy_magic_19_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X560 VOUT+.t121 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 bgr_9_0.1st_Vout_1.t30 bgr_9_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X562 GNDA.t197 GNDA.t216 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X563 GNDA.t292 VDDA.t268 VDDA.t270 VDDA.t269 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X564 a_6810_23838.t0 a_6930_22564.t0 GNDA.t75 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X565 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t4 two_stage_opamp_dummy_magic_19_0.Y.t48 GNDA.t129 VDDA.t184 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X566 VOUT+.t122 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X567 GNDA.t199 GNDA.t215 bgr_9_0.Vin-.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X568 VOUT+.t123 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X569 bgr_9_0.1st_Vout_2.t30 bgr_9_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 VOUT+.t124 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X571 GNDA.t164 bgr_9_0.NFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_19_0.V_err_gate.t2 GNDA.t163 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X572 bgr_9_0.Vin-.t4 bgr_9_0.V_TOP.t39 VDDA.t26 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X573 a_12530_23988.t1 a_12410_22380.t0 GNDA.t306 sky130_fd_pr__res_xhigh_po_0p35 l=6
X574 two_stage_opamp_dummy_magic_19_0.Vb3.t7 bgr_9_0.NFET_GATE_10uA.t19 GNDA.t162 GNDA.t161 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X575 two_stage_opamp_dummy_magic_19_0.VD4.t28 two_stage_opamp_dummy_magic_19_0.Vb3.t21 VDDA.t210 VDDA.t209 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X576 bgr_9_0.1st_Vout_2.t31 bgr_9_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X577 VOUT-.t118 two_stage_opamp_dummy_magic_19_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X578 VDDA.t129 bgr_9_0.V_mir2.t2 bgr_9_0.V_mir2.t3 VDDA.t128 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X579 VOUT+.t125 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X580 bgr_9_0.1st_Vout_1.t31 bgr_9_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X581 bgr_9_0.1st_Vout_2.t32 bgr_9_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X582 bgr_9_0.V_p_1.t10 VDDA.t413 GNDA.t152 GNDA.t151 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X583 VDDA.t208 two_stage_opamp_dummy_magic_19_0.Vb3.t22 two_stage_opamp_dummy_magic_19_0.VD3.t30 VDDA.t207 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X584 VDDA.t267 VDDA.t265 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t14 VDDA.t266 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X585 VOUT+.t126 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X586 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t13 bgr_9_0.PFET_GATE_10uA.t22 VDDA.t194 VDDA.t193 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X587 VOUT-.t119 two_stage_opamp_dummy_magic_19_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X588 VOUT-.t120 two_stage_opamp_dummy_magic_19_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X589 a_13180_23838.t1 a_13060_22630.t0 GNDA.t65 sky130_fd_pr__res_xhigh_po_0p35 l=4
X590 VDDA.t115 two_stage_opamp_dummy_magic_19_0.X.t46 VOUT-.t4 VDDA.t114 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X591 VOUT+.t127 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X592 a_14330_5524.t1 two_stage_opamp_dummy_magic_19_0.V_tot.t1 GNDA.t132 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X593 VOUT+.t128 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X594 VOUT+.t129 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X595 two_stage_opamp_dummy_magic_19_0.VD2.t9 VIN+.t9 two_stage_opamp_dummy_magic_19_0.V_source.t10 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X596 two_stage_opamp_dummy_magic_19_0.VD1.t6 two_stage_opamp_dummy_magic_19_0.Vb1.t28 two_stage_opamp_dummy_magic_19_0.X.t6 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X597 bgr_9_0.V_p_1.t6 bgr_9_0.Vin+.t9 bgr_9_0.1st_Vout_1.t8 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X598 VDDA.t132 bgr_9_0.V_mir1.t22 bgr_9_0.1st_Vout_1.t0 VDDA.t131 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X599 bgr_9_0.V_TOP.t40 VDDA.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X600 two_stage_opamp_dummy_magic_19_0.VD4.t27 two_stage_opamp_dummy_magic_19_0.Vb3.t23 VDDA.t206 VDDA.t205 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X601 two_stage_opamp_dummy_magic_19_0.Vb2_2.t1 two_stage_opamp_dummy_magic_19_0.Vb2.t1 two_stage_opamp_dummy_magic_19_0.Vb2.t2 two_stage_opamp_dummy_magic_19_0.Vb2_2.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X602 VOUT-.t121 two_stage_opamp_dummy_magic_19_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X603 VOUT-.t122 two_stage_opamp_dummy_magic_19_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X604 VOUT-.t123 two_stage_opamp_dummy_magic_19_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X605 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t1 two_stage_opamp_dummy_magic_19_0.X.t47 VDDA.t39 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X606 VOUT-.t124 two_stage_opamp_dummy_magic_19_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X607 VDDA.t49 two_stage_opamp_dummy_magic_19_0.Y.t49 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t2 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X608 GNDA.t219 GNDA.t217 two_stage_opamp_dummy_magic_19_0.VD1.t19 GNDA.t218 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X609 VOUT+.t130 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X610 VOUT+.t131 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X611 VDDA.t80 bgr_9_0.PFET_GATE_10uA.t23 bgr_9_0.V_CUR_REF_REG.t1 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X612 VOUT-.t17 two_stage_opamp_dummy_magic_19_0.X.t48 VDDA.t377 VDDA.t376 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X613 GNDA.t52 two_stage_opamp_dummy_magic_19_0.X.t49 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t5 VDDA.t65 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X614 bgr_9_0.V_TOP.t41 VDDA.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X615 bgr_9_0.V_p_1.t5 bgr_9_0.Vin+.t10 bgr_9_0.1st_Vout_1.t7 GNDA.t95 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X616 VDDA.t264 VDDA.t262 bgr_9_0.V_TOP.t8 VDDA.t263 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X617 VOUT-.t125 two_stage_opamp_dummy_magic_19_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X618 two_stage_opamp_dummy_magic_19_0.Vb2.t3 bgr_9_0.NFET_GATE_10uA.t20 GNDA.t160 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X619 GNDA.t158 bgr_9_0.NFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t11 GNDA.t157 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X620 VOUT-.t126 two_stage_opamp_dummy_magic_19_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X621 VOUT-.t127 two_stage_opamp_dummy_magic_19_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X622 two_stage_opamp_dummy_magic_19_0.VD3.t36 VDDA.t259 VDDA.t261 VDDA.t260 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X623 VDDA.t258 VDDA.t256 VOUT+.t15 VDDA.t257 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X624 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t12 bgr_9_0.NFET_GATE_10uA.t22 GNDA.t156 GNDA.t155 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X625 bgr_9_0.V_TOP.t42 VDDA.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X626 VOUT-.t6 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t7 GNDA.t107 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X627 bgr_9_0.V_TOP.t43 VDDA.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X628 VOUT-.t128 two_stage_opamp_dummy_magic_19_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X629 two_stage_opamp_dummy_magic_19_0.Vb1.t4 two_stage_opamp_dummy_magic_19_0.Vb1.t3 two_stage_opamp_dummy_magic_19_0.Vb1_2.t1 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X630 VOUT-.t129 two_stage_opamp_dummy_magic_19_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X631 VDDA.t186 bgr_9_0.V_mir2.t22 bgr_9_0.1st_Vout_2.t7 VDDA.t185 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X632 two_stage_opamp_dummy_magic_19_0.VD4.t3 two_stage_opamp_dummy_magic_19_0.Vb2.t30 two_stage_opamp_dummy_magic_19_0.Y.t5 two_stage_opamp_dummy_magic_19_0.VD4.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X633 two_stage_opamp_dummy_magic_19_0.Y.t14 two_stage_opamp_dummy_magic_19_0.Vb1.t29 two_stage_opamp_dummy_magic_19_0.VD2.t5 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X634 VOUT-.t130 two_stage_opamp_dummy_magic_19_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X635 VDDA.t150 bgr_9_0.1st_Vout_1.t32 bgr_9_0.V_TOP.t5 VDDA.t149 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X636 VOUT+.t132 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X637 VOUT-.t131 two_stage_opamp_dummy_magic_19_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X638 VOUT-.t132 two_stage_opamp_dummy_magic_19_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X639 GNDA.t213 GNDA.t211 two_stage_opamp_dummy_magic_19_0.V_source.t38 GNDA.t212 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X640 a_5420_5524.t0 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t0 GNDA.t64 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X641 VOUT+.t133 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X642 VOUT+.t134 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X643 VDDA.t255 VDDA.t253 GNDA.t293 VDDA.t254 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X644 bgr_9_0.V_TOP.t44 VDDA.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X645 VOUT-.t15 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t8 GNDA.t299 GNDA.t298 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X646 two_stage_opamp_dummy_magic_19_0.VD3.t29 two_stage_opamp_dummy_magic_19_0.Vb3.t24 VDDA.t204 VDDA.t203 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X647 VOUT-.t133 two_stage_opamp_dummy_magic_19_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X648 VDDA.t18 two_stage_opamp_dummy_magic_19_0.X.t50 VOUT-.t0 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X649 two_stage_opamp_dummy_magic_19_0.VD3.t1 two_stage_opamp_dummy_magic_19_0.Vb2.t31 two_stage_opamp_dummy_magic_19_0.X.t20 two_stage_opamp_dummy_magic_19_0.VD3.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X650 bgr_9_0.V_TOP.t45 VDDA.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X651 bgr_9_0.V_mir2.t1 bgr_9_0.V_mir2.t0 VDDA.t95 VDDA.t94 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X652 VDDA.t127 bgr_9_0.V_mir1.t3 bgr_9_0.V_mir1.t4 VDDA.t126 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X653 two_stage_opamp_dummy_magic_19_0.Vb1.t11 VDDA.t250 VDDA.t252 VDDA.t251 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X654 VOUT-.t134 two_stage_opamp_dummy_magic_19_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X655 two_stage_opamp_dummy_magic_19_0.VD1.t5 two_stage_opamp_dummy_magic_19_0.Vb1.t30 two_stage_opamp_dummy_magic_19_0.X.t15 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X656 VOUT-.t135 two_stage_opamp_dummy_magic_19_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X657 VOUT-.t136 two_stage_opamp_dummy_magic_19_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X658 bgr_9_0.V_mir2.t14 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t11 bgr_9_0.V_p_2.t0 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X659 VOUT+.t135 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X660 VOUT+.t136 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X661 bgr_9_0.PFET_GATE_10uA.t7 VDDA.t414 GNDA.t313 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X662 VOUT+.t137 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X663 bgr_9_0.1st_Vout_1.t33 bgr_9_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X664 two_stage_opamp_dummy_magic_19_0.VD3.t28 two_stage_opamp_dummy_magic_19_0.Vb3.t25 VDDA.t202 VDDA.t201 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X665 VOUT-.t137 two_stage_opamp_dummy_magic_19_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X666 VDDA.t45 bgr_9_0.V_TOP.t46 bgr_9_0.Vin-.t3 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X667 VDDA.t237 GNDA.t208 GNDA.t210 GNDA.t209 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X668 VDDA.t16 two_stage_opamp_dummy_magic_19_0.Y.t50 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t1 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X669 VOUT+.t138 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X670 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t0 a_5820_2720.t0 GNDA.t126 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X671 two_stage_opamp_dummy_magic_19_0.V_source.t13 VIN-.t9 two_stage_opamp_dummy_magic_19_0.VD1.t16 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X672 VOUT-.t138 two_stage_opamp_dummy_magic_19_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X673 bgr_9_0.PFET_GATE_10uA.t1 bgr_9_0.1st_Vout_2.t33 VDDA.t77 VDDA.t76 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X674 VOUT-.t14 two_stage_opamp_dummy_magic_19_0.X.t51 VDDA.t373 VDDA.t372 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X675 GNDA.t31 two_stage_opamp_dummy_magic_19_0.X.t52 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t4 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X676 VOUT+.t139 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X677 VDDA.t75 bgr_9_0.PFET_GATE_10uA.t24 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t1 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X678 VDDA.t5 two_stage_opamp_dummy_magic_19_0.Y.t51 VOUT+.t0 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X679 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t13 VDDA.t247 VDDA.t249 VDDA.t248 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X680 GNDA.t207 GNDA.t206 two_stage_opamp_dummy_magic_19_0.V_p_mir.t2 GNDA.t143 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X681 VOUT-.t139 two_stage_opamp_dummy_magic_19_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X682 VDDA.t188 two_stage_opamp_dummy_magic_19_0.Y.t52 VOUT+.t12 VDDA.t187 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X683 VDDA.t200 two_stage_opamp_dummy_magic_19_0.Vb3.t26 two_stage_opamp_dummy_magic_19_0.VD4.t26 VDDA.t199 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X684 VOUT-.t140 two_stage_opamp_dummy_magic_19_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X685 VOUT+.t140 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X686 VDDA.t152 bgr_9_0.1st_Vout_2.t34 bgr_9_0.PFET_GATE_10uA.t0 VDDA.t151 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X687 VOUT+.t141 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X688 VOUT+.t142 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X689 GNDA.t205 GNDA.t203 VOUT+.t13 GNDA.t204 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X690 two_stage_opamp_dummy_magic_19_0.Y.t21 GNDA.t200 GNDA.t202 GNDA.t201 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X691 VOUT+.t143 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X692 VOUT+.t144 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X693 bgr_9_0.1st_Vout_1.t34 bgr_9_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X694 GNDA.t111 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t24 two_stage_opamp_dummy_magic_19_0.V_source.t22 GNDA.t110 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X695 bgr_9_0.1st_Vout_2.t35 bgr_9_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X696 VOUT-.t141 two_stage_opamp_dummy_magic_19_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X697 GNDA.t113 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t25 two_stage_opamp_dummy_magic_19_0.V_source.t21 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X698 bgr_9_0.V_mir2.t13 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t12 bgr_9_0.V_p_2.t1 GNDA.t63 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X699 two_stage_opamp_dummy_magic_19_0.VD3.t27 two_stage_opamp_dummy_magic_19_0.Vb3.t27 VDDA.t198 VDDA.t197 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X700 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t11 bgr_9_0.NFET_GATE_10uA.t23 GNDA.t154 GNDA.t153 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X701 VOUT-.t142 two_stage_opamp_dummy_magic_19_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X702 VOUT-.t143 two_stage_opamp_dummy_magic_19_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X703 GNDA.t199 GNDA.t198 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X704 VOUT-.t144 two_stage_opamp_dummy_magic_19_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X705 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t3 two_stage_opamp_dummy_magic_19_0.X.t53 GNDA.t122 VDDA.t170 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X706 VOUT+.t145 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X707 bgr_9_0.1st_Vout_1.t35 bgr_9_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X708 VOUT-.t145 two_stage_opamp_dummy_magic_19_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X709 VDDA.t89 bgr_9_0.1st_Vout_1.t36 bgr_9_0.V_TOP.t1 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X710 GNDA.t80 two_stage_opamp_dummy_magic_19_0.Y.t53 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t3 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X711 GNDA.t314 VDDA.t415 bgr_9_0.V_TOP.t7 GNDA.t289 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X712 bgr_9_0.V_TOP.t47 VDDA.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X713 two_stage_opamp_dummy_magic_19_0.VD2.t15 VIN+.t10 two_stage_opamp_dummy_magic_19_0.V_source.t18 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X714 VOUT-.t146 two_stage_opamp_dummy_magic_19_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X715 VDDA.t108 bgr_9_0.V_TOP.t48 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t3 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X716 VDDA.t246 VDDA.t244 two_stage_opamp_dummy_magic_19_0.VD4.t36 VDDA.t245 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X717 two_stage_opamp_dummy_magic_19_0.V_err_gate.t0 two_stage_opamp_dummy_magic_19_0.V_tot.t5 two_stage_opamp_dummy_magic_19_0.V_err_mir_p.t0 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X718 VOUT+.t146 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X719 VOUT+.t147 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X720 VOUT+.t148 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X721 VOUT-.t147 two_stage_opamp_dummy_magic_19_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X722 two_stage_opamp_dummy_magic_19_0.Vb2_2.t5 two_stage_opamp_dummy_magic_19_0.Vb2_2.t3 two_stage_opamp_dummy_magic_19_0.Vb2_2.t5 two_stage_opamp_dummy_magic_19_0.Vb2_2.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X723 two_stage_opamp_dummy_magic_19_0.Y.t12 two_stage_opamp_dummy_magic_19_0.VD4.t20 two_stage_opamp_dummy_magic_19_0.VD4.t22 two_stage_opamp_dummy_magic_19_0.VD4.t21 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X724 two_stage_opamp_dummy_magic_19_0.VD1.t4 two_stage_opamp_dummy_magic_19_0.Vb1.t31 two_stage_opamp_dummy_magic_19_0.X.t24 GNDA.t102 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X725 VOUT-.t148 two_stage_opamp_dummy_magic_19_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X726 bgr_9_0.V_mir2.t12 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t13 bgr_9_0.V_p_2.t2 GNDA.t78 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X727 two_stage_opamp_dummy_magic_19_0.VD2.t12 two_stage_opamp_dummy_magic_19_0.Vb1.t32 two_stage_opamp_dummy_magic_19_0.Y.t18 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X728 VOUT+.t149 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X729 VOUT+.t150 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X730 VOUT-.t149 two_stage_opamp_dummy_magic_19_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X731 VOUT+.t151 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X732 VOUT-.t150 two_stage_opamp_dummy_magic_19_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X733 VOUT-.t151 two_stage_opamp_dummy_magic_19_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X734 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t0 two_stage_opamp_dummy_magic_19_0.X.t54 VDDA.t78 GNDA.t69 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X735 VOUT+.t152 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X736 VOUT-.t152 two_stage_opamp_dummy_magic_19_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X737 GNDA.t105 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t9 VOUT-.t5 GNDA.t104 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X738 VOUT-.t153 two_stage_opamp_dummy_magic_19_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X739 VDDA.t196 two_stage_opamp_dummy_magic_19_0.Vb3.t28 two_stage_opamp_dummy_magic_19_0.VD3.t26 VDDA.t195 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X740 two_stage_opamp_dummy_magic_19_0.V_source.t12 VIN-.t10 two_stage_opamp_dummy_magic_19_0.VD1.t15 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X741 bgr_9_0.V_TOP.t49 VDDA.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X742 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t1 VDDA.t241 VDDA.t243 VDDA.t242 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X743 two_stage_opamp_dummy_magic_19_0.X.t9 two_stage_opamp_dummy_magic_19_0.VD3.t20 two_stage_opamp_dummy_magic_19_0.VD3.t22 two_stage_opamp_dummy_magic_19_0.VD3.t21 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X744 VOUT+.t153 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X745 VDDA.t166 two_stage_opamp_dummy_magic_19_0.Y.t54 VOUT+.t9 VDDA.t165 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X746 VOUT-.t154 two_stage_opamp_dummy_magic_19_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X747 VOUT+.t154 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X748 VOUT-.t155 two_stage_opamp_dummy_magic_19_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X749 bgr_9_0.1st_Vout_2.t36 bgr_9_0.cap_res2.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X750 two_stage_opamp_dummy_magic_19_0.V_source.t20 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t26 GNDA.t10 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X751 GNDA.t12 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t27 two_stage_opamp_dummy_magic_19_0.V_p_mir.t0 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X752 VDDA.t401 bgr_9_0.V_mir1.t1 bgr_9_0.V_mir1.t2 VDDA.t400 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X753 VOUT+.t155 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X754 two_stage_opamp_dummy_magic_19_0.Y.t6 two_stage_opamp_dummy_magic_19_0.Vb2.t32 two_stage_opamp_dummy_magic_19_0.VD4.t1 two_stage_opamp_dummy_magic_19_0.VD4.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X755 VOUT+.t156 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X756 VOUT-.t156 two_stage_opamp_dummy_magic_19_0.cap_res_X.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 bgr_9_0.NFET_GATE_10uA.n19 bgr_9_0.NFET_GATE_10uA.t1 384.967
R1 bgr_9_0.NFET_GATE_10uA.n10 bgr_9_0.NFET_GATE_10uA.t10 369.534
R2 bgr_9_0.NFET_GATE_10uA.n9 bgr_9_0.NFET_GATE_10uA.t22 369.534
R3 bgr_9_0.NFET_GATE_10uA.n7 bgr_9_0.NFET_GATE_10uA.t7 369.534
R4 bgr_9_0.NFET_GATE_10uA.n4 bgr_9_0.NFET_GATE_10uA.t16 369.534
R5 bgr_9_0.NFET_GATE_10uA.n1 bgr_9_0.NFET_GATE_10uA.t12 369.534
R6 bgr_9_0.NFET_GATE_10uA.t1 bgr_9_0.NFET_GATE_10uA.n18 369.534
R7 bgr_9_0.NFET_GATE_10uA bgr_9_0.NFET_GATE_10uA.n20 366.147
R8 bgr_9_0.NFET_GATE_10uA.n12 bgr_9_0.NFET_GATE_10uA.t9 192.8
R9 bgr_9_0.NFET_GATE_10uA.n11 bgr_9_0.NFET_GATE_10uA.t17 192.8
R10 bgr_9_0.NFET_GATE_10uA.n10 bgr_9_0.NFET_GATE_10uA.t23 192.8
R11 bgr_9_0.NFET_GATE_10uA.n9 bgr_9_0.NFET_GATE_10uA.t11 192.8
R12 bgr_9_0.NFET_GATE_10uA.n7 bgr_9_0.NFET_GATE_10uA.t20 192.8
R13 bgr_9_0.NFET_GATE_10uA.n4 bgr_9_0.NFET_GATE_10uA.t21 192.8
R14 bgr_9_0.NFET_GATE_10uA.n5 bgr_9_0.NFET_GATE_10uA.t8 192.8
R15 bgr_9_0.NFET_GATE_10uA.n6 bgr_9_0.NFET_GATE_10uA.t15 192.8
R16 bgr_9_0.NFET_GATE_10uA.n3 bgr_9_0.NFET_GATE_10uA.t19 192.8
R17 bgr_9_0.NFET_GATE_10uA.n2 bgr_9_0.NFET_GATE_10uA.t5 192.8
R18 bgr_9_0.NFET_GATE_10uA.n1 bgr_9_0.NFET_GATE_10uA.t13 192.8
R19 bgr_9_0.NFET_GATE_10uA.n18 bgr_9_0.NFET_GATE_10uA.t18 192.8
R20 bgr_9_0.NFET_GATE_10uA.n17 bgr_9_0.NFET_GATE_10uA.t6 192.8
R21 bgr_9_0.NFET_GATE_10uA.n16 bgr_9_0.NFET_GATE_10uA.t14 192.8
R22 bgr_9_0.NFET_GATE_10uA.n12 bgr_9_0.NFET_GATE_10uA.n11 176.733
R23 bgr_9_0.NFET_GATE_10uA.n11 bgr_9_0.NFET_GATE_10uA.n10 176.733
R24 bgr_9_0.NFET_GATE_10uA.n5 bgr_9_0.NFET_GATE_10uA.n4 176.733
R25 bgr_9_0.NFET_GATE_10uA.n6 bgr_9_0.NFET_GATE_10uA.n5 176.733
R26 bgr_9_0.NFET_GATE_10uA.n3 bgr_9_0.NFET_GATE_10uA.n2 176.733
R27 bgr_9_0.NFET_GATE_10uA.n2 bgr_9_0.NFET_GATE_10uA.n1 176.733
R28 bgr_9_0.NFET_GATE_10uA.n18 bgr_9_0.NFET_GATE_10uA.n17 176.733
R29 bgr_9_0.NFET_GATE_10uA.n17 bgr_9_0.NFET_GATE_10uA.n16 176.733
R30 bgr_9_0.NFET_GATE_10uA.n14 bgr_9_0.NFET_GATE_10uA.n13 169.852
R31 bgr_9_0.NFET_GATE_10uA.n14 bgr_9_0.NFET_GATE_10uA.n8 169.852
R32 bgr_9_0.NFET_GATE_10uA.n15 bgr_9_0.NFET_GATE_10uA.n14 166.133
R33 bgr_9_0.NFET_GATE_10uA.n19 bgr_9_0.NFET_GATE_10uA.n0 132.5
R34 bgr_9_0.NFET_GATE_10uA.n13 bgr_9_0.NFET_GATE_10uA.n12 56.2338
R35 bgr_9_0.NFET_GATE_10uA.n13 bgr_9_0.NFET_GATE_10uA.n9 56.2338
R36 bgr_9_0.NFET_GATE_10uA.n8 bgr_9_0.NFET_GATE_10uA.n7 56.2338
R37 bgr_9_0.NFET_GATE_10uA.n8 bgr_9_0.NFET_GATE_10uA.n6 56.2338
R38 bgr_9_0.NFET_GATE_10uA.n15 bgr_9_0.NFET_GATE_10uA.n3 56.2338
R39 bgr_9_0.NFET_GATE_10uA.n16 bgr_9_0.NFET_GATE_10uA.n15 56.2338
R40 bgr_9_0.NFET_GATE_10uA.n20 bgr_9_0.NFET_GATE_10uA.t3 39.4005
R41 bgr_9_0.NFET_GATE_10uA.n20 bgr_9_0.NFET_GATE_10uA.t4 39.4005
R42 bgr_9_0.NFET_GATE_10uA bgr_9_0.NFET_GATE_10uA.n19 30.6442
R43 bgr_9_0.NFET_GATE_10uA.n0 bgr_9_0.NFET_GATE_10uA.t0 24.0005
R44 bgr_9_0.NFET_GATE_10uA.n0 bgr_9_0.NFET_GATE_10uA.t2 24.0005
R45 two_stage_opamp_dummy_magic_19_0.Vb3.n23 two_stage_opamp_dummy_magic_19_0.Vb3.t12 650.511
R46 two_stage_opamp_dummy_magic_19_0.Vb3.n19 two_stage_opamp_dummy_magic_19_0.Vb3.t23 611.739
R47 two_stage_opamp_dummy_magic_19_0.Vb3.n14 two_stage_opamp_dummy_magic_19_0.Vb3.t15 611.739
R48 two_stage_opamp_dummy_magic_19_0.Vb3.n8 two_stage_opamp_dummy_magic_19_0.Vb3.t11 611.739
R49 two_stage_opamp_dummy_magic_19_0.Vb3.n6 two_stage_opamp_dummy_magic_19_0.Vb3.t28 611.739
R50 two_stage_opamp_dummy_magic_19_0.Vb3.n21 two_stage_opamp_dummy_magic_19_0.Vb3.t10 463.925
R51 two_stage_opamp_dummy_magic_19_0.Vb3.n13 two_stage_opamp_dummy_magic_19_0.Vb3.t16 463.925
R52 two_stage_opamp_dummy_magic_19_0.Vb3.n22 two_stage_opamp_dummy_magic_19_0.Vb3.n21 446.728
R53 two_stage_opamp_dummy_magic_19_0.Vb3.n22 two_stage_opamp_dummy_magic_19_0.Vb3.n13 446.166
R54 two_stage_opamp_dummy_magic_19_0.Vb3.n19 two_stage_opamp_dummy_magic_19_0.Vb3.t18 421.75
R55 two_stage_opamp_dummy_magic_19_0.Vb3.n20 two_stage_opamp_dummy_magic_19_0.Vb3.t14 421.75
R56 two_stage_opamp_dummy_magic_19_0.Vb3.n14 two_stage_opamp_dummy_magic_19_0.Vb3.t19 421.75
R57 two_stage_opamp_dummy_magic_19_0.Vb3.n15 two_stage_opamp_dummy_magic_19_0.Vb3.t17 421.75
R58 two_stage_opamp_dummy_magic_19_0.Vb3.n16 two_stage_opamp_dummy_magic_19_0.Vb3.t21 421.75
R59 two_stage_opamp_dummy_magic_19_0.Vb3.n17 two_stage_opamp_dummy_magic_19_0.Vb3.t26 421.75
R60 two_stage_opamp_dummy_magic_19_0.Vb3.n18 two_stage_opamp_dummy_magic_19_0.Vb3.t8 421.75
R61 two_stage_opamp_dummy_magic_19_0.Vb3.n8 two_stage_opamp_dummy_magic_19_0.Vb3.t9 421.75
R62 two_stage_opamp_dummy_magic_19_0.Vb3.n9 two_stage_opamp_dummy_magic_19_0.Vb3.t27 421.75
R63 two_stage_opamp_dummy_magic_19_0.Vb3.n10 two_stage_opamp_dummy_magic_19_0.Vb3.t22 421.75
R64 two_stage_opamp_dummy_magic_19_0.Vb3.n11 two_stage_opamp_dummy_magic_19_0.Vb3.t24 421.75
R65 two_stage_opamp_dummy_magic_19_0.Vb3.n12 two_stage_opamp_dummy_magic_19_0.Vb3.t20 421.75
R66 two_stage_opamp_dummy_magic_19_0.Vb3.n6 two_stage_opamp_dummy_magic_19_0.Vb3.t25 421.75
R67 two_stage_opamp_dummy_magic_19_0.Vb3.n7 two_stage_opamp_dummy_magic_19_0.Vb3.t13 421.75
R68 two_stage_opamp_dummy_magic_19_0.Vb3.n20 two_stage_opamp_dummy_magic_19_0.Vb3.n19 167.094
R69 two_stage_opamp_dummy_magic_19_0.Vb3.n15 two_stage_opamp_dummy_magic_19_0.Vb3.n14 167.094
R70 two_stage_opamp_dummy_magic_19_0.Vb3.n16 two_stage_opamp_dummy_magic_19_0.Vb3.n15 167.094
R71 two_stage_opamp_dummy_magic_19_0.Vb3.n17 two_stage_opamp_dummy_magic_19_0.Vb3.n16 167.094
R72 two_stage_opamp_dummy_magic_19_0.Vb3.n18 two_stage_opamp_dummy_magic_19_0.Vb3.n17 167.094
R73 two_stage_opamp_dummy_magic_19_0.Vb3.n9 two_stage_opamp_dummy_magic_19_0.Vb3.n8 167.094
R74 two_stage_opamp_dummy_magic_19_0.Vb3.n10 two_stage_opamp_dummy_magic_19_0.Vb3.n9 167.094
R75 two_stage_opamp_dummy_magic_19_0.Vb3.n11 two_stage_opamp_dummy_magic_19_0.Vb3.n10 167.094
R76 two_stage_opamp_dummy_magic_19_0.Vb3.n12 two_stage_opamp_dummy_magic_19_0.Vb3.n11 167.094
R77 two_stage_opamp_dummy_magic_19_0.Vb3.n7 two_stage_opamp_dummy_magic_19_0.Vb3.n6 167.094
R78 two_stage_opamp_dummy_magic_19_0.Vb3.n21 two_stage_opamp_dummy_magic_19_0.Vb3.n20 147.814
R79 two_stage_opamp_dummy_magic_19_0.Vb3.n21 two_stage_opamp_dummy_magic_19_0.Vb3.n18 147.814
R80 two_stage_opamp_dummy_magic_19_0.Vb3.n13 two_stage_opamp_dummy_magic_19_0.Vb3.n12 147.814
R81 two_stage_opamp_dummy_magic_19_0.Vb3.n13 two_stage_opamp_dummy_magic_19_0.Vb3.n7 147.814
R82 two_stage_opamp_dummy_magic_19_0.Vb3.n2 two_stage_opamp_dummy_magic_19_0.Vb3.n1 145.262
R83 two_stage_opamp_dummy_magic_19_0.Vb3.n2 two_stage_opamp_dummy_magic_19_0.Vb3.n0 145.262
R84 two_stage_opamp_dummy_magic_19_0.Vb3.n4 two_stage_opamp_dummy_magic_19_0.Vb3.n3 140.201
R85 two_stage_opamp_dummy_magic_19_0.Vb3.n24 two_stage_opamp_dummy_magic_19_0.Vb3.n5 73.1484
R86 bgr_9_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_19_0.Vb3.n24 48.0943
R87 bgr_9_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_19_0.Vb3.n4 41.063
R88 two_stage_opamp_dummy_magic_19_0.Vb3.n3 two_stage_opamp_dummy_magic_19_0.Vb3.t6 24.0005
R89 two_stage_opamp_dummy_magic_19_0.Vb3.n3 two_stage_opamp_dummy_magic_19_0.Vb3.t4 24.0005
R90 two_stage_opamp_dummy_magic_19_0.Vb3.n1 two_stage_opamp_dummy_magic_19_0.Vb3.t5 24.0005
R91 two_stage_opamp_dummy_magic_19_0.Vb3.n1 two_stage_opamp_dummy_magic_19_0.Vb3.t0 24.0005
R92 two_stage_opamp_dummy_magic_19_0.Vb3.n0 two_stage_opamp_dummy_magic_19_0.Vb3.t3 24.0005
R93 two_stage_opamp_dummy_magic_19_0.Vb3.n0 two_stage_opamp_dummy_magic_19_0.Vb3.t7 24.0005
R94 two_stage_opamp_dummy_magic_19_0.Vb3.n23 two_stage_opamp_dummy_magic_19_0.Vb3.n22 13.7349
R95 two_stage_opamp_dummy_magic_19_0.Vb3.n5 two_stage_opamp_dummy_magic_19_0.Vb3.t2 11.2576
R96 two_stage_opamp_dummy_magic_19_0.Vb3.n5 two_stage_opamp_dummy_magic_19_0.Vb3.t1 11.2576
R97 two_stage_opamp_dummy_magic_19_0.Vb3.n4 two_stage_opamp_dummy_magic_19_0.Vb3.n2 4.5005
R98 two_stage_opamp_dummy_magic_19_0.Vb3.n24 two_stage_opamp_dummy_magic_19_0.Vb3.n23 1.438
R99 GNDA.n2088 GNDA.n52 89432.2
R100 GNDA.n2086 GNDA.n52 87364.4
R101 GNDA.n2160 GNDA.n41 21966.8
R102 GNDA.n2210 GNDA.n7 21966.8
R103 GNDA.n2092 GNDA.n43 14422.9
R104 GNDA.n2211 GNDA.n2210 14422.9
R105 GNDA.n51 GNDA.n50 13528.5
R106 GNDA.n2091 GNDA.n44 13525
R107 GNDA.n49 GNDA.n5 13200
R108 GNDA.n2093 GNDA.n5 12089.3
R109 GNDA.n2212 GNDA.n5 12089.3
R110 GNDA.n2086 GNDA.n2085 11953.3
R111 GNDA.n2085 GNDA.n53 11949.5
R112 GNDA.n50 GNDA.n49 11178.4
R113 GNDA.n118 GNDA.n53 10235.4
R114 GNDA.n50 GNDA.n6 9632.43
R115 GNDA.n47 GNDA.n6 9001.83
R116 GNDA.n2089 GNDA.n2088 8675.66
R117 GNDA.n2087 GNDA.n46 7809.38
R118 GNDA.n2211 GNDA.n6 7750.87
R119 GNDA.n118 GNDA.n46 7720.41
R120 GNDA.n2092 GNDA.n2091 7550.39
R121 GNDA.n2091 GNDA.n2090 6585.23
R122 GNDA.n52 GNDA.n45 5523.81
R123 GNDA.n51 GNDA.n44 4710.92
R124 GNDA.n2087 GNDA.n2086 4106.67
R125 GNDA.n49 GNDA.n44 3989.43
R126 GNDA.n2085 GNDA.n2084 3974.19
R127 GNDA.n120 GNDA.n53 3962.24
R128 GNDA.n47 GNDA.t294 3393.05
R129 GNDA.n2089 GNDA.n46 3166.19
R130 GNDA.n2090 GNDA.n43 2972.3
R131 GNDA.n2090 GNDA.n45 2522.64
R132 GNDA.n2089 GNDA.n51 2313.14
R133 GNDA.n2212 GNDA.n2211 1986.41
R134 GNDA.n2093 GNDA.n2092 1986.41
R135 GNDA.t132 GNDA.n41 1966.49
R136 GNDA.n2088 GNDA.n2087 1863.53
R137 GNDA.n2090 GNDA.n2089 1697.99
R138 GNDA.n2089 GNDA.n48 1647.44
R139 GNDA.n119 GNDA.n48 1397
R140 GNDA.n1913 GNDA.n1912 1336.64
R141 GNDA.t149 GNDA.n120 1225.15
R142 GNDA.n1522 GNDA.n136 1221.08
R143 GNDA.n1806 GNDA.n148 1214.72
R144 GNDA.n1813 GNDA.n1806 1214.72
R145 GNDA.n1814 GNDA.n1813 1214.72
R146 GNDA.n1814 GNDA.n1802 1214.72
R147 GNDA.n1820 GNDA.n1802 1214.72
R148 GNDA.n1822 GNDA.n1798 1214.72
R149 GNDA.n1828 GNDA.n1798 1214.72
R150 GNDA.n1828 GNDA.n1794 1214.72
R151 GNDA.n1834 GNDA.n1794 1214.72
R152 GNDA.n1835 GNDA.n1834 1214.72
R153 GNDA.n1091 GNDA.n1090 1214.72
R154 GNDA.n1090 GNDA.n1089 1214.72
R155 GNDA.n1089 GNDA.n1052 1214.72
R156 GNDA.n1083 GNDA.n1052 1214.72
R157 GNDA.n1083 GNDA.n1082 1214.72
R158 GNDA.n1079 GNDA.n1060 1214.72
R159 GNDA.n1066 GNDA.n1060 1214.72
R160 GNDA.n1072 GNDA.n1066 1214.72
R161 GNDA.n1072 GNDA.n1071 1214.72
R162 GNDA.n1071 GNDA.n1070 1214.72
R163 GNDA.n2058 GNDA.n2057 1185.07
R164 GNDA.n2057 GNDA.n81 1185.07
R165 GNDA.n120 GNDA.n119 937.1
R166 GNDA.n43 GNDA.t145 927.827
R167 GNDA.n119 GNDA.n118 832.433
R168 GNDA.n1820 GNDA.t199 823.313
R169 GNDA.n1082 GNDA.t199 823.313
R170 GNDA.t96 GNDA.n45 744.481
R171 GNDA.n2111 GNDA.t264 739.701
R172 GNDA.n2095 GNDA.t254 739.701
R173 GNDA.n2205 GNDA.t281 739.701
R174 GNDA.n2207 GNDA.t208 739.701
R175 GNDA.t145 GNDA.n41 726.957
R176 GNDA.n1955 GNDA.n1954 669.307
R177 GNDA.n2135 GNDA.t211 659.367
R178 GNDA.n2114 GNDA.t223 659.367
R179 GNDA.n2147 GNDA.t206 659.367
R180 GNDA.n2172 GNDA.t262 659.367
R181 GNDA.n2168 GNDA.t240 659.367
R182 GNDA.n2177 GNDA.t287 659.367
R183 GNDA.t85 GNDA.n117 585
R184 GNDA.n1520 GNDA.n1519 585
R185 GNDA.n1527 GNDA.n1526 585
R186 GNDA.n1528 GNDA.n1527 585
R187 GNDA.n1517 GNDA.n1516 585
R188 GNDA.n1529 GNDA.n1517 585
R189 GNDA.n1532 GNDA.n1531 585
R190 GNDA.n1531 GNDA.n1530 585
R191 GNDA.n1533 GNDA.n1515 585
R192 GNDA.n1518 GNDA.n1515 585
R193 GNDA.n1535 GNDA.n1534 585
R194 GNDA.n1535 GNDA.n89 585
R195 GNDA.n1536 GNDA.n1514 585
R196 GNDA.n1536 GNDA.n88 585
R197 GNDA.n1539 GNDA.n1538 585
R198 GNDA.n1538 GNDA.n1537 585
R199 GNDA.n1540 GNDA.n1512 585
R200 GNDA.n1512 GNDA.n1511 585
R201 GNDA.n1542 GNDA.n1541 585
R202 GNDA.n1543 GNDA.n1542 585
R203 GNDA.n1513 GNDA.n1510 585
R204 GNDA.n1544 GNDA.n1510 585
R205 GNDA.n1546 GNDA.n1508 585
R206 GNDA.n1546 GNDA.n1545 585
R207 GNDA.n1523 GNDA.n1522 585
R208 GNDA.n679 GNDA.n678 585
R209 GNDA.n673 GNDA.n487 585
R210 GNDA.n677 GNDA.n487 585
R211 GNDA.n675 GNDA.n674 585
R212 GNDA.n676 GNDA.n675 585
R213 GNDA.n672 GNDA.n489 585
R214 GNDA.n489 GNDA.n488 585
R215 GNDA.n671 GNDA.n670 585
R216 GNDA.n670 GNDA.n669 585
R217 GNDA.n667 GNDA.n490 585
R218 GNDA.n668 GNDA.n667 585
R219 GNDA.n666 GNDA.n492 585
R220 GNDA.n666 GNDA.n665 585
R221 GNDA.n660 GNDA.n491 585
R222 GNDA.n664 GNDA.n491 585
R223 GNDA.n662 GNDA.n661 585
R224 GNDA.n663 GNDA.n662 585
R225 GNDA.n659 GNDA.n494 585
R226 GNDA.n494 GNDA.n493 585
R227 GNDA.n658 GNDA.n657 585
R228 GNDA.n657 GNDA.n656 585
R229 GNDA.n654 GNDA.n495 585
R230 GNDA.n655 GNDA.n654 585
R231 GNDA.n681 GNDA.n486 585
R232 GNDA.n1889 GNDA.n174 585
R233 GNDA.n1888 GNDA.n1887 585
R234 GNDA.n1892 GNDA.n1891 585
R235 GNDA.n1891 GNDA.n1890 585
R236 GNDA.n1893 GNDA.n172 585
R237 GNDA.n172 GNDA.n171 585
R238 GNDA.n1895 GNDA.n1894 585
R239 GNDA.n1896 GNDA.n1895 585
R240 GNDA.n170 GNDA.n169 585
R241 GNDA.n1897 GNDA.n170 585
R242 GNDA.n1900 GNDA.n1899 585
R243 GNDA.n1899 GNDA.n1898 585
R244 GNDA.n1901 GNDA.n168 585
R245 GNDA.n168 GNDA.n167 585
R246 GNDA.n1903 GNDA.n1902 585
R247 GNDA.n1904 GNDA.n1903 585
R248 GNDA.n166 GNDA.n165 585
R249 GNDA.n1905 GNDA.n166 585
R250 GNDA.n1908 GNDA.n1907 585
R251 GNDA.n1907 GNDA.n1906 585
R252 GNDA.n1909 GNDA.n164 585
R253 GNDA.n164 GNDA.n163 585
R254 GNDA.n1911 GNDA.n1910 585
R255 GNDA.n1912 GNDA.n1911 585
R256 GNDA.n1836 GNDA.n1793 585
R257 GNDA.n1836 GNDA.n1835 585
R258 GNDA.n1832 GNDA.n1792 585
R259 GNDA.n1834 GNDA.n1792 585
R260 GNDA.n1831 GNDA.n1830 585
R261 GNDA.n1830 GNDA.n1794 585
R262 GNDA.n1829 GNDA.n1796 585
R263 GNDA.n1829 GNDA.n1828 585
R264 GNDA.n1825 GNDA.n1797 585
R265 GNDA.n1798 GNDA.n1797 585
R266 GNDA.n1824 GNDA.n1823 585
R267 GNDA.n1823 GNDA.n1822 585
R268 GNDA.n1821 GNDA.n1800 585
R269 GNDA.n1821 GNDA.n1820 585
R270 GNDA.n1817 GNDA.n1801 585
R271 GNDA.n1802 GNDA.n1801 585
R272 GNDA.n1816 GNDA.n1815 585
R273 GNDA.n1815 GNDA.n1814 585
R274 GNDA.n1805 GNDA.n1804 585
R275 GNDA.n1813 GNDA.n1805 585
R276 GNDA.n1810 GNDA.n1809 585
R277 GNDA.n1809 GNDA.n1806 585
R278 GNDA.n1808 GNDA.n1807 585
R279 GNDA.n1808 GNDA.n148 585
R280 GNDA.n1807 GNDA.n150 585
R281 GNDA.n150 GNDA.n148 585
R282 GNDA.n1811 GNDA.n1810 585
R283 GNDA.n1811 GNDA.n1806 585
R284 GNDA.n1812 GNDA.n1804 585
R285 GNDA.n1813 GNDA.n1812 585
R286 GNDA.n1816 GNDA.n1803 585
R287 GNDA.n1814 GNDA.n1803 585
R288 GNDA.n1818 GNDA.n1817 585
R289 GNDA.n1818 GNDA.n1802 585
R290 GNDA.n1819 GNDA.n1800 585
R291 GNDA.n1820 GNDA.n1819 585
R292 GNDA.n1824 GNDA.n1799 585
R293 GNDA.n1822 GNDA.n1799 585
R294 GNDA.n1826 GNDA.n1825 585
R295 GNDA.n1826 GNDA.n1798 585
R296 GNDA.n1827 GNDA.n1796 585
R297 GNDA.n1828 GNDA.n1827 585
R298 GNDA.n1831 GNDA.n1795 585
R299 GNDA.n1795 GNDA.n1794 585
R300 GNDA.n1833 GNDA.n1832 585
R301 GNDA.n1834 GNDA.n1833 585
R302 GNDA.n1793 GNDA.n253 585
R303 GNDA.n1835 GNDA.n253 585
R304 GNDA.n571 GNDA.n570 585
R305 GNDA.n573 GNDA.n561 585
R306 GNDA.n574 GNDA.n560 585
R307 GNDA.n577 GNDA.n559 585
R308 GNDA.n578 GNDA.n558 585
R309 GNDA.n581 GNDA.n557 585
R310 GNDA.n582 GNDA.n556 585
R311 GNDA.n585 GNDA.n555 585
R312 GNDA.n586 GNDA.n554 585
R313 GNDA.n587 GNDA.n553 585
R314 GNDA.n562 GNDA.n545 585
R315 GNDA.n592 GNDA.n509 585
R316 GNDA.n592 GNDA.n591 585
R317 GNDA.n547 GNDA.n545 585
R318 GNDA.n588 GNDA.n587 585
R319 GNDA.n589 GNDA.n588 585
R320 GNDA.n586 GNDA.n552 585
R321 GNDA.n585 GNDA.n584 585
R322 GNDA.n583 GNDA.n582 585
R323 GNDA.n581 GNDA.n580 585
R324 GNDA.n579 GNDA.n578 585
R325 GNDA.n577 GNDA.n576 585
R326 GNDA.n575 GNDA.n574 585
R327 GNDA.n573 GNDA.n572 585
R328 GNDA.n571 GNDA.n372 585
R329 GNDA.n589 GNDA.n372 585
R330 GNDA.n1595 GNDA.n1594 585
R331 GNDA.n1491 GNDA.n1490 585
R332 GNDA.n1493 GNDA.n1492 585
R333 GNDA.n1587 GNDA.n1586 585
R334 GNDA.n1585 GNDA.n1584 585
R335 GNDA.n1583 GNDA.n1497 585
R336 GNDA.n1496 GNDA.n1495 585
R337 GNDA.n1577 GNDA.n1576 585
R338 GNDA.n1575 GNDA.n1574 585
R339 GNDA.n1573 GNDA.n1500 585
R340 GNDA.n1499 GNDA.n379 585
R341 GNDA.n1711 GNDA.n376 585
R342 GNDA.n1568 GNDA.n376 585
R343 GNDA.n1570 GNDA.n1499 585
R344 GNDA.n1573 GNDA.n1572 585
R345 GNDA.n1574 GNDA.n1498 585
R346 GNDA.n1578 GNDA.n1577 585
R347 GNDA.n1580 GNDA.n1495 585
R348 GNDA.n1583 GNDA.n1582 585
R349 GNDA.n1584 GNDA.n1494 585
R350 GNDA.n1588 GNDA.n1587 585
R351 GNDA.n1590 GNDA.n1493 585
R352 GNDA.n1591 GNDA.n1490 585
R353 GNDA.n1594 GNDA.n1593 585
R354 GNDA.n1678 GNDA.n394 585
R355 GNDA.n1676 GNDA.n1675 585
R356 GNDA.n396 GNDA.n395 585
R357 GNDA.n1323 GNDA.n1322 585
R358 GNDA.n1328 GNDA.n1320 585
R359 GNDA.n1329 GNDA.n1318 585
R360 GNDA.n1330 GNDA.n1317 585
R361 GNDA.n1315 GNDA.n1313 585
R362 GNDA.n1335 GNDA.n1312 585
R363 GNDA.n1336 GNDA.n1310 585
R364 GNDA.n1309 GNDA.n1281 585
R365 GNDA.n1341 GNDA.n1279 585
R366 GNDA.n1341 GNDA.n1340 585
R367 GNDA.n1338 GNDA.n1281 585
R368 GNDA.n1337 GNDA.n1336 585
R369 GNDA.n1335 GNDA.n1334 585
R370 GNDA.n1333 GNDA.n1313 585
R371 GNDA.n1331 GNDA.n1330 585
R372 GNDA.n1329 GNDA.n1314 585
R373 GNDA.n1328 GNDA.n1327 585
R374 GNDA.n1325 GNDA.n1323 585
R375 GNDA.n397 GNDA.n396 585
R376 GNDA.n1675 GNDA.n1674 585
R377 GNDA.n1672 GNDA.n394 585
R378 GNDA.n1720 GNDA.n365 585
R379 GNDA.n1721 GNDA.n356 585
R380 GNDA.n1724 GNDA.n355 585
R381 GNDA.n1725 GNDA.n354 585
R382 GNDA.n1728 GNDA.n353 585
R383 GNDA.n1729 GNDA.n352 585
R384 GNDA.n1732 GNDA.n351 585
R385 GNDA.n1734 GNDA.n350 585
R386 GNDA.n1735 GNDA.n349 585
R387 GNDA.n1736 GNDA.n348 585
R388 GNDA.n357 GNDA.n339 585
R389 GNDA.n1742 GNDA.n338 585
R390 GNDA.n1742 GNDA.n1741 585
R391 GNDA.n341 GNDA.n339 585
R392 GNDA.n1737 GNDA.n1736 585
R393 GNDA.n1735 GNDA.n347 585
R394 GNDA.n1734 GNDA.n1733 585
R395 GNDA.n1732 GNDA.n1731 585
R396 GNDA.n1730 GNDA.n1729 585
R397 GNDA.n1728 GNDA.n1727 585
R398 GNDA.n1726 GNDA.n1725 585
R399 GNDA.n1724 GNDA.n1723 585
R400 GNDA.n1722 GNDA.n1721 585
R401 GNDA.n1720 GNDA.n1719 585
R402 GNDA.n1068 GNDA.n335 585
R403 GNDA.n1070 GNDA.n1068 585
R404 GNDA.n1067 GNDA.n1064 585
R405 GNDA.n1071 GNDA.n1067 585
R406 GNDA.n1074 GNDA.n1063 585
R407 GNDA.n1072 GNDA.n1063 585
R408 GNDA.n1075 GNDA.n1062 585
R409 GNDA.n1066 GNDA.n1062 585
R410 GNDA.n1076 GNDA.n1058 585
R411 GNDA.n1060 GNDA.n1058 585
R412 GNDA.n1080 GNDA.n1059 585
R413 GNDA.n1080 GNDA.n1079 585
R414 GNDA.n1081 GNDA.n1056 585
R415 GNDA.n1082 GNDA.n1081 585
R416 GNDA.n1085 GNDA.n1055 585
R417 GNDA.n1083 GNDA.n1055 585
R418 GNDA.n1086 GNDA.n1054 585
R419 GNDA.n1054 GNDA.n1052 585
R420 GNDA.n1087 GNDA.n1051 585
R421 GNDA.n1089 GNDA.n1051 585
R422 GNDA.n1050 GNDA.n1033 585
R423 GNDA.n1090 GNDA.n1050 585
R424 GNDA.n1093 GNDA.n1031 585
R425 GNDA.n1091 GNDA.n1031 585
R426 GNDA.n1093 GNDA.n1092 585
R427 GNDA.n1092 GNDA.n1091 585
R428 GNDA.n1049 GNDA.n1033 585
R429 GNDA.n1090 GNDA.n1049 585
R430 GNDA.n1088 GNDA.n1087 585
R431 GNDA.n1089 GNDA.n1088 585
R432 GNDA.n1086 GNDA.n1053 585
R433 GNDA.n1053 GNDA.n1052 585
R434 GNDA.n1085 GNDA.n1084 585
R435 GNDA.n1084 GNDA.n1083 585
R436 GNDA.n1057 GNDA.n1056 585
R437 GNDA.n1082 GNDA.n1057 585
R438 GNDA.n1078 GNDA.n1059 585
R439 GNDA.n1079 GNDA.n1078 585
R440 GNDA.n1077 GNDA.n1076 585
R441 GNDA.n1077 GNDA.n1060 585
R442 GNDA.n1075 GNDA.n1061 585
R443 GNDA.n1066 GNDA.n1061 585
R444 GNDA.n1074 GNDA.n1073 585
R445 GNDA.n1073 GNDA.n1072 585
R446 GNDA.n1065 GNDA.n1064 585
R447 GNDA.n1071 GNDA.n1065 585
R448 GNDA.n1069 GNDA.n335 585
R449 GNDA.n1070 GNDA.n1069 585
R450 GNDA.n1096 GNDA.n1095 585
R451 GNDA.n1097 GNDA.n1096 585
R452 GNDA.n1029 GNDA.n1028 585
R453 GNDA.n1098 GNDA.n1029 585
R454 GNDA.n1101 GNDA.n1100 585
R455 GNDA.n1100 GNDA.n1099 585
R456 GNDA.n1102 GNDA.n1027 585
R457 GNDA.n1027 GNDA.n1026 585
R458 GNDA.n1104 GNDA.n1103 585
R459 GNDA.n1105 GNDA.n1104 585
R460 GNDA.n1025 GNDA.n1024 585
R461 GNDA.n1106 GNDA.n1025 585
R462 GNDA.n1109 GNDA.n1108 585
R463 GNDA.n1108 GNDA.n1107 585
R464 GNDA.n1110 GNDA.n1023 585
R465 GNDA.n1023 GNDA.n1022 585
R466 GNDA.n1112 GNDA.n1111 585
R467 GNDA.n1113 GNDA.n1112 585
R468 GNDA.n1020 GNDA.n1019 585
R469 GNDA.n1114 GNDA.n1020 585
R470 GNDA.n1117 GNDA.n1116 585
R471 GNDA.n1116 GNDA.n1115 585
R472 GNDA.n1118 GNDA.n1018 585
R473 GNDA.n1021 GNDA.n1018 585
R474 GNDA.n147 GNDA.n146 585
R475 GNDA.n1938 GNDA.n147 585
R476 GNDA.n1941 GNDA.n1940 585
R477 GNDA.n1940 GNDA.n1939 585
R478 GNDA.n1942 GNDA.n145 585
R479 GNDA.n145 GNDA.n144 585
R480 GNDA.n1944 GNDA.n1943 585
R481 GNDA.n1945 GNDA.n1944 585
R482 GNDA.n143 GNDA.n141 585
R483 GNDA.n1946 GNDA.n143 585
R484 GNDA.n1949 GNDA.n1948 585
R485 GNDA.n1948 GNDA.n1947 585
R486 GNDA.n142 GNDA.n140 585
R487 GNDA.n1038 GNDA.n142 585
R488 GNDA.n1041 GNDA.n1040 585
R489 GNDA.n1040 GNDA.n1039 585
R490 GNDA.n1042 GNDA.n1036 585
R491 GNDA.n1036 GNDA.n1035 585
R492 GNDA.n1044 GNDA.n1043 585
R493 GNDA.n1045 GNDA.n1044 585
R494 GNDA.n1037 GNDA.n1034 585
R495 GNDA.n1046 GNDA.n1034 585
R496 GNDA.n1048 GNDA.n1032 585
R497 GNDA.n1048 GNDA.n1047 585
R498 GNDA.n162 GNDA.n161 585
R499 GNDA.n1913 GNDA.n162 585
R500 GNDA.n1916 GNDA.n1915 585
R501 GNDA.n1915 GNDA.n1914 585
R502 GNDA.n1917 GNDA.n160 585
R503 GNDA.n160 GNDA.n159 585
R504 GNDA.n1919 GNDA.n1918 585
R505 GNDA.n1920 GNDA.n1919 585
R506 GNDA.n158 GNDA.n157 585
R507 GNDA.n1921 GNDA.n158 585
R508 GNDA.n1924 GNDA.n1923 585
R509 GNDA.n1923 GNDA.n1922 585
R510 GNDA.n1925 GNDA.n156 585
R511 GNDA.n156 GNDA.n155 585
R512 GNDA.n1927 GNDA.n1926 585
R513 GNDA.n1928 GNDA.n1927 585
R514 GNDA.n154 GNDA.n153 585
R515 GNDA.n1929 GNDA.n154 585
R516 GNDA.n1932 GNDA.n1931 585
R517 GNDA.n1931 GNDA.n1930 585
R518 GNDA.n1933 GNDA.n151 585
R519 GNDA.n151 GNDA.n149 585
R520 GNDA.n1935 GNDA.n1934 585
R521 GNDA.n1936 GNDA.n1935 585
R522 GNDA.n1953 GNDA.n139 585
R523 GNDA.n1952 GNDA.n1951 585
R524 GNDA.n1952 GNDA.t199 585
R525 GNDA.n645 GNDA.n336 585
R526 GNDA.n644 GNDA.n643 585
R527 GNDA.n642 GNDA.n602 585
R528 GNDA.n641 GNDA.n640 585
R529 GNDA.n639 GNDA.n638 585
R530 GNDA.n637 GNDA.n636 585
R531 GNDA.n635 GNDA.n634 585
R532 GNDA.n633 GNDA.n632 585
R533 GNDA.n631 GNDA.n630 585
R534 GNDA.n629 GNDA.n628 585
R535 GNDA.n627 GNDA.n626 585
R536 GNDA.n625 GNDA.n624 585
R537 GNDA.n595 GNDA.n594 585
R538 GNDA.n528 GNDA.n508 585
R539 GNDA.n527 GNDA.n526 585
R540 GNDA.n525 GNDA.n524 585
R541 GNDA.n523 GNDA.n522 585
R542 GNDA.n521 GNDA.n520 585
R543 GNDA.n519 GNDA.n518 585
R544 GNDA.n517 GNDA.n516 585
R545 GNDA.n515 GNDA.n514 585
R546 GNDA.n513 GNDA.n512 585
R547 GNDA.n511 GNDA.n510 585
R548 GNDA.n340 GNDA.n337 585
R549 GNDA.n653 GNDA.n652 585
R550 GNDA.n651 GNDA.n650 585
R551 GNDA.n649 GNDA.n497 585
R552 GNDA.n529 GNDA.n498 585
R553 GNDA.n531 GNDA.n530 585
R554 GNDA.n533 GNDA.n532 585
R555 GNDA.n535 GNDA.n534 585
R556 GNDA.n537 GNDA.n536 585
R557 GNDA.n539 GNDA.n538 585
R558 GNDA.n541 GNDA.n540 585
R559 GNDA.n543 GNDA.n542 585
R560 GNDA.n546 GNDA.n544 585
R561 GNDA.n1744 GNDA.n257 585
R562 GNDA.n1838 GNDA.n257 585
R563 GNDA.n1239 GNDA.n1119 585
R564 GNDA.n1237 GNDA.n1236 585
R565 GNDA.n1122 GNDA.n1120 585
R566 GNDA.n1231 GNDA.n1230 585
R567 GNDA.n1228 GNDA.n1227 585
R568 GNDA.n1150 GNDA.n1127 585
R569 GNDA.n1153 GNDA.n1152 585
R570 GNDA.n1156 GNDA.n1148 585
R571 GNDA.n1162 GNDA.n1161 585
R572 GNDA.n1164 GNDA.n1147 585
R573 GNDA.n1168 GNDA.n1167 585
R574 GNDA.n1165 GNDA.n334 585
R575 GNDA.n1837 GNDA.n254 585
R576 GNDA.n1838 GNDA.n1837 585
R577 GNDA.n1744 GNDA.n256 585
R578 GNDA.n1838 GNDA.n256 585
R579 GNDA.n1748 GNDA.n1747 585
R580 GNDA.n1749 GNDA.n271 585
R581 GNDA.n1759 GNDA.n1758 585
R582 GNDA.n1761 GNDA.n270 585
R583 GNDA.n1764 GNDA.n1763 585
R584 GNDA.n1765 GNDA.n266 585
R585 GNDA.n1774 GNDA.n1773 585
R586 GNDA.n1776 GNDA.n265 585
R587 GNDA.n1779 GNDA.n1778 585
R588 GNDA.n1780 GNDA.n259 585
R589 GNDA.n1789 GNDA.n1788 585
R590 GNDA.n1791 GNDA.n258 585
R591 GNDA.n1839 GNDA.n254 585
R592 GNDA.n1839 GNDA.n1838 585
R593 GNDA.n1842 GNDA.n1841 585
R594 GNDA.n1843 GNDA.n189 585
R595 GNDA.n1853 GNDA.n1852 585
R596 GNDA.n1855 GNDA.n188 585
R597 GNDA.n1858 GNDA.n1857 585
R598 GNDA.n1859 GNDA.n184 585
R599 GNDA.n1868 GNDA.n1867 585
R600 GNDA.n1870 GNDA.n183 585
R601 GNDA.n1873 GNDA.n1872 585
R602 GNDA.n1874 GNDA.n177 585
R603 GNDA.n1883 GNDA.n1882 585
R604 GNDA.n1885 GNDA.n175 585
R605 GNDA.n1344 GNDA.n1343 585
R606 GNDA.n1346 GNDA.n1277 585
R607 GNDA.n1348 GNDA.n1347 585
R608 GNDA.n1349 GNDA.n1276 585
R609 GNDA.n1351 GNDA.n1350 585
R610 GNDA.n1353 GNDA.n1274 585
R611 GNDA.n1355 GNDA.n1354 585
R612 GNDA.n1356 GNDA.n1273 585
R613 GNDA.n1358 GNDA.n1357 585
R614 GNDA.n1360 GNDA.n1271 585
R615 GNDA.n1362 GNDA.n1361 585
R616 GNDA.n1363 GNDA.n1270 585
R617 GNDA.n1713 GNDA.n1712 585
R618 GNDA.n1288 GNDA.n377 585
R619 GNDA.n1290 GNDA.n1289 585
R620 GNDA.n1292 GNDA.n1286 585
R621 GNDA.n1294 GNDA.n1293 585
R622 GNDA.n1295 GNDA.n1285 585
R623 GNDA.n1297 GNDA.n1296 585
R624 GNDA.n1299 GNDA.n1283 585
R625 GNDA.n1301 GNDA.n1300 585
R626 GNDA.n1302 GNDA.n1282 585
R627 GNDA.n1304 GNDA.n1303 585
R628 GNDA.n1306 GNDA.n1280 585
R629 GNDA.n1548 GNDA.n1547 585
R630 GNDA.n1549 GNDA.n1507 585
R631 GNDA.n1551 GNDA.n1550 585
R632 GNDA.n1553 GNDA.n1505 585
R633 GNDA.n1555 GNDA.n1554 585
R634 GNDA.n1556 GNDA.n1504 585
R635 GNDA.n1558 GNDA.n1557 585
R636 GNDA.n1560 GNDA.n1502 585
R637 GNDA.n1562 GNDA.n1561 585
R638 GNDA.n1563 GNDA.n1501 585
R639 GNDA.n1565 GNDA.n1564 585
R640 GNDA.n1567 GNDA.n375 585
R641 GNDA.n370 GNDA.n368 585
R642 GNDA.n1717 GNDA.n370 585
R643 GNDA.n1011 GNDA.n449 585
R644 GNDA.n1009 GNDA.n1008 585
R645 GNDA.n898 GNDA.n453 585
R646 GNDA.n1004 GNDA.n1003 585
R647 GNDA.n900 GNDA.n897 585
R648 GNDA.n926 GNDA.n925 585
R649 GNDA.n928 GNDA.n927 585
R650 GNDA.n931 GNDA.n930 585
R651 GNDA.n929 GNDA.n919 585
R652 GNDA.n940 GNDA.n939 585
R653 GNDA.n942 GNDA.n941 585
R654 GNDA.n944 GNDA.n943 585
R655 GNDA.n1715 GNDA.n371 585
R656 GNDA.n1717 GNDA.n371 585
R657 GNDA.n1718 GNDA.n368 585
R658 GNDA.n1718 GNDA.n1717 585
R659 GNDA.n778 GNDA.n367 585
R660 GNDA.n891 GNDA.n890 585
R661 GNDA.n780 GNDA.n777 585
R662 GNDA.n885 GNDA.n884 585
R663 GNDA.n883 GNDA.n882 585
R664 GNDA.n808 GNDA.n784 585
R665 GNDA.n810 GNDA.n809 585
R666 GNDA.n815 GNDA.n814 585
R667 GNDA.n813 GNDA.n806 585
R668 GNDA.n821 GNDA.n820 585
R669 GNDA.n823 GNDA.n822 585
R670 GNDA.n804 GNDA.n803 585
R671 GNDA.n1716 GNDA.n1715 585
R672 GNDA.n1717 GNDA.n1716 585
R673 GNDA.n460 GNDA.n373 585
R674 GNDA.n770 GNDA.n769 585
R675 GNDA.n462 GNDA.n459 585
R676 GNDA.n764 GNDA.n763 585
R677 GNDA.n762 GNDA.n761 585
R678 GNDA.n687 GNDA.n466 585
R679 GNDA.n689 GNDA.n688 585
R680 GNDA.n694 GNDA.n693 585
R681 GNDA.n692 GNDA.n685 585
R682 GNDA.n700 GNDA.n699 585
R683 GNDA.n702 GNDA.n701 585
R684 GNDA.n683 GNDA.n682 585
R685 GNDA.n1365 GNDA.n1364 585
R686 GNDA.n1367 GNDA.n1269 585
R687 GNDA.n1370 GNDA.n1369 585
R688 GNDA.n1371 GNDA.n1268 585
R689 GNDA.n1373 GNDA.n1372 585
R690 GNDA.n1375 GNDA.n1267 585
R691 GNDA.n1378 GNDA.n1377 585
R692 GNDA.n1379 GNDA.n1266 585
R693 GNDA.n1381 GNDA.n1380 585
R694 GNDA.n1383 GNDA.n1265 585
R695 GNDA.n1384 GNDA.n437 585
R696 GNDA.n1264 GNDA.n436 585
R697 GNDA.n623 GNDA.n622 585
R698 GNDA.n621 GNDA.n620 585
R699 GNDA.n619 GNDA.n618 585
R700 GNDA.n617 GNDA.n616 585
R701 GNDA.n615 GNDA.n614 585
R702 GNDA.n613 GNDA.n612 585
R703 GNDA.n611 GNDA.n610 585
R704 GNDA.n609 GNDA.n608 585
R705 GNDA.n607 GNDA.n606 585
R706 GNDA.n605 GNDA.n604 585
R707 GNDA.n603 GNDA.n450 585
R708 GNDA.n1264 GNDA.n1014 585
R709 GNDA.n1262 GNDA.n1261 585
R710 GNDA.n1260 GNDA.n1017 585
R711 GNDA.n1259 GNDA.n1016 585
R712 GNDA.n1264 GNDA.n1016 585
R713 GNDA.n1258 GNDA.n1257 585
R714 GNDA.n1256 GNDA.n1255 585
R715 GNDA.n1254 GNDA.n1253 585
R716 GNDA.n1252 GNDA.n1251 585
R717 GNDA.n1250 GNDA.n1249 585
R718 GNDA.n1248 GNDA.n1247 585
R719 GNDA.n1246 GNDA.n1245 585
R720 GNDA.n1244 GNDA.n1243 585
R721 GNDA.n1242 GNDA.n1241 585
R722 GNDA.n1241 GNDA.n1240 585
R723 GNDA.n435 GNDA.n434 585
R724 GNDA.n1682 GNDA.n1681 585
R725 GNDA.n1708 GNDA.n1707 585
R726 GNDA.n1694 GNDA.n386 585
R727 GNDA.n1691 GNDA.n1690 585
R728 GNDA.n1964 GNDA.n1963 585
R729 GNDA.n1679 GNDA.n393 585
R730 GNDA.n1680 GNDA.n1679 585
R731 GNDA.n1441 GNDA.n1440 585
R732 GNDA.n1442 GNDA.n1441 585
R733 GNDA.n427 GNDA.n425 585
R734 GNDA.n1443 GNDA.n427 585
R735 GNDA.n1468 GNDA.n1467 585
R736 GNDA.n1467 GNDA.n1466 585
R737 GNDA.n1446 GNDA.n428 585
R738 GNDA.n1465 GNDA.n428 585
R739 GNDA.n1463 GNDA.n1462 585
R740 GNDA.n1464 GNDA.n1463 585
R741 GNDA.n1458 GNDA.n1445 585
R742 GNDA.n1445 GNDA.n1444 585
R743 GNDA.n1452 GNDA.n1451 585
R744 GNDA.n1451 GNDA.n1450 585
R745 GNDA.n1453 GNDA.n401 585
R746 GNDA.n1449 GNDA.n401 585
R747 GNDA.n1476 GNDA.n1475 585
R748 GNDA.n1477 GNDA.n1476 585
R749 GNDA.n403 GNDA.n400 585
R750 GNDA.n1478 GNDA.n400 585
R751 GNDA.n1482 GNDA.n1481 585
R752 GNDA.n1481 GNDA.n1480 585
R753 GNDA.n1484 GNDA.n392 585
R754 GNDA.n1479 GNDA.n392 585
R755 GNDA.n1596 GNDA.n1489 585
R756 GNDA.n1598 GNDA.n1596 585
R757 GNDA.n1671 GNDA.n393 585
R758 GNDA.n1671 GNDA.n389 585
R759 GNDA.n1670 GNDA.n1668 585
R760 GNDA.n1670 GNDA.n1669 585
R761 GNDA.n79 GNDA.n77 585
R762 GNDA.n2059 GNDA.n79 585
R763 GNDA.n2074 GNDA.n2073 585
R764 GNDA.n2073 GNDA.n2072 585
R765 GNDA.n2061 GNDA.n80 585
R766 GNDA.n2071 GNDA.n80 585
R767 GNDA.n2069 GNDA.n2068 585
R768 GNDA.n2070 GNDA.n2069 585
R769 GNDA.n2064 GNDA.n54 585
R770 GNDA.n2060 GNDA.n54 585
R771 GNDA.n2082 GNDA.n2081 585
R772 GNDA.n2083 GNDA.n2082 585
R773 GNDA.n56 GNDA.n55 585
R774 GNDA.n1601 GNDA.n55 585
R775 GNDA.n1606 GNDA.n1605 585
R776 GNDA.n1607 GNDA.n1606 585
R777 GNDA.n1488 GNDA.n1487 585
R778 GNDA.n1608 GNDA.n1488 585
R779 GNDA.n1611 GNDA.n1610 585
R780 GNDA.n1610 GNDA.n1609 585
R781 GNDA.n1600 GNDA.n1597 585
R782 GNDA.n1600 GNDA.n1599 585
R783 GNDA.n1489 GNDA.n122 585
R784 GNDA.n1689 GNDA.n122 585
R785 GNDA.n2026 GNDA.n2025 585
R786 GNDA.n2027 GNDA.n2026 585
R787 GNDA.n115 GNDA.n113 585
R788 GNDA.n2028 GNDA.n115 585
R789 GNDA.n2043 GNDA.n2042 585
R790 GNDA.n2042 GNDA.n2041 585
R791 GNDA.n2030 GNDA.n116 585
R792 GNDA.n2040 GNDA.n116 585
R793 GNDA.n2038 GNDA.n2037 585
R794 GNDA.n2039 GNDA.n2038 585
R795 GNDA.n2033 GNDA.n90 585
R796 GNDA.n2029 GNDA.n90 585
R797 GNDA.n2051 GNDA.n2050 585
R798 GNDA.n2052 GNDA.n2051 585
R799 GNDA.n92 GNDA.n91 585
R800 GNDA.n128 GNDA.n91 585
R801 GNDA.n133 GNDA.n132 585
R802 GNDA.n134 GNDA.n133 585
R803 GNDA.n126 GNDA.n125 585
R804 GNDA.n135 GNDA.n126 585
R805 GNDA.n1968 GNDA.n1967 585
R806 GNDA.n1967 GNDA.n1966 585
R807 GNDA.n1521 GNDA.n127 585
R808 GNDA.n1965 GNDA.n127 585
R809 GNDA.n2100 GNDA.t193 514.768
R810 GNDA.n2194 GNDA.t284 514.768
R811 GNDA.n2200 GNDA.t203 514.768
R812 GNDA.n2106 GNDA.t257 514.768
R813 GNDA.n1835 GNDA.t199 512.884
R814 GNDA.n1070 GNDA.t199 512.884
R815 GNDA.n2140 GNDA.t217 508.743
R816 GNDA.n2150 GNDA.t227 508.743
R817 GNDA.n2188 GNDA.t269 508.743
R818 GNDA.n2190 GNDA.t279 508.743
R819 GNDA.n2162 GNDA.t220 508.743
R820 GNDA.n2165 GNDA.t236 508.743
R821 GNDA.n2182 GNDA.t275 508.743
R822 GNDA.n2180 GNDA.t200 508.743
R823 GNDA.n1 GNDA.t260 508.743
R824 GNDA.n2220 GNDA.t267 508.743
R825 GNDA.n28 GNDA.t238 498.7
R826 GNDA.n2176 GNDA.t277 498.7
R827 GNDA.n2109 GNDA.n42 445.375
R828 GNDA.n2203 GNDA.n2192 445.375
R829 GNDA.n2170 GNDA.n27 431.902
R830 GNDA.n2184 GNDA.n22 431.902
R831 GNDA.n433 GNDA.t244 409.067
R832 GNDA.n1683 GNDA.t251 409.067
R833 GNDA.n1706 GNDA.t272 409.067
R834 GNDA.n1695 GNDA.t230 409.067
R835 GNDA.n1692 GNDA.t247 409.067
R836 GNDA.n1962 GNDA.t233 409.067
R837 GNDA.n1822 GNDA.t199 391.411
R838 GNDA.n1079 GNDA.t199 391.411
R839 GNDA.n2160 GNDA.t218 364.418
R840 GNDA.t228 GNDA.n27 364.418
R841 GNDA.t143 GNDA.n2170 364.418
R842 GNDA.t15 GNDA.n22 364.418
R843 GNDA.t270 GNDA.n2184 364.418
R844 GNDA.t201 GNDA.n7 364.418
R845 GNDA.n385 GNDA.t199 172.876
R846 GNDA.n1709 GNDA.t199 172.876
R847 GNDA.n388 GNDA.t199 172.615
R848 GNDA.t199 GNDA.n87 172.615
R849 GNDA.n48 GNDA.n47 309.122
R850 GNDA.n2171 GNDA.n26 299.443
R851 GNDA.t7 GNDA.t228 296.933
R852 GNDA.t304 GNDA.t49 296.933
R853 GNDA.n2139 GNDA.n42 296.158
R854 GNDA.n2152 GNDA.n2151 296.158
R855 GNDA.n2187 GNDA.n2186 296.158
R856 GNDA.n2192 GNDA.n2191 296.158
R857 GNDA.n2161 GNDA.n2160 296.158
R858 GNDA.n2164 GNDA.n27 296.158
R859 GNDA.n2145 GNDA.n2144 296.158
R860 GNDA.n2175 GNDA.n2174 296.158
R861 GNDA.n2184 GNDA.n2183 296.158
R862 GNDA.n2179 GNDA.n7 296.158
R863 GNDA.n2219 GNDA.n2218 296.158
R864 GNDA.t67 GNDA.t199 294.625
R865 GNDA.n1264 GNDA.n442 264.301
R866 GNDA.n1525 GNDA.n1524 264.301
R867 GNDA.n680 GNDA.n485 264.301
R868 GNDA.n1886 GNDA.n173 264.301
R869 GNDA.n1387 GNDA.n1386 264.301
R870 GNDA.n1013 GNDA.n1012 264.301
R871 GNDA.n1096 GNDA.n1031 259.416
R872 GNDA.n645 GNDA.n338 259.416
R873 GNDA.n1344 GNDA.n1279 259.416
R874 GNDA.n1712 GNDA.n1711 259.416
R875 GNDA.n595 GNDA.n509 259.416
R876 GNDA.n1808 GNDA.n147 259.416
R877 GNDA.n654 GNDA.n653 259.416
R878 GNDA.n1547 GNDA.n1546 259.416
R879 GNDA.n1911 GNDA.n162 259.416
R880 GNDA.n1205 GNDA.n1144 258.334
R881 GNDA.n981 GNDA.n979 258.334
R882 GNDA.n1422 GNDA.n1421 258.334
R883 GNDA.n1650 GNDA.n1649 258.334
R884 GNDA.n860 GNDA.n801 258.334
R885 GNDA.n319 GNDA.n277 258.334
R886 GNDA.n739 GNDA.n483 258.334
R887 GNDA.n2007 GNDA.n2006 258.334
R888 GNDA.n237 GNDA.n195 258.334
R889 GNDA.n569 GNDA.n568 254.34
R890 GNDA.n568 GNDA.n567 254.34
R891 GNDA.n568 GNDA.n566 254.34
R892 GNDA.n568 GNDA.n565 254.34
R893 GNDA.n568 GNDA.n564 254.34
R894 GNDA.n568 GNDA.n563 254.34
R895 GNDA.n590 GNDA.n589 254.34
R896 GNDA.n589 GNDA.n548 254.34
R897 GNDA.n589 GNDA.n549 254.34
R898 GNDA.n589 GNDA.n550 254.34
R899 GNDA.n589 GNDA.n551 254.34
R900 GNDA.n1709 GNDA.n384 254.34
R901 GNDA.n1709 GNDA.n383 254.34
R902 GNDA.n1709 GNDA.n382 254.34
R903 GNDA.n1709 GNDA.n381 254.34
R904 GNDA.n1709 GNDA.n380 254.34
R905 GNDA.n1710 GNDA.n1709 254.34
R906 GNDA.n1569 GNDA.n87 254.34
R907 GNDA.n1571 GNDA.n87 254.34
R908 GNDA.n1579 GNDA.n87 254.34
R909 GNDA.n1581 GNDA.n87 254.34
R910 GNDA.n1589 GNDA.n87 254.34
R911 GNDA.n1592 GNDA.n87 254.34
R912 GNDA.n1677 GNDA.n385 254.34
R913 GNDA.n1321 GNDA.n385 254.34
R914 GNDA.n1319 GNDA.n385 254.34
R915 GNDA.n1316 GNDA.n385 254.34
R916 GNDA.n1311 GNDA.n385 254.34
R917 GNDA.n1308 GNDA.n385 254.34
R918 GNDA.n1339 GNDA.n388 254.34
R919 GNDA.n1307 GNDA.n388 254.34
R920 GNDA.n1332 GNDA.n388 254.34
R921 GNDA.n1326 GNDA.n388 254.34
R922 GNDA.n1324 GNDA.n388 254.34
R923 GNDA.n1673 GNDA.n388 254.34
R924 GNDA.n364 GNDA.n363 254.34
R925 GNDA.n363 GNDA.n362 254.34
R926 GNDA.n363 GNDA.n361 254.34
R927 GNDA.n363 GNDA.n360 254.34
R928 GNDA.n363 GNDA.n359 254.34
R929 GNDA.n363 GNDA.n358 254.34
R930 GNDA.n1740 GNDA.n1739 254.34
R931 GNDA.n1739 GNDA.n1738 254.34
R932 GNDA.n1739 GNDA.n346 254.34
R933 GNDA.n1739 GNDA.n345 254.34
R934 GNDA.n1739 GNDA.n344 254.34
R935 GNDA.n1739 GNDA.n343 254.34
R936 GNDA.n647 GNDA.n646 254.34
R937 GNDA.n647 GNDA.n601 254.34
R938 GNDA.n647 GNDA.n600 254.34
R939 GNDA.n647 GNDA.n599 254.34
R940 GNDA.n647 GNDA.n598 254.34
R941 GNDA.n647 GNDA.n597 254.34
R942 GNDA.n647 GNDA.n596 254.34
R943 GNDA.n647 GNDA.n507 254.34
R944 GNDA.n647 GNDA.n506 254.34
R945 GNDA.n647 GNDA.n505 254.34
R946 GNDA.n647 GNDA.n504 254.34
R947 GNDA.n647 GNDA.n503 254.34
R948 GNDA.n647 GNDA.n496 254.34
R949 GNDA.n648 GNDA.n647 254.34
R950 GNDA.n647 GNDA.n502 254.34
R951 GNDA.n647 GNDA.n501 254.34
R952 GNDA.n647 GNDA.n500 254.34
R953 GNDA.n647 GNDA.n499 254.34
R954 GNDA.n1238 GNDA.n176 254.34
R955 GNDA.n1229 GNDA.n176 254.34
R956 GNDA.n1126 GNDA.n176 254.34
R957 GNDA.n1151 GNDA.n176 254.34
R958 GNDA.n1163 GNDA.n176 254.34
R959 GNDA.n1166 GNDA.n176 254.34
R960 GNDA.n1746 GNDA.n176 254.34
R961 GNDA.n1760 GNDA.n176 254.34
R962 GNDA.n1762 GNDA.n176 254.34
R963 GNDA.n1775 GNDA.n176 254.34
R964 GNDA.n1777 GNDA.n176 254.34
R965 GNDA.n1790 GNDA.n176 254.34
R966 GNDA.n1840 GNDA.n176 254.34
R967 GNDA.n1854 GNDA.n176 254.34
R968 GNDA.n1856 GNDA.n176 254.34
R969 GNDA.n1869 GNDA.n176 254.34
R970 GNDA.n1871 GNDA.n176 254.34
R971 GNDA.n1884 GNDA.n176 254.34
R972 GNDA.n1345 GNDA.n387 254.34
R973 GNDA.n1278 GNDA.n387 254.34
R974 GNDA.n1352 GNDA.n387 254.34
R975 GNDA.n1275 GNDA.n387 254.34
R976 GNDA.n1359 GNDA.n387 254.34
R977 GNDA.n1272 GNDA.n387 254.34
R978 GNDA.n387 GNDA.n378 254.34
R979 GNDA.n1291 GNDA.n387 254.34
R980 GNDA.n1287 GNDA.n387 254.34
R981 GNDA.n1298 GNDA.n387 254.34
R982 GNDA.n1284 GNDA.n387 254.34
R983 GNDA.n1305 GNDA.n387 254.34
R984 GNDA.n1509 GNDA.n387 254.34
R985 GNDA.n1552 GNDA.n387 254.34
R986 GNDA.n1506 GNDA.n387 254.34
R987 GNDA.n1559 GNDA.n387 254.34
R988 GNDA.n1503 GNDA.n387 254.34
R989 GNDA.n1566 GNDA.n387 254.34
R990 GNDA.n1007 GNDA.n1006 254.34
R991 GNDA.n1006 GNDA.n1005 254.34
R992 GNDA.n1006 GNDA.n896 254.34
R993 GNDA.n1006 GNDA.n895 254.34
R994 GNDA.n1006 GNDA.n894 254.34
R995 GNDA.n1006 GNDA.n893 254.34
R996 GNDA.n1006 GNDA.n892 254.34
R997 GNDA.n1006 GNDA.n776 254.34
R998 GNDA.n1006 GNDA.n775 254.34
R999 GNDA.n1006 GNDA.n774 254.34
R1000 GNDA.n1006 GNDA.n773 254.34
R1001 GNDA.n1006 GNDA.n772 254.34
R1002 GNDA.n1006 GNDA.n771 254.34
R1003 GNDA.n1006 GNDA.n458 254.34
R1004 GNDA.n1006 GNDA.n457 254.34
R1005 GNDA.n1006 GNDA.n456 254.34
R1006 GNDA.n1006 GNDA.n455 254.34
R1007 GNDA.n1006 GNDA.n454 254.34
R1008 GNDA.n1366 GNDA.n1264 254.34
R1009 GNDA.n1368 GNDA.n1264 254.34
R1010 GNDA.n1374 GNDA.n1264 254.34
R1011 GNDA.n1376 GNDA.n1264 254.34
R1012 GNDA.n1382 GNDA.n1264 254.34
R1013 GNDA.n1385 GNDA.n1264 254.34
R1014 GNDA.n1264 GNDA.n443 254.34
R1015 GNDA.n1264 GNDA.n444 254.34
R1016 GNDA.n1264 GNDA.n445 254.34
R1017 GNDA.n1264 GNDA.n446 254.34
R1018 GNDA.n1264 GNDA.n447 254.34
R1019 GNDA.n1264 GNDA.n448 254.34
R1020 GNDA.n1264 GNDA.n1263 254.34
R1021 GNDA.n1264 GNDA.n438 254.34
R1022 GNDA.n1264 GNDA.n439 254.34
R1023 GNDA.n1264 GNDA.n440 254.34
R1024 GNDA.n1264 GNDA.n441 254.34
R1025 GNDA.n1954 GNDA.t199 250.349
R1026 GNDA.n1262 GNDA.n1018 249.663
R1027 GNDA.n624 GNDA.n623 249.663
R1028 GNDA.n1365 GNDA.n1270 249.663
R1029 GNDA.n1340 GNDA.n1306 249.663
R1030 GNDA.n1741 GNDA.n340 249.663
R1031 GNDA.n1092 GNDA.n1048 249.663
R1032 GNDA.n591 GNDA.n546 249.663
R1033 GNDA.n1568 GNDA.n1567 249.663
R1034 GNDA.n1935 GNDA.n150 249.663
R1035 GNDA.n2158 GNDA.n2094 201.192
R1036 GNDA.n2214 GNDA.n4 201.192
R1037 GNDA.n2146 GNDA.n2145 197.133
R1038 GNDA.n2174 GNDA.n2173 197.133
R1039 GNDA.n2170 GNDA.n2169 197.133
R1040 GNDA.n25 GNDA.n22 197.133
R1041 GNDA.n1953 GNDA.n1952 197
R1042 GNDA.n1165 GNDA.n257 197
R1043 GNDA.n943 GNDA.n370 197
R1044 GNDA.n1679 GNDA.n392 197
R1045 GNDA.n1600 GNDA.n1596 197
R1046 GNDA.n803 GNDA.n371 197
R1047 GNDA.n1837 GNDA.n1791 197
R1048 GNDA.n682 GNDA.n681 197
R1049 GNDA.n1523 GNDA.n127 197
R1050 GNDA.n1887 GNDA.n1885 197
R1051 GNDA.n2054 GNDA.n2053 195
R1052 GNDA.n1448 GNDA.n83 195
R1053 GNDA.n1240 GNDA.n1239 187.249
R1054 GNDA.n1014 GNDA.n449 187.249
R1055 GNDA.n1441 GNDA.n436 187.249
R1056 GNDA.n1671 GNDA.n1670 187.249
R1057 GNDA.n1718 GNDA.n367 187.249
R1058 GNDA.n1747 GNDA.n256 187.249
R1059 GNDA.n1716 GNDA.n373 187.249
R1060 GNDA.n2026 GNDA.n122 187.249
R1061 GNDA.n1841 GNDA.n1839 187.249
R1062 GNDA.n1207 GNDA.n1144 185
R1063 GNDA.n1222 GNDA.n1221 185
R1064 GNDA.n1220 GNDA.n1145 185
R1065 GNDA.n1219 GNDA.n1218 185
R1066 GNDA.n1217 GNDA.n1216 185
R1067 GNDA.n1215 GNDA.n1214 185
R1068 GNDA.n1213 GNDA.n1212 185
R1069 GNDA.n1211 GNDA.n1210 185
R1070 GNDA.n1209 GNDA.n1208 185
R1071 GNDA.n1190 GNDA.n1189 185
R1072 GNDA.n1192 GNDA.n1191 185
R1073 GNDA.n1194 GNDA.n1193 185
R1074 GNDA.n1196 GNDA.n1195 185
R1075 GNDA.n1198 GNDA.n1197 185
R1076 GNDA.n1200 GNDA.n1199 185
R1077 GNDA.n1202 GNDA.n1201 185
R1078 GNDA.n1204 GNDA.n1203 185
R1079 GNDA.n1206 GNDA.n1205 185
R1080 GNDA.n1172 GNDA.n1171 185
R1081 GNDA.n1174 GNDA.n1173 185
R1082 GNDA.n1176 GNDA.n1175 185
R1083 GNDA.n1178 GNDA.n1177 185
R1084 GNDA.n1180 GNDA.n1179 185
R1085 GNDA.n1182 GNDA.n1181 185
R1086 GNDA.n1184 GNDA.n1183 185
R1087 GNDA.n1186 GNDA.n1185 185
R1088 GNDA.n1188 GNDA.n1187 185
R1089 GNDA.n1170 GNDA.n1169 185
R1090 GNDA.n1160 GNDA.n1159 185
R1091 GNDA.n1158 GNDA.n1157 185
R1092 GNDA.n1155 GNDA.n1154 185
R1093 GNDA.n1149 GNDA.n1129 185
R1094 GNDA.n1226 GNDA.n1225 185
R1095 GNDA.n1128 GNDA.n1125 185
R1096 GNDA.n1233 GNDA.n1232 185
R1097 GNDA.n1235 GNDA.n1234 185
R1098 GNDA.n982 GNDA.n981 185
R1099 GNDA.n983 GNDA.n905 185
R1100 GNDA.n985 GNDA.n984 185
R1101 GNDA.n987 GNDA.n904 185
R1102 GNDA.n990 GNDA.n989 185
R1103 GNDA.n991 GNDA.n903 185
R1104 GNDA.n993 GNDA.n992 185
R1105 GNDA.n995 GNDA.n902 185
R1106 GNDA.n996 GNDA.n451 185
R1107 GNDA.n963 GNDA.n910 185
R1108 GNDA.n966 GNDA.n965 185
R1109 GNDA.n967 GNDA.n909 185
R1110 GNDA.n969 GNDA.n968 185
R1111 GNDA.n971 GNDA.n908 185
R1112 GNDA.n974 GNDA.n973 185
R1113 GNDA.n975 GNDA.n907 185
R1114 GNDA.n977 GNDA.n976 185
R1115 GNDA.n979 GNDA.n906 185
R1116 GNDA.n947 GNDA.n946 185
R1117 GNDA.n949 GNDA.n915 185
R1118 GNDA.n951 GNDA.n950 185
R1119 GNDA.n952 GNDA.n914 185
R1120 GNDA.n954 GNDA.n953 185
R1121 GNDA.n956 GNDA.n912 185
R1122 GNDA.n958 GNDA.n957 185
R1123 GNDA.n959 GNDA.n911 185
R1124 GNDA.n961 GNDA.n960 185
R1125 GNDA.n918 GNDA.n917 185
R1126 GNDA.n938 GNDA.n937 185
R1127 GNDA.n935 GNDA.n920 185
R1128 GNDA.n933 GNDA.n932 185
R1129 GNDA.n924 GNDA.n922 185
R1130 GNDA.n923 GNDA.n901 185
R1131 GNDA.n1002 GNDA.n1001 185
R1132 GNDA.n999 GNDA.n899 185
R1133 GNDA.n998 GNDA.n452 185
R1134 GNDA.n1423 GNDA.n1422 185
R1135 GNDA.n1425 GNDA.n1424 185
R1136 GNDA.n1427 GNDA.n1426 185
R1137 GNDA.n1429 GNDA.n1428 185
R1138 GNDA.n1431 GNDA.n1430 185
R1139 GNDA.n1433 GNDA.n1432 185
R1140 GNDA.n1435 GNDA.n1434 185
R1141 GNDA.n1437 GNDA.n1436 185
R1142 GNDA.n1438 GNDA.n423 185
R1143 GNDA.n1405 GNDA.n1404 185
R1144 GNDA.n1407 GNDA.n1406 185
R1145 GNDA.n1409 GNDA.n1408 185
R1146 GNDA.n1411 GNDA.n1410 185
R1147 GNDA.n1413 GNDA.n1412 185
R1148 GNDA.n1415 GNDA.n1414 185
R1149 GNDA.n1417 GNDA.n1416 185
R1150 GNDA.n1419 GNDA.n1418 185
R1151 GNDA.n1421 GNDA.n1420 185
R1152 GNDA.n415 GNDA.n398 185
R1153 GNDA.n1389 GNDA.n1388 185
R1154 GNDA.n1391 GNDA.n1390 185
R1155 GNDA.n1393 GNDA.n1392 185
R1156 GNDA.n1395 GNDA.n1394 185
R1157 GNDA.n1397 GNDA.n1396 185
R1158 GNDA.n1399 GNDA.n1398 185
R1159 GNDA.n1401 GNDA.n1400 185
R1160 GNDA.n1403 GNDA.n1402 185
R1161 GNDA.n405 GNDA.n399 185
R1162 GNDA.n1474 GNDA.n1473 185
R1163 GNDA.n404 GNDA.n402 185
R1164 GNDA.n1455 GNDA.n1454 185
R1165 GNDA.n1457 GNDA.n1456 185
R1166 GNDA.n1461 GNDA.n1460 185
R1167 GNDA.n1459 GNDA.n1447 185
R1168 GNDA.n426 GNDA.n424 185
R1169 GNDA.n1470 GNDA.n1469 185
R1170 GNDA.n1651 GNDA.n1650 185
R1171 GNDA.n1653 GNDA.n1652 185
R1172 GNDA.n1655 GNDA.n1654 185
R1173 GNDA.n1657 GNDA.n1656 185
R1174 GNDA.n1659 GNDA.n1658 185
R1175 GNDA.n1661 GNDA.n1660 185
R1176 GNDA.n1663 GNDA.n1662 185
R1177 GNDA.n1665 GNDA.n1664 185
R1178 GNDA.n1666 GNDA.n75 185
R1179 GNDA.n1633 GNDA.n1632 185
R1180 GNDA.n1635 GNDA.n1634 185
R1181 GNDA.n1637 GNDA.n1636 185
R1182 GNDA.n1639 GNDA.n1638 185
R1183 GNDA.n1641 GNDA.n1640 185
R1184 GNDA.n1643 GNDA.n1642 185
R1185 GNDA.n1645 GNDA.n1644 185
R1186 GNDA.n1647 GNDA.n1646 185
R1187 GNDA.n1649 GNDA.n1648 185
R1188 GNDA.n1615 GNDA.n1614 185
R1189 GNDA.n1617 GNDA.n1616 185
R1190 GNDA.n1619 GNDA.n1618 185
R1191 GNDA.n1621 GNDA.n1620 185
R1192 GNDA.n1623 GNDA.n1622 185
R1193 GNDA.n1625 GNDA.n1624 185
R1194 GNDA.n1627 GNDA.n1626 185
R1195 GNDA.n1629 GNDA.n1628 185
R1196 GNDA.n1631 GNDA.n1630 185
R1197 GNDA.n1613 GNDA.n1612 185
R1198 GNDA.n1604 GNDA.n1603 185
R1199 GNDA.n1602 GNDA.n58 185
R1200 GNDA.n2080 GNDA.n2079 185
R1201 GNDA.n2063 GNDA.n57 185
R1202 GNDA.n2067 GNDA.n2066 185
R1203 GNDA.n2065 GNDA.n2062 185
R1204 GNDA.n78 GNDA.n76 185
R1205 GNDA.n2076 GNDA.n2075 185
R1206 GNDA.n862 GNDA.n801 185
R1207 GNDA.n877 GNDA.n876 185
R1208 GNDA.n875 GNDA.n802 185
R1209 GNDA.n874 GNDA.n873 185
R1210 GNDA.n872 GNDA.n871 185
R1211 GNDA.n870 GNDA.n869 185
R1212 GNDA.n868 GNDA.n867 185
R1213 GNDA.n866 GNDA.n865 185
R1214 GNDA.n864 GNDA.n863 185
R1215 GNDA.n845 GNDA.n844 185
R1216 GNDA.n847 GNDA.n846 185
R1217 GNDA.n849 GNDA.n848 185
R1218 GNDA.n851 GNDA.n850 185
R1219 GNDA.n853 GNDA.n852 185
R1220 GNDA.n855 GNDA.n854 185
R1221 GNDA.n857 GNDA.n856 185
R1222 GNDA.n859 GNDA.n858 185
R1223 GNDA.n861 GNDA.n860 185
R1224 GNDA.n827 GNDA.n826 185
R1225 GNDA.n829 GNDA.n828 185
R1226 GNDA.n831 GNDA.n830 185
R1227 GNDA.n833 GNDA.n832 185
R1228 GNDA.n835 GNDA.n834 185
R1229 GNDA.n837 GNDA.n836 185
R1230 GNDA.n839 GNDA.n838 185
R1231 GNDA.n841 GNDA.n840 185
R1232 GNDA.n843 GNDA.n842 185
R1233 GNDA.n825 GNDA.n824 185
R1234 GNDA.n819 GNDA.n818 185
R1235 GNDA.n817 GNDA.n816 185
R1236 GNDA.n812 GNDA.n811 185
R1237 GNDA.n807 GNDA.n786 185
R1238 GNDA.n881 GNDA.n880 185
R1239 GNDA.n785 GNDA.n783 185
R1240 GNDA.n887 GNDA.n886 185
R1241 GNDA.n889 GNDA.n888 185
R1242 GNDA.n319 GNDA.n318 185
R1243 GNDA.n321 GNDA.n276 185
R1244 GNDA.n324 GNDA.n323 185
R1245 GNDA.n325 GNDA.n275 185
R1246 GNDA.n327 GNDA.n326 185
R1247 GNDA.n329 GNDA.n274 185
R1248 GNDA.n332 GNDA.n331 185
R1249 GNDA.n333 GNDA.n273 185
R1250 GNDA.n1752 GNDA.n1751 185
R1251 GNDA.n301 GNDA.n281 185
R1252 GNDA.n303 GNDA.n302 185
R1253 GNDA.n305 GNDA.n280 185
R1254 GNDA.n308 GNDA.n307 185
R1255 GNDA.n309 GNDA.n279 185
R1256 GNDA.n311 GNDA.n310 185
R1257 GNDA.n313 GNDA.n278 185
R1258 GNDA.n316 GNDA.n315 185
R1259 GNDA.n317 GNDA.n277 185
R1260 GNDA.n1786 GNDA.n1785 185
R1261 GNDA.n286 GNDA.n261 185
R1262 GNDA.n288 GNDA.n287 185
R1263 GNDA.n290 GNDA.n284 185
R1264 GNDA.n292 GNDA.n291 185
R1265 GNDA.n293 GNDA.n283 185
R1266 GNDA.n295 GNDA.n294 185
R1267 GNDA.n297 GNDA.n282 185
R1268 GNDA.n300 GNDA.n299 185
R1269 GNDA.n1784 GNDA.n260 185
R1270 GNDA.n1782 GNDA.n1781 185
R1271 GNDA.n264 GNDA.n263 185
R1272 GNDA.n1772 GNDA.n1771 185
R1273 GNDA.n1769 GNDA.n267 185
R1274 GNDA.n1767 GNDA.n1766 185
R1275 GNDA.n269 GNDA.n268 185
R1276 GNDA.n1757 GNDA.n1756 185
R1277 GNDA.n1754 GNDA.n272 185
R1278 GNDA.n741 GNDA.n483 185
R1279 GNDA.n756 GNDA.n755 185
R1280 GNDA.n754 GNDA.n484 185
R1281 GNDA.n753 GNDA.n752 185
R1282 GNDA.n751 GNDA.n750 185
R1283 GNDA.n749 GNDA.n748 185
R1284 GNDA.n747 GNDA.n746 185
R1285 GNDA.n745 GNDA.n744 185
R1286 GNDA.n743 GNDA.n742 185
R1287 GNDA.n724 GNDA.n723 185
R1288 GNDA.n726 GNDA.n725 185
R1289 GNDA.n728 GNDA.n727 185
R1290 GNDA.n730 GNDA.n729 185
R1291 GNDA.n732 GNDA.n731 185
R1292 GNDA.n734 GNDA.n733 185
R1293 GNDA.n736 GNDA.n735 185
R1294 GNDA.n738 GNDA.n737 185
R1295 GNDA.n740 GNDA.n739 185
R1296 GNDA.n706 GNDA.n705 185
R1297 GNDA.n708 GNDA.n707 185
R1298 GNDA.n710 GNDA.n709 185
R1299 GNDA.n712 GNDA.n711 185
R1300 GNDA.n714 GNDA.n713 185
R1301 GNDA.n716 GNDA.n715 185
R1302 GNDA.n718 GNDA.n717 185
R1303 GNDA.n720 GNDA.n719 185
R1304 GNDA.n722 GNDA.n721 185
R1305 GNDA.n704 GNDA.n703 185
R1306 GNDA.n698 GNDA.n697 185
R1307 GNDA.n696 GNDA.n695 185
R1308 GNDA.n691 GNDA.n690 185
R1309 GNDA.n686 GNDA.n468 185
R1310 GNDA.n760 GNDA.n759 185
R1311 GNDA.n467 GNDA.n465 185
R1312 GNDA.n766 GNDA.n765 185
R1313 GNDA.n768 GNDA.n767 185
R1314 GNDA.n2008 GNDA.n2007 185
R1315 GNDA.n2010 GNDA.n2009 185
R1316 GNDA.n2012 GNDA.n2011 185
R1317 GNDA.n2014 GNDA.n2013 185
R1318 GNDA.n2016 GNDA.n2015 185
R1319 GNDA.n2018 GNDA.n2017 185
R1320 GNDA.n2020 GNDA.n2019 185
R1321 GNDA.n2022 GNDA.n2021 185
R1322 GNDA.n2023 GNDA.n111 185
R1323 GNDA.n1990 GNDA.n1989 185
R1324 GNDA.n1992 GNDA.n1991 185
R1325 GNDA.n1994 GNDA.n1993 185
R1326 GNDA.n1996 GNDA.n1995 185
R1327 GNDA.n1998 GNDA.n1997 185
R1328 GNDA.n2000 GNDA.n1999 185
R1329 GNDA.n2002 GNDA.n2001 185
R1330 GNDA.n2004 GNDA.n2003 185
R1331 GNDA.n2006 GNDA.n2005 185
R1332 GNDA.n1972 GNDA.n1971 185
R1333 GNDA.n1974 GNDA.n1973 185
R1334 GNDA.n1976 GNDA.n1975 185
R1335 GNDA.n1978 GNDA.n1977 185
R1336 GNDA.n1980 GNDA.n1979 185
R1337 GNDA.n1982 GNDA.n1981 185
R1338 GNDA.n1984 GNDA.n1983 185
R1339 GNDA.n1986 GNDA.n1985 185
R1340 GNDA.n1988 GNDA.n1987 185
R1341 GNDA.n1970 GNDA.n1969 185
R1342 GNDA.n131 GNDA.n130 185
R1343 GNDA.n129 GNDA.n94 185
R1344 GNDA.n2049 GNDA.n2048 185
R1345 GNDA.n2032 GNDA.n93 185
R1346 GNDA.n2036 GNDA.n2035 185
R1347 GNDA.n2034 GNDA.n2031 185
R1348 GNDA.n114 GNDA.n112 185
R1349 GNDA.n2045 GNDA.n2044 185
R1350 GNDA.n237 GNDA.n236 185
R1351 GNDA.n239 GNDA.n194 185
R1352 GNDA.n242 GNDA.n241 185
R1353 GNDA.n243 GNDA.n193 185
R1354 GNDA.n245 GNDA.n244 185
R1355 GNDA.n247 GNDA.n192 185
R1356 GNDA.n250 GNDA.n249 185
R1357 GNDA.n251 GNDA.n191 185
R1358 GNDA.n1846 GNDA.n1845 185
R1359 GNDA.n219 GNDA.n199 185
R1360 GNDA.n221 GNDA.n220 185
R1361 GNDA.n223 GNDA.n198 185
R1362 GNDA.n226 GNDA.n225 185
R1363 GNDA.n227 GNDA.n197 185
R1364 GNDA.n229 GNDA.n228 185
R1365 GNDA.n231 GNDA.n196 185
R1366 GNDA.n234 GNDA.n233 185
R1367 GNDA.n235 GNDA.n195 185
R1368 GNDA.n1880 GNDA.n1879 185
R1369 GNDA.n204 GNDA.n179 185
R1370 GNDA.n206 GNDA.n205 185
R1371 GNDA.n208 GNDA.n202 185
R1372 GNDA.n210 GNDA.n209 185
R1373 GNDA.n211 GNDA.n201 185
R1374 GNDA.n213 GNDA.n212 185
R1375 GNDA.n215 GNDA.n200 185
R1376 GNDA.n218 GNDA.n217 185
R1377 GNDA.n1878 GNDA.n178 185
R1378 GNDA.n1876 GNDA.n1875 185
R1379 GNDA.n182 GNDA.n181 185
R1380 GNDA.n1866 GNDA.n1865 185
R1381 GNDA.n1863 GNDA.n185 185
R1382 GNDA.n1861 GNDA.n1860 185
R1383 GNDA.n187 GNDA.n186 185
R1384 GNDA.n1851 GNDA.n1850 185
R1385 GNDA.n1848 GNDA.n190 185
R1386 GNDA.n1097 GNDA.n1030 183.948
R1387 GNDA.n1938 GNDA.n1937 183.948
R1388 GNDA.n1047 GNDA.n1030 180.013
R1389 GNDA.n1937 GNDA.n1936 180.013
R1390 GNDA.n1017 GNDA.n1016 175.546
R1391 GNDA.n1257 GNDA.n1016 175.546
R1392 GNDA.n1255 GNDA.n1254 175.546
R1393 GNDA.n1251 GNDA.n1250 175.546
R1394 GNDA.n1247 GNDA.n1246 175.546
R1395 GNDA.n1243 GNDA.n1242 175.546
R1396 GNDA.n1116 GNDA.n1018 175.546
R1397 GNDA.n1116 GNDA.n1020 175.546
R1398 GNDA.n1112 GNDA.n1020 175.546
R1399 GNDA.n1112 GNDA.n1023 175.546
R1400 GNDA.n1108 GNDA.n1023 175.546
R1401 GNDA.n1108 GNDA.n1025 175.546
R1402 GNDA.n1104 GNDA.n1025 175.546
R1403 GNDA.n1104 GNDA.n1027 175.546
R1404 GNDA.n1100 GNDA.n1027 175.546
R1405 GNDA.n1100 GNDA.n1029 175.546
R1406 GNDA.n1096 GNDA.n1029 175.546
R1407 GNDA.n1237 GNDA.n1120 175.546
R1408 GNDA.n1230 GNDA.n1228 175.546
R1409 GNDA.n1152 GNDA.n1150 175.546
R1410 GNDA.n1162 GNDA.n1148 175.546
R1411 GNDA.n1167 GNDA.n1164 175.546
R1412 GNDA.n1050 GNDA.n1031 175.546
R1413 GNDA.n1051 GNDA.n1050 175.546
R1414 GNDA.n1054 GNDA.n1051 175.546
R1415 GNDA.n1055 GNDA.n1054 175.546
R1416 GNDA.n1081 GNDA.n1055 175.546
R1417 GNDA.n1081 GNDA.n1080 175.546
R1418 GNDA.n1080 GNDA.n1058 175.546
R1419 GNDA.n1062 GNDA.n1058 175.546
R1420 GNDA.n1063 GNDA.n1062 175.546
R1421 GNDA.n1067 GNDA.n1063 175.546
R1422 GNDA.n1068 GNDA.n1067 175.546
R1423 GNDA.n620 GNDA.n619 175.546
R1424 GNDA.n616 GNDA.n615 175.546
R1425 GNDA.n612 GNDA.n611 175.546
R1426 GNDA.n608 GNDA.n607 175.546
R1427 GNDA.n604 GNDA.n603 175.546
R1428 GNDA.n628 GNDA.n627 175.546
R1429 GNDA.n632 GNDA.n631 175.546
R1430 GNDA.n636 GNDA.n635 175.546
R1431 GNDA.n640 GNDA.n639 175.546
R1432 GNDA.n644 GNDA.n602 175.546
R1433 GNDA.n1008 GNDA.n453 175.546
R1434 GNDA.n1004 GNDA.n897 175.546
R1435 GNDA.n927 GNDA.n926 175.546
R1436 GNDA.n930 GNDA.n929 175.546
R1437 GNDA.n941 GNDA.n940 175.546
R1438 GNDA.n357 GNDA.n348 175.546
R1439 GNDA.n350 GNDA.n349 175.546
R1440 GNDA.n352 GNDA.n351 175.546
R1441 GNDA.n354 GNDA.n353 175.546
R1442 GNDA.n356 GNDA.n355 175.546
R1443 GNDA.n1369 GNDA.n1367 175.546
R1444 GNDA.n1373 GNDA.n1268 175.546
R1445 GNDA.n1377 GNDA.n1375 175.546
R1446 GNDA.n1381 GNDA.n1266 175.546
R1447 GNDA.n1384 GNDA.n1383 175.546
R1448 GNDA.n1361 GNDA.n1360 175.546
R1449 GNDA.n1358 GNDA.n1273 175.546
R1450 GNDA.n1354 GNDA.n1353 175.546
R1451 GNDA.n1351 GNDA.n1276 175.546
R1452 GNDA.n1347 GNDA.n1346 175.546
R1453 GNDA.n1441 GNDA.n427 175.546
R1454 GNDA.n1467 GNDA.n427 175.546
R1455 GNDA.n1467 GNDA.n428 175.546
R1456 GNDA.n1463 GNDA.n428 175.546
R1457 GNDA.n1463 GNDA.n1445 175.546
R1458 GNDA.n1451 GNDA.n1445 175.546
R1459 GNDA.n1451 GNDA.n401 175.546
R1460 GNDA.n1476 GNDA.n401 175.546
R1461 GNDA.n1476 GNDA.n400 175.546
R1462 GNDA.n1481 GNDA.n400 175.546
R1463 GNDA.n1481 GNDA.n392 175.546
R1464 GNDA.n1310 GNDA.n1309 175.546
R1465 GNDA.n1315 GNDA.n1312 175.546
R1466 GNDA.n1318 GNDA.n1317 175.546
R1467 GNDA.n1322 GNDA.n1320 175.546
R1468 GNDA.n1676 GNDA.n395 175.546
R1469 GNDA.n1338 GNDA.n1337 175.546
R1470 GNDA.n1334 GNDA.n1333 175.546
R1471 GNDA.n1331 GNDA.n1314 175.546
R1472 GNDA.n1327 GNDA.n1325 175.546
R1473 GNDA.n1674 GNDA.n397 175.546
R1474 GNDA.n1304 GNDA.n1282 175.546
R1475 GNDA.n1300 GNDA.n1299 175.546
R1476 GNDA.n1297 GNDA.n1285 175.546
R1477 GNDA.n1293 GNDA.n1292 175.546
R1478 GNDA.n1290 GNDA.n1288 175.546
R1479 GNDA.n1670 GNDA.n79 175.546
R1480 GNDA.n2073 GNDA.n79 175.546
R1481 GNDA.n2073 GNDA.n80 175.546
R1482 GNDA.n2069 GNDA.n80 175.546
R1483 GNDA.n2069 GNDA.n54 175.546
R1484 GNDA.n2082 GNDA.n54 175.546
R1485 GNDA.n2082 GNDA.n55 175.546
R1486 GNDA.n1606 GNDA.n55 175.546
R1487 GNDA.n1606 GNDA.n1488 175.546
R1488 GNDA.n1610 GNDA.n1488 175.546
R1489 GNDA.n1610 GNDA.n1600 175.546
R1490 GNDA.n1500 GNDA.n379 175.546
R1491 GNDA.n1576 GNDA.n1575 175.546
R1492 GNDA.n1497 GNDA.n1496 175.546
R1493 GNDA.n1586 GNDA.n1585 175.546
R1494 GNDA.n1492 GNDA.n1491 175.546
R1495 GNDA.n1737 GNDA.n341 175.546
R1496 GNDA.n1733 GNDA.n347 175.546
R1497 GNDA.n1731 GNDA.n1730 175.546
R1498 GNDA.n1727 GNDA.n1726 175.546
R1499 GNDA.n1723 GNDA.n1722 175.546
R1500 GNDA.n512 GNDA.n511 175.546
R1501 GNDA.n516 GNDA.n515 175.546
R1502 GNDA.n520 GNDA.n519 175.546
R1503 GNDA.n524 GNDA.n523 175.546
R1504 GNDA.n526 GNDA.n508 175.546
R1505 GNDA.n891 GNDA.n777 175.546
R1506 GNDA.n884 GNDA.n883 175.546
R1507 GNDA.n809 GNDA.n808 175.546
R1508 GNDA.n814 GNDA.n813 175.546
R1509 GNDA.n822 GNDA.n821 175.546
R1510 GNDA.n562 GNDA.n553 175.546
R1511 GNDA.n555 GNDA.n554 175.546
R1512 GNDA.n557 GNDA.n556 175.546
R1513 GNDA.n559 GNDA.n558 175.546
R1514 GNDA.n561 GNDA.n560 175.546
R1515 GNDA.n1092 GNDA.n1049 175.546
R1516 GNDA.n1088 GNDA.n1049 175.546
R1517 GNDA.n1088 GNDA.n1053 175.546
R1518 GNDA.n1084 GNDA.n1053 175.546
R1519 GNDA.n1084 GNDA.n1057 175.546
R1520 GNDA.n1078 GNDA.n1057 175.546
R1521 GNDA.n1078 GNDA.n1077 175.546
R1522 GNDA.n1077 GNDA.n1061 175.546
R1523 GNDA.n1073 GNDA.n1061 175.546
R1524 GNDA.n1073 GNDA.n1065 175.546
R1525 GNDA.n1069 GNDA.n1065 175.546
R1526 GNDA.n1048 GNDA.n1034 175.546
R1527 GNDA.n1044 GNDA.n1034 175.546
R1528 GNDA.n1044 GNDA.n1036 175.546
R1529 GNDA.n1040 GNDA.n1036 175.546
R1530 GNDA.n1040 GNDA.n142 175.546
R1531 GNDA.n1948 GNDA.n142 175.546
R1532 GNDA.n1948 GNDA.n143 175.546
R1533 GNDA.n1944 GNDA.n143 175.546
R1534 GNDA.n1944 GNDA.n145 175.546
R1535 GNDA.n1940 GNDA.n145 175.546
R1536 GNDA.n1940 GNDA.n147 175.546
R1537 GNDA.n1759 GNDA.n271 175.546
R1538 GNDA.n1763 GNDA.n1761 175.546
R1539 GNDA.n1774 GNDA.n266 175.546
R1540 GNDA.n1778 GNDA.n1776 175.546
R1541 GNDA.n1789 GNDA.n259 175.546
R1542 GNDA.n1809 GNDA.n1808 175.546
R1543 GNDA.n1809 GNDA.n1805 175.546
R1544 GNDA.n1815 GNDA.n1805 175.546
R1545 GNDA.n1815 GNDA.n1801 175.546
R1546 GNDA.n1821 GNDA.n1801 175.546
R1547 GNDA.n1823 GNDA.n1821 175.546
R1548 GNDA.n1823 GNDA.n1797 175.546
R1549 GNDA.n1829 GNDA.n1797 175.546
R1550 GNDA.n1830 GNDA.n1829 175.546
R1551 GNDA.n1830 GNDA.n1792 175.546
R1552 GNDA.n1836 GNDA.n1792 175.546
R1553 GNDA.n588 GNDA.n547 175.546
R1554 GNDA.n588 GNDA.n552 175.546
R1555 GNDA.n584 GNDA.n583 175.546
R1556 GNDA.n580 GNDA.n579 175.546
R1557 GNDA.n576 GNDA.n575 175.546
R1558 GNDA.n572 GNDA.n372 175.546
R1559 GNDA.n542 GNDA.n541 175.546
R1560 GNDA.n538 GNDA.n537 175.546
R1561 GNDA.n534 GNDA.n533 175.546
R1562 GNDA.n530 GNDA.n498 175.546
R1563 GNDA.n650 GNDA.n649 175.546
R1564 GNDA.n770 GNDA.n459 175.546
R1565 GNDA.n763 GNDA.n762 175.546
R1566 GNDA.n688 GNDA.n687 175.546
R1567 GNDA.n693 GNDA.n692 175.546
R1568 GNDA.n701 GNDA.n700 175.546
R1569 GNDA.n657 GNDA.n654 175.546
R1570 GNDA.n657 GNDA.n494 175.546
R1571 GNDA.n662 GNDA.n494 175.546
R1572 GNDA.n662 GNDA.n491 175.546
R1573 GNDA.n666 GNDA.n491 175.546
R1574 GNDA.n667 GNDA.n666 175.546
R1575 GNDA.n670 GNDA.n667 175.546
R1576 GNDA.n670 GNDA.n489 175.546
R1577 GNDA.n675 GNDA.n489 175.546
R1578 GNDA.n675 GNDA.n487 175.546
R1579 GNDA.n679 GNDA.n487 175.546
R1580 GNDA.n1572 GNDA.n1570 175.546
R1581 GNDA.n1578 GNDA.n1498 175.546
R1582 GNDA.n1582 GNDA.n1580 175.546
R1583 GNDA.n1588 GNDA.n1494 175.546
R1584 GNDA.n1591 GNDA.n1590 175.546
R1585 GNDA.n1565 GNDA.n1501 175.546
R1586 GNDA.n1561 GNDA.n1560 175.546
R1587 GNDA.n1558 GNDA.n1504 175.546
R1588 GNDA.n1554 GNDA.n1553 175.546
R1589 GNDA.n1551 GNDA.n1507 175.546
R1590 GNDA.n2026 GNDA.n115 175.546
R1591 GNDA.n2042 GNDA.n115 175.546
R1592 GNDA.n2042 GNDA.n116 175.546
R1593 GNDA.n2038 GNDA.n116 175.546
R1594 GNDA.n2038 GNDA.n90 175.546
R1595 GNDA.n2051 GNDA.n90 175.546
R1596 GNDA.n2051 GNDA.n91 175.546
R1597 GNDA.n133 GNDA.n91 175.546
R1598 GNDA.n133 GNDA.n126 175.546
R1599 GNDA.n1967 GNDA.n126 175.546
R1600 GNDA.n1967 GNDA.n127 175.546
R1601 GNDA.n1546 GNDA.n1510 175.546
R1602 GNDA.n1542 GNDA.n1510 175.546
R1603 GNDA.n1542 GNDA.n1512 175.546
R1604 GNDA.n1538 GNDA.n1512 175.546
R1605 GNDA.n1538 GNDA.n1536 175.546
R1606 GNDA.n1536 GNDA.n1535 175.546
R1607 GNDA.n1535 GNDA.n1515 175.546
R1608 GNDA.n1531 GNDA.n1515 175.546
R1609 GNDA.n1531 GNDA.n1517 175.546
R1610 GNDA.n1527 GNDA.n1517 175.546
R1611 GNDA.n1527 GNDA.n1520 175.546
R1612 GNDA.n1811 GNDA.n150 175.546
R1613 GNDA.n1812 GNDA.n1811 175.546
R1614 GNDA.n1812 GNDA.n1803 175.546
R1615 GNDA.n1818 GNDA.n1803 175.546
R1616 GNDA.n1819 GNDA.n1818 175.546
R1617 GNDA.n1819 GNDA.n1799 175.546
R1618 GNDA.n1826 GNDA.n1799 175.546
R1619 GNDA.n1827 GNDA.n1826 175.546
R1620 GNDA.n1827 GNDA.n1795 175.546
R1621 GNDA.n1833 GNDA.n1795 175.546
R1622 GNDA.n1833 GNDA.n253 175.546
R1623 GNDA.n1935 GNDA.n151 175.546
R1624 GNDA.n1931 GNDA.n151 175.546
R1625 GNDA.n1931 GNDA.n154 175.546
R1626 GNDA.n1927 GNDA.n154 175.546
R1627 GNDA.n1927 GNDA.n156 175.546
R1628 GNDA.n1923 GNDA.n156 175.546
R1629 GNDA.n1923 GNDA.n158 175.546
R1630 GNDA.n1919 GNDA.n158 175.546
R1631 GNDA.n1919 GNDA.n160 175.546
R1632 GNDA.n1915 GNDA.n160 175.546
R1633 GNDA.n1915 GNDA.n162 175.546
R1634 GNDA.n1853 GNDA.n189 175.546
R1635 GNDA.n1857 GNDA.n1855 175.546
R1636 GNDA.n1868 GNDA.n184 175.546
R1637 GNDA.n1872 GNDA.n1870 175.546
R1638 GNDA.n1883 GNDA.n177 175.546
R1639 GNDA.n1911 GNDA.n164 175.546
R1640 GNDA.n1907 GNDA.n164 175.546
R1641 GNDA.n1907 GNDA.n166 175.546
R1642 GNDA.n1903 GNDA.n166 175.546
R1643 GNDA.n1903 GNDA.n168 175.546
R1644 GNDA.n1899 GNDA.n168 175.546
R1645 GNDA.n1899 GNDA.n170 175.546
R1646 GNDA.n1895 GNDA.n170 175.546
R1647 GNDA.n1895 GNDA.n172 175.546
R1648 GNDA.n1891 GNDA.n172 175.546
R1649 GNDA.n1891 GNDA.n174 175.546
R1650 GNDA.n363 GNDA.n342 173.881
R1651 GNDA.n568 GNDA.t199 172.876
R1652 GNDA.n589 GNDA.t199 172.615
R1653 GNDA.n1739 GNDA.n342 171.624
R1654 GNDA.n1171 GNDA.n1170 163.333
R1655 GNDA.n947 GNDA.n917 163.333
R1656 GNDA.n415 GNDA.n405 163.333
R1657 GNDA.n1614 GNDA.n1613 163.333
R1658 GNDA.n826 GNDA.n825 163.333
R1659 GNDA.n1785 GNDA.n1784 163.333
R1660 GNDA.n705 GNDA.n704 163.333
R1661 GNDA.n1971 GNDA.n1970 163.333
R1662 GNDA.n1879 GNDA.n1878 163.333
R1663 GNDA.n1203 GNDA.n1202 150
R1664 GNDA.n1199 GNDA.n1198 150
R1665 GNDA.n1195 GNDA.n1194 150
R1666 GNDA.n1191 GNDA.n1190 150
R1667 GNDA.n1187 GNDA.n1186 150
R1668 GNDA.n1183 GNDA.n1182 150
R1669 GNDA.n1179 GNDA.n1178 150
R1670 GNDA.n1175 GNDA.n1174 150
R1671 GNDA.n1234 GNDA.n1233 150
R1672 GNDA.n1225 GNDA.n1128 150
R1673 GNDA.n1154 GNDA.n1129 150
R1674 GNDA.n1159 GNDA.n1158 150
R1675 GNDA.n1222 GNDA.n1145 150
R1676 GNDA.n1218 GNDA.n1217 150
R1677 GNDA.n1214 GNDA.n1213 150
R1678 GNDA.n1210 GNDA.n1209 150
R1679 GNDA.n977 GNDA.n907 150
R1680 GNDA.n973 GNDA.n971 150
R1681 GNDA.n969 GNDA.n909 150
R1682 GNDA.n965 GNDA.n963 150
R1683 GNDA.n961 GNDA.n911 150
R1684 GNDA.n957 GNDA.n956 150
R1685 GNDA.n954 GNDA.n914 150
R1686 GNDA.n950 GNDA.n949 150
R1687 GNDA.n999 GNDA.n998 150
R1688 GNDA.n1001 GNDA.n901 150
R1689 GNDA.n933 GNDA.n922 150
R1690 GNDA.n937 GNDA.n935 150
R1691 GNDA.n985 GNDA.n905 150
R1692 GNDA.n989 GNDA.n987 150
R1693 GNDA.n993 GNDA.n903 150
R1694 GNDA.n996 GNDA.n995 150
R1695 GNDA.n1418 GNDA.n1417 150
R1696 GNDA.n1414 GNDA.n1413 150
R1697 GNDA.n1410 GNDA.n1409 150
R1698 GNDA.n1406 GNDA.n1405 150
R1699 GNDA.n1402 GNDA.n1401 150
R1700 GNDA.n1398 GNDA.n1397 150
R1701 GNDA.n1394 GNDA.n1393 150
R1702 GNDA.n1390 GNDA.n1389 150
R1703 GNDA.n1470 GNDA.n424 150
R1704 GNDA.n1460 GNDA.n1459 150
R1705 GNDA.n1456 GNDA.n1455 150
R1706 GNDA.n1473 GNDA.n404 150
R1707 GNDA.n1426 GNDA.n1425 150
R1708 GNDA.n1430 GNDA.n1429 150
R1709 GNDA.n1434 GNDA.n1433 150
R1710 GNDA.n1436 GNDA.n423 150
R1711 GNDA.n1646 GNDA.n1645 150
R1712 GNDA.n1642 GNDA.n1641 150
R1713 GNDA.n1638 GNDA.n1637 150
R1714 GNDA.n1634 GNDA.n1633 150
R1715 GNDA.n1630 GNDA.n1629 150
R1716 GNDA.n1626 GNDA.n1625 150
R1717 GNDA.n1622 GNDA.n1621 150
R1718 GNDA.n1618 GNDA.n1617 150
R1719 GNDA.n2076 GNDA.n76 150
R1720 GNDA.n2066 GNDA.n2065 150
R1721 GNDA.n2079 GNDA.n57 150
R1722 GNDA.n1603 GNDA.n58 150
R1723 GNDA.n1654 GNDA.n1653 150
R1724 GNDA.n1658 GNDA.n1657 150
R1725 GNDA.n1662 GNDA.n1661 150
R1726 GNDA.n1664 GNDA.n75 150
R1727 GNDA.n858 GNDA.n857 150
R1728 GNDA.n854 GNDA.n853 150
R1729 GNDA.n850 GNDA.n849 150
R1730 GNDA.n846 GNDA.n845 150
R1731 GNDA.n842 GNDA.n841 150
R1732 GNDA.n838 GNDA.n837 150
R1733 GNDA.n834 GNDA.n833 150
R1734 GNDA.n830 GNDA.n829 150
R1735 GNDA.n888 GNDA.n887 150
R1736 GNDA.n880 GNDA.n785 150
R1737 GNDA.n811 GNDA.n786 150
R1738 GNDA.n818 GNDA.n817 150
R1739 GNDA.n877 GNDA.n802 150
R1740 GNDA.n873 GNDA.n872 150
R1741 GNDA.n869 GNDA.n868 150
R1742 GNDA.n865 GNDA.n864 150
R1743 GNDA.n315 GNDA.n313 150
R1744 GNDA.n311 GNDA.n279 150
R1745 GNDA.n307 GNDA.n305 150
R1746 GNDA.n303 GNDA.n281 150
R1747 GNDA.n299 GNDA.n297 150
R1748 GNDA.n295 GNDA.n283 150
R1749 GNDA.n291 GNDA.n290 150
R1750 GNDA.n288 GNDA.n286 150
R1751 GNDA.n1756 GNDA.n1754 150
R1752 GNDA.n1767 GNDA.n268 150
R1753 GNDA.n1771 GNDA.n1769 150
R1754 GNDA.n1782 GNDA.n263 150
R1755 GNDA.n323 GNDA.n321 150
R1756 GNDA.n327 GNDA.n275 150
R1757 GNDA.n331 GNDA.n329 150
R1758 GNDA.n1752 GNDA.n273 150
R1759 GNDA.n737 GNDA.n736 150
R1760 GNDA.n733 GNDA.n732 150
R1761 GNDA.n729 GNDA.n728 150
R1762 GNDA.n725 GNDA.n724 150
R1763 GNDA.n721 GNDA.n720 150
R1764 GNDA.n717 GNDA.n716 150
R1765 GNDA.n713 GNDA.n712 150
R1766 GNDA.n709 GNDA.n708 150
R1767 GNDA.n767 GNDA.n766 150
R1768 GNDA.n759 GNDA.n467 150
R1769 GNDA.n690 GNDA.n468 150
R1770 GNDA.n697 GNDA.n696 150
R1771 GNDA.n756 GNDA.n484 150
R1772 GNDA.n752 GNDA.n751 150
R1773 GNDA.n748 GNDA.n747 150
R1774 GNDA.n744 GNDA.n743 150
R1775 GNDA.n2003 GNDA.n2002 150
R1776 GNDA.n1999 GNDA.n1998 150
R1777 GNDA.n1995 GNDA.n1994 150
R1778 GNDA.n1991 GNDA.n1990 150
R1779 GNDA.n1987 GNDA.n1986 150
R1780 GNDA.n1983 GNDA.n1982 150
R1781 GNDA.n1979 GNDA.n1978 150
R1782 GNDA.n1975 GNDA.n1974 150
R1783 GNDA.n2045 GNDA.n112 150
R1784 GNDA.n2035 GNDA.n2034 150
R1785 GNDA.n2048 GNDA.n93 150
R1786 GNDA.n130 GNDA.n94 150
R1787 GNDA.n2011 GNDA.n2010 150
R1788 GNDA.n2015 GNDA.n2014 150
R1789 GNDA.n2019 GNDA.n2018 150
R1790 GNDA.n2021 GNDA.n111 150
R1791 GNDA.n233 GNDA.n231 150
R1792 GNDA.n229 GNDA.n197 150
R1793 GNDA.n225 GNDA.n223 150
R1794 GNDA.n221 GNDA.n199 150
R1795 GNDA.n217 GNDA.n215 150
R1796 GNDA.n213 GNDA.n201 150
R1797 GNDA.n209 GNDA.n208 150
R1798 GNDA.n206 GNDA.n204 150
R1799 GNDA.n1850 GNDA.n1848 150
R1800 GNDA.n1861 GNDA.n186 150
R1801 GNDA.n1865 GNDA.n1863 150
R1802 GNDA.n1876 GNDA.n181 150
R1803 GNDA.n241 GNDA.n239 150
R1804 GNDA.n245 GNDA.n193 150
R1805 GNDA.n249 GNDA.n247 150
R1806 GNDA.n1846 GNDA.n191 150
R1807 GNDA.n2110 GNDA.n2109 148.017
R1808 GNDA.n2097 GNDA.n2096 148.017
R1809 GNDA.n2204 GNDA.n2203 148.017
R1810 GNDA.n2209 GNDA.n2208 148.017
R1811 GNDA.t44 GNDA.t96 147.84
R1812 GNDA.n432 GNDA.n431 144.701
R1813 GNDA.n430 GNDA.n429 144.701
R1814 GNDA.n391 GNDA.n390 144.701
R1815 GNDA.n1704 GNDA.n1703 144.701
R1816 GNDA.n1702 GNDA.n1701 144.701
R1817 GNDA.n1700 GNDA.n1699 144.701
R1818 GNDA.n1698 GNDA.n1697 144.701
R1819 GNDA.n1688 GNDA.n1687 144.701
R1820 GNDA.n1686 GNDA.n1685 144.701
R1821 GNDA.n138 GNDA.n137 144.701
R1822 GNDA.t66 GNDA.t311 144.321
R1823 GNDA.t151 GNDA.t307 139.041
R1824 GNDA.n1013 GNDA.n448 132.721
R1825 GNDA.n1386 GNDA.n1385 132.721
R1826 GNDA.n1068 GNDA.n257 124.832
R1827 GNDA.n370 GNDA.n365 124.832
R1828 GNDA.n1679 GNDA.n1678 124.832
R1829 GNDA.n1672 GNDA.n1671 124.832
R1830 GNDA.n1596 GNDA.n1595 124.832
R1831 GNDA.n1719 GNDA.n1718 124.832
R1832 GNDA.n570 GNDA.n371 124.832
R1833 GNDA.n1069 GNDA.n256 124.832
R1834 GNDA.n1837 GNDA.n1836 124.832
R1835 GNDA.n1716 GNDA.n372 124.832
R1836 GNDA.n1593 GNDA.n122 124.832
R1837 GNDA.n1839 GNDA.n253 124.832
R1838 GNDA.n32 GNDA.n30 124.465
R1839 GNDA.n12 GNDA.n10 124.465
R1840 GNDA.n38 GNDA.n37 123.903
R1841 GNDA.n36 GNDA.n35 123.903
R1842 GNDA.n34 GNDA.n33 123.903
R1843 GNDA.n32 GNDA.n31 123.903
R1844 GNDA.n18 GNDA.n17 123.903
R1845 GNDA.n16 GNDA.n15 123.903
R1846 GNDA.n14 GNDA.n13 123.903
R1847 GNDA.n12 GNDA.n11 123.903
R1848 GNDA.n117 GNDA.t86 122.189
R1849 GNDA.n39 GNDA.n29 119.403
R1850 GNDA.n19 GNDA.n9 119.403
R1851 GNDA.n434 GNDA.t246 116.501
R1852 GNDA.n1682 GNDA.t253 116.501
R1853 GNDA.n1707 GNDA.t274 116.501
R1854 GNDA.n1694 GNDA.t232 116.501
R1855 GNDA.n1691 GNDA.t249 116.501
R1856 GNDA.n1963 GNDA.t235 116.501
R1857 GNDA.n84 GNDA.t308 116.073
R1858 GNDA.n1957 GNDA.t89 115.105
R1859 GNDA.n84 GNDA.t312 114.635
R1860 GNDA.n1956 GNDA.t119 114.635
R1861 GNDA.t218 GNDA.n42 103.665
R1862 GNDA.n2192 GNDA.t201 103.665
R1863 GNDA.t231 GNDA.n1598 101.942
R1864 GNDA.n387 GNDA.t199 47.6748
R1865 GNDA.n1545 GNDA.t199 98.9756
R1866 GNDA.n1669 GNDA.n389 98.8538
R1867 GNDA.n2028 GNDA.n2027 92.6754
R1868 GNDA.t310 GNDA.t132 92.1471
R1869 GNDA.t303 GNDA.t310 92.1471
R1870 GNDA.t127 GNDA.t303 92.1471
R1871 GNDA.t120 GNDA.t128 92.1471
R1872 GNDA.t252 GNDA.n1479 90.616
R1873 GNDA.n655 GNDA.t90 89.6052
R1874 GNDA.n1115 GNDA.n1021 88.5317
R1875 GNDA.n1115 GNDA.n1114 88.5317
R1876 GNDA.n1114 GNDA.n1113 88.5317
R1877 GNDA.n1113 GNDA.n1022 88.5317
R1878 GNDA.n1107 GNDA.n1022 88.5317
R1879 GNDA.n1106 GNDA.n1105 88.5317
R1880 GNDA.n1105 GNDA.n1026 88.5317
R1881 GNDA.n1099 GNDA.n1026 88.5317
R1882 GNDA.n1099 GNDA.n1098 88.5317
R1883 GNDA.n1098 GNDA.n1097 88.5317
R1884 GNDA.n1047 GNDA.n1046 88.5317
R1885 GNDA.n1046 GNDA.n1045 88.5317
R1886 GNDA.n1045 GNDA.n1035 88.5317
R1887 GNDA.n1039 GNDA.n1035 88.5317
R1888 GNDA.n1039 GNDA.n1038 88.5317
R1889 GNDA.n1947 GNDA.n1946 88.5317
R1890 GNDA.n1946 GNDA.n1945 88.5317
R1891 GNDA.n1945 GNDA.n144 88.5317
R1892 GNDA.n1939 GNDA.n144 88.5317
R1893 GNDA.n1939 GNDA.n1938 88.5317
R1894 GNDA.n1936 GNDA.n149 88.5317
R1895 GNDA.n1930 GNDA.n149 88.5317
R1896 GNDA.n1930 GNDA.n1929 88.5317
R1897 GNDA.n1929 GNDA.n1928 88.5317
R1898 GNDA.n1928 GNDA.n155 88.5317
R1899 GNDA.n1922 GNDA.n1921 88.5317
R1900 GNDA.n1921 GNDA.n1920 88.5317
R1901 GNDA.n1920 GNDA.n159 88.5317
R1902 GNDA.n1914 GNDA.n159 88.5317
R1903 GNDA.n1914 GNDA.n1913 88.5317
R1904 GNDA.n2097 GNDA.t120 88.3077
R1905 GNDA.t83 GNDA.t121 84.4682
R1906 GNDA.t53 GNDA.t101 84.4682
R1907 GNDA.t93 GNDA.t69 84.4682
R1908 GNDA.t81 GNDA.t123 84.4682
R1909 GNDA.t54 GNDA.t41 84.4682
R1910 GNDA.t143 GNDA.t13 84.4682
R1911 GNDA.t94 GNDA.t15 84.4682
R1912 GNDA.t305 GNDA.t42 84.4682
R1913 GNDA.t33 GNDA.t48 84.4682
R1914 GNDA.t146 GNDA.t100 84.4682
R1915 GNDA.t98 GNDA.t99 84.4682
R1916 GNDA.t45 GNDA.t91 84.4682
R1917 GNDA.n2070 GNDA.t171 84.4377
R1918 GNDA.n1954 GNDA.n1953 84.306
R1919 GNDA.t22 GNDA.t67 82.3782
R1920 GNDA.t85 GNDA.t68 82.3782
R1921 GNDA.n1937 GNDA.n148 80.9821
R1922 GNDA.n1091 GNDA.n1030 80.9821
R1923 GNDA.t255 GNDA.t194 80.6288
R1924 GNDA.t258 GNDA.t265 80.6288
R1925 GNDA.t282 GNDA.t204 80.6288
R1926 GNDA.t285 GNDA.t209 80.6288
R1927 GNDA.n1601 GNDA.t161 80.3188
R1928 GNDA.t228 GNDA.t114 76.7893
R1929 GNDA.t9 GNDA.t270 76.7893
R1930 GNDA.n342 GNDA.t199 76.3879
R1931 GNDA.n1263 GNDA.n1262 76.3222
R1932 GNDA.n1257 GNDA.n438 76.3222
R1933 GNDA.n1254 GNDA.n439 76.3222
R1934 GNDA.n1250 GNDA.n440 76.3222
R1935 GNDA.n1246 GNDA.n441 76.3222
R1936 GNDA.n1239 GNDA.n1238 76.3222
R1937 GNDA.n1229 GNDA.n1120 76.3222
R1938 GNDA.n1228 GNDA.n1126 76.3222
R1939 GNDA.n1152 GNDA.n1151 76.3222
R1940 GNDA.n1163 GNDA.n1162 76.3222
R1941 GNDA.n1167 GNDA.n1166 76.3222
R1942 GNDA.n623 GNDA.n443 76.3222
R1943 GNDA.n619 GNDA.n444 76.3222
R1944 GNDA.n615 GNDA.n445 76.3222
R1945 GNDA.n611 GNDA.n446 76.3222
R1946 GNDA.n607 GNDA.n447 76.3222
R1947 GNDA.n603 GNDA.n448 76.3222
R1948 GNDA.n627 GNDA.n597 76.3222
R1949 GNDA.n631 GNDA.n598 76.3222
R1950 GNDA.n635 GNDA.n599 76.3222
R1951 GNDA.n639 GNDA.n600 76.3222
R1952 GNDA.n602 GNDA.n601 76.3222
R1953 GNDA.n646 GNDA.n645 76.3222
R1954 GNDA.n1007 GNDA.n449 76.3222
R1955 GNDA.n1005 GNDA.n453 76.3222
R1956 GNDA.n897 GNDA.n896 76.3222
R1957 GNDA.n927 GNDA.n895 76.3222
R1958 GNDA.n929 GNDA.n894 76.3222
R1959 GNDA.n941 GNDA.n893 76.3222
R1960 GNDA.n358 GNDA.n338 76.3222
R1961 GNDA.n359 GNDA.n348 76.3222
R1962 GNDA.n360 GNDA.n350 76.3222
R1963 GNDA.n361 GNDA.n352 76.3222
R1964 GNDA.n362 GNDA.n354 76.3222
R1965 GNDA.n364 GNDA.n356 76.3222
R1966 GNDA.n1366 GNDA.n1365 76.3222
R1967 GNDA.n1369 GNDA.n1368 76.3222
R1968 GNDA.n1374 GNDA.n1373 76.3222
R1969 GNDA.n1377 GNDA.n1376 76.3222
R1970 GNDA.n1382 GNDA.n1381 76.3222
R1971 GNDA.n1385 GNDA.n1384 76.3222
R1972 GNDA.n1361 GNDA.n1272 76.3222
R1973 GNDA.n1359 GNDA.n1358 76.3222
R1974 GNDA.n1354 GNDA.n1275 76.3222
R1975 GNDA.n1352 GNDA.n1351 76.3222
R1976 GNDA.n1347 GNDA.n1278 76.3222
R1977 GNDA.n1345 GNDA.n1344 76.3222
R1978 GNDA.n1308 GNDA.n1279 76.3222
R1979 GNDA.n1311 GNDA.n1310 76.3222
R1980 GNDA.n1316 GNDA.n1315 76.3222
R1981 GNDA.n1319 GNDA.n1318 76.3222
R1982 GNDA.n1322 GNDA.n1321 76.3222
R1983 GNDA.n1677 GNDA.n1676 76.3222
R1984 GNDA.n1340 GNDA.n1339 76.3222
R1985 GNDA.n1337 GNDA.n1307 76.3222
R1986 GNDA.n1333 GNDA.n1332 76.3222
R1987 GNDA.n1326 GNDA.n1314 76.3222
R1988 GNDA.n1325 GNDA.n1324 76.3222
R1989 GNDA.n1674 GNDA.n1673 76.3222
R1990 GNDA.n1305 GNDA.n1304 76.3222
R1991 GNDA.n1300 GNDA.n1284 76.3222
R1992 GNDA.n1298 GNDA.n1297 76.3222
R1993 GNDA.n1293 GNDA.n1287 76.3222
R1994 GNDA.n1291 GNDA.n1290 76.3222
R1995 GNDA.n1712 GNDA.n378 76.3222
R1996 GNDA.n1711 GNDA.n1710 76.3222
R1997 GNDA.n1500 GNDA.n380 76.3222
R1998 GNDA.n1576 GNDA.n381 76.3222
R1999 GNDA.n1497 GNDA.n382 76.3222
R2000 GNDA.n1586 GNDA.n383 76.3222
R2001 GNDA.n1491 GNDA.n384 76.3222
R2002 GNDA.n1741 GNDA.n1740 76.3222
R2003 GNDA.n1738 GNDA.n1737 76.3222
R2004 GNDA.n1733 GNDA.n346 76.3222
R2005 GNDA.n1730 GNDA.n345 76.3222
R2006 GNDA.n1726 GNDA.n344 76.3222
R2007 GNDA.n1722 GNDA.n343 76.3222
R2008 GNDA.n511 GNDA.n503 76.3222
R2009 GNDA.n515 GNDA.n504 76.3222
R2010 GNDA.n519 GNDA.n505 76.3222
R2011 GNDA.n523 GNDA.n506 76.3222
R2012 GNDA.n526 GNDA.n507 76.3222
R2013 GNDA.n596 GNDA.n595 76.3222
R2014 GNDA.n892 GNDA.n367 76.3222
R2015 GNDA.n777 GNDA.n776 76.3222
R2016 GNDA.n883 GNDA.n775 76.3222
R2017 GNDA.n809 GNDA.n774 76.3222
R2018 GNDA.n813 GNDA.n773 76.3222
R2019 GNDA.n822 GNDA.n772 76.3222
R2020 GNDA.n563 GNDA.n509 76.3222
R2021 GNDA.n564 GNDA.n553 76.3222
R2022 GNDA.n565 GNDA.n555 76.3222
R2023 GNDA.n566 GNDA.n557 76.3222
R2024 GNDA.n567 GNDA.n559 76.3222
R2025 GNDA.n569 GNDA.n561 76.3222
R2026 GNDA.n1747 GNDA.n1746 76.3222
R2027 GNDA.n1760 GNDA.n1759 76.3222
R2028 GNDA.n1763 GNDA.n1762 76.3222
R2029 GNDA.n1775 GNDA.n1774 76.3222
R2030 GNDA.n1778 GNDA.n1777 76.3222
R2031 GNDA.n1790 GNDA.n1789 76.3222
R2032 GNDA.n591 GNDA.n590 76.3222
R2033 GNDA.n552 GNDA.n548 76.3222
R2034 GNDA.n583 GNDA.n549 76.3222
R2035 GNDA.n579 GNDA.n550 76.3222
R2036 GNDA.n575 GNDA.n551 76.3222
R2037 GNDA.n542 GNDA.n499 76.3222
R2038 GNDA.n538 GNDA.n500 76.3222
R2039 GNDA.n534 GNDA.n501 76.3222
R2040 GNDA.n530 GNDA.n502 76.3222
R2041 GNDA.n649 GNDA.n648 76.3222
R2042 GNDA.n653 GNDA.n496 76.3222
R2043 GNDA.n771 GNDA.n373 76.3222
R2044 GNDA.n459 GNDA.n458 76.3222
R2045 GNDA.n762 GNDA.n457 76.3222
R2046 GNDA.n688 GNDA.n456 76.3222
R2047 GNDA.n692 GNDA.n455 76.3222
R2048 GNDA.n701 GNDA.n454 76.3222
R2049 GNDA.n1569 GNDA.n1568 76.3222
R2050 GNDA.n1572 GNDA.n1571 76.3222
R2051 GNDA.n1579 GNDA.n1578 76.3222
R2052 GNDA.n1582 GNDA.n1581 76.3222
R2053 GNDA.n1589 GNDA.n1588 76.3222
R2054 GNDA.n1592 GNDA.n1591 76.3222
R2055 GNDA.n1566 GNDA.n1565 76.3222
R2056 GNDA.n1561 GNDA.n1503 76.3222
R2057 GNDA.n1559 GNDA.n1558 76.3222
R2058 GNDA.n1554 GNDA.n1506 76.3222
R2059 GNDA.n1552 GNDA.n1551 76.3222
R2060 GNDA.n1547 GNDA.n1509 76.3222
R2061 GNDA.n1841 GNDA.n1840 76.3222
R2062 GNDA.n1854 GNDA.n1853 76.3222
R2063 GNDA.n1857 GNDA.n1856 76.3222
R2064 GNDA.n1869 GNDA.n1868 76.3222
R2065 GNDA.n1872 GNDA.n1871 76.3222
R2066 GNDA.n1884 GNDA.n1883 76.3222
R2067 GNDA.n570 GNDA.n569 76.3222
R2068 GNDA.n567 GNDA.n560 76.3222
R2069 GNDA.n566 GNDA.n558 76.3222
R2070 GNDA.n565 GNDA.n556 76.3222
R2071 GNDA.n564 GNDA.n554 76.3222
R2072 GNDA.n563 GNDA.n562 76.3222
R2073 GNDA.n590 GNDA.n547 76.3222
R2074 GNDA.n584 GNDA.n548 76.3222
R2075 GNDA.n580 GNDA.n549 76.3222
R2076 GNDA.n576 GNDA.n550 76.3222
R2077 GNDA.n572 GNDA.n551 76.3222
R2078 GNDA.n1595 GNDA.n384 76.3222
R2079 GNDA.n1492 GNDA.n383 76.3222
R2080 GNDA.n1585 GNDA.n382 76.3222
R2081 GNDA.n1496 GNDA.n381 76.3222
R2082 GNDA.n1575 GNDA.n380 76.3222
R2083 GNDA.n1710 GNDA.n379 76.3222
R2084 GNDA.n1570 GNDA.n1569 76.3222
R2085 GNDA.n1571 GNDA.n1498 76.3222
R2086 GNDA.n1580 GNDA.n1579 76.3222
R2087 GNDA.n1581 GNDA.n1494 76.3222
R2088 GNDA.n1590 GNDA.n1589 76.3222
R2089 GNDA.n1593 GNDA.n1592 76.3222
R2090 GNDA.n1678 GNDA.n1677 76.3222
R2091 GNDA.n1321 GNDA.n395 76.3222
R2092 GNDA.n1320 GNDA.n1319 76.3222
R2093 GNDA.n1317 GNDA.n1316 76.3222
R2094 GNDA.n1312 GNDA.n1311 76.3222
R2095 GNDA.n1309 GNDA.n1308 76.3222
R2096 GNDA.n1339 GNDA.n1338 76.3222
R2097 GNDA.n1334 GNDA.n1307 76.3222
R2098 GNDA.n1332 GNDA.n1331 76.3222
R2099 GNDA.n1327 GNDA.n1326 76.3222
R2100 GNDA.n1324 GNDA.n397 76.3222
R2101 GNDA.n1673 GNDA.n1672 76.3222
R2102 GNDA.n365 GNDA.n364 76.3222
R2103 GNDA.n362 GNDA.n355 76.3222
R2104 GNDA.n361 GNDA.n353 76.3222
R2105 GNDA.n360 GNDA.n351 76.3222
R2106 GNDA.n359 GNDA.n349 76.3222
R2107 GNDA.n358 GNDA.n357 76.3222
R2108 GNDA.n1740 GNDA.n341 76.3222
R2109 GNDA.n1738 GNDA.n347 76.3222
R2110 GNDA.n1731 GNDA.n346 76.3222
R2111 GNDA.n1727 GNDA.n345 76.3222
R2112 GNDA.n1723 GNDA.n344 76.3222
R2113 GNDA.n1719 GNDA.n343 76.3222
R2114 GNDA.n646 GNDA.n644 76.3222
R2115 GNDA.n640 GNDA.n601 76.3222
R2116 GNDA.n636 GNDA.n600 76.3222
R2117 GNDA.n632 GNDA.n599 76.3222
R2118 GNDA.n628 GNDA.n598 76.3222
R2119 GNDA.n624 GNDA.n597 76.3222
R2120 GNDA.n596 GNDA.n508 76.3222
R2121 GNDA.n524 GNDA.n507 76.3222
R2122 GNDA.n520 GNDA.n506 76.3222
R2123 GNDA.n516 GNDA.n505 76.3222
R2124 GNDA.n512 GNDA.n504 76.3222
R2125 GNDA.n503 GNDA.n340 76.3222
R2126 GNDA.n650 GNDA.n496 76.3222
R2127 GNDA.n648 GNDA.n498 76.3222
R2128 GNDA.n533 GNDA.n502 76.3222
R2129 GNDA.n537 GNDA.n501 76.3222
R2130 GNDA.n541 GNDA.n500 76.3222
R2131 GNDA.n546 GNDA.n499 76.3222
R2132 GNDA.n1238 GNDA.n1237 76.3222
R2133 GNDA.n1230 GNDA.n1229 76.3222
R2134 GNDA.n1150 GNDA.n1126 76.3222
R2135 GNDA.n1151 GNDA.n1148 76.3222
R2136 GNDA.n1164 GNDA.n1163 76.3222
R2137 GNDA.n1166 GNDA.n1165 76.3222
R2138 GNDA.n1746 GNDA.n271 76.3222
R2139 GNDA.n1761 GNDA.n1760 76.3222
R2140 GNDA.n1762 GNDA.n266 76.3222
R2141 GNDA.n1776 GNDA.n1775 76.3222
R2142 GNDA.n1777 GNDA.n259 76.3222
R2143 GNDA.n1791 GNDA.n1790 76.3222
R2144 GNDA.n1840 GNDA.n189 76.3222
R2145 GNDA.n1855 GNDA.n1854 76.3222
R2146 GNDA.n1856 GNDA.n184 76.3222
R2147 GNDA.n1870 GNDA.n1869 76.3222
R2148 GNDA.n1871 GNDA.n177 76.3222
R2149 GNDA.n1885 GNDA.n1884 76.3222
R2150 GNDA.n1346 GNDA.n1345 76.3222
R2151 GNDA.n1278 GNDA.n1276 76.3222
R2152 GNDA.n1353 GNDA.n1352 76.3222
R2153 GNDA.n1275 GNDA.n1273 76.3222
R2154 GNDA.n1360 GNDA.n1359 76.3222
R2155 GNDA.n1272 GNDA.n1270 76.3222
R2156 GNDA.n1288 GNDA.n378 76.3222
R2157 GNDA.n1292 GNDA.n1291 76.3222
R2158 GNDA.n1287 GNDA.n1285 76.3222
R2159 GNDA.n1299 GNDA.n1298 76.3222
R2160 GNDA.n1284 GNDA.n1282 76.3222
R2161 GNDA.n1306 GNDA.n1305 76.3222
R2162 GNDA.n1509 GNDA.n1507 76.3222
R2163 GNDA.n1553 GNDA.n1552 76.3222
R2164 GNDA.n1506 GNDA.n1504 76.3222
R2165 GNDA.n1560 GNDA.n1559 76.3222
R2166 GNDA.n1503 GNDA.n1501 76.3222
R2167 GNDA.n1567 GNDA.n1566 76.3222
R2168 GNDA.n1008 GNDA.n1007 76.3222
R2169 GNDA.n1005 GNDA.n1004 76.3222
R2170 GNDA.n926 GNDA.n896 76.3222
R2171 GNDA.n930 GNDA.n895 76.3222
R2172 GNDA.n940 GNDA.n894 76.3222
R2173 GNDA.n943 GNDA.n893 76.3222
R2174 GNDA.n892 GNDA.n891 76.3222
R2175 GNDA.n884 GNDA.n776 76.3222
R2176 GNDA.n808 GNDA.n775 76.3222
R2177 GNDA.n814 GNDA.n774 76.3222
R2178 GNDA.n821 GNDA.n773 76.3222
R2179 GNDA.n803 GNDA.n772 76.3222
R2180 GNDA.n771 GNDA.n770 76.3222
R2181 GNDA.n763 GNDA.n458 76.3222
R2182 GNDA.n687 GNDA.n457 76.3222
R2183 GNDA.n693 GNDA.n456 76.3222
R2184 GNDA.n700 GNDA.n455 76.3222
R2185 GNDA.n682 GNDA.n454 76.3222
R2186 GNDA.n1367 GNDA.n1366 76.3222
R2187 GNDA.n1368 GNDA.n1268 76.3222
R2188 GNDA.n1375 GNDA.n1374 76.3222
R2189 GNDA.n1376 GNDA.n1266 76.3222
R2190 GNDA.n1383 GNDA.n1382 76.3222
R2191 GNDA.n620 GNDA.n443 76.3222
R2192 GNDA.n616 GNDA.n444 76.3222
R2193 GNDA.n612 GNDA.n445 76.3222
R2194 GNDA.n608 GNDA.n446 76.3222
R2195 GNDA.n604 GNDA.n447 76.3222
R2196 GNDA.n1263 GNDA.n1017 76.3222
R2197 GNDA.n1255 GNDA.n438 76.3222
R2198 GNDA.n1251 GNDA.n439 76.3222
R2199 GNDA.n1247 GNDA.n440 76.3222
R2200 GNDA.n1243 GNDA.n441 76.3222
R2201 GNDA.n1190 GNDA.n1134 74.5978
R2202 GNDA.n1187 GNDA.n1134 74.5978
R2203 GNDA.n963 GNDA.n962 74.5978
R2204 GNDA.n962 GNDA.n961 74.5978
R2205 GNDA.n1405 GNDA.n411 74.5978
R2206 GNDA.n1402 GNDA.n411 74.5978
R2207 GNDA.n1633 GNDA.n64 74.5978
R2208 GNDA.n1630 GNDA.n64 74.5978
R2209 GNDA.n845 GNDA.n791 74.5978
R2210 GNDA.n842 GNDA.n791 74.5978
R2211 GNDA.n298 GNDA.n281 74.5978
R2212 GNDA.n299 GNDA.n298 74.5978
R2213 GNDA.n724 GNDA.n473 74.5978
R2214 GNDA.n721 GNDA.n473 74.5978
R2215 GNDA.n1990 GNDA.n100 74.5978
R2216 GNDA.n1987 GNDA.n100 74.5978
R2217 GNDA.n216 GNDA.n199 74.5978
R2218 GNDA.n217 GNDA.n216 74.5978
R2219 GNDA.t177 GNDA.n1608 74.1404
R2220 GNDA.t7 GNDA.t148 72.9499
R2221 GNDA.n2072 GNDA.t173 70.0216
R2222 GNDA.n121 GNDA.t149 69.4695
R2223 GNDA.n1234 GNDA.n1123 69.3109
R2224 GNDA.n1209 GNDA.n1123 69.3109
R2225 GNDA.n998 GNDA.n997 69.3109
R2226 GNDA.n997 GNDA.n996 69.3109
R2227 GNDA.n1471 GNDA.n1470 69.3109
R2228 GNDA.n1471 GNDA.n423 69.3109
R2229 GNDA.n2077 GNDA.n2076 69.3109
R2230 GNDA.n2077 GNDA.n75 69.3109
R2231 GNDA.n888 GNDA.n781 69.3109
R2232 GNDA.n864 GNDA.n781 69.3109
R2233 GNDA.n1754 GNDA.n1753 69.3109
R2234 GNDA.n1753 GNDA.n1752 69.3109
R2235 GNDA.n767 GNDA.n463 69.3109
R2236 GNDA.n743 GNDA.n463 69.3109
R2237 GNDA.n2046 GNDA.n2045 69.3109
R2238 GNDA.n2046 GNDA.n111 69.3109
R2239 GNDA.n1848 GNDA.n1847 69.3109
R2240 GNDA.n1847 GNDA.n1846 69.3109
R2241 GNDA.t214 GNDA.n1223 65.8183
R2242 GNDA.t214 GNDA.n1143 65.8183
R2243 GNDA.t214 GNDA.n1142 65.8183
R2244 GNDA.t214 GNDA.n1141 65.8183
R2245 GNDA.t214 GNDA.n1132 65.8183
R2246 GNDA.t214 GNDA.n1139 65.8183
R2247 GNDA.t214 GNDA.n1130 65.8183
R2248 GNDA.t214 GNDA.n1140 65.8183
R2249 GNDA.t214 GNDA.n1138 65.8183
R2250 GNDA.t214 GNDA.n1137 65.8183
R2251 GNDA.t214 GNDA.n1136 65.8183
R2252 GNDA.t214 GNDA.n1135 65.8183
R2253 GNDA.t214 GNDA.n1133 65.8183
R2254 GNDA.t214 GNDA.n1131 65.8183
R2255 GNDA.n1224 GNDA.t214 65.8183
R2256 GNDA.t214 GNDA.n1124 65.8183
R2257 GNDA.n980 GNDA.t242 65.8183
R2258 GNDA.n986 GNDA.t242 65.8183
R2259 GNDA.n988 GNDA.t242 65.8183
R2260 GNDA.n994 GNDA.t242 65.8183
R2261 GNDA.n964 GNDA.t242 65.8183
R2262 GNDA.n970 GNDA.t242 65.8183
R2263 GNDA.n972 GNDA.t242 65.8183
R2264 GNDA.n978 GNDA.t242 65.8183
R2265 GNDA.n948 GNDA.t242 65.8183
R2266 GNDA.n916 GNDA.t242 65.8183
R2267 GNDA.n955 GNDA.t242 65.8183
R2268 GNDA.n913 GNDA.t242 65.8183
R2269 GNDA.n936 GNDA.t242 65.8183
R2270 GNDA.n934 GNDA.t242 65.8183
R2271 GNDA.n921 GNDA.t242 65.8183
R2272 GNDA.n1000 GNDA.t242 65.8183
R2273 GNDA.t243 GNDA.n422 65.8183
R2274 GNDA.t243 GNDA.n421 65.8183
R2275 GNDA.t243 GNDA.n420 65.8183
R2276 GNDA.t243 GNDA.n419 65.8183
R2277 GNDA.t243 GNDA.n410 65.8183
R2278 GNDA.t243 GNDA.n417 65.8183
R2279 GNDA.t243 GNDA.n407 65.8183
R2280 GNDA.t243 GNDA.n418 65.8183
R2281 GNDA.t243 GNDA.n416 65.8183
R2282 GNDA.t243 GNDA.n414 65.8183
R2283 GNDA.t243 GNDA.n413 65.8183
R2284 GNDA.t243 GNDA.n412 65.8183
R2285 GNDA.n1472 GNDA.t243 65.8183
R2286 GNDA.t243 GNDA.n409 65.8183
R2287 GNDA.t243 GNDA.n408 65.8183
R2288 GNDA.t243 GNDA.n406 65.8183
R2289 GNDA.t216 GNDA.n74 65.8183
R2290 GNDA.t216 GNDA.n73 65.8183
R2291 GNDA.t216 GNDA.n72 65.8183
R2292 GNDA.t216 GNDA.n71 65.8183
R2293 GNDA.t216 GNDA.n62 65.8183
R2294 GNDA.t216 GNDA.n69 65.8183
R2295 GNDA.t216 GNDA.n60 65.8183
R2296 GNDA.t216 GNDA.n70 65.8183
R2297 GNDA.t216 GNDA.n68 65.8183
R2298 GNDA.t216 GNDA.n67 65.8183
R2299 GNDA.t216 GNDA.n66 65.8183
R2300 GNDA.t216 GNDA.n65 65.8183
R2301 GNDA.t216 GNDA.n63 65.8183
R2302 GNDA.n2078 GNDA.t216 65.8183
R2303 GNDA.t216 GNDA.n61 65.8183
R2304 GNDA.t216 GNDA.n59 65.8183
R2305 GNDA.t215 GNDA.n878 65.8183
R2306 GNDA.t215 GNDA.n800 65.8183
R2307 GNDA.t215 GNDA.n799 65.8183
R2308 GNDA.t215 GNDA.n798 65.8183
R2309 GNDA.t215 GNDA.n789 65.8183
R2310 GNDA.t215 GNDA.n796 65.8183
R2311 GNDA.t215 GNDA.n787 65.8183
R2312 GNDA.t215 GNDA.n797 65.8183
R2313 GNDA.t215 GNDA.n795 65.8183
R2314 GNDA.t215 GNDA.n794 65.8183
R2315 GNDA.t215 GNDA.n793 65.8183
R2316 GNDA.t215 GNDA.n792 65.8183
R2317 GNDA.t215 GNDA.n790 65.8183
R2318 GNDA.t215 GNDA.n788 65.8183
R2319 GNDA.n879 GNDA.t215 65.8183
R2320 GNDA.t215 GNDA.n782 65.8183
R2321 GNDA.n320 GNDA.t198 65.8183
R2322 GNDA.n322 GNDA.t198 65.8183
R2323 GNDA.n328 GNDA.t198 65.8183
R2324 GNDA.n330 GNDA.t198 65.8183
R2325 GNDA.n304 GNDA.t198 65.8183
R2326 GNDA.n306 GNDA.t198 65.8183
R2327 GNDA.n312 GNDA.t198 65.8183
R2328 GNDA.n314 GNDA.t198 65.8183
R2329 GNDA.t198 GNDA.n262 65.8183
R2330 GNDA.n289 GNDA.t198 65.8183
R2331 GNDA.n285 GNDA.t198 65.8183
R2332 GNDA.n296 GNDA.t198 65.8183
R2333 GNDA.n1783 GNDA.t198 65.8183
R2334 GNDA.n1770 GNDA.t198 65.8183
R2335 GNDA.n1768 GNDA.t198 65.8183
R2336 GNDA.n1755 GNDA.t198 65.8183
R2337 GNDA.t250 GNDA.n757 65.8183
R2338 GNDA.t250 GNDA.n482 65.8183
R2339 GNDA.t250 GNDA.n481 65.8183
R2340 GNDA.t250 GNDA.n480 65.8183
R2341 GNDA.t250 GNDA.n471 65.8183
R2342 GNDA.t250 GNDA.n478 65.8183
R2343 GNDA.t250 GNDA.n469 65.8183
R2344 GNDA.t250 GNDA.n479 65.8183
R2345 GNDA.t250 GNDA.n477 65.8183
R2346 GNDA.t250 GNDA.n476 65.8183
R2347 GNDA.t250 GNDA.n475 65.8183
R2348 GNDA.t250 GNDA.n474 65.8183
R2349 GNDA.t250 GNDA.n472 65.8183
R2350 GNDA.t250 GNDA.n470 65.8183
R2351 GNDA.n758 GNDA.t250 65.8183
R2352 GNDA.t250 GNDA.n464 65.8183
R2353 GNDA.t196 GNDA.n110 65.8183
R2354 GNDA.t196 GNDA.n109 65.8183
R2355 GNDA.t196 GNDA.n108 65.8183
R2356 GNDA.t196 GNDA.n107 65.8183
R2357 GNDA.t196 GNDA.n98 65.8183
R2358 GNDA.t196 GNDA.n105 65.8183
R2359 GNDA.t196 GNDA.n96 65.8183
R2360 GNDA.t196 GNDA.n106 65.8183
R2361 GNDA.t196 GNDA.n104 65.8183
R2362 GNDA.t196 GNDA.n103 65.8183
R2363 GNDA.t196 GNDA.n102 65.8183
R2364 GNDA.t196 GNDA.n101 65.8183
R2365 GNDA.t196 GNDA.n99 65.8183
R2366 GNDA.n2047 GNDA.t196 65.8183
R2367 GNDA.t196 GNDA.n97 65.8183
R2368 GNDA.t196 GNDA.n95 65.8183
R2369 GNDA.n238 GNDA.t222 65.8183
R2370 GNDA.n240 GNDA.t222 65.8183
R2371 GNDA.n246 GNDA.t222 65.8183
R2372 GNDA.n248 GNDA.t222 65.8183
R2373 GNDA.n222 GNDA.t222 65.8183
R2374 GNDA.n224 GNDA.t222 65.8183
R2375 GNDA.n230 GNDA.t222 65.8183
R2376 GNDA.n232 GNDA.t222 65.8183
R2377 GNDA.t222 GNDA.n180 65.8183
R2378 GNDA.n207 GNDA.t222 65.8183
R2379 GNDA.n203 GNDA.t222 65.8183
R2380 GNDA.n214 GNDA.t222 65.8183
R2381 GNDA.n1877 GNDA.t222 65.8183
R2382 GNDA.n1864 GNDA.t222 65.8183
R2383 GNDA.n1862 GNDA.t222 65.8183
R2384 GNDA.n1849 GNDA.t222 65.8183
R2385 GNDA.t218 GNDA.t0 65.7614
R2386 GNDA.t51 GNDA.t309 65.7614
R2387 GNDA.t309 GNDA.t77 65.7614
R2388 GNDA.t11 GNDA.t2 65.7614
R2389 GNDA.t15 GNDA.t11 65.7614
R2390 GNDA.t73 GNDA.t27 65.7614
R2391 GNDA.t27 GNDA.t38 65.7614
R2392 GNDA.t38 GNDA.t39 65.7614
R2393 GNDA.t201 GNDA.t8 65.7614
R2394 GNDA.t121 GNDA.t298 65.271
R2395 GNDA.t104 GNDA.t54 65.271
R2396 GNDA.n2145 GNDA.t138 65.271
R2397 GNDA.n2174 GNDA.t61 65.271
R2398 GNDA.t42 GNDA.t18 65.271
R2399 GNDA.t28 GNDA.t45 65.271
R2400 GNDA.n486 GNDA.t199 65.0078
R2401 GNDA.n1466 GNDA.t167 63.8432
R2402 GNDA.n2071 GNDA.t189 63.8432
R2403 GNDA.n2039 GNDA.t183 63.8432
R2404 GNDA.t126 GNDA.t133 62.9326
R2405 GNDA.t21 GNDA.t64 62.9326
R2406 GNDA.t88 GNDA.t21 62.9326
R2407 GNDA.n2139 GNDA.t219 62.2505
R2408 GNDA.n2151 GNDA.t229 62.2505
R2409 GNDA.n2187 GNDA.t271 62.2505
R2410 GNDA.n2191 GNDA.t280 62.2505
R2411 GNDA.n2161 GNDA.t221 62.2505
R2412 GNDA.n2164 GNDA.t237 62.2505
R2413 GNDA.n2144 GNDA.t239 62.2505
R2414 GNDA.n2175 GNDA.t278 62.2505
R2415 GNDA.n2183 GNDA.t276 62.2505
R2416 GNDA.n2179 GNDA.t202 62.2505
R2417 GNDA.n26 GNDA.t261 62.2505
R2418 GNDA.n2219 GNDA.t268 62.2505
R2419 GNDA.n2210 GNDA.n2209 61.4316
R2420 GNDA.t102 GNDA.n2156 59.7836
R2421 GNDA.t20 GNDA.n2155 59.7836
R2422 GNDA.t34 GNDA.n2154 59.7836
R2423 GNDA.t118 GNDA.n2153 59.7836
R2424 GNDA.n2216 GNDA.t55 59.7836
R2425 GNDA.n2215 GNDA.t6 59.7836
R2426 GNDA.n2185 GNDA.t49 59.7836
R2427 GNDA.n2217 GNDA.t76 59.7836
R2428 GNDA.t43 GNDA.n2157 59.7836
R2429 GNDA.t169 GNDA.n1449 59.7243
R2430 GNDA.n1607 GNDA.t191 59.7243
R2431 GNDA.n135 GNDA.t181 59.7243
R2432 GNDA.n2193 GNDA.n8 59.2425
R2433 GNDA.n2202 GNDA.n2201 59.2425
R2434 GNDA.n2108 GNDA.n2107 59.2425
R2435 GNDA.n2099 GNDA.n2098 59.2425
R2436 GNDA.t24 GNDA.n1442 58.6946
R2437 GNDA.n1464 GNDA.t95 58.6946
R2438 GNDA.t131 GNDA.n1477 58.6946
R2439 GNDA.t214 GNDA.n1123 57.8461
R2440 GNDA.n997 GNDA.t242 57.8461
R2441 GNDA.t243 GNDA.n1471 57.8461
R2442 GNDA.t216 GNDA.n2077 57.8461
R2443 GNDA.t215 GNDA.n781 57.8461
R2444 GNDA.n1753 GNDA.t198 57.8461
R2445 GNDA.t250 GNDA.n463 57.8461
R2446 GNDA.t196 GNDA.n2046 57.8461
R2447 GNDA.n1847 GNDA.t222 57.8461
R2448 GNDA.n2098 GNDA.t255 57.5921
R2449 GNDA.n2108 GNDA.t265 57.5921
R2450 GNDA.n2152 GNDA.t138 57.5921
R2451 GNDA.n2186 GNDA.t61 57.5921
R2452 GNDA.n2218 GNDA.t304 57.5921
R2453 GNDA.n2202 GNDA.t282 57.5921
R2454 GNDA.t209 GNDA.n8 57.5921
R2455 GNDA.t300 GNDA.t157 56.6352
R2456 GNDA.n2058 GNDA.t273 56.6352
R2457 GNDA.t74 GNDA.t153 56.6352
R2458 GNDA.n1242 GNDA.n442 56.3995
R2459 GNDA.n1240 GNDA.n442 56.3995
R2460 GNDA.n680 GNDA.n679 56.3995
R2461 GNDA.n1524 GNDA.n1520 56.3995
R2462 GNDA.n1524 GNDA.n1523 56.3995
R2463 GNDA.n681 GNDA.n680 56.3995
R2464 GNDA.n1886 GNDA.n174 56.3995
R2465 GNDA.n1887 GNDA.n1886 56.3995
R2466 GNDA.n1386 GNDA.n436 56.3995
R2467 GNDA.n1014 GNDA.n1013 56.3995
R2468 GNDA.n1681 GNDA.n1680 55.6055
R2469 GNDA.t214 GNDA.n1134 55.2026
R2470 GNDA.n962 GNDA.t242 55.2026
R2471 GNDA.t243 GNDA.n411 55.2026
R2472 GNDA.t216 GNDA.n64 55.2026
R2473 GNDA.t215 GNDA.n791 55.2026
R2474 GNDA.n298 GNDA.t198 55.2026
R2475 GNDA.t250 GNDA.n473 55.2026
R2476 GNDA.t196 GNDA.n100 55.2026
R2477 GNDA.n216 GNDA.t222 55.2026
R2478 GNDA.n1599 GNDA.n81 54.5757
R2479 GNDA.n1690 GNDA.n1689 54.5757
R2480 GNDA.t79 GNDA.n2040 54.5757
R2481 GNDA.n128 GNDA.t50 54.5757
R2482 GNDA.t30 GNDA.n1965 54.5757
R2483 GNDA.t175 GNDA.n1607 53.546
R2484 GNDA.n1205 GNDA.n1140 53.3664
R2485 GNDA.n1202 GNDA.n1130 53.3664
R2486 GNDA.n1198 GNDA.n1139 53.3664
R2487 GNDA.n1194 GNDA.n1132 53.3664
R2488 GNDA.n1183 GNDA.n1135 53.3664
R2489 GNDA.n1179 GNDA.n1136 53.3664
R2490 GNDA.n1175 GNDA.n1137 53.3664
R2491 GNDA.n1171 GNDA.n1138 53.3664
R2492 GNDA.n1233 GNDA.n1124 53.3664
R2493 GNDA.n1225 GNDA.n1224 53.3664
R2494 GNDA.n1154 GNDA.n1131 53.3664
R2495 GNDA.n1159 GNDA.n1133 53.3664
R2496 GNDA.n1223 GNDA.n1222 53.3664
R2497 GNDA.n1145 GNDA.n1143 53.3664
R2498 GNDA.n1217 GNDA.n1142 53.3664
R2499 GNDA.n1213 GNDA.n1141 53.3664
R2500 GNDA.n1223 GNDA.n1144 53.3664
R2501 GNDA.n1218 GNDA.n1143 53.3664
R2502 GNDA.n1214 GNDA.n1142 53.3664
R2503 GNDA.n1210 GNDA.n1141 53.3664
R2504 GNDA.n1191 GNDA.n1132 53.3664
R2505 GNDA.n1195 GNDA.n1139 53.3664
R2506 GNDA.n1199 GNDA.n1130 53.3664
R2507 GNDA.n1203 GNDA.n1140 53.3664
R2508 GNDA.n1174 GNDA.n1138 53.3664
R2509 GNDA.n1178 GNDA.n1137 53.3664
R2510 GNDA.n1182 GNDA.n1136 53.3664
R2511 GNDA.n1186 GNDA.n1135 53.3664
R2512 GNDA.n1170 GNDA.n1133 53.3664
R2513 GNDA.n1158 GNDA.n1131 53.3664
R2514 GNDA.n1224 GNDA.n1129 53.3664
R2515 GNDA.n1128 GNDA.n1124 53.3664
R2516 GNDA.n979 GNDA.n978 53.3664
R2517 GNDA.n972 GNDA.n907 53.3664
R2518 GNDA.n971 GNDA.n970 53.3664
R2519 GNDA.n964 GNDA.n909 53.3664
R2520 GNDA.n957 GNDA.n913 53.3664
R2521 GNDA.n955 GNDA.n954 53.3664
R2522 GNDA.n950 GNDA.n916 53.3664
R2523 GNDA.n948 GNDA.n947 53.3664
R2524 GNDA.n1000 GNDA.n999 53.3664
R2525 GNDA.n921 GNDA.n901 53.3664
R2526 GNDA.n934 GNDA.n933 53.3664
R2527 GNDA.n937 GNDA.n936 53.3664
R2528 GNDA.n980 GNDA.n905 53.3664
R2529 GNDA.n986 GNDA.n985 53.3664
R2530 GNDA.n989 GNDA.n988 53.3664
R2531 GNDA.n994 GNDA.n993 53.3664
R2532 GNDA.n981 GNDA.n980 53.3664
R2533 GNDA.n987 GNDA.n986 53.3664
R2534 GNDA.n988 GNDA.n903 53.3664
R2535 GNDA.n995 GNDA.n994 53.3664
R2536 GNDA.n965 GNDA.n964 53.3664
R2537 GNDA.n970 GNDA.n969 53.3664
R2538 GNDA.n973 GNDA.n972 53.3664
R2539 GNDA.n978 GNDA.n977 53.3664
R2540 GNDA.n949 GNDA.n948 53.3664
R2541 GNDA.n916 GNDA.n914 53.3664
R2542 GNDA.n956 GNDA.n955 53.3664
R2543 GNDA.n913 GNDA.n911 53.3664
R2544 GNDA.n936 GNDA.n917 53.3664
R2545 GNDA.n935 GNDA.n934 53.3664
R2546 GNDA.n922 GNDA.n921 53.3664
R2547 GNDA.n1001 GNDA.n1000 53.3664
R2548 GNDA.n1421 GNDA.n418 53.3664
R2549 GNDA.n1417 GNDA.n407 53.3664
R2550 GNDA.n1413 GNDA.n417 53.3664
R2551 GNDA.n1409 GNDA.n410 53.3664
R2552 GNDA.n1398 GNDA.n412 53.3664
R2553 GNDA.n1394 GNDA.n413 53.3664
R2554 GNDA.n1390 GNDA.n414 53.3664
R2555 GNDA.n416 GNDA.n415 53.3664
R2556 GNDA.n424 GNDA.n406 53.3664
R2557 GNDA.n1460 GNDA.n408 53.3664
R2558 GNDA.n1455 GNDA.n409 53.3664
R2559 GNDA.n1473 GNDA.n1472 53.3664
R2560 GNDA.n1425 GNDA.n422 53.3664
R2561 GNDA.n1426 GNDA.n421 53.3664
R2562 GNDA.n1430 GNDA.n420 53.3664
R2563 GNDA.n1434 GNDA.n419 53.3664
R2564 GNDA.n1422 GNDA.n422 53.3664
R2565 GNDA.n1429 GNDA.n421 53.3664
R2566 GNDA.n1433 GNDA.n420 53.3664
R2567 GNDA.n1436 GNDA.n419 53.3664
R2568 GNDA.n1406 GNDA.n410 53.3664
R2569 GNDA.n1410 GNDA.n417 53.3664
R2570 GNDA.n1414 GNDA.n407 53.3664
R2571 GNDA.n1418 GNDA.n418 53.3664
R2572 GNDA.n1389 GNDA.n416 53.3664
R2573 GNDA.n1393 GNDA.n414 53.3664
R2574 GNDA.n1397 GNDA.n413 53.3664
R2575 GNDA.n1401 GNDA.n412 53.3664
R2576 GNDA.n1472 GNDA.n405 53.3664
R2577 GNDA.n409 GNDA.n404 53.3664
R2578 GNDA.n1456 GNDA.n408 53.3664
R2579 GNDA.n1459 GNDA.n406 53.3664
R2580 GNDA.n1649 GNDA.n70 53.3664
R2581 GNDA.n1645 GNDA.n60 53.3664
R2582 GNDA.n1641 GNDA.n69 53.3664
R2583 GNDA.n1637 GNDA.n62 53.3664
R2584 GNDA.n1626 GNDA.n65 53.3664
R2585 GNDA.n1622 GNDA.n66 53.3664
R2586 GNDA.n1618 GNDA.n67 53.3664
R2587 GNDA.n1614 GNDA.n68 53.3664
R2588 GNDA.n76 GNDA.n59 53.3664
R2589 GNDA.n2066 GNDA.n61 53.3664
R2590 GNDA.n2079 GNDA.n2078 53.3664
R2591 GNDA.n1603 GNDA.n63 53.3664
R2592 GNDA.n1653 GNDA.n74 53.3664
R2593 GNDA.n1654 GNDA.n73 53.3664
R2594 GNDA.n1658 GNDA.n72 53.3664
R2595 GNDA.n1662 GNDA.n71 53.3664
R2596 GNDA.n1650 GNDA.n74 53.3664
R2597 GNDA.n1657 GNDA.n73 53.3664
R2598 GNDA.n1661 GNDA.n72 53.3664
R2599 GNDA.n1664 GNDA.n71 53.3664
R2600 GNDA.n1634 GNDA.n62 53.3664
R2601 GNDA.n1638 GNDA.n69 53.3664
R2602 GNDA.n1642 GNDA.n60 53.3664
R2603 GNDA.n1646 GNDA.n70 53.3664
R2604 GNDA.n1617 GNDA.n68 53.3664
R2605 GNDA.n1621 GNDA.n67 53.3664
R2606 GNDA.n1625 GNDA.n66 53.3664
R2607 GNDA.n1629 GNDA.n65 53.3664
R2608 GNDA.n1613 GNDA.n63 53.3664
R2609 GNDA.n2078 GNDA.n58 53.3664
R2610 GNDA.n61 GNDA.n57 53.3664
R2611 GNDA.n2065 GNDA.n59 53.3664
R2612 GNDA.n860 GNDA.n797 53.3664
R2613 GNDA.n857 GNDA.n787 53.3664
R2614 GNDA.n853 GNDA.n796 53.3664
R2615 GNDA.n849 GNDA.n789 53.3664
R2616 GNDA.n838 GNDA.n792 53.3664
R2617 GNDA.n834 GNDA.n793 53.3664
R2618 GNDA.n830 GNDA.n794 53.3664
R2619 GNDA.n826 GNDA.n795 53.3664
R2620 GNDA.n887 GNDA.n782 53.3664
R2621 GNDA.n880 GNDA.n879 53.3664
R2622 GNDA.n811 GNDA.n788 53.3664
R2623 GNDA.n818 GNDA.n790 53.3664
R2624 GNDA.n878 GNDA.n877 53.3664
R2625 GNDA.n802 GNDA.n800 53.3664
R2626 GNDA.n872 GNDA.n799 53.3664
R2627 GNDA.n868 GNDA.n798 53.3664
R2628 GNDA.n878 GNDA.n801 53.3664
R2629 GNDA.n873 GNDA.n800 53.3664
R2630 GNDA.n869 GNDA.n799 53.3664
R2631 GNDA.n865 GNDA.n798 53.3664
R2632 GNDA.n846 GNDA.n789 53.3664
R2633 GNDA.n850 GNDA.n796 53.3664
R2634 GNDA.n854 GNDA.n787 53.3664
R2635 GNDA.n858 GNDA.n797 53.3664
R2636 GNDA.n829 GNDA.n795 53.3664
R2637 GNDA.n833 GNDA.n794 53.3664
R2638 GNDA.n837 GNDA.n793 53.3664
R2639 GNDA.n841 GNDA.n792 53.3664
R2640 GNDA.n825 GNDA.n790 53.3664
R2641 GNDA.n817 GNDA.n788 53.3664
R2642 GNDA.n879 GNDA.n786 53.3664
R2643 GNDA.n785 GNDA.n782 53.3664
R2644 GNDA.n314 GNDA.n277 53.3664
R2645 GNDA.n313 GNDA.n312 53.3664
R2646 GNDA.n306 GNDA.n279 53.3664
R2647 GNDA.n305 GNDA.n304 53.3664
R2648 GNDA.n296 GNDA.n295 53.3664
R2649 GNDA.n291 GNDA.n285 53.3664
R2650 GNDA.n289 GNDA.n288 53.3664
R2651 GNDA.n1785 GNDA.n262 53.3664
R2652 GNDA.n1756 GNDA.n1755 53.3664
R2653 GNDA.n1768 GNDA.n1767 53.3664
R2654 GNDA.n1771 GNDA.n1770 53.3664
R2655 GNDA.n1783 GNDA.n1782 53.3664
R2656 GNDA.n321 GNDA.n320 53.3664
R2657 GNDA.n323 GNDA.n322 53.3664
R2658 GNDA.n328 GNDA.n327 53.3664
R2659 GNDA.n331 GNDA.n330 53.3664
R2660 GNDA.n320 GNDA.n319 53.3664
R2661 GNDA.n322 GNDA.n275 53.3664
R2662 GNDA.n329 GNDA.n328 53.3664
R2663 GNDA.n330 GNDA.n273 53.3664
R2664 GNDA.n304 GNDA.n303 53.3664
R2665 GNDA.n307 GNDA.n306 53.3664
R2666 GNDA.n312 GNDA.n311 53.3664
R2667 GNDA.n315 GNDA.n314 53.3664
R2668 GNDA.n286 GNDA.n262 53.3664
R2669 GNDA.n290 GNDA.n289 53.3664
R2670 GNDA.n285 GNDA.n283 53.3664
R2671 GNDA.n297 GNDA.n296 53.3664
R2672 GNDA.n1784 GNDA.n1783 53.3664
R2673 GNDA.n1770 GNDA.n263 53.3664
R2674 GNDA.n1769 GNDA.n1768 53.3664
R2675 GNDA.n1755 GNDA.n268 53.3664
R2676 GNDA.n739 GNDA.n479 53.3664
R2677 GNDA.n736 GNDA.n469 53.3664
R2678 GNDA.n732 GNDA.n478 53.3664
R2679 GNDA.n728 GNDA.n471 53.3664
R2680 GNDA.n717 GNDA.n474 53.3664
R2681 GNDA.n713 GNDA.n475 53.3664
R2682 GNDA.n709 GNDA.n476 53.3664
R2683 GNDA.n705 GNDA.n477 53.3664
R2684 GNDA.n766 GNDA.n464 53.3664
R2685 GNDA.n759 GNDA.n758 53.3664
R2686 GNDA.n690 GNDA.n470 53.3664
R2687 GNDA.n697 GNDA.n472 53.3664
R2688 GNDA.n757 GNDA.n756 53.3664
R2689 GNDA.n484 GNDA.n482 53.3664
R2690 GNDA.n751 GNDA.n481 53.3664
R2691 GNDA.n747 GNDA.n480 53.3664
R2692 GNDA.n757 GNDA.n483 53.3664
R2693 GNDA.n752 GNDA.n482 53.3664
R2694 GNDA.n748 GNDA.n481 53.3664
R2695 GNDA.n744 GNDA.n480 53.3664
R2696 GNDA.n725 GNDA.n471 53.3664
R2697 GNDA.n729 GNDA.n478 53.3664
R2698 GNDA.n733 GNDA.n469 53.3664
R2699 GNDA.n737 GNDA.n479 53.3664
R2700 GNDA.n708 GNDA.n477 53.3664
R2701 GNDA.n712 GNDA.n476 53.3664
R2702 GNDA.n716 GNDA.n475 53.3664
R2703 GNDA.n720 GNDA.n474 53.3664
R2704 GNDA.n704 GNDA.n472 53.3664
R2705 GNDA.n696 GNDA.n470 53.3664
R2706 GNDA.n758 GNDA.n468 53.3664
R2707 GNDA.n467 GNDA.n464 53.3664
R2708 GNDA.n2006 GNDA.n106 53.3664
R2709 GNDA.n2002 GNDA.n96 53.3664
R2710 GNDA.n1998 GNDA.n105 53.3664
R2711 GNDA.n1994 GNDA.n98 53.3664
R2712 GNDA.n1983 GNDA.n101 53.3664
R2713 GNDA.n1979 GNDA.n102 53.3664
R2714 GNDA.n1975 GNDA.n103 53.3664
R2715 GNDA.n1971 GNDA.n104 53.3664
R2716 GNDA.n112 GNDA.n95 53.3664
R2717 GNDA.n2035 GNDA.n97 53.3664
R2718 GNDA.n2048 GNDA.n2047 53.3664
R2719 GNDA.n130 GNDA.n99 53.3664
R2720 GNDA.n2010 GNDA.n110 53.3664
R2721 GNDA.n2011 GNDA.n109 53.3664
R2722 GNDA.n2015 GNDA.n108 53.3664
R2723 GNDA.n2019 GNDA.n107 53.3664
R2724 GNDA.n2007 GNDA.n110 53.3664
R2725 GNDA.n2014 GNDA.n109 53.3664
R2726 GNDA.n2018 GNDA.n108 53.3664
R2727 GNDA.n2021 GNDA.n107 53.3664
R2728 GNDA.n1991 GNDA.n98 53.3664
R2729 GNDA.n1995 GNDA.n105 53.3664
R2730 GNDA.n1999 GNDA.n96 53.3664
R2731 GNDA.n2003 GNDA.n106 53.3664
R2732 GNDA.n1974 GNDA.n104 53.3664
R2733 GNDA.n1978 GNDA.n103 53.3664
R2734 GNDA.n1982 GNDA.n102 53.3664
R2735 GNDA.n1986 GNDA.n101 53.3664
R2736 GNDA.n1970 GNDA.n99 53.3664
R2737 GNDA.n2047 GNDA.n94 53.3664
R2738 GNDA.n97 GNDA.n93 53.3664
R2739 GNDA.n2034 GNDA.n95 53.3664
R2740 GNDA.n232 GNDA.n195 53.3664
R2741 GNDA.n231 GNDA.n230 53.3664
R2742 GNDA.n224 GNDA.n197 53.3664
R2743 GNDA.n223 GNDA.n222 53.3664
R2744 GNDA.n214 GNDA.n213 53.3664
R2745 GNDA.n209 GNDA.n203 53.3664
R2746 GNDA.n207 GNDA.n206 53.3664
R2747 GNDA.n1879 GNDA.n180 53.3664
R2748 GNDA.n1850 GNDA.n1849 53.3664
R2749 GNDA.n1862 GNDA.n1861 53.3664
R2750 GNDA.n1865 GNDA.n1864 53.3664
R2751 GNDA.n1877 GNDA.n1876 53.3664
R2752 GNDA.n239 GNDA.n238 53.3664
R2753 GNDA.n241 GNDA.n240 53.3664
R2754 GNDA.n246 GNDA.n245 53.3664
R2755 GNDA.n249 GNDA.n248 53.3664
R2756 GNDA.n238 GNDA.n237 53.3664
R2757 GNDA.n240 GNDA.n193 53.3664
R2758 GNDA.n247 GNDA.n246 53.3664
R2759 GNDA.n248 GNDA.n191 53.3664
R2760 GNDA.n222 GNDA.n221 53.3664
R2761 GNDA.n225 GNDA.n224 53.3664
R2762 GNDA.n230 GNDA.n229 53.3664
R2763 GNDA.n233 GNDA.n232 53.3664
R2764 GNDA.n204 GNDA.n180 53.3664
R2765 GNDA.n208 GNDA.n207 53.3664
R2766 GNDA.n203 GNDA.n201 53.3664
R2767 GNDA.n215 GNDA.n214 53.3664
R2768 GNDA.n1878 GNDA.n1877 53.3664
R2769 GNDA.n1864 GNDA.n181 53.3664
R2770 GNDA.n1863 GNDA.n1862 53.3664
R2771 GNDA.n1849 GNDA.n186 53.3664
R2772 GNDA.n1912 GNDA.n163 52.7091
R2773 GNDA.n1906 GNDA.n163 52.7091
R2774 GNDA.n1906 GNDA.n1905 52.7091
R2775 GNDA.n1905 GNDA.n1904 52.7091
R2776 GNDA.n1904 GNDA.n167 52.7091
R2777 GNDA.n1898 GNDA.n1897 52.7091
R2778 GNDA.n1897 GNDA.n1896 52.7091
R2779 GNDA.n1896 GNDA.n171 52.7091
R2780 GNDA.n1890 GNDA.n171 52.7091
R2781 GNDA.n1890 GNDA.n1889 52.7091
R2782 GNDA.n1889 GNDA.n1888 52.7091
R2783 GNDA.n1888 GNDA.t103 52.7091
R2784 GNDA.n656 GNDA.n655 52.7091
R2785 GNDA.n656 GNDA.n493 52.7091
R2786 GNDA.n663 GNDA.n493 52.7091
R2787 GNDA.n664 GNDA.n663 52.7091
R2788 GNDA.n665 GNDA.n664 52.7091
R2789 GNDA.n669 GNDA.n668 52.7091
R2790 GNDA.n669 GNDA.n488 52.7091
R2791 GNDA.n676 GNDA.n488 52.7091
R2792 GNDA.n677 GNDA.n676 52.7091
R2793 GNDA.n678 GNDA.n677 52.7091
R2794 GNDA.n678 GNDA.n486 52.7091
R2795 GNDA.n1545 GNDA.n1544 52.7091
R2796 GNDA.n1544 GNDA.n1543 52.7091
R2797 GNDA.n1543 GNDA.n1511 52.7091
R2798 GNDA.n1537 GNDA.n1511 52.7091
R2799 GNDA.n1537 GNDA.n88 52.7091
R2800 GNDA.n1518 GNDA.n89 52.7091
R2801 GNDA.n1530 GNDA.n1518 52.7091
R2802 GNDA.n1530 GNDA.n1529 52.7091
R2803 GNDA.n1529 GNDA.n1528 52.7091
R2804 GNDA.n1528 GNDA.n1519 52.7091
R2805 GNDA.n1522 GNDA.n1519 52.7091
R2806 GNDA.t199 GNDA.n1708 51.4866
R2807 GNDA.t199 GNDA.n386 51.4866
R2808 GNDA.n2056 GNDA.n83 51.0266
R2809 GNDA.n2159 GNDA.t51 50.8162
R2810 GNDA.t39 GNDA.n2213 50.8162
R2811 GNDA.n2171 GNDA.t143 50.8162
R2812 GNDA.t101 GNDA.t301 49.9132
R2813 GNDA.t106 GNDA.t81 49.9132
R2814 GNDA.t48 GNDA.t295 49.9132
R2815 GNDA.t134 GNDA.t98 49.9132
R2816 GNDA.t163 GNDA.n2071 49.4271
R2817 GNDA.n1689 GNDA.t71 48.3974
R2818 GNDA.n647 GNDA.t199 47.6748
R2819 GNDA.n1680 GNDA.t289 47.3677
R2820 GNDA.n2055 GNDA.n2054 46.9641
R2821 GNDA.t130 GNDA.t245 46.338
R2822 GNDA.t234 GNDA.t63 46.338
R2823 GNDA.n1107 GNDA.t199 46.2335
R2824 GNDA.n1038 GNDA.t199 46.2335
R2825 GNDA.t199 GNDA.n155 46.2335
R2826 GNDA.n2098 GNDA.n2097 46.0738
R2827 GNDA.n2109 GNDA.n2108 46.0738
R2828 GNDA.n2203 GNDA.n2202 46.0738
R2829 GNDA.n2209 GNDA.n8 46.0738
R2830 GNDA.t77 GNDA.n2158 44.838
R2831 GNDA.n2214 GNDA.t73 44.838
R2832 GNDA.t294 GNDA.t25 44.0529
R2833 GNDA.t245 GNDA.n1443 43.2488
R2834 GNDA.n2072 GNDA.t163 43.2488
R2835 GNDA.n2040 GNDA.t179 43.2488
R2836 GNDA.t199 GNDA.n1106 42.2987
R2837 GNDA.n1947 GNDA.t199 42.2987
R2838 GNDA.n1922 GNDA.t199 42.2987
R2839 GNDA.t65 GNDA.t44 42.2405
R2840 GNDA.t311 GNDA.t65 42.2405
R2841 GNDA.t306 GNDA.t66 42.2405
R2842 GNDA.t307 GNDA.t306 42.2405
R2843 GNDA.n2060 GNDA.t26 42.2191
R2844 GNDA.t199 GNDA.t289 41.1894
R2845 GNDA.t199 GNDA.t71 41.1894
R2846 GNDA.n2159 GNDA.n2093 40.5993
R2847 GNDA.n2213 GNDA.n2212 40.5993
R2848 GNDA.n2054 GNDA.t150 40.4338
R2849 GNDA.n2054 GNDA.t313 40.4338
R2850 GNDA.n2094 GNDA.t213 40.4338
R2851 GNDA.n4 GNDA.t226 40.4338
R2852 GNDA.n2146 GNDA.t207 40.4338
R2853 GNDA.n2173 GNDA.t263 40.4338
R2854 GNDA.n2169 GNDA.t241 40.4338
R2855 GNDA.n25 GNDA.t288 40.4338
R2856 GNDA.n1477 GNDA.t159 39.1299
R2857 GNDA.n2084 GNDA.n2083 39.1299
R2858 GNDA.n1608 GNDA.t175 39.1299
R2859 GNDA.n1966 GNDA.t234 39.1299
R2860 GNDA.n82 GNDA.t152 38.6076
R2861 GNDA.n82 GNDA.t314 38.6076
R2862 GNDA.n1708 GNDA.n389 38.1002
R2863 GNDA.n1609 GNDA.n81 38.1002
R2864 GNDA.n2052 GNDA.t50 38.1002
R2865 GNDA.n1966 GNDA.t30 38.1002
R2866 GNDA.n2134 GNDA.n2133 37.5297
R2867 GNDA.n2132 GNDA.n2131 37.5297
R2868 GNDA.n2130 GNDA.n2129 37.5297
R2869 GNDA.n2128 GNDA.n2127 37.5297
R2870 GNDA.n2126 GNDA.n2125 37.5297
R2871 GNDA.n2124 GNDA.n2123 37.5297
R2872 GNDA.n2122 GNDA.n2121 37.5297
R2873 GNDA.n2120 GNDA.n2119 37.5297
R2874 GNDA.n2118 GNDA.n2117 37.5297
R2875 GNDA.n2116 GNDA.n2115 37.5297
R2876 GNDA.n2143 GNDA.n2142 37.5297
R2877 GNDA.n24 GNDA.n23 37.5297
R2878 GNDA.n1598 GNDA.n386 37.0705
R2879 GNDA.t185 GNDA.t199 36.0408
R2880 GNDA.t199 GNDA.t165 36.0408
R2881 GNDA.t199 GNDA.n167 35.7252
R2882 GNDA.n665 GNDA.t199 35.7252
R2883 GNDA.t199 GNDA.n88 35.7252
R2884 GNDA.t301 GNDA.t93 34.5555
R2885 GNDA.t69 GNDA.t106 34.5555
R2886 GNDA.t295 GNDA.t146 34.5555
R2887 GNDA.t100 GNDA.t134 34.5555
R2888 GNDA.n1443 GNDA.t24 33.9813
R2889 GNDA.n1444 GNDA.t95 33.9813
R2890 GNDA.n2059 GNDA.n2058 33.9813
R2891 GNDA.n1450 GNDA.t169 32.9516
R2892 GNDA.t191 GNDA.n1601 32.9516
R2893 GNDA.t181 GNDA.n134 32.9516
R2894 GNDA.n255 GNDA.t199 32.9056
R2895 GNDA.n369 GNDA.t199 32.9056
R2896 GNDA.n1959 GNDA.n117 32.3063
R2897 GNDA.n2110 GNDA.t266 31.1255
R2898 GNDA.n2096 GNDA.t256 31.1255
R2899 GNDA.n2204 GNDA.t283 31.1255
R2900 GNDA.n2208 GNDA.t210 31.1255
R2901 GNDA.t128 GNDA.t127 30.716
R2902 GNDA.n2224 GNDA.n0 29.8047
R2903 GNDA.t167 GNDA.n1465 28.8327
R2904 GNDA.t189 GNDA.n2070 28.8327
R2905 GNDA.t183 GNDA.n2029 28.8327
R2906 GNDA.n1465 GNDA.t300 27.803
R2907 GNDA.n1449 GNDA.t1 27.803
R2908 GNDA.n1479 GNDA.t87 27.803
R2909 GNDA.n1207 GNDA.n1206 27.5561
R2910 GNDA.n982 GNDA.n906 27.5561
R2911 GNDA.n1423 GNDA.n1420 27.5561
R2912 GNDA.n1651 GNDA.n1648 27.5561
R2913 GNDA.n862 GNDA.n861 27.5561
R2914 GNDA.n318 GNDA.n317 27.5561
R2915 GNDA.n741 GNDA.n740 27.5561
R2916 GNDA.n2008 GNDA.n2005 27.5561
R2917 GNDA.n236 GNDA.n235 27.5561
R2918 GNDA.t114 GNDA.n2152 26.8766
R2919 GNDA.n2186 GNDA.t9 26.8766
R2920 GNDA.n1189 GNDA.n1188 26.6672
R2921 GNDA.n960 GNDA.n910 26.6672
R2922 GNDA.n1404 GNDA.n1403 26.6672
R2923 GNDA.n1632 GNDA.n1631 26.6672
R2924 GNDA.n844 GNDA.n843 26.6672
R2925 GNDA.n301 GNDA.n300 26.6672
R2926 GNDA.n723 GNDA.n722 26.6672
R2927 GNDA.n1989 GNDA.n1988 26.6672
R2928 GNDA.n219 GNDA.n218 26.6672
R2929 GNDA.t1 GNDA.t159 25.7435
R2930 GNDA.t179 GNDA.t78 25.7435
R2931 GNDA.n431 GNDA.t168 24.0005
R2932 GNDA.n431 GNDA.t158 24.0005
R2933 GNDA.n429 GNDA.t186 24.0005
R2934 GNDA.n429 GNDA.t170 24.0005
R2935 GNDA.n390 GNDA.t160 24.0005
R2936 GNDA.n390 GNDA.t188 24.0005
R2937 GNDA.n1703 GNDA.t174 24.0005
R2938 GNDA.n1703 GNDA.t164 24.0005
R2939 GNDA.n1701 GNDA.t190 24.0005
R2940 GNDA.n1701 GNDA.t172 24.0005
R2941 GNDA.n1699 GNDA.t162 24.0005
R2942 GNDA.n1699 GNDA.t192 24.0005
R2943 GNDA.n1697 GNDA.t176 24.0005
R2944 GNDA.n1697 GNDA.t178 24.0005
R2945 GNDA.n1687 GNDA.t156 24.0005
R2946 GNDA.n1687 GNDA.t180 24.0005
R2947 GNDA.n1685 GNDA.t184 24.0005
R2948 GNDA.n1685 GNDA.t166 24.0005
R2949 GNDA.n137 GNDA.t154 24.0005
R2950 GNDA.n137 GNDA.t182 24.0005
R2951 GNDA.n2027 GNDA.t140 23.6841
R2952 GNDA.t78 GNDA.n2039 23.6841
R2953 GNDA.n134 GNDA.t74 23.6841
R2954 GNDA.n1683 GNDA.n1682 23.1624
R2955 GNDA.n1707 GNDA.n1706 23.1624
R2956 GNDA.n1695 GNDA.n1694 23.1624
R2957 GNDA.n1692 GNDA.n1691 23.1624
R2958 GNDA.n1963 GNDA.n1962 23.1624
R2959 GNDA.n434 GNDA.n433 23.1624
R2960 GNDA.t173 GNDA.n2059 22.6544
R2961 GNDA.n2041 GNDA.t155 22.6544
R2962 GNDA.n1956 GNDA.n1955 21.0192
R2963 GNDA.t64 GNDA.t126 20.9779
R2964 GNDA.n2158 GNDA.t43 20.9249
R2965 GNDA.t6 GNDA.n2214 20.9249
R2966 GNDA.n1448 GNDA.t199 20.5949
R2967 GNDA.t23 GNDA.n1448 20.5949
R2968 GNDA.n1681 GNDA.t87 20.5949
R2969 GNDA.n1690 GNDA.t140 20.5949
R2970 GNDA.n2053 GNDA.t32 20.5949
R2971 GNDA.n2053 GNDA.t199 20.5949
R2972 GNDA.n1015 GNDA.t199 19.9378
R2973 GNDA.n37 GNDA.t297 19.7005
R2974 GNDA.n37 GNDA.t315 19.7005
R2975 GNDA.n35 GNDA.t316 19.7005
R2976 GNDA.n35 GNDA.t31 19.7005
R2977 GNDA.n33 GNDA.t84 19.7005
R2978 GNDA.n33 GNDA.t52 19.7005
R2979 GNDA.n31 GNDA.t122 19.7005
R2980 GNDA.n31 GNDA.t97 19.7005
R2981 GNDA.n30 GNDA.t293 19.7005
R2982 GNDA.n30 GNDA.t82 19.7005
R2983 GNDA.n29 GNDA.t40 19.7005
R2984 GNDA.n29 GNDA.t292 19.7005
R2985 GNDA.n17 GNDA.t35 19.7005
R2986 GNDA.n17 GNDA.t92 19.7005
R2987 GNDA.n15 GNDA.t17 19.7005
R2988 GNDA.n15 GNDA.t37 19.7005
R2989 GNDA.n13 GNDA.t147 19.7005
R2990 GNDA.n13 GNDA.t36 19.7005
R2991 GNDA.n11 GNDA.t46 19.7005
R2992 GNDA.n11 GNDA.t47 19.7005
R2993 GNDA.n10 GNDA.t129 19.7005
R2994 GNDA.n10 GNDA.t291 19.7005
R2995 GNDA.n9 GNDA.t290 19.7005
R2996 GNDA.n9 GNDA.t80 19.7005
R2997 GNDA.n1021 GNDA.t199 19.6741
R2998 GNDA.t298 GNDA.t53 19.1977
R2999 GNDA.t123 GNDA.t104 19.1977
R3000 GNDA.n2145 GNDA.t13 19.1977
R3001 GNDA.n2174 GNDA.t94 19.1977
R3002 GNDA.n2218 GNDA.t116 19.1977
R3003 GNDA.t18 GNDA.t33 19.1977
R3004 GNDA.t99 GNDA.t28 19.1977
R3005 GNDA.n2224 GNDA.n2223 19.008
R3006 GNDA.t25 GNDA.t88 18.8801
R3007 GNDA.n1951 GNDA.n1950 18.5605
R3008 GNDA.n1478 GNDA.t187 18.5355
R3009 GNDA.n1609 GNDA.t177 18.5355
R3010 GNDA.n2210 GNDA.t133 18.3557
R3011 GNDA GNDA.n85 18.1546
R3012 GNDA.n652 GNDA.n495 17.5843
R3013 GNDA.n1548 GNDA.n1508 17.5843
R3014 GNDA.n1910 GNDA.n161 17.5843
R3015 GNDA.n435 GNDA.t199 17.5058
R3016 GNDA.n1964 GNDA.n136 17.5058
R3017 GNDA.t85 GNDA.n121 17.1379
R3018 GNDA.n1898 GNDA.t199 16.9844
R3019 GNDA.n668 GNDA.t199 16.9844
R3020 GNDA.t199 GNDA.n89 16.9844
R3021 GNDA.n1261 GNDA.n1118 16.9379
R3022 GNDA.n625 GNDA.n622 16.9379
R3023 GNDA.n1364 GNDA.n1363 16.9379
R3024 GNDA.n593 GNDA.n254 16.7709
R3025 GNDA.n1715 GNDA.n1714 16.7709
R3026 GNDA.n1342 GNDA.n368 16.7709
R3027 GNDA.n1744 GNDA.n1743 16.7709
R3028 GNDA.n20 GNDA.n19 16.4693
R3029 GNDA.n1221 GNDA.n1207 16.0005
R3030 GNDA.n1221 GNDA.n1220 16.0005
R3031 GNDA.n1220 GNDA.n1219 16.0005
R3032 GNDA.n1219 GNDA.n1216 16.0005
R3033 GNDA.n1216 GNDA.n1215 16.0005
R3034 GNDA.n1215 GNDA.n1212 16.0005
R3035 GNDA.n1212 GNDA.n1211 16.0005
R3036 GNDA.n1211 GNDA.n1208 16.0005
R3037 GNDA.n1206 GNDA.n1204 16.0005
R3038 GNDA.n1204 GNDA.n1201 16.0005
R3039 GNDA.n1201 GNDA.n1200 16.0005
R3040 GNDA.n1200 GNDA.n1197 16.0005
R3041 GNDA.n1197 GNDA.n1196 16.0005
R3042 GNDA.n1196 GNDA.n1193 16.0005
R3043 GNDA.n1193 GNDA.n1192 16.0005
R3044 GNDA.n1192 GNDA.n1189 16.0005
R3045 GNDA.n1188 GNDA.n1185 16.0005
R3046 GNDA.n1185 GNDA.n1184 16.0005
R3047 GNDA.n1184 GNDA.n1181 16.0005
R3048 GNDA.n1181 GNDA.n1180 16.0005
R3049 GNDA.n1180 GNDA.n1177 16.0005
R3050 GNDA.n1177 GNDA.n1176 16.0005
R3051 GNDA.n1176 GNDA.n1173 16.0005
R3052 GNDA.n1173 GNDA.n1172 16.0005
R3053 GNDA.n983 GNDA.n982 16.0005
R3054 GNDA.n984 GNDA.n983 16.0005
R3055 GNDA.n984 GNDA.n904 16.0005
R3056 GNDA.n990 GNDA.n904 16.0005
R3057 GNDA.n991 GNDA.n990 16.0005
R3058 GNDA.n992 GNDA.n991 16.0005
R3059 GNDA.n992 GNDA.n902 16.0005
R3060 GNDA.n902 GNDA.n451 16.0005
R3061 GNDA.n976 GNDA.n906 16.0005
R3062 GNDA.n976 GNDA.n975 16.0005
R3063 GNDA.n975 GNDA.n974 16.0005
R3064 GNDA.n974 GNDA.n908 16.0005
R3065 GNDA.n968 GNDA.n908 16.0005
R3066 GNDA.n968 GNDA.n967 16.0005
R3067 GNDA.n967 GNDA.n966 16.0005
R3068 GNDA.n966 GNDA.n910 16.0005
R3069 GNDA.n960 GNDA.n959 16.0005
R3070 GNDA.n959 GNDA.n958 16.0005
R3071 GNDA.n958 GNDA.n912 16.0005
R3072 GNDA.n953 GNDA.n912 16.0005
R3073 GNDA.n953 GNDA.n952 16.0005
R3074 GNDA.n952 GNDA.n951 16.0005
R3075 GNDA.n951 GNDA.n915 16.0005
R3076 GNDA.n946 GNDA.n915 16.0005
R3077 GNDA.n1424 GNDA.n1423 16.0005
R3078 GNDA.n1427 GNDA.n1424 16.0005
R3079 GNDA.n1428 GNDA.n1427 16.0005
R3080 GNDA.n1431 GNDA.n1428 16.0005
R3081 GNDA.n1432 GNDA.n1431 16.0005
R3082 GNDA.n1435 GNDA.n1432 16.0005
R3083 GNDA.n1437 GNDA.n1435 16.0005
R3084 GNDA.n1438 GNDA.n1437 16.0005
R3085 GNDA.n1420 GNDA.n1419 16.0005
R3086 GNDA.n1419 GNDA.n1416 16.0005
R3087 GNDA.n1416 GNDA.n1415 16.0005
R3088 GNDA.n1415 GNDA.n1412 16.0005
R3089 GNDA.n1412 GNDA.n1411 16.0005
R3090 GNDA.n1411 GNDA.n1408 16.0005
R3091 GNDA.n1408 GNDA.n1407 16.0005
R3092 GNDA.n1407 GNDA.n1404 16.0005
R3093 GNDA.n1403 GNDA.n1400 16.0005
R3094 GNDA.n1400 GNDA.n1399 16.0005
R3095 GNDA.n1399 GNDA.n1396 16.0005
R3096 GNDA.n1396 GNDA.n1395 16.0005
R3097 GNDA.n1395 GNDA.n1392 16.0005
R3098 GNDA.n1392 GNDA.n1391 16.0005
R3099 GNDA.n1391 GNDA.n1388 16.0005
R3100 GNDA.n1388 GNDA.n398 16.0005
R3101 GNDA.n1652 GNDA.n1651 16.0005
R3102 GNDA.n1655 GNDA.n1652 16.0005
R3103 GNDA.n1656 GNDA.n1655 16.0005
R3104 GNDA.n1659 GNDA.n1656 16.0005
R3105 GNDA.n1660 GNDA.n1659 16.0005
R3106 GNDA.n1663 GNDA.n1660 16.0005
R3107 GNDA.n1665 GNDA.n1663 16.0005
R3108 GNDA.n1666 GNDA.n1665 16.0005
R3109 GNDA.n1648 GNDA.n1647 16.0005
R3110 GNDA.n1647 GNDA.n1644 16.0005
R3111 GNDA.n1644 GNDA.n1643 16.0005
R3112 GNDA.n1643 GNDA.n1640 16.0005
R3113 GNDA.n1640 GNDA.n1639 16.0005
R3114 GNDA.n1639 GNDA.n1636 16.0005
R3115 GNDA.n1636 GNDA.n1635 16.0005
R3116 GNDA.n1635 GNDA.n1632 16.0005
R3117 GNDA.n1631 GNDA.n1628 16.0005
R3118 GNDA.n1628 GNDA.n1627 16.0005
R3119 GNDA.n1627 GNDA.n1624 16.0005
R3120 GNDA.n1624 GNDA.n1623 16.0005
R3121 GNDA.n1623 GNDA.n1620 16.0005
R3122 GNDA.n1620 GNDA.n1619 16.0005
R3123 GNDA.n1619 GNDA.n1616 16.0005
R3124 GNDA.n1616 GNDA.n1615 16.0005
R3125 GNDA.n876 GNDA.n862 16.0005
R3126 GNDA.n876 GNDA.n875 16.0005
R3127 GNDA.n875 GNDA.n874 16.0005
R3128 GNDA.n874 GNDA.n871 16.0005
R3129 GNDA.n871 GNDA.n870 16.0005
R3130 GNDA.n870 GNDA.n867 16.0005
R3131 GNDA.n867 GNDA.n866 16.0005
R3132 GNDA.n866 GNDA.n863 16.0005
R3133 GNDA.n861 GNDA.n859 16.0005
R3134 GNDA.n859 GNDA.n856 16.0005
R3135 GNDA.n856 GNDA.n855 16.0005
R3136 GNDA.n855 GNDA.n852 16.0005
R3137 GNDA.n852 GNDA.n851 16.0005
R3138 GNDA.n851 GNDA.n848 16.0005
R3139 GNDA.n848 GNDA.n847 16.0005
R3140 GNDA.n847 GNDA.n844 16.0005
R3141 GNDA.n843 GNDA.n840 16.0005
R3142 GNDA.n840 GNDA.n839 16.0005
R3143 GNDA.n839 GNDA.n836 16.0005
R3144 GNDA.n836 GNDA.n835 16.0005
R3145 GNDA.n835 GNDA.n832 16.0005
R3146 GNDA.n832 GNDA.n831 16.0005
R3147 GNDA.n831 GNDA.n828 16.0005
R3148 GNDA.n828 GNDA.n827 16.0005
R3149 GNDA.n318 GNDA.n276 16.0005
R3150 GNDA.n324 GNDA.n276 16.0005
R3151 GNDA.n325 GNDA.n324 16.0005
R3152 GNDA.n326 GNDA.n325 16.0005
R3153 GNDA.n326 GNDA.n274 16.0005
R3154 GNDA.n332 GNDA.n274 16.0005
R3155 GNDA.n333 GNDA.n332 16.0005
R3156 GNDA.n1751 GNDA.n333 16.0005
R3157 GNDA.n317 GNDA.n316 16.0005
R3158 GNDA.n316 GNDA.n278 16.0005
R3159 GNDA.n310 GNDA.n278 16.0005
R3160 GNDA.n310 GNDA.n309 16.0005
R3161 GNDA.n309 GNDA.n308 16.0005
R3162 GNDA.n308 GNDA.n280 16.0005
R3163 GNDA.n302 GNDA.n280 16.0005
R3164 GNDA.n302 GNDA.n301 16.0005
R3165 GNDA.n300 GNDA.n282 16.0005
R3166 GNDA.n294 GNDA.n282 16.0005
R3167 GNDA.n294 GNDA.n293 16.0005
R3168 GNDA.n293 GNDA.n292 16.0005
R3169 GNDA.n292 GNDA.n284 16.0005
R3170 GNDA.n287 GNDA.n284 16.0005
R3171 GNDA.n287 GNDA.n261 16.0005
R3172 GNDA.n1786 GNDA.n261 16.0005
R3173 GNDA.n1955 GNDA.n139 16.0005
R3174 GNDA.n1951 GNDA.n139 16.0005
R3175 GNDA.n755 GNDA.n741 16.0005
R3176 GNDA.n755 GNDA.n754 16.0005
R3177 GNDA.n754 GNDA.n753 16.0005
R3178 GNDA.n753 GNDA.n750 16.0005
R3179 GNDA.n750 GNDA.n749 16.0005
R3180 GNDA.n749 GNDA.n746 16.0005
R3181 GNDA.n746 GNDA.n745 16.0005
R3182 GNDA.n745 GNDA.n742 16.0005
R3183 GNDA.n740 GNDA.n738 16.0005
R3184 GNDA.n738 GNDA.n735 16.0005
R3185 GNDA.n735 GNDA.n734 16.0005
R3186 GNDA.n734 GNDA.n731 16.0005
R3187 GNDA.n731 GNDA.n730 16.0005
R3188 GNDA.n730 GNDA.n727 16.0005
R3189 GNDA.n727 GNDA.n726 16.0005
R3190 GNDA.n726 GNDA.n723 16.0005
R3191 GNDA.n722 GNDA.n719 16.0005
R3192 GNDA.n719 GNDA.n718 16.0005
R3193 GNDA.n718 GNDA.n715 16.0005
R3194 GNDA.n715 GNDA.n714 16.0005
R3195 GNDA.n714 GNDA.n711 16.0005
R3196 GNDA.n711 GNDA.n710 16.0005
R3197 GNDA.n710 GNDA.n707 16.0005
R3198 GNDA.n707 GNDA.n706 16.0005
R3199 GNDA.n2009 GNDA.n2008 16.0005
R3200 GNDA.n2012 GNDA.n2009 16.0005
R3201 GNDA.n2013 GNDA.n2012 16.0005
R3202 GNDA.n2016 GNDA.n2013 16.0005
R3203 GNDA.n2017 GNDA.n2016 16.0005
R3204 GNDA.n2020 GNDA.n2017 16.0005
R3205 GNDA.n2022 GNDA.n2020 16.0005
R3206 GNDA.n2023 GNDA.n2022 16.0005
R3207 GNDA.n2005 GNDA.n2004 16.0005
R3208 GNDA.n2004 GNDA.n2001 16.0005
R3209 GNDA.n2001 GNDA.n2000 16.0005
R3210 GNDA.n2000 GNDA.n1997 16.0005
R3211 GNDA.n1997 GNDA.n1996 16.0005
R3212 GNDA.n1996 GNDA.n1993 16.0005
R3213 GNDA.n1993 GNDA.n1992 16.0005
R3214 GNDA.n1992 GNDA.n1989 16.0005
R3215 GNDA.n1988 GNDA.n1985 16.0005
R3216 GNDA.n1985 GNDA.n1984 16.0005
R3217 GNDA.n1984 GNDA.n1981 16.0005
R3218 GNDA.n1981 GNDA.n1980 16.0005
R3219 GNDA.n1980 GNDA.n1977 16.0005
R3220 GNDA.n1977 GNDA.n1976 16.0005
R3221 GNDA.n1976 GNDA.n1973 16.0005
R3222 GNDA.n1973 GNDA.n1972 16.0005
R3223 GNDA.n236 GNDA.n194 16.0005
R3224 GNDA.n242 GNDA.n194 16.0005
R3225 GNDA.n243 GNDA.n242 16.0005
R3226 GNDA.n244 GNDA.n243 16.0005
R3227 GNDA.n244 GNDA.n192 16.0005
R3228 GNDA.n250 GNDA.n192 16.0005
R3229 GNDA.n251 GNDA.n250 16.0005
R3230 GNDA.n1845 GNDA.n251 16.0005
R3231 GNDA.n235 GNDA.n234 16.0005
R3232 GNDA.n234 GNDA.n196 16.0005
R3233 GNDA.n228 GNDA.n196 16.0005
R3234 GNDA.n228 GNDA.n227 16.0005
R3235 GNDA.n227 GNDA.n226 16.0005
R3236 GNDA.n226 GNDA.n198 16.0005
R3237 GNDA.n220 GNDA.n198 16.0005
R3238 GNDA.n220 GNDA.n219 16.0005
R3239 GNDA.n218 GNDA.n200 16.0005
R3240 GNDA.n212 GNDA.n200 16.0005
R3241 GNDA.n212 GNDA.n211 16.0005
R3242 GNDA.n211 GNDA.n210 16.0005
R3243 GNDA.n210 GNDA.n202 16.0005
R3244 GNDA.n205 GNDA.n202 16.0005
R3245 GNDA.n205 GNDA.n179 16.0005
R3246 GNDA.n1880 GNDA.n179 16.0005
R3247 GNDA.n2102 GNDA.n2101 15.8233
R3248 GNDA.n2196 GNDA.n2195 15.8233
R3249 GNDA.t187 GNDA.t131 15.4463
R3250 GNDA.t155 GNDA.t79 15.4463
R3251 GNDA.t0 GNDA.n2159 14.9467
R3252 GNDA.n2213 GNDA.t8 14.9467
R3253 GNDA.t2 GNDA.n2171 14.9467
R3254 GNDA.n255 GNDA.n176 14.555
R3255 GNDA.n1006 GNDA.n369 14.555
R3256 GNDA.n433 GNDA.n432 14.363
R3257 GNDA.n1684 GNDA.n1683 13.8005
R3258 GNDA.n1706 GNDA.n1705 13.8005
R3259 GNDA.n1696 GNDA.n1695 13.8005
R3260 GNDA.n1693 GNDA.n1692 13.8005
R3261 GNDA.n1962 GNDA.n1961 13.8005
R3262 GNDA.n2055 GNDA.n86 12.7542
R3263 GNDA.n2099 GNDA.t195 12.6791
R3264 GNDA.n2193 GNDA.t286 12.6791
R3265 GNDA.n2201 GNDA.t205 12.6791
R3266 GNDA.n2107 GNDA.t259 12.6791
R3267 GNDA.n1444 GNDA.t185 12.3572
R3268 GNDA.n2083 GNDA.t161 12.3572
R3269 GNDA.t153 GNDA.n128 12.3572
R3270 GNDA.n2057 GNDA.n2056 12.2193
R3271 GNDA.n2190 GNDA.n2189 12.1151
R3272 GNDA.n40 GNDA.n39 11.7193
R3273 GNDA.t75 GNDA.t103 11.7135
R3274 GNDA.n1261 GNDA.n1260 11.6369
R3275 GNDA.n1260 GNDA.n1259 11.6369
R3276 GNDA.n1259 GNDA.n1258 11.6369
R3277 GNDA.n1258 GNDA.n1256 11.6369
R3278 GNDA.n1256 GNDA.n1253 11.6369
R3279 GNDA.n1253 GNDA.n1252 11.6369
R3280 GNDA.n1252 GNDA.n1249 11.6369
R3281 GNDA.n1249 GNDA.n1248 11.6369
R3282 GNDA.n1248 GNDA.n1245 11.6369
R3283 GNDA.n1245 GNDA.n1244 11.6369
R3284 GNDA.n1118 GNDA.n1117 11.6369
R3285 GNDA.n1117 GNDA.n1019 11.6369
R3286 GNDA.n1111 GNDA.n1019 11.6369
R3287 GNDA.n1111 GNDA.n1110 11.6369
R3288 GNDA.n1110 GNDA.n1109 11.6369
R3289 GNDA.n1109 GNDA.n1024 11.6369
R3290 GNDA.n1103 GNDA.n1024 11.6369
R3291 GNDA.n1103 GNDA.n1102 11.6369
R3292 GNDA.n1102 GNDA.n1101 11.6369
R3293 GNDA.n1101 GNDA.n1028 11.6369
R3294 GNDA.n1095 GNDA.n1028 11.6369
R3295 GNDA.n622 GNDA.n621 11.6369
R3296 GNDA.n621 GNDA.n618 11.6369
R3297 GNDA.n618 GNDA.n617 11.6369
R3298 GNDA.n617 GNDA.n614 11.6369
R3299 GNDA.n614 GNDA.n613 11.6369
R3300 GNDA.n613 GNDA.n610 11.6369
R3301 GNDA.n610 GNDA.n609 11.6369
R3302 GNDA.n609 GNDA.n606 11.6369
R3303 GNDA.n606 GNDA.n605 11.6369
R3304 GNDA.n605 GNDA.n450 11.6369
R3305 GNDA.n626 GNDA.n625 11.6369
R3306 GNDA.n629 GNDA.n626 11.6369
R3307 GNDA.n630 GNDA.n629 11.6369
R3308 GNDA.n633 GNDA.n630 11.6369
R3309 GNDA.n634 GNDA.n633 11.6369
R3310 GNDA.n637 GNDA.n634 11.6369
R3311 GNDA.n638 GNDA.n637 11.6369
R3312 GNDA.n641 GNDA.n638 11.6369
R3313 GNDA.n642 GNDA.n641 11.6369
R3314 GNDA.n643 GNDA.n642 11.6369
R3315 GNDA.n643 GNDA.n336 11.6369
R3316 GNDA.n1364 GNDA.n1269 11.6369
R3317 GNDA.n1370 GNDA.n1269 11.6369
R3318 GNDA.n1371 GNDA.n1370 11.6369
R3319 GNDA.n1372 GNDA.n1371 11.6369
R3320 GNDA.n1372 GNDA.n1267 11.6369
R3321 GNDA.n1378 GNDA.n1267 11.6369
R3322 GNDA.n1379 GNDA.n1378 11.6369
R3323 GNDA.n1380 GNDA.n1379 11.6369
R3324 GNDA.n1380 GNDA.n1265 11.6369
R3325 GNDA.n1265 GNDA.n437 11.6369
R3326 GNDA.n510 GNDA.n337 11.6369
R3327 GNDA.n513 GNDA.n510 11.6369
R3328 GNDA.n514 GNDA.n513 11.6369
R3329 GNDA.n517 GNDA.n514 11.6369
R3330 GNDA.n518 GNDA.n517 11.6369
R3331 GNDA.n521 GNDA.n518 11.6369
R3332 GNDA.n522 GNDA.n521 11.6369
R3333 GNDA.n525 GNDA.n522 11.6369
R3334 GNDA.n527 GNDA.n525 11.6369
R3335 GNDA.n528 GNDA.n527 11.6369
R3336 GNDA.n594 GNDA.n528 11.6369
R3337 GNDA.n544 GNDA.n543 11.6369
R3338 GNDA.n543 GNDA.n540 11.6369
R3339 GNDA.n540 GNDA.n539 11.6369
R3340 GNDA.n539 GNDA.n536 11.6369
R3341 GNDA.n536 GNDA.n535 11.6369
R3342 GNDA.n535 GNDA.n532 11.6369
R3343 GNDA.n532 GNDA.n531 11.6369
R3344 GNDA.n531 GNDA.n529 11.6369
R3345 GNDA.n529 GNDA.n497 11.6369
R3346 GNDA.n651 GNDA.n497 11.6369
R3347 GNDA.n652 GNDA.n651 11.6369
R3348 GNDA.n658 GNDA.n495 11.6369
R3349 GNDA.n659 GNDA.n658 11.6369
R3350 GNDA.n661 GNDA.n659 11.6369
R3351 GNDA.n661 GNDA.n660 11.6369
R3352 GNDA.n660 GNDA.n492 11.6369
R3353 GNDA.n492 GNDA.n490 11.6369
R3354 GNDA.n671 GNDA.n490 11.6369
R3355 GNDA.n672 GNDA.n671 11.6369
R3356 GNDA.n674 GNDA.n672 11.6369
R3357 GNDA.n674 GNDA.n673 11.6369
R3358 GNDA.n1564 GNDA.n375 11.6369
R3359 GNDA.n1564 GNDA.n1563 11.6369
R3360 GNDA.n1563 GNDA.n1562 11.6369
R3361 GNDA.n1562 GNDA.n1502 11.6369
R3362 GNDA.n1557 GNDA.n1502 11.6369
R3363 GNDA.n1557 GNDA.n1556 11.6369
R3364 GNDA.n1556 GNDA.n1555 11.6369
R3365 GNDA.n1555 GNDA.n1505 11.6369
R3366 GNDA.n1550 GNDA.n1505 11.6369
R3367 GNDA.n1550 GNDA.n1549 11.6369
R3368 GNDA.n1549 GNDA.n1548 11.6369
R3369 GNDA.n1513 GNDA.n1508 11.6369
R3370 GNDA.n1541 GNDA.n1513 11.6369
R3371 GNDA.n1541 GNDA.n1540 11.6369
R3372 GNDA.n1540 GNDA.n1539 11.6369
R3373 GNDA.n1539 GNDA.n1514 11.6369
R3374 GNDA.n1534 GNDA.n1514 11.6369
R3375 GNDA.n1534 GNDA.n1533 11.6369
R3376 GNDA.n1533 GNDA.n1532 11.6369
R3377 GNDA.n1532 GNDA.n1516 11.6369
R3378 GNDA.n1526 GNDA.n1516 11.6369
R3379 GNDA.n1910 GNDA.n1909 11.6369
R3380 GNDA.n1909 GNDA.n1908 11.6369
R3381 GNDA.n1908 GNDA.n165 11.6369
R3382 GNDA.n1902 GNDA.n165 11.6369
R3383 GNDA.n1902 GNDA.n1901 11.6369
R3384 GNDA.n1901 GNDA.n1900 11.6369
R3385 GNDA.n1900 GNDA.n169 11.6369
R3386 GNDA.n1894 GNDA.n169 11.6369
R3387 GNDA.n1894 GNDA.n1893 11.6369
R3388 GNDA.n1893 GNDA.n1892 11.6369
R3389 GNDA.n1934 GNDA.n1933 11.6369
R3390 GNDA.n1933 GNDA.n1932 11.6369
R3391 GNDA.n1932 GNDA.n153 11.6369
R3392 GNDA.n1926 GNDA.n153 11.6369
R3393 GNDA.n1926 GNDA.n1925 11.6369
R3394 GNDA.n1925 GNDA.n1924 11.6369
R3395 GNDA.n1924 GNDA.n157 11.6369
R3396 GNDA.n1918 GNDA.n157 11.6369
R3397 GNDA.n1918 GNDA.n1917 11.6369
R3398 GNDA.n1917 GNDA.n1916 11.6369
R3399 GNDA.n1916 GNDA.n161 11.6369
R3400 GNDA.n1037 GNDA.n1032 11.6369
R3401 GNDA.n1043 GNDA.n1037 11.6369
R3402 GNDA.n1043 GNDA.n1042 11.6369
R3403 GNDA.n1042 GNDA.n1041 11.6369
R3404 GNDA.n1041 GNDA.n140 11.6369
R3405 GNDA.n1949 GNDA.n141 11.6369
R3406 GNDA.n1943 GNDA.n141 11.6369
R3407 GNDA.n1943 GNDA.n1942 11.6369
R3408 GNDA.n1942 GNDA.n1941 11.6369
R3409 GNDA.n1941 GNDA.n146 11.6369
R3410 GNDA.n1303 GNDA.n1280 11.6369
R3411 GNDA.n1303 GNDA.n1302 11.6369
R3412 GNDA.n1302 GNDA.n1301 11.6369
R3413 GNDA.n1301 GNDA.n1283 11.6369
R3414 GNDA.n1296 GNDA.n1283 11.6369
R3415 GNDA.n1296 GNDA.n1295 11.6369
R3416 GNDA.n1295 GNDA.n1294 11.6369
R3417 GNDA.n1294 GNDA.n1286 11.6369
R3418 GNDA.n1289 GNDA.n1286 11.6369
R3419 GNDA.n1289 GNDA.n377 11.6369
R3420 GNDA.n1713 GNDA.n377 11.6369
R3421 GNDA.n1363 GNDA.n1362 11.6369
R3422 GNDA.n1362 GNDA.n1271 11.6369
R3423 GNDA.n1357 GNDA.n1271 11.6369
R3424 GNDA.n1357 GNDA.n1356 11.6369
R3425 GNDA.n1356 GNDA.n1355 11.6369
R3426 GNDA.n1355 GNDA.n1274 11.6369
R3427 GNDA.n1350 GNDA.n1274 11.6369
R3428 GNDA.n1350 GNDA.n1349 11.6369
R3429 GNDA.n1349 GNDA.n1348 11.6369
R3430 GNDA.n1348 GNDA.n1277 11.6369
R3431 GNDA.n1343 GNDA.n1277 11.6369
R3432 GNDA.n1961 GNDA.n1960 11.3792
R3433 GNDA.n2104 GNDA.n2103 11.3233
R3434 GNDA.n2198 GNDA.n2197 11.3233
R3435 GNDA.n20 GNDA.n3 10.8286
R3436 GNDA.t90 GNDA.t75 9.95658
R3437 GNDA.n1958 GNDA.n0 9.75668
R3438 GNDA.n2133 GNDA.t125 9.6005
R3439 GNDA.n2133 GNDA.t113 9.6005
R3440 GNDA.n2131 GNDA.t57 9.6005
R3441 GNDA.n2131 GNDA.t111 9.6005
R3442 GNDA.n2129 GNDA.t5 9.6005
R3443 GNDA.n2129 GNDA.t115 9.6005
R3444 GNDA.n2127 GNDA.t139 9.6005
R3445 GNDA.n2127 GNDA.t14 9.6005
R3446 GNDA.n2125 GNDA.t144 9.6005
R3447 GNDA.n2125 GNDA.t60 9.6005
R3448 GNDA.n2123 GNDA.t109 9.6005
R3449 GNDA.n2123 GNDA.t16 9.6005
R3450 GNDA.n2121 GNDA.t108 9.6005
R3451 GNDA.n2121 GNDA.t62 9.6005
R3452 GNDA.n2119 GNDA.t10 9.6005
R3453 GNDA.n2119 GNDA.t137 9.6005
R3454 GNDA.n2117 GNDA.t117 9.6005
R3455 GNDA.n2117 GNDA.t142 9.6005
R3456 GNDA.n2115 GNDA.t59 9.6005
R3457 GNDA.n2115 GNDA.t225 9.6005
R3458 GNDA.n2142 GNDA.t3 9.6005
R3459 GNDA.n2142 GNDA.t12 9.6005
R3460 GNDA.n23 GNDA.t72 9.6005
R3461 GNDA.n23 GNDA.t70 9.6005
R3462 GNDA.n2181 GNDA.n2180 8.79217
R3463 GNDA.n2112 GNDA.n2095 8.67238
R3464 GNDA.n2207 GNDA.n2206 8.67238
R3465 GNDA.n1838 GNDA.n255 8.60107
R3466 GNDA.n1717 GNDA.n369 8.60107
R3467 GNDA.t157 GNDA.n1464 8.23827
R3468 GNDA.t171 GNDA.n2060 8.23827
R3469 GNDA.t165 GNDA.n2052 8.23827
R3470 GNDA.n2141 GNDA.n2140 8.11508
R3471 GNDA.n2150 GNDA.n2149 8.11508
R3472 GNDA.n2189 GNDA.n2188 8.11508
R3473 GNDA.t228 GNDA.t4 7.67938
R3474 GNDA.t49 GNDA.t116 7.67938
R3475 GNDA.n85 GNDA.n84 7.56675
R3476 GNDA.n1958 GNDA.n1957 7.56675
R3477 GNDA.n2198 GNDA.n3 7.53175
R3478 GNDA.n2104 GNDA.n2 7.53175
R3479 GNDA.n2137 GNDA.n2136 7.5005
R3480 GNDA.t67 GNDA.n1478 7.20855
R3481 GNDA.n2029 GNDA.t32 7.20855
R3482 GNDA.t63 GNDA.n135 7.20855
R3483 GNDA.n1965 GNDA.n1964 7.20855
R3484 GNDA.n2222 GNDA.n2 6.78175
R3485 GNDA.n1095 GNDA.n1094 6.72373
R3486 GNDA.n1743 GNDA.n336 6.72373
R3487 GNDA.n594 GNDA.n593 6.72373
R3488 GNDA.n152 GNDA.n146 6.72373
R3489 GNDA.n1714 GNDA.n1713 6.72373
R3490 GNDA.n1343 GNDA.n1342 6.72373
R3491 GNDA.n2137 GNDA.n2 6.688
R3492 GNDA.n1743 GNDA.n337 6.20656
R3493 GNDA.n593 GNDA.n544 6.20656
R3494 GNDA.n1714 GNDA.n375 6.20656
R3495 GNDA.n1934 GNDA.n152 6.20656
R3496 GNDA.n1094 GNDA.n1032 6.20656
R3497 GNDA.n1342 GNDA.n1280 6.20656
R3498 GNDA.t26 GNDA.t199 6.17883
R3499 GNDA.n1950 GNDA.n140 6.07727
R3500 GNDA.t76 GNDA.n2216 5.97926
R3501 GNDA.t55 GNDA.n2215 5.97926
R3502 GNDA.n2156 GNDA.t20 5.97926
R3503 GNDA.n2155 GNDA.t34 5.97926
R3504 GNDA.n2154 GNDA.t118 5.97926
R3505 GNDA.n2153 GNDA.t7 5.97926
R3506 GNDA.n2157 GNDA.t102 5.97926
R3507 GNDA.t270 GNDA.n2185 5.97926
R3508 GNDA.t304 GNDA.n2217 5.97926
R3509 GNDA.n85 GNDA.n0 5.737
R3510 GNDA.n2196 GNDA.n2194 5.6255
R3511 GNDA.n2200 GNDA.n2199 5.6255
R3512 GNDA.n2106 GNDA.n2105 5.6255
R3513 GNDA.n2102 GNDA.n2100 5.6255
R3514 GNDA.n2113 GNDA.n2112 5.60318
R3515 GNDA.n2206 GNDA.n20 5.60318
R3516 GNDA.n1950 GNDA.n1949 5.5601
R3517 GNDA.n1172 GNDA.n1146 5.51161
R3518 GNDA.n946 GNDA.n945 5.51161
R3519 GNDA.n1483 GNDA.n398 5.51161
R3520 GNDA.n1615 GNDA.n1486 5.51161
R3521 GNDA.n827 GNDA.n805 5.51161
R3522 GNDA.n1787 GNDA.n1786 5.51161
R3523 GNDA.n706 GNDA.n684 5.51161
R3524 GNDA.n1972 GNDA.n124 5.51161
R3525 GNDA.n1881 GNDA.n1880 5.51161
R3526 GNDA.n2141 GNDA.n2138 5.46925
R3527 GNDA.n2163 GNDA.n40 5.46925
R3528 GNDA.n683 GNDA.n485 5.1717
R3529 GNDA.n1525 GNDA.n1521 5.1717
R3530 GNDA.n175 GNDA.n173 5.1717
R3531 GNDA.n2084 GNDA.t199 5.14911
R3532 GNDA.t68 GNDA.t248 5.14911
R3533 GNDA.n39 GNDA.n38 5.063
R3534 GNDA.n19 GNDA.n18 5.063
R3535 GNDA.n1241 GNDA.n1119 4.9157
R3536 GNDA.n1012 GNDA.n1011 4.9157
R3537 GNDA.n1440 GNDA.n1387 4.9157
R3538 GNDA.n2163 GNDA.n2162 4.79217
R3539 GNDA.n2166 GNDA.n2165 4.79217
R3540 GNDA.n2182 GNDA.n2181 4.79217
R3541 GNDA.n2116 GNDA.n2114 4.71925
R3542 GNDA.n2221 GNDA.n3 4.71925
R3543 GNDA.n2221 GNDA.n2220 4.70883
R3544 GNDA.n2112 GNDA.n2111 4.67238
R3545 GNDA.n2206 GNDA.n2205 4.67238
R3546 GNDA.n2113 GNDA.n40 4.563
R3547 GNDA.n2136 GNDA.n2135 4.5005
R3548 GNDA.n2172 GNDA.n21 4.5005
R3549 GNDA.n2148 GNDA.n2147 4.5005
R3550 GNDA.n2178 GNDA.n2177 4.5005
R3551 GNDA.n2168 GNDA.n2167 4.5005
R3552 GNDA.n2199 GNDA.n2198 4.5005
R3553 GNDA.n2223 GNDA.n2222 4.5005
R3554 GNDA.n2105 GNDA.n2104 4.5005
R3555 GNDA.n1810 GNDA.n1807 4.26717
R3556 GNDA.n1810 GNDA.n1804 4.26717
R3557 GNDA.n1816 GNDA.n1804 4.26717
R3558 GNDA.n1817 GNDA.n1816 4.26717
R3559 GNDA.n1817 GNDA.n1800 4.26717
R3560 GNDA.n1824 GNDA.n1800 4.26717
R3561 GNDA.n1825 GNDA.n1824 4.26717
R3562 GNDA.n1825 GNDA.n1796 4.26717
R3563 GNDA.n1831 GNDA.n1796 4.26717
R3564 GNDA.n1832 GNDA.n1831 4.26717
R3565 GNDA.n1832 GNDA.n1793 4.26717
R3566 GNDA.n592 GNDA.n545 4.26717
R3567 GNDA.n587 GNDA.n545 4.26717
R3568 GNDA.n587 GNDA.n586 4.26717
R3569 GNDA.n586 GNDA.n585 4.26717
R3570 GNDA.n585 GNDA.n582 4.26717
R3571 GNDA.n582 GNDA.n581 4.26717
R3572 GNDA.n581 GNDA.n578 4.26717
R3573 GNDA.n578 GNDA.n577 4.26717
R3574 GNDA.n577 GNDA.n574 4.26717
R3575 GNDA.n574 GNDA.n573 4.26717
R3576 GNDA.n573 GNDA.n571 4.26717
R3577 GNDA.n1499 GNDA.n376 4.26717
R3578 GNDA.n1573 GNDA.n1499 4.26717
R3579 GNDA.n1574 GNDA.n1573 4.26717
R3580 GNDA.n1577 GNDA.n1574 4.26717
R3581 GNDA.n1577 GNDA.n1495 4.26717
R3582 GNDA.n1583 GNDA.n1495 4.26717
R3583 GNDA.n1584 GNDA.n1583 4.26717
R3584 GNDA.n1587 GNDA.n1584 4.26717
R3585 GNDA.n1587 GNDA.n1493 4.26717
R3586 GNDA.n1493 GNDA.n1490 4.26717
R3587 GNDA.n1594 GNDA.n1490 4.26717
R3588 GNDA.n1341 GNDA.n1281 4.26717
R3589 GNDA.n1336 GNDA.n1281 4.26717
R3590 GNDA.n1336 GNDA.n1335 4.26717
R3591 GNDA.n1335 GNDA.n1313 4.26717
R3592 GNDA.n1330 GNDA.n1313 4.26717
R3593 GNDA.n1330 GNDA.n1329 4.26717
R3594 GNDA.n1329 GNDA.n1328 4.26717
R3595 GNDA.n1328 GNDA.n1323 4.26717
R3596 GNDA.n1323 GNDA.n396 4.26717
R3597 GNDA.n1675 GNDA.n396 4.26717
R3598 GNDA.n1675 GNDA.n394 4.26717
R3599 GNDA.n1742 GNDA.n339 4.26717
R3600 GNDA.n1736 GNDA.n339 4.26717
R3601 GNDA.n1736 GNDA.n1735 4.26717
R3602 GNDA.n1735 GNDA.n1734 4.26717
R3603 GNDA.n1734 GNDA.n1732 4.26717
R3604 GNDA.n1732 GNDA.n1729 4.26717
R3605 GNDA.n1729 GNDA.n1728 4.26717
R3606 GNDA.n1728 GNDA.n1725 4.26717
R3607 GNDA.n1725 GNDA.n1724 4.26717
R3608 GNDA.n1724 GNDA.n1721 4.26717
R3609 GNDA.n1721 GNDA.n1720 4.26717
R3610 GNDA.n1093 GNDA.n1033 4.26717
R3611 GNDA.n1087 GNDA.n1033 4.26717
R3612 GNDA.n1087 GNDA.n1086 4.26717
R3613 GNDA.n1086 GNDA.n1085 4.26717
R3614 GNDA.n1085 GNDA.n1056 4.26717
R3615 GNDA.n1059 GNDA.n1056 4.26717
R3616 GNDA.n1076 GNDA.n1059 4.26717
R3617 GNDA.n1076 GNDA.n1075 4.26717
R3618 GNDA.n1075 GNDA.n1074 4.26717
R3619 GNDA.n1074 GNDA.n1064 4.26717
R3620 GNDA.n1064 GNDA.n335 4.26717
R3621 GNDA GNDA.n2224 4.2117
R3622 GNDA.n2056 GNDA.n2055 4.063
R3623 GNDA.n2149 GNDA.n2141 4.0005
R3624 GNDA.n2166 GNDA.n2163 4.0005
R3625 GNDA.n1807 GNDA.n152 3.93531
R3626 GNDA.n593 GNDA.n592 3.93531
R3627 GNDA.n1714 GNDA.n376 3.93531
R3628 GNDA.n1342 GNDA.n1341 3.93531
R3629 GNDA.n1743 GNDA.n1742 3.93531
R3630 GNDA.n1094 GNDA.n1093 3.93531
R3631 GNDA.t194 GNDA.t83 3.83994
R3632 GNDA.t41 GNDA.t258 3.83994
R3633 GNDA.t4 GNDA.t148 3.83994
R3634 GNDA.t204 GNDA.t305 3.83994
R3635 GNDA.t91 GNDA.t285 3.83994
R3636 GNDA.n1236 GNDA.n1235 3.7893
R3637 GNDA.n1232 GNDA.n1122 3.7893
R3638 GNDA.n1231 GNDA.n1125 3.7893
R3639 GNDA.n1227 GNDA.n1226 3.7893
R3640 GNDA.n1149 GNDA.n1127 3.7893
R3641 GNDA.n1157 GNDA.n1156 3.7893
R3642 GNDA.n1161 GNDA.n1160 3.7893
R3643 GNDA.n1169 GNDA.n1147 3.7893
R3644 GNDA.n1009 GNDA.n452 3.7893
R3645 GNDA.n899 GNDA.n898 3.7893
R3646 GNDA.n1003 GNDA.n1002 3.7893
R3647 GNDA.n923 GNDA.n900 3.7893
R3648 GNDA.n925 GNDA.n924 3.7893
R3649 GNDA.n931 GNDA.n920 3.7893
R3650 GNDA.n938 GNDA.n919 3.7893
R3651 GNDA.n939 GNDA.n918 3.7893
R3652 GNDA.n1469 GNDA.n425 3.7893
R3653 GNDA.n1468 GNDA.n426 3.7893
R3654 GNDA.n1447 GNDA.n1446 3.7893
R3655 GNDA.n1462 GNDA.n1461 3.7893
R3656 GNDA.n1458 GNDA.n1457 3.7893
R3657 GNDA.n1453 GNDA.n402 3.7893
R3658 GNDA.n1475 GNDA.n1474 3.7893
R3659 GNDA.n403 GNDA.n399 3.7893
R3660 GNDA.n2075 GNDA.n77 3.7893
R3661 GNDA.n2074 GNDA.n78 3.7893
R3662 GNDA.n2062 GNDA.n2061 3.7893
R3663 GNDA.n2068 GNDA.n2067 3.7893
R3664 GNDA.n2064 GNDA.n2063 3.7893
R3665 GNDA.n1602 GNDA.n56 3.7893
R3666 GNDA.n1605 GNDA.n1604 3.7893
R3667 GNDA.n1612 GNDA.n1487 3.7893
R3668 GNDA.n890 GNDA.n889 3.7893
R3669 GNDA.n886 GNDA.n780 3.7893
R3670 GNDA.n885 GNDA.n783 3.7893
R3671 GNDA.n882 GNDA.n881 3.7893
R3672 GNDA.n807 GNDA.n784 3.7893
R3673 GNDA.n816 GNDA.n815 3.7893
R3674 GNDA.n819 GNDA.n806 3.7893
R3675 GNDA.n824 GNDA.n820 3.7893
R3676 GNDA.n1749 GNDA.n272 3.7893
R3677 GNDA.n1758 GNDA.n1757 3.7893
R3678 GNDA.n270 GNDA.n269 3.7893
R3679 GNDA.n1766 GNDA.n1764 3.7893
R3680 GNDA.n1765 GNDA.n267 3.7893
R3681 GNDA.n265 GNDA.n264 3.7893
R3682 GNDA.n1781 GNDA.n1779 3.7893
R3683 GNDA.n1780 GNDA.n260 3.7893
R3684 GNDA.n769 GNDA.n768 3.7893
R3685 GNDA.n765 GNDA.n462 3.7893
R3686 GNDA.n764 GNDA.n465 3.7893
R3687 GNDA.n761 GNDA.n760 3.7893
R3688 GNDA.n686 GNDA.n466 3.7893
R3689 GNDA.n695 GNDA.n694 3.7893
R3690 GNDA.n698 GNDA.n685 3.7893
R3691 GNDA.n703 GNDA.n699 3.7893
R3692 GNDA.n2044 GNDA.n113 3.7893
R3693 GNDA.n2043 GNDA.n114 3.7893
R3694 GNDA.n2031 GNDA.n2030 3.7893
R3695 GNDA.n2037 GNDA.n2036 3.7893
R3696 GNDA.n2033 GNDA.n2032 3.7893
R3697 GNDA.n129 GNDA.n92 3.7893
R3698 GNDA.n132 GNDA.n131 3.7893
R3699 GNDA.n1969 GNDA.n125 3.7893
R3700 GNDA.n1843 GNDA.n190 3.7893
R3701 GNDA.n1852 GNDA.n1851 3.7893
R3702 GNDA.n188 GNDA.n187 3.7893
R3703 GNDA.n1860 GNDA.n1858 3.7893
R3704 GNDA.n1859 GNDA.n185 3.7893
R3705 GNDA.n183 GNDA.n182 3.7893
R3706 GNDA.n1875 GNDA.n1873 3.7893
R3707 GNDA.n1874 GNDA.n178 3.7893
R3708 GNDA.n1155 GNDA 3.7381
R3709 GNDA.n932 GNDA 3.7381
R3710 GNDA.n1454 GNDA 3.7381
R3711 GNDA GNDA.n2080 3.7381
R3712 GNDA.n812 GNDA 3.7381
R3713 GNDA GNDA.n1772 3.7381
R3714 GNDA.n691 GNDA 3.7381
R3715 GNDA GNDA.n2049 3.7381
R3716 GNDA GNDA.n1866 3.7381
R3717 GNDA.n2140 GNDA.n2139 3.55883
R3718 GNDA.n2151 GNDA.n2150 3.55883
R3719 GNDA.n2188 GNDA.n2187 3.55883
R3720 GNDA.n2191 GNDA.n2190 3.55883
R3721 GNDA.n2162 GNDA.n2161 3.55883
R3722 GNDA.n2165 GNDA.n2164 3.55883
R3723 GNDA.n2183 GNDA.n2182 3.55883
R3724 GNDA.n2180 GNDA.n2179 3.55883
R3725 GNDA.n26 GNDA.n1 3.55883
R3726 GNDA.n2220 GNDA.n2219 3.55883
R3727 GNDA.n2144 GNDA.n28 3.538
R3728 GNDA.n2176 GNDA.n2175 3.538
R3729 GNDA.n1960 GNDA.n1958 3.51962
R3730 GNDA.n2101 GNDA.t299 3.42907
R3731 GNDA.n2101 GNDA.t302 3.42907
R3732 GNDA.n2103 GNDA.t107 3.42907
R3733 GNDA.n2103 GNDA.t105 3.42907
R3734 GNDA.n2195 GNDA.t135 3.42907
R3735 GNDA.n2195 GNDA.t29 3.42907
R3736 GNDA.n2197 GNDA.t19 3.42907
R3737 GNDA.n2197 GNDA.t296 3.42907
R3738 GNDA.n136 GNDA.n121 3.16665
R3739 GNDA.n1442 GNDA.n435 3.08966
R3740 GNDA.n1466 GNDA.t130 3.08966
R3741 GNDA.n1450 GNDA.t23 3.08966
R3742 GNDA.n1480 GNDA.t22 3.08966
R3743 GNDA.n2041 GNDA.t85 3.08966
R3744 GNDA.n2138 GNDA.n2137 2.96925
R3745 GNDA.n1121 GNDA.n1119 2.6629
R3746 GNDA.n1745 GNDA.n334 2.6629
R3747 GNDA.n1011 GNDA.n1010 2.6629
R3748 GNDA.n944 GNDA.n366 2.6629
R3749 GNDA.n1440 GNDA.n1439 2.6629
R3750 GNDA.n1485 GNDA.n1484 2.6629
R3751 GNDA.n1668 GNDA.n1667 2.6629
R3752 GNDA.n1597 GNDA.n123 2.6629
R3753 GNDA.n779 GNDA.n778 2.6629
R3754 GNDA.n804 GNDA.n374 2.6629
R3755 GNDA.n1750 GNDA.n1748 2.6629
R3756 GNDA.n258 GNDA.n252 2.6629
R3757 GNDA.n461 GNDA.n460 2.6629
R3758 GNDA.n2025 GNDA.n2024 2.6629
R3759 GNDA.n1844 GNDA.n1842 2.6629
R3760 GNDA.n1146 GNDA.n334 2.4581
R3761 GNDA.n945 GNDA.n944 2.4581
R3762 GNDA.n1484 GNDA.n1483 2.4581
R3763 GNDA.n1668 GNDA.n1485 2.4581
R3764 GNDA.n1597 GNDA.n1486 2.4581
R3765 GNDA.n778 GNDA.n366 2.4581
R3766 GNDA.n805 GNDA.n804 2.4581
R3767 GNDA.n1748 GNDA.n1745 2.4581
R3768 GNDA.n1787 GNDA.n258 2.4581
R3769 GNDA.n460 GNDA.n374 2.4581
R3770 GNDA.n684 GNDA.n683 2.4581
R3771 GNDA.n2025 GNDA.n123 2.4581
R3772 GNDA.n1521 GNDA.n124 2.4581
R3773 GNDA.n1842 GNDA.n252 2.4581
R3774 GNDA.n1881 GNDA.n175 2.4581
R3775 GNDA.n2135 GNDA.n2094 2.19633
R3776 GNDA.n2114 GNDA.n4 2.19633
R3777 GNDA.n2147 GNDA.n2146 2.19633
R3778 GNDA.n2173 GNDA.n2172 2.19633
R3779 GNDA.n2169 GNDA.n2168 2.19633
R3780 GNDA.n2177 GNDA.n25 2.19633
R3781 GNDA.n1793 GNDA.n252 2.18124
R3782 GNDA.n571 GNDA.n374 2.18124
R3783 GNDA.n1594 GNDA.n123 2.18124
R3784 GNDA.n1485 GNDA.n394 2.18124
R3785 GNDA.n1720 GNDA.n366 2.18124
R3786 GNDA.n1745 GNDA.n335 2.18124
R3787 GNDA.n1168 GNDA.n1146 2.1509
R3788 GNDA.n945 GNDA.n942 2.1509
R3789 GNDA.n1483 GNDA.n1482 2.1509
R3790 GNDA.n1611 GNDA.n1486 2.1509
R3791 GNDA.n823 GNDA.n805 2.1509
R3792 GNDA.n1788 GNDA.n1787 2.1509
R3793 GNDA.n702 GNDA.n684 2.1509
R3794 GNDA.n1968 GNDA.n124 2.1509
R3795 GNDA.n1882 GNDA.n1881 2.1509
R3796 GNDA.n1208 GNDA.n1121 2.13383
R3797 GNDA.n1010 GNDA.n451 2.13383
R3798 GNDA.n1439 GNDA.n1438 2.13383
R3799 GNDA.n1667 GNDA.n1666 2.13383
R3800 GNDA.n863 GNDA.n779 2.13383
R3801 GNDA.n1751 GNDA.n1750 2.13383
R3802 GNDA.n742 GNDA.n461 2.13383
R3803 GNDA.n2024 GNDA.n2023 2.13383
R3804 GNDA.n1845 GNDA.n1844 2.13383
R3805 GNDA.n86 GNDA 2.09787
R3806 GNDA.n254 GNDA.n252 2.08643
R3807 GNDA.n1715 GNDA.n374 2.08643
R3808 GNDA.n1489 GNDA.n123 2.08643
R3809 GNDA.n1485 GNDA.n393 2.08643
R3810 GNDA.n368 GNDA.n366 2.08643
R3811 GNDA.n1745 GNDA.n1744 2.08643
R3812 GNDA.n2194 GNDA.n2193 2.07331
R3813 GNDA.n2201 GNDA.n2200 2.07331
R3814 GNDA.n2107 GNDA.n2106 2.07331
R3815 GNDA.n2100 GNDA.n2099 2.07331
R3816 GNDA.n1480 GNDA.t252 2.05994
R3817 GNDA.n1669 GNDA.t273 2.05994
R3818 GNDA.n1599 GNDA.t231 2.05994
R3819 GNDA.t248 GNDA.n2028 2.05994
R3820 GNDA.n1236 GNDA.n1121 1.9461
R3821 GNDA.n1010 GNDA.n1009 1.9461
R3822 GNDA.n1439 GNDA.n425 1.9461
R3823 GNDA.n1667 GNDA.n77 1.9461
R3824 GNDA.n890 GNDA.n779 1.9461
R3825 GNDA.n1750 GNDA.n1749 1.9461
R3826 GNDA.n769 GNDA.n461 1.9461
R3827 GNDA.n2024 GNDA.n113 1.9461
R3828 GNDA.n1844 GNDA.n1843 1.9461
R3829 GNDA.n2222 GNDA.n2221 1.938
R3830 GNDA.n2111 GNDA.n2110 1.913
R3831 GNDA.n2096 GNDA.n2095 1.913
R3832 GNDA.n2205 GNDA.n2204 1.913
R3833 GNDA.n2208 GNDA.n2207 1.913
R3834 GNDA.n1957 GNDA.n1956 1.90675
R3835 GNDA.n1015 GNDA.t151 1.83728
R3836 GNDA.n2156 GNDA.t124 1.54702
R3837 GNDA.n2155 GNDA.t112 1.54702
R3838 GNDA.n2154 GNDA.t56 1.54702
R3839 GNDA.n2153 GNDA.t110 1.54702
R3840 GNDA.n2216 GNDA.t58 1.54702
R3841 GNDA.n2215 GNDA.t224 1.54702
R3842 GNDA.n2157 GNDA.t212 1.54702
R3843 GNDA.n2185 GNDA.t136 1.54702
R3844 GNDA.n2217 GNDA.t141 1.54702
R3845 GNDA.n1244 GNDA.n1241 1.47392
R3846 GNDA.n1012 GNDA.n450 1.47392
R3847 GNDA.n1387 GNDA.n437 1.47392
R3848 GNDA.n673 GNDA.n485 1.47392
R3849 GNDA.n1526 GNDA.n1525 1.47392
R3850 GNDA.n1892 GNDA.n173 1.47392
R3851 GNDA.n2199 GNDA.n2196 1.1255
R3852 GNDA.n2105 GNDA.n2102 1.1255
R3853 GNDA.n1696 GNDA.n1693 0.96925
R3854 GNDA.n1705 GNDA.n1684 0.96925
R3855 GNDA.n2138 GNDA.n2113 0.922375
R3856 GNDA.n83 GNDA.n82 0.914368
R3857 GNDA.n2189 GNDA.n21 0.8755
R3858 GNDA.n2149 GNDA.n2148 0.8755
R3859 GNDA.n2181 GNDA.n2178 0.8755
R3860 GNDA.n2167 GNDA.n2166 0.8755
R3861 GNDA.n1235 GNDA.n1122 0.8197
R3862 GNDA.n1232 GNDA.n1231 0.8197
R3863 GNDA.n1227 GNDA.n1125 0.8197
R3864 GNDA.n1226 GNDA.n1127 0.8197
R3865 GNDA.n1156 GNDA.n1155 0.8197
R3866 GNDA.n1161 GNDA.n1157 0.8197
R3867 GNDA.n1160 GNDA.n1147 0.8197
R3868 GNDA.n1169 GNDA.n1168 0.8197
R3869 GNDA.n898 GNDA.n452 0.8197
R3870 GNDA.n1003 GNDA.n899 0.8197
R3871 GNDA.n1002 GNDA.n900 0.8197
R3872 GNDA.n925 GNDA.n923 0.8197
R3873 GNDA.n932 GNDA.n931 0.8197
R3874 GNDA.n920 GNDA.n919 0.8197
R3875 GNDA.n939 GNDA.n938 0.8197
R3876 GNDA.n942 GNDA.n918 0.8197
R3877 GNDA.n1469 GNDA.n1468 0.8197
R3878 GNDA.n1446 GNDA.n426 0.8197
R3879 GNDA.n1462 GNDA.n1447 0.8197
R3880 GNDA.n1461 GNDA.n1458 0.8197
R3881 GNDA.n1454 GNDA.n1453 0.8197
R3882 GNDA.n1475 GNDA.n402 0.8197
R3883 GNDA.n1474 GNDA.n403 0.8197
R3884 GNDA.n1482 GNDA.n399 0.8197
R3885 GNDA.n2075 GNDA.n2074 0.8197
R3886 GNDA.n2061 GNDA.n78 0.8197
R3887 GNDA.n2068 GNDA.n2062 0.8197
R3888 GNDA.n2067 GNDA.n2064 0.8197
R3889 GNDA.n2080 GNDA.n56 0.8197
R3890 GNDA.n1605 GNDA.n1602 0.8197
R3891 GNDA.n1604 GNDA.n1487 0.8197
R3892 GNDA.n1612 GNDA.n1611 0.8197
R3893 GNDA.n889 GNDA.n780 0.8197
R3894 GNDA.n886 GNDA.n885 0.8197
R3895 GNDA.n882 GNDA.n783 0.8197
R3896 GNDA.n881 GNDA.n784 0.8197
R3897 GNDA.n815 GNDA.n812 0.8197
R3898 GNDA.n816 GNDA.n806 0.8197
R3899 GNDA.n820 GNDA.n819 0.8197
R3900 GNDA.n824 GNDA.n823 0.8197
R3901 GNDA.n1758 GNDA.n272 0.8197
R3902 GNDA.n1757 GNDA.n270 0.8197
R3903 GNDA.n1764 GNDA.n269 0.8197
R3904 GNDA.n1766 GNDA.n1765 0.8197
R3905 GNDA.n1772 GNDA.n265 0.8197
R3906 GNDA.n1779 GNDA.n264 0.8197
R3907 GNDA.n1781 GNDA.n1780 0.8197
R3908 GNDA.n1788 GNDA.n260 0.8197
R3909 GNDA.n768 GNDA.n462 0.8197
R3910 GNDA.n765 GNDA.n764 0.8197
R3911 GNDA.n761 GNDA.n465 0.8197
R3912 GNDA.n760 GNDA.n466 0.8197
R3913 GNDA.n694 GNDA.n691 0.8197
R3914 GNDA.n695 GNDA.n685 0.8197
R3915 GNDA.n699 GNDA.n698 0.8197
R3916 GNDA.n703 GNDA.n702 0.8197
R3917 GNDA.n2044 GNDA.n2043 0.8197
R3918 GNDA.n2030 GNDA.n114 0.8197
R3919 GNDA.n2037 GNDA.n2031 0.8197
R3920 GNDA.n2036 GNDA.n2033 0.8197
R3921 GNDA.n2049 GNDA.n92 0.8197
R3922 GNDA.n132 GNDA.n129 0.8197
R3923 GNDA.n131 GNDA.n125 0.8197
R3924 GNDA.n1969 GNDA.n1968 0.8197
R3925 GNDA.n1852 GNDA.n190 0.8197
R3926 GNDA.n1851 GNDA.n188 0.8197
R3927 GNDA.n1858 GNDA.n187 0.8197
R3928 GNDA.n1860 GNDA.n1859 0.8197
R3929 GNDA.n1866 GNDA.n183 0.8197
R3930 GNDA.n1873 GNDA.n182 0.8197
R3931 GNDA.n1875 GNDA.n1874 0.8197
R3932 GNDA.n1882 GNDA.n178 0.8197
R3933 GNDA.n1264 GNDA.n1015 0.575776
R3934 GNDA GNDA.n1149 0.5637
R3935 GNDA.n924 GNDA 0.5637
R3936 GNDA.n1457 GNDA 0.5637
R3937 GNDA.n2063 GNDA 0.5637
R3938 GNDA GNDA.n807 0.5637
R3939 GNDA.n267 GNDA 0.5637
R3940 GNDA GNDA.n686 0.5637
R3941 GNDA.n2032 GNDA 0.5637
R3942 GNDA.n185 GNDA 0.5637
R3943 GNDA.n1961 GNDA.n138 0.563
R3944 GNDA.n1686 GNDA.n138 0.563
R3945 GNDA.n1688 GNDA.n1686 0.563
R3946 GNDA.n1693 GNDA.n1688 0.563
R3947 GNDA.n1698 GNDA.n1696 0.563
R3948 GNDA.n1700 GNDA.n1698 0.563
R3949 GNDA.n1702 GNDA.n1700 0.563
R3950 GNDA.n1704 GNDA.n1702 0.563
R3951 GNDA.n1705 GNDA.n1704 0.563
R3952 GNDA.n1684 GNDA.n391 0.563
R3953 GNDA.n430 GNDA.n391 0.563
R3954 GNDA.n432 GNDA.n430 0.563
R3955 GNDA.n2118 GNDA.n2116 0.563
R3956 GNDA.n2120 GNDA.n2118 0.563
R3957 GNDA.n2122 GNDA.n2120 0.563
R3958 GNDA.n2124 GNDA.n2122 0.563
R3959 GNDA.n2126 GNDA.n2124 0.563
R3960 GNDA.n2128 GNDA.n2126 0.563
R3961 GNDA.n2130 GNDA.n2128 0.563
R3962 GNDA.n2132 GNDA.n2130 0.563
R3963 GNDA.n2134 GNDA.n2132 0.563
R3964 GNDA.n2136 GNDA.n2134 0.563
R3965 GNDA.n2143 GNDA.n21 0.563
R3966 GNDA.n2148 GNDA.n2143 0.563
R3967 GNDA.n2178 GNDA.n24 0.563
R3968 GNDA.n2167 GNDA.n24 0.563
R3969 GNDA.n34 GNDA.n32 0.563
R3970 GNDA.n36 GNDA.n34 0.563
R3971 GNDA.n38 GNDA.n36 0.563
R3972 GNDA.n14 GNDA.n12 0.563
R3973 GNDA.n16 GNDA.n14 0.563
R3974 GNDA.n18 GNDA.n16 0.563
R3975 GNDA.n2168 GNDA.n28 0.5005
R3976 GNDA.n2177 GNDA.n2176 0.5005
R3977 GNDA.n1959 GNDA.n86 0.276625
R3978 GNDA.n1153 GNDA 0.2565
R3979 GNDA.n928 GNDA 0.2565
R3980 GNDA.n1452 GNDA 0.2565
R3981 GNDA.n2081 GNDA 0.2565
R3982 GNDA.n810 GNDA 0.2565
R3983 GNDA.n1773 GNDA 0.2565
R3984 GNDA.n689 GNDA 0.2565
R3985 GNDA.n2050 GNDA 0.2565
R3986 GNDA.n1867 GNDA 0.2565
R3987 GNDA.n1960 GNDA.n1959 0.22375
R3988 GNDA.n2223 GNDA.n1 0.208833
R3989 GNDA GNDA.n1153 0.0517
R3990 GNDA GNDA.n928 0.0517
R3991 GNDA GNDA.n1452 0.0517
R3992 GNDA.n2081 GNDA 0.0517
R3993 GNDA GNDA.n810 0.0517
R3994 GNDA.n1773 GNDA 0.0517
R3995 GNDA GNDA.n689 0.0517
R3996 GNDA.n2050 GNDA 0.0517
R3997 GNDA.n1867 GNDA 0.0517
R3998 VDDA.n103 VDDA.t274 1221.7
R3999 VDDA.n106 VDDA.t256 1221.7
R4000 VDDA.n39 VDDA.t327 1221.7
R4001 VDDA.n42 VDDA.t339 1221.7
R4002 VDDA.n51 VDDA.t303 755.768
R4003 VDDA.n55 VDDA.t312 755.768
R4004 VDDA.n48 VDDA.t271 755.768
R4005 VDDA.n60 VDDA.t351 755.768
R4006 VDDA.n71 VDDA.t300 698.095
R4007 VDDA.n5 VDDA.t315 698.095
R4008 VDDA.n188 VDDA.t355 683.365
R4009 VDDA.n119 VDDA.t297 661.375
R4010 VDDA.n122 VDDA.t345 661.375
R4011 VDDA.n69 VDDA.t244 661.375
R4012 VDDA.n7 VDDA.t259 661.375
R4013 VDDA.t322 VDDA.n179 660
R4014 VDDA.n180 VDDA.t295 660
R4015 VDDA.t263 VDDA.n157 660
R4016 VDDA.n158 VDDA.t284 660
R4017 VDDA.t319 VDDA.n187 643.037
R4018 VDDA.t266 VDDA.n253 643.037
R4019 VDDA.n254 VDDA.t334 643.037
R4020 VDDA.t331 VDDA.n236 643.037
R4021 VDDA.n237 VDDA.t248 643.037
R4022 VDDA.t307 VDDA.n228 643.037
R4023 VDDA.n229 VDDA.t343 643.037
R4024 VDDA.n212 VDDA.t336 611.909
R4025 VDDA.n222 VDDA.t348 601.867
R4026 VDDA.n247 VDDA.t286 601.867
R4027 VDDA.n89 VDDA.t324 581.436
R4028 VDDA.n25 VDDA.t253 581.436
R4029 VDDA.n210 VDDA.t250 579.775
R4030 VDDA.n91 VDDA.t309 579.034
R4031 VDDA.n27 VDDA.t268 579.034
R4032 VDDA.t278 VDDA.t279 565.923
R4033 VDDA.n115 VDDA.t277 461.026
R4034 VDDA.n112 VDDA.t290 456.526
R4035 VDDA.n186 VDDA.t318 413.084
R4036 VDDA.n189 VDDA.t354 413.084
R4037 VDDA.n252 VDDA.t265 409.067
R4038 VDDA.n255 VDDA.t333 409.067
R4039 VDDA.n235 VDDA.t330 409.067
R4040 VDDA.n227 VDDA.t306 409.067
R4041 VDDA.n230 VDDA.t342 409.067
R4042 VDDA.t76 VDDA.t322 407.144
R4043 VDDA.t378 VDDA.t76 407.144
R4044 VDDA.t90 VDDA.t378 407.144
R4045 VDDA.t0 VDDA.t90 407.144
R4046 VDDA.t94 VDDA.t0 407.144
R4047 VDDA.t119 VDDA.t94 407.144
R4048 VDDA.t402 VDDA.t119 407.144
R4049 VDDA.t161 VDDA.t402 407.144
R4050 VDDA.t72 VDDA.t161 407.144
R4051 VDDA.t367 VDDA.t72 407.144
R4052 VDDA.t2 VDDA.t367 407.144
R4053 VDDA.t153 VDDA.t2 407.144
R4054 VDDA.t390 VDDA.t153 407.144
R4055 VDDA.t185 VDDA.t390 407.144
R4056 VDDA.t191 VDDA.t185 407.144
R4057 VDDA.t128 VDDA.t191 407.144
R4058 VDDA.t140 VDDA.t128 407.144
R4059 VDDA.t151 VDDA.t140 407.144
R4060 VDDA.t295 VDDA.t151 407.144
R4061 VDDA.t133 VDDA.t263 407.144
R4062 VDDA.t172 VDDA.t133 407.144
R4063 VDDA.t9 VDDA.t172 407.144
R4064 VDDA.t131 VDDA.t9 407.144
R4065 VDDA.t382 VDDA.t131 407.144
R4066 VDDA.t88 VDDA.t382 407.144
R4067 VDDA.t105 VDDA.t88 407.144
R4068 VDDA.t126 VDDA.t105 407.144
R4069 VDDA.t147 VDDA.t126 407.144
R4070 VDDA.t145 VDDA.t147 407.144
R4071 VDDA.t59 VDDA.t145 407.144
R4072 VDDA.t149 VDDA.t59 407.144
R4073 VDDA.t174 VDDA.t149 407.144
R4074 VDDA.t400 VDDA.t174 407.144
R4075 VDDA.t388 VDDA.t400 407.144
R4076 VDDA.t380 VDDA.t388 407.144
R4077 VDDA.t57 VDDA.t380 407.144
R4078 VDDA.t396 VDDA.t57 407.144
R4079 VDDA.t284 VDDA.t396 407.144
R4080 VDDA.n111 VDDA.t291 397.784
R4081 VDDA.n238 VDDA.t247 390.322
R4082 VDDA.t19 VDDA.t319 373.214
R4083 VDDA.t386 VDDA.t19 373.214
R4084 VDDA.t355 VDDA.t386 373.214
R4085 VDDA.t163 VDDA.t266 373.214
R4086 VDDA.t363 VDDA.t163 373.214
R4087 VDDA.t193 VDDA.t363 373.214
R4088 VDDA.t6 VDDA.t193 373.214
R4089 VDDA.t334 VDDA.t6 373.214
R4090 VDDA.t99 VDDA.t331 373.214
R4091 VDDA.t74 VDDA.t99 373.214
R4092 VDDA.t408 VDDA.t74 373.214
R4093 VDDA.t41 VDDA.t408 373.214
R4094 VDDA.t248 VDDA.t41 373.214
R4095 VDDA.t365 VDDA.t307 373.214
R4096 VDDA.t79 VDDA.t365 373.214
R4097 VDDA.t343 VDDA.t79 373.214
R4098 VDDA.n208 VDDA.t241 360.868
R4099 VDDA.n191 VDDA.t280 360.868
R4100 VDDA.n159 VDDA.t283 358.858
R4101 VDDA.n137 VDDA.n136 347.104
R4102 VDDA.n162 VDDA.n161 347.104
R4103 VDDA.n164 VDDA.n163 347.104
R4104 VDDA.n166 VDDA.n165 347.104
R4105 VDDA.n168 VDDA.n167 347.104
R4106 VDDA.n170 VDDA.n169 347.104
R4107 VDDA.n172 VDDA.n171 347.104
R4108 VDDA.n174 VDDA.n173 347.104
R4109 VDDA.n176 VDDA.n175 347.104
R4110 VDDA.n139 VDDA.n138 347.104
R4111 VDDA.n141 VDDA.n140 347.104
R4112 VDDA.n143 VDDA.n142 347.104
R4113 VDDA.n145 VDDA.n144 347.104
R4114 VDDA.n147 VDDA.n146 347.104
R4115 VDDA.n149 VDDA.n148 347.104
R4116 VDDA.n151 VDDA.n150 347.104
R4117 VDDA.n153 VDDA.n152 347.104
R4118 VDDA.n155 VDDA.n154 347.104
R4119 VDDA.n224 VDDA.n223 345.127
R4120 VDDA.n233 VDDA.n232 345.127
R4121 VDDA.n226 VDDA.n225 345.127
R4122 VDDA.n219 VDDA.n218 344.7
R4123 VDDA.n250 VDDA.n249 344.7
R4124 VDDA.n90 VDDA.t310 343.882
R4125 VDDA.t325 VDDA.n89 343.882
R4126 VDDA.t254 VDDA.n25 343.882
R4127 VDDA.n26 VDDA.t269 343.882
R4128 VDDA.n213 VDDA.t337 341.188
R4129 VDDA.t251 VDDA.n211 341.188
R4130 VDDA.t349 VDDA.n245 341.188
R4131 VDDA.n246 VDDA.t287 341.188
R4132 VDDA.n236 VDDA.t332 332.267
R4133 VDDA.n237 VDDA.t249 332.267
R4134 VDDA.n228 VDDA.t308 332.267
R4135 VDDA.n229 VDDA.t344 332.267
R4136 VDDA.n253 VDDA.t267 332.084
R4137 VDDA.n254 VDDA.t335 332.084
R4138 VDDA.n179 VDDA.t323 331.901
R4139 VDDA.n180 VDDA.t296 331.901
R4140 VDDA.n157 VDDA.t264 331.901
R4141 VDDA.n158 VDDA.t285 331.901
R4142 VDDA.n187 VDDA.t320 331.901
R4143 VDDA.n188 VDDA.t356 331.901
R4144 VDDA.n59 VDDA.t352 284.921
R4145 VDDA.n50 VDDA.t304 284.921
R4146 VDDA.t242 VDDA.n184 280.798
R4147 VDDA.n185 VDDA.t281 280.798
R4148 VDDA.t398 VDDA.t278 259.091
R4149 VDDA.t291 VDDA.t398 259.091
R4150 VDDA.t281 VDDA.t159 240.845
R4151 VDDA.t159 VDDA.t392 240.845
R4152 VDDA.t392 VDDA.t61 240.845
R4153 VDDA.t61 VDDA.t44 240.845
R4154 VDDA.t44 VDDA.t122 240.845
R4155 VDDA.t122 VDDA.t179 240.845
R4156 VDDA.t179 VDDA.t155 240.845
R4157 VDDA.t155 VDDA.t81 240.845
R4158 VDDA.t81 VDDA.t124 240.845
R4159 VDDA.t124 VDDA.t157 240.845
R4160 VDDA.t157 VDDA.t83 240.845
R4161 VDDA.t83 VDDA.t85 240.845
R4162 VDDA.t85 VDDA.t25 240.845
R4163 VDDA.t25 VDDA.t404 240.845
R4164 VDDA.t404 VDDA.t176 240.845
R4165 VDDA.t176 VDDA.t107 240.845
R4166 VDDA.t107 VDDA.t242 240.845
R4167 VDDA.t272 VDDA.n58 221.121
R4168 VDDA.n58 VDDA.t313 221.121
R4169 VDDA.t310 VDDA.t92 217.708
R4170 VDDA.t92 VDDA.t31 217.708
R4171 VDDA.t31 VDDA.t117 217.708
R4172 VDDA.t117 VDDA.t8 217.708
R4173 VDDA.t8 VDDA.t37 217.708
R4174 VDDA.t37 VDDA.t190 217.708
R4175 VDDA.t190 VDDA.t32 217.708
R4176 VDDA.t32 VDDA.t50 217.708
R4177 VDDA.t50 VDDA.t51 217.708
R4178 VDDA.t51 VDDA.t184 217.708
R4179 VDDA.t184 VDDA.t325 217.708
R4180 VDDA.t98 VDDA.t254 217.708
R4181 VDDA.t170 VDDA.t98 217.708
R4182 VDDA.t130 VDDA.t170 217.708
R4183 VDDA.t102 VDDA.t130 217.708
R4184 VDDA.t65 VDDA.t102 217.708
R4185 VDDA.t411 VDDA.t65 217.708
R4186 VDDA.t11 VDDA.t411 217.708
R4187 VDDA.t369 VDDA.t11 217.708
R4188 VDDA.t410 VDDA.t369 217.708
R4189 VDDA.t38 VDDA.t410 217.708
R4190 VDDA.t269 VDDA.t38 217.708
R4191 VDDA.t337 VDDA.t20 217.708
R4192 VDDA.t20 VDDA.t251 217.708
R4193 VDDA.t361 VDDA.t349 217.708
R4194 VDDA.t142 VDDA.t361 217.708
R4195 VDDA.t357 VDDA.t142 217.708
R4196 VDDA.t359 VDDA.t357 217.708
R4197 VDDA.t287 VDDA.t359 217.708
R4198 VDDA.t298 VDDA.n120 213.131
R4199 VDDA.n121 VDDA.t346 213.131
R4200 VDDA.t245 VDDA.n70 213.131
R4201 VDDA.n6 VDDA.t260 213.131
R4202 VDDA.n71 VDDA.t301 211.625
R4203 VDDA.t316 VDDA.n5 211.625
R4204 VDDA.n221 VDDA.n220 190.534
R4205 VDDA.n242 VDDA.n241 190.534
R4206 VDDA.n244 VDDA.n243 190.534
R4207 VDDA.n215 VDDA.n214 186.034
R4208 VDDA.t352 VDDA.t48 180.173
R4209 VDDA.t48 VDDA.t12 180.173
R4210 VDDA.t12 VDDA.t55 180.173
R4211 VDDA.t55 VDDA.t35 180.173
R4212 VDDA.t35 VDDA.t272 180.173
R4213 VDDA.t47 VDDA.t313 180.173
R4214 VDDA.t14 VDDA.t47 180.173
R4215 VDDA.t103 VDDA.t14 180.173
R4216 VDDA.t36 VDDA.t103 180.173
R4217 VDDA.t304 VDDA.t36 180.173
R4218 VDDA.n178 VDDA.t321 179.43
R4219 VDDA.n156 VDDA.t262 179.43
R4220 VDDA.n181 VDDA.t294 179.358
R4221 VDDA.n132 VDDA.t413 169.55
R4222 VDDA.n111 VDDA.t293 168.139
R4223 VDDA.n134 VDDA.t412 165.8
R4224 VDDA.n133 VDDA.t414 165.8
R4225 VDDA.n132 VDDA.t415 165.8
R4226 VDDA.n114 VDDA.n113 153.576
R4227 VDDA.n193 VDDA.n192 147.792
R4228 VDDA.n195 VDDA.n194 147.792
R4229 VDDA.n197 VDDA.n196 147.792
R4230 VDDA.n199 VDDA.n198 147.792
R4231 VDDA.n201 VDDA.n200 147.792
R4232 VDDA.n203 VDDA.n202 147.792
R4233 VDDA.n205 VDDA.n204 147.792
R4234 VDDA.n207 VDDA.n206 147.792
R4235 VDDA.t227 VDDA.t298 146.155
R4236 VDDA.t346 VDDA.t227 146.155
R4237 VDDA.t205 VDDA.t245 146.155
R4238 VDDA.t215 VDDA.t205 146.155
R4239 VDDA.t223 VDDA.t215 146.155
R4240 VDDA.t231 VDDA.t223 146.155
R4241 VDDA.t235 VDDA.t231 146.155
R4242 VDDA.t199 VDDA.t235 146.155
R4243 VDDA.t209 VDDA.t199 146.155
R4244 VDDA.t217 VDDA.t209 146.155
R4245 VDDA.t213 VDDA.t217 146.155
R4246 VDDA.t221 VDDA.t213 146.155
R4247 VDDA.t301 VDDA.t221 146.155
R4248 VDDA.t229 VDDA.t316 146.155
R4249 VDDA.t233 VDDA.t229 146.155
R4250 VDDA.t197 VDDA.t233 146.155
R4251 VDDA.t207 VDDA.t197 146.155
R4252 VDDA.t203 VDDA.t207 146.155
R4253 VDDA.t211 VDDA.t203 146.155
R4254 VDDA.t219 VDDA.t211 146.155
R4255 VDDA.t225 VDDA.t219 146.155
R4256 VDDA.t201 VDDA.t225 146.155
R4257 VDDA.t195 VDDA.t201 146.155
R4258 VDDA.t260 VDDA.t195 146.155
R4259 VDDA.n90 VDDA.t311 136.701
R4260 VDDA.n89 VDDA.t326 136.701
R4261 VDDA.n25 VDDA.t255 136.701
R4262 VDDA.n26 VDDA.t270 136.701
R4263 VDDA.t338 VDDA.n213 136.701
R4264 VDDA.n211 VDDA.t252 136.701
R4265 VDDA.n245 VDDA.t350 136.701
R4266 VDDA.n246 VDDA.t289 136.701
R4267 VDDA.n105 VDDA.t257 122.829
R4268 VDDA.t275 VDDA.n104 122.829
R4269 VDDA.t328 VDDA.n40 122.829
R4270 VDDA.n41 VDDA.t340 122.829
R4271 VDDA.n56 VDDA.t314 113.26
R4272 VDDA.n47 VDDA.t273 113.26
R4273 VDDA.n59 VDDA.t353 113.26
R4274 VDDA.n50 VDDA.t305 113.26
R4275 VDDA.n46 VDDA.n45 104.322
R4276 VDDA.n53 VDDA.n52 104.322
R4277 VDDA.n193 VDDA.n191 99.2005
R4278 VDDA.n208 VDDA.n207 99.2005
R4279 VDDA.n195 VDDA.n193 96.0005
R4280 VDDA.n197 VDDA.n195 96.0005
R4281 VDDA.n199 VDDA.n197 96.0005
R4282 VDDA.n201 VDDA.n199 96.0005
R4283 VDDA.n203 VDDA.n201 96.0005
R4284 VDDA.n205 VDDA.n203 96.0005
R4285 VDDA.n207 VDDA.n205 96.0005
R4286 VDDA.n185 VDDA.t282 86.2588
R4287 VDDA.n184 VDDA.t243 86.2588
R4288 VDDA.t257 VDDA.t112 81.6411
R4289 VDDA.t112 VDDA.t187 81.6411
R4290 VDDA.t187 VDDA.t136 81.6411
R4291 VDDA.t136 VDDA.t4 81.6411
R4292 VDDA.t4 VDDA.t110 81.6411
R4293 VDDA.t110 VDDA.t165 81.6411
R4294 VDDA.t165 VDDA.t384 81.6411
R4295 VDDA.t384 VDDA.t33 81.6411
R4296 VDDA.t33 VDDA.t29 81.6411
R4297 VDDA.t29 VDDA.t52 81.6411
R4298 VDDA.t52 VDDA.t275 81.6411
R4299 VDDA.t376 VDDA.t328 81.6411
R4300 VDDA.t70 VDDA.t376 81.6411
R4301 VDDA.t372 VDDA.t70 81.6411
R4302 VDDA.t68 VDDA.t372 81.6411
R4303 VDDA.t370 VDDA.t68 81.6411
R4304 VDDA.t114 VDDA.t370 81.6411
R4305 VDDA.t96 VDDA.t114 81.6411
R4306 VDDA.t17 VDDA.t96 81.6411
R4307 VDDA.t374 VDDA.t17 81.6411
R4308 VDDA.t167 VDDA.t374 81.6411
R4309 VDDA.t340 VDDA.t167 81.6411
R4310 VDDA.n120 VDDA.t299 76.2576
R4311 VDDA.n121 VDDA.t347 76.2576
R4312 VDDA.n70 VDDA.t246 76.2576
R4313 VDDA.n71 VDDA.t302 76.2576
R4314 VDDA.n5 VDDA.t317 76.2576
R4315 VDDA.n6 VDDA.t261 76.2576
R4316 VDDA.n118 VDDA.n117 71.388
R4317 VDDA.n66 VDDA.n65 71.388
R4318 VDDA.n68 VDDA.n67 71.388
R4319 VDDA.n73 VDDA.n72 71.388
R4320 VDDA.n75 VDDA.n74 71.388
R4321 VDDA.n2 VDDA.n1 71.388
R4322 VDDA.n4 VDDA.n3 71.388
R4323 VDDA.n9 VDDA.n8 71.388
R4324 VDDA.n11 VDDA.n10 71.388
R4325 VDDA.n77 VDDA.n64 66.888
R4326 VDDA.n13 VDDA.n0 66.888
R4327 VDDA.n58 VDDA.n57 61.6672
R4328 VDDA.n105 VDDA.t258 40.9789
R4329 VDDA.n104 VDDA.t276 40.9789
R4330 VDDA.n40 VDDA.t329 40.9789
R4331 VDDA.n41 VDDA.t341 40.9789
R4332 VDDA.n94 VDDA.n93 40.8685
R4333 VDDA.n96 VDDA.n95 40.8685
R4334 VDDA.n98 VDDA.n97 40.8685
R4335 VDDA.n100 VDDA.n99 40.8685
R4336 VDDA.n102 VDDA.n101 40.8685
R4337 VDDA.n30 VDDA.n29 40.8685
R4338 VDDA.n32 VDDA.n31 40.8685
R4339 VDDA.n34 VDDA.n33 40.8685
R4340 VDDA.n36 VDDA.n35 40.8685
R4341 VDDA.n38 VDDA.n37 40.8685
R4342 VDDA.n136 VDDA.t141 39.4005
R4343 VDDA.n136 VDDA.t152 39.4005
R4344 VDDA.n161 VDDA.t192 39.4005
R4345 VDDA.n161 VDDA.t129 39.4005
R4346 VDDA.n163 VDDA.t391 39.4005
R4347 VDDA.n163 VDDA.t186 39.4005
R4348 VDDA.n165 VDDA.t3 39.4005
R4349 VDDA.n165 VDDA.t154 39.4005
R4350 VDDA.n167 VDDA.t73 39.4005
R4351 VDDA.n167 VDDA.t368 39.4005
R4352 VDDA.n169 VDDA.t403 39.4005
R4353 VDDA.n169 VDDA.t162 39.4005
R4354 VDDA.n171 VDDA.t95 39.4005
R4355 VDDA.n171 VDDA.t120 39.4005
R4356 VDDA.n173 VDDA.t91 39.4005
R4357 VDDA.n173 VDDA.t1 39.4005
R4358 VDDA.n175 VDDA.t77 39.4005
R4359 VDDA.n175 VDDA.t379 39.4005
R4360 VDDA.n138 VDDA.t58 39.4005
R4361 VDDA.n138 VDDA.t397 39.4005
R4362 VDDA.n140 VDDA.t389 39.4005
R4363 VDDA.n140 VDDA.t381 39.4005
R4364 VDDA.n142 VDDA.t175 39.4005
R4365 VDDA.n142 VDDA.t401 39.4005
R4366 VDDA.n144 VDDA.t60 39.4005
R4367 VDDA.n144 VDDA.t150 39.4005
R4368 VDDA.n146 VDDA.t148 39.4005
R4369 VDDA.n146 VDDA.t146 39.4005
R4370 VDDA.n148 VDDA.t106 39.4005
R4371 VDDA.n148 VDDA.t127 39.4005
R4372 VDDA.n150 VDDA.t383 39.4005
R4373 VDDA.n150 VDDA.t89 39.4005
R4374 VDDA.n152 VDDA.t10 39.4005
R4375 VDDA.n152 VDDA.t132 39.4005
R4376 VDDA.n154 VDDA.t134 39.4005
R4377 VDDA.n154 VDDA.t173 39.4005
R4378 VDDA.n218 VDDA.t194 39.4005
R4379 VDDA.n218 VDDA.t7 39.4005
R4380 VDDA.n249 VDDA.t164 39.4005
R4381 VDDA.n249 VDDA.t364 39.4005
R4382 VDDA.n223 VDDA.t409 39.4005
R4383 VDDA.n223 VDDA.t42 39.4005
R4384 VDDA.n232 VDDA.t100 39.4005
R4385 VDDA.n232 VDDA.t75 39.4005
R4386 VDDA.n225 VDDA.t366 39.4005
R4387 VDDA.n225 VDDA.t80 39.4005
R4388 VDDA.n211 VDDA.n210 36.5719
R4389 VDDA.n213 VDDA.n212 36.5719
R4390 VDDA.n247 VDDA.n246 36.5719
R4391 VDDA.n245 VDDA.n222 36.5719
R4392 VDDA.n208 VDDA.n184 35.0481
R4393 VDDA.n191 VDDA.n185 35.0481
R4394 VDDA.n80 VDDA.n78 30.1005
R4395 VDDA.n16 VDDA.n14 30.1005
R4396 VDDA.n88 VDDA.n87 29.538
R4397 VDDA.n86 VDDA.n85 29.538
R4398 VDDA.n84 VDDA.n83 29.538
R4399 VDDA.n82 VDDA.n81 29.538
R4400 VDDA.n80 VDDA.n79 29.538
R4401 VDDA.n24 VDDA.n23 29.538
R4402 VDDA.n22 VDDA.n21 29.538
R4403 VDDA.n20 VDDA.n19 29.538
R4404 VDDA.n18 VDDA.n17 29.538
R4405 VDDA.n16 VDDA.n15 29.538
R4406 VDDA.n131 VDDA.n125 27.9413
R4407 VDDA.n255 VDDA.n254 27.2462
R4408 VDDA.n253 VDDA.n252 27.2462
R4409 VDDA.n238 VDDA.n237 27.2462
R4410 VDDA.n236 VDDA.n235 27.2462
R4411 VDDA.n230 VDDA.n229 27.2462
R4412 VDDA.n228 VDDA.n227 27.2462
R4413 VDDA.n156 VDDA.n155 26.5117
R4414 VDDA.n182 VDDA.n181 25.8913
R4415 VDDA.n178 VDDA.n177 25.8867
R4416 VDDA.n159 VDDA.n158 25.2957
R4417 VDDA.n187 VDDA.n186 25.2957
R4418 VDDA.n113 VDDA.t399 21.8894
R4419 VDDA.n113 VDDA.t292 21.8894
R4420 VDDA.n125 VDDA.n124 20.883
R4421 VDDA.n131 VDDA.t28 19.9244
R4422 VDDA.n214 VDDA.t338 19.7005
R4423 VDDA.n214 VDDA.t21 19.7005
R4424 VDDA.n220 VDDA.t360 19.7005
R4425 VDDA.n220 VDDA.t288 19.7005
R4426 VDDA.n241 VDDA.t143 19.7005
R4427 VDDA.n241 VDDA.t358 19.7005
R4428 VDDA.t350 VDDA.n244 19.7005
R4429 VDDA.n244 VDDA.t362 19.7005
R4430 VDDA.n216 VDDA.n208 16.3005
R4431 VDDA.n45 VDDA.t13 15.7605
R4432 VDDA.n45 VDDA.t56 15.7605
R4433 VDDA.n52 VDDA.t15 15.7605
R4434 VDDA.n52 VDDA.t104 15.7605
R4435 VDDA.n191 VDDA.n190 15.6443
R4436 VDDA.n190 VDDA.n186 15.488
R4437 VDDA.n189 VDDA.n188 14.9338
R4438 VDDA.n210 VDDA.n209 14.363
R4439 VDDA.n227 VDDA.n226 14.2693
R4440 VDDA.n190 VDDA.n189 14.238
R4441 VDDA.n212 VDDA.n209 14.0818
R4442 VDDA.n160 VDDA.n159 14.0713
R4443 VDDA.n252 VDDA.n251 13.8005
R4444 VDDA.n240 VDDA.n222 13.8005
R4445 VDDA.n235 VDDA.n234 13.8005
R4446 VDDA.n231 VDDA.n230 13.8005
R4447 VDDA.n239 VDDA.n238 13.8005
R4448 VDDA.n248 VDDA.n247 13.8005
R4449 VDDA.n256 VDDA.n255 13.8005
R4450 VDDA.n192 VDDA.t160 13.1338
R4451 VDDA.n192 VDDA.t393 13.1338
R4452 VDDA.n194 VDDA.t62 13.1338
R4453 VDDA.n194 VDDA.t45 13.1338
R4454 VDDA.n196 VDDA.t123 13.1338
R4455 VDDA.n196 VDDA.t180 13.1338
R4456 VDDA.n198 VDDA.t156 13.1338
R4457 VDDA.n198 VDDA.t82 13.1338
R4458 VDDA.n200 VDDA.t125 13.1338
R4459 VDDA.n200 VDDA.t158 13.1338
R4460 VDDA.n202 VDDA.t84 13.1338
R4461 VDDA.n202 VDDA.t86 13.1338
R4462 VDDA.n204 VDDA.t26 13.1338
R4463 VDDA.n204 VDDA.t405 13.1338
R4464 VDDA.n206 VDDA.t177 13.1338
R4465 VDDA.n206 VDDA.t108 13.1338
R4466 VDDA.n179 VDDA.n178 12.6486
R4467 VDDA.n157 VDDA.n156 12.6486
R4468 VDDA.n181 VDDA.n180 12.6436
R4469 VDDA.n257 VDDA.n256 11.4105
R4470 VDDA.n135 VDDA.n134 11.348
R4471 VDDA.t299 VDDA.n118 11.2576
R4472 VDDA.n118 VDDA.t228 11.2576
R4473 VDDA.n65 VDDA.t224 11.2576
R4474 VDDA.n65 VDDA.t232 11.2576
R4475 VDDA.n67 VDDA.t206 11.2576
R4476 VDDA.n67 VDDA.t216 11.2576
R4477 VDDA.n72 VDDA.t214 11.2576
R4478 VDDA.n72 VDDA.t222 11.2576
R4479 VDDA.n74 VDDA.t210 11.2576
R4480 VDDA.n74 VDDA.t218 11.2576
R4481 VDDA.n64 VDDA.t236 11.2576
R4482 VDDA.n64 VDDA.t200 11.2576
R4483 VDDA.n1 VDDA.t198 11.2576
R4484 VDDA.n1 VDDA.t208 11.2576
R4485 VDDA.n3 VDDA.t230 11.2576
R4486 VDDA.n3 VDDA.t234 11.2576
R4487 VDDA.n8 VDDA.t202 11.2576
R4488 VDDA.n8 VDDA.t196 11.2576
R4489 VDDA.n10 VDDA.t220 11.2576
R4490 VDDA.n10 VDDA.t226 11.2576
R4491 VDDA.n0 VDDA.t204 11.2576
R4492 VDDA.n0 VDDA.t212 11.2576
R4493 VDDA.n92 VDDA.n88 10.8443
R4494 VDDA.n28 VDDA.n24 10.8443
R4495 VDDA.n92 VDDA.n91 10.3755
R4496 VDDA.n28 VDDA.n27 10.3755
R4497 VDDA.n217 VDDA.n216 9.7855
R4498 VDDA.n183 VDDA.n182 8.973
R4499 VDDA.n109 VDDA.n108 8.8755
R4500 VDDA.n62 VDDA.n61 8.688
R4501 VDDA.n63 VDDA.n62 8.3755
R4502 VDDA.n109 VDDA.n77 8.1255
R4503 VDDA.n63 VDDA.n13 8.1255
R4504 VDDA.n87 VDDA.t240 8.0005
R4505 VDDA.n87 VDDA.t387 8.0005
R4506 VDDA.n85 VDDA.t40 8.0005
R4507 VDDA.n85 VDDA.t16 8.0005
R4508 VDDA.n83 VDDA.t54 8.0005
R4509 VDDA.n83 VDDA.t189 8.0005
R4510 VDDA.n81 VDDA.t139 8.0005
R4511 VDDA.n81 VDDA.t135 8.0005
R4512 VDDA.n79 VDDA.t138 8.0005
R4513 VDDA.n79 VDDA.t49 8.0005
R4514 VDDA.n78 VDDA.t116 8.0005
R4515 VDDA.n78 VDDA.t237 8.0005
R4516 VDDA.n23 VDDA.t39 8.0005
R4517 VDDA.n23 VDDA.t239 8.0005
R4518 VDDA.n21 VDDA.t171 8.0005
R4519 VDDA.n21 VDDA.t67 8.0005
R4520 VDDA.n19 VDDA.t78 8.0005
R4521 VDDA.n19 VDDA.t93 8.0005
R4522 VDDA.n17 VDDA.t144 8.0005
R4523 VDDA.n17 VDDA.t118 8.0005
R4524 VDDA.n15 VDDA.t169 8.0005
R4525 VDDA.n15 VDDA.t66 8.0005
R4526 VDDA.n14 VDDA.t238 8.0005
R4527 VDDA.n14 VDDA.t101 8.0005
R4528 VDDA.n73 VDDA.n71 7.013
R4529 VDDA.n5 VDDA.n4 7.013
R4530 VDDA.n93 VDDA.t113 6.56717
R4531 VDDA.n93 VDDA.t188 6.56717
R4532 VDDA.n95 VDDA.t137 6.56717
R4533 VDDA.n95 VDDA.t5 6.56717
R4534 VDDA.n97 VDDA.t111 6.56717
R4535 VDDA.n97 VDDA.t166 6.56717
R4536 VDDA.n99 VDDA.t385 6.56717
R4537 VDDA.n99 VDDA.t34 6.56717
R4538 VDDA.n101 VDDA.t30 6.56717
R4539 VDDA.n101 VDDA.t53 6.56717
R4540 VDDA.n29 VDDA.t375 6.56717
R4541 VDDA.n29 VDDA.t168 6.56717
R4542 VDDA.n31 VDDA.t97 6.56717
R4543 VDDA.n31 VDDA.t18 6.56717
R4544 VDDA.n33 VDDA.t371 6.56717
R4545 VDDA.n33 VDDA.t115 6.56717
R4546 VDDA.n35 VDDA.t373 6.56717
R4547 VDDA.n35 VDDA.t69 6.56717
R4548 VDDA.n37 VDDA.t377 6.56717
R4549 VDDA.n37 VDDA.t71 6.56717
R4550 VDDA.n116 VDDA.n110 6.563
R4551 VDDA.n110 VDDA.n109 6.5005
R4552 VDDA.n110 VDDA.n63 6.5005
R4553 VDDA.n108 VDDA.n107 5.8755
R4554 VDDA.n44 VDDA.n43 5.8755
R4555 VDDA.n53 VDDA.n51 5.40675
R4556 VDDA.n124 VDDA.n123 5.28175
R4557 VDDA.n116 VDDA.n115 5.28175
R4558 VDDA.n69 VDDA.n68 5.1255
R4559 VDDA.n9 VDDA.n7 5.1255
R4560 VDDA.n103 VDDA.n102 5.063
R4561 VDDA.n39 VDDA.n38 5.063
R4562 VDDA.n108 VDDA.n92 4.96925
R4563 VDDA.n44 VDDA.n28 4.96925
R4564 VDDA.n119 VDDA.n117 4.7505
R4565 VDDA.n114 VDDA.n112 4.7505
R4566 VDDA.n216 VDDA.n215 4.7505
R4567 VDDA.n135 VDDA.n131 4.5595
R4568 VDDA.n123 VDDA.n122 4.5005
R4569 VDDA.n107 VDDA.n106 4.5005
R4570 VDDA.n77 VDDA.n76 4.5005
R4571 VDDA.n55 VDDA.n54 4.5005
R4572 VDDA.n49 VDDA.n48 4.5005
R4573 VDDA.n61 VDDA.n60 4.5005
R4574 VDDA.n43 VDDA.n42 4.5005
R4575 VDDA.n13 VDDA.n12 4.5005
R4576 VDDA.n215 VDDA.n209 4.5005
R4577 VDDA.n133 VDDA.n132 4.3755
R4578 VDDA.n134 VDDA.n133 3.7505
R4579 VDDA.n258 VDDA.n257 3.71013
R4580 VDDA.n112 VDDA.n111 2.8255
R4581 VDDA.n240 VDDA.n239 2.78175
R4582 VDDA.n251 VDDA.n248 2.78175
R4583 VDDA.n91 VDDA.n90 2.40217
R4584 VDDA.n27 VDDA.n26 2.40217
R4585 VDDA.n56 VDDA.n55 2.32133
R4586 VDDA.n48 VDDA.n47 2.32133
R4587 VDDA.n60 VDDA.n59 2.32133
R4588 VDDA.n51 VDDA.n50 2.32133
R4589 VDDA.n258 VDDA.n125 2.1343
R4590 VDDA.n57 VDDA.n47 2.13383
R4591 VDDA.n57 VDDA.n56 2.13383
R4592 VDDA VDDA.n258 2.0779
R4593 VDDA.n234 VDDA.n231 2.063
R4594 VDDA.n106 VDDA.n105 1.95675
R4595 VDDA.n104 VDDA.n103 1.95675
R4596 VDDA.n42 VDDA.n41 1.95675
R4597 VDDA.n40 VDDA.n39 1.95675
R4598 VDDA.n122 VDDA.n121 1.888
R4599 VDDA.n120 VDDA.n119 1.888
R4600 VDDA.n70 VDDA.n69 1.888
R4601 VDDA.n7 VDDA.n6 1.888
R4602 VDDA.n177 VDDA.n160 1.8755
R4603 VDDA.n124 VDDA.n116 0.938
R4604 VDDA.n54 VDDA.n53 0.90675
R4605 VDDA.n49 VDDA.n46 0.90675
R4606 VDDA.n61 VDDA.n46 0.90675
R4607 VDDA.n183 VDDA.n135 0.840625
R4608 VDDA.n217 VDDA.n183 0.74075
R4609 VDDA.n231 VDDA.n226 0.65675
R4610 VDDA.n123 VDDA.n117 0.6255
R4611 VDDA.n115 VDDA.n114 0.6255
R4612 VDDA.n76 VDDA.n75 0.6255
R4613 VDDA.n75 VDDA.n73 0.6255
R4614 VDDA.n68 VDDA.n66 0.6255
R4615 VDDA.n76 VDDA.n66 0.6255
R4616 VDDA.n12 VDDA.n11 0.6255
R4617 VDDA.n11 VDDA.n9 0.6255
R4618 VDDA.n4 VDDA.n2 0.6255
R4619 VDDA.n12 VDDA.n2 0.6255
R4620 VDDA.n155 VDDA.n153 0.6255
R4621 VDDA.n153 VDDA.n151 0.6255
R4622 VDDA.n151 VDDA.n149 0.6255
R4623 VDDA.n149 VDDA.n147 0.6255
R4624 VDDA.n147 VDDA.n145 0.6255
R4625 VDDA.n145 VDDA.n143 0.6255
R4626 VDDA.n143 VDDA.n141 0.6255
R4627 VDDA.n141 VDDA.n139 0.6255
R4628 VDDA.n160 VDDA.n139 0.6255
R4629 VDDA.n177 VDDA.n176 0.6255
R4630 VDDA.n176 VDDA.n174 0.6255
R4631 VDDA.n174 VDDA.n172 0.6255
R4632 VDDA.n172 VDDA.n170 0.6255
R4633 VDDA.n170 VDDA.n168 0.6255
R4634 VDDA.n168 VDDA.n166 0.6255
R4635 VDDA.n166 VDDA.n164 0.6255
R4636 VDDA.n164 VDDA.n162 0.6255
R4637 VDDA.n162 VDDA.n137 0.6255
R4638 VDDA.n182 VDDA.n137 0.6255
R4639 VDDA.n102 VDDA.n100 0.563
R4640 VDDA.n100 VDDA.n98 0.563
R4641 VDDA.n98 VDDA.n96 0.563
R4642 VDDA.n96 VDDA.n94 0.563
R4643 VDDA.n107 VDDA.n94 0.563
R4644 VDDA.n82 VDDA.n80 0.563
R4645 VDDA.n84 VDDA.n82 0.563
R4646 VDDA.n86 VDDA.n84 0.563
R4647 VDDA.n88 VDDA.n86 0.563
R4648 VDDA.n38 VDDA.n36 0.563
R4649 VDDA.n36 VDDA.n34 0.563
R4650 VDDA.n34 VDDA.n32 0.563
R4651 VDDA.n32 VDDA.n30 0.563
R4652 VDDA.n43 VDDA.n30 0.563
R4653 VDDA.n18 VDDA.n16 0.563
R4654 VDDA.n20 VDDA.n18 0.563
R4655 VDDA.n22 VDDA.n20 0.563
R4656 VDDA.n24 VDDA.n22 0.563
R4657 VDDA.n234 VDDA.n233 0.563
R4658 VDDA.n233 VDDA.n224 0.563
R4659 VDDA.n239 VDDA.n224 0.563
R4660 VDDA.n243 VDDA.n242 0.563
R4661 VDDA.n242 VDDA.n221 0.563
R4662 VDDA.n251 VDDA.n250 0.563
R4663 VDDA.n250 VDDA.n219 0.563
R4664 VDDA.n256 VDDA.n219 0.563
R4665 VDDA VDDA.n217 0.41175
R4666 VDDA.n54 VDDA.n49 0.3755
R4667 VDDA.n62 VDDA.n44 0.3755
R4668 VDDA.n243 VDDA.n240 0.28175
R4669 VDDA.n248 VDDA.n221 0.28175
R4670 VDDA.t46 VDDA.t27 0.1603
R4671 VDDA.t183 VDDA.t87 0.1603
R4672 VDDA.t109 VDDA.t22 0.1603
R4673 VDDA.t178 VDDA.t64 0.1603
R4674 VDDA.t407 VDDA.t394 0.1603
R4675 VDDA.n127 VDDA.t395 0.159278
R4676 VDDA.n128 VDDA.t181 0.159278
R4677 VDDA.n129 VDDA.t24 0.159278
R4678 VDDA.n130 VDDA.t63 0.159278
R4679 VDDA.n130 VDDA.t406 0.1368
R4680 VDDA.n130 VDDA.t46 0.1368
R4681 VDDA.n129 VDDA.t23 0.1368
R4682 VDDA.n129 VDDA.t183 0.1368
R4683 VDDA.n128 VDDA.t121 0.1368
R4684 VDDA.n128 VDDA.t109 0.1368
R4685 VDDA.n127 VDDA.t43 0.1368
R4686 VDDA.n127 VDDA.t178 0.1368
R4687 VDDA.n126 VDDA.t182 0.1368
R4688 VDDA.n126 VDDA.t407 0.1368
R4689 VDDA.n257 VDDA 0.135625
R4690 VDDA.t395 VDDA.n126 0.00152174
R4691 VDDA.t181 VDDA.n127 0.00152174
R4692 VDDA.t24 VDDA.n128 0.00152174
R4693 VDDA.t63 VDDA.n129 0.00152174
R4694 VDDA.t28 VDDA.n130 0.00152174
R4695 bgr_9_0.V_TOP.n0 bgr_9_0.V_TOP.t29 369.534
R4696 bgr_9_0.V_TOP.n23 bgr_9_0.V_TOP.n21 345.389
R4697 bgr_9_0.V_TOP.n19 bgr_9_0.V_TOP.n18 344.7
R4698 bgr_9_0.V_TOP.n23 bgr_9_0.V_TOP.n22 344.7
R4699 bgr_9_0.V_TOP.n27 bgr_9_0.V_TOP.n26 344.7
R4700 bgr_9_0.V_TOP.n29 bgr_9_0.V_TOP.n28 344.7
R4701 bgr_9_0.V_TOP.n24 bgr_9_0.V_TOP.n20 340.2
R4702 bgr_9_0.V_TOP.n39 bgr_9_0.V_TOP.n38 224.934
R4703 bgr_9_0.V_TOP.n38 bgr_9_0.V_TOP.n37 224.934
R4704 bgr_9_0.V_TOP.n37 bgr_9_0.V_TOP.n36 224.934
R4705 bgr_9_0.V_TOP.n36 bgr_9_0.V_TOP.n35 224.934
R4706 bgr_9_0.V_TOP.n35 bgr_9_0.V_TOP.n34 224.934
R4707 bgr_9_0.V_TOP.n34 bgr_9_0.V_TOP.n33 224.934
R4708 bgr_9_0.V_TOP.n33 bgr_9_0.V_TOP.n32 224.934
R4709 bgr_9_0.V_TOP.n1 bgr_9_0.V_TOP.n0 224.934
R4710 bgr_9_0.V_TOP.n2 bgr_9_0.V_TOP.n1 224.934
R4711 bgr_9_0.V_TOP.n3 bgr_9_0.V_TOP.n2 224.934
R4712 bgr_9_0.V_TOP.n4 bgr_9_0.V_TOP.n3 224.934
R4713 bgr_9_0.V_TOP.n5 bgr_9_0.V_TOP.n4 224.934
R4714 bgr_9_0.V_TOP bgr_9_0.V_TOP.t48 214.222
R4715 bgr_9_0.V_TOP.n31 bgr_9_0.V_TOP.n30 163.175
R4716 bgr_9_0.V_TOP.n39 bgr_9_0.V_TOP.t24 144.601
R4717 bgr_9_0.V_TOP.n38 bgr_9_0.V_TOP.t33 144.601
R4718 bgr_9_0.V_TOP.n37 bgr_9_0.V_TOP.t39 144.601
R4719 bgr_9_0.V_TOP.n36 bgr_9_0.V_TOP.t16 144.601
R4720 bgr_9_0.V_TOP.n35 bgr_9_0.V_TOP.t15 144.601
R4721 bgr_9_0.V_TOP.n34 bgr_9_0.V_TOP.t28 144.601
R4722 bgr_9_0.V_TOP.n33 bgr_9_0.V_TOP.t38 144.601
R4723 bgr_9_0.V_TOP.n32 bgr_9_0.V_TOP.t14 144.601
R4724 bgr_9_0.V_TOP.n0 bgr_9_0.V_TOP.t30 144.601
R4725 bgr_9_0.V_TOP.n1 bgr_9_0.V_TOP.t18 144.601
R4726 bgr_9_0.V_TOP.n2 bgr_9_0.V_TOP.t46 144.601
R4727 bgr_9_0.V_TOP.n3 bgr_9_0.V_TOP.t37 144.601
R4728 bgr_9_0.V_TOP.n4 bgr_9_0.V_TOP.t26 144.601
R4729 bgr_9_0.V_TOP.n5 bgr_9_0.V_TOP.t27 144.601
R4730 bgr_9_0.V_TOP.n30 bgr_9_0.V_TOP.t7 111.397
R4731 bgr_9_0.V_TOP.n17 bgr_9_0.V_TOP.t3 108.424
R4732 bgr_9_0.V_TOP bgr_9_0.V_TOP.n39 69.6227
R4733 bgr_9_0.V_TOP.n32 bgr_9_0.V_TOP.n31 69.6227
R4734 bgr_9_0.V_TOP.n31 bgr_9_0.V_TOP.n5 69.6227
R4735 bgr_9_0.V_TOP.n18 bgr_9_0.V_TOP.t8 39.4005
R4736 bgr_9_0.V_TOP.n18 bgr_9_0.V_TOP.t4 39.4005
R4737 bgr_9_0.V_TOP.n20 bgr_9_0.V_TOP.t1 39.4005
R4738 bgr_9_0.V_TOP.n20 bgr_9_0.V_TOP.t2 39.4005
R4739 bgr_9_0.V_TOP.n22 bgr_9_0.V_TOP.t12 39.4005
R4740 bgr_9_0.V_TOP.n22 bgr_9_0.V_TOP.t11 39.4005
R4741 bgr_9_0.V_TOP.n21 bgr_9_0.V_TOP.t10 39.4005
R4742 bgr_9_0.V_TOP.n21 bgr_9_0.V_TOP.t0 39.4005
R4743 bgr_9_0.V_TOP.n26 bgr_9_0.V_TOP.t5 39.4005
R4744 bgr_9_0.V_TOP.n26 bgr_9_0.V_TOP.t6 39.4005
R4745 bgr_9_0.V_TOP.n28 bgr_9_0.V_TOP.t13 39.4005
R4746 bgr_9_0.V_TOP.n28 bgr_9_0.V_TOP.t9 39.4005
R4747 bgr_9_0.V_TOP.n17 bgr_9_0.V_TOP.n16 37.1479
R4748 bgr_9_0.V_TOP.n19 bgr_9_0.V_TOP.n17 27.8371
R4749 bgr_9_0.V_TOP.n24 bgr_9_0.V_TOP.n23 8.313
R4750 bgr_9_0.V_TOP.n30 bgr_9_0.V_TOP.n29 5.188
R4751 bgr_9_0.V_TOP.n6 bgr_9_0.V_TOP.t31 4.8295
R4752 bgr_9_0.V_TOP.n7 bgr_9_0.V_TOP.t22 4.8295
R4753 bgr_9_0.V_TOP.n8 bgr_9_0.V_TOP.t20 4.8295
R4754 bgr_9_0.V_TOP.n9 bgr_9_0.V_TOP.t45 4.8295
R4755 bgr_9_0.V_TOP.n10 bgr_9_0.V_TOP.t42 4.8295
R4756 bgr_9_0.V_TOP.n11 bgr_9_0.V_TOP.t36 4.8295
R4757 bgr_9_0.V_TOP.n12 bgr_9_0.V_TOP.t17 4.8295
R4758 bgr_9_0.V_TOP.n13 bgr_9_0.V_TOP.t43 4.8295
R4759 bgr_9_0.V_TOP.n14 bgr_9_0.V_TOP.t34 4.8295
R4760 bgr_9_0.V_TOP.n6 bgr_9_0.V_TOP.t35 4.5005
R4761 bgr_9_0.V_TOP.n7 bgr_9_0.V_TOP.t32 4.5005
R4762 bgr_9_0.V_TOP.n8 bgr_9_0.V_TOP.t25 4.5005
R4763 bgr_9_0.V_TOP.n9 bgr_9_0.V_TOP.t21 4.5005
R4764 bgr_9_0.V_TOP.n10 bgr_9_0.V_TOP.t49 4.5005
R4765 bgr_9_0.V_TOP.n11 bgr_9_0.V_TOP.t44 4.5005
R4766 bgr_9_0.V_TOP.n12 bgr_9_0.V_TOP.t23 4.5005
R4767 bgr_9_0.V_TOP.n13 bgr_9_0.V_TOP.t19 4.5005
R4768 bgr_9_0.V_TOP.n16 bgr_9_0.V_TOP.t40 4.5005
R4769 bgr_9_0.V_TOP.n15 bgr_9_0.V_TOP.t47 4.5005
R4770 bgr_9_0.V_TOP.n14 bgr_9_0.V_TOP.t41 4.5005
R4771 bgr_9_0.V_TOP.n25 bgr_9_0.V_TOP.n24 4.5005
R4772 bgr_9_0.V_TOP.n29 bgr_9_0.V_TOP.n27 2.1255
R4773 bgr_9_0.V_TOP.n27 bgr_9_0.V_TOP.n25 2.1255
R4774 bgr_9_0.V_TOP.n25 bgr_9_0.V_TOP.n19 2.1255
R4775 bgr_9_0.V_TOP.n7 bgr_9_0.V_TOP.n6 0.3295
R4776 bgr_9_0.V_TOP.n9 bgr_9_0.V_TOP.n8 0.3295
R4777 bgr_9_0.V_TOP.n11 bgr_9_0.V_TOP.n10 0.3295
R4778 bgr_9_0.V_TOP.n13 bgr_9_0.V_TOP.n12 0.3295
R4779 bgr_9_0.V_TOP.n16 bgr_9_0.V_TOP.n15 0.3295
R4780 bgr_9_0.V_TOP.n15 bgr_9_0.V_TOP.n14 0.3295
R4781 bgr_9_0.V_TOP.n9 bgr_9_0.V_TOP.n7 0.2825
R4782 bgr_9_0.V_TOP.n11 bgr_9_0.V_TOP.n9 0.2825
R4783 bgr_9_0.V_TOP.n13 bgr_9_0.V_TOP.n11 0.2825
R4784 bgr_9_0.V_TOP.n14 bgr_9_0.V_TOP.n13 0.2825
R4785 VOUT-.n91 VOUT-.t7 112.159
R4786 VOUT-.n4 VOUT-.n2 41.431
R4787 VOUT-.n9 VOUT-.n1 41.431
R4788 VOUT-.n8 VOUT-.n7 40.8685
R4789 VOUT-.n6 VOUT-.n5 40.8685
R4790 VOUT-.n4 VOUT-.n3 40.8685
R4791 VOUT-.n10 VOUT-.n0 36.3685
R4792 VOUT-.n88 VOUT-.n86 16.9483
R4793 VOUT-.n90 VOUT-.n89 15.8233
R4794 VOUT-.n88 VOUT-.n87 15.8233
R4795 VOUT-.n85 VOUT-.n10 15.063
R4796 VOUT-.n85 VOUT-.n84 11.5649
R4797 VOUT- VOUT-.n85 9.5005
R4798 VOUT-.n7 VOUT-.t1 6.56717
R4799 VOUT-.n7 VOUT-.t13 6.56717
R4800 VOUT-.n5 VOUT-.t4 6.56717
R4801 VOUT-.n5 VOUT-.t3 6.56717
R4802 VOUT-.n3 VOUT-.t0 6.56717
R4803 VOUT-.n3 VOUT-.t16 6.56717
R4804 VOUT-.n2 VOUT-.t8 6.56717
R4805 VOUT-.n2 VOUT-.t12 6.56717
R4806 VOUT-.n1 VOUT-.t11 6.56717
R4807 VOUT-.n1 VOUT-.t17 6.56717
R4808 VOUT-.n0 VOUT-.t2 6.56717
R4809 VOUT-.n0 VOUT-.t14 6.56717
R4810 VOUT-.n39 VOUT-.t68 4.8295
R4811 VOUT-.n47 VOUT-.t66 4.8295
R4812 VOUT-.n45 VOUT-.t115 4.8295
R4813 VOUT-.n43 VOUT-.t150 4.8295
R4814 VOUT-.n42 VOUT-.t132 4.8295
R4815 VOUT-.n41 VOUT-.t29 4.8295
R4816 VOUT-.n59 VOUT-.t125 4.8295
R4817 VOUT-.n60 VOUT-.t73 4.8295
R4818 VOUT-.n61 VOUT-.t23 4.8295
R4819 VOUT-.n62 VOUT-.t109 4.8295
R4820 VOUT-.n63 VOUT-.t76 4.8295
R4821 VOUT-.n64 VOUT-.t44 4.8295
R4822 VOUT-.n66 VOUT-.t37 4.8295
R4823 VOUT-.n67 VOUT-.t143 4.8295
R4824 VOUT-.n69 VOUT-.t70 4.8295
R4825 VOUT-.n70 VOUT-.t39 4.8295
R4826 VOUT-.n72 VOUT-.t32 4.8295
R4827 VOUT-.n73 VOUT-.t138 4.8295
R4828 VOUT-.n75 VOUT-.t131 4.8295
R4829 VOUT-.n76 VOUT-.t101 4.8295
R4830 VOUT-.n78 VOUT-.t28 4.8295
R4831 VOUT-.n79 VOUT-.t133 4.8295
R4832 VOUT-.n11 VOUT-.t26 4.8295
R4833 VOUT-.n13 VOUT-.t36 4.8295
R4834 VOUT-.n24 VOUT-.t140 4.8295
R4835 VOUT-.n25 VOUT-.t111 4.8295
R4836 VOUT-.n27 VOUT-.t41 4.8295
R4837 VOUT-.n28 VOUT-.t151 4.8295
R4838 VOUT-.n30 VOUT-.t80 4.8295
R4839 VOUT-.n31 VOUT-.t51 4.8295
R4840 VOUT-.n33 VOUT-.t49 4.8295
R4841 VOUT-.n34 VOUT-.t19 4.8295
R4842 VOUT-.n36 VOUT-.t85 4.8295
R4843 VOUT-.n37 VOUT-.t55 4.8295
R4844 VOUT-.n81 VOUT-.t124 4.8295
R4845 VOUT-.n49 VOUT-.t91 4.8154
R4846 VOUT-.n50 VOUT-.t69 4.8154
R4847 VOUT-.n51 VOUT-.t107 4.8154
R4848 VOUT-.n49 VOUT-.t31 4.806
R4849 VOUT-.n50 VOUT-.t149 4.806
R4850 VOUT-.n51 VOUT-.t50 4.806
R4851 VOUT-.n52 VOUT-.t144 4.806
R4852 VOUT-.n52 VOUT-.t83 4.806
R4853 VOUT-.n53 VOUT-.t120 4.806
R4854 VOUT-.n54 VOUT-.t104 4.806
R4855 VOUT-.n55 VOUT-.t137 4.806
R4856 VOUT-.n56 VOUT-.t35 4.806
R4857 VOUT-.n57 VOUT-.t156 4.806
R4858 VOUT-.n14 VOUT-.t71 4.806
R4859 VOUT-.n14 VOUT-.t113 4.806
R4860 VOUT-.n15 VOUT-.t114 4.806
R4861 VOUT-.n15 VOUT-.t24 4.806
R4862 VOUT-.n16 VOUT-.t65 4.806
R4863 VOUT-.n16 VOUT-.t62 4.806
R4864 VOUT-.n17 VOUT-.t154 4.806
R4865 VOUT-.n17 VOUT-.t95 4.806
R4866 VOUT-.n18 VOUT-.t105 4.806
R4867 VOUT-.n18 VOUT-.t126 4.806
R4868 VOUT-.n19 VOUT-.t141 4.806
R4869 VOUT-.n19 VOUT-.t38 4.806
R4870 VOUT-.n20 VOUT-.t92 4.806
R4871 VOUT-.n20 VOUT-.t74 4.806
R4872 VOUT-.n21 VOUT-.t42 4.806
R4873 VOUT-.n22 VOUT-.t82 4.806
R4874 VOUT-.n39 VOUT-.t86 4.5005
R4875 VOUT-.n40 VOUT-.t54 4.5005
R4876 VOUT-.n47 VOUT-.t77 4.5005
R4877 VOUT-.n48 VOUT-.t43 4.5005
R4878 VOUT-.n45 VOUT-.t58 4.5005
R4879 VOUT-.n46 VOUT-.t22 4.5005
R4880 VOUT-.n43 VOUT-.t94 4.5005
R4881 VOUT-.n44 VOUT-.t61 4.5005
R4882 VOUT-.n42 VOUT-.t99 4.5005
R4883 VOUT-.n41 VOUT-.t52 4.5005
R4884 VOUT-.n58 VOUT-.t155 4.5005
R4885 VOUT-.n57 VOUT-.t116 4.5005
R4886 VOUT-.n56 VOUT-.t136 4.5005
R4887 VOUT-.n55 VOUT-.t100 4.5005
R4888 VOUT-.n54 VOUT-.t64 4.5005
R4889 VOUT-.n53 VOUT-.t81 4.5005
R4890 VOUT-.n52 VOUT-.t45 4.5005
R4891 VOUT-.n51 VOUT-.t146 4.5005
R4892 VOUT-.n50 VOUT-.t108 4.5005
R4893 VOUT-.n49 VOUT-.t130 4.5005
R4894 VOUT-.n59 VOUT-.t152 4.5005
R4895 VOUT-.n60 VOUT-.t112 4.5005
R4896 VOUT-.n61 VOUT-.t47 4.5005
R4897 VOUT-.n62 VOUT-.t147 4.5005
R4898 VOUT-.n63 VOUT-.t27 4.5005
R4899 VOUT-.n65 VOUT-.t128 4.5005
R4900 VOUT-.n64 VOUT-.t97 4.5005
R4901 VOUT-.n66 VOUT-.t123 4.5005
R4902 VOUT-.n68 VOUT-.t88 4.5005
R4903 VOUT-.n67 VOUT-.t57 4.5005
R4904 VOUT-.n69 VOUT-.t20 4.5005
R4905 VOUT-.n71 VOUT-.t121 4.5005
R4906 VOUT-.n70 VOUT-.t87 4.5005
R4907 VOUT-.n72 VOUT-.t118 4.5005
R4908 VOUT-.n74 VOUT-.t84 4.5005
R4909 VOUT-.n73 VOUT-.t53 4.5005
R4910 VOUT-.n75 VOUT-.t79 4.5005
R4911 VOUT-.n77 VOUT-.t48 4.5005
R4912 VOUT-.n76 VOUT-.t153 4.5005
R4913 VOUT-.n78 VOUT-.t117 4.5005
R4914 VOUT-.n80 VOUT-.t78 4.5005
R4915 VOUT-.n79 VOUT-.t46 4.5005
R4916 VOUT-.n11 VOUT-.t119 4.5005
R4917 VOUT-.n12 VOUT-.t33 4.5005
R4918 VOUT-.n13 VOUT-.t122 4.5005
R4919 VOUT-.n23 VOUT-.t90 4.5005
R4920 VOUT-.n22 VOUT-.t56 4.5005
R4921 VOUT-.n21 VOUT-.t142 4.5005
R4922 VOUT-.n20 VOUT-.t110 4.5005
R4923 VOUT-.n19 VOUT-.t72 4.5005
R4924 VOUT-.n18 VOUT-.t25 4.5005
R4925 VOUT-.n17 VOUT-.t127 4.5005
R4926 VOUT-.n16 VOUT-.t93 4.5005
R4927 VOUT-.n15 VOUT-.t60 4.5005
R4928 VOUT-.n14 VOUT-.t148 4.5005
R4929 VOUT-.n24 VOUT-.t89 4.5005
R4930 VOUT-.n26 VOUT-.t59 4.5005
R4931 VOUT-.n25 VOUT-.t21 4.5005
R4932 VOUT-.n27 VOUT-.t129 4.5005
R4933 VOUT-.n29 VOUT-.t98 4.5005
R4934 VOUT-.n28 VOUT-.t63 4.5005
R4935 VOUT-.n30 VOUT-.t30 4.5005
R4936 VOUT-.n32 VOUT-.t134 4.5005
R4937 VOUT-.n31 VOUT-.t103 4.5005
R4938 VOUT-.n33 VOUT-.t135 4.5005
R4939 VOUT-.n35 VOUT-.t102 4.5005
R4940 VOUT-.n34 VOUT-.t67 4.5005
R4941 VOUT-.n36 VOUT-.t34 4.5005
R4942 VOUT-.n38 VOUT-.t139 4.5005
R4943 VOUT-.n37 VOUT-.t106 4.5005
R4944 VOUT-.n81 VOUT-.t75 4.5005
R4945 VOUT-.n82 VOUT-.t40 4.5005
R4946 VOUT-.n83 VOUT-.t145 4.5005
R4947 VOUT-.n84 VOUT-.t96 4.5005
R4948 VOUT-.n10 VOUT-.n9 4.5005
R4949 VOUT-.n89 VOUT-.t10 3.42907
R4950 VOUT-.n89 VOUT-.t15 3.42907
R4951 VOUT-.n87 VOUT-.t18 3.42907
R4952 VOUT-.n87 VOUT-.t6 3.42907
R4953 VOUT-.n86 VOUT-.t5 3.42907
R4954 VOUT-.n86 VOUT-.t9 3.42907
R4955 VOUT-.n91 VOUT-.n90 1.30519
R4956 VOUT-.n90 VOUT-.n88 1.1255
R4957 VOUT- VOUT-.n91 0.742688
R4958 VOUT-.n6 VOUT-.n4 0.563
R4959 VOUT-.n8 VOUT-.n6 0.563
R4960 VOUT-.n9 VOUT-.n8 0.563
R4961 VOUT-.n40 VOUT-.n39 0.3295
R4962 VOUT-.n48 VOUT-.n47 0.3295
R4963 VOUT-.n46 VOUT-.n45 0.3295
R4964 VOUT-.n44 VOUT-.n43 0.3295
R4965 VOUT-.n58 VOUT-.n41 0.3295
R4966 VOUT-.n58 VOUT-.n57 0.3295
R4967 VOUT-.n57 VOUT-.n56 0.3295
R4968 VOUT-.n56 VOUT-.n55 0.3295
R4969 VOUT-.n55 VOUT-.n54 0.3295
R4970 VOUT-.n54 VOUT-.n53 0.3295
R4971 VOUT-.n53 VOUT-.n52 0.3295
R4972 VOUT-.n52 VOUT-.n51 0.3295
R4973 VOUT-.n51 VOUT-.n50 0.3295
R4974 VOUT-.n50 VOUT-.n49 0.3295
R4975 VOUT-.n60 VOUT-.n59 0.3295
R4976 VOUT-.n62 VOUT-.n61 0.3295
R4977 VOUT-.n65 VOUT-.n63 0.3295
R4978 VOUT-.n65 VOUT-.n64 0.3295
R4979 VOUT-.n68 VOUT-.n66 0.3295
R4980 VOUT-.n68 VOUT-.n67 0.3295
R4981 VOUT-.n71 VOUT-.n69 0.3295
R4982 VOUT-.n71 VOUT-.n70 0.3295
R4983 VOUT-.n74 VOUT-.n72 0.3295
R4984 VOUT-.n74 VOUT-.n73 0.3295
R4985 VOUT-.n77 VOUT-.n75 0.3295
R4986 VOUT-.n77 VOUT-.n76 0.3295
R4987 VOUT-.n80 VOUT-.n78 0.3295
R4988 VOUT-.n80 VOUT-.n79 0.3295
R4989 VOUT-.n12 VOUT-.n11 0.3295
R4990 VOUT-.n23 VOUT-.n13 0.3295
R4991 VOUT-.n23 VOUT-.n22 0.3295
R4992 VOUT-.n22 VOUT-.n21 0.3295
R4993 VOUT-.n21 VOUT-.n20 0.3295
R4994 VOUT-.n20 VOUT-.n19 0.3295
R4995 VOUT-.n19 VOUT-.n18 0.3295
R4996 VOUT-.n18 VOUT-.n17 0.3295
R4997 VOUT-.n17 VOUT-.n16 0.3295
R4998 VOUT-.n16 VOUT-.n15 0.3295
R4999 VOUT-.n15 VOUT-.n14 0.3295
R5000 VOUT-.n26 VOUT-.n24 0.3295
R5001 VOUT-.n26 VOUT-.n25 0.3295
R5002 VOUT-.n29 VOUT-.n27 0.3295
R5003 VOUT-.n29 VOUT-.n28 0.3295
R5004 VOUT-.n32 VOUT-.n30 0.3295
R5005 VOUT-.n32 VOUT-.n31 0.3295
R5006 VOUT-.n35 VOUT-.n33 0.3295
R5007 VOUT-.n35 VOUT-.n34 0.3295
R5008 VOUT-.n38 VOUT-.n36 0.3295
R5009 VOUT-.n38 VOUT-.n37 0.3295
R5010 VOUT-.n82 VOUT-.n81 0.3295
R5011 VOUT-.n83 VOUT-.n82 0.3295
R5012 VOUT-.n84 VOUT-.n83 0.3295
R5013 VOUT-.n53 VOUT-.n48 0.306
R5014 VOUT-.n54 VOUT-.n46 0.306
R5015 VOUT-.n55 VOUT-.n44 0.306
R5016 VOUT-.n56 VOUT-.n42 0.306
R5017 VOUT-.n58 VOUT-.n40 0.2825
R5018 VOUT-.n60 VOUT-.n58 0.2825
R5019 VOUT-.n62 VOUT-.n60 0.2825
R5020 VOUT-.n65 VOUT-.n62 0.2825
R5021 VOUT-.n68 VOUT-.n65 0.2825
R5022 VOUT-.n71 VOUT-.n68 0.2825
R5023 VOUT-.n74 VOUT-.n71 0.2825
R5024 VOUT-.n77 VOUT-.n74 0.2825
R5025 VOUT-.n80 VOUT-.n77 0.2825
R5026 VOUT-.n23 VOUT-.n12 0.2825
R5027 VOUT-.n26 VOUT-.n23 0.2825
R5028 VOUT-.n29 VOUT-.n26 0.2825
R5029 VOUT-.n32 VOUT-.n29 0.2825
R5030 VOUT-.n35 VOUT-.n32 0.2825
R5031 VOUT-.n38 VOUT-.n35 0.2825
R5032 VOUT-.n82 VOUT-.n38 0.2825
R5033 VOUT-.n82 VOUT-.n80 0.2825
R5034 two_stage_opamp_dummy_magic_19_0.cap_res_X two_stage_opamp_dummy_magic_19_0.cap_res_X.t138 49.197
R5035 two_stage_opamp_dummy_magic_19_0.cap_res_X two_stage_opamp_dummy_magic_19_0.cap_res_X.t6 0.87
R5036 two_stage_opamp_dummy_magic_19_0.cap_res_X.t26 two_stage_opamp_dummy_magic_19_0.cap_res_X.t65 0.1603
R5037 two_stage_opamp_dummy_magic_19_0.cap_res_X.t48 two_stage_opamp_dummy_magic_19_0.cap_res_X.t87 0.1603
R5038 two_stage_opamp_dummy_magic_19_0.cap_res_X.t10 two_stage_opamp_dummy_magic_19_0.cap_res_X.t49 0.1603
R5039 two_stage_opamp_dummy_magic_19_0.cap_res_X.t111 two_stage_opamp_dummy_magic_19_0.cap_res_X.t12 0.1603
R5040 two_stage_opamp_dummy_magic_19_0.cap_res_X.t79 two_stage_opamp_dummy_magic_19_0.cap_res_X.t90 0.1603
R5041 two_stage_opamp_dummy_magic_19_0.cap_res_X.t113 two_stage_opamp_dummy_magic_19_0.cap_res_X.t79 0.1603
R5042 two_stage_opamp_dummy_magic_19_0.cap_res_X.t75 two_stage_opamp_dummy_magic_19_0.cap_res_X.t113 0.1603
R5043 two_stage_opamp_dummy_magic_19_0.cap_res_X.t98 two_stage_opamp_dummy_magic_19_0.cap_res_X.t41 0.1603
R5044 two_stage_opamp_dummy_magic_19_0.cap_res_X.t134 two_stage_opamp_dummy_magic_19_0.cap_res_X.t98 0.1603
R5045 two_stage_opamp_dummy_magic_19_0.cap_res_X.t92 two_stage_opamp_dummy_magic_19_0.cap_res_X.t134 0.1603
R5046 two_stage_opamp_dummy_magic_19_0.cap_res_X.t104 two_stage_opamp_dummy_magic_19_0.cap_res_X.t127 0.1603
R5047 two_stage_opamp_dummy_magic_19_0.cap_res_X.t70 two_stage_opamp_dummy_magic_19_0.cap_res_X.t88 0.1603
R5048 two_stage_opamp_dummy_magic_19_0.cap_res_X.t4 two_stage_opamp_dummy_magic_19_0.cap_res_X.t31 0.1603
R5049 two_stage_opamp_dummy_magic_19_0.cap_res_X.t109 two_stage_opamp_dummy_magic_19_0.cap_res_X.t133 0.1603
R5050 two_stage_opamp_dummy_magic_19_0.cap_res_X.t59 two_stage_opamp_dummy_magic_19_0.cap_res_X.t112 0.1603
R5051 two_stage_opamp_dummy_magic_19_0.cap_res_X.t129 two_stage_opamp_dummy_magic_19_0.cap_res_X.t80 0.1603
R5052 two_stage_opamp_dummy_magic_19_0.cap_res_X.t99 two_stage_opamp_dummy_magic_19_0.cap_res_X.t13 0.1603
R5053 two_stage_opamp_dummy_magic_19_0.cap_res_X.t33 two_stage_opamp_dummy_magic_19_0.cap_res_X.t119 0.1603
R5054 two_stage_opamp_dummy_magic_19_0.cap_res_X.t69 two_stage_opamp_dummy_magic_19_0.cap_res_X.t117 0.1603
R5055 two_stage_opamp_dummy_magic_19_0.cap_res_X.t136 two_stage_opamp_dummy_magic_19_0.cap_res_X.t86 0.1603
R5056 two_stage_opamp_dummy_magic_19_0.cap_res_X.t103 two_stage_opamp_dummy_magic_19_0.cap_res_X.t18 0.1603
R5057 two_stage_opamp_dummy_magic_19_0.cap_res_X.t38 two_stage_opamp_dummy_magic_19_0.cap_res_X.t124 0.1603
R5058 two_stage_opamp_dummy_magic_19_0.cap_res_X.t3 two_stage_opamp_dummy_magic_19_0.cap_res_X.t55 0.1603
R5059 two_stage_opamp_dummy_magic_19_0.cap_res_X.t77 two_stage_opamp_dummy_magic_19_0.cap_res_X.t25 0.1603
R5060 two_stage_opamp_dummy_magic_19_0.cap_res_X.t110 two_stage_opamp_dummy_magic_19_0.cap_res_X.t23 0.1603
R5061 two_stage_opamp_dummy_magic_19_0.cap_res_X.t39 two_stage_opamp_dummy_magic_19_0.cap_res_X.t128 0.1603
R5062 two_stage_opamp_dummy_magic_19_0.cap_res_X.t11 two_stage_opamp_dummy_magic_19_0.cap_res_X.t60 0.1603
R5063 two_stage_opamp_dummy_magic_19_0.cap_res_X.t81 two_stage_opamp_dummy_magic_19_0.cap_res_X.t32 0.1603
R5064 two_stage_opamp_dummy_magic_19_0.cap_res_X.t50 two_stage_opamp_dummy_magic_19_0.cap_res_X.t101 0.1603
R5065 two_stage_opamp_dummy_magic_19_0.cap_res_X.t122 two_stage_opamp_dummy_magic_19_0.cap_res_X.t71 0.1603
R5066 two_stage_opamp_dummy_magic_19_0.cap_res_X.t89 two_stage_opamp_dummy_magic_19_0.cap_res_X.t137 0.1603
R5067 two_stage_opamp_dummy_magic_19_0.cap_res_X.t21 two_stage_opamp_dummy_magic_19_0.cap_res_X.t107 0.1603
R5068 two_stage_opamp_dummy_magic_19_0.cap_res_X.t53 two_stage_opamp_dummy_magic_19_0.cap_res_X.t105 0.1603
R5069 two_stage_opamp_dummy_magic_19_0.cap_res_X.t126 two_stage_opamp_dummy_magic_19_0.cap_res_X.t76 0.1603
R5070 two_stage_opamp_dummy_magic_19_0.cap_res_X.t93 two_stage_opamp_dummy_magic_19_0.cap_res_X.t5 0.1603
R5071 two_stage_opamp_dummy_magic_19_0.cap_res_X.t27 two_stage_opamp_dummy_magic_19_0.cap_res_X.t115 0.1603
R5072 two_stage_opamp_dummy_magic_19_0.cap_res_X.t135 two_stage_opamp_dummy_magic_19_0.cap_res_X.t45 0.1603
R5073 two_stage_opamp_dummy_magic_19_0.cap_res_X.t67 two_stage_opamp_dummy_magic_19_0.cap_res_X.t16 0.1603
R5074 two_stage_opamp_dummy_magic_19_0.cap_res_X.t8 two_stage_opamp_dummy_magic_19_0.cap_res_X.t85 0.1603
R5075 two_stage_opamp_dummy_magic_19_0.cap_res_X.t96 two_stage_opamp_dummy_magic_19_0.cap_res_X.t42 0.1603
R5076 two_stage_opamp_dummy_magic_19_0.cap_res_X.t63 two_stage_opamp_dummy_magic_19_0.cap_res_X.t91 0.1603
R5077 two_stage_opamp_dummy_magic_19_0.cap_res_X.t29 two_stage_opamp_dummy_magic_19_0.cap_res_X.t2 0.1603
R5078 two_stage_opamp_dummy_magic_19_0.cap_res_X.t131 two_stage_opamp_dummy_magic_19_0.cap_res_X.t51 0.1603
R5079 two_stage_opamp_dummy_magic_19_0.cap_res_X.t84 two_stage_opamp_dummy_magic_19_0.cap_res_X.t15 0.1603
R5080 two_stage_opamp_dummy_magic_19_0.cap_res_X.t46 two_stage_opamp_dummy_magic_19_0.cap_res_X.t64 0.1603
R5081 two_stage_opamp_dummy_magic_19_0.cap_res_X.t14 two_stage_opamp_dummy_magic_19_0.cap_res_X.t114 0.1603
R5082 two_stage_opamp_dummy_magic_19_0.cap_res_X.t100 two_stage_opamp_dummy_magic_19_0.cap_res_X.t74 0.1603
R5083 two_stage_opamp_dummy_magic_19_0.cap_res_X.t34 two_stage_opamp_dummy_magic_19_0.cap_res_X.t120 0.1603
R5084 two_stage_opamp_dummy_magic_19_0.cap_res_X.t37 two_stage_opamp_dummy_magic_19_0.cap_res_X.t130 0.1603
R5085 two_stage_opamp_dummy_magic_19_0.cap_res_X.t57 two_stage_opamp_dummy_magic_19_0.cap_res_X.t24 0.1603
R5086 two_stage_opamp_dummy_magic_19_0.cap_res_X.t20 two_stage_opamp_dummy_magic_19_0.cap_res_X.t57 0.1603
R5087 two_stage_opamp_dummy_magic_19_0.cap_res_X.t95 two_stage_opamp_dummy_magic_19_0.cap_res_X.t56 0.1603
R5088 two_stage_opamp_dummy_magic_19_0.cap_res_X.t62 two_stage_opamp_dummy_magic_19_0.cap_res_X.t95 0.1603
R5089 two_stage_opamp_dummy_magic_19_0.cap_res_X.t6 two_stage_opamp_dummy_magic_19_0.cap_res_X.t62 0.1603
R5090 two_stage_opamp_dummy_magic_19_0.cap_res_X.n28 two_stage_opamp_dummy_magic_19_0.cap_res_X.t125 0.159278
R5091 two_stage_opamp_dummy_magic_19_0.cap_res_X.n29 two_stage_opamp_dummy_magic_19_0.cap_res_X.t7 0.159278
R5092 two_stage_opamp_dummy_magic_19_0.cap_res_X.n30 two_stage_opamp_dummy_magic_19_0.cap_res_X.t106 0.159278
R5093 two_stage_opamp_dummy_magic_19_0.cap_res_X.n31 two_stage_opamp_dummy_magic_19_0.cap_res_X.t73 0.159278
R5094 two_stage_opamp_dummy_magic_19_0.cap_res_X.n32 two_stage_opamp_dummy_magic_19_0.cap_res_X.t36 0.159278
R5095 two_stage_opamp_dummy_magic_19_0.cap_res_X.n33 two_stage_opamp_dummy_magic_19_0.cap_res_X.t52 0.159278
R5096 two_stage_opamp_dummy_magic_19_0.cap_res_X.n25 two_stage_opamp_dummy_magic_19_0.cap_res_X.t102 0.159278
R5097 two_stage_opamp_dummy_magic_19_0.cap_res_X.n0 two_stage_opamp_dummy_magic_19_0.cap_res_X.t43 0.159278
R5098 two_stage_opamp_dummy_magic_19_0.cap_res_X.n1 two_stage_opamp_dummy_magic_19_0.cap_res_X.t132 0.159278
R5099 two_stage_opamp_dummy_magic_19_0.cap_res_X.n2 two_stage_opamp_dummy_magic_19_0.cap_res_X.t94 0.159278
R5100 two_stage_opamp_dummy_magic_19_0.cap_res_X.n3 two_stage_opamp_dummy_magic_19_0.cap_res_X.t61 0.159278
R5101 two_stage_opamp_dummy_magic_19_0.cap_res_X.n4 two_stage_opamp_dummy_magic_19_0.cap_res_X.t30 0.159278
R5102 two_stage_opamp_dummy_magic_19_0.cap_res_X.n5 two_stage_opamp_dummy_magic_19_0.cap_res_X.t118 0.159278
R5103 two_stage_opamp_dummy_magic_19_0.cap_res_X.n6 two_stage_opamp_dummy_magic_19_0.cap_res_X.t82 0.159278
R5104 two_stage_opamp_dummy_magic_19_0.cap_res_X.t66 two_stage_opamp_dummy_magic_19_0.cap_res_X.n9 0.159278
R5105 two_stage_opamp_dummy_magic_19_0.cap_res_X.t97 two_stage_opamp_dummy_magic_19_0.cap_res_X.n10 0.159278
R5106 two_stage_opamp_dummy_magic_19_0.cap_res_X.t58 two_stage_opamp_dummy_magic_19_0.cap_res_X.n11 0.159278
R5107 two_stage_opamp_dummy_magic_19_0.cap_res_X.t22 two_stage_opamp_dummy_magic_19_0.cap_res_X.n12 0.159278
R5108 two_stage_opamp_dummy_magic_19_0.cap_res_X.t54 two_stage_opamp_dummy_magic_19_0.cap_res_X.n13 0.159278
R5109 two_stage_opamp_dummy_magic_19_0.cap_res_X.t17 two_stage_opamp_dummy_magic_19_0.cap_res_X.n14 0.159278
R5110 two_stage_opamp_dummy_magic_19_0.cap_res_X.t116 two_stage_opamp_dummy_magic_19_0.cap_res_X.n15 0.159278
R5111 two_stage_opamp_dummy_magic_19_0.cap_res_X.t78 two_stage_opamp_dummy_magic_19_0.cap_res_X.n16 0.159278
R5112 two_stage_opamp_dummy_magic_19_0.cap_res_X.t108 two_stage_opamp_dummy_magic_19_0.cap_res_X.n17 0.159278
R5113 two_stage_opamp_dummy_magic_19_0.cap_res_X.t72 two_stage_opamp_dummy_magic_19_0.cap_res_X.n18 0.159278
R5114 two_stage_opamp_dummy_magic_19_0.cap_res_X.t35 two_stage_opamp_dummy_magic_19_0.cap_res_X.n19 0.159278
R5115 two_stage_opamp_dummy_magic_19_0.cap_res_X.t68 two_stage_opamp_dummy_magic_19_0.cap_res_X.n20 0.159278
R5116 two_stage_opamp_dummy_magic_19_0.cap_res_X.t28 two_stage_opamp_dummy_magic_19_0.cap_res_X.n21 0.159278
R5117 two_stage_opamp_dummy_magic_19_0.cap_res_X.t9 two_stage_opamp_dummy_magic_19_0.cap_res_X.n22 0.159278
R5118 two_stage_opamp_dummy_magic_19_0.cap_res_X.t44 two_stage_opamp_dummy_magic_19_0.cap_res_X.n23 0.159278
R5119 two_stage_opamp_dummy_magic_19_0.cap_res_X.t1 two_stage_opamp_dummy_magic_19_0.cap_res_X.n24 0.159278
R5120 two_stage_opamp_dummy_magic_19_0.cap_res_X.n26 two_stage_opamp_dummy_magic_19_0.cap_res_X.t0 0.159278
R5121 two_stage_opamp_dummy_magic_19_0.cap_res_X.n27 two_stage_opamp_dummy_magic_19_0.cap_res_X.t121 0.159278
R5122 two_stage_opamp_dummy_magic_19_0.cap_res_X.n34 two_stage_opamp_dummy_magic_19_0.cap_res_X.t19 0.159278
R5123 two_stage_opamp_dummy_magic_19_0.cap_res_X.t102 two_stage_opamp_dummy_magic_19_0.cap_res_X.t70 0.137822
R5124 two_stage_opamp_dummy_magic_19_0.cap_res_X.n25 two_stage_opamp_dummy_magic_19_0.cap_res_X.t104 0.1368
R5125 two_stage_opamp_dummy_magic_19_0.cap_res_X.n24 two_stage_opamp_dummy_magic_19_0.cap_res_X.t83 0.1368
R5126 two_stage_opamp_dummy_magic_19_0.cap_res_X.n24 two_stage_opamp_dummy_magic_19_0.cap_res_X.t4 0.1368
R5127 two_stage_opamp_dummy_magic_19_0.cap_res_X.n23 two_stage_opamp_dummy_magic_19_0.cap_res_X.t47 0.1368
R5128 two_stage_opamp_dummy_magic_19_0.cap_res_X.n23 two_stage_opamp_dummy_magic_19_0.cap_res_X.t109 0.1368
R5129 two_stage_opamp_dummy_magic_19_0.cap_res_X.n22 two_stage_opamp_dummy_magic_19_0.cap_res_X.t59 0.1368
R5130 two_stage_opamp_dummy_magic_19_0.cap_res_X.n22 two_stage_opamp_dummy_magic_19_0.cap_res_X.t129 0.1368
R5131 two_stage_opamp_dummy_magic_19_0.cap_res_X.n21 two_stage_opamp_dummy_magic_19_0.cap_res_X.t99 0.1368
R5132 two_stage_opamp_dummy_magic_19_0.cap_res_X.n21 two_stage_opamp_dummy_magic_19_0.cap_res_X.t33 0.1368
R5133 two_stage_opamp_dummy_magic_19_0.cap_res_X.n20 two_stage_opamp_dummy_magic_19_0.cap_res_X.t69 0.1368
R5134 two_stage_opamp_dummy_magic_19_0.cap_res_X.n20 two_stage_opamp_dummy_magic_19_0.cap_res_X.t136 0.1368
R5135 two_stage_opamp_dummy_magic_19_0.cap_res_X.n19 two_stage_opamp_dummy_magic_19_0.cap_res_X.t103 0.1368
R5136 two_stage_opamp_dummy_magic_19_0.cap_res_X.n19 two_stage_opamp_dummy_magic_19_0.cap_res_X.t38 0.1368
R5137 two_stage_opamp_dummy_magic_19_0.cap_res_X.n18 two_stage_opamp_dummy_magic_19_0.cap_res_X.t3 0.1368
R5138 two_stage_opamp_dummy_magic_19_0.cap_res_X.n18 two_stage_opamp_dummy_magic_19_0.cap_res_X.t77 0.1368
R5139 two_stage_opamp_dummy_magic_19_0.cap_res_X.n17 two_stage_opamp_dummy_magic_19_0.cap_res_X.t110 0.1368
R5140 two_stage_opamp_dummy_magic_19_0.cap_res_X.n17 two_stage_opamp_dummy_magic_19_0.cap_res_X.t39 0.1368
R5141 two_stage_opamp_dummy_magic_19_0.cap_res_X.n16 two_stage_opamp_dummy_magic_19_0.cap_res_X.t11 0.1368
R5142 two_stage_opamp_dummy_magic_19_0.cap_res_X.n16 two_stage_opamp_dummy_magic_19_0.cap_res_X.t81 0.1368
R5143 two_stage_opamp_dummy_magic_19_0.cap_res_X.n15 two_stage_opamp_dummy_magic_19_0.cap_res_X.t50 0.1368
R5144 two_stage_opamp_dummy_magic_19_0.cap_res_X.n15 two_stage_opamp_dummy_magic_19_0.cap_res_X.t122 0.1368
R5145 two_stage_opamp_dummy_magic_19_0.cap_res_X.n14 two_stage_opamp_dummy_magic_19_0.cap_res_X.t89 0.1368
R5146 two_stage_opamp_dummy_magic_19_0.cap_res_X.n14 two_stage_opamp_dummy_magic_19_0.cap_res_X.t21 0.1368
R5147 two_stage_opamp_dummy_magic_19_0.cap_res_X.n13 two_stage_opamp_dummy_magic_19_0.cap_res_X.t53 0.1368
R5148 two_stage_opamp_dummy_magic_19_0.cap_res_X.n13 two_stage_opamp_dummy_magic_19_0.cap_res_X.t126 0.1368
R5149 two_stage_opamp_dummy_magic_19_0.cap_res_X.n12 two_stage_opamp_dummy_magic_19_0.cap_res_X.t93 0.1368
R5150 two_stage_opamp_dummy_magic_19_0.cap_res_X.n12 two_stage_opamp_dummy_magic_19_0.cap_res_X.t27 0.1368
R5151 two_stage_opamp_dummy_magic_19_0.cap_res_X.n11 two_stage_opamp_dummy_magic_19_0.cap_res_X.t135 0.1368
R5152 two_stage_opamp_dummy_magic_19_0.cap_res_X.n11 two_stage_opamp_dummy_magic_19_0.cap_res_X.t67 0.1368
R5153 two_stage_opamp_dummy_magic_19_0.cap_res_X.n10 two_stage_opamp_dummy_magic_19_0.cap_res_X.t34 0.1368
R5154 two_stage_opamp_dummy_magic_19_0.cap_res_X.n9 two_stage_opamp_dummy_magic_19_0.cap_res_X.t37 0.1368
R5155 two_stage_opamp_dummy_magic_19_0.cap_res_X.n29 two_stage_opamp_dummy_magic_19_0.cap_res_X.n28 0.1133
R5156 two_stage_opamp_dummy_magic_19_0.cap_res_X.n30 two_stage_opamp_dummy_magic_19_0.cap_res_X.n29 0.1133
R5157 two_stage_opamp_dummy_magic_19_0.cap_res_X.n31 two_stage_opamp_dummy_magic_19_0.cap_res_X.n30 0.1133
R5158 two_stage_opamp_dummy_magic_19_0.cap_res_X.n32 two_stage_opamp_dummy_magic_19_0.cap_res_X.n31 0.1133
R5159 two_stage_opamp_dummy_magic_19_0.cap_res_X.n33 two_stage_opamp_dummy_magic_19_0.cap_res_X.n32 0.1133
R5160 two_stage_opamp_dummy_magic_19_0.cap_res_X.n1 two_stage_opamp_dummy_magic_19_0.cap_res_X.n0 0.1133
R5161 two_stage_opamp_dummy_magic_19_0.cap_res_X.n2 two_stage_opamp_dummy_magic_19_0.cap_res_X.n1 0.1133
R5162 two_stage_opamp_dummy_magic_19_0.cap_res_X.n3 two_stage_opamp_dummy_magic_19_0.cap_res_X.n2 0.1133
R5163 two_stage_opamp_dummy_magic_19_0.cap_res_X.n4 two_stage_opamp_dummy_magic_19_0.cap_res_X.n3 0.1133
R5164 two_stage_opamp_dummy_magic_19_0.cap_res_X.n5 two_stage_opamp_dummy_magic_19_0.cap_res_X.n4 0.1133
R5165 two_stage_opamp_dummy_magic_19_0.cap_res_X.n6 two_stage_opamp_dummy_magic_19_0.cap_res_X.n5 0.1133
R5166 two_stage_opamp_dummy_magic_19_0.cap_res_X.n7 two_stage_opamp_dummy_magic_19_0.cap_res_X.n6 0.1133
R5167 two_stage_opamp_dummy_magic_19_0.cap_res_X.n8 two_stage_opamp_dummy_magic_19_0.cap_res_X.n7 0.1133
R5168 two_stage_opamp_dummy_magic_19_0.cap_res_X.n10 two_stage_opamp_dummy_magic_19_0.cap_res_X.n8 0.1133
R5169 two_stage_opamp_dummy_magic_19_0.cap_res_X.n26 two_stage_opamp_dummy_magic_19_0.cap_res_X.n25 0.1133
R5170 two_stage_opamp_dummy_magic_19_0.cap_res_X.n27 two_stage_opamp_dummy_magic_19_0.cap_res_X.n26 0.1133
R5171 two_stage_opamp_dummy_magic_19_0.cap_res_X.n34 two_stage_opamp_dummy_magic_19_0.cap_res_X.n27 0.1133
R5172 two_stage_opamp_dummy_magic_19_0.cap_res_X.n34 two_stage_opamp_dummy_magic_19_0.cap_res_X.n33 0.1133
R5173 two_stage_opamp_dummy_magic_19_0.cap_res_X.n28 two_stage_opamp_dummy_magic_19_0.cap_res_X.t26 0.00152174
R5174 two_stage_opamp_dummy_magic_19_0.cap_res_X.n29 two_stage_opamp_dummy_magic_19_0.cap_res_X.t48 0.00152174
R5175 two_stage_opamp_dummy_magic_19_0.cap_res_X.n30 two_stage_opamp_dummy_magic_19_0.cap_res_X.t10 0.00152174
R5176 two_stage_opamp_dummy_magic_19_0.cap_res_X.n31 two_stage_opamp_dummy_magic_19_0.cap_res_X.t111 0.00152174
R5177 two_stage_opamp_dummy_magic_19_0.cap_res_X.n32 two_stage_opamp_dummy_magic_19_0.cap_res_X.t75 0.00152174
R5178 two_stage_opamp_dummy_magic_19_0.cap_res_X.n33 two_stage_opamp_dummy_magic_19_0.cap_res_X.t92 0.00152174
R5179 two_stage_opamp_dummy_magic_19_0.cap_res_X.n0 two_stage_opamp_dummy_magic_19_0.cap_res_X.t8 0.00152174
R5180 two_stage_opamp_dummy_magic_19_0.cap_res_X.n1 two_stage_opamp_dummy_magic_19_0.cap_res_X.t96 0.00152174
R5181 two_stage_opamp_dummy_magic_19_0.cap_res_X.n2 two_stage_opamp_dummy_magic_19_0.cap_res_X.t63 0.00152174
R5182 two_stage_opamp_dummy_magic_19_0.cap_res_X.n3 two_stage_opamp_dummy_magic_19_0.cap_res_X.t29 0.00152174
R5183 two_stage_opamp_dummy_magic_19_0.cap_res_X.n4 two_stage_opamp_dummy_magic_19_0.cap_res_X.t131 0.00152174
R5184 two_stage_opamp_dummy_magic_19_0.cap_res_X.n5 two_stage_opamp_dummy_magic_19_0.cap_res_X.t84 0.00152174
R5185 two_stage_opamp_dummy_magic_19_0.cap_res_X.n6 two_stage_opamp_dummy_magic_19_0.cap_res_X.t46 0.00152174
R5186 two_stage_opamp_dummy_magic_19_0.cap_res_X.n7 two_stage_opamp_dummy_magic_19_0.cap_res_X.t14 0.00152174
R5187 two_stage_opamp_dummy_magic_19_0.cap_res_X.n8 two_stage_opamp_dummy_magic_19_0.cap_res_X.t100 0.00152174
R5188 two_stage_opamp_dummy_magic_19_0.cap_res_X.n9 two_stage_opamp_dummy_magic_19_0.cap_res_X.t123 0.00152174
R5189 two_stage_opamp_dummy_magic_19_0.cap_res_X.n10 two_stage_opamp_dummy_magic_19_0.cap_res_X.t66 0.00152174
R5190 two_stage_opamp_dummy_magic_19_0.cap_res_X.n11 two_stage_opamp_dummy_magic_19_0.cap_res_X.t97 0.00152174
R5191 two_stage_opamp_dummy_magic_19_0.cap_res_X.n12 two_stage_opamp_dummy_magic_19_0.cap_res_X.t58 0.00152174
R5192 two_stage_opamp_dummy_magic_19_0.cap_res_X.n13 two_stage_opamp_dummy_magic_19_0.cap_res_X.t22 0.00152174
R5193 two_stage_opamp_dummy_magic_19_0.cap_res_X.n14 two_stage_opamp_dummy_magic_19_0.cap_res_X.t54 0.00152174
R5194 two_stage_opamp_dummy_magic_19_0.cap_res_X.n15 two_stage_opamp_dummy_magic_19_0.cap_res_X.t17 0.00152174
R5195 two_stage_opamp_dummy_magic_19_0.cap_res_X.n16 two_stage_opamp_dummy_magic_19_0.cap_res_X.t116 0.00152174
R5196 two_stage_opamp_dummy_magic_19_0.cap_res_X.n17 two_stage_opamp_dummy_magic_19_0.cap_res_X.t78 0.00152174
R5197 two_stage_opamp_dummy_magic_19_0.cap_res_X.n18 two_stage_opamp_dummy_magic_19_0.cap_res_X.t108 0.00152174
R5198 two_stage_opamp_dummy_magic_19_0.cap_res_X.n19 two_stage_opamp_dummy_magic_19_0.cap_res_X.t72 0.00152174
R5199 two_stage_opamp_dummy_magic_19_0.cap_res_X.n20 two_stage_opamp_dummy_magic_19_0.cap_res_X.t35 0.00152174
R5200 two_stage_opamp_dummy_magic_19_0.cap_res_X.n21 two_stage_opamp_dummy_magic_19_0.cap_res_X.t68 0.00152174
R5201 two_stage_opamp_dummy_magic_19_0.cap_res_X.n22 two_stage_opamp_dummy_magic_19_0.cap_res_X.t28 0.00152174
R5202 two_stage_opamp_dummy_magic_19_0.cap_res_X.n23 two_stage_opamp_dummy_magic_19_0.cap_res_X.t9 0.00152174
R5203 two_stage_opamp_dummy_magic_19_0.cap_res_X.n24 two_stage_opamp_dummy_magic_19_0.cap_res_X.t44 0.00152174
R5204 two_stage_opamp_dummy_magic_19_0.cap_res_X.n25 two_stage_opamp_dummy_magic_19_0.cap_res_X.t1 0.00152174
R5205 two_stage_opamp_dummy_magic_19_0.cap_res_X.n26 two_stage_opamp_dummy_magic_19_0.cap_res_X.t40 0.00152174
R5206 two_stage_opamp_dummy_magic_19_0.cap_res_X.n27 two_stage_opamp_dummy_magic_19_0.cap_res_X.t20 0.00152174
R5207 two_stage_opamp_dummy_magic_19_0.cap_res_X.t56 two_stage_opamp_dummy_magic_19_0.cap_res_X.n34 0.00152174
R5208 two_stage_opamp_dummy_magic_19_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_19_0.err_amp_mir.t5 573.044
R5209 two_stage_opamp_dummy_magic_19_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_19_0.err_amp_mir.t1 433.8
R5210 two_stage_opamp_dummy_magic_19_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_19_0.err_amp_mir.n1 163.978
R5211 two_stage_opamp_dummy_magic_19_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_19_0.err_amp_mir.n0 110.843
R5212 two_stage_opamp_dummy_magic_19_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_19_0.err_amp_mir.n2 33.0088
R5213 two_stage_opamp_dummy_magic_19_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_19_0.err_amp_mir.t0 15.7605
R5214 two_stage_opamp_dummy_magic_19_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_19_0.err_amp_mir.t4 15.7605
R5215 two_stage_opamp_dummy_magic_19_0.err_amp_mir.t2 two_stage_opamp_dummy_magic_19_0.err_amp_mir.n3 9.6005
R5216 two_stage_opamp_dummy_magic_19_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_19_0.err_amp_mir.t3 9.6005
R5217 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t25 610.534
R5218 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t13 610.534
R5219 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t27 488.428
R5220 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t16 488.428
R5221 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t9 433.8
R5222 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t18 433.8
R5223 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t26 433.8
R5224 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t15 433.8
R5225 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t22 433.8
R5226 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t11 433.8
R5227 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t23 433.8
R5228 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t14 433.8
R5229 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t21 433.8
R5230 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t10 433.8
R5231 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t19 433.8
R5232 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t8 433.8
R5233 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t17 433.8
R5234 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t24 433.8
R5235 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t12 433.8
R5236 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t20 433.8
R5237 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n22 321.914
R5238 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n0 264.63
R5239 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n7 176.733
R5240 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n8 176.733
R5241 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n9 176.733
R5242 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n10 176.733
R5243 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n11 176.733
R5244 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n12 176.733
R5245 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n13 176.733
R5246 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n14 176.733
R5247 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n15 176.733
R5248 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n16 176.733
R5249 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n17 176.733
R5250 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n18 176.733
R5251 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n19 176.733
R5252 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n20 176.733
R5253 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n23 161.3
R5254 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n1 117.001
R5255 bgr_9_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_19_0.V_tail_gate.n2 73.188
R5256 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n4 59.5797
R5257 bgr_9_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_19_0.V_tail_gate.n25 59.1277
R5258 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n6 56.2338
R5259 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n21 56.2338
R5260 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n3 50.0172
R5261 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t6 19.7005
R5262 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t0 19.7005
R5263 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t4 19.7005
R5264 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t5 19.7005
R5265 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t1 16.0005
R5266 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t7 16.0005
R5267 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t3 16.0005
R5268 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t2 16.0005
R5269 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n5 5.15154
R5270 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n24 5.07342
R5271 two_stage_opamp_dummy_magic_19_0.V_source.n1 two_stage_opamp_dummy_magic_19_0.V_source.t19 84.0067
R5272 two_stage_opamp_dummy_magic_19_0.V_source.n12 two_stage_opamp_dummy_magic_19_0.V_source.n10 54.8505
R5273 two_stage_opamp_dummy_magic_19_0.V_source.n5 two_stage_opamp_dummy_magic_19_0.V_source.n3 54.8505
R5274 two_stage_opamp_dummy_magic_19_0.V_source.n18 two_stage_opamp_dummy_magic_19_0.V_source.n17 54.288
R5275 two_stage_opamp_dummy_magic_19_0.V_source.n16 two_stage_opamp_dummy_magic_19_0.V_source.n15 54.288
R5276 two_stage_opamp_dummy_magic_19_0.V_source.n14 two_stage_opamp_dummy_magic_19_0.V_source.n13 54.288
R5277 two_stage_opamp_dummy_magic_19_0.V_source.n12 two_stage_opamp_dummy_magic_19_0.V_source.n11 54.288
R5278 two_stage_opamp_dummy_magic_19_0.V_source.n9 two_stage_opamp_dummy_magic_19_0.V_source.n8 54.288
R5279 two_stage_opamp_dummy_magic_19_0.V_source.n7 two_stage_opamp_dummy_magic_19_0.V_source.n6 54.288
R5280 two_stage_opamp_dummy_magic_19_0.V_source.n5 two_stage_opamp_dummy_magic_19_0.V_source.n4 54.288
R5281 two_stage_opamp_dummy_magic_19_0.V_source.n20 two_stage_opamp_dummy_magic_19_0.V_source.n2 49.7672
R5282 two_stage_opamp_dummy_magic_19_0.V_source.n28 two_stage_opamp_dummy_magic_19_0.V_source.n26 38.0713
R5283 two_stage_opamp_dummy_magic_19_0.V_source.n36 two_stage_opamp_dummy_magic_19_0.V_source.n35 37.5088
R5284 two_stage_opamp_dummy_magic_19_0.V_source.n34 two_stage_opamp_dummy_magic_19_0.V_source.n33 37.5088
R5285 two_stage_opamp_dummy_magic_19_0.V_source.n32 two_stage_opamp_dummy_magic_19_0.V_source.n31 37.5088
R5286 two_stage_opamp_dummy_magic_19_0.V_source.n30 two_stage_opamp_dummy_magic_19_0.V_source.n29 37.5088
R5287 two_stage_opamp_dummy_magic_19_0.V_source.n28 two_stage_opamp_dummy_magic_19_0.V_source.n27 37.5088
R5288 two_stage_opamp_dummy_magic_19_0.V_source.n25 two_stage_opamp_dummy_magic_19_0.V_source.n24 37.5088
R5289 two_stage_opamp_dummy_magic_19_0.V_source.n1 two_stage_opamp_dummy_magic_19_0.V_source.n0 37.5088
R5290 two_stage_opamp_dummy_magic_19_0.V_source.n38 two_stage_opamp_dummy_magic_19_0.V_source.n37 37.5088
R5291 two_stage_opamp_dummy_magic_19_0.V_source.n22 two_stage_opamp_dummy_magic_19_0.V_source.n21 32.988
R5292 two_stage_opamp_dummy_magic_19_0.V_source.n17 two_stage_opamp_dummy_magic_19_0.V_source.t6 16.0005
R5293 two_stage_opamp_dummy_magic_19_0.V_source.n17 two_stage_opamp_dummy_magic_19_0.V_source.t39 16.0005
R5294 two_stage_opamp_dummy_magic_19_0.V_source.n15 two_stage_opamp_dummy_magic_19_0.V_source.t10 16.0005
R5295 two_stage_opamp_dummy_magic_19_0.V_source.n15 two_stage_opamp_dummy_magic_19_0.V_source.t7 16.0005
R5296 two_stage_opamp_dummy_magic_19_0.V_source.n13 two_stage_opamp_dummy_magic_19_0.V_source.t1 16.0005
R5297 two_stage_opamp_dummy_magic_19_0.V_source.n13 two_stage_opamp_dummy_magic_19_0.V_source.t9 16.0005
R5298 two_stage_opamp_dummy_magic_19_0.V_source.n11 two_stage_opamp_dummy_magic_19_0.V_source.t3 16.0005
R5299 two_stage_opamp_dummy_magic_19_0.V_source.n11 two_stage_opamp_dummy_magic_19_0.V_source.t15 16.0005
R5300 two_stage_opamp_dummy_magic_19_0.V_source.n10 two_stage_opamp_dummy_magic_19_0.V_source.t18 16.0005
R5301 two_stage_opamp_dummy_magic_19_0.V_source.n10 two_stage_opamp_dummy_magic_19_0.V_source.t2 16.0005
R5302 two_stage_opamp_dummy_magic_19_0.V_source.n8 two_stage_opamp_dummy_magic_19_0.V_source.t8 16.0005
R5303 two_stage_opamp_dummy_magic_19_0.V_source.n8 two_stage_opamp_dummy_magic_19_0.V_source.t11 16.0005
R5304 two_stage_opamp_dummy_magic_19_0.V_source.n6 two_stage_opamp_dummy_magic_19_0.V_source.t5 16.0005
R5305 two_stage_opamp_dummy_magic_19_0.V_source.n6 two_stage_opamp_dummy_magic_19_0.V_source.t14 16.0005
R5306 two_stage_opamp_dummy_magic_19_0.V_source.n4 two_stage_opamp_dummy_magic_19_0.V_source.t40 16.0005
R5307 two_stage_opamp_dummy_magic_19_0.V_source.n4 two_stage_opamp_dummy_magic_19_0.V_source.t12 16.0005
R5308 two_stage_opamp_dummy_magic_19_0.V_source.n3 two_stage_opamp_dummy_magic_19_0.V_source.t0 16.0005
R5309 two_stage_opamp_dummy_magic_19_0.V_source.n3 two_stage_opamp_dummy_magic_19_0.V_source.t13 16.0005
R5310 two_stage_opamp_dummy_magic_19_0.V_source.n2 two_stage_opamp_dummy_magic_19_0.V_source.t16 16.0005
R5311 two_stage_opamp_dummy_magic_19_0.V_source.n2 two_stage_opamp_dummy_magic_19_0.V_source.t4 16.0005
R5312 two_stage_opamp_dummy_magic_19_0.V_source.n35 two_stage_opamp_dummy_magic_19_0.V_source.t35 9.6005
R5313 two_stage_opamp_dummy_magic_19_0.V_source.n35 two_stage_opamp_dummy_magic_19_0.V_source.t25 9.6005
R5314 two_stage_opamp_dummy_magic_19_0.V_source.n33 two_stage_opamp_dummy_magic_19_0.V_source.t31 9.6005
R5315 two_stage_opamp_dummy_magic_19_0.V_source.n33 two_stage_opamp_dummy_magic_19_0.V_source.t23 9.6005
R5316 two_stage_opamp_dummy_magic_19_0.V_source.n31 two_stage_opamp_dummy_magic_19_0.V_source.t34 9.6005
R5317 two_stage_opamp_dummy_magic_19_0.V_source.n31 two_stage_opamp_dummy_magic_19_0.V_source.t24 9.6005
R5318 two_stage_opamp_dummy_magic_19_0.V_source.n29 two_stage_opamp_dummy_magic_19_0.V_source.t30 9.6005
R5319 two_stage_opamp_dummy_magic_19_0.V_source.n29 two_stage_opamp_dummy_magic_19_0.V_source.t20 9.6005
R5320 two_stage_opamp_dummy_magic_19_0.V_source.n27 two_stage_opamp_dummy_magic_19_0.V_source.t28 9.6005
R5321 two_stage_opamp_dummy_magic_19_0.V_source.n27 two_stage_opamp_dummy_magic_19_0.V_source.t36 9.6005
R5322 two_stage_opamp_dummy_magic_19_0.V_source.n26 two_stage_opamp_dummy_magic_19_0.V_source.t26 9.6005
R5323 two_stage_opamp_dummy_magic_19_0.V_source.n26 two_stage_opamp_dummy_magic_19_0.V_source.t32 9.6005
R5324 two_stage_opamp_dummy_magic_19_0.V_source.n24 two_stage_opamp_dummy_magic_19_0.V_source.t22 9.6005
R5325 two_stage_opamp_dummy_magic_19_0.V_source.n24 two_stage_opamp_dummy_magic_19_0.V_source.t29 9.6005
R5326 two_stage_opamp_dummy_magic_19_0.V_source.n21 two_stage_opamp_dummy_magic_19_0.V_source.t21 9.6005
R5327 two_stage_opamp_dummy_magic_19_0.V_source.n21 two_stage_opamp_dummy_magic_19_0.V_source.t33 9.6005
R5328 two_stage_opamp_dummy_magic_19_0.V_source.n0 two_stage_opamp_dummy_magic_19_0.V_source.t38 9.6005
R5329 two_stage_opamp_dummy_magic_19_0.V_source.n0 two_stage_opamp_dummy_magic_19_0.V_source.t17 9.6005
R5330 two_stage_opamp_dummy_magic_19_0.V_source.t37 two_stage_opamp_dummy_magic_19_0.V_source.n38 9.6005
R5331 two_stage_opamp_dummy_magic_19_0.V_source.n38 two_stage_opamp_dummy_magic_19_0.V_source.t27 9.6005
R5332 two_stage_opamp_dummy_magic_19_0.V_source.n22 two_stage_opamp_dummy_magic_19_0.V_source.n20 4.67758
R5333 two_stage_opamp_dummy_magic_19_0.V_source.n19 two_stage_opamp_dummy_magic_19_0.V_source.n18 4.6255
R5334 two_stage_opamp_dummy_magic_19_0.V_source.n20 two_stage_opamp_dummy_magic_19_0.V_source.n19 4.5005
R5335 two_stage_opamp_dummy_magic_19_0.V_source.n23 two_stage_opamp_dummy_magic_19_0.V_source.n22 4.5005
R5336 two_stage_opamp_dummy_magic_19_0.V_source.n30 two_stage_opamp_dummy_magic_19_0.V_source.n28 0.563
R5337 two_stage_opamp_dummy_magic_19_0.V_source.n32 two_stage_opamp_dummy_magic_19_0.V_source.n30 0.563
R5338 two_stage_opamp_dummy_magic_19_0.V_source.n34 two_stage_opamp_dummy_magic_19_0.V_source.n32 0.563
R5339 two_stage_opamp_dummy_magic_19_0.V_source.n36 two_stage_opamp_dummy_magic_19_0.V_source.n34 0.563
R5340 two_stage_opamp_dummy_magic_19_0.V_source.n37 two_stage_opamp_dummy_magic_19_0.V_source.n36 0.563
R5341 two_stage_opamp_dummy_magic_19_0.V_source.n14 two_stage_opamp_dummy_magic_19_0.V_source.n12 0.563
R5342 two_stage_opamp_dummy_magic_19_0.V_source.n16 two_stage_opamp_dummy_magic_19_0.V_source.n14 0.563
R5343 two_stage_opamp_dummy_magic_19_0.V_source.n18 two_stage_opamp_dummy_magic_19_0.V_source.n16 0.563
R5344 two_stage_opamp_dummy_magic_19_0.V_source.n7 two_stage_opamp_dummy_magic_19_0.V_source.n5 0.563
R5345 two_stage_opamp_dummy_magic_19_0.V_source.n9 two_stage_opamp_dummy_magic_19_0.V_source.n7 0.563
R5346 two_stage_opamp_dummy_magic_19_0.V_source.n19 two_stage_opamp_dummy_magic_19_0.V_source.n9 0.563
R5347 two_stage_opamp_dummy_magic_19_0.V_source.n23 two_stage_opamp_dummy_magic_19_0.V_source.n1 0.563
R5348 two_stage_opamp_dummy_magic_19_0.V_source.n25 two_stage_opamp_dummy_magic_19_0.V_source.n23 0.563
R5349 two_stage_opamp_dummy_magic_19_0.V_source.n37 two_stage_opamp_dummy_magic_19_0.V_source.n25 0.563
R5350 VOUT+.n5 VOUT+.t10 112.159
R5351 VOUT+.n15 VOUT+.n14 41.431
R5352 VOUT+.n9 VOUT+.n7 41.431
R5353 VOUT+.n13 VOUT+.n12 40.8685
R5354 VOUT+.n11 VOUT+.n10 40.8685
R5355 VOUT+.n9 VOUT+.n8 40.8685
R5356 VOUT+.n16 VOUT+.n6 36.3685
R5357 VOUT+.n2 VOUT+.n0 16.9483
R5358 VOUT+.n4 VOUT+.n3 15.8233
R5359 VOUT+.n2 VOUT+.n1 15.8233
R5360 VOUT+.n91 VOUT+.n16 15.063
R5361 VOUT+.n91 VOUT+.n90 11.5649
R5362 VOUT+ VOUT+.n91 9.28175
R5363 VOUT+.n14 VOUT+.t5 6.56717
R5364 VOUT+.n14 VOUT+.t16 6.56717
R5365 VOUT+.n12 VOUT+.t9 6.56717
R5366 VOUT+.n12 VOUT+.t18 6.56717
R5367 VOUT+.n10 VOUT+.t0 6.56717
R5368 VOUT+.n10 VOUT+.t6 6.56717
R5369 VOUT+.n8 VOUT+.t12 6.56717
R5370 VOUT+.n8 VOUT+.t8 6.56717
R5371 VOUT+.n7 VOUT+.t15 6.56717
R5372 VOUT+.n7 VOUT+.t7 6.56717
R5373 VOUT+.n6 VOUT+.t4 6.56717
R5374 VOUT+.n6 VOUT+.t3 6.56717
R5375 VOUT+.n45 VOUT+.t56 4.8295
R5376 VOUT+.n47 VOUT+.t105 4.8295
R5377 VOUT+.n48 VOUT+.t29 4.8295
R5378 VOUT+.n50 VOUT+.t60 4.8295
R5379 VOUT+.n52 VOUT+.t115 4.8295
R5380 VOUT+.n63 VOUT+.t20 4.8295
R5381 VOUT+.n66 VOUT+.t31 4.8295
R5382 VOUT+.n65 VOUT+.t121 4.8295
R5383 VOUT+.n68 VOUT+.t67 4.8295
R5384 VOUT+.n67 VOUT+.t152 4.8295
R5385 VOUT+.n69 VOUT+.t131 4.8295
R5386 VOUT+.n70 VOUT+.t118 4.8295
R5387 VOUT+.n72 VOUT+.t89 4.8295
R5388 VOUT+.n73 VOUT+.t76 4.8295
R5389 VOUT+.n75 VOUT+.t127 4.8295
R5390 VOUT+.n76 VOUT+.t110 4.8295
R5391 VOUT+.n78 VOUT+.t84 4.8295
R5392 VOUT+.n79 VOUT+.t68 4.8295
R5393 VOUT+.n81 VOUT+.t42 4.8295
R5394 VOUT+.n82 VOUT+.t30 4.8295
R5395 VOUT+.n84 VOUT+.t81 4.8295
R5396 VOUT+.n85 VOUT+.t64 4.8295
R5397 VOUT+.n17 VOUT+.t150 4.8295
R5398 VOUT+.n28 VOUT+.t75 4.8295
R5399 VOUT+.n30 VOUT+.t54 4.8295
R5400 VOUT+.n31 VOUT+.t34 4.8295
R5401 VOUT+.n33 VOUT+.t95 4.8295
R5402 VOUT+.n34 VOUT+.t79 4.8295
R5403 VOUT+.n36 VOUT+.t134 4.8295
R5404 VOUT+.n37 VOUT+.t122 4.8295
R5405 VOUT+.n39 VOUT+.t102 4.8295
R5406 VOUT+.n40 VOUT+.t82 4.8295
R5407 VOUT+.n42 VOUT+.t137 4.8295
R5408 VOUT+.n43 VOUT+.t126 4.8295
R5409 VOUT+.n87 VOUT+.t28 4.8295
R5410 VOUT+.n56 VOUT+.t57 4.8154
R5411 VOUT+.n55 VOUT+.t33 4.8154
R5412 VOUT+.n54 VOUT+.t77 4.8154
R5413 VOUT+.n62 VOUT+.t116 4.806
R5414 VOUT+.n61 VOUT+.t147 4.806
R5415 VOUT+.n60 VOUT+.t43 4.806
R5416 VOUT+.n59 VOUT+.t83 4.806
R5417 VOUT+.n58 VOUT+.t63 4.806
R5418 VOUT+.n57 VOUT+.t26 4.806
R5419 VOUT+.n57 VOUT+.t103 4.806
R5420 VOUT+.n56 VOUT+.t135 4.806
R5421 VOUT+.n55 VOUT+.t120 4.806
R5422 VOUT+.n54 VOUT+.t155 4.806
R5423 VOUT+.n27 VOUT+.t91 4.806
R5424 VOUT+.n26 VOUT+.t38 4.806
R5425 VOUT+.n25 VOUT+.t130 4.806
R5426 VOUT+.n25 VOUT+.t90 4.806
R5427 VOUT+.n24 VOUT+.t80 4.806
R5428 VOUT+.n24 VOUT+.t128 4.806
R5429 VOUT+.n23 VOUT+.t124 4.806
R5430 VOUT+.n23 VOUT+.t32 4.806
R5431 VOUT+.n22 VOUT+.t70 4.806
R5432 VOUT+.n22 VOUT+.t73 4.806
R5433 VOUT+.n21 VOUT+.t23 4.806
R5434 VOUT+.n21 VOUT+.t108 4.806
R5435 VOUT+.n20 VOUT+.t62 4.806
R5436 VOUT+.n20 VOUT+.t19 4.806
R5437 VOUT+.n19 VOUT+.t151 4.806
R5438 VOUT+.n19 VOUT+.t49 4.806
R5439 VOUT+.n46 VOUT+.t132 4.5005
R5440 VOUT+.n45 VOUT+.t96 4.5005
R5441 VOUT+.n47 VOUT+.t69 4.5005
R5442 VOUT+.n48 VOUT+.t139 4.5005
R5443 VOUT+.n49 VOUT+.t109 4.5005
R5444 VOUT+.n50 VOUT+.t37 4.5005
R5445 VOUT+.n51 VOUT+.t144 4.5005
R5446 VOUT+.n52 VOUT+.t21 4.5005
R5447 VOUT+.n53 VOUT+.t125 4.5005
R5448 VOUT+.n54 VOUT+.t119 4.5005
R5449 VOUT+.n55 VOUT+.t78 4.5005
R5450 VOUT+.n56 VOUT+.t97 4.5005
R5451 VOUT+.n57 VOUT+.t61 4.5005
R5452 VOUT+.n58 VOUT+.t27 4.5005
R5453 VOUT+.n59 VOUT+.t41 4.5005
R5454 VOUT+.n60 VOUT+.t145 4.5005
R5455 VOUT+.n61 VOUT+.t113 4.5005
R5456 VOUT+.n62 VOUT+.t72 4.5005
R5457 VOUT+.n64 VOUT+.t92 4.5005
R5458 VOUT+.n63 VOUT+.t55 4.5005
R5459 VOUT+.n66 VOUT+.t50 4.5005
R5460 VOUT+.n65 VOUT+.t156 4.5005
R5461 VOUT+.n68 VOUT+.t86 4.5005
R5462 VOUT+.n67 VOUT+.t47 4.5005
R5463 VOUT+.n69 VOUT+.t94 4.5005
R5464 VOUT+.n71 VOUT+.t39 4.5005
R5465 VOUT+.n70 VOUT+.t146 4.5005
R5466 VOUT+.n72 VOUT+.t53 4.5005
R5467 VOUT+.n74 VOUT+.t142 4.5005
R5468 VOUT+.n73 VOUT+.t112 4.5005
R5469 VOUT+.n75 VOUT+.t88 4.5005
R5470 VOUT+.n77 VOUT+.t35 4.5005
R5471 VOUT+.n76 VOUT+.t140 4.5005
R5472 VOUT+.n78 VOUT+.t46 4.5005
R5473 VOUT+.n80 VOUT+.t136 4.5005
R5474 VOUT+.n79 VOUT+.t104 4.5005
R5475 VOUT+.n81 VOUT+.t149 4.5005
R5476 VOUT+.n83 VOUT+.t99 4.5005
R5477 VOUT+.n82 VOUT+.t65 4.5005
R5478 VOUT+.n84 VOUT+.t40 4.5005
R5479 VOUT+.n86 VOUT+.t133 4.5005
R5480 VOUT+.n85 VOUT+.t98 4.5005
R5481 VOUT+.n18 VOUT+.t45 4.5005
R5482 VOUT+.n17 VOUT+.t101 4.5005
R5483 VOUT+.n19 VOUT+.t85 4.5005
R5484 VOUT+.n20 VOUT+.t48 4.5005
R5485 VOUT+.n21 VOUT+.t138 4.5005
R5486 VOUT+.n22 VOUT+.t107 4.5005
R5487 VOUT+.n23 VOUT+.t71 4.5005
R5488 VOUT+.n24 VOUT+.t25 4.5005
R5489 VOUT+.n25 VOUT+.t129 4.5005
R5490 VOUT+.n26 VOUT+.t87 4.5005
R5491 VOUT+.n27 VOUT+.t52 4.5005
R5492 VOUT+.n29 VOUT+.t141 4.5005
R5493 VOUT+.n28 VOUT+.t111 4.5005
R5494 VOUT+.n30 VOUT+.t24 4.5005
R5495 VOUT+.n32 VOUT+.t114 4.5005
R5496 VOUT+.n31 VOUT+.t74 4.5005
R5497 VOUT+.n33 VOUT+.t59 4.5005
R5498 VOUT+.n35 VOUT+.t148 4.5005
R5499 VOUT+.n34 VOUT+.t117 4.5005
R5500 VOUT+.n36 VOUT+.t100 4.5005
R5501 VOUT+.n38 VOUT+.t44 4.5005
R5502 VOUT+.n37 VOUT+.t153 4.5005
R5503 VOUT+.n39 VOUT+.t66 4.5005
R5504 VOUT+.n41 VOUT+.t154 4.5005
R5505 VOUT+.n40 VOUT+.t123 4.5005
R5506 VOUT+.n42 VOUT+.t106 4.5005
R5507 VOUT+.n44 VOUT+.t51 4.5005
R5508 VOUT+.n43 VOUT+.t22 4.5005
R5509 VOUT+.n90 VOUT+.t36 4.5005
R5510 VOUT+.n89 VOUT+.t143 4.5005
R5511 VOUT+.n88 VOUT+.t93 4.5005
R5512 VOUT+.n87 VOUT+.t58 4.5005
R5513 VOUT+.n16 VOUT+.n15 4.5005
R5514 VOUT+.n3 VOUT+.t2 3.42907
R5515 VOUT+.n3 VOUT+.t14 3.42907
R5516 VOUT+.n1 VOUT+.t17 3.42907
R5517 VOUT+.n1 VOUT+.t11 3.42907
R5518 VOUT+.n0 VOUT+.t13 3.42907
R5519 VOUT+.n0 VOUT+.t1 3.42907
R5520 VOUT+.n5 VOUT+.n4 1.30519
R5521 VOUT+.n4 VOUT+.n2 1.1255
R5522 VOUT+ VOUT+.n5 0.961438
R5523 VOUT+.n11 VOUT+.n9 0.563
R5524 VOUT+.n13 VOUT+.n11 0.563
R5525 VOUT+.n15 VOUT+.n13 0.563
R5526 VOUT+.n46 VOUT+.n45 0.3295
R5527 VOUT+.n49 VOUT+.n48 0.3295
R5528 VOUT+.n51 VOUT+.n50 0.3295
R5529 VOUT+.n53 VOUT+.n52 0.3295
R5530 VOUT+.n55 VOUT+.n54 0.3295
R5531 VOUT+.n56 VOUT+.n55 0.3295
R5532 VOUT+.n57 VOUT+.n56 0.3295
R5533 VOUT+.n58 VOUT+.n57 0.3295
R5534 VOUT+.n59 VOUT+.n58 0.3295
R5535 VOUT+.n60 VOUT+.n59 0.3295
R5536 VOUT+.n61 VOUT+.n60 0.3295
R5537 VOUT+.n62 VOUT+.n61 0.3295
R5538 VOUT+.n64 VOUT+.n62 0.3295
R5539 VOUT+.n64 VOUT+.n63 0.3295
R5540 VOUT+.n66 VOUT+.n65 0.3295
R5541 VOUT+.n68 VOUT+.n67 0.3295
R5542 VOUT+.n71 VOUT+.n69 0.3295
R5543 VOUT+.n71 VOUT+.n70 0.3295
R5544 VOUT+.n74 VOUT+.n72 0.3295
R5545 VOUT+.n74 VOUT+.n73 0.3295
R5546 VOUT+.n77 VOUT+.n75 0.3295
R5547 VOUT+.n77 VOUT+.n76 0.3295
R5548 VOUT+.n80 VOUT+.n78 0.3295
R5549 VOUT+.n80 VOUT+.n79 0.3295
R5550 VOUT+.n83 VOUT+.n81 0.3295
R5551 VOUT+.n83 VOUT+.n82 0.3295
R5552 VOUT+.n86 VOUT+.n84 0.3295
R5553 VOUT+.n86 VOUT+.n85 0.3295
R5554 VOUT+.n18 VOUT+.n17 0.3295
R5555 VOUT+.n20 VOUT+.n19 0.3295
R5556 VOUT+.n21 VOUT+.n20 0.3295
R5557 VOUT+.n22 VOUT+.n21 0.3295
R5558 VOUT+.n23 VOUT+.n22 0.3295
R5559 VOUT+.n24 VOUT+.n23 0.3295
R5560 VOUT+.n25 VOUT+.n24 0.3295
R5561 VOUT+.n26 VOUT+.n25 0.3295
R5562 VOUT+.n27 VOUT+.n26 0.3295
R5563 VOUT+.n29 VOUT+.n27 0.3295
R5564 VOUT+.n29 VOUT+.n28 0.3295
R5565 VOUT+.n32 VOUT+.n30 0.3295
R5566 VOUT+.n32 VOUT+.n31 0.3295
R5567 VOUT+.n35 VOUT+.n33 0.3295
R5568 VOUT+.n35 VOUT+.n34 0.3295
R5569 VOUT+.n38 VOUT+.n36 0.3295
R5570 VOUT+.n38 VOUT+.n37 0.3295
R5571 VOUT+.n41 VOUT+.n39 0.3295
R5572 VOUT+.n41 VOUT+.n40 0.3295
R5573 VOUT+.n44 VOUT+.n42 0.3295
R5574 VOUT+.n44 VOUT+.n43 0.3295
R5575 VOUT+.n90 VOUT+.n89 0.3295
R5576 VOUT+.n89 VOUT+.n88 0.3295
R5577 VOUT+.n88 VOUT+.n87 0.3295
R5578 VOUT+.n61 VOUT+.n47 0.306
R5579 VOUT+.n60 VOUT+.n49 0.306
R5580 VOUT+.n59 VOUT+.n51 0.306
R5581 VOUT+.n58 VOUT+.n53 0.306
R5582 VOUT+.n64 VOUT+.n46 0.2825
R5583 VOUT+.n66 VOUT+.n64 0.2825
R5584 VOUT+.n68 VOUT+.n66 0.2825
R5585 VOUT+.n71 VOUT+.n68 0.2825
R5586 VOUT+.n74 VOUT+.n71 0.2825
R5587 VOUT+.n77 VOUT+.n74 0.2825
R5588 VOUT+.n80 VOUT+.n77 0.2825
R5589 VOUT+.n83 VOUT+.n80 0.2825
R5590 VOUT+.n86 VOUT+.n83 0.2825
R5591 VOUT+.n29 VOUT+.n18 0.2825
R5592 VOUT+.n32 VOUT+.n29 0.2825
R5593 VOUT+.n35 VOUT+.n32 0.2825
R5594 VOUT+.n38 VOUT+.n35 0.2825
R5595 VOUT+.n41 VOUT+.n38 0.2825
R5596 VOUT+.n44 VOUT+.n41 0.2825
R5597 VOUT+.n88 VOUT+.n44 0.2825
R5598 VOUT+.n88 VOUT+.n86 0.2825
R5599 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t127 50.3211
R5600 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t101 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t136 0.1603
R5601 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t60 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t100 0.1603
R5602 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t35 0.1603
R5603 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t109 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t4 0.1603
R5604 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t10 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t38 0.1603
R5605 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t62 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t25 0.1603
R5606 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t80 0.1603
R5607 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t103 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t67 0.1603
R5608 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t46 0.1603
R5609 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t68 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t29 0.1603
R5610 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t52 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t88 0.1603
R5611 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t110 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t72 0.1603
R5612 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t91 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t126 0.1603
R5613 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t7 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t114 0.1603
R5614 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t58 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t92 0.1603
R5615 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t116 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t75 0.1603
R5616 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t98 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t128 0.1603
R5617 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t13 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t120 0.1603
R5618 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t134 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t30 0.1603
R5619 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t50 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t19 0.1603
R5620 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t33 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t74 0.1603
R5621 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t90 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t54 0.1603
R5622 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t3 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t34 0.1603
R5623 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t56 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t22 0.1603
R5624 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t39 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t77 0.1603
R5625 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t97 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t61 0.1603
R5626 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t82 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t122 0.1603
R5627 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t132 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t102 0.1603
R5628 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t45 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t81 0.1603
R5629 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t71 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t5 0.1603
R5630 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t108 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t94 0.1603
R5631 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t18 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t133 0.1603
R5632 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t49 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t86 0.1603
R5633 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t85 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t32 0.1603
R5634 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t131 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t76 0.1603
R5635 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t27 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t26 0.1603
R5636 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t69 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t118 0.1603
R5637 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t104 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t65 0.1603
R5638 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t55 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t6 0.1603
R5639 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t87 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t51 0.1603
R5640 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t43 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t87 0.1603
R5641 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t37 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t79 0.1603
R5642 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t78 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t123 0.1603
R5643 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t99 0.1603
R5644 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t95 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t130 0.1603
R5645 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t135 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t41 0.1603
R5646 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t31 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t135 0.1603
R5647 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t129 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t31 0.1603
R5648 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t119 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t96 0.1603
R5649 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t12 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t119 0.1603
R5650 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t115 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t12 0.1603
R5651 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t47 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t11 0.1603
R5652 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t17 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t47 0.1603
R5653 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t127 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t17 0.1603
R5654 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t24 0.159278
R5655 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t107 0.159278
R5656 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t137 0.159278
R5657 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t48 0.159278
R5658 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t83 0.159278
R5659 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t124 0.159278
R5660 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t28 0.159278
R5661 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t66 0.159278
R5662 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t15 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n15 0.159278
R5663 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t42 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n16 0.159278
R5664 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t8 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n17 0.159278
R5665 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t112 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n18 0.159278
R5666 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t2 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n19 0.159278
R5667 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t105 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n20 0.159278
R5668 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t63 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n21 0.159278
R5669 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t23 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n22 0.159278
R5670 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t57 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n23 0.159278
R5671 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t20 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n24 0.159278
R5672 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t121 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n25 0.159278
R5673 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t14 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n26 0.159278
R5674 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t117 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n27 0.159278
R5675 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t70 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n28 0.159278
R5676 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t106 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n29 0.159278
R5677 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t64 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n30 0.159278
R5678 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t40 0.159278
R5679 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t9 0.159278
R5680 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t1 0.159278
R5681 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t36 0.159278
R5682 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t21 0.159278
R5683 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t53 0.159278
R5684 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t93 0.159278
R5685 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t73 0.159278
R5686 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t113 0.159278
R5687 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t24 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t60 0.137822
R5688 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t101 0.1368
R5689 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t0 0.1368
R5690 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t125 0.1368
R5691 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t109 0.1368
R5692 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t89 0.1368
R5693 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t10 0.1368
R5694 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t62 0.1368
R5695 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t44 0.1368
R5696 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t103 0.1368
R5697 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t16 0.1368
R5698 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t68 0.1368
R5699 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t52 0.1368
R5700 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t110 0.1368
R5701 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t91 0.1368
R5702 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t7 0.1368
R5703 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t58 0.1368
R5704 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t116 0.1368
R5705 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t98 0.1368
R5706 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t13 0.1368
R5707 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t134 0.1368
R5708 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t50 0.1368
R5709 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t33 0.1368
R5710 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t90 0.1368
R5711 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t3 0.1368
R5712 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t56 0.1368
R5713 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t39 0.1368
R5714 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t97 0.1368
R5715 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t82 0.1368
R5716 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t132 0.1368
R5717 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t45 0.1368
R5718 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t55 0.1368
R5719 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n6 0.1133
R5720 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n7 0.1133
R5721 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n8 0.1133
R5722 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n9 0.1133
R5723 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n10 0.1133
R5724 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n11 0.1133
R5725 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n12 0.1133
R5726 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n13 0.1133
R5727 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n14 0.1133
R5728 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n31 0.1133
R5729 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n32 0.1133
R5730 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n0 0.1133
R5731 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n1 0.1133
R5732 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n2 0.1133
R5733 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n3 0.1133
R5734 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n4 0.1133
R5735 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n5 0.1133
R5736 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n33 0.1133
R5737 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t71 0.00152174
R5738 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t108 0.00152174
R5739 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t18 0.00152174
R5740 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t49 0.00152174
R5741 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t85 0.00152174
R5742 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t131 0.00152174
R5743 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t27 0.00152174
R5744 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t69 0.00152174
R5745 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t104 0.00152174
R5746 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t111 0.00152174
R5747 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t15 0.00152174
R5748 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t42 0.00152174
R5749 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t8 0.00152174
R5750 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t112 0.00152174
R5751 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t2 0.00152174
R5752 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t105 0.00152174
R5753 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t63 0.00152174
R5754 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t23 0.00152174
R5755 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t57 0.00152174
R5756 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t20 0.00152174
R5757 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t121 0.00152174
R5758 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t14 0.00152174
R5759 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t117 0.00152174
R5760 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t70 0.00152174
R5761 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t106 0.00152174
R5762 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t64 0.00152174
R5763 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t84 0.00152174
R5764 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t43 0.00152174
R5765 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t37 0.00152174
R5766 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t78 0.00152174
R5767 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t59 0.00152174
R5768 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t95 0.00152174
R5769 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t129 0.00152174
R5770 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t115 0.00152174
R5771 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t11 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n34 0.00152174
R5772 two_stage_opamp_dummy_magic_19_0.X.n57 two_stage_opamp_dummy_magic_19_0.X.t48 1172.87
R5773 two_stage_opamp_dummy_magic_19_0.X.n53 two_stage_opamp_dummy_magic_19_0.X.t43 1172.87
R5774 two_stage_opamp_dummy_magic_19_0.X.n57 two_stage_opamp_dummy_magic_19_0.X.t35 996.134
R5775 two_stage_opamp_dummy_magic_19_0.X.n58 two_stage_opamp_dummy_magic_19_0.X.t51 996.134
R5776 two_stage_opamp_dummy_magic_19_0.X.n59 two_stage_opamp_dummy_magic_19_0.X.t39 996.134
R5777 two_stage_opamp_dummy_magic_19_0.X.n60 two_stage_opamp_dummy_magic_19_0.X.t31 996.134
R5778 two_stage_opamp_dummy_magic_19_0.X.n56 two_stage_opamp_dummy_magic_19_0.X.t46 996.134
R5779 two_stage_opamp_dummy_magic_19_0.X.n55 two_stage_opamp_dummy_magic_19_0.X.t33 996.134
R5780 two_stage_opamp_dummy_magic_19_0.X.n54 two_stage_opamp_dummy_magic_19_0.X.t50 996.134
R5781 two_stage_opamp_dummy_magic_19_0.X.n53 two_stage_opamp_dummy_magic_19_0.X.t28 996.134
R5782 two_stage_opamp_dummy_magic_19_0.X.n45 two_stage_opamp_dummy_magic_19_0.X.t25 690.867
R5783 two_stage_opamp_dummy_magic_19_0.X.n42 two_stage_opamp_dummy_magic_19_0.X.t47 690.867
R5784 two_stage_opamp_dummy_magic_19_0.X.n36 two_stage_opamp_dummy_magic_19_0.X.t36 530.201
R5785 two_stage_opamp_dummy_magic_19_0.X.n33 two_stage_opamp_dummy_magic_19_0.X.t30 530.201
R5786 two_stage_opamp_dummy_magic_19_0.X.n49 two_stage_opamp_dummy_magic_19_0.X.t54 514.134
R5787 two_stage_opamp_dummy_magic_19_0.X.n48 two_stage_opamp_dummy_magic_19_0.X.t37 514.134
R5788 two_stage_opamp_dummy_magic_19_0.X.n47 two_stage_opamp_dummy_magic_19_0.X.t44 514.134
R5789 two_stage_opamp_dummy_magic_19_0.X.n46 two_stage_opamp_dummy_magic_19_0.X.t29 514.134
R5790 two_stage_opamp_dummy_magic_19_0.X.n45 two_stage_opamp_dummy_magic_19_0.X.t42 514.134
R5791 two_stage_opamp_dummy_magic_19_0.X.n42 two_stage_opamp_dummy_magic_19_0.X.t32 514.134
R5792 two_stage_opamp_dummy_magic_19_0.X.n43 two_stage_opamp_dummy_magic_19_0.X.t27 514.134
R5793 two_stage_opamp_dummy_magic_19_0.X.n44 two_stage_opamp_dummy_magic_19_0.X.t41 514.134
R5794 two_stage_opamp_dummy_magic_19_0.X.n62 two_stage_opamp_dummy_magic_19_0.X.n61 424.875
R5795 two_stage_opamp_dummy_magic_19_0.X.n36 two_stage_opamp_dummy_magic_19_0.X.t53 353.467
R5796 two_stage_opamp_dummy_magic_19_0.X.n37 two_stage_opamp_dummy_magic_19_0.X.t40 353.467
R5797 two_stage_opamp_dummy_magic_19_0.X.n38 two_stage_opamp_dummy_magic_19_0.X.t26 353.467
R5798 two_stage_opamp_dummy_magic_19_0.X.n39 two_stage_opamp_dummy_magic_19_0.X.t49 353.467
R5799 two_stage_opamp_dummy_magic_19_0.X.n40 two_stage_opamp_dummy_magic_19_0.X.t34 353.467
R5800 two_stage_opamp_dummy_magic_19_0.X.n35 two_stage_opamp_dummy_magic_19_0.X.t52 353.467
R5801 two_stage_opamp_dummy_magic_19_0.X.n34 two_stage_opamp_dummy_magic_19_0.X.t38 353.467
R5802 two_stage_opamp_dummy_magic_19_0.X.n33 two_stage_opamp_dummy_magic_19_0.X.t45 353.467
R5803 two_stage_opamp_dummy_magic_19_0.X.n56 two_stage_opamp_dummy_magic_19_0.X.n55 176.733
R5804 two_stage_opamp_dummy_magic_19_0.X.n55 two_stage_opamp_dummy_magic_19_0.X.n54 176.733
R5805 two_stage_opamp_dummy_magic_19_0.X.n54 two_stage_opamp_dummy_magic_19_0.X.n53 176.733
R5806 two_stage_opamp_dummy_magic_19_0.X.n58 two_stage_opamp_dummy_magic_19_0.X.n57 176.733
R5807 two_stage_opamp_dummy_magic_19_0.X.n59 two_stage_opamp_dummy_magic_19_0.X.n58 176.733
R5808 two_stage_opamp_dummy_magic_19_0.X.n60 two_stage_opamp_dummy_magic_19_0.X.n59 176.733
R5809 two_stage_opamp_dummy_magic_19_0.X.n35 two_stage_opamp_dummy_magic_19_0.X.n34 176.733
R5810 two_stage_opamp_dummy_magic_19_0.X.n34 two_stage_opamp_dummy_magic_19_0.X.n33 176.733
R5811 two_stage_opamp_dummy_magic_19_0.X.n37 two_stage_opamp_dummy_magic_19_0.X.n36 176.733
R5812 two_stage_opamp_dummy_magic_19_0.X.n38 two_stage_opamp_dummy_magic_19_0.X.n37 176.733
R5813 two_stage_opamp_dummy_magic_19_0.X.n39 two_stage_opamp_dummy_magic_19_0.X.n38 176.733
R5814 two_stage_opamp_dummy_magic_19_0.X.n40 two_stage_opamp_dummy_magic_19_0.X.n39 176.733
R5815 two_stage_opamp_dummy_magic_19_0.X.n44 two_stage_opamp_dummy_magic_19_0.X.n43 176.733
R5816 two_stage_opamp_dummy_magic_19_0.X.n43 two_stage_opamp_dummy_magic_19_0.X.n42 176.733
R5817 two_stage_opamp_dummy_magic_19_0.X.n46 two_stage_opamp_dummy_magic_19_0.X.n45 176.733
R5818 two_stage_opamp_dummy_magic_19_0.X.n47 two_stage_opamp_dummy_magic_19_0.X.n46 176.733
R5819 two_stage_opamp_dummy_magic_19_0.X.n48 two_stage_opamp_dummy_magic_19_0.X.n47 176.733
R5820 two_stage_opamp_dummy_magic_19_0.X.n49 two_stage_opamp_dummy_magic_19_0.X.n48 176.733
R5821 two_stage_opamp_dummy_magic_19_0.X.n52 two_stage_opamp_dummy_magic_19_0.X.n51 174.769
R5822 two_stage_opamp_dummy_magic_19_0.X.n51 two_stage_opamp_dummy_magic_19_0.X.n41 162.675
R5823 two_stage_opamp_dummy_magic_19_0.X.n51 two_stage_opamp_dummy_magic_19_0.X.n50 162.675
R5824 two_stage_opamp_dummy_magic_19_0.X.n6 two_stage_opamp_dummy_magic_19_0.X.n4 72.013
R5825 two_stage_opamp_dummy_magic_19_0.X.n3 two_stage_opamp_dummy_magic_19_0.X.n1 72.013
R5826 two_stage_opamp_dummy_magic_19_0.X.n8 two_stage_opamp_dummy_magic_19_0.X.n7 71.388
R5827 two_stage_opamp_dummy_magic_19_0.X.n6 two_stage_opamp_dummy_magic_19_0.X.n5 71.388
R5828 two_stage_opamp_dummy_magic_19_0.X.n3 two_stage_opamp_dummy_magic_19_0.X.n2 71.388
R5829 two_stage_opamp_dummy_magic_19_0.X.n10 two_stage_opamp_dummy_magic_19_0.X.n0 66.888
R5830 two_stage_opamp_dummy_magic_19_0.X.n61 two_stage_opamp_dummy_magic_19_0.X.n56 56.2338
R5831 two_stage_opamp_dummy_magic_19_0.X.n61 two_stage_opamp_dummy_magic_19_0.X.n60 56.2338
R5832 two_stage_opamp_dummy_magic_19_0.X.n41 two_stage_opamp_dummy_magic_19_0.X.n35 56.2338
R5833 two_stage_opamp_dummy_magic_19_0.X.n41 two_stage_opamp_dummy_magic_19_0.X.n40 56.2338
R5834 two_stage_opamp_dummy_magic_19_0.X.n50 two_stage_opamp_dummy_magic_19_0.X.n44 56.2338
R5835 two_stage_opamp_dummy_magic_19_0.X.n50 two_stage_opamp_dummy_magic_19_0.X.n49 56.2338
R5836 two_stage_opamp_dummy_magic_19_0.X.t17 two_stage_opamp_dummy_magic_19_0.X.n62 49.8023
R5837 two_stage_opamp_dummy_magic_19_0.X.n14 two_stage_opamp_dummy_magic_19_0.X.n13 49.3505
R5838 two_stage_opamp_dummy_magic_19_0.X.n17 two_stage_opamp_dummy_magic_19_0.X.n16 49.3505
R5839 two_stage_opamp_dummy_magic_19_0.X.n20 two_stage_opamp_dummy_magic_19_0.X.n19 49.3505
R5840 two_stage_opamp_dummy_magic_19_0.X.n24 two_stage_opamp_dummy_magic_19_0.X.n23 49.3505
R5841 two_stage_opamp_dummy_magic_19_0.X.n27 two_stage_opamp_dummy_magic_19_0.X.n26 49.3505
R5842 two_stage_opamp_dummy_magic_19_0.X.n30 two_stage_opamp_dummy_magic_19_0.X.n29 49.3505
R5843 two_stage_opamp_dummy_magic_19_0.X.n32 two_stage_opamp_dummy_magic_19_0.X.n10 17.688
R5844 two_stage_opamp_dummy_magic_19_0.X.n13 two_stage_opamp_dummy_magic_19_0.X.t0 16.0005
R5845 two_stage_opamp_dummy_magic_19_0.X.n13 two_stage_opamp_dummy_magic_19_0.X.t19 16.0005
R5846 two_stage_opamp_dummy_magic_19_0.X.n16 two_stage_opamp_dummy_magic_19_0.X.t5 16.0005
R5847 two_stage_opamp_dummy_magic_19_0.X.n16 two_stage_opamp_dummy_magic_19_0.X.t14 16.0005
R5848 two_stage_opamp_dummy_magic_19_0.X.n19 two_stage_opamp_dummy_magic_19_0.X.t24 16.0005
R5849 two_stage_opamp_dummy_magic_19_0.X.n19 two_stage_opamp_dummy_magic_19_0.X.t1 16.0005
R5850 two_stage_opamp_dummy_magic_19_0.X.n23 two_stage_opamp_dummy_magic_19_0.X.t15 16.0005
R5851 two_stage_opamp_dummy_magic_19_0.X.n23 two_stage_opamp_dummy_magic_19_0.X.t16 16.0005
R5852 two_stage_opamp_dummy_magic_19_0.X.n26 two_stage_opamp_dummy_magic_19_0.X.t6 16.0005
R5853 two_stage_opamp_dummy_magic_19_0.X.n26 two_stage_opamp_dummy_magic_19_0.X.t23 16.0005
R5854 two_stage_opamp_dummy_magic_19_0.X.n29 two_stage_opamp_dummy_magic_19_0.X.t18 16.0005
R5855 two_stage_opamp_dummy_magic_19_0.X.n29 two_stage_opamp_dummy_magic_19_0.X.t4 16.0005
R5856 two_stage_opamp_dummy_magic_19_0.X.n7 two_stage_opamp_dummy_magic_19_0.X.t20 11.2576
R5857 two_stage_opamp_dummy_magic_19_0.X.n7 two_stage_opamp_dummy_magic_19_0.X.t8 11.2576
R5858 two_stage_opamp_dummy_magic_19_0.X.n5 two_stage_opamp_dummy_magic_19_0.X.t7 11.2576
R5859 two_stage_opamp_dummy_magic_19_0.X.n5 two_stage_opamp_dummy_magic_19_0.X.t11 11.2576
R5860 two_stage_opamp_dummy_magic_19_0.X.n4 two_stage_opamp_dummy_magic_19_0.X.t10 11.2576
R5861 two_stage_opamp_dummy_magic_19_0.X.n4 two_stage_opamp_dummy_magic_19_0.X.t9 11.2576
R5862 two_stage_opamp_dummy_magic_19_0.X.n2 two_stage_opamp_dummy_magic_19_0.X.t2 11.2576
R5863 two_stage_opamp_dummy_magic_19_0.X.n2 two_stage_opamp_dummy_magic_19_0.X.t22 11.2576
R5864 two_stage_opamp_dummy_magic_19_0.X.n1 two_stage_opamp_dummy_magic_19_0.X.t12 11.2576
R5865 two_stage_opamp_dummy_magic_19_0.X.n1 two_stage_opamp_dummy_magic_19_0.X.t21 11.2576
R5866 two_stage_opamp_dummy_magic_19_0.X.n0 two_stage_opamp_dummy_magic_19_0.X.t13 11.2576
R5867 two_stage_opamp_dummy_magic_19_0.X.n0 two_stage_opamp_dummy_magic_19_0.X.t3 11.2576
R5868 two_stage_opamp_dummy_magic_19_0.X.n62 two_stage_opamp_dummy_magic_19_0.X.n52 7.09425
R5869 two_stage_opamp_dummy_magic_19_0.X.n32 two_stage_opamp_dummy_magic_19_0.X.n31 6.3755
R5870 two_stage_opamp_dummy_magic_19_0.X.n15 two_stage_opamp_dummy_magic_19_0.X.n14 5.71404
R5871 two_stage_opamp_dummy_magic_19_0.X.n30 two_stage_opamp_dummy_magic_19_0.X.n28 5.71404
R5872 two_stage_opamp_dummy_magic_19_0.X.n18 two_stage_opamp_dummy_magic_19_0.X.n14 5.5005
R5873 two_stage_opamp_dummy_magic_19_0.X.n17 two_stage_opamp_dummy_magic_19_0.X.n15 5.10988
R5874 two_stage_opamp_dummy_magic_19_0.X.n20 two_stage_opamp_dummy_magic_19_0.X.n12 5.10988
R5875 two_stage_opamp_dummy_magic_19_0.X.n25 two_stage_opamp_dummy_magic_19_0.X.n24 5.10988
R5876 two_stage_opamp_dummy_magic_19_0.X.n28 two_stage_opamp_dummy_magic_19_0.X.n27 5.10988
R5877 two_stage_opamp_dummy_magic_19_0.X.n18 two_stage_opamp_dummy_magic_19_0.X.n17 4.938
R5878 two_stage_opamp_dummy_magic_19_0.X.n21 two_stage_opamp_dummy_magic_19_0.X.n20 4.938
R5879 two_stage_opamp_dummy_magic_19_0.X.n24 two_stage_opamp_dummy_magic_19_0.X.n22 4.938
R5880 two_stage_opamp_dummy_magic_19_0.X.n27 two_stage_opamp_dummy_magic_19_0.X.n11 4.938
R5881 two_stage_opamp_dummy_magic_19_0.X.n31 two_stage_opamp_dummy_magic_19_0.X.n30 4.938
R5882 two_stage_opamp_dummy_magic_19_0.X.n10 two_stage_opamp_dummy_magic_19_0.X.n9 4.5005
R5883 two_stage_opamp_dummy_magic_19_0.X.n52 two_stage_opamp_dummy_magic_19_0.X.n32 1.03175
R5884 two_stage_opamp_dummy_magic_19_0.X.n8 two_stage_opamp_dummy_magic_19_0.X.n6 0.6255
R5885 two_stage_opamp_dummy_magic_19_0.X.n9 two_stage_opamp_dummy_magic_19_0.X.n8 0.6255
R5886 two_stage_opamp_dummy_magic_19_0.X.n9 two_stage_opamp_dummy_magic_19_0.X.n3 0.6255
R5887 two_stage_opamp_dummy_magic_19_0.X.n28 two_stage_opamp_dummy_magic_19_0.X.n25 0.604667
R5888 two_stage_opamp_dummy_magic_19_0.X.n25 two_stage_opamp_dummy_magic_19_0.X.n12 0.604667
R5889 two_stage_opamp_dummy_magic_19_0.X.n15 two_stage_opamp_dummy_magic_19_0.X.n12 0.604667
R5890 two_stage_opamp_dummy_magic_19_0.X.n21 two_stage_opamp_dummy_magic_19_0.X.n18 0.563
R5891 two_stage_opamp_dummy_magic_19_0.X.n22 two_stage_opamp_dummy_magic_19_0.X.n21 0.563
R5892 two_stage_opamp_dummy_magic_19_0.X.n22 two_stage_opamp_dummy_magic_19_0.X.n11 0.563
R5893 two_stage_opamp_dummy_magic_19_0.X.n31 two_stage_opamp_dummy_magic_19_0.X.n11 0.563
R5894 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n0 150.451
R5895 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n1 140.201
R5896 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t10 118.861
R5897 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n2 37.4067
R5898 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n12 33.83
R5899 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n3 30.038
R5900 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n10 29.4755
R5901 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n8 29.4755
R5902 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n6 29.4755
R5903 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n4 29.4755
R5904 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t11 24.0005
R5905 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t12 24.0005
R5906 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t13 24.0005
R5907 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t14 24.0005
R5908 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t9 8.0005
R5909 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t3 8.0005
R5910 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t7 8.0005
R5911 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t2 8.0005
R5912 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t5 8.0005
R5913 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t0 8.0005
R5914 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t4 8.0005
R5915 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t8 8.0005
R5916 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t6 8.0005
R5917 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t1 8.0005
R5918 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n11 5.6255
R5919 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n5 0.563
R5920 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n7 0.563
R5921 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n9 0.563
R5922 bgr_9_0.V_CMFB_S2 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n13 0.047375
R5923 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t11 688.859
R5924 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t8 651.384
R5925 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t9 648.072
R5926 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n2 514.134
R5927 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n4 214.056
R5928 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t7 174.726
R5929 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t13 174.726
R5930 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t10 174.726
R5931 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t12 174.726
R5932 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n6 173.149
R5933 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n9 168.774
R5934 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n7 168.774
R5935 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n1 128.534
R5936 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n3 128.534
R5937 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t0 125.736
R5938 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n11 46.6411
R5939 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t3 13.1338
R5940 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t1 13.1338
R5941 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t6 13.1338
R5942 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t4 13.1338
R5943 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t2 13.1338
R5944 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t5 13.1338
R5945 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n10 10.0317
R5946 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n8 4.3755
R5947 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n5 3.03175
R5948 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n0 1.53175
R5949 two_stage_opamp_dummy_magic_19_0.err_amp_out.n1 two_stage_opamp_dummy_magic_19_0.err_amp_out.t4 857.505
R5950 two_stage_opamp_dummy_magic_19_0.err_amp_out.n1 two_stage_opamp_dummy_magic_19_0.err_amp_out.n0 105.519
R5951 two_stage_opamp_dummy_magic_19_0.err_amp_out.n2 two_stage_opamp_dummy_magic_19_0.err_amp_out.n1 39.4984
R5952 two_stage_opamp_dummy_magic_19_0.err_amp_out.n0 two_stage_opamp_dummy_magic_19_0.err_amp_out.t3 15.7605
R5953 two_stage_opamp_dummy_magic_19_0.err_amp_out.n0 two_stage_opamp_dummy_magic_19_0.err_amp_out.t0 15.7605
R5954 two_stage_opamp_dummy_magic_19_0.err_amp_out.n2 two_stage_opamp_dummy_magic_19_0.err_amp_out.t2 9.6005
R5955 two_stage_opamp_dummy_magic_19_0.err_amp_out.t1 two_stage_opamp_dummy_magic_19_0.err_amp_out.n2 9.6005
R5956 bgr_9_0.Vin+.n3 bgr_9_0.Vin+.n2 526.183
R5957 bgr_9_0.Vin+.n1 bgr_9_0.Vin+.n0 514.134
R5958 bgr_9_0.Vin+.n0 bgr_9_0.Vin+.t8 303.259
R5959 bgr_9_0.Vin+.n5 bgr_9_0.Vin+.n3 227.169
R5960 bgr_9_0.Vin+.n0 bgr_9_0.Vin+.t9 174.726
R5961 bgr_9_0.Vin+.n1 bgr_9_0.Vin+.t6 174.726
R5962 bgr_9_0.Vin+.n2 bgr_9_0.Vin+.t10 174.726
R5963 bgr_9_0.Vin+.n7 bgr_9_0.Vin+.n6 167.993
R5964 bgr_9_0.Vin+.n5 bgr_9_0.Vin+.n4 167.993
R5965 bgr_9_0.Vin+.t0 bgr_9_0.Vin+.n8 158.989
R5966 bgr_9_0.Vin+.n2 bgr_9_0.Vin+.n1 128.534
R5967 bgr_9_0.Vin+.n8 bgr_9_0.Vin+.t1 119.067
R5968 bgr_9_0.Vin+.n3 bgr_9_0.Vin+.t7 96.4005
R5969 bgr_9_0.Vin+.n8 bgr_9_0.Vin+.n7 35.0317
R5970 bgr_9_0.Vin+.n6 bgr_9_0.Vin+.t2 13.1338
R5971 bgr_9_0.Vin+.n6 bgr_9_0.Vin+.t5 13.1338
R5972 bgr_9_0.Vin+.n4 bgr_9_0.Vin+.t4 13.1338
R5973 bgr_9_0.Vin+.n4 bgr_9_0.Vin+.t3 13.1338
R5974 bgr_9_0.Vin+.n7 bgr_9_0.Vin+.n5 2.1255
R5975 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n0 344.837
R5976 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n1 344.274
R5977 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n3 292.5
R5978 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n5 124.403
R5979 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n12 123.84
R5980 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n10 123.84
R5981 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n8 123.84
R5982 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n6 123.84
R5983 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t15 120.43
R5984 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n2 52.3363
R5985 bgr_9_0.V_CMFB_S1 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n4 52.1563
R5986 bgr_9_0.V_CMFB_S1 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n14 41.1227
R5987 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t0 39.4005
R5988 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t13 39.4005
R5989 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t1 39.4005
R5990 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t16 39.4005
R5991 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t14 39.4005
R5992 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t2 39.4005
R5993 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t9 19.7005
R5994 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t3 19.7005
R5995 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t7 19.7005
R5996 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t12 19.7005
R5997 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t5 19.7005
R5998 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t10 19.7005
R5999 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t4 19.7005
R6000 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t8 19.7005
R6001 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t6 19.7005
R6002 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t11 19.7005
R6003 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n13 5.90675
R6004 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n7 0.563
R6005 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n9 0.563
R6006 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n11 0.563
R6007 bgr_9_0.V_mir1.n13 bgr_9_0.V_mir1.n12 330.901
R6008 bgr_9_0.V_mir1.n4 bgr_9_0.V_mir1.n3 330.901
R6009 bgr_9_0.V_mir1.n20 bgr_9_0.V_mir1.n19 330.901
R6010 bgr_9_0.V_mir1.n16 bgr_9_0.V_mir1.t19 310.488
R6011 bgr_9_0.V_mir1.n9 bgr_9_0.V_mir1.t21 310.488
R6012 bgr_9_0.V_mir1.n0 bgr_9_0.V_mir1.t20 310.488
R6013 bgr_9_0.V_mir1.n7 bgr_9_0.V_mir1.t15 278.312
R6014 bgr_9_0.V_mir1.n7 bgr_9_0.V_mir1.n6 228.939
R6015 bgr_9_0.V_mir1.n8 bgr_9_0.V_mir1.n5 224.439
R6016 bgr_9_0.V_mir1.n18 bgr_9_0.V_mir1.t7 184.097
R6017 bgr_9_0.V_mir1.n11 bgr_9_0.V_mir1.t3 184.097
R6018 bgr_9_0.V_mir1.n2 bgr_9_0.V_mir1.t1 184.097
R6019 bgr_9_0.V_mir1.n17 bgr_9_0.V_mir1.n16 167.094
R6020 bgr_9_0.V_mir1.n10 bgr_9_0.V_mir1.n9 167.094
R6021 bgr_9_0.V_mir1.n1 bgr_9_0.V_mir1.n0 167.094
R6022 bgr_9_0.V_mir1.n13 bgr_9_0.V_mir1.n11 152
R6023 bgr_9_0.V_mir1.n4 bgr_9_0.V_mir1.n2 152
R6024 bgr_9_0.V_mir1.n19 bgr_9_0.V_mir1.n18 152
R6025 bgr_9_0.V_mir1.n16 bgr_9_0.V_mir1.t22 120.501
R6026 bgr_9_0.V_mir1.n17 bgr_9_0.V_mir1.t11 120.501
R6027 bgr_9_0.V_mir1.n9 bgr_9_0.V_mir1.t17 120.501
R6028 bgr_9_0.V_mir1.n10 bgr_9_0.V_mir1.t9 120.501
R6029 bgr_9_0.V_mir1.n0 bgr_9_0.V_mir1.t18 120.501
R6030 bgr_9_0.V_mir1.n1 bgr_9_0.V_mir1.t5 120.501
R6031 bgr_9_0.V_mir1.n6 bgr_9_0.V_mir1.t0 48.0005
R6032 bgr_9_0.V_mir1.n6 bgr_9_0.V_mir1.t14 48.0005
R6033 bgr_9_0.V_mir1.n5 bgr_9_0.V_mir1.t13 48.0005
R6034 bgr_9_0.V_mir1.n5 bgr_9_0.V_mir1.t16 48.0005
R6035 bgr_9_0.V_mir1.n18 bgr_9_0.V_mir1.n17 40.7027
R6036 bgr_9_0.V_mir1.n11 bgr_9_0.V_mir1.n10 40.7027
R6037 bgr_9_0.V_mir1.n2 bgr_9_0.V_mir1.n1 40.7027
R6038 bgr_9_0.V_mir1.n12 bgr_9_0.V_mir1.t4 39.4005
R6039 bgr_9_0.V_mir1.n12 bgr_9_0.V_mir1.t10 39.4005
R6040 bgr_9_0.V_mir1.n3 bgr_9_0.V_mir1.t2 39.4005
R6041 bgr_9_0.V_mir1.n3 bgr_9_0.V_mir1.t6 39.4005
R6042 bgr_9_0.V_mir1.n20 bgr_9_0.V_mir1.t8 39.4005
R6043 bgr_9_0.V_mir1.t12 bgr_9_0.V_mir1.n20 39.4005
R6044 bgr_9_0.V_mir1.n15 bgr_9_0.V_mir1.n4 15.8005
R6045 bgr_9_0.V_mir1.n19 bgr_9_0.V_mir1.n15 15.8005
R6046 bgr_9_0.V_mir1.n14 bgr_9_0.V_mir1.n13 9.3005
R6047 bgr_9_0.V_mir1.n8 bgr_9_0.V_mir1.n7 5.8755
R6048 bgr_9_0.V_mir1.n15 bgr_9_0.V_mir1.n14 4.5005
R6049 bgr_9_0.V_mir1.n14 bgr_9_0.V_mir1.n8 0.78175
R6050 bgr_9_0.1st_Vout_1 bgr_9_0.1st_Vout_1.t13 354.854
R6051 bgr_9_0.1st_Vout_1.n5 bgr_9_0.1st_Vout_1.t21 346.8
R6052 bgr_9_0.1st_Vout_1.n20 bgr_9_0.1st_Vout_1.n19 344.95
R6053 bgr_9_0.1st_Vout_1.n7 bgr_9_0.1st_Vout_1.n6 344.95
R6054 bgr_9_0.1st_Vout_1.n15 bgr_9_0.1st_Vout_1.n14 340.45
R6055 bgr_9_0.1st_Vout_1.n11 bgr_9_0.1st_Vout_1.t10 275.909
R6056 bgr_9_0.1st_Vout_1.n11 bgr_9_0.1st_Vout_1.n10 227.909
R6057 bgr_9_0.1st_Vout_1.n13 bgr_9_0.1st_Vout_1.n12 222.034
R6058 bgr_9_0.1st_Vout_1.n17 bgr_9_0.1st_Vout_1.t22 184.097
R6059 bgr_9_0.1st_Vout_1.n17 bgr_9_0.1st_Vout_1.t32 184.097
R6060 bgr_9_0.1st_Vout_1.n8 bgr_9_0.1st_Vout_1.t16 184.097
R6061 bgr_9_0.1st_Vout_1.n8 bgr_9_0.1st_Vout_1.t36 184.097
R6062 bgr_9_0.1st_Vout_1.n18 bgr_9_0.1st_Vout_1.n17 166.05
R6063 bgr_9_0.1st_Vout_1.n9 bgr_9_0.1st_Vout_1.n8 166.05
R6064 bgr_9_0.1st_Vout_1.n5 bgr_9_0.1st_Vout_1.n4 54.2759
R6065 bgr_9_0.1st_Vout_1.n12 bgr_9_0.1st_Vout_1.t7 48.0005
R6066 bgr_9_0.1st_Vout_1.n12 bgr_9_0.1st_Vout_1.t6 48.0005
R6067 bgr_9_0.1st_Vout_1.n10 bgr_9_0.1st_Vout_1.t8 48.0005
R6068 bgr_9_0.1st_Vout_1.n10 bgr_9_0.1st_Vout_1.t9 48.0005
R6069 bgr_9_0.1st_Vout_1.n19 bgr_9_0.1st_Vout_1.t4 39.4005
R6070 bgr_9_0.1st_Vout_1.n19 bgr_9_0.1st_Vout_1.t2 39.4005
R6071 bgr_9_0.1st_Vout_1.n6 bgr_9_0.1st_Vout_1.t0 39.4005
R6072 bgr_9_0.1st_Vout_1.n6 bgr_9_0.1st_Vout_1.t3 39.4005
R6073 bgr_9_0.1st_Vout_1.n14 bgr_9_0.1st_Vout_1.t5 39.4005
R6074 bgr_9_0.1st_Vout_1.n14 bgr_9_0.1st_Vout_1.t1 39.4005
R6075 bgr_9_0.1st_Vout_1.n0 bgr_9_0.1st_Vout_1.t11 4.8295
R6076 bgr_9_0.1st_Vout_1.n0 bgr_9_0.1st_Vout_1.t29 4.8295
R6077 bgr_9_0.1st_Vout_1.n2 bgr_9_0.1st_Vout_1.t31 4.8295
R6078 bgr_9_0.1st_Vout_1.n1 bgr_9_0.1st_Vout_1.t20 4.8295
R6079 bgr_9_0.1st_Vout_1.n2 bgr_9_0.1st_Vout_1.t24 4.8295
R6080 bgr_9_0.1st_Vout_1.n2 bgr_9_0.1st_Vout_1.t14 4.8295
R6081 bgr_9_0.1st_Vout_1.n3 bgr_9_0.1st_Vout_1.t30 4.8295
R6082 bgr_9_0.1st_Vout_1.n3 bgr_9_0.1st_Vout_1.t18 4.8295
R6083 bgr_9_0.1st_Vout_1.n3 bgr_9_0.1st_Vout_1.t23 4.8295
R6084 bgr_9_0.1st_Vout_1.n0 bgr_9_0.1st_Vout_1.t15 4.5005
R6085 bgr_9_0.1st_Vout_1.n0 bgr_9_0.1st_Vout_1.t35 4.5005
R6086 bgr_9_0.1st_Vout_1.n2 bgr_9_0.1st_Vout_1.t34 4.5005
R6087 bgr_9_0.1st_Vout_1.n1 bgr_9_0.1st_Vout_1.t28 4.5005
R6088 bgr_9_0.1st_Vout_1.n2 bgr_9_0.1st_Vout_1.t27 4.5005
R6089 bgr_9_0.1st_Vout_1.n2 bgr_9_0.1st_Vout_1.t19 4.5005
R6090 bgr_9_0.1st_Vout_1.n3 bgr_9_0.1st_Vout_1.t33 4.5005
R6091 bgr_9_0.1st_Vout_1.n3 bgr_9_0.1st_Vout_1.t26 4.5005
R6092 bgr_9_0.1st_Vout_1.n3 bgr_9_0.1st_Vout_1.t25 4.5005
R6093 bgr_9_0.1st_Vout_1.n4 bgr_9_0.1st_Vout_1.t17 4.5005
R6094 bgr_9_0.1st_Vout_1.n4 bgr_9_0.1st_Vout_1.t12 4.5005
R6095 bgr_9_0.1st_Vout_1.n13 bgr_9_0.1st_Vout_1.n11 4.5005
R6096 bgr_9_0.1st_Vout_1.n16 bgr_9_0.1st_Vout_1.n15 4.5005
R6097 bgr_9_0.1st_Vout_1.n20 bgr_9_0.1st_Vout_1.n18 1.3755
R6098 bgr_9_0.1st_Vout_1.n16 bgr_9_0.1st_Vout_1.n9 1.3755
R6099 bgr_9_0.1st_Vout_1.n7 bgr_9_0.1st_Vout_1.n5 1.188
R6100 bgr_9_0.1st_Vout_1.n3 bgr_9_0.1st_Vout_1.n2 0.8935
R6101 bgr_9_0.1st_Vout_1.n2 bgr_9_0.1st_Vout_1.n0 0.8935
R6102 bgr_9_0.1st_Vout_1.n15 bgr_9_0.1st_Vout_1.n13 0.78175
R6103 bgr_9_0.1st_Vout_1.n4 bgr_9_0.1st_Vout_1.n3 0.6585
R6104 bgr_9_0.1st_Vout_1.n2 bgr_9_0.1st_Vout_1.n1 0.6585
R6105 bgr_9_0.1st_Vout_1.n18 bgr_9_0.1st_Vout_1.n16 0.6255
R6106 bgr_9_0.1st_Vout_1.n9 bgr_9_0.1st_Vout_1.n7 0.6255
R6107 bgr_9_0.1st_Vout_1 bgr_9_0.1st_Vout_1.n20 0.438
R6108 bgr_9_0.1st_Vout_2.n1 bgr_9_0.1st_Vout_2.t33 355.293
R6109 bgr_9_0.1st_Vout_2.n0 bgr_9_0.1st_Vout_2.t34 346.8
R6110 bgr_9_0.1st_Vout_2.n0 bgr_9_0.1st_Vout_2.n10 344.95
R6111 bgr_9_0.1st_Vout_2.n1 bgr_9_0.1st_Vout_2.n8 344.95
R6112 bgr_9_0.1st_Vout_2.n12 bgr_9_0.1st_Vout_2.n3 340.45
R6113 bgr_9_0.1st_Vout_2.n6 bgr_9_0.1st_Vout_2.t0 275.909
R6114 bgr_9_0.1st_Vout_2.n6 bgr_9_0.1st_Vout_2.n5 227.909
R6115 bgr_9_0.1st_Vout_2.n3 bgr_9_0.1st_Vout_2.n7 222.034
R6116 bgr_9_0.1st_Vout_2.n11 bgr_9_0.1st_Vout_2.t16 184.097
R6117 bgr_9_0.1st_Vout_2.n11 bgr_9_0.1st_Vout_2.t27 184.097
R6118 bgr_9_0.1st_Vout_2.n9 bgr_9_0.1st_Vout_2.t13 184.097
R6119 bgr_9_0.1st_Vout_2.n9 bgr_9_0.1st_Vout_2.t24 184.097
R6120 bgr_9_0.1st_Vout_2.n0 bgr_9_0.1st_Vout_2.n11 166.05
R6121 bgr_9_0.1st_Vout_2.n1 bgr_9_0.1st_Vout_2.n9 166.05
R6122 bgr_9_0.1st_Vout_2.n0 bgr_9_0.1st_Vout_2.n4 52.9634
R6123 bgr_9_0.1st_Vout_2.n7 bgr_9_0.1st_Vout_2.t1 48.0005
R6124 bgr_9_0.1st_Vout_2.n7 bgr_9_0.1st_Vout_2.t2 48.0005
R6125 bgr_9_0.1st_Vout_2.n5 bgr_9_0.1st_Vout_2.t8 48.0005
R6126 bgr_9_0.1st_Vout_2.n5 bgr_9_0.1st_Vout_2.t4 48.0005
R6127 bgr_9_0.1st_Vout_2.n10 bgr_9_0.1st_Vout_2.t7 39.4005
R6128 bgr_9_0.1st_Vout_2.n10 bgr_9_0.1st_Vout_2.t9 39.4005
R6129 bgr_9_0.1st_Vout_2.n8 bgr_9_0.1st_Vout_2.t10 39.4005
R6130 bgr_9_0.1st_Vout_2.n8 bgr_9_0.1st_Vout_2.t5 39.4005
R6131 bgr_9_0.1st_Vout_2.n12 bgr_9_0.1st_Vout_2.t6 39.4005
R6132 bgr_9_0.1st_Vout_2.t3 bgr_9_0.1st_Vout_2.n12 39.4005
R6133 bgr_9_0.1st_Vout_2.n3 bgr_9_0.1st_Vout_2.n1 5.28175
R6134 bgr_9_0.1st_Vout_2.n1 bgr_9_0.1st_Vout_2.n0 5.188
R6135 bgr_9_0.1st_Vout_2.n2 bgr_9_0.1st_Vout_2.t17 4.8295
R6136 bgr_9_0.1st_Vout_2.n2 bgr_9_0.1st_Vout_2.t35 4.8295
R6137 bgr_9_0.1st_Vout_2.n2 bgr_9_0.1st_Vout_2.t11 4.8295
R6138 bgr_9_0.1st_Vout_2.n2 bgr_9_0.1st_Vout_2.t26 4.8295
R6139 bgr_9_0.1st_Vout_2.n2 bgr_9_0.1st_Vout_2.t30 4.8295
R6140 bgr_9_0.1st_Vout_2.n2 bgr_9_0.1st_Vout_2.t19 4.8295
R6141 bgr_9_0.1st_Vout_2.n4 bgr_9_0.1st_Vout_2.t36 4.8295
R6142 bgr_9_0.1st_Vout_2.n4 bgr_9_0.1st_Vout_2.t25 4.8295
R6143 bgr_9_0.1st_Vout_2.n4 bgr_9_0.1st_Vout_2.t18 4.8295
R6144 bgr_9_0.1st_Vout_2.n2 bgr_9_0.1st_Vout_2.t12 4.5005
R6145 bgr_9_0.1st_Vout_2.n2 bgr_9_0.1st_Vout_2.t32 4.5005
R6146 bgr_9_0.1st_Vout_2.n2 bgr_9_0.1st_Vout_2.t31 4.5005
R6147 bgr_9_0.1st_Vout_2.n2 bgr_9_0.1st_Vout_2.t23 4.5005
R6148 bgr_9_0.1st_Vout_2.n2 bgr_9_0.1st_Vout_2.t22 4.5005
R6149 bgr_9_0.1st_Vout_2.n2 bgr_9_0.1st_Vout_2.t15 4.5005
R6150 bgr_9_0.1st_Vout_2.n4 bgr_9_0.1st_Vout_2.t29 4.5005
R6151 bgr_9_0.1st_Vout_2.n4 bgr_9_0.1st_Vout_2.t21 4.5005
R6152 bgr_9_0.1st_Vout_2.n4 bgr_9_0.1st_Vout_2.t28 4.5005
R6153 bgr_9_0.1st_Vout_2.n4 bgr_9_0.1st_Vout_2.t20 4.5005
R6154 bgr_9_0.1st_Vout_2.n4 bgr_9_0.1st_Vout_2.t14 4.5005
R6155 bgr_9_0.1st_Vout_2.n3 bgr_9_0.1st_Vout_2.n6 4.5005
R6156 bgr_9_0.1st_Vout_2.n4 bgr_9_0.1st_Vout_2.n2 3.1025
R6157 bgr_9_0.cap_res2.t20 bgr_9_0.cap_res2.t17 121.245
R6158 bgr_9_0.cap_res2.t12 bgr_9_0.cap_res2.t6 0.1603
R6159 bgr_9_0.cap_res2.t5 bgr_9_0.cap_res2.t0 0.1603
R6160 bgr_9_0.cap_res2.t10 bgr_9_0.cap_res2.t4 0.1603
R6161 bgr_9_0.cap_res2.t3 bgr_9_0.cap_res2.t19 0.1603
R6162 bgr_9_0.cap_res2.t18 bgr_9_0.cap_res2.t15 0.1603
R6163 bgr_9_0.cap_res2.n1 bgr_9_0.cap_res2.t2 0.159278
R6164 bgr_9_0.cap_res2.n2 bgr_9_0.cap_res2.t9 0.159278
R6165 bgr_9_0.cap_res2.n3 bgr_9_0.cap_res2.t16 0.159278
R6166 bgr_9_0.cap_res2.n4 bgr_9_0.cap_res2.t11 0.159278
R6167 bgr_9_0.cap_res2.n4 bgr_9_0.cap_res2.t14 0.1368
R6168 bgr_9_0.cap_res2.n4 bgr_9_0.cap_res2.t12 0.1368
R6169 bgr_9_0.cap_res2.n3 bgr_9_0.cap_res2.t8 0.1368
R6170 bgr_9_0.cap_res2.n3 bgr_9_0.cap_res2.t5 0.1368
R6171 bgr_9_0.cap_res2.n2 bgr_9_0.cap_res2.t13 0.1368
R6172 bgr_9_0.cap_res2.n2 bgr_9_0.cap_res2.t10 0.1368
R6173 bgr_9_0.cap_res2.n1 bgr_9_0.cap_res2.t7 0.1368
R6174 bgr_9_0.cap_res2.n1 bgr_9_0.cap_res2.t3 0.1368
R6175 bgr_9_0.cap_res2.n0 bgr_9_0.cap_res2.t1 0.1368
R6176 bgr_9_0.cap_res2.n0 bgr_9_0.cap_res2.t18 0.1368
R6177 bgr_9_0.cap_res2.t2 bgr_9_0.cap_res2.n0 0.00152174
R6178 bgr_9_0.cap_res2.t9 bgr_9_0.cap_res2.n1 0.00152174
R6179 bgr_9_0.cap_res2.t16 bgr_9_0.cap_res2.n2 0.00152174
R6180 bgr_9_0.cap_res2.t11 bgr_9_0.cap_res2.n3 0.00152174
R6181 bgr_9_0.cap_res2.t17 bgr_9_0.cap_res2.n4 0.00152174
R6182 two_stage_opamp_dummy_magic_19_0.Vb2.n21 two_stage_opamp_dummy_magic_19_0.Vb2.t16 650.273
R6183 two_stage_opamp_dummy_magic_19_0.Vb2.n1 two_stage_opamp_dummy_magic_19_0.Vb2.t1 650.273
R6184 two_stage_opamp_dummy_magic_19_0.Vb2.n16 two_stage_opamp_dummy_magic_19_0.Vb2.t23 611.739
R6185 two_stage_opamp_dummy_magic_19_0.Vb2.n11 two_stage_opamp_dummy_magic_19_0.Vb2.t12 611.739
R6186 two_stage_opamp_dummy_magic_19_0.Vb2.n5 two_stage_opamp_dummy_magic_19_0.Vb2.t24 611.739
R6187 two_stage_opamp_dummy_magic_19_0.Vb2.n3 two_stage_opamp_dummy_magic_19_0.Vb2.t13 611.739
R6188 two_stage_opamp_dummy_magic_19_0.Vb2.n18 two_stage_opamp_dummy_magic_19_0.Vb2.t14 463.925
R6189 two_stage_opamp_dummy_magic_19_0.Vb2.n10 two_stage_opamp_dummy_magic_19_0.Vb2.t22 463.925
R6190 two_stage_opamp_dummy_magic_19_0.Vb2.n2 two_stage_opamp_dummy_magic_19_0.Vb2.t28 445.423
R6191 two_stage_opamp_dummy_magic_19_0.Vb2.n16 two_stage_opamp_dummy_magic_19_0.Vb2.t27 421.75
R6192 two_stage_opamp_dummy_magic_19_0.Vb2.n17 two_stage_opamp_dummy_magic_19_0.Vb2.t20 421.75
R6193 two_stage_opamp_dummy_magic_19_0.Vb2.n11 two_stage_opamp_dummy_magic_19_0.Vb2.t18 421.75
R6194 two_stage_opamp_dummy_magic_19_0.Vb2.n12 two_stage_opamp_dummy_magic_19_0.Vb2.t25 421.75
R6195 two_stage_opamp_dummy_magic_19_0.Vb2.n13 two_stage_opamp_dummy_magic_19_0.Vb2.t29 421.75
R6196 two_stage_opamp_dummy_magic_19_0.Vb2.n14 two_stage_opamp_dummy_magic_19_0.Vb2.t30 421.75
R6197 two_stage_opamp_dummy_magic_19_0.Vb2.n15 two_stage_opamp_dummy_magic_19_0.Vb2.t32 421.75
R6198 two_stage_opamp_dummy_magic_19_0.Vb2.n5 two_stage_opamp_dummy_magic_19_0.Vb2.t17 421.75
R6199 two_stage_opamp_dummy_magic_19_0.Vb2.n6 two_stage_opamp_dummy_magic_19_0.Vb2.t21 421.75
R6200 two_stage_opamp_dummy_magic_19_0.Vb2.n7 two_stage_opamp_dummy_magic_19_0.Vb2.t15 421.75
R6201 two_stage_opamp_dummy_magic_19_0.Vb2.n8 two_stage_opamp_dummy_magic_19_0.Vb2.t11 421.75
R6202 two_stage_opamp_dummy_magic_19_0.Vb2.n9 two_stage_opamp_dummy_magic_19_0.Vb2.t31 421.75
R6203 two_stage_opamp_dummy_magic_19_0.Vb2.n3 two_stage_opamp_dummy_magic_19_0.Vb2.t19 421.75
R6204 two_stage_opamp_dummy_magic_19_0.Vb2.n4 two_stage_opamp_dummy_magic_19_0.Vb2.t26 421.75
R6205 two_stage_opamp_dummy_magic_19_0.Vb2.n19 two_stage_opamp_dummy_magic_19_0.Vb2.n10 331.226
R6206 two_stage_opamp_dummy_magic_19_0.Vb2.n19 two_stage_opamp_dummy_magic_19_0.Vb2.n18 330.663
R6207 two_stage_opamp_dummy_magic_19_0.Vb2.n1 two_stage_opamp_dummy_magic_19_0.Vb2.n0 170.793
R6208 two_stage_opamp_dummy_magic_19_0.Vb2.n17 two_stage_opamp_dummy_magic_19_0.Vb2.n16 167.094
R6209 two_stage_opamp_dummy_magic_19_0.Vb2.n12 two_stage_opamp_dummy_magic_19_0.Vb2.n11 167.094
R6210 two_stage_opamp_dummy_magic_19_0.Vb2.n13 two_stage_opamp_dummy_magic_19_0.Vb2.n12 167.094
R6211 two_stage_opamp_dummy_magic_19_0.Vb2.n14 two_stage_opamp_dummy_magic_19_0.Vb2.n13 167.094
R6212 two_stage_opamp_dummy_magic_19_0.Vb2.n15 two_stage_opamp_dummy_magic_19_0.Vb2.n14 167.094
R6213 two_stage_opamp_dummy_magic_19_0.Vb2.n6 two_stage_opamp_dummy_magic_19_0.Vb2.n5 167.094
R6214 two_stage_opamp_dummy_magic_19_0.Vb2.n7 two_stage_opamp_dummy_magic_19_0.Vb2.n6 167.094
R6215 two_stage_opamp_dummy_magic_19_0.Vb2.n8 two_stage_opamp_dummy_magic_19_0.Vb2.n7 167.094
R6216 two_stage_opamp_dummy_magic_19_0.Vb2.n9 two_stage_opamp_dummy_magic_19_0.Vb2.n8 167.094
R6217 two_stage_opamp_dummy_magic_19_0.Vb2.n4 two_stage_opamp_dummy_magic_19_0.Vb2.n3 167.094
R6218 two_stage_opamp_dummy_magic_19_0.Vb2.n18 two_stage_opamp_dummy_magic_19_0.Vb2.n17 147.814
R6219 two_stage_opamp_dummy_magic_19_0.Vb2.n18 two_stage_opamp_dummy_magic_19_0.Vb2.n15 147.814
R6220 two_stage_opamp_dummy_magic_19_0.Vb2.n10 two_stage_opamp_dummy_magic_19_0.Vb2.n9 147.814
R6221 two_stage_opamp_dummy_magic_19_0.Vb2.n10 two_stage_opamp_dummy_magic_19_0.Vb2.n4 147.814
R6222 two_stage_opamp_dummy_magic_19_0.Vb2.n27 two_stage_opamp_dummy_magic_19_0.Vb2.n26 146.482
R6223 two_stage_opamp_dummy_magic_19_0.Vb2.n25 two_stage_opamp_dummy_magic_19_0.Vb2.n24 145.232
R6224 two_stage_opamp_dummy_magic_19_0.Vb2.n23 two_stage_opamp_dummy_magic_19_0.Vb2.n22 145.232
R6225 two_stage_opamp_dummy_magic_19_0.Vb2.n28 two_stage_opamp_dummy_magic_19_0.Vb2.n27 145.232
R6226 two_stage_opamp_dummy_magic_19_0.Vb2.n23 two_stage_opamp_dummy_magic_19_0.Vb2.n21 61.3224
R6227 two_stage_opamp_dummy_magic_19_0.Vb2.n26 two_stage_opamp_dummy_magic_19_0.Vb2.t7 24.0005
R6228 two_stage_opamp_dummy_magic_19_0.Vb2.n26 two_stage_opamp_dummy_magic_19_0.Vb2.t9 24.0005
R6229 two_stage_opamp_dummy_magic_19_0.Vb2.n24 two_stage_opamp_dummy_magic_19_0.Vb2.t5 24.0005
R6230 two_stage_opamp_dummy_magic_19_0.Vb2.n24 two_stage_opamp_dummy_magic_19_0.Vb2.t3 24.0005
R6231 two_stage_opamp_dummy_magic_19_0.Vb2.n22 two_stage_opamp_dummy_magic_19_0.Vb2.t10 24.0005
R6232 two_stage_opamp_dummy_magic_19_0.Vb2.n22 two_stage_opamp_dummy_magic_19_0.Vb2.t4 24.0005
R6233 two_stage_opamp_dummy_magic_19_0.Vb2.n28 two_stage_opamp_dummy_magic_19_0.Vb2.t6 24.0005
R6234 two_stage_opamp_dummy_magic_19_0.Vb2.t8 two_stage_opamp_dummy_magic_19_0.Vb2.n28 24.0005
R6235 two_stage_opamp_dummy_magic_19_0.Vb2.n20 two_stage_opamp_dummy_magic_19_0.Vb2.n19 12.8443
R6236 two_stage_opamp_dummy_magic_19_0.Vb2.n0 two_stage_opamp_dummy_magic_19_0.Vb2.t2 11.2576
R6237 two_stage_opamp_dummy_magic_19_0.Vb2.n0 two_stage_opamp_dummy_magic_19_0.Vb2.t0 11.2576
R6238 two_stage_opamp_dummy_magic_19_0.Vb2.n27 two_stage_opamp_dummy_magic_19_0.Vb2.n25 7.563
R6239 two_stage_opamp_dummy_magic_19_0.Vb2.n21 two_stage_opamp_dummy_magic_19_0.Vb2.n20 4.55362
R6240 two_stage_opamp_dummy_magic_19_0.Vb2.n2 two_stage_opamp_dummy_magic_19_0.Vb2.n1 2.84425
R6241 two_stage_opamp_dummy_magic_19_0.Vb2.n25 two_stage_opamp_dummy_magic_19_0.Vb2.n23 1.2505
R6242 two_stage_opamp_dummy_magic_19_0.Vb2.n20 two_stage_opamp_dummy_magic_19_0.Vb2.n2 0.928625
R6243 two_stage_opamp_dummy_magic_19_0.VD3.n16 two_stage_opamp_dummy_magic_19_0.VD3.t23 652.076
R6244 two_stage_opamp_dummy_magic_19_0.VD3.n19 two_stage_opamp_dummy_magic_19_0.VD3.t20 652.076
R6245 two_stage_opamp_dummy_magic_19_0.VD3.t24 two_stage_opamp_dummy_magic_19_0.VD3.n17 211.625
R6246 two_stage_opamp_dummy_magic_19_0.VD3.n18 two_stage_opamp_dummy_magic_19_0.VD3.t21 211.625
R6247 two_stage_opamp_dummy_magic_19_0.VD3.t4 two_stage_opamp_dummy_magic_19_0.VD3.t24 146.155
R6248 two_stage_opamp_dummy_magic_19_0.VD3.t12 two_stage_opamp_dummy_magic_19_0.VD3.t4 146.155
R6249 two_stage_opamp_dummy_magic_19_0.VD3.t8 two_stage_opamp_dummy_magic_19_0.VD3.t12 146.155
R6250 two_stage_opamp_dummy_magic_19_0.VD3.t14 two_stage_opamp_dummy_magic_19_0.VD3.t8 146.155
R6251 two_stage_opamp_dummy_magic_19_0.VD3.t18 two_stage_opamp_dummy_magic_19_0.VD3.t14 146.155
R6252 two_stage_opamp_dummy_magic_19_0.VD3.t0 two_stage_opamp_dummy_magic_19_0.VD3.t18 146.155
R6253 two_stage_opamp_dummy_magic_19_0.VD3.t6 two_stage_opamp_dummy_magic_19_0.VD3.t0 146.155
R6254 two_stage_opamp_dummy_magic_19_0.VD3.t2 two_stage_opamp_dummy_magic_19_0.VD3.t6 146.155
R6255 two_stage_opamp_dummy_magic_19_0.VD3.t10 two_stage_opamp_dummy_magic_19_0.VD3.t2 146.155
R6256 two_stage_opamp_dummy_magic_19_0.VD3.t16 two_stage_opamp_dummy_magic_19_0.VD3.t10 146.155
R6257 two_stage_opamp_dummy_magic_19_0.VD3.t21 two_stage_opamp_dummy_magic_19_0.VD3.t16 146.155
R6258 two_stage_opamp_dummy_magic_19_0.VD3.n17 two_stage_opamp_dummy_magic_19_0.VD3.t25 76.2576
R6259 two_stage_opamp_dummy_magic_19_0.VD3.n18 two_stage_opamp_dummy_magic_19_0.VD3.t22 76.2576
R6260 two_stage_opamp_dummy_magic_19_0.VD3.n4 two_stage_opamp_dummy_magic_19_0.VD3.n2 72.013
R6261 two_stage_opamp_dummy_magic_19_0.VD3.n1 two_stage_opamp_dummy_magic_19_0.VD3.n0 71.388
R6262 two_stage_opamp_dummy_magic_19_0.VD3.n14 two_stage_opamp_dummy_magic_19_0.VD3.n13 71.388
R6263 two_stage_opamp_dummy_magic_19_0.VD3.n21 two_stage_opamp_dummy_magic_19_0.VD3.n20 71.388
R6264 two_stage_opamp_dummy_magic_19_0.VD3.n23 two_stage_opamp_dummy_magic_19_0.VD3.n22 71.388
R6265 two_stage_opamp_dummy_magic_19_0.VD3.n12 two_stage_opamp_dummy_magic_19_0.VD3.n11 71.388
R6266 two_stage_opamp_dummy_magic_19_0.VD3.n10 two_stage_opamp_dummy_magic_19_0.VD3.n9 71.388
R6267 two_stage_opamp_dummy_magic_19_0.VD3.n8 two_stage_opamp_dummy_magic_19_0.VD3.n7 71.388
R6268 two_stage_opamp_dummy_magic_19_0.VD3.n6 two_stage_opamp_dummy_magic_19_0.VD3.n5 71.388
R6269 two_stage_opamp_dummy_magic_19_0.VD3.n4 two_stage_opamp_dummy_magic_19_0.VD3.n3 71.388
R6270 two_stage_opamp_dummy_magic_19_0.VD3.n25 two_stage_opamp_dummy_magic_19_0.VD3.n24 71.388
R6271 two_stage_opamp_dummy_magic_19_0.VD3.n19 two_stage_opamp_dummy_magic_19_0.VD3.n18 46.0195
R6272 two_stage_opamp_dummy_magic_19_0.VD3.n17 two_stage_opamp_dummy_magic_19_0.VD3.n16 46.0195
R6273 two_stage_opamp_dummy_magic_19_0.VD3.n21 two_stage_opamp_dummy_magic_19_0.VD3.n19 14.4255
R6274 two_stage_opamp_dummy_magic_19_0.VD3.n15 two_stage_opamp_dummy_magic_19_0.VD3.n12 14.1567
R6275 two_stage_opamp_dummy_magic_19_0.VD3.n16 two_stage_opamp_dummy_magic_19_0.VD3.n15 13.8005
R6276 two_stage_opamp_dummy_magic_19_0.VD3.n0 two_stage_opamp_dummy_magic_19_0.VD3.t9 11.2576
R6277 two_stage_opamp_dummy_magic_19_0.VD3.n0 two_stage_opamp_dummy_magic_19_0.VD3.t15 11.2576
R6278 two_stage_opamp_dummy_magic_19_0.VD3.n13 two_stage_opamp_dummy_magic_19_0.VD3.t5 11.2576
R6279 two_stage_opamp_dummy_magic_19_0.VD3.n13 two_stage_opamp_dummy_magic_19_0.VD3.t13 11.2576
R6280 two_stage_opamp_dummy_magic_19_0.VD3.n20 two_stage_opamp_dummy_magic_19_0.VD3.t11 11.2576
R6281 two_stage_opamp_dummy_magic_19_0.VD3.n20 two_stage_opamp_dummy_magic_19_0.VD3.t17 11.2576
R6282 two_stage_opamp_dummy_magic_19_0.VD3.n22 two_stage_opamp_dummy_magic_19_0.VD3.t7 11.2576
R6283 two_stage_opamp_dummy_magic_19_0.VD3.n22 two_stage_opamp_dummy_magic_19_0.VD3.t3 11.2576
R6284 two_stage_opamp_dummy_magic_19_0.VD3.n11 two_stage_opamp_dummy_magic_19_0.VD3.t26 11.2576
R6285 two_stage_opamp_dummy_magic_19_0.VD3.n11 two_stage_opamp_dummy_magic_19_0.VD3.t36 11.2576
R6286 two_stage_opamp_dummy_magic_19_0.VD3.n9 two_stage_opamp_dummy_magic_19_0.VD3.t33 11.2576
R6287 two_stage_opamp_dummy_magic_19_0.VD3.n9 two_stage_opamp_dummy_magic_19_0.VD3.t28 11.2576
R6288 two_stage_opamp_dummy_magic_19_0.VD3.n7 two_stage_opamp_dummy_magic_19_0.VD3.t31 11.2576
R6289 two_stage_opamp_dummy_magic_19_0.VD3.n7 two_stage_opamp_dummy_magic_19_0.VD3.t32 11.2576
R6290 two_stage_opamp_dummy_magic_19_0.VD3.n5 two_stage_opamp_dummy_magic_19_0.VD3.t30 11.2576
R6291 two_stage_opamp_dummy_magic_19_0.VD3.n5 two_stage_opamp_dummy_magic_19_0.VD3.t29 11.2576
R6292 two_stage_opamp_dummy_magic_19_0.VD3.n3 two_stage_opamp_dummy_magic_19_0.VD3.t35 11.2576
R6293 two_stage_opamp_dummy_magic_19_0.VD3.n3 two_stage_opamp_dummy_magic_19_0.VD3.t27 11.2576
R6294 two_stage_opamp_dummy_magic_19_0.VD3.n2 two_stage_opamp_dummy_magic_19_0.VD3.t37 11.2576
R6295 two_stage_opamp_dummy_magic_19_0.VD3.n2 two_stage_opamp_dummy_magic_19_0.VD3.t34 11.2576
R6296 two_stage_opamp_dummy_magic_19_0.VD3.t19 two_stage_opamp_dummy_magic_19_0.VD3.n25 11.2576
R6297 two_stage_opamp_dummy_magic_19_0.VD3.n25 two_stage_opamp_dummy_magic_19_0.VD3.t1 11.2576
R6298 two_stage_opamp_dummy_magic_19_0.VD3.n24 two_stage_opamp_dummy_magic_19_0.VD3.n23 0.6255
R6299 two_stage_opamp_dummy_magic_19_0.VD3.n23 two_stage_opamp_dummy_magic_19_0.VD3.n21 0.6255
R6300 two_stage_opamp_dummy_magic_19_0.VD3.n6 two_stage_opamp_dummy_magic_19_0.VD3.n4 0.6255
R6301 two_stage_opamp_dummy_magic_19_0.VD3.n8 two_stage_opamp_dummy_magic_19_0.VD3.n6 0.6255
R6302 two_stage_opamp_dummy_magic_19_0.VD3.n10 two_stage_opamp_dummy_magic_19_0.VD3.n8 0.6255
R6303 two_stage_opamp_dummy_magic_19_0.VD3.n12 two_stage_opamp_dummy_magic_19_0.VD3.n10 0.6255
R6304 two_stage_opamp_dummy_magic_19_0.VD3.n15 two_stage_opamp_dummy_magic_19_0.VD3.n14 0.6255
R6305 two_stage_opamp_dummy_magic_19_0.VD3.n14 two_stage_opamp_dummy_magic_19_0.VD3.n1 0.6255
R6306 two_stage_opamp_dummy_magic_19_0.VD3.n24 two_stage_opamp_dummy_magic_19_0.VD3.n1 0.6255
R6307 two_stage_opamp_dummy_magic_19_0.Y.n57 two_stage_opamp_dummy_magic_19_0.Y.t36 1172.87
R6308 two_stage_opamp_dummy_magic_19_0.Y.n53 two_stage_opamp_dummy_magic_19_0.Y.t30 1172.87
R6309 two_stage_opamp_dummy_magic_19_0.Y.n57 two_stage_opamp_dummy_magic_19_0.Y.t52 996.134
R6310 two_stage_opamp_dummy_magic_19_0.Y.n58 two_stage_opamp_dummy_magic_19_0.Y.t46 996.134
R6311 two_stage_opamp_dummy_magic_19_0.Y.n59 two_stage_opamp_dummy_magic_19_0.Y.t51 996.134
R6312 two_stage_opamp_dummy_magic_19_0.Y.n60 two_stage_opamp_dummy_magic_19_0.Y.t37 996.134
R6313 two_stage_opamp_dummy_magic_19_0.Y.n56 two_stage_opamp_dummy_magic_19_0.Y.t54 996.134
R6314 two_stage_opamp_dummy_magic_19_0.Y.n55 two_stage_opamp_dummy_magic_19_0.Y.t40 996.134
R6315 two_stage_opamp_dummy_magic_19_0.Y.n54 two_stage_opamp_dummy_magic_19_0.Y.t26 996.134
R6316 two_stage_opamp_dummy_magic_19_0.Y.n53 two_stage_opamp_dummy_magic_19_0.Y.t43 996.134
R6317 two_stage_opamp_dummy_magic_19_0.Y.n47 two_stage_opamp_dummy_magic_19_0.Y.t41 690.867
R6318 two_stage_opamp_dummy_magic_19_0.Y.n42 two_stage_opamp_dummy_magic_19_0.Y.t35 690.867
R6319 two_stage_opamp_dummy_magic_19_0.Y.n38 two_stage_opamp_dummy_magic_19_0.Y.t53 530.201
R6320 two_stage_opamp_dummy_magic_19_0.Y.n33 two_stage_opamp_dummy_magic_19_0.Y.t48 530.201
R6321 two_stage_opamp_dummy_magic_19_0.Y.n49 two_stage_opamp_dummy_magic_19_0.Y.t27 514.134
R6322 two_stage_opamp_dummy_magic_19_0.Y.n48 two_stage_opamp_dummy_magic_19_0.Y.t50 514.134
R6323 two_stage_opamp_dummy_magic_19_0.Y.n47 two_stage_opamp_dummy_magic_19_0.Y.t28 514.134
R6324 two_stage_opamp_dummy_magic_19_0.Y.n42 two_stage_opamp_dummy_magic_19_0.Y.t49 514.134
R6325 two_stage_opamp_dummy_magic_19_0.Y.n43 two_stage_opamp_dummy_magic_19_0.Y.t33 514.134
R6326 two_stage_opamp_dummy_magic_19_0.Y.n44 two_stage_opamp_dummy_magic_19_0.Y.t47 514.134
R6327 two_stage_opamp_dummy_magic_19_0.Y.n45 two_stage_opamp_dummy_magic_19_0.Y.t31 514.134
R6328 two_stage_opamp_dummy_magic_19_0.Y.n46 two_stage_opamp_dummy_magic_19_0.Y.t44 514.134
R6329 two_stage_opamp_dummy_magic_19_0.Y.n62 two_stage_opamp_dummy_magic_19_0.Y.n61 424.875
R6330 two_stage_opamp_dummy_magic_19_0.Y.n38 two_stage_opamp_dummy_magic_19_0.Y.t39 353.467
R6331 two_stage_opamp_dummy_magic_19_0.Y.n39 two_stage_opamp_dummy_magic_19_0.Y.t34 353.467
R6332 two_stage_opamp_dummy_magic_19_0.Y.n40 two_stage_opamp_dummy_magic_19_0.Y.t38 353.467
R6333 two_stage_opamp_dummy_magic_19_0.Y.n37 two_stage_opamp_dummy_magic_19_0.Y.t25 353.467
R6334 two_stage_opamp_dummy_magic_19_0.Y.n36 two_stage_opamp_dummy_magic_19_0.Y.t42 353.467
R6335 two_stage_opamp_dummy_magic_19_0.Y.n35 two_stage_opamp_dummy_magic_19_0.Y.t29 353.467
R6336 two_stage_opamp_dummy_magic_19_0.Y.n34 two_stage_opamp_dummy_magic_19_0.Y.t45 353.467
R6337 two_stage_opamp_dummy_magic_19_0.Y.n33 two_stage_opamp_dummy_magic_19_0.Y.t32 353.467
R6338 two_stage_opamp_dummy_magic_19_0.Y.n56 two_stage_opamp_dummy_magic_19_0.Y.n55 176.733
R6339 two_stage_opamp_dummy_magic_19_0.Y.n55 two_stage_opamp_dummy_magic_19_0.Y.n54 176.733
R6340 two_stage_opamp_dummy_magic_19_0.Y.n54 two_stage_opamp_dummy_magic_19_0.Y.n53 176.733
R6341 two_stage_opamp_dummy_magic_19_0.Y.n58 two_stage_opamp_dummy_magic_19_0.Y.n57 176.733
R6342 two_stage_opamp_dummy_magic_19_0.Y.n59 two_stage_opamp_dummy_magic_19_0.Y.n58 176.733
R6343 two_stage_opamp_dummy_magic_19_0.Y.n60 two_stage_opamp_dummy_magic_19_0.Y.n59 176.733
R6344 two_stage_opamp_dummy_magic_19_0.Y.n37 two_stage_opamp_dummy_magic_19_0.Y.n36 176.733
R6345 two_stage_opamp_dummy_magic_19_0.Y.n36 two_stage_opamp_dummy_magic_19_0.Y.n35 176.733
R6346 two_stage_opamp_dummy_magic_19_0.Y.n35 two_stage_opamp_dummy_magic_19_0.Y.n34 176.733
R6347 two_stage_opamp_dummy_magic_19_0.Y.n34 two_stage_opamp_dummy_magic_19_0.Y.n33 176.733
R6348 two_stage_opamp_dummy_magic_19_0.Y.n39 two_stage_opamp_dummy_magic_19_0.Y.n38 176.733
R6349 two_stage_opamp_dummy_magic_19_0.Y.n40 two_stage_opamp_dummy_magic_19_0.Y.n39 176.733
R6350 two_stage_opamp_dummy_magic_19_0.Y.n46 two_stage_opamp_dummy_magic_19_0.Y.n45 176.733
R6351 two_stage_opamp_dummy_magic_19_0.Y.n45 two_stage_opamp_dummy_magic_19_0.Y.n44 176.733
R6352 two_stage_opamp_dummy_magic_19_0.Y.n44 two_stage_opamp_dummy_magic_19_0.Y.n43 176.733
R6353 two_stage_opamp_dummy_magic_19_0.Y.n43 two_stage_opamp_dummy_magic_19_0.Y.n42 176.733
R6354 two_stage_opamp_dummy_magic_19_0.Y.n48 two_stage_opamp_dummy_magic_19_0.Y.n47 176.733
R6355 two_stage_opamp_dummy_magic_19_0.Y.n49 two_stage_opamp_dummy_magic_19_0.Y.n48 176.733
R6356 two_stage_opamp_dummy_magic_19_0.Y.n52 two_stage_opamp_dummy_magic_19_0.Y.n51 174.769
R6357 two_stage_opamp_dummy_magic_19_0.Y.n51 two_stage_opamp_dummy_magic_19_0.Y.n41 162.675
R6358 two_stage_opamp_dummy_magic_19_0.Y.n51 two_stage_opamp_dummy_magic_19_0.Y.n50 162.675
R6359 two_stage_opamp_dummy_magic_19_0.Y.n8 two_stage_opamp_dummy_magic_19_0.Y.n6 72.013
R6360 two_stage_opamp_dummy_magic_19_0.Y.n3 two_stage_opamp_dummy_magic_19_0.Y.n1 72.013
R6361 two_stage_opamp_dummy_magic_19_0.Y.n8 two_stage_opamp_dummy_magic_19_0.Y.n7 71.388
R6362 two_stage_opamp_dummy_magic_19_0.Y.n5 two_stage_opamp_dummy_magic_19_0.Y.n4 71.388
R6363 two_stage_opamp_dummy_magic_19_0.Y.n3 two_stage_opamp_dummy_magic_19_0.Y.n2 71.388
R6364 two_stage_opamp_dummy_magic_19_0.Y.n10 two_stage_opamp_dummy_magic_19_0.Y.n0 66.888
R6365 two_stage_opamp_dummy_magic_19_0.Y.n61 two_stage_opamp_dummy_magic_19_0.Y.n56 56.2338
R6366 two_stage_opamp_dummy_magic_19_0.Y.n61 two_stage_opamp_dummy_magic_19_0.Y.n60 56.2338
R6367 two_stage_opamp_dummy_magic_19_0.Y.n41 two_stage_opamp_dummy_magic_19_0.Y.n37 56.2338
R6368 two_stage_opamp_dummy_magic_19_0.Y.n41 two_stage_opamp_dummy_magic_19_0.Y.n40 56.2338
R6369 two_stage_opamp_dummy_magic_19_0.Y.n50 two_stage_opamp_dummy_magic_19_0.Y.n46 56.2338
R6370 two_stage_opamp_dummy_magic_19_0.Y.n50 two_stage_opamp_dummy_magic_19_0.Y.n49 56.2338
R6371 two_stage_opamp_dummy_magic_19_0.Y.t11 two_stage_opamp_dummy_magic_19_0.Y.n62 49.8031
R6372 two_stage_opamp_dummy_magic_19_0.Y.n14 two_stage_opamp_dummy_magic_19_0.Y.n13 49.3505
R6373 two_stage_opamp_dummy_magic_19_0.Y.n17 two_stage_opamp_dummy_magic_19_0.Y.n16 49.3505
R6374 two_stage_opamp_dummy_magic_19_0.Y.n20 two_stage_opamp_dummy_magic_19_0.Y.n19 49.3505
R6375 two_stage_opamp_dummy_magic_19_0.Y.n24 two_stage_opamp_dummy_magic_19_0.Y.n23 49.3505
R6376 two_stage_opamp_dummy_magic_19_0.Y.n27 two_stage_opamp_dummy_magic_19_0.Y.n26 49.3505
R6377 two_stage_opamp_dummy_magic_19_0.Y.n30 two_stage_opamp_dummy_magic_19_0.Y.n29 49.3505
R6378 two_stage_opamp_dummy_magic_19_0.Y.n32 two_stage_opamp_dummy_magic_19_0.Y.n10 17.688
R6379 two_stage_opamp_dummy_magic_19_0.Y.n13 two_stage_opamp_dummy_magic_19_0.Y.t22 16.0005
R6380 two_stage_opamp_dummy_magic_19_0.Y.n13 two_stage_opamp_dummy_magic_19_0.Y.t19 16.0005
R6381 two_stage_opamp_dummy_magic_19_0.Y.n16 two_stage_opamp_dummy_magic_19_0.Y.t23 16.0005
R6382 two_stage_opamp_dummy_magic_19_0.Y.n16 two_stage_opamp_dummy_magic_19_0.Y.t17 16.0005
R6383 two_stage_opamp_dummy_magic_19_0.Y.n19 two_stage_opamp_dummy_magic_19_0.Y.t16 16.0005
R6384 two_stage_opamp_dummy_magic_19_0.Y.n19 two_stage_opamp_dummy_magic_19_0.Y.t20 16.0005
R6385 two_stage_opamp_dummy_magic_19_0.Y.n23 two_stage_opamp_dummy_magic_19_0.Y.t18 16.0005
R6386 two_stage_opamp_dummy_magic_19_0.Y.n23 two_stage_opamp_dummy_magic_19_0.Y.t24 16.0005
R6387 two_stage_opamp_dummy_magic_19_0.Y.n26 two_stage_opamp_dummy_magic_19_0.Y.t13 16.0005
R6388 two_stage_opamp_dummy_magic_19_0.Y.n26 two_stage_opamp_dummy_magic_19_0.Y.t14 16.0005
R6389 two_stage_opamp_dummy_magic_19_0.Y.n29 two_stage_opamp_dummy_magic_19_0.Y.t0 16.0005
R6390 two_stage_opamp_dummy_magic_19_0.Y.n29 two_stage_opamp_dummy_magic_19_0.Y.t21 16.0005
R6391 two_stage_opamp_dummy_magic_19_0.Y.n7 two_stage_opamp_dummy_magic_19_0.Y.t9 11.2576
R6392 two_stage_opamp_dummy_magic_19_0.Y.n7 two_stage_opamp_dummy_magic_19_0.Y.t4 11.2576
R6393 two_stage_opamp_dummy_magic_19_0.Y.n6 two_stage_opamp_dummy_magic_19_0.Y.t2 11.2576
R6394 two_stage_opamp_dummy_magic_19_0.Y.n6 two_stage_opamp_dummy_magic_19_0.Y.t12 11.2576
R6395 two_stage_opamp_dummy_magic_19_0.Y.n4 two_stage_opamp_dummy_magic_19_0.Y.t7 11.2576
R6396 two_stage_opamp_dummy_magic_19_0.Y.n4 two_stage_opamp_dummy_magic_19_0.Y.t6 11.2576
R6397 two_stage_opamp_dummy_magic_19_0.Y.n2 two_stage_opamp_dummy_magic_19_0.Y.t8 11.2576
R6398 two_stage_opamp_dummy_magic_19_0.Y.n2 two_stage_opamp_dummy_magic_19_0.Y.t1 11.2576
R6399 two_stage_opamp_dummy_magic_19_0.Y.n1 two_stage_opamp_dummy_magic_19_0.Y.t15 11.2576
R6400 two_stage_opamp_dummy_magic_19_0.Y.n1 two_stage_opamp_dummy_magic_19_0.Y.t10 11.2576
R6401 two_stage_opamp_dummy_magic_19_0.Y.n0 two_stage_opamp_dummy_magic_19_0.Y.t5 11.2576
R6402 two_stage_opamp_dummy_magic_19_0.Y.n0 two_stage_opamp_dummy_magic_19_0.Y.t3 11.2576
R6403 two_stage_opamp_dummy_magic_19_0.Y.n62 two_stage_opamp_dummy_magic_19_0.Y.n52 7.09425
R6404 two_stage_opamp_dummy_magic_19_0.Y.n32 two_stage_opamp_dummy_magic_19_0.Y.n31 6.3755
R6405 two_stage_opamp_dummy_magic_19_0.Y.n15 two_stage_opamp_dummy_magic_19_0.Y.n14 5.71404
R6406 two_stage_opamp_dummy_magic_19_0.Y.n30 two_stage_opamp_dummy_magic_19_0.Y.n28 5.71404
R6407 two_stage_opamp_dummy_magic_19_0.Y.n18 two_stage_opamp_dummy_magic_19_0.Y.n14 5.5005
R6408 two_stage_opamp_dummy_magic_19_0.Y.n17 two_stage_opamp_dummy_magic_19_0.Y.n15 5.10988
R6409 two_stage_opamp_dummy_magic_19_0.Y.n20 two_stage_opamp_dummy_magic_19_0.Y.n12 5.10988
R6410 two_stage_opamp_dummy_magic_19_0.Y.n25 two_stage_opamp_dummy_magic_19_0.Y.n24 5.10988
R6411 two_stage_opamp_dummy_magic_19_0.Y.n28 two_stage_opamp_dummy_magic_19_0.Y.n27 5.10988
R6412 two_stage_opamp_dummy_magic_19_0.Y.n18 two_stage_opamp_dummy_magic_19_0.Y.n17 4.938
R6413 two_stage_opamp_dummy_magic_19_0.Y.n21 two_stage_opamp_dummy_magic_19_0.Y.n20 4.938
R6414 two_stage_opamp_dummy_magic_19_0.Y.n24 two_stage_opamp_dummy_magic_19_0.Y.n22 4.938
R6415 two_stage_opamp_dummy_magic_19_0.Y.n27 two_stage_opamp_dummy_magic_19_0.Y.n11 4.938
R6416 two_stage_opamp_dummy_magic_19_0.Y.n31 two_stage_opamp_dummy_magic_19_0.Y.n30 4.938
R6417 two_stage_opamp_dummy_magic_19_0.Y.n10 two_stage_opamp_dummy_magic_19_0.Y.n9 4.5005
R6418 two_stage_opamp_dummy_magic_19_0.Y.n52 two_stage_opamp_dummy_magic_19_0.Y.n32 1.03175
R6419 two_stage_opamp_dummy_magic_19_0.Y.n9 two_stage_opamp_dummy_magic_19_0.Y.n8 0.6255
R6420 two_stage_opamp_dummy_magic_19_0.Y.n5 two_stage_opamp_dummy_magic_19_0.Y.n3 0.6255
R6421 two_stage_opamp_dummy_magic_19_0.Y.n9 two_stage_opamp_dummy_magic_19_0.Y.n5 0.6255
R6422 two_stage_opamp_dummy_magic_19_0.Y.n28 two_stage_opamp_dummy_magic_19_0.Y.n25 0.604667
R6423 two_stage_opamp_dummy_magic_19_0.Y.n25 two_stage_opamp_dummy_magic_19_0.Y.n12 0.604667
R6424 two_stage_opamp_dummy_magic_19_0.Y.n15 two_stage_opamp_dummy_magic_19_0.Y.n12 0.604667
R6425 two_stage_opamp_dummy_magic_19_0.Y.n21 two_stage_opamp_dummy_magic_19_0.Y.n18 0.563
R6426 two_stage_opamp_dummy_magic_19_0.Y.n22 two_stage_opamp_dummy_magic_19_0.Y.n21 0.563
R6427 two_stage_opamp_dummy_magic_19_0.Y.n22 two_stage_opamp_dummy_magic_19_0.Y.n11 0.563
R6428 two_stage_opamp_dummy_magic_19_0.Y.n31 two_stage_opamp_dummy_magic_19_0.Y.n11 0.563
R6429 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n0 345.264
R6430 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n1 344.7
R6431 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n3 292.5
R6432 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n5 124.403
R6433 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n12 123.84
R6434 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n10 123.84
R6435 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n8 123.84
R6436 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n6 123.84
R6437 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t1 120.43
R6438 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n2 52.763
R6439 bgr_9_0.V_CMFB_S3 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n4 51.7297
R6440 bgr_9_0.V_CMFB_S3 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n14 41.1227
R6441 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t14 39.4005
R6442 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t2 39.4005
R6443 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t16 39.4005
R6444 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t13 39.4005
R6445 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t0 39.4005
R6446 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t15 39.4005
R6447 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t10 19.7005
R6448 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t4 19.7005
R6449 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t11 19.7005
R6450 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t5 19.7005
R6451 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t12 19.7005
R6452 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t6 19.7005
R6453 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t9 19.7005
R6454 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t8 19.7005
R6455 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t3 19.7005
R6456 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t7 19.7005
R6457 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n13 5.90675
R6458 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n7 0.563
R6459 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n9 0.563
R6460 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n11 0.563
R6461 bgr_9_0.V_CUR_REF_REG.n4 bgr_9_0.V_CUR_REF_REG.n3 526.183
R6462 bgr_9_0.V_CUR_REF_REG.n2 bgr_9_0.V_CUR_REF_REG.n1 514.134
R6463 bgr_9_0.V_CUR_REF_REG.n5 bgr_9_0.V_CUR_REF_REG.n0 378.053
R6464 bgr_9_0.V_CUR_REF_REG.n1 bgr_9_0.V_CUR_REF_REG.t5 303.259
R6465 bgr_9_0.V_CUR_REF_REG.n5 bgr_9_0.V_CUR_REF_REG.n4 210.169
R6466 bgr_9_0.V_CUR_REF_REG.n1 bgr_9_0.V_CUR_REF_REG.t3 174.726
R6467 bgr_9_0.V_CUR_REF_REG.n2 bgr_9_0.V_CUR_REF_REG.t7 174.726
R6468 bgr_9_0.V_CUR_REF_REG.n3 bgr_9_0.V_CUR_REF_REG.t4 174.726
R6469 bgr_9_0.V_CUR_REF_REG.t0 bgr_9_0.V_CUR_REF_REG.n5 153.474
R6470 bgr_9_0.V_CUR_REF_REG.n3 bgr_9_0.V_CUR_REF_REG.n2 128.534
R6471 bgr_9_0.V_CUR_REF_REG.n4 bgr_9_0.V_CUR_REF_REG.t6 96.4005
R6472 bgr_9_0.V_CUR_REF_REG.n0 bgr_9_0.V_CUR_REF_REG.t1 39.4005
R6473 bgr_9_0.V_CUR_REF_REG.n0 bgr_9_0.V_CUR_REF_REG.t2 39.4005
R6474 bgr_9_0.V_p_2.n6 bgr_9_0.V_p_2.n5 263.933
R6475 bgr_9_0.V_p_2.n2 bgr_9_0.V_p_2.n0 263.933
R6476 bgr_9_0.V_p_2.n2 bgr_9_0.V_p_2.n1 206.333
R6477 bgr_9_0.V_p_2.n4 bgr_9_0.V_p_2.n3 206.333
R6478 bgr_9_0.V_p_2.n7 bgr_9_0.V_p_2.n6 206.333
R6479 bgr_9_0.V_p_2.n4 bgr_9_0.V_p_2.t10 134.474
R6480 bgr_9_0.V_p_2.n4 bgr_9_0.V_p_2.n2 57.6005
R6481 bgr_9_0.V_p_2.n6 bgr_9_0.V_p_2.n4 57.6005
R6482 bgr_9_0.V_p_2.n5 bgr_9_0.V_p_2.t0 48.0005
R6483 bgr_9_0.V_p_2.n5 bgr_9_0.V_p_2.t7 48.0005
R6484 bgr_9_0.V_p_2.n0 bgr_9_0.V_p_2.t1 48.0005
R6485 bgr_9_0.V_p_2.n0 bgr_9_0.V_p_2.t6 48.0005
R6486 bgr_9_0.V_p_2.n1 bgr_9_0.V_p_2.t8 48.0005
R6487 bgr_9_0.V_p_2.n1 bgr_9_0.V_p_2.t3 48.0005
R6488 bgr_9_0.V_p_2.n3 bgr_9_0.V_p_2.t2 48.0005
R6489 bgr_9_0.V_p_2.n3 bgr_9_0.V_p_2.t5 48.0005
R6490 bgr_9_0.V_p_2.t9 bgr_9_0.V_p_2.n7 48.0005
R6491 bgr_9_0.V_p_2.n7 bgr_9_0.V_p_2.t4 48.0005
R6492 a_7460_23988.t0 a_7460_23988.t1 178.133
R6493 two_stage_opamp_dummy_magic_19_0.VD2.n8 two_stage_opamp_dummy_magic_19_0.VD2.n6 54.8765
R6494 two_stage_opamp_dummy_magic_19_0.VD2.n5 two_stage_opamp_dummy_magic_19_0.VD2.n3 54.839
R6495 two_stage_opamp_dummy_magic_19_0.VD2.n12 two_stage_opamp_dummy_magic_19_0.VD2.n10 54.788
R6496 two_stage_opamp_dummy_magic_19_0.VD2.n16 two_stage_opamp_dummy_magic_19_0.VD2.n14 54.788
R6497 two_stage_opamp_dummy_magic_19_0.VD2.n8 two_stage_opamp_dummy_magic_19_0.VD2.n7 54.2724
R6498 two_stage_opamp_dummy_magic_19_0.VD2.n5 two_stage_opamp_dummy_magic_19_0.VD2.n4 54.2724
R6499 two_stage_opamp_dummy_magic_19_0.VD2.n16 two_stage_opamp_dummy_magic_19_0.VD2.n15 54.2255
R6500 two_stage_opamp_dummy_magic_19_0.VD2.n1 two_stage_opamp_dummy_magic_19_0.VD2.n17 54.2255
R6501 two_stage_opamp_dummy_magic_19_0.VD2.n0 two_stage_opamp_dummy_magic_19_0.VD2.n13 54.2255
R6502 two_stage_opamp_dummy_magic_19_0.VD2.n12 two_stage_opamp_dummy_magic_19_0.VD2.n11 54.2255
R6503 two_stage_opamp_dummy_magic_19_0.VD2 two_stage_opamp_dummy_magic_19_0.VD2.n2 49.7724
R6504 two_stage_opamp_dummy_magic_19_0.VD2.n15 two_stage_opamp_dummy_magic_19_0.VD2.t14 16.0005
R6505 two_stage_opamp_dummy_magic_19_0.VD2.n15 two_stage_opamp_dummy_magic_19_0.VD2.t15 16.0005
R6506 two_stage_opamp_dummy_magic_19_0.VD2.n17 two_stage_opamp_dummy_magic_19_0.VD2.t8 16.0005
R6507 two_stage_opamp_dummy_magic_19_0.VD2.n17 two_stage_opamp_dummy_magic_19_0.VD2.t3 16.0005
R6508 two_stage_opamp_dummy_magic_19_0.VD2.n7 two_stage_opamp_dummy_magic_19_0.VD2.t21 16.0005
R6509 two_stage_opamp_dummy_magic_19_0.VD2.n7 two_stage_opamp_dummy_magic_19_0.VD2.t4 16.0005
R6510 two_stage_opamp_dummy_magic_19_0.VD2.n6 two_stage_opamp_dummy_magic_19_0.VD2.t5 16.0005
R6511 two_stage_opamp_dummy_magic_19_0.VD2.n6 two_stage_opamp_dummy_magic_19_0.VD2.t1 16.0005
R6512 two_stage_opamp_dummy_magic_19_0.VD2.n4 two_stage_opamp_dummy_magic_19_0.VD2.t11 16.0005
R6513 two_stage_opamp_dummy_magic_19_0.VD2.n4 two_stage_opamp_dummy_magic_19_0.VD2.t10 16.0005
R6514 two_stage_opamp_dummy_magic_19_0.VD2.n3 two_stage_opamp_dummy_magic_19_0.VD2.t13 16.0005
R6515 two_stage_opamp_dummy_magic_19_0.VD2.n3 two_stage_opamp_dummy_magic_19_0.VD2.t19 16.0005
R6516 two_stage_opamp_dummy_magic_19_0.VD2.n2 two_stage_opamp_dummy_magic_19_0.VD2.t16 16.0005
R6517 two_stage_opamp_dummy_magic_19_0.VD2.n2 two_stage_opamp_dummy_magic_19_0.VD2.t12 16.0005
R6518 two_stage_opamp_dummy_magic_19_0.VD2.n13 two_stage_opamp_dummy_magic_19_0.VD2.t7 16.0005
R6519 two_stage_opamp_dummy_magic_19_0.VD2.n13 two_stage_opamp_dummy_magic_19_0.VD2.t0 16.0005
R6520 two_stage_opamp_dummy_magic_19_0.VD2.n11 two_stage_opamp_dummy_magic_19_0.VD2.t20 16.0005
R6521 two_stage_opamp_dummy_magic_19_0.VD2.n11 two_stage_opamp_dummy_magic_19_0.VD2.t9 16.0005
R6522 two_stage_opamp_dummy_magic_19_0.VD2.n10 two_stage_opamp_dummy_magic_19_0.VD2.t17 16.0005
R6523 two_stage_opamp_dummy_magic_19_0.VD2.n10 two_stage_opamp_dummy_magic_19_0.VD2.t6 16.0005
R6524 two_stage_opamp_dummy_magic_19_0.VD2.n14 two_stage_opamp_dummy_magic_19_0.VD2.t2 16.0005
R6525 two_stage_opamp_dummy_magic_19_0.VD2.n14 two_stage_opamp_dummy_magic_19_0.VD2.t18 16.0005
R6526 two_stage_opamp_dummy_magic_19_0.VD2 two_stage_opamp_dummy_magic_19_0.VD2.n9 4.94321
R6527 two_stage_opamp_dummy_magic_19_0.VD2 two_stage_opamp_dummy_magic_19_0.VD2.n1 4.813
R6528 two_stage_opamp_dummy_magic_19_0.VD2.n9 two_stage_opamp_dummy_magic_19_0.VD2.n8 0.604667
R6529 two_stage_opamp_dummy_magic_19_0.VD2.n9 two_stage_opamp_dummy_magic_19_0.VD2.n5 0.604667
R6530 two_stage_opamp_dummy_magic_19_0.VD2.n0 two_stage_opamp_dummy_magic_19_0.VD2.n12 0.563
R6531 two_stage_opamp_dummy_magic_19_0.VD2.n1 two_stage_opamp_dummy_magic_19_0.VD2.n16 0.563
R6532 two_stage_opamp_dummy_magic_19_0.VD2.n1 two_stage_opamp_dummy_magic_19_0.VD2.n0 0.46925
R6533 two_stage_opamp_dummy_magic_19_0.V_err_gate.n2 two_stage_opamp_dummy_magic_19_0.V_err_gate.t6 479.322
R6534 two_stage_opamp_dummy_magic_19_0.V_err_gate.n2 two_stage_opamp_dummy_magic_19_0.V_err_gate.t8 479.322
R6535 two_stage_opamp_dummy_magic_19_0.V_err_gate.n6 two_stage_opamp_dummy_magic_19_0.V_err_gate.t9 479.322
R6536 two_stage_opamp_dummy_magic_19_0.V_err_gate.n6 two_stage_opamp_dummy_magic_19_0.V_err_gate.t7 479.322
R6537 two_stage_opamp_dummy_magic_19_0.V_err_gate two_stage_opamp_dummy_magic_19_0.V_err_gate.n0 180.637
R6538 two_stage_opamp_dummy_magic_19_0.V_err_gate.n3 two_stage_opamp_dummy_magic_19_0.V_err_gate.n2 165.8
R6539 two_stage_opamp_dummy_magic_19_0.V_err_gate two_stage_opamp_dummy_magic_19_0.V_err_gate.n6 165.8
R6540 two_stage_opamp_dummy_magic_19_0.V_err_gate.n3 two_stage_opamp_dummy_magic_19_0.V_err_gate.n1 104.957
R6541 two_stage_opamp_dummy_magic_19_0.V_err_gate.n5 two_stage_opamp_dummy_magic_19_0.V_err_gate.n4 104.3
R6542 two_stage_opamp_dummy_magic_19_0.V_err_gate.n0 two_stage_opamp_dummy_magic_19_0.V_err_gate.t2 24.0005
R6543 two_stage_opamp_dummy_magic_19_0.V_err_gate.n0 two_stage_opamp_dummy_magic_19_0.V_err_gate.t3 24.0005
R6544 two_stage_opamp_dummy_magic_19_0.V_err_gate.n4 two_stage_opamp_dummy_magic_19_0.V_err_gate.t4 15.7605
R6545 two_stage_opamp_dummy_magic_19_0.V_err_gate.n4 two_stage_opamp_dummy_magic_19_0.V_err_gate.t0 15.7605
R6546 two_stage_opamp_dummy_magic_19_0.V_err_gate.n1 two_stage_opamp_dummy_magic_19_0.V_err_gate.t1 15.7605
R6547 two_stage_opamp_dummy_magic_19_0.V_err_gate.n1 two_stage_opamp_dummy_magic_19_0.V_err_gate.t5 15.7605
R6548 two_stage_opamp_dummy_magic_19_0.V_err_gate two_stage_opamp_dummy_magic_19_0.V_err_gate.n5 1.71925
R6549 two_stage_opamp_dummy_magic_19_0.V_err_gate.n5 two_stage_opamp_dummy_magic_19_0.V_err_gate.n3 0.65675
R6550 two_stage_opamp_dummy_magic_19_0.V_err_mir_p two_stage_opamp_dummy_magic_19_0.V_err_mir_p.n0 109.197
R6551 two_stage_opamp_dummy_magic_19_0.V_err_mir_p two_stage_opamp_dummy_magic_19_0.V_err_mir_p.n1 99.5713
R6552 two_stage_opamp_dummy_magic_19_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_19_0.V_err_mir_p.t0 15.7605
R6553 two_stage_opamp_dummy_magic_19_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_19_0.V_err_mir_p.t1 15.7605
R6554 two_stage_opamp_dummy_magic_19_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_19_0.V_err_mir_p.t2 15.7605
R6555 two_stage_opamp_dummy_magic_19_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_19_0.V_err_mir_p.t3 15.7605
R6556 two_stage_opamp_dummy_magic_19_0.Vb1.n16 two_stage_opamp_dummy_magic_19_0.Vb1.t20 449.868
R6557 two_stage_opamp_dummy_magic_19_0.Vb1.n10 two_stage_opamp_dummy_magic_19_0.Vb1.t26 449.868
R6558 two_stage_opamp_dummy_magic_19_0.Vb1.n3 two_stage_opamp_dummy_magic_19_0.Vb1.t12 449.868
R6559 two_stage_opamp_dummy_magic_19_0.Vb1.n1 two_stage_opamp_dummy_magic_19_0.Vb1.t18 449.868
R6560 two_stage_opamp_dummy_magic_19_0.Vb1.n23 two_stage_opamp_dummy_magic_19_0.Vb1.t5 449.868
R6561 two_stage_opamp_dummy_magic_19_0.Vb1.n22 two_stage_opamp_dummy_magic_19_0.Vb1.t3 449.868
R6562 two_stage_opamp_dummy_magic_19_0.Vb1.n19 two_stage_opamp_dummy_magic_19_0.Vb1.n9 335.248
R6563 two_stage_opamp_dummy_magic_19_0.Vb1.n19 two_stage_opamp_dummy_magic_19_0.Vb1.n18 326.467
R6564 two_stage_opamp_dummy_magic_19_0.Vb1.n16 two_stage_opamp_dummy_magic_19_0.Vb1.t29 273.134
R6565 two_stage_opamp_dummy_magic_19_0.Vb1.n17 two_stage_opamp_dummy_magic_19_0.Vb1.t14 273.134
R6566 two_stage_opamp_dummy_magic_19_0.Vb1.n15 two_stage_opamp_dummy_magic_19_0.Vb1.t25 273.134
R6567 two_stage_opamp_dummy_magic_19_0.Vb1.n14 two_stage_opamp_dummy_magic_19_0.Vb1.t32 273.134
R6568 two_stage_opamp_dummy_magic_19_0.Vb1.n13 two_stage_opamp_dummy_magic_19_0.Vb1.t22 273.134
R6569 two_stage_opamp_dummy_magic_19_0.Vb1.n12 two_stage_opamp_dummy_magic_19_0.Vb1.t17 273.134
R6570 two_stage_opamp_dummy_magic_19_0.Vb1.n11 two_stage_opamp_dummy_magic_19_0.Vb1.t27 273.134
R6571 two_stage_opamp_dummy_magic_19_0.Vb1.n10 two_stage_opamp_dummy_magic_19_0.Vb1.t16 273.134
R6572 two_stage_opamp_dummy_magic_19_0.Vb1.n3 two_stage_opamp_dummy_magic_19_0.Vb1.t23 273.134
R6573 two_stage_opamp_dummy_magic_19_0.Vb1.n4 two_stage_opamp_dummy_magic_19_0.Vb1.t13 273.134
R6574 two_stage_opamp_dummy_magic_19_0.Vb1.n5 two_stage_opamp_dummy_magic_19_0.Vb1.t24 273.134
R6575 two_stage_opamp_dummy_magic_19_0.Vb1.n6 two_stage_opamp_dummy_magic_19_0.Vb1.t31 273.134
R6576 two_stage_opamp_dummy_magic_19_0.Vb1.n7 two_stage_opamp_dummy_magic_19_0.Vb1.t21 273.134
R6577 two_stage_opamp_dummy_magic_19_0.Vb1.n8 two_stage_opamp_dummy_magic_19_0.Vb1.t30 273.134
R6578 two_stage_opamp_dummy_magic_19_0.Vb1.n2 two_stage_opamp_dummy_magic_19_0.Vb1.t19 273.134
R6579 two_stage_opamp_dummy_magic_19_0.Vb1.n1 two_stage_opamp_dummy_magic_19_0.Vb1.t28 273.134
R6580 two_stage_opamp_dummy_magic_19_0.Vb1.n23 two_stage_opamp_dummy_magic_19_0.Vb1.t1 273.134
R6581 two_stage_opamp_dummy_magic_19_0.Vb1.n22 two_stage_opamp_dummy_magic_19_0.Vb1.t7 273.134
R6582 bgr_9_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_19_0.Vb1.n0 202.94
R6583 two_stage_opamp_dummy_magic_19_0.Vb1.n11 two_stage_opamp_dummy_magic_19_0.Vb1.n10 176.733
R6584 two_stage_opamp_dummy_magic_19_0.Vb1.n12 two_stage_opamp_dummy_magic_19_0.Vb1.n11 176.733
R6585 two_stage_opamp_dummy_magic_19_0.Vb1.n13 two_stage_opamp_dummy_magic_19_0.Vb1.n12 176.733
R6586 two_stage_opamp_dummy_magic_19_0.Vb1.n14 two_stage_opamp_dummy_magic_19_0.Vb1.n13 176.733
R6587 two_stage_opamp_dummy_magic_19_0.Vb1.n15 two_stage_opamp_dummy_magic_19_0.Vb1.n14 176.733
R6588 two_stage_opamp_dummy_magic_19_0.Vb1.n17 two_stage_opamp_dummy_magic_19_0.Vb1.n16 176.733
R6589 two_stage_opamp_dummy_magic_19_0.Vb1.n2 two_stage_opamp_dummy_magic_19_0.Vb1.n1 176.733
R6590 two_stage_opamp_dummy_magic_19_0.Vb1.n8 two_stage_opamp_dummy_magic_19_0.Vb1.n7 176.733
R6591 two_stage_opamp_dummy_magic_19_0.Vb1.n7 two_stage_opamp_dummy_magic_19_0.Vb1.n6 176.733
R6592 two_stage_opamp_dummy_magic_19_0.Vb1.n6 two_stage_opamp_dummy_magic_19_0.Vb1.n5 176.733
R6593 two_stage_opamp_dummy_magic_19_0.Vb1.n5 two_stage_opamp_dummy_magic_19_0.Vb1.n4 176.733
R6594 two_stage_opamp_dummy_magic_19_0.Vb1.n4 two_stage_opamp_dummy_magic_19_0.Vb1.n3 176.733
R6595 two_stage_opamp_dummy_magic_19_0.Vb1.n21 two_stage_opamp_dummy_magic_19_0.Vb1.t15 167.925
R6596 two_stage_opamp_dummy_magic_19_0.Vb1.n26 two_stage_opamp_dummy_magic_19_0.Vb1.n24 161.3
R6597 two_stage_opamp_dummy_magic_19_0.Vb1.n18 two_stage_opamp_dummy_magic_19_0.Vb1.n17 96.4005
R6598 two_stage_opamp_dummy_magic_19_0.Vb1.n9 two_stage_opamp_dummy_magic_19_0.Vb1.n2 96.4005
R6599 two_stage_opamp_dummy_magic_19_0.Vb1.n18 two_stage_opamp_dummy_magic_19_0.Vb1.n15 80.3338
R6600 two_stage_opamp_dummy_magic_19_0.Vb1.n9 two_stage_opamp_dummy_magic_19_0.Vb1.n8 80.3338
R6601 two_stage_opamp_dummy_magic_19_0.Vb1.n21 two_stage_opamp_dummy_magic_19_0.Vb1.n20 54.288
R6602 two_stage_opamp_dummy_magic_19_0.Vb1.n29 two_stage_opamp_dummy_magic_19_0.Vb1.n28 54.288
R6603 two_stage_opamp_dummy_magic_19_0.Vb1.n26 two_stage_opamp_dummy_magic_19_0.Vb1.n25 49.788
R6604 bgr_9_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_19_0.Vb1.n30 45.5943
R6605 two_stage_opamp_dummy_magic_19_0.Vb1.n24 two_stage_opamp_dummy_magic_19_0.Vb1.n23 45.5227
R6606 two_stage_opamp_dummy_magic_19_0.Vb1.n24 two_stage_opamp_dummy_magic_19_0.Vb1.n22 45.5227
R6607 two_stage_opamp_dummy_magic_19_0.Vb1.n30 two_stage_opamp_dummy_magic_19_0.Vb1.n29 25.2193
R6608 two_stage_opamp_dummy_magic_19_0.Vb1.n0 two_stage_opamp_dummy_magic_19_0.Vb1.t0 19.7005
R6609 two_stage_opamp_dummy_magic_19_0.Vb1.n0 two_stage_opamp_dummy_magic_19_0.Vb1.t11 19.7005
R6610 two_stage_opamp_dummy_magic_19_0.Vb1.n25 two_stage_opamp_dummy_magic_19_0.Vb1.t8 16.0005
R6611 two_stage_opamp_dummy_magic_19_0.Vb1.n25 two_stage_opamp_dummy_magic_19_0.Vb1.t2 16.0005
R6612 two_stage_opamp_dummy_magic_19_0.Vb1.n20 two_stage_opamp_dummy_magic_19_0.Vb1.t9 16.0005
R6613 two_stage_opamp_dummy_magic_19_0.Vb1.n20 two_stage_opamp_dummy_magic_19_0.Vb1.t4 16.0005
R6614 two_stage_opamp_dummy_magic_19_0.Vb1.n28 two_stage_opamp_dummy_magic_19_0.Vb1.t6 16.0005
R6615 two_stage_opamp_dummy_magic_19_0.Vb1.n28 two_stage_opamp_dummy_magic_19_0.Vb1.t10 16.0005
R6616 two_stage_opamp_dummy_magic_19_0.Vb1.n27 two_stage_opamp_dummy_magic_19_0.Vb1.n26 4.5005
R6617 two_stage_opamp_dummy_magic_19_0.Vb1.n30 two_stage_opamp_dummy_magic_19_0.Vb1.n19 1.39112
R6618 two_stage_opamp_dummy_magic_19_0.Vb1.n27 two_stage_opamp_dummy_magic_19_0.Vb1.n21 0.563
R6619 two_stage_opamp_dummy_magic_19_0.Vb1.n29 two_stage_opamp_dummy_magic_19_0.Vb1.n27 0.563
R6620 two_stage_opamp_dummy_magic_19_0.VD1.n6 two_stage_opamp_dummy_magic_19_0.VD1.n4 54.8765
R6621 two_stage_opamp_dummy_magic_19_0.VD1.n3 two_stage_opamp_dummy_magic_19_0.VD1.n1 54.8765
R6622 two_stage_opamp_dummy_magic_19_0.VD1.n16 two_stage_opamp_dummy_magic_19_0.VD1.n14 54.788
R6623 two_stage_opamp_dummy_magic_19_0.VD1.n11 two_stage_opamp_dummy_magic_19_0.VD1.n9 54.788
R6624 two_stage_opamp_dummy_magic_19_0.VD1.n6 two_stage_opamp_dummy_magic_19_0.VD1.n5 54.2724
R6625 two_stage_opamp_dummy_magic_19_0.VD1.n3 two_stage_opamp_dummy_magic_19_0.VD1.n2 54.2724
R6626 two_stage_opamp_dummy_magic_19_0.VD1.n18 two_stage_opamp_dummy_magic_19_0.VD1.n17 54.2255
R6627 two_stage_opamp_dummy_magic_19_0.VD1.n16 two_stage_opamp_dummy_magic_19_0.VD1.n15 54.2255
R6628 two_stage_opamp_dummy_magic_19_0.VD1.n13 two_stage_opamp_dummy_magic_19_0.VD1.n12 54.2255
R6629 two_stage_opamp_dummy_magic_19_0.VD1.n11 two_stage_opamp_dummy_magic_19_0.VD1.n10 54.2255
R6630 two_stage_opamp_dummy_magic_19_0.VD1.n8 two_stage_opamp_dummy_magic_19_0.VD1.n0 49.7724
R6631 two_stage_opamp_dummy_magic_19_0.VD1.n5 two_stage_opamp_dummy_magic_19_0.VD1.t7 16.0005
R6632 two_stage_opamp_dummy_magic_19_0.VD1.n5 two_stage_opamp_dummy_magic_19_0.VD1.t12 16.0005
R6633 two_stage_opamp_dummy_magic_19_0.VD1.n0 two_stage_opamp_dummy_magic_19_0.VD1.t9 16.0005
R6634 two_stage_opamp_dummy_magic_19_0.VD1.n0 two_stage_opamp_dummy_magic_19_0.VD1.t4 16.0005
R6635 two_stage_opamp_dummy_magic_19_0.VD1.n17 two_stage_opamp_dummy_magic_19_0.VD1.t17 16.0005
R6636 two_stage_opamp_dummy_magic_19_0.VD1.n17 two_stage_opamp_dummy_magic_19_0.VD1.t3 16.0005
R6637 two_stage_opamp_dummy_magic_19_0.VD1.n15 two_stage_opamp_dummy_magic_19_0.VD1.t14 16.0005
R6638 two_stage_opamp_dummy_magic_19_0.VD1.n15 two_stage_opamp_dummy_magic_19_0.VD1.t18 16.0005
R6639 two_stage_opamp_dummy_magic_19_0.VD1.n14 two_stage_opamp_dummy_magic_19_0.VD1.t1 16.0005
R6640 two_stage_opamp_dummy_magic_19_0.VD1.n14 two_stage_opamp_dummy_magic_19_0.VD1.t20 16.0005
R6641 two_stage_opamp_dummy_magic_19_0.VD1.n12 two_stage_opamp_dummy_magic_19_0.VD1.t15 16.0005
R6642 two_stage_opamp_dummy_magic_19_0.VD1.n12 two_stage_opamp_dummy_magic_19_0.VD1.t2 16.0005
R6643 two_stage_opamp_dummy_magic_19_0.VD1.n10 two_stage_opamp_dummy_magic_19_0.VD1.t16 16.0005
R6644 two_stage_opamp_dummy_magic_19_0.VD1.n10 two_stage_opamp_dummy_magic_19_0.VD1.t21 16.0005
R6645 two_stage_opamp_dummy_magic_19_0.VD1.n9 two_stage_opamp_dummy_magic_19_0.VD1.t19 16.0005
R6646 two_stage_opamp_dummy_magic_19_0.VD1.n9 two_stage_opamp_dummy_magic_19_0.VD1.t0 16.0005
R6647 two_stage_opamp_dummy_magic_19_0.VD1.n2 two_stage_opamp_dummy_magic_19_0.VD1.t10 16.0005
R6648 two_stage_opamp_dummy_magic_19_0.VD1.n2 two_stage_opamp_dummy_magic_19_0.VD1.t5 16.0005
R6649 two_stage_opamp_dummy_magic_19_0.VD1.n1 two_stage_opamp_dummy_magic_19_0.VD1.t11 16.0005
R6650 two_stage_opamp_dummy_magic_19_0.VD1.n1 two_stage_opamp_dummy_magic_19_0.VD1.t6 16.0005
R6651 two_stage_opamp_dummy_magic_19_0.VD1.n4 two_stage_opamp_dummy_magic_19_0.VD1.t8 16.0005
R6652 two_stage_opamp_dummy_magic_19_0.VD1.n4 two_stage_opamp_dummy_magic_19_0.VD1.t13 16.0005
R6653 two_stage_opamp_dummy_magic_19_0.VD1 two_stage_opamp_dummy_magic_19_0.VD1.n19 4.813
R6654 two_stage_opamp_dummy_magic_19_0.VD1.n8 two_stage_opamp_dummy_magic_19_0.VD1.n7 4.5005
R6655 two_stage_opamp_dummy_magic_19_0.VD1.n7 two_stage_opamp_dummy_magic_19_0.VD1.n3 0.604667
R6656 two_stage_opamp_dummy_magic_19_0.VD1.n7 two_stage_opamp_dummy_magic_19_0.VD1.n6 0.604667
R6657 two_stage_opamp_dummy_magic_19_0.VD1.n18 two_stage_opamp_dummy_magic_19_0.VD1.n16 0.563
R6658 two_stage_opamp_dummy_magic_19_0.VD1.n13 two_stage_opamp_dummy_magic_19_0.VD1.n11 0.563
R6659 two_stage_opamp_dummy_magic_19_0.VD1 two_stage_opamp_dummy_magic_19_0.VD1.n8 0.443208
R6660 two_stage_opamp_dummy_magic_19_0.VD1.n19 two_stage_opamp_dummy_magic_19_0.VD1.n18 0.234875
R6661 two_stage_opamp_dummy_magic_19_0.VD1.n19 two_stage_opamp_dummy_magic_19_0.VD1.n13 0.234875
R6662 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t4 525.38
R6663 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t5 525.38
R6664 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t8 525.38
R6665 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t9 525.38
R6666 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n6 328.476
R6667 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n2 328.476
R6668 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t6 281.168
R6669 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t2 281.168
R6670 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t3 281.168
R6671 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t7 281.168
R6672 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t1 115.388
R6673 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t0 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n7 115.388
R6674 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n5 89.9738
R6675 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n4 89.9738
R6676 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n1 89.9738
R6677 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n0 89.9738
R6678 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n3 39.2505
R6679 a_6930_22564.t0 a_6930_22564.t1 178.133
R6680 bgr_9_0.PFET_GATE_10uA.n16 bgr_9_0.PFET_GATE_10uA.t18 565.114
R6681 bgr_9_0.PFET_GATE_10uA.n19 bgr_9_0.PFET_GATE_10uA.t15 530.201
R6682 bgr_9_0.PFET_GATE_10uA.n21 bgr_9_0.PFET_GATE_10uA.t14 409.7
R6683 bgr_9_0.PFET_GATE_10uA.n6 bgr_9_0.PFET_GATE_10uA.t12 369.534
R6684 bgr_9_0.PFET_GATE_10uA.n5 bgr_9_0.PFET_GATE_10uA.t11 369.534
R6685 bgr_9_0.PFET_GATE_10uA.n2 bgr_9_0.PFET_GATE_10uA.t20 369.534
R6686 bgr_9_0.PFET_GATE_10uA.n1 bgr_9_0.PFET_GATE_10uA.t19 369.534
R6687 bgr_9_0.PFET_GATE_10uA.n19 bgr_9_0.PFET_GATE_10uA.t21 353.467
R6688 bgr_9_0.PFET_GATE_10uA.n20 bgr_9_0.PFET_GATE_10uA.t10 353.467
R6689 bgr_9_0.PFET_GATE_10uA.n10 bgr_9_0.PFET_GATE_10uA.n8 346.825
R6690 bgr_9_0.PFET_GATE_10uA.n12 bgr_9_0.PFET_GATE_10uA.n11 344.7
R6691 bgr_9_0.PFET_GATE_10uA.n10 bgr_9_0.PFET_GATE_10uA.n9 344.7
R6692 bgr_9_0.PFET_GATE_10uA.n15 bgr_9_0.PFET_GATE_10uA.n14 340.2
R6693 bgr_9_0.PFET_GATE_10uA.n0 bgr_9_0.PFET_GATE_10uA.t17 325.351
R6694 bgr_9_0.PFET_GATE_10uA.n4 bgr_9_0.PFET_GATE_10uA.n0 202.364
R6695 bgr_9_0.PFET_GATE_10uA.n6 bgr_9_0.PFET_GATE_10uA.t22 192.8
R6696 bgr_9_0.PFET_GATE_10uA.n5 bgr_9_0.PFET_GATE_10uA.t16 192.8
R6697 bgr_9_0.PFET_GATE_10uA.n2 bgr_9_0.PFET_GATE_10uA.t13 192.8
R6698 bgr_9_0.PFET_GATE_10uA.n1 bgr_9_0.PFET_GATE_10uA.t24 192.8
R6699 bgr_9_0.PFET_GATE_10uA.n0 bgr_9_0.PFET_GATE_10uA.t23 192.8
R6700 bgr_9_0.PFET_GATE_10uA.n20 bgr_9_0.PFET_GATE_10uA.n19 176.733
R6701 bgr_9_0.PFET_GATE_10uA.n18 bgr_9_0.PFET_GATE_10uA.n7 168.166
R6702 bgr_9_0.PFET_GATE_10uA bgr_9_0.PFET_GATE_10uA.n21 166.071
R6703 bgr_9_0.PFET_GATE_10uA.n4 bgr_9_0.PFET_GATE_10uA.n3 166.071
R6704 bgr_9_0.PFET_GATE_10uA.n16 bgr_9_0.PFET_GATE_10uA.t6 137.386
R6705 bgr_9_0.PFET_GATE_10uA.n13 bgr_9_0.PFET_GATE_10uA.t7 116.584
R6706 bgr_9_0.PFET_GATE_10uA.n7 bgr_9_0.PFET_GATE_10uA.n6 56.2338
R6707 bgr_9_0.PFET_GATE_10uA.n7 bgr_9_0.PFET_GATE_10uA.n5 56.2338
R6708 bgr_9_0.PFET_GATE_10uA.n21 bgr_9_0.PFET_GATE_10uA.n20 56.2338
R6709 bgr_9_0.PFET_GATE_10uA.n3 bgr_9_0.PFET_GATE_10uA.n2 56.2338
R6710 bgr_9_0.PFET_GATE_10uA.n3 bgr_9_0.PFET_GATE_10uA.n1 56.2338
R6711 bgr_9_0.PFET_GATE_10uA.n14 bgr_9_0.PFET_GATE_10uA.t9 39.4005
R6712 bgr_9_0.PFET_GATE_10uA.n14 bgr_9_0.PFET_GATE_10uA.t1 39.4005
R6713 bgr_9_0.PFET_GATE_10uA.n11 bgr_9_0.PFET_GATE_10uA.t3 39.4005
R6714 bgr_9_0.PFET_GATE_10uA.n11 bgr_9_0.PFET_GATE_10uA.t5 39.4005
R6715 bgr_9_0.PFET_GATE_10uA.n9 bgr_9_0.PFET_GATE_10uA.t2 39.4005
R6716 bgr_9_0.PFET_GATE_10uA.n9 bgr_9_0.PFET_GATE_10uA.t4 39.4005
R6717 bgr_9_0.PFET_GATE_10uA.n8 bgr_9_0.PFET_GATE_10uA.t0 39.4005
R6718 bgr_9_0.PFET_GATE_10uA.n8 bgr_9_0.PFET_GATE_10uA.t8 39.4005
R6719 bgr_9_0.PFET_GATE_10uA.n18 bgr_9_0.PFET_GATE_10uA.n17 27.5005
R6720 bgr_9_0.PFET_GATE_10uA.n17 bgr_9_0.PFET_GATE_10uA.n15 9.53175
R6721 bgr_9_0.PFET_GATE_10uA bgr_9_0.PFET_GATE_10uA.n4 5.2505
R6722 bgr_9_0.PFET_GATE_10uA.n15 bgr_9_0.PFET_GATE_10uA.n13 4.5005
R6723 bgr_9_0.PFET_GATE_10uA bgr_9_0.PFET_GATE_10uA.n18 2.34425
R6724 bgr_9_0.PFET_GATE_10uA.n12 bgr_9_0.PFET_GATE_10uA.n10 2.1255
R6725 bgr_9_0.PFET_GATE_10uA.n13 bgr_9_0.PFET_GATE_10uA.n12 2.1255
R6726 bgr_9_0.PFET_GATE_10uA.n17 bgr_9_0.PFET_GATE_10uA.n16 1.78175
R6727 bgr_9_0.cap_res1.t0 bgr_9_0.cap_res1.t10 121.245
R6728 bgr_9_0.cap_res1.t16 bgr_9_0.cap_res1.t19 0.1603
R6729 bgr_9_0.cap_res1.t9 bgr_9_0.cap_res1.t15 0.1603
R6730 bgr_9_0.cap_res1.t14 bgr_9_0.cap_res1.t18 0.1603
R6731 bgr_9_0.cap_res1.t7 bgr_9_0.cap_res1.t13 0.1603
R6732 bgr_9_0.cap_res1.t1 bgr_9_0.cap_res1.t6 0.1603
R6733 bgr_9_0.cap_res1.n1 bgr_9_0.cap_res1.t17 0.159278
R6734 bgr_9_0.cap_res1.n2 bgr_9_0.cap_res1.t2 0.159278
R6735 bgr_9_0.cap_res1.n3 bgr_9_0.cap_res1.t8 0.159278
R6736 bgr_9_0.cap_res1.n4 bgr_9_0.cap_res1.t3 0.159278
R6737 bgr_9_0.cap_res1.n4 bgr_9_0.cap_res1.t16 0.1368
R6738 bgr_9_0.cap_res1.n4 bgr_9_0.cap_res1.t12 0.1368
R6739 bgr_9_0.cap_res1.n3 bgr_9_0.cap_res1.t9 0.1368
R6740 bgr_9_0.cap_res1.n3 bgr_9_0.cap_res1.t5 0.1368
R6741 bgr_9_0.cap_res1.n2 bgr_9_0.cap_res1.t14 0.1368
R6742 bgr_9_0.cap_res1.n2 bgr_9_0.cap_res1.t11 0.1368
R6743 bgr_9_0.cap_res1.n1 bgr_9_0.cap_res1.t7 0.1368
R6744 bgr_9_0.cap_res1.n1 bgr_9_0.cap_res1.t4 0.1368
R6745 bgr_9_0.cap_res1.n0 bgr_9_0.cap_res1.t1 0.1368
R6746 bgr_9_0.cap_res1.n0 bgr_9_0.cap_res1.t20 0.1368
R6747 bgr_9_0.cap_res1.t17 bgr_9_0.cap_res1.n0 0.00152174
R6748 bgr_9_0.cap_res1.t2 bgr_9_0.cap_res1.n1 0.00152174
R6749 bgr_9_0.cap_res1.t8 bgr_9_0.cap_res1.n2 0.00152174
R6750 bgr_9_0.cap_res1.t3 bgr_9_0.cap_res1.n3 0.00152174
R6751 bgr_9_0.cap_res1.t10 bgr_9_0.cap_res1.n4 0.00152174
R6752 bgr_9_0.V_mir2.n13 bgr_9_0.V_mir2.n12 330.901
R6753 bgr_9_0.V_mir2.n8 bgr_9_0.V_mir2.n7 330.901
R6754 bgr_9_0.V_mir2.n20 bgr_9_0.V_mir2.n19 330.901
R6755 bgr_9_0.V_mir2.n16 bgr_9_0.V_mir2.t21 310.488
R6756 bgr_9_0.V_mir2.n9 bgr_9_0.V_mir2.t22 310.488
R6757 bgr_9_0.V_mir2.n4 bgr_9_0.V_mir2.t20 310.488
R6758 bgr_9_0.V_mir2.n2 bgr_9_0.V_mir2.t14 278.312
R6759 bgr_9_0.V_mir2.n2 bgr_9_0.V_mir2.n1 228.939
R6760 bgr_9_0.V_mir2.n3 bgr_9_0.V_mir2.n0 224.439
R6761 bgr_9_0.V_mir2.n18 bgr_9_0.V_mir2.t10 184.097
R6762 bgr_9_0.V_mir2.n11 bgr_9_0.V_mir2.t8 184.097
R6763 bgr_9_0.V_mir2.n6 bgr_9_0.V_mir2.t0 184.097
R6764 bgr_9_0.V_mir2.n17 bgr_9_0.V_mir2.n16 167.094
R6765 bgr_9_0.V_mir2.n10 bgr_9_0.V_mir2.n9 167.094
R6766 bgr_9_0.V_mir2.n5 bgr_9_0.V_mir2.n4 167.094
R6767 bgr_9_0.V_mir2.n13 bgr_9_0.V_mir2.n11 152
R6768 bgr_9_0.V_mir2.n8 bgr_9_0.V_mir2.n6 152
R6769 bgr_9_0.V_mir2.n19 bgr_9_0.V_mir2.n18 152
R6770 bgr_9_0.V_mir2.n16 bgr_9_0.V_mir2.t19 120.501
R6771 bgr_9_0.V_mir2.n17 bgr_9_0.V_mir2.t6 120.501
R6772 bgr_9_0.V_mir2.n9 bgr_9_0.V_mir2.t18 120.501
R6773 bgr_9_0.V_mir2.n10 bgr_9_0.V_mir2.t2 120.501
R6774 bgr_9_0.V_mir2.n4 bgr_9_0.V_mir2.t17 120.501
R6775 bgr_9_0.V_mir2.n5 bgr_9_0.V_mir2.t4 120.501
R6776 bgr_9_0.V_mir2.n1 bgr_9_0.V_mir2.t16 48.0005
R6777 bgr_9_0.V_mir2.n1 bgr_9_0.V_mir2.t12 48.0005
R6778 bgr_9_0.V_mir2.n0 bgr_9_0.V_mir2.t15 48.0005
R6779 bgr_9_0.V_mir2.n0 bgr_9_0.V_mir2.t13 48.0005
R6780 bgr_9_0.V_mir2.n18 bgr_9_0.V_mir2.n17 40.7027
R6781 bgr_9_0.V_mir2.n11 bgr_9_0.V_mir2.n10 40.7027
R6782 bgr_9_0.V_mir2.n6 bgr_9_0.V_mir2.n5 40.7027
R6783 bgr_9_0.V_mir2.n12 bgr_9_0.V_mir2.t3 39.4005
R6784 bgr_9_0.V_mir2.n12 bgr_9_0.V_mir2.t9 39.4005
R6785 bgr_9_0.V_mir2.n7 bgr_9_0.V_mir2.t5 39.4005
R6786 bgr_9_0.V_mir2.n7 bgr_9_0.V_mir2.t1 39.4005
R6787 bgr_9_0.V_mir2.n20 bgr_9_0.V_mir2.t7 39.4005
R6788 bgr_9_0.V_mir2.t11 bgr_9_0.V_mir2.n20 39.4005
R6789 bgr_9_0.V_mir2.n14 bgr_9_0.V_mir2.n13 15.8005
R6790 bgr_9_0.V_mir2.n14 bgr_9_0.V_mir2.n8 15.8005
R6791 bgr_9_0.V_mir2.n19 bgr_9_0.V_mir2.n15 9.3005
R6792 bgr_9_0.V_mir2.n3 bgr_9_0.V_mir2.n2 5.8755
R6793 bgr_9_0.V_mir2.n15 bgr_9_0.V_mir2.n14 4.5005
R6794 bgr_9_0.V_mir2.n15 bgr_9_0.V_mir2.n3 0.78175
R6795 bgr_9_0.Vin-.n7 bgr_9_0.Vin-.t12 688.859
R6796 bgr_9_0.Vin-.n9 bgr_9_0.Vin-.n8 514.134
R6797 bgr_9_0.Vin-.n6 bgr_9_0.Vin-.n5 356.95
R6798 bgr_9_0.Vin-.n11 bgr_9_0.Vin-.n10 213.4
R6799 bgr_9_0.Vin-.n7 bgr_9_0.Vin-.t8 174.726
R6800 bgr_9_0.Vin-.n8 bgr_9_0.Vin-.t10 174.726
R6801 bgr_9_0.Vin-.n9 bgr_9_0.Vin-.t9 174.726
R6802 bgr_9_0.Vin-.n10 bgr_9_0.Vin-.t11 174.726
R6803 bgr_9_0.Vin-.n4 bgr_9_0.Vin-.n2 172.585
R6804 bgr_9_0.Vin-.n4 bgr_9_0.Vin-.n3 168.21
R6805 bgr_9_0.Vin-.n8 bgr_9_0.Vin-.n7 128.534
R6806 bgr_9_0.Vin-.n10 bgr_9_0.Vin-.n9 128.534
R6807 bgr_9_0.Vin-.n12 bgr_9_0.Vin-.t1 119.099
R6808 bgr_9_0.Vin-.n16 bgr_9_0.Vin-.n15 83.5719
R6809 bgr_9_0.Vin-.n1 bgr_9_0.Vin-.n0 83.5719
R6810 bgr_9_0.Vin-.n19 bgr_9_0.Vin-.n1 73.8495
R6811 bgr_9_0.Vin-.t2 bgr_9_0.Vin-.n14 65.0341
R6812 bgr_9_0.Vin-.n5 bgr_9_0.Vin-.t0 39.4005
R6813 bgr_9_0.Vin-.n5 bgr_9_0.Vin-.t7 39.4005
R6814 bgr_9_0.Vin-.n13 bgr_9_0.Vin-.n12 28.813
R6815 bgr_9_0.Vin-.n15 bgr_9_0.Vin-.n1 26.074
R6816 bgr_9_0.Vin-.n12 bgr_9_0.Vin-.n11 16.188
R6817 bgr_9_0.Vin-.n3 bgr_9_0.Vin-.t3 13.1338
R6818 bgr_9_0.Vin-.n3 bgr_9_0.Vin-.t5 13.1338
R6819 bgr_9_0.Vin-.n2 bgr_9_0.Vin-.t6 13.1338
R6820 bgr_9_0.Vin-.n2 bgr_9_0.Vin-.t4 13.1338
R6821 bgr_9_0.Vin-.n11 bgr_9_0.Vin-.n6 11.2193
R6822 bgr_9_0.Vin-.n6 bgr_9_0.Vin-.n4 3.8755
R6823 bgr_9_0.Vin-.n16 bgr_9_0.Vin-.n14 1.56483
R6824 bgr_9_0.Vin-.n18 bgr_9_0.Vin-.n17 1.5505
R6825 bgr_9_0.Vin-.n17 bgr_9_0.Vin-.n0 0.885803
R6826 bgr_9_0.Vin-.n17 bgr_9_0.Vin-.n16 0.77514
R6827 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_9_0.Vin-.n0 0.756696
R6828 bgr_9_0.Vin-.n19 bgr_9_0.Vin-.n18 0.711459
R6829 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_9_0.Vin-.n19 0.576566
R6830 bgr_9_0.Vin-.n14 bgr_9_0.Vin-.n13 0.531499
R6831 bgr_9_0.Vin-.n15 bgr_9_0.Vin-.t2 0.290206
R6832 bgr_9_0.Vin-.n18 bgr_9_0.Vin-.n13 0.00817857
R6833 a_5820_2720.t0 a_5820_2720.t1 169.905
R6834 bgr_9_0.V_p_1.n2 bgr_9_0.V_p_1.n0 263.933
R6835 bgr_9_0.V_p_1.n6 bgr_9_0.V_p_1.n4 263.933
R6836 bgr_9_0.V_p_1.n2 bgr_9_0.V_p_1.n1 206.333
R6837 bgr_9_0.V_p_1.n7 bgr_9_0.V_p_1.n3 206.333
R6838 bgr_9_0.V_p_1.n6 bgr_9_0.V_p_1.n5 206.333
R6839 bgr_9_0.V_p_1 bgr_9_0.V_p_1.t10 120.677
R6840 bgr_9_0.V_p_1.n7 bgr_9_0.V_p_1.n2 57.6005
R6841 bgr_9_0.V_p_1.n7 bgr_9_0.V_p_1.n6 57.6005
R6842 bgr_9_0.V_p_1.n0 bgr_9_0.V_p_1.t8 48.0005
R6843 bgr_9_0.V_p_1.n0 bgr_9_0.V_p_1.t1 48.0005
R6844 bgr_9_0.V_p_1.n1 bgr_9_0.V_p_1.t3 48.0005
R6845 bgr_9_0.V_p_1.n1 bgr_9_0.V_p_1.t5 48.0005
R6846 bgr_9_0.V_p_1.n3 bgr_9_0.V_p_1.t9 48.0005
R6847 bgr_9_0.V_p_1.n3 bgr_9_0.V_p_1.t2 48.0005
R6848 bgr_9_0.V_p_1.n4 bgr_9_0.V_p_1.t7 48.0005
R6849 bgr_9_0.V_p_1.n4 bgr_9_0.V_p_1.t0 48.0005
R6850 bgr_9_0.V_p_1.n5 bgr_9_0.V_p_1.t4 48.0005
R6851 bgr_9_0.V_p_1.n5 bgr_9_0.V_p_1.t6 48.0005
R6852 bgr_9_0.V_p_1 bgr_9_0.V_p_1.n7 13.7338
R6853 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t5 661.375
R6854 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t2 661.375
R6855 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n5 213.131
R6856 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t6 213.131
R6857 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t0 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t3 146.155
R6858 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t0 146.155
R6859 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n0 78.7265
R6860 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t4 76.2576
R6861 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n6 76.2576
R6862 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n2 71.388
R6863 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t1 11.2576
R6864 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t7 11.2576
R6865 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t9 11.2576
R6866 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.t10 11.2576
R6867 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n3 5.1255
R6868 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n1 4.7505
R6869 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n4 1.888
R6870 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_19_0.Vb2_Vb3.n1 1.888
R6871 VIN-.n8 VIN-.t1 635.702
R6872 VIN-.n2 VIN-.t2 449.868
R6873 VIN-.n0 VIN-.t4 449.868
R6874 VIN-.n8 VIN-.n7 310.401
R6875 VIN-.n7 VIN-.t10 273.134
R6876 VIN-.n2 VIN-.t7 273.134
R6877 VIN-.n3 VIN-.t3 273.134
R6878 VIN-.n4 VIN-.t8 273.134
R6879 VIN-.n5 VIN-.t0 273.134
R6880 VIN-.n6 VIN-.t6 273.134
R6881 VIN-.n1 VIN-.t5 273.134
R6882 VIN-.n0 VIN-.t9 273.134
R6883 VIN-.n1 VIN-.n0 176.733
R6884 VIN-.n7 VIN-.n1 176.733
R6885 VIN-.n7 VIN-.n6 176.733
R6886 VIN-.n6 VIN-.n5 176.733
R6887 VIN-.n5 VIN-.n4 176.733
R6888 VIN-.n4 VIN-.n3 176.733
R6889 VIN-.n3 VIN-.n2 176.733
R6890 VIN- VIN-.n8 1.60988
R6891 two_stage_opamp_dummy_magic_19_0.Vb1_2.n1 two_stage_opamp_dummy_magic_19_0.Vb1_2.t0 71.6942
R6892 two_stage_opamp_dummy_magic_19_0.Vb1_2.n1 two_stage_opamp_dummy_magic_19_0.Vb1_2.n0 54.8505
R6893 two_stage_opamp_dummy_magic_19_0.Vb1_2.n2 two_stage_opamp_dummy_magic_19_0.Vb1_2.n1 54.288
R6894 two_stage_opamp_dummy_magic_19_0.Vb1_2.n0 two_stage_opamp_dummy_magic_19_0.Vb1_2.t4 16.0005
R6895 two_stage_opamp_dummy_magic_19_0.Vb1_2.n0 two_stage_opamp_dummy_magic_19_0.Vb1_2.t2 16.0005
R6896 two_stage_opamp_dummy_magic_19_0.Vb1_2.n2 two_stage_opamp_dummy_magic_19_0.Vb1_2.t1 16.0005
R6897 two_stage_opamp_dummy_magic_19_0.Vb1_2.t3 two_stage_opamp_dummy_magic_19_0.Vb1_2.n2 16.0005
R6898 two_stage_opamp_dummy_magic_19_0.VD4.n21 two_stage_opamp_dummy_magic_19_0.VD4.t23 652.076
R6899 two_stage_opamp_dummy_magic_19_0.VD4.n24 two_stage_opamp_dummy_magic_19_0.VD4.t20 652.076
R6900 two_stage_opamp_dummy_magic_19_0.VD4.t24 two_stage_opamp_dummy_magic_19_0.VD4.n22 211.625
R6901 two_stage_opamp_dummy_magic_19_0.VD4.n23 two_stage_opamp_dummy_magic_19_0.VD4.t21 211.625
R6902 two_stage_opamp_dummy_magic_19_0.VD4.t10 two_stage_opamp_dummy_magic_19_0.VD4.t24 146.155
R6903 two_stage_opamp_dummy_magic_19_0.VD4.t6 two_stage_opamp_dummy_magic_19_0.VD4.t10 146.155
R6904 two_stage_opamp_dummy_magic_19_0.VD4.t12 two_stage_opamp_dummy_magic_19_0.VD4.t6 146.155
R6905 two_stage_opamp_dummy_magic_19_0.VD4.t16 two_stage_opamp_dummy_magic_19_0.VD4.t12 146.155
R6906 two_stage_opamp_dummy_magic_19_0.VD4.t0 two_stage_opamp_dummy_magic_19_0.VD4.t16 146.155
R6907 two_stage_opamp_dummy_magic_19_0.VD4.t2 two_stage_opamp_dummy_magic_19_0.VD4.t0 146.155
R6908 two_stage_opamp_dummy_magic_19_0.VD4.t4 two_stage_opamp_dummy_magic_19_0.VD4.t2 146.155
R6909 two_stage_opamp_dummy_magic_19_0.VD4.t8 two_stage_opamp_dummy_magic_19_0.VD4.t4 146.155
R6910 two_stage_opamp_dummy_magic_19_0.VD4.t14 two_stage_opamp_dummy_magic_19_0.VD4.t8 146.155
R6911 two_stage_opamp_dummy_magic_19_0.VD4.t18 two_stage_opamp_dummy_magic_19_0.VD4.t14 146.155
R6912 two_stage_opamp_dummy_magic_19_0.VD4.t21 two_stage_opamp_dummy_magic_19_0.VD4.t18 146.155
R6913 two_stage_opamp_dummy_magic_19_0.VD4.n22 two_stage_opamp_dummy_magic_19_0.VD4.t25 76.2576
R6914 two_stage_opamp_dummy_magic_19_0.VD4.n23 two_stage_opamp_dummy_magic_19_0.VD4.t22 76.2576
R6915 two_stage_opamp_dummy_magic_19_0.VD4.n2 two_stage_opamp_dummy_magic_19_0.VD4.n0 72.013
R6916 two_stage_opamp_dummy_magic_19_0.VD4.n14 two_stage_opamp_dummy_magic_19_0.VD4.n13 71.388
R6917 two_stage_opamp_dummy_magic_19_0.VD4.n16 two_stage_opamp_dummy_magic_19_0.VD4.n15 71.388
R6918 two_stage_opamp_dummy_magic_19_0.VD4.n18 two_stage_opamp_dummy_magic_19_0.VD4.n17 71.388
R6919 two_stage_opamp_dummy_magic_19_0.VD4.n20 two_stage_opamp_dummy_magic_19_0.VD4.n19 71.388
R6920 two_stage_opamp_dummy_magic_19_0.VD4.n10 two_stage_opamp_dummy_magic_19_0.VD4.n9 71.388
R6921 two_stage_opamp_dummy_magic_19_0.VD4.n8 two_stage_opamp_dummy_magic_19_0.VD4.n7 71.388
R6922 two_stage_opamp_dummy_magic_19_0.VD4.n6 two_stage_opamp_dummy_magic_19_0.VD4.n5 71.388
R6923 two_stage_opamp_dummy_magic_19_0.VD4.n4 two_stage_opamp_dummy_magic_19_0.VD4.n3 71.388
R6924 two_stage_opamp_dummy_magic_19_0.VD4.n2 two_stage_opamp_dummy_magic_19_0.VD4.n1 71.388
R6925 two_stage_opamp_dummy_magic_19_0.VD4.n12 two_stage_opamp_dummy_magic_19_0.VD4.n11 71.388
R6926 two_stage_opamp_dummy_magic_19_0.VD4.n24 two_stage_opamp_dummy_magic_19_0.VD4.n23 46.0195
R6927 two_stage_opamp_dummy_magic_19_0.VD4.n22 two_stage_opamp_dummy_magic_19_0.VD4.n21 46.0195
R6928 two_stage_opamp_dummy_magic_19_0.VD4.n21 two_stage_opamp_dummy_magic_19_0.VD4.n20 14.4255
R6929 two_stage_opamp_dummy_magic_19_0.VD4.n25 two_stage_opamp_dummy_magic_19_0.VD4.n24 13.8005
R6930 two_stage_opamp_dummy_magic_19_0.VD4.n13 two_stage_opamp_dummy_magic_19_0.VD4.t5 11.2576
R6931 two_stage_opamp_dummy_magic_19_0.VD4.n13 two_stage_opamp_dummy_magic_19_0.VD4.t9 11.2576
R6932 two_stage_opamp_dummy_magic_19_0.VD4.n15 two_stage_opamp_dummy_magic_19_0.VD4.t1 11.2576
R6933 two_stage_opamp_dummy_magic_19_0.VD4.n15 two_stage_opamp_dummy_magic_19_0.VD4.t3 11.2576
R6934 two_stage_opamp_dummy_magic_19_0.VD4.n17 two_stage_opamp_dummy_magic_19_0.VD4.t13 11.2576
R6935 two_stage_opamp_dummy_magic_19_0.VD4.n17 two_stage_opamp_dummy_magic_19_0.VD4.t17 11.2576
R6936 two_stage_opamp_dummy_magic_19_0.VD4.n19 two_stage_opamp_dummy_magic_19_0.VD4.t11 11.2576
R6937 two_stage_opamp_dummy_magic_19_0.VD4.n19 two_stage_opamp_dummy_magic_19_0.VD4.t7 11.2576
R6938 two_stage_opamp_dummy_magic_19_0.VD4.n9 two_stage_opamp_dummy_magic_19_0.VD4.t36 11.2576
R6939 two_stage_opamp_dummy_magic_19_0.VD4.n9 two_stage_opamp_dummy_magic_19_0.VD4.t27 11.2576
R6940 two_stage_opamp_dummy_magic_19_0.VD4.n7 two_stage_opamp_dummy_magic_19_0.VD4.t30 11.2576
R6941 two_stage_opamp_dummy_magic_19_0.VD4.n7 two_stage_opamp_dummy_magic_19_0.VD4.t33 11.2576
R6942 two_stage_opamp_dummy_magic_19_0.VD4.n5 two_stage_opamp_dummy_magic_19_0.VD4.t34 11.2576
R6943 two_stage_opamp_dummy_magic_19_0.VD4.n5 two_stage_opamp_dummy_magic_19_0.VD4.t35 11.2576
R6944 two_stage_opamp_dummy_magic_19_0.VD4.n3 two_stage_opamp_dummy_magic_19_0.VD4.t26 11.2576
R6945 two_stage_opamp_dummy_magic_19_0.VD4.n3 two_stage_opamp_dummy_magic_19_0.VD4.t28 11.2576
R6946 two_stage_opamp_dummy_magic_19_0.VD4.n1 two_stage_opamp_dummy_magic_19_0.VD4.t31 11.2576
R6947 two_stage_opamp_dummy_magic_19_0.VD4.n1 two_stage_opamp_dummy_magic_19_0.VD4.t29 11.2576
R6948 two_stage_opamp_dummy_magic_19_0.VD4.n0 two_stage_opamp_dummy_magic_19_0.VD4.t32 11.2576
R6949 two_stage_opamp_dummy_magic_19_0.VD4.n0 two_stage_opamp_dummy_magic_19_0.VD4.t37 11.2576
R6950 two_stage_opamp_dummy_magic_19_0.VD4.n11 two_stage_opamp_dummy_magic_19_0.VD4.t15 11.2576
R6951 two_stage_opamp_dummy_magic_19_0.VD4.n11 two_stage_opamp_dummy_magic_19_0.VD4.t19 11.2576
R6952 two_stage_opamp_dummy_magic_19_0.VD4.n26 two_stage_opamp_dummy_magic_19_0.VD4.n10 8.21925
R6953 two_stage_opamp_dummy_magic_19_0.VD4.n26 two_stage_opamp_dummy_magic_19_0.VD4.n25 5.8755
R6954 two_stage_opamp_dummy_magic_19_0.VD4.n4 two_stage_opamp_dummy_magic_19_0.VD4.n2 0.6255
R6955 two_stage_opamp_dummy_magic_19_0.VD4.n6 two_stage_opamp_dummy_magic_19_0.VD4.n4 0.6255
R6956 two_stage_opamp_dummy_magic_19_0.VD4.n8 two_stage_opamp_dummy_magic_19_0.VD4.n6 0.6255
R6957 two_stage_opamp_dummy_magic_19_0.VD4.n10 two_stage_opamp_dummy_magic_19_0.VD4.n8 0.6255
R6958 two_stage_opamp_dummy_magic_19_0.VD4.n25 two_stage_opamp_dummy_magic_19_0.VD4.n12 0.6255
R6959 two_stage_opamp_dummy_magic_19_0.VD4.n20 two_stage_opamp_dummy_magic_19_0.VD4.n18 0.6255
R6960 two_stage_opamp_dummy_magic_19_0.VD4.n18 two_stage_opamp_dummy_magic_19_0.VD4.n16 0.6255
R6961 two_stage_opamp_dummy_magic_19_0.VD4.n16 two_stage_opamp_dummy_magic_19_0.VD4.n14 0.6255
R6962 two_stage_opamp_dummy_magic_19_0.VD4.n14 two_stage_opamp_dummy_magic_19_0.VD4.n12 0.6255
R6963 two_stage_opamp_dummy_magic_19_0.VD4 two_stage_opamp_dummy_magic_19_0.VD4.n26 0.063
R6964 VIN+.n8 VIN+.t7 635.702
R6965 VIN+.n5 VIN+.t4 449.868
R6966 VIN+.n0 VIN+.t8 449.868
R6967 VIN+.n8 VIN+.n7 310.401
R6968 VIN+.n7 VIN+.t6 273.134
R6969 VIN+.n5 VIN+.t10 273.134
R6970 VIN+.n6 VIN+.t1 273.134
R6971 VIN+.n4 VIN+.t0 273.134
R6972 VIN+.n3 VIN+.t5 273.134
R6973 VIN+.n2 VIN+.t3 273.134
R6974 VIN+.n1 VIN+.t9 273.134
R6975 VIN+.n0 VIN+.t2 273.134
R6976 VIN+.n1 VIN+.n0 176.733
R6977 VIN+.n2 VIN+.n1 176.733
R6978 VIN+.n3 VIN+.n2 176.733
R6979 VIN+.n4 VIN+.n3 176.733
R6980 VIN+.n7 VIN+.n4 176.733
R6981 VIN+.n7 VIN+.n6 176.733
R6982 VIN+.n6 VIN+.n5 176.733
R6983 VIN+ VIN+.n8 1.60988
R6984 bgr_9_0.START_UP.n4 bgr_9_0.START_UP.t6 238.322
R6985 bgr_9_0.START_UP.n4 bgr_9_0.START_UP.t7 238.322
R6986 bgr_9_0.START_UP.n3 bgr_9_0.START_UP.n1 175.118
R6987 bgr_9_0.START_UP.n3 bgr_9_0.START_UP.n2 168.493
R6988 bgr_9_0.START_UP.n5 bgr_9_0.START_UP.n4 166.925
R6989 bgr_9_0.START_UP.n0 bgr_9_0.START_UP.t1 116.501
R6990 bgr_9_0.START_UP.n0 bgr_9_0.START_UP.t0 82.7823
R6991 bgr_9_0.START_UP bgr_9_0.START_UP.n0 35.8817
R6992 bgr_9_0.START_UP bgr_9_0.START_UP.n5 13.4693
R6993 bgr_9_0.START_UP.n1 bgr_9_0.START_UP.t2 13.1338
R6994 bgr_9_0.START_UP.n1 bgr_9_0.START_UP.t4 13.1338
R6995 bgr_9_0.START_UP.n2 bgr_9_0.START_UP.t3 13.1338
R6996 bgr_9_0.START_UP.n2 bgr_9_0.START_UP.t5 13.1338
R6997 bgr_9_0.START_UP.n5 bgr_9_0.START_UP.n3 4.21925
R6998 a_14170_2720.t0 a_14170_2720.t1 169.905
R6999 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n0 150.451
R7000 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n1 140.201
R7001 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t0 118.861
R7002 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n2 37.4067
R7003 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n12 33.83
R7004 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n3 30.038
R7005 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n10 29.4755
R7006 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n8 29.4755
R7007 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n6 29.4755
R7008 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n4 29.4755
R7009 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t13 24.0005
R7010 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t11 24.0005
R7011 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t14 24.0005
R7012 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t12 24.0005
R7013 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t2 8.0005
R7014 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t6 8.0005
R7015 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t3 8.0005
R7016 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t7 8.0005
R7017 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t4 8.0005
R7018 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t8 8.0005
R7019 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t1 8.0005
R7020 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t10 8.0005
R7021 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t5 8.0005
R7022 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t9 8.0005
R7023 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n11 5.6255
R7024 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n5 0.563
R7025 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n7 0.563
R7026 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n9 0.563
R7027 bgr_9_0.V_CMFB_S4 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n13 0.047375
R7028 two_stage_opamp_dummy_magic_19_0.V_err_p.n1 two_stage_opamp_dummy_magic_19_0.V_err_p.n0 208.829
R7029 two_stage_opamp_dummy_magic_19_0.V_err_p.n0 two_stage_opamp_dummy_magic_19_0.V_err_p.t1 15.7605
R7030 two_stage_opamp_dummy_magic_19_0.V_err_p.n0 two_stage_opamp_dummy_magic_19_0.V_err_p.t0 15.7605
R7031 two_stage_opamp_dummy_magic_19_0.V_err_p.n1 two_stage_opamp_dummy_magic_19_0.V_err_p.t3 15.7605
R7032 two_stage_opamp_dummy_magic_19_0.V_err_p.t2 two_stage_opamp_dummy_magic_19_0.V_err_p.n1 15.7605
R7033 two_stage_opamp_dummy_magic_19_0.V_p_mir.n2 two_stage_opamp_dummy_magic_19_0.V_p_mir.n0 60.064
R7034 two_stage_opamp_dummy_magic_19_0.V_p_mir.n2 two_stage_opamp_dummy_magic_19_0.V_p_mir.n1 42.8213
R7035 two_stage_opamp_dummy_magic_19_0.V_p_mir.n3 two_stage_opamp_dummy_magic_19_0.V_p_mir.n2 33.2588
R7036 two_stage_opamp_dummy_magic_19_0.V_p_mir.n0 two_stage_opamp_dummy_magic_19_0.V_p_mir.t5 16.0005
R7037 two_stage_opamp_dummy_magic_19_0.V_p_mir.n0 two_stage_opamp_dummy_magic_19_0.V_p_mir.t4 16.0005
R7038 two_stage_opamp_dummy_magic_19_0.V_p_mir.n1 two_stage_opamp_dummy_magic_19_0.V_p_mir.t0 9.6005
R7039 two_stage_opamp_dummy_magic_19_0.V_p_mir.n1 two_stage_opamp_dummy_magic_19_0.V_p_mir.t3 9.6005
R7040 two_stage_opamp_dummy_magic_19_0.V_p_mir.n3 two_stage_opamp_dummy_magic_19_0.V_p_mir.t2 9.6005
R7041 two_stage_opamp_dummy_magic_19_0.V_p_mir.t1 two_stage_opamp_dummy_magic_19_0.V_p_mir.n3 9.6005
R7042 bgr_9_0.START_UP_NFET1 bgr_9_0.START_UP_NFET1.t0 147.275
R7043 a_12530_23988.t0 a_12530_23988.t1 178.133
R7044 two_stage_opamp_dummy_magic_19_0.V_tot.n2 two_stage_opamp_dummy_magic_19_0.V_tot.t5 648.384
R7045 two_stage_opamp_dummy_magic_19_0.V_tot.n1 two_stage_opamp_dummy_magic_19_0.V_tot.t4 648.384
R7046 two_stage_opamp_dummy_magic_19_0.V_tot.t0 two_stage_opamp_dummy_magic_19_0.V_tot.n3 116.546
R7047 two_stage_opamp_dummy_magic_19_0.V_tot.n0 two_stage_opamp_dummy_magic_19_0.V_tot.t3 116.546
R7048 two_stage_opamp_dummy_magic_19_0.V_tot.n3 two_stage_opamp_dummy_magic_19_0.V_tot.t2 107.328
R7049 two_stage_opamp_dummy_magic_19_0.V_tot.n0 two_stage_opamp_dummy_magic_19_0.V_tot.t1 107.328
R7050 two_stage_opamp_dummy_magic_19_0.V_tot.n3 two_stage_opamp_dummy_magic_19_0.V_tot.n2 35.3494
R7051 two_stage_opamp_dummy_magic_19_0.V_tot.n1 two_stage_opamp_dummy_magic_19_0.V_tot.n0 35.3181
R7052 two_stage_opamp_dummy_magic_19_0.V_tot.n2 two_stage_opamp_dummy_magic_19_0.V_tot.n1 1.59425
R7053 a_7580_22380.t0 a_7580_22380.t1 178.133
R7054 a_14330_5524.t0 a_14330_5524.t1 262.248
R7055 a_6810_23838.t0 a_6810_23838.t1 178.133
R7056 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 195.608
R7057 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 83.5719
R7058 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 83.5719
R7059 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 83.5719
R7060 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 83.5719
R7061 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 83.5719
R7062 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 83.5719
R7063 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 83.5719
R7064 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 83.5719
R7065 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 83.5719
R7066 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 83.5719
R7067 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 83.5719
R7068 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 83.5719
R7069 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 83.5719
R7070 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 83.5719
R7071 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 83.5719
R7072 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 83.5719
R7073 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 83.5719
R7074 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 83.5719
R7075 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 83.5719
R7076 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 83.5719
R7077 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R7078 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 83.5719
R7079 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 73.8495
R7080 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 73.8495
R7081 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 73.3165
R7082 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 73.3165
R7083 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 73.3165
R7084 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 73.3165
R7085 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 73.3165
R7086 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 73.3165
R7087 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 73.19
R7088 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 73.19
R7089 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 73.19
R7090 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 73.19
R7091 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 73.19
R7092 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 73.19
R7093 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 65.0299
R7094 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 65.0299
R7095 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 26.074
R7096 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 26.074
R7097 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 26.074
R7098 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 26.074
R7099 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 26.074
R7100 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 26.074
R7101 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 26.074
R7102 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 26.074
R7103 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 25.7843
R7104 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 25.7843
R7105 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 25.7843
R7106 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 25.7843
R7107 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 25.7843
R7108 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 25.7843
R7109 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R7110 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R7111 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R7112 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R7113 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R7114 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R7115 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R7116 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 9.3005
R7117 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R7118 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R7119 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R7120 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R7121 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 9.3005
R7122 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 9.3005
R7123 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R7124 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R7125 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R7126 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R7127 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R7128 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R7129 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R7130 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R7131 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R7132 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R7133 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R7134 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 9.3005
R7135 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 9.3005
R7136 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 9.3005
R7137 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R7138 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R7139 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R7140 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 9.3005
R7141 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R7142 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R7143 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R7144 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 9.3005
R7145 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R7146 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R7147 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R7148 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R7149 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R7150 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R7151 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R7152 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R7153 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R7154 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R7155 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R7156 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R7157 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 9.3005
R7158 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 9.3005
R7159 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R7160 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R7161 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R7162 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R7163 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 4.64654
R7164 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 4.64654
R7165 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 4.64654
R7166 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 4.64654
R7167 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 4.64654
R7168 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 4.64654
R7169 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 4.64654
R7170 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 4.64654
R7171 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 4.64654
R7172 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 2.36206
R7173 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 2.36206
R7174 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 2.36206
R7175 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 2.36206
R7176 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 2.19742
R7177 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 2.19742
R7178 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 2.19742
R7179 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 2.19742
R7180 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 1.56363
R7181 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.56363
R7182 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 1.5505
R7183 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R7184 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 1.5505
R7185 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 1.5505
R7186 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 1.5505
R7187 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 1.5505
R7188 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 1.5505
R7189 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 1.5505
R7190 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 1.5505
R7191 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 1.5505
R7192 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 1.5505
R7193 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 1.5505
R7194 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 1.5505
R7195 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 1.5505
R7196 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 1.5505
R7197 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 1.5505
R7198 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 1.5505
R7199 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 1.5505
R7200 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.25468
R7201 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 1.25468
R7202 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.25468
R7203 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.25468
R7204 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 1.25468
R7205 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 1.25468
R7206 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 1.19225
R7207 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 1.19225
R7208 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 1.19225
R7209 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 1.19225
R7210 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 1.19225
R7211 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.19225
R7212 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 1.07024
R7213 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 1.07024
R7214 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 1.07024
R7215 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 1.07024
R7216 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 1.07024
R7217 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.07024
R7218 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.0237
R7219 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 1.0237
R7220 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.0237
R7221 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.0237
R7222 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 1.0237
R7223 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 1.0237
R7224 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.885803
R7225 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 0.885803
R7226 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 0.885803
R7227 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 0.885803
R7228 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.885803
R7229 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.885803
R7230 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 0.885803
R7231 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.885803
R7232 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 0.812055
R7233 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 0.812055
R7234 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.77514
R7235 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.77514
R7236 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 0.77514
R7237 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.77514
R7238 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.77514
R7239 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 0.77514
R7240 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 0.77514
R7241 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 0.77514
R7242 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.756696
R7243 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R7244 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.756696
R7245 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 0.756696
R7246 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R7247 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.756696
R7248 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R7249 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.756696
R7250 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 0.711459
R7251 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.711459
R7252 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.647417
R7253 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 0.647417
R7254 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.590702
R7255 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 0.590702
R7256 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.590702
R7257 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 0.590702
R7258 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.590702
R7259 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 0.590702
R7260 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.576566
R7261 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.576566
R7262 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 0.530034
R7263 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 0.530034
R7264 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 0.290206
R7265 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 0.290206
R7266 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 0.290206
R7267 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 0.290206
R7268 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 0.290206
R7269 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 0.290206
R7270 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 0.290206
R7271 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 0.290206
R7272 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R7273 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R7274 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R7275 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.203382
R7276 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R7277 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 0.203382
R7278 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 0.154071
R7279 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 0.154071
R7280 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 0.154071
R7281 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 0.154071
R7282 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 0.137464
R7283 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 0.137464
R7284 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 0.134964
R7285 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 0.134964
R7286 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R7287 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 0.0183571
R7288 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R7289 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R7290 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 0.0183571
R7291 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R7292 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R7293 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 0.0183571
R7294 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0183571
R7295 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R7296 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R7297 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R7298 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R7299 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 0.0183571
R7300 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R7301 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R7302 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 0.0183571
R7303 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0183571
R7304 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0106786
R7305 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0106786
R7306 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.0106786
R7307 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 0.00992001
R7308 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 0.00992001
R7309 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R7310 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 0.00992001
R7311 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R7312 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R7313 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R7314 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 0.00992001
R7315 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 0.00992001
R7316 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 0.00992001
R7317 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R7318 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 0.00992001
R7319 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R7320 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R7321 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R7322 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R7323 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 0.00992001
R7324 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R7325 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.00817857
R7326 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00817857
R7327 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 0.00817857
R7328 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 0.00817857
R7329 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.00817857
R7330 a_12410_22380.t0 a_12410_22380.t1 178.133
R7331 a_13060_22630.t0 a_13060_22630.t1 178.133
R7332 a_5420_5524.t0 a_5420_5524.t1 262.248
R7333 a_14450_5524.t0 a_14450_5524.t1 169.905
R7334 two_stage_opamp_dummy_magic_19_0.Vb2_2.n2 two_stage_opamp_dummy_magic_19_0.Vb2_2.t3 661.375
R7335 two_stage_opamp_dummy_magic_19_0.Vb2_2.n4 two_stage_opamp_dummy_magic_19_0.Vb2_2.t6 661.375
R7336 two_stage_opamp_dummy_magic_19_0.Vb2_2.t4 two_stage_opamp_dummy_magic_19_0.Vb2_2.n0 213.131
R7337 two_stage_opamp_dummy_magic_19_0.Vb2_2.n3 two_stage_opamp_dummy_magic_19_0.Vb2_2.t7 213.131
R7338 two_stage_opamp_dummy_magic_19_0.Vb2_2.n2 two_stage_opamp_dummy_magic_19_0.Vb2_2.n1 162.132
R7339 two_stage_opamp_dummy_magic_19_0.Vb2_2.t0 two_stage_opamp_dummy_magic_19_0.Vb2_2.t4 146.155
R7340 two_stage_opamp_dummy_magic_19_0.Vb2_2.t7 two_stage_opamp_dummy_magic_19_0.Vb2_2.t0 146.155
R7341 two_stage_opamp_dummy_magic_19_0.Vb2_2.t5 two_stage_opamp_dummy_magic_19_0.Vb2_2.n0 76.2576
R7342 two_stage_opamp_dummy_magic_19_0.Vb2_2.n3 two_stage_opamp_dummy_magic_19_0.Vb2_2.t8 76.2576
R7343 two_stage_opamp_dummy_magic_19_0.Vb2_2.n6 two_stage_opamp_dummy_magic_19_0.Vb2_2.n5 71.388
R7344 two_stage_opamp_dummy_magic_19_0.Vb2_2.n1 two_stage_opamp_dummy_magic_19_0.Vb2_2.t9 21.8894
R7345 two_stage_opamp_dummy_magic_19_0.Vb2_2.n1 two_stage_opamp_dummy_magic_19_0.Vb2_2.t2 21.8894
R7346 two_stage_opamp_dummy_magic_19_0.Vb2_2.t5 two_stage_opamp_dummy_magic_19_0.Vb2_2.n6 11.2576
R7347 two_stage_opamp_dummy_magic_19_0.Vb2_2.n6 two_stage_opamp_dummy_magic_19_0.Vb2_2.t1 11.2576
R7348 two_stage_opamp_dummy_magic_19_0.Vb2_2.n5 two_stage_opamp_dummy_magic_19_0.Vb2_2.n4 5.1255
R7349 two_stage_opamp_dummy_magic_19_0.Vb2_2.n5 two_stage_opamp_dummy_magic_19_0.Vb2_2.n2 4.7505
R7350 two_stage_opamp_dummy_magic_19_0.Vb2_2.n4 two_stage_opamp_dummy_magic_19_0.Vb2_2.n3 1.888
R7351 two_stage_opamp_dummy_magic_19_0.Vb2_2.n2 two_stage_opamp_dummy_magic_19_0.Vb2_2.n0 1.888
R7352 a_5540_5524.t0 a_5540_5524.t1 169.905
R7353 a_13180_23838.t0 a_13180_23838.t1 178.133
C0 bgr_9_0.START_UP two_stage_opamp_dummy_magic_19_0.V_err_amp_ref 1.36583f
C1 bgr_9_0.V_TOP bgr_9_0.1st_Vout_1 2.48388f
C2 bgr_9_0.NFET_GATE_10uA bgr_9_0.START_UP_NFET1 0.351171f
C3 bgr_9_0.NFET_GATE_10uA bgr_9_0.1st_Vout_1 0.03875f
C4 bgr_9_0.START_UP_NFET1 bgr_9_0.START_UP 0.145663f
C5 two_stage_opamp_dummy_magic_19_0.V_err_gate bgr_9_0.1st_Vout_1 0.041119f
C6 bgr_9_0.START_UP bgr_9_0.1st_Vout_1 0.044074f
C7 two_stage_opamp_dummy_magic_19_0.V_err_mir_p VDDA 1.13437f
C8 bgr_9_0.V_p_1 bgr_9_0.1st_Vout_1 0.311617f
C9 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref VDDA 2.82258f
C10 m1_4880_3600# m2_4880_3600# 0.016063f
C11 two_stage_opamp_dummy_magic_19_0.cap_res_X VOUT+ 0.037134f
C12 two_stage_opamp_dummy_magic_19_0.V_err_gate two_stage_opamp_dummy_magic_19_0.cap_res_X 0.33348f
C13 bgr_9_0.V_TOP bgr_9_0.PFET_GATE_10uA 0.212258f
C14 bgr_9_0.START_UP_NFET1 VDDA 0.151315f
C15 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter VDDA 0.046803f
C16 two_stage_opamp_dummy_magic_19_0.cap_res_X VOUT- 51.024498f
C17 two_stage_opamp_dummy_magic_19_0.VD4 VOUT+ 0.040325f
C18 bgr_9_0.NFET_GATE_10uA bgr_9_0.PFET_GATE_10uA 0.011067f
C19 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref two_stage_opamp_dummy_magic_19_0.V_err_mir_p 0.059807f
C20 bgr_9_0.1st_Vout_1 VDDA 0.920268f
C21 two_stage_opamp_dummy_magic_19_0.V_err_gate bgr_9_0.PFET_GATE_10uA 0.091127f
C22 bgr_9_0.V_TOP bgr_9_0.NFET_GATE_10uA 0.049214f
C23 two_stage_opamp_dummy_magic_19_0.VD2 VIN+ 0.88084f
C24 bgr_9_0.V_TOP two_stage_opamp_dummy_magic_19_0.V_err_gate 0.08195f
C25 two_stage_opamp_dummy_magic_19_0.cap_res_X VDDA 0.445525f
C26 bgr_9_0.V_TOP bgr_9_0.START_UP 0.792764f
C27 two_stage_opamp_dummy_magic_19_0.VD1 VIN- 0.880738f
C28 two_stage_opamp_dummy_magic_19_0.VD1 VDDA 0.012732f
C29 bgr_9_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_19_0.V_err_gate 3.51904f
C30 two_stage_opamp_dummy_magic_19_0.VD2 VDDA 0.012624f
C31 bgr_9_0.NFET_GATE_10uA bgr_9_0.START_UP 1.64125f
C32 two_stage_opamp_dummy_magic_19_0.VD4 VDDA 7.98282f
C33 bgr_9_0.PFET_GATE_10uA VDDA 8.3027f
C34 VOUT+ VOUT- 0.397591f
C35 two_stage_opamp_dummy_magic_19_0.V_err_gate VOUT- 0.038042f
C36 bgr_9_0.START_UP bgr_9_0.V_p_1 0.038571f
C37 bgr_9_0.V_TOP VDDA 13.5266f
C38 two_stage_opamp_dummy_magic_19_0.VD4 two_stage_opamp_dummy_magic_19_0.V_err_mir_p 0.019941f
C39 two_stage_opamp_dummy_magic_19_0.VD4 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref 0.044858f
C40 bgr_9_0.NFET_GATE_10uA VDDA 0.214466f
C41 bgr_9_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_19_0.V_err_amp_ref 1.67029f
C42 VDDA VOUT+ 12.271099f
C43 two_stage_opamp_dummy_magic_19_0.V_err_gate VDDA 2.70518f
C44 bgr_9_0.START_UP VDDA 1.08377f
C45 bgr_9_0.START_UP_NFET1 bgr_9_0.PFET_GATE_10uA 0.0108f
C46 bgr_9_0.V_TOP two_stage_opamp_dummy_magic_19_0.V_err_amp_ref 0.583702f
C47 VDDA VOUT- 12.274099f
C48 bgr_9_0.V_p_1 VDDA 0.417418f
C49 two_stage_opamp_dummy_magic_19_0.V_err_gate two_stage_opamp_dummy_magic_19_0.V_err_mir_p 0.885274f
C50 VIN+ VIN- 0.120537f
C51 bgr_9_0.V_TOP bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.055802f
C52 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref VOUT+ 0.038959f
C53 two_stage_opamp_dummy_magic_19_0.V_err_gate two_stage_opamp_dummy_magic_19_0.V_err_amp_ref 0.841328f
C54 VIN- GNDA 2.45458f
C55 VIN+ GNDA 2.45147f
C56 VOUT- GNDA 17.659557f
C57 VOUT+ GNDA 17.69017f
C58 VDDA GNDA 0.123135p
C59 m2_4880_3600# GNDA 0.052359f $ **FLOATING
C60 m1_4880_3600# GNDA 0.059483f $ **FLOATING
C61 two_stage_opamp_dummy_magic_19_0.cap_res_X GNDA 32.93443f
C62 two_stage_opamp_dummy_magic_19_0.VD1 GNDA 1.314036f
C63 two_stage_opamp_dummy_magic_19_0.VD2 GNDA 1.668806f
C64 two_stage_opamp_dummy_magic_19_0.V_err_mir_p GNDA 0.060575f
C65 bgr_9_0.1st_Vout_1 GNDA 7.806533f
C66 bgr_9_0.V_p_1 GNDA 0.763998f
C67 bgr_9_0.START_UP GNDA 5.883708f
C68 bgr_9_0.START_UP_NFET1 GNDA 4.30721f
C69 two_stage_opamp_dummy_magic_19_0.V_err_gate GNDA 9.14163f
C70 bgr_9_0.NFET_GATE_10uA GNDA 7.21764f
C71 bgr_9_0.V_TOP GNDA 9.886665f
C72 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA 17.900902f
C73 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref GNDA 7.10432f
C74 bgr_9_0.PFET_GATE_10uA GNDA 6.290109f
C75 two_stage_opamp_dummy_magic_19_0.VD4 GNDA 4.745979f
C76 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t14 GNDA 0.026064f
C77 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t12 GNDA 0.026064f
C78 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n0 GNDA 0.093973f
C79 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t13 GNDA 0.026064f
C80 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t11 GNDA 0.026064f
C81 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n1 GNDA 0.078548f
C82 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n2 GNDA 1.53645f
C83 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t0 GNDA 0.319725f
C84 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t5 GNDA 0.078193f
C85 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t9 GNDA 0.078193f
C86 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n3 GNDA 0.259679f
C87 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t1 GNDA 0.078193f
C88 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t10 GNDA 0.078193f
C89 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n4 GNDA 0.25098f
C90 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n5 GNDA 0.938516f
C91 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t4 GNDA 0.078193f
C92 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t8 GNDA 0.078193f
C93 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n6 GNDA 0.25098f
C94 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n7 GNDA 0.482729f
C95 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t3 GNDA 0.078193f
C96 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t7 GNDA 0.078193f
C97 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n8 GNDA 0.25098f
C98 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n9 GNDA 0.482729f
C99 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t2 GNDA 0.078193f
C100 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.t6 GNDA 0.078193f
C101 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n10 GNDA 0.25098f
C102 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n11 GNDA 0.572912f
C103 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n12 GNDA 1.84331f
C104 two_stage_opamp_dummy_magic_19_0.V_CMFB_S4.n13 GNDA 2.28828f
C105 bgr_9_0.V_CMFB_S4 GNDA 0.013032f
C106 bgr_9_0.START_UP.t0 GNDA 1.11411f
C107 bgr_9_0.START_UP.t1 GNDA 0.031262f
C108 bgr_9_0.START_UP.n0 GNDA 0.717543f
C109 bgr_9_0.START_UP.t2 GNDA 0.027731f
C110 bgr_9_0.START_UP.t4 GNDA 0.027731f
C111 bgr_9_0.START_UP.n1 GNDA 0.104651f
C112 bgr_9_0.START_UP.t3 GNDA 0.027731f
C113 bgr_9_0.START_UP.t5 GNDA 0.027731f
C114 bgr_9_0.START_UP.n2 GNDA 0.096735f
C115 bgr_9_0.START_UP.n3 GNDA 0.471093f
C116 bgr_9_0.START_UP.t7 GNDA 0.010421f
C117 bgr_9_0.START_UP.t6 GNDA 0.010421f
C118 bgr_9_0.START_UP.n4 GNDA 0.029418f
C119 bgr_9_0.START_UP.n5 GNDA 0.270117f
C120 two_stage_opamp_dummy_magic_19_0.VD4.t32 GNDA 0.058707f
C121 two_stage_opamp_dummy_magic_19_0.VD4.t37 GNDA 0.058707f
C122 two_stage_opamp_dummy_magic_19_0.VD4.n0 GNDA 0.150855f
C123 two_stage_opamp_dummy_magic_19_0.VD4.t31 GNDA 0.058707f
C124 two_stage_opamp_dummy_magic_19_0.VD4.t29 GNDA 0.058707f
C125 two_stage_opamp_dummy_magic_19_0.VD4.n1 GNDA 0.147477f
C126 two_stage_opamp_dummy_magic_19_0.VD4.n2 GNDA 0.788587f
C127 two_stage_opamp_dummy_magic_19_0.VD4.t26 GNDA 0.058707f
C128 two_stage_opamp_dummy_magic_19_0.VD4.t28 GNDA 0.058707f
C129 two_stage_opamp_dummy_magic_19_0.VD4.n3 GNDA 0.147477f
C130 two_stage_opamp_dummy_magic_19_0.VD4.n4 GNDA 0.402692f
C131 two_stage_opamp_dummy_magic_19_0.VD4.t34 GNDA 0.058707f
C132 two_stage_opamp_dummy_magic_19_0.VD4.t35 GNDA 0.058707f
C133 two_stage_opamp_dummy_magic_19_0.VD4.n5 GNDA 0.147477f
C134 two_stage_opamp_dummy_magic_19_0.VD4.n6 GNDA 0.402692f
C135 two_stage_opamp_dummy_magic_19_0.VD4.t30 GNDA 0.058707f
C136 two_stage_opamp_dummy_magic_19_0.VD4.t33 GNDA 0.058707f
C137 two_stage_opamp_dummy_magic_19_0.VD4.n7 GNDA 0.147477f
C138 two_stage_opamp_dummy_magic_19_0.VD4.n8 GNDA 0.402692f
C139 two_stage_opamp_dummy_magic_19_0.VD4.t36 GNDA 0.058707f
C140 two_stage_opamp_dummy_magic_19_0.VD4.t27 GNDA 0.058707f
C141 two_stage_opamp_dummy_magic_19_0.VD4.n9 GNDA 0.147477f
C142 two_stage_opamp_dummy_magic_19_0.VD4.n10 GNDA 0.495479f
C143 two_stage_opamp_dummy_magic_19_0.VD4.t15 GNDA 0.058707f
C144 two_stage_opamp_dummy_magic_19_0.VD4.t19 GNDA 0.058707f
C145 two_stage_opamp_dummy_magic_19_0.VD4.n11 GNDA 0.147477f
C146 two_stage_opamp_dummy_magic_19_0.VD4.n12 GNDA 0.402692f
C147 two_stage_opamp_dummy_magic_19_0.VD4.t22 GNDA 0.208829f
C148 two_stage_opamp_dummy_magic_19_0.VD4.t23 GNDA 0.102932f
C149 two_stage_opamp_dummy_magic_19_0.VD4.t5 GNDA 0.058707f
C150 two_stage_opamp_dummy_magic_19_0.VD4.t9 GNDA 0.058707f
C151 two_stage_opamp_dummy_magic_19_0.VD4.n13 GNDA 0.147477f
C152 two_stage_opamp_dummy_magic_19_0.VD4.n14 GNDA 0.402692f
C153 two_stage_opamp_dummy_magic_19_0.VD4.t1 GNDA 0.058707f
C154 two_stage_opamp_dummy_magic_19_0.VD4.t3 GNDA 0.058707f
C155 two_stage_opamp_dummy_magic_19_0.VD4.n15 GNDA 0.147477f
C156 two_stage_opamp_dummy_magic_19_0.VD4.n16 GNDA 0.402692f
C157 two_stage_opamp_dummy_magic_19_0.VD4.t13 GNDA 0.058707f
C158 two_stage_opamp_dummy_magic_19_0.VD4.t17 GNDA 0.058707f
C159 two_stage_opamp_dummy_magic_19_0.VD4.n17 GNDA 0.147477f
C160 two_stage_opamp_dummy_magic_19_0.VD4.n18 GNDA 0.402692f
C161 two_stage_opamp_dummy_magic_19_0.VD4.t11 GNDA 0.058707f
C162 two_stage_opamp_dummy_magic_19_0.VD4.t7 GNDA 0.058707f
C163 two_stage_opamp_dummy_magic_19_0.VD4.n19 GNDA 0.147477f
C164 two_stage_opamp_dummy_magic_19_0.VD4.n20 GNDA 0.458507f
C165 two_stage_opamp_dummy_magic_19_0.VD4.n21 GNDA 0.158682f
C166 two_stage_opamp_dummy_magic_19_0.VD4.t25 GNDA 0.208829f
C167 two_stage_opamp_dummy_magic_19_0.VD4.n22 GNDA 0.373261f
C168 two_stage_opamp_dummy_magic_19_0.VD4.t24 GNDA 0.497708f
C169 two_stage_opamp_dummy_magic_19_0.VD4.t10 GNDA 0.392499f
C170 two_stage_opamp_dummy_magic_19_0.VD4.t6 GNDA 0.392499f
C171 two_stage_opamp_dummy_magic_19_0.VD4.t12 GNDA 0.392499f
C172 two_stage_opamp_dummy_magic_19_0.VD4.t16 GNDA 0.392499f
C173 two_stage_opamp_dummy_magic_19_0.VD4.t0 GNDA 0.392499f
C174 two_stage_opamp_dummy_magic_19_0.VD4.t2 GNDA 0.392499f
C175 two_stage_opamp_dummy_magic_19_0.VD4.t4 GNDA 0.392499f
C176 two_stage_opamp_dummy_magic_19_0.VD4.t8 GNDA 0.392499f
C177 two_stage_opamp_dummy_magic_19_0.VD4.t14 GNDA 0.392499f
C178 two_stage_opamp_dummy_magic_19_0.VD4.t18 GNDA 0.392499f
C179 two_stage_opamp_dummy_magic_19_0.VD4.t21 GNDA 0.497708f
C180 two_stage_opamp_dummy_magic_19_0.VD4.n23 GNDA 0.373261f
C181 two_stage_opamp_dummy_magic_19_0.VD4.t20 GNDA 0.102932f
C182 two_stage_opamp_dummy_magic_19_0.VD4.n24 GNDA 0.156154f
C183 two_stage_opamp_dummy_magic_19_0.VD4.n25 GNDA 0.138141f
C184 two_stage_opamp_dummy_magic_19_0.VD4.n26 GNDA 0.17127f
C185 bgr_9_0.Vin-.n0 GNDA 0.070741f
C186 bgr_9_0.Vin-.n1 GNDA 0.320657f
C187 bgr_9_0.Vin-.t6 GNDA 0.027487f
C188 bgr_9_0.Vin-.t4 GNDA 0.027487f
C189 bgr_9_0.Vin-.n2 GNDA 0.099751f
C190 bgr_9_0.Vin-.t3 GNDA 0.027487f
C191 bgr_9_0.Vin-.t5 GNDA 0.027487f
C192 bgr_9_0.Vin-.n3 GNDA 0.09553f
C193 bgr_9_0.Vin-.n4 GNDA 0.383788f
C194 bgr_9_0.Vin-.n5 GNDA 0.028037f
C195 bgr_9_0.Vin-.n6 GNDA 0.371517f
C196 bgr_9_0.Vin-.t12 GNDA 0.022665f
C197 bgr_9_0.Vin-.n7 GNDA 0.026583f
C198 bgr_9_0.Vin-.n8 GNDA 0.021761f
C199 bgr_9_0.Vin-.n9 GNDA 0.021761f
C200 bgr_9_0.Vin-.n10 GNDA 0.037011f
C201 bgr_9_0.Vin-.n11 GNDA 0.505034f
C202 bgr_9_0.Vin-.t1 GNDA 0.120899f
C203 bgr_9_0.Vin-.n12 GNDA 0.678321f
C204 bgr_9_0.Vin-.n13 GNDA 1.08827f
C205 bgr_9_0.Vin-.n14 GNDA 0.478045f
C206 bgr_9_0.Vin-.t2 GNDA 0.265362f
C207 bgr_9_0.Vin-.n15 GNDA 0.070872f
C208 bgr_9_0.Vin-.n16 GNDA 0.121299f
C209 bgr_9_0.Vin-.n17 GNDA 0.071536f
C210 bgr_9_0.Vin-.n18 GNDA 0.587286f
C211 bgr_9_0.Vin-.n19 GNDA 0.363325f
C212 bgr_9_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter GNDA 0.087772f
C213 bgr_9_0.V_mir2.t7 GNDA 0.019293f
C214 bgr_9_0.V_mir2.n0 GNDA 0.025223f
C215 bgr_9_0.V_mir2.t14 GNDA 0.041163f
C216 bgr_9_0.V_mir2.n1 GNDA 0.027381f
C217 bgr_9_0.V_mir2.n2 GNDA 0.451535f
C218 bgr_9_0.V_mir2.n3 GNDA 0.146338f
C219 bgr_9_0.V_mir2.t4 GNDA 0.023151f
C220 bgr_9_0.V_mir2.t17 GNDA 0.023151f
C221 bgr_9_0.V_mir2.t20 GNDA 0.037369f
C222 bgr_9_0.V_mir2.n4 GNDA 0.041731f
C223 bgr_9_0.V_mir2.n5 GNDA 0.028507f
C224 bgr_9_0.V_mir2.t0 GNDA 0.02939f
C225 bgr_9_0.V_mir2.n6 GNDA 0.044354f
C226 bgr_9_0.V_mir2.t5 GNDA 0.019293f
C227 bgr_9_0.V_mir2.t1 GNDA 0.019293f
C228 bgr_9_0.V_mir2.n7 GNDA 0.044322f
C229 bgr_9_0.V_mir2.n8 GNDA 0.109787f
C230 bgr_9_0.V_mir2.t2 GNDA 0.023151f
C231 bgr_9_0.V_mir2.t18 GNDA 0.023151f
C232 bgr_9_0.V_mir2.t22 GNDA 0.037369f
C233 bgr_9_0.V_mir2.n9 GNDA 0.041731f
C234 bgr_9_0.V_mir2.n10 GNDA 0.028507f
C235 bgr_9_0.V_mir2.t8 GNDA 0.02939f
C236 bgr_9_0.V_mir2.n11 GNDA 0.044354f
C237 bgr_9_0.V_mir2.t3 GNDA 0.019293f
C238 bgr_9_0.V_mir2.t9 GNDA 0.019293f
C239 bgr_9_0.V_mir2.n12 GNDA 0.044322f
C240 bgr_9_0.V_mir2.n13 GNDA 0.110886f
C241 bgr_9_0.V_mir2.n14 GNDA 0.381359f
C242 bgr_9_0.V_mir2.n15 GNDA 0.051125f
C243 bgr_9_0.V_mir2.t6 GNDA 0.023151f
C244 bgr_9_0.V_mir2.t19 GNDA 0.023151f
C245 bgr_9_0.V_mir2.t21 GNDA 0.037369f
C246 bgr_9_0.V_mir2.n16 GNDA 0.041731f
C247 bgr_9_0.V_mir2.n17 GNDA 0.028507f
C248 bgr_9_0.V_mir2.t10 GNDA 0.02939f
C249 bgr_9_0.V_mir2.n18 GNDA 0.044354f
C250 bgr_9_0.V_mir2.n19 GNDA 0.084938f
C251 bgr_9_0.V_mir2.n20 GNDA 0.044322f
C252 bgr_9_0.V_mir2.t11 GNDA 0.019293f
C253 bgr_9_0.cap_res1.t12 GNDA 0.332137f
C254 bgr_9_0.cap_res1.t19 GNDA 0.349634f
C255 bgr_9_0.cap_res1.t16 GNDA 0.350901f
C256 bgr_9_0.cap_res1.t5 GNDA 0.332137f
C257 bgr_9_0.cap_res1.t15 GNDA 0.349634f
C258 bgr_9_0.cap_res1.t9 GNDA 0.350901f
C259 bgr_9_0.cap_res1.t11 GNDA 0.332137f
C260 bgr_9_0.cap_res1.t18 GNDA 0.349634f
C261 bgr_9_0.cap_res1.t14 GNDA 0.350901f
C262 bgr_9_0.cap_res1.t4 GNDA 0.332137f
C263 bgr_9_0.cap_res1.t13 GNDA 0.349634f
C264 bgr_9_0.cap_res1.t7 GNDA 0.350901f
C265 bgr_9_0.cap_res1.t20 GNDA 0.332137f
C266 bgr_9_0.cap_res1.t6 GNDA 0.349634f
C267 bgr_9_0.cap_res1.t1 GNDA 0.350901f
C268 bgr_9_0.cap_res1.n0 GNDA 0.23436f
C269 bgr_9_0.cap_res1.t17 GNDA 0.186633f
C270 bgr_9_0.cap_res1.n1 GNDA 0.254286f
C271 bgr_9_0.cap_res1.t2 GNDA 0.186633f
C272 bgr_9_0.cap_res1.n2 GNDA 0.254286f
C273 bgr_9_0.cap_res1.t8 GNDA 0.186633f
C274 bgr_9_0.cap_res1.n3 GNDA 0.254286f
C275 bgr_9_0.cap_res1.t3 GNDA 0.186633f
C276 bgr_9_0.cap_res1.n4 GNDA 0.254286f
C277 bgr_9_0.cap_res1.t10 GNDA 0.355331f
C278 bgr_9_0.cap_res1.t0 GNDA 0.083274f
C279 bgr_9_0.PFET_GATE_10uA.t23 GNDA 0.020877f
C280 bgr_9_0.PFET_GATE_10uA.t17 GNDA 0.030909f
C281 bgr_9_0.PFET_GATE_10uA.n0 GNDA 0.066443f
C282 bgr_9_0.PFET_GATE_10uA.t24 GNDA 0.020877f
C283 bgr_9_0.PFET_GATE_10uA.t19 GNDA 0.030861f
C284 bgr_9_0.PFET_GATE_10uA.n1 GNDA 0.034006f
C285 bgr_9_0.PFET_GATE_10uA.t13 GNDA 0.020877f
C286 bgr_9_0.PFET_GATE_10uA.t20 GNDA 0.030861f
C287 bgr_9_0.PFET_GATE_10uA.n2 GNDA 0.034006f
C288 bgr_9_0.PFET_GATE_10uA.n3 GNDA 0.031726f
C289 bgr_9_0.PFET_GATE_10uA.n4 GNDA 0.656762f
C290 bgr_9_0.PFET_GATE_10uA.t16 GNDA 0.020877f
C291 bgr_9_0.PFET_GATE_10uA.t11 GNDA 0.030861f
C292 bgr_9_0.PFET_GATE_10uA.n5 GNDA 0.034006f
C293 bgr_9_0.PFET_GATE_10uA.t22 GNDA 0.020877f
C294 bgr_9_0.PFET_GATE_10uA.t12 GNDA 0.030861f
C295 bgr_9_0.PFET_GATE_10uA.n6 GNDA 0.034006f
C296 bgr_9_0.PFET_GATE_10uA.n7 GNDA 0.034115f
C297 bgr_9_0.PFET_GATE_10uA.t7 GNDA 0.311852f
C298 bgr_9_0.PFET_GATE_10uA.t0 GNDA 0.021412f
C299 bgr_9_0.PFET_GATE_10uA.t8 GNDA 0.021412f
C300 bgr_9_0.PFET_GATE_10uA.n8 GNDA 0.054804f
C301 bgr_9_0.PFET_GATE_10uA.t2 GNDA 0.021412f
C302 bgr_9_0.PFET_GATE_10uA.t4 GNDA 0.021412f
C303 bgr_9_0.PFET_GATE_10uA.n9 GNDA 0.053412f
C304 bgr_9_0.PFET_GATE_10uA.n10 GNDA 0.521294f
C305 bgr_9_0.PFET_GATE_10uA.t3 GNDA 0.021412f
C306 bgr_9_0.PFET_GATE_10uA.t5 GNDA 0.021412f
C307 bgr_9_0.PFET_GATE_10uA.n11 GNDA 0.053412f
C308 bgr_9_0.PFET_GATE_10uA.n12 GNDA 0.295602f
C309 bgr_9_0.PFET_GATE_10uA.n13 GNDA 0.604578f
C310 bgr_9_0.PFET_GATE_10uA.t9 GNDA 0.021412f
C311 bgr_9_0.PFET_GATE_10uA.t1 GNDA 0.021412f
C312 bgr_9_0.PFET_GATE_10uA.n14 GNDA 0.051768f
C313 bgr_9_0.PFET_GATE_10uA.n15 GNDA 0.275557f
C314 bgr_9_0.PFET_GATE_10uA.t6 GNDA 0.471424f
C315 bgr_9_0.PFET_GATE_10uA.t18 GNDA 0.062678f
C316 bgr_9_0.PFET_GATE_10uA.n16 GNDA 1.9454f
C317 bgr_9_0.PFET_GATE_10uA.n17 GNDA 0.775485f
C318 bgr_9_0.PFET_GATE_10uA.n18 GNDA 0.759978f
C319 bgr_9_0.PFET_GATE_10uA.t10 GNDA 0.044965f
C320 bgr_9_0.PFET_GATE_10uA.t21 GNDA 0.044965f
C321 bgr_9_0.PFET_GATE_10uA.t15 GNDA 0.0546f
C322 bgr_9_0.PFET_GATE_10uA.n19 GNDA 0.0546f
C323 bgr_9_0.PFET_GATE_10uA.n20 GNDA 0.031143f
C324 bgr_9_0.PFET_GATE_10uA.t14 GNDA 0.048358f
C325 bgr_9_0.PFET_GATE_10uA.n21 GNDA 0.053053f
C326 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t1 GNDA 0.116135f
C327 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t7 GNDA 0.293601f
C328 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t9 GNDA 0.348459f
C329 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n0 GNDA 0.179119f
C330 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t3 GNDA 0.293601f
C331 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t8 GNDA 0.348459f
C332 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n1 GNDA 0.179119f
C333 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n2 GNDA 0.026022f
C334 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n3 GNDA 0.615485f
C335 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t2 GNDA 0.293601f
C336 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t5 GNDA 0.348459f
C337 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n4 GNDA 0.179119f
C338 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t6 GNDA 0.293601f
C339 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t4 GNDA 0.348459f
C340 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n5 GNDA 0.179119f
C341 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n6 GNDA 0.026022f
C342 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.n7 GNDA 0.615484f
C343 two_stage_opamp_dummy_magic_19_0.V_b_2nd_stage.t0 GNDA 0.116135f
C344 two_stage_opamp_dummy_magic_19_0.VD1.t9 GNDA 0.044491f
C345 two_stage_opamp_dummy_magic_19_0.VD1.t4 GNDA 0.044491f
C346 two_stage_opamp_dummy_magic_19_0.VD1.n0 GNDA 0.098712f
C347 two_stage_opamp_dummy_magic_19_0.VD1.t11 GNDA 0.044491f
C348 two_stage_opamp_dummy_magic_19_0.VD1.t6 GNDA 0.044491f
C349 two_stage_opamp_dummy_magic_19_0.VD1.n1 GNDA 0.126567f
C350 two_stage_opamp_dummy_magic_19_0.VD1.t10 GNDA 0.044491f
C351 two_stage_opamp_dummy_magic_19_0.VD1.t5 GNDA 0.044491f
C352 two_stage_opamp_dummy_magic_19_0.VD1.n2 GNDA 0.122991f
C353 two_stage_opamp_dummy_magic_19_0.VD1.n3 GNDA 0.666968f
C354 two_stage_opamp_dummy_magic_19_0.VD1.t8 GNDA 0.044491f
C355 two_stage_opamp_dummy_magic_19_0.VD1.t13 GNDA 0.044491f
C356 two_stage_opamp_dummy_magic_19_0.VD1.n4 GNDA 0.126567f
C357 two_stage_opamp_dummy_magic_19_0.VD1.t7 GNDA 0.044491f
C358 two_stage_opamp_dummy_magic_19_0.VD1.t12 GNDA 0.044491f
C359 two_stage_opamp_dummy_magic_19_0.VD1.n5 GNDA 0.122991f
C360 two_stage_opamp_dummy_magic_19_0.VD1.n6 GNDA 0.666968f
C361 two_stage_opamp_dummy_magic_19_0.VD1.n7 GNDA 0.077119f
C362 two_stage_opamp_dummy_magic_19_0.VD1.n8 GNDA 0.329663f
C363 two_stage_opamp_dummy_magic_19_0.VD1.t19 GNDA 0.044491f
C364 two_stage_opamp_dummy_magic_19_0.VD1.t0 GNDA 0.044491f
C365 two_stage_opamp_dummy_magic_19_0.VD1.n9 GNDA 0.12611f
C366 two_stage_opamp_dummy_magic_19_0.VD1.t16 GNDA 0.044491f
C367 two_stage_opamp_dummy_magic_19_0.VD1.t21 GNDA 0.044491f
C368 two_stage_opamp_dummy_magic_19_0.VD1.n10 GNDA 0.122664f
C369 two_stage_opamp_dummy_magic_19_0.VD1.n11 GNDA 0.688514f
C370 two_stage_opamp_dummy_magic_19_0.VD1.t15 GNDA 0.044491f
C371 two_stage_opamp_dummy_magic_19_0.VD1.t2 GNDA 0.044491f
C372 two_stage_opamp_dummy_magic_19_0.VD1.n12 GNDA 0.122664f
C373 two_stage_opamp_dummy_magic_19_0.VD1.n13 GNDA 0.339751f
C374 two_stage_opamp_dummy_magic_19_0.VD1.t1 GNDA 0.044491f
C375 two_stage_opamp_dummy_magic_19_0.VD1.t20 GNDA 0.044491f
C376 two_stage_opamp_dummy_magic_19_0.VD1.n14 GNDA 0.12611f
C377 two_stage_opamp_dummy_magic_19_0.VD1.t14 GNDA 0.044491f
C378 two_stage_opamp_dummy_magic_19_0.VD1.t18 GNDA 0.044491f
C379 two_stage_opamp_dummy_magic_19_0.VD1.n15 GNDA 0.122664f
C380 two_stage_opamp_dummy_magic_19_0.VD1.n16 GNDA 0.688514f
C381 two_stage_opamp_dummy_magic_19_0.VD1.t17 GNDA 0.044491f
C382 two_stage_opamp_dummy_magic_19_0.VD1.t3 GNDA 0.044491f
C383 two_stage_opamp_dummy_magic_19_0.VD1.n17 GNDA 0.122664f
C384 two_stage_opamp_dummy_magic_19_0.VD1.n18 GNDA 0.339751f
C385 two_stage_opamp_dummy_magic_19_0.VD1.n19 GNDA 0.054339f
C386 two_stage_opamp_dummy_magic_19_0.Vb1.t0 GNDA 0.011823f
C387 two_stage_opamp_dummy_magic_19_0.Vb1.t11 GNDA 0.011823f
C388 two_stage_opamp_dummy_magic_19_0.Vb1.n0 GNDA 0.043357f
C389 two_stage_opamp_dummy_magic_19_0.Vb1.t18 GNDA 0.011789f
C390 two_stage_opamp_dummy_magic_19_0.Vb1.n1 GNDA 0.012818f
C391 two_stage_opamp_dummy_magic_19_0.Vb1.t12 GNDA 0.011789f
C392 two_stage_opamp_dummy_magic_19_0.Vb1.n3 GNDA 0.012818f
C393 two_stage_opamp_dummy_magic_19_0.Vb1.n9 GNDA 0.012267f
C394 two_stage_opamp_dummy_magic_19_0.Vb1.t26 GNDA 0.011789f
C395 two_stage_opamp_dummy_magic_19_0.Vb1.n10 GNDA 0.012818f
C396 two_stage_opamp_dummy_magic_19_0.Vb1.t20 GNDA 0.011789f
C397 two_stage_opamp_dummy_magic_19_0.Vb1.n16 GNDA 0.012818f
C398 two_stage_opamp_dummy_magic_19_0.Vb1.n19 GNDA 0.223636f
C399 two_stage_opamp_dummy_magic_19_0.Vb1.t15 GNDA 0.277108f
C400 two_stage_opamp_dummy_magic_19_0.Vb1.n20 GNDA 0.024723f
C401 two_stage_opamp_dummy_magic_19_0.Vb1.n21 GNDA 0.133851f
C402 two_stage_opamp_dummy_magic_19_0.Vb1.t3 GNDA 0.011789f
C403 two_stage_opamp_dummy_magic_19_0.Vb1.n22 GNDA 0.01212f
C404 two_stage_opamp_dummy_magic_19_0.Vb1.t5 GNDA 0.011789f
C405 two_stage_opamp_dummy_magic_19_0.Vb1.n23 GNDA 0.01212f
C406 two_stage_opamp_dummy_magic_19_0.Vb1.n25 GNDA 0.019691f
C407 two_stage_opamp_dummy_magic_19_0.Vb1.n26 GNDA 0.069619f
C408 two_stage_opamp_dummy_magic_19_0.Vb1.n27 GNDA 0.017735f
C409 two_stage_opamp_dummy_magic_19_0.Vb1.n28 GNDA 0.024723f
C410 two_stage_opamp_dummy_magic_19_0.Vb1.n29 GNDA 0.249517f
C411 two_stage_opamp_dummy_magic_19_0.Vb1.n30 GNDA 0.442758f
C412 bgr_9_0.VB1_CUR_BIAS GNDA 0.456948f
C413 two_stage_opamp_dummy_magic_19_0.V_err_gate.t2 GNDA 0.027098f
C414 two_stage_opamp_dummy_magic_19_0.V_err_gate.t3 GNDA 0.027098f
C415 two_stage_opamp_dummy_magic_19_0.V_err_gate.n0 GNDA 0.401617f
C416 two_stage_opamp_dummy_magic_19_0.V_err_gate.t1 GNDA 0.067744f
C417 two_stage_opamp_dummy_magic_19_0.V_err_gate.t5 GNDA 0.067744f
C418 two_stage_opamp_dummy_magic_19_0.V_err_gate.n1 GNDA 0.16347f
C419 two_stage_opamp_dummy_magic_19_0.V_err_gate.t8 GNDA 0.075647f
C420 two_stage_opamp_dummy_magic_19_0.V_err_gate.t6 GNDA 0.075647f
C421 two_stage_opamp_dummy_magic_19_0.V_err_gate.n2 GNDA 0.113628f
C422 two_stage_opamp_dummy_magic_19_0.V_err_gate.n3 GNDA 0.659577f
C423 two_stage_opamp_dummy_magic_19_0.V_err_gate.t4 GNDA 0.067744f
C424 two_stage_opamp_dummy_magic_19_0.V_err_gate.t0 GNDA 0.067744f
C425 two_stage_opamp_dummy_magic_19_0.V_err_gate.n4 GNDA 0.160398f
C426 two_stage_opamp_dummy_magic_19_0.V_err_gate.n5 GNDA 0.557689f
C427 two_stage_opamp_dummy_magic_19_0.V_err_gate.t7 GNDA 0.075647f
C428 two_stage_opamp_dummy_magic_19_0.V_err_gate.t9 GNDA 0.075647f
C429 two_stage_opamp_dummy_magic_19_0.V_err_gate.n6 GNDA 0.113628f
C430 two_stage_opamp_dummy_magic_19_0.VD2.n0 GNDA 0.339511f
C431 two_stage_opamp_dummy_magic_19_0.VD2.n1 GNDA 0.393812f
C432 two_stage_opamp_dummy_magic_19_0.VD2.t16 GNDA 0.04446f
C433 two_stage_opamp_dummy_magic_19_0.VD2.t12 GNDA 0.04446f
C434 two_stage_opamp_dummy_magic_19_0.VD2.n2 GNDA 0.098642f
C435 two_stage_opamp_dummy_magic_19_0.VD2.t13 GNDA 0.04446f
C436 two_stage_opamp_dummy_magic_19_0.VD2.t19 GNDA 0.04446f
C437 two_stage_opamp_dummy_magic_19_0.VD2.n3 GNDA 0.126282f
C438 two_stage_opamp_dummy_magic_19_0.VD2.t11 GNDA 0.04446f
C439 two_stage_opamp_dummy_magic_19_0.VD2.t10 GNDA 0.04446f
C440 two_stage_opamp_dummy_magic_19_0.VD2.n4 GNDA 0.122904f
C441 two_stage_opamp_dummy_magic_19_0.VD2.n5 GNDA 0.671139f
C442 two_stage_opamp_dummy_magic_19_0.VD2.t5 GNDA 0.04446f
C443 two_stage_opamp_dummy_magic_19_0.VD2.t1 GNDA 0.04446f
C444 two_stage_opamp_dummy_magic_19_0.VD2.n6 GNDA 0.126478f
C445 two_stage_opamp_dummy_magic_19_0.VD2.t21 GNDA 0.04446f
C446 two_stage_opamp_dummy_magic_19_0.VD2.t4 GNDA 0.04446f
C447 two_stage_opamp_dummy_magic_19_0.VD2.n7 GNDA 0.122904f
C448 two_stage_opamp_dummy_magic_19_0.VD2.n8 GNDA 0.666497f
C449 two_stage_opamp_dummy_magic_19_0.VD2.n9 GNDA 0.077064f
C450 two_stage_opamp_dummy_magic_19_0.VD2.t17 GNDA 0.04446f
C451 two_stage_opamp_dummy_magic_19_0.VD2.t6 GNDA 0.04446f
C452 two_stage_opamp_dummy_magic_19_0.VD2.n10 GNDA 0.126021f
C453 two_stage_opamp_dummy_magic_19_0.VD2.t20 GNDA 0.04446f
C454 two_stage_opamp_dummy_magic_19_0.VD2.t9 GNDA 0.04446f
C455 two_stage_opamp_dummy_magic_19_0.VD2.n11 GNDA 0.122578f
C456 two_stage_opamp_dummy_magic_19_0.VD2.n12 GNDA 0.688028f
C457 two_stage_opamp_dummy_magic_19_0.VD2.t7 GNDA 0.04446f
C458 two_stage_opamp_dummy_magic_19_0.VD2.t0 GNDA 0.04446f
C459 two_stage_opamp_dummy_magic_19_0.VD2.n13 GNDA 0.122578f
C460 two_stage_opamp_dummy_magic_19_0.VD2.t2 GNDA 0.04446f
C461 two_stage_opamp_dummy_magic_19_0.VD2.t18 GNDA 0.04446f
C462 two_stage_opamp_dummy_magic_19_0.VD2.n14 GNDA 0.126021f
C463 two_stage_opamp_dummy_magic_19_0.VD2.t14 GNDA 0.04446f
C464 two_stage_opamp_dummy_magic_19_0.VD2.t15 GNDA 0.04446f
C465 two_stage_opamp_dummy_magic_19_0.VD2.n15 GNDA 0.122578f
C466 two_stage_opamp_dummy_magic_19_0.VD2.n16 GNDA 0.688028f
C467 two_stage_opamp_dummy_magic_19_0.VD2.t8 GNDA 0.04446f
C468 two_stage_opamp_dummy_magic_19_0.VD2.t3 GNDA 0.04446f
C469 two_stage_opamp_dummy_magic_19_0.VD2.n17 GNDA 0.122578f
C470 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t0 GNDA 0.015138f
C471 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t15 GNDA 0.015138f
C472 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n0 GNDA 0.037962f
C473 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t16 GNDA 0.015138f
C474 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t13 GNDA 0.015138f
C475 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n1 GNDA 0.037762f
C476 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n2 GNDA 0.335688f
C477 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t14 GNDA 0.015138f
C478 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t2 GNDA 0.015138f
C479 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n3 GNDA 0.030276f
C480 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n4 GNDA 0.05628f
C481 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t1 GNDA 0.190995f
C482 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t3 GNDA 0.030276f
C483 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t7 GNDA 0.030276f
C484 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n5 GNDA 0.0707f
C485 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t9 GNDA 0.030276f
C486 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t8 GNDA 0.030276f
C487 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n6 GNDA 0.069684f
C488 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n7 GNDA 0.459076f
C489 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t12 GNDA 0.030276f
C490 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t6 GNDA 0.030276f
C491 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n8 GNDA 0.069684f
C492 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n9 GNDA 0.235344f
C493 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t11 GNDA 0.030276f
C494 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t5 GNDA 0.030276f
C495 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n10 GNDA 0.069684f
C496 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n11 GNDA 0.235344f
C497 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t10 GNDA 0.030276f
C498 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.t4 GNDA 0.030276f
C499 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n12 GNDA 0.069684f
C500 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n13 GNDA 0.297878f
C501 two_stage_opamp_dummy_magic_19_0.V_CMFB_S3.n14 GNDA 1.29708f
C502 bgr_9_0.V_CMFB_S3 GNDA 0.843286f
C503 two_stage_opamp_dummy_magic_19_0.Y.t5 GNDA 0.063779f
C504 two_stage_opamp_dummy_magic_19_0.Y.t3 GNDA 0.063779f
C505 two_stage_opamp_dummy_magic_19_0.Y.n0 GNDA 0.134708f
C506 two_stage_opamp_dummy_magic_19_0.Y.t15 GNDA 0.063779f
C507 two_stage_opamp_dummy_magic_19_0.Y.t10 GNDA 0.063779f
C508 two_stage_opamp_dummy_magic_19_0.Y.n1 GNDA 0.163887f
C509 two_stage_opamp_dummy_magic_19_0.Y.t8 GNDA 0.063779f
C510 two_stage_opamp_dummy_magic_19_0.Y.t1 GNDA 0.063779f
C511 two_stage_opamp_dummy_magic_19_0.Y.n2 GNDA 0.160217f
C512 two_stage_opamp_dummy_magic_19_0.Y.n3 GNDA 0.856711f
C513 two_stage_opamp_dummy_magic_19_0.Y.t7 GNDA 0.063779f
C514 two_stage_opamp_dummy_magic_19_0.Y.t6 GNDA 0.063779f
C515 two_stage_opamp_dummy_magic_19_0.Y.n4 GNDA 0.160217f
C516 two_stage_opamp_dummy_magic_19_0.Y.n5 GNDA 0.437479f
C517 two_stage_opamp_dummy_magic_19_0.Y.t2 GNDA 0.063779f
C518 two_stage_opamp_dummy_magic_19_0.Y.t12 GNDA 0.063779f
C519 two_stage_opamp_dummy_magic_19_0.Y.n6 GNDA 0.163887f
C520 two_stage_opamp_dummy_magic_19_0.Y.t9 GNDA 0.063779f
C521 two_stage_opamp_dummy_magic_19_0.Y.t4 GNDA 0.063779f
C522 two_stage_opamp_dummy_magic_19_0.Y.n7 GNDA 0.160217f
C523 two_stage_opamp_dummy_magic_19_0.Y.n8 GNDA 0.856711f
C524 two_stage_opamp_dummy_magic_19_0.Y.n9 GNDA 0.058312f
C525 two_stage_opamp_dummy_magic_19_0.Y.n10 GNDA 0.662444f
C526 two_stage_opamp_dummy_magic_19_0.Y.n11 GNDA 0.059027f
C527 two_stage_opamp_dummy_magic_19_0.Y.n12 GNDA 0.053999f
C528 two_stage_opamp_dummy_magic_19_0.Y.t22 GNDA 0.027334f
C529 two_stage_opamp_dummy_magic_19_0.Y.t19 GNDA 0.027334f
C530 two_stage_opamp_dummy_magic_19_0.Y.n13 GNDA 0.059475f
C531 two_stage_opamp_dummy_magic_19_0.Y.n14 GNDA 0.243865f
C532 two_stage_opamp_dummy_magic_19_0.Y.n15 GNDA 0.09088f
C533 two_stage_opamp_dummy_magic_19_0.Y.t23 GNDA 0.027334f
C534 two_stage_opamp_dummy_magic_19_0.Y.t17 GNDA 0.027334f
C535 two_stage_opamp_dummy_magic_19_0.Y.n16 GNDA 0.059475f
C536 two_stage_opamp_dummy_magic_19_0.Y.n17 GNDA 0.234771f
C537 two_stage_opamp_dummy_magic_19_0.Y.n18 GNDA 0.100566f
C538 two_stage_opamp_dummy_magic_19_0.Y.t16 GNDA 0.027334f
C539 two_stage_opamp_dummy_magic_19_0.Y.t20 GNDA 0.027334f
C540 two_stage_opamp_dummy_magic_19_0.Y.n19 GNDA 0.059475f
C541 two_stage_opamp_dummy_magic_19_0.Y.n20 GNDA 0.234771f
C542 two_stage_opamp_dummy_magic_19_0.Y.n21 GNDA 0.059027f
C543 two_stage_opamp_dummy_magic_19_0.Y.n22 GNDA 0.059027f
C544 two_stage_opamp_dummy_magic_19_0.Y.t18 GNDA 0.027334f
C545 two_stage_opamp_dummy_magic_19_0.Y.t24 GNDA 0.027334f
C546 two_stage_opamp_dummy_magic_19_0.Y.n23 GNDA 0.059475f
C547 two_stage_opamp_dummy_magic_19_0.Y.n24 GNDA 0.234771f
C548 two_stage_opamp_dummy_magic_19_0.Y.n25 GNDA 0.053999f
C549 two_stage_opamp_dummy_magic_19_0.Y.t13 GNDA 0.027334f
C550 two_stage_opamp_dummy_magic_19_0.Y.t14 GNDA 0.027334f
C551 two_stage_opamp_dummy_magic_19_0.Y.n26 GNDA 0.059475f
C552 two_stage_opamp_dummy_magic_19_0.Y.n27 GNDA 0.234771f
C553 two_stage_opamp_dummy_magic_19_0.Y.n28 GNDA 0.09088f
C554 two_stage_opamp_dummy_magic_19_0.Y.t0 GNDA 0.027334f
C555 two_stage_opamp_dummy_magic_19_0.Y.t21 GNDA 0.027334f
C556 two_stage_opamp_dummy_magic_19_0.Y.n29 GNDA 0.059475f
C557 two_stage_opamp_dummy_magic_19_0.Y.n30 GNDA 0.239132f
C558 two_stage_opamp_dummy_magic_19_0.Y.n31 GNDA 0.153891f
C559 two_stage_opamp_dummy_magic_19_0.Y.n32 GNDA 0.433668f
C560 two_stage_opamp_dummy_magic_19_0.Y.t25 GNDA 0.038267f
C561 two_stage_opamp_dummy_magic_19_0.Y.t42 GNDA 0.038267f
C562 two_stage_opamp_dummy_magic_19_0.Y.t29 GNDA 0.038267f
C563 two_stage_opamp_dummy_magic_19_0.Y.t45 GNDA 0.038267f
C564 two_stage_opamp_dummy_magic_19_0.Y.t32 GNDA 0.038267f
C565 two_stage_opamp_dummy_magic_19_0.Y.t48 GNDA 0.046467f
C566 two_stage_opamp_dummy_magic_19_0.Y.n33 GNDA 0.046467f
C567 two_stage_opamp_dummy_magic_19_0.Y.n34 GNDA 0.030067f
C568 two_stage_opamp_dummy_magic_19_0.Y.n35 GNDA 0.030067f
C569 two_stage_opamp_dummy_magic_19_0.Y.n36 GNDA 0.030067f
C570 two_stage_opamp_dummy_magic_19_0.Y.n37 GNDA 0.024942f
C571 two_stage_opamp_dummy_magic_19_0.Y.t38 GNDA 0.038267f
C572 two_stage_opamp_dummy_magic_19_0.Y.t34 GNDA 0.038267f
C573 two_stage_opamp_dummy_magic_19_0.Y.t39 GNDA 0.038267f
C574 two_stage_opamp_dummy_magic_19_0.Y.t53 GNDA 0.046467f
C575 two_stage_opamp_dummy_magic_19_0.Y.n38 GNDA 0.046467f
C576 two_stage_opamp_dummy_magic_19_0.Y.n39 GNDA 0.030067f
C577 two_stage_opamp_dummy_magic_19_0.Y.n40 GNDA 0.024942f
C578 two_stage_opamp_dummy_magic_19_0.Y.n41 GNDA 0.020627f
C579 two_stage_opamp_dummy_magic_19_0.Y.t44 GNDA 0.058767f
C580 two_stage_opamp_dummy_magic_19_0.Y.t31 GNDA 0.058767f
C581 two_stage_opamp_dummy_magic_19_0.Y.t47 GNDA 0.058767f
C582 two_stage_opamp_dummy_magic_19_0.Y.t33 GNDA 0.058767f
C583 two_stage_opamp_dummy_magic_19_0.Y.t49 GNDA 0.058767f
C584 two_stage_opamp_dummy_magic_19_0.Y.t35 GNDA 0.066809f
C585 two_stage_opamp_dummy_magic_19_0.Y.n42 GNDA 0.060293f
C586 two_stage_opamp_dummy_magic_19_0.Y.n43 GNDA 0.036901f
C587 two_stage_opamp_dummy_magic_19_0.Y.n44 GNDA 0.036901f
C588 two_stage_opamp_dummy_magic_19_0.Y.n45 GNDA 0.036901f
C589 two_stage_opamp_dummy_magic_19_0.Y.n46 GNDA 0.031775f
C590 two_stage_opamp_dummy_magic_19_0.Y.t27 GNDA 0.058767f
C591 two_stage_opamp_dummy_magic_19_0.Y.t50 GNDA 0.058767f
C592 two_stage_opamp_dummy_magic_19_0.Y.t28 GNDA 0.058767f
C593 two_stage_opamp_dummy_magic_19_0.Y.t41 GNDA 0.066809f
C594 two_stage_opamp_dummy_magic_19_0.Y.n47 GNDA 0.060293f
C595 two_stage_opamp_dummy_magic_19_0.Y.n48 GNDA 0.036901f
C596 two_stage_opamp_dummy_magic_19_0.Y.n49 GNDA 0.031775f
C597 two_stage_opamp_dummy_magic_19_0.Y.n50 GNDA 0.020627f
C598 two_stage_opamp_dummy_magic_19_0.Y.n51 GNDA 0.060216f
C599 two_stage_opamp_dummy_magic_19_0.Y.n52 GNDA 0.468971f
C600 two_stage_opamp_dummy_magic_19_0.Y.t54 GNDA 0.120268f
C601 two_stage_opamp_dummy_magic_19_0.Y.t40 GNDA 0.120268f
C602 two_stage_opamp_dummy_magic_19_0.Y.t26 GNDA 0.120268f
C603 two_stage_opamp_dummy_magic_19_0.Y.t43 GNDA 0.120268f
C604 two_stage_opamp_dummy_magic_19_0.Y.t30 GNDA 0.128094f
C605 two_stage_opamp_dummy_magic_19_0.Y.n53 GNDA 0.101509f
C606 two_stage_opamp_dummy_magic_19_0.Y.n54 GNDA 0.057401f
C607 two_stage_opamp_dummy_magic_19_0.Y.n55 GNDA 0.057401f
C608 two_stage_opamp_dummy_magic_19_0.Y.n56 GNDA 0.052276f
C609 two_stage_opamp_dummy_magic_19_0.Y.t37 GNDA 0.120268f
C610 two_stage_opamp_dummy_magic_19_0.Y.t51 GNDA 0.120268f
C611 two_stage_opamp_dummy_magic_19_0.Y.t46 GNDA 0.120268f
C612 two_stage_opamp_dummy_magic_19_0.Y.t52 GNDA 0.120268f
C613 two_stage_opamp_dummy_magic_19_0.Y.t36 GNDA 0.128094f
C614 two_stage_opamp_dummy_magic_19_0.Y.n57 GNDA 0.101509f
C615 two_stage_opamp_dummy_magic_19_0.Y.n58 GNDA 0.057401f
C616 two_stage_opamp_dummy_magic_19_0.Y.n59 GNDA 0.057401f
C617 two_stage_opamp_dummy_magic_19_0.Y.n60 GNDA 0.052276f
C618 two_stage_opamp_dummy_magic_19_0.Y.n61 GNDA 0.046271f
C619 two_stage_opamp_dummy_magic_19_0.Y.n62 GNDA 1.00986f
C620 two_stage_opamp_dummy_magic_19_0.Y.t11 GNDA 0.878241f
C621 two_stage_opamp_dummy_magic_19_0.VD3.t1 GNDA 0.058707f
C622 two_stage_opamp_dummy_magic_19_0.VD3.t9 GNDA 0.058707f
C623 two_stage_opamp_dummy_magic_19_0.VD3.t15 GNDA 0.058707f
C624 two_stage_opamp_dummy_magic_19_0.VD3.n0 GNDA 0.147477f
C625 two_stage_opamp_dummy_magic_19_0.VD3.n1 GNDA 0.402692f
C626 two_stage_opamp_dummy_magic_19_0.VD3.t22 GNDA 0.208829f
C627 two_stage_opamp_dummy_magic_19_0.VD3.t23 GNDA 0.102932f
C628 two_stage_opamp_dummy_magic_19_0.VD3.t37 GNDA 0.058707f
C629 two_stage_opamp_dummy_magic_19_0.VD3.t34 GNDA 0.058707f
C630 two_stage_opamp_dummy_magic_19_0.VD3.n2 GNDA 0.150855f
C631 two_stage_opamp_dummy_magic_19_0.VD3.t35 GNDA 0.058707f
C632 two_stage_opamp_dummy_magic_19_0.VD3.t27 GNDA 0.058707f
C633 two_stage_opamp_dummy_magic_19_0.VD3.n3 GNDA 0.147477f
C634 two_stage_opamp_dummy_magic_19_0.VD3.n4 GNDA 0.788587f
C635 two_stage_opamp_dummy_magic_19_0.VD3.t30 GNDA 0.058707f
C636 two_stage_opamp_dummy_magic_19_0.VD3.t29 GNDA 0.058707f
C637 two_stage_opamp_dummy_magic_19_0.VD3.n5 GNDA 0.147477f
C638 two_stage_opamp_dummy_magic_19_0.VD3.n6 GNDA 0.402692f
C639 two_stage_opamp_dummy_magic_19_0.VD3.t31 GNDA 0.058707f
C640 two_stage_opamp_dummy_magic_19_0.VD3.t32 GNDA 0.058707f
C641 two_stage_opamp_dummy_magic_19_0.VD3.n7 GNDA 0.147477f
C642 two_stage_opamp_dummy_magic_19_0.VD3.n8 GNDA 0.402692f
C643 two_stage_opamp_dummy_magic_19_0.VD3.t33 GNDA 0.058707f
C644 two_stage_opamp_dummy_magic_19_0.VD3.t28 GNDA 0.058707f
C645 two_stage_opamp_dummy_magic_19_0.VD3.n9 GNDA 0.147477f
C646 two_stage_opamp_dummy_magic_19_0.VD3.n10 GNDA 0.402692f
C647 two_stage_opamp_dummy_magic_19_0.VD3.t26 GNDA 0.058707f
C648 two_stage_opamp_dummy_magic_19_0.VD3.t36 GNDA 0.058707f
C649 two_stage_opamp_dummy_magic_19_0.VD3.n11 GNDA 0.147477f
C650 two_stage_opamp_dummy_magic_19_0.VD3.n12 GNDA 0.569977f
C651 two_stage_opamp_dummy_magic_19_0.VD3.t5 GNDA 0.058707f
C652 two_stage_opamp_dummy_magic_19_0.VD3.t13 GNDA 0.058707f
C653 two_stage_opamp_dummy_magic_19_0.VD3.n13 GNDA 0.147477f
C654 two_stage_opamp_dummy_magic_19_0.VD3.n14 GNDA 0.402692f
C655 two_stage_opamp_dummy_magic_19_0.VD3.n15 GNDA 0.241623f
C656 two_stage_opamp_dummy_magic_19_0.VD3.n16 GNDA 0.156154f
C657 two_stage_opamp_dummy_magic_19_0.VD3.t25 GNDA 0.208829f
C658 two_stage_opamp_dummy_magic_19_0.VD3.n17 GNDA 0.373262f
C659 two_stage_opamp_dummy_magic_19_0.VD3.t24 GNDA 0.497708f
C660 two_stage_opamp_dummy_magic_19_0.VD3.t4 GNDA 0.392499f
C661 two_stage_opamp_dummy_magic_19_0.VD3.t12 GNDA 0.392499f
C662 two_stage_opamp_dummy_magic_19_0.VD3.t8 GNDA 0.392499f
C663 two_stage_opamp_dummy_magic_19_0.VD3.t14 GNDA 0.392499f
C664 two_stage_opamp_dummy_magic_19_0.VD3.t18 GNDA 0.392499f
C665 two_stage_opamp_dummy_magic_19_0.VD3.t0 GNDA 0.392499f
C666 two_stage_opamp_dummy_magic_19_0.VD3.t6 GNDA 0.392499f
C667 two_stage_opamp_dummy_magic_19_0.VD3.t2 GNDA 0.392499f
C668 two_stage_opamp_dummy_magic_19_0.VD3.t10 GNDA 0.392499f
C669 two_stage_opamp_dummy_magic_19_0.VD3.t16 GNDA 0.392499f
C670 two_stage_opamp_dummy_magic_19_0.VD3.t21 GNDA 0.497708f
C671 two_stage_opamp_dummy_magic_19_0.VD3.n18 GNDA 0.373262f
C672 two_stage_opamp_dummy_magic_19_0.VD3.t20 GNDA 0.102932f
C673 two_stage_opamp_dummy_magic_19_0.VD3.n19 GNDA 0.158682f
C674 two_stage_opamp_dummy_magic_19_0.VD3.t11 GNDA 0.058707f
C675 two_stage_opamp_dummy_magic_19_0.VD3.t17 GNDA 0.058707f
C676 two_stage_opamp_dummy_magic_19_0.VD3.n20 GNDA 0.147477f
C677 two_stage_opamp_dummy_magic_19_0.VD3.n21 GNDA 0.458507f
C678 two_stage_opamp_dummy_magic_19_0.VD3.t7 GNDA 0.058707f
C679 two_stage_opamp_dummy_magic_19_0.VD3.t3 GNDA 0.058707f
C680 two_stage_opamp_dummy_magic_19_0.VD3.n22 GNDA 0.147477f
C681 two_stage_opamp_dummy_magic_19_0.VD3.n23 GNDA 0.402692f
C682 two_stage_opamp_dummy_magic_19_0.VD3.n24 GNDA 0.402692f
C683 two_stage_opamp_dummy_magic_19_0.VD3.n25 GNDA 0.147477f
C684 two_stage_opamp_dummy_magic_19_0.VD3.t19 GNDA 0.058707f
C685 two_stage_opamp_dummy_magic_19_0.Vb2.t2 GNDA 0.030271f
C686 two_stage_opamp_dummy_magic_19_0.Vb2.t0 GNDA 0.030271f
C687 two_stage_opamp_dummy_magic_19_0.Vb2.n0 GNDA 0.053397f
C688 two_stage_opamp_dummy_magic_19_0.Vb2.t1 GNDA 0.052349f
C689 two_stage_opamp_dummy_magic_19_0.Vb2.n1 GNDA 0.145198f
C690 two_stage_opamp_dummy_magic_19_0.Vb2.t28 GNDA 0.030909f
C691 two_stage_opamp_dummy_magic_19_0.Vb2.n2 GNDA 0.092586f
C692 two_stage_opamp_dummy_magic_19_0.Vb2.t26 GNDA 0.042811f
C693 two_stage_opamp_dummy_magic_19_0.Vb2.t19 GNDA 0.042811f
C694 two_stage_opamp_dummy_magic_19_0.Vb2.t13 GNDA 0.049404f
C695 two_stage_opamp_dummy_magic_19_0.Vb2.n3 GNDA 0.040111f
C696 two_stage_opamp_dummy_magic_19_0.Vb2.n4 GNDA 0.02417f
C697 two_stage_opamp_dummy_magic_19_0.Vb2.t31 GNDA 0.042811f
C698 two_stage_opamp_dummy_magic_19_0.Vb2.t11 GNDA 0.042811f
C699 two_stage_opamp_dummy_magic_19_0.Vb2.t15 GNDA 0.042811f
C700 two_stage_opamp_dummy_magic_19_0.Vb2.t21 GNDA 0.042811f
C701 two_stage_opamp_dummy_magic_19_0.Vb2.t17 GNDA 0.042811f
C702 two_stage_opamp_dummy_magic_19_0.Vb2.t24 GNDA 0.049404f
C703 two_stage_opamp_dummy_magic_19_0.Vb2.n5 GNDA 0.040111f
C704 two_stage_opamp_dummy_magic_19_0.Vb2.n6 GNDA 0.024649f
C705 two_stage_opamp_dummy_magic_19_0.Vb2.n7 GNDA 0.024649f
C706 two_stage_opamp_dummy_magic_19_0.Vb2.n8 GNDA 0.024649f
C707 two_stage_opamp_dummy_magic_19_0.Vb2.n9 GNDA 0.02417f
C708 two_stage_opamp_dummy_magic_19_0.Vb2.t22 GNDA 0.044325f
C709 two_stage_opamp_dummy_magic_19_0.Vb2.n10 GNDA 0.039367f
C710 two_stage_opamp_dummy_magic_19_0.Vb2.t32 GNDA 0.042811f
C711 two_stage_opamp_dummy_magic_19_0.Vb2.t30 GNDA 0.042811f
C712 two_stage_opamp_dummy_magic_19_0.Vb2.t29 GNDA 0.042811f
C713 two_stage_opamp_dummy_magic_19_0.Vb2.t25 GNDA 0.042811f
C714 two_stage_opamp_dummy_magic_19_0.Vb2.t18 GNDA 0.042811f
C715 two_stage_opamp_dummy_magic_19_0.Vb2.t12 GNDA 0.049404f
C716 two_stage_opamp_dummy_magic_19_0.Vb2.n11 GNDA 0.040111f
C717 two_stage_opamp_dummy_magic_19_0.Vb2.n12 GNDA 0.024649f
C718 two_stage_opamp_dummy_magic_19_0.Vb2.n13 GNDA 0.024649f
C719 two_stage_opamp_dummy_magic_19_0.Vb2.n14 GNDA 0.024649f
C720 two_stage_opamp_dummy_magic_19_0.Vb2.n15 GNDA 0.02417f
C721 two_stage_opamp_dummy_magic_19_0.Vb2.t20 GNDA 0.042811f
C722 two_stage_opamp_dummy_magic_19_0.Vb2.t27 GNDA 0.042811f
C723 two_stage_opamp_dummy_magic_19_0.Vb2.t23 GNDA 0.049404f
C724 two_stage_opamp_dummy_magic_19_0.Vb2.n16 GNDA 0.040111f
C725 two_stage_opamp_dummy_magic_19_0.Vb2.n17 GNDA 0.02417f
C726 two_stage_opamp_dummy_magic_19_0.Vb2.t14 GNDA 0.044325f
C727 two_stage_opamp_dummy_magic_19_0.Vb2.n18 GNDA 0.039171f
C728 two_stage_opamp_dummy_magic_19_0.Vb2.n19 GNDA 0.306521f
C729 two_stage_opamp_dummy_magic_19_0.Vb2.n20 GNDA 0.151435f
C730 two_stage_opamp_dummy_magic_19_0.Vb2.t16 GNDA 0.052349f
C731 two_stage_opamp_dummy_magic_19_0.Vb2.n21 GNDA 0.70951f
C732 two_stage_opamp_dummy_magic_19_0.Vb2.n22 GNDA 0.028446f
C733 two_stage_opamp_dummy_magic_19_0.Vb2.n23 GNDA 0.793734f
C734 two_stage_opamp_dummy_magic_19_0.Vb2.n24 GNDA 0.028446f
C735 two_stage_opamp_dummy_magic_19_0.Vb2.n25 GNDA 0.200747f
C736 two_stage_opamp_dummy_magic_19_0.Vb2.n26 GNDA 0.029281f
C737 two_stage_opamp_dummy_magic_19_0.Vb2.n27 GNDA 0.297738f
C738 two_stage_opamp_dummy_magic_19_0.Vb2.n28 GNDA 0.028446f
C739 bgr_9_0.cap_res2.t6 GNDA 0.358835f
C740 bgr_9_0.cap_res2.t12 GNDA 0.360135f
C741 bgr_9_0.cap_res2.t14 GNDA 0.340877f
C742 bgr_9_0.cap_res2.t0 GNDA 0.358835f
C743 bgr_9_0.cap_res2.t5 GNDA 0.360135f
C744 bgr_9_0.cap_res2.t8 GNDA 0.340877f
C745 bgr_9_0.cap_res2.t4 GNDA 0.358835f
C746 bgr_9_0.cap_res2.t10 GNDA 0.360135f
C747 bgr_9_0.cap_res2.t13 GNDA 0.340877f
C748 bgr_9_0.cap_res2.t19 GNDA 0.358835f
C749 bgr_9_0.cap_res2.t3 GNDA 0.360135f
C750 bgr_9_0.cap_res2.t7 GNDA 0.340877f
C751 bgr_9_0.cap_res2.t15 GNDA 0.358835f
C752 bgr_9_0.cap_res2.t18 GNDA 0.360135f
C753 bgr_9_0.cap_res2.t1 GNDA 0.340877f
C754 bgr_9_0.cap_res2.n0 GNDA 0.240527f
C755 bgr_9_0.cap_res2.t2 GNDA 0.191544f
C756 bgr_9_0.cap_res2.n1 GNDA 0.260978f
C757 bgr_9_0.cap_res2.t9 GNDA 0.191544f
C758 bgr_9_0.cap_res2.n2 GNDA 0.260978f
C759 bgr_9_0.cap_res2.t16 GNDA 0.191544f
C760 bgr_9_0.cap_res2.n3 GNDA 0.260978f
C761 bgr_9_0.cap_res2.t11 GNDA 0.191544f
C762 bgr_9_0.cap_res2.n4 GNDA 0.260978f
C763 bgr_9_0.cap_res2.t17 GNDA 0.364682f
C764 bgr_9_0.cap_res2.t20 GNDA 0.085466f
C765 bgr_9_0.1st_Vout_2.n0 GNDA 0.722974f
C766 bgr_9_0.1st_Vout_2.n1 GNDA 0.237543f
C767 bgr_9_0.1st_Vout_2.n2 GNDA 1.43086f
C768 bgr_9_0.1st_Vout_2.n3 GNDA 0.104357f
C769 bgr_9_0.1st_Vout_2.n4 GNDA 1.45767f
C770 bgr_9_0.1st_Vout_2.n5 GNDA 0.010417f
C771 bgr_9_0.1st_Vout_2.t0 GNDA 0.015189f
C772 bgr_9_0.1st_Vout_2.n6 GNDA 0.157567f
C773 bgr_9_0.1st_Vout_2.t33 GNDA 0.017308f
C774 bgr_9_0.1st_Vout_2.n8 GNDA 0.018209f
C775 bgr_9_0.1st_Vout_2.t24 GNDA 0.010986f
C776 bgr_9_0.1st_Vout_2.t13 GNDA 0.010986f
C777 bgr_9_0.1st_Vout_2.n9 GNDA 0.024439f
C778 bgr_9_0.1st_Vout_2.t28 GNDA 0.288462f
C779 bgr_9_0.1st_Vout_2.t17 GNDA 0.293375f
C780 bgr_9_0.1st_Vout_2.t12 GNDA 0.288462f
C781 bgr_9_0.1st_Vout_2.t32 GNDA 0.288462f
C782 bgr_9_0.1st_Vout_2.t35 GNDA 0.293375f
C783 bgr_9_0.1st_Vout_2.t11 GNDA 0.293375f
C784 bgr_9_0.1st_Vout_2.t31 GNDA 0.288462f
C785 bgr_9_0.1st_Vout_2.t23 GNDA 0.288462f
C786 bgr_9_0.1st_Vout_2.t26 GNDA 0.293375f
C787 bgr_9_0.1st_Vout_2.t30 GNDA 0.293375f
C788 bgr_9_0.1st_Vout_2.t22 GNDA 0.288462f
C789 bgr_9_0.1st_Vout_2.t15 GNDA 0.288462f
C790 bgr_9_0.1st_Vout_2.t19 GNDA 0.293375f
C791 bgr_9_0.1st_Vout_2.t36 GNDA 0.293375f
C792 bgr_9_0.1st_Vout_2.t29 GNDA 0.288462f
C793 bgr_9_0.1st_Vout_2.t21 GNDA 0.288462f
C794 bgr_9_0.1st_Vout_2.t25 GNDA 0.293375f
C795 bgr_9_0.1st_Vout_2.t18 GNDA 0.293375f
C796 bgr_9_0.1st_Vout_2.t14 GNDA 0.288462f
C797 bgr_9_0.1st_Vout_2.t20 GNDA 0.288462f
C798 bgr_9_0.1st_Vout_2.t34 GNDA 0.018845f
C799 bgr_9_0.1st_Vout_2.n10 GNDA 0.018209f
C800 bgr_9_0.1st_Vout_2.t27 GNDA 0.010986f
C801 bgr_9_0.1st_Vout_2.t16 GNDA 0.010986f
C802 bgr_9_0.1st_Vout_2.n11 GNDA 0.024439f
C803 bgr_9_0.1st_Vout_2.n12 GNDA 0.017468f
C804 bgr_9_0.1st_Vout_1.n0 GNDA 0.538712f
C805 bgr_9_0.1st_Vout_1.n1 GNDA 0.236313f
C806 bgr_9_0.1st_Vout_1.n2 GNDA 0.973284f
C807 bgr_9_0.1st_Vout_1.n3 GNDA 0.907198f
C808 bgr_9_0.1st_Vout_1.n4 GNDA 0.891647f
C809 bgr_9_0.1st_Vout_1.t11 GNDA 0.358463f
C810 bgr_9_0.1st_Vout_1.t15 GNDA 0.35246f
C811 bgr_9_0.1st_Vout_1.t29 GNDA 0.358463f
C812 bgr_9_0.1st_Vout_1.t35 GNDA 0.35246f
C813 bgr_9_0.1st_Vout_1.t31 GNDA 0.358463f
C814 bgr_9_0.1st_Vout_1.t34 GNDA 0.35246f
C815 bgr_9_0.1st_Vout_1.t20 GNDA 0.358463f
C816 bgr_9_0.1st_Vout_1.t28 GNDA 0.35246f
C817 bgr_9_0.1st_Vout_1.t24 GNDA 0.358463f
C818 bgr_9_0.1st_Vout_1.t27 GNDA 0.35246f
C819 bgr_9_0.1st_Vout_1.t14 GNDA 0.358463f
C820 bgr_9_0.1st_Vout_1.t19 GNDA 0.35246f
C821 bgr_9_0.1st_Vout_1.t30 GNDA 0.358463f
C822 bgr_9_0.1st_Vout_1.t33 GNDA 0.35246f
C823 bgr_9_0.1st_Vout_1.t18 GNDA 0.358463f
C824 bgr_9_0.1st_Vout_1.t26 GNDA 0.35246f
C825 bgr_9_0.1st_Vout_1.t23 GNDA 0.358463f
C826 bgr_9_0.1st_Vout_1.t25 GNDA 0.35246f
C827 bgr_9_0.1st_Vout_1.t17 GNDA 0.35246f
C828 bgr_9_0.1st_Vout_1.t12 GNDA 0.35246f
C829 bgr_9_0.1st_Vout_1.t21 GNDA 0.023025f
C830 bgr_9_0.1st_Vout_1.n5 GNDA 0.715456f
C831 bgr_9_0.1st_Vout_1.n6 GNDA 0.022249f
C832 bgr_9_0.1st_Vout_1.n7 GNDA 0.104637f
C833 bgr_9_0.1st_Vout_1.t36 GNDA 0.013423f
C834 bgr_9_0.1st_Vout_1.t16 GNDA 0.013423f
C835 bgr_9_0.1st_Vout_1.n8 GNDA 0.029862f
C836 bgr_9_0.1st_Vout_1.n9 GNDA 0.082514f
C837 bgr_9_0.1st_Vout_1.t10 GNDA 0.018559f
C838 bgr_9_0.1st_Vout_1.n10 GNDA 0.012728f
C839 bgr_9_0.1st_Vout_1.n11 GNDA 0.192525f
C840 bgr_9_0.1st_Vout_1.n12 GNDA 0.011517f
C841 bgr_9_0.1st_Vout_1.n13 GNDA 0.048842f
C842 bgr_9_0.1st_Vout_1.n14 GNDA 0.021343f
C843 bgr_9_0.1st_Vout_1.n15 GNDA 0.078667f
C844 bgr_9_0.1st_Vout_1.n16 GNDA 0.038771f
C845 bgr_9_0.1st_Vout_1.t32 GNDA 0.013423f
C846 bgr_9_0.1st_Vout_1.t22 GNDA 0.013423f
C847 bgr_9_0.1st_Vout_1.n17 GNDA 0.029862f
C848 bgr_9_0.1st_Vout_1.n18 GNDA 0.082514f
C849 bgr_9_0.1st_Vout_1.n19 GNDA 0.022249f
C850 bgr_9_0.1st_Vout_1.n20 GNDA 0.104637f
C851 bgr_9_0.1st_Vout_1.t13 GNDA 0.021069f
C852 bgr_9_0.V_mir1.t8 GNDA 0.019293f
C853 bgr_9_0.V_mir1.t1 GNDA 0.02939f
C854 bgr_9_0.V_mir1.t5 GNDA 0.023151f
C855 bgr_9_0.V_mir1.t18 GNDA 0.023151f
C856 bgr_9_0.V_mir1.t20 GNDA 0.037369f
C857 bgr_9_0.V_mir1.n0 GNDA 0.041731f
C858 bgr_9_0.V_mir1.n1 GNDA 0.028507f
C859 bgr_9_0.V_mir1.n2 GNDA 0.044354f
C860 bgr_9_0.V_mir1.t2 GNDA 0.019293f
C861 bgr_9_0.V_mir1.t6 GNDA 0.019293f
C862 bgr_9_0.V_mir1.n3 GNDA 0.044322f
C863 bgr_9_0.V_mir1.n4 GNDA 0.109787f
C864 bgr_9_0.V_mir1.n5 GNDA 0.025223f
C865 bgr_9_0.V_mir1.t15 GNDA 0.041163f
C866 bgr_9_0.V_mir1.n6 GNDA 0.027381f
C867 bgr_9_0.V_mir1.n7 GNDA 0.451535f
C868 bgr_9_0.V_mir1.n8 GNDA 0.146338f
C869 bgr_9_0.V_mir1.t3 GNDA 0.02939f
C870 bgr_9_0.V_mir1.t9 GNDA 0.023151f
C871 bgr_9_0.V_mir1.t17 GNDA 0.023151f
C872 bgr_9_0.V_mir1.t21 GNDA 0.037369f
C873 bgr_9_0.V_mir1.n9 GNDA 0.041731f
C874 bgr_9_0.V_mir1.n10 GNDA 0.028507f
C875 bgr_9_0.V_mir1.n11 GNDA 0.044354f
C876 bgr_9_0.V_mir1.t4 GNDA 0.019293f
C877 bgr_9_0.V_mir1.t10 GNDA 0.019293f
C878 bgr_9_0.V_mir1.n12 GNDA 0.044322f
C879 bgr_9_0.V_mir1.n13 GNDA 0.084938f
C880 bgr_9_0.V_mir1.n14 GNDA 0.051125f
C881 bgr_9_0.V_mir1.n15 GNDA 0.381359f
C882 bgr_9_0.V_mir1.t7 GNDA 0.02939f
C883 bgr_9_0.V_mir1.t11 GNDA 0.023151f
C884 bgr_9_0.V_mir1.t22 GNDA 0.023151f
C885 bgr_9_0.V_mir1.t19 GNDA 0.037369f
C886 bgr_9_0.V_mir1.n16 GNDA 0.041731f
C887 bgr_9_0.V_mir1.n17 GNDA 0.028507f
C888 bgr_9_0.V_mir1.n18 GNDA 0.044354f
C889 bgr_9_0.V_mir1.n19 GNDA 0.110886f
C890 bgr_9_0.V_mir1.n20 GNDA 0.044322f
C891 bgr_9_0.V_mir1.t12 GNDA 0.019293f
C892 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t14 GNDA 0.015138f
C893 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t2 GNDA 0.015138f
C894 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n0 GNDA 0.037946f
C895 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t1 GNDA 0.015138f
C896 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t16 GNDA 0.015138f
C897 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n1 GNDA 0.037745f
C898 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n2 GNDA 0.335479f
C899 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t0 GNDA 0.015138f
C900 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t13 GNDA 0.015138f
C901 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n3 GNDA 0.030276f
C902 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n4 GNDA 0.056304f
C903 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t15 GNDA 0.190995f
C904 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t6 GNDA 0.030276f
C905 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t11 GNDA 0.030276f
C906 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n5 GNDA 0.0707f
C907 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t4 GNDA 0.030276f
C908 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t8 GNDA 0.030276f
C909 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n6 GNDA 0.069684f
C910 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n7 GNDA 0.459076f
C911 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t5 GNDA 0.030276f
C912 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t10 GNDA 0.030276f
C913 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n8 GNDA 0.069684f
C914 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n9 GNDA 0.235344f
C915 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t7 GNDA 0.030276f
C916 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t12 GNDA 0.030276f
C917 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n10 GNDA 0.069684f
C918 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n11 GNDA 0.235344f
C919 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t9 GNDA 0.030276f
C920 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.t3 GNDA 0.030276f
C921 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n12 GNDA 0.069684f
C922 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n13 GNDA 0.297878f
C923 two_stage_opamp_dummy_magic_19_0.V_CMFB_S1.n14 GNDA 1.29708f
C924 bgr_9_0.V_CMFB_S1 GNDA 0.843505f
C925 bgr_9_0.Vin+.t7 GNDA 0.010641f
C926 bgr_9_0.Vin+.t8 GNDA 0.025236f
C927 bgr_9_0.Vin+.t9 GNDA 0.016404f
C928 bgr_9_0.Vin+.n0 GNDA 0.054125f
C929 bgr_9_0.Vin+.t6 GNDA 0.016404f
C930 bgr_9_0.Vin+.n1 GNDA 0.042119f
C931 bgr_9_0.Vin+.t10 GNDA 0.016404f
C932 bgr_9_0.Vin+.n2 GNDA 0.042687f
C933 bgr_9_0.Vin+.n3 GNDA 0.130116f
C934 bgr_9_0.Vin+.t4 GNDA 0.053203f
C935 bgr_9_0.Vin+.t3 GNDA 0.053203f
C936 bgr_9_0.Vin+.n4 GNDA 0.183813f
C937 bgr_9_0.Vin+.n5 GNDA 1.26385f
C938 bgr_9_0.Vin+.t2 GNDA 0.053203f
C939 bgr_9_0.Vin+.t5 GNDA 0.053203f
C940 bgr_9_0.Vin+.n6 GNDA 0.183813f
C941 bgr_9_0.Vin+.n7 GNDA 1.0517f
C942 bgr_9_0.Vin+.t1 GNDA 0.233821f
C943 bgr_9_0.Vin+.n8 GNDA 1.743f
C944 bgr_9_0.Vin+.t0 GNDA 0.173052f
C945 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t8 GNDA 0.066721f
C946 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t9 GNDA 0.065264f
C947 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n0 GNDA 0.49991f
C948 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t0 GNDA 0.309512f
C949 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t11 GNDA 0.047746f
C950 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t7 GNDA 0.017854f
C951 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n1 GNDA 0.056f
C952 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t13 GNDA 0.017854f
C953 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n2 GNDA 0.045842f
C954 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t10 GNDA 0.017854f
C955 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n3 GNDA 0.045842f
C956 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t12 GNDA 0.017854f
C957 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n4 GNDA 0.079873f
C958 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n5 GNDA 1.61828f
C959 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t2 GNDA 0.057905f
C960 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t5 GNDA 0.057905f
C961 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n6 GNDA 0.212469f
C962 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t6 GNDA 0.057905f
C963 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t4 GNDA 0.057905f
C964 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n7 GNDA 0.202767f
C965 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n8 GNDA 0.88956f
C966 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t3 GNDA 0.057905f
C967 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.t1 GNDA 0.057905f
C968 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n9 GNDA 0.202767f
C969 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n10 GNDA 0.639717f
C970 two_stage_opamp_dummy_magic_19_0.V_err_amp_ref.n11 GNDA 1.3379f
C971 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t13 GNDA 0.025582f
C972 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t14 GNDA 0.025582f
C973 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n0 GNDA 0.092232f
C974 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t11 GNDA 0.025582f
C975 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t12 GNDA 0.025582f
C976 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n1 GNDA 0.077093f
C977 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n2 GNDA 1.508f
C978 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t10 GNDA 0.313805f
C979 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t6 GNDA 0.076745f
C980 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t1 GNDA 0.076745f
C981 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n3 GNDA 0.25487f
C982 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t4 GNDA 0.076745f
C983 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t8 GNDA 0.076745f
C984 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n4 GNDA 0.246333f
C985 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n5 GNDA 0.921136f
C986 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t5 GNDA 0.076745f
C987 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t0 GNDA 0.076745f
C988 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n6 GNDA 0.246333f
C989 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n7 GNDA 0.47379f
C990 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t7 GNDA 0.076745f
C991 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t2 GNDA 0.076745f
C992 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n8 GNDA 0.246333f
C993 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n9 GNDA 0.47379f
C994 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t9 GNDA 0.076745f
C995 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.t3 GNDA 0.076745f
C996 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n10 GNDA 0.246333f
C997 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n11 GNDA 0.562302f
C998 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n12 GNDA 1.80918f
C999 two_stage_opamp_dummy_magic_19_0.V_CMFB_S2.n13 GNDA 2.24591f
C1000 bgr_9_0.V_CMFB_S2 GNDA 0.012791f
C1001 two_stage_opamp_dummy_magic_19_0.X.t13 GNDA 0.063779f
C1002 two_stage_opamp_dummy_magic_19_0.X.t3 GNDA 0.063779f
C1003 two_stage_opamp_dummy_magic_19_0.X.n0 GNDA 0.134708f
C1004 two_stage_opamp_dummy_magic_19_0.X.t12 GNDA 0.063779f
C1005 two_stage_opamp_dummy_magic_19_0.X.t21 GNDA 0.063779f
C1006 two_stage_opamp_dummy_magic_19_0.X.n1 GNDA 0.163887f
C1007 two_stage_opamp_dummy_magic_19_0.X.t2 GNDA 0.063779f
C1008 two_stage_opamp_dummy_magic_19_0.X.t22 GNDA 0.063779f
C1009 two_stage_opamp_dummy_magic_19_0.X.n2 GNDA 0.160217f
C1010 two_stage_opamp_dummy_magic_19_0.X.n3 GNDA 0.856711f
C1011 two_stage_opamp_dummy_magic_19_0.X.t10 GNDA 0.063779f
C1012 two_stage_opamp_dummy_magic_19_0.X.t9 GNDA 0.063779f
C1013 two_stage_opamp_dummy_magic_19_0.X.n4 GNDA 0.163887f
C1014 two_stage_opamp_dummy_magic_19_0.X.t7 GNDA 0.063779f
C1015 two_stage_opamp_dummy_magic_19_0.X.t11 GNDA 0.063779f
C1016 two_stage_opamp_dummy_magic_19_0.X.n5 GNDA 0.160217f
C1017 two_stage_opamp_dummy_magic_19_0.X.n6 GNDA 0.856711f
C1018 two_stage_opamp_dummy_magic_19_0.X.t20 GNDA 0.063779f
C1019 two_stage_opamp_dummy_magic_19_0.X.t8 GNDA 0.063779f
C1020 two_stage_opamp_dummy_magic_19_0.X.n7 GNDA 0.160217f
C1021 two_stage_opamp_dummy_magic_19_0.X.n8 GNDA 0.437479f
C1022 two_stage_opamp_dummy_magic_19_0.X.n9 GNDA 0.058312f
C1023 two_stage_opamp_dummy_magic_19_0.X.n10 GNDA 0.662444f
C1024 two_stage_opamp_dummy_magic_19_0.X.n11 GNDA 0.059027f
C1025 two_stage_opamp_dummy_magic_19_0.X.n12 GNDA 0.053999f
C1026 two_stage_opamp_dummy_magic_19_0.X.t0 GNDA 0.027334f
C1027 two_stage_opamp_dummy_magic_19_0.X.t19 GNDA 0.027334f
C1028 two_stage_opamp_dummy_magic_19_0.X.n13 GNDA 0.059475f
C1029 two_stage_opamp_dummy_magic_19_0.X.n14 GNDA 0.243865f
C1030 two_stage_opamp_dummy_magic_19_0.X.n15 GNDA 0.09088f
C1031 two_stage_opamp_dummy_magic_19_0.X.t5 GNDA 0.027334f
C1032 two_stage_opamp_dummy_magic_19_0.X.t14 GNDA 0.027334f
C1033 two_stage_opamp_dummy_magic_19_0.X.n16 GNDA 0.059475f
C1034 two_stage_opamp_dummy_magic_19_0.X.n17 GNDA 0.234771f
C1035 two_stage_opamp_dummy_magic_19_0.X.n18 GNDA 0.100566f
C1036 two_stage_opamp_dummy_magic_19_0.X.t24 GNDA 0.027334f
C1037 two_stage_opamp_dummy_magic_19_0.X.t1 GNDA 0.027334f
C1038 two_stage_opamp_dummy_magic_19_0.X.n19 GNDA 0.059475f
C1039 two_stage_opamp_dummy_magic_19_0.X.n20 GNDA 0.234771f
C1040 two_stage_opamp_dummy_magic_19_0.X.n21 GNDA 0.059027f
C1041 two_stage_opamp_dummy_magic_19_0.X.n22 GNDA 0.059027f
C1042 two_stage_opamp_dummy_magic_19_0.X.t15 GNDA 0.027334f
C1043 two_stage_opamp_dummy_magic_19_0.X.t16 GNDA 0.027334f
C1044 two_stage_opamp_dummy_magic_19_0.X.n23 GNDA 0.059475f
C1045 two_stage_opamp_dummy_magic_19_0.X.n24 GNDA 0.234771f
C1046 two_stage_opamp_dummy_magic_19_0.X.n25 GNDA 0.053999f
C1047 two_stage_opamp_dummy_magic_19_0.X.t6 GNDA 0.027334f
C1048 two_stage_opamp_dummy_magic_19_0.X.t23 GNDA 0.027334f
C1049 two_stage_opamp_dummy_magic_19_0.X.n26 GNDA 0.059475f
C1050 two_stage_opamp_dummy_magic_19_0.X.n27 GNDA 0.234771f
C1051 two_stage_opamp_dummy_magic_19_0.X.n28 GNDA 0.09088f
C1052 two_stage_opamp_dummy_magic_19_0.X.t18 GNDA 0.027334f
C1053 two_stage_opamp_dummy_magic_19_0.X.t4 GNDA 0.027334f
C1054 two_stage_opamp_dummy_magic_19_0.X.n29 GNDA 0.059475f
C1055 two_stage_opamp_dummy_magic_19_0.X.n30 GNDA 0.239132f
C1056 two_stage_opamp_dummy_magic_19_0.X.n31 GNDA 0.153891f
C1057 two_stage_opamp_dummy_magic_19_0.X.n32 GNDA 0.433668f
C1058 two_stage_opamp_dummy_magic_19_0.X.t52 GNDA 0.038267f
C1059 two_stage_opamp_dummy_magic_19_0.X.t38 GNDA 0.038267f
C1060 two_stage_opamp_dummy_magic_19_0.X.t45 GNDA 0.038267f
C1061 two_stage_opamp_dummy_magic_19_0.X.t30 GNDA 0.046467f
C1062 two_stage_opamp_dummy_magic_19_0.X.n33 GNDA 0.046467f
C1063 two_stage_opamp_dummy_magic_19_0.X.n34 GNDA 0.030067f
C1064 two_stage_opamp_dummy_magic_19_0.X.n35 GNDA 0.024942f
C1065 two_stage_opamp_dummy_magic_19_0.X.t34 GNDA 0.038267f
C1066 two_stage_opamp_dummy_magic_19_0.X.t49 GNDA 0.038267f
C1067 two_stage_opamp_dummy_magic_19_0.X.t26 GNDA 0.038267f
C1068 two_stage_opamp_dummy_magic_19_0.X.t40 GNDA 0.038267f
C1069 two_stage_opamp_dummy_magic_19_0.X.t53 GNDA 0.038267f
C1070 two_stage_opamp_dummy_magic_19_0.X.t36 GNDA 0.046467f
C1071 two_stage_opamp_dummy_magic_19_0.X.n36 GNDA 0.046467f
C1072 two_stage_opamp_dummy_magic_19_0.X.n37 GNDA 0.030067f
C1073 two_stage_opamp_dummy_magic_19_0.X.n38 GNDA 0.030067f
C1074 two_stage_opamp_dummy_magic_19_0.X.n39 GNDA 0.030067f
C1075 two_stage_opamp_dummy_magic_19_0.X.n40 GNDA 0.024942f
C1076 two_stage_opamp_dummy_magic_19_0.X.n41 GNDA 0.020627f
C1077 two_stage_opamp_dummy_magic_19_0.X.t41 GNDA 0.058767f
C1078 two_stage_opamp_dummy_magic_19_0.X.t27 GNDA 0.058767f
C1079 two_stage_opamp_dummy_magic_19_0.X.t32 GNDA 0.058767f
C1080 two_stage_opamp_dummy_magic_19_0.X.t47 GNDA 0.066809f
C1081 two_stage_opamp_dummy_magic_19_0.X.n42 GNDA 0.060293f
C1082 two_stage_opamp_dummy_magic_19_0.X.n43 GNDA 0.036901f
C1083 two_stage_opamp_dummy_magic_19_0.X.n44 GNDA 0.031775f
C1084 two_stage_opamp_dummy_magic_19_0.X.t54 GNDA 0.058767f
C1085 two_stage_opamp_dummy_magic_19_0.X.t37 GNDA 0.058767f
C1086 two_stage_opamp_dummy_magic_19_0.X.t44 GNDA 0.058767f
C1087 two_stage_opamp_dummy_magic_19_0.X.t29 GNDA 0.058767f
C1088 two_stage_opamp_dummy_magic_19_0.X.t42 GNDA 0.058767f
C1089 two_stage_opamp_dummy_magic_19_0.X.t25 GNDA 0.066809f
C1090 two_stage_opamp_dummy_magic_19_0.X.n45 GNDA 0.060293f
C1091 two_stage_opamp_dummy_magic_19_0.X.n46 GNDA 0.036901f
C1092 two_stage_opamp_dummy_magic_19_0.X.n47 GNDA 0.036901f
C1093 two_stage_opamp_dummy_magic_19_0.X.n48 GNDA 0.036901f
C1094 two_stage_opamp_dummy_magic_19_0.X.n49 GNDA 0.031775f
C1095 two_stage_opamp_dummy_magic_19_0.X.n50 GNDA 0.020627f
C1096 two_stage_opamp_dummy_magic_19_0.X.n51 GNDA 0.060216f
C1097 two_stage_opamp_dummy_magic_19_0.X.n52 GNDA 0.468971f
C1098 two_stage_opamp_dummy_magic_19_0.X.t46 GNDA 0.120268f
C1099 two_stage_opamp_dummy_magic_19_0.X.t33 GNDA 0.120268f
C1100 two_stage_opamp_dummy_magic_19_0.X.t50 GNDA 0.120268f
C1101 two_stage_opamp_dummy_magic_19_0.X.t28 GNDA 0.120268f
C1102 two_stage_opamp_dummy_magic_19_0.X.t43 GNDA 0.128094f
C1103 two_stage_opamp_dummy_magic_19_0.X.n53 GNDA 0.101509f
C1104 two_stage_opamp_dummy_magic_19_0.X.n54 GNDA 0.057401f
C1105 two_stage_opamp_dummy_magic_19_0.X.n55 GNDA 0.057401f
C1106 two_stage_opamp_dummy_magic_19_0.X.n56 GNDA 0.052276f
C1107 two_stage_opamp_dummy_magic_19_0.X.t31 GNDA 0.120268f
C1108 two_stage_opamp_dummy_magic_19_0.X.t39 GNDA 0.120268f
C1109 two_stage_opamp_dummy_magic_19_0.X.t51 GNDA 0.120268f
C1110 two_stage_opamp_dummy_magic_19_0.X.t35 GNDA 0.120268f
C1111 two_stage_opamp_dummy_magic_19_0.X.t48 GNDA 0.128094f
C1112 two_stage_opamp_dummy_magic_19_0.X.n57 GNDA 0.101509f
C1113 two_stage_opamp_dummy_magic_19_0.X.n58 GNDA 0.057401f
C1114 two_stage_opamp_dummy_magic_19_0.X.n59 GNDA 0.057401f
C1115 two_stage_opamp_dummy_magic_19_0.X.n60 GNDA 0.052276f
C1116 two_stage_opamp_dummy_magic_19_0.X.n61 GNDA 0.046271f
C1117 two_stage_opamp_dummy_magic_19_0.X.n62 GNDA 1.00986f
C1118 two_stage_opamp_dummy_magic_19_0.X.t17 GNDA 0.878237f
C1119 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t1 GNDA 0.345142f
C1120 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t79 GNDA 0.346293f
C1121 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t37 GNDA 0.186001f
C1122 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n0 GNDA 0.198613f
C1123 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t36 GNDA 0.345142f
C1124 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t123 GNDA 0.346293f
C1125 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t78 GNDA 0.186001f
C1126 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n1 GNDA 0.217197f
C1127 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t21 GNDA 0.345142f
C1128 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t99 GNDA 0.346293f
C1129 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t59 GNDA 0.186001f
C1130 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n2 GNDA 0.217197f
C1131 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t53 GNDA 0.345142f
C1132 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t130 GNDA 0.346293f
C1133 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t95 GNDA 0.186001f
C1134 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n3 GNDA 0.217197f
C1135 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t93 GNDA 0.345142f
C1136 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t41 GNDA 0.346293f
C1137 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t135 GNDA 0.364878f
C1138 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t31 GNDA 0.364878f
C1139 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t129 GNDA 0.186001f
C1140 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n4 GNDA 0.217197f
C1141 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t73 GNDA 0.345142f
C1142 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t96 GNDA 0.346293f
C1143 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t119 GNDA 0.364878f
C1144 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t12 GNDA 0.364878f
C1145 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t115 GNDA 0.186001f
C1146 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n5 GNDA 0.217197f
C1147 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t136 GNDA 0.346293f
C1148 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t101 GNDA 0.347548f
C1149 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t100 GNDA 0.346293f
C1150 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t60 GNDA 0.349008f
C1151 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t24 GNDA 0.379597f
C1152 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t125 GNDA 0.328964f
C1153 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t35 GNDA 0.346293f
C1154 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t0 GNDA 0.347548f
C1155 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t89 GNDA 0.328964f
C1156 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t4 GNDA 0.346293f
C1157 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t109 GNDA 0.347548f
C1158 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t25 GNDA 0.346293f
C1159 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t62 GNDA 0.347548f
C1160 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t38 GNDA 0.346293f
C1161 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t10 GNDA 0.347548f
C1162 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t67 GNDA 0.346293f
C1163 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t103 GNDA 0.347548f
C1164 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t80 GNDA 0.346293f
C1165 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t44 GNDA 0.347548f
C1166 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t29 GNDA 0.346293f
C1167 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t68 GNDA 0.347548f
C1168 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t46 GNDA 0.346293f
C1169 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t16 GNDA 0.347548f
C1170 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t72 GNDA 0.346293f
C1171 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t110 GNDA 0.347548f
C1172 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t88 GNDA 0.346293f
C1173 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t52 GNDA 0.347548f
C1174 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t114 GNDA 0.346293f
C1175 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t7 GNDA 0.347548f
C1176 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t126 GNDA 0.346293f
C1177 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t91 GNDA 0.347548f
C1178 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t75 GNDA 0.346293f
C1179 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t116 GNDA 0.347548f
C1180 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t92 GNDA 0.346293f
C1181 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t58 GNDA 0.347548f
C1182 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t120 GNDA 0.346293f
C1183 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t13 GNDA 0.347548f
C1184 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t128 GNDA 0.346293f
C1185 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t98 GNDA 0.347548f
C1186 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t19 GNDA 0.346293f
C1187 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t50 GNDA 0.347548f
C1188 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t30 GNDA 0.346293f
C1189 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t134 GNDA 0.347548f
C1190 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t54 GNDA 0.346293f
C1191 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t90 GNDA 0.347548f
C1192 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t74 GNDA 0.346293f
C1193 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t33 GNDA 0.347548f
C1194 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t22 GNDA 0.346293f
C1195 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t56 GNDA 0.347548f
C1196 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t34 GNDA 0.346293f
C1197 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t3 GNDA 0.347548f
C1198 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t61 GNDA 0.346293f
C1199 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t97 GNDA 0.347548f
C1200 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t77 GNDA 0.346293f
C1201 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t39 GNDA 0.347548f
C1202 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t102 GNDA 0.346293f
C1203 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t132 GNDA 0.347548f
C1204 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t122 GNDA 0.346293f
C1205 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t82 GNDA 0.347548f
C1206 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t107 GNDA 0.345142f
C1207 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t5 GNDA 0.346293f
C1208 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t71 GNDA 0.186001f
C1209 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n6 GNDA 0.198613f
C1210 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t137 GNDA 0.345142f
C1211 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t94 GNDA 0.346293f
C1212 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t108 GNDA 0.186001f
C1213 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n7 GNDA 0.217197f
C1214 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t48 GNDA 0.345142f
C1215 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t133 GNDA 0.346293f
C1216 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t18 GNDA 0.186001f
C1217 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n8 GNDA 0.217197f
C1218 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t83 GNDA 0.345142f
C1219 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t86 GNDA 0.346293f
C1220 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t49 GNDA 0.186001f
C1221 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n9 GNDA 0.217197f
C1222 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t124 GNDA 0.345142f
C1223 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t32 GNDA 0.346293f
C1224 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t85 GNDA 0.186001f
C1225 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n10 GNDA 0.217197f
C1226 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t28 GNDA 0.345142f
C1227 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t76 GNDA 0.346293f
C1228 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t131 GNDA 0.186001f
C1229 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n11 GNDA 0.217197f
C1230 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t66 GNDA 0.345142f
C1231 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t26 GNDA 0.346293f
C1232 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t27 GNDA 0.186001f
C1233 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n12 GNDA 0.217197f
C1234 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t118 GNDA 0.346293f
C1235 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t69 GNDA 0.186001f
C1236 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n13 GNDA 0.197462f
C1237 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t65 GNDA 0.346293f
C1238 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t104 GNDA 0.186001f
C1239 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n14 GNDA 0.197462f
C1240 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t81 GNDA 0.346293f
C1241 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t45 GNDA 0.347548f
C1242 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t6 GNDA 0.346293f
C1243 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t55 GNDA 0.347548f
C1244 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t111 GNDA 0.167416f
C1245 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n15 GNDA 0.215942f
C1246 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t15 GNDA 0.18485f
C1247 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n16 GNDA 0.234527f
C1248 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t42 GNDA 0.18485f
C1249 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n17 GNDA 0.251856f
C1250 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t8 GNDA 0.18485f
C1251 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n18 GNDA 0.251856f
C1252 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t112 GNDA 0.18485f
C1253 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n19 GNDA 0.251856f
C1254 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t2 GNDA 0.18485f
C1255 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n20 GNDA 0.251856f
C1256 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t105 GNDA 0.18485f
C1257 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n21 GNDA 0.251856f
C1258 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t63 GNDA 0.18485f
C1259 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n22 GNDA 0.251856f
C1260 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t23 GNDA 0.18485f
C1261 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n23 GNDA 0.251856f
C1262 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t57 GNDA 0.18485f
C1263 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n24 GNDA 0.251856f
C1264 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t20 GNDA 0.18485f
C1265 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n25 GNDA 0.251856f
C1266 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t121 GNDA 0.18485f
C1267 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n26 GNDA 0.251856f
C1268 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t14 GNDA 0.18485f
C1269 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n27 GNDA 0.251856f
C1270 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t117 GNDA 0.18485f
C1271 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n28 GNDA 0.251856f
C1272 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t70 GNDA 0.18485f
C1273 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n29 GNDA 0.251856f
C1274 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t106 GNDA 0.18485f
C1275 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n30 GNDA 0.251856f
C1276 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t64 GNDA 0.18485f
C1277 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n31 GNDA 0.234527f
C1278 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t40 GNDA 0.345142f
C1279 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t84 GNDA 0.167416f
C1280 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n32 GNDA 0.217197f
C1281 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t9 GNDA 0.345142f
C1282 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t51 GNDA 0.346293f
C1283 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t87 GNDA 0.364878f
C1284 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t43 GNDA 0.186001f
C1285 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n33 GNDA 0.217197f
C1286 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t113 GNDA 0.345142f
C1287 two_stage_opamp_dummy_magic_19_0.cap_res_Y.n34 GNDA 0.217197f
C1288 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t11 GNDA 0.186001f
C1289 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t47 GNDA 0.364878f
C1290 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t17 GNDA 0.364878f
C1291 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t127 GNDA 0.730561f
C1292 two_stage_opamp_dummy_magic_19_0.cap_res_Y.t138 GNDA 0.29977f
C1293 VOUT+.t13 GNDA 0.053328f
C1294 VOUT+.t1 GNDA 0.053328f
C1295 VOUT+.n0 GNDA 0.249232f
C1296 VOUT+.t17 GNDA 0.053328f
C1297 VOUT+.t11 GNDA 0.053328f
C1298 VOUT+.n1 GNDA 0.23402f
C1299 VOUT+.n2 GNDA 0.455316f
C1300 VOUT+.t2 GNDA 0.053328f
C1301 VOUT+.t14 GNDA 0.053328f
C1302 VOUT+.n3 GNDA 0.23402f
C1303 VOUT+.n4 GNDA 0.243524f
C1304 VOUT+.t10 GNDA 0.088718f
C1305 VOUT+.n5 GNDA 0.093346f
C1306 VOUT+.t4 GNDA 0.045709f
C1307 VOUT+.t3 GNDA 0.045709f
C1308 VOUT+.n6 GNDA 0.102649f
C1309 VOUT+.t15 GNDA 0.045709f
C1310 VOUT+.t7 GNDA 0.045709f
C1311 VOUT+.n7 GNDA 0.136517f
C1312 VOUT+.t12 GNDA 0.045709f
C1313 VOUT+.t8 GNDA 0.045709f
C1314 VOUT+.n8 GNDA 0.132953f
C1315 VOUT+.n9 GNDA 0.526637f
C1316 VOUT+.t0 GNDA 0.045709f
C1317 VOUT+.t6 GNDA 0.045709f
C1318 VOUT+.n10 GNDA 0.132953f
C1319 VOUT+.n11 GNDA 0.267766f
C1320 VOUT+.t9 GNDA 0.045709f
C1321 VOUT+.t18 GNDA 0.045709f
C1322 VOUT+.n12 GNDA 0.132953f
C1323 VOUT+.n13 GNDA 0.267766f
C1324 VOUT+.t5 GNDA 0.045709f
C1325 VOUT+.t16 GNDA 0.045709f
C1326 VOUT+.n14 GNDA 0.136517f
C1327 VOUT+.n15 GNDA 0.281725f
C1328 VOUT+.n16 GNDA 0.356093f
C1329 VOUT+.t45 GNDA 0.30473f
C1330 VOUT+.t150 GNDA 0.30992f
C1331 VOUT+.t101 GNDA 0.30473f
C1332 VOUT+.n17 GNDA 0.204311f
C1333 VOUT+.n18 GNDA 0.133319f
C1334 VOUT+.t91 GNDA 0.30927f
C1335 VOUT+.t38 GNDA 0.30927f
C1336 VOUT+.t130 GNDA 0.30927f
C1337 VOUT+.t90 GNDA 0.30927f
C1338 VOUT+.t80 GNDA 0.30927f
C1339 VOUT+.t128 GNDA 0.30927f
C1340 VOUT+.t124 GNDA 0.30927f
C1341 VOUT+.t32 GNDA 0.30927f
C1342 VOUT+.t70 GNDA 0.30927f
C1343 VOUT+.t73 GNDA 0.30927f
C1344 VOUT+.t23 GNDA 0.30927f
C1345 VOUT+.t108 GNDA 0.30927f
C1346 VOUT+.t62 GNDA 0.30927f
C1347 VOUT+.t19 GNDA 0.30927f
C1348 VOUT+.t151 GNDA 0.30927f
C1349 VOUT+.t49 GNDA 0.30927f
C1350 VOUT+.t85 GNDA 0.30473f
C1351 VOUT+.n19 GNDA 0.33374f
C1352 VOUT+.t48 GNDA 0.30473f
C1353 VOUT+.n20 GNDA 0.390877f
C1354 VOUT+.t138 GNDA 0.30473f
C1355 VOUT+.n21 GNDA 0.390877f
C1356 VOUT+.t107 GNDA 0.30473f
C1357 VOUT+.n22 GNDA 0.390877f
C1358 VOUT+.t71 GNDA 0.30473f
C1359 VOUT+.n23 GNDA 0.390877f
C1360 VOUT+.t25 GNDA 0.30473f
C1361 VOUT+.n24 GNDA 0.390877f
C1362 VOUT+.t129 GNDA 0.30473f
C1363 VOUT+.n25 GNDA 0.390877f
C1364 VOUT+.t87 GNDA 0.30473f
C1365 VOUT+.n26 GNDA 0.262098f
C1366 VOUT+.t52 GNDA 0.30473f
C1367 VOUT+.n27 GNDA 0.262098f
C1368 VOUT+.t141 GNDA 0.30473f
C1369 VOUT+.t75 GNDA 0.30992f
C1370 VOUT+.t111 GNDA 0.30473f
C1371 VOUT+.n28 GNDA 0.204311f
C1372 VOUT+.n29 GNDA 0.247593f
C1373 VOUT+.t54 GNDA 0.30992f
C1374 VOUT+.t24 GNDA 0.30473f
C1375 VOUT+.n30 GNDA 0.204311f
C1376 VOUT+.t114 GNDA 0.30473f
C1377 VOUT+.t34 GNDA 0.30992f
C1378 VOUT+.t74 GNDA 0.30473f
C1379 VOUT+.n31 GNDA 0.204311f
C1380 VOUT+.n32 GNDA 0.247593f
C1381 VOUT+.t95 GNDA 0.30992f
C1382 VOUT+.t59 GNDA 0.30473f
C1383 VOUT+.n33 GNDA 0.204311f
C1384 VOUT+.t148 GNDA 0.30473f
C1385 VOUT+.t79 GNDA 0.30992f
C1386 VOUT+.t117 GNDA 0.30473f
C1387 VOUT+.n34 GNDA 0.204311f
C1388 VOUT+.n35 GNDA 0.247593f
C1389 VOUT+.t134 GNDA 0.30992f
C1390 VOUT+.t100 GNDA 0.30473f
C1391 VOUT+.n36 GNDA 0.204311f
C1392 VOUT+.t44 GNDA 0.30473f
C1393 VOUT+.t122 GNDA 0.30992f
C1394 VOUT+.t153 GNDA 0.30473f
C1395 VOUT+.n37 GNDA 0.204311f
C1396 VOUT+.n38 GNDA 0.247593f
C1397 VOUT+.t102 GNDA 0.30992f
C1398 VOUT+.t66 GNDA 0.30473f
C1399 VOUT+.n39 GNDA 0.204311f
C1400 VOUT+.t154 GNDA 0.30473f
C1401 VOUT+.t82 GNDA 0.30992f
C1402 VOUT+.t123 GNDA 0.30473f
C1403 VOUT+.n40 GNDA 0.204311f
C1404 VOUT+.n41 GNDA 0.247593f
C1405 VOUT+.t137 GNDA 0.30992f
C1406 VOUT+.t106 GNDA 0.30473f
C1407 VOUT+.n42 GNDA 0.204311f
C1408 VOUT+.t51 GNDA 0.30473f
C1409 VOUT+.t126 GNDA 0.30992f
C1410 VOUT+.t22 GNDA 0.30473f
C1411 VOUT+.n43 GNDA 0.204311f
C1412 VOUT+.n44 GNDA 0.247593f
C1413 VOUT+.t132 GNDA 0.30473f
C1414 VOUT+.t56 GNDA 0.30992f
C1415 VOUT+.t96 GNDA 0.30473f
C1416 VOUT+.n45 GNDA 0.204311f
C1417 VOUT+.n46 GNDA 0.133319f
C1418 VOUT+.t116 GNDA 0.30927f
C1419 VOUT+.t105 GNDA 0.30992f
C1420 VOUT+.t69 GNDA 0.30473f
C1421 VOUT+.n47 GNDA 0.19955f
C1422 VOUT+.t147 GNDA 0.30927f
C1423 VOUT+.t29 GNDA 0.30992f
C1424 VOUT+.t139 GNDA 0.30473f
C1425 VOUT+.n48 GNDA 0.204311f
C1426 VOUT+.t109 GNDA 0.30473f
C1427 VOUT+.n49 GNDA 0.128558f
C1428 VOUT+.t43 GNDA 0.30927f
C1429 VOUT+.t60 GNDA 0.30992f
C1430 VOUT+.t37 GNDA 0.30473f
C1431 VOUT+.n50 GNDA 0.204311f
C1432 VOUT+.t144 GNDA 0.30473f
C1433 VOUT+.n51 GNDA 0.128558f
C1434 VOUT+.t83 GNDA 0.30927f
C1435 VOUT+.t115 GNDA 0.30992f
C1436 VOUT+.t21 GNDA 0.30473f
C1437 VOUT+.n52 GNDA 0.204311f
C1438 VOUT+.t125 GNDA 0.30473f
C1439 VOUT+.n53 GNDA 0.128558f
C1440 VOUT+.t63 GNDA 0.30927f
C1441 VOUT+.t26 GNDA 0.30927f
C1442 VOUT+.t103 GNDA 0.30927f
C1443 VOUT+.t57 GNDA 0.309525f
C1444 VOUT+.t135 GNDA 0.30927f
C1445 VOUT+.t33 GNDA 0.309525f
C1446 VOUT+.t120 GNDA 0.30927f
C1447 VOUT+.t77 GNDA 0.309525f
C1448 VOUT+.t155 GNDA 0.30927f
C1449 VOUT+.t119 GNDA 0.30473f
C1450 VOUT+.n54 GNDA 0.337294f
C1451 VOUT+.t78 GNDA 0.30473f
C1452 VOUT+.n55 GNDA 0.394431f
C1453 VOUT+.t97 GNDA 0.30473f
C1454 VOUT+.n56 GNDA 0.394431f
C1455 VOUT+.t61 GNDA 0.30473f
C1456 VOUT+.n57 GNDA 0.390877f
C1457 VOUT+.t27 GNDA 0.30473f
C1458 VOUT+.n58 GNDA 0.323996f
C1459 VOUT+.t41 GNDA 0.30473f
C1460 VOUT+.n59 GNDA 0.323996f
C1461 VOUT+.t145 GNDA 0.30473f
C1462 VOUT+.n60 GNDA 0.323996f
C1463 VOUT+.t113 GNDA 0.30473f
C1464 VOUT+.n61 GNDA 0.323996f
C1465 VOUT+.t72 GNDA 0.30473f
C1466 VOUT+.n62 GNDA 0.262098f
C1467 VOUT+.t92 GNDA 0.30473f
C1468 VOUT+.t20 GNDA 0.30992f
C1469 VOUT+.t55 GNDA 0.30473f
C1470 VOUT+.n63 GNDA 0.204311f
C1471 VOUT+.n64 GNDA 0.247593f
C1472 VOUT+.t31 GNDA 0.30992f
C1473 VOUT+.t50 GNDA 0.30473f
C1474 VOUT+.t121 GNDA 0.30992f
C1475 VOUT+.t156 GNDA 0.30473f
C1476 VOUT+.n65 GNDA 0.204311f
C1477 VOUT+.n66 GNDA 0.318585f
C1478 VOUT+.t67 GNDA 0.30992f
C1479 VOUT+.t86 GNDA 0.30473f
C1480 VOUT+.t152 GNDA 0.30992f
C1481 VOUT+.t47 GNDA 0.30473f
C1482 VOUT+.n67 GNDA 0.204311f
C1483 VOUT+.n68 GNDA 0.318585f
C1484 VOUT+.t131 GNDA 0.30992f
C1485 VOUT+.t94 GNDA 0.30473f
C1486 VOUT+.n69 GNDA 0.204311f
C1487 VOUT+.t39 GNDA 0.30473f
C1488 VOUT+.t118 GNDA 0.30992f
C1489 VOUT+.t146 GNDA 0.30473f
C1490 VOUT+.n70 GNDA 0.204311f
C1491 VOUT+.n71 GNDA 0.247593f
C1492 VOUT+.t89 GNDA 0.30992f
C1493 VOUT+.t53 GNDA 0.30473f
C1494 VOUT+.n72 GNDA 0.204311f
C1495 VOUT+.t142 GNDA 0.30473f
C1496 VOUT+.t76 GNDA 0.30992f
C1497 VOUT+.t112 GNDA 0.30473f
C1498 VOUT+.n73 GNDA 0.204311f
C1499 VOUT+.n74 GNDA 0.247593f
C1500 VOUT+.t127 GNDA 0.30992f
C1501 VOUT+.t88 GNDA 0.30473f
C1502 VOUT+.n75 GNDA 0.204311f
C1503 VOUT+.t35 GNDA 0.30473f
C1504 VOUT+.t110 GNDA 0.30992f
C1505 VOUT+.t140 GNDA 0.30473f
C1506 VOUT+.n76 GNDA 0.204311f
C1507 VOUT+.n77 GNDA 0.247593f
C1508 VOUT+.t84 GNDA 0.30992f
C1509 VOUT+.t46 GNDA 0.30473f
C1510 VOUT+.n78 GNDA 0.204311f
C1511 VOUT+.t136 GNDA 0.30473f
C1512 VOUT+.t68 GNDA 0.30992f
C1513 VOUT+.t104 GNDA 0.30473f
C1514 VOUT+.n79 GNDA 0.204311f
C1515 VOUT+.n80 GNDA 0.247593f
C1516 VOUT+.t42 GNDA 0.30992f
C1517 VOUT+.t149 GNDA 0.30473f
C1518 VOUT+.n81 GNDA 0.204311f
C1519 VOUT+.t99 GNDA 0.30473f
C1520 VOUT+.t30 GNDA 0.30992f
C1521 VOUT+.t65 GNDA 0.30473f
C1522 VOUT+.n82 GNDA 0.204311f
C1523 VOUT+.n83 GNDA 0.247593f
C1524 VOUT+.t81 GNDA 0.30992f
C1525 VOUT+.t40 GNDA 0.30473f
C1526 VOUT+.n84 GNDA 0.204311f
C1527 VOUT+.t133 GNDA 0.30473f
C1528 VOUT+.t64 GNDA 0.30992f
C1529 VOUT+.t98 GNDA 0.30473f
C1530 VOUT+.n85 GNDA 0.204311f
C1531 VOUT+.n86 GNDA 0.247593f
C1532 VOUT+.t28 GNDA 0.30992f
C1533 VOUT+.t58 GNDA 0.30473f
C1534 VOUT+.n87 GNDA 0.204311f
C1535 VOUT+.t93 GNDA 0.30473f
C1536 VOUT+.n88 GNDA 0.247593f
C1537 VOUT+.t143 GNDA 0.30473f
C1538 VOUT+.n89 GNDA 0.133319f
C1539 VOUT+.t36 GNDA 0.30473f
C1540 VOUT+.n90 GNDA 0.19441f
C1541 VOUT+.n91 GNDA 0.226601f
C1542 two_stage_opamp_dummy_magic_19_0.V_source.t27 GNDA 0.02347f
C1543 two_stage_opamp_dummy_magic_19_0.V_source.t19 GNDA 0.087069f
C1544 two_stage_opamp_dummy_magic_19_0.V_source.t38 GNDA 0.02347f
C1545 two_stage_opamp_dummy_magic_19_0.V_source.t17 GNDA 0.02347f
C1546 two_stage_opamp_dummy_magic_19_0.V_source.n0 GNDA 0.070305f
C1547 two_stage_opamp_dummy_magic_19_0.V_source.n1 GNDA 0.412007f
C1548 two_stage_opamp_dummy_magic_19_0.V_source.t16 GNDA 0.014082f
C1549 two_stage_opamp_dummy_magic_19_0.V_source.t4 GNDA 0.014082f
C1550 two_stage_opamp_dummy_magic_19_0.V_source.n2 GNDA 0.031237f
C1551 two_stage_opamp_dummy_magic_19_0.V_source.t0 GNDA 0.014082f
C1552 two_stage_opamp_dummy_magic_19_0.V_source.t13 GNDA 0.014082f
C1553 two_stage_opamp_dummy_magic_19_0.V_source.n3 GNDA 0.04039f
C1554 two_stage_opamp_dummy_magic_19_0.V_source.t40 GNDA 0.014082f
C1555 two_stage_opamp_dummy_magic_19_0.V_source.t12 GNDA 0.014082f
C1556 two_stage_opamp_dummy_magic_19_0.V_source.n4 GNDA 0.039262f
C1557 two_stage_opamp_dummy_magic_19_0.V_source.n5 GNDA 0.225457f
C1558 two_stage_opamp_dummy_magic_19_0.V_source.t5 GNDA 0.014082f
C1559 two_stage_opamp_dummy_magic_19_0.V_source.t14 GNDA 0.014082f
C1560 two_stage_opamp_dummy_magic_19_0.V_source.n6 GNDA 0.039262f
C1561 two_stage_opamp_dummy_magic_19_0.V_source.n7 GNDA 0.116578f
C1562 two_stage_opamp_dummy_magic_19_0.V_source.t8 GNDA 0.014082f
C1563 two_stage_opamp_dummy_magic_19_0.V_source.t11 GNDA 0.014082f
C1564 two_stage_opamp_dummy_magic_19_0.V_source.n8 GNDA 0.039262f
C1565 two_stage_opamp_dummy_magic_19_0.V_source.n9 GNDA 0.116578f
C1566 two_stage_opamp_dummy_magic_19_0.V_source.t18 GNDA 0.014082f
C1567 two_stage_opamp_dummy_magic_19_0.V_source.t2 GNDA 0.014082f
C1568 two_stage_opamp_dummy_magic_19_0.V_source.n10 GNDA 0.04039f
C1569 two_stage_opamp_dummy_magic_19_0.V_source.t3 GNDA 0.014082f
C1570 two_stage_opamp_dummy_magic_19_0.V_source.t15 GNDA 0.014082f
C1571 two_stage_opamp_dummy_magic_19_0.V_source.n11 GNDA 0.039262f
C1572 two_stage_opamp_dummy_magic_19_0.V_source.n12 GNDA 0.225457f
C1573 two_stage_opamp_dummy_magic_19_0.V_source.t1 GNDA 0.014082f
C1574 two_stage_opamp_dummy_magic_19_0.V_source.t9 GNDA 0.014082f
C1575 two_stage_opamp_dummy_magic_19_0.V_source.n13 GNDA 0.039262f
C1576 two_stage_opamp_dummy_magic_19_0.V_source.n14 GNDA 0.116578f
C1577 two_stage_opamp_dummy_magic_19_0.V_source.t10 GNDA 0.014082f
C1578 two_stage_opamp_dummy_magic_19_0.V_source.t7 GNDA 0.014082f
C1579 two_stage_opamp_dummy_magic_19_0.V_source.n15 GNDA 0.039262f
C1580 two_stage_opamp_dummy_magic_19_0.V_source.n16 GNDA 0.116578f
C1581 two_stage_opamp_dummy_magic_19_0.V_source.t6 GNDA 0.014082f
C1582 two_stage_opamp_dummy_magic_19_0.V_source.t39 GNDA 0.014082f
C1583 two_stage_opamp_dummy_magic_19_0.V_source.n17 GNDA 0.039262f
C1584 two_stage_opamp_dummy_magic_19_0.V_source.n18 GNDA 0.1776f
C1585 two_stage_opamp_dummy_magic_19_0.V_source.n19 GNDA 0.089186f
C1586 two_stage_opamp_dummy_magic_19_0.V_source.n20 GNDA 0.172952f
C1587 two_stage_opamp_dummy_magic_19_0.V_source.t21 GNDA 0.02347f
C1588 two_stage_opamp_dummy_magic_19_0.V_source.t33 GNDA 0.02347f
C1589 two_stage_opamp_dummy_magic_19_0.V_source.n21 GNDA 0.052352f
C1590 two_stage_opamp_dummy_magic_19_0.V_source.n22 GNDA 0.225532f
C1591 two_stage_opamp_dummy_magic_19_0.V_source.n23 GNDA 0.028164f
C1592 two_stage_opamp_dummy_magic_19_0.V_source.t22 GNDA 0.02347f
C1593 two_stage_opamp_dummy_magic_19_0.V_source.t29 GNDA 0.02347f
C1594 two_stage_opamp_dummy_magic_19_0.V_source.n24 GNDA 0.070305f
C1595 two_stage_opamp_dummy_magic_19_0.V_source.n25 GNDA 0.159231f
C1596 two_stage_opamp_dummy_magic_19_0.V_source.t26 GNDA 0.02347f
C1597 two_stage_opamp_dummy_magic_19_0.V_source.t32 GNDA 0.02347f
C1598 two_stage_opamp_dummy_magic_19_0.V_source.n26 GNDA 0.072561f
C1599 two_stage_opamp_dummy_magic_19_0.V_source.t28 GNDA 0.02347f
C1600 two_stage_opamp_dummy_magic_19_0.V_source.t36 GNDA 0.02347f
C1601 two_stage_opamp_dummy_magic_19_0.V_source.n27 GNDA 0.070305f
C1602 two_stage_opamp_dummy_magic_19_0.V_source.n28 GNDA 0.309635f
C1603 two_stage_opamp_dummy_magic_19_0.V_source.t30 GNDA 0.02347f
C1604 two_stage_opamp_dummy_magic_19_0.V_source.t20 GNDA 0.02347f
C1605 two_stage_opamp_dummy_magic_19_0.V_source.n29 GNDA 0.070305f
C1606 two_stage_opamp_dummy_magic_19_0.V_source.n30 GNDA 0.159231f
C1607 two_stage_opamp_dummy_magic_19_0.V_source.t34 GNDA 0.02347f
C1608 two_stage_opamp_dummy_magic_19_0.V_source.t24 GNDA 0.02347f
C1609 two_stage_opamp_dummy_magic_19_0.V_source.n31 GNDA 0.070305f
C1610 two_stage_opamp_dummy_magic_19_0.V_source.n32 GNDA 0.159231f
C1611 two_stage_opamp_dummy_magic_19_0.V_source.t31 GNDA 0.02347f
C1612 two_stage_opamp_dummy_magic_19_0.V_source.t23 GNDA 0.02347f
C1613 two_stage_opamp_dummy_magic_19_0.V_source.n33 GNDA 0.070305f
C1614 two_stage_opamp_dummy_magic_19_0.V_source.n34 GNDA 0.159231f
C1615 two_stage_opamp_dummy_magic_19_0.V_source.t35 GNDA 0.02347f
C1616 two_stage_opamp_dummy_magic_19_0.V_source.t25 GNDA 0.02347f
C1617 two_stage_opamp_dummy_magic_19_0.V_source.n35 GNDA 0.070305f
C1618 two_stage_opamp_dummy_magic_19_0.V_source.n36 GNDA 0.159231f
C1619 two_stage_opamp_dummy_magic_19_0.V_source.n37 GNDA 0.159231f
C1620 two_stage_opamp_dummy_magic_19_0.V_source.n38 GNDA 0.070305f
C1621 two_stage_opamp_dummy_magic_19_0.V_source.t37 GNDA 0.02347f
C1622 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t4 GNDA 0.013327f
C1623 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t5 GNDA 0.013327f
C1624 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n0 GNDA 0.069778f
C1625 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t6 GNDA 0.013327f
C1626 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t0 GNDA 0.013327f
C1627 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n1 GNDA 0.026655f
C1628 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n2 GNDA 0.109409f
C1629 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n3 GNDA 0.0225f
C1630 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n4 GNDA 0.037659f
C1631 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n5 GNDA 0.197494f
C1632 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t20 GNDA 0.017742f
C1633 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t13 GNDA 0.020708f
C1634 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n6 GNDA 0.01765f
C1635 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t9 GNDA 0.017742f
C1636 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t18 GNDA 0.017742f
C1637 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t26 GNDA 0.017742f
C1638 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t15 GNDA 0.017742f
C1639 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t22 GNDA 0.017742f
C1640 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t11 GNDA 0.017742f
C1641 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t23 GNDA 0.017742f
C1642 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t14 GNDA 0.017742f
C1643 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t21 GNDA 0.017742f
C1644 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t10 GNDA 0.017742f
C1645 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t19 GNDA 0.017742f
C1646 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t8 GNDA 0.017742f
C1647 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t17 GNDA 0.017742f
C1648 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t24 GNDA 0.017742f
C1649 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t12 GNDA 0.017742f
C1650 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t25 GNDA 0.020708f
C1651 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n7 GNDA 0.019524f
C1652 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n8 GNDA 0.012245f
C1653 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n9 GNDA 0.012245f
C1654 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n10 GNDA 0.012245f
C1655 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n11 GNDA 0.012245f
C1656 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n12 GNDA 0.012245f
C1657 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n13 GNDA 0.012245f
C1658 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n14 GNDA 0.012245f
C1659 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n15 GNDA 0.012245f
C1660 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n16 GNDA 0.012245f
C1661 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n17 GNDA 0.012245f
C1662 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n18 GNDA 0.012245f
C1663 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n19 GNDA 0.012245f
C1664 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n20 GNDA 0.012245f
C1665 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n21 GNDA 0.01037f
C1666 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n22 GNDA 0.017109f
C1667 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t16 GNDA 0.018743f
C1668 two_stage_opamp_dummy_magic_19_0.V_tail_gate.t27 GNDA 0.018743f
C1669 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n23 GNDA 0.025948f
C1670 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n24 GNDA 0.177369f
C1671 two_stage_opamp_dummy_magic_19_0.V_tail_gate.n25 GNDA 0.428127f
C1672 bgr_9_0.TAIL_CUR_MIR_BIAS GNDA 0.525154f
C1673 two_stage_opamp_dummy_magic_19_0.cap_res_X.t127 GNDA 0.346251f
C1674 two_stage_opamp_dummy_magic_19_0.cap_res_X.t104 GNDA 0.347506f
C1675 two_stage_opamp_dummy_magic_19_0.cap_res_X.t88 GNDA 0.346251f
C1676 two_stage_opamp_dummy_magic_19_0.cap_res_X.t70 GNDA 0.348966f
C1677 two_stage_opamp_dummy_magic_19_0.cap_res_X.t102 GNDA 0.379551f
C1678 two_stage_opamp_dummy_magic_19_0.cap_res_X.t31 GNDA 0.346251f
C1679 two_stage_opamp_dummy_magic_19_0.cap_res_X.t4 GNDA 0.347506f
C1680 two_stage_opamp_dummy_magic_19_0.cap_res_X.t83 GNDA 0.328924f
C1681 two_stage_opamp_dummy_magic_19_0.cap_res_X.t133 GNDA 0.346251f
C1682 two_stage_opamp_dummy_magic_19_0.cap_res_X.t109 GNDA 0.347506f
C1683 two_stage_opamp_dummy_magic_19_0.cap_res_X.t47 GNDA 0.328924f
C1684 two_stage_opamp_dummy_magic_19_0.cap_res_X.t80 GNDA 0.346251f
C1685 two_stage_opamp_dummy_magic_19_0.cap_res_X.t129 GNDA 0.347506f
C1686 two_stage_opamp_dummy_magic_19_0.cap_res_X.t112 GNDA 0.346251f
C1687 two_stage_opamp_dummy_magic_19_0.cap_res_X.t59 GNDA 0.347506f
C1688 two_stage_opamp_dummy_magic_19_0.cap_res_X.t119 GNDA 0.346251f
C1689 two_stage_opamp_dummy_magic_19_0.cap_res_X.t33 GNDA 0.347506f
C1690 two_stage_opamp_dummy_magic_19_0.cap_res_X.t13 GNDA 0.346251f
C1691 two_stage_opamp_dummy_magic_19_0.cap_res_X.t99 GNDA 0.347506f
C1692 two_stage_opamp_dummy_magic_19_0.cap_res_X.t86 GNDA 0.346251f
C1693 two_stage_opamp_dummy_magic_19_0.cap_res_X.t136 GNDA 0.347506f
C1694 two_stage_opamp_dummy_magic_19_0.cap_res_X.t117 GNDA 0.346251f
C1695 two_stage_opamp_dummy_magic_19_0.cap_res_X.t69 GNDA 0.347506f
C1696 two_stage_opamp_dummy_magic_19_0.cap_res_X.t124 GNDA 0.346251f
C1697 two_stage_opamp_dummy_magic_19_0.cap_res_X.t38 GNDA 0.347506f
C1698 two_stage_opamp_dummy_magic_19_0.cap_res_X.t18 GNDA 0.346251f
C1699 two_stage_opamp_dummy_magic_19_0.cap_res_X.t103 GNDA 0.347506f
C1700 two_stage_opamp_dummy_magic_19_0.cap_res_X.t25 GNDA 0.346251f
C1701 two_stage_opamp_dummy_magic_19_0.cap_res_X.t77 GNDA 0.347506f
C1702 two_stage_opamp_dummy_magic_19_0.cap_res_X.t55 GNDA 0.346251f
C1703 two_stage_opamp_dummy_magic_19_0.cap_res_X.t3 GNDA 0.347506f
C1704 two_stage_opamp_dummy_magic_19_0.cap_res_X.t128 GNDA 0.346251f
C1705 two_stage_opamp_dummy_magic_19_0.cap_res_X.t39 GNDA 0.347506f
C1706 two_stage_opamp_dummy_magic_19_0.cap_res_X.t23 GNDA 0.346251f
C1707 two_stage_opamp_dummy_magic_19_0.cap_res_X.t110 GNDA 0.347506f
C1708 two_stage_opamp_dummy_magic_19_0.cap_res_X.t32 GNDA 0.346251f
C1709 two_stage_opamp_dummy_magic_19_0.cap_res_X.t81 GNDA 0.347506f
C1710 two_stage_opamp_dummy_magic_19_0.cap_res_X.t60 GNDA 0.346251f
C1711 two_stage_opamp_dummy_magic_19_0.cap_res_X.t11 GNDA 0.347506f
C1712 two_stage_opamp_dummy_magic_19_0.cap_res_X.t71 GNDA 0.346251f
C1713 two_stage_opamp_dummy_magic_19_0.cap_res_X.t122 GNDA 0.347506f
C1714 two_stage_opamp_dummy_magic_19_0.cap_res_X.t101 GNDA 0.346251f
C1715 two_stage_opamp_dummy_magic_19_0.cap_res_X.t50 GNDA 0.347506f
C1716 two_stage_opamp_dummy_magic_19_0.cap_res_X.t107 GNDA 0.346251f
C1717 two_stage_opamp_dummy_magic_19_0.cap_res_X.t21 GNDA 0.347506f
C1718 two_stage_opamp_dummy_magic_19_0.cap_res_X.t137 GNDA 0.346251f
C1719 two_stage_opamp_dummy_magic_19_0.cap_res_X.t89 GNDA 0.347506f
C1720 two_stage_opamp_dummy_magic_19_0.cap_res_X.t76 GNDA 0.346251f
C1721 two_stage_opamp_dummy_magic_19_0.cap_res_X.t126 GNDA 0.347506f
C1722 two_stage_opamp_dummy_magic_19_0.cap_res_X.t105 GNDA 0.346251f
C1723 two_stage_opamp_dummy_magic_19_0.cap_res_X.t53 GNDA 0.347506f
C1724 two_stage_opamp_dummy_magic_19_0.cap_res_X.t115 GNDA 0.346251f
C1725 two_stage_opamp_dummy_magic_19_0.cap_res_X.t27 GNDA 0.347506f
C1726 two_stage_opamp_dummy_magic_19_0.cap_res_X.t5 GNDA 0.346251f
C1727 two_stage_opamp_dummy_magic_19_0.cap_res_X.t93 GNDA 0.347506f
C1728 two_stage_opamp_dummy_magic_19_0.cap_res_X.t16 GNDA 0.346251f
C1729 two_stage_opamp_dummy_magic_19_0.cap_res_X.t67 GNDA 0.347506f
C1730 two_stage_opamp_dummy_magic_19_0.cap_res_X.t45 GNDA 0.346251f
C1731 two_stage_opamp_dummy_magic_19_0.cap_res_X.t135 GNDA 0.347506f
C1732 two_stage_opamp_dummy_magic_19_0.cap_res_X.t120 GNDA 0.346251f
C1733 two_stage_opamp_dummy_magic_19_0.cap_res_X.t34 GNDA 0.347506f
C1734 two_stage_opamp_dummy_magic_19_0.cap_res_X.t43 GNDA 0.3451f
C1735 two_stage_opamp_dummy_magic_19_0.cap_res_X.t85 GNDA 0.346251f
C1736 two_stage_opamp_dummy_magic_19_0.cap_res_X.t8 GNDA 0.185978f
C1737 two_stage_opamp_dummy_magic_19_0.cap_res_X.n0 GNDA 0.198589f
C1738 two_stage_opamp_dummy_magic_19_0.cap_res_X.t132 GNDA 0.3451f
C1739 two_stage_opamp_dummy_magic_19_0.cap_res_X.t42 GNDA 0.346251f
C1740 two_stage_opamp_dummy_magic_19_0.cap_res_X.t96 GNDA 0.185978f
C1741 two_stage_opamp_dummy_magic_19_0.cap_res_X.n1 GNDA 0.217171f
C1742 two_stage_opamp_dummy_magic_19_0.cap_res_X.t94 GNDA 0.3451f
C1743 two_stage_opamp_dummy_magic_19_0.cap_res_X.t91 GNDA 0.346251f
C1744 two_stage_opamp_dummy_magic_19_0.cap_res_X.t63 GNDA 0.185978f
C1745 two_stage_opamp_dummy_magic_19_0.cap_res_X.n2 GNDA 0.217171f
C1746 two_stage_opamp_dummy_magic_19_0.cap_res_X.t61 GNDA 0.3451f
C1747 two_stage_opamp_dummy_magic_19_0.cap_res_X.t2 GNDA 0.346251f
C1748 two_stage_opamp_dummy_magic_19_0.cap_res_X.t29 GNDA 0.185978f
C1749 two_stage_opamp_dummy_magic_19_0.cap_res_X.n3 GNDA 0.217171f
C1750 two_stage_opamp_dummy_magic_19_0.cap_res_X.t30 GNDA 0.3451f
C1751 two_stage_opamp_dummy_magic_19_0.cap_res_X.t51 GNDA 0.346251f
C1752 two_stage_opamp_dummy_magic_19_0.cap_res_X.t131 GNDA 0.185978f
C1753 two_stage_opamp_dummy_magic_19_0.cap_res_X.n4 GNDA 0.217171f
C1754 two_stage_opamp_dummy_magic_19_0.cap_res_X.t118 GNDA 0.3451f
C1755 two_stage_opamp_dummy_magic_19_0.cap_res_X.t15 GNDA 0.346251f
C1756 two_stage_opamp_dummy_magic_19_0.cap_res_X.t84 GNDA 0.185978f
C1757 two_stage_opamp_dummy_magic_19_0.cap_res_X.n5 GNDA 0.217171f
C1758 two_stage_opamp_dummy_magic_19_0.cap_res_X.t82 GNDA 0.3451f
C1759 two_stage_opamp_dummy_magic_19_0.cap_res_X.t64 GNDA 0.346251f
C1760 two_stage_opamp_dummy_magic_19_0.cap_res_X.t46 GNDA 0.185978f
C1761 two_stage_opamp_dummy_magic_19_0.cap_res_X.n6 GNDA 0.217171f
C1762 two_stage_opamp_dummy_magic_19_0.cap_res_X.t114 GNDA 0.346251f
C1763 two_stage_opamp_dummy_magic_19_0.cap_res_X.t14 GNDA 0.185978f
C1764 two_stage_opamp_dummy_magic_19_0.cap_res_X.n7 GNDA 0.197438f
C1765 two_stage_opamp_dummy_magic_19_0.cap_res_X.t74 GNDA 0.346251f
C1766 two_stage_opamp_dummy_magic_19_0.cap_res_X.t100 GNDA 0.185978f
C1767 two_stage_opamp_dummy_magic_19_0.cap_res_X.n8 GNDA 0.197438f
C1768 two_stage_opamp_dummy_magic_19_0.cap_res_X.t130 GNDA 0.346251f
C1769 two_stage_opamp_dummy_magic_19_0.cap_res_X.t37 GNDA 0.347506f
C1770 two_stage_opamp_dummy_magic_19_0.cap_res_X.t123 GNDA 0.167396f
C1771 two_stage_opamp_dummy_magic_19_0.cap_res_X.n9 GNDA 0.215916f
C1772 two_stage_opamp_dummy_magic_19_0.cap_res_X.t66 GNDA 0.184828f
C1773 two_stage_opamp_dummy_magic_19_0.cap_res_X.n10 GNDA 0.234498f
C1774 two_stage_opamp_dummy_magic_19_0.cap_res_X.t97 GNDA 0.184828f
C1775 two_stage_opamp_dummy_magic_19_0.cap_res_X.n11 GNDA 0.251826f
C1776 two_stage_opamp_dummy_magic_19_0.cap_res_X.t58 GNDA 0.184828f
C1777 two_stage_opamp_dummy_magic_19_0.cap_res_X.n12 GNDA 0.251826f
C1778 two_stage_opamp_dummy_magic_19_0.cap_res_X.t22 GNDA 0.184828f
C1779 two_stage_opamp_dummy_magic_19_0.cap_res_X.n13 GNDA 0.251826f
C1780 two_stage_opamp_dummy_magic_19_0.cap_res_X.t54 GNDA 0.184828f
C1781 two_stage_opamp_dummy_magic_19_0.cap_res_X.n14 GNDA 0.251826f
C1782 two_stage_opamp_dummy_magic_19_0.cap_res_X.t17 GNDA 0.184828f
C1783 two_stage_opamp_dummy_magic_19_0.cap_res_X.n15 GNDA 0.251826f
C1784 two_stage_opamp_dummy_magic_19_0.cap_res_X.t116 GNDA 0.184828f
C1785 two_stage_opamp_dummy_magic_19_0.cap_res_X.n16 GNDA 0.251826f
C1786 two_stage_opamp_dummy_magic_19_0.cap_res_X.t78 GNDA 0.184828f
C1787 two_stage_opamp_dummy_magic_19_0.cap_res_X.n17 GNDA 0.251826f
C1788 two_stage_opamp_dummy_magic_19_0.cap_res_X.t108 GNDA 0.184828f
C1789 two_stage_opamp_dummy_magic_19_0.cap_res_X.n18 GNDA 0.251826f
C1790 two_stage_opamp_dummy_magic_19_0.cap_res_X.t72 GNDA 0.184828f
C1791 two_stage_opamp_dummy_magic_19_0.cap_res_X.n19 GNDA 0.251826f
C1792 two_stage_opamp_dummy_magic_19_0.cap_res_X.t35 GNDA 0.184828f
C1793 two_stage_opamp_dummy_magic_19_0.cap_res_X.n20 GNDA 0.251826f
C1794 two_stage_opamp_dummy_magic_19_0.cap_res_X.t68 GNDA 0.184828f
C1795 two_stage_opamp_dummy_magic_19_0.cap_res_X.n21 GNDA 0.251826f
C1796 two_stage_opamp_dummy_magic_19_0.cap_res_X.t28 GNDA 0.184828f
C1797 two_stage_opamp_dummy_magic_19_0.cap_res_X.n22 GNDA 0.251826f
C1798 two_stage_opamp_dummy_magic_19_0.cap_res_X.t9 GNDA 0.184828f
C1799 two_stage_opamp_dummy_magic_19_0.cap_res_X.n23 GNDA 0.251826f
C1800 two_stage_opamp_dummy_magic_19_0.cap_res_X.t44 GNDA 0.184828f
C1801 two_stage_opamp_dummy_magic_19_0.cap_res_X.n24 GNDA 0.251826f
C1802 two_stage_opamp_dummy_magic_19_0.cap_res_X.t1 GNDA 0.184828f
C1803 two_stage_opamp_dummy_magic_19_0.cap_res_X.n25 GNDA 0.234498f
C1804 two_stage_opamp_dummy_magic_19_0.cap_res_X.t0 GNDA 0.3451f
C1805 two_stage_opamp_dummy_magic_19_0.cap_res_X.t40 GNDA 0.167396f
C1806 two_stage_opamp_dummy_magic_19_0.cap_res_X.n26 GNDA 0.217171f
C1807 two_stage_opamp_dummy_magic_19_0.cap_res_X.t121 GNDA 0.3451f
C1808 two_stage_opamp_dummy_magic_19_0.cap_res_X.t24 GNDA 0.346251f
C1809 two_stage_opamp_dummy_magic_19_0.cap_res_X.t57 GNDA 0.364834f
C1810 two_stage_opamp_dummy_magic_19_0.cap_res_X.t20 GNDA 0.185978f
C1811 two_stage_opamp_dummy_magic_19_0.cap_res_X.n27 GNDA 0.217171f
C1812 two_stage_opamp_dummy_magic_19_0.cap_res_X.t125 GNDA 0.3451f
C1813 two_stage_opamp_dummy_magic_19_0.cap_res_X.t65 GNDA 0.346251f
C1814 two_stage_opamp_dummy_magic_19_0.cap_res_X.t26 GNDA 0.185978f
C1815 two_stage_opamp_dummy_magic_19_0.cap_res_X.n28 GNDA 0.198589f
C1816 two_stage_opamp_dummy_magic_19_0.cap_res_X.t7 GNDA 0.3451f
C1817 two_stage_opamp_dummy_magic_19_0.cap_res_X.t87 GNDA 0.346251f
C1818 two_stage_opamp_dummy_magic_19_0.cap_res_X.t48 GNDA 0.185978f
C1819 two_stage_opamp_dummy_magic_19_0.cap_res_X.n29 GNDA 0.217171f
C1820 two_stage_opamp_dummy_magic_19_0.cap_res_X.t106 GNDA 0.3451f
C1821 two_stage_opamp_dummy_magic_19_0.cap_res_X.t49 GNDA 0.346251f
C1822 two_stage_opamp_dummy_magic_19_0.cap_res_X.t10 GNDA 0.185978f
C1823 two_stage_opamp_dummy_magic_19_0.cap_res_X.n30 GNDA 0.217171f
C1824 two_stage_opamp_dummy_magic_19_0.cap_res_X.t73 GNDA 0.3451f
C1825 two_stage_opamp_dummy_magic_19_0.cap_res_X.t12 GNDA 0.346251f
C1826 two_stage_opamp_dummy_magic_19_0.cap_res_X.t111 GNDA 0.185978f
C1827 two_stage_opamp_dummy_magic_19_0.cap_res_X.n31 GNDA 0.217171f
C1828 two_stage_opamp_dummy_magic_19_0.cap_res_X.t36 GNDA 0.3451f
C1829 two_stage_opamp_dummy_magic_19_0.cap_res_X.t90 GNDA 0.346251f
C1830 two_stage_opamp_dummy_magic_19_0.cap_res_X.t79 GNDA 0.364834f
C1831 two_stage_opamp_dummy_magic_19_0.cap_res_X.t113 GNDA 0.364834f
C1832 two_stage_opamp_dummy_magic_19_0.cap_res_X.t75 GNDA 0.185978f
C1833 two_stage_opamp_dummy_magic_19_0.cap_res_X.n32 GNDA 0.217171f
C1834 two_stage_opamp_dummy_magic_19_0.cap_res_X.t52 GNDA 0.3451f
C1835 two_stage_opamp_dummy_magic_19_0.cap_res_X.t41 GNDA 0.346251f
C1836 two_stage_opamp_dummy_magic_19_0.cap_res_X.t98 GNDA 0.364834f
C1837 two_stage_opamp_dummy_magic_19_0.cap_res_X.t134 GNDA 0.364834f
C1838 two_stage_opamp_dummy_magic_19_0.cap_res_X.t92 GNDA 0.185978f
C1839 two_stage_opamp_dummy_magic_19_0.cap_res_X.n33 GNDA 0.217171f
C1840 two_stage_opamp_dummy_magic_19_0.cap_res_X.t19 GNDA 0.3451f
C1841 two_stage_opamp_dummy_magic_19_0.cap_res_X.n34 GNDA 0.217171f
C1842 two_stage_opamp_dummy_magic_19_0.cap_res_X.t56 GNDA 0.185978f
C1843 two_stage_opamp_dummy_magic_19_0.cap_res_X.t95 GNDA 0.364834f
C1844 two_stage_opamp_dummy_magic_19_0.cap_res_X.t62 GNDA 0.364834f
C1845 two_stage_opamp_dummy_magic_19_0.cap_res_X.t6 GNDA 0.430822f
C1846 two_stage_opamp_dummy_magic_19_0.cap_res_X.t138 GNDA 0.292647f
C1847 VOUT-.t2 GNDA 0.045709f
C1848 VOUT-.t14 GNDA 0.045709f
C1849 VOUT-.n0 GNDA 0.102649f
C1850 VOUT-.t11 GNDA 0.045709f
C1851 VOUT-.t17 GNDA 0.045709f
C1852 VOUT-.n1 GNDA 0.136516f
C1853 VOUT-.t8 GNDA 0.045709f
C1854 VOUT-.t12 GNDA 0.045709f
C1855 VOUT-.n2 GNDA 0.136516f
C1856 VOUT-.t0 GNDA 0.045709f
C1857 VOUT-.t16 GNDA 0.045709f
C1858 VOUT-.n3 GNDA 0.132953f
C1859 VOUT-.n4 GNDA 0.526637f
C1860 VOUT-.t4 GNDA 0.045709f
C1861 VOUT-.t3 GNDA 0.045709f
C1862 VOUT-.n5 GNDA 0.132953f
C1863 VOUT-.n6 GNDA 0.267766f
C1864 VOUT-.t1 GNDA 0.045709f
C1865 VOUT-.t13 GNDA 0.045709f
C1866 VOUT-.n7 GNDA 0.132953f
C1867 VOUT-.n8 GNDA 0.267766f
C1868 VOUT-.n9 GNDA 0.281725f
C1869 VOUT-.n10 GNDA 0.356093f
C1870 VOUT-.t26 GNDA 0.30992f
C1871 VOUT-.t119 GNDA 0.30473f
C1872 VOUT-.n11 GNDA 0.204311f
C1873 VOUT-.t33 GNDA 0.30473f
C1874 VOUT-.n12 GNDA 0.133319f
C1875 VOUT-.t36 GNDA 0.30992f
C1876 VOUT-.t122 GNDA 0.30473f
C1877 VOUT-.n13 GNDA 0.204311f
C1878 VOUT-.t90 GNDA 0.30473f
C1879 VOUT-.t82 GNDA 0.30927f
C1880 VOUT-.t42 GNDA 0.30927f
C1881 VOUT-.t92 GNDA 0.30927f
C1882 VOUT-.t74 GNDA 0.30927f
C1883 VOUT-.t141 GNDA 0.30927f
C1884 VOUT-.t38 GNDA 0.30927f
C1885 VOUT-.t105 GNDA 0.30927f
C1886 VOUT-.t126 GNDA 0.30927f
C1887 VOUT-.t154 GNDA 0.30927f
C1888 VOUT-.t95 GNDA 0.30927f
C1889 VOUT-.t65 GNDA 0.30927f
C1890 VOUT-.t62 GNDA 0.30927f
C1891 VOUT-.t114 GNDA 0.30927f
C1892 VOUT-.t24 GNDA 0.30927f
C1893 VOUT-.t71 GNDA 0.30927f
C1894 VOUT-.t113 GNDA 0.30927f
C1895 VOUT-.t148 GNDA 0.30473f
C1896 VOUT-.n14 GNDA 0.33374f
C1897 VOUT-.t60 GNDA 0.30473f
C1898 VOUT-.n15 GNDA 0.390877f
C1899 VOUT-.t93 GNDA 0.30473f
C1900 VOUT-.n16 GNDA 0.390877f
C1901 VOUT-.t127 GNDA 0.30473f
C1902 VOUT-.n17 GNDA 0.390877f
C1903 VOUT-.t25 GNDA 0.30473f
C1904 VOUT-.n18 GNDA 0.390877f
C1905 VOUT-.t72 GNDA 0.30473f
C1906 VOUT-.n19 GNDA 0.390877f
C1907 VOUT-.t110 GNDA 0.30473f
C1908 VOUT-.n20 GNDA 0.390877f
C1909 VOUT-.t142 GNDA 0.30473f
C1910 VOUT-.n21 GNDA 0.262098f
C1911 VOUT-.t56 GNDA 0.30473f
C1912 VOUT-.n22 GNDA 0.262098f
C1913 VOUT-.n23 GNDA 0.247593f
C1914 VOUT-.t140 GNDA 0.30992f
C1915 VOUT-.t89 GNDA 0.30473f
C1916 VOUT-.n24 GNDA 0.204311f
C1917 VOUT-.t59 GNDA 0.30473f
C1918 VOUT-.t111 GNDA 0.30992f
C1919 VOUT-.t21 GNDA 0.30473f
C1920 VOUT-.n25 GNDA 0.204311f
C1921 VOUT-.n26 GNDA 0.247593f
C1922 VOUT-.t41 GNDA 0.30992f
C1923 VOUT-.t129 GNDA 0.30473f
C1924 VOUT-.n27 GNDA 0.204311f
C1925 VOUT-.t98 GNDA 0.30473f
C1926 VOUT-.t151 GNDA 0.30992f
C1927 VOUT-.t63 GNDA 0.30473f
C1928 VOUT-.n28 GNDA 0.204311f
C1929 VOUT-.n29 GNDA 0.247593f
C1930 VOUT-.t80 GNDA 0.30992f
C1931 VOUT-.t30 GNDA 0.30473f
C1932 VOUT-.n30 GNDA 0.204311f
C1933 VOUT-.t134 GNDA 0.30473f
C1934 VOUT-.t51 GNDA 0.30992f
C1935 VOUT-.t103 GNDA 0.30473f
C1936 VOUT-.n31 GNDA 0.204311f
C1937 VOUT-.n32 GNDA 0.247593f
C1938 VOUT-.t49 GNDA 0.30992f
C1939 VOUT-.t135 GNDA 0.30473f
C1940 VOUT-.n33 GNDA 0.204311f
C1941 VOUT-.t102 GNDA 0.30473f
C1942 VOUT-.t19 GNDA 0.30992f
C1943 VOUT-.t67 GNDA 0.30473f
C1944 VOUT-.n34 GNDA 0.204311f
C1945 VOUT-.n35 GNDA 0.247593f
C1946 VOUT-.t85 GNDA 0.30992f
C1947 VOUT-.t34 GNDA 0.30473f
C1948 VOUT-.n36 GNDA 0.204311f
C1949 VOUT-.t139 GNDA 0.30473f
C1950 VOUT-.t55 GNDA 0.30992f
C1951 VOUT-.t106 GNDA 0.30473f
C1952 VOUT-.n37 GNDA 0.204311f
C1953 VOUT-.n38 GNDA 0.247593f
C1954 VOUT-.t68 GNDA 0.30992f
C1955 VOUT-.t86 GNDA 0.30473f
C1956 VOUT-.n39 GNDA 0.204311f
C1957 VOUT-.t54 GNDA 0.30473f
C1958 VOUT-.n40 GNDA 0.133319f
C1959 VOUT-.t29 GNDA 0.30992f
C1960 VOUT-.t52 GNDA 0.30473f
C1961 VOUT-.n41 GNDA 0.204311f
C1962 VOUT-.t155 GNDA 0.30473f
C1963 VOUT-.t156 GNDA 0.30927f
C1964 VOUT-.t132 GNDA 0.30992f
C1965 VOUT-.t99 GNDA 0.30473f
C1966 VOUT-.n42 GNDA 0.19955f
C1967 VOUT-.t35 GNDA 0.30927f
C1968 VOUT-.t150 GNDA 0.30992f
C1969 VOUT-.t94 GNDA 0.30473f
C1970 VOUT-.n43 GNDA 0.204311f
C1971 VOUT-.t61 GNDA 0.30473f
C1972 VOUT-.n44 GNDA 0.128558f
C1973 VOUT-.t137 GNDA 0.30927f
C1974 VOUT-.t115 GNDA 0.30992f
C1975 VOUT-.t58 GNDA 0.30473f
C1976 VOUT-.n45 GNDA 0.204311f
C1977 VOUT-.t22 GNDA 0.30473f
C1978 VOUT-.n46 GNDA 0.128558f
C1979 VOUT-.t104 GNDA 0.30927f
C1980 VOUT-.t66 GNDA 0.30992f
C1981 VOUT-.t77 GNDA 0.30473f
C1982 VOUT-.n47 GNDA 0.204311f
C1983 VOUT-.t43 GNDA 0.30473f
C1984 VOUT-.n48 GNDA 0.128558f
C1985 VOUT-.t120 GNDA 0.30927f
C1986 VOUT-.t144 GNDA 0.30927f
C1987 VOUT-.t83 GNDA 0.30927f
C1988 VOUT-.t107 GNDA 0.309525f
C1989 VOUT-.t50 GNDA 0.30927f
C1990 VOUT-.t69 GNDA 0.309525f
C1991 VOUT-.t149 GNDA 0.30927f
C1992 VOUT-.t91 GNDA 0.309525f
C1993 VOUT-.t31 GNDA 0.30927f
C1994 VOUT-.t130 GNDA 0.30473f
C1995 VOUT-.n49 GNDA 0.337294f
C1996 VOUT-.t108 GNDA 0.30473f
C1997 VOUT-.n50 GNDA 0.394431f
C1998 VOUT-.t146 GNDA 0.30473f
C1999 VOUT-.n51 GNDA 0.394431f
C2000 VOUT-.t45 GNDA 0.30473f
C2001 VOUT-.n52 GNDA 0.390877f
C2002 VOUT-.t81 GNDA 0.30473f
C2003 VOUT-.n53 GNDA 0.323996f
C2004 VOUT-.t64 GNDA 0.30473f
C2005 VOUT-.n54 GNDA 0.323996f
C2006 VOUT-.t100 GNDA 0.30473f
C2007 VOUT-.n55 GNDA 0.323996f
C2008 VOUT-.t136 GNDA 0.30473f
C2009 VOUT-.n56 GNDA 0.323996f
C2010 VOUT-.t116 GNDA 0.30473f
C2011 VOUT-.n57 GNDA 0.262098f
C2012 VOUT-.n58 GNDA 0.247593f
C2013 VOUT-.t125 GNDA 0.30992f
C2014 VOUT-.t152 GNDA 0.30473f
C2015 VOUT-.n59 GNDA 0.204311f
C2016 VOUT-.t112 GNDA 0.30473f
C2017 VOUT-.t73 GNDA 0.30992f
C2018 VOUT-.n60 GNDA 0.318585f
C2019 VOUT-.t23 GNDA 0.30992f
C2020 VOUT-.t47 GNDA 0.30473f
C2021 VOUT-.n61 GNDA 0.204311f
C2022 VOUT-.t147 GNDA 0.30473f
C2023 VOUT-.t109 GNDA 0.30992f
C2024 VOUT-.n62 GNDA 0.318585f
C2025 VOUT-.t76 GNDA 0.30992f
C2026 VOUT-.t27 GNDA 0.30473f
C2027 VOUT-.n63 GNDA 0.204311f
C2028 VOUT-.t128 GNDA 0.30473f
C2029 VOUT-.t44 GNDA 0.30992f
C2030 VOUT-.t97 GNDA 0.30473f
C2031 VOUT-.n64 GNDA 0.204311f
C2032 VOUT-.n65 GNDA 0.247593f
C2033 VOUT-.t37 GNDA 0.30992f
C2034 VOUT-.t123 GNDA 0.30473f
C2035 VOUT-.n66 GNDA 0.204311f
C2036 VOUT-.t88 GNDA 0.30473f
C2037 VOUT-.t143 GNDA 0.30992f
C2038 VOUT-.t57 GNDA 0.30473f
C2039 VOUT-.n67 GNDA 0.204311f
C2040 VOUT-.n68 GNDA 0.247593f
C2041 VOUT-.t70 GNDA 0.30992f
C2042 VOUT-.t20 GNDA 0.30473f
C2043 VOUT-.n69 GNDA 0.204311f
C2044 VOUT-.t121 GNDA 0.30473f
C2045 VOUT-.t39 GNDA 0.30992f
C2046 VOUT-.t87 GNDA 0.30473f
C2047 VOUT-.n70 GNDA 0.204311f
C2048 VOUT-.n71 GNDA 0.247593f
C2049 VOUT-.t32 GNDA 0.30992f
C2050 VOUT-.t118 GNDA 0.30473f
C2051 VOUT-.n72 GNDA 0.204311f
C2052 VOUT-.t84 GNDA 0.30473f
C2053 VOUT-.t138 GNDA 0.30992f
C2054 VOUT-.t53 GNDA 0.30473f
C2055 VOUT-.n73 GNDA 0.204311f
C2056 VOUT-.n74 GNDA 0.247593f
C2057 VOUT-.t131 GNDA 0.30992f
C2058 VOUT-.t79 GNDA 0.30473f
C2059 VOUT-.n75 GNDA 0.204311f
C2060 VOUT-.t48 GNDA 0.30473f
C2061 VOUT-.t101 GNDA 0.30992f
C2062 VOUT-.t153 GNDA 0.30473f
C2063 VOUT-.n76 GNDA 0.204311f
C2064 VOUT-.n77 GNDA 0.247593f
C2065 VOUT-.t28 GNDA 0.30992f
C2066 VOUT-.t117 GNDA 0.30473f
C2067 VOUT-.n78 GNDA 0.204311f
C2068 VOUT-.t78 GNDA 0.30473f
C2069 VOUT-.t133 GNDA 0.30992f
C2070 VOUT-.t46 GNDA 0.30473f
C2071 VOUT-.n79 GNDA 0.204311f
C2072 VOUT-.n80 GNDA 0.247593f
C2073 VOUT-.t124 GNDA 0.30992f
C2074 VOUT-.t75 GNDA 0.30473f
C2075 VOUT-.n81 GNDA 0.204311f
C2076 VOUT-.t40 GNDA 0.30473f
C2077 VOUT-.n82 GNDA 0.247593f
C2078 VOUT-.t145 GNDA 0.30473f
C2079 VOUT-.n83 GNDA 0.133319f
C2080 VOUT-.t96 GNDA 0.30473f
C2081 VOUT-.n84 GNDA 0.19441f
C2082 VOUT-.n85 GNDA 0.227911f
C2083 VOUT-.t5 GNDA 0.053328f
C2084 VOUT-.t9 GNDA 0.053328f
C2085 VOUT-.n86 GNDA 0.249232f
C2086 VOUT-.t18 GNDA 0.053328f
C2087 VOUT-.t6 GNDA 0.053328f
C2088 VOUT-.n87 GNDA 0.23402f
C2089 VOUT-.n88 GNDA 0.455316f
C2090 VOUT-.t10 GNDA 0.053328f
C2091 VOUT-.t15 GNDA 0.053328f
C2092 VOUT-.n89 GNDA 0.23402f
C2093 VOUT-.n90 GNDA 0.243523f
C2094 VOUT-.t7 GNDA 0.088718f
C2095 VOUT-.n91 GNDA 0.090646f
C2096 bgr_9_0.V_TOP.t24 GNDA 0.097271f
C2097 bgr_9_0.V_TOP.t33 GNDA 0.097271f
C2098 bgr_9_0.V_TOP.t39 GNDA 0.097271f
C2099 bgr_9_0.V_TOP.t16 GNDA 0.097271f
C2100 bgr_9_0.V_TOP.t15 GNDA 0.097271f
C2101 bgr_9_0.V_TOP.t28 GNDA 0.097271f
C2102 bgr_9_0.V_TOP.t38 GNDA 0.097271f
C2103 bgr_9_0.V_TOP.t14 GNDA 0.097271f
C2104 bgr_9_0.V_TOP.t27 GNDA 0.097271f
C2105 bgr_9_0.V_TOP.t26 GNDA 0.097271f
C2106 bgr_9_0.V_TOP.t37 GNDA 0.097271f
C2107 bgr_9_0.V_TOP.t46 GNDA 0.097271f
C2108 bgr_9_0.V_TOP.t18 GNDA 0.097271f
C2109 bgr_9_0.V_TOP.t30 GNDA 0.097271f
C2110 bgr_9_0.V_TOP.t29 GNDA 0.127158f
C2111 bgr_9_0.V_TOP.n0 GNDA 0.071091f
C2112 bgr_9_0.V_TOP.n1 GNDA 0.051878f
C2113 bgr_9_0.V_TOP.n2 GNDA 0.051878f
C2114 bgr_9_0.V_TOP.n3 GNDA 0.051878f
C2115 bgr_9_0.V_TOP.n4 GNDA 0.051878f
C2116 bgr_9_0.V_TOP.n5 GNDA 0.048377f
C2117 bgr_9_0.V_TOP.t7 GNDA 0.126138f
C2118 bgr_9_0.V_TOP.t40 GNDA 0.370558f
C2119 bgr_9_0.V_TOP.t31 GNDA 0.37687f
C2120 bgr_9_0.V_TOP.t35 GNDA 0.370558f
C2121 bgr_9_0.V_TOP.n6 GNDA 0.248447f
C2122 bgr_9_0.V_TOP.t32 GNDA 0.370558f
C2123 bgr_9_0.V_TOP.t22 GNDA 0.37687f
C2124 bgr_9_0.V_TOP.n7 GNDA 0.317927f
C2125 bgr_9_0.V_TOP.t20 GNDA 0.37687f
C2126 bgr_9_0.V_TOP.t25 GNDA 0.370558f
C2127 bgr_9_0.V_TOP.n8 GNDA 0.248447f
C2128 bgr_9_0.V_TOP.t21 GNDA 0.370558f
C2129 bgr_9_0.V_TOP.t45 GNDA 0.37687f
C2130 bgr_9_0.V_TOP.n9 GNDA 0.387406f
C2131 bgr_9_0.V_TOP.t42 GNDA 0.37687f
C2132 bgr_9_0.V_TOP.t49 GNDA 0.370558f
C2133 bgr_9_0.V_TOP.n10 GNDA 0.248447f
C2134 bgr_9_0.V_TOP.t44 GNDA 0.370558f
C2135 bgr_9_0.V_TOP.t36 GNDA 0.37687f
C2136 bgr_9_0.V_TOP.n11 GNDA 0.387406f
C2137 bgr_9_0.V_TOP.t17 GNDA 0.37687f
C2138 bgr_9_0.V_TOP.t23 GNDA 0.370558f
C2139 bgr_9_0.V_TOP.n12 GNDA 0.248447f
C2140 bgr_9_0.V_TOP.t19 GNDA 0.370558f
C2141 bgr_9_0.V_TOP.t43 GNDA 0.37687f
C2142 bgr_9_0.V_TOP.n13 GNDA 0.387406f
C2143 bgr_9_0.V_TOP.t34 GNDA 0.37687f
C2144 bgr_9_0.V_TOP.t41 GNDA 0.370558f
C2145 bgr_9_0.V_TOP.n14 GNDA 0.317927f
C2146 bgr_9_0.V_TOP.t47 GNDA 0.370558f
C2147 bgr_9_0.V_TOP.n15 GNDA 0.162119f
C2148 bgr_9_0.V_TOP.n16 GNDA 0.554811f
C2149 bgr_9_0.V_TOP.t3 GNDA 0.104243f
C2150 bgr_9_0.V_TOP.n17 GNDA 0.73814f
C2151 bgr_9_0.V_TOP.n18 GNDA 0.023109f
C2152 bgr_9_0.V_TOP.n19 GNDA 0.422529f
C2153 bgr_9_0.V_TOP.n20 GNDA 0.022398f
C2154 bgr_9_0.V_TOP.n21 GNDA 0.023262f
C2155 bgr_9_0.V_TOP.n22 GNDA 0.023109f
C2156 bgr_9_0.V_TOP.n23 GNDA 0.213681f
C2157 bgr_9_0.V_TOP.n24 GNDA 0.129796f
C2158 bgr_9_0.V_TOP.n25 GNDA 0.074112f
C2159 bgr_9_0.V_TOP.n26 GNDA 0.023109f
C2160 bgr_9_0.V_TOP.n27 GNDA 0.127893f
C2161 bgr_9_0.V_TOP.n28 GNDA 0.023109f
C2162 bgr_9_0.V_TOP.n29 GNDA 0.126677f
C2163 bgr_9_0.V_TOP.n30 GNDA 0.277504f
C2164 bgr_9_0.V_TOP.n31 GNDA 0.019602f
C2165 bgr_9_0.V_TOP.n32 GNDA 0.048377f
C2166 bgr_9_0.V_TOP.n33 GNDA 0.051878f
C2167 bgr_9_0.V_TOP.n34 GNDA 0.051878f
C2168 bgr_9_0.V_TOP.n35 GNDA 0.051878f
C2169 bgr_9_0.V_TOP.n36 GNDA 0.051878f
C2170 bgr_9_0.V_TOP.n37 GNDA 0.051878f
C2171 bgr_9_0.V_TOP.n38 GNDA 0.051878f
C2172 bgr_9_0.V_TOP.n39 GNDA 0.048377f
C2173 bgr_9_0.V_TOP.t48 GNDA 0.112091f
C2174 VDDA.t204 GNDA 0.029949f
C2175 VDDA.t212 GNDA 0.029949f
C2176 VDDA.n0 GNDA 0.063256f
C2177 VDDA.t198 GNDA 0.029949f
C2178 VDDA.t208 GNDA 0.029949f
C2179 VDDA.n1 GNDA 0.075235f
C2180 VDDA.n2 GNDA 0.205432f
C2181 VDDA.t315 GNDA 0.057468f
C2182 VDDA.t317 GNDA 0.106534f
C2183 VDDA.t230 GNDA 0.029949f
C2184 VDDA.t234 GNDA 0.029949f
C2185 VDDA.n3 GNDA 0.075235f
C2186 VDDA.n4 GNDA 0.244164f
C2187 VDDA.n5 GNDA 0.43585f
C2188 VDDA.t316 GNDA 0.253905f
C2189 VDDA.t229 GNDA 0.200232f
C2190 VDDA.t233 GNDA 0.200232f
C2191 VDDA.t197 GNDA 0.200232f
C2192 VDDA.t207 GNDA 0.200232f
C2193 VDDA.t203 GNDA 0.200232f
C2194 VDDA.t211 GNDA 0.200232f
C2195 VDDA.t219 GNDA 0.200232f
C2196 VDDA.t225 GNDA 0.200232f
C2197 VDDA.t201 GNDA 0.200232f
C2198 VDDA.t195 GNDA 0.200232f
C2199 VDDA.t260 GNDA 0.255285f
C2200 VDDA.t261 GNDA 0.106534f
C2201 VDDA.n6 GNDA 0.340751f
C2202 VDDA.t259 GNDA 0.053036f
C2203 VDDA.n7 GNDA 0.113716f
C2204 VDDA.t202 GNDA 0.029949f
C2205 VDDA.t196 GNDA 0.029949f
C2206 VDDA.n8 GNDA 0.075235f
C2207 VDDA.n9 GNDA 0.223465f
C2208 VDDA.t220 GNDA 0.029949f
C2209 VDDA.t226 GNDA 0.029949f
C2210 VDDA.n10 GNDA 0.075235f
C2211 VDDA.n11 GNDA 0.205432f
C2212 VDDA.n12 GNDA 0.027382f
C2213 VDDA.n13 GNDA 0.23219f
C2214 VDDA.t238 GNDA 0.025671f
C2215 VDDA.t101 GNDA 0.025671f
C2216 VDDA.n14 GNDA 0.086154f
C2217 VDDA.t169 GNDA 0.025671f
C2218 VDDA.t66 GNDA 0.025671f
C2219 VDDA.n15 GNDA 0.083248f
C2220 VDDA.n16 GNDA 0.314065f
C2221 VDDA.t144 GNDA 0.025671f
C2222 VDDA.t118 GNDA 0.025671f
C2223 VDDA.n17 GNDA 0.083248f
C2224 VDDA.n18 GNDA 0.16148f
C2225 VDDA.t78 GNDA 0.025671f
C2226 VDDA.t93 GNDA 0.025671f
C2227 VDDA.n19 GNDA 0.083248f
C2228 VDDA.n20 GNDA 0.16148f
C2229 VDDA.t171 GNDA 0.025671f
C2230 VDDA.t67 GNDA 0.025671f
C2231 VDDA.n21 GNDA 0.083248f
C2232 VDDA.n22 GNDA 0.16148f
C2233 VDDA.t39 GNDA 0.025671f
C2234 VDDA.t239 GNDA 0.025671f
C2235 VDDA.n23 GNDA 0.083248f
C2236 VDDA.n24 GNDA 0.23931f
C2237 VDDA.t268 GNDA 0.025774f
C2238 VDDA.t270 GNDA 0.061056f
C2239 VDDA.t253 GNDA 0.026078f
C2240 VDDA.t255 GNDA 0.061056f
C2241 VDDA.n25 GNDA 0.260694f
C2242 VDDA.t254 GNDA 0.15211f
C2243 VDDA.t98 GNDA 0.112951f
C2244 VDDA.t170 GNDA 0.112951f
C2245 VDDA.t130 GNDA 0.112951f
C2246 VDDA.t102 GNDA 0.112951f
C2247 VDDA.t65 GNDA 0.112951f
C2248 VDDA.t411 GNDA 0.112951f
C2249 VDDA.t11 GNDA 0.112951f
C2250 VDDA.t369 GNDA 0.112951f
C2251 VDDA.t410 GNDA 0.112951f
C2252 VDDA.t38 GNDA 0.112951f
C2253 VDDA.t269 GNDA 0.15211f
C2254 VDDA.n26 GNDA 0.187188f
C2255 VDDA.n27 GNDA 0.118307f
C2256 VDDA.n28 GNDA 0.221235f
C2257 VDDA.t375 GNDA 0.051342f
C2258 VDDA.t168 GNDA 0.051342f
C2259 VDDA.n29 GNDA 0.149335f
C2260 VDDA.n30 GNDA 0.300759f
C2261 VDDA.t339 GNDA 0.062544f
C2262 VDDA.t329 GNDA 0.180684f
C2263 VDDA.t327 GNDA 0.062544f
C2264 VDDA.t97 GNDA 0.051342f
C2265 VDDA.t18 GNDA 0.051342f
C2266 VDDA.n31 GNDA 0.149335f
C2267 VDDA.n32 GNDA 0.300759f
C2268 VDDA.t371 GNDA 0.051342f
C2269 VDDA.t115 GNDA 0.051342f
C2270 VDDA.n33 GNDA 0.149335f
C2271 VDDA.n34 GNDA 0.300759f
C2272 VDDA.t373 GNDA 0.051342f
C2273 VDDA.t69 GNDA 0.051342f
C2274 VDDA.n35 GNDA 0.149335f
C2275 VDDA.n36 GNDA 0.300759f
C2276 VDDA.t377 GNDA 0.051342f
C2277 VDDA.t71 GNDA 0.051342f
C2278 VDDA.n37 GNDA 0.149335f
C2279 VDDA.n38 GNDA 0.318253f
C2280 VDDA.n39 GNDA 0.133198f
C2281 VDDA.n40 GNDA 0.603628f
C2282 VDDA.t328 GNDA 0.391455f
C2283 VDDA.t376 GNDA 0.301204f
C2284 VDDA.t70 GNDA 0.301204f
C2285 VDDA.t372 GNDA 0.301204f
C2286 VDDA.t68 GNDA 0.301204f
C2287 VDDA.t370 GNDA 0.301204f
C2288 VDDA.t114 GNDA 0.301204f
C2289 VDDA.t96 GNDA 0.301204f
C2290 VDDA.t17 GNDA 0.301204f
C2291 VDDA.t374 GNDA 0.301204f
C2292 VDDA.t167 GNDA 0.301204f
C2293 VDDA.t340 GNDA 0.391455f
C2294 VDDA.t341 GNDA 0.180684f
C2295 VDDA.n41 GNDA 0.603628f
C2296 VDDA.n42 GNDA 0.131011f
C2297 VDDA.n43 GNDA 0.06039f
C2298 VDDA.n44 GNDA 0.09064f
C2299 VDDA.t13 GNDA 0.021392f
C2300 VDDA.t56 GNDA 0.021392f
C2301 VDDA.n45 GNDA 0.051019f
C2302 VDDA.n46 GNDA 0.176596f
C2303 VDDA.t351 GNDA 0.031741f
C2304 VDDA.t313 GNDA 0.151992f
C2305 VDDA.t273 GNDA 0.076639f
C2306 VDDA.n47 GNDA 0.098967f
C2307 VDDA.t312 GNDA 0.031741f
C2308 VDDA.t271 GNDA 0.031741f
C2309 VDDA.n48 GNDA 0.103484f
C2310 VDDA.n49 GNDA 0.02781f
C2311 VDDA.t303 GNDA 0.031741f
C2312 VDDA.t305 GNDA 0.076639f
C2313 VDDA.t47 GNDA 0.136483f
C2314 VDDA.t14 GNDA 0.136483f
C2315 VDDA.t103 GNDA 0.136483f
C2316 VDDA.t36 GNDA 0.136483f
C2317 VDDA.t304 GNDA 0.18361f
C2318 VDDA.n50 GNDA 0.236669f
C2319 VDDA.n51 GNDA 0.107572f
C2320 VDDA.t15 GNDA 0.021392f
C2321 VDDA.t104 GNDA 0.021392f
C2322 VDDA.n52 GNDA 0.051019f
C2323 VDDA.n53 GNDA 0.196895f
C2324 VDDA.n54 GNDA 0.02781f
C2325 VDDA.n55 GNDA 0.103484f
C2326 VDDA.t314 GNDA 0.076639f
C2327 VDDA.n56 GNDA 0.098967f
C2328 VDDA.n57 GNDA 0.039362f
C2329 VDDA.n58 GNDA 0.124717f
C2330 VDDA.t272 GNDA 0.151992f
C2331 VDDA.t35 GNDA 0.136483f
C2332 VDDA.t55 GNDA 0.136483f
C2333 VDDA.t12 GNDA 0.136483f
C2334 VDDA.t48 GNDA 0.136483f
C2335 VDDA.t352 GNDA 0.18361f
C2336 VDDA.t353 GNDA 0.076639f
C2337 VDDA.n59 GNDA 0.236669f
C2338 VDDA.n60 GNDA 0.103484f
C2339 VDDA.n61 GNDA 0.115909f
C2340 VDDA.n62 GNDA 0.136807f
C2341 VDDA.n63 GNDA 0.210837f
C2342 VDDA.t236 GNDA 0.029949f
C2343 VDDA.t200 GNDA 0.029949f
C2344 VDDA.n64 GNDA 0.063256f
C2345 VDDA.t224 GNDA 0.029949f
C2346 VDDA.t232 GNDA 0.029949f
C2347 VDDA.n65 GNDA 0.075235f
C2348 VDDA.n66 GNDA 0.205432f
C2349 VDDA.t300 GNDA 0.057468f
C2350 VDDA.t302 GNDA 0.106534f
C2351 VDDA.t246 GNDA 0.106534f
C2352 VDDA.t244 GNDA 0.053036f
C2353 VDDA.t206 GNDA 0.029949f
C2354 VDDA.t216 GNDA 0.029949f
C2355 VDDA.n67 GNDA 0.075235f
C2356 VDDA.n68 GNDA 0.223465f
C2357 VDDA.n69 GNDA 0.113716f
C2358 VDDA.n70 GNDA 0.340751f
C2359 VDDA.t245 GNDA 0.255285f
C2360 VDDA.t205 GNDA 0.200232f
C2361 VDDA.t215 GNDA 0.200232f
C2362 VDDA.t223 GNDA 0.200232f
C2363 VDDA.t231 GNDA 0.200232f
C2364 VDDA.t235 GNDA 0.200232f
C2365 VDDA.t199 GNDA 0.200232f
C2366 VDDA.t209 GNDA 0.200232f
C2367 VDDA.t217 GNDA 0.200232f
C2368 VDDA.t213 GNDA 0.200232f
C2369 VDDA.t221 GNDA 0.200232f
C2370 VDDA.t301 GNDA 0.253905f
C2371 VDDA.n71 GNDA 0.43585f
C2372 VDDA.t214 GNDA 0.029949f
C2373 VDDA.t222 GNDA 0.029949f
C2374 VDDA.n72 GNDA 0.075235f
C2375 VDDA.n73 GNDA 0.244164f
C2376 VDDA.t210 GNDA 0.029949f
C2377 VDDA.t218 GNDA 0.029949f
C2378 VDDA.n74 GNDA 0.075235f
C2379 VDDA.n75 GNDA 0.205432f
C2380 VDDA.n76 GNDA 0.027382f
C2381 VDDA.n77 GNDA 0.23219f
C2382 VDDA.t116 GNDA 0.025671f
C2383 VDDA.t237 GNDA 0.025671f
C2384 VDDA.n78 GNDA 0.086154f
C2385 VDDA.t138 GNDA 0.025671f
C2386 VDDA.t49 GNDA 0.025671f
C2387 VDDA.n79 GNDA 0.083248f
C2388 VDDA.n80 GNDA 0.314065f
C2389 VDDA.t139 GNDA 0.025671f
C2390 VDDA.t135 GNDA 0.025671f
C2391 VDDA.n81 GNDA 0.083248f
C2392 VDDA.n82 GNDA 0.16148f
C2393 VDDA.t54 GNDA 0.025671f
C2394 VDDA.t189 GNDA 0.025671f
C2395 VDDA.n83 GNDA 0.083248f
C2396 VDDA.n84 GNDA 0.16148f
C2397 VDDA.t40 GNDA 0.025671f
C2398 VDDA.t16 GNDA 0.025671f
C2399 VDDA.n85 GNDA 0.083248f
C2400 VDDA.n86 GNDA 0.16148f
C2401 VDDA.t240 GNDA 0.025671f
C2402 VDDA.t387 GNDA 0.025671f
C2403 VDDA.n87 GNDA 0.083248f
C2404 VDDA.n88 GNDA 0.23931f
C2405 VDDA.t309 GNDA 0.025774f
C2406 VDDA.t324 GNDA 0.026078f
C2407 VDDA.t326 GNDA 0.061056f
C2408 VDDA.n89 GNDA 0.260694f
C2409 VDDA.t325 GNDA 0.15211f
C2410 VDDA.t184 GNDA 0.112951f
C2411 VDDA.t51 GNDA 0.112951f
C2412 VDDA.t50 GNDA 0.112951f
C2413 VDDA.t32 GNDA 0.112951f
C2414 VDDA.t190 GNDA 0.112951f
C2415 VDDA.t37 GNDA 0.112951f
C2416 VDDA.t8 GNDA 0.112951f
C2417 VDDA.t117 GNDA 0.112951f
C2418 VDDA.t31 GNDA 0.112951f
C2419 VDDA.t92 GNDA 0.112951f
C2420 VDDA.t310 GNDA 0.15211f
C2421 VDDA.t311 GNDA 0.061056f
C2422 VDDA.n90 GNDA 0.187188f
C2423 VDDA.n91 GNDA 0.118307f
C2424 VDDA.n92 GNDA 0.221235f
C2425 VDDA.t113 GNDA 0.051342f
C2426 VDDA.t188 GNDA 0.051342f
C2427 VDDA.n93 GNDA 0.149335f
C2428 VDDA.n94 GNDA 0.300759f
C2429 VDDA.t256 GNDA 0.062544f
C2430 VDDA.t276 GNDA 0.180684f
C2431 VDDA.t274 GNDA 0.062544f
C2432 VDDA.t137 GNDA 0.051342f
C2433 VDDA.t5 GNDA 0.051342f
C2434 VDDA.n95 GNDA 0.149335f
C2435 VDDA.n96 GNDA 0.300759f
C2436 VDDA.t111 GNDA 0.051342f
C2437 VDDA.t166 GNDA 0.051342f
C2438 VDDA.n97 GNDA 0.149335f
C2439 VDDA.n98 GNDA 0.300759f
C2440 VDDA.t385 GNDA 0.051342f
C2441 VDDA.t34 GNDA 0.051342f
C2442 VDDA.n99 GNDA 0.149335f
C2443 VDDA.n100 GNDA 0.300759f
C2444 VDDA.t30 GNDA 0.051342f
C2445 VDDA.t53 GNDA 0.051342f
C2446 VDDA.n101 GNDA 0.149335f
C2447 VDDA.n102 GNDA 0.318253f
C2448 VDDA.n103 GNDA 0.133198f
C2449 VDDA.n104 GNDA 0.603628f
C2450 VDDA.t275 GNDA 0.391455f
C2451 VDDA.t52 GNDA 0.301204f
C2452 VDDA.t29 GNDA 0.301204f
C2453 VDDA.t33 GNDA 0.301204f
C2454 VDDA.t384 GNDA 0.301204f
C2455 VDDA.t165 GNDA 0.301204f
C2456 VDDA.t110 GNDA 0.301204f
C2457 VDDA.t4 GNDA 0.301204f
C2458 VDDA.t136 GNDA 0.301204f
C2459 VDDA.t187 GNDA 0.301204f
C2460 VDDA.t112 GNDA 0.301204f
C2461 VDDA.t257 GNDA 0.391455f
C2462 VDDA.t258 GNDA 0.180684f
C2463 VDDA.n105 GNDA 0.603628f
C2464 VDDA.n106 GNDA 0.131011f
C2465 VDDA.n107 GNDA 0.06039f
C2466 VDDA.n108 GNDA 0.181849f
C2467 VDDA.n109 GNDA 0.21618f
C2468 VDDA.n110 GNDA 0.200892f
C2469 VDDA.t290 GNDA 0.03219f
C2470 VDDA.t293 GNDA 0.055595f
C2471 VDDA.t279 GNDA 0.137921f
C2472 VDDA.t278 GNDA 0.183819f
C2473 VDDA.t398 GNDA 0.112951f
C2474 VDDA.t291 GNDA 0.149021f
C2475 VDDA.n111 GNDA 0.167387f
C2476 VDDA.n112 GNDA 0.08522f
C2477 VDDA.t399 GNDA 0.015403f
C2478 VDDA.t292 GNDA 0.015403f
C2479 VDDA.n113 GNDA 0.034437f
C2480 VDDA.n114 GNDA 0.125622f
C2481 VDDA.t277 GNDA 0.032602f
C2482 VDDA.n115 GNDA 0.090686f
C2483 VDDA.n116 GNDA 0.082274f
C2484 VDDA.n117 GNDA 0.21489f
C2485 VDDA.t345 GNDA 0.053036f
C2486 VDDA.t228 GNDA 0.029949f
C2487 VDDA.n118 GNDA 0.075235f
C2488 VDDA.t299 GNDA 0.136483f
C2489 VDDA.t297 GNDA 0.053036f
C2490 VDDA.n119 GNDA 0.112023f
C2491 VDDA.n120 GNDA 0.340751f
C2492 VDDA.t298 GNDA 0.255285f
C2493 VDDA.t227 GNDA 0.200232f
C2494 VDDA.t346 GNDA 0.255285f
C2495 VDDA.t347 GNDA 0.106534f
C2496 VDDA.n121 GNDA 0.340751f
C2497 VDDA.n122 GNDA 0.111212f
C2498 VDDA.n123 GNDA 0.048843f
C2499 VDDA.n124 GNDA 0.242807f
C2500 VDDA.n125 GNDA 4.59792f
C2501 VDDA.t27 GNDA 0.478332f
C2502 VDDA.t46 GNDA 0.480066f
C2503 VDDA.t406 GNDA 0.454395f
C2504 VDDA.t87 GNDA 0.478332f
C2505 VDDA.t183 GNDA 0.480066f
C2506 VDDA.t23 GNDA 0.454395f
C2507 VDDA.t22 GNDA 0.478332f
C2508 VDDA.t109 GNDA 0.480066f
C2509 VDDA.t121 GNDA 0.454395f
C2510 VDDA.t64 GNDA 0.478332f
C2511 VDDA.t178 GNDA 0.480066f
C2512 VDDA.t43 GNDA 0.454395f
C2513 VDDA.t394 GNDA 0.478332f
C2514 VDDA.t407 GNDA 0.480066f
C2515 VDDA.t182 GNDA 0.454395f
C2516 VDDA.n126 GNDA 0.320627f
C2517 VDDA.t395 GNDA 0.255332f
C2518 VDDA.n127 GNDA 0.347887f
C2519 VDDA.t181 GNDA 0.255332f
C2520 VDDA.n128 GNDA 0.347887f
C2521 VDDA.t24 GNDA 0.255332f
C2522 VDDA.n129 GNDA 0.347887f
C2523 VDDA.t63 GNDA 0.255332f
C2524 VDDA.n130 GNDA 0.347887f
C2525 VDDA.t28 GNDA 0.447299f
C2526 VDDA.n131 GNDA 3.97243f
C2527 VDDA.t413 GNDA 1.0849f
C2528 VDDA.t415 GNDA 1.08296f
C2529 VDDA.n132 GNDA 0.231496f
C2530 VDDA.t414 GNDA 1.08311f
C2531 VDDA.n133 GNDA 0.147379f
C2532 VDDA.t412 GNDA 1.08311f
C2533 VDDA.n134 GNDA 0.232411f
C2534 VDDA.n135 GNDA 0.870778f
C2535 VDDA.n136 GNDA 0.021559f
C2536 VDDA.n137 GNDA 0.087114f
C2537 VDDA.t296 GNDA 0.03118f
C2538 VDDA.n138 GNDA 0.021559f
C2539 VDDA.n139 GNDA 0.087114f
C2540 VDDA.t285 GNDA 0.03118f
C2541 VDDA.n140 GNDA 0.021559f
C2542 VDDA.n141 GNDA 0.087114f
C2543 VDDA.n142 GNDA 0.021559f
C2544 VDDA.n143 GNDA 0.087114f
C2545 VDDA.n144 GNDA 0.021559f
C2546 VDDA.n145 GNDA 0.087114f
C2547 VDDA.n146 GNDA 0.021559f
C2548 VDDA.n147 GNDA 0.087114f
C2549 VDDA.n148 GNDA 0.021559f
C2550 VDDA.n149 GNDA 0.087114f
C2551 VDDA.n150 GNDA 0.021559f
C2552 VDDA.n151 GNDA 0.087114f
C2553 VDDA.n152 GNDA 0.021559f
C2554 VDDA.n153 GNDA 0.087114f
C2555 VDDA.n154 GNDA 0.021559f
C2556 VDDA.n155 GNDA 0.141816f
C2557 VDDA.t262 GNDA 0.032106f
C2558 VDDA.n156 GNDA 0.020661f
C2559 VDDA.t264 GNDA 0.03118f
C2560 VDDA.n157 GNDA 0.114786f
C2561 VDDA.t263 GNDA 0.098256f
C2562 VDDA.t133 GNDA 0.071878f
C2563 VDDA.t172 GNDA 0.071878f
C2564 VDDA.t9 GNDA 0.071878f
C2565 VDDA.t131 GNDA 0.071878f
C2566 VDDA.t382 GNDA 0.071878f
C2567 VDDA.t88 GNDA 0.071878f
C2568 VDDA.t105 GNDA 0.071878f
C2569 VDDA.t126 GNDA 0.071878f
C2570 VDDA.t147 GNDA 0.071878f
C2571 VDDA.t145 GNDA 0.071878f
C2572 VDDA.t59 GNDA 0.071878f
C2573 VDDA.t149 GNDA 0.071878f
C2574 VDDA.t174 GNDA 0.071878f
C2575 VDDA.t400 GNDA 0.071878f
C2576 VDDA.t388 GNDA 0.071878f
C2577 VDDA.t380 GNDA 0.071878f
C2578 VDDA.t57 GNDA 0.071878f
C2579 VDDA.t396 GNDA 0.071878f
C2580 VDDA.t284 GNDA 0.099935f
C2581 VDDA.n158 GNDA 0.095579f
C2582 VDDA.t283 GNDA 0.021181f
C2583 VDDA.n159 GNDA 0.03558f
C2584 VDDA.n160 GNDA 0.063741f
C2585 VDDA.n161 GNDA 0.021559f
C2586 VDDA.n162 GNDA 0.087114f
C2587 VDDA.n163 GNDA 0.021559f
C2588 VDDA.n164 GNDA 0.087114f
C2589 VDDA.n165 GNDA 0.021559f
C2590 VDDA.n166 GNDA 0.087114f
C2591 VDDA.n167 GNDA 0.021559f
C2592 VDDA.n168 GNDA 0.087114f
C2593 VDDA.n169 GNDA 0.021559f
C2594 VDDA.n170 GNDA 0.087114f
C2595 VDDA.n171 GNDA 0.021559f
C2596 VDDA.n172 GNDA 0.087114f
C2597 VDDA.n173 GNDA 0.021559f
C2598 VDDA.n174 GNDA 0.087114f
C2599 VDDA.n175 GNDA 0.021559f
C2600 VDDA.n176 GNDA 0.087114f
C2601 VDDA.n177 GNDA 0.079981f
C2602 VDDA.t321 GNDA 0.032106f
C2603 VDDA.n178 GNDA 0.01934f
C2604 VDDA.t323 GNDA 0.03118f
C2605 VDDA.n179 GNDA 0.114786f
C2606 VDDA.t322 GNDA 0.098256f
C2607 VDDA.t76 GNDA 0.071878f
C2608 VDDA.t378 GNDA 0.071878f
C2609 VDDA.t90 GNDA 0.071878f
C2610 VDDA.t0 GNDA 0.071878f
C2611 VDDA.t94 GNDA 0.071878f
C2612 VDDA.t119 GNDA 0.071878f
C2613 VDDA.t402 GNDA 0.071878f
C2614 VDDA.t161 GNDA 0.071878f
C2615 VDDA.t72 GNDA 0.071878f
C2616 VDDA.t367 GNDA 0.071878f
C2617 VDDA.t2 GNDA 0.071878f
C2618 VDDA.t153 GNDA 0.071878f
C2619 VDDA.t390 GNDA 0.071878f
C2620 VDDA.t185 GNDA 0.071878f
C2621 VDDA.t191 GNDA 0.071878f
C2622 VDDA.t128 GNDA 0.071878f
C2623 VDDA.t140 GNDA 0.071878f
C2624 VDDA.t151 GNDA 0.071878f
C2625 VDDA.t295 GNDA 0.098256f
C2626 VDDA.n180 GNDA 0.115013f
C2627 VDDA.t294 GNDA 0.032093f
C2628 VDDA.n181 GNDA 0.019337f
C2629 VDDA.n182 GNDA 0.163967f
C2630 VDDA.n183 GNDA 0.284822f
C2631 VDDA.t243 GNDA 0.090958f
C2632 VDDA.n184 GNDA 0.25893f
C2633 VDDA.t242 GNDA 0.295166f
C2634 VDDA.t107 GNDA 0.273394f
C2635 VDDA.t176 GNDA 0.273394f
C2636 VDDA.t404 GNDA 0.273394f
C2637 VDDA.t25 GNDA 0.273394f
C2638 VDDA.t85 GNDA 0.273394f
C2639 VDDA.t83 GNDA 0.273394f
C2640 VDDA.t157 GNDA 0.273394f
C2641 VDDA.t124 GNDA 0.273394f
C2642 VDDA.t81 GNDA 0.273394f
C2643 VDDA.t155 GNDA 0.273394f
C2644 VDDA.t179 GNDA 0.273394f
C2645 VDDA.t122 GNDA 0.273394f
C2646 VDDA.t44 GNDA 0.273394f
C2647 VDDA.t61 GNDA 0.273394f
C2648 VDDA.t392 GNDA 0.273394f
C2649 VDDA.t159 GNDA 0.273394f
C2650 VDDA.t281 GNDA 0.295166f
C2651 VDDA.t282 GNDA 0.090958f
C2652 VDDA.n185 GNDA 0.25893f
C2653 VDDA.t280 GNDA 0.122409f
C2654 VDDA.t318 GNDA 0.016222f
C2655 VDDA.n186 GNDA 0.042612f
C2656 VDDA.t320 GNDA 0.03118f
C2657 VDDA.n187 GNDA 0.089664f
C2658 VDDA.t319 GNDA 0.09387f
C2659 VDDA.t19 GNDA 0.065888f
C2660 VDDA.t386 GNDA 0.065888f
C2661 VDDA.t355 GNDA 0.097272f
C2662 VDDA.t356 GNDA 0.034951f
C2663 VDDA.n188 GNDA 0.102665f
C2664 VDDA.t354 GNDA 0.016222f
C2665 VDDA.n189 GNDA 0.035693f
C2666 VDDA.n190 GNDA 0.166462f
C2667 VDDA.n191 GNDA 0.098432f
C2668 VDDA.t160 GNDA 0.025671f
C2669 VDDA.t393 GNDA 0.025671f
C2670 VDDA.n192 GNDA 0.081495f
C2671 VDDA.n193 GNDA 0.080824f
C2672 VDDA.t62 GNDA 0.025671f
C2673 VDDA.t45 GNDA 0.025671f
C2674 VDDA.n194 GNDA 0.081495f
C2675 VDDA.n195 GNDA 0.080231f
C2676 VDDA.t123 GNDA 0.025671f
C2677 VDDA.t180 GNDA 0.025671f
C2678 VDDA.n196 GNDA 0.081495f
C2679 VDDA.n197 GNDA 0.080231f
C2680 VDDA.t156 GNDA 0.025671f
C2681 VDDA.t82 GNDA 0.025671f
C2682 VDDA.n198 GNDA 0.081495f
C2683 VDDA.n199 GNDA 0.080231f
C2684 VDDA.t125 GNDA 0.025671f
C2685 VDDA.t158 GNDA 0.025671f
C2686 VDDA.n200 GNDA 0.081495f
C2687 VDDA.n201 GNDA 0.080231f
C2688 VDDA.t84 GNDA 0.025671f
C2689 VDDA.t86 GNDA 0.025671f
C2690 VDDA.n202 GNDA 0.081495f
C2691 VDDA.n203 GNDA 0.080231f
C2692 VDDA.t26 GNDA 0.025671f
C2693 VDDA.t405 GNDA 0.025671f
C2694 VDDA.n204 GNDA 0.081495f
C2695 VDDA.n205 GNDA 0.080231f
C2696 VDDA.t177 GNDA 0.025671f
C2697 VDDA.t108 GNDA 0.025671f
C2698 VDDA.n206 GNDA 0.081495f
C2699 VDDA.n207 GNDA 0.080824f
C2700 VDDA.t241 GNDA 0.122409f
C2701 VDDA.n208 GNDA 0.10146f
C2702 VDDA.n209 GNDA 0.074152f
C2703 VDDA.t252 GNDA 0.061056f
C2704 VDDA.t250 GNDA 0.024614f
C2705 VDDA.n210 GNDA 0.04832f
C2706 VDDA.n211 GNDA 0.167065f
C2707 VDDA.t251 GNDA 0.151213f
C2708 VDDA.t20 GNDA 0.112951f
C2709 VDDA.t337 GNDA 0.151213f
C2710 VDDA.t336 GNDA 0.025195f
C2711 VDDA.n212 GNDA 0.048391f
C2712 VDDA.n213 GNDA 0.167065f
C2713 VDDA.t338 GNDA 0.07817f
C2714 VDDA.t21 GNDA 0.017114f
C2715 VDDA.n214 GNDA 0.050879f
C2716 VDDA.n215 GNDA 0.079231f
C2717 VDDA.n216 GNDA 0.214111f
C2718 VDDA.n217 GNDA 0.232385f
C2719 VDDA.n218 GNDA 0.021345f
C2720 VDDA.n219 GNDA 0.075348f
C2721 VDDA.t335 GNDA 0.031197f
C2722 VDDA.t267 GNDA 0.031197f
C2723 VDDA.t265 GNDA 0.016852f
C2724 VDDA.t360 GNDA 0.017114f
C2725 VDDA.t288 GNDA 0.017114f
C2726 VDDA.n220 GNDA 0.052365f
C2727 VDDA.n221 GNDA 0.083262f
C2728 VDDA.t289 GNDA 0.061056f
C2729 VDDA.t348 GNDA 0.025868f
C2730 VDDA.n222 GNDA 0.049999f
C2731 VDDA.t362 GNDA 0.017114f
C2732 VDDA.n223 GNDA 0.021354f
C2733 VDDA.n224 GNDA 0.075339f
C2734 VDDA.t249 GNDA 0.031213f
C2735 VDDA.t332 GNDA 0.031213f
C2736 VDDA.t330 GNDA 0.016852f
C2737 VDDA.n225 GNDA 0.021354f
C2738 VDDA.n226 GNDA 0.102056f
C2739 VDDA.t344 GNDA 0.031213f
C2740 VDDA.t308 GNDA 0.031213f
C2741 VDDA.t306 GNDA 0.016852f
C2742 VDDA.n227 GNDA 0.035565f
C2743 VDDA.n228 GNDA 0.089072f
C2744 VDDA.t307 GNDA 0.09387f
C2745 VDDA.t365 GNDA 0.065888f
C2746 VDDA.t79 GNDA 0.065888f
C2747 VDDA.t343 GNDA 0.09387f
C2748 VDDA.n229 GNDA 0.089072f
C2749 VDDA.t342 GNDA 0.016852f
C2750 VDDA.n230 GNDA 0.034658f
C2751 VDDA.n231 GNDA 0.056718f
C2752 VDDA.n232 GNDA 0.021354f
C2753 VDDA.n233 GNDA 0.075339f
C2754 VDDA.n234 GNDA 0.055434f
C2755 VDDA.n235 GNDA 0.034658f
C2756 VDDA.n236 GNDA 0.089072f
C2757 VDDA.t331 GNDA 0.09387f
C2758 VDDA.t99 GNDA 0.065888f
C2759 VDDA.t74 GNDA 0.065888f
C2760 VDDA.t408 GNDA 0.065888f
C2761 VDDA.t41 GNDA 0.065888f
C2762 VDDA.t248 GNDA 0.09387f
C2763 VDDA.n237 GNDA 0.089072f
C2764 VDDA.t247 GNDA 0.017386f
C2765 VDDA.n238 GNDA 0.035193f
C2766 VDDA.n239 GNDA 0.065274f
C2767 VDDA.n240 GNDA 0.061424f
C2768 VDDA.t143 GNDA 0.017114f
C2769 VDDA.t358 GNDA 0.017114f
C2770 VDDA.n241 GNDA 0.052365f
C2771 VDDA.n242 GNDA 0.087113f
C2772 VDDA.n243 GNDA 0.083262f
C2773 VDDA.n244 GNDA 0.052365f
C2774 VDDA.t350 GNDA 0.07817f
C2775 VDDA.n245 GNDA 0.167065f
C2776 VDDA.t349 GNDA 0.151213f
C2777 VDDA.t361 GNDA 0.112951f
C2778 VDDA.t142 GNDA 0.112951f
C2779 VDDA.t357 GNDA 0.112951f
C2780 VDDA.t359 GNDA 0.112951f
C2781 VDDA.t287 GNDA 0.151213f
C2782 VDDA.n246 GNDA 0.167065f
C2783 VDDA.t286 GNDA 0.025868f
C2784 VDDA.n247 GNDA 0.049999f
C2785 VDDA.n248 GNDA 0.061424f
C2786 VDDA.n249 GNDA 0.021345f
C2787 VDDA.n250 GNDA 0.075348f
C2788 VDDA.n251 GNDA 0.065274f
C2789 VDDA.n252 GNDA 0.034658f
C2790 VDDA.n253 GNDA 0.089088f
C2791 VDDA.t266 GNDA 0.09387f
C2792 VDDA.t163 GNDA 0.065888f
C2793 VDDA.t363 GNDA 0.065888f
C2794 VDDA.t193 GNDA 0.065888f
C2795 VDDA.t6 GNDA 0.065888f
C2796 VDDA.t334 GNDA 0.09387f
C2797 VDDA.n254 GNDA 0.089088f
C2798 VDDA.t333 GNDA 0.016852f
C2799 VDDA.n255 GNDA 0.034658f
C2800 VDDA.n256 GNDA 0.173039f
C2801 VDDA.n257 GNDA 0.202015f
C2802 VDDA.n258 GNDA 0.963064f
C2803 two_stage_opamp_dummy_magic_19_0.Vb3.t3 GNDA 0.014009f
C2804 two_stage_opamp_dummy_magic_19_0.Vb3.t7 GNDA 0.014009f
C2805 two_stage_opamp_dummy_magic_19_0.Vb3.n0 GNDA 0.044923f
C2806 two_stage_opamp_dummy_magic_19_0.Vb3.t5 GNDA 0.014009f
C2807 two_stage_opamp_dummy_magic_19_0.Vb3.t0 GNDA 0.014009f
C2808 two_stage_opamp_dummy_magic_19_0.Vb3.n1 GNDA 0.044923f
C2809 two_stage_opamp_dummy_magic_19_0.Vb3.n2 GNDA 0.249171f
C2810 two_stage_opamp_dummy_magic_19_0.Vb3.t6 GNDA 0.014009f
C2811 two_stage_opamp_dummy_magic_19_0.Vb3.t4 GNDA 0.014009f
C2812 two_stage_opamp_dummy_magic_19_0.Vb3.n3 GNDA 0.042218f
C2813 two_stage_opamp_dummy_magic_19_0.Vb3.n4 GNDA 0.753572f
C2814 two_stage_opamp_dummy_magic_19_0.Vb3.t2 GNDA 0.049031f
C2815 two_stage_opamp_dummy_magic_19_0.Vb3.t1 GNDA 0.049031f
C2816 two_stage_opamp_dummy_magic_19_0.Vb3.n5 GNDA 0.133207f
C2817 two_stage_opamp_dummy_magic_19_0.Vb3.t13 GNDA 0.069344f
C2818 two_stage_opamp_dummy_magic_19_0.Vb3.t25 GNDA 0.069344f
C2819 two_stage_opamp_dummy_magic_19_0.Vb3.t28 GNDA 0.080023f
C2820 two_stage_opamp_dummy_magic_19_0.Vb3.n6 GNDA 0.06497f
C2821 two_stage_opamp_dummy_magic_19_0.Vb3.n7 GNDA 0.039149f
C2822 two_stage_opamp_dummy_magic_19_0.Vb3.t20 GNDA 0.069344f
C2823 two_stage_opamp_dummy_magic_19_0.Vb3.t24 GNDA 0.069344f
C2824 two_stage_opamp_dummy_magic_19_0.Vb3.t22 GNDA 0.069344f
C2825 two_stage_opamp_dummy_magic_19_0.Vb3.t27 GNDA 0.069344f
C2826 two_stage_opamp_dummy_magic_19_0.Vb3.t9 GNDA 0.069344f
C2827 two_stage_opamp_dummy_magic_19_0.Vb3.t11 GNDA 0.080023f
C2828 two_stage_opamp_dummy_magic_19_0.Vb3.n8 GNDA 0.06497f
C2829 two_stage_opamp_dummy_magic_19_0.Vb3.n9 GNDA 0.039926f
C2830 two_stage_opamp_dummy_magic_19_0.Vb3.n10 GNDA 0.039926f
C2831 two_stage_opamp_dummy_magic_19_0.Vb3.n11 GNDA 0.039926f
C2832 two_stage_opamp_dummy_magic_19_0.Vb3.n12 GNDA 0.039149f
C2833 two_stage_opamp_dummy_magic_19_0.Vb3.t16 GNDA 0.071796f
C2834 two_stage_opamp_dummy_magic_19_0.Vb3.n13 GNDA 0.073333f
C2835 two_stage_opamp_dummy_magic_19_0.Vb3.t8 GNDA 0.069344f
C2836 two_stage_opamp_dummy_magic_19_0.Vb3.t26 GNDA 0.069344f
C2837 two_stage_opamp_dummy_magic_19_0.Vb3.t21 GNDA 0.069344f
C2838 two_stage_opamp_dummy_magic_19_0.Vb3.t17 GNDA 0.069344f
C2839 two_stage_opamp_dummy_magic_19_0.Vb3.t19 GNDA 0.069344f
C2840 two_stage_opamp_dummy_magic_19_0.Vb3.t15 GNDA 0.080023f
C2841 two_stage_opamp_dummy_magic_19_0.Vb3.n14 GNDA 0.06497f
C2842 two_stage_opamp_dummy_magic_19_0.Vb3.n15 GNDA 0.039926f
C2843 two_stage_opamp_dummy_magic_19_0.Vb3.n16 GNDA 0.039926f
C2844 two_stage_opamp_dummy_magic_19_0.Vb3.n17 GNDA 0.039926f
C2845 two_stage_opamp_dummy_magic_19_0.Vb3.n18 GNDA 0.039149f
C2846 two_stage_opamp_dummy_magic_19_0.Vb3.t14 GNDA 0.069344f
C2847 two_stage_opamp_dummy_magic_19_0.Vb3.t18 GNDA 0.069344f
C2848 two_stage_opamp_dummy_magic_19_0.Vb3.t23 GNDA 0.080023f
C2849 two_stage_opamp_dummy_magic_19_0.Vb3.n19 GNDA 0.06497f
C2850 two_stage_opamp_dummy_magic_19_0.Vb3.n20 GNDA 0.039149f
C2851 two_stage_opamp_dummy_magic_19_0.Vb3.t10 GNDA 0.071796f
C2852 two_stage_opamp_dummy_magic_19_0.Vb3.n21 GNDA 0.07397f
C2853 two_stage_opamp_dummy_magic_19_0.Vb3.n22 GNDA 1.13237f
C2854 two_stage_opamp_dummy_magic_19_0.Vb3.t12 GNDA 0.085002f
C2855 two_stage_opamp_dummy_magic_19_0.Vb3.n23 GNDA 0.295485f
C2856 two_stage_opamp_dummy_magic_19_0.Vb3.n24 GNDA 1.03141f
C2857 bgr_9_0.VB3_CUR_BIAS GNDA 1.56776f
C2858 bgr_9_0.NFET_GATE_10uA.t0 GNDA 0.01675f
C2859 bgr_9_0.NFET_GATE_10uA.t2 GNDA 0.01675f
C2860 bgr_9_0.NFET_GATE_10uA.n0 GNDA 0.047154f
C2861 bgr_9_0.NFET_GATE_10uA.t18 GNDA 0.016332f
C2862 bgr_9_0.NFET_GATE_10uA.t6 GNDA 0.016332f
C2863 bgr_9_0.NFET_GATE_10uA.t14 GNDA 0.016332f
C2864 bgr_9_0.NFET_GATE_10uA.t19 GNDA 0.016332f
C2865 bgr_9_0.NFET_GATE_10uA.t5 GNDA 0.016332f
C2866 bgr_9_0.NFET_GATE_10uA.t13 GNDA 0.016332f
C2867 bgr_9_0.NFET_GATE_10uA.t12 GNDA 0.024143f
C2868 bgr_9_0.NFET_GATE_10uA.n1 GNDA 0.029878f
C2869 bgr_9_0.NFET_GATE_10uA.n2 GNDA 0.021357f
C2870 bgr_9_0.NFET_GATE_10uA.n3 GNDA 0.018081f
C2871 bgr_9_0.NFET_GATE_10uA.t15 GNDA 0.016332f
C2872 bgr_9_0.NFET_GATE_10uA.t8 GNDA 0.016332f
C2873 bgr_9_0.NFET_GATE_10uA.t21 GNDA 0.016332f
C2874 bgr_9_0.NFET_GATE_10uA.t16 GNDA 0.024143f
C2875 bgr_9_0.NFET_GATE_10uA.n4 GNDA 0.029878f
C2876 bgr_9_0.NFET_GATE_10uA.n5 GNDA 0.021357f
C2877 bgr_9_0.NFET_GATE_10uA.n6 GNDA 0.018081f
C2878 bgr_9_0.NFET_GATE_10uA.t20 GNDA 0.016332f
C2879 bgr_9_0.NFET_GATE_10uA.t7 GNDA 0.024143f
C2880 bgr_9_0.NFET_GATE_10uA.n7 GNDA 0.026602f
C2881 bgr_9_0.NFET_GATE_10uA.n8 GNDA 0.029239f
C2882 bgr_9_0.NFET_GATE_10uA.t11 GNDA 0.016332f
C2883 bgr_9_0.NFET_GATE_10uA.t22 GNDA 0.024143f
C2884 bgr_9_0.NFET_GATE_10uA.n9 GNDA 0.026602f
C2885 bgr_9_0.NFET_GATE_10uA.t9 GNDA 0.016332f
C2886 bgr_9_0.NFET_GATE_10uA.t17 GNDA 0.016332f
C2887 bgr_9_0.NFET_GATE_10uA.t23 GNDA 0.016332f
C2888 bgr_9_0.NFET_GATE_10uA.t10 GNDA 0.024143f
C2889 bgr_9_0.NFET_GATE_10uA.n10 GNDA 0.029878f
C2890 bgr_9_0.NFET_GATE_10uA.n11 GNDA 0.021357f
C2891 bgr_9_0.NFET_GATE_10uA.n12 GNDA 0.018081f
C2892 bgr_9_0.NFET_GATE_10uA.n13 GNDA 0.029239f
C2893 bgr_9_0.NFET_GATE_10uA.n14 GNDA 0.67829f
C2894 bgr_9_0.NFET_GATE_10uA.n15 GNDA 0.024928f
C2895 bgr_9_0.NFET_GATE_10uA.n16 GNDA 0.018081f
C2896 bgr_9_0.NFET_GATE_10uA.n17 GNDA 0.021357f
C2897 bgr_9_0.NFET_GATE_10uA.n18 GNDA 0.029878f
C2898 bgr_9_0.NFET_GATE_10uA.t1 GNDA 0.038251f
C2899 bgr_9_0.NFET_GATE_10uA.n19 GNDA 0.366443f
C2900 bgr_9_0.NFET_GATE_10uA.t3 GNDA 0.01675f
C2901 bgr_9_0.NFET_GATE_10uA.t4 GNDA 0.01675f
C2902 bgr_9_0.NFET_GATE_10uA.n20 GNDA 0.069531f
.ends

