** sch_path: /foss/designs/my_design/projects/ASU/EEE572/schematic/tb_OPAMP_OL_AC_3.sch
**.subckt tb_OPAMP_OL_AC_3
V1 VDD GND 1.8
V2 VIN_P DC_BIAS 0 AC 1
V3 DC_BIAS GND 0.7
C1 AMP_OUT GND 1p m=1
C2 net1 GND 1Meg m=1
L6 AMP_OUT net1 100Meg m=1
x2 VDD AMP_OUT net1 VIN_P GND opamp_bandgap_5
**** begin user architecture code
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt



.options method=gear
.options wnflag=1
.options savecurrents

.control

  * let start_DC = 0.5
  * let stop_DC = 1.3
  * dowhile start_DC <= stop_DC
    * alter V3 dc = start_DC
    save v(amp_out) v(ph(amp_out)) v(DC_BIAS) v(VIN_P)
    ac dec 20 1k 10G
    remzerovec
    * echo $&start_DC
    write tb_OPAMP_OL_AC_3.raw
    set appendwrite
    * reset
    * let start_DC = start_DC + 0.1

  * end

.endc



**** end user architecture code
**.ends

* expanding   symbol:  opamp_bandgap_5.sym # of pins=5
** sym_path: /foss/designs/my_design/projects/ASU/EEE572/schematic/opamp_bandgap_5.sym
** sch_path: /foss/designs/my_design/projects/ASU/EEE572/schematic/opamp_bandgap_5.sch
.subckt opamp_bandgap_5 VDDA Vout Vin- Vin+ GNDA
*.ipin Vin+
*.opin Vout
*.ipin Vin-
*.ipin GNDA
*.ipin VDDA
XM1 V_p V_mirror GNDA GNDA sky130_fd_pr__nfet_01v8 L=5 W=2.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 V_mirror Vin+ V_p GNDA sky130_fd_pr__nfet_01v8 L=0.5 W=12 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vout Vin- V_p GNDA sky130_fd_pr__nfet_01v8 L=0.5 W=12 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 V_mirror V_mirror VDDA VDDA sky130_fd_pr__pfet_01v8 L=0.5 W=12 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
XM6 Vout V_mirror VDDA VDDA sky130_fd_pr__pfet_01v8 L=0.5 W=12 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
.ends

.GLOBAL GND
.GLOBAL VDD
.end
