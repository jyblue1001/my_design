** sch_path: /foss/designs/my_design/projects/pll/divider/xschem_ngspice/tb_xcp_FF_divide3.sch
**.subckt tb_xcp_FF_divide3
VDD VDD GND 1.8
V3 CK GND pulse(0 1.8 0ps 8.34ps 8.34ps 200.16ps 417ps)
x1 VDD C A C CK GND xcp_FF
**** begin user architecture code



.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

.option method=gear
.option wnflag=1
* .option savecurrents

.save
+@m.x1.xm1.msky130_fd_pr__nfet_01v8[gm]
+@m.x1.xm2.msky130_fd_pr__nfet_01v8[gm]
+@m.x1.xm3.msky130_fd_pr__pfet_01v8[gm]
+@m.x1.xm4.msky130_fd_pr__pfet_01v8[gm]
+@m.x1.xm5.msky130_fd_pr__nfet_01v8[gm]
+@m.x2.xm1.msky130_fd_pr__nfet_01v8[gm]
+@m.x2.xm2.msky130_fd_pr__nfet_01v8[gm]
+@m.x2.xm3.msky130_fd_pr__pfet_01v8[gm]
+@m.x2.xm4.msky130_fd_pr__pfet_01v8[gm]
+@m.x2.xm5.msky130_fd_pr__nfet_01v8[gm]
+@v.x1.vmeas
+@v.x1.vmeas1
+@v.x1.vmeas2
+@v.x5.vmeas
+@v.x5.vmeas1
+@v.x5.vmeas2


*.ic v(b)=0

.control

  save v(a) v(a_b) v(b) v(b_b) v(c) v(ck)
  * save all
  *tran 0.1n 1u
  tran 0.2p 10n
  *ac dec 20 1 1T
  remzerovec
  write tb_xcp_FF_divide3.raw
  set appendwrite

.endc




.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/my_design/projects/pll/divider/xschem_ngspice/xcp_FF.sym # of pins=6
** sym_path: /foss/designs/my_design/projects/pll/divider/xschem_ngspice/xcp_FF.sym
** sch_path: /foss/designs/my_design/projects/pll/divider/xschem_ngspice/xcp_FF.sch
.subckt xcp_FF VDDA D Q Q_b CK GNDA
*.ipin VDDA
*.opin Q
*.ipin CK
*.ipin GNDA
*.ipin D
*.opin Q_b
x1 VDDA A_b A net1 D CK GNDA xcp_latch
x2 VDDA Q_b Q A_b A net2 GNDA xcp_latch
x3 CK VGND VNB VPB VPWR net2 sky130_fd_sc_hd__inv_1
x4 D VGND VNB VPB VPWR net1 sky130_fd_sc_hd__inv_1
.ends


* expanding   symbol:  /foss/designs/my_design/projects/pll/divider/xschem_ngspice/xcp_latch.sym # of pins=7
** sym_path: /foss/designs/my_design/projects/pll/divider/xschem_ngspice/xcp_latch.sym
** sch_path: /foss/designs/my_design/projects/pll/divider/xschem_ngspice/xcp_latch.sch
.subckt xcp_latch VDDA Q_b Q D_b D CK GNDA
*.ipin D
*.opin Q
*.ipin D_b
*.ipin CK
*.opin Q_b
*.ipin VDDA
*.ipin GNDA
XM5 net1 CK GNDA GNDA sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 net3 D V_common GNDA sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net2 D_b V_common GNDA sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vmeas V_common net1 0
.save i(vmeas)
Vmeas1 Q_b net3 0
.save i(vmeas1)
Vmeas2 Q net2 0
.save i(vmeas2)
XM3 Q_b Q VDDA VDDA sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 Q Q_b VDDA VDDA sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
