* PEX produced on Wed Jul  9 08:05:41 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr.ext - technology: sky130A

.subckt bgr VDDA ERR_AMP_REF V_CMFB_S3 VB1_CUR_BIAS TAIL_CUR_MIR_BIAS V_CMFB_S1 ERR_AMP_CUR_BIAS
+ VB3_CUR_BIAS V_CMFB_S4 V_CMFB_S2 VB2_CUR_BIAS GNDA
X0 1st_Vout_2.t11 cap_res2.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1 GNDA.t75 NFET_GATE_10uA.t5 V_CMFB_S2.t3 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X2 V_mir2.t14 V_mir2.t13 VDDA.t130 VDDA.t129 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X3 VB2_CUR_BIAS.t5 NFET_GATE_10uA.t6 GNDA.t73 GNDA.t72 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X4 a_38570_n6530.t1 a_38690_n7778.t1 GNDA.t9 sky130_fd_pr__res_xhigh_po_0p35 l=4.2
X5 GNDA.t104 GNDA.t102 V_CMFB_S2.t0 GNDA.t103 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X6 1st_Vout_1.t11 cap_res1.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 GNDA.t71 NFET_GATE_10uA.t7 V_CMFB_S4.t2 GNDA.t70 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X8 V_p_1.t10 Vin+.t6 1st_Vout_1.t8 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X9 VB2_CUR_BIAS.t4 NFET_GATE_10uA.t8 GNDA.t69 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X10 V_p_2.t4 ERR_AMP_REF.t7 V_mir2.t16 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X11 1st_Vout_1.t12 cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 GNDA.t29 START_UP_NFET1.t0 START_UP_NFET1.t1 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X13 VDDA.t178 VDDA.t176 V_CMFB_S1.t4 VDDA.t177 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X14 V_TOP.t13 START_UP.t6 Vin-.t7 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X15 V_CMFB_S3.t5 VDDA.t173 VDDA.t175 VDDA.t174 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X16 GNDA.t67 NFET_GATE_10uA.t9 VB3_CUR_BIAS.t4 GNDA.t66 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X17 VB3_CUR_BIAS.t3 NFET_GATE_10uA.t10 GNDA.t65 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X18 NFET_GATE_10uA.t0 GNDA.t99 GNDA.t101 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X19 1st_Vout_1.t13 cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 GNDA.t63 NFET_GATE_10uA.t2 NFET_GATE_10uA.t3 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X21 1st_Vout_2.t7 V_mir2.t17 VDDA.t128 VDDA.t127 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X22 V_p_1.t0 Vin-.t8 V_mir1.t16 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X23 V_p_2.t10 VDDA.t214 GNDA.t18 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X24 1st_Vout_2.t12 cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 V_CUR_REF_REG.t0 a_32320_n7778.t1 GNDA.t20 sky130_fd_pr__res_xhigh_po_0p35 l=4
X26 VB2_CUR_BIAS.t7 GNDA.t96 GNDA.t98 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X27 1st_Vout_2.t13 cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X28 1st_Vout_2.t14 cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X29 VDDA.t187 V_TOP.t14 ERR_AMP_REF.t6 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X30 1st_Vout_2.t15 cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 VDDA.t92 PFET_GATE_10uA.t10 V_CMFB_S1.t2 VDDA.t91 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X32 1st_Vout_2.t16 cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 VB2_CUR_BIAS.t3 NFET_GATE_10uA.t11 GNDA.t61 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X34 1st_Vout_1.t14 cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 VDDA.t76 PFET_GATE_10uA.t11 VB1_CUR_BIAS.t1 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X36 VDDA.t172 VDDA.t170 VB1_CUR_BIAS.t3 VDDA.t171 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X37 1st_Vout_2.t17 cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 1st_Vout_2.t18 cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 1st_Vout_1.t15 cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 VDDA.t189 V_mir1.t10 V_mir1.t11 VDDA.t188 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X41 Vin+.t3 V_TOP.t15 VDDA.t45 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X42 1st_Vout_1.t16 cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 V_TOP.t16 VDDA.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 V_mir1.t15 Vin-.t9 V_p_1.t1 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X45 1st_Vout_1.t17 cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 1st_Vout_1.t18 cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 TAIL_CUR_MIR_BIAS.t7 PFET_GATE_10uA.t12 VDDA.t31 VDDA.t30 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X48 VDDA.t126 V_mir2.t3 V_mir2.t4 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X49 V_TOP.t17 VDDA.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 ERR_AMP_REF.t4 VDDA.t167 VDDA.t169 VDDA.t168 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X51 V_mir1.t14 Vin-.t10 V_p_1.t2 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X52 1st_Vout_1.t4 V_mir1.t17 VDDA.t60 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X53 V_TOP.t18 VDDA.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X54 1st_Vout_2.t19 cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 V_CMFB_S3.t3 PFET_GATE_10uA.t13 VDDA.t100 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X56 VDDA.t22 V_TOP.t19 Vin+.t2 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X57 V_TOP.t20 VDDA.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X58 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 Vin+.t0 GNDA.t1 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X59 VDDA.t193 PFET_GATE_10uA.t14 NFET_GATE_10uA.t4 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X60 PFET_GATE_10uA.t9 1st_Vout_2.t20 VDDA.t213 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X61 1st_Vout_1.t9 Vin+.t7 V_p_1.t9 GNDA.t109 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X62 VDDA.t124 V_mir2.t18 1st_Vout_2.t0 VDDA.t123 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X63 GNDA.t95 GNDA.t93 VB3_CUR_BIAS.t5 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X64 TAIL_CUR_MIR_BIAS.t6 PFET_GATE_10uA.t15 VDDA.t49 VDDA.t48 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X65 VDDA.t211 1st_Vout_2.t21 PFET_GATE_10uA.t8 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X66 V_p_1.t8 Vin+.t8 1st_Vout_1.t10 GNDA.t111 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X67 V_CMFB_S3.t2 PFET_GATE_10uA.t16 VDDA.t66 VDDA.t65 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X68 VDDA.t166 VDDA.t164 V_TOP.t5 VDDA.t165 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X69 V_CMFB_S2.t2 NFET_GATE_10uA.t12 GNDA.t59 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X70 V_CMFB_S2.t1 NFET_GATE_10uA.t13 GNDA.t57 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X71 V_CMFB_S1.t0 PFET_GATE_10uA.t17 VDDA.t29 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X72 Vin+.t1 a_38040_n7928.t0 GNDA.t7 sky130_fd_pr__res_xhigh_po_0p35 l=6
X73 1st_Vout_1.t7 V_mir1.t18 VDDA.t104 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X74 TAIL_CUR_MIR_BIAS.t5 PFET_GATE_10uA.t18 VDDA.t24 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X75 V_mir1.t9 V_mir1.t8 VDDA.t36 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X76 V_TOP.t21 VDDA.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X77 GNDA.t105 VDDA.t215 PFET_GATE_10uA.t1 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X78 VDDA.t15 1st_Vout_1.t19 V_TOP.t11 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X79 PFET_GATE_10uA.t7 1st_Vout_2.t22 VDDA.t209 VDDA.t208 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X80 V_p_2.t3 ERR_AMP_REF.t8 V_mir2.t1 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X81 V_TOP.t1 VDDA.t216 GNDA.t106 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X82 V_TOP.t22 VDDA.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 VB3_CUR_BIAS.t2 NFET_GATE_10uA.t14 GNDA.t55 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X84 GNDA.t53 NFET_GATE_10uA.t15 ERR_AMP_CUR_BIAS.t1 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X85 VDDA.t38 V_mir1.t19 1st_Vout_1.t1 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X86 V_p_1.t7 Vin+.t9 1st_Vout_1.t2 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X87 1st_Vout_2.t23 cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 1st_Vout_2.t24 cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 V_CMFB_S1.t3 VDDA.t161 VDDA.t163 VDDA.t162 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X90 VDDA.t122 V_mir2.t19 1st_Vout_2.t9 VDDA.t121 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X91 1st_Vout_2.t25 cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X92 VDDA.t207 1st_Vout_2.t26 PFET_GATE_10uA.t6 VDDA.t206 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X93 V_p_2.t5 V_CUR_REF_REG.t3 1st_Vout_2.t2 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X94 1st_Vout_1.t20 cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 NFET_GATE_10uA.t1 VDDA.t158 VDDA.t160 VDDA.t159 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X96 TAIL_CUR_MIR_BIAS.t4 PFET_GATE_10uA.t19 VDDA.t74 VDDA.t73 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X97 V_TOP.t4 VDDA.t155 VDDA.t157 VDDA.t156 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X98 1st_Vout_2.t27 cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X99 V_CUR_REF_REG.t2 PFET_GATE_10uA.t20 VDDA.t201 VDDA.t200 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X100 1st_Vout_1.t21 cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X101 V_TOP.t23 VDDA.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X102 V_CMFB_S4.t1 NFET_GATE_10uA.t16 GNDA.t51 GNDA.t50 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X103 V_mir2.t6 V_mir2.t5 VDDA.t120 VDDA.t119 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X104 1st_Vout_1.t22 cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 GNDA.t49 NFET_GATE_10uA.t17 V_CMFB_S4.t0 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X106 1st_Vout_2.t1 V_mir2.t20 VDDA.t118 VDDA.t117 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X107 1st_Vout_1.t23 cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 GNDA.t77 GNDA.t91 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X109 V_TOP.t24 VDDA.t199 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X110 1st_Vout_2.t28 cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 Vin-.t0 a_32970_n7928.t0 GNDA.t11 sky130_fd_pr__res_xhigh_po_0p35 l=6
X112 GNDA.t77 GNDA.t90 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X113 VDDA.t154 VDDA.t152 V_TOP.t3 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=0.45 pd=2.9 as=0.2 ps=1.4 w=1 l=0.15
X114 VDDA.t52 V_TOP.t25 Vin-.t3 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X115 V_TOP.t26 VDDA.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X116 a_32440_n6570.t0 a_32320_n7778.t0 GNDA.t0 sky130_fd_pr__res_xhigh_po_0p35 l=4
X117 GNDA.t77 GNDA.t92 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X118 ERR_AMP_REF.t5 V_TOP.t27 VDDA.t182 VDDA.t181 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X119 VDDA.t84 V_mir1.t20 1st_Vout_1.t5 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X120 1st_Vout_2.t10 V_CUR_REF_REG.t4 V_p_2.t9 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X121 VDDA.t6 V_mir1.t6 V_mir1.t7 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X122 Vin+.t5 V_TOP.t28 VDDA.t185 VDDA.t184 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X123 V_mir1.t13 Vin-.t11 V_p_1.t4 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X124 V_TOP.t29 VDDA.t198 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 a_38570_n6530.t0 GNDA.t10 GNDA.t9 sky130_fd_pr__res_xhigh_po_0p35 l=4.2
X126 a_33090_n6320.t0 GNDA.t16 GNDA.t15 sky130_fd_pr__res_xhigh_po_0p35 l=6
X127 V_mir1.t5 V_mir1.t4 VDDA.t98 VDDA.t97 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X128 VDDA.t151 VDDA.t149 PFET_GATE_10uA.t3 VDDA.t150 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X129 GNDA.t14 VDDA.t217 V_p_1.t5 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X130 V_CMFB_S1.t1 PFET_GATE_10uA.t21 VDDA.t64 VDDA.t63 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X131 Vin-.t6 START_UP.t7 V_TOP.t12 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X132 V_TOP.t10 1st_Vout_1.t24 VDDA.t54 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X133 V_mir2.t15 ERR_AMP_REF.t9 V_p_2.t2 GNDA.t107 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X134 Vin-.t4 V_TOP.t30 VDDA.t57 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X135 a_37920_n6320.t0 GNDA.t8 GNDA.t7 sky130_fd_pr__res_xhigh_po_0p35 l=6
X136 V_mir2.t8 V_mir2.t7 VDDA.t116 VDDA.t115 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X137 PFET_GATE_10uA.t0 cap_res2.t0 GNDA.t12 sky130_fd_pr__res_high_po_0p35 l=2.05
X138 VDDA.t11 V_TOP.t31 START_UP.t0 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X139 1st_Vout_2.t8 V_mir2.t21 VDDA.t114 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X140 V_TOP.t32 VDDA.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X141 VDDA.t205 1st_Vout_2.t29 PFET_GATE_10uA.t5 VDDA.t204 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X142 V_TOP.t0 cap_res1.t0 GNDA.t30 sky130_fd_pr__res_high_po_0p35 l=2.05
X143 V_TOP.t33 VDDA.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 VDDA.t4 V_TOP.t34 ERR_AMP_REF.t1 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X145 VDDA.t112 V_mir2.t11 V_mir2.t12 VDDA.t111 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X146 VDDA.t90 PFET_GATE_10uA.t22 TAIL_CUR_MIR_BIAS.t3 VDDA.t89 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X147 V_TOP.t35 VDDA.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 1st_Vout_2.t30 cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 GNDA.t47 NFET_GATE_10uA.t18 VB2_CUR_BIAS.t2 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X150 V_TOP.t36 VDDA.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 VDDA.t80 V_TOP.t37 START_UP.t1 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X152 VB1_CUR_BIAS.t2 VDDA.t146 VDDA.t148 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X153 VB1_CUR_BIAS.t0 PFET_GATE_10uA.t23 VDDA.t86 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X154 GNDA.t89 GNDA.t87 VB2_CUR_BIAS.t6 GNDA.t88 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X155 VDDA.t145 VDDA.t143 V_CMFB_S3.t4 VDDA.t144 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X156 START_UP_NFET1.t1 START_UP.t4 START_UP.t5 GNDA.t110 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X157 1st_Vout_1.t25 cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 PFET_GATE_10uA.t2 VDDA.t140 VDDA.t142 VDDA.t141 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X159 1st_Vout_2.t31 cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X160 V_p_1.t3 Vin-.t12 V_mir1.t12 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X161 V_p_2.t7 V_CUR_REF_REG.t5 1st_Vout_2.t4 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X162 START_UP.t3 V_TOP.t38 VDDA.t96 VDDA.t95 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X163 1st_Vout_1.t26 cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 V_TOP.t39 VDDA.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 VB3_CUR_BIAS.t1 NFET_GATE_10uA.t19 GNDA.t45 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X166 1st_Vout_1.t27 cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X167 GNDA.t43 NFET_GATE_10uA.t20 VB3_CUR_BIAS.t0 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X168 ERR_AMP_CUR_BIAS.t0 NFET_GATE_10uA.t21 GNDA.t41 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X169 VDDA.t62 PFET_GATE_10uA.t24 TAIL_CUR_MIR_BIAS.t2 VDDA.t61 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X170 ERR_AMP_REF.t0 V_TOP.t40 VDDA.t2 VDDA.t1 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X171 V_TOP.t9 1st_Vout_1.t28 VDDA.t180 VDDA.t179 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X172 V_p_2.t1 ERR_AMP_REF.t10 V_mir2.t2 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X173 1st_Vout_1.t29 cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 1st_Vout_1.t0 V_mir1.t21 VDDA.t9 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X175 ERR_AMP_REF.t2 a_38690_n7778.t0 GNDA.t9 sky130_fd_pr__res_xhigh_po_0p35 l=4.2
X176 START_UP.t2 V_TOP.t41 VDDA.t94 VDDA.t93 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X177 VDDA.t88 V_mir1.t2 V_mir1.t3 VDDA.t87 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X178 GNDA.t39 NFET_GATE_10uA.t22 VB2_CUR_BIAS.t1 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X179 GNDA.t77 GNDA.t85 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X180 VDDA.t18 PFET_GATE_10uA.t25 V_CMFB_S3.t0 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X181 GNDA.t77 GNDA.t86 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X182 VDDA.t78 1st_Vout_1.t30 V_TOP.t8 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X183 V_TOP.t2 VDDA.t137 VDDA.t139 VDDA.t138 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X184 VDDA.t110 V_mir2.t9 V_mir2.t10 VDDA.t109 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X185 GNDA.t37 NFET_GATE_10uA.t23 VB2_CUR_BIAS.t0 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X186 V_CMFB_S4.t3 GNDA.t82 GNDA.t84 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X187 VDDA.t33 V_TOP.t42 Vin-.t1 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X188 1st_Vout_1.t31 cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 VDDA.t108 V_mir2.t22 1st_Vout_2.t6 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X190 a_33090_n6320.t1 a_32970_n7928.t1 GNDA.t34 sky130_fd_pr__res_xhigh_po_0p35 l=6
X191 GNDA.t77 GNDA.t79 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X192 VDDA.t68 PFET_GATE_10uA.t26 TAIL_CUR_MIR_BIAS.t1 VDDA.t67 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X193 VDDA.t82 V_TOP.t43 Vin+.t4 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X194 PFET_GATE_10uA.t4 1st_Vout_2.t32 VDDA.t203 VDDA.t202 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X195 1st_Vout_2.t33 cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 V_TOP.t44 VDDA.t183 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 VDDA.t40 PFET_GATE_10uA.t27 V_CMFB_S3.t1 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X198 1st_Vout_2.t34 cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 1st_Vout_1.t3 Vin+.t10 V_p_1.t6 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X200 V_mir2.t0 ERR_AMP_REF.t11 V_p_2.t0 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X201 VDDA.t191 PFET_GATE_10uA.t28 V_CMFB_S1.t5 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X202 V_TOP.t7 1st_Vout_1.t32 VDDA.t197 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X203 1st_Vout_2.t35 cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X204 Vin-.t2 V_TOP.t45 VDDA.t42 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X205 1st_Vout_1.t33 cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X206 GNDA.t77 GNDA.t76 Vin-.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X207 VDDA.t47 PFET_GATE_10uA.t29 TAIL_CUR_MIR_BIAS.t0 VDDA.t46 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X208 VDDA.t136 VDDA.t134 V_CUR_REF_REG.t1 VDDA.t135 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X209 1st_Vout_2.t3 V_CUR_REF_REG.t6 V_p_2.t6 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X210 1st_Vout_1.t34 cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 1st_Vout_1.t35 cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 a_37920_n6320.t1 a_38040_n7928.t1 GNDA.t7 sky130_fd_pr__res_xhigh_po_0p35 l=6
X213 GNDA.t81 GNDA.t80 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X214 VDDA.t195 1st_Vout_1.t36 V_TOP.t6 VDDA.t194 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X215 V_TOP.t46 VDDA.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 1st_Vout_2.t5 V_CUR_REF_REG.t7 V_p_2.t8 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X217 VDDA.t133 VDDA.t131 ERR_AMP_REF.t3 VDDA.t132 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X218 VDDA.t102 V_mir1.t22 1st_Vout_1.t6 VDDA.t101 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X219 V_TOP.t47 VDDA.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X220 GNDA.t77 GNDA.t78 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X221 V_TOP.t48 VDDA.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 1st_Vout_2.t36 cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 a_32440_n6570.t1 GNDA.t6 GNDA.t5 sky130_fd_pr__res_xhigh_po_0p35 l=4
X224 V_TOP.t49 VDDA.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X225 V_mir1.t1 V_mir1.t0 VDDA.t106 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
R0 1st_Vout_2 1st_Vout_2.t29 354.854
R1 1st_Vout_2.n0 1st_Vout_2.t22 346.8
R2 1st_Vout_2 1st_Vout_2.n11 339.522
R3 1st_Vout_2.n0 1st_Vout_2.n4 339.522
R4 1st_Vout_2.n2 1st_Vout_2.n6 335.022
R5 1st_Vout_2.n8 1st_Vout_2.t3 275.909
R6 1st_Vout_2.n8 1st_Vout_2.n7 227.909
R7 1st_Vout_2.n2 1st_Vout_2.n9 222.034
R8 1st_Vout_2.n10 1st_Vout_2.t32 184.097
R9 1st_Vout_2.n10 1st_Vout_2.t21 184.097
R10 1st_Vout_2.n5 1st_Vout_2.t20 184.097
R11 1st_Vout_2.n5 1st_Vout_2.t26 184.097
R12 1st_Vout_2 1st_Vout_2.n10 166.05
R13 1st_Vout_2.n0 1st_Vout_2.n5 166.05
R14 1st_Vout_2.n0 1st_Vout_2.n3 52.9634
R15 1st_Vout_2.n9 1st_Vout_2.t2 48.0005
R16 1st_Vout_2.n9 1st_Vout_2.t5 48.0005
R17 1st_Vout_2.n7 1st_Vout_2.t4 48.0005
R18 1st_Vout_2.n7 1st_Vout_2.t10 48.0005
R19 1st_Vout_2.n6 1st_Vout_2.t9 39.4005
R20 1st_Vout_2.n6 1st_Vout_2.t1 39.4005
R21 1st_Vout_2.n4 1st_Vout_2.t6 39.4005
R22 1st_Vout_2.n4 1st_Vout_2.t8 39.4005
R23 1st_Vout_2.n11 1st_Vout_2.t0 39.4005
R24 1st_Vout_2.n11 1st_Vout_2.t7 39.4005
R25 1st_Vout_2 1st_Vout_2.n0 5.6255
R26 1st_Vout_2 1st_Vout_2.n2 5.28175
R27 1st_Vout_2.n1 1st_Vout_2.t27 4.8295
R28 1st_Vout_2.n1 1st_Vout_2.t11 4.8295
R29 1st_Vout_2.n1 1st_Vout_2.t18 4.8295
R30 1st_Vout_2.n1 1st_Vout_2.t31 4.8295
R31 1st_Vout_2.n1 1st_Vout_2.t35 4.8295
R32 1st_Vout_2.n1 1st_Vout_2.t24 4.8295
R33 1st_Vout_2.n3 1st_Vout_2.t16 4.8295
R34 1st_Vout_2.n3 1st_Vout_2.t30 4.8295
R35 1st_Vout_2.n3 1st_Vout_2.t28 4.8295
R36 1st_Vout_2.n2 1st_Vout_2.n8 4.5005
R37 1st_Vout_2.n1 1st_Vout_2.t25 4.5005
R38 1st_Vout_2.n1 1st_Vout_2.t23 4.5005
R39 1st_Vout_2.n1 1st_Vout_2.t17 4.5005
R40 1st_Vout_2.n1 1st_Vout_2.t15 4.5005
R41 1st_Vout_2.n1 1st_Vout_2.t34 4.5005
R42 1st_Vout_2.n1 1st_Vout_2.t33 4.5005
R43 1st_Vout_2.n3 1st_Vout_2.t13 4.5005
R44 1st_Vout_2.n3 1st_Vout_2.t12 4.5005
R45 1st_Vout_2.n3 1st_Vout_2.t19 4.5005
R46 1st_Vout_2.n3 1st_Vout_2.t36 4.5005
R47 1st_Vout_2.n3 1st_Vout_2.t14 4.5005
R48 1st_Vout_2.n3 1st_Vout_2.n1 3.1025
R49 cap_res2 cap_res2.t0 121.05
R50 cap_res2 cap_res2.t12 0.194375
R51 cap_res2.t1 cap_res2.t17 0.1603
R52 cap_res2.t19 cap_res2.t6 0.1603
R53 cap_res2.t4 cap_res2.t10 0.1603
R54 cap_res2.t16 cap_res2.t5 0.1603
R55 cap_res2.t11 cap_res2.t20 0.1603
R56 cap_res2.n1 cap_res2.t9 0.159278
R57 cap_res2.n2 cap_res2.t14 0.159278
R58 cap_res2.n3 cap_res2.t3 0.159278
R59 cap_res2.n4 cap_res2.t18 0.159278
R60 cap_res2.n4 cap_res2.t1 0.1368
R61 cap_res2.n4 cap_res2.t7 0.1368
R62 cap_res2.n3 cap_res2.t19 0.1368
R63 cap_res2.n3 cap_res2.t15 0.1368
R64 cap_res2.n2 cap_res2.t4 0.1368
R65 cap_res2.n2 cap_res2.t2 0.1368
R66 cap_res2.n1 cap_res2.t16 0.1368
R67 cap_res2.n1 cap_res2.t13 0.1368
R68 cap_res2.n0 cap_res2.t11 0.1368
R69 cap_res2.n0 cap_res2.t8 0.1368
R70 cap_res2.t9 cap_res2.n0 0.00152174
R71 cap_res2.t14 cap_res2.n1 0.00152174
R72 cap_res2.t3 cap_res2.n2 0.00152174
R73 cap_res2.t18 cap_res2.n3 0.00152174
R74 cap_res2.t12 cap_res2.n4 0.00152174
R75 NFET_GATE_10uA.n19 NFET_GATE_10uA.n0 397.197
R76 NFET_GATE_10uA.n19 NFET_GATE_10uA.t2 384.967
R77 NFET_GATE_10uA.n10 NFET_GATE_10uA.t22 369.534
R78 NFET_GATE_10uA.n9 NFET_GATE_10uA.t13 369.534
R79 NFET_GATE_10uA.n7 NFET_GATE_10uA.t17 369.534
R80 NFET_GATE_10uA.n4 NFET_GATE_10uA.t8 369.534
R81 NFET_GATE_10uA.n1 NFET_GATE_10uA.t19 369.534
R82 NFET_GATE_10uA.t2 NFET_GATE_10uA.n18 369.534
R83 NFET_GATE_10uA.n10 NFET_GATE_10uA.t12 192.8
R84 NFET_GATE_10uA.n11 NFET_GATE_10uA.t5 192.8
R85 NFET_GATE_10uA.n12 NFET_GATE_10uA.t6 192.8
R86 NFET_GATE_10uA.n9 NFET_GATE_10uA.t18 192.8
R87 NFET_GATE_10uA.n7 NFET_GATE_10uA.t11 192.8
R88 NFET_GATE_10uA.n6 NFET_GATE_10uA.t23 192.8
R89 NFET_GATE_10uA.n5 NFET_GATE_10uA.t16 192.8
R90 NFET_GATE_10uA.n4 NFET_GATE_10uA.t7 192.8
R91 NFET_GATE_10uA.n3 NFET_GATE_10uA.t20 192.8
R92 NFET_GATE_10uA.n2 NFET_GATE_10uA.t14 192.8
R93 NFET_GATE_10uA.n1 NFET_GATE_10uA.t9 192.8
R94 NFET_GATE_10uA.n18 NFET_GATE_10uA.t21 192.8
R95 NFET_GATE_10uA.n17 NFET_GATE_10uA.t15 192.8
R96 NFET_GATE_10uA.n16 NFET_GATE_10uA.t10 192.8
R97 NFET_GATE_10uA.n12 NFET_GATE_10uA.n11 176.733
R98 NFET_GATE_10uA.n11 NFET_GATE_10uA.n10 176.733
R99 NFET_GATE_10uA.n5 NFET_GATE_10uA.n4 176.733
R100 NFET_GATE_10uA.n6 NFET_GATE_10uA.n5 176.733
R101 NFET_GATE_10uA.n2 NFET_GATE_10uA.n1 176.733
R102 NFET_GATE_10uA.n3 NFET_GATE_10uA.n2 176.733
R103 NFET_GATE_10uA.n17 NFET_GATE_10uA.n16 176.733
R104 NFET_GATE_10uA.n18 NFET_GATE_10uA.n17 176.733
R105 NFET_GATE_10uA.n14 NFET_GATE_10uA.n13 169.852
R106 NFET_GATE_10uA.n14 NFET_GATE_10uA.n8 169.852
R107 NFET_GATE_10uA.n15 NFET_GATE_10uA.n14 166.133
R108 NFET_GATE_10uA.n20 NFET_GATE_10uA.n19 126.876
R109 NFET_GATE_10uA.n13 NFET_GATE_10uA.n12 56.2338
R110 NFET_GATE_10uA.n13 NFET_GATE_10uA.n9 56.2338
R111 NFET_GATE_10uA.n8 NFET_GATE_10uA.n7 56.2338
R112 NFET_GATE_10uA.n8 NFET_GATE_10uA.n6 56.2338
R113 NFET_GATE_10uA.n15 NFET_GATE_10uA.n3 56.2338
R114 NFET_GATE_10uA.n16 NFET_GATE_10uA.n15 56.2338
R115 NFET_GATE_10uA.n0 NFET_GATE_10uA.t4 39.4005
R116 NFET_GATE_10uA.n0 NFET_GATE_10uA.t1 39.4005
R117 NFET_GATE_10uA.n20 NFET_GATE_10uA.t3 24.0005
R118 NFET_GATE_10uA.t0 NFET_GATE_10uA.n20 24.0005
R119 V_CMFB_S2.n2 V_CMFB_S2.n0 144.827
R120 V_CMFB_S2.n2 V_CMFB_S2.n1 134.577
R121 V_CMFB_S2 V_CMFB_S2.n2 37.563
R122 V_CMFB_S2.n1 V_CMFB_S2.t3 24.0005
R123 V_CMFB_S2.n1 V_CMFB_S2.t2 24.0005
R124 V_CMFB_S2.n0 V_CMFB_S2.t0 24.0005
R125 V_CMFB_S2.n0 V_CMFB_S2.t1 24.0005
R126 GNDA.n2035 GNDA.n2034 9343.35
R127 GNDA.n2035 GNDA.n16 9291.68
R128 GNDA.n2037 GNDA.n2035 8202.33
R129 GNDA.n1363 GNDA.n1207 1367.21
R130 GNDA.n2034 GNDA.t13 1311.87
R131 GNDA.n1819 GNDA.n1816 1185.07
R132 GNDA.n1819 GNDA.n1818 1185.07
R133 GNDA.n1496 GNDA.n16 1104.89
R134 GNDA.n1829 GNDA.n1828 686.717
R135 GNDA.n1617 GNDA.n1616 686.717
R136 GNDA.n1613 GNDA.n1602 686.717
R137 GNDA.n1821 GNDA.n192 686.717
R138 GNDA.n211 GNDA.n207 669.307
R139 GNDA.n1496 GNDA.n1495 585.003
R140 GNDA.n1701 GNDA.n1700 585.001
R141 GNDA.n1722 GNDA.n1721 585.001
R142 GNDA.n1716 GNDA.n199 585.001
R143 GNDA.n1919 GNDA.n1918 585.001
R144 GNDA.n1913 GNDA.n1912 585.001
R145 GNDA.n137 GNDA.n17 585.001
R146 GNDA.n935 GNDA.n20 585
R147 GNDA.n959 GNDA.n808 585
R148 GNDA.n957 GNDA.n956 585
R149 GNDA.n955 GNDA.n810 585
R150 GNDA.n954 GNDA.n953 585
R151 GNDA.n951 GNDA.n811 585
R152 GNDA.n949 GNDA.n948 585
R153 GNDA.n947 GNDA.n812 585
R154 GNDA.n946 GNDA.n945 585
R155 GNDA.n943 GNDA.n813 585
R156 GNDA.n941 GNDA.n940 585
R157 GNDA.n939 GNDA.n814 585
R158 GNDA.n2012 GNDA.n2011 585
R159 GNDA.n2013 GNDA.n27 585
R160 GNDA.n2015 GNDA.n2014 585
R161 GNDA.n2017 GNDA.n25 585
R162 GNDA.n2019 GNDA.n2018 585
R163 GNDA.n2020 GNDA.n24 585
R164 GNDA.n2022 GNDA.n2021 585
R165 GNDA.n2024 GNDA.n22 585
R166 GNDA.n2026 GNDA.n2025 585
R167 GNDA.n2027 GNDA.n21 585
R168 GNDA.n2029 GNDA.n2028 585
R169 GNDA.n1342 GNDA.n1341 585
R170 GNDA.n1341 GNDA.n1340 585
R171 GNDA.n1342 GNDA.n1218 585
R172 GNDA.n1218 GNDA.n1217 585
R173 GNDA.n1344 GNDA.n1343 585
R174 GNDA.n1345 GNDA.n1344 585
R175 GNDA.n1216 GNDA.n1215 585
R176 GNDA.n1346 GNDA.n1216 585
R177 GNDA.n1350 GNDA.n1349 585
R178 GNDA.n1349 GNDA.n1348 585
R179 GNDA.n1351 GNDA.n1214 585
R180 GNDA.n1347 GNDA.n1214 585
R181 GNDA.n1353 GNDA.n1352 585
R182 GNDA.n1353 GNDA.n1201 585
R183 GNDA.n1354 GNDA.n1213 585
R184 GNDA.n1354 GNDA.n1202 585
R185 GNDA.n1357 GNDA.n1356 585
R186 GNDA.n1356 GNDA.n1355 585
R187 GNDA.n1358 GNDA.n1212 585
R188 GNDA.n1212 GNDA.n1211 585
R189 GNDA.n1360 GNDA.n1359 585
R190 GNDA.n1361 GNDA.n1360 585
R191 GNDA.n1210 GNDA.n1209 585
R192 GNDA.n1362 GNDA.n1210 585
R193 GNDA.n1365 GNDA.n1364 585
R194 GNDA.n1364 GNDA.n1363 585
R195 GNDA.n529 GNDA.n528 585
R196 GNDA.n528 GNDA.n49 585
R197 GNDA.n529 GNDA.n527 585
R198 GNDA.n527 GNDA.n526 585
R199 GNDA.n467 GNDA.n466 585
R200 GNDA.n525 GNDA.n467 585
R201 GNDA.n523 GNDA.n522 585
R202 GNDA.n524 GNDA.n523 585
R203 GNDA.n521 GNDA.n469 585
R204 GNDA.n469 GNDA.n468 585
R205 GNDA.n520 GNDA.n519 585
R206 GNDA.n519 GNDA.n518 585
R207 GNDA.n517 GNDA.n470 585
R208 GNDA.n517 GNDA.n56 585
R209 GNDA.n516 GNDA.n515 585
R210 GNDA.n516 GNDA.n57 585
R211 GNDA.n514 GNDA.n471 585
R212 GNDA.n474 GNDA.n471 585
R213 GNDA.n513 GNDA.n512 585
R214 GNDA.n512 GNDA.n511 585
R215 GNDA.n473 GNDA.n472 585
R216 GNDA.n510 GNDA.n473 585
R217 GNDA.n508 GNDA.n507 585
R218 GNDA.n509 GNDA.n508 585
R219 GNDA.n506 GNDA.n476 585
R220 GNDA.n476 GNDA.n475 585
R221 GNDA.n1502 GNDA.n1500 585
R222 GNDA.n1554 GNDA.n1502 585
R223 GNDA.n1552 GNDA.n1551 585
R224 GNDA.n1553 GNDA.n1552 585
R225 GNDA.n1550 GNDA.n1504 585
R226 GNDA.n1504 GNDA.n1503 585
R227 GNDA.n1549 GNDA.n1548 585
R228 GNDA.n1548 GNDA.n1547 585
R229 GNDA.n1546 GNDA.n1505 585
R230 GNDA.n1546 GNDA.n63 585
R231 GNDA.n1545 GNDA.n1544 585
R232 GNDA.n1545 GNDA.n64 585
R233 GNDA.n1543 GNDA.n1506 585
R234 GNDA.n1509 GNDA.n1506 585
R235 GNDA.n1542 GNDA.n1541 585
R236 GNDA.n1541 GNDA.n1540 585
R237 GNDA.n1508 GNDA.n1507 585
R238 GNDA.n1539 GNDA.n1508 585
R239 GNDA.n1537 GNDA.n1536 585
R240 GNDA.n1538 GNDA.n1537 585
R241 GNDA.n1535 GNDA.n1510 585
R242 GNDA.n1510 GNDA.n50 585
R243 GNDA.n170 GNDA.n18 585
R244 GNDA.n1848 GNDA.n18 585
R245 GNDA.n1851 GNDA.n1850 585
R246 GNDA.n1850 GNDA.n1849 585
R247 GNDA.n173 GNDA.n172 585
R248 GNDA.n1847 GNDA.n173 585
R249 GNDA.n1845 GNDA.n1844 585
R250 GNDA.n1846 GNDA.n1845 585
R251 GNDA.n1839 GNDA.n174 585
R252 GNDA.n1831 GNDA.n174 585
R253 GNDA.n1834 GNDA.n1833 585
R254 GNDA.n1833 GNDA.n1832 585
R255 GNDA.n176 GNDA.n175 585
R256 GNDA.n191 GNDA.n176 585
R257 GNDA.n189 GNDA.n188 585
R258 GNDA.n190 GNDA.n189 585
R259 GNDA.n183 GNDA.n181 585
R260 GNDA.n181 GNDA.n180 585
R261 GNDA.n177 GNDA.n149 585
R262 GNDA.n179 GNDA.n177 585
R263 GNDA.n1907 GNDA.n147 585
R264 GNDA.n178 GNDA.n147 585
R265 GNDA.n1910 GNDA.n1909 585
R266 GNDA.n1911 GNDA.n1910 585
R267 GNDA.n2033 GNDA.n2032 585
R268 GNDA.n1606 GNDA.n1604 585
R269 GNDA.n1610 GNDA.n1603 585
R270 GNDA.n1618 GNDA.n1603 585
R271 GNDA.n1609 GNDA.n1608 585
R272 GNDA.n196 GNDA.n194 585
R273 GNDA.n1826 GNDA.n193 585
R274 GNDA.n1830 GNDA.n193 585
R275 GNDA.n1824 GNDA.n1823 585
R276 GNDA.n621 GNDA.n620 585
R277 GNDA.n618 GNDA.n617 585
R278 GNDA.n616 GNDA.n615 585
R279 GNDA.n590 GNDA.n440 585
R280 GNDA.n596 GNDA.n595 585
R281 GNDA.n598 GNDA.n589 585
R282 GNDA.n600 GNDA.n599 585
R283 GNDA.n586 GNDA.n585 585
R284 GNDA.n606 GNDA.n605 585
R285 GNDA.n609 GNDA.n608 585
R286 GNDA.n584 GNDA.n463 585
R287 GNDA.n582 GNDA.n581 585
R288 GNDA.n745 GNDA.n744 585
R289 GNDA.n742 GNDA.n741 585
R290 GNDA.n627 GNDA.n626 585
R291 GNDA.n735 GNDA.n734 585
R292 GNDA.n732 GNDA.n731 585
R293 GNDA.n721 GNDA.n720 585
R294 GNDA.n723 GNDA.n722 585
R295 GNDA.n718 GNDA.n634 585
R296 GNDA.n717 GNDA.n716 585
R297 GNDA.n707 GNDA.n636 585
R298 GNDA.n709 GNDA.n708 585
R299 GNDA.n705 GNDA.n704 585
R300 GNDA.n934 GNDA.n815 585
R301 GNDA.n932 GNDA.n931 585
R302 GNDA.n851 GNDA.n816 585
R303 GNDA.n849 GNDA.n848 585
R304 GNDA.n861 GNDA.n860 585
R305 GNDA.n863 GNDA.n846 585
R306 GNDA.n865 GNDA.n864 585
R307 GNDA.n842 GNDA.n841 585
R308 GNDA.n872 GNDA.n871 585
R309 GNDA.n875 GNDA.n874 585
R310 GNDA.n840 GNDA.n836 585
R311 GNDA.n838 GNDA.n746 585
R312 GNDA.n1512 GNDA.n1511 585
R313 GNDA.n1514 GNDA.n1513 585
R314 GNDA.n1516 GNDA.n1515 585
R315 GNDA.n1518 GNDA.n1517 585
R316 GNDA.n1520 GNDA.n1519 585
R317 GNDA.n1522 GNDA.n1521 585
R318 GNDA.n1524 GNDA.n1523 585
R319 GNDA.n1526 GNDA.n1525 585
R320 GNDA.n1528 GNDA.n1527 585
R321 GNDA.n1530 GNDA.n1529 585
R322 GNDA.n1532 GNDA.n1531 585
R323 GNDA.n1534 GNDA.n1533 585
R324 GNDA.n1960 GNDA.n1959 585
R325 GNDA.n1962 GNDA.n1961 585
R326 GNDA.n1964 GNDA.n1963 585
R327 GNDA.n1966 GNDA.n1965 585
R328 GNDA.n1968 GNDA.n1967 585
R329 GNDA.n1970 GNDA.n1969 585
R330 GNDA.n1972 GNDA.n1971 585
R331 GNDA.n1974 GNDA.n1973 585
R332 GNDA.n1976 GNDA.n1975 585
R333 GNDA.n1978 GNDA.n1977 585
R334 GNDA.n1980 GNDA.n1979 585
R335 GNDA.n1982 GNDA.n1981 585
R336 GNDA.n2010 GNDA.n28 585
R337 GNDA.n99 GNDA.n30 585
R338 GNDA.n101 GNDA.n100 585
R339 GNDA.n103 GNDA.n102 585
R340 GNDA.n105 GNDA.n104 585
R341 GNDA.n107 GNDA.n106 585
R342 GNDA.n109 GNDA.n108 585
R343 GNDA.n111 GNDA.n110 585
R344 GNDA.n113 GNDA.n112 585
R345 GNDA.n115 GNDA.n114 585
R346 GNDA.n117 GNDA.n116 585
R347 GNDA.n119 GNDA.n118 585
R348 GNDA.n1276 GNDA.n1049 585
R349 GNDA.n1279 GNDA.n1278 585
R350 GNDA.n1275 GNDA.n1245 585
R351 GNDA.n1273 GNDA.n1272 585
R352 GNDA.n1267 GNDA.n1246 585
R353 GNDA.n1262 GNDA.n1261 585
R354 GNDA.n1259 GNDA.n1247 585
R355 GNDA.n1257 GNDA.n1256 585
R356 GNDA.n1251 GNDA.n1249 585
R357 GNDA.n1222 GNDA.n1220 585
R358 GNDA.n1336 GNDA.n1335 585
R359 GNDA.n1338 GNDA.n1219 585
R360 GNDA.n485 GNDA.n421 585
R361 GNDA.n487 GNDA.n483 585
R362 GNDA.n489 GNDA.n488 585
R363 GNDA.n490 GNDA.n482 585
R364 GNDA.n492 GNDA.n491 585
R365 GNDA.n494 GNDA.n480 585
R366 GNDA.n496 GNDA.n495 585
R367 GNDA.n497 GNDA.n479 585
R368 GNDA.n499 GNDA.n498 585
R369 GNDA.n501 GNDA.n478 585
R370 GNDA.n502 GNDA.n477 585
R371 GNDA.n505 GNDA.n504 585
R372 GNDA.n798 GNDA.n797 585
R373 GNDA.n795 GNDA.n771 585
R374 GNDA.n794 GNDA.n793 585
R375 GNDA.n792 GNDA.n791 585
R376 GNDA.n790 GNDA.n773 585
R377 GNDA.n788 GNDA.n787 585
R378 GNDA.n786 GNDA.n774 585
R379 GNDA.n785 GNDA.n784 585
R380 GNDA.n782 GNDA.n775 585
R381 GNDA.n780 GNDA.n779 585
R382 GNDA.n778 GNDA.n777 585
R383 GNDA.n424 GNDA.n420 585
R384 GNDA.n961 GNDA.n960 585
R385 GNDA.n962 GNDA.n807 585
R386 GNDA.n964 GNDA.n963 585
R387 GNDA.n966 GNDA.n805 585
R388 GNDA.n968 GNDA.n967 585
R389 GNDA.n969 GNDA.n804 585
R390 GNDA.n971 GNDA.n970 585
R391 GNDA.n973 GNDA.n802 585
R392 GNDA.n975 GNDA.n974 585
R393 GNDA.n976 GNDA.n801 585
R394 GNDA.n978 GNDA.n977 585
R395 GNDA.n980 GNDA.n800 585
R396 GNDA.n1389 GNDA.n1388 585
R397 GNDA.n1388 GNDA.n1387 585
R398 GNDA.n1186 GNDA.n1185 585
R399 GNDA.n1386 GNDA.n1186 585
R400 GNDA.n1384 GNDA.n1383 585
R401 GNDA.n1385 GNDA.n1384 585
R402 GNDA.n1382 GNDA.n1188 585
R403 GNDA.n1188 GNDA.n1187 585
R404 GNDA.n1381 GNDA.n1380 585
R405 GNDA.n1380 GNDA.n1379 585
R406 GNDA.n1190 GNDA.n1189 585
R407 GNDA.n1378 GNDA.n1190 585
R408 GNDA.n1376 GNDA.n1375 585
R409 GNDA.n1377 GNDA.n1376 585
R410 GNDA.n1374 GNDA.n1204 585
R411 GNDA.n1204 GNDA.n1203 585
R412 GNDA.n1373 GNDA.n1372 585
R413 GNDA.n1372 GNDA.n1371 585
R414 GNDA.n1206 GNDA.n1205 585
R415 GNDA.n1370 GNDA.n1206 585
R416 GNDA.n1368 GNDA.n1367 585
R417 GNDA.n1369 GNDA.n1368 585
R418 GNDA.n1366 GNDA.n1208 585
R419 GNDA.n1208 GNDA.n1207 585
R420 GNDA.n396 GNDA.n395 585
R421 GNDA.n395 GNDA.n52 585
R422 GNDA.n397 GNDA.n242 585
R423 GNDA.n242 GNDA.n241 585
R424 GNDA.n399 GNDA.n398 585
R425 GNDA.n400 GNDA.n399 585
R426 GNDA.n240 GNDA.n239 585
R427 GNDA.n401 GNDA.n240 585
R428 GNDA.n404 GNDA.n403 585
R429 GNDA.n403 GNDA.n402 585
R430 GNDA.n405 GNDA.n238 585
R431 GNDA.n238 GNDA.n55 585
R432 GNDA.n407 GNDA.n406 585
R433 GNDA.n407 GNDA.n54 585
R434 GNDA.n408 GNDA.n237 585
R435 GNDA.n409 GNDA.n408 585
R436 GNDA.n412 GNDA.n411 585
R437 GNDA.n411 GNDA.n410 585
R438 GNDA.n413 GNDA.n236 585
R439 GNDA.n236 GNDA.n235 585
R440 GNDA.n415 GNDA.n414 585
R441 GNDA.n416 GNDA.n415 585
R442 GNDA.n220 GNDA.n217 585
R443 GNDA.n417 GNDA.n220 585
R444 GNDA.n394 GNDA.n243 585
R445 GNDA.n394 GNDA.n20 585
R446 GNDA.n393 GNDA.n244 585
R447 GNDA.n391 GNDA.n390 585
R448 GNDA.n389 GNDA.n245 585
R449 GNDA.n388 GNDA.n387 585
R450 GNDA.n385 GNDA.n246 585
R451 GNDA.n383 GNDA.n382 585
R452 GNDA.n381 GNDA.n247 585
R453 GNDA.n380 GNDA.n379 585
R454 GNDA.n377 GNDA.n248 585
R455 GNDA.n375 GNDA.n374 585
R456 GNDA.n370 GNDA.n250 585
R457 GNDA.n368 GNDA.n367 585
R458 GNDA.n287 GNDA.n251 585
R459 GNDA.n285 GNDA.n284 585
R460 GNDA.n297 GNDA.n296 585
R461 GNDA.n299 GNDA.n282 585
R462 GNDA.n301 GNDA.n300 585
R463 GNDA.n278 GNDA.n277 585
R464 GNDA.n308 GNDA.n307 585
R465 GNDA.n311 GNDA.n310 585
R466 GNDA.n276 GNDA.n271 585
R467 GNDA.n274 GNDA.n273 585
R468 GNDA.n373 GNDA.n372 585
R469 GNDA.n373 GNDA.n249 585
R470 GNDA.n1074 GNDA.n232 585
R471 GNDA.n1109 GNDA.n1108 585
R472 GNDA.n1106 GNDA.n1076 585
R473 GNDA.n1104 GNDA.n1103 585
R474 GNDA.n1098 GNDA.n1077 585
R475 GNDA.n1093 GNDA.n1092 585
R476 GNDA.n1090 GNDA.n1078 585
R477 GNDA.n1088 GNDA.n1087 585
R478 GNDA.n1082 GNDA.n1080 585
R479 GNDA.n1052 GNDA.n1051 585
R480 GNDA.n1166 GNDA.n1165 585
R481 GNDA.n1169 GNDA.n1168 585
R482 GNDA.n1435 GNDA.n233 585
R483 GNDA.n1435 GNDA.n1434 585
R484 GNDA.n1472 GNDA.n219 585
R485 GNDA.n1461 GNDA.n218 585
R486 GNDA.n1462 GNDA.n221 585
R487 GNDA.n1465 GNDA.n1464 585
R488 GNDA.n1459 GNDA.n223 585
R489 GNDA.n1457 GNDA.n1456 585
R490 GNDA.n225 GNDA.n224 585
R491 GNDA.n1450 GNDA.n1449 585
R492 GNDA.n1447 GNDA.n227 585
R493 GNDA.n1445 GNDA.n1444 585
R494 GNDA.n229 GNDA.n228 585
R495 GNDA.n1438 GNDA.n1437 585
R496 GNDA.n418 GNDA.n233 585
R497 GNDA.n1434 GNDA.n418 585
R498 GNDA.n1439 GNDA.n1438 585
R499 GNDA.n1441 GNDA.n229 585
R500 GNDA.n1444 GNDA.n1443 585
R501 GNDA.n227 GNDA.n226 585
R502 GNDA.n1451 GNDA.n1450 585
R503 GNDA.n1453 GNDA.n225 585
R504 GNDA.n1456 GNDA.n1455 585
R505 GNDA.n223 GNDA.n222 585
R506 GNDA.n1466 GNDA.n1465 585
R507 GNDA.n1468 GNDA.n221 585
R508 GNDA.n1469 GNDA.n218 585
R509 GNDA.n1472 GNDA.n1471 585
R510 GNDA.n1006 GNDA.n623 585
R511 GNDA.n1009 GNDA.n623 585
R512 GNDA.n983 GNDA.n770 585
R513 GNDA.n984 GNDA.n768 585
R514 GNDA.n985 GNDA.n767 585
R515 GNDA.n765 GNDA.n763 585
R516 GNDA.n991 GNDA.n762 585
R517 GNDA.n992 GNDA.n760 585
R518 GNDA.n993 GNDA.n759 585
R519 GNDA.n757 GNDA.n755 585
R520 GNDA.n998 GNDA.n754 585
R521 GNDA.n999 GNDA.n752 585
R522 GNDA.n751 GNDA.n748 585
R523 GNDA.n1004 GNDA.n747 585
R524 GNDA.n1007 GNDA.n1006 585
R525 GNDA.n1009 GNDA.n1007 585
R526 GNDA.n1004 GNDA.n1003 585
R527 GNDA.n1001 GNDA.n748 585
R528 GNDA.n1000 GNDA.n999 585
R529 GNDA.n998 GNDA.n997 585
R530 GNDA.n996 GNDA.n755 585
R531 GNDA.n994 GNDA.n993 585
R532 GNDA.n992 GNDA.n756 585
R533 GNDA.n991 GNDA.n990 585
R534 GNDA.n988 GNDA.n763 585
R535 GNDA.n986 GNDA.n985 585
R536 GNDA.n984 GNDA.n764 585
R537 GNDA.n983 GNDA.n982 585
R538 GNDA.n1921 GNDA.n132 585
R539 GNDA.n1921 GNDA.n1920 585
R540 GNDA.n1958 GNDA.n1957 585
R541 GNDA.n1946 GNDA.n98 585
R542 GNDA.n1947 GNDA.n120 585
R543 GNDA.n1950 GNDA.n1949 585
R544 GNDA.n1945 GNDA.n122 585
R545 GNDA.n1943 GNDA.n1942 585
R546 GNDA.n124 GNDA.n123 585
R547 GNDA.n1936 GNDA.n1935 585
R548 GNDA.n1933 GNDA.n126 585
R549 GNDA.n1931 GNDA.n1930 585
R550 GNDA.n128 GNDA.n127 585
R551 GNDA.n1924 GNDA.n1923 585
R552 GNDA.n145 GNDA.n132 585
R553 GNDA.n146 GNDA.n145 585
R554 GNDA.n1925 GNDA.n1924 585
R555 GNDA.n1927 GNDA.n128 585
R556 GNDA.n1930 GNDA.n1929 585
R557 GNDA.n126 GNDA.n125 585
R558 GNDA.n1937 GNDA.n1936 585
R559 GNDA.n1939 GNDA.n124 585
R560 GNDA.n1942 GNDA.n1941 585
R561 GNDA.n122 GNDA.n121 585
R562 GNDA.n1951 GNDA.n1950 585
R563 GNDA.n1953 GNDA.n120 585
R564 GNDA.n1954 GNDA.n98 585
R565 GNDA.n1957 GNDA.n1956 585
R566 GNDA.n1747 GNDA.n131 585
R567 GNDA.n133 GNDA.n131 585
R568 GNDA.n9 GNDA.n6 585
R569 GNDA.n1817 GNDA.n6 585
R570 GNDA.n2053 GNDA.n2052 585
R571 GNDA.n2054 GNDA.n2053 585
R572 GNDA.n7 GNDA.n5 585
R573 GNDA.n2055 GNDA.n5 585
R574 GNDA.n2058 GNDA.n2057 585
R575 GNDA.n2057 GNDA.n2056 585
R576 GNDA.n11 GNDA.n4 585
R577 GNDA.n2036 GNDA.n4 585
R578 GNDA.n2040 GNDA.n2039 585
R579 GNDA.n2039 GNDA.n2038 585
R580 GNDA.n15 GNDA.n14 585
R581 GNDA.n1805 GNDA.n15 585
R582 GNDA.n1808 GNDA.n1807 585
R583 GNDA.n1807 GNDA.n1806 585
R584 GNDA.n1733 GNDA.n1730 585
R585 GNDA.n1804 GNDA.n1730 585
R586 GNDA.n1814 GNDA.n1813 585
R587 GNDA.n1815 GNDA.n1814 585
R588 GNDA.n1731 GNDA.n1729 585
R589 GNDA.n1729 GNDA.n1728 585
R590 GNDA.n1580 GNDA.n200 585
R591 GNDA.n1636 GNDA.n200 585
R592 GNDA.n1639 GNDA.n1638 585
R593 GNDA.n1638 GNDA.n1637 585
R594 GNDA.n1583 GNDA.n1582 585
R595 GNDA.n1635 GNDA.n1583 585
R596 GNDA.n1633 GNDA.n1632 585
R597 GNDA.n1634 GNDA.n1633 585
R598 GNDA.n1627 GNDA.n1584 585
R599 GNDA.n1619 GNDA.n1584 585
R600 GNDA.n1622 GNDA.n1621 585
R601 GNDA.n1621 GNDA.n1620 585
R602 GNDA.n1586 GNDA.n1585 585
R603 GNDA.n1601 GNDA.n1586 585
R604 GNDA.n1599 GNDA.n1598 585
R605 GNDA.n1600 GNDA.n1599 585
R606 GNDA.n1593 GNDA.n1591 585
R607 GNDA.n1591 GNDA.n1590 585
R608 GNDA.n1587 GNDA.n1559 585
R609 GNDA.n1589 GNDA.n1587 585
R610 GNDA.n1695 GNDA.n1499 585
R611 GNDA.n1588 GNDA.n1499 585
R612 GNDA.n1698 GNDA.n1697 585
R613 GNDA.n1699 GNDA.n1698 585
R614 GNDA.n1557 GNDA.n1501 585
R615 GNDA.n1501 GNDA.n1497 585
R616 GNDA.n1557 GNDA.n1556 585
R617 GNDA.n1556 GNDA.n1555 585
R618 GNDA.n1725 GNDA.n1724 585
R619 GNDA.n1724 GNDA.n1723 585
R620 GNDA.n1984 GNDA.n94 585
R621 GNDA.n1985 GNDA.n92 585
R622 GNDA.n1988 GNDA.n91 585
R623 GNDA.n1989 GNDA.n89 585
R624 GNDA.n1992 GNDA.n88 585
R625 GNDA.n1993 GNDA.n86 585
R626 GNDA.n1996 GNDA.n85 585
R627 GNDA.n1997 GNDA.n83 585
R628 GNDA.n2000 GNDA.n82 585
R629 GNDA.n2002 GNDA.n80 585
R630 GNDA.n2003 GNDA.n79 585
R631 GNDA.n2004 GNDA.n77 585
R632 GNDA.n1726 GNDA.n1725 585
R633 GNDA.n1727 GNDA.n1726 585
R634 GNDA.n2005 GNDA.n2004 585
R635 GNDA.n2003 GNDA.n74 585
R636 GNDA.n2002 GNDA.n2001 585
R637 GNDA.n2000 GNDA.n1999 585
R638 GNDA.n1998 GNDA.n1997 585
R639 GNDA.n1996 GNDA.n1995 585
R640 GNDA.n1994 GNDA.n1993 585
R641 GNDA.n1992 GNDA.n1991 585
R642 GNDA.n1990 GNDA.n1989 585
R643 GNDA.n1988 GNDA.n1987 585
R644 GNDA.n1986 GNDA.n1985 585
R645 GNDA.n1984 GNDA.n1983 585
R646 GNDA.n1010 GNDA.n622 585
R647 GNDA.n1010 GNDA.n1009 585
R648 GNDA.n1047 GNDA.n423 585
R649 GNDA.n1036 GNDA.n422 585
R650 GNDA.n1037 GNDA.n425 585
R651 GNDA.n1040 GNDA.n1039 585
R652 GNDA.n1034 GNDA.n427 585
R653 GNDA.n1032 GNDA.n1031 585
R654 GNDA.n429 GNDA.n428 585
R655 GNDA.n1025 GNDA.n1024 585
R656 GNDA.n1022 GNDA.n431 585
R657 GNDA.n1020 GNDA.n1019 585
R658 GNDA.n433 GNDA.n432 585
R659 GNDA.n1013 GNDA.n1012 585
R660 GNDA.n1008 GNDA.n622 585
R661 GNDA.n1009 GNDA.n1008 585
R662 GNDA.n1014 GNDA.n1013 585
R663 GNDA.n1016 GNDA.n433 585
R664 GNDA.n1019 GNDA.n1018 585
R665 GNDA.n431 GNDA.n430 585
R666 GNDA.n1026 GNDA.n1025 585
R667 GNDA.n1028 GNDA.n429 585
R668 GNDA.n1031 GNDA.n1030 585
R669 GNDA.n427 GNDA.n426 585
R670 GNDA.n1041 GNDA.n1040 585
R671 GNDA.n1043 GNDA.n425 585
R672 GNDA.n1044 GNDA.n422 585
R673 GNDA.n1047 GNDA.n1046 585
R674 GNDA.n1432 GNDA.n234 585
R675 GNDA.n1434 GNDA.n234 585
R676 GNDA.n1409 GNDA.n1184 585
R677 GNDA.n1410 GNDA.n1183 585
R678 GNDA.n1411 GNDA.n1182 585
R679 GNDA.n1197 GNDA.n1180 585
R680 GNDA.n1417 GNDA.n1179 585
R681 GNDA.n1418 GNDA.n1178 585
R682 GNDA.n1419 GNDA.n1177 585
R683 GNDA.n1194 GNDA.n1175 585
R684 GNDA.n1424 GNDA.n1174 585
R685 GNDA.n1425 GNDA.n1173 585
R686 GNDA.n1191 GNDA.n1171 585
R687 GNDA.n1430 GNDA.n1170 585
R688 GNDA.n1433 GNDA.n1432 585
R689 GNDA.n1434 GNDA.n1433 585
R690 GNDA.n1430 GNDA.n1429 585
R691 GNDA.n1427 GNDA.n1171 585
R692 GNDA.n1426 GNDA.n1425 585
R693 GNDA.n1424 GNDA.n1423 585
R694 GNDA.n1422 GNDA.n1175 585
R695 GNDA.n1420 GNDA.n1419 585
R696 GNDA.n1418 GNDA.n1176 585
R697 GNDA.n1417 GNDA.n1416 585
R698 GNDA.n1414 GNDA.n1180 585
R699 GNDA.n1412 GNDA.n1411 585
R700 GNDA.n1410 GNDA.n1181 585
R701 GNDA.n1409 GNDA.n1408 585
R702 GNDA.n1474 GNDA.n216 585
R703 GNDA.n216 GNDA.n215 585
R704 GNDA.n1476 GNDA.n1475 585
R705 GNDA.n1477 GNDA.n1476 585
R706 GNDA.n214 GNDA.n213 585
R707 GNDA.n1478 GNDA.n214 585
R708 GNDA.n1481 GNDA.n1480 585
R709 GNDA.n1480 GNDA.n1479 585
R710 GNDA.n1482 GNDA.n210 585
R711 GNDA.n210 GNDA.n208 585
R712 GNDA.n1484 GNDA.n1483 585
R713 GNDA.n1485 GNDA.n1484 585
R714 GNDA.n1396 GNDA.n209 585
R715 GNDA.n209 GNDA.n206 585
R716 GNDA.n1399 GNDA.n1398 585
R717 GNDA.n1398 GNDA.n1397 585
R718 GNDA.n1400 GNDA.n1394 585
R719 GNDA.n1394 GNDA.n1393 585
R720 GNDA.n1402 GNDA.n1401 585
R721 GNDA.n1403 GNDA.n1402 585
R722 GNDA.n1395 GNDA.n1391 585
R723 GNDA.n1404 GNDA.n1391 585
R724 GNDA.n1406 GNDA.n1392 585
R725 GNDA.n1406 GNDA.n1405 585
R726 GNDA.n203 GNDA.n202 585
R727 GNDA.n1487 GNDA.n1486 585
R728 GNDA.n1486 GNDA.t77 585
R729 GNDA.n1702 GNDA.t87 409.067
R730 GNDA.n1720 GNDA.t82 409.067
R731 GNDA.n1717 GNDA.t93 409.067
R732 GNDA.n1917 GNDA.t99 409.067
R733 GNDA.n1914 GNDA.t102 409.067
R734 GNDA.n138 GNDA.t96 409.067
R735 GNDA.n134 GNDA.n65 370.214
R736 GNDA.n68 GNDA.n67 370.214
R737 GNDA.n134 GNDA.n66 365.957
R738 GNDA.n2007 GNDA.n68 365.957
R739 GNDA.t77 GNDA.n204 172.876
R740 GNDA.t77 GNDA.n66 327.661
R741 GNDA.t77 GNDA.n2007 327.661
R742 GNDA.t77 GNDA.n59 172.876
R743 GNDA.t77 GNDA.n61 172.876
R744 GNDA.t77 GNDA.n53 172.876
R745 GNDA.t77 GNDA.n1200 172.615
R746 GNDA.t77 GNDA.n65 323.404
R747 GNDA.t77 GNDA.n67 323.404
R748 GNDA.t77 GNDA.n58 172.615
R749 GNDA.t77 GNDA.n60 172.615
R750 GNDA.t77 GNDA.n205 172.615
R751 GNDA.t77 GNDA.n50 274.089
R752 GNDA.n371 GNDA.n20 263.904
R753 GNDA.n938 GNDA.n937 263.904
R754 GNDA.n2031 GNDA.n19 263.904
R755 GNDA.n1408 GNDA.n1406 257.466
R756 GNDA.n1983 GNDA.n1982 257.466
R757 GNDA.n1046 GNDA.n424 257.466
R758 GNDA.n1956 GNDA.n119 257.466
R759 GNDA.n982 GNDA.n980 257.466
R760 GNDA.n1533 GNDA.n1510 257.466
R761 GNDA.n504 GNDA.n476 257.466
R762 GNDA.n1364 GNDA.n1208 257.466
R763 GNDA.n1471 GNDA.n220 257.466
R764 GNDA.n958 GNDA.n20 254.34
R765 GNDA.n952 GNDA.n20 254.34
R766 GNDA.n950 GNDA.n20 254.34
R767 GNDA.n944 GNDA.n20 254.34
R768 GNDA.n942 GNDA.n20 254.34
R769 GNDA.n936 GNDA.n20 254.34
R770 GNDA.n29 GNDA.n20 254.34
R771 GNDA.n2016 GNDA.n20 254.34
R772 GNDA.n26 GNDA.n20 254.34
R773 GNDA.n2023 GNDA.n20 254.34
R774 GNDA.n23 GNDA.n20 254.34
R775 GNDA.n2030 GNDA.n20 254.34
R776 GNDA.n436 GNDA.n48 254.34
R777 GNDA.n439 GNDA.n48 254.34
R778 GNDA.n597 GNDA.n48 254.34
R779 GNDA.n588 GNDA.n48 254.34
R780 GNDA.n607 GNDA.n48 254.34
R781 GNDA.n583 GNDA.n48 254.34
R782 GNDA.n743 GNDA.n48 254.34
R783 GNDA.n733 GNDA.n48 254.34
R784 GNDA.n631 GNDA.n48 254.34
R785 GNDA.n719 GNDA.n48 254.34
R786 GNDA.n635 GNDA.n48 254.34
R787 GNDA.n706 GNDA.n48 254.34
R788 GNDA.n933 GNDA.n48 254.34
R789 GNDA.n847 GNDA.n48 254.34
R790 GNDA.n862 GNDA.n48 254.34
R791 GNDA.n845 GNDA.n48 254.34
R792 GNDA.n873 GNDA.n48 254.34
R793 GNDA.n839 GNDA.n48 254.34
R794 GNDA.n2008 GNDA.n47 254.34
R795 GNDA.n2008 GNDA.n46 254.34
R796 GNDA.n2008 GNDA.n45 254.34
R797 GNDA.n2008 GNDA.n44 254.34
R798 GNDA.n2008 GNDA.n43 254.34
R799 GNDA.n2008 GNDA.n42 254.34
R800 GNDA.n2008 GNDA.n41 254.34
R801 GNDA.n2008 GNDA.n40 254.34
R802 GNDA.n2008 GNDA.n39 254.34
R803 GNDA.n2008 GNDA.n38 254.34
R804 GNDA.n2008 GNDA.n37 254.34
R805 GNDA.n2008 GNDA.n36 254.34
R806 GNDA.n2009 GNDA.n2008 254.34
R807 GNDA.n2008 GNDA.n35 254.34
R808 GNDA.n2008 GNDA.n34 254.34
R809 GNDA.n2008 GNDA.n33 254.34
R810 GNDA.n2008 GNDA.n32 254.34
R811 GNDA.n2008 GNDA.n31 254.34
R812 GNDA.n1277 GNDA.n51 254.34
R813 GNDA.n1274 GNDA.n51 254.34
R814 GNDA.n1260 GNDA.n51 254.34
R815 GNDA.n1258 GNDA.n51 254.34
R816 GNDA.n1248 GNDA.n51 254.34
R817 GNDA.n1337 GNDA.n51 254.34
R818 GNDA.n486 GNDA.n62 254.34
R819 GNDA.n484 GNDA.n62 254.34
R820 GNDA.n493 GNDA.n62 254.34
R821 GNDA.n481 GNDA.n62 254.34
R822 GNDA.n500 GNDA.n62 254.34
R823 GNDA.n503 GNDA.n62 254.34
R824 GNDA.n796 GNDA.n62 254.34
R825 GNDA.n772 GNDA.n62 254.34
R826 GNDA.n789 GNDA.n62 254.34
R827 GNDA.n783 GNDA.n62 254.34
R828 GNDA.n781 GNDA.n62 254.34
R829 GNDA.n776 GNDA.n62 254.34
R830 GNDA.n809 GNDA.n62 254.34
R831 GNDA.n965 GNDA.n62 254.34
R832 GNDA.n806 GNDA.n62 254.34
R833 GNDA.n972 GNDA.n62 254.34
R834 GNDA.n803 GNDA.n62 254.34
R835 GNDA.n979 GNDA.n62 254.34
R836 GNDA.n392 GNDA.n20 254.34
R837 GNDA.n386 GNDA.n20 254.34
R838 GNDA.n384 GNDA.n20 254.34
R839 GNDA.n378 GNDA.n20 254.34
R840 GNDA.n376 GNDA.n20 254.34
R841 GNDA.n369 GNDA.n51 254.34
R842 GNDA.n283 GNDA.n51 254.34
R843 GNDA.n298 GNDA.n51 254.34
R844 GNDA.n281 GNDA.n51 254.34
R845 GNDA.n309 GNDA.n51 254.34
R846 GNDA.n275 GNDA.n51 254.34
R847 GNDA.n1107 GNDA.n51 254.34
R848 GNDA.n1105 GNDA.n51 254.34
R849 GNDA.n1091 GNDA.n51 254.34
R850 GNDA.n1089 GNDA.n51 254.34
R851 GNDA.n1079 GNDA.n51 254.34
R852 GNDA.n1167 GNDA.n51 254.34
R853 GNDA.n1460 GNDA.n205 254.34
R854 GNDA.n1463 GNDA.n205 254.34
R855 GNDA.n1458 GNDA.n205 254.34
R856 GNDA.n1448 GNDA.n205 254.34
R857 GNDA.n1446 GNDA.n205 254.34
R858 GNDA.n1436 GNDA.n205 254.34
R859 GNDA.n1440 GNDA.n53 254.34
R860 GNDA.n1442 GNDA.n53 254.34
R861 GNDA.n1452 GNDA.n53 254.34
R862 GNDA.n1454 GNDA.n53 254.34
R863 GNDA.n1467 GNDA.n53 254.34
R864 GNDA.n1470 GNDA.n53 254.34
R865 GNDA.n769 GNDA.n58 254.34
R866 GNDA.n766 GNDA.n58 254.34
R867 GNDA.n761 GNDA.n58 254.34
R868 GNDA.n758 GNDA.n58 254.34
R869 GNDA.n753 GNDA.n58 254.34
R870 GNDA.n750 GNDA.n58 254.34
R871 GNDA.n1002 GNDA.n59 254.34
R872 GNDA.n749 GNDA.n59 254.34
R873 GNDA.n995 GNDA.n59 254.34
R874 GNDA.n989 GNDA.n59 254.34
R875 GNDA.n987 GNDA.n59 254.34
R876 GNDA.n981 GNDA.n59 254.34
R877 GNDA.n97 GNDA.n65 254.34
R878 GNDA.n1948 GNDA.n65 254.34
R879 GNDA.n1944 GNDA.n65 254.34
R880 GNDA.n1934 GNDA.n65 254.34
R881 GNDA.n1932 GNDA.n65 254.34
R882 GNDA.n1922 GNDA.n65 254.34
R883 GNDA.n1926 GNDA.n66 254.34
R884 GNDA.n1928 GNDA.n66 254.34
R885 GNDA.n1938 GNDA.n66 254.34
R886 GNDA.n1940 GNDA.n66 254.34
R887 GNDA.n1952 GNDA.n66 254.34
R888 GNDA.n1955 GNDA.n66 254.34
R889 GNDA.n93 GNDA.n67 254.34
R890 GNDA.n90 GNDA.n67 254.34
R891 GNDA.n87 GNDA.n67 254.34
R892 GNDA.n84 GNDA.n67 254.34
R893 GNDA.n81 GNDA.n67 254.34
R894 GNDA.n78 GNDA.n67 254.34
R895 GNDA.n2007 GNDA.n2006 254.34
R896 GNDA.n2007 GNDA.n73 254.34
R897 GNDA.n2007 GNDA.n72 254.34
R898 GNDA.n2007 GNDA.n71 254.34
R899 GNDA.n2007 GNDA.n70 254.34
R900 GNDA.n2007 GNDA.n69 254.34
R901 GNDA.n1035 GNDA.n60 254.34
R902 GNDA.n1038 GNDA.n60 254.34
R903 GNDA.n1033 GNDA.n60 254.34
R904 GNDA.n1023 GNDA.n60 254.34
R905 GNDA.n1021 GNDA.n60 254.34
R906 GNDA.n1011 GNDA.n60 254.34
R907 GNDA.n1015 GNDA.n61 254.34
R908 GNDA.n1017 GNDA.n61 254.34
R909 GNDA.n1027 GNDA.n61 254.34
R910 GNDA.n1029 GNDA.n61 254.34
R911 GNDA.n1042 GNDA.n61 254.34
R912 GNDA.n1045 GNDA.n61 254.34
R913 GNDA.n1200 GNDA.n1199 254.34
R914 GNDA.n1200 GNDA.n1198 254.34
R915 GNDA.n1200 GNDA.n1196 254.34
R916 GNDA.n1200 GNDA.n1195 254.34
R917 GNDA.n1200 GNDA.n1193 254.34
R918 GNDA.n1200 GNDA.n1192 254.34
R919 GNDA.n1428 GNDA.n204 254.34
R920 GNDA.n1172 GNDA.n204 254.34
R921 GNDA.n1421 GNDA.n204 254.34
R922 GNDA.n1415 GNDA.n204 254.34
R923 GNDA.n1413 GNDA.n204 254.34
R924 GNDA.n1407 GNDA.n204 254.34
R925 GNDA.n219 GNDA.n216 251.614
R926 GNDA.n1959 GNDA.n1958 251.614
R927 GNDA.n797 GNDA.n770 251.614
R928 GNDA.n2011 GNDA.n2010 251.614
R929 GNDA.n960 GNDA.n959 251.614
R930 GNDA.n1511 GNDA.n94 251.614
R931 GNDA.n485 GNDA.n423 251.614
R932 GNDA.n1388 GNDA.n1184 251.614
R933 GNDA.n395 GNDA.n394 251.614
R934 GNDA.t77 GNDA.n207 250.349
R935 GNDA.n475 GNDA.t7 248.139
R936 GNDA.n194 GNDA.n193 246.25
R937 GNDA.n1823 GNDA.n193 246.25
R938 GNDA.n1604 GNDA.n1603 246.25
R939 GNDA.n1608 GNDA.n1603 246.25
R940 GNDA.n1618 GNDA.n1617 241.643
R941 GNDA.n1618 GNDA.n1602 241.643
R942 GNDA.n1830 GNDA.n1829 241.643
R943 GNDA.n1830 GNDA.n192 241.643
R944 GNDA.t20 GNDA.t30 224.626
R945 GNDA.n1642 GNDA.n1641 221.667
R946 GNDA.n1112 GNDA.n1111 221.667
R947 GNDA.n739 GNDA.n628 221.667
R948 GNDA.n1854 GNDA.n1853 221.667
R949 GNDA.n928 GNDA.n819 221.667
R950 GNDA.n451 GNDA.n442 221.667
R951 GNDA.n1282 GNDA.n1281 221.667
R952 GNDA.n364 GNDA.n254 221.667
R953 GNDA.n2050 GNDA.n10 221.667
R954 GNDA.t11 GNDA.t5 219.279
R955 GNDA.n20 GNDA.t15 215
R956 GNDA.t17 GNDA.n1496 205.945
R957 GNDA.n1486 GNDA.n203 197
R958 GNDA.n1168 GNDA.n419 195.049
R959 GNDA.n1729 GNDA.n75 195.049
R960 GNDA.n705 GNDA.n434 195.049
R961 GNDA.n1910 GNDA.n129 195.049
R962 GNDA.n838 GNDA.n624 195.049
R963 GNDA.n1698 GNDA.n1498 195.049
R964 GNDA.n582 GNDA.n465 195.049
R965 GNDA.n1339 GNDA.n1338 195.049
R966 GNDA.n274 GNDA.n230 195.049
R967 GNDA.n1435 GNDA.n232 187.249
R968 GNDA.n1921 GNDA.n131 187.249
R969 GNDA.n744 GNDA.n623 187.249
R970 GNDA.n2032 GNDA.n18 187.249
R971 GNDA.n935 GNDA.n934 187.249
R972 GNDA.n1724 GNDA.n200 187.249
R973 GNDA.n1010 GNDA.n621 187.249
R974 GNDA.n1276 GNDA.n234 187.249
R975 GNDA.n372 GNDA.n370 187.249
R976 GNDA.n1659 GNDA.n1658 185
R977 GNDA.n1657 GNDA.n1656 185
R978 GNDA.n1655 GNDA.n1654 185
R979 GNDA.n1653 GNDA.n1652 185
R980 GNDA.n1651 GNDA.n1650 185
R981 GNDA.n1649 GNDA.n1648 185
R982 GNDA.n1647 GNDA.n1646 185
R983 GNDA.n1645 GNDA.n1644 185
R984 GNDA.n1643 GNDA.n1642 185
R985 GNDA.n1661 GNDA.n1660 185
R986 GNDA.n1662 GNDA.n1569 185
R987 GNDA.t92 GNDA.n1569 185
R988 GNDA.n1664 GNDA.n1663 185
R989 GNDA.n1666 GNDA.n1665 185
R990 GNDA.n1668 GNDA.n1667 185
R991 GNDA.n1670 GNDA.n1669 185
R992 GNDA.n1672 GNDA.n1671 185
R993 GNDA.n1674 GNDA.n1673 185
R994 GNDA.n1676 GNDA.n1675 185
R995 GNDA.n1560 GNDA.n1558 185
R996 GNDA.n1691 GNDA.n1690 185
R997 GNDA.n1689 GNDA.n1579 185
R998 GNDA.n1688 GNDA.n1687 185
R999 GNDA.n1686 GNDA.n1685 185
R1000 GNDA.n1684 GNDA.n1683 185
R1001 GNDA.n1682 GNDA.n1681 185
R1002 GNDA.n1680 GNDA.n1679 185
R1003 GNDA.n1678 GNDA.n1677 185
R1004 GNDA.n1129 GNDA.n1128 185
R1005 GNDA.n1127 GNDA.n1126 185
R1006 GNDA.n1125 GNDA.n1124 185
R1007 GNDA.n1123 GNDA.n1122 185
R1008 GNDA.n1121 GNDA.n1120 185
R1009 GNDA.n1119 GNDA.n1118 185
R1010 GNDA.n1117 GNDA.n1116 185
R1011 GNDA.n1115 GNDA.n1114 185
R1012 GNDA.n1113 GNDA.n1112 185
R1013 GNDA.n1131 GNDA.n1130 185
R1014 GNDA.n1132 GNDA.n1062 185
R1015 GNDA.t80 GNDA.n1062 185
R1016 GNDA.n1134 GNDA.n1133 185
R1017 GNDA.n1136 GNDA.n1135 185
R1018 GNDA.n1138 GNDA.n1137 185
R1019 GNDA.n1140 GNDA.n1139 185
R1020 GNDA.n1142 GNDA.n1141 185
R1021 GNDA.n1144 GNDA.n1143 185
R1022 GNDA.n1146 GNDA.n1145 185
R1023 GNDA.n1073 GNDA.n1053 185
R1024 GNDA.n1161 GNDA.n1160 185
R1025 GNDA.n1159 GNDA.n1072 185
R1026 GNDA.n1158 GNDA.n1157 185
R1027 GNDA.n1156 GNDA.n1155 185
R1028 GNDA.n1154 GNDA.n1153 185
R1029 GNDA.n1152 GNDA.n1151 185
R1030 GNDA.n1150 GNDA.n1149 185
R1031 GNDA.n1148 GNDA.n1147 185
R1032 GNDA.n666 GNDA.n646 185
R1033 GNDA.n665 GNDA.n664 185
R1034 GNDA.n663 GNDA.n662 185
R1035 GNDA.n661 GNDA.n648 185
R1036 GNDA.n659 GNDA.n658 185
R1037 GNDA.n657 GNDA.n649 185
R1038 GNDA.n656 GNDA.n655 185
R1039 GNDA.n653 GNDA.n651 185
R1040 GNDA.n650 GNDA.n628 185
R1041 GNDA.n669 GNDA.n668 185
R1042 GNDA.n670 GNDA.n645 185
R1043 GNDA.n645 GNDA.t76 185
R1044 GNDA.n672 GNDA.n671 185
R1045 GNDA.n674 GNDA.n644 185
R1046 GNDA.n677 GNDA.n676 185
R1047 GNDA.n678 GNDA.n643 185
R1048 GNDA.n680 GNDA.n679 185
R1049 GNDA.n682 GNDA.n642 185
R1050 GNDA.n685 GNDA.n684 185
R1051 GNDA.n702 GNDA.n637 185
R1052 GNDA.n701 GNDA.n700 185
R1053 GNDA.n698 GNDA.n638 185
R1054 GNDA.n696 GNDA.n695 185
R1055 GNDA.n694 GNDA.n639 185
R1056 GNDA.n693 GNDA.n692 185
R1057 GNDA.n690 GNDA.n640 185
R1058 GNDA.n688 GNDA.n687 185
R1059 GNDA.n686 GNDA.n641 185
R1060 GNDA.n740 GNDA.n739 185
R1061 GNDA.n737 GNDA.n736 185
R1062 GNDA.n630 GNDA.n629 185
R1063 GNDA.n730 GNDA.n729 185
R1064 GNDA.n727 GNDA.n632 185
R1065 GNDA.n725 GNDA.n724 185
R1066 GNDA.n715 GNDA.n633 185
R1067 GNDA.n714 GNDA.n713 185
R1068 GNDA.n711 GNDA.n710 185
R1069 GNDA.n711 GNDA.t76 185
R1070 GNDA.n1828 GNDA.n1827 185
R1071 GNDA.n1827 GNDA.n1826 185
R1072 GNDA.n1821 GNDA.n195 185
R1073 GNDA.n1828 GNDA.n195 185
R1074 GNDA.n1616 GNDA.n1615 185
R1075 GNDA.n1613 GNDA.n1612 185
R1076 GNDA.n1871 GNDA.n1870 185
R1077 GNDA.n1869 GNDA.n1868 185
R1078 GNDA.n1867 GNDA.n1866 185
R1079 GNDA.n1865 GNDA.n1864 185
R1080 GNDA.n1863 GNDA.n1862 185
R1081 GNDA.n1861 GNDA.n1860 185
R1082 GNDA.n1859 GNDA.n1858 185
R1083 GNDA.n1857 GNDA.n1856 185
R1084 GNDA.n1855 GNDA.n1854 185
R1085 GNDA.n1873 GNDA.n1872 185
R1086 GNDA.n1874 GNDA.n159 185
R1087 GNDA.t79 GNDA.n159 185
R1088 GNDA.n1876 GNDA.n1875 185
R1089 GNDA.n1878 GNDA.n1877 185
R1090 GNDA.n1880 GNDA.n1879 185
R1091 GNDA.n1882 GNDA.n1881 185
R1092 GNDA.n1884 GNDA.n1883 185
R1093 GNDA.n1886 GNDA.n1885 185
R1094 GNDA.n1888 GNDA.n1887 185
R1095 GNDA.n150 GNDA.n148 185
R1096 GNDA.n1903 GNDA.n1902 185
R1097 GNDA.n1901 GNDA.n169 185
R1098 GNDA.n1900 GNDA.n1899 185
R1099 GNDA.n1898 GNDA.n1897 185
R1100 GNDA.n1896 GNDA.n1895 185
R1101 GNDA.n1894 GNDA.n1893 185
R1102 GNDA.n1892 GNDA.n1891 185
R1103 GNDA.n1890 GNDA.n1889 185
R1104 GNDA.n1853 GNDA.n1852 185
R1105 GNDA.n1843 GNDA.n1842 185
R1106 GNDA.n1841 GNDA.n1840 185
R1107 GNDA.n1838 GNDA.n1837 185
R1108 GNDA.n1836 GNDA.n1835 185
R1109 GNDA.n187 GNDA.n186 185
R1110 GNDA.n185 GNDA.n184 185
R1111 GNDA.n182 GNDA.n151 185
R1112 GNDA.n1906 GNDA.n1905 185
R1113 GNDA.n1905 GNDA.t79 185
R1114 GNDA.n914 GNDA.n824 185
R1115 GNDA.n916 GNDA.n915 185
R1116 GNDA.n918 GNDA.n822 185
R1117 GNDA.n920 GNDA.n919 185
R1118 GNDA.n921 GNDA.n821 185
R1119 GNDA.n923 GNDA.n922 185
R1120 GNDA.n925 GNDA.n820 185
R1121 GNDA.n926 GNDA.n818 185
R1122 GNDA.n929 GNDA.n928 185
R1123 GNDA.n913 GNDA.n912 185
R1124 GNDA.n910 GNDA.n825 185
R1125 GNDA.n910 GNDA.t85 185
R1126 GNDA.n909 GNDA.n826 185
R1127 GNDA.n907 GNDA.n906 185
R1128 GNDA.n905 GNDA.n827 185
R1129 GNDA.n904 GNDA.n903 185
R1130 GNDA.n901 GNDA.n828 185
R1131 GNDA.n899 GNDA.n898 185
R1132 GNDA.n897 GNDA.n829 185
R1133 GNDA.n880 GNDA.n879 185
R1134 GNDA.n881 GNDA.n833 185
R1135 GNDA.n883 GNDA.n882 185
R1136 GNDA.n885 GNDA.n832 185
R1137 GNDA.n888 GNDA.n887 185
R1138 GNDA.n889 GNDA.n831 185
R1139 GNDA.n891 GNDA.n890 185
R1140 GNDA.n893 GNDA.n830 185
R1141 GNDA.n896 GNDA.n895 185
R1142 GNDA.n819 GNDA.n817 185
R1143 GNDA.n853 GNDA.n852 185
R1144 GNDA.n859 GNDA.n858 185
R1145 GNDA.n856 GNDA.n855 185
R1146 GNDA.n854 GNDA.n844 185
R1147 GNDA.n867 GNDA.n866 185
R1148 GNDA.n870 GNDA.n869 185
R1149 GNDA.n837 GNDA.n835 185
R1150 GNDA.n877 GNDA.n876 185
R1151 GNDA.n877 GNDA.t85 185
R1152 GNDA.n545 GNDA.n544 185
R1153 GNDA.n543 GNDA.n542 185
R1154 GNDA.n541 GNDA.n540 185
R1155 GNDA.n539 GNDA.n538 185
R1156 GNDA.n537 GNDA.n536 185
R1157 GNDA.n535 GNDA.n534 185
R1158 GNDA.n533 GNDA.n532 185
R1159 GNDA.n531 GNDA.n530 185
R1160 GNDA.n451 GNDA.n437 185
R1161 GNDA.n547 GNDA.n546 185
R1162 GNDA.n548 GNDA.n449 185
R1163 GNDA.t91 GNDA.n449 185
R1164 GNDA.n550 GNDA.n549 185
R1165 GNDA.n552 GNDA.n551 185
R1166 GNDA.n554 GNDA.n553 185
R1167 GNDA.n556 GNDA.n555 185
R1168 GNDA.n558 GNDA.n557 185
R1169 GNDA.n560 GNDA.n559 185
R1170 GNDA.n562 GNDA.n561 185
R1171 GNDA.n579 GNDA.n461 185
R1172 GNDA.n578 GNDA.n577 185
R1173 GNDA.n576 GNDA.n575 185
R1174 GNDA.n574 GNDA.n573 185
R1175 GNDA.n572 GNDA.n571 185
R1176 GNDA.n570 GNDA.n569 185
R1177 GNDA.n568 GNDA.n567 185
R1178 GNDA.n566 GNDA.n565 185
R1179 GNDA.n564 GNDA.n563 185
R1180 GNDA.n442 GNDA.n438 185
R1181 GNDA.n614 GNDA.n613 185
R1182 GNDA.n594 GNDA.n441 185
R1183 GNDA.n593 GNDA.n592 185
R1184 GNDA.n591 GNDA.n587 185
R1185 GNDA.n602 GNDA.n601 185
R1186 GNDA.n604 GNDA.n603 185
R1187 GNDA.n464 GNDA.n462 185
R1188 GNDA.n611 GNDA.n610 185
R1189 GNDA.t91 GNDA.n611 185
R1190 GNDA.n1299 GNDA.n1298 185
R1191 GNDA.n1297 GNDA.n1296 185
R1192 GNDA.n1295 GNDA.n1294 185
R1193 GNDA.n1293 GNDA.n1292 185
R1194 GNDA.n1291 GNDA.n1290 185
R1195 GNDA.n1289 GNDA.n1288 185
R1196 GNDA.n1287 GNDA.n1286 185
R1197 GNDA.n1285 GNDA.n1284 185
R1198 GNDA.n1283 GNDA.n1282 185
R1199 GNDA.n1301 GNDA.n1300 185
R1200 GNDA.n1302 GNDA.n1232 185
R1201 GNDA.t90 GNDA.n1232 185
R1202 GNDA.n1304 GNDA.n1303 185
R1203 GNDA.n1306 GNDA.n1305 185
R1204 GNDA.n1308 GNDA.n1307 185
R1205 GNDA.n1310 GNDA.n1309 185
R1206 GNDA.n1312 GNDA.n1311 185
R1207 GNDA.n1314 GNDA.n1313 185
R1208 GNDA.n1316 GNDA.n1315 185
R1209 GNDA.n1243 GNDA.n1223 185
R1210 GNDA.n1331 GNDA.n1330 185
R1211 GNDA.n1329 GNDA.n1242 185
R1212 GNDA.n1328 GNDA.n1327 185
R1213 GNDA.n1326 GNDA.n1325 185
R1214 GNDA.n1324 GNDA.n1323 185
R1215 GNDA.n1322 GNDA.n1321 185
R1216 GNDA.n1320 GNDA.n1319 185
R1217 GNDA.n1318 GNDA.n1317 185
R1218 GNDA.n1281 GNDA.n1280 185
R1219 GNDA.n1271 GNDA.n1270 185
R1220 GNDA.n1269 GNDA.n1268 185
R1221 GNDA.n1266 GNDA.n1265 185
R1222 GNDA.n1264 GNDA.n1263 185
R1223 GNDA.n1255 GNDA.n1254 185
R1224 GNDA.n1253 GNDA.n1252 185
R1225 GNDA.n1250 GNDA.n1224 185
R1226 GNDA.n1334 GNDA.n1333 185
R1227 GNDA.n1333 GNDA.t90 185
R1228 GNDA.n350 GNDA.n259 185
R1229 GNDA.n352 GNDA.n351 185
R1230 GNDA.n354 GNDA.n257 185
R1231 GNDA.n356 GNDA.n355 185
R1232 GNDA.n357 GNDA.n256 185
R1233 GNDA.n359 GNDA.n358 185
R1234 GNDA.n361 GNDA.n255 185
R1235 GNDA.n362 GNDA.n253 185
R1236 GNDA.n365 GNDA.n364 185
R1237 GNDA.n349 GNDA.n348 185
R1238 GNDA.n346 GNDA.n260 185
R1239 GNDA.n346 GNDA.t86 185
R1240 GNDA.n345 GNDA.n261 185
R1241 GNDA.n343 GNDA.n342 185
R1242 GNDA.n341 GNDA.n262 185
R1243 GNDA.n340 GNDA.n339 185
R1244 GNDA.n337 GNDA.n263 185
R1245 GNDA.n335 GNDA.n334 185
R1246 GNDA.n333 GNDA.n264 185
R1247 GNDA.n316 GNDA.n315 185
R1248 GNDA.n317 GNDA.n268 185
R1249 GNDA.n319 GNDA.n318 185
R1250 GNDA.n321 GNDA.n267 185
R1251 GNDA.n324 GNDA.n323 185
R1252 GNDA.n325 GNDA.n266 185
R1253 GNDA.n327 GNDA.n326 185
R1254 GNDA.n329 GNDA.n265 185
R1255 GNDA.n332 GNDA.n331 185
R1256 GNDA.n254 GNDA.n252 185
R1257 GNDA.n289 GNDA.n288 185
R1258 GNDA.n295 GNDA.n294 185
R1259 GNDA.n292 GNDA.n291 185
R1260 GNDA.n290 GNDA.n280 185
R1261 GNDA.n303 GNDA.n302 185
R1262 GNDA.n306 GNDA.n305 185
R1263 GNDA.n272 GNDA.n270 185
R1264 GNDA.n313 GNDA.n312 185
R1265 GNDA.n313 GNDA.t86 185
R1266 GNDA.n1111 GNDA.n1110 185
R1267 GNDA.n1102 GNDA.n1101 185
R1268 GNDA.n1100 GNDA.n1099 185
R1269 GNDA.n1097 GNDA.n1096 185
R1270 GNDA.n1095 GNDA.n1094 185
R1271 GNDA.n1086 GNDA.n1085 185
R1272 GNDA.n1084 GNDA.n1083 185
R1273 GNDA.n1081 GNDA.n1054 185
R1274 GNDA.n1164 GNDA.n1163 185
R1275 GNDA.n1163 GNDA.t80 185
R1276 GNDA.n1765 GNDA.n1743 185
R1277 GNDA.n1764 GNDA.n1763 185
R1278 GNDA.n1762 GNDA.n1761 185
R1279 GNDA.n1760 GNDA.n1745 185
R1280 GNDA.n1758 GNDA.n1757 185
R1281 GNDA.n1756 GNDA.n1746 185
R1282 GNDA.n1755 GNDA.n1754 185
R1283 GNDA.n1752 GNDA.n1750 185
R1284 GNDA.n1749 GNDA.n10 185
R1285 GNDA.n1768 GNDA.n1767 185
R1286 GNDA.n1769 GNDA.n1742 185
R1287 GNDA.n1742 GNDA.t78 185
R1288 GNDA.n1771 GNDA.n1770 185
R1289 GNDA.n1773 GNDA.n1741 185
R1290 GNDA.n1776 GNDA.n1775 185
R1291 GNDA.n1777 GNDA.n1740 185
R1292 GNDA.n1779 GNDA.n1778 185
R1293 GNDA.n1781 GNDA.n1739 185
R1294 GNDA.n1784 GNDA.n1783 185
R1295 GNDA.n1801 GNDA.n1800 185
R1296 GNDA.n1799 GNDA.n1798 185
R1297 GNDA.n1797 GNDA.n1735 185
R1298 GNDA.n1795 GNDA.n1794 185
R1299 GNDA.n1793 GNDA.n1736 185
R1300 GNDA.n1792 GNDA.n1791 185
R1301 GNDA.n1789 GNDA.n1737 185
R1302 GNDA.n1787 GNDA.n1786 185
R1303 GNDA.n1785 GNDA.n1738 185
R1304 GNDA.n2051 GNDA.n2050 185
R1305 GNDA.n2048 GNDA.n8 185
R1306 GNDA.n2047 GNDA.n3 185
R1307 GNDA.n2045 GNDA.n2 185
R1308 GNDA.n2044 GNDA.n12 185
R1309 GNDA.n2042 GNDA.n2041 185
R1310 GNDA.n1803 GNDA.n13 185
R1311 GNDA.n1810 GNDA.n1809 185
R1312 GNDA.n1812 GNDA.n1811 185
R1313 GNDA.n1811 GNDA.t78 185
R1314 GNDA.n1641 GNDA.n1640 185
R1315 GNDA.n1631 GNDA.n1630 185
R1316 GNDA.n1629 GNDA.n1628 185
R1317 GNDA.n1626 GNDA.n1625 185
R1318 GNDA.n1624 GNDA.n1623 185
R1319 GNDA.n1597 GNDA.n1596 185
R1320 GNDA.n1595 GNDA.n1594 185
R1321 GNDA.n1592 GNDA.n1561 185
R1322 GNDA.n1694 GNDA.n1693 185
R1323 GNDA.n1693 GNDA.t92 185
R1324 GNDA.n1405 GNDA.t77 183.948
R1325 GNDA.t77 GNDA.n417 183.948
R1326 GNDA.t77 GNDA.n49 180.023
R1327 GNDA.n1387 GNDA.t77 180.013
R1328 GNDA.t77 GNDA.n215 180.013
R1329 GNDA.n1445 GNDA.n228 175.546
R1330 GNDA.n1449 GNDA.n1447 175.546
R1331 GNDA.n1457 GNDA.n224 175.546
R1332 GNDA.n1464 GNDA.n1459 175.546
R1333 GNDA.n1462 GNDA.n1461 175.546
R1334 GNDA.n1406 GNDA.n1391 175.546
R1335 GNDA.n1402 GNDA.n1391 175.546
R1336 GNDA.n1402 GNDA.n1394 175.546
R1337 GNDA.n1398 GNDA.n1394 175.546
R1338 GNDA.n1398 GNDA.n209 175.546
R1339 GNDA.n1484 GNDA.n209 175.546
R1340 GNDA.n1484 GNDA.n210 175.546
R1341 GNDA.n1480 GNDA.n210 175.546
R1342 GNDA.n1480 GNDA.n214 175.546
R1343 GNDA.n1476 GNDA.n214 175.546
R1344 GNDA.n1476 GNDA.n216 175.546
R1345 GNDA.n1427 GNDA.n1426 175.546
R1346 GNDA.n1423 GNDA.n1422 175.546
R1347 GNDA.n1420 GNDA.n1176 175.546
R1348 GNDA.n1416 GNDA.n1414 175.546
R1349 GNDA.n1412 GNDA.n1181 175.546
R1350 GNDA.n1166 GNDA.n1051 175.546
R1351 GNDA.n1088 GNDA.n1080 175.546
R1352 GNDA.n1092 GNDA.n1090 175.546
R1353 GNDA.n1104 GNDA.n1077 175.546
R1354 GNDA.n1108 GNDA.n1106 175.546
R1355 GNDA.n2001 GNDA.n74 175.546
R1356 GNDA.n1999 GNDA.n1998 175.546
R1357 GNDA.n1995 GNDA.n1994 175.546
R1358 GNDA.n1991 GNDA.n1990 175.546
R1359 GNDA.n1987 GNDA.n1986 175.546
R1360 GNDA.n1814 GNDA.n1729 175.546
R1361 GNDA.n1814 GNDA.n1730 175.546
R1362 GNDA.n1807 GNDA.n1730 175.546
R1363 GNDA.n1807 GNDA.n15 175.546
R1364 GNDA.n2039 GNDA.n15 175.546
R1365 GNDA.n2039 GNDA.n4 175.546
R1366 GNDA.n2057 GNDA.n4 175.546
R1367 GNDA.n2057 GNDA.n5 175.546
R1368 GNDA.n2053 GNDA.n5 175.546
R1369 GNDA.n2053 GNDA.n6 175.546
R1370 GNDA.n131 GNDA.n6 175.546
R1371 GNDA.n1931 GNDA.n127 175.546
R1372 GNDA.n1935 GNDA.n1933 175.546
R1373 GNDA.n1943 GNDA.n123 175.546
R1374 GNDA.n1949 GNDA.n1945 175.546
R1375 GNDA.n1947 GNDA.n1946 175.546
R1376 GNDA.n1979 GNDA.n1978 175.546
R1377 GNDA.n1975 GNDA.n1974 175.546
R1378 GNDA.n1971 GNDA.n1970 175.546
R1379 GNDA.n1967 GNDA.n1966 175.546
R1380 GNDA.n1963 GNDA.n1962 175.546
R1381 GNDA.n752 GNDA.n751 175.546
R1382 GNDA.n757 GNDA.n754 175.546
R1383 GNDA.n760 GNDA.n759 175.546
R1384 GNDA.n765 GNDA.n762 175.546
R1385 GNDA.n768 GNDA.n767 175.546
R1386 GNDA.n780 GNDA.n777 175.546
R1387 GNDA.n784 GNDA.n782 175.546
R1388 GNDA.n788 GNDA.n774 175.546
R1389 GNDA.n791 GNDA.n790 175.546
R1390 GNDA.n795 GNDA.n794 175.546
R1391 GNDA.n1018 GNDA.n1016 175.546
R1392 GNDA.n1026 GNDA.n430 175.546
R1393 GNDA.n1030 GNDA.n1028 175.546
R1394 GNDA.n1041 GNDA.n426 175.546
R1395 GNDA.n1044 GNDA.n1043 175.546
R1396 GNDA.n708 GNDA.n707 175.546
R1397 GNDA.n718 GNDA.n717 175.546
R1398 GNDA.n722 GNDA.n721 175.546
R1399 GNDA.n734 GNDA.n732 175.546
R1400 GNDA.n742 GNDA.n626 175.546
R1401 GNDA.n1910 GNDA.n147 175.546
R1402 GNDA.n177 GNDA.n147 175.546
R1403 GNDA.n181 GNDA.n177 175.546
R1404 GNDA.n189 GNDA.n181 175.546
R1405 GNDA.n189 GNDA.n176 175.546
R1406 GNDA.n1833 GNDA.n176 175.546
R1407 GNDA.n1833 GNDA.n174 175.546
R1408 GNDA.n1845 GNDA.n174 175.546
R1409 GNDA.n1845 GNDA.n173 175.546
R1410 GNDA.n1850 GNDA.n173 175.546
R1411 GNDA.n1850 GNDA.n18 175.546
R1412 GNDA.n1929 GNDA.n1927 175.546
R1413 GNDA.n1937 GNDA.n125 175.546
R1414 GNDA.n1941 GNDA.n1939 175.546
R1415 GNDA.n1951 GNDA.n121 175.546
R1416 GNDA.n1954 GNDA.n1953 175.546
R1417 GNDA.n116 GNDA.n115 175.546
R1418 GNDA.n112 GNDA.n111 175.546
R1419 GNDA.n108 GNDA.n107 175.546
R1420 GNDA.n104 GNDA.n103 175.546
R1421 GNDA.n100 GNDA.n30 175.546
R1422 GNDA.n2029 GNDA.n21 175.546
R1423 GNDA.n2025 GNDA.n2024 175.546
R1424 GNDA.n2022 GNDA.n24 175.546
R1425 GNDA.n2018 GNDA.n2017 175.546
R1426 GNDA.n2015 GNDA.n27 175.546
R1427 GNDA.n941 GNDA.n814 175.546
R1428 GNDA.n945 GNDA.n943 175.546
R1429 GNDA.n949 GNDA.n812 175.546
R1430 GNDA.n953 GNDA.n951 175.546
R1431 GNDA.n957 GNDA.n810 175.546
R1432 GNDA.n978 GNDA.n801 175.546
R1433 GNDA.n974 GNDA.n973 175.546
R1434 GNDA.n971 GNDA.n804 175.546
R1435 GNDA.n967 GNDA.n966 175.546
R1436 GNDA.n964 GNDA.n807 175.546
R1437 GNDA.n1001 GNDA.n1000 175.546
R1438 GNDA.n997 GNDA.n996 175.546
R1439 GNDA.n994 GNDA.n756 175.546
R1440 GNDA.n990 GNDA.n988 175.546
R1441 GNDA.n986 GNDA.n764 175.546
R1442 GNDA.n874 GNDA.n840 175.546
R1443 GNDA.n872 GNDA.n841 175.546
R1444 GNDA.n864 GNDA.n863 175.546
R1445 GNDA.n861 GNDA.n848 175.546
R1446 GNDA.n932 GNDA.n816 175.546
R1447 GNDA.n1698 GNDA.n1499 175.546
R1448 GNDA.n1587 GNDA.n1499 175.546
R1449 GNDA.n1591 GNDA.n1587 175.546
R1450 GNDA.n1599 GNDA.n1591 175.546
R1451 GNDA.n1599 GNDA.n1586 175.546
R1452 GNDA.n1621 GNDA.n1586 175.546
R1453 GNDA.n1621 GNDA.n1584 175.546
R1454 GNDA.n1633 GNDA.n1584 175.546
R1455 GNDA.n1633 GNDA.n1583 175.546
R1456 GNDA.n1638 GNDA.n1583 175.546
R1457 GNDA.n1638 GNDA.n200 175.546
R1458 GNDA.n80 GNDA.n79 175.546
R1459 GNDA.n83 GNDA.n82 175.546
R1460 GNDA.n86 GNDA.n85 175.546
R1461 GNDA.n89 GNDA.n88 175.546
R1462 GNDA.n92 GNDA.n91 175.546
R1463 GNDA.n1531 GNDA.n1530 175.546
R1464 GNDA.n1527 GNDA.n1526 175.546
R1465 GNDA.n1523 GNDA.n1522 175.546
R1466 GNDA.n1519 GNDA.n1518 175.546
R1467 GNDA.n1515 GNDA.n1514 175.546
R1468 GNDA.n1556 GNDA.n1502 175.546
R1469 GNDA.n1552 GNDA.n1502 175.546
R1470 GNDA.n1552 GNDA.n1504 175.546
R1471 GNDA.n1548 GNDA.n1504 175.546
R1472 GNDA.n1548 GNDA.n1546 175.546
R1473 GNDA.n1546 GNDA.n1545 175.546
R1474 GNDA.n1545 GNDA.n1506 175.546
R1475 GNDA.n1541 GNDA.n1506 175.546
R1476 GNDA.n1541 GNDA.n1508 175.546
R1477 GNDA.n1537 GNDA.n1508 175.546
R1478 GNDA.n1537 GNDA.n1510 175.546
R1479 GNDA.n1020 GNDA.n432 175.546
R1480 GNDA.n1024 GNDA.n1022 175.546
R1481 GNDA.n1032 GNDA.n428 175.546
R1482 GNDA.n1039 GNDA.n1034 175.546
R1483 GNDA.n1037 GNDA.n1036 175.546
R1484 GNDA.n502 GNDA.n501 175.546
R1485 GNDA.n499 GNDA.n479 175.546
R1486 GNDA.n495 GNDA.n494 175.546
R1487 GNDA.n492 GNDA.n482 175.546
R1488 GNDA.n488 GNDA.n487 175.546
R1489 GNDA.n527 GNDA.n467 175.546
R1490 GNDA.n523 GNDA.n467 175.546
R1491 GNDA.n523 GNDA.n469 175.546
R1492 GNDA.n519 GNDA.n469 175.546
R1493 GNDA.n519 GNDA.n517 175.546
R1494 GNDA.n517 GNDA.n516 175.546
R1495 GNDA.n516 GNDA.n471 175.546
R1496 GNDA.n512 GNDA.n471 175.546
R1497 GNDA.n512 GNDA.n473 175.546
R1498 GNDA.n508 GNDA.n473 175.546
R1499 GNDA.n508 GNDA.n476 175.546
R1500 GNDA.n608 GNDA.n584 175.546
R1501 GNDA.n606 GNDA.n585 175.546
R1502 GNDA.n599 GNDA.n598 175.546
R1503 GNDA.n596 GNDA.n590 175.546
R1504 GNDA.n617 GNDA.n616 175.546
R1505 GNDA.n1191 GNDA.n1173 175.546
R1506 GNDA.n1194 GNDA.n1174 175.546
R1507 GNDA.n1178 GNDA.n1177 175.546
R1508 GNDA.n1197 GNDA.n1179 175.546
R1509 GNDA.n1183 GNDA.n1182 175.546
R1510 GNDA.n1368 GNDA.n1208 175.546
R1511 GNDA.n1368 GNDA.n1206 175.546
R1512 GNDA.n1372 GNDA.n1206 175.546
R1513 GNDA.n1372 GNDA.n1204 175.546
R1514 GNDA.n1376 GNDA.n1204 175.546
R1515 GNDA.n1376 GNDA.n1190 175.546
R1516 GNDA.n1380 GNDA.n1190 175.546
R1517 GNDA.n1380 GNDA.n1188 175.546
R1518 GNDA.n1384 GNDA.n1188 175.546
R1519 GNDA.n1384 GNDA.n1186 175.546
R1520 GNDA.n1388 GNDA.n1186 175.546
R1521 GNDA.n1344 GNDA.n1218 175.546
R1522 GNDA.n1344 GNDA.n1216 175.546
R1523 GNDA.n1349 GNDA.n1216 175.546
R1524 GNDA.n1349 GNDA.n1214 175.546
R1525 GNDA.n1353 GNDA.n1214 175.546
R1526 GNDA.n1354 GNDA.n1353 175.546
R1527 GNDA.n1356 GNDA.n1354 175.546
R1528 GNDA.n1356 GNDA.n1212 175.546
R1529 GNDA.n1360 GNDA.n1212 175.546
R1530 GNDA.n1360 GNDA.n1210 175.546
R1531 GNDA.n1364 GNDA.n1210 175.546
R1532 GNDA.n1336 GNDA.n1220 175.546
R1533 GNDA.n1257 GNDA.n1249 175.546
R1534 GNDA.n1261 GNDA.n1259 175.546
R1535 GNDA.n1273 GNDA.n1246 175.546
R1536 GNDA.n1278 GNDA.n1275 175.546
R1537 GNDA.n1443 GNDA.n1441 175.546
R1538 GNDA.n1451 GNDA.n226 175.546
R1539 GNDA.n1455 GNDA.n1453 175.546
R1540 GNDA.n1466 GNDA.n222 175.546
R1541 GNDA.n1469 GNDA.n1468 175.546
R1542 GNDA.n310 GNDA.n276 175.546
R1543 GNDA.n308 GNDA.n277 175.546
R1544 GNDA.n300 GNDA.n299 175.546
R1545 GNDA.n297 GNDA.n284 175.546
R1546 GNDA.n368 GNDA.n251 175.546
R1547 GNDA.n375 GNDA.n249 175.546
R1548 GNDA.n379 GNDA.n377 175.546
R1549 GNDA.n383 GNDA.n247 175.546
R1550 GNDA.n387 GNDA.n385 175.546
R1551 GNDA.n391 GNDA.n245 175.546
R1552 GNDA.n394 GNDA.n393 175.546
R1553 GNDA.n415 GNDA.n220 175.546
R1554 GNDA.n415 GNDA.n236 175.546
R1555 GNDA.n411 GNDA.n236 175.546
R1556 GNDA.n411 GNDA.n408 175.546
R1557 GNDA.n408 GNDA.n407 175.546
R1558 GNDA.n407 GNDA.n238 175.546
R1559 GNDA.n403 GNDA.n238 175.546
R1560 GNDA.n403 GNDA.n240 175.546
R1561 GNDA.n399 GNDA.n240 175.546
R1562 GNDA.n399 GNDA.n242 175.546
R1563 GNDA.n395 GNDA.n242 175.546
R1564 GNDA.n1693 GNDA.n1560 163.333
R1565 GNDA.n1163 GNDA.n1053 163.333
R1566 GNDA.n711 GNDA.n637 163.333
R1567 GNDA.n1905 GNDA.n150 163.333
R1568 GNDA.n879 GNDA.n877 163.333
R1569 GNDA.n611 GNDA.n461 163.333
R1570 GNDA.n1333 GNDA.n1223 163.333
R1571 GNDA.n315 GNDA.n313 163.333
R1572 GNDA.n1811 GNDA.n1801 163.333
R1573 GNDA.n1693 GNDA.n1561 150
R1574 GNDA.n1596 GNDA.n1595 150
R1575 GNDA.n1625 GNDA.n1624 150
R1576 GNDA.n1630 GNDA.n1629 150
R1577 GNDA.n1691 GNDA.n1579 150
R1578 GNDA.n1687 GNDA.n1686 150
R1579 GNDA.n1683 GNDA.n1682 150
R1580 GNDA.n1679 GNDA.n1678 150
R1581 GNDA.n1675 GNDA.n1674 150
R1582 GNDA.n1671 GNDA.n1670 150
R1583 GNDA.n1667 GNDA.n1666 150
R1584 GNDA.n1663 GNDA.n1569 150
R1585 GNDA.n1660 GNDA.n1569 150
R1586 GNDA.n1646 GNDA.n1645 150
R1587 GNDA.n1650 GNDA.n1649 150
R1588 GNDA.n1654 GNDA.n1653 150
R1589 GNDA.n1658 GNDA.n1657 150
R1590 GNDA.n1163 GNDA.n1054 150
R1591 GNDA.n1085 GNDA.n1084 150
R1592 GNDA.n1096 GNDA.n1095 150
R1593 GNDA.n1101 GNDA.n1100 150
R1594 GNDA.n1161 GNDA.n1072 150
R1595 GNDA.n1157 GNDA.n1156 150
R1596 GNDA.n1153 GNDA.n1152 150
R1597 GNDA.n1149 GNDA.n1148 150
R1598 GNDA.n1145 GNDA.n1144 150
R1599 GNDA.n1141 GNDA.n1140 150
R1600 GNDA.n1137 GNDA.n1136 150
R1601 GNDA.n1133 GNDA.n1062 150
R1602 GNDA.n1130 GNDA.n1062 150
R1603 GNDA.n1116 GNDA.n1115 150
R1604 GNDA.n1120 GNDA.n1119 150
R1605 GNDA.n1124 GNDA.n1123 150
R1606 GNDA.n1128 GNDA.n1127 150
R1607 GNDA.n713 GNDA.n711 150
R1608 GNDA.n725 GNDA.n633 150
R1609 GNDA.n729 GNDA.n727 150
R1610 GNDA.n737 GNDA.n629 150
R1611 GNDA.n700 GNDA.n698 150
R1612 GNDA.n696 GNDA.n639 150
R1613 GNDA.n692 GNDA.n690 150
R1614 GNDA.n688 GNDA.n641 150
R1615 GNDA.n684 GNDA.n682 150
R1616 GNDA.n680 GNDA.n643 150
R1617 GNDA.n676 GNDA.n674 150
R1618 GNDA.n672 GNDA.n645 150
R1619 GNDA.n668 GNDA.n645 150
R1620 GNDA.n655 GNDA.n653 150
R1621 GNDA.n659 GNDA.n649 150
R1622 GNDA.n662 GNDA.n661 150
R1623 GNDA.n666 GNDA.n665 150
R1624 GNDA.n1905 GNDA.n151 150
R1625 GNDA.n186 GNDA.n185 150
R1626 GNDA.n1837 GNDA.n1836 150
R1627 GNDA.n1842 GNDA.n1841 150
R1628 GNDA.n1903 GNDA.n169 150
R1629 GNDA.n1899 GNDA.n1898 150
R1630 GNDA.n1895 GNDA.n1894 150
R1631 GNDA.n1891 GNDA.n1890 150
R1632 GNDA.n1887 GNDA.n1886 150
R1633 GNDA.n1883 GNDA.n1882 150
R1634 GNDA.n1879 GNDA.n1878 150
R1635 GNDA.n1875 GNDA.n159 150
R1636 GNDA.n1872 GNDA.n159 150
R1637 GNDA.n1858 GNDA.n1857 150
R1638 GNDA.n1862 GNDA.n1861 150
R1639 GNDA.n1866 GNDA.n1865 150
R1640 GNDA.n1870 GNDA.n1869 150
R1641 GNDA.n877 GNDA.n835 150
R1642 GNDA.n869 GNDA.n867 150
R1643 GNDA.n856 GNDA.n854 150
R1644 GNDA.n858 GNDA.n853 150
R1645 GNDA.n883 GNDA.n833 150
R1646 GNDA.n887 GNDA.n885 150
R1647 GNDA.n891 GNDA.n831 150
R1648 GNDA.n895 GNDA.n893 150
R1649 GNDA.n899 GNDA.n829 150
R1650 GNDA.n903 GNDA.n901 150
R1651 GNDA.n907 GNDA.n827 150
R1652 GNDA.n910 GNDA.n909 150
R1653 GNDA.n912 GNDA.n910 150
R1654 GNDA.n926 GNDA.n925 150
R1655 GNDA.n923 GNDA.n821 150
R1656 GNDA.n919 GNDA.n918 150
R1657 GNDA.n916 GNDA.n824 150
R1658 GNDA.n611 GNDA.n462 150
R1659 GNDA.n603 GNDA.n602 150
R1660 GNDA.n592 GNDA.n591 150
R1661 GNDA.n613 GNDA.n441 150
R1662 GNDA.n577 GNDA.n576 150
R1663 GNDA.n573 GNDA.n572 150
R1664 GNDA.n569 GNDA.n568 150
R1665 GNDA.n565 GNDA.n564 150
R1666 GNDA.n561 GNDA.n560 150
R1667 GNDA.n557 GNDA.n556 150
R1668 GNDA.n553 GNDA.n552 150
R1669 GNDA.n549 GNDA.n449 150
R1670 GNDA.n546 GNDA.n449 150
R1671 GNDA.n532 GNDA.n531 150
R1672 GNDA.n536 GNDA.n535 150
R1673 GNDA.n540 GNDA.n539 150
R1674 GNDA.n544 GNDA.n543 150
R1675 GNDA.n1333 GNDA.n1224 150
R1676 GNDA.n1254 GNDA.n1253 150
R1677 GNDA.n1265 GNDA.n1264 150
R1678 GNDA.n1270 GNDA.n1269 150
R1679 GNDA.n1331 GNDA.n1242 150
R1680 GNDA.n1327 GNDA.n1326 150
R1681 GNDA.n1323 GNDA.n1322 150
R1682 GNDA.n1319 GNDA.n1318 150
R1683 GNDA.n1315 GNDA.n1314 150
R1684 GNDA.n1311 GNDA.n1310 150
R1685 GNDA.n1307 GNDA.n1306 150
R1686 GNDA.n1303 GNDA.n1232 150
R1687 GNDA.n1300 GNDA.n1232 150
R1688 GNDA.n1286 GNDA.n1285 150
R1689 GNDA.n1290 GNDA.n1289 150
R1690 GNDA.n1294 GNDA.n1293 150
R1691 GNDA.n1298 GNDA.n1297 150
R1692 GNDA.n313 GNDA.n270 150
R1693 GNDA.n305 GNDA.n303 150
R1694 GNDA.n292 GNDA.n290 150
R1695 GNDA.n294 GNDA.n289 150
R1696 GNDA.n319 GNDA.n268 150
R1697 GNDA.n323 GNDA.n321 150
R1698 GNDA.n327 GNDA.n266 150
R1699 GNDA.n331 GNDA.n329 150
R1700 GNDA.n335 GNDA.n264 150
R1701 GNDA.n339 GNDA.n337 150
R1702 GNDA.n343 GNDA.n262 150
R1703 GNDA.n346 GNDA.n345 150
R1704 GNDA.n348 GNDA.n346 150
R1705 GNDA.n362 GNDA.n361 150
R1706 GNDA.n359 GNDA.n256 150
R1707 GNDA.n355 GNDA.n354 150
R1708 GNDA.n352 GNDA.n259 150
R1709 GNDA.n1811 GNDA.n1810 150
R1710 GNDA.n2042 GNDA.n13 150
R1711 GNDA.n2045 GNDA.n2044 150
R1712 GNDA.n2048 GNDA.n2047 150
R1713 GNDA.n1798 GNDA.n1797 150
R1714 GNDA.n1795 GNDA.n1736 150
R1715 GNDA.n1791 GNDA.n1789 150
R1716 GNDA.n1787 GNDA.n1738 150
R1717 GNDA.n1783 GNDA.n1781 150
R1718 GNDA.n1779 GNDA.n1740 150
R1719 GNDA.n1775 GNDA.n1773 150
R1720 GNDA.n1771 GNDA.n1742 150
R1721 GNDA.n1767 GNDA.n1742 150
R1722 GNDA.n1754 GNDA.n1752 150
R1723 GNDA.n1758 GNDA.n1746 150
R1724 GNDA.n1761 GNDA.n1760 150
R1725 GNDA.n1765 GNDA.n1764 150
R1726 GNDA.n1555 GNDA.n1554 145.964
R1727 GNDA.n1554 GNDA.n1553 145.964
R1728 GNDA.n1553 GNDA.n1503 145.964
R1729 GNDA.n1547 GNDA.n1503 145.964
R1730 GNDA.n1547 GNDA.n63 145.964
R1731 GNDA.n1509 GNDA.n64 145.964
R1732 GNDA.n1540 GNDA.n1509 145.964
R1733 GNDA.n1540 GNDA.n1539 145.964
R1734 GNDA.n1539 GNDA.n1538 145.964
R1735 GNDA.n1538 GNDA.n50 145.964
R1736 GNDA.n526 GNDA.n49 145.964
R1737 GNDA.n526 GNDA.n525 145.964
R1738 GNDA.n525 GNDA.n524 145.964
R1739 GNDA.n524 GNDA.n468 145.964
R1740 GNDA.n518 GNDA.n468 145.964
R1741 GNDA.n518 GNDA.n56 145.964
R1742 GNDA.n474 GNDA.n57 145.964
R1743 GNDA.n511 GNDA.n474 145.964
R1744 GNDA.n511 GNDA.n510 145.964
R1745 GNDA.n510 GNDA.n509 145.964
R1746 GNDA.n509 GNDA.n475 145.964
R1747 GNDA.n1340 GNDA.t12 145.964
R1748 GNDA.n1340 GNDA.n1217 145.964
R1749 GNDA.n1345 GNDA.n1217 145.964
R1750 GNDA.n1346 GNDA.n1345 145.964
R1751 GNDA.n1348 GNDA.n1346 145.964
R1752 GNDA.n1348 GNDA.n1347 145.964
R1753 GNDA.n1347 GNDA.n1201 145.964
R1754 GNDA.n1355 GNDA.n1202 145.964
R1755 GNDA.n1355 GNDA.n1211 145.964
R1756 GNDA.n1361 GNDA.n1211 145.964
R1757 GNDA.n1362 GNDA.n1361 145.964
R1758 GNDA.n1363 GNDA.n1362 145.964
R1759 GNDA.n1705 GNDA.n1704 139.077
R1760 GNDA.n1707 GNDA.n1706 139.077
R1761 GNDA.n1709 GNDA.n1708 139.077
R1762 GNDA.n1715 GNDA.n1714 139.077
R1763 GNDA.n1713 GNDA.n1712 139.077
R1764 GNDA.n1711 GNDA.n1710 139.077
R1765 GNDA.n136 GNDA.n135 139.077
R1766 GNDA.n144 GNDA.n143 139.077
R1767 GNDA.n142 GNDA.n141 139.077
R1768 GNDA.n140 GNDA.n139 139.077
R1769 GNDA.n1495 GNDA.t29 135.69
R1770 GNDA.n1827 GNDA.n197 134.268
R1771 GNDA.n197 GNDA.n195 134.268
R1772 GNDA.n2031 GNDA.n2030 133.517
R1773 GNDA.n937 GNDA.n936 133.517
R1774 GNDA.n1721 GNDA.t84 130.001
R1775 GNDA.n1716 GNDA.t95 130.001
R1776 GNDA.n1918 GNDA.t101 130.001
R1777 GNDA.n1913 GNDA.t104 130.001
R1778 GNDA.n137 GNDA.t98 130.001
R1779 GNDA.n1701 GNDA.t89 130.001
R1780 GNDA.n1437 GNDA.n1435 126.782
R1781 GNDA.n1923 GNDA.n1921 126.782
R1782 GNDA.n747 GNDA.n623 126.782
R1783 GNDA.n1724 GNDA.n77 126.782
R1784 GNDA.n1012 GNDA.n1010 126.782
R1785 GNDA.n1170 GNDA.n234 126.782
R1786 GNDA.n1429 GNDA.n419 124.832
R1787 GNDA.n2005 GNDA.n75 124.832
R1788 GNDA.n1014 GNDA.n434 124.832
R1789 GNDA.n1925 GNDA.n129 124.832
R1790 GNDA.n1003 GNDA.n624 124.832
R1791 GNDA.n1556 GNDA.n1498 124.832
R1792 GNDA.n527 GNDA.n465 124.832
R1793 GNDA.n1339 GNDA.n1218 124.832
R1794 GNDA.n1439 GNDA.n230 124.832
R1795 GNDA.n1491 GNDA.t16 115.948
R1796 GNDA.n1489 GNDA.t10 115.105
R1797 GNDA.n1488 GNDA.t8 114.635
R1798 GNDA.n1491 GNDA.t6 114.635
R1799 GNDA.n1 GNDA.n48 14.555
R1800 GNDA.n0 GNDA.n51 14.555
R1801 GNDA.t94 GNDA.n1727 101.942
R1802 GNDA.n1823 GNDA.n192 101.718
R1803 GNDA.n1608 GNDA.n1602 101.718
R1804 GNDA.n1617 GNDA.n1604 101.718
R1805 GNDA.n1829 GNDA.n194 101.718
R1806 GNDA.t77 GNDA.n64 98.9316
R1807 GNDA.t77 GNDA.n57 98.9316
R1808 GNDA.t77 GNDA.n1202 98.9316
R1809 GNDA.n1920 GNDA.n133 98.8538
R1810 GNDA.n1700 GNDA.n1497 96.7943
R1811 GNDA.n2033 GNDA.n17 95.7646
R1812 GNDA.n1637 GNDA.n1636 92.6754
R1813 GNDA.n1827 GNDA.n1822 91.069
R1814 GNDA.n1825 GNDA.n195 91.069
R1815 GNDA.n1615 GNDA.n1607 91.069
R1816 GNDA.n1615 GNDA.n1614 91.069
R1817 GNDA.n1612 GNDA.n1605 91.069
R1818 GNDA.n1612 GNDA.n1611 91.069
R1819 GNDA.n1911 GNDA.t103 90.616
R1820 GNDA.n1369 GNDA.n1207 88.5317
R1821 GNDA.n1370 GNDA.n1369 88.5317
R1822 GNDA.n1371 GNDA.n1370 88.5317
R1823 GNDA.n1371 GNDA.n1203 88.5317
R1824 GNDA.n1377 GNDA.n1203 88.5317
R1825 GNDA.n1379 GNDA.n1378 88.5317
R1826 GNDA.n1379 GNDA.n1187 88.5317
R1827 GNDA.n1385 GNDA.n1187 88.5317
R1828 GNDA.n1386 GNDA.n1385 88.5317
R1829 GNDA.n1387 GNDA.n1386 88.5317
R1830 GNDA.n1405 GNDA.n1404 88.5317
R1831 GNDA.n1404 GNDA.n1403 88.5317
R1832 GNDA.n1403 GNDA.n1393 88.5317
R1833 GNDA.n1397 GNDA.n1393 88.5317
R1834 GNDA.n1397 GNDA.n206 88.5317
R1835 GNDA.n1485 GNDA.n208 88.5317
R1836 GNDA.n1479 GNDA.n208 88.5317
R1837 GNDA.n1479 GNDA.n1478 88.5317
R1838 GNDA.n1478 GNDA.n1477 88.5317
R1839 GNDA.n1477 GNDA.n215 88.5317
R1840 GNDA.n417 GNDA.n416 88.5317
R1841 GNDA.n416 GNDA.n235 88.5317
R1842 GNDA.n410 GNDA.n235 88.5317
R1843 GNDA.n410 GNDA.n409 88.5317
R1844 GNDA.n409 GNDA.n54 88.5317
R1845 GNDA.n402 GNDA.n55 88.5317
R1846 GNDA.n402 GNDA.n401 88.5317
R1847 GNDA.n401 GNDA.n400 88.5317
R1848 GNDA.n400 GNDA.n241 88.5317
R1849 GNDA.n241 GNDA.n52 88.5317
R1850 GNDA.n2056 GNDA.t64 84.4377
R1851 GNDA.n207 GNDA.n203 84.306
R1852 GNDA.t24 GNDA.t28 82.3782
R1853 GNDA.t110 GNDA.t109 82.3782
R1854 GNDA.n1805 GNDA.t42 80.3188
R1855 GNDA.n1436 GNDA.n228 76.3222
R1856 GNDA.n1447 GNDA.n1446 76.3222
R1857 GNDA.n1448 GNDA.n224 76.3222
R1858 GNDA.n1459 GNDA.n1458 76.3222
R1859 GNDA.n1463 GNDA.n1462 76.3222
R1860 GNDA.n1460 GNDA.n219 76.3222
R1861 GNDA.n1429 GNDA.n1428 76.3222
R1862 GNDA.n1426 GNDA.n1172 76.3222
R1863 GNDA.n1422 GNDA.n1421 76.3222
R1864 GNDA.n1415 GNDA.n1176 76.3222
R1865 GNDA.n1414 GNDA.n1413 76.3222
R1866 GNDA.n1407 GNDA.n1181 76.3222
R1867 GNDA.n1167 GNDA.n1166 76.3222
R1868 GNDA.n1080 GNDA.n1079 76.3222
R1869 GNDA.n1090 GNDA.n1089 76.3222
R1870 GNDA.n1091 GNDA.n1077 76.3222
R1871 GNDA.n1106 GNDA.n1105 76.3222
R1872 GNDA.n1107 GNDA.n232 76.3222
R1873 GNDA.n2006 GNDA.n2005 76.3222
R1874 GNDA.n2001 GNDA.n73 76.3222
R1875 GNDA.n1998 GNDA.n72 76.3222
R1876 GNDA.n1994 GNDA.n71 76.3222
R1877 GNDA.n1990 GNDA.n70 76.3222
R1878 GNDA.n1986 GNDA.n69 76.3222
R1879 GNDA.n1922 GNDA.n127 76.3222
R1880 GNDA.n1933 GNDA.n1932 76.3222
R1881 GNDA.n1934 GNDA.n123 76.3222
R1882 GNDA.n1945 GNDA.n1944 76.3222
R1883 GNDA.n1948 GNDA.n1947 76.3222
R1884 GNDA.n1958 GNDA.n97 76.3222
R1885 GNDA.n1979 GNDA.n36 76.3222
R1886 GNDA.n1975 GNDA.n37 76.3222
R1887 GNDA.n1971 GNDA.n38 76.3222
R1888 GNDA.n1967 GNDA.n39 76.3222
R1889 GNDA.n1963 GNDA.n40 76.3222
R1890 GNDA.n1959 GNDA.n41 76.3222
R1891 GNDA.n751 GNDA.n750 76.3222
R1892 GNDA.n754 GNDA.n753 76.3222
R1893 GNDA.n759 GNDA.n758 76.3222
R1894 GNDA.n762 GNDA.n761 76.3222
R1895 GNDA.n767 GNDA.n766 76.3222
R1896 GNDA.n770 GNDA.n769 76.3222
R1897 GNDA.n777 GNDA.n776 76.3222
R1898 GNDA.n782 GNDA.n781 76.3222
R1899 GNDA.n783 GNDA.n774 76.3222
R1900 GNDA.n790 GNDA.n789 76.3222
R1901 GNDA.n794 GNDA.n772 76.3222
R1902 GNDA.n797 GNDA.n796 76.3222
R1903 GNDA.n1015 GNDA.n1014 76.3222
R1904 GNDA.n1018 GNDA.n1017 76.3222
R1905 GNDA.n1027 GNDA.n1026 76.3222
R1906 GNDA.n1030 GNDA.n1029 76.3222
R1907 GNDA.n1042 GNDA.n1041 76.3222
R1908 GNDA.n1045 GNDA.n1044 76.3222
R1909 GNDA.n708 GNDA.n706 76.3222
R1910 GNDA.n717 GNDA.n635 76.3222
R1911 GNDA.n722 GNDA.n719 76.3222
R1912 GNDA.n732 GNDA.n631 76.3222
R1913 GNDA.n733 GNDA.n626 76.3222
R1914 GNDA.n744 GNDA.n743 76.3222
R1915 GNDA.n1926 GNDA.n1925 76.3222
R1916 GNDA.n1929 GNDA.n1928 76.3222
R1917 GNDA.n1938 GNDA.n1937 76.3222
R1918 GNDA.n1941 GNDA.n1940 76.3222
R1919 GNDA.n1952 GNDA.n1951 76.3222
R1920 GNDA.n1955 GNDA.n1954 76.3222
R1921 GNDA.n116 GNDA.n31 76.3222
R1922 GNDA.n112 GNDA.n32 76.3222
R1923 GNDA.n108 GNDA.n33 76.3222
R1924 GNDA.n104 GNDA.n34 76.3222
R1925 GNDA.n100 GNDA.n35 76.3222
R1926 GNDA.n2010 GNDA.n2009 76.3222
R1927 GNDA.n2030 GNDA.n2029 76.3222
R1928 GNDA.n2025 GNDA.n23 76.3222
R1929 GNDA.n2023 GNDA.n2022 76.3222
R1930 GNDA.n2018 GNDA.n26 76.3222
R1931 GNDA.n2016 GNDA.n2015 76.3222
R1932 GNDA.n2011 GNDA.n29 76.3222
R1933 GNDA.n936 GNDA.n814 76.3222
R1934 GNDA.n943 GNDA.n942 76.3222
R1935 GNDA.n944 GNDA.n812 76.3222
R1936 GNDA.n951 GNDA.n950 76.3222
R1937 GNDA.n952 GNDA.n810 76.3222
R1938 GNDA.n959 GNDA.n958 76.3222
R1939 GNDA.n979 GNDA.n978 76.3222
R1940 GNDA.n974 GNDA.n803 76.3222
R1941 GNDA.n972 GNDA.n971 76.3222
R1942 GNDA.n967 GNDA.n806 76.3222
R1943 GNDA.n965 GNDA.n964 76.3222
R1944 GNDA.n960 GNDA.n809 76.3222
R1945 GNDA.n1003 GNDA.n1002 76.3222
R1946 GNDA.n1000 GNDA.n749 76.3222
R1947 GNDA.n996 GNDA.n995 76.3222
R1948 GNDA.n989 GNDA.n756 76.3222
R1949 GNDA.n988 GNDA.n987 76.3222
R1950 GNDA.n981 GNDA.n764 76.3222
R1951 GNDA.n840 GNDA.n839 76.3222
R1952 GNDA.n873 GNDA.n872 76.3222
R1953 GNDA.n864 GNDA.n845 76.3222
R1954 GNDA.n862 GNDA.n861 76.3222
R1955 GNDA.n847 GNDA.n816 76.3222
R1956 GNDA.n934 GNDA.n933 76.3222
R1957 GNDA.n958 GNDA.n957 76.3222
R1958 GNDA.n953 GNDA.n952 76.3222
R1959 GNDA.n950 GNDA.n949 76.3222
R1960 GNDA.n945 GNDA.n944 76.3222
R1961 GNDA.n942 GNDA.n941 76.3222
R1962 GNDA.n29 GNDA.n27 76.3222
R1963 GNDA.n2017 GNDA.n2016 76.3222
R1964 GNDA.n26 GNDA.n24 76.3222
R1965 GNDA.n2024 GNDA.n2023 76.3222
R1966 GNDA.n23 GNDA.n21 76.3222
R1967 GNDA.n79 GNDA.n78 76.3222
R1968 GNDA.n82 GNDA.n81 76.3222
R1969 GNDA.n85 GNDA.n84 76.3222
R1970 GNDA.n88 GNDA.n87 76.3222
R1971 GNDA.n91 GNDA.n90 76.3222
R1972 GNDA.n94 GNDA.n93 76.3222
R1973 GNDA.n1531 GNDA.n42 76.3222
R1974 GNDA.n1527 GNDA.n43 76.3222
R1975 GNDA.n1523 GNDA.n44 76.3222
R1976 GNDA.n1519 GNDA.n45 76.3222
R1977 GNDA.n1515 GNDA.n46 76.3222
R1978 GNDA.n1511 GNDA.n47 76.3222
R1979 GNDA.n1011 GNDA.n432 76.3222
R1980 GNDA.n1022 GNDA.n1021 76.3222
R1981 GNDA.n1023 GNDA.n428 76.3222
R1982 GNDA.n1034 GNDA.n1033 76.3222
R1983 GNDA.n1038 GNDA.n1037 76.3222
R1984 GNDA.n1035 GNDA.n423 76.3222
R1985 GNDA.n503 GNDA.n502 76.3222
R1986 GNDA.n500 GNDA.n499 76.3222
R1987 GNDA.n495 GNDA.n481 76.3222
R1988 GNDA.n493 GNDA.n492 76.3222
R1989 GNDA.n488 GNDA.n484 76.3222
R1990 GNDA.n486 GNDA.n485 76.3222
R1991 GNDA.n584 GNDA.n583 76.3222
R1992 GNDA.n607 GNDA.n606 76.3222
R1993 GNDA.n599 GNDA.n588 76.3222
R1994 GNDA.n597 GNDA.n596 76.3222
R1995 GNDA.n616 GNDA.n439 76.3222
R1996 GNDA.n621 GNDA.n436 76.3222
R1997 GNDA.n1192 GNDA.n1191 76.3222
R1998 GNDA.n1193 GNDA.n1174 76.3222
R1999 GNDA.n1195 GNDA.n1177 76.3222
R2000 GNDA.n1196 GNDA.n1179 76.3222
R2001 GNDA.n1198 GNDA.n1182 76.3222
R2002 GNDA.n1199 GNDA.n1184 76.3222
R2003 GNDA.n1337 GNDA.n1336 76.3222
R2004 GNDA.n1249 GNDA.n1248 76.3222
R2005 GNDA.n1259 GNDA.n1258 76.3222
R2006 GNDA.n1260 GNDA.n1246 76.3222
R2007 GNDA.n1275 GNDA.n1274 76.3222
R2008 GNDA.n1277 GNDA.n1276 76.3222
R2009 GNDA.n617 GNDA.n436 76.3222
R2010 GNDA.n590 GNDA.n439 76.3222
R2011 GNDA.n598 GNDA.n597 76.3222
R2012 GNDA.n588 GNDA.n585 76.3222
R2013 GNDA.n608 GNDA.n607 76.3222
R2014 GNDA.n583 GNDA.n582 76.3222
R2015 GNDA.n743 GNDA.n742 76.3222
R2016 GNDA.n734 GNDA.n733 76.3222
R2017 GNDA.n721 GNDA.n631 76.3222
R2018 GNDA.n719 GNDA.n718 76.3222
R2019 GNDA.n707 GNDA.n635 76.3222
R2020 GNDA.n706 GNDA.n705 76.3222
R2021 GNDA.n933 GNDA.n932 76.3222
R2022 GNDA.n848 GNDA.n847 76.3222
R2023 GNDA.n863 GNDA.n862 76.3222
R2024 GNDA.n845 GNDA.n841 76.3222
R2025 GNDA.n874 GNDA.n873 76.3222
R2026 GNDA.n839 GNDA.n838 76.3222
R2027 GNDA.n1514 GNDA.n47 76.3222
R2028 GNDA.n1518 GNDA.n46 76.3222
R2029 GNDA.n1522 GNDA.n45 76.3222
R2030 GNDA.n1526 GNDA.n44 76.3222
R2031 GNDA.n1530 GNDA.n43 76.3222
R2032 GNDA.n1533 GNDA.n42 76.3222
R2033 GNDA.n1962 GNDA.n41 76.3222
R2034 GNDA.n1966 GNDA.n40 76.3222
R2035 GNDA.n1970 GNDA.n39 76.3222
R2036 GNDA.n1974 GNDA.n38 76.3222
R2037 GNDA.n1978 GNDA.n37 76.3222
R2038 GNDA.n1982 GNDA.n36 76.3222
R2039 GNDA.n2009 GNDA.n30 76.3222
R2040 GNDA.n103 GNDA.n35 76.3222
R2041 GNDA.n107 GNDA.n34 76.3222
R2042 GNDA.n111 GNDA.n33 76.3222
R2043 GNDA.n115 GNDA.n32 76.3222
R2044 GNDA.n119 GNDA.n31 76.3222
R2045 GNDA.n1278 GNDA.n1277 76.3222
R2046 GNDA.n1274 GNDA.n1273 76.3222
R2047 GNDA.n1261 GNDA.n1260 76.3222
R2048 GNDA.n1258 GNDA.n1257 76.3222
R2049 GNDA.n1248 GNDA.n1220 76.3222
R2050 GNDA.n1338 GNDA.n1337 76.3222
R2051 GNDA.n487 GNDA.n486 76.3222
R2052 GNDA.n484 GNDA.n482 76.3222
R2053 GNDA.n494 GNDA.n493 76.3222
R2054 GNDA.n481 GNDA.n479 76.3222
R2055 GNDA.n501 GNDA.n500 76.3222
R2056 GNDA.n504 GNDA.n503 76.3222
R2057 GNDA.n796 GNDA.n795 76.3222
R2058 GNDA.n791 GNDA.n772 76.3222
R2059 GNDA.n789 GNDA.n788 76.3222
R2060 GNDA.n784 GNDA.n783 76.3222
R2061 GNDA.n781 GNDA.n780 76.3222
R2062 GNDA.n776 GNDA.n424 76.3222
R2063 GNDA.n809 GNDA.n807 76.3222
R2064 GNDA.n966 GNDA.n965 76.3222
R2065 GNDA.n806 GNDA.n804 76.3222
R2066 GNDA.n973 GNDA.n972 76.3222
R2067 GNDA.n803 GNDA.n801 76.3222
R2068 GNDA.n980 GNDA.n979 76.3222
R2069 GNDA.n1440 GNDA.n1439 76.3222
R2070 GNDA.n1443 GNDA.n1442 76.3222
R2071 GNDA.n1452 GNDA.n1451 76.3222
R2072 GNDA.n1455 GNDA.n1454 76.3222
R2073 GNDA.n1467 GNDA.n1466 76.3222
R2074 GNDA.n1470 GNDA.n1469 76.3222
R2075 GNDA.n276 GNDA.n275 76.3222
R2076 GNDA.n309 GNDA.n308 76.3222
R2077 GNDA.n300 GNDA.n281 76.3222
R2078 GNDA.n298 GNDA.n297 76.3222
R2079 GNDA.n283 GNDA.n251 76.3222
R2080 GNDA.n370 GNDA.n369 76.3222
R2081 GNDA.n376 GNDA.n375 76.3222
R2082 GNDA.n379 GNDA.n378 76.3222
R2083 GNDA.n384 GNDA.n383 76.3222
R2084 GNDA.n387 GNDA.n386 76.3222
R2085 GNDA.n392 GNDA.n391 76.3222
R2086 GNDA.n393 GNDA.n392 76.3222
R2087 GNDA.n386 GNDA.n245 76.3222
R2088 GNDA.n385 GNDA.n384 76.3222
R2089 GNDA.n378 GNDA.n247 76.3222
R2090 GNDA.n377 GNDA.n376 76.3222
R2091 GNDA.n369 GNDA.n368 76.3222
R2092 GNDA.n284 GNDA.n283 76.3222
R2093 GNDA.n299 GNDA.n298 76.3222
R2094 GNDA.n281 GNDA.n277 76.3222
R2095 GNDA.n310 GNDA.n309 76.3222
R2096 GNDA.n275 GNDA.n274 76.3222
R2097 GNDA.n1108 GNDA.n1107 76.3222
R2098 GNDA.n1105 GNDA.n1104 76.3222
R2099 GNDA.n1092 GNDA.n1091 76.3222
R2100 GNDA.n1089 GNDA.n1088 76.3222
R2101 GNDA.n1079 GNDA.n1051 76.3222
R2102 GNDA.n1168 GNDA.n1167 76.3222
R2103 GNDA.n1461 GNDA.n1460 76.3222
R2104 GNDA.n1464 GNDA.n1463 76.3222
R2105 GNDA.n1458 GNDA.n1457 76.3222
R2106 GNDA.n1449 GNDA.n1448 76.3222
R2107 GNDA.n1446 GNDA.n1445 76.3222
R2108 GNDA.n1437 GNDA.n1436 76.3222
R2109 GNDA.n1441 GNDA.n1440 76.3222
R2110 GNDA.n1442 GNDA.n226 76.3222
R2111 GNDA.n1453 GNDA.n1452 76.3222
R2112 GNDA.n1454 GNDA.n222 76.3222
R2113 GNDA.n1468 GNDA.n1467 76.3222
R2114 GNDA.n1471 GNDA.n1470 76.3222
R2115 GNDA.n769 GNDA.n768 76.3222
R2116 GNDA.n766 GNDA.n765 76.3222
R2117 GNDA.n761 GNDA.n760 76.3222
R2118 GNDA.n758 GNDA.n757 76.3222
R2119 GNDA.n753 GNDA.n752 76.3222
R2120 GNDA.n750 GNDA.n747 76.3222
R2121 GNDA.n1002 GNDA.n1001 76.3222
R2122 GNDA.n997 GNDA.n749 76.3222
R2123 GNDA.n995 GNDA.n994 76.3222
R2124 GNDA.n990 GNDA.n989 76.3222
R2125 GNDA.n987 GNDA.n986 76.3222
R2126 GNDA.n982 GNDA.n981 76.3222
R2127 GNDA.n1946 GNDA.n97 76.3222
R2128 GNDA.n1949 GNDA.n1948 76.3222
R2129 GNDA.n1944 GNDA.n1943 76.3222
R2130 GNDA.n1935 GNDA.n1934 76.3222
R2131 GNDA.n1932 GNDA.n1931 76.3222
R2132 GNDA.n1923 GNDA.n1922 76.3222
R2133 GNDA.n1927 GNDA.n1926 76.3222
R2134 GNDA.n1928 GNDA.n125 76.3222
R2135 GNDA.n1939 GNDA.n1938 76.3222
R2136 GNDA.n1940 GNDA.n121 76.3222
R2137 GNDA.n1953 GNDA.n1952 76.3222
R2138 GNDA.n1956 GNDA.n1955 76.3222
R2139 GNDA.n93 GNDA.n92 76.3222
R2140 GNDA.n90 GNDA.n89 76.3222
R2141 GNDA.n87 GNDA.n86 76.3222
R2142 GNDA.n84 GNDA.n83 76.3222
R2143 GNDA.n81 GNDA.n80 76.3222
R2144 GNDA.n78 GNDA.n77 76.3222
R2145 GNDA.n2006 GNDA.n74 76.3222
R2146 GNDA.n1999 GNDA.n73 76.3222
R2147 GNDA.n1995 GNDA.n72 76.3222
R2148 GNDA.n1991 GNDA.n71 76.3222
R2149 GNDA.n1987 GNDA.n70 76.3222
R2150 GNDA.n1983 GNDA.n69 76.3222
R2151 GNDA.n1036 GNDA.n1035 76.3222
R2152 GNDA.n1039 GNDA.n1038 76.3222
R2153 GNDA.n1033 GNDA.n1032 76.3222
R2154 GNDA.n1024 GNDA.n1023 76.3222
R2155 GNDA.n1021 GNDA.n1020 76.3222
R2156 GNDA.n1012 GNDA.n1011 76.3222
R2157 GNDA.n1016 GNDA.n1015 76.3222
R2158 GNDA.n1017 GNDA.n430 76.3222
R2159 GNDA.n1028 GNDA.n1027 76.3222
R2160 GNDA.n1029 GNDA.n426 76.3222
R2161 GNDA.n1043 GNDA.n1042 76.3222
R2162 GNDA.n1046 GNDA.n1045 76.3222
R2163 GNDA.n1199 GNDA.n1183 76.3222
R2164 GNDA.n1198 GNDA.n1197 76.3222
R2165 GNDA.n1196 GNDA.n1178 76.3222
R2166 GNDA.n1195 GNDA.n1194 76.3222
R2167 GNDA.n1193 GNDA.n1173 76.3222
R2168 GNDA.n1192 GNDA.n1170 76.3222
R2169 GNDA.n1428 GNDA.n1427 76.3222
R2170 GNDA.n1423 GNDA.n1172 76.3222
R2171 GNDA.n1421 GNDA.n1420 76.3222
R2172 GNDA.n1416 GNDA.n1415 76.3222
R2173 GNDA.n1413 GNDA.n1412 76.3222
R2174 GNDA.n1408 GNDA.n1407 76.3222
R2175 GNDA.n1660 GNDA.n1570 76.062
R2176 GNDA.n1658 GNDA.n1570 76.062
R2177 GNDA.n1130 GNDA.n1063 76.062
R2178 GNDA.n1128 GNDA.n1063 76.062
R2179 GNDA.n668 GNDA.n667 76.062
R2180 GNDA.n667 GNDA.n666 76.062
R2181 GNDA.n1872 GNDA.n160 76.062
R2182 GNDA.n1870 GNDA.n160 76.062
R2183 GNDA.n912 GNDA.n911 76.062
R2184 GNDA.n911 GNDA.n824 76.062
R2185 GNDA.n546 GNDA.n450 76.062
R2186 GNDA.n544 GNDA.n450 76.062
R2187 GNDA.n1300 GNDA.n1233 76.062
R2188 GNDA.n1298 GNDA.n1233 76.062
R2189 GNDA.n348 GNDA.n347 76.062
R2190 GNDA.n347 GNDA.n259 76.062
R2191 GNDA.n1767 GNDA.n1766 76.062
R2192 GNDA.n1766 GNDA.n1765 76.062
R2193 GNDA.n1678 GNDA.n1575 74.5978
R2194 GNDA.n1675 GNDA.n1575 74.5978
R2195 GNDA.n1148 GNDA.n1068 74.5978
R2196 GNDA.n1145 GNDA.n1068 74.5978
R2197 GNDA.n683 GNDA.n641 74.5978
R2198 GNDA.n684 GNDA.n683 74.5978
R2199 GNDA.n1890 GNDA.n165 74.5978
R2200 GNDA.n1887 GNDA.n165 74.5978
R2201 GNDA.n895 GNDA.n894 74.5978
R2202 GNDA.n894 GNDA.n829 74.5978
R2203 GNDA.n564 GNDA.n456 74.5978
R2204 GNDA.n561 GNDA.n456 74.5978
R2205 GNDA.n1318 GNDA.n1238 74.5978
R2206 GNDA.n1315 GNDA.n1238 74.5978
R2207 GNDA.n331 GNDA.n330 74.5978
R2208 GNDA.n330 GNDA.n264 74.5978
R2209 GNDA.n1782 GNDA.n1738 74.5978
R2210 GNDA.n1783 GNDA.n1782 74.5978
R2211 GNDA.n1804 GNDA.t44 74.1404
R2212 GNDA.n2054 GNDA.t62 70.0216
R2213 GNDA.t92 GNDA.n1574 65.8183
R2214 GNDA.t92 GNDA.n1573 65.8183
R2215 GNDA.t92 GNDA.n1572 65.8183
R2216 GNDA.t92 GNDA.n1571 65.8183
R2217 GNDA.t92 GNDA.n1567 65.8183
R2218 GNDA.t92 GNDA.n1565 65.8183
R2219 GNDA.t92 GNDA.n1563 65.8183
R2220 GNDA.t92 GNDA.n1692 65.8183
R2221 GNDA.t92 GNDA.n1578 65.8183
R2222 GNDA.t92 GNDA.n1577 65.8183
R2223 GNDA.t92 GNDA.n1576 65.8183
R2224 GNDA.t80 GNDA.n1067 65.8183
R2225 GNDA.t80 GNDA.n1066 65.8183
R2226 GNDA.t80 GNDA.n1065 65.8183
R2227 GNDA.t80 GNDA.n1064 65.8183
R2228 GNDA.t80 GNDA.n1060 65.8183
R2229 GNDA.t80 GNDA.n1058 65.8183
R2230 GNDA.t80 GNDA.n1056 65.8183
R2231 GNDA.t80 GNDA.n1162 65.8183
R2232 GNDA.t80 GNDA.n1071 65.8183
R2233 GNDA.t80 GNDA.n1070 65.8183
R2234 GNDA.t80 GNDA.n1069 65.8183
R2235 GNDA.n647 GNDA.t76 65.8183
R2236 GNDA.n660 GNDA.t76 65.8183
R2237 GNDA.n654 GNDA.t76 65.8183
R2238 GNDA.n652 GNDA.t76 65.8183
R2239 GNDA.n673 GNDA.t76 65.8183
R2240 GNDA.n675 GNDA.t76 65.8183
R2241 GNDA.n681 GNDA.t76 65.8183
R2242 GNDA.n699 GNDA.t76 65.8183
R2243 GNDA.n697 GNDA.t76 65.8183
R2244 GNDA.n691 GNDA.t76 65.8183
R2245 GNDA.n689 GNDA.t76 65.8183
R2246 GNDA.n738 GNDA.t76 65.8183
R2247 GNDA.n728 GNDA.t76 65.8183
R2248 GNDA.n726 GNDA.t76 65.8183
R2249 GNDA.n712 GNDA.t76 65.8183
R2250 GNDA.t79 GNDA.n164 65.8183
R2251 GNDA.t79 GNDA.n163 65.8183
R2252 GNDA.t79 GNDA.n162 65.8183
R2253 GNDA.t79 GNDA.n161 65.8183
R2254 GNDA.t79 GNDA.n157 65.8183
R2255 GNDA.t79 GNDA.n155 65.8183
R2256 GNDA.t79 GNDA.n153 65.8183
R2257 GNDA.t79 GNDA.n1904 65.8183
R2258 GNDA.t79 GNDA.n168 65.8183
R2259 GNDA.t79 GNDA.n167 65.8183
R2260 GNDA.t79 GNDA.n166 65.8183
R2261 GNDA.t79 GNDA.n158 65.8183
R2262 GNDA.t79 GNDA.n156 65.8183
R2263 GNDA.t79 GNDA.n154 65.8183
R2264 GNDA.t79 GNDA.n152 65.8183
R2265 GNDA.n917 GNDA.t85 65.8183
R2266 GNDA.n823 GNDA.t85 65.8183
R2267 GNDA.n924 GNDA.t85 65.8183
R2268 GNDA.n927 GNDA.t85 65.8183
R2269 GNDA.n908 GNDA.t85 65.8183
R2270 GNDA.n902 GNDA.t85 65.8183
R2271 GNDA.n900 GNDA.t85 65.8183
R2272 GNDA.n878 GNDA.t85 65.8183
R2273 GNDA.n884 GNDA.t85 65.8183
R2274 GNDA.n886 GNDA.t85 65.8183
R2275 GNDA.n892 GNDA.t85 65.8183
R2276 GNDA.n850 GNDA.t85 65.8183
R2277 GNDA.n857 GNDA.t85 65.8183
R2278 GNDA.n843 GNDA.t85 65.8183
R2279 GNDA.n868 GNDA.t85 65.8183
R2280 GNDA.t91 GNDA.n455 65.8183
R2281 GNDA.t91 GNDA.n454 65.8183
R2282 GNDA.t91 GNDA.n453 65.8183
R2283 GNDA.t91 GNDA.n452 65.8183
R2284 GNDA.t91 GNDA.n448 65.8183
R2285 GNDA.t91 GNDA.n446 65.8183
R2286 GNDA.t91 GNDA.n444 65.8183
R2287 GNDA.t91 GNDA.n460 65.8183
R2288 GNDA.t91 GNDA.n459 65.8183
R2289 GNDA.t91 GNDA.n458 65.8183
R2290 GNDA.t91 GNDA.n457 65.8183
R2291 GNDA.n612 GNDA.t91 65.8183
R2292 GNDA.t91 GNDA.n447 65.8183
R2293 GNDA.t91 GNDA.n445 65.8183
R2294 GNDA.t91 GNDA.n443 65.8183
R2295 GNDA.t90 GNDA.n1237 65.8183
R2296 GNDA.t90 GNDA.n1236 65.8183
R2297 GNDA.t90 GNDA.n1235 65.8183
R2298 GNDA.t90 GNDA.n1234 65.8183
R2299 GNDA.t90 GNDA.n1230 65.8183
R2300 GNDA.t90 GNDA.n1228 65.8183
R2301 GNDA.t90 GNDA.n1226 65.8183
R2302 GNDA.t90 GNDA.n1332 65.8183
R2303 GNDA.t90 GNDA.n1241 65.8183
R2304 GNDA.t90 GNDA.n1240 65.8183
R2305 GNDA.t90 GNDA.n1239 65.8183
R2306 GNDA.t90 GNDA.n1231 65.8183
R2307 GNDA.t90 GNDA.n1229 65.8183
R2308 GNDA.t90 GNDA.n1227 65.8183
R2309 GNDA.t90 GNDA.n1225 65.8183
R2310 GNDA.n353 GNDA.t86 65.8183
R2311 GNDA.n258 GNDA.t86 65.8183
R2312 GNDA.n360 GNDA.t86 65.8183
R2313 GNDA.n363 GNDA.t86 65.8183
R2314 GNDA.n344 GNDA.t86 65.8183
R2315 GNDA.n338 GNDA.t86 65.8183
R2316 GNDA.n336 GNDA.t86 65.8183
R2317 GNDA.n314 GNDA.t86 65.8183
R2318 GNDA.n320 GNDA.t86 65.8183
R2319 GNDA.n322 GNDA.t86 65.8183
R2320 GNDA.n328 GNDA.t86 65.8183
R2321 GNDA.n286 GNDA.t86 65.8183
R2322 GNDA.n293 GNDA.t86 65.8183
R2323 GNDA.n279 GNDA.t86 65.8183
R2324 GNDA.n304 GNDA.t86 65.8183
R2325 GNDA.t80 GNDA.n1061 65.8183
R2326 GNDA.t80 GNDA.n1059 65.8183
R2327 GNDA.t80 GNDA.n1057 65.8183
R2328 GNDA.t80 GNDA.n1055 65.8183
R2329 GNDA.n1744 GNDA.t78 65.8183
R2330 GNDA.n1759 GNDA.t78 65.8183
R2331 GNDA.n1753 GNDA.t78 65.8183
R2332 GNDA.n1751 GNDA.t78 65.8183
R2333 GNDA.n1772 GNDA.t78 65.8183
R2334 GNDA.n1774 GNDA.t78 65.8183
R2335 GNDA.n1780 GNDA.t78 65.8183
R2336 GNDA.n1734 GNDA.t78 65.8183
R2337 GNDA.n1796 GNDA.t78 65.8183
R2338 GNDA.n1790 GNDA.t78 65.8183
R2339 GNDA.n1788 GNDA.t78 65.8183
R2340 GNDA.n2049 GNDA.t78 65.8183
R2341 GNDA.n2046 GNDA.t78 65.8183
R2342 GNDA.n2043 GNDA.t78 65.8183
R2343 GNDA.n1802 GNDA.t78 65.8183
R2344 GNDA.t92 GNDA.n1568 65.8183
R2345 GNDA.t92 GNDA.n1566 65.8183
R2346 GNDA.t92 GNDA.n1564 65.8183
R2347 GNDA.t92 GNDA.n1562 65.8183
R2348 GNDA.t15 GNDA.t34 64.1794
R2349 GNDA.t34 GNDA.t11 64.1794
R2350 GNDA.t5 GNDA.t0 64.1794
R2351 GNDA.t36 GNDA.n1619 63.8432
R2352 GNDA.t52 GNDA.n2055 63.8432
R2353 GNDA.n1847 GNDA.t38 63.8432
R2354 GNDA.n1555 GNDA.n16 61.6297
R2355 GNDA.n1 GNDA.t77 32.9056
R2356 GNDA.n0 GNDA.t77 32.9056
R2357 GNDA.t68 GNDA.n1589 59.7243
R2358 GNDA.n1806 GNDA.t54 59.7243
R2359 GNDA.t72 GNDA.n190 59.7243
R2360 GNDA.n180 GNDA.t2 58.6946
R2361 GNDA.t27 GNDA.n1831 58.6946
R2362 GNDA.t111 GNDA.n1848 58.6946
R2363 GNDA.n2034 GNDA.t0 58.2964
R2364 GNDA.n372 GNDA.n371 57.1945
R2365 GNDA.n371 GNDA.n249 57.1945
R2366 GNDA.n937 GNDA.n935 57.1945
R2367 GNDA.n2032 GNDA.n2031 57.1945
R2368 GNDA.t107 GNDA.t70 56.6352
R2369 GNDA.n1818 GNDA.t100 56.6352
R2370 GNDA.t58 GNDA.t31 56.6352
R2371 GNDA.n1912 GNDA.n146 55.6055
R2372 GNDA.t92 GNDA.n1575 55.2026
R2373 GNDA.t80 GNDA.n1068 55.2026
R2374 GNDA.n683 GNDA.t76 55.2026
R2375 GNDA.t79 GNDA.n165 55.2026
R2376 GNDA.n894 GNDA.t85 55.2026
R2377 GNDA.t91 GNDA.n456 55.2026
R2378 GNDA.t90 GNDA.n1238 55.2026
R2379 GNDA.n330 GNDA.t86 55.2026
R2380 GNDA.n1782 GNDA.t78 55.2026
R2381 GNDA.n1699 GNDA.t23 54.5757
R2382 GNDA.t22 GNDA.n1600 54.5757
R2383 GNDA.t4 GNDA.n1634 54.5757
R2384 GNDA.n1723 GNDA.n1722 54.5757
R2385 GNDA.n1816 GNDA.n1728 54.5757
R2386 GNDA.t92 GNDA.n1570 54.4705
R2387 GNDA.t80 GNDA.n1063 54.4705
R2388 GNDA.n667 GNDA.t76 54.4705
R2389 GNDA.t79 GNDA.n160 54.4705
R2390 GNDA.n911 GNDA.t85 54.4705
R2391 GNDA.t91 GNDA.n450 54.4705
R2392 GNDA.t90 GNDA.n1233 54.4705
R2393 GNDA.n347 GNDA.t86 54.4705
R2394 GNDA.n1766 GNDA.t78 54.4705
R2395 GNDA.n1806 GNDA.t66 53.546
R2396 GNDA.n1562 GNDA.n1561 53.3664
R2397 GNDA.n1596 GNDA.n1564 53.3664
R2398 GNDA.n1625 GNDA.n1566 53.3664
R2399 GNDA.n1630 GNDA.n1568 53.3664
R2400 GNDA.n1692 GNDA.n1560 53.3664
R2401 GNDA.n1579 GNDA.n1578 53.3664
R2402 GNDA.n1686 GNDA.n1577 53.3664
R2403 GNDA.n1682 GNDA.n1576 53.3664
R2404 GNDA.n1674 GNDA.n1563 53.3664
R2405 GNDA.n1670 GNDA.n1565 53.3664
R2406 GNDA.n1666 GNDA.n1567 53.3664
R2407 GNDA.n1645 GNDA.n1571 53.3664
R2408 GNDA.n1649 GNDA.n1572 53.3664
R2409 GNDA.n1653 GNDA.n1573 53.3664
R2410 GNDA.n1657 GNDA.n1574 53.3664
R2411 GNDA.n1654 GNDA.n1574 53.3664
R2412 GNDA.n1650 GNDA.n1573 53.3664
R2413 GNDA.n1646 GNDA.n1572 53.3664
R2414 GNDA.n1642 GNDA.n1571 53.3664
R2415 GNDA.n1663 GNDA.n1567 53.3664
R2416 GNDA.n1667 GNDA.n1565 53.3664
R2417 GNDA.n1671 GNDA.n1563 53.3664
R2418 GNDA.n1692 GNDA.n1691 53.3664
R2419 GNDA.n1687 GNDA.n1578 53.3664
R2420 GNDA.n1683 GNDA.n1577 53.3664
R2421 GNDA.n1679 GNDA.n1576 53.3664
R2422 GNDA.n1055 GNDA.n1054 53.3664
R2423 GNDA.n1085 GNDA.n1057 53.3664
R2424 GNDA.n1096 GNDA.n1059 53.3664
R2425 GNDA.n1101 GNDA.n1061 53.3664
R2426 GNDA.n1162 GNDA.n1053 53.3664
R2427 GNDA.n1072 GNDA.n1071 53.3664
R2428 GNDA.n1156 GNDA.n1070 53.3664
R2429 GNDA.n1152 GNDA.n1069 53.3664
R2430 GNDA.n1144 GNDA.n1056 53.3664
R2431 GNDA.n1140 GNDA.n1058 53.3664
R2432 GNDA.n1136 GNDA.n1060 53.3664
R2433 GNDA.n1115 GNDA.n1064 53.3664
R2434 GNDA.n1119 GNDA.n1065 53.3664
R2435 GNDA.n1123 GNDA.n1066 53.3664
R2436 GNDA.n1127 GNDA.n1067 53.3664
R2437 GNDA.n1124 GNDA.n1067 53.3664
R2438 GNDA.n1120 GNDA.n1066 53.3664
R2439 GNDA.n1116 GNDA.n1065 53.3664
R2440 GNDA.n1112 GNDA.n1064 53.3664
R2441 GNDA.n1133 GNDA.n1060 53.3664
R2442 GNDA.n1137 GNDA.n1058 53.3664
R2443 GNDA.n1141 GNDA.n1056 53.3664
R2444 GNDA.n1162 GNDA.n1161 53.3664
R2445 GNDA.n1157 GNDA.n1071 53.3664
R2446 GNDA.n1153 GNDA.n1070 53.3664
R2447 GNDA.n1149 GNDA.n1069 53.3664
R2448 GNDA.n713 GNDA.n712 53.3664
R2449 GNDA.n726 GNDA.n725 53.3664
R2450 GNDA.n729 GNDA.n728 53.3664
R2451 GNDA.n738 GNDA.n737 53.3664
R2452 GNDA.n699 GNDA.n637 53.3664
R2453 GNDA.n698 GNDA.n697 53.3664
R2454 GNDA.n691 GNDA.n639 53.3664
R2455 GNDA.n690 GNDA.n689 53.3664
R2456 GNDA.n682 GNDA.n681 53.3664
R2457 GNDA.n675 GNDA.n643 53.3664
R2458 GNDA.n674 GNDA.n673 53.3664
R2459 GNDA.n653 GNDA.n652 53.3664
R2460 GNDA.n654 GNDA.n649 53.3664
R2461 GNDA.n661 GNDA.n660 53.3664
R2462 GNDA.n665 GNDA.n647 53.3664
R2463 GNDA.n662 GNDA.n647 53.3664
R2464 GNDA.n660 GNDA.n659 53.3664
R2465 GNDA.n655 GNDA.n654 53.3664
R2466 GNDA.n652 GNDA.n628 53.3664
R2467 GNDA.n673 GNDA.n672 53.3664
R2468 GNDA.n676 GNDA.n675 53.3664
R2469 GNDA.n681 GNDA.n680 53.3664
R2470 GNDA.n700 GNDA.n699 53.3664
R2471 GNDA.n697 GNDA.n696 53.3664
R2472 GNDA.n692 GNDA.n691 53.3664
R2473 GNDA.n689 GNDA.n688 53.3664
R2474 GNDA.n739 GNDA.n738 53.3664
R2475 GNDA.n728 GNDA.n629 53.3664
R2476 GNDA.n727 GNDA.n726 53.3664
R2477 GNDA.n712 GNDA.n633 53.3664
R2478 GNDA.n152 GNDA.n151 53.3664
R2479 GNDA.n186 GNDA.n154 53.3664
R2480 GNDA.n1837 GNDA.n156 53.3664
R2481 GNDA.n1842 GNDA.n158 53.3664
R2482 GNDA.n1904 GNDA.n150 53.3664
R2483 GNDA.n169 GNDA.n168 53.3664
R2484 GNDA.n1898 GNDA.n167 53.3664
R2485 GNDA.n1894 GNDA.n166 53.3664
R2486 GNDA.n1886 GNDA.n153 53.3664
R2487 GNDA.n1882 GNDA.n155 53.3664
R2488 GNDA.n1878 GNDA.n157 53.3664
R2489 GNDA.n1857 GNDA.n161 53.3664
R2490 GNDA.n1861 GNDA.n162 53.3664
R2491 GNDA.n1865 GNDA.n163 53.3664
R2492 GNDA.n1869 GNDA.n164 53.3664
R2493 GNDA.n1866 GNDA.n164 53.3664
R2494 GNDA.n1862 GNDA.n163 53.3664
R2495 GNDA.n1858 GNDA.n162 53.3664
R2496 GNDA.n1854 GNDA.n161 53.3664
R2497 GNDA.n1875 GNDA.n157 53.3664
R2498 GNDA.n1879 GNDA.n155 53.3664
R2499 GNDA.n1883 GNDA.n153 53.3664
R2500 GNDA.n1904 GNDA.n1903 53.3664
R2501 GNDA.n1899 GNDA.n168 53.3664
R2502 GNDA.n1895 GNDA.n167 53.3664
R2503 GNDA.n1891 GNDA.n166 53.3664
R2504 GNDA.n1853 GNDA.n158 53.3664
R2505 GNDA.n1841 GNDA.n156 53.3664
R2506 GNDA.n1836 GNDA.n154 53.3664
R2507 GNDA.n185 GNDA.n152 53.3664
R2508 GNDA.n868 GNDA.n835 53.3664
R2509 GNDA.n867 GNDA.n843 53.3664
R2510 GNDA.n857 GNDA.n856 53.3664
R2511 GNDA.n853 GNDA.n850 53.3664
R2512 GNDA.n879 GNDA.n878 53.3664
R2513 GNDA.n884 GNDA.n883 53.3664
R2514 GNDA.n887 GNDA.n886 53.3664
R2515 GNDA.n892 GNDA.n891 53.3664
R2516 GNDA.n900 GNDA.n899 53.3664
R2517 GNDA.n903 GNDA.n902 53.3664
R2518 GNDA.n908 GNDA.n907 53.3664
R2519 GNDA.n927 GNDA.n926 53.3664
R2520 GNDA.n924 GNDA.n923 53.3664
R2521 GNDA.n919 GNDA.n823 53.3664
R2522 GNDA.n917 GNDA.n916 53.3664
R2523 GNDA.n918 GNDA.n917 53.3664
R2524 GNDA.n823 GNDA.n821 53.3664
R2525 GNDA.n925 GNDA.n924 53.3664
R2526 GNDA.n928 GNDA.n927 53.3664
R2527 GNDA.n909 GNDA.n908 53.3664
R2528 GNDA.n902 GNDA.n827 53.3664
R2529 GNDA.n901 GNDA.n900 53.3664
R2530 GNDA.n878 GNDA.n833 53.3664
R2531 GNDA.n885 GNDA.n884 53.3664
R2532 GNDA.n886 GNDA.n831 53.3664
R2533 GNDA.n893 GNDA.n892 53.3664
R2534 GNDA.n850 GNDA.n819 53.3664
R2535 GNDA.n858 GNDA.n857 53.3664
R2536 GNDA.n854 GNDA.n843 53.3664
R2537 GNDA.n869 GNDA.n868 53.3664
R2538 GNDA.n462 GNDA.n443 53.3664
R2539 GNDA.n602 GNDA.n445 53.3664
R2540 GNDA.n592 GNDA.n447 53.3664
R2541 GNDA.n613 GNDA.n612 53.3664
R2542 GNDA.n461 GNDA.n460 53.3664
R2543 GNDA.n576 GNDA.n459 53.3664
R2544 GNDA.n572 GNDA.n458 53.3664
R2545 GNDA.n568 GNDA.n457 53.3664
R2546 GNDA.n560 GNDA.n444 53.3664
R2547 GNDA.n556 GNDA.n446 53.3664
R2548 GNDA.n552 GNDA.n448 53.3664
R2549 GNDA.n531 GNDA.n452 53.3664
R2550 GNDA.n535 GNDA.n453 53.3664
R2551 GNDA.n539 GNDA.n454 53.3664
R2552 GNDA.n543 GNDA.n455 53.3664
R2553 GNDA.n540 GNDA.n455 53.3664
R2554 GNDA.n536 GNDA.n454 53.3664
R2555 GNDA.n532 GNDA.n453 53.3664
R2556 GNDA.n452 GNDA.n451 53.3664
R2557 GNDA.n549 GNDA.n448 53.3664
R2558 GNDA.n553 GNDA.n446 53.3664
R2559 GNDA.n557 GNDA.n444 53.3664
R2560 GNDA.n577 GNDA.n460 53.3664
R2561 GNDA.n573 GNDA.n459 53.3664
R2562 GNDA.n569 GNDA.n458 53.3664
R2563 GNDA.n565 GNDA.n457 53.3664
R2564 GNDA.n612 GNDA.n442 53.3664
R2565 GNDA.n447 GNDA.n441 53.3664
R2566 GNDA.n591 GNDA.n445 53.3664
R2567 GNDA.n603 GNDA.n443 53.3664
R2568 GNDA.n1225 GNDA.n1224 53.3664
R2569 GNDA.n1254 GNDA.n1227 53.3664
R2570 GNDA.n1265 GNDA.n1229 53.3664
R2571 GNDA.n1270 GNDA.n1231 53.3664
R2572 GNDA.n1332 GNDA.n1223 53.3664
R2573 GNDA.n1242 GNDA.n1241 53.3664
R2574 GNDA.n1326 GNDA.n1240 53.3664
R2575 GNDA.n1322 GNDA.n1239 53.3664
R2576 GNDA.n1314 GNDA.n1226 53.3664
R2577 GNDA.n1310 GNDA.n1228 53.3664
R2578 GNDA.n1306 GNDA.n1230 53.3664
R2579 GNDA.n1285 GNDA.n1234 53.3664
R2580 GNDA.n1289 GNDA.n1235 53.3664
R2581 GNDA.n1293 GNDA.n1236 53.3664
R2582 GNDA.n1297 GNDA.n1237 53.3664
R2583 GNDA.n1294 GNDA.n1237 53.3664
R2584 GNDA.n1290 GNDA.n1236 53.3664
R2585 GNDA.n1286 GNDA.n1235 53.3664
R2586 GNDA.n1282 GNDA.n1234 53.3664
R2587 GNDA.n1303 GNDA.n1230 53.3664
R2588 GNDA.n1307 GNDA.n1228 53.3664
R2589 GNDA.n1311 GNDA.n1226 53.3664
R2590 GNDA.n1332 GNDA.n1331 53.3664
R2591 GNDA.n1327 GNDA.n1241 53.3664
R2592 GNDA.n1323 GNDA.n1240 53.3664
R2593 GNDA.n1319 GNDA.n1239 53.3664
R2594 GNDA.n1281 GNDA.n1231 53.3664
R2595 GNDA.n1269 GNDA.n1229 53.3664
R2596 GNDA.n1264 GNDA.n1227 53.3664
R2597 GNDA.n1253 GNDA.n1225 53.3664
R2598 GNDA.n304 GNDA.n270 53.3664
R2599 GNDA.n303 GNDA.n279 53.3664
R2600 GNDA.n293 GNDA.n292 53.3664
R2601 GNDA.n289 GNDA.n286 53.3664
R2602 GNDA.n315 GNDA.n314 53.3664
R2603 GNDA.n320 GNDA.n319 53.3664
R2604 GNDA.n323 GNDA.n322 53.3664
R2605 GNDA.n328 GNDA.n327 53.3664
R2606 GNDA.n336 GNDA.n335 53.3664
R2607 GNDA.n339 GNDA.n338 53.3664
R2608 GNDA.n344 GNDA.n343 53.3664
R2609 GNDA.n363 GNDA.n362 53.3664
R2610 GNDA.n360 GNDA.n359 53.3664
R2611 GNDA.n355 GNDA.n258 53.3664
R2612 GNDA.n353 GNDA.n352 53.3664
R2613 GNDA.n354 GNDA.n353 53.3664
R2614 GNDA.n258 GNDA.n256 53.3664
R2615 GNDA.n361 GNDA.n360 53.3664
R2616 GNDA.n364 GNDA.n363 53.3664
R2617 GNDA.n345 GNDA.n344 53.3664
R2618 GNDA.n338 GNDA.n262 53.3664
R2619 GNDA.n337 GNDA.n336 53.3664
R2620 GNDA.n314 GNDA.n268 53.3664
R2621 GNDA.n321 GNDA.n320 53.3664
R2622 GNDA.n322 GNDA.n266 53.3664
R2623 GNDA.n329 GNDA.n328 53.3664
R2624 GNDA.n286 GNDA.n254 53.3664
R2625 GNDA.n294 GNDA.n293 53.3664
R2626 GNDA.n290 GNDA.n279 53.3664
R2627 GNDA.n305 GNDA.n304 53.3664
R2628 GNDA.n1111 GNDA.n1061 53.3664
R2629 GNDA.n1100 GNDA.n1059 53.3664
R2630 GNDA.n1095 GNDA.n1057 53.3664
R2631 GNDA.n1084 GNDA.n1055 53.3664
R2632 GNDA.n1810 GNDA.n1802 53.3664
R2633 GNDA.n2043 GNDA.n2042 53.3664
R2634 GNDA.n2046 GNDA.n2045 53.3664
R2635 GNDA.n2049 GNDA.n2048 53.3664
R2636 GNDA.n1801 GNDA.n1734 53.3664
R2637 GNDA.n1797 GNDA.n1796 53.3664
R2638 GNDA.n1790 GNDA.n1736 53.3664
R2639 GNDA.n1789 GNDA.n1788 53.3664
R2640 GNDA.n1781 GNDA.n1780 53.3664
R2641 GNDA.n1774 GNDA.n1740 53.3664
R2642 GNDA.n1773 GNDA.n1772 53.3664
R2643 GNDA.n1752 GNDA.n1751 53.3664
R2644 GNDA.n1753 GNDA.n1746 53.3664
R2645 GNDA.n1760 GNDA.n1759 53.3664
R2646 GNDA.n1764 GNDA.n1744 53.3664
R2647 GNDA.n1761 GNDA.n1744 53.3664
R2648 GNDA.n1759 GNDA.n1758 53.3664
R2649 GNDA.n1754 GNDA.n1753 53.3664
R2650 GNDA.n1751 GNDA.n10 53.3664
R2651 GNDA.n1772 GNDA.n1771 53.3664
R2652 GNDA.n1775 GNDA.n1774 53.3664
R2653 GNDA.n1780 GNDA.n1779 53.3664
R2654 GNDA.n1798 GNDA.n1734 53.3664
R2655 GNDA.n1796 GNDA.n1795 53.3664
R2656 GNDA.n1791 GNDA.n1790 53.3664
R2657 GNDA.n1788 GNDA.n1787 53.3664
R2658 GNDA.n2050 GNDA.n2049 53.3664
R2659 GNDA.n2047 GNDA.n2046 53.3664
R2660 GNDA.n2044 GNDA.n2043 53.3664
R2661 GNDA.n1802 GNDA.n13 53.3664
R2662 GNDA.n1641 GNDA.n1568 53.3664
R2663 GNDA.n1629 GNDA.n1566 53.3664
R2664 GNDA.n1624 GNDA.n1564 53.3664
R2665 GNDA.n1595 GNDA.n1562 53.3664
R2666 GNDA.n199 GNDA.n68 51.4866
R2667 GNDA.n1919 GNDA.n134 51.4866
R2668 GNDA.n2055 GNDA.t40 49.4271
R2669 GNDA.n1723 GNDA.t21 48.3974
R2670 GNDA.n2008 GNDA.t77 47.6748
R2671 GNDA.t77 GNDA.n62 47.6748
R2672 GNDA.n146 GNDA.t32 47.3677
R2673 GNDA.t77 GNDA.n63 47.0333
R2674 GNDA.t77 GNDA.n56 47.0333
R2675 GNDA.t77 GNDA.n1201 47.0333
R2676 GNDA.t33 GNDA.t88 46.338
R2677 GNDA.t97 GNDA.t19 46.338
R2678 GNDA.n1378 GNDA.t77 46.2335
R2679 GNDA.t77 GNDA.n1485 46.2335
R2680 GNDA.t77 GNDA.n55 46.2335
R2681 GNDA.n1634 GNDA.t60 43.2488
R2682 GNDA.t40 GNDA.n2054 43.2488
R2683 GNDA.n1849 GNDA.t97 43.2488
R2684 GNDA.t77 GNDA.n1377 42.2987
R2685 GNDA.t77 GNDA.n206 42.2987
R2686 GNDA.t77 GNDA.n54 42.2987
R2687 GNDA.t1 GNDA.n2036 42.2191
R2688 GNDA.t21 GNDA.n68 41.1894
R2689 GNDA.t32 GNDA.n134 41.1894
R2690 GNDA.t77 GNDA.n20 40.6472
R2691 GNDA.n1821 GNDA.n1820 39.3903
R2692 GNDA.t88 GNDA.n1588 39.1299
R2693 GNDA.t66 GNDA.n1804 39.1299
R2694 GNDA.n2038 GNDA.n2037 39.1299
R2695 GNDA.n180 GNDA.t46 39.1299
R2696 GNDA.n1588 GNDA.t23 38.1002
R2697 GNDA.n1601 GNDA.t22 38.1002
R2698 GNDA.n1816 GNDA.n1815 38.1002
R2699 GNDA.n1920 GNDA.n1919 38.1002
R2700 GNDA.n1727 GNDA.n199 37.0705
R2701 GNDA.t77 GNDA.t50 36.0408
R2702 GNDA.t74 GNDA.t77 36.0408
R2703 GNDA.n1613 GNDA.n198 35.3278
R2704 GNDA.n1818 GNDA.n1817 33.9813
R2705 GNDA.n1832 GNDA.t27 33.9813
R2706 GNDA.n1849 GNDA.t111 33.9813
R2707 GNDA.n1590 GNDA.t68 32.9516
R2708 GNDA.t54 GNDA.n1805 32.9516
R2709 GNDA.n191 GNDA.t72 32.9516
R2710 GNDA.n1495 GNDA.n1494 32.3063
R2711 GNDA.n1620 GNDA.t36 28.8327
R2712 GNDA.n2056 GNDA.t52 28.8327
R2713 GNDA.t38 GNDA.n1846 28.8327
R2714 GNDA.t26 GNDA.n1911 27.803
R2715 GNDA.n190 GNDA.t3 27.803
R2716 GNDA.n1846 GNDA.t31 27.803
R2717 GNDA.n1661 GNDA.n1659 27.5561
R2718 GNDA.n1131 GNDA.n1129 27.5561
R2719 GNDA.n669 GNDA.n646 27.5561
R2720 GNDA.n1873 GNDA.n1871 27.5561
R2721 GNDA.n914 GNDA.n913 27.5561
R2722 GNDA.n547 GNDA.n545 27.5561
R2723 GNDA.n1301 GNDA.n1299 27.5561
R2724 GNDA.n350 GNDA.n349 27.5561
R2725 GNDA.n1768 GNDA.n1743 27.5561
R2726 GNDA.n1009 GNDA.n1 8.60107
R2727 GNDA.n1434 GNDA.n0 8.60107
R2728 GNDA.n1677 GNDA.n1676 26.6672
R2729 GNDA.n1147 GNDA.n1146 26.6672
R2730 GNDA.n686 GNDA.n685 26.6672
R2731 GNDA.n1889 GNDA.n1888 26.6672
R2732 GNDA.n897 GNDA.n896 26.6672
R2733 GNDA.n563 GNDA.n562 26.6672
R2734 GNDA.n1317 GNDA.n1316 26.6672
R2735 GNDA.n333 GNDA.n332 26.6672
R2736 GNDA.n1785 GNDA.n1784 26.6672
R2737 GNDA.t77 GNDA.t7 25.9496
R2738 GNDA.t112 GNDA.t60 25.7435
R2739 GNDA.t46 GNDA.t3 25.7435
R2740 GNDA.n197 GNDA.n196 25.3679
R2741 GNDA.n1704 GNDA.t69 24.0005
R2742 GNDA.n1704 GNDA.t71 24.0005
R2743 GNDA.n1706 GNDA.t51 24.0005
R2744 GNDA.n1706 GNDA.t37 24.0005
R2745 GNDA.n1708 GNDA.t61 24.0005
R2746 GNDA.n1708 GNDA.t49 24.0005
R2747 GNDA.n1714 GNDA.t45 24.0005
R2748 GNDA.n1714 GNDA.t67 24.0005
R2749 GNDA.n1712 GNDA.t55 24.0005
R2750 GNDA.n1712 GNDA.t43 24.0005
R2751 GNDA.n1710 GNDA.t65 24.0005
R2752 GNDA.n1710 GNDA.t53 24.0005
R2753 GNDA.n135 GNDA.t41 24.0005
R2754 GNDA.n135 GNDA.t63 24.0005
R2755 GNDA.n143 GNDA.t57 24.0005
R2756 GNDA.n143 GNDA.t47 24.0005
R2757 GNDA.n141 GNDA.t73 24.0005
R2758 GNDA.n141 GNDA.t75 24.0005
R2759 GNDA.n139 GNDA.t59 24.0005
R2760 GNDA.n139 GNDA.t39 24.0005
R2761 GNDA.n1590 GNDA.t107 23.6841
R2762 GNDA.n1619 GNDA.t112 23.6841
R2763 GNDA.n1636 GNDA.t35 23.6841
R2764 GNDA.t77 GNDA.t9 22.706
R2765 GNDA.n1635 GNDA.t48 22.6544
R2766 GNDA.n1817 GNDA.t62 22.6544
R2767 GNDA.n1488 GNDA.n1487 21.0192
R2768 GNDA.n1721 GNDA.n1720 20.8233
R2769 GNDA.n1717 GNDA.n1716 20.8233
R2770 GNDA.n1918 GNDA.n1917 20.8233
R2771 GNDA.n1914 GNDA.n1913 20.8233
R2772 GNDA.n138 GNDA.n137 20.8233
R2773 GNDA.n1702 GNDA.n1701 20.8233
R2774 GNDA.n1618 GNDA.t77 20.5949
R2775 GNDA.t25 GNDA.n1618 20.5949
R2776 GNDA.n1722 GNDA.t35 20.5949
R2777 GNDA.n1912 GNDA.t26 20.5949
R2778 GNDA.n1830 GNDA.t108 20.5949
R2779 GNDA.t77 GNDA.n1830 20.5949
R2780 GNDA.t77 GNDA.n52 19.6741
R2781 GNDA.n212 GNDA.n211 18.5605
R2782 GNDA.n1815 GNDA.t44 18.5355
R2783 GNDA.t56 GNDA.n179 18.5355
R2784 GNDA GNDA.n1492 18.1546
R2785 GNDA.n1535 GNDA.n1534 17.455
R2786 GNDA.n506 GNDA.n505 17.455
R2787 GNDA.n1366 GNDA.n1365 17.455
R2788 GNDA.n2012 GNDA.n28 17.0672
R2789 GNDA.n961 GNDA.n808 17.0672
R2790 GNDA.n396 GNDA.n243 17.0672
R2791 GNDA.n799 GNDA.n233 16.7235
R2792 GNDA.n1006 GNDA.n96 16.7235
R2793 GNDA.n622 GNDA.n95 16.7235
R2794 GNDA.n1432 GNDA.n1048 16.7235
R2795 GNDA.n1644 GNDA.n1643 16.0005
R2796 GNDA.n1647 GNDA.n1644 16.0005
R2797 GNDA.n1648 GNDA.n1647 16.0005
R2798 GNDA.n1651 GNDA.n1648 16.0005
R2799 GNDA.n1652 GNDA.n1651 16.0005
R2800 GNDA.n1655 GNDA.n1652 16.0005
R2801 GNDA.n1656 GNDA.n1655 16.0005
R2802 GNDA.n1659 GNDA.n1656 16.0005
R2803 GNDA.n1676 GNDA.n1673 16.0005
R2804 GNDA.n1673 GNDA.n1672 16.0005
R2805 GNDA.n1672 GNDA.n1669 16.0005
R2806 GNDA.n1669 GNDA.n1668 16.0005
R2807 GNDA.n1668 GNDA.n1665 16.0005
R2808 GNDA.n1665 GNDA.n1664 16.0005
R2809 GNDA.n1664 GNDA.n1662 16.0005
R2810 GNDA.n1662 GNDA.n1661 16.0005
R2811 GNDA.n1690 GNDA.n1558 16.0005
R2812 GNDA.n1690 GNDA.n1689 16.0005
R2813 GNDA.n1689 GNDA.n1688 16.0005
R2814 GNDA.n1688 GNDA.n1685 16.0005
R2815 GNDA.n1685 GNDA.n1684 16.0005
R2816 GNDA.n1684 GNDA.n1681 16.0005
R2817 GNDA.n1681 GNDA.n1680 16.0005
R2818 GNDA.n1680 GNDA.n1677 16.0005
R2819 GNDA.n1114 GNDA.n1113 16.0005
R2820 GNDA.n1117 GNDA.n1114 16.0005
R2821 GNDA.n1118 GNDA.n1117 16.0005
R2822 GNDA.n1121 GNDA.n1118 16.0005
R2823 GNDA.n1122 GNDA.n1121 16.0005
R2824 GNDA.n1125 GNDA.n1122 16.0005
R2825 GNDA.n1126 GNDA.n1125 16.0005
R2826 GNDA.n1129 GNDA.n1126 16.0005
R2827 GNDA.n1146 GNDA.n1143 16.0005
R2828 GNDA.n1143 GNDA.n1142 16.0005
R2829 GNDA.n1142 GNDA.n1139 16.0005
R2830 GNDA.n1139 GNDA.n1138 16.0005
R2831 GNDA.n1138 GNDA.n1135 16.0005
R2832 GNDA.n1135 GNDA.n1134 16.0005
R2833 GNDA.n1134 GNDA.n1132 16.0005
R2834 GNDA.n1132 GNDA.n1131 16.0005
R2835 GNDA.n1160 GNDA.n1073 16.0005
R2836 GNDA.n1160 GNDA.n1159 16.0005
R2837 GNDA.n1159 GNDA.n1158 16.0005
R2838 GNDA.n1158 GNDA.n1155 16.0005
R2839 GNDA.n1155 GNDA.n1154 16.0005
R2840 GNDA.n1154 GNDA.n1151 16.0005
R2841 GNDA.n1151 GNDA.n1150 16.0005
R2842 GNDA.n1150 GNDA.n1147 16.0005
R2843 GNDA.n651 GNDA.n650 16.0005
R2844 GNDA.n656 GNDA.n651 16.0005
R2845 GNDA.n657 GNDA.n656 16.0005
R2846 GNDA.n658 GNDA.n657 16.0005
R2847 GNDA.n658 GNDA.n648 16.0005
R2848 GNDA.n663 GNDA.n648 16.0005
R2849 GNDA.n664 GNDA.n663 16.0005
R2850 GNDA.n664 GNDA.n646 16.0005
R2851 GNDA.n685 GNDA.n642 16.0005
R2852 GNDA.n679 GNDA.n642 16.0005
R2853 GNDA.n679 GNDA.n678 16.0005
R2854 GNDA.n678 GNDA.n677 16.0005
R2855 GNDA.n677 GNDA.n644 16.0005
R2856 GNDA.n671 GNDA.n644 16.0005
R2857 GNDA.n671 GNDA.n670 16.0005
R2858 GNDA.n670 GNDA.n669 16.0005
R2859 GNDA.n702 GNDA.n701 16.0005
R2860 GNDA.n701 GNDA.n638 16.0005
R2861 GNDA.n695 GNDA.n638 16.0005
R2862 GNDA.n695 GNDA.n694 16.0005
R2863 GNDA.n694 GNDA.n693 16.0005
R2864 GNDA.n693 GNDA.n640 16.0005
R2865 GNDA.n687 GNDA.n640 16.0005
R2866 GNDA.n687 GNDA.n686 16.0005
R2867 GNDA.n1856 GNDA.n1855 16.0005
R2868 GNDA.n1859 GNDA.n1856 16.0005
R2869 GNDA.n1860 GNDA.n1859 16.0005
R2870 GNDA.n1863 GNDA.n1860 16.0005
R2871 GNDA.n1864 GNDA.n1863 16.0005
R2872 GNDA.n1867 GNDA.n1864 16.0005
R2873 GNDA.n1868 GNDA.n1867 16.0005
R2874 GNDA.n1871 GNDA.n1868 16.0005
R2875 GNDA.n1888 GNDA.n1885 16.0005
R2876 GNDA.n1885 GNDA.n1884 16.0005
R2877 GNDA.n1884 GNDA.n1881 16.0005
R2878 GNDA.n1881 GNDA.n1880 16.0005
R2879 GNDA.n1880 GNDA.n1877 16.0005
R2880 GNDA.n1877 GNDA.n1876 16.0005
R2881 GNDA.n1876 GNDA.n1874 16.0005
R2882 GNDA.n1874 GNDA.n1873 16.0005
R2883 GNDA.n1902 GNDA.n148 16.0005
R2884 GNDA.n1902 GNDA.n1901 16.0005
R2885 GNDA.n1901 GNDA.n1900 16.0005
R2886 GNDA.n1900 GNDA.n1897 16.0005
R2887 GNDA.n1897 GNDA.n1896 16.0005
R2888 GNDA.n1896 GNDA.n1893 16.0005
R2889 GNDA.n1893 GNDA.n1892 16.0005
R2890 GNDA.n1892 GNDA.n1889 16.0005
R2891 GNDA.n929 GNDA.n818 16.0005
R2892 GNDA.n820 GNDA.n818 16.0005
R2893 GNDA.n922 GNDA.n820 16.0005
R2894 GNDA.n922 GNDA.n921 16.0005
R2895 GNDA.n921 GNDA.n920 16.0005
R2896 GNDA.n920 GNDA.n822 16.0005
R2897 GNDA.n915 GNDA.n822 16.0005
R2898 GNDA.n915 GNDA.n914 16.0005
R2899 GNDA.n898 GNDA.n897 16.0005
R2900 GNDA.n898 GNDA.n828 16.0005
R2901 GNDA.n904 GNDA.n828 16.0005
R2902 GNDA.n905 GNDA.n904 16.0005
R2903 GNDA.n906 GNDA.n905 16.0005
R2904 GNDA.n906 GNDA.n826 16.0005
R2905 GNDA.n826 GNDA.n825 16.0005
R2906 GNDA.n913 GNDA.n825 16.0005
R2907 GNDA.n881 GNDA.n880 16.0005
R2908 GNDA.n882 GNDA.n881 16.0005
R2909 GNDA.n882 GNDA.n832 16.0005
R2910 GNDA.n888 GNDA.n832 16.0005
R2911 GNDA.n889 GNDA.n888 16.0005
R2912 GNDA.n890 GNDA.n889 16.0005
R2913 GNDA.n890 GNDA.n830 16.0005
R2914 GNDA.n896 GNDA.n830 16.0005
R2915 GNDA.n530 GNDA.n437 16.0005
R2916 GNDA.n533 GNDA.n530 16.0005
R2917 GNDA.n534 GNDA.n533 16.0005
R2918 GNDA.n537 GNDA.n534 16.0005
R2919 GNDA.n538 GNDA.n537 16.0005
R2920 GNDA.n541 GNDA.n538 16.0005
R2921 GNDA.n542 GNDA.n541 16.0005
R2922 GNDA.n545 GNDA.n542 16.0005
R2923 GNDA.n562 GNDA.n559 16.0005
R2924 GNDA.n559 GNDA.n558 16.0005
R2925 GNDA.n558 GNDA.n555 16.0005
R2926 GNDA.n555 GNDA.n554 16.0005
R2927 GNDA.n554 GNDA.n551 16.0005
R2928 GNDA.n551 GNDA.n550 16.0005
R2929 GNDA.n550 GNDA.n548 16.0005
R2930 GNDA.n548 GNDA.n547 16.0005
R2931 GNDA.n579 GNDA.n578 16.0005
R2932 GNDA.n578 GNDA.n575 16.0005
R2933 GNDA.n575 GNDA.n574 16.0005
R2934 GNDA.n574 GNDA.n571 16.0005
R2935 GNDA.n571 GNDA.n570 16.0005
R2936 GNDA.n570 GNDA.n567 16.0005
R2937 GNDA.n567 GNDA.n566 16.0005
R2938 GNDA.n566 GNDA.n563 16.0005
R2939 GNDA.n1284 GNDA.n1283 16.0005
R2940 GNDA.n1287 GNDA.n1284 16.0005
R2941 GNDA.n1288 GNDA.n1287 16.0005
R2942 GNDA.n1291 GNDA.n1288 16.0005
R2943 GNDA.n1292 GNDA.n1291 16.0005
R2944 GNDA.n1295 GNDA.n1292 16.0005
R2945 GNDA.n1296 GNDA.n1295 16.0005
R2946 GNDA.n1299 GNDA.n1296 16.0005
R2947 GNDA.n1316 GNDA.n1313 16.0005
R2948 GNDA.n1313 GNDA.n1312 16.0005
R2949 GNDA.n1312 GNDA.n1309 16.0005
R2950 GNDA.n1309 GNDA.n1308 16.0005
R2951 GNDA.n1308 GNDA.n1305 16.0005
R2952 GNDA.n1305 GNDA.n1304 16.0005
R2953 GNDA.n1304 GNDA.n1302 16.0005
R2954 GNDA.n1302 GNDA.n1301 16.0005
R2955 GNDA.n1330 GNDA.n1243 16.0005
R2956 GNDA.n1330 GNDA.n1329 16.0005
R2957 GNDA.n1329 GNDA.n1328 16.0005
R2958 GNDA.n1328 GNDA.n1325 16.0005
R2959 GNDA.n1325 GNDA.n1324 16.0005
R2960 GNDA.n1324 GNDA.n1321 16.0005
R2961 GNDA.n1321 GNDA.n1320 16.0005
R2962 GNDA.n1320 GNDA.n1317 16.0005
R2963 GNDA.n365 GNDA.n253 16.0005
R2964 GNDA.n255 GNDA.n253 16.0005
R2965 GNDA.n358 GNDA.n255 16.0005
R2966 GNDA.n358 GNDA.n357 16.0005
R2967 GNDA.n357 GNDA.n356 16.0005
R2968 GNDA.n356 GNDA.n257 16.0005
R2969 GNDA.n351 GNDA.n257 16.0005
R2970 GNDA.n351 GNDA.n350 16.0005
R2971 GNDA.n334 GNDA.n333 16.0005
R2972 GNDA.n334 GNDA.n263 16.0005
R2973 GNDA.n340 GNDA.n263 16.0005
R2974 GNDA.n341 GNDA.n340 16.0005
R2975 GNDA.n342 GNDA.n341 16.0005
R2976 GNDA.n342 GNDA.n261 16.0005
R2977 GNDA.n261 GNDA.n260 16.0005
R2978 GNDA.n349 GNDA.n260 16.0005
R2979 GNDA.n317 GNDA.n316 16.0005
R2980 GNDA.n318 GNDA.n317 16.0005
R2981 GNDA.n318 GNDA.n267 16.0005
R2982 GNDA.n324 GNDA.n267 16.0005
R2983 GNDA.n325 GNDA.n324 16.0005
R2984 GNDA.n326 GNDA.n325 16.0005
R2985 GNDA.n326 GNDA.n265 16.0005
R2986 GNDA.n332 GNDA.n265 16.0005
R2987 GNDA.n1750 GNDA.n1749 16.0005
R2988 GNDA.n1755 GNDA.n1750 16.0005
R2989 GNDA.n1756 GNDA.n1755 16.0005
R2990 GNDA.n1757 GNDA.n1756 16.0005
R2991 GNDA.n1757 GNDA.n1745 16.0005
R2992 GNDA.n1762 GNDA.n1745 16.0005
R2993 GNDA.n1763 GNDA.n1762 16.0005
R2994 GNDA.n1763 GNDA.n1743 16.0005
R2995 GNDA.n1784 GNDA.n1739 16.0005
R2996 GNDA.n1778 GNDA.n1739 16.0005
R2997 GNDA.n1778 GNDA.n1777 16.0005
R2998 GNDA.n1777 GNDA.n1776 16.0005
R2999 GNDA.n1776 GNDA.n1741 16.0005
R3000 GNDA.n1770 GNDA.n1741 16.0005
R3001 GNDA.n1770 GNDA.n1769 16.0005
R3002 GNDA.n1769 GNDA.n1768 16.0005
R3003 GNDA.n1800 GNDA.n1799 16.0005
R3004 GNDA.n1799 GNDA.n1735 16.0005
R3005 GNDA.n1794 GNDA.n1735 16.0005
R3006 GNDA.n1794 GNDA.n1793 16.0005
R3007 GNDA.n1793 GNDA.n1792 16.0005
R3008 GNDA.n1792 GNDA.n1737 16.0005
R3009 GNDA.n1786 GNDA.n1737 16.0005
R3010 GNDA.n1786 GNDA.n1785 16.0005
R3011 GNDA.n211 GNDA.n202 16.0005
R3012 GNDA.n1487 GNDA.n202 16.0005
R3013 GNDA.n1492 GNDA.n1490 15.4932
R3014 GNDA.t48 GNDA.t4 15.4463
R3015 GNDA.t2 GNDA.t56 15.4463
R3016 GNDA.n140 GNDA.n138 14.363
R3017 GNDA.n1720 GNDA.n1719 13.8005
R3018 GNDA.n1718 GNDA.n1717 13.8005
R3019 GNDA.n1917 GNDA.n1916 13.8005
R3020 GNDA.n1915 GNDA.n1914 13.8005
R3021 GNDA.n1703 GNDA.n1702 13.8005
R3022 GNDA.n1493 GNDA.n198 12.7542
R3023 GNDA.n1600 GNDA.t70 12.3572
R3024 GNDA.n2038 GNDA.t42 12.3572
R3025 GNDA.n1832 GNDA.t74 12.3572
R3026 GNDA.n1820 GNDA.n1819 12.2193
R3027 GNDA.n778 GNDA.n420 11.6369
R3028 GNDA.n779 GNDA.n778 11.6369
R3029 GNDA.n779 GNDA.n775 11.6369
R3030 GNDA.n785 GNDA.n775 11.6369
R3031 GNDA.n786 GNDA.n785 11.6369
R3032 GNDA.n787 GNDA.n786 11.6369
R3033 GNDA.n787 GNDA.n773 11.6369
R3034 GNDA.n792 GNDA.n773 11.6369
R3035 GNDA.n793 GNDA.n792 11.6369
R3036 GNDA.n793 GNDA.n771 11.6369
R3037 GNDA.n798 GNDA.n771 11.6369
R3038 GNDA.n1981 GNDA.n1980 11.6369
R3039 GNDA.n1980 GNDA.n1977 11.6369
R3040 GNDA.n1977 GNDA.n1976 11.6369
R3041 GNDA.n1976 GNDA.n1973 11.6369
R3042 GNDA.n1973 GNDA.n1972 11.6369
R3043 GNDA.n1972 GNDA.n1969 11.6369
R3044 GNDA.n1969 GNDA.n1968 11.6369
R3045 GNDA.n1968 GNDA.n1965 11.6369
R3046 GNDA.n1965 GNDA.n1964 11.6369
R3047 GNDA.n1964 GNDA.n1961 11.6369
R3048 GNDA.n1961 GNDA.n1960 11.6369
R3049 GNDA.n118 GNDA.n117 11.6369
R3050 GNDA.n117 GNDA.n114 11.6369
R3051 GNDA.n114 GNDA.n113 11.6369
R3052 GNDA.n113 GNDA.n110 11.6369
R3053 GNDA.n110 GNDA.n109 11.6369
R3054 GNDA.n109 GNDA.n106 11.6369
R3055 GNDA.n106 GNDA.n105 11.6369
R3056 GNDA.n105 GNDA.n102 11.6369
R3057 GNDA.n102 GNDA.n101 11.6369
R3058 GNDA.n101 GNDA.n99 11.6369
R3059 GNDA.n99 GNDA.n28 11.6369
R3060 GNDA.n2028 GNDA.n2027 11.6369
R3061 GNDA.n2027 GNDA.n2026 11.6369
R3062 GNDA.n2026 GNDA.n22 11.6369
R3063 GNDA.n2021 GNDA.n22 11.6369
R3064 GNDA.n2021 GNDA.n2020 11.6369
R3065 GNDA.n2020 GNDA.n2019 11.6369
R3066 GNDA.n2019 GNDA.n25 11.6369
R3067 GNDA.n2014 GNDA.n25 11.6369
R3068 GNDA.n2014 GNDA.n2013 11.6369
R3069 GNDA.n2013 GNDA.n2012 11.6369
R3070 GNDA.n977 GNDA.n800 11.6369
R3071 GNDA.n977 GNDA.n976 11.6369
R3072 GNDA.n976 GNDA.n975 11.6369
R3073 GNDA.n975 GNDA.n802 11.6369
R3074 GNDA.n970 GNDA.n802 11.6369
R3075 GNDA.n970 GNDA.n969 11.6369
R3076 GNDA.n969 GNDA.n968 11.6369
R3077 GNDA.n968 GNDA.n805 11.6369
R3078 GNDA.n963 GNDA.n805 11.6369
R3079 GNDA.n963 GNDA.n962 11.6369
R3080 GNDA.n962 GNDA.n961 11.6369
R3081 GNDA.n940 GNDA.n939 11.6369
R3082 GNDA.n940 GNDA.n813 11.6369
R3083 GNDA.n946 GNDA.n813 11.6369
R3084 GNDA.n947 GNDA.n946 11.6369
R3085 GNDA.n948 GNDA.n947 11.6369
R3086 GNDA.n948 GNDA.n811 11.6369
R3087 GNDA.n954 GNDA.n811 11.6369
R3088 GNDA.n955 GNDA.n954 11.6369
R3089 GNDA.n956 GNDA.n955 11.6369
R3090 GNDA.n956 GNDA.n808 11.6369
R3091 GNDA.n1534 GNDA.n1532 11.6369
R3092 GNDA.n1532 GNDA.n1529 11.6369
R3093 GNDA.n1529 GNDA.n1528 11.6369
R3094 GNDA.n1528 GNDA.n1525 11.6369
R3095 GNDA.n1525 GNDA.n1524 11.6369
R3096 GNDA.n1524 GNDA.n1521 11.6369
R3097 GNDA.n1521 GNDA.n1520 11.6369
R3098 GNDA.n1520 GNDA.n1517 11.6369
R3099 GNDA.n1517 GNDA.n1516 11.6369
R3100 GNDA.n1516 GNDA.n1513 11.6369
R3101 GNDA.n1513 GNDA.n1512 11.6369
R3102 GNDA.n1551 GNDA.n1500 11.6369
R3103 GNDA.n1551 GNDA.n1550 11.6369
R3104 GNDA.n1550 GNDA.n1549 11.6369
R3105 GNDA.n1549 GNDA.n1505 11.6369
R3106 GNDA.n1544 GNDA.n1505 11.6369
R3107 GNDA.n1544 GNDA.n1543 11.6369
R3108 GNDA.n1543 GNDA.n1542 11.6369
R3109 GNDA.n1542 GNDA.n1507 11.6369
R3110 GNDA.n1536 GNDA.n1507 11.6369
R3111 GNDA.n1536 GNDA.n1535 11.6369
R3112 GNDA.n505 GNDA.n477 11.6369
R3113 GNDA.n478 GNDA.n477 11.6369
R3114 GNDA.n498 GNDA.n478 11.6369
R3115 GNDA.n498 GNDA.n497 11.6369
R3116 GNDA.n497 GNDA.n496 11.6369
R3117 GNDA.n496 GNDA.n480 11.6369
R3118 GNDA.n491 GNDA.n480 11.6369
R3119 GNDA.n491 GNDA.n490 11.6369
R3120 GNDA.n490 GNDA.n489 11.6369
R3121 GNDA.n489 GNDA.n483 11.6369
R3122 GNDA.n483 GNDA.n421 11.6369
R3123 GNDA.n522 GNDA.n466 11.6369
R3124 GNDA.n522 GNDA.n521 11.6369
R3125 GNDA.n521 GNDA.n520 11.6369
R3126 GNDA.n520 GNDA.n470 11.6369
R3127 GNDA.n515 GNDA.n470 11.6369
R3128 GNDA.n515 GNDA.n514 11.6369
R3129 GNDA.n514 GNDA.n513 11.6369
R3130 GNDA.n513 GNDA.n472 11.6369
R3131 GNDA.n507 GNDA.n472 11.6369
R3132 GNDA.n507 GNDA.n506 11.6369
R3133 GNDA.n1367 GNDA.n1366 11.6369
R3134 GNDA.n1367 GNDA.n1205 11.6369
R3135 GNDA.n1373 GNDA.n1205 11.6369
R3136 GNDA.n1374 GNDA.n1373 11.6369
R3137 GNDA.n1375 GNDA.n1374 11.6369
R3138 GNDA.n1375 GNDA.n1189 11.6369
R3139 GNDA.n1381 GNDA.n1189 11.6369
R3140 GNDA.n1382 GNDA.n1381 11.6369
R3141 GNDA.n1383 GNDA.n1382 11.6369
R3142 GNDA.n1383 GNDA.n1185 11.6369
R3143 GNDA.n1389 GNDA.n1185 11.6369
R3144 GNDA.n1343 GNDA.n1215 11.6369
R3145 GNDA.n1350 GNDA.n1215 11.6369
R3146 GNDA.n1351 GNDA.n1350 11.6369
R3147 GNDA.n1352 GNDA.n1351 11.6369
R3148 GNDA.n1352 GNDA.n1213 11.6369
R3149 GNDA.n1357 GNDA.n1213 11.6369
R3150 GNDA.n1358 GNDA.n1357 11.6369
R3151 GNDA.n1359 GNDA.n1358 11.6369
R3152 GNDA.n1359 GNDA.n1209 11.6369
R3153 GNDA.n1365 GNDA.n1209 11.6369
R3154 GNDA.n414 GNDA.n217 11.6369
R3155 GNDA.n414 GNDA.n413 11.6369
R3156 GNDA.n413 GNDA.n412 11.6369
R3157 GNDA.n412 GNDA.n237 11.6369
R3158 GNDA.n406 GNDA.n237 11.6369
R3159 GNDA.n406 GNDA.n405 11.6369
R3160 GNDA.n405 GNDA.n404 11.6369
R3161 GNDA.n404 GNDA.n239 11.6369
R3162 GNDA.n398 GNDA.n239 11.6369
R3163 GNDA.n398 GNDA.n397 11.6369
R3164 GNDA.n397 GNDA.n396 11.6369
R3165 GNDA.n374 GNDA.n248 11.6369
R3166 GNDA.n380 GNDA.n248 11.6369
R3167 GNDA.n381 GNDA.n380 11.6369
R3168 GNDA.n382 GNDA.n381 11.6369
R3169 GNDA.n382 GNDA.n246 11.6369
R3170 GNDA.n388 GNDA.n246 11.6369
R3171 GNDA.n389 GNDA.n388 11.6369
R3172 GNDA.n390 GNDA.n389 11.6369
R3173 GNDA.n390 GNDA.n244 11.6369
R3174 GNDA.n244 GNDA.n243 11.6369
R3175 GNDA.n1395 GNDA.n1392 11.6369
R3176 GNDA.n1401 GNDA.n1395 11.6369
R3177 GNDA.n1401 GNDA.n1400 11.6369
R3178 GNDA.n1400 GNDA.n1399 11.6369
R3179 GNDA.n1399 GNDA.n1396 11.6369
R3180 GNDA.n1483 GNDA.n1482 11.6369
R3181 GNDA.n1482 GNDA.n1481 11.6369
R3182 GNDA.n1481 GNDA.n213 11.6369
R3183 GNDA.n1475 GNDA.n213 11.6369
R3184 GNDA.n1475 GNDA.n1474 11.6369
R3185 GNDA.n1703 GNDA.n201 11.3792
R3186 GNDA.t12 GNDA.t9 11.3532
R3187 GNDA.n1612 GNDA.t105 9.6005
R3188 GNDA.n1615 GNDA.t18 9.6005
R3189 GNDA.n195 GNDA.t106 9.6005
R3190 GNDA.n1827 GNDA.t14 9.6005
R3191 GNDA.t50 GNDA.n1601 8.23827
R3192 GNDA.n2036 GNDA.t64 8.23827
R3193 GNDA.n1831 GNDA.t58 8.23827
R3194 GNDA.n1490 GNDA.n1489 7.56675
R3195 GNDA.n1492 GNDA.n1491 7.56675
R3196 GNDA.n1700 GNDA.n1699 7.20855
R3197 GNDA.n1589 GNDA.t33 7.20855
R3198 GNDA.n1620 GNDA.t25 7.20855
R3199 GNDA.n179 GNDA.t110 7.20855
R3200 GNDA.t13 GNDA.n2033 7.20855
R3201 GNDA.n1048 GNDA.n420 6.72373
R3202 GNDA.n1981 GNDA.n95 6.72373
R3203 GNDA.n118 GNDA.n96 6.72373
R3204 GNDA.n800 GNDA.n799 6.72373
R3205 GNDA.n1473 GNDA.n217 6.72373
R3206 GNDA.n1392 GNDA.n1390 6.72373
R3207 GNDA.n799 GNDA.n798 6.20656
R3208 GNDA.n1960 GNDA.n96 6.20656
R3209 GNDA.n1512 GNDA.n95 6.20656
R3210 GNDA.n1048 GNDA.n421 6.20656
R3211 GNDA.n1390 GNDA.n1389 6.20656
R3212 GNDA.n1474 GNDA.n1473 6.20656
R3213 GNDA.n1497 GNDA.t17 6.17883
R3214 GNDA.t77 GNDA.t1 6.17883
R3215 GNDA.n1483 GNDA.n212 6.07727
R3216 GNDA.n2034 GNDA.t20 5.88357
R3217 GNDA.n1828 GNDA.n196 5.81868
R3218 GNDA.n1826 GNDA.n196 5.81868
R3219 GNDA.n1396 GNDA.n212 5.5601
R3220 GNDA.n1696 GNDA.n1558 5.51161
R3221 GNDA.n1073 GNDA.n1050 5.51161
R3222 GNDA.n703 GNDA.n702 5.51161
R3223 GNDA.n1908 GNDA.n148 5.51161
R3224 GNDA.n880 GNDA.n834 5.51161
R3225 GNDA.n580 GNDA.n579 5.51161
R3226 GNDA.n1243 GNDA.n1221 5.51161
R3227 GNDA.n316 GNDA.n269 5.51161
R3228 GNDA.n1800 GNDA.n1732 5.51161
R3229 GNDA.n581 GNDA.n529 5.1717
R3230 GNDA.n1342 GNDA.n1219 5.1717
R3231 GNDA.n1697 GNDA.n1557 5.1717
R3232 GNDA.t83 GNDA.t24 5.14911
R3233 GNDA.n2037 GNDA.t77 5.14911
R3234 GNDA.n170 GNDA.n19 4.9157
R3235 GNDA.n938 GNDA.n815 4.9157
R3236 GNDA.n373 GNDA.n250 4.9157
R3237 GNDA.n1438 GNDA.n229 4.26717
R3238 GNDA.n1444 GNDA.n229 4.26717
R3239 GNDA.n1444 GNDA.n227 4.26717
R3240 GNDA.n1450 GNDA.n227 4.26717
R3241 GNDA.n1450 GNDA.n225 4.26717
R3242 GNDA.n1456 GNDA.n225 4.26717
R3243 GNDA.n1456 GNDA.n223 4.26717
R3244 GNDA.n1465 GNDA.n223 4.26717
R3245 GNDA.n1465 GNDA.n221 4.26717
R3246 GNDA.n221 GNDA.n218 4.26717
R3247 GNDA.n1472 GNDA.n218 4.26717
R3248 GNDA.n1004 GNDA.n748 4.26717
R3249 GNDA.n999 GNDA.n748 4.26717
R3250 GNDA.n999 GNDA.n998 4.26717
R3251 GNDA.n998 GNDA.n755 4.26717
R3252 GNDA.n993 GNDA.n755 4.26717
R3253 GNDA.n993 GNDA.n992 4.26717
R3254 GNDA.n992 GNDA.n991 4.26717
R3255 GNDA.n991 GNDA.n763 4.26717
R3256 GNDA.n985 GNDA.n763 4.26717
R3257 GNDA.n985 GNDA.n984 4.26717
R3258 GNDA.n984 GNDA.n983 4.26717
R3259 GNDA.n1924 GNDA.n128 4.26717
R3260 GNDA.n1930 GNDA.n128 4.26717
R3261 GNDA.n1930 GNDA.n126 4.26717
R3262 GNDA.n1936 GNDA.n126 4.26717
R3263 GNDA.n1936 GNDA.n124 4.26717
R3264 GNDA.n1942 GNDA.n124 4.26717
R3265 GNDA.n1942 GNDA.n122 4.26717
R3266 GNDA.n1950 GNDA.n122 4.26717
R3267 GNDA.n1950 GNDA.n120 4.26717
R3268 GNDA.n120 GNDA.n98 4.26717
R3269 GNDA.n1957 GNDA.n98 4.26717
R3270 GNDA.n2004 GNDA.n2003 4.26717
R3271 GNDA.n2003 GNDA.n2002 4.26717
R3272 GNDA.n2002 GNDA.n2000 4.26717
R3273 GNDA.n2000 GNDA.n1997 4.26717
R3274 GNDA.n1997 GNDA.n1996 4.26717
R3275 GNDA.n1996 GNDA.n1993 4.26717
R3276 GNDA.n1993 GNDA.n1992 4.26717
R3277 GNDA.n1992 GNDA.n1989 4.26717
R3278 GNDA.n1989 GNDA.n1988 4.26717
R3279 GNDA.n1988 GNDA.n1985 4.26717
R3280 GNDA.n1985 GNDA.n1984 4.26717
R3281 GNDA.n1013 GNDA.n433 4.26717
R3282 GNDA.n1019 GNDA.n433 4.26717
R3283 GNDA.n1019 GNDA.n431 4.26717
R3284 GNDA.n1025 GNDA.n431 4.26717
R3285 GNDA.n1025 GNDA.n429 4.26717
R3286 GNDA.n1031 GNDA.n429 4.26717
R3287 GNDA.n1031 GNDA.n427 4.26717
R3288 GNDA.n1040 GNDA.n427 4.26717
R3289 GNDA.n1040 GNDA.n425 4.26717
R3290 GNDA.n425 GNDA.n422 4.26717
R3291 GNDA.n1047 GNDA.n422 4.26717
R3292 GNDA.n1430 GNDA.n1171 4.26717
R3293 GNDA.n1425 GNDA.n1171 4.26717
R3294 GNDA.n1425 GNDA.n1424 4.26717
R3295 GNDA.n1424 GNDA.n1175 4.26717
R3296 GNDA.n1419 GNDA.n1175 4.26717
R3297 GNDA.n1419 GNDA.n1418 4.26717
R3298 GNDA.n1418 GNDA.n1417 4.26717
R3299 GNDA.n1417 GNDA.n1180 4.26717
R3300 GNDA.n1411 GNDA.n1180 4.26717
R3301 GNDA.n1411 GNDA.n1410 4.26717
R3302 GNDA.n1410 GNDA.n1409 4.26717
R3303 GNDA.n1820 GNDA.n198 4.063
R3304 GNDA.n1473 GNDA.n1472 3.98272
R3305 GNDA.n983 GNDA.n799 3.98272
R3306 GNDA.n1957 GNDA.n96 3.98272
R3307 GNDA.n1984 GNDA.n95 3.98272
R3308 GNDA.n1048 GNDA.n1047 3.98272
R3309 GNDA.n1409 GNDA.n1390 3.98272
R3310 GNDA.n710 GNDA.n636 3.7893
R3311 GNDA.n716 GNDA.n714 3.7893
R3312 GNDA.n715 GNDA.n634 3.7893
R3313 GNDA.n724 GNDA.n723 3.7893
R3314 GNDA.n720 GNDA.n632 3.7893
R3315 GNDA.n735 GNDA.n630 3.7893
R3316 GNDA.n736 GNDA.n627 3.7893
R3317 GNDA.n741 GNDA.n740 3.7893
R3318 GNDA.n1906 GNDA.n149 3.7893
R3319 GNDA.n183 GNDA.n182 3.7893
R3320 GNDA.n188 GNDA.n184 3.7893
R3321 GNDA.n187 GNDA.n175 3.7893
R3322 GNDA.n1835 GNDA.n1834 3.7893
R3323 GNDA.n1844 GNDA.n1840 3.7893
R3324 GNDA.n1843 GNDA.n172 3.7893
R3325 GNDA.n1852 GNDA.n1851 3.7893
R3326 GNDA.n876 GNDA.n875 3.7893
R3327 GNDA.n871 GNDA.n837 3.7893
R3328 GNDA.n870 GNDA.n842 3.7893
R3329 GNDA.n866 GNDA.n865 3.7893
R3330 GNDA.n846 GNDA.n844 3.7893
R3331 GNDA.n859 GNDA.n849 3.7893
R3332 GNDA.n852 GNDA.n851 3.7893
R3333 GNDA.n931 GNDA.n817 3.7893
R3334 GNDA.n610 GNDA.n609 3.7893
R3335 GNDA.n605 GNDA.n464 3.7893
R3336 GNDA.n604 GNDA.n586 3.7893
R3337 GNDA.n601 GNDA.n600 3.7893
R3338 GNDA.n589 GNDA.n587 3.7893
R3339 GNDA.n594 GNDA.n440 3.7893
R3340 GNDA.n615 GNDA.n614 3.7893
R3341 GNDA.n618 GNDA.n438 3.7893
R3342 GNDA.n1334 GNDA.n1222 3.7893
R3343 GNDA.n1251 GNDA.n1250 3.7893
R3344 GNDA.n1256 GNDA.n1252 3.7893
R3345 GNDA.n1255 GNDA.n1247 3.7893
R3346 GNDA.n1263 GNDA.n1262 3.7893
R3347 GNDA.n1272 GNDA.n1268 3.7893
R3348 GNDA.n1271 GNDA.n1245 3.7893
R3349 GNDA.n1280 GNDA.n1279 3.7893
R3350 GNDA.n312 GNDA.n311 3.7893
R3351 GNDA.n307 GNDA.n272 3.7893
R3352 GNDA.n306 GNDA.n278 3.7893
R3353 GNDA.n302 GNDA.n301 3.7893
R3354 GNDA.n282 GNDA.n280 3.7893
R3355 GNDA.n295 GNDA.n285 3.7893
R3356 GNDA.n288 GNDA.n287 3.7893
R3357 GNDA.n367 GNDA.n252 3.7893
R3358 GNDA.n1164 GNDA.n1052 3.7893
R3359 GNDA.n1082 GNDA.n1081 3.7893
R3360 GNDA.n1087 GNDA.n1083 3.7893
R3361 GNDA.n1086 GNDA.n1078 3.7893
R3362 GNDA.n1094 GNDA.n1093 3.7893
R3363 GNDA.n1103 GNDA.n1099 3.7893
R3364 GNDA.n1102 GNDA.n1076 3.7893
R3365 GNDA.n1110 GNDA.n1109 3.7893
R3366 GNDA.n1812 GNDA.n1733 3.7893
R3367 GNDA.n1809 GNDA.n1808 3.7893
R3368 GNDA.n1803 GNDA.n14 3.7893
R3369 GNDA.n2041 GNDA.n2040 3.7893
R3370 GNDA.n12 GNDA.n11 3.7893
R3371 GNDA.n7 GNDA.n3 3.7893
R3372 GNDA.n2052 GNDA.n8 3.7893
R3373 GNDA.n2051 GNDA.n9 3.7893
R3374 GNDA.n1694 GNDA.n1559 3.7893
R3375 GNDA.n1593 GNDA.n1592 3.7893
R3376 GNDA.n1598 GNDA.n1594 3.7893
R3377 GNDA.n1597 GNDA.n1585 3.7893
R3378 GNDA.n1623 GNDA.n1622 3.7893
R3379 GNDA.n1632 GNDA.n1628 3.7893
R3380 GNDA.n1631 GNDA.n1582 3.7893
R3381 GNDA.n1640 GNDA.n1639 3.7893
R3382 GNDA.n1490 GNDA.n201 3.51962
R3383 GNDA.t28 GNDA.n1635 3.08966
R3384 GNDA.t109 GNDA.n178 3.08966
R3385 GNDA.t108 GNDA.n191 3.08966
R3386 GNDA.t19 GNDA.n1847 3.08966
R3387 GNDA.n1848 GNDA.n17 3.08966
R3388 GNDA.n731 GNDA 2.9189
R3389 GNDA.n1839 GNDA 2.9189
R3390 GNDA.n860 GNDA 2.9189
R3391 GNDA.n595 GNDA 2.9189
R3392 GNDA.n1267 GNDA 2.9189
R3393 GNDA.n296 GNDA 2.9189
R3394 GNDA.n1098 GNDA 2.9189
R3395 GNDA GNDA.n2058 2.9189
R3396 GNDA.n1627 GNDA 2.9189
R3397 GNDA.n1825 GNDA.n1824 2.86505
R3398 GNDA.n1824 GNDA.n1822 2.86505
R3399 GNDA.n1822 GNDA.n1821 2.86505
R3400 GNDA.n1826 GNDA.n1825 2.86505
R3401 GNDA.n1606 GNDA.n1605 2.86505
R3402 GNDA.n1607 GNDA.n1606 2.86505
R3403 GNDA.n1611 GNDA.n1609 2.86505
R3404 GNDA.n1614 GNDA.n1609 2.86505
R3405 GNDA.n1610 GNDA.n1607 2.86505
R3406 GNDA.n1614 GNDA.n1613 2.86505
R3407 GNDA.n1616 GNDA.n1605 2.86505
R3408 GNDA.n1611 GNDA.n1610 2.86505
R3409 GNDA.n704 GNDA.n435 2.6629
R3410 GNDA.n745 GNDA.n625 2.6629
R3411 GNDA.n1909 GNDA.n130 2.6629
R3412 GNDA.n171 GNDA.n170 2.6629
R3413 GNDA.n1005 GNDA.n746 2.6629
R3414 GNDA.n930 GNDA.n815 2.6629
R3415 GNDA.n620 GNDA.n619 2.6629
R3416 GNDA.n1244 GNDA.n1049 2.6629
R3417 GNDA.n273 GNDA.n231 2.6629
R3418 GNDA.n366 GNDA.n250 2.6629
R3419 GNDA.n1431 GNDA.n1169 2.6629
R3420 GNDA.n1075 GNDA.n1074 2.6629
R3421 GNDA.n1731 GNDA.n76 2.6629
R3422 GNDA.n1748 GNDA.n1747 2.6629
R3423 GNDA.n1581 GNDA.n1580 2.6629
R3424 GNDA.n704 GNDA.n703 2.4581
R3425 GNDA.n1005 GNDA.n745 2.4581
R3426 GNDA.n1909 GNDA.n1908 2.4581
R3427 GNDA.n834 GNDA.n746 2.4581
R3428 GNDA.n581 GNDA.n580 2.4581
R3429 GNDA.n620 GNDA.n435 2.4581
R3430 GNDA.n1221 GNDA.n1219 2.4581
R3431 GNDA.n1431 GNDA.n1049 2.4581
R3432 GNDA.n273 GNDA.n269 2.4581
R3433 GNDA.n1169 GNDA.n1050 2.4581
R3434 GNDA.n1074 GNDA.n231 2.4581
R3435 GNDA.n1732 GNDA.n1731 2.4581
R3436 GNDA.n1747 GNDA.n130 2.4581
R3437 GNDA.n1697 GNDA.n1696 2.4581
R3438 GNDA.n1580 GNDA.n76 2.4581
R3439 GNDA.n1438 GNDA.n231 2.18124
R3440 GNDA.n1005 GNDA.n1004 2.18124
R3441 GNDA.n1924 GNDA.n130 2.18124
R3442 GNDA.n2004 GNDA.n76 2.18124
R3443 GNDA.n1013 GNDA.n435 2.18124
R3444 GNDA.n1431 GNDA.n1430 2.18124
R3445 GNDA.n709 GNDA.n703 2.1509
R3446 GNDA.n1908 GNDA.n1907 2.1509
R3447 GNDA.n836 GNDA.n834 2.1509
R3448 GNDA.n580 GNDA.n463 2.1509
R3449 GNDA.n1335 GNDA.n1221 2.1509
R3450 GNDA.n271 GNDA.n269 2.1509
R3451 GNDA.n1165 GNDA.n1050 2.1509
R3452 GNDA.n1813 GNDA.n1732 2.1509
R3453 GNDA.n1696 GNDA.n1695 2.1509
R3454 GNDA.n1643 GNDA.n1581 2.13383
R3455 GNDA.n1113 GNDA.n1075 2.13383
R3456 GNDA.n650 GNDA.n625 2.13383
R3457 GNDA.n1855 GNDA.n171 2.13383
R3458 GNDA.n930 GNDA.n929 2.13383
R3459 GNDA.n619 GNDA.n437 2.13383
R3460 GNDA.n1283 GNDA.n1244 2.13383
R3461 GNDA.n366 GNDA.n365 2.13383
R3462 GNDA.n1749 GNDA.n1748 2.13383
R3463 GNDA.n1493 GNDA 2.09787
R3464 GNDA.n233 GNDA.n231 2.08643
R3465 GNDA.n1006 GNDA.n1005 2.08643
R3466 GNDA.n132 GNDA.n130 2.08643
R3467 GNDA.n1725 GNDA.n76 2.08643
R3468 GNDA.n622 GNDA.n435 2.08643
R3469 GNDA.n1432 GNDA.n1431 2.08643
R3470 GNDA.n1637 GNDA.t83 2.05994
R3471 GNDA.n1728 GNDA.t94 2.05994
R3472 GNDA.t100 GNDA.n133 2.05994
R3473 GNDA.n178 GNDA.t103 2.05994
R3474 GNDA.n1433 GNDA.n419 1.951
R3475 GNDA.n1726 GNDA.n75 1.951
R3476 GNDA.n1008 GNDA.n434 1.951
R3477 GNDA.n145 GNDA.n129 1.951
R3478 GNDA.n1007 GNDA.n624 1.951
R3479 GNDA.n1501 GNDA.n1498 1.951
R3480 GNDA.n528 GNDA.n465 1.951
R3481 GNDA.n1341 GNDA.n1339 1.951
R3482 GNDA.n418 GNDA.n230 1.951
R3483 GNDA.n741 GNDA.n625 1.9461
R3484 GNDA.n1851 GNDA.n171 1.9461
R3485 GNDA.n931 GNDA.n930 1.9461
R3486 GNDA.n619 GNDA.n618 1.9461
R3487 GNDA.n1279 GNDA.n1244 1.9461
R3488 GNDA.n367 GNDA.n366 1.9461
R3489 GNDA.n1109 GNDA.n1075 1.9461
R3490 GNDA.n1748 GNDA.n9 1.9461
R3491 GNDA.n1639 GNDA.n1581 1.9461
R3492 GNDA.n1489 GNDA.n1488 1.90675
R3493 GNDA.n2028 GNDA.n19 1.52512
R3494 GNDA.n939 GNDA.n938 1.52512
R3495 GNDA.n374 GNDA.n373 1.52512
R3496 GNDA.n1557 GNDA.n1500 1.42272
R3497 GNDA.n529 GNDA.n466 1.42272
R3498 GNDA.n1343 GNDA.n1342 1.42272
R3499 GNDA.n1916 GNDA.n1915 0.96925
R3500 GNDA.n1719 GNDA.n1718 0.96925
R3501 GNDA GNDA.n730 0.8709
R3502 GNDA GNDA.n1838 0.8709
R3503 GNDA.n855 GNDA 0.8709
R3504 GNDA GNDA.n593 0.8709
R3505 GNDA GNDA.n1266 0.8709
R3506 GNDA.n291 GNDA 0.8709
R3507 GNDA GNDA.n1097 0.8709
R3508 GNDA GNDA.n2 0.8709
R3509 GNDA GNDA.n1626 0.8709
R3510 GNDA.n710 GNDA.n709 0.8197
R3511 GNDA.n714 GNDA.n636 0.8197
R3512 GNDA.n716 GNDA.n715 0.8197
R3513 GNDA.n724 GNDA.n634 0.8197
R3514 GNDA.n723 GNDA.n632 0.8197
R3515 GNDA.n731 GNDA.n630 0.8197
R3516 GNDA.n736 GNDA.n735 0.8197
R3517 GNDA.n740 GNDA.n627 0.8197
R3518 GNDA.n1907 GNDA.n1906 0.8197
R3519 GNDA.n182 GNDA.n149 0.8197
R3520 GNDA.n184 GNDA.n183 0.8197
R3521 GNDA.n188 GNDA.n187 0.8197
R3522 GNDA.n1835 GNDA.n175 0.8197
R3523 GNDA.n1840 GNDA.n1839 0.8197
R3524 GNDA.n1844 GNDA.n1843 0.8197
R3525 GNDA.n1852 GNDA.n172 0.8197
R3526 GNDA.n876 GNDA.n836 0.8197
R3527 GNDA.n875 GNDA.n837 0.8197
R3528 GNDA.n871 GNDA.n870 0.8197
R3529 GNDA.n866 GNDA.n842 0.8197
R3530 GNDA.n865 GNDA.n844 0.8197
R3531 GNDA.n860 GNDA.n859 0.8197
R3532 GNDA.n852 GNDA.n849 0.8197
R3533 GNDA.n851 GNDA.n817 0.8197
R3534 GNDA.n610 GNDA.n463 0.8197
R3535 GNDA.n609 GNDA.n464 0.8197
R3536 GNDA.n605 GNDA.n604 0.8197
R3537 GNDA.n601 GNDA.n586 0.8197
R3538 GNDA.n600 GNDA.n587 0.8197
R3539 GNDA.n595 GNDA.n594 0.8197
R3540 GNDA.n614 GNDA.n440 0.8197
R3541 GNDA.n615 GNDA.n438 0.8197
R3542 GNDA.n1335 GNDA.n1334 0.8197
R3543 GNDA.n1250 GNDA.n1222 0.8197
R3544 GNDA.n1252 GNDA.n1251 0.8197
R3545 GNDA.n1256 GNDA.n1255 0.8197
R3546 GNDA.n1263 GNDA.n1247 0.8197
R3547 GNDA.n1268 GNDA.n1267 0.8197
R3548 GNDA.n1272 GNDA.n1271 0.8197
R3549 GNDA.n1280 GNDA.n1245 0.8197
R3550 GNDA.n312 GNDA.n271 0.8197
R3551 GNDA.n311 GNDA.n272 0.8197
R3552 GNDA.n307 GNDA.n306 0.8197
R3553 GNDA.n302 GNDA.n278 0.8197
R3554 GNDA.n301 GNDA.n280 0.8197
R3555 GNDA.n296 GNDA.n295 0.8197
R3556 GNDA.n288 GNDA.n285 0.8197
R3557 GNDA.n287 GNDA.n252 0.8197
R3558 GNDA.n1165 GNDA.n1164 0.8197
R3559 GNDA.n1081 GNDA.n1052 0.8197
R3560 GNDA.n1083 GNDA.n1082 0.8197
R3561 GNDA.n1087 GNDA.n1086 0.8197
R3562 GNDA.n1094 GNDA.n1078 0.8197
R3563 GNDA.n1099 GNDA.n1098 0.8197
R3564 GNDA.n1103 GNDA.n1102 0.8197
R3565 GNDA.n1110 GNDA.n1076 0.8197
R3566 GNDA.n1813 GNDA.n1812 0.8197
R3567 GNDA.n1809 GNDA.n1733 0.8197
R3568 GNDA.n1808 GNDA.n1803 0.8197
R3569 GNDA.n2041 GNDA.n14 0.8197
R3570 GNDA.n2040 GNDA.n12 0.8197
R3571 GNDA.n2058 GNDA.n3 0.8197
R3572 GNDA.n8 GNDA.n7 0.8197
R3573 GNDA.n2052 GNDA.n2051 0.8197
R3574 GNDA.n1695 GNDA.n1694 0.8197
R3575 GNDA.n1592 GNDA.n1559 0.8197
R3576 GNDA.n1594 GNDA.n1593 0.8197
R3577 GNDA.n1598 GNDA.n1597 0.8197
R3578 GNDA.n1623 GNDA.n1585 0.8197
R3579 GNDA.n1628 GNDA.n1627 0.8197
R3580 GNDA.n1632 GNDA.n1631 0.8197
R3581 GNDA.n1640 GNDA.n1582 0.8197
R3582 GNDA.n142 GNDA.n140 0.563
R3583 GNDA.n144 GNDA.n142 0.563
R3584 GNDA.n1915 GNDA.n144 0.563
R3585 GNDA.n1916 GNDA.n136 0.563
R3586 GNDA.n1711 GNDA.n136 0.563
R3587 GNDA.n1713 GNDA.n1711 0.563
R3588 GNDA.n1715 GNDA.n1713 0.563
R3589 GNDA.n1718 GNDA.n1715 0.563
R3590 GNDA.n1719 GNDA.n1709 0.563
R3591 GNDA.n1709 GNDA.n1707 0.563
R3592 GNDA.n1707 GNDA.n1705 0.563
R3593 GNDA.n1705 GNDA.n1703 0.563
R3594 GNDA.n720 GNDA 0.5125
R3595 GNDA.n1834 GNDA 0.5125
R3596 GNDA GNDA.n846 0.5125
R3597 GNDA GNDA.n589 0.5125
R3598 GNDA.n1262 GNDA 0.5125
R3599 GNDA GNDA.n282 0.5125
R3600 GNDA.n1093 GNDA 0.5125
R3601 GNDA.n11 GNDA 0.5125
R3602 GNDA.n1622 GNDA 0.5125
R3603 GNDA.n730 GNDA 0.3077
R3604 GNDA.n1838 GNDA 0.3077
R3605 GNDA.n855 GNDA 0.3077
R3606 GNDA.n593 GNDA 0.3077
R3607 GNDA.n1266 GNDA 0.3077
R3608 GNDA.n291 GNDA 0.3077
R3609 GNDA.n1097 GNDA 0.3077
R3610 GNDA GNDA.n2 0.3077
R3611 GNDA.n1626 GNDA 0.3077
R3612 GNDA.n1494 GNDA.n1493 0.276625
R3613 GNDA.n1494 GNDA.n201 0.22375
R3614 V_mir2.n5 V_mir2.n1 325.473
R3615 V_mir2.n10 V_mir2.n6 325.471
R3616 V_mir2.n19 V_mir2.n18 325.471
R3617 V_mir2.n15 V_mir2.t21 310.488
R3618 V_mir2.n7 V_mir2.t20 310.488
R3619 V_mir2.n2 V_mir2.t17 310.488
R3620 V_mir2.n13 V_mir2.t1 278.312
R3621 V_mir2.n13 V_mir2.n12 228.939
R3622 V_mir2.n0 V_mir2.n11 224.439
R3623 V_mir2.n17 V_mir2.t3 184.097
R3624 V_mir2.n9 V_mir2.t9 184.097
R3625 V_mir2.n4 V_mir2.t11 184.097
R3626 V_mir2.n16 V_mir2.n15 167.094
R3627 V_mir2.n8 V_mir2.n7 167.094
R3628 V_mir2.n3 V_mir2.n2 167.094
R3629 V_mir2.n10 V_mir2.n9 152
R3630 V_mir2.n5 V_mir2.n4 152
R3631 V_mir2.n18 V_mir2.n17 152
R3632 V_mir2.n15 V_mir2.t22 120.501
R3633 V_mir2.n16 V_mir2.t13 120.501
R3634 V_mir2.n7 V_mir2.t19 120.501
R3635 V_mir2.n8 V_mir2.t7 120.501
R3636 V_mir2.n2 V_mir2.t18 120.501
R3637 V_mir2.n3 V_mir2.t5 120.501
R3638 V_mir2.n12 V_mir2.t16 48.0005
R3639 V_mir2.n12 V_mir2.t0 48.0005
R3640 V_mir2.n11 V_mir2.t2 48.0005
R3641 V_mir2.n11 V_mir2.t15 48.0005
R3642 V_mir2.n17 V_mir2.n16 40.7027
R3643 V_mir2.n9 V_mir2.n8 40.7027
R3644 V_mir2.n4 V_mir2.n3 40.7027
R3645 V_mir2.n6 V_mir2.t10 39.4005
R3646 V_mir2.n6 V_mir2.t8 39.4005
R3647 V_mir2.n1 V_mir2.t12 39.4005
R3648 V_mir2.n1 V_mir2.t6 39.4005
R3649 V_mir2.t4 V_mir2.n19 39.4005
R3650 V_mir2.n19 V_mir2.t14 39.4005
R3651 V_mir2.n14 V_mir2.n5 15.8005
R3652 V_mir2.n18 V_mir2.n14 15.8005
R3653 V_mir2.n0 V_mir2.n10 9.3005
R3654 V_mir2.n0 V_mir2.n13 5.8755
R3655 V_mir2.n14 V_mir2.n0 5.28175
R3656 VDDA.n129 VDDA.t153 676.966
R3657 VDDA.n90 VDDA.t165 660.001
R3658 VDDA.n26 VDDA.t135 645.231
R3659 VDDA.t159 VDDA.n25 645.231
R3660 VDDA.t171 VDDA.n164 643.038
R3661 VDDA.n165 VDDA.t147 643.038
R3662 VDDA.t138 VDDA.n128 643.038
R3663 VDDA.n32 VDDA.t144 643.037
R3664 VDDA.t174 VDDA.n31 643.037
R3665 VDDA.n20 VDDA.t177 643.037
R3666 VDDA.t162 VDDA.n19 643.037
R3667 VDDA.n150 VDDA.n105 587.407
R3668 VDDA.n152 VDDA.n151 587.407
R3669 VDDA.n144 VDDA.n143 587.407
R3670 VDDA.n136 VDDA.n135 587.407
R3671 VDDA.n156 VDDA.n150 585
R3672 VDDA.n155 VDDA.n151 585
R3673 VDDA.n143 VDDA.n142 585
R3674 VDDA.n139 VDDA.n135 585
R3675 VDDA.n98 VDDA.t150 540.818
R3676 VDDA.t141 VDDA.n97 540.818
R3677 VDDA.t156 VDDA.n89 540.818
R3678 VDDA.n163 VDDA.t170 419.108
R3679 VDDA.n166 VDDA.t146 419.108
R3680 VDDA.n127 VDDA.t137 413.084
R3681 VDDA.n130 VDDA.t152 413.084
R3682 VDDA.n30 VDDA.t173 409.067
R3683 VDDA.n33 VDDA.t143 409.067
R3684 VDDA.n24 VDDA.t158 409.067
R3685 VDDA.n27 VDDA.t134 409.067
R3686 VDDA.n18 VDDA.t161 409.067
R3687 VDDA.t150 VDDA.t208 407.144
R3688 VDDA.t208 VDDA.t125 407.144
R3689 VDDA.t125 VDDA.t129 407.144
R3690 VDDA.t129 VDDA.t107 407.144
R3691 VDDA.t107 VDDA.t113 407.144
R3692 VDDA.t113 VDDA.t206 407.144
R3693 VDDA.t206 VDDA.t212 407.144
R3694 VDDA.t212 VDDA.t109 407.144
R3695 VDDA.t109 VDDA.t115 407.144
R3696 VDDA.t115 VDDA.t121 407.144
R3697 VDDA.t121 VDDA.t117 407.144
R3698 VDDA.t117 VDDA.t210 407.144
R3699 VDDA.t210 VDDA.t202 407.144
R3700 VDDA.t202 VDDA.t111 407.144
R3701 VDDA.t111 VDDA.t119 407.144
R3702 VDDA.t119 VDDA.t123 407.144
R3703 VDDA.t123 VDDA.t127 407.144
R3704 VDDA.t127 VDDA.t204 407.144
R3705 VDDA.t204 VDDA.t141 407.144
R3706 VDDA.t165 VDDA.t196 407.144
R3707 VDDA.t196 VDDA.t101 407.144
R3708 VDDA.t101 VDDA.t8 407.144
R3709 VDDA.t8 VDDA.t5 407.144
R3710 VDDA.t5 VDDA.t35 407.144
R3711 VDDA.t35 VDDA.t194 407.144
R3712 VDDA.t194 VDDA.t179 407.144
R3713 VDDA.t179 VDDA.t83 407.144
R3714 VDDA.t83 VDDA.t103 407.144
R3715 VDDA.t103 VDDA.t188 407.144
R3716 VDDA.t188 VDDA.t105 407.144
R3717 VDDA.t105 VDDA.t77 407.144
R3718 VDDA.t77 VDDA.t53 407.144
R3719 VDDA.t53 VDDA.t37 407.144
R3720 VDDA.t37 VDDA.t59 407.144
R3721 VDDA.t59 VDDA.t87 407.144
R3722 VDDA.t87 VDDA.t97 407.144
R3723 VDDA.t97 VDDA.t14 407.144
R3724 VDDA.t14 VDDA.t156 407.144
R3725 VDDA.n21 VDDA.t176 390.322
R3726 VDDA.t140 VDDA.n50 379.582
R3727 VDDA.t155 VDDA.n69 379.582
R3728 VDDA.t149 VDDA.n99 379.277
R3729 VDDA.t144 VDDA.t99 373.214
R3730 VDDA.t99 VDDA.t17 373.214
R3731 VDDA.t17 VDDA.t65 373.214
R3732 VDDA.t65 VDDA.t39 373.214
R3733 VDDA.t39 VDDA.t174 373.214
R3734 VDDA.t135 VDDA.t200 373.214
R3735 VDDA.t200 VDDA.t89 373.214
R3736 VDDA.t89 VDDA.t30 373.214
R3737 VDDA.t30 VDDA.t61 373.214
R3738 VDDA.t61 VDDA.t48 373.214
R3739 VDDA.t48 VDDA.t67 373.214
R3740 VDDA.t67 VDDA.t23 373.214
R3741 VDDA.t23 VDDA.t46 373.214
R3742 VDDA.t46 VDDA.t73 373.214
R3743 VDDA.t73 VDDA.t192 373.214
R3744 VDDA.t192 VDDA.t159 373.214
R3745 VDDA.t177 VDDA.t63 373.214
R3746 VDDA.t63 VDDA.t91 373.214
R3747 VDDA.t91 VDDA.t28 373.214
R3748 VDDA.t28 VDDA.t190 373.214
R3749 VDDA.t190 VDDA.t162 373.214
R3750 VDDA.t85 VDDA.t171 373.214
R3751 VDDA.t75 VDDA.t85 373.214
R3752 VDDA.t147 VDDA.t75 373.214
R3753 VDDA.t153 VDDA.t34 373.214
R3754 VDDA.t34 VDDA.t13 373.214
R3755 VDDA.t13 VDDA.t138 373.214
R3756 VDDA.n133 VDDA.t167 360.868
R3757 VDDA.n161 VDDA.t131 360.868
R3758 VDDA.n100 VDDA.t149 358.858
R3759 VDDA.n94 VDDA.t140 358.858
R3760 VDDA.n91 VDDA.t164 358.858
R3761 VDDA.n86 VDDA.t155 358.858
R3762 VDDA.n26 VDDA.t136 354.154
R3763 VDDA.n25 VDDA.t160 354.154
R3764 VDDA.n165 VDDA.t148 354.065
R3765 VDDA.n128 VDDA.t139 354.065
R3766 VDDA.n90 VDDA.t166 354.065
R3767 VDDA.n164 VDDA.t172 354.063
R3768 VDDA.n49 VDDA.t151 351.793
R3769 VDDA.n95 VDDA.t142 351.793
R3770 VDDA.n87 VDDA.t157 351.793
R3771 VDDA.n129 VDDA.t154 347.224
R3772 VDDA.n15 VDDA.n14 345.127
R3773 VDDA.n17 VDDA.n16 345.127
R3774 VDDA.n1 VDDA.n0 344.7
R3775 VDDA.n3 VDDA.n2 344.7
R3776 VDDA.n47 VDDA.n46 341.676
R3777 VDDA.n52 VDDA.n51 341.676
R3778 VDDA.n54 VDDA.n53 341.676
R3779 VDDA.n56 VDDA.n55 341.676
R3780 VDDA.n58 VDDA.n57 341.676
R3781 VDDA.n60 VDDA.n59 341.676
R3782 VDDA.n62 VDDA.n61 341.676
R3783 VDDA.n64 VDDA.n63 341.676
R3784 VDDA.n66 VDDA.n65 341.676
R3785 VDDA.n68 VDDA.n67 341.676
R3786 VDDA.n71 VDDA.n70 341.676
R3787 VDDA.n73 VDDA.n72 341.676
R3788 VDDA.n75 VDDA.n74 341.676
R3789 VDDA.n77 VDDA.n76 341.676
R3790 VDDA.n79 VDDA.n78 341.676
R3791 VDDA.n81 VDDA.n80 341.676
R3792 VDDA.n83 VDDA.n82 341.676
R3793 VDDA.n85 VDDA.n84 341.676
R3794 VDDA.n5 VDDA.n4 339.272
R3795 VDDA.n7 VDDA.n6 339.272
R3796 VDDA.n9 VDDA.n8 339.272
R3797 VDDA.n11 VDDA.n10 339.272
R3798 VDDA.n13 VDDA.n12 339.272
R3799 VDDA.n169 VDDA.n168 334.772
R3800 VDDA.n20 VDDA.t178 332.267
R3801 VDDA.n19 VDDA.t163 332.267
R3802 VDDA.n32 VDDA.t145 332.084
R3803 VDDA.n31 VDDA.t175 332.084
R3804 VDDA.t132 VDDA.t181 251.471
R3805 VDDA.t181 VDDA.t10 251.471
R3806 VDDA.t10 VDDA.t95 251.471
R3807 VDDA.t95 VDDA.t32 251.471
R3808 VDDA.t32 VDDA.t41 251.471
R3809 VDDA.t41 VDDA.t21 251.471
R3810 VDDA.t21 VDDA.t184 251.471
R3811 VDDA.t184 VDDA.t3 251.471
R3812 VDDA.t3 VDDA.t1 251.471
R3813 VDDA.t1 VDDA.t81 251.471
R3814 VDDA.t81 VDDA.t44 251.471
R3815 VDDA.t44 VDDA.t51 251.471
R3816 VDDA.t51 VDDA.t56 251.471
R3817 VDDA.t56 VDDA.t79 251.471
R3818 VDDA.t79 VDDA.t93 251.471
R3819 VDDA.t93 VDDA.t186 251.471
R3820 VDDA.t186 VDDA.t168 251.471
R3821 VDDA.n160 VDDA.n159 238.367
R3822 VDDA.n98 VDDA.n48 238.367
R3823 VDDA.n99 VDDA.n98 238.367
R3824 VDDA.n97 VDDA.n50 238.367
R3825 VDDA.n97 VDDA.n96 238.367
R3826 VDDA.n89 VDDA.n69 238.367
R3827 VDDA.n89 VDDA.n88 238.367
R3828 VDDA.n158 VDDA.t132 237.5
R3829 VDDA.t168 VDDA.n147 237.5
R3830 VDDA.n152 VDDA.n108 190.333
R3831 VDDA.n136 VDDA.n111 190.333
R3832 VDDA.n149 VDDA.n106 185
R3833 VDDA.n157 VDDA.n156 185
R3834 VDDA.n158 VDDA.n157 185
R3835 VDDA.n155 VDDA.n148 185
R3836 VDDA.n154 VDDA.n153 185
R3837 VDDA.n158 VDDA.n108 185
R3838 VDDA.n146 VDDA.n145 185
R3839 VDDA.n147 VDDA.n146 185
R3840 VDDA.n134 VDDA.n112 185
R3841 VDDA.n142 VDDA.n141 185
R3842 VDDA.n140 VDDA.n139 185
R3843 VDDA.n138 VDDA.n137 185
R3844 VDDA.n147 VDDA.n111 185
R3845 VDDA.n104 VDDA.n103 168.435
R3846 VDDA.n114 VDDA.n113 168.435
R3847 VDDA.n116 VDDA.n115 168.435
R3848 VDDA.n118 VDDA.n117 168.435
R3849 VDDA.n120 VDDA.n119 168.435
R3850 VDDA.n122 VDDA.n121 168.435
R3851 VDDA.n124 VDDA.n123 168.435
R3852 VDDA.n126 VDDA.n125 168.435
R3853 VDDA.n157 VDDA.n106 150
R3854 VDDA.n157 VDDA.n148 150
R3855 VDDA.n153 VDDA.n108 150
R3856 VDDA.n146 VDDA.n112 150
R3857 VDDA.n141 VDDA.n140 150
R3858 VDDA.n137 VDDA.n111 150
R3859 VDDA.t133 VDDA.n150 123.126
R3860 VDDA.n151 VDDA.t133 123.126
R3861 VDDA.n143 VDDA.t169 123.126
R3862 VDDA.n135 VDDA.t169 123.126
R3863 VDDA.n159 VDDA.n158 65.8183
R3864 VDDA.n158 VDDA.n107 65.8183
R3865 VDDA.n147 VDDA.n109 65.8183
R3866 VDDA.n147 VDDA.n110 65.8183
R3867 VDDA.n42 VDDA.t216 59.5681
R3868 VDDA.n43 VDDA.t215 59.5681
R3869 VDDA.n148 VDDA.n107 53.3664
R3870 VDDA.n159 VDDA.n106 53.3664
R3871 VDDA.n153 VDDA.n107 53.3664
R3872 VDDA.n112 VDDA.n109 53.3664
R3873 VDDA.n140 VDDA.n110 53.3664
R3874 VDDA.n141 VDDA.n109 53.3664
R3875 VDDA.n137 VDDA.n110 53.3664
R3876 VDDA.n42 VDDA.t217 52.3887
R3877 VDDA.n44 VDDA.t214 48.9557
R3878 VDDA.n0 VDDA.t100 39.4005
R3879 VDDA.n0 VDDA.t18 39.4005
R3880 VDDA.n2 VDDA.t66 39.4005
R3881 VDDA.n2 VDDA.t40 39.4005
R3882 VDDA.n4 VDDA.t201 39.4005
R3883 VDDA.n4 VDDA.t90 39.4005
R3884 VDDA.n6 VDDA.t31 39.4005
R3885 VDDA.n6 VDDA.t62 39.4005
R3886 VDDA.n8 VDDA.t49 39.4005
R3887 VDDA.n8 VDDA.t68 39.4005
R3888 VDDA.n10 VDDA.t24 39.4005
R3889 VDDA.n10 VDDA.t47 39.4005
R3890 VDDA.n12 VDDA.t74 39.4005
R3891 VDDA.n12 VDDA.t193 39.4005
R3892 VDDA.n14 VDDA.t64 39.4005
R3893 VDDA.n14 VDDA.t92 39.4005
R3894 VDDA.n16 VDDA.t29 39.4005
R3895 VDDA.n16 VDDA.t191 39.4005
R3896 VDDA.n168 VDDA.t86 39.4005
R3897 VDDA.n168 VDDA.t76 39.4005
R3898 VDDA.n46 VDDA.t209 39.4005
R3899 VDDA.n46 VDDA.t126 39.4005
R3900 VDDA.n51 VDDA.t130 39.4005
R3901 VDDA.n51 VDDA.t108 39.4005
R3902 VDDA.n53 VDDA.t114 39.4005
R3903 VDDA.n53 VDDA.t207 39.4005
R3904 VDDA.n55 VDDA.t213 39.4005
R3905 VDDA.n55 VDDA.t110 39.4005
R3906 VDDA.n57 VDDA.t116 39.4005
R3907 VDDA.n57 VDDA.t122 39.4005
R3908 VDDA.n59 VDDA.t118 39.4005
R3909 VDDA.n59 VDDA.t211 39.4005
R3910 VDDA.n61 VDDA.t203 39.4005
R3911 VDDA.n61 VDDA.t112 39.4005
R3912 VDDA.n63 VDDA.t120 39.4005
R3913 VDDA.n63 VDDA.t124 39.4005
R3914 VDDA.n65 VDDA.t128 39.4005
R3915 VDDA.n65 VDDA.t205 39.4005
R3916 VDDA.n67 VDDA.t197 39.4005
R3917 VDDA.n67 VDDA.t102 39.4005
R3918 VDDA.n70 VDDA.t9 39.4005
R3919 VDDA.n70 VDDA.t6 39.4005
R3920 VDDA.n72 VDDA.t36 39.4005
R3921 VDDA.n72 VDDA.t195 39.4005
R3922 VDDA.n74 VDDA.t180 39.4005
R3923 VDDA.n74 VDDA.t84 39.4005
R3924 VDDA.n76 VDDA.t104 39.4005
R3925 VDDA.n76 VDDA.t189 39.4005
R3926 VDDA.n78 VDDA.t106 39.4005
R3927 VDDA.n78 VDDA.t78 39.4005
R3928 VDDA.n80 VDDA.t54 39.4005
R3929 VDDA.n80 VDDA.t38 39.4005
R3930 VDDA.n82 VDDA.t60 39.4005
R3931 VDDA.n82 VDDA.t88 39.4005
R3932 VDDA.n84 VDDA.t98 39.4005
R3933 VDDA.n84 VDDA.t15 39.4005
R3934 VDDA.n41 VDDA.n35 33.7847
R3935 VDDA.n33 VDDA.n32 27.2462
R3936 VDDA.n31 VDDA.n30 27.2462
R3937 VDDA.n21 VDDA.n20 27.2462
R3938 VDDA.n19 VDDA.n18 27.2462
R3939 VDDA.n164 VDDA.n163 25.087
R3940 VDDA.n166 VDDA.n165 25.087
R3941 VDDA.n27 VDDA.n26 25.0384
R3942 VDDA.n25 VDDA.n24 25.0384
R3943 VDDA.n128 VDDA.n127 22.9536
R3944 VDDA.n91 VDDA.n90 22.9536
R3945 VDDA.n161 VDDA.n160 22.8576
R3946 VDDA.n145 VDDA.n133 22.8576
R3947 VDDA.n100 VDDA.n48 20.7243
R3948 VDDA.n96 VDDA.n94 20.7243
R3949 VDDA.n88 VDDA.n86 20.7243
R3950 VDDA.n130 VDDA.n129 20.4312
R3951 VDDA.n41 VDDA.t198 19.9244
R3952 VDDA.n131 VDDA.n127 15.488
R3953 VDDA.n86 VDDA.n85 14.6963
R3954 VDDA.n18 VDDA.n17 14.363
R3955 VDDA.n167 VDDA.n166 14.363
R3956 VDDA.n167 VDDA.n163 14.363
R3957 VDDA.n131 VDDA.n130 14.238
R3958 VDDA.n94 VDDA.n93 14.0713
R3959 VDDA.n101 VDDA.n100 14.0713
R3960 VDDA.n92 VDDA.n91 14.0713
R3961 VDDA.n30 VDDA.n29 13.8005
R3962 VDDA.n24 VDDA.n23 13.8005
R3963 VDDA.n22 VDDA.n21 13.8005
R3964 VDDA.n28 VDDA.n27 13.8005
R3965 VDDA.n34 VDDA.n33 13.8005
R3966 VDDA.n133 VDDA.n132 13.8005
R3967 VDDA.n162 VDDA.n161 13.8005
R3968 VDDA.n103 VDDA.t182 13.1338
R3969 VDDA.n103 VDDA.t11 13.1338
R3970 VDDA.n113 VDDA.t96 13.1338
R3971 VDDA.n113 VDDA.t33 13.1338
R3972 VDDA.n115 VDDA.t42 13.1338
R3973 VDDA.n115 VDDA.t22 13.1338
R3974 VDDA.n117 VDDA.t185 13.1338
R3975 VDDA.n117 VDDA.t4 13.1338
R3976 VDDA.n119 VDDA.t2 13.1338
R3977 VDDA.n119 VDDA.t82 13.1338
R3978 VDDA.n121 VDDA.t45 13.1338
R3979 VDDA.n121 VDDA.t52 13.1338
R3980 VDDA.n123 VDDA.t57 13.1338
R3981 VDDA.n123 VDDA.t80 13.1338
R3982 VDDA.n125 VDDA.t94 13.1338
R3983 VDDA.n125 VDDA.t187 13.1338
R3984 VDDA.n35 VDDA.n34 11.4105
R3985 VDDA.n45 VDDA.n44 11.1572
R3986 VDDA.n171 VDDA.n170 9.7855
R3987 VDDA.n156 VDDA.n149 9.14336
R3988 VDDA.n156 VDDA.n155 9.14336
R3989 VDDA.n155 VDDA.n154 9.14336
R3990 VDDA.n142 VDDA.n134 9.14336
R3991 VDDA.n142 VDDA.n139 9.14336
R3992 VDDA.n139 VDDA.n138 9.14336
R3993 VDDA.n102 VDDA.n101 8.973
R3994 VDDA.n160 VDDA.n105 5.33286
R3995 VDDA.n145 VDDA.n144 5.33286
R3996 VDDA.n170 VDDA.n169 5.0005
R3997 VDDA.n45 VDDA.n41 4.5595
R3998 VDDA.n99 VDDA.n49 4.54311
R3999 VDDA.n49 VDDA.n48 4.54311
R4000 VDDA.n95 VDDA.n50 4.54311
R4001 VDDA.n96 VDDA.n95 4.54311
R4002 VDDA.n87 VDDA.n69 4.54311
R4003 VDDA.n88 VDDA.n87 4.54311
R4004 VDDA.n169 VDDA.n167 4.5005
R4005 VDDA.n43 VDDA.n42 4.12334
R4006 VDDA.n149 VDDA.n105 3.75335
R4007 VDDA.n154 VDDA.n152 3.75335
R4008 VDDA.n144 VDDA.n134 3.75335
R4009 VDDA.n138 VDDA.n136 3.75335
R4010 VDDA.n44 VDDA.n43 3.43377
R4011 VDDA.n170 VDDA.n162 2.5005
R4012 VDDA.n93 VDDA.n92 1.8755
R4013 VDDA.n132 VDDA.n131 1.84425
R4014 VDDA.n23 VDDA.n22 1.813
R4015 VDDA.n29 VDDA.n28 1.813
R4016 VDDA.n132 VDDA.n126 1.0005
R4017 VDDA.n126 VDDA.n124 1.0005
R4018 VDDA.n124 VDDA.n122 1.0005
R4019 VDDA.n122 VDDA.n120 1.0005
R4020 VDDA.n120 VDDA.n118 1.0005
R4021 VDDA.n118 VDDA.n116 1.0005
R4022 VDDA.n116 VDDA.n114 1.0005
R4023 VDDA.n114 VDDA.n104 1.0005
R4024 VDDA.n162 VDDA.n104 1.0005
R4025 VDDA.n102 VDDA.n45 0.840625
R4026 VDDA.n171 VDDA.n102 0.74075
R4027 VDDA.n85 VDDA.n83 0.6255
R4028 VDDA.n83 VDDA.n81 0.6255
R4029 VDDA.n81 VDDA.n79 0.6255
R4030 VDDA.n79 VDDA.n77 0.6255
R4031 VDDA.n77 VDDA.n75 0.6255
R4032 VDDA.n75 VDDA.n73 0.6255
R4033 VDDA.n73 VDDA.n71 0.6255
R4034 VDDA.n71 VDDA.n68 0.6255
R4035 VDDA.n92 VDDA.n68 0.6255
R4036 VDDA.n93 VDDA.n66 0.6255
R4037 VDDA.n66 VDDA.n64 0.6255
R4038 VDDA.n64 VDDA.n62 0.6255
R4039 VDDA.n62 VDDA.n60 0.6255
R4040 VDDA.n60 VDDA.n58 0.6255
R4041 VDDA.n58 VDDA.n56 0.6255
R4042 VDDA.n56 VDDA.n54 0.6255
R4043 VDDA.n54 VDDA.n52 0.6255
R4044 VDDA.n52 VDDA.n47 0.6255
R4045 VDDA.n101 VDDA.n47 0.6255
R4046 VDDA.n17 VDDA.n15 0.563
R4047 VDDA.n22 VDDA.n15 0.563
R4048 VDDA.n23 VDDA.n13 0.563
R4049 VDDA.n13 VDDA.n11 0.563
R4050 VDDA.n11 VDDA.n9 0.563
R4051 VDDA.n9 VDDA.n7 0.563
R4052 VDDA.n7 VDDA.n5 0.563
R4053 VDDA.n28 VDDA.n5 0.563
R4054 VDDA.n29 VDDA.n3 0.563
R4055 VDDA.n3 VDDA.n1 0.563
R4056 VDDA.n34 VDDA.n1 0.563
R4057 VDDA VDDA.n171 0.41175
R4058 VDDA.t71 VDDA.t20 0.1603
R4059 VDDA.t12 VDDA.t58 0.1603
R4060 VDDA.t19 VDDA.t55 0.1603
R4061 VDDA.t72 VDDA.t27 0.1603
R4062 VDDA.t50 VDDA.t199 0.1603
R4063 VDDA.n37 VDDA.t25 0.159278
R4064 VDDA.n38 VDDA.t16 0.159278
R4065 VDDA.n39 VDDA.t43 0.159278
R4066 VDDA.n40 VDDA.t7 0.159278
R4067 VDDA.n40 VDDA.t71 0.1368
R4068 VDDA.n40 VDDA.t183 0.1368
R4069 VDDA.n39 VDDA.t12 0.1368
R4070 VDDA.n39 VDDA.t0 0.1368
R4071 VDDA.n38 VDDA.t19 0.1368
R4072 VDDA.n38 VDDA.t26 0.1368
R4073 VDDA.n37 VDDA.t72 0.1368
R4074 VDDA.n37 VDDA.t69 0.1368
R4075 VDDA.n36 VDDA.t50 0.1368
R4076 VDDA.n36 VDDA.t70 0.1368
R4077 VDDA VDDA.n35 0.135625
R4078 VDDA.t25 VDDA.n36 0.00152174
R4079 VDDA.t16 VDDA.n37 0.00152174
R4080 VDDA.t43 VDDA.n38 0.00152174
R4081 VDDA.t7 VDDA.n39 0.00152174
R4082 VDDA.t198 VDDA.n40 0.00152174
R4083 VB2_CUR_BIAS.n2 VB2_CUR_BIAS.n0 140.857
R4084 VB2_CUR_BIAS.n6 VB2_CUR_BIAS.n5 139.608
R4085 VB2_CUR_BIAS.n4 VB2_CUR_BIAS.n3 139.607
R4086 VB2_CUR_BIAS.n2 VB2_CUR_BIAS.n1 139.607
R4087 VB2_CUR_BIAS VB2_CUR_BIAS.n6 29.688
R4088 VB2_CUR_BIAS.n5 VB2_CUR_BIAS.t1 24.0005
R4089 VB2_CUR_BIAS.n5 VB2_CUR_BIAS.t7 24.0005
R4090 VB2_CUR_BIAS.n3 VB2_CUR_BIAS.t2 24.0005
R4091 VB2_CUR_BIAS.n3 VB2_CUR_BIAS.t5 24.0005
R4092 VB2_CUR_BIAS.n1 VB2_CUR_BIAS.t0 24.0005
R4093 VB2_CUR_BIAS.n1 VB2_CUR_BIAS.t3 24.0005
R4094 VB2_CUR_BIAS.n0 VB2_CUR_BIAS.t6 24.0005
R4095 VB2_CUR_BIAS.n0 VB2_CUR_BIAS.t4 24.0005
R4096 VB2_CUR_BIAS.n4 VB2_CUR_BIAS.n2 7.563
R4097 VB2_CUR_BIAS.n6 VB2_CUR_BIAS.n4 1.2505
R4098 a_38570_n6530.t0 a_38570_n6530.t1 178.133
R4099 a_38690_n7778.t0 a_38690_n7778.t1 178.133
R4100 1st_Vout_1.n12 1st_Vout_1.t32 355.293
R4101 1st_Vout_1.n0 1st_Vout_1.t19 346.8
R4102 1st_Vout_1.n1 1st_Vout_1.n5 339.522
R4103 1st_Vout_1.n13 1st_Vout_1.n12 339.522
R4104 1st_Vout_1.n3 1st_Vout_1.n7 335.022
R4105 1st_Vout_1.n9 1st_Vout_1.t10 275.909
R4106 1st_Vout_1.n9 1st_Vout_1.n8 227.909
R4107 1st_Vout_1.n3 1st_Vout_1.n10 222.034
R4108 1st_Vout_1.n11 1st_Vout_1.t28 184.097
R4109 1st_Vout_1.n11 1st_Vout_1.t36 184.097
R4110 1st_Vout_1.n6 1st_Vout_1.t24 184.097
R4111 1st_Vout_1.n6 1st_Vout_1.t30 184.097
R4112 1st_Vout_1.n1 1st_Vout_1.n11 166.05
R4113 1st_Vout_1.n1 1st_Vout_1.n6 166.05
R4114 1st_Vout_1.n0 1st_Vout_1.n4 54.2759
R4115 1st_Vout_1.n10 1st_Vout_1.t8 48.0005
R4116 1st_Vout_1.n10 1st_Vout_1.t3 48.0005
R4117 1st_Vout_1.n8 1st_Vout_1.t2 48.0005
R4118 1st_Vout_1.n8 1st_Vout_1.t9 48.0005
R4119 1st_Vout_1.n7 1st_Vout_1.t5 39.4005
R4120 1st_Vout_1.n7 1st_Vout_1.t7 39.4005
R4121 1st_Vout_1.n5 1st_Vout_1.t1 39.4005
R4122 1st_Vout_1.n5 1st_Vout_1.t4 39.4005
R4123 1st_Vout_1.n13 1st_Vout_1.t6 39.4005
R4124 1st_Vout_1.t0 1st_Vout_1.n13 39.4005
R4125 1st_Vout_1.n1 1st_Vout_1.n3 5.28175
R4126 1st_Vout_1.n2 1st_Vout_1.t23 4.8295
R4127 1st_Vout_1.n2 1st_Vout_1.t11 4.8295
R4128 1st_Vout_1.n2 1st_Vout_1.t18 4.8295
R4129 1st_Vout_1.n2 1st_Vout_1.t27 4.8295
R4130 1st_Vout_1.n2 1st_Vout_1.t34 4.8295
R4131 1st_Vout_1.n2 1st_Vout_1.t20 4.8295
R4132 1st_Vout_1.n4 1st_Vout_1.t15 4.8295
R4133 1st_Vout_1.n4 1st_Vout_1.t25 4.8295
R4134 1st_Vout_1.n4 1st_Vout_1.t31 4.8295
R4135 1st_Vout_1.n3 1st_Vout_1.n9 4.5005
R4136 1st_Vout_1.n2 1st_Vout_1.t21 4.5005
R4137 1st_Vout_1.n2 1st_Vout_1.t12 4.5005
R4138 1st_Vout_1.n2 1st_Vout_1.t16 4.5005
R4139 1st_Vout_1.n2 1st_Vout_1.t29 4.5005
R4140 1st_Vout_1.n2 1st_Vout_1.t33 4.5005
R4141 1st_Vout_1.n2 1st_Vout_1.t22 4.5005
R4142 1st_Vout_1.n4 1st_Vout_1.t14 4.5005
R4143 1st_Vout_1.n4 1st_Vout_1.t26 4.5005
R4144 1st_Vout_1.n4 1st_Vout_1.t17 4.5005
R4145 1st_Vout_1.n4 1st_Vout_1.t35 4.5005
R4146 1st_Vout_1.n4 1st_Vout_1.t13 4.5005
R4147 1st_Vout_1.n1 1st_Vout_1.n0 3.188
R4148 1st_Vout_1.n4 1st_Vout_1.n2 3.1025
R4149 1st_Vout_1.n12 1st_Vout_1.n1 2.0005
R4150 cap_res1.t0 cap_res1.t18 121.245
R4151 cap_res1.t1 cap_res1.t14 0.1603
R4152 cap_res1.t17 cap_res1.t16 0.1603
R4153 cap_res1.t3 cap_res1.t2 0.1603
R4154 cap_res1.t15 cap_res1.t13 0.1603
R4155 cap_res1.t11 cap_res1.t9 0.1603
R4156 cap_res1.n1 cap_res1.t19 0.159278
R4157 cap_res1.n2 cap_res1.t5 0.159278
R4158 cap_res1.n3 cap_res1.t10 0.159278
R4159 cap_res1.n4 cap_res1.t7 0.159278
R4160 cap_res1.n4 cap_res1.t4 0.1368
R4161 cap_res1.n4 cap_res1.t1 0.1368
R4162 cap_res1.n3 cap_res1.t8 0.1368
R4163 cap_res1.n3 cap_res1.t17 0.1368
R4164 cap_res1.n2 cap_res1.t12 0.1368
R4165 cap_res1.n2 cap_res1.t3 0.1368
R4166 cap_res1.n1 cap_res1.t6 0.1368
R4167 cap_res1.n1 cap_res1.t15 0.1368
R4168 cap_res1.n0 cap_res1.t20 0.1368
R4169 cap_res1.n0 cap_res1.t11 0.1368
R4170 cap_res1.t19 cap_res1.n0 0.00152174
R4171 cap_res1.t5 cap_res1.n1 0.00152174
R4172 cap_res1.t10 cap_res1.n2 0.00152174
R4173 cap_res1.t7 cap_res1.n3 0.00152174
R4174 cap_res1.t18 cap_res1.n4 0.00152174
R4175 V_CMFB_S4.n2 V_CMFB_S4.n0 144.827
R4176 V_CMFB_S4.n2 V_CMFB_S4.n1 134.577
R4177 V_CMFB_S4 V_CMFB_S4.n2 37.563
R4178 V_CMFB_S4.n1 V_CMFB_S4.t2 24.0005
R4179 V_CMFB_S4.n1 V_CMFB_S4.t1 24.0005
R4180 V_CMFB_S4.n0 V_CMFB_S4.t0 24.0005
R4181 V_CMFB_S4.n0 V_CMFB_S4.t3 24.0005
R4182 Vin+.n3 Vin+.n2 526.183
R4183 Vin+.n1 Vin+.n0 514.134
R4184 Vin+.n0 Vin+.t9 303.259
R4185 Vin+.n5 Vin+.n3 227.169
R4186 Vin+.n0 Vin+.t7 174.726
R4187 Vin+.n1 Vin+.t6 174.726
R4188 Vin+.n2 Vin+.t10 174.726
R4189 Vin+.n5 Vin+.n4 168.435
R4190 Vin+.n7 Vin+.n6 168.435
R4191 Vin+.t0 Vin+.n8 158.989
R4192 Vin+.n2 Vin+.n1 128.534
R4193 Vin+.n8 Vin+.t1 119.067
R4194 Vin+.n3 Vin+.t8 96.4005
R4195 Vin+.n8 Vin+.n7 35.0317
R4196 Vin+.n6 Vin+.t2 13.1338
R4197 Vin+.n6 Vin+.t5 13.1338
R4198 Vin+.n4 Vin+.t4 13.1338
R4199 Vin+.n4 Vin+.t3 13.1338
R4200 Vin+.n7 Vin+.n5 2.1255
R4201 V_p_1.n1 V_p_1.n2 229.562
R4202 V_p_1.n1 V_p_1.n5 228.939
R4203 V_p_1.n0 V_p_1.n4 228.939
R4204 V_p_1.n0 V_p_1.n3 228.939
R4205 V_p_1.n6 V_p_1.n1 228.938
R4206 V_p_1.n0 V_p_1.t5 98.7282
R4207 V_p_1.n5 V_p_1.t1 48.0005
R4208 V_p_1.n5 V_p_1.t10 48.0005
R4209 V_p_1.n4 V_p_1.t6 48.0005
R4210 V_p_1.n4 V_p_1.t3 48.0005
R4211 V_p_1.n3 V_p_1.t2 48.0005
R4212 V_p_1.n3 V_p_1.t8 48.0005
R4213 V_p_1.n2 V_p_1.t4 48.0005
R4214 V_p_1.n2 V_p_1.t7 48.0005
R4215 V_p_1.t9 V_p_1.n6 48.0005
R4216 V_p_1.n6 V_p_1.t0 48.0005
R4217 V_p_1.n1 V_p_1.n0 1.8755
R4218 ERR_AMP_REF.n0 ERR_AMP_REF.t8 688.859
R4219 ERR_AMP_REF.n2 ERR_AMP_REF.n1 514.134
R4220 ERR_AMP_REF.n4 ERR_AMP_REF.n3 214.056
R4221 ERR_AMP_REF.n0 ERR_AMP_REF.t11 174.726
R4222 ERR_AMP_REF.n1 ERR_AMP_REF.t7 174.726
R4223 ERR_AMP_REF.n2 ERR_AMP_REF.t9 174.726
R4224 ERR_AMP_REF.n3 ERR_AMP_REF.t10 174.726
R4225 ERR_AMP_REF.n7 ERR_AMP_REF.n5 173.591
R4226 ERR_AMP_REF.n9 ERR_AMP_REF.n8 169.215
R4227 ERR_AMP_REF.n7 ERR_AMP_REF.n6 169.215
R4228 ERR_AMP_REF.n1 ERR_AMP_REF.n0 128.534
R4229 ERR_AMP_REF.n3 ERR_AMP_REF.n2 128.534
R4230 ERR_AMP_REF.n4 ERR_AMP_REF.t2 125.817
R4231 ERR_AMP_REF.n8 ERR_AMP_REF.t3 13.1338
R4232 ERR_AMP_REF.n8 ERR_AMP_REF.t5 13.1338
R4233 ERR_AMP_REF.n6 ERR_AMP_REF.t1 13.1338
R4234 ERR_AMP_REF.n6 ERR_AMP_REF.t0 13.1338
R4235 ERR_AMP_REF.n5 ERR_AMP_REF.t6 13.1338
R4236 ERR_AMP_REF.n5 ERR_AMP_REF.t4 13.1338
R4237 ERR_AMP_REF.n10 ERR_AMP_REF.n9 10.0317
R4238 ERR_AMP_REF ERR_AMP_REF.n10 8.09425
R4239 ERR_AMP_REF.n9 ERR_AMP_REF.n7 4.3755
R4240 ERR_AMP_REF.n10 ERR_AMP_REF.n4 3.03175
R4241 V_p_2.n1 V_p_2.n4 229.562
R4242 V_p_2.n1 V_p_2.n5 228.939
R4243 V_p_2.n0 V_p_2.n3 228.939
R4244 V_p_2.n0 V_p_2.n2 228.939
R4245 V_p_2.n6 V_p_2.n0 228.938
R4246 V_p_2.n0 V_p_2.t10 98.7282
R4247 V_p_2.n5 V_p_2.t0 48.0005
R4248 V_p_2.n5 V_p_2.t7 48.0005
R4249 V_p_2.n4 V_p_2.t9 48.0005
R4250 V_p_2.n4 V_p_2.t3 48.0005
R4251 V_p_2.n3 V_p_2.t2 48.0005
R4252 V_p_2.n3 V_p_2.t5 48.0005
R4253 V_p_2.n2 V_p_2.t6 48.0005
R4254 V_p_2.n2 V_p_2.t1 48.0005
R4255 V_p_2.n6 V_p_2.t8 48.0005
R4256 V_p_2.t4 V_p_2.n6 48.0005
R4257 V_p_2.n0 V_p_2.n1 1.8755
R4258 START_UP_NFET1.t1 START_UP_NFET1.t0 178.194
R4259 V_CMFB_S1.n2 V_CMFB_S1.n0 344.837
R4260 V_CMFB_S1.n2 V_CMFB_S1.n1 344.274
R4261 V_CMFB_S1.n4 V_CMFB_S1.n3 292.5
R4262 V_CMFB_S1.n4 V_CMFB_S1.n2 52.3363
R4263 V_CMFB_S1 V_CMFB_S1.n4 52.1563
R4264 V_CMFB_S1.n3 V_CMFB_S1.t4 39.4005
R4265 V_CMFB_S1.n3 V_CMFB_S1.t1 39.4005
R4266 V_CMFB_S1.n1 V_CMFB_S1.t2 39.4005
R4267 V_CMFB_S1.n1 V_CMFB_S1.t0 39.4005
R4268 V_CMFB_S1.n0 V_CMFB_S1.t5 39.4005
R4269 V_CMFB_S1.n0 V_CMFB_S1.t3 39.4005
R4270 START_UP.n1 START_UP.t7 238.322
R4271 START_UP.n1 START_UP.t6 238.322
R4272 START_UP.n5 START_UP.n4 175.558
R4273 START_UP.n4 START_UP.n3 168.935
R4274 START_UP.n2 START_UP.n1 166.925
R4275 START_UP.n0 START_UP.t5 130.001
R4276 START_UP.n0 START_UP.t4 81.7084
R4277 START_UP.n2 START_UP.n0 50.4177
R4278 START_UP.n3 START_UP.t1 13.1338
R4279 START_UP.n3 START_UP.t2 13.1338
R4280 START_UP.t0 START_UP.n5 13.1338
R4281 START_UP.n5 START_UP.t3 13.1338
R4282 START_UP.n4 START_UP.n2 4.21925
R4283 Vin-.n7 Vin-.t11 688.859
R4284 Vin-.n9 Vin-.n8 514.134
R4285 Vin-.n6 Vin-.n5 351.522
R4286 Vin-.n11 Vin-.n10 213.4
R4287 Vin-.n7 Vin-.t8 174.726
R4288 Vin-.n8 Vin-.t9 174.726
R4289 Vin-.n9 Vin-.t12 174.726
R4290 Vin-.n10 Vin-.t10 174.726
R4291 Vin-.n4 Vin-.n2 173.029
R4292 Vin-.n4 Vin-.n3 168.654
R4293 Vin-.n8 Vin-.n7 128.534
R4294 Vin-.n10 Vin-.n9 128.534
R4295 Vin-.n12 Vin-.t0 119.099
R4296 Vin-.n1 Vin-.n0 83.5719
R4297 Vin-.n17 Vin-.n1 73.682
R4298 Vin-.n5 Vin-.t7 39.4005
R4299 Vin-.n5 Vin-.t6 39.4005
R4300 Vin-.n14 Vin-.t5 36.6632
R4301 Vin-.n13 Vin-.n12 28.813
R4302 Vin-.t5 Vin-.n1 25.7843
R4303 Vin-.n12 Vin-.n11 16.188
R4304 Vin-.n3 Vin-.t3 13.1338
R4305 Vin-.n3 Vin-.t4 13.1338
R4306 Vin-.n2 Vin-.t1 13.1338
R4307 Vin-.n2 Vin-.t2 13.1338
R4308 Vin-.n11 Vin-.n6 11.2193
R4309 Vin-.n6 Vin-.n4 3.8755
R4310 Vin-.n15 Vin-.n14 1.80777
R4311 Vin-.n16 Vin-.n15 1.5505
R4312 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter Vin-.n17 1.07742
R4313 Vin-.n14 Vin-.n13 1.04793
R4314 Vin-.n17 Vin-.n16 0.763532
R4315 Vin-.n15 Vin-.n0 0.590702
R4316 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter Vin-.n0 0.498483
R4317 Vin-.n16 Vin-.n13 0.0106786
R4318 V_TOP.n0 V_TOP.t14 369.534
R4319 V_TOP.n22 V_TOP.n20 339.961
R4320 V_TOP.n19 V_TOP.n18 339.272
R4321 V_TOP.n27 V_TOP.n26 339.272
R4322 V_TOP.n29 V_TOP.n28 339.272
R4323 V_TOP.n22 V_TOP.n21 339.272
R4324 V_TOP.n24 V_TOP.n23 334.772
R4325 V_TOP.n1 V_TOP.n0 224.934
R4326 V_TOP.n2 V_TOP.n1 224.934
R4327 V_TOP.n3 V_TOP.n2 224.934
R4328 V_TOP.n4 V_TOP.n3 224.934
R4329 V_TOP.n5 V_TOP.n4 224.934
R4330 V_TOP.n39 V_TOP.n38 224.934
R4331 V_TOP.n38 V_TOP.n37 224.934
R4332 V_TOP.n37 V_TOP.n36 224.934
R4333 V_TOP.n36 V_TOP.n35 224.934
R4334 V_TOP.n35 V_TOP.n34 224.934
R4335 V_TOP.n34 V_TOP.n33 224.934
R4336 V_TOP.n33 V_TOP.n32 224.934
R4337 V_TOP V_TOP.t27 214.222
R4338 V_TOP.n31 V_TOP.n30 163.175
R4339 V_TOP.n0 V_TOP.t41 144.601
R4340 V_TOP.n1 V_TOP.t37 144.601
R4341 V_TOP.n2 V_TOP.t30 144.601
R4342 V_TOP.n3 V_TOP.t25 144.601
R4343 V_TOP.n4 V_TOP.t15 144.601
R4344 V_TOP.n5 V_TOP.t43 144.601
R4345 V_TOP.n39 V_TOP.t31 144.601
R4346 V_TOP.n38 V_TOP.t38 144.601
R4347 V_TOP.n37 V_TOP.t42 144.601
R4348 V_TOP.n36 V_TOP.t45 144.601
R4349 V_TOP.n35 V_TOP.t19 144.601
R4350 V_TOP.n34 V_TOP.t28 144.601
R4351 V_TOP.n33 V_TOP.t34 144.601
R4352 V_TOP.n32 V_TOP.t40 144.601
R4353 V_TOP.n17 V_TOP.t0 108.424
R4354 V_TOP.n30 V_TOP.t1 95.447
R4355 V_TOP.n31 V_TOP.n5 69.6227
R4356 V_TOP V_TOP.n39 69.6227
R4357 V_TOP.n32 V_TOP.n31 69.6227
R4358 V_TOP.n18 V_TOP.t11 39.4005
R4359 V_TOP.n18 V_TOP.t4 39.4005
R4360 V_TOP.n23 V_TOP.t8 39.4005
R4361 V_TOP.n23 V_TOP.t10 39.4005
R4362 V_TOP.n21 V_TOP.t3 39.4005
R4363 V_TOP.n21 V_TOP.t13 39.4005
R4364 V_TOP.n20 V_TOP.t12 39.4005
R4365 V_TOP.n20 V_TOP.t2 39.4005
R4366 V_TOP.n26 V_TOP.t6 39.4005
R4367 V_TOP.n26 V_TOP.t9 39.4005
R4368 V_TOP.n28 V_TOP.t5 39.4005
R4369 V_TOP.n28 V_TOP.t7 39.4005
R4370 V_TOP.n17 V_TOP.n16 37.1479
R4371 V_TOP.n19 V_TOP.n17 27.8371
R4372 V_TOP.n24 V_TOP.n22 8.313
R4373 V_TOP.n30 V_TOP.n29 5.188
R4374 V_TOP.n7 V_TOP.t49 4.8295
R4375 V_TOP.n6 V_TOP.t24 4.8295
R4376 V_TOP.n9 V_TOP.t36 4.8295
R4377 V_TOP.n8 V_TOP.t18 4.8295
R4378 V_TOP.n11 V_TOP.t22 4.8295
R4379 V_TOP.n10 V_TOP.t46 4.8295
R4380 V_TOP.n13 V_TOP.t33 4.8295
R4381 V_TOP.n12 V_TOP.t16 4.8295
R4382 V_TOP.n14 V_TOP.t44 4.8295
R4383 V_TOP.n7 V_TOP.t47 4.5005
R4384 V_TOP.n6 V_TOP.t26 4.5005
R4385 V_TOP.n9 V_TOP.t35 4.5005
R4386 V_TOP.n8 V_TOP.t20 4.5005
R4387 V_TOP.n11 V_TOP.t21 4.5005
R4388 V_TOP.n10 V_TOP.t48 4.5005
R4389 V_TOP.n13 V_TOP.t32 4.5005
R4390 V_TOP.n12 V_TOP.t17 4.5005
R4391 V_TOP.n14 V_TOP.t29 4.5005
R4392 V_TOP.n15 V_TOP.t39 4.5005
R4393 V_TOP.n16 V_TOP.t23 4.5005
R4394 V_TOP.n25 V_TOP.n24 4.5005
R4395 V_TOP.n29 V_TOP.n27 2.1255
R4396 V_TOP.n27 V_TOP.n25 2.1255
R4397 V_TOP.n25 V_TOP.n19 2.1255
R4398 V_TOP.n7 V_TOP.n6 0.3295
R4399 V_TOP.n9 V_TOP.n8 0.3295
R4400 V_TOP.n11 V_TOP.n10 0.3295
R4401 V_TOP.n13 V_TOP.n12 0.3295
R4402 V_TOP.n15 V_TOP.n14 0.3295
R4403 V_TOP.n16 V_TOP.n15 0.3295
R4404 V_TOP.n9 V_TOP.n7 0.2825
R4405 V_TOP.n11 V_TOP.n9 0.2825
R4406 V_TOP.n13 V_TOP.n11 0.2825
R4407 V_TOP.n14 V_TOP.n13 0.2825
R4408 V_CMFB_S3.n2 V_CMFB_S3.n0 345.264
R4409 V_CMFB_S3.n2 V_CMFB_S3.n1 344.7
R4410 V_CMFB_S3.n4 V_CMFB_S3.n3 292.5
R4411 V_CMFB_S3.n4 V_CMFB_S3.n2 52.763
R4412 V_CMFB_S3 V_CMFB_S3.n4 51.7297
R4413 V_CMFB_S3.n3 V_CMFB_S3.t1 39.4005
R4414 V_CMFB_S3.n3 V_CMFB_S3.t5 39.4005
R4415 V_CMFB_S3.n1 V_CMFB_S3.t0 39.4005
R4416 V_CMFB_S3.n1 V_CMFB_S3.t2 39.4005
R4417 V_CMFB_S3.n0 V_CMFB_S3.t4 39.4005
R4418 V_CMFB_S3.n0 V_CMFB_S3.t3 39.4005
R4419 VB3_CUR_BIAS.n2 VB3_CUR_BIAS.n1 139.639
R4420 VB3_CUR_BIAS.n2 VB3_CUR_BIAS.n0 139.638
R4421 VB3_CUR_BIAS.n4 VB3_CUR_BIAS.n3 134.577
R4422 VB3_CUR_BIAS VB3_CUR_BIAS.n4 41.063
R4423 VB3_CUR_BIAS.n3 VB3_CUR_BIAS.t4 24.0005
R4424 VB3_CUR_BIAS.n3 VB3_CUR_BIAS.t2 24.0005
R4425 VB3_CUR_BIAS.n1 VB3_CUR_BIAS.t0 24.0005
R4426 VB3_CUR_BIAS.n1 VB3_CUR_BIAS.t3 24.0005
R4427 VB3_CUR_BIAS.n0 VB3_CUR_BIAS.t5 24.0005
R4428 VB3_CUR_BIAS.n0 VB3_CUR_BIAS.t1 24.0005
R4429 VB3_CUR_BIAS.n4 VB3_CUR_BIAS.n2 4.5005
R4430 V_mir1.n9 V_mir1.n5 325.473
R4431 V_mir1.n4 V_mir1.n0 325.471
R4432 V_mir1.n20 V_mir1.n19 325.471
R4433 V_mir1.n16 V_mir1.t20 310.488
R4434 V_mir1.n6 V_mir1.t19 310.488
R4435 V_mir1.n1 V_mir1.t22 310.488
R4436 V_mir1.n13 V_mir1.t13 278.312
R4437 V_mir1.n13 V_mir1.n12 228.939
R4438 V_mir1.n14 V_mir1.n11 224.439
R4439 V_mir1.n18 V_mir1.t0 184.097
R4440 V_mir1.n8 V_mir1.t4 184.097
R4441 V_mir1.n3 V_mir1.t8 184.097
R4442 V_mir1.n17 V_mir1.n16 167.094
R4443 V_mir1.n7 V_mir1.n6 167.094
R4444 V_mir1.n2 V_mir1.n1 167.094
R4445 V_mir1.n9 V_mir1.n8 152
R4446 V_mir1.n4 V_mir1.n3 152
R4447 V_mir1.n19 V_mir1.n18 152
R4448 V_mir1.n16 V_mir1.t18 120.501
R4449 V_mir1.n17 V_mir1.t10 120.501
R4450 V_mir1.n6 V_mir1.t17 120.501
R4451 V_mir1.n7 V_mir1.t2 120.501
R4452 V_mir1.n1 V_mir1.t21 120.501
R4453 V_mir1.n2 V_mir1.t6 120.501
R4454 V_mir1.n12 V_mir1.t16 48.0005
R4455 V_mir1.n12 V_mir1.t15 48.0005
R4456 V_mir1.n11 V_mir1.t12 48.0005
R4457 V_mir1.n11 V_mir1.t14 48.0005
R4458 V_mir1.n18 V_mir1.n17 40.7027
R4459 V_mir1.n8 V_mir1.n7 40.7027
R4460 V_mir1.n3 V_mir1.n2 40.7027
R4461 V_mir1.n5 V_mir1.t3 39.4005
R4462 V_mir1.n5 V_mir1.t5 39.4005
R4463 V_mir1.n0 V_mir1.t7 39.4005
R4464 V_mir1.n0 V_mir1.t9 39.4005
R4465 V_mir1.t11 V_mir1.n20 39.4005
R4466 V_mir1.n20 V_mir1.t1 39.4005
R4467 V_mir1.n10 V_mir1.n9 15.8005
R4468 V_mir1.n10 V_mir1.n4 15.8005
R4469 V_mir1.n19 V_mir1.n15 9.3005
R4470 V_mir1.n14 V_mir1.n13 5.8755
R4471 V_mir1.n15 V_mir1.n10 4.5005
R4472 V_mir1.n15 V_mir1.n14 0.78175
R4473 V_CUR_REF_REG.n4 V_CUR_REF_REG.n3 526.183
R4474 V_CUR_REF_REG.n2 V_CUR_REF_REG.n1 514.134
R4475 V_CUR_REF_REG.n5 V_CUR_REF_REG.n0 360.586
R4476 V_CUR_REF_REG.n1 V_CUR_REF_REG.t4 303.259
R4477 V_CUR_REF_REG.n5 V_CUR_REF_REG.n4 210.169
R4478 V_CUR_REF_REG.n1 V_CUR_REF_REG.t5 174.726
R4479 V_CUR_REF_REG.n2 V_CUR_REF_REG.t7 174.726
R4480 V_CUR_REF_REG.n3 V_CUR_REF_REG.t3 174.726
R4481 V_CUR_REF_REG.t0 V_CUR_REF_REG.n5 153.474
R4482 V_CUR_REF_REG.n3 V_CUR_REF_REG.n2 128.534
R4483 V_CUR_REF_REG.n4 V_CUR_REF_REG.t6 96.4005
R4484 V_CUR_REF_REG.n0 V_CUR_REF_REG.t1 39.4005
R4485 V_CUR_REF_REG.n0 V_CUR_REF_REG.t2 39.4005
R4486 a_32320_n7778.t0 a_32320_n7778.t1 178.133
R4487 PFET_GATE_10uA.n21 PFET_GATE_10uA.t14 369.534
R4488 PFET_GATE_10uA.n18 PFET_GATE_10uA.t20 369.534
R4489 PFET_GATE_10uA.n16 PFET_GATE_10uA.t28 369.534
R4490 PFET_GATE_10uA.n15 PFET_GATE_10uA.t21 369.534
R4491 PFET_GATE_10uA.n1 PFET_GATE_10uA.t27 369.534
R4492 PFET_GATE_10uA.n0 PFET_GATE_10uA.t13 369.534
R4493 PFET_GATE_10uA.n7 PFET_GATE_10uA.n5 341.397
R4494 PFET_GATE_10uA.n9 PFET_GATE_10uA.n8 339.272
R4495 PFET_GATE_10uA.n7 PFET_GATE_10uA.n6 339.272
R4496 PFET_GATE_10uA.n12 PFET_GATE_10uA.n11 334.772
R4497 PFET_GATE_10uA.n3 PFET_GATE_10uA.t11 238.322
R4498 PFET_GATE_10uA.n3 PFET_GATE_10uA.t23 238.322
R4499 PFET_GATE_10uA.n21 PFET_GATE_10uA.t19 192.8
R4500 PFET_GATE_10uA.n22 PFET_GATE_10uA.t29 192.8
R4501 PFET_GATE_10uA.n23 PFET_GATE_10uA.t18 192.8
R4502 PFET_GATE_10uA.n24 PFET_GATE_10uA.t26 192.8
R4503 PFET_GATE_10uA.n25 PFET_GATE_10uA.t15 192.8
R4504 PFET_GATE_10uA.n20 PFET_GATE_10uA.t24 192.8
R4505 PFET_GATE_10uA.n19 PFET_GATE_10uA.t12 192.8
R4506 PFET_GATE_10uA.n18 PFET_GATE_10uA.t22 192.8
R4507 PFET_GATE_10uA.n16 PFET_GATE_10uA.t17 192.8
R4508 PFET_GATE_10uA.n15 PFET_GATE_10uA.t10 192.8
R4509 PFET_GATE_10uA.n1 PFET_GATE_10uA.t16 192.8
R4510 PFET_GATE_10uA.n0 PFET_GATE_10uA.t25 192.8
R4511 PFET_GATE_10uA.n25 PFET_GATE_10uA.n24 176.733
R4512 PFET_GATE_10uA.n24 PFET_GATE_10uA.n23 176.733
R4513 PFET_GATE_10uA.n23 PFET_GATE_10uA.n22 176.733
R4514 PFET_GATE_10uA.n22 PFET_GATE_10uA.n21 176.733
R4515 PFET_GATE_10uA.n19 PFET_GATE_10uA.n18 176.733
R4516 PFET_GATE_10uA.n20 PFET_GATE_10uA.n19 176.733
R4517 PFET_GATE_10uA PFET_GATE_10uA.n17 171.321
R4518 PFET_GATE_10uA.n14 PFET_GATE_10uA.n2 168.166
R4519 PFET_GATE_10uA.n4 PFET_GATE_10uA.n3 167.519
R4520 PFET_GATE_10uA PFET_GATE_10uA.n26 166.071
R4521 PFET_GATE_10uA.n4 PFET_GATE_10uA.t0 137.48
R4522 PFET_GATE_10uA.n10 PFET_GATE_10uA.t1 100.635
R4523 PFET_GATE_10uA.n26 PFET_GATE_10uA.n25 56.2338
R4524 PFET_GATE_10uA.n26 PFET_GATE_10uA.n20 56.2338
R4525 PFET_GATE_10uA.n17 PFET_GATE_10uA.n16 56.2338
R4526 PFET_GATE_10uA.n17 PFET_GATE_10uA.n15 56.2338
R4527 PFET_GATE_10uA.n2 PFET_GATE_10uA.n1 56.2338
R4528 PFET_GATE_10uA.n2 PFET_GATE_10uA.n0 56.2338
R4529 PFET_GATE_10uA.n11 PFET_GATE_10uA.t5 39.4005
R4530 PFET_GATE_10uA.n11 PFET_GATE_10uA.t2 39.4005
R4531 PFET_GATE_10uA.n8 PFET_GATE_10uA.t8 39.4005
R4532 PFET_GATE_10uA.n8 PFET_GATE_10uA.t4 39.4005
R4533 PFET_GATE_10uA.n6 PFET_GATE_10uA.t6 39.4005
R4534 PFET_GATE_10uA.n6 PFET_GATE_10uA.t9 39.4005
R4535 PFET_GATE_10uA.n5 PFET_GATE_10uA.t3 39.4005
R4536 PFET_GATE_10uA.n5 PFET_GATE_10uA.t7 39.4005
R4537 PFET_GATE_10uA.n14 PFET_GATE_10uA.n13 27.5005
R4538 PFET_GATE_10uA.n13 PFET_GATE_10uA.n12 9.53175
R4539 PFET_GATE_10uA.n12 PFET_GATE_10uA.n10 4.5005
R4540 PFET_GATE_10uA PFET_GATE_10uA.n14 2.34425
R4541 PFET_GATE_10uA.n9 PFET_GATE_10uA.n7 2.1255
R4542 PFET_GATE_10uA.n10 PFET_GATE_10uA.n9 2.1255
R4543 PFET_GATE_10uA.n13 PFET_GATE_10uA.n4 1.688
R4544 VB1_CUR_BIAS.n2 VB1_CUR_BIAS.n0 339.961
R4545 VB1_CUR_BIAS.n2 VB1_CUR_BIAS.n1 339.272
R4546 VB1_CUR_BIAS.n1 VB1_CUR_BIAS.t3 39.4005
R4547 VB1_CUR_BIAS.n1 VB1_CUR_BIAS.t0 39.4005
R4548 VB1_CUR_BIAS.n0 VB1_CUR_BIAS.t1 39.4005
R4549 VB1_CUR_BIAS.n0 VB1_CUR_BIAS.t2 39.4005
R4550 VB1_CUR_BIAS VB1_CUR_BIAS.n2 12.1255
R4551 TAIL_CUR_MIR_BIAS.n4 TAIL_CUR_MIR_BIAS.n3 339.836
R4552 TAIL_CUR_MIR_BIAS.n2 TAIL_CUR_MIR_BIAS.n0 339.834
R4553 TAIL_CUR_MIR_BIAS.n2 TAIL_CUR_MIR_BIAS.n1 339.272
R4554 TAIL_CUR_MIR_BIAS.n6 TAIL_CUR_MIR_BIAS.n5 287.264
R4555 TAIL_CUR_MIR_BIAS.n6 TAIL_CUR_MIR_BIAS.n4 52.01
R4556 TAIL_CUR_MIR_BIAS TAIL_CUR_MIR_BIAS.n6 51.6642
R4557 TAIL_CUR_MIR_BIAS.n5 TAIL_CUR_MIR_BIAS.t1 39.4005
R4558 TAIL_CUR_MIR_BIAS.n5 TAIL_CUR_MIR_BIAS.t5 39.4005
R4559 TAIL_CUR_MIR_BIAS.n3 TAIL_CUR_MIR_BIAS.t0 39.4005
R4560 TAIL_CUR_MIR_BIAS.n3 TAIL_CUR_MIR_BIAS.t4 39.4005
R4561 TAIL_CUR_MIR_BIAS.n1 TAIL_CUR_MIR_BIAS.t2 39.4005
R4562 TAIL_CUR_MIR_BIAS.n1 TAIL_CUR_MIR_BIAS.t6 39.4005
R4563 TAIL_CUR_MIR_BIAS.n0 TAIL_CUR_MIR_BIAS.t3 39.4005
R4564 TAIL_CUR_MIR_BIAS.n0 TAIL_CUR_MIR_BIAS.t7 39.4005
R4565 TAIL_CUR_MIR_BIAS.n4 TAIL_CUR_MIR_BIAS.n2 0.563
R4566 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 195.608
R4567 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 83.5719
R4568 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 83.5719
R4569 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 83.5719
R4570 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 83.5719
R4571 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 83.5719
R4572 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 83.5719
R4573 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 83.5719
R4574 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 83.5719
R4575 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 83.5719
R4576 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 83.5719
R4577 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 83.5719
R4578 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 83.5719
R4579 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 83.5719
R4580 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 83.5719
R4581 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 83.5719
R4582 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 83.5719
R4583 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 83.5719
R4584 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 83.5719
R4585 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 83.5719
R4586 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R4587 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 73.682
R4588 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 73.682
R4589 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 73.3165
R4590 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 73.3165
R4591 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 73.3165
R4592 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 73.3165
R4593 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 73.3165
R4594 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 73.3165
R4595 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 73.19
R4596 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 73.19
R4597 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 73.19
R4598 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 73.19
R4599 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 73.19
R4600 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 73.19
R4601 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 36.6632
R4602 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 36.6632
R4603 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 26.074
R4604 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 26.074
R4605 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 26.074
R4606 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 26.074
R4607 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 26.074
R4608 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 26.074
R4609 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 25.7843
R4610 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 25.7843
R4611 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 25.7843
R4612 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 25.7843
R4613 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 25.7843
R4614 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 25.7843
R4615 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 25.7843
R4616 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 25.7843
R4617 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 9.3005
R4618 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 9.3005
R4619 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 9.3005
R4620 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 9.3005
R4621 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 9.3005
R4622 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 9.3005
R4623 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 9.3005
R4624 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 9.3005
R4625 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 9.3005
R4626 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 9.3005
R4627 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 9.3005
R4628 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 9.3005
R4629 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 9.3005
R4630 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 9.3005
R4631 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 9.3005
R4632 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 9.3005
R4633 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 9.3005
R4634 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 9.3005
R4635 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 9.3005
R4636 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R4637 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 9.3005
R4638 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 9.3005
R4639 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 9.3005
R4640 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 9.3005
R4641 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R4642 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 9.3005
R4643 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R4644 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R4645 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 9.3005
R4646 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 9.3005
R4647 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R4648 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R4649 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R4650 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 9.3005
R4651 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R4652 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 9.3005
R4653 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R4654 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R4655 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 9.3005
R4656 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 9.3005
R4657 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R4658 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R4659 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 9.3005
R4660 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R4661 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R4662 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R4663 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 9.3005
R4664 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 9.3005
R4665 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 9.3005
R4666 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R4667 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R4668 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 9.3005
R4669 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 9.3005
R4670 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 9.3005
R4671 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 4.64654
R4672 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 4.64654
R4673 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 4.64654
R4674 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 4.64654
R4675 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 4.64654
R4676 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 4.64654
R4677 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 4.64654
R4678 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 4.64654
R4679 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 4.64654
R4680 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 2.36206
R4681 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 2.36206
R4682 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 2.36206
R4683 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 2.36206
R4684 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 2.19742
R4685 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 2.19742
R4686 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 2.19742
R4687 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 2.19742
R4688 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 1.80777
R4689 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 1.80777
R4690 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 1.5505
R4691 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R4692 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 1.5505
R4693 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 1.5505
R4694 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 1.5505
R4695 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 1.5505
R4696 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 1.5505
R4697 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 1.5505
R4698 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 1.5505
R4699 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 1.5505
R4700 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 1.5505
R4701 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 1.5505
R4702 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 1.5505
R4703 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 1.5505
R4704 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 1.5505
R4705 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 1.5505
R4706 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 1.5505
R4707 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 1.5505
R4708 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 1.19225
R4709 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 1.19225
R4710 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 1.19225
R4711 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 1.19225
R4712 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 1.19225
R4713 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 1.19225
R4714 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 1.07742
R4715 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 1.07742
R4716 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 1.07024
R4717 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 1.07024
R4718 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 1.07024
R4719 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 1.07024
R4720 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 1.07024
R4721 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.07024
R4722 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.04793
R4723 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 1.04793
R4724 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 1.0237
R4725 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 1.0237
R4726 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 1.0237
R4727 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 1.0237
R4728 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 1.0237
R4729 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.0237
R4730 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 0.959578
R4731 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 0.959578
R4732 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.959578
R4733 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.959578
R4734 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 0.959578
R4735 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 0.959578
R4736 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 0.885803
R4737 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.885803
R4738 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 0.885803
R4739 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.885803
R4740 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 0.885803
R4741 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 0.885803
R4742 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 0.812055
R4743 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 0.812055
R4744 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 0.77514
R4745 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 0.77514
R4746 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 0.77514
R4747 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.77514
R4748 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.77514
R4749 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 0.77514
R4750 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 0.763532
R4751 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 0.763532
R4752 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.756696
R4753 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R4754 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R4755 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.756696
R4756 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R4757 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 0.756696
R4758 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.647417
R4759 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.647417
R4760 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 0.590702
R4761 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.590702
R4762 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 0.590702
R4763 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 0.590702
R4764 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 0.590702
R4765 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.590702
R4766 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 0.590702
R4767 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.590702
R4768 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.498483
R4769 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.498483
R4770 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 0.498483
R4771 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 0.498483
R4772 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.498483
R4773 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.498483
R4774 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.498483
R4775 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.498483
R4776 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 0.290206
R4777 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 0.290206
R4778 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 0.290206
R4779 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 0.290206
R4780 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.290206
R4781 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 0.290206
R4782 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 0.154071
R4783 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 0.154071
R4784 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 0.154071
R4785 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 0.154071
R4786 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 0.137464
R4787 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 0.137464
R4788 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 0.134964
R4789 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 0.134964
R4790 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R4791 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 0.0183571
R4792 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R4793 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R4794 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 0.0183571
R4795 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R4796 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R4797 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 0.0183571
R4798 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 0.0183571
R4799 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.0183571
R4800 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.0183571
R4801 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.0183571
R4802 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.0183571
R4803 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 0.0183571
R4804 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 0.0183571
R4805 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 0.0183571
R4806 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 0.0183571
R4807 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.0183571
R4808 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0106786
R4809 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 0.0106786
R4810 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 0.0106786
R4811 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 0.0106786
R4812 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 0.0106786
R4813 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 0.00992001
R4814 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 0.00992001
R4815 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 0.00992001
R4816 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 0.00992001
R4817 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 0.00992001
R4818 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 0.00992001
R4819 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 0.00992001
R4820 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 0.00992001
R4821 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 0.00992001
R4822 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 0.00992001
R4823 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 0.00992001
R4824 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R4825 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.00992001
R4826 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.00992001
R4827 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.00992001
R4828 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.00992001
R4829 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 0.00992001
R4830 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.00992001
R4831 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00817857
R4832 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00817857
R4833 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 0.00817857
R4834 a_38040_n7928.t0 a_38040_n7928.t1 178.133
R4835 ERR_AMP_CUR_BIAS ERR_AMP_CUR_BIAS.n0 175.172
R4836 ERR_AMP_CUR_BIAS.n0 ERR_AMP_CUR_BIAS.t1 24.0005
R4837 ERR_AMP_CUR_BIAS.n0 ERR_AMP_CUR_BIAS.t0 24.0005
R4838 a_32970_n7928.t0 a_32970_n7928.t1 178.133
R4839 a_32440_n6570.t0 a_32440_n6570.t1 178.133
R4840 a_33090_n6320.t0 a_33090_n6320.t1 178.133
R4841 a_37920_n6320.t0 a_37920_n6320.t1 178.133
C0 PFET_GATE_10uA VDDA 7.95837f
C1 1st_Vout_2 V_TOP 0.073737f
C2 PFET_GATE_10uA 1st_Vout_2 1.49161f
C3 PFET_GATE_10uA m2_36240_n160# 0.012f
C4 PFET_GATE_10uA V_CMFB_S3 0.35671f
C5 PFET_GATE_10uA V_CMFB_S1 0.215745f
C6 ERR_AMP_REF V_TOP 0.583702f
C7 PFET_GATE_10uA ERR_AMP_REF 1.67646f
C8 VB2_CUR_BIAS V_CMFB_S4 0.559002f
C9 PFET_GATE_10uA TAIL_CUR_MIR_BIAS 0.268567f
C10 PFET_GATE_10uA V_CMFB_S4 0.137571f
C11 PFET_GATE_10uA VB1_CUR_BIAS 0.254932f
C12 VDDA VB3_CUR_BIAS 0.183389f
C13 ERR_AMP_CUR_BIAS VB3_CUR_BIAS 0.051953f
C14 cap_res2 V_TOP 0.01893f
C15 VB3_CUR_BIAS 1st_Vout_2 0.042806f
C16 PFET_GATE_10uA cap_res2 0.012589f
C17 VB2_CUR_BIAS m1_35560_n3690# 0.08176f
C18 VB2_CUR_BIAS V_TOP 0.936691f
C19 VB3_CUR_BIAS ERR_AMP_REF 0.414647f
C20 PFET_GATE_10uA V_TOP 0.221314f
C21 VDDA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.046803f
C22 VB3_CUR_BIAS V_CMFB_S4 0.818388f
C23 V_CMFB_S2 VDDA 0.029799f
C24 V_CMFB_S2 ERR_AMP_CUR_BIAS 0.063017f
C25 ERR_AMP_CUR_BIAS VDDA 0.016199f
C26 VDDA 1st_Vout_2 1.51114f
C27 VDDA V_CMFB_S3 0.776564f
C28 VB3_CUR_BIAS m1_35560_n3690# 0.177673f
C29 VB2_CUR_BIAS VB3_CUR_BIAS 0.361534f
C30 1st_Vout_2 m2_36240_n160# 0.075543f
C31 VDDA V_CMFB_S1 0.776027f
C32 PFET_GATE_10uA VB3_CUR_BIAS 1.13473f
C33 VDDA ERR_AMP_REF 1.49115f
C34 1st_Vout_2 ERR_AMP_REF 0.670862f
C35 VDDA TAIL_CUR_MIR_BIAS 0.978678f
C36 VDDA V_CMFB_S4 0.23294f
C37 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter m1_35560_n3690# 0.013969f
C38 TAIL_CUR_MIR_BIAS V_CMFB_S3 0.018569f
C39 VDDA VB1_CUR_BIAS 0.616356f
C40 VB2_CUR_BIAS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.01158f
C41 V_CMFB_S4 1st_Vout_2 1.40961f
C42 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter V_TOP 0.055802f
C43 V_CMFB_S1 TAIL_CUR_MIR_BIAS 0.024906f
C44 V_CMFB_S3 VB1_CUR_BIAS 0.017903f
C45 VDDA cap_res2 1.06737f
C46 VB2_CUR_BIAS V_CMFB_S2 1.66154f
C47 cap_res2 1st_Vout_2 7.78906f
C48 m2_34880_n160# V_TOP 0.012f
C49 V_CMFB_S2 V_TOP 0.503779f
C50 V_CMFB_S4 ERR_AMP_REF 0.03827f
C51 ERR_AMP_REF VB1_CUR_BIAS 0.201706f
C52 VB2_CUR_BIAS VDDA 0.010405f
C53 ERR_AMP_CUR_BIAS m1_35560_n3690# 0.091711f
C54 VB2_CUR_BIAS ERR_AMP_CUR_BIAS 1.86165f
C55 VDDA V_TOP 13.237201f
C56 ERR_AMP_CUR_BIAS V_TOP 0.08195f
C57 V_CMFB_S4 GNDA 3.39226f
C58 VB3_CUR_BIAS GNDA 2.27736f
C59 ERR_AMP_CUR_BIAS GNDA 4.35357f
C60 V_CMFB_S2 GNDA 2.64383f
C61 VB2_CUR_BIAS GNDA 2.85457f
C62 VB1_CUR_BIAS GNDA 0.758311f
C63 ERR_AMP_REF GNDA 3.981564f
C64 V_CMFB_S3 GNDA 0.548687f
C65 TAIL_CUR_MIR_BIAS GNDA 0.571451f
C66 V_CMFB_S1 GNDA 0.590703f
C67 VDDA GNDA 73.76033f
C68 m2_36240_n160# GNDA 0.010002f $ **FLOATING
C69 m2_34880_n160# GNDA 0.0105f $ **FLOATING
C70 m1_35560_n3690# GNDA 0.259273f $ **FLOATING
C71 cap_res2 GNDA 6.744387f
C72 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA 17.895401f
C73 1st_Vout_2 GNDA 8.099878f
C74 V_TOP GNDA 9.96016f
C75 PFET_GATE_10uA GNDA 6.795063f
C76 ERR_AMP_CUR_BIAS.t1 GNDA 0.029966f
C77 ERR_AMP_CUR_BIAS.t0 GNDA 0.029966f
C78 ERR_AMP_CUR_BIAS.n0 GNDA 0.458302f
C79 PFET_GATE_10uA.t25 GNDA 0.020856f
C80 PFET_GATE_10uA.t13 GNDA 0.030831f
C81 PFET_GATE_10uA.n0 GNDA 0.033972f
C82 PFET_GATE_10uA.t16 GNDA 0.020856f
C83 PFET_GATE_10uA.t27 GNDA 0.030831f
C84 PFET_GATE_10uA.n1 GNDA 0.033972f
C85 PFET_GATE_10uA.n2 GNDA 0.034081f
C86 PFET_GATE_10uA.t0 GNDA 0.464967f
C87 PFET_GATE_10uA.t23 GNDA 0.024114f
C88 PFET_GATE_10uA.t11 GNDA 0.024114f
C89 PFET_GATE_10uA.n3 GNDA 0.069715f
C90 PFET_GATE_10uA.n4 GNDA 1.91969f
C91 PFET_GATE_10uA.t3 GNDA 0.021391f
C92 PFET_GATE_10uA.t7 GNDA 0.021391f
C93 PFET_GATE_10uA.n5 GNDA 0.054673f
C94 PFET_GATE_10uA.t6 GNDA 0.021391f
C95 PFET_GATE_10uA.t9 GNDA 0.021391f
C96 PFET_GATE_10uA.n6 GNDA 0.05326f
C97 PFET_GATE_10uA.n7 GNDA 0.520952f
C98 PFET_GATE_10uA.t8 GNDA 0.021391f
C99 PFET_GATE_10uA.t4 GNDA 0.021391f
C100 PFET_GATE_10uA.n8 GNDA 0.05326f
C101 PFET_GATE_10uA.n9 GNDA 0.295408f
C102 PFET_GATE_10uA.t1 GNDA 0.312465f
C103 PFET_GATE_10uA.n10 GNDA 0.603055f
C104 PFET_GATE_10uA.t5 GNDA 0.021391f
C105 PFET_GATE_10uA.t2 GNDA 0.021391f
C106 PFET_GATE_10uA.n11 GNDA 0.05159f
C107 PFET_GATE_10uA.n12 GNDA 0.27541f
C108 PFET_GATE_10uA.n13 GNDA 0.771508f
C109 PFET_GATE_10uA.n14 GNDA 0.759224f
C110 PFET_GATE_10uA.t10 GNDA 0.020856f
C111 PFET_GATE_10uA.t21 GNDA 0.030831f
C112 PFET_GATE_10uA.n15 GNDA 0.033972f
C113 PFET_GATE_10uA.t17 GNDA 0.020856f
C114 PFET_GATE_10uA.t28 GNDA 0.030831f
C115 PFET_GATE_10uA.n16 GNDA 0.033972f
C116 PFET_GATE_10uA.n17 GNDA 0.040878f
C117 PFET_GATE_10uA.t24 GNDA 0.020856f
C118 PFET_GATE_10uA.t12 GNDA 0.020856f
C119 PFET_GATE_10uA.t22 GNDA 0.020856f
C120 PFET_GATE_10uA.t20 GNDA 0.030831f
C121 PFET_GATE_10uA.n18 GNDA 0.038154f
C122 PFET_GATE_10uA.n19 GNDA 0.027273f
C123 PFET_GATE_10uA.n20 GNDA 0.023091f
C124 PFET_GATE_10uA.t15 GNDA 0.020856f
C125 PFET_GATE_10uA.t26 GNDA 0.020856f
C126 PFET_GATE_10uA.t18 GNDA 0.020856f
C127 PFET_GATE_10uA.t29 GNDA 0.020856f
C128 PFET_GATE_10uA.t19 GNDA 0.020856f
C129 PFET_GATE_10uA.t14 GNDA 0.030831f
C130 PFET_GATE_10uA.n21 GNDA 0.038154f
C131 PFET_GATE_10uA.n22 GNDA 0.027273f
C132 PFET_GATE_10uA.n23 GNDA 0.027273f
C133 PFET_GATE_10uA.n24 GNDA 0.027273f
C134 PFET_GATE_10uA.n25 GNDA 0.023091f
C135 PFET_GATE_10uA.n26 GNDA 0.031695f
C136 V_mir1.t1 GNDA 0.019293f
C137 V_mir1.t7 GNDA 0.019293f
C138 V_mir1.t9 GNDA 0.019293f
C139 V_mir1.n0 GNDA 0.044166f
C140 V_mir1.t6 GNDA 0.023151f
C141 V_mir1.t21 GNDA 0.023151f
C142 V_mir1.t22 GNDA 0.037369f
C143 V_mir1.n1 GNDA 0.041731f
C144 V_mir1.n2 GNDA 0.028507f
C145 V_mir1.t8 GNDA 0.02939f
C146 V_mir1.n3 GNDA 0.044354f
C147 V_mir1.n4 GNDA 0.109943f
C148 V_mir1.t3 GNDA 0.019293f
C149 V_mir1.t5 GNDA 0.019293f
C150 V_mir1.n5 GNDA 0.044166f
C151 V_mir1.t2 GNDA 0.023151f
C152 V_mir1.t17 GNDA 0.023151f
C153 V_mir1.t19 GNDA 0.037369f
C154 V_mir1.n6 GNDA 0.041731f
C155 V_mir1.n7 GNDA 0.028507f
C156 V_mir1.t4 GNDA 0.02939f
C157 V_mir1.n8 GNDA 0.044354f
C158 V_mir1.n9 GNDA 0.111042f
C159 V_mir1.n10 GNDA 0.381359f
C160 V_mir1.n11 GNDA 0.025223f
C161 V_mir1.t13 GNDA 0.041163f
C162 V_mir1.n12 GNDA 0.027381f
C163 V_mir1.n13 GNDA 0.451535f
C164 V_mir1.n14 GNDA 0.146338f
C165 V_mir1.n15 GNDA 0.051125f
C166 V_mir1.t10 GNDA 0.023151f
C167 V_mir1.t18 GNDA 0.023151f
C168 V_mir1.t20 GNDA 0.037369f
C169 V_mir1.n16 GNDA 0.041731f
C170 V_mir1.n17 GNDA 0.028507f
C171 V_mir1.t0 GNDA 0.02939f
C172 V_mir1.n18 GNDA 0.044354f
C173 V_mir1.n19 GNDA 0.085095f
C174 V_mir1.n20 GNDA 0.044166f
C175 V_mir1.t11 GNDA 0.019293f
C176 V_TOP.t27 GNDA 0.109989f
C177 V_TOP.t31 GNDA 0.095448f
C178 V_TOP.t38 GNDA 0.095448f
C179 V_TOP.t42 GNDA 0.095448f
C180 V_TOP.t45 GNDA 0.095448f
C181 V_TOP.t19 GNDA 0.095448f
C182 V_TOP.t28 GNDA 0.095448f
C183 V_TOP.t34 GNDA 0.095448f
C184 V_TOP.t40 GNDA 0.095448f
C185 V_TOP.t43 GNDA 0.095448f
C186 V_TOP.t15 GNDA 0.095448f
C187 V_TOP.t25 GNDA 0.095448f
C188 V_TOP.t30 GNDA 0.095448f
C189 V_TOP.t37 GNDA 0.095448f
C190 V_TOP.t41 GNDA 0.095448f
C191 V_TOP.t14 GNDA 0.124774f
C192 V_TOP.n0 GNDA 0.069758f
C193 V_TOP.n1 GNDA 0.050905f
C194 V_TOP.n2 GNDA 0.050905f
C195 V_TOP.n3 GNDA 0.050905f
C196 V_TOP.n4 GNDA 0.050905f
C197 V_TOP.n5 GNDA 0.04747f
C198 V_TOP.t1 GNDA 0.122745f
C199 V_TOP.t49 GNDA 0.369803f
C200 V_TOP.t47 GNDA 0.36361f
C201 V_TOP.t24 GNDA 0.369803f
C202 V_TOP.t26 GNDA 0.36361f
C203 V_TOP.n6 GNDA 0.243789f
C204 V_TOP.n7 GNDA 0.311966f
C205 V_TOP.t36 GNDA 0.369803f
C206 V_TOP.t35 GNDA 0.36361f
C207 V_TOP.t18 GNDA 0.369803f
C208 V_TOP.t20 GNDA 0.36361f
C209 V_TOP.n8 GNDA 0.243789f
C210 V_TOP.n9 GNDA 0.380143f
C211 V_TOP.t22 GNDA 0.369803f
C212 V_TOP.t21 GNDA 0.36361f
C213 V_TOP.t46 GNDA 0.369803f
C214 V_TOP.t48 GNDA 0.36361f
C215 V_TOP.n10 GNDA 0.243789f
C216 V_TOP.n11 GNDA 0.380143f
C217 V_TOP.t33 GNDA 0.369803f
C218 V_TOP.t32 GNDA 0.36361f
C219 V_TOP.t16 GNDA 0.369803f
C220 V_TOP.t17 GNDA 0.36361f
C221 V_TOP.n12 GNDA 0.243789f
C222 V_TOP.n13 GNDA 0.380143f
C223 V_TOP.t44 GNDA 0.369803f
C224 V_TOP.t29 GNDA 0.36361f
C225 V_TOP.n14 GNDA 0.311966f
C226 V_TOP.t39 GNDA 0.36361f
C227 V_TOP.n15 GNDA 0.159079f
C228 V_TOP.t23 GNDA 0.36361f
C229 V_TOP.n16 GNDA 0.544408f
C230 V_TOP.t0 GNDA 0.102288f
C231 V_TOP.n17 GNDA 0.724299f
C232 V_TOP.n18 GNDA 0.022634f
C233 V_TOP.n19 GNDA 0.414649f
C234 V_TOP.n20 GNDA 0.022786f
C235 V_TOP.n21 GNDA 0.022634f
C236 V_TOP.n22 GNDA 0.209756f
C237 V_TOP.n23 GNDA 0.021924f
C238 V_TOP.n24 GNDA 0.127416f
C239 V_TOP.n25 GNDA 0.072722f
C240 V_TOP.n26 GNDA 0.022634f
C241 V_TOP.n27 GNDA 0.125537f
C242 V_TOP.n28 GNDA 0.022634f
C243 V_TOP.n29 GNDA 0.124344f
C244 V_TOP.n30 GNDA 0.273328f
C245 V_TOP.n31 GNDA 0.019234f
C246 V_TOP.n32 GNDA 0.04747f
C247 V_TOP.n33 GNDA 0.050905f
C248 V_TOP.n34 GNDA 0.050905f
C249 V_TOP.n35 GNDA 0.050905f
C250 V_TOP.n36 GNDA 0.050905f
C251 V_TOP.n37 GNDA 0.050905f
C252 V_TOP.n38 GNDA 0.050905f
C253 V_TOP.n39 GNDA 0.04747f
C254 Vin-.n0 GNDA 0.046236f
C255 Vin-.n1 GNDA 0.316004f
C256 Vin-.t1 GNDA 0.027101f
C257 Vin-.t2 GNDA 0.027101f
C258 Vin-.n2 GNDA 0.094346f
C259 Vin-.t3 GNDA 0.027101f
C260 Vin-.t4 GNDA 0.027101f
C261 Vin-.n3 GNDA 0.090091f
C262 Vin-.n4 GNDA 0.386489f
C263 Vin-.n5 GNDA 0.027681f
C264 Vin-.n6 GNDA 0.366254f
C265 Vin-.t11 GNDA 0.022346f
C266 Vin-.n7 GNDA 0.026209f
C267 Vin-.n8 GNDA 0.021455f
C268 Vin-.n9 GNDA 0.021455f
C269 Vin-.n10 GNDA 0.036491f
C270 Vin-.n11 GNDA 0.497932f
C271 Vin-.t0 GNDA 0.117924f
C272 Vin-.n12 GNDA 0.65583f
C273 Vin-.n13 GNDA 1.33843f
C274 Vin-.t5 GNDA 0.32907f
C275 Vin-.n14 GNDA 0.294079f
C276 Vin-.n15 GNDA 0.122514f
C277 Vin-.n16 GNDA 0.578948f
C278 Vin-.n17 GNDA 0.368244f
C279 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter GNDA 0.082077f
C280 START_UP.t3 GNDA 0.026778f
C281 START_UP.t4 GNDA 1.06745f
C282 START_UP.t5 GNDA 0.02806f
C283 START_UP.n0 GNDA 0.801406f
C284 START_UP.t6 GNDA 0.010062f
C285 START_UP.t7 GNDA 0.010062f
C286 START_UP.n1 GNDA 0.028407f
C287 START_UP.n2 GNDA 0.498066f
C288 START_UP.t1 GNDA 0.026778f
C289 START_UP.t2 GNDA 0.026778f
C290 START_UP.n3 GNDA 0.08937f
C291 START_UP.n4 GNDA 0.462855f
C292 START_UP.n5 GNDA 0.097147f
C293 START_UP.t0 GNDA 0.026778f
C294 ERR_AMP_REF.t2 GNDA 0.145472f
C295 ERR_AMP_REF.t8 GNDA 0.022696f
C296 ERR_AMP_REF.n0 GNDA 0.02662f
C297 ERR_AMP_REF.n1 GNDA 0.021791f
C298 ERR_AMP_REF.n2 GNDA 0.021791f
C299 ERR_AMP_REF.n3 GNDA 0.037771f
C300 ERR_AMP_REF.n4 GNDA 0.757207f
C301 ERR_AMP_REF.t6 GNDA 0.027525f
C302 ERR_AMP_REF.t4 GNDA 0.027525f
C303 ERR_AMP_REF.n5 GNDA 0.096943f
C304 ERR_AMP_REF.t1 GNDA 0.027525f
C305 ERR_AMP_REF.t0 GNDA 0.027525f
C306 ERR_AMP_REF.n6 GNDA 0.092238f
C307 ERR_AMP_REF.n7 GNDA 0.431057f
C308 ERR_AMP_REF.t3 GNDA 0.027525f
C309 ERR_AMP_REF.t5 GNDA 0.027525f
C310 ERR_AMP_REF.n8 GNDA 0.092238f
C311 ERR_AMP_REF.n9 GNDA 0.308239f
C312 ERR_AMP_REF.n10 GNDA 0.226163f
C313 Vin+.t8 GNDA 0.010696f
C314 Vin+.t9 GNDA 0.025367f
C315 Vin+.t7 GNDA 0.01649f
C316 Vin+.n0 GNDA 0.054406f
C317 Vin+.t6 GNDA 0.01649f
C318 Vin+.n1 GNDA 0.042338f
C319 Vin+.t10 GNDA 0.01649f
C320 Vin+.n2 GNDA 0.042909f
C321 Vin+.n3 GNDA 0.130793f
C322 Vin+.t4 GNDA 0.05348f
C323 Vin+.t3 GNDA 0.05348f
C324 Vin+.n4 GNDA 0.176679f
C325 Vin+.n5 GNDA 1.27851f
C326 Vin+.t2 GNDA 0.05348f
C327 Vin+.t5 GNDA 0.05348f
C328 Vin+.n6 GNDA 0.17668f
C329 Vin+.n7 GNDA 1.06525f
C330 Vin+.t1 GNDA 0.232527f
C331 Vin+.n8 GNDA 1.7265f
C332 Vin+.t0 GNDA 0.173951f
C333 cap_res1.t14 GNDA 0.349187f
C334 cap_res1.t1 GNDA 0.350452f
C335 cap_res1.t4 GNDA 0.331712f
C336 cap_res1.t16 GNDA 0.349187f
C337 cap_res1.t17 GNDA 0.350452f
C338 cap_res1.t8 GNDA 0.331712f
C339 cap_res1.t2 GNDA 0.349187f
C340 cap_res1.t3 GNDA 0.350452f
C341 cap_res1.t12 GNDA 0.331712f
C342 cap_res1.t13 GNDA 0.349187f
C343 cap_res1.t15 GNDA 0.350452f
C344 cap_res1.t6 GNDA 0.331712f
C345 cap_res1.t9 GNDA 0.349187f
C346 cap_res1.t11 GNDA 0.350452f
C347 cap_res1.t20 GNDA 0.331712f
C348 cap_res1.n0 GNDA 0.23406f
C349 cap_res1.t19 GNDA 0.186395f
C350 cap_res1.n1 GNDA 0.253961f
C351 cap_res1.t5 GNDA 0.186395f
C352 cap_res1.n2 GNDA 0.253961f
C353 cap_res1.t10 GNDA 0.186395f
C354 cap_res1.n3 GNDA 0.253961f
C355 cap_res1.t7 GNDA 0.186395f
C356 cap_res1.n4 GNDA 0.253961f
C357 cap_res1.t18 GNDA 0.363549f
C358 cap_res1.t0 GNDA 0.08421f
C359 1st_Vout_1.n0 GNDA 0.715456f
C360 1st_Vout_1.n1 GNDA 0.308472f
C361 1st_Vout_1.n2 GNDA 1.74831f
C362 1st_Vout_1.n3 GNDA 0.127561f
C363 1st_Vout_1.n4 GNDA 1.79885f
C364 1st_Vout_1.t32 GNDA 0.021148f
C365 1st_Vout_1.t17 GNDA 0.35246f
C366 1st_Vout_1.t23 GNDA 0.358463f
C367 1st_Vout_1.t21 GNDA 0.35246f
C368 1st_Vout_1.t12 GNDA 0.35246f
C369 1st_Vout_1.t11 GNDA 0.358463f
C370 1st_Vout_1.t18 GNDA 0.358463f
C371 1st_Vout_1.t16 GNDA 0.35246f
C372 1st_Vout_1.t29 GNDA 0.35246f
C373 1st_Vout_1.t27 GNDA 0.358463f
C374 1st_Vout_1.t34 GNDA 0.358463f
C375 1st_Vout_1.t33 GNDA 0.35246f
C376 1st_Vout_1.t22 GNDA 0.35246f
C377 1st_Vout_1.t20 GNDA 0.358463f
C378 1st_Vout_1.t15 GNDA 0.358463f
C379 1st_Vout_1.t14 GNDA 0.35246f
C380 1st_Vout_1.t26 GNDA 0.35246f
C381 1st_Vout_1.t25 GNDA 0.358463f
C382 1st_Vout_1.t31 GNDA 0.358463f
C383 1st_Vout_1.t13 GNDA 0.35246f
C384 1st_Vout_1.t35 GNDA 0.35246f
C385 1st_Vout_1.t19 GNDA 0.023025f
C386 1st_Vout_1.n5 GNDA 0.022212f
C387 1st_Vout_1.t30 GNDA 0.013423f
C388 1st_Vout_1.t24 GNDA 0.013423f
C389 1st_Vout_1.n6 GNDA 0.029862f
C390 1st_Vout_1.n7 GNDA 0.021291f
C391 1st_Vout_1.n8 GNDA 0.012728f
C392 1st_Vout_1.t10 GNDA 0.018559f
C393 1st_Vout_1.n9 GNDA 0.192525f
C394 1st_Vout_1.n10 GNDA 0.011517f
C395 1st_Vout_1.t36 GNDA 0.013423f
C396 1st_Vout_1.t28 GNDA 0.013423f
C397 1st_Vout_1.n11 GNDA 0.029862f
C398 1st_Vout_1.n12 GNDA 0.168997f
C399 1st_Vout_1.n13 GNDA 0.022212f
C400 VDDA.n1 GNDA 0.034117f
C401 VDDA.t145 GNDA 0.014126f
C402 VDDA.n3 GNDA 0.034117f
C403 VDDA.n5 GNDA 0.034135f
C404 VDDA.n7 GNDA 0.034135f
C405 VDDA.n9 GNDA 0.034135f
C406 VDDA.n11 GNDA 0.034135f
C407 VDDA.n13 GNDA 0.034135f
C408 VDDA.n15 GNDA 0.034113f
C409 VDDA.t178 GNDA 0.014133f
C410 VDDA.n17 GNDA 0.046689f
C411 VDDA.n18 GNDA 0.016205f
C412 VDDA.t163 GNDA 0.014133f
C413 VDDA.n19 GNDA 0.040331f
C414 VDDA.t162 GNDA 0.042504f
C415 VDDA.t190 GNDA 0.029834f
C416 VDDA.t28 GNDA 0.029834f
C417 VDDA.t91 GNDA 0.029834f
C418 VDDA.t63 GNDA 0.029834f
C419 VDDA.t177 GNDA 0.042504f
C420 VDDA.n20 GNDA 0.040331f
C421 VDDA.n21 GNDA 0.015935f
C422 VDDA.n22 GNDA 0.02355f
C423 VDDA.n23 GNDA 0.02355f
C424 VDDA.n24 GNDA 0.015075f
C425 VDDA.t160 GNDA 0.013543f
C426 VDDA.n25 GNDA 0.04143f
C427 VDDA.t159 GNDA 0.042612f
C428 VDDA.t192 GNDA 0.029834f
C429 VDDA.t73 GNDA 0.029834f
C430 VDDA.t46 GNDA 0.029834f
C431 VDDA.t23 GNDA 0.029834f
C432 VDDA.t67 GNDA 0.029834f
C433 VDDA.t48 GNDA 0.029834f
C434 VDDA.t61 GNDA 0.029834f
C435 VDDA.t30 GNDA 0.029834f
C436 VDDA.t89 GNDA 0.029834f
C437 VDDA.t200 GNDA 0.029834f
C438 VDDA.t135 GNDA 0.042612f
C439 VDDA.t136 GNDA 0.013543f
C440 VDDA.n26 GNDA 0.04143f
C441 VDDA.n27 GNDA 0.015075f
C442 VDDA.n28 GNDA 0.02355f
C443 VDDA.n29 GNDA 0.02355f
C444 VDDA.n30 GNDA 0.015693f
C445 VDDA.t175 GNDA 0.014126f
C446 VDDA.n31 GNDA 0.040338f
C447 VDDA.t174 GNDA 0.042504f
C448 VDDA.t39 GNDA 0.029834f
C449 VDDA.t65 GNDA 0.029834f
C450 VDDA.t17 GNDA 0.029834f
C451 VDDA.t99 GNDA 0.029834f
C452 VDDA.t144 GNDA 0.042504f
C453 VDDA.n32 GNDA 0.040338f
C454 VDDA.n33 GNDA 0.015693f
C455 VDDA.n34 GNDA 0.07835f
C456 VDDA.n35 GNDA 1.68458f
C457 VDDA.t183 GNDA 0.205746f
C458 VDDA.t20 GNDA 0.216585f
C459 VDDA.t71 GNDA 0.217369f
C460 VDDA.t0 GNDA 0.205746f
C461 VDDA.t58 GNDA 0.216585f
C462 VDDA.t12 GNDA 0.217369f
C463 VDDA.t26 GNDA 0.205746f
C464 VDDA.t55 GNDA 0.216585f
C465 VDDA.t19 GNDA 0.217369f
C466 VDDA.t69 GNDA 0.205746f
C467 VDDA.t27 GNDA 0.216585f
C468 VDDA.t72 GNDA 0.217369f
C469 VDDA.t70 GNDA 0.205746f
C470 VDDA.t199 GNDA 0.216585f
C471 VDDA.t50 GNDA 0.217369f
C472 VDDA.n36 GNDA 0.145177f
C473 VDDA.t25 GNDA 0.115612f
C474 VDDA.n37 GNDA 0.15752f
C475 VDDA.t16 GNDA 0.115612f
C476 VDDA.n38 GNDA 0.15752f
C477 VDDA.t43 GNDA 0.115612f
C478 VDDA.n39 GNDA 0.15752f
C479 VDDA.t7 GNDA 0.115612f
C480 VDDA.n40 GNDA 0.15752f
C481 VDDA.t198 GNDA 0.202533f
C482 VDDA.n41 GNDA 2.08495f
C483 VDDA.t214 GNDA 0.428342f
C484 VDDA.t217 GNDA 0.439174f
C485 VDDA.t216 GNDA 0.456352f
C486 VDDA.n42 GNDA 0.305709f
C487 VDDA.t215 GNDA 0.45653f
C488 VDDA.n43 GNDA 0.150128f
C489 VDDA.n44 GNDA 0.218222f
C490 VDDA.n45 GNDA 0.398338f
C491 VDDA.n47 GNDA 0.039461f
C492 VDDA.n48 GNDA 0.016386f
C493 VDDA.t151 GNDA 0.013477f
C494 VDDA.n50 GNDA 0.025833f
C495 VDDA.t140 GNDA 0.014303f
C496 VDDA.n52 GNDA 0.039461f
C497 VDDA.n54 GNDA 0.039461f
C498 VDDA.n56 GNDA 0.039461f
C499 VDDA.n58 GNDA 0.039461f
C500 VDDA.n60 GNDA 0.039461f
C501 VDDA.n62 GNDA 0.039461f
C502 VDDA.n64 GNDA 0.039461f
C503 VDDA.n66 GNDA 0.039461f
C504 VDDA.n68 GNDA 0.039461f
C505 VDDA.n69 GNDA 0.025833f
C506 VDDA.t155 GNDA 0.014303f
C507 VDDA.n71 GNDA 0.039461f
C508 VDDA.n73 GNDA 0.039461f
C509 VDDA.n75 GNDA 0.039461f
C510 VDDA.n77 GNDA 0.039461f
C511 VDDA.n79 GNDA 0.039461f
C512 VDDA.n81 GNDA 0.039461f
C513 VDDA.n83 GNDA 0.039461f
C514 VDDA.n85 GNDA 0.056708f
C515 VDDA.n86 GNDA 0.015024f
C516 VDDA.t157 GNDA 0.013477f
C517 VDDA.n88 GNDA 0.016386f
C518 VDDA.n89 GNDA 0.047759f
C519 VDDA.t156 GNDA 0.040209f
C520 VDDA.t14 GNDA 0.032546f
C521 VDDA.t97 GNDA 0.032546f
C522 VDDA.t87 GNDA 0.032546f
C523 VDDA.t59 GNDA 0.032546f
C524 VDDA.t37 GNDA 0.032546f
C525 VDDA.t53 GNDA 0.032546f
C526 VDDA.t77 GNDA 0.032546f
C527 VDDA.t105 GNDA 0.032546f
C528 VDDA.t188 GNDA 0.032546f
C529 VDDA.t103 GNDA 0.032546f
C530 VDDA.t83 GNDA 0.032546f
C531 VDDA.t179 GNDA 0.032546f
C532 VDDA.t194 GNDA 0.032546f
C533 VDDA.t35 GNDA 0.032546f
C534 VDDA.t5 GNDA 0.032546f
C535 VDDA.t8 GNDA 0.032546f
C536 VDDA.t101 GNDA 0.032546f
C537 VDDA.t196 GNDA 0.032546f
C538 VDDA.t165 GNDA 0.049644f
C539 VDDA.t166 GNDA 0.013571f
C540 VDDA.n90 GNDA 0.070687f
C541 VDDA.n91 GNDA 0.01585f
C542 VDDA.n92 GNDA 0.028862f
C543 VDDA.n93 GNDA 0.028862f
C544 VDDA.n94 GNDA 0.014258f
C545 VDDA.t142 GNDA 0.013477f
C546 VDDA.n96 GNDA 0.016386f
C547 VDDA.n97 GNDA 0.047759f
C548 VDDA.t141 GNDA 0.040209f
C549 VDDA.t204 GNDA 0.032546f
C550 VDDA.t127 GNDA 0.032546f
C551 VDDA.t123 GNDA 0.032546f
C552 VDDA.t119 GNDA 0.032546f
C553 VDDA.t111 GNDA 0.032546f
C554 VDDA.t202 GNDA 0.032546f
C555 VDDA.t210 GNDA 0.032546f
C556 VDDA.t117 GNDA 0.032546f
C557 VDDA.t121 GNDA 0.032546f
C558 VDDA.t115 GNDA 0.032546f
C559 VDDA.t109 GNDA 0.032546f
C560 VDDA.t212 GNDA 0.032546f
C561 VDDA.t206 GNDA 0.032546f
C562 VDDA.t113 GNDA 0.032546f
C563 VDDA.t107 GNDA 0.032546f
C564 VDDA.t129 GNDA 0.032546f
C565 VDDA.t125 GNDA 0.032546f
C566 VDDA.t208 GNDA 0.032546f
C567 VDDA.t150 GNDA 0.040209f
C568 VDDA.n98 GNDA 0.047759f
C569 VDDA.n99 GNDA 0.025937f
C570 VDDA.t149 GNDA 0.014295f
C571 VDDA.n100 GNDA 0.014258f
C572 VDDA.n101 GNDA 0.066888f
C573 VDDA.n102 GNDA 0.128965f
C574 VDDA.t182 GNDA 0.011623f
C575 VDDA.t11 GNDA 0.011623f
C576 VDDA.n103 GNDA 0.0384f
C577 VDDA.n104 GNDA 0.049551f
C578 VDDA.t167 GNDA 0.055426f
C579 VDDA.t96 GNDA 0.011623f
C580 VDDA.t33 GNDA 0.011623f
C581 VDDA.n113 GNDA 0.0384f
C582 VDDA.n114 GNDA 0.049551f
C583 VDDA.t42 GNDA 0.011623f
C584 VDDA.t22 GNDA 0.011623f
C585 VDDA.n115 GNDA 0.0384f
C586 VDDA.n116 GNDA 0.049551f
C587 VDDA.t185 GNDA 0.011623f
C588 VDDA.t4 GNDA 0.011623f
C589 VDDA.n117 GNDA 0.0384f
C590 VDDA.n118 GNDA 0.049551f
C591 VDDA.t2 GNDA 0.011623f
C592 VDDA.t82 GNDA 0.011623f
C593 VDDA.n119 GNDA 0.0384f
C594 VDDA.n120 GNDA 0.049551f
C595 VDDA.t45 GNDA 0.011623f
C596 VDDA.t52 GNDA 0.011623f
C597 VDDA.n121 GNDA 0.0384f
C598 VDDA.n122 GNDA 0.049551f
C599 VDDA.t57 GNDA 0.011623f
C600 VDDA.t80 GNDA 0.011623f
C601 VDDA.n123 GNDA 0.0384f
C602 VDDA.n124 GNDA 0.049551f
C603 VDDA.t94 GNDA 0.011623f
C604 VDDA.t187 GNDA 0.011623f
C605 VDDA.n125 GNDA 0.0384f
C606 VDDA.n126 GNDA 0.049551f
C607 VDDA.n127 GNDA 0.019033f
C608 VDDA.t139 GNDA 0.013571f
C609 VDDA.n128 GNDA 0.067892f
C610 VDDA.t138 GNDA 0.047014f
C611 VDDA.t13 GNDA 0.029834f
C612 VDDA.t34 GNDA 0.029834f
C613 VDDA.t153 GNDA 0.048049f
C614 VDDA.t154 GNDA 0.015469f
C615 VDDA.n129 GNDA 0.071105f
C616 VDDA.n130 GNDA 0.018888f
C617 VDDA.n131 GNDA 0.056819f
C618 VDDA.n132 GNDA 0.026456f
C619 VDDA.n133 GNDA 0.0207f
C620 VDDA.n134 GNDA 0.013561f
C621 VDDA.n135 GNDA 0.013479f
C622 VDDA.n136 GNDA 0.019629f
C623 VDDA.n138 GNDA 0.013561f
C624 VDDA.n139 GNDA 0.013561f
C625 VDDA.n142 GNDA 0.013561f
C626 VDDA.n143 GNDA 0.013479f
C627 VDDA.n145 GNDA 0.015368f
C628 VDDA.n147 GNDA 0.10868f
C629 VDDA.t168 GNDA 0.115266f
C630 VDDA.t186 GNDA 0.11856f
C631 VDDA.t93 GNDA 0.11856f
C632 VDDA.t79 GNDA 0.11856f
C633 VDDA.t56 GNDA 0.11856f
C634 VDDA.t51 GNDA 0.11856f
C635 VDDA.t44 GNDA 0.11856f
C636 VDDA.t81 GNDA 0.11856f
C637 VDDA.t1 GNDA 0.11856f
C638 VDDA.t3 GNDA 0.11856f
C639 VDDA.t184 GNDA 0.11856f
C640 VDDA.t21 GNDA 0.11856f
C641 VDDA.t41 GNDA 0.11856f
C642 VDDA.t32 GNDA 0.11856f
C643 VDDA.t95 GNDA 0.11856f
C644 VDDA.t10 GNDA 0.11856f
C645 VDDA.t181 GNDA 0.11856f
C646 VDDA.t132 GNDA 0.115266f
C647 VDDA.n149 GNDA 0.013561f
C648 VDDA.n150 GNDA 0.013479f
C649 VDDA.n151 GNDA 0.013479f
C650 VDDA.n152 GNDA 0.019629f
C651 VDDA.n154 GNDA 0.013561f
C652 VDDA.n155 GNDA 0.013561f
C653 VDDA.n156 GNDA 0.013561f
C654 VDDA.n158 GNDA 0.10868f
C655 VDDA.n160 GNDA 0.017103f
C656 VDDA.t131 GNDA 0.055426f
C657 VDDA.n161 GNDA 0.0207f
C658 VDDA.n162 GNDA 0.030524f
C659 VDDA.n163 GNDA 0.015289f
C660 VDDA.t172 GNDA 0.013571f
C661 VDDA.n164 GNDA 0.06751f
C662 VDDA.t171 GNDA 0.047014f
C663 VDDA.t85 GNDA 0.029834f
C664 VDDA.t75 GNDA 0.029834f
C665 VDDA.t147 GNDA 0.047014f
C666 VDDA.t148 GNDA 0.013571f
C667 VDDA.n165 GNDA 0.06751f
C668 VDDA.n166 GNDA 0.015289f
C669 VDDA.n167 GNDA 0.036776f
C670 VDDA.n169 GNDA 0.03281f
C671 VDDA.n170 GNDA 0.076182f
C672 VDDA.n171 GNDA 0.105222f
C673 V_mir2.n0 GNDA 0.197463f
C674 V_mir2.t14 GNDA 0.019293f
C675 V_mir2.t12 GNDA 0.019293f
C676 V_mir2.t6 GNDA 0.019293f
C677 V_mir2.n1 GNDA 0.044166f
C678 V_mir2.t11 GNDA 0.02939f
C679 V_mir2.t5 GNDA 0.023151f
C680 V_mir2.t18 GNDA 0.023151f
C681 V_mir2.t17 GNDA 0.037369f
C682 V_mir2.n2 GNDA 0.041731f
C683 V_mir2.n3 GNDA 0.028507f
C684 V_mir2.n4 GNDA 0.044354f
C685 V_mir2.n5 GNDA 0.109943f
C686 V_mir2.t10 GNDA 0.019293f
C687 V_mir2.t8 GNDA 0.019293f
C688 V_mir2.n6 GNDA 0.044166f
C689 V_mir2.t9 GNDA 0.02939f
C690 V_mir2.t7 GNDA 0.023151f
C691 V_mir2.t19 GNDA 0.023151f
C692 V_mir2.t20 GNDA 0.037369f
C693 V_mir2.n7 GNDA 0.041731f
C694 V_mir2.n8 GNDA 0.028507f
C695 V_mir2.n9 GNDA 0.044354f
C696 V_mir2.n10 GNDA 0.085095f
C697 V_mir2.n11 GNDA 0.025223f
C698 V_mir2.t1 GNDA 0.041163f
C699 V_mir2.n12 GNDA 0.027381f
C700 V_mir2.n13 GNDA 0.451535f
C701 V_mir2.n14 GNDA 0.381359f
C702 V_mir2.t3 GNDA 0.02939f
C703 V_mir2.t13 GNDA 0.023151f
C704 V_mir2.t22 GNDA 0.023151f
C705 V_mir2.t21 GNDA 0.037369f
C706 V_mir2.n15 GNDA 0.041731f
C707 V_mir2.n16 GNDA 0.028507f
C708 V_mir2.n17 GNDA 0.044354f
C709 V_mir2.n18 GNDA 0.111042f
C710 V_mir2.n19 GNDA 0.044166f
C711 V_mir2.t4 GNDA 0.019293f
C712 NFET_GATE_10uA.t3 GNDA 0.01496f
C713 NFET_GATE_10uA.t4 GNDA 0.01496f
C714 NFET_GATE_10uA.t1 GNDA 0.01496f
C715 NFET_GATE_10uA.n0 GNDA 0.216655f
C716 NFET_GATE_10uA.t21 GNDA 0.014586f
C717 NFET_GATE_10uA.t15 GNDA 0.014586f
C718 NFET_GATE_10uA.t10 GNDA 0.014586f
C719 NFET_GATE_10uA.t20 GNDA 0.014586f
C720 NFET_GATE_10uA.t14 GNDA 0.014586f
C721 NFET_GATE_10uA.t9 GNDA 0.014586f
C722 NFET_GATE_10uA.t19 GNDA 0.021563f
C723 NFET_GATE_10uA.n1 GNDA 0.026685f
C724 NFET_GATE_10uA.n2 GNDA 0.019075f
C725 NFET_GATE_10uA.n3 GNDA 0.016149f
C726 NFET_GATE_10uA.t23 GNDA 0.014586f
C727 NFET_GATE_10uA.t16 GNDA 0.014586f
C728 NFET_GATE_10uA.t7 GNDA 0.014586f
C729 NFET_GATE_10uA.t8 GNDA 0.021563f
C730 NFET_GATE_10uA.n4 GNDA 0.026685f
C731 NFET_GATE_10uA.n5 GNDA 0.019075f
C732 NFET_GATE_10uA.n6 GNDA 0.016149f
C733 NFET_GATE_10uA.t11 GNDA 0.014586f
C734 NFET_GATE_10uA.t17 GNDA 0.021563f
C735 NFET_GATE_10uA.n7 GNDA 0.02376f
C736 NFET_GATE_10uA.n8 GNDA 0.026114f
C737 NFET_GATE_10uA.t18 GNDA 0.014586f
C738 NFET_GATE_10uA.t13 GNDA 0.021563f
C739 NFET_GATE_10uA.n9 GNDA 0.02376f
C740 NFET_GATE_10uA.t6 GNDA 0.014586f
C741 NFET_GATE_10uA.t5 GNDA 0.014586f
C742 NFET_GATE_10uA.t12 GNDA 0.014586f
C743 NFET_GATE_10uA.t22 GNDA 0.021563f
C744 NFET_GATE_10uA.n10 GNDA 0.026685f
C745 NFET_GATE_10uA.n11 GNDA 0.019075f
C746 NFET_GATE_10uA.n12 GNDA 0.016149f
C747 NFET_GATE_10uA.n13 GNDA 0.026114f
C748 NFET_GATE_10uA.n14 GNDA 0.605807f
C749 NFET_GATE_10uA.n15 GNDA 0.022264f
C750 NFET_GATE_10uA.n16 GNDA 0.016149f
C751 NFET_GATE_10uA.n17 GNDA 0.019075f
C752 NFET_GATE_10uA.n18 GNDA 0.026685f
C753 NFET_GATE_10uA.t2 GNDA 0.034164f
C754 NFET_GATE_10uA.n19 GNDA 1.85977f
C755 NFET_GATE_10uA.n20 GNDA 0.042091f
C756 NFET_GATE_10uA.t0 GNDA 0.01496f
C757 cap_res2.t7 GNDA 0.340442f
C758 cap_res2.t17 GNDA 0.358376f
C759 cap_res2.t1 GNDA 0.359675f
C760 cap_res2.t15 GNDA 0.340442f
C761 cap_res2.t6 GNDA 0.358376f
C762 cap_res2.t19 GNDA 0.359675f
C763 cap_res2.t2 GNDA 0.340442f
C764 cap_res2.t10 GNDA 0.358376f
C765 cap_res2.t4 GNDA 0.359675f
C766 cap_res2.t13 GNDA 0.340442f
C767 cap_res2.t5 GNDA 0.358376f
C768 cap_res2.t16 GNDA 0.359675f
C769 cap_res2.t8 GNDA 0.340442f
C770 cap_res2.t20 GNDA 0.358376f
C771 cap_res2.t11 GNDA 0.359675f
C772 cap_res2.n0 GNDA 0.24022f
C773 cap_res2.t9 GNDA 0.1913f
C774 cap_res2.n1 GNDA 0.260644f
C775 cap_res2.t14 GNDA 0.1913f
C776 cap_res2.n2 GNDA 0.260644f
C777 cap_res2.t3 GNDA 0.1913f
C778 cap_res2.n3 GNDA 0.260644f
C779 cap_res2.t18 GNDA 0.1913f
C780 cap_res2.n4 GNDA 0.260644f
C781 cap_res2.t12 GNDA 0.179319f
C782 cap_res2.t0 GNDA 0.086116f
C783 1st_Vout_2.n0 GNDA 0.723004f
C784 1st_Vout_2.n1 GNDA 1.43086f
C785 1st_Vout_2.n2 GNDA 0.104399f
C786 1st_Vout_2.n3 GNDA 1.45767f
C787 1st_Vout_2.t27 GNDA 0.293375f
C788 1st_Vout_2.t25 GNDA 0.288462f
C789 1st_Vout_2.t11 GNDA 0.293375f
C790 1st_Vout_2.t23 GNDA 0.288462f
C791 1st_Vout_2.t18 GNDA 0.293375f
C792 1st_Vout_2.t17 GNDA 0.288462f
C793 1st_Vout_2.t31 GNDA 0.293375f
C794 1st_Vout_2.t15 GNDA 0.288462f
C795 1st_Vout_2.t35 GNDA 0.293375f
C796 1st_Vout_2.t34 GNDA 0.288462f
C797 1st_Vout_2.t24 GNDA 0.293375f
C798 1st_Vout_2.t33 GNDA 0.288462f
C799 1st_Vout_2.t16 GNDA 0.293375f
C800 1st_Vout_2.t13 GNDA 0.288462f
C801 1st_Vout_2.t30 GNDA 0.293375f
C802 1st_Vout_2.t12 GNDA 0.288462f
C803 1st_Vout_2.t28 GNDA 0.293375f
C804 1st_Vout_2.t19 GNDA 0.288462f
C805 1st_Vout_2.t36 GNDA 0.288462f
C806 1st_Vout_2.t14 GNDA 0.288462f
C807 1st_Vout_2.t22 GNDA 0.018845f
C808 1st_Vout_2.n4 GNDA 0.018179f
C809 1st_Vout_2.t26 GNDA 0.010986f
C810 1st_Vout_2.t20 GNDA 0.010986f
C811 1st_Vout_2.n5 GNDA 0.024439f
C812 1st_Vout_2.n6 GNDA 0.017425f
C813 1st_Vout_2.t3 GNDA 0.015189f
C814 1st_Vout_2.n7 GNDA 0.010417f
C815 1st_Vout_2.n8 GNDA 0.157567f
C816 1st_Vout_2.t21 GNDA 0.010986f
C817 1st_Vout_2.t32 GNDA 0.010986f
C818 1st_Vout_2.n10 GNDA 0.024439f
C819 1st_Vout_2.n11 GNDA 0.018179f
C820 1st_Vout_2.t29 GNDA 0.017243f
.ends

