magic
tech sky130A
timestamp 1738055258
<< nwell >>
rect 885 150 2005 1565
<< nmos >>
rect 1185 -225 1200 -125
rect 1350 -225 1365 -125
rect 1515 -225 1530 -125
rect 1680 -225 1695 -125
rect 1845 -325 1860 -125
rect 1615 -970 1665 -470
rect 1815 -970 1865 -470
<< pmos >>
rect 1115 510 1165 1510
rect 1315 510 1365 1510
rect 1185 175 1200 375
rect 1350 175 1365 375
rect 1515 175 1530 375
rect 1680 175 1695 375
rect 1845 175 1860 575
<< ndiff >>
rect 1135 -140 1185 -125
rect 1135 -210 1150 -140
rect 1170 -210 1185 -140
rect 1135 -225 1185 -210
rect 1200 -140 1250 -125
rect 1200 -210 1215 -140
rect 1235 -210 1250 -140
rect 1200 -225 1250 -210
rect 1300 -140 1350 -125
rect 1300 -210 1315 -140
rect 1335 -210 1350 -140
rect 1300 -225 1350 -210
rect 1365 -140 1415 -125
rect 1365 -210 1380 -140
rect 1400 -210 1415 -140
rect 1365 -225 1415 -210
rect 1465 -140 1515 -125
rect 1465 -210 1480 -140
rect 1500 -210 1515 -140
rect 1465 -225 1515 -210
rect 1530 -140 1580 -125
rect 1530 -210 1545 -140
rect 1565 -210 1580 -140
rect 1530 -225 1580 -210
rect 1630 -140 1680 -125
rect 1630 -210 1645 -140
rect 1665 -210 1680 -140
rect 1630 -225 1680 -210
rect 1695 -140 1745 -125
rect 1695 -210 1710 -140
rect 1730 -210 1745 -140
rect 1695 -225 1745 -210
rect 1795 -140 1845 -125
rect 1795 -310 1810 -140
rect 1830 -310 1845 -140
rect 1795 -325 1845 -310
rect 1860 -140 1910 -125
rect 1860 -310 1875 -140
rect 1895 -310 1910 -140
rect 1860 -325 1910 -310
rect 1565 -485 1615 -470
rect 1565 -955 1580 -485
rect 1600 -955 1615 -485
rect 1565 -970 1615 -955
rect 1665 -485 1715 -470
rect 1665 -955 1680 -485
rect 1700 -955 1715 -485
rect 1665 -970 1715 -955
rect 1765 -485 1815 -470
rect 1765 -955 1780 -485
rect 1800 -955 1815 -485
rect 1765 -970 1815 -955
rect 1865 -485 1915 -470
rect 1865 -955 1880 -485
rect 1900 -955 1915 -485
rect 1865 -970 1915 -955
<< pdiff >>
rect 1065 1495 1115 1510
rect 1065 525 1080 1495
rect 1100 525 1115 1495
rect 1065 510 1115 525
rect 1165 1495 1215 1510
rect 1165 525 1180 1495
rect 1200 525 1215 1495
rect 1165 510 1215 525
rect 1265 1495 1315 1510
rect 1265 525 1280 1495
rect 1300 525 1315 1495
rect 1265 510 1315 525
rect 1365 1495 1415 1510
rect 1365 525 1380 1495
rect 1400 525 1415 1495
rect 1365 510 1415 525
rect 1795 560 1845 575
rect 1135 360 1185 375
rect 1135 190 1150 360
rect 1170 190 1185 360
rect 1135 175 1185 190
rect 1200 360 1250 375
rect 1200 190 1215 360
rect 1235 190 1250 360
rect 1200 175 1250 190
rect 1300 360 1350 375
rect 1300 190 1315 360
rect 1335 190 1350 360
rect 1300 175 1350 190
rect 1365 360 1415 375
rect 1365 190 1380 360
rect 1400 190 1415 360
rect 1365 175 1415 190
rect 1465 360 1515 375
rect 1465 190 1480 360
rect 1500 190 1515 360
rect 1465 175 1515 190
rect 1530 360 1580 375
rect 1530 190 1545 360
rect 1565 190 1580 360
rect 1530 175 1580 190
rect 1630 360 1680 375
rect 1630 190 1645 360
rect 1665 190 1680 360
rect 1630 175 1680 190
rect 1695 360 1745 375
rect 1695 190 1710 360
rect 1730 190 1745 360
rect 1695 175 1745 190
rect 1795 190 1810 560
rect 1830 190 1845 560
rect 1795 175 1845 190
rect 1860 560 1910 575
rect 1860 190 1875 560
rect 1895 190 1910 560
rect 1860 175 1910 190
<< ndiffc >>
rect 1150 -210 1170 -140
rect 1215 -210 1235 -140
rect 1315 -210 1335 -140
rect 1380 -210 1400 -140
rect 1480 -210 1500 -140
rect 1545 -210 1565 -140
rect 1645 -210 1665 -140
rect 1710 -210 1730 -140
rect 1810 -310 1830 -140
rect 1875 -310 1895 -140
rect 1580 -955 1600 -485
rect 1680 -955 1700 -485
rect 1780 -955 1800 -485
rect 1880 -955 1900 -485
<< pdiffc >>
rect 1080 525 1100 1495
rect 1180 525 1200 1495
rect 1280 525 1300 1495
rect 1380 525 1400 1495
rect 1150 190 1170 360
rect 1215 190 1235 360
rect 1315 190 1335 360
rect 1380 190 1400 360
rect 1480 190 1500 360
rect 1545 190 1565 360
rect 1645 190 1665 360
rect 1710 190 1730 360
rect 1810 190 1830 560
rect 1875 190 1895 560
<< psubdiff >>
rect 1225 -320 1325 -305
rect 1225 -340 1240 -320
rect 1310 -340 1325 -320
rect 1225 -355 1325 -340
rect 1725 -370 1825 -355
rect 1725 -390 1740 -370
rect 1810 -390 1825 -370
rect 1725 -405 1825 -390
rect 1970 -660 2020 -645
rect 1970 -680 1985 -660
rect 2005 -680 2020 -660
rect 1970 -695 2020 -680
<< nsubdiff >>
rect 1595 685 1795 700
rect 1595 665 1610 685
rect 1780 665 1795 685
rect 1595 650 1795 665
<< psubdiffcont >>
rect 1240 -340 1310 -320
rect 1740 -390 1810 -370
rect 1985 -680 2005 -660
<< nsubdiffcont >>
rect 1610 665 1780 685
<< poly >>
rect 1320 1555 1360 1560
rect 1320 1535 1330 1555
rect 1350 1535 1360 1555
rect 1320 1525 1360 1535
rect 1115 1510 1165 1525
rect 1315 1510 1365 1525
rect 1845 575 1860 590
rect 1115 500 1165 510
rect 1315 500 1365 510
rect 1115 475 1365 500
rect 720 390 1200 405
rect 735 -55 750 390
rect 1185 375 1200 390
rect 1350 375 1365 390
rect 1515 375 1530 390
rect 1680 375 1695 390
rect 1185 160 1200 175
rect 1350 85 1365 175
rect 1515 165 1530 175
rect 1680 165 1695 175
rect 1515 160 1695 165
rect 1845 160 1860 175
rect 1480 145 1695 160
rect 1805 150 2105 160
rect 1805 145 2075 150
rect 1480 125 1495 145
rect 1515 125 1530 145
rect 1480 110 1530 125
rect 1805 125 1820 145
rect 1840 125 1860 145
rect 1805 110 1860 125
rect 2065 130 2075 145
rect 2095 130 2105 150
rect 2065 120 2105 130
rect 800 70 1640 85
rect 1590 50 1605 70
rect 1625 50 1640 70
rect 1590 35 1640 50
rect 1350 10 1400 25
rect 1350 -10 1365 10
rect 1385 5 1400 10
rect 1385 -10 1860 5
rect 1350 -25 1400 -10
rect 735 -70 1530 -55
rect 1185 -125 1200 -110
rect 1350 -125 1365 -110
rect 1515 -125 1530 -70
rect 1590 -75 1640 -60
rect 1590 -95 1605 -75
rect 1625 -95 1640 -75
rect 1590 -110 1695 -95
rect 1680 -125 1695 -110
rect 1845 -125 1860 -10
rect 1185 -235 1200 -225
rect 1350 -235 1365 -225
rect 1185 -240 1365 -235
rect 1515 -240 1530 -225
rect 1680 -240 1695 -225
rect 1150 -250 1365 -240
rect 1150 -255 1200 -250
rect 1150 -275 1165 -255
rect 1185 -275 1200 -255
rect 1150 -290 1200 -275
rect 2065 -320 2105 -310
rect 1845 -335 1860 -325
rect 2065 -335 2075 -320
rect 1845 -340 2075 -335
rect 2095 -340 2105 -320
rect 1845 -350 2105 -340
rect 1615 -470 1665 -455
rect 1815 -470 1865 -455
rect 1615 -980 1665 -970
rect 1815 -980 1865 -970
rect 1615 -990 1865 -980
rect 1615 -995 1830 -990
rect 1820 -1010 1830 -995
rect 1850 -995 1865 -990
rect 1850 -1010 1860 -995
rect 1820 -1020 1860 -1010
<< polycont >>
rect 1330 1535 1350 1555
rect 1495 125 1515 145
rect 1820 125 1840 145
rect 2075 130 2095 150
rect 1605 50 1625 70
rect 1365 -10 1385 10
rect 1605 -95 1625 -75
rect 1165 -275 1185 -255
rect 2075 -340 2095 -320
rect 1830 -1010 1850 -990
<< xpolycontact >>
rect 2070 528 2105 748
rect 2070 210 2105 430
rect 975 -705 1195 -420
rect 1230 -705 1450 -420
rect 2070 -640 2105 -420
rect 2070 -930 2105 -710
<< xpolyres >>
rect 2070 430 2105 528
rect 1195 -705 1230 -420
rect 2070 -710 2105 -640
<< locali >>
rect 1320 1555 1360 1560
rect 1320 1550 1330 1555
rect 905 1535 1330 1550
rect 1350 1545 1360 1555
rect 1350 1535 1400 1545
rect 905 1530 1400 1535
rect 905 -420 925 1530
rect 1320 1525 1400 1530
rect 1320 1520 1360 1525
rect 1380 1505 1400 1525
rect 1065 1495 1110 1505
rect 1065 525 1080 1495
rect 1100 525 1110 1495
rect 1065 515 1110 525
rect 1170 1495 1215 1505
rect 1170 525 1180 1495
rect 1200 525 1215 1495
rect 1170 515 1215 525
rect 1265 1495 1310 1505
rect 1265 525 1280 1495
rect 1300 525 1310 1495
rect 1265 515 1310 525
rect 1370 1495 1415 1505
rect 1370 525 1380 1495
rect 1400 525 1415 1495
rect 2125 1080 2175 1090
rect 2125 1070 2135 1080
rect 2085 1050 2135 1070
rect 2165 1050 2175 1080
rect 2085 748 2105 1050
rect 2125 1040 2175 1050
rect 1600 685 1790 695
rect 1370 515 1415 525
rect 1495 665 1610 685
rect 1780 665 1830 685
rect 1080 410 1100 515
rect 1180 485 1200 515
rect 1280 485 1300 515
rect 1495 485 1515 665
rect 1180 465 1515 485
rect 1080 390 1335 410
rect 1215 370 1235 390
rect 1315 370 1335 390
rect 1545 370 1565 665
rect 1600 655 1790 665
rect 1645 370 1665 655
rect 1810 570 1830 665
rect 1795 560 1840 570
rect 1135 360 1180 370
rect 1135 190 1150 360
rect 1170 190 1180 360
rect 1135 180 1180 190
rect 1205 360 1250 370
rect 1205 190 1215 360
rect 1235 190 1250 360
rect 1205 180 1250 190
rect 1300 360 1345 370
rect 1300 190 1315 360
rect 1335 190 1345 360
rect 1300 180 1345 190
rect 1370 360 1415 370
rect 1370 190 1380 360
rect 1400 190 1415 360
rect 1370 180 1415 190
rect 1465 360 1510 370
rect 1465 190 1480 360
rect 1500 190 1510 360
rect 1465 180 1510 190
rect 1535 360 1580 370
rect 1535 190 1545 360
rect 1565 190 1580 360
rect 1535 180 1580 190
rect 1630 360 1675 370
rect 1630 190 1645 360
rect 1665 190 1675 360
rect 1630 180 1675 190
rect 1700 360 1745 370
rect 1700 190 1710 360
rect 1730 190 1745 360
rect 1700 180 1745 190
rect 1795 190 1810 560
rect 1830 190 1840 560
rect 1795 180 1840 190
rect 1865 560 1910 570
rect 1865 190 1875 560
rect 1895 190 1910 560
rect 1865 180 1910 190
rect 1150 -130 1170 180
rect 1380 25 1400 180
rect 1350 10 1400 25
rect 1350 -10 1365 10
rect 1385 -10 1400 10
rect 1350 -25 1400 -10
rect 1380 -130 1400 -25
rect 1480 160 1500 180
rect 1710 160 1730 180
rect 1480 145 1530 160
rect 1480 125 1495 145
rect 1515 125 1530 145
rect 1480 110 1530 125
rect 1710 145 1855 160
rect 1710 140 1820 145
rect 1480 -130 1500 110
rect 1590 70 1640 85
rect 1590 50 1605 70
rect 1625 50 1640 70
rect 1590 35 1640 50
rect 1590 -60 1610 35
rect 1590 -75 1640 -60
rect 1590 -95 1605 -75
rect 1625 -95 1640 -75
rect 1590 -110 1640 -95
rect 1710 -130 1730 140
rect 1805 125 1820 140
rect 1840 125 1855 145
rect 1805 110 1855 125
rect 1875 30 1895 180
rect 2070 160 2090 210
rect 2065 150 2105 160
rect 2065 130 2075 150
rect 2095 130 2105 150
rect 2065 120 2105 130
rect 2125 115 2180 125
rect 2125 80 2135 115
rect 2170 80 2180 115
rect 2125 70 2180 80
rect 2125 30 2145 70
rect 1875 10 2285 30
rect 2265 -10 2285 10
rect 2265 -30 3285 -10
rect 2265 -50 2285 -30
rect 1875 -70 2285 -50
rect 1875 -130 1895 -70
rect 2125 -125 2145 -70
rect 1135 -140 1180 -130
rect 1135 -210 1150 -140
rect 1170 -210 1180 -140
rect 1135 -220 1180 -210
rect 1205 -140 1250 -130
rect 1205 -210 1215 -140
rect 1235 -210 1250 -140
rect 1205 -220 1250 -210
rect 1150 -240 1170 -220
rect 1150 -255 1200 -240
rect 1150 -275 1165 -255
rect 1185 -275 1200 -255
rect 1150 -290 1200 -275
rect 1230 -310 1250 -220
rect 1300 -140 1345 -130
rect 1300 -210 1315 -140
rect 1335 -210 1345 -140
rect 1300 -220 1345 -210
rect 1370 -140 1415 -130
rect 1370 -210 1380 -140
rect 1400 -210 1415 -140
rect 1370 -220 1415 -210
rect 1465 -140 1510 -130
rect 1465 -210 1480 -140
rect 1500 -210 1510 -140
rect 1465 -220 1510 -210
rect 1535 -140 1580 -130
rect 1535 -210 1545 -140
rect 1565 -210 1580 -140
rect 1535 -220 1580 -210
rect 1630 -140 1675 -130
rect 1630 -210 1645 -140
rect 1665 -210 1675 -140
rect 1630 -220 1675 -210
rect 1700 -140 1745 -130
rect 1700 -210 1710 -140
rect 1730 -210 1745 -140
rect 1700 -220 1745 -210
rect 1795 -140 1840 -130
rect 1300 -310 1320 -220
rect 1230 -320 1320 -310
rect 1230 -340 1240 -320
rect 1310 -340 1320 -320
rect 1545 -315 1565 -220
rect 1645 -315 1665 -220
rect 1545 -335 1665 -315
rect 1795 -310 1810 -140
rect 1830 -310 1840 -140
rect 1795 -320 1840 -310
rect 1865 -140 1910 -130
rect 1865 -310 1875 -140
rect 1895 -310 1910 -140
rect 2125 -135 2180 -125
rect 2125 -170 2135 -135
rect 2170 -170 2180 -135
rect 2125 -180 2180 -170
rect 1865 -320 1910 -310
rect 2065 -320 2105 -310
rect 1230 -350 1320 -340
rect 905 -440 975 -420
rect 1580 -475 1600 -335
rect 1800 -360 1820 -320
rect 2065 -340 2075 -320
rect 2095 -340 2105 -320
rect 2065 -350 2105 -340
rect 1730 -370 1820 -360
rect 1730 -380 1740 -370
rect 1695 -390 1740 -380
rect 1810 -390 1820 -370
rect 1695 -400 1820 -390
rect 1695 -475 1715 -400
rect 1780 -475 1800 -400
rect 2085 -420 2105 -350
rect 1430 -985 1450 -705
rect 1565 -485 1610 -475
rect 1565 -955 1580 -485
rect 1600 -955 1610 -485
rect 1565 -965 1610 -955
rect 1670 -485 1715 -475
rect 1670 -955 1680 -485
rect 1700 -955 1715 -485
rect 1670 -965 1715 -955
rect 1765 -485 1810 -475
rect 1765 -955 1780 -485
rect 1800 -955 1810 -485
rect 1765 -965 1810 -955
rect 1870 -485 1915 -475
rect 1870 -955 1880 -485
rect 1900 -955 1915 -485
rect 1975 -660 2015 -650
rect 1975 -680 1985 -660
rect 2005 -680 2015 -660
rect 1975 -690 2015 -680
rect 1870 -965 1915 -955
rect 1820 -985 1860 -980
rect 1880 -985 1900 -965
rect 1430 -990 1900 -985
rect 1430 -1005 1830 -990
rect 1820 -1010 1830 -1005
rect 1850 -1005 1900 -990
rect 1850 -1010 1860 -1005
rect 1820 -1020 1860 -1010
rect 2085 -1105 2105 -930
rect 2125 -1105 2175 -1095
rect 2085 -1125 2135 -1105
rect 2125 -1135 2135 -1125
rect 2165 -1135 2175 -1105
rect 2125 -1145 2175 -1135
<< viali >>
rect 1180 525 1200 1495
rect 1280 525 1300 1495
rect 2135 1050 2165 1080
rect 1610 665 1780 685
rect 1545 190 1565 360
rect 1645 190 1665 360
rect 1810 190 1830 560
rect 2135 80 2170 115
rect 1215 -210 1235 -140
rect 1315 -210 1335 -140
rect 1240 -340 1310 -320
rect 1810 -310 1830 -140
rect 2135 -170 2170 -135
rect 1740 -390 1810 -370
rect 1680 -955 1700 -485
rect 1780 -955 1800 -485
rect 2135 -1135 2165 -1105
<< metal1 >>
rect 855 1495 2025 1565
rect 855 525 1180 1495
rect 1200 525 1280 1495
rect 1300 685 2025 1495
rect 2125 1080 2175 1090
rect 2125 1050 2135 1080
rect 2165 1050 2175 1080
rect 2125 1040 2175 1050
rect 1300 665 1610 685
rect 1780 665 2025 685
rect 1300 560 2025 665
rect 1300 525 1810 560
rect 855 360 1810 525
rect 855 190 1545 360
rect 1565 190 1645 360
rect 1665 190 1810 360
rect 1830 190 2025 560
rect 855 150 2025 190
rect 2125 115 2180 125
rect 2125 80 2135 115
rect 2170 80 2180 115
rect 2125 70 2180 80
rect 955 -140 1955 -85
rect 955 -210 1215 -140
rect 1235 -210 1315 -140
rect 1335 -210 1810 -140
rect 955 -310 1810 -210
rect 1830 -310 1955 -140
rect 2125 -135 2180 -125
rect 2125 -170 2135 -135
rect 2170 -170 2180 -135
rect 2125 -180 2180 -170
rect 955 -320 1955 -310
rect 955 -340 1240 -320
rect 1310 -340 1955 -320
rect 955 -370 1955 -340
rect 955 -390 1740 -370
rect 1810 -390 1955 -370
rect 955 -485 1955 -390
rect 955 -745 1680 -485
rect 1510 -795 1680 -745
rect 1515 -955 1680 -795
rect 1700 -955 1780 -485
rect 1800 -955 1955 -485
rect 1515 -1025 1955 -955
rect 2125 -1105 2175 -1095
rect 2125 -1135 2135 -1105
rect 2165 -1135 2175 -1105
rect 2125 -1145 2175 -1135
<< via1 >>
rect 2135 1050 2165 1080
rect 2135 80 2170 115
rect 2135 -170 2170 -135
rect 2135 -1135 2165 -1105
<< metal2 >>
rect 2125 1080 2175 1090
rect 2125 1050 2135 1080
rect 2165 1050 2175 1080
rect 2125 1040 2175 1050
rect 2125 115 2180 125
rect 2125 80 2135 115
rect 2170 80 2180 115
rect 2125 70 2180 80
rect 2125 -135 2180 -125
rect 2125 -170 2135 -135
rect 2170 -170 2180 -135
rect 2125 -180 2180 -170
rect 2125 -1105 2175 -1095
rect 2125 -1135 2135 -1105
rect 2165 -1135 2175 -1105
rect 2125 -1145 2175 -1135
<< via2 >>
rect 2135 1050 2165 1080
rect 2135 80 2170 115
rect 2135 -170 2170 -135
rect 2135 -1135 2165 -1105
<< metal3 >>
rect 2125 1085 2175 1090
rect 2125 1080 3330 1085
rect 2125 1050 2135 1080
rect 2165 1050 3330 1080
rect 2125 1040 3330 1050
rect 2125 115 2180 125
rect 2125 80 2135 115
rect 2170 80 2180 115
rect 2125 70 2180 80
rect 2300 55 3330 1040
rect 2125 -135 2180 -125
rect 2125 -170 2135 -135
rect 2170 -170 2180 -135
rect 2125 -180 2180 -170
rect 2300 -1095 3330 -110
rect 2125 -1105 3330 -1095
rect 2125 -1135 2135 -1105
rect 2165 -1135 3330 -1105
rect 2125 -1140 3330 -1135
rect 2125 -1145 2175 -1140
<< via3 >>
rect 2135 80 2170 115
rect 2135 -170 2170 -135
<< mimcap >>
rect 2315 115 3315 1070
rect 2315 80 2325 115
rect 2360 80 3315 115
rect 2315 70 3315 80
rect 2315 -135 3315 -125
rect 2315 -170 2325 -135
rect 2360 -170 3315 -135
rect 2315 -1125 3315 -170
<< mimcapcontact >>
rect 2325 80 2360 115
rect 2325 -170 2360 -135
<< metal4 >>
rect 2125 115 2365 125
rect 2125 80 2135 115
rect 2170 80 2325 115
rect 2360 80 2365 115
rect 2125 70 2365 80
rect 2125 -135 2365 -125
rect 2125 -170 2135 -135
rect 2170 -170 2325 -135
rect 2360 -170 2365 -135
rect 2125 -180 2365 -170
<< labels >>
flabel metal1 855 795 855 795 7 FreeSans 400 0 0 0 VDDA
flabel metal1 955 -360 955 -360 7 FreeSans 400 0 0 0 GNDA
flabel locali 3285 -20 3285 -20 3 FreeSans 400 0 0 0 VOUT
flabel poly 800 80 800 80 7 FreeSans 400 0 0 0 VIN-
flabel poly 720 400 720 400 7 FreeSans 400 0 0 0 VIN+
<< end >>
